** sch_path: /foss/designs/Analog_FA23_SP24/flashADC/xschem/resistorDivider_v0p0p1.sch
.lib /foss/pdks/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.include /foss/pdks/sky130A/libs.ref/sky130_fd_sc_hd/spice/sky130_fd_sc_hd.spice

.subckt resistorDivider_v0p0p1 VFS V1 V2 V3 V4 V5 V6 V7 V8 V9 V10 V11 V12 V13 V14 V15 V16 VL GND
*.PININFO VFS:I V1:O V2:O V3:O V4:O V5:O V6:O V7:O V8:O V9:O V10:O V11:O V12:O V13:O V14:O V15:O V16:O VL:I GND:I
XR1 VL V1 GND sky130_fd_pr__res_xhigh_po_5p73 L=2.677 mult=8 m=8
XR2 V1 V2 GND sky130_fd_pr__res_xhigh_po_5p73 L=2.677 mult=8 m=8
XR3 V2 V3 GND sky130_fd_pr__res_xhigh_po_5p73 L=2.677 mult=8 m=8
XR4 V3 V4 GND sky130_fd_pr__res_xhigh_po_5p73 L=2.677 mult=8 m=8
XR5 V4 V5 GND sky130_fd_pr__res_xhigh_po_5p73 L=2.677 mult=8 m=8
XR6 V5 V6 GND sky130_fd_pr__res_xhigh_po_5p73 L=2.677 mult=8 m=8
XR7 V6 V7 GND sky130_fd_pr__res_xhigh_po_5p73 L=2.677 mult=8 m=8
XR8 V7 V8 GND sky130_fd_pr__res_xhigh_po_5p73 L=2.677 mult=8 m=8
XR9 V8 V9 GND sky130_fd_pr__res_xhigh_po_5p73 L=2.677 mult=8 m=8
XR10 V9 V10 GND sky130_fd_pr__res_xhigh_po_5p73 L=2.677 mult=8 m=8
XR11 V10 V11 GND sky130_fd_pr__res_xhigh_po_5p73 L=2.677 mult=8 m=8
XR12 V11 V12 GND sky130_fd_pr__res_xhigh_po_5p73 L=2.677 mult=8 m=8
XR13 V12 V13 GND sky130_fd_pr__res_xhigh_po_5p73 L=2.677 mult=8 m=8
XR14 V13 V14 GND sky130_fd_pr__res_xhigh_po_5p73 L=2.677 mult=8 m=8
XR15 V14 V15 GND sky130_fd_pr__res_xhigh_po_5p73 L=2.677 mult=8 m=8
XR16 V15 V16 GND sky130_fd_pr__res_xhigh_po_5p73 L=2.677 mult=8 m=8
XR17 V16 VFS GND sky130_fd_pr__res_xhigh_po_5p73 L=2.677 mult=8 m=8
.ends
.GLOBAL GND
.end
