magic
tech sky130A
magscale 1 2
timestamp 1709390584
<< pwell >>
rect -739 -29232 739 29232
<< psubdiff >>
rect -703 29162 -607 29196
rect 607 29162 703 29196
rect -703 29100 -669 29162
rect 669 29100 703 29162
rect -703 -29162 -669 -29100
rect 669 -29162 703 -29100
rect -703 -29196 -607 -29162
rect 607 -29196 703 -29162
<< psubdiffcont >>
rect -607 29162 607 29196
rect -703 -29100 -669 29100
rect 669 -29100 703 29100
rect -607 -29196 607 -29162
<< xpolycontact >>
rect -573 28634 573 29066
rect -573 -29066 573 -28634
<< xpolyres >>
rect -573 -28634 573 28634
<< locali >>
rect -703 29162 -607 29196
rect 607 29162 703 29196
rect -703 29100 -669 29162
rect 669 29100 703 29162
rect -703 -29162 -669 -29100
rect 669 -29162 703 -29100
rect -703 -29196 -607 -29162
rect 607 -29196 703 -29162
<< viali >>
rect -557 28651 557 29048
rect -557 -29048 557 -28651
<< metal1 >>
rect -569 29048 569 29054
rect -569 28651 -557 29048
rect 557 28651 569 29048
rect -569 28645 569 28651
rect -569 -28651 569 -28645
rect -569 -29048 -557 -28651
rect 557 -29048 569 -28651
rect -569 -29054 569 -29048
<< properties >>
string FIXED_BBOX -686 -29179 686 29179
string gencell sky130_fd_pr__res_xhigh_po_5p73
string library sky130
string parameters w 5.730 l 286.5 m 1 nx 1 wmin 5.730 lmin 0.50 rho 2000 val 100.065k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 5.730 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
