magic
tech sky130A
magscale 1 2
timestamp 1713626893
<< nwell >>
rect -1410 6040 5250 10790
<< locali >>
rect -4070 10060 -3410 10180
rect 7180 10060 7840 10180
rect -4040 8717 -3860 8750
rect -4040 8683 -4039 8717
rect -4005 8683 -3967 8717
rect -3933 8683 -3895 8717
rect -3861 8683 -3860 8717
rect -4040 8650 -3860 8683
rect -3620 8717 -3440 8750
rect -3620 8683 -3619 8717
rect -3585 8683 -3547 8717
rect -3513 8683 -3475 8717
rect -3441 8683 -3440 8717
rect -3620 8650 -3440 8683
rect 7210 8717 7390 8750
rect 7210 8683 7211 8717
rect 7245 8683 7283 8717
rect 7317 8683 7355 8717
rect 7389 8683 7390 8717
rect 7210 8650 7390 8683
rect 7630 8717 7810 8750
rect 7630 8683 7631 8717
rect 7665 8683 7703 8717
rect 7737 8683 7775 8717
rect 7809 8683 7810 8717
rect 7630 8650 7810 8683
rect 900 7639 1470 7670
rect 900 7461 916 7639
rect 1454 7461 1470 7639
rect 900 7430 1470 7461
rect 2370 7639 2940 7670
rect 2370 7461 2386 7639
rect 2924 7461 2940 7639
rect 2370 7430 2940 7461
<< viali >>
rect -4039 8683 -4005 8717
rect -3967 8683 -3933 8717
rect -3895 8683 -3861 8717
rect -3619 8683 -3585 8717
rect -3547 8683 -3513 8717
rect -3475 8683 -3441 8717
rect 7211 8683 7245 8717
rect 7283 8683 7317 8717
rect 7355 8683 7389 8717
rect 7631 8683 7665 8717
rect 7703 8683 7737 8717
rect 7775 8683 7809 8717
rect 916 7461 1454 7639
rect 2386 7461 2924 7639
<< metal1 >>
rect -5050 10230 -4610 11420
rect -5940 10201 -4610 10230
rect -5940 10149 -5801 10201
rect -5749 10149 -4610 10201
rect -5940 10091 -4610 10149
rect -5940 10039 -5911 10091
rect -5859 10039 -4610 10091
rect -5940 10010 -4610 10039
rect -5050 8810 -4610 10010
rect -2620 10150 -2180 11430
rect 1240 10917 2620 10980
rect 1240 10673 1283 10917
rect 1527 10673 2333 10917
rect 2577 10673 2620 10917
rect 1240 10640 2620 10673
rect -1410 10530 5250 10580
rect -1410 10150 -1330 10530
rect -1290 10441 -1200 10450
rect -1290 10389 -1271 10441
rect -1219 10389 -1200 10441
rect -1290 10380 -1200 10389
rect -970 10441 -880 10450
rect -970 10389 -951 10441
rect -899 10389 -880 10441
rect -970 10380 -880 10389
rect -660 10441 -570 10450
rect -660 10389 -641 10441
rect -589 10389 -570 10441
rect -660 10380 -570 10389
rect -340 10441 -250 10450
rect -340 10389 -321 10441
rect -269 10389 -250 10441
rect -340 10380 -250 10389
rect -30 10441 60 10450
rect -30 10389 -11 10441
rect 41 10389 60 10441
rect -30 10380 60 10389
rect 290 10441 380 10450
rect 290 10389 309 10441
rect 361 10389 380 10441
rect 290 10380 380 10389
rect 610 10441 700 10450
rect 610 10389 629 10441
rect 681 10389 700 10441
rect 610 10380 700 10389
rect 920 10441 1010 10450
rect 920 10389 939 10441
rect 991 10389 1010 10441
rect 920 10380 1010 10389
rect 1240 10441 1330 10450
rect 1240 10389 1259 10441
rect 1311 10389 1330 10441
rect 1240 10380 1330 10389
rect 1560 10441 1650 10450
rect 1560 10389 1579 10441
rect 1631 10389 1650 10441
rect 1560 10380 1650 10389
rect 1870 10441 1960 10450
rect 1870 10389 1889 10441
rect 1941 10389 1960 10441
rect 1870 10380 1960 10389
rect 2190 10441 2280 10450
rect 2190 10389 2209 10441
rect 2261 10389 2280 10441
rect 2190 10380 2280 10389
rect 2500 10441 2590 10450
rect 2500 10389 2519 10441
rect 2571 10389 2590 10441
rect 2500 10380 2590 10389
rect 2820 10441 2910 10450
rect 2820 10389 2839 10441
rect 2891 10389 2910 10441
rect 2820 10380 2910 10389
rect 3140 10441 3230 10450
rect 3140 10389 3159 10441
rect 3211 10389 3230 10441
rect 3140 10380 3230 10389
rect 3450 10441 3540 10450
rect 3450 10389 3469 10441
rect 3521 10389 3540 10441
rect 3450 10380 3540 10389
rect 3770 10441 3860 10450
rect 3770 10389 3789 10441
rect 3841 10389 3860 10441
rect 3770 10380 3860 10389
rect 4080 10441 4170 10450
rect 4080 10389 4099 10441
rect 4151 10389 4170 10441
rect 4080 10380 4170 10389
rect 4400 10441 4490 10450
rect 4400 10389 4419 10441
rect 4471 10389 4490 10441
rect 4400 10380 4490 10389
rect 4720 10441 4810 10450
rect 4720 10389 4739 10441
rect 4791 10389 4810 10441
rect 4720 10380 4810 10389
rect 5030 10441 5120 10450
rect 5030 10389 5049 10441
rect 5101 10389 5120 10441
rect 5030 10380 5120 10389
rect -2620 9860 -1330 10150
rect -1290 10201 -1200 10210
rect -1290 10149 -1271 10201
rect -1219 10149 -1200 10201
rect -1290 10140 -1200 10149
rect -970 10201 -880 10210
rect -970 10149 -951 10201
rect -899 10149 -880 10201
rect -970 10140 -880 10149
rect -660 10201 -570 10210
rect -660 10149 -641 10201
rect -589 10149 -570 10201
rect -660 10140 -570 10149
rect -340 10201 -250 10210
rect -340 10149 -321 10201
rect -269 10149 -250 10201
rect -340 10140 -250 10149
rect -30 10201 60 10210
rect -30 10149 -11 10201
rect 41 10149 60 10201
rect -30 10140 60 10149
rect 290 10201 380 10210
rect 290 10149 309 10201
rect 361 10149 380 10201
rect 290 10140 380 10149
rect 610 10201 700 10210
rect 610 10149 629 10201
rect 681 10149 700 10201
rect 610 10140 700 10149
rect 920 10201 1010 10210
rect 920 10149 939 10201
rect 991 10149 1010 10201
rect 920 10140 1010 10149
rect 1240 10201 1330 10210
rect 1240 10149 1259 10201
rect 1311 10149 1330 10201
rect 1240 10140 1330 10149
rect 1560 10201 1650 10210
rect 1560 10149 1579 10201
rect 1631 10149 1650 10201
rect 1560 10140 1650 10149
rect 1870 10201 1960 10210
rect 1870 10149 1889 10201
rect 1941 10149 1960 10201
rect 1870 10140 1960 10149
rect 2190 10201 2280 10210
rect 2190 10149 2209 10201
rect 2261 10149 2280 10201
rect 2190 10140 2280 10149
rect 2500 10201 2590 10210
rect 2500 10149 2519 10201
rect 2571 10149 2590 10201
rect 2500 10140 2590 10149
rect 2820 10201 2910 10210
rect 2820 10149 2839 10201
rect 2891 10149 2910 10201
rect 2820 10140 2910 10149
rect 3140 10201 3230 10210
rect 3140 10149 3159 10201
rect 3211 10149 3230 10201
rect 3140 10140 3230 10149
rect 3450 10201 3540 10210
rect 3450 10149 3469 10201
rect 3521 10149 3540 10201
rect 3450 10140 3540 10149
rect 3770 10201 3860 10210
rect 3770 10149 3789 10201
rect 3841 10149 3860 10201
rect 3770 10140 3860 10149
rect 4080 10201 4170 10210
rect 4080 10149 4099 10201
rect 4151 10149 4170 10201
rect 4080 10140 4170 10149
rect 4400 10201 4490 10210
rect 4400 10149 4419 10201
rect 4471 10149 4490 10201
rect 4400 10140 4490 10149
rect 4720 10201 4810 10210
rect 4720 10149 4739 10201
rect 4791 10149 4810 10201
rect 4720 10140 4810 10149
rect 5030 10201 5120 10210
rect 5030 10149 5049 10201
rect 5101 10149 5120 10201
rect 5030 10140 5120 10149
rect 5170 10150 5250 10530
rect 6020 10150 6450 11420
rect -2620 8810 -2180 9860
rect -1410 9450 -1330 9860
rect 5170 9860 6450 10150
rect -1130 9831 -1040 9840
rect -1130 9779 -1111 9831
rect -1059 9779 -1040 9831
rect -1130 9770 -1040 9779
rect -820 9831 -730 9840
rect -820 9779 -801 9831
rect -749 9779 -730 9831
rect -820 9770 -730 9779
rect -500 9831 -410 9840
rect -500 9779 -481 9831
rect -429 9779 -410 9831
rect -500 9770 -410 9779
rect -180 9831 -90 9840
rect -180 9779 -161 9831
rect -109 9779 -90 9831
rect -180 9770 -90 9779
rect 130 9831 220 9840
rect 130 9779 149 9831
rect 201 9779 220 9831
rect 130 9770 220 9779
rect 450 9831 540 9840
rect 450 9779 469 9831
rect 521 9779 540 9831
rect 450 9770 540 9779
rect 760 9831 850 9840
rect 760 9779 779 9831
rect 831 9779 850 9831
rect 760 9770 850 9779
rect 1080 9831 1170 9840
rect 1080 9779 1099 9831
rect 1151 9779 1170 9831
rect 1080 9770 1170 9779
rect 1400 9831 1490 9840
rect 1400 9779 1419 9831
rect 1471 9779 1490 9831
rect 1400 9770 1490 9779
rect 1710 9831 1800 9840
rect 1710 9779 1729 9831
rect 1781 9779 1800 9831
rect 1710 9770 1800 9779
rect 2030 9831 2120 9840
rect 2030 9779 2049 9831
rect 2101 9779 2120 9831
rect 2030 9770 2120 9779
rect 2350 9831 2440 9840
rect 2350 9779 2369 9831
rect 2421 9779 2440 9831
rect 2350 9770 2440 9779
rect 2660 9831 2750 9840
rect 2660 9779 2679 9831
rect 2731 9779 2750 9831
rect 2660 9770 2750 9779
rect 2980 9831 3070 9840
rect 2980 9779 2999 9831
rect 3051 9779 3070 9831
rect 2980 9770 3070 9779
rect 3290 9831 3380 9840
rect 3290 9779 3309 9831
rect 3361 9779 3380 9831
rect 3290 9770 3380 9779
rect 3610 9831 3700 9840
rect 3610 9779 3629 9831
rect 3681 9779 3700 9831
rect 3610 9770 3700 9779
rect 3930 9831 4020 9840
rect 3930 9779 3949 9831
rect 4001 9779 4020 9831
rect 3930 9770 4020 9779
rect 4240 9831 4330 9840
rect 4240 9779 4259 9831
rect 4311 9779 4330 9831
rect 4240 9770 4330 9779
rect 4560 9831 4650 9840
rect 4560 9779 4579 9831
rect 4631 9779 4650 9831
rect 4560 9770 4650 9779
rect 4880 9831 4970 9840
rect 4880 9779 4899 9831
rect 4951 9779 4970 9831
rect 4880 9770 4970 9779
rect -1130 9591 -1040 9600
rect -1130 9539 -1111 9591
rect -1059 9539 -1040 9591
rect -1130 9530 -1040 9539
rect -820 9591 -730 9600
rect -820 9539 -801 9591
rect -749 9539 -730 9591
rect -820 9530 -730 9539
rect -500 9591 -410 9600
rect -500 9539 -481 9591
rect -429 9539 -410 9591
rect -500 9530 -410 9539
rect -180 9591 -90 9600
rect -180 9539 -161 9591
rect -109 9539 -90 9591
rect -180 9530 -90 9539
rect 130 9591 220 9600
rect 130 9539 149 9591
rect 201 9539 220 9591
rect 130 9530 220 9539
rect 450 9591 540 9600
rect 450 9539 469 9591
rect 521 9539 540 9591
rect 450 9530 540 9539
rect 760 9591 850 9600
rect 760 9539 779 9591
rect 831 9539 850 9591
rect 760 9530 850 9539
rect 1080 9591 1170 9600
rect 1080 9539 1099 9591
rect 1151 9539 1170 9591
rect 1080 9530 1170 9539
rect 1400 9591 1490 9600
rect 1400 9539 1419 9591
rect 1471 9539 1490 9591
rect 1400 9530 1490 9539
rect 1710 9591 1800 9600
rect 1710 9539 1729 9591
rect 1781 9539 1800 9591
rect 1710 9530 1800 9539
rect 2030 9591 2120 9600
rect 2030 9539 2049 9591
rect 2101 9539 2120 9591
rect 2030 9530 2120 9539
rect 2350 9591 2440 9600
rect 2350 9539 2369 9591
rect 2421 9539 2440 9591
rect 2350 9530 2440 9539
rect 2660 9591 2750 9600
rect 2660 9539 2679 9591
rect 2731 9539 2750 9591
rect 2660 9530 2750 9539
rect 2980 9591 3070 9600
rect 2980 9539 2999 9591
rect 3051 9539 3070 9591
rect 2980 9530 3070 9539
rect 3290 9591 3380 9600
rect 3290 9539 3309 9591
rect 3361 9539 3380 9591
rect 3290 9530 3380 9539
rect 3610 9591 3700 9600
rect 3610 9539 3629 9591
rect 3681 9539 3700 9591
rect 3610 9530 3700 9539
rect 3930 9591 4020 9600
rect 3930 9539 3949 9591
rect 4001 9539 4020 9591
rect 3930 9530 4020 9539
rect 4240 9591 4330 9600
rect 4240 9539 4259 9591
rect 4311 9539 4330 9591
rect 4240 9530 4330 9539
rect 4560 9591 4650 9600
rect 4560 9539 4579 9591
rect 4631 9539 4650 9591
rect 4560 9530 4650 9539
rect 4880 9591 4970 9600
rect 4880 9539 4899 9591
rect 4951 9539 4970 9591
rect 4880 9530 4970 9539
rect 5170 9450 5250 9860
rect -1410 9416 5250 9450
rect -1410 9400 -146 9416
rect -200 9364 -146 9400
rect -94 9400 3914 9416
rect -94 9364 -40 9400
rect -200 9340 -40 9364
rect 3860 9364 3914 9400
rect 3966 9400 5250 9416
rect 3966 9364 4020 9400
rect 1020 9277 2810 9350
rect 3860 9340 4020 9364
rect 1020 9033 1283 9277
rect 1527 9033 2333 9277
rect 2577 9033 2810 9277
rect 1020 8960 2810 9033
rect 90 8860 3740 8910
rect -4052 8726 -3848 8756
rect -4052 8674 -4040 8726
rect -3988 8674 -3976 8726
rect -3924 8674 -3912 8726
rect -3860 8674 -3848 8726
rect -4052 8644 -3848 8674
rect -3632 8726 -3428 8756
rect -3632 8674 -3620 8726
rect -3568 8674 -3556 8726
rect -3504 8674 -3492 8726
rect -3440 8674 -3428 8726
rect -3632 8644 -3428 8674
rect 90 7780 170 8860
rect 210 8771 300 8780
rect 210 8719 229 8771
rect 281 8719 300 8771
rect 210 8710 300 8719
rect 530 8771 620 8780
rect 530 8719 549 8771
rect 601 8719 620 8771
rect 530 8710 620 8719
rect 840 8771 930 8780
rect 840 8719 859 8771
rect 911 8719 930 8771
rect 840 8710 930 8719
rect 1160 8771 1250 8780
rect 1160 8719 1179 8771
rect 1231 8719 1250 8771
rect 1160 8710 1250 8719
rect 1480 8771 1570 8780
rect 1480 8719 1499 8771
rect 1551 8719 1570 8771
rect 1480 8710 1570 8719
rect 1790 8771 1880 8780
rect 1790 8719 1809 8771
rect 1861 8719 1880 8771
rect 1790 8710 1880 8719
rect 2110 8771 2200 8780
rect 2110 8719 2129 8771
rect 2181 8719 2200 8771
rect 2110 8710 2200 8719
rect 2430 8771 2520 8780
rect 2430 8719 2449 8771
rect 2501 8719 2520 8771
rect 2430 8710 2520 8719
rect 2740 8771 2830 8780
rect 2740 8719 2759 8771
rect 2811 8719 2830 8771
rect 2740 8710 2830 8719
rect 3060 8771 3150 8780
rect 3060 8719 3079 8771
rect 3131 8719 3150 8771
rect 3060 8710 3150 8719
rect 3370 8771 3460 8780
rect 3370 8719 3389 8771
rect 3441 8719 3460 8771
rect 3370 8710 3460 8719
rect 210 8561 300 8570
rect 210 8509 229 8561
rect 281 8509 300 8561
rect 210 8500 300 8509
rect 530 8561 620 8570
rect 530 8509 549 8561
rect 601 8509 620 8561
rect 530 8500 620 8509
rect 840 8561 930 8570
rect 840 8509 859 8561
rect 911 8509 930 8561
rect 840 8500 930 8509
rect 1160 8561 1250 8570
rect 1160 8509 1179 8561
rect 1231 8509 1250 8561
rect 1160 8500 1250 8509
rect 1480 8561 1570 8570
rect 1480 8509 1499 8561
rect 1551 8509 1570 8561
rect 1480 8500 1570 8509
rect 1790 8561 1880 8570
rect 1790 8509 1809 8561
rect 1861 8509 1880 8561
rect 1790 8500 1880 8509
rect 2110 8561 2200 8570
rect 2110 8509 2129 8561
rect 2181 8509 2200 8561
rect 2110 8500 2200 8509
rect 2430 8561 2520 8570
rect 2430 8509 2449 8561
rect 2501 8509 2520 8561
rect 2430 8500 2520 8509
rect 2740 8561 2830 8570
rect 2740 8509 2759 8561
rect 2811 8509 2830 8561
rect 2740 8500 2830 8509
rect 3060 8561 3150 8570
rect 3060 8509 3079 8561
rect 3131 8509 3150 8561
rect 3060 8500 3150 8509
rect 3370 8561 3460 8570
rect 3370 8509 3389 8561
rect 3441 8509 3460 8561
rect 3370 8500 3460 8509
rect 370 8131 460 8140
rect 370 8079 389 8131
rect 441 8079 460 8131
rect 370 8070 460 8079
rect 690 8131 780 8140
rect 690 8079 709 8131
rect 761 8079 780 8131
rect 690 8070 780 8079
rect 1000 8131 1090 8140
rect 1000 8079 1019 8131
rect 1071 8079 1090 8131
rect 1000 8070 1090 8079
rect 1320 8131 1410 8140
rect 1320 8079 1339 8131
rect 1391 8079 1410 8131
rect 1320 8070 1410 8079
rect 1640 8131 1730 8140
rect 1640 8079 1659 8131
rect 1711 8079 1730 8131
rect 1640 8070 1730 8079
rect 1950 8131 2040 8140
rect 1950 8079 1969 8131
rect 2021 8079 2040 8131
rect 1950 8070 2040 8079
rect 2270 8131 2360 8140
rect 2270 8079 2289 8131
rect 2341 8079 2360 8131
rect 2270 8070 2360 8079
rect 2580 8131 2670 8140
rect 2580 8079 2599 8131
rect 2651 8079 2670 8131
rect 2580 8070 2670 8079
rect 2900 8131 2990 8140
rect 2900 8079 2919 8131
rect 2971 8079 2990 8131
rect 2900 8070 2990 8079
rect 3220 8131 3310 8140
rect 3220 8079 3239 8131
rect 3291 8079 3310 8131
rect 3220 8070 3310 8079
rect 3530 8131 3620 8140
rect 3530 8079 3549 8131
rect 3601 8079 3620 8131
rect 3530 8070 3620 8079
rect 370 7921 460 7930
rect 370 7869 389 7921
rect 441 7869 460 7921
rect 370 7860 460 7869
rect 690 7921 780 7930
rect 690 7869 709 7921
rect 761 7869 780 7921
rect 690 7860 780 7869
rect 1000 7921 1090 7930
rect 1000 7869 1019 7921
rect 1071 7869 1090 7921
rect 1000 7860 1090 7869
rect 1320 7921 1410 7930
rect 1320 7869 1339 7921
rect 1391 7869 1410 7921
rect 1320 7860 1410 7869
rect 1640 7921 1730 7930
rect 1640 7869 1659 7921
rect 1711 7869 1730 7921
rect 1640 7860 1730 7869
rect 1950 7921 2040 7930
rect 1950 7869 1969 7921
rect 2021 7869 2040 7921
rect 1950 7860 2040 7869
rect 2270 7921 2360 7930
rect 2270 7869 2289 7921
rect 2341 7869 2360 7921
rect 2270 7860 2360 7869
rect 2580 7921 2670 7930
rect 2580 7869 2599 7921
rect 2651 7869 2670 7921
rect 2580 7860 2670 7869
rect 2900 7921 2990 7930
rect 2900 7869 2919 7921
rect 2971 7869 2990 7921
rect 2900 7860 2990 7869
rect 3220 7921 3310 7930
rect 3220 7869 3239 7921
rect 3291 7869 3310 7921
rect 3220 7860 3310 7869
rect 3530 7921 3620 7930
rect 3530 7869 3549 7921
rect 3601 7869 3620 7921
rect 3530 7860 3620 7869
rect 3660 7780 3740 8860
rect 6020 8810 6450 9860
rect 8450 10230 8890 11420
rect 8450 10201 9780 10230
rect 8450 10149 9589 10201
rect 9641 10149 9780 10201
rect 8450 10091 9780 10149
rect 8450 10039 9699 10091
rect 9751 10039 9780 10091
rect 8450 10010 9780 10039
rect 8450 8810 8890 10010
rect 7198 8726 7402 8756
rect 7198 8674 7210 8726
rect 7262 8674 7274 8726
rect 7326 8674 7338 8726
rect 7390 8674 7402 8726
rect 7198 8644 7402 8674
rect 7618 8726 7822 8756
rect 7618 8674 7630 8726
rect 7682 8674 7694 8726
rect 7746 8674 7758 8726
rect 7810 8674 7822 8726
rect 7618 8644 7822 8674
rect 90 7730 3740 7780
rect 280 7370 550 7730
rect 1030 7676 1310 7680
rect 888 7672 1482 7676
rect 888 7639 1048 7672
rect 1292 7639 1482 7672
rect 888 7461 916 7639
rect 1454 7461 1482 7639
rect 888 7428 1048 7461
rect 1292 7428 1482 7461
rect 888 7424 1482 7428
rect 1030 7420 1310 7424
rect 1780 7370 2050 7730
rect 2530 7676 2810 7680
rect 2358 7672 2952 7676
rect 2358 7639 2548 7672
rect 2792 7639 2952 7672
rect 2358 7461 2386 7639
rect 2924 7461 2952 7639
rect 2358 7428 2548 7461
rect 2792 7428 2952 7461
rect 2358 7424 2952 7428
rect 2530 7420 2810 7424
rect 3280 7370 3550 7730
rect 280 7320 3550 7370
rect 210 7221 300 7230
rect 210 7169 229 7221
rect 281 7169 300 7221
rect 210 7160 300 7169
rect 530 7221 620 7230
rect 530 7169 549 7221
rect 601 7169 620 7221
rect 530 7160 620 7169
rect 210 7011 300 7020
rect 210 6959 229 7011
rect 281 6959 300 7011
rect 210 6950 300 6959
rect 530 7011 620 7020
rect 530 6959 549 7011
rect 601 6959 620 7011
rect 530 6950 620 6959
rect 700 6600 760 7320
rect 840 7221 930 7230
rect 840 7169 859 7221
rect 911 7169 930 7221
rect 840 7160 930 7169
rect 840 7011 930 7020
rect 840 6959 859 7011
rect 911 6959 930 7011
rect 840 6950 930 6959
rect 1020 6600 1080 7320
rect 1160 7221 1250 7230
rect 1160 7169 1179 7221
rect 1231 7169 1250 7221
rect 1160 7160 1250 7169
rect 1480 7221 1570 7230
rect 1480 7169 1499 7221
rect 1551 7169 1570 7221
rect 1480 7160 1570 7169
rect 1790 7221 1880 7230
rect 1790 7169 1809 7221
rect 1861 7169 1880 7221
rect 1790 7160 1880 7169
rect 2110 7221 2200 7230
rect 2110 7169 2129 7221
rect 2181 7169 2200 7221
rect 2110 7160 2200 7169
rect 2420 7221 2510 7230
rect 2420 7169 2439 7221
rect 2491 7169 2510 7221
rect 2420 7160 2510 7169
rect 2740 7221 2830 7230
rect 2740 7169 2759 7221
rect 2811 7169 2830 7221
rect 2740 7160 2830 7169
rect 1160 7011 1250 7020
rect 1160 6959 1179 7011
rect 1231 6959 1250 7011
rect 1160 6950 1250 6959
rect 1480 7011 1570 7020
rect 1480 6959 1499 7011
rect 1551 6959 1570 7011
rect 1480 6950 1570 6959
rect 1790 7011 1880 7020
rect 1790 6959 1809 7011
rect 1861 6959 1880 7011
rect 1790 6950 1880 6959
rect 2110 7011 2200 7020
rect 2110 6959 2129 7011
rect 2181 6959 2200 7011
rect 2110 6950 2200 6959
rect 2420 7011 2510 7020
rect 2420 6959 2439 7011
rect 2491 6959 2510 7011
rect 2420 6950 2510 6959
rect 2740 7011 2830 7020
rect 2740 6959 2759 7011
rect 2811 6959 2830 7011
rect 2740 6950 2830 6959
rect 2910 6600 2970 7320
rect 3060 7221 3150 7230
rect 3060 7169 3079 7221
rect 3131 7169 3150 7221
rect 3060 7160 3150 7169
rect 3060 7011 3150 7020
rect 3060 6959 3079 7011
rect 3131 6959 3150 7011
rect 3060 6950 3150 6959
rect 3230 6600 3290 7320
rect 3370 7221 3460 7230
rect 3370 7169 3389 7221
rect 3441 7169 3460 7221
rect 3370 7160 3460 7169
rect 3370 7011 3460 7020
rect 3370 6959 3389 7011
rect 3441 6959 3460 7011
rect 3370 6950 3460 6959
rect 370 6591 460 6600
rect 370 6539 389 6591
rect 441 6539 460 6591
rect 370 6530 460 6539
rect 690 6591 780 6600
rect 690 6539 709 6591
rect 761 6539 780 6591
rect 690 6530 780 6539
rect 1000 6591 1090 6600
rect 1000 6539 1019 6591
rect 1071 6539 1090 6591
rect 1000 6530 1090 6539
rect 1320 6591 1410 6600
rect 1320 6539 1339 6591
rect 1391 6539 1410 6591
rect 1320 6530 1410 6539
rect 1630 6591 1720 6600
rect 1630 6539 1649 6591
rect 1701 6539 1720 6591
rect 1630 6530 1720 6539
rect 1950 6591 2040 6600
rect 1950 6539 1969 6591
rect 2021 6539 2040 6591
rect 1950 6530 2040 6539
rect 2270 6591 2360 6600
rect 2270 6539 2289 6591
rect 2341 6539 2360 6591
rect 2270 6530 2360 6539
rect 2580 6591 2670 6600
rect 2580 6539 2599 6591
rect 2651 6539 2670 6591
rect 2580 6530 2670 6539
rect 2900 6591 2990 6600
rect 2900 6539 2919 6591
rect 2971 6539 2990 6591
rect 2900 6530 2990 6539
rect 3210 6591 3300 6600
rect 3210 6539 3229 6591
rect 3281 6539 3300 6591
rect 3210 6530 3300 6539
rect 3530 6591 3620 6600
rect 3530 6539 3549 6591
rect 3601 6539 3620 6591
rect 3530 6530 3620 6539
rect 700 6390 760 6530
rect 1020 6390 1080 6530
rect 2910 6390 2970 6530
rect 3230 6390 3290 6530
rect 370 6381 460 6390
rect 370 6329 389 6381
rect 441 6329 460 6381
rect 370 6320 460 6329
rect 690 6381 780 6390
rect 690 6329 709 6381
rect 761 6329 780 6381
rect 690 6320 780 6329
rect 1000 6381 1090 6390
rect 1000 6329 1019 6381
rect 1071 6329 1090 6381
rect 1000 6320 1090 6329
rect 1320 6381 1410 6390
rect 1320 6329 1339 6381
rect 1391 6329 1410 6381
rect 1320 6320 1410 6329
rect 1630 6381 1720 6390
rect 1630 6329 1649 6381
rect 1701 6329 1720 6381
rect 1630 6320 1720 6329
rect 1950 6381 2040 6390
rect 1950 6329 1969 6381
rect 2021 6329 2040 6381
rect 1950 6320 2040 6329
rect 2270 6381 2360 6390
rect 2270 6329 2289 6381
rect 2341 6329 2360 6381
rect 2270 6320 2360 6329
rect 2580 6381 2670 6390
rect 2580 6329 2599 6381
rect 2651 6329 2670 6381
rect 2580 6320 2670 6329
rect 2900 6381 2990 6390
rect 2900 6329 2919 6381
rect 2971 6329 2990 6381
rect 2900 6320 2990 6329
rect 3210 6381 3300 6390
rect 3210 6329 3229 6381
rect 3281 6329 3300 6381
rect 3210 6320 3300 6329
rect 3530 6381 3620 6390
rect 3530 6329 3549 6381
rect 3601 6329 3620 6381
rect 3530 6320 3620 6329
rect 700 6240 760 6320
rect 1020 6240 1080 6320
rect 2910 6240 2970 6320
rect 3230 6240 3290 6320
rect 280 6190 3550 6240
rect 1130 5740 2690 5790
rect 1130 4680 1210 5740
rect 1310 5661 1400 5670
rect 1310 5609 1329 5661
rect 1381 5609 1400 5661
rect 1310 5600 1400 5609
rect 1630 5661 1720 5670
rect 1630 5609 1649 5661
rect 1701 5609 1720 5661
rect 1630 5600 1720 5609
rect 1940 5661 2030 5670
rect 1940 5609 1959 5661
rect 2011 5609 2030 5661
rect 1940 5600 2030 5609
rect 2260 5661 2350 5670
rect 2260 5609 2279 5661
rect 2331 5609 2350 5661
rect 2260 5600 2350 5609
rect 1310 5371 1400 5380
rect 1310 5319 1329 5371
rect 1381 5319 1400 5371
rect 1310 5310 1400 5319
rect 1630 5371 1720 5380
rect 1630 5319 1649 5371
rect 1701 5319 1720 5371
rect 1630 5310 1720 5319
rect 1940 5371 2030 5380
rect 1940 5319 1959 5371
rect 2011 5319 2030 5371
rect 1940 5310 2030 5319
rect 2260 5371 2350 5380
rect 2260 5319 2279 5371
rect 2331 5319 2350 5371
rect 2260 5310 2350 5319
rect 1470 5101 1560 5110
rect 1470 5049 1489 5101
rect 1541 5049 1560 5101
rect 1470 5040 1560 5049
rect 1780 5101 1870 5110
rect 1780 5049 1799 5101
rect 1851 5049 1870 5101
rect 1780 5040 1870 5049
rect 2100 5101 2190 5110
rect 2100 5049 2119 5101
rect 2171 5049 2190 5101
rect 2100 5040 2190 5049
rect 2420 5101 2510 5110
rect 2420 5049 2439 5101
rect 2491 5049 2510 5101
rect 2420 5040 2510 5049
rect 1470 4811 1560 4820
rect 1470 4759 1489 4811
rect 1541 4759 1560 4811
rect 1470 4750 1560 4759
rect 1780 4811 1870 4820
rect 1780 4759 1799 4811
rect 1851 4759 1870 4811
rect 1780 4750 1870 4759
rect 2100 4811 2190 4820
rect 2100 4759 2119 4811
rect 2171 4759 2190 4811
rect 2100 4750 2190 4759
rect 2420 4811 2510 4820
rect 2420 4759 2439 4811
rect 2491 4759 2510 4811
rect 2420 4750 2510 4759
rect 2610 4680 2690 5740
rect 1130 4630 2690 4680
rect 1770 4572 2050 4580
rect 1770 4328 1788 4572
rect 2032 4328 2050 4572
rect 1770 4320 2050 4328
rect 1130 4220 2690 4270
rect 1130 3160 1210 4220
rect 1310 4141 1400 4150
rect 1310 4089 1329 4141
rect 1381 4089 1400 4141
rect 1310 4080 1400 4089
rect 1630 4141 1720 4150
rect 1630 4089 1649 4141
rect 1701 4089 1720 4141
rect 1630 4080 1720 4089
rect 1940 4141 2030 4150
rect 1940 4089 1959 4141
rect 2011 4089 2030 4141
rect 1940 4080 2030 4089
rect 2260 4141 2350 4150
rect 2260 4089 2279 4141
rect 2331 4089 2350 4141
rect 2260 4080 2350 4089
rect 1310 3851 1400 3860
rect 1310 3799 1329 3851
rect 1381 3799 1400 3851
rect 1310 3790 1400 3799
rect 1630 3851 1720 3860
rect 1630 3799 1649 3851
rect 1701 3799 1720 3851
rect 1630 3790 1720 3799
rect 1940 3851 2030 3860
rect 1940 3799 1959 3851
rect 2011 3799 2030 3851
rect 1940 3790 2030 3799
rect 2260 3851 2350 3860
rect 2260 3799 2279 3851
rect 2331 3799 2350 3851
rect 2260 3790 2350 3799
rect 1470 3581 1560 3590
rect 1470 3529 1489 3581
rect 1541 3529 1560 3581
rect 1470 3520 1560 3529
rect 1780 3581 1870 3590
rect 1780 3529 1799 3581
rect 1851 3529 1870 3581
rect 1780 3520 1870 3529
rect 2100 3581 2190 3590
rect 2100 3529 2119 3581
rect 2171 3529 2190 3581
rect 2100 3520 2190 3529
rect 2420 3581 2510 3590
rect 2420 3529 2439 3581
rect 2491 3529 2510 3581
rect 2420 3520 2510 3529
rect 1470 3291 1560 3300
rect 1470 3239 1489 3291
rect 1541 3239 1560 3291
rect 1470 3230 1560 3239
rect 1780 3291 1870 3300
rect 1780 3239 1799 3291
rect 1851 3239 1870 3291
rect 1780 3230 1870 3239
rect 2100 3291 2190 3300
rect 2100 3239 2119 3291
rect 2171 3239 2190 3291
rect 2100 3230 2190 3239
rect 2420 3291 2510 3300
rect 2420 3239 2439 3291
rect 2491 3239 2510 3291
rect 2420 3230 2510 3239
rect 2610 3160 2690 4220
rect 1130 3110 2690 3160
rect 1770 3052 2050 3060
rect 1770 2808 1788 3052
rect 2032 2808 2050 3052
rect 1770 2800 2050 2808
rect -490 2751 -360 2780
rect -490 2750 -451 2751
rect -500 2700 -451 2750
rect -490 2699 -451 2700
rect -399 2750 -360 2751
rect -240 2751 -110 2780
rect -240 2750 -201 2751
rect -399 2700 -201 2750
rect -399 2699 -360 2700
rect -490 2670 -360 2699
rect -240 2699 -201 2700
rect -149 2750 -110 2751
rect 3910 2751 4040 2780
rect 3910 2750 3949 2751
rect -149 2700 3949 2750
rect -149 2699 -110 2700
rect -240 2670 -110 2699
rect 3910 2699 3949 2700
rect 4001 2750 4040 2751
rect 4160 2751 4290 2780
rect 4160 2750 4199 2751
rect 4001 2700 4199 2750
rect 4001 2699 4040 2700
rect 3910 2670 4040 2699
rect 4160 2699 4199 2700
rect 4251 2750 4290 2751
rect 4251 2700 4300 2750
rect 4251 2699 4290 2700
rect 4160 2670 4290 2699
rect 320 2621 410 2630
rect 320 2569 339 2621
rect 391 2569 410 2621
rect 320 2560 410 2569
rect 840 2621 930 2630
rect 840 2569 859 2621
rect 911 2569 930 2621
rect 840 2560 930 2569
rect 1350 2621 1440 2630
rect 1350 2569 1369 2621
rect 1421 2569 1440 2621
rect 1350 2560 1440 2569
rect 1870 2621 1960 2630
rect 1870 2569 1889 2621
rect 1941 2569 1960 2621
rect 1870 2560 1960 2569
rect 2380 2621 2470 2630
rect 2380 2569 2399 2621
rect 2451 2569 2470 2621
rect 2380 2560 2470 2569
rect 2900 2621 2990 2630
rect 2900 2569 2919 2621
rect 2971 2569 2990 2621
rect 2900 2560 2990 2569
rect 3420 2621 3510 2630
rect 3420 2569 3439 2621
rect 3491 2569 3510 2621
rect 3420 2560 3510 2569
rect 320 2441 410 2450
rect 320 2389 339 2441
rect 391 2389 410 2441
rect 320 2380 410 2389
rect 840 2441 930 2450
rect 840 2389 859 2441
rect 911 2389 930 2441
rect 840 2380 930 2389
rect 1350 2441 1440 2450
rect 1350 2389 1369 2441
rect 1421 2389 1440 2441
rect 1350 2380 1440 2389
rect 1870 2441 1960 2450
rect 1870 2389 1889 2441
rect 1941 2389 1960 2441
rect 1870 2380 1960 2389
rect 2380 2441 2470 2450
rect 2380 2389 2399 2441
rect 2451 2389 2470 2441
rect 2380 2380 2470 2389
rect 2900 2441 2990 2450
rect 2900 2389 2919 2441
rect 2971 2389 2990 2441
rect 2900 2380 2990 2389
rect 3420 2441 3510 2450
rect 3420 2389 3439 2441
rect 3491 2389 3510 2441
rect 3420 2380 3510 2389
rect 580 1951 670 1960
rect 580 1899 599 1951
rect 651 1899 670 1951
rect 580 1890 670 1899
rect 1090 1951 1180 1960
rect 1090 1899 1109 1951
rect 1161 1899 1180 1951
rect 1090 1890 1180 1899
rect 1610 1951 1700 1960
rect 1610 1899 1629 1951
rect 1681 1899 1700 1951
rect 1610 1890 1700 1899
rect 2130 1951 2220 1960
rect 2130 1899 2149 1951
rect 2201 1899 2220 1951
rect 2130 1890 2220 1899
rect 2640 1951 2730 1960
rect 2640 1899 2659 1951
rect 2711 1899 2730 1951
rect 2640 1890 2730 1899
rect 3160 1951 3250 1960
rect 3160 1899 3179 1951
rect 3231 1899 3250 1951
rect 3160 1890 3250 1899
rect 580 1771 670 1780
rect 580 1719 599 1771
rect 651 1719 670 1771
rect 580 1710 670 1719
rect 1090 1771 1180 1780
rect 1090 1719 1109 1771
rect 1161 1719 1180 1771
rect 1090 1710 1180 1719
rect 1610 1771 1700 1780
rect 1610 1719 1629 1771
rect 1681 1719 1700 1771
rect 1610 1710 1700 1719
rect 2130 1771 2220 1780
rect 2130 1719 2149 1771
rect 2201 1719 2220 1771
rect 2130 1710 2220 1719
rect 2640 1771 2730 1780
rect 2640 1719 2659 1771
rect 2711 1719 2730 1771
rect 2640 1710 2730 1719
rect 3160 1771 3250 1780
rect 3160 1719 3179 1771
rect 3231 1719 3250 1771
rect 3160 1710 3250 1719
rect -490 1641 -360 1670
rect -490 1640 -451 1641
rect -500 1590 -451 1640
rect -490 1589 -451 1590
rect -399 1640 -360 1641
rect -240 1641 -110 1670
rect -240 1640 -201 1641
rect -399 1590 -201 1640
rect -399 1589 -360 1590
rect -490 1560 -360 1589
rect -240 1589 -201 1590
rect -149 1640 -110 1641
rect 3910 1641 4040 1670
rect 3910 1640 3949 1641
rect -149 1590 3949 1640
rect -149 1589 -110 1590
rect -240 1560 -110 1589
rect 3910 1589 3949 1590
rect 4001 1640 4040 1641
rect 4160 1641 4290 1670
rect 4160 1640 4199 1641
rect 4001 1590 4199 1640
rect 4001 1589 4040 1590
rect 3910 1560 4040 1589
rect 4160 1589 4199 1590
rect 4251 1640 4290 1641
rect 4251 1590 4300 1640
rect 4251 1589 4290 1590
rect 4160 1560 4290 1589
rect 1780 1537 2050 1540
rect 1780 1293 1793 1537
rect 2037 1293 2050 1537
rect 1780 1280 2050 1293
rect -490 1231 -360 1260
rect -490 1230 -451 1231
rect -500 1180 -451 1230
rect -490 1179 -451 1180
rect -399 1230 -360 1231
rect -240 1231 -110 1260
rect -240 1230 -201 1231
rect -399 1180 -201 1230
rect -399 1179 -360 1180
rect -490 1150 -360 1179
rect -240 1179 -201 1180
rect -149 1230 -110 1231
rect 3910 1231 4040 1260
rect 3910 1230 3949 1231
rect -149 1180 3949 1230
rect -149 1179 -110 1180
rect -240 1150 -110 1179
rect 3910 1179 3949 1180
rect 4001 1230 4040 1231
rect 4160 1231 4290 1260
rect 4160 1230 4199 1231
rect 4001 1180 4199 1230
rect 4001 1179 4040 1180
rect 3910 1150 4040 1179
rect 4160 1179 4199 1180
rect 4251 1230 4290 1231
rect 4251 1180 4300 1230
rect 4251 1179 4290 1180
rect 4160 1150 4290 1179
rect 60 1101 150 1110
rect 60 1049 79 1101
rect 131 1049 150 1101
rect 60 1040 150 1049
rect 580 1101 670 1110
rect 580 1049 599 1101
rect 651 1049 670 1101
rect 580 1040 670 1049
rect 1090 1101 1180 1110
rect 1090 1049 1109 1101
rect 1161 1049 1180 1101
rect 1090 1040 1180 1049
rect 1610 1101 1700 1110
rect 1610 1049 1629 1101
rect 1681 1049 1700 1101
rect 1610 1040 1700 1049
rect 2120 1101 2210 1110
rect 2120 1049 2139 1101
rect 2191 1049 2210 1101
rect 2120 1040 2210 1049
rect 2640 1101 2730 1110
rect 2640 1049 2659 1101
rect 2711 1049 2730 1101
rect 2640 1040 2730 1049
rect 3160 1101 3250 1110
rect 3160 1049 3179 1101
rect 3231 1049 3250 1101
rect 3160 1040 3250 1049
rect 3670 1101 3760 1110
rect 3670 1049 3689 1101
rect 3741 1049 3760 1101
rect 3670 1040 3760 1049
rect 60 921 150 930
rect 60 869 79 921
rect 131 869 150 921
rect 60 860 150 869
rect 580 921 670 930
rect 580 869 599 921
rect 651 869 670 921
rect 580 860 670 869
rect 1090 921 1180 930
rect 1090 869 1109 921
rect 1161 869 1180 921
rect 1090 860 1180 869
rect 1610 921 1700 930
rect 1610 869 1629 921
rect 1681 869 1700 921
rect 1610 860 1700 869
rect 2120 921 2210 930
rect 2120 869 2139 921
rect 2191 869 2210 921
rect 2120 860 2210 869
rect 2640 921 2730 930
rect 2640 869 2659 921
rect 2711 869 2730 921
rect 2640 860 2730 869
rect 3160 921 3250 930
rect 3160 869 3179 921
rect 3231 869 3250 921
rect 3160 860 3250 869
rect 3670 921 3760 930
rect 3670 869 3689 921
rect 3741 869 3760 921
rect 3670 860 3760 869
rect 320 431 410 440
rect 320 379 339 431
rect 391 379 410 431
rect 320 370 410 379
rect 830 431 920 440
rect 830 379 849 431
rect 901 379 920 431
rect 830 370 920 379
rect 1350 431 1440 440
rect 1350 379 1369 431
rect 1421 379 1440 431
rect 1350 370 1440 379
rect 1870 431 1960 440
rect 1870 379 1889 431
rect 1941 379 1960 431
rect 1870 370 1960 379
rect 2380 431 2470 440
rect 2380 379 2399 431
rect 2451 379 2470 431
rect 2380 370 2470 379
rect 2900 431 2990 440
rect 2900 379 2919 431
rect 2971 379 2990 431
rect 2900 370 2990 379
rect 3410 431 3500 440
rect 3410 379 3429 431
rect 3481 379 3500 431
rect 3410 370 3500 379
rect 320 251 410 260
rect 320 199 339 251
rect 391 199 410 251
rect 320 190 410 199
rect 830 251 920 260
rect 830 199 849 251
rect 901 199 920 251
rect 830 190 920 199
rect 1350 251 1440 260
rect 1350 199 1369 251
rect 1421 199 1440 251
rect 1350 190 1440 199
rect 1870 251 1960 260
rect 1870 199 1889 251
rect 1941 199 1960 251
rect 1870 190 1960 199
rect 2380 251 2470 260
rect 2380 199 2399 251
rect 2451 199 2470 251
rect 2380 190 2470 199
rect 2900 251 2990 260
rect 2900 199 2919 251
rect 2971 199 2990 251
rect 2900 190 2990 199
rect 3410 251 3500 260
rect 3410 199 3429 251
rect 3481 199 3500 251
rect 3410 190 3500 199
rect -490 121 -360 150
rect -490 120 -451 121
rect -500 70 -451 120
rect -490 69 -451 70
rect -399 120 -360 121
rect -240 121 -110 150
rect -240 120 -201 121
rect -399 70 -201 120
rect -399 69 -360 70
rect -490 40 -360 69
rect -240 69 -201 70
rect -149 120 -110 121
rect 3910 121 4040 150
rect 3910 120 3949 121
rect -149 70 3949 120
rect -149 69 -110 70
rect -240 40 -110 69
rect 3910 69 3949 70
rect 4001 120 4040 121
rect 4160 121 4290 150
rect 4160 120 4199 121
rect 4001 70 4199 120
rect 4001 69 4040 70
rect 3910 40 4040 69
rect 4160 69 4199 70
rect 4251 120 4290 121
rect 4251 70 4300 120
rect 4251 69 4290 70
rect 4160 40 4290 69
rect 1780 7 2050 10
rect 1780 -237 1793 7
rect 2037 -237 2050 7
rect 1780 -240 2050 -237
<< via1 >>
rect -5801 10149 -5749 10201
rect -5911 10039 -5859 10091
rect 1283 10673 1527 10917
rect 2333 10673 2577 10917
rect -1271 10389 -1219 10441
rect -951 10389 -899 10441
rect -641 10389 -589 10441
rect -321 10389 -269 10441
rect -11 10389 41 10441
rect 309 10389 361 10441
rect 629 10389 681 10441
rect 939 10389 991 10441
rect 1259 10389 1311 10441
rect 1579 10389 1631 10441
rect 1889 10389 1941 10441
rect 2209 10389 2261 10441
rect 2519 10389 2571 10441
rect 2839 10389 2891 10441
rect 3159 10389 3211 10441
rect 3469 10389 3521 10441
rect 3789 10389 3841 10441
rect 4099 10389 4151 10441
rect 4419 10389 4471 10441
rect 4739 10389 4791 10441
rect 5049 10389 5101 10441
rect -1271 10149 -1219 10201
rect -951 10149 -899 10201
rect -641 10149 -589 10201
rect -321 10149 -269 10201
rect -11 10149 41 10201
rect 309 10149 361 10201
rect 629 10149 681 10201
rect 939 10149 991 10201
rect 1259 10149 1311 10201
rect 1579 10149 1631 10201
rect 1889 10149 1941 10201
rect 2209 10149 2261 10201
rect 2519 10149 2571 10201
rect 2839 10149 2891 10201
rect 3159 10149 3211 10201
rect 3469 10149 3521 10201
rect 3789 10149 3841 10201
rect 4099 10149 4151 10201
rect 4419 10149 4471 10201
rect 4739 10149 4791 10201
rect 5049 10149 5101 10201
rect -1111 9779 -1059 9831
rect -801 9779 -749 9831
rect -481 9779 -429 9831
rect -161 9779 -109 9831
rect 149 9779 201 9831
rect 469 9779 521 9831
rect 779 9779 831 9831
rect 1099 9779 1151 9831
rect 1419 9779 1471 9831
rect 1729 9779 1781 9831
rect 2049 9779 2101 9831
rect 2369 9779 2421 9831
rect 2679 9779 2731 9831
rect 2999 9779 3051 9831
rect 3309 9779 3361 9831
rect 3629 9779 3681 9831
rect 3949 9779 4001 9831
rect 4259 9779 4311 9831
rect 4579 9779 4631 9831
rect 4899 9779 4951 9831
rect -1111 9539 -1059 9591
rect -801 9539 -749 9591
rect -481 9539 -429 9591
rect -161 9539 -109 9591
rect 149 9539 201 9591
rect 469 9539 521 9591
rect 779 9539 831 9591
rect 1099 9539 1151 9591
rect 1419 9539 1471 9591
rect 1729 9539 1781 9591
rect 2049 9539 2101 9591
rect 2369 9539 2421 9591
rect 2679 9539 2731 9591
rect 2999 9539 3051 9591
rect 3309 9539 3361 9591
rect 3629 9539 3681 9591
rect 3949 9539 4001 9591
rect 4259 9539 4311 9591
rect 4579 9539 4631 9591
rect 4899 9539 4951 9591
rect -146 9364 -94 9416
rect 3914 9364 3966 9416
rect 1283 9033 1527 9277
rect 2333 9033 2577 9277
rect -4040 8717 -3988 8726
rect -4040 8683 -4039 8717
rect -4039 8683 -4005 8717
rect -4005 8683 -3988 8717
rect -4040 8674 -3988 8683
rect -3976 8717 -3924 8726
rect -3976 8683 -3967 8717
rect -3967 8683 -3933 8717
rect -3933 8683 -3924 8717
rect -3976 8674 -3924 8683
rect -3912 8717 -3860 8726
rect -3912 8683 -3895 8717
rect -3895 8683 -3861 8717
rect -3861 8683 -3860 8717
rect -3912 8674 -3860 8683
rect -3620 8717 -3568 8726
rect -3620 8683 -3619 8717
rect -3619 8683 -3585 8717
rect -3585 8683 -3568 8717
rect -3620 8674 -3568 8683
rect -3556 8717 -3504 8726
rect -3556 8683 -3547 8717
rect -3547 8683 -3513 8717
rect -3513 8683 -3504 8717
rect -3556 8674 -3504 8683
rect -3492 8717 -3440 8726
rect -3492 8683 -3475 8717
rect -3475 8683 -3441 8717
rect -3441 8683 -3440 8717
rect -3492 8674 -3440 8683
rect 229 8719 281 8771
rect 549 8719 601 8771
rect 859 8719 911 8771
rect 1179 8719 1231 8771
rect 1499 8719 1551 8771
rect 1809 8719 1861 8771
rect 2129 8719 2181 8771
rect 2449 8719 2501 8771
rect 2759 8719 2811 8771
rect 3079 8719 3131 8771
rect 3389 8719 3441 8771
rect 229 8509 281 8561
rect 549 8509 601 8561
rect 859 8509 911 8561
rect 1179 8509 1231 8561
rect 1499 8509 1551 8561
rect 1809 8509 1861 8561
rect 2129 8509 2181 8561
rect 2449 8509 2501 8561
rect 2759 8509 2811 8561
rect 3079 8509 3131 8561
rect 3389 8509 3441 8561
rect 389 8079 441 8131
rect 709 8079 761 8131
rect 1019 8079 1071 8131
rect 1339 8079 1391 8131
rect 1659 8079 1711 8131
rect 1969 8079 2021 8131
rect 2289 8079 2341 8131
rect 2599 8079 2651 8131
rect 2919 8079 2971 8131
rect 3239 8079 3291 8131
rect 3549 8079 3601 8131
rect 389 7869 441 7921
rect 709 7869 761 7921
rect 1019 7869 1071 7921
rect 1339 7869 1391 7921
rect 1659 7869 1711 7921
rect 1969 7869 2021 7921
rect 2289 7869 2341 7921
rect 2599 7869 2651 7921
rect 2919 7869 2971 7921
rect 3239 7869 3291 7921
rect 3549 7869 3601 7921
rect 9589 10149 9641 10201
rect 9699 10039 9751 10091
rect 7210 8717 7262 8726
rect 7210 8683 7211 8717
rect 7211 8683 7245 8717
rect 7245 8683 7262 8717
rect 7210 8674 7262 8683
rect 7274 8717 7326 8726
rect 7274 8683 7283 8717
rect 7283 8683 7317 8717
rect 7317 8683 7326 8717
rect 7274 8674 7326 8683
rect 7338 8717 7390 8726
rect 7338 8683 7355 8717
rect 7355 8683 7389 8717
rect 7389 8683 7390 8717
rect 7338 8674 7390 8683
rect 7630 8717 7682 8726
rect 7630 8683 7631 8717
rect 7631 8683 7665 8717
rect 7665 8683 7682 8717
rect 7630 8674 7682 8683
rect 7694 8717 7746 8726
rect 7694 8683 7703 8717
rect 7703 8683 7737 8717
rect 7737 8683 7746 8717
rect 7694 8674 7746 8683
rect 7758 8717 7810 8726
rect 7758 8683 7775 8717
rect 7775 8683 7809 8717
rect 7809 8683 7810 8717
rect 7758 8674 7810 8683
rect 1048 7639 1292 7672
rect 1048 7461 1292 7639
rect 1048 7428 1292 7461
rect 2548 7639 2792 7672
rect 2548 7461 2792 7639
rect 2548 7428 2792 7461
rect 229 7169 281 7221
rect 549 7169 601 7221
rect 229 6959 281 7011
rect 549 6959 601 7011
rect 859 7169 911 7221
rect 859 6959 911 7011
rect 1179 7169 1231 7221
rect 1499 7169 1551 7221
rect 1809 7169 1861 7221
rect 2129 7169 2181 7221
rect 2439 7169 2491 7221
rect 2759 7169 2811 7221
rect 1179 6959 1231 7011
rect 1499 6959 1551 7011
rect 1809 6959 1861 7011
rect 2129 6959 2181 7011
rect 2439 6959 2491 7011
rect 2759 6959 2811 7011
rect 3079 7169 3131 7221
rect 3079 6959 3131 7011
rect 3389 7169 3441 7221
rect 3389 6959 3441 7011
rect 389 6539 441 6591
rect 709 6539 761 6591
rect 1019 6539 1071 6591
rect 1339 6539 1391 6591
rect 1649 6539 1701 6591
rect 1969 6539 2021 6591
rect 2289 6539 2341 6591
rect 2599 6539 2651 6591
rect 2919 6539 2971 6591
rect 3229 6539 3281 6591
rect 3549 6539 3601 6591
rect 389 6329 441 6381
rect 709 6329 761 6381
rect 1019 6329 1071 6381
rect 1339 6329 1391 6381
rect 1649 6329 1701 6381
rect 1969 6329 2021 6381
rect 2289 6329 2341 6381
rect 2599 6329 2651 6381
rect 2919 6329 2971 6381
rect 3229 6329 3281 6381
rect 3549 6329 3601 6381
rect 1329 5609 1381 5661
rect 1649 5609 1701 5661
rect 1959 5609 2011 5661
rect 2279 5609 2331 5661
rect 1329 5319 1381 5371
rect 1649 5319 1701 5371
rect 1959 5319 2011 5371
rect 2279 5319 2331 5371
rect 1489 5049 1541 5101
rect 1799 5049 1851 5101
rect 2119 5049 2171 5101
rect 2439 5049 2491 5101
rect 1489 4759 1541 4811
rect 1799 4759 1851 4811
rect 2119 4759 2171 4811
rect 2439 4759 2491 4811
rect 1788 4328 2032 4572
rect 1329 4089 1381 4141
rect 1649 4089 1701 4141
rect 1959 4089 2011 4141
rect 2279 4089 2331 4141
rect 1329 3799 1381 3851
rect 1649 3799 1701 3851
rect 1959 3799 2011 3851
rect 2279 3799 2331 3851
rect 1489 3529 1541 3581
rect 1799 3529 1851 3581
rect 2119 3529 2171 3581
rect 2439 3529 2491 3581
rect 1489 3239 1541 3291
rect 1799 3239 1851 3291
rect 2119 3239 2171 3291
rect 2439 3239 2491 3291
rect 1788 2808 2032 3052
rect -451 2699 -399 2751
rect -201 2699 -149 2751
rect 3949 2699 4001 2751
rect 4199 2699 4251 2751
rect 339 2569 391 2621
rect 859 2569 911 2621
rect 1369 2569 1421 2621
rect 1889 2569 1941 2621
rect 2399 2569 2451 2621
rect 2919 2569 2971 2621
rect 3439 2569 3491 2621
rect 339 2389 391 2441
rect 859 2389 911 2441
rect 1369 2389 1421 2441
rect 1889 2389 1941 2441
rect 2399 2389 2451 2441
rect 2919 2389 2971 2441
rect 3439 2389 3491 2441
rect 599 1899 651 1951
rect 1109 1899 1161 1951
rect 1629 1899 1681 1951
rect 2149 1899 2201 1951
rect 2659 1899 2711 1951
rect 3179 1899 3231 1951
rect 599 1719 651 1771
rect 1109 1719 1161 1771
rect 1629 1719 1681 1771
rect 2149 1719 2201 1771
rect 2659 1719 2711 1771
rect 3179 1719 3231 1771
rect -451 1589 -399 1641
rect -201 1589 -149 1641
rect 3949 1589 4001 1641
rect 4199 1589 4251 1641
rect 1793 1293 2037 1537
rect -451 1179 -399 1231
rect -201 1179 -149 1231
rect 3949 1179 4001 1231
rect 4199 1179 4251 1231
rect 79 1049 131 1101
rect 599 1049 651 1101
rect 1109 1049 1161 1101
rect 1629 1049 1681 1101
rect 2139 1049 2191 1101
rect 2659 1049 2711 1101
rect 3179 1049 3231 1101
rect 3689 1049 3741 1101
rect 79 869 131 921
rect 599 869 651 921
rect 1109 869 1161 921
rect 1629 869 1681 921
rect 2139 869 2191 921
rect 2659 869 2711 921
rect 3179 869 3231 921
rect 3689 869 3741 921
rect 339 379 391 431
rect 849 379 901 431
rect 1369 379 1421 431
rect 1889 379 1941 431
rect 2399 379 2451 431
rect 2919 379 2971 431
rect 3429 379 3481 431
rect 339 199 391 251
rect 849 199 901 251
rect 1369 199 1421 251
rect 1889 199 1941 251
rect 2399 199 2451 251
rect 2919 199 2971 251
rect 3429 199 3481 251
rect -451 69 -399 121
rect -201 69 -149 121
rect 3949 69 4001 121
rect 4199 69 4251 121
rect 1793 -237 2037 7
<< metal2 >>
rect 1270 10917 1540 10940
rect 1270 10673 1283 10917
rect 1527 10673 1540 10917
rect 1270 10650 1540 10673
rect 2320 10917 2590 10940
rect 2320 10673 2333 10917
rect 2577 10673 2590 10917
rect 2320 10650 2590 10673
rect -1280 10443 -1210 10460
rect -1280 10387 -1273 10443
rect -1217 10387 -1210 10443
rect -1280 10370 -1210 10387
rect -960 10443 -890 10460
rect -960 10387 -953 10443
rect -897 10387 -890 10443
rect -960 10370 -890 10387
rect -650 10443 -580 10460
rect -650 10387 -643 10443
rect -587 10387 -580 10443
rect -650 10370 -580 10387
rect -330 10443 -260 10460
rect -330 10387 -323 10443
rect -267 10387 -260 10443
rect -330 10370 -260 10387
rect -20 10443 50 10460
rect -20 10387 -13 10443
rect 43 10387 50 10443
rect -20 10370 50 10387
rect 300 10443 370 10460
rect 300 10387 307 10443
rect 363 10387 370 10443
rect 300 10370 370 10387
rect 620 10443 690 10460
rect 620 10387 627 10443
rect 683 10387 690 10443
rect 620 10370 690 10387
rect 930 10443 1000 10460
rect 930 10387 937 10443
rect 993 10387 1000 10443
rect 930 10370 1000 10387
rect 1250 10443 1320 10460
rect 1250 10387 1257 10443
rect 1313 10387 1320 10443
rect 1250 10370 1320 10387
rect 1570 10443 1640 10460
rect 1570 10387 1577 10443
rect 1633 10387 1640 10443
rect 1570 10370 1640 10387
rect 1880 10443 1950 10460
rect 1880 10387 1887 10443
rect 1943 10387 1950 10443
rect 1880 10370 1950 10387
rect 2200 10443 2270 10460
rect 2200 10387 2207 10443
rect 2263 10387 2270 10443
rect 2200 10370 2270 10387
rect 2510 10443 2580 10460
rect 2510 10387 2517 10443
rect 2573 10387 2580 10443
rect 2510 10370 2580 10387
rect 2830 10443 2900 10460
rect 2830 10387 2837 10443
rect 2893 10387 2900 10443
rect 2830 10370 2900 10387
rect 3150 10443 3220 10460
rect 3150 10387 3157 10443
rect 3213 10387 3220 10443
rect 3150 10370 3220 10387
rect 3460 10443 3530 10460
rect 3460 10387 3467 10443
rect 3523 10387 3530 10443
rect 3460 10370 3530 10387
rect 3780 10443 3850 10460
rect 3780 10387 3787 10443
rect 3843 10387 3850 10443
rect 3780 10370 3850 10387
rect 4090 10443 4160 10460
rect 4090 10387 4097 10443
rect 4153 10387 4160 10443
rect 4090 10370 4160 10387
rect 4410 10443 4480 10460
rect 4410 10387 4417 10443
rect 4473 10387 4480 10443
rect 4410 10370 4480 10387
rect 4730 10443 4800 10460
rect 4730 10387 4737 10443
rect 4793 10387 4800 10443
rect 4730 10370 4800 10387
rect 5040 10443 5110 10460
rect 5040 10387 5047 10443
rect 5103 10387 5110 10443
rect 5040 10370 5110 10387
rect -5940 10203 -5720 10230
rect -5940 10147 -5803 10203
rect -5747 10147 -5720 10203
rect -5940 10093 -5720 10147
rect -1280 10203 -1210 10220
rect -1280 10147 -1273 10203
rect -1217 10147 -1210 10203
rect -1280 10130 -1210 10147
rect -960 10203 -890 10220
rect -960 10147 -953 10203
rect -897 10147 -890 10203
rect -960 10130 -890 10147
rect -650 10203 -580 10220
rect -650 10147 -643 10203
rect -587 10147 -580 10203
rect -650 10130 -580 10147
rect -330 10203 -260 10220
rect -330 10147 -323 10203
rect -267 10147 -260 10203
rect -330 10130 -260 10147
rect -20 10203 50 10220
rect -20 10147 -13 10203
rect 43 10147 50 10203
rect -20 10130 50 10147
rect 300 10203 370 10220
rect 300 10147 307 10203
rect 363 10147 370 10203
rect 300 10130 370 10147
rect 620 10203 690 10220
rect 620 10147 627 10203
rect 683 10147 690 10203
rect 620 10130 690 10147
rect 930 10203 1000 10220
rect 930 10147 937 10203
rect 993 10147 1000 10203
rect 930 10130 1000 10147
rect 1250 10203 1320 10220
rect 1250 10147 1257 10203
rect 1313 10147 1320 10203
rect 1250 10130 1320 10147
rect 1570 10203 1640 10220
rect 1570 10147 1577 10203
rect 1633 10147 1640 10203
rect 1570 10130 1640 10147
rect 1880 10203 1950 10220
rect 1880 10147 1887 10203
rect 1943 10147 1950 10203
rect 1880 10130 1950 10147
rect 2200 10203 2270 10220
rect 2200 10147 2207 10203
rect 2263 10147 2270 10203
rect 2200 10130 2270 10147
rect 2510 10203 2580 10220
rect 2510 10147 2517 10203
rect 2573 10147 2580 10203
rect 2510 10130 2580 10147
rect 2830 10203 2900 10220
rect 2830 10147 2837 10203
rect 2893 10147 2900 10203
rect 2830 10130 2900 10147
rect 3150 10203 3220 10220
rect 3150 10147 3157 10203
rect 3213 10147 3220 10203
rect 3150 10130 3220 10147
rect 3460 10203 3530 10220
rect 3460 10147 3467 10203
rect 3523 10147 3530 10203
rect 3460 10130 3530 10147
rect 3780 10203 3850 10220
rect 3780 10147 3787 10203
rect 3843 10147 3850 10203
rect 3780 10130 3850 10147
rect 4090 10203 4160 10220
rect 4090 10147 4097 10203
rect 4153 10147 4160 10203
rect 4090 10130 4160 10147
rect 4410 10203 4480 10220
rect 4410 10147 4417 10203
rect 4473 10147 4480 10203
rect 4410 10130 4480 10147
rect 4730 10203 4800 10220
rect 4730 10147 4737 10203
rect 4793 10147 4800 10203
rect 4730 10130 4800 10147
rect 5040 10203 5110 10220
rect 5040 10147 5047 10203
rect 5103 10147 5110 10203
rect 5040 10130 5110 10147
rect 9560 10203 9780 10230
rect 9560 10147 9587 10203
rect 9643 10147 9780 10203
rect -5940 10037 -5913 10093
rect -5857 10037 -5720 10093
rect -5940 10010 -5720 10037
rect 9560 10093 9780 10147
rect 9560 10037 9697 10093
rect 9753 10037 9780 10093
rect 9560 10010 9780 10037
rect -1150 9833 -1020 9850
rect -1150 9777 -1113 9833
rect -1057 9777 -1020 9833
rect -1150 9593 -1020 9777
rect -810 9833 -740 9850
rect -810 9777 -803 9833
rect -747 9777 -740 9833
rect -810 9760 -740 9777
rect -490 9833 -420 9850
rect -490 9777 -483 9833
rect -427 9777 -420 9833
rect -490 9760 -420 9777
rect -170 9833 -100 9850
rect -170 9777 -163 9833
rect -107 9777 -100 9833
rect -170 9760 -100 9777
rect 140 9833 210 9850
rect 140 9777 147 9833
rect 203 9777 210 9833
rect 140 9760 210 9777
rect 460 9833 530 9850
rect 460 9777 467 9833
rect 523 9777 530 9833
rect 460 9760 530 9777
rect 770 9833 840 9850
rect 770 9777 777 9833
rect 833 9777 840 9833
rect 770 9760 840 9777
rect 1090 9833 1160 9850
rect 1090 9777 1097 9833
rect 1153 9777 1160 9833
rect 1090 9760 1160 9777
rect 1410 9833 1480 9850
rect 1410 9777 1417 9833
rect 1473 9777 1480 9833
rect 1410 9760 1480 9777
rect 1720 9833 1790 9850
rect 1720 9777 1727 9833
rect 1783 9777 1790 9833
rect 1720 9760 1790 9777
rect 2040 9833 2110 9850
rect 2040 9777 2047 9833
rect 2103 9777 2110 9833
rect 2040 9760 2110 9777
rect 2360 9833 2430 9850
rect 2360 9777 2367 9833
rect 2423 9777 2430 9833
rect 2360 9760 2430 9777
rect 2670 9833 2740 9850
rect 2670 9777 2677 9833
rect 2733 9777 2740 9833
rect 2670 9760 2740 9777
rect 2990 9833 3060 9850
rect 2990 9777 2997 9833
rect 3053 9777 3060 9833
rect 2990 9760 3060 9777
rect 3300 9833 3370 9850
rect 3300 9777 3307 9833
rect 3363 9777 3370 9833
rect 3300 9760 3370 9777
rect 3620 9833 3690 9850
rect 3620 9777 3627 9833
rect 3683 9777 3690 9833
rect 3620 9760 3690 9777
rect 3940 9833 4010 9850
rect 3940 9777 3947 9833
rect 4003 9777 4010 9833
rect 3940 9760 4010 9777
rect 4250 9833 4320 9850
rect 4250 9777 4257 9833
rect 4313 9777 4320 9833
rect 4250 9760 4320 9777
rect 4570 9833 4640 9850
rect 4570 9777 4577 9833
rect 4633 9777 4640 9833
rect 4570 9760 4640 9777
rect 4860 9833 4990 9850
rect 4860 9777 4897 9833
rect 4953 9777 4990 9833
rect -1150 9537 -1113 9593
rect -1057 9537 -1020 9593
rect -1150 9223 -1020 9537
rect -810 9593 -740 9610
rect -810 9537 -803 9593
rect -747 9537 -740 9593
rect -810 9520 -740 9537
rect -490 9593 -420 9610
rect -490 9537 -483 9593
rect -427 9537 -420 9593
rect -490 9520 -420 9537
rect -170 9593 -100 9610
rect -170 9537 -163 9593
rect -107 9537 -100 9593
rect -170 9520 -100 9537
rect 140 9593 210 9610
rect 140 9537 147 9593
rect 203 9537 210 9593
rect 140 9520 210 9537
rect 460 9593 530 9610
rect 460 9537 467 9593
rect 523 9537 530 9593
rect 460 9520 530 9537
rect 770 9593 840 9610
rect 770 9537 777 9593
rect 833 9537 840 9593
rect 770 9520 840 9537
rect 1090 9593 1160 9610
rect 1090 9537 1097 9593
rect 1153 9537 1160 9593
rect 1090 9520 1160 9537
rect 1410 9593 1480 9610
rect 1410 9537 1417 9593
rect 1473 9537 1480 9593
rect 1410 9520 1480 9537
rect 1720 9593 1790 9610
rect 1720 9537 1727 9593
rect 1783 9537 1790 9593
rect 1720 9520 1790 9537
rect 2040 9593 2110 9610
rect 2040 9537 2047 9593
rect 2103 9537 2110 9593
rect 2040 9520 2110 9537
rect 2360 9593 2430 9610
rect 2360 9537 2367 9593
rect 2423 9537 2430 9593
rect 2360 9520 2430 9537
rect 2670 9593 2740 9610
rect 2670 9537 2677 9593
rect 2733 9537 2740 9593
rect 2670 9520 2740 9537
rect 2990 9593 3060 9610
rect 2990 9537 2997 9593
rect 3053 9537 3060 9593
rect 2990 9520 3060 9537
rect 3300 9593 3370 9610
rect 3300 9537 3307 9593
rect 3363 9537 3370 9593
rect 3300 9520 3370 9537
rect 3620 9593 3690 9610
rect 3620 9537 3627 9593
rect 3683 9537 3690 9593
rect 3620 9520 3690 9537
rect 3940 9593 4010 9610
rect 3940 9537 3947 9593
rect 4003 9537 4010 9593
rect 3940 9520 4010 9537
rect 4250 9593 4320 9610
rect 4250 9537 4257 9593
rect 4313 9537 4320 9593
rect 4250 9520 4320 9537
rect 4570 9593 4640 9610
rect 4570 9537 4577 9593
rect 4633 9537 4640 9593
rect 4570 9520 4640 9537
rect 4860 9593 4990 9777
rect 4860 9537 4897 9593
rect 4953 9537 4990 9593
rect -1150 9167 -1113 9223
rect -1057 9167 -1020 9223
rect -4040 8728 -3860 8760
rect -4040 8726 -4018 8728
rect -3962 8726 -3938 8728
rect -3882 8726 -3860 8728
rect -4040 8672 -4018 8674
rect -3962 8672 -3938 8674
rect -3882 8672 -3860 8674
rect -4040 8640 -3860 8672
rect -3620 8728 -3440 8760
rect -3620 8726 -3598 8728
rect -3542 8726 -3518 8728
rect -3462 8726 -3440 8728
rect -3620 8672 -3598 8674
rect -3542 8672 -3518 8674
rect -3462 8672 -3440 8674
rect -3620 8640 -3440 8672
rect -1150 2613 -1020 9167
rect -200 9416 -40 9450
rect -200 9364 -146 9416
rect -94 9364 -40 9416
rect -200 8118 -40 9364
rect 3860 9416 4020 9450
rect 3860 9364 3914 9416
rect 3966 9364 4020 9416
rect 1270 9277 1540 9300
rect 1270 9033 1283 9277
rect 1527 9033 1540 9277
rect 1270 9010 1540 9033
rect 2320 9277 2590 9300
rect 2320 9033 2333 9277
rect 2577 9033 2590 9277
rect 2320 9010 2590 9033
rect 220 8773 290 8790
rect 220 8717 227 8773
rect 283 8717 290 8773
rect 220 8700 290 8717
rect 540 8773 610 8790
rect 540 8717 547 8773
rect 603 8717 610 8773
rect 540 8700 610 8717
rect 850 8773 920 8790
rect 850 8717 857 8773
rect 913 8717 920 8773
rect 850 8700 920 8717
rect 1170 8773 1240 8790
rect 1170 8717 1177 8773
rect 1233 8717 1240 8773
rect 1170 8700 1240 8717
rect 1490 8773 1560 8790
rect 1490 8717 1497 8773
rect 1553 8717 1560 8773
rect 1490 8700 1560 8717
rect 1800 8773 1870 8790
rect 1800 8717 1807 8773
rect 1863 8717 1870 8773
rect 1800 8700 1870 8717
rect 2120 8773 2190 8790
rect 2120 8717 2127 8773
rect 2183 8717 2190 8773
rect 2120 8700 2190 8717
rect 2440 8773 2510 8790
rect 2440 8717 2447 8773
rect 2503 8717 2510 8773
rect 2440 8700 2510 8717
rect 2750 8773 2820 8790
rect 2750 8717 2757 8773
rect 2813 8717 2820 8773
rect 2750 8700 2820 8717
rect 3070 8773 3140 8790
rect 3070 8717 3077 8773
rect 3133 8717 3140 8773
rect 3070 8700 3140 8717
rect 3380 8773 3450 8790
rect 3380 8717 3387 8773
rect 3443 8717 3450 8773
rect 3380 8700 3450 8717
rect 220 8563 290 8580
rect 220 8507 227 8563
rect 283 8507 290 8563
rect 220 8490 290 8507
rect 540 8563 610 8580
rect 540 8507 547 8563
rect 603 8507 610 8563
rect 540 8490 610 8507
rect 850 8563 920 8580
rect 850 8507 857 8563
rect 913 8507 920 8563
rect 850 8490 920 8507
rect 1170 8563 1240 8580
rect 1170 8507 1177 8563
rect 1233 8507 1240 8563
rect 1170 8490 1240 8507
rect 1490 8563 1560 8580
rect 1490 8507 1497 8563
rect 1553 8507 1560 8563
rect 1490 8490 1560 8507
rect 1800 8563 1870 8580
rect 1800 8507 1807 8563
rect 1863 8507 1870 8563
rect 1800 8490 1870 8507
rect 2120 8563 2190 8580
rect 2120 8507 2127 8563
rect 2183 8507 2190 8563
rect 2120 8490 2190 8507
rect 2440 8563 2510 8580
rect 2440 8507 2447 8563
rect 2503 8507 2510 8563
rect 2440 8490 2510 8507
rect 2750 8563 2820 8580
rect 2750 8507 2757 8563
rect 2813 8507 2820 8563
rect 2750 8490 2820 8507
rect 3070 8563 3140 8580
rect 3070 8507 3077 8563
rect 3133 8507 3140 8563
rect 3070 8490 3140 8507
rect 3380 8563 3450 8580
rect 3380 8507 3387 8563
rect 3443 8507 3450 8563
rect 3380 8490 3450 8507
rect -200 8062 -148 8118
rect -92 8062 -40 8118
rect -200 7938 -40 8062
rect 380 8133 450 8150
rect 380 8077 387 8133
rect 443 8077 450 8133
rect 380 8060 450 8077
rect 700 8133 770 8150
rect 700 8077 707 8133
rect 763 8077 770 8133
rect 700 8060 770 8077
rect 1010 8133 1080 8150
rect 1010 8077 1017 8133
rect 1073 8077 1080 8133
rect 1010 8060 1080 8077
rect 1330 8133 1400 8150
rect 1330 8077 1337 8133
rect 1393 8077 1400 8133
rect 1330 8060 1400 8077
rect 1650 8133 1720 8150
rect 1650 8077 1657 8133
rect 1713 8077 1720 8133
rect 1650 8060 1720 8077
rect 1960 8133 2030 8150
rect 1960 8077 1967 8133
rect 2023 8077 2030 8133
rect 1960 8060 2030 8077
rect 2280 8133 2350 8150
rect 2280 8077 2287 8133
rect 2343 8077 2350 8133
rect 2280 8060 2350 8077
rect 2590 8133 2660 8150
rect 2590 8077 2597 8133
rect 2653 8077 2660 8133
rect 2590 8060 2660 8077
rect 2910 8133 2980 8150
rect 2910 8077 2917 8133
rect 2973 8077 2980 8133
rect 2910 8060 2980 8077
rect 3230 8133 3300 8150
rect 3230 8077 3237 8133
rect 3293 8077 3300 8133
rect 3230 8060 3300 8077
rect 3540 8133 3610 8150
rect 3540 8077 3547 8133
rect 3603 8077 3610 8133
rect 3540 8060 3610 8077
rect 3860 8118 4020 9364
rect 3860 8062 3912 8118
rect 3968 8062 4020 8118
rect -200 7882 -148 7938
rect -92 7882 -40 7938
rect -200 5628 -40 7882
rect 380 7923 450 7940
rect 380 7867 387 7923
rect 443 7867 450 7923
rect 380 7850 450 7867
rect 700 7923 770 7940
rect 700 7867 707 7923
rect 763 7867 770 7923
rect 700 7850 770 7867
rect 1010 7923 1080 7940
rect 1010 7867 1017 7923
rect 1073 7867 1080 7923
rect 1010 7850 1080 7867
rect 1330 7923 1400 7940
rect 1330 7867 1337 7923
rect 1393 7867 1400 7923
rect 1330 7850 1400 7867
rect 1650 7923 1720 7940
rect 1650 7867 1657 7923
rect 1713 7867 1720 7923
rect 1650 7850 1720 7867
rect 1960 7923 2030 7940
rect 1960 7867 1967 7923
rect 2023 7867 2030 7923
rect 1960 7850 2030 7867
rect 2280 7923 2350 7940
rect 2280 7867 2287 7923
rect 2343 7867 2350 7923
rect 2280 7850 2350 7867
rect 2590 7923 2660 7940
rect 2590 7867 2597 7923
rect 2653 7867 2660 7923
rect 2590 7850 2660 7867
rect 2910 7923 2980 7940
rect 2910 7867 2917 7923
rect 2973 7867 2980 7923
rect 2910 7850 2980 7867
rect 3230 7923 3300 7940
rect 3230 7867 3237 7923
rect 3293 7867 3300 7923
rect 3230 7850 3300 7867
rect 3540 7923 3610 7940
rect 3540 7867 3547 7923
rect 3603 7867 3610 7923
rect 3540 7850 3610 7867
rect 3860 7938 4020 8062
rect 3860 7882 3912 7938
rect 3968 7882 4020 7938
rect 1040 7672 1300 7690
rect 1040 7428 1048 7672
rect 1292 7428 1300 7672
rect 1040 7410 1300 7428
rect 2540 7672 2800 7690
rect 2540 7428 2548 7672
rect 2792 7428 2800 7672
rect 2540 7410 2800 7428
rect 220 7223 290 7240
rect 220 7167 227 7223
rect 283 7167 290 7223
rect 220 7150 290 7167
rect 540 7223 610 7240
rect 540 7167 547 7223
rect 603 7167 610 7223
rect 540 7150 610 7167
rect 850 7223 920 7240
rect 850 7167 857 7223
rect 913 7167 920 7223
rect 850 7150 920 7167
rect 1170 7223 1240 7240
rect 1170 7167 1177 7223
rect 1233 7167 1240 7223
rect 1170 7150 1240 7167
rect 1490 7223 1560 7240
rect 1490 7167 1497 7223
rect 1553 7167 1560 7223
rect 1490 7150 1560 7167
rect 1800 7223 1870 7240
rect 1800 7167 1807 7223
rect 1863 7167 1870 7223
rect 1800 7150 1870 7167
rect 2120 7223 2190 7240
rect 2120 7167 2127 7223
rect 2183 7167 2190 7223
rect 2120 7150 2190 7167
rect 2430 7223 2500 7240
rect 2430 7167 2437 7223
rect 2493 7167 2500 7223
rect 2430 7150 2500 7167
rect 2750 7223 2820 7240
rect 2750 7167 2757 7223
rect 2813 7167 2820 7223
rect 2750 7150 2820 7167
rect 3070 7223 3140 7240
rect 3070 7167 3077 7223
rect 3133 7167 3140 7223
rect 3070 7150 3140 7167
rect 3380 7223 3450 7240
rect 3380 7167 3387 7223
rect 3443 7167 3450 7223
rect 3380 7150 3450 7167
rect 220 7013 290 7030
rect 220 6957 227 7013
rect 283 6957 290 7013
rect 220 6940 290 6957
rect 540 7013 610 7030
rect 540 6957 547 7013
rect 603 6957 610 7013
rect 540 6940 610 6957
rect 850 7013 920 7030
rect 850 6957 857 7013
rect 913 6957 920 7013
rect 850 6940 920 6957
rect 1170 7013 1240 7030
rect 1170 6957 1177 7013
rect 1233 6957 1240 7013
rect 1170 6940 1240 6957
rect 1490 7013 1560 7030
rect 1490 6957 1497 7013
rect 1553 6957 1560 7013
rect 1490 6940 1560 6957
rect 1800 7013 1870 7030
rect 1800 6957 1807 7013
rect 1863 6957 1870 7013
rect 1800 6940 1870 6957
rect 2120 7013 2190 7030
rect 2120 6957 2127 7013
rect 2183 6957 2190 7013
rect 2120 6940 2190 6957
rect 2430 7013 2500 7030
rect 2430 6957 2437 7013
rect 2493 6957 2500 7013
rect 2430 6940 2500 6957
rect 2750 7013 2820 7030
rect 2750 6957 2757 7013
rect 2813 6957 2820 7013
rect 2750 6940 2820 6957
rect 3070 7013 3140 7030
rect 3070 6957 3077 7013
rect 3133 6957 3140 7013
rect 3070 6940 3140 6957
rect 3380 7013 3450 7030
rect 3380 6957 3387 7013
rect 3443 6957 3450 7013
rect 3380 6940 3450 6957
rect 380 6593 450 6610
rect 380 6537 387 6593
rect 443 6537 450 6593
rect 380 6520 450 6537
rect 670 6593 800 6610
rect 670 6537 707 6593
rect 763 6537 800 6593
rect 380 6383 450 6400
rect 380 6327 387 6383
rect 443 6327 450 6383
rect 380 6310 450 6327
rect 670 6383 800 6537
rect 1010 6593 1080 6610
rect 1010 6537 1017 6593
rect 1073 6537 1080 6593
rect 1010 6520 1080 6537
rect 1330 6593 1400 6610
rect 1330 6537 1337 6593
rect 1393 6537 1400 6593
rect 1330 6520 1400 6537
rect 1640 6593 1710 6610
rect 1640 6537 1647 6593
rect 1703 6537 1710 6593
rect 1640 6520 1710 6537
rect 1960 6593 2030 6610
rect 1960 6537 1967 6593
rect 2023 6537 2030 6593
rect 1960 6520 2030 6537
rect 2280 6593 2350 6610
rect 2280 6537 2287 6593
rect 2343 6537 2350 6593
rect 2280 6520 2350 6537
rect 2590 6593 2660 6610
rect 2590 6537 2597 6593
rect 2653 6537 2660 6593
rect 2590 6520 2660 6537
rect 2910 6593 2980 6610
rect 2910 6537 2917 6593
rect 2973 6537 2980 6593
rect 2910 6520 2980 6537
rect 3190 6593 3320 6610
rect 3190 6537 3227 6593
rect 3283 6537 3320 6593
rect 670 6327 707 6383
rect 763 6327 800 6383
rect -200 5572 -148 5628
rect -92 5572 -40 5628
rect -200 5408 -40 5572
rect -200 5352 -148 5408
rect -92 5352 -40 5408
rect -200 5300 -40 5352
rect 40 5068 200 5120
rect 40 5012 92 5068
rect 148 5012 200 5068
rect 40 4848 200 5012
rect 40 4792 92 4848
rect 148 4792 200 4848
rect 40 4108 200 4792
rect 40 4052 92 4108
rect 148 4052 200 4108
rect 40 3888 200 4052
rect 40 3832 92 3888
rect 148 3832 200 3888
rect -1150 2557 -1113 2613
rect -1057 2557 -1020 2613
rect -1150 2453 -1020 2557
rect -1150 2397 -1113 2453
rect -1057 2397 -1020 2453
rect -1150 2370 -1020 2397
rect -500 2751 -100 2900
rect -500 2699 -451 2751
rect -399 2699 -201 2751
rect -149 2699 -100 2751
rect -500 1641 -100 2699
rect -500 1589 -451 1641
rect -399 1589 -201 1641
rect -149 1589 -100 1641
rect -500 1231 -100 1589
rect -500 1179 -451 1231
rect -399 1179 -201 1231
rect -149 1179 -100 1231
rect -500 121 -100 1179
rect 40 1103 200 3832
rect 670 3563 800 6327
rect 1010 6383 1080 6400
rect 1010 6327 1017 6383
rect 1073 6327 1080 6383
rect 1010 6310 1080 6327
rect 1330 6383 1400 6400
rect 1330 6327 1337 6383
rect 1393 6327 1400 6383
rect 1330 6310 1400 6327
rect 1640 6383 1710 6400
rect 1640 6327 1647 6383
rect 1703 6327 1710 6383
rect 1640 6310 1710 6327
rect 1960 6383 2030 6400
rect 1960 6327 1967 6383
rect 2023 6327 2030 6383
rect 1960 6310 2030 6327
rect 2280 6383 2350 6400
rect 2280 6327 2287 6383
rect 2343 6327 2350 6383
rect 2280 6310 2350 6327
rect 2590 6383 2660 6400
rect 2590 6327 2597 6383
rect 2653 6327 2660 6383
rect 2590 6310 2660 6327
rect 2910 6383 2980 6400
rect 2910 6327 2917 6383
rect 2973 6327 2980 6383
rect 2910 6310 2980 6327
rect 3190 6383 3320 6537
rect 3540 6593 3610 6610
rect 3540 6537 3547 6593
rect 3603 6537 3610 6593
rect 3540 6520 3610 6537
rect 3190 6327 3227 6383
rect 3283 6327 3320 6383
rect 1320 5663 1390 5680
rect 1320 5607 1327 5663
rect 1383 5607 1390 5663
rect 1320 5590 1390 5607
rect 1640 5663 1710 5680
rect 1640 5607 1647 5663
rect 1703 5607 1710 5663
rect 1640 5590 1710 5607
rect 1950 5663 2020 5680
rect 1950 5607 1957 5663
rect 2013 5607 2020 5663
rect 1950 5590 2020 5607
rect 2270 5663 2340 5680
rect 2270 5607 2277 5663
rect 2333 5607 2340 5663
rect 2270 5590 2340 5607
rect 1320 5373 1390 5390
rect 1320 5317 1327 5373
rect 1383 5317 1390 5373
rect 1320 5300 1390 5317
rect 1640 5373 1710 5390
rect 1640 5317 1647 5373
rect 1703 5317 1710 5373
rect 1640 5300 1710 5317
rect 1950 5373 2020 5390
rect 1950 5317 1957 5373
rect 2013 5317 2020 5373
rect 1950 5300 2020 5317
rect 2270 5373 2340 5390
rect 2270 5317 2277 5373
rect 2333 5317 2340 5373
rect 2270 5300 2340 5317
rect 1480 5103 1550 5120
rect 1480 5047 1487 5103
rect 1543 5047 1550 5103
rect 1480 5030 1550 5047
rect 1790 5103 1860 5120
rect 1790 5047 1797 5103
rect 1853 5047 1860 5103
rect 1790 5030 1860 5047
rect 2110 5103 2180 5120
rect 2110 5047 2117 5103
rect 2173 5047 2180 5103
rect 2110 5030 2180 5047
rect 2430 5103 2500 5120
rect 2430 5047 2437 5103
rect 2493 5047 2500 5103
rect 2430 5030 2500 5047
rect 1480 4813 1550 4830
rect 1480 4757 1487 4813
rect 1543 4757 1550 4813
rect 1480 4740 1550 4757
rect 1790 4813 1860 4830
rect 1790 4757 1797 4813
rect 1853 4757 1860 4813
rect 1790 4740 1860 4757
rect 2110 4813 2180 4830
rect 2110 4757 2117 4813
rect 2173 4757 2180 4813
rect 2110 4740 2180 4757
rect 2430 4813 2500 4830
rect 2430 4757 2437 4813
rect 2493 4757 2500 4813
rect 2430 4740 2500 4757
rect 1780 4572 2040 4590
rect 1780 4328 1788 4572
rect 2032 4328 2040 4572
rect 1780 4310 2040 4328
rect 1320 4143 1390 4160
rect 1320 4087 1327 4143
rect 1383 4087 1390 4143
rect 1320 4070 1390 4087
rect 1640 4143 1710 4160
rect 1640 4087 1647 4143
rect 1703 4087 1710 4143
rect 1640 4070 1710 4087
rect 1950 4143 2020 4160
rect 1950 4087 1957 4143
rect 2013 4087 2020 4143
rect 1950 4070 2020 4087
rect 2270 4143 2340 4160
rect 2270 4087 2277 4143
rect 2333 4087 2340 4143
rect 2270 4070 2340 4087
rect 1320 3853 1390 3870
rect 1320 3797 1327 3853
rect 1383 3797 1390 3853
rect 1320 3780 1390 3797
rect 1640 3853 1710 3870
rect 1640 3797 1647 3853
rect 1703 3797 1710 3853
rect 1640 3780 1710 3797
rect 1950 3853 2020 3870
rect 1950 3797 1957 3853
rect 2013 3797 2020 3853
rect 1950 3780 2020 3797
rect 2270 3853 2340 3870
rect 2270 3797 2277 3853
rect 2333 3797 2340 3853
rect 2270 3780 2340 3797
rect 670 3507 707 3563
rect 763 3507 800 3563
rect 1480 3583 1550 3600
rect 1480 3527 1487 3583
rect 1543 3527 1550 3583
rect 1480 3510 1550 3527
rect 1790 3583 1860 3600
rect 1790 3527 1797 3583
rect 1853 3527 1860 3583
rect 1790 3510 1860 3527
rect 2110 3583 2180 3600
rect 2110 3527 2117 3583
rect 2173 3527 2180 3583
rect 2110 3510 2180 3527
rect 2430 3583 2500 3600
rect 2430 3527 2437 3583
rect 2493 3527 2500 3583
rect 2430 3510 2500 3527
rect 3190 3563 3320 6327
rect 3540 6383 3610 6400
rect 3540 6327 3547 6383
rect 3603 6327 3610 6383
rect 3540 6310 3610 6327
rect 3860 5628 4020 7882
rect 3860 5572 3912 5628
rect 3968 5572 4020 5628
rect 3860 5408 4020 5572
rect 3860 5352 3912 5408
rect 3968 5352 4020 5408
rect 3860 5300 4020 5352
rect 4860 9223 4990 9537
rect 4860 9167 4897 9223
rect 4953 9167 4990 9223
rect 670 3313 800 3507
rect 670 3257 707 3313
rect 763 3257 800 3313
rect 3190 3507 3227 3563
rect 3283 3507 3320 3563
rect 3190 3313 3320 3507
rect 670 3220 800 3257
rect 1480 3293 1550 3310
rect 1480 3237 1487 3293
rect 1543 3237 1550 3293
rect 1480 3220 1550 3237
rect 1790 3293 1860 3310
rect 1790 3237 1797 3293
rect 1853 3237 1860 3293
rect 1790 3220 1860 3237
rect 2110 3293 2180 3310
rect 2110 3237 2117 3293
rect 2173 3237 2180 3293
rect 2110 3220 2180 3237
rect 2430 3293 2500 3310
rect 2430 3237 2437 3293
rect 2493 3237 2500 3293
rect 2430 3220 2500 3237
rect 3190 3257 3227 3313
rect 3283 3257 3320 3313
rect 3190 3220 3320 3257
rect 3620 5068 3780 5120
rect 3620 5012 3672 5068
rect 3728 5012 3780 5068
rect 3620 4848 3780 5012
rect 3620 4792 3672 4848
rect 3728 4792 3780 4848
rect 3620 4108 3780 4792
rect 3620 4052 3672 4108
rect 3728 4052 3780 4108
rect 3620 3888 3780 4052
rect 3620 3832 3672 3888
rect 3728 3832 3780 3888
rect 1780 3052 2040 3070
rect 1780 2808 1788 3052
rect 2032 2808 2040 3052
rect 1780 2790 2040 2808
rect 330 2623 400 2640
rect 330 2567 337 2623
rect 393 2567 400 2623
rect 330 2550 400 2567
rect 850 2623 920 2640
rect 850 2567 857 2623
rect 913 2567 920 2623
rect 850 2550 920 2567
rect 1360 2623 1430 2640
rect 1360 2567 1367 2623
rect 1423 2567 1430 2623
rect 1360 2550 1430 2567
rect 1880 2623 1950 2640
rect 1880 2567 1887 2623
rect 1943 2567 1950 2623
rect 1880 2550 1950 2567
rect 2390 2623 2460 2640
rect 2390 2567 2397 2623
rect 2453 2567 2460 2623
rect 2390 2550 2460 2567
rect 2910 2623 2980 2640
rect 2910 2567 2917 2623
rect 2973 2567 2980 2623
rect 2910 2550 2980 2567
rect 3430 2623 3500 2640
rect 3430 2567 3437 2623
rect 3493 2567 3500 2623
rect 3430 2550 3500 2567
rect 330 2443 400 2460
rect 330 2387 337 2443
rect 393 2387 400 2443
rect 330 2370 400 2387
rect 850 2443 920 2460
rect 850 2387 857 2443
rect 913 2387 920 2443
rect 850 2370 920 2387
rect 1360 2443 1430 2460
rect 1360 2387 1367 2443
rect 1423 2387 1430 2443
rect 1360 2370 1430 2387
rect 1880 2443 1950 2460
rect 1880 2387 1887 2443
rect 1943 2387 1950 2443
rect 1880 2370 1950 2387
rect 2390 2443 2460 2460
rect 2390 2387 2397 2443
rect 2453 2387 2460 2443
rect 2390 2370 2460 2387
rect 2910 2443 2980 2460
rect 2910 2387 2917 2443
rect 2973 2387 2980 2443
rect 2910 2370 2980 2387
rect 3430 2443 3500 2460
rect 3430 2387 3437 2443
rect 3493 2387 3500 2443
rect 3430 2370 3500 2387
rect 590 1953 660 1970
rect 590 1897 597 1953
rect 653 1897 660 1953
rect 590 1880 660 1897
rect 1100 1953 1170 1970
rect 1100 1897 1107 1953
rect 1163 1897 1170 1953
rect 1100 1880 1170 1897
rect 1620 1953 1690 1970
rect 1620 1897 1627 1953
rect 1683 1897 1690 1953
rect 1620 1880 1690 1897
rect 2140 1953 2210 1970
rect 2140 1897 2147 1953
rect 2203 1897 2210 1953
rect 2140 1880 2210 1897
rect 2650 1953 2720 1970
rect 2650 1897 2657 1953
rect 2713 1897 2720 1953
rect 2650 1880 2720 1897
rect 3170 1953 3240 1970
rect 3170 1897 3177 1953
rect 3233 1897 3240 1953
rect 3170 1880 3240 1897
rect 590 1773 660 1790
rect 590 1717 597 1773
rect 653 1717 660 1773
rect 590 1700 660 1717
rect 1100 1773 1170 1790
rect 1100 1717 1107 1773
rect 1163 1717 1170 1773
rect 1100 1700 1170 1717
rect 1620 1773 1690 1790
rect 1620 1717 1627 1773
rect 1683 1717 1690 1773
rect 1620 1700 1690 1717
rect 2140 1773 2210 1790
rect 2140 1717 2147 1773
rect 2203 1717 2210 1773
rect 2140 1700 2210 1717
rect 2650 1773 2720 1790
rect 2650 1717 2657 1773
rect 2713 1717 2720 1773
rect 2650 1700 2720 1717
rect 3170 1773 3240 1790
rect 3170 1717 3177 1773
rect 3233 1717 3240 1773
rect 3170 1700 3240 1717
rect 1790 1537 2040 1550
rect 1790 1293 1793 1537
rect 2037 1293 2040 1537
rect 1790 1280 2040 1293
rect 40 1047 77 1103
rect 133 1047 200 1103
rect 40 923 200 1047
rect 590 1103 660 1120
rect 590 1047 597 1103
rect 653 1047 660 1103
rect 590 1030 660 1047
rect 1100 1103 1170 1120
rect 1100 1047 1107 1103
rect 1163 1047 1170 1103
rect 1100 1030 1170 1047
rect 1620 1103 1690 1120
rect 1620 1047 1627 1103
rect 1683 1047 1690 1103
rect 1620 1030 1690 1047
rect 2130 1103 2200 1120
rect 2130 1047 2137 1103
rect 2193 1047 2200 1103
rect 2130 1030 2200 1047
rect 2650 1103 2720 1120
rect 2650 1047 2657 1103
rect 2713 1047 2720 1103
rect 2650 1030 2720 1047
rect 3170 1103 3240 1120
rect 3170 1047 3177 1103
rect 3233 1047 3240 1103
rect 3170 1030 3240 1047
rect 3620 1103 3780 3832
rect 3620 1047 3687 1103
rect 3743 1047 3780 1103
rect 40 867 77 923
rect 133 867 200 923
rect 40 850 200 867
rect 590 923 660 940
rect 590 867 597 923
rect 653 867 660 923
rect 590 850 660 867
rect 1100 923 1170 940
rect 1100 867 1107 923
rect 1163 867 1170 923
rect 1100 850 1170 867
rect 1620 923 1690 940
rect 1620 867 1627 923
rect 1683 867 1690 923
rect 1620 850 1690 867
rect 2130 923 2200 940
rect 2130 867 2137 923
rect 2193 867 2200 923
rect 2130 850 2200 867
rect 2650 923 2720 940
rect 2650 867 2657 923
rect 2713 867 2720 923
rect 2650 850 2720 867
rect 3170 923 3240 940
rect 3170 867 3177 923
rect 3233 867 3240 923
rect 3170 850 3240 867
rect 3620 923 3780 1047
rect 3620 867 3687 923
rect 3743 867 3780 923
rect 3620 850 3780 867
rect 3900 2751 4300 2900
rect 3900 2699 3949 2751
rect 4001 2699 4199 2751
rect 4251 2699 4300 2751
rect 3900 1641 4300 2699
rect 4860 2613 4990 9167
rect 7210 8728 7390 8760
rect 7210 8726 7232 8728
rect 7288 8726 7312 8728
rect 7368 8726 7390 8728
rect 7210 8672 7232 8674
rect 7288 8672 7312 8674
rect 7368 8672 7390 8674
rect 7210 8640 7390 8672
rect 7630 8728 7810 8760
rect 7630 8726 7652 8728
rect 7708 8726 7732 8728
rect 7788 8726 7810 8728
rect 7630 8672 7652 8674
rect 7708 8672 7732 8674
rect 7788 8672 7810 8674
rect 7630 8640 7810 8672
rect 4860 2557 4897 2613
rect 4953 2557 4990 2613
rect 4860 2453 4990 2557
rect 4860 2397 4897 2453
rect 4953 2397 4990 2453
rect 4860 2370 4990 2397
rect 3900 1589 3949 1641
rect 4001 1589 4199 1641
rect 4251 1589 4300 1641
rect 3900 1231 4300 1589
rect 3900 1179 3949 1231
rect 4001 1179 4199 1231
rect 4251 1179 4300 1231
rect 330 433 400 450
rect 330 377 337 433
rect 393 377 400 433
rect 330 360 400 377
rect 840 433 910 450
rect 840 377 847 433
rect 903 377 910 433
rect 840 360 910 377
rect 1360 433 1430 450
rect 1360 377 1367 433
rect 1423 377 1430 433
rect 1360 360 1430 377
rect 1880 433 1950 450
rect 1880 377 1887 433
rect 1943 377 1950 433
rect 1880 360 1950 377
rect 2390 433 2460 450
rect 2390 377 2397 433
rect 2453 377 2460 433
rect 2390 360 2460 377
rect 2910 433 2980 450
rect 2910 377 2917 433
rect 2973 377 2980 433
rect 2910 360 2980 377
rect 3420 433 3490 450
rect 3420 377 3427 433
rect 3483 377 3490 433
rect 3420 360 3490 377
rect 330 253 400 270
rect 330 197 337 253
rect 393 197 400 253
rect 330 180 400 197
rect 840 253 910 270
rect 840 197 847 253
rect 903 197 910 253
rect 840 180 910 197
rect 1360 253 1430 270
rect 1360 197 1367 253
rect 1423 197 1430 253
rect 1360 180 1430 197
rect 1880 253 1950 270
rect 1880 197 1887 253
rect 1943 197 1950 253
rect 1880 180 1950 197
rect 2390 253 2460 270
rect 2390 197 2397 253
rect 2453 197 2460 253
rect 2390 180 2460 197
rect 2910 253 2980 270
rect 2910 197 2917 253
rect 2973 197 2980 253
rect 2910 180 2980 197
rect 3420 253 3490 270
rect 3420 197 3427 253
rect 3483 197 3490 253
rect 3420 180 3490 197
rect -500 69 -451 121
rect -399 69 -201 121
rect -149 69 -100 121
rect -500 -100 -100 69
rect 3900 121 4300 1179
rect 3900 69 3949 121
rect 4001 69 4199 121
rect 4251 69 4300 121
rect 1790 7 2040 20
rect 1790 -237 1793 7
rect 2037 -237 2040 7
rect 3900 -100 4300 69
rect 1790 -250 2040 -237
<< via2 >>
rect 1297 10687 1513 10903
rect 2347 10687 2563 10903
rect -1273 10441 -1217 10443
rect -1273 10389 -1271 10441
rect -1271 10389 -1219 10441
rect -1219 10389 -1217 10441
rect -1273 10387 -1217 10389
rect -953 10441 -897 10443
rect -953 10389 -951 10441
rect -951 10389 -899 10441
rect -899 10389 -897 10441
rect -953 10387 -897 10389
rect -643 10441 -587 10443
rect -643 10389 -641 10441
rect -641 10389 -589 10441
rect -589 10389 -587 10441
rect -643 10387 -587 10389
rect -323 10441 -267 10443
rect -323 10389 -321 10441
rect -321 10389 -269 10441
rect -269 10389 -267 10441
rect -323 10387 -267 10389
rect -13 10441 43 10443
rect -13 10389 -11 10441
rect -11 10389 41 10441
rect 41 10389 43 10441
rect -13 10387 43 10389
rect 307 10441 363 10443
rect 307 10389 309 10441
rect 309 10389 361 10441
rect 361 10389 363 10441
rect 307 10387 363 10389
rect 627 10441 683 10443
rect 627 10389 629 10441
rect 629 10389 681 10441
rect 681 10389 683 10441
rect 627 10387 683 10389
rect 937 10441 993 10443
rect 937 10389 939 10441
rect 939 10389 991 10441
rect 991 10389 993 10441
rect 937 10387 993 10389
rect 1257 10441 1313 10443
rect 1257 10389 1259 10441
rect 1259 10389 1311 10441
rect 1311 10389 1313 10441
rect 1257 10387 1313 10389
rect 1577 10441 1633 10443
rect 1577 10389 1579 10441
rect 1579 10389 1631 10441
rect 1631 10389 1633 10441
rect 1577 10387 1633 10389
rect 1887 10441 1943 10443
rect 1887 10389 1889 10441
rect 1889 10389 1941 10441
rect 1941 10389 1943 10441
rect 1887 10387 1943 10389
rect 2207 10441 2263 10443
rect 2207 10389 2209 10441
rect 2209 10389 2261 10441
rect 2261 10389 2263 10441
rect 2207 10387 2263 10389
rect 2517 10441 2573 10443
rect 2517 10389 2519 10441
rect 2519 10389 2571 10441
rect 2571 10389 2573 10441
rect 2517 10387 2573 10389
rect 2837 10441 2893 10443
rect 2837 10389 2839 10441
rect 2839 10389 2891 10441
rect 2891 10389 2893 10441
rect 2837 10387 2893 10389
rect 3157 10441 3213 10443
rect 3157 10389 3159 10441
rect 3159 10389 3211 10441
rect 3211 10389 3213 10441
rect 3157 10387 3213 10389
rect 3467 10441 3523 10443
rect 3467 10389 3469 10441
rect 3469 10389 3521 10441
rect 3521 10389 3523 10441
rect 3467 10387 3523 10389
rect 3787 10441 3843 10443
rect 3787 10389 3789 10441
rect 3789 10389 3841 10441
rect 3841 10389 3843 10441
rect 3787 10387 3843 10389
rect 4097 10441 4153 10443
rect 4097 10389 4099 10441
rect 4099 10389 4151 10441
rect 4151 10389 4153 10441
rect 4097 10387 4153 10389
rect 4417 10441 4473 10443
rect 4417 10389 4419 10441
rect 4419 10389 4471 10441
rect 4471 10389 4473 10441
rect 4417 10387 4473 10389
rect 4737 10441 4793 10443
rect 4737 10389 4739 10441
rect 4739 10389 4791 10441
rect 4791 10389 4793 10441
rect 4737 10387 4793 10389
rect 5047 10441 5103 10443
rect 5047 10389 5049 10441
rect 5049 10389 5101 10441
rect 5101 10389 5103 10441
rect 5047 10387 5103 10389
rect -5803 10201 -5747 10203
rect -5803 10149 -5801 10201
rect -5801 10149 -5749 10201
rect -5749 10149 -5747 10201
rect -5803 10147 -5747 10149
rect -1273 10201 -1217 10203
rect -1273 10149 -1271 10201
rect -1271 10149 -1219 10201
rect -1219 10149 -1217 10201
rect -1273 10147 -1217 10149
rect -953 10201 -897 10203
rect -953 10149 -951 10201
rect -951 10149 -899 10201
rect -899 10149 -897 10201
rect -953 10147 -897 10149
rect -643 10201 -587 10203
rect -643 10149 -641 10201
rect -641 10149 -589 10201
rect -589 10149 -587 10201
rect -643 10147 -587 10149
rect -323 10201 -267 10203
rect -323 10149 -321 10201
rect -321 10149 -269 10201
rect -269 10149 -267 10201
rect -323 10147 -267 10149
rect -13 10201 43 10203
rect -13 10149 -11 10201
rect -11 10149 41 10201
rect 41 10149 43 10201
rect -13 10147 43 10149
rect 307 10201 363 10203
rect 307 10149 309 10201
rect 309 10149 361 10201
rect 361 10149 363 10201
rect 307 10147 363 10149
rect 627 10201 683 10203
rect 627 10149 629 10201
rect 629 10149 681 10201
rect 681 10149 683 10201
rect 627 10147 683 10149
rect 937 10201 993 10203
rect 937 10149 939 10201
rect 939 10149 991 10201
rect 991 10149 993 10201
rect 937 10147 993 10149
rect 1257 10201 1313 10203
rect 1257 10149 1259 10201
rect 1259 10149 1311 10201
rect 1311 10149 1313 10201
rect 1257 10147 1313 10149
rect 1577 10201 1633 10203
rect 1577 10149 1579 10201
rect 1579 10149 1631 10201
rect 1631 10149 1633 10201
rect 1577 10147 1633 10149
rect 1887 10201 1943 10203
rect 1887 10149 1889 10201
rect 1889 10149 1941 10201
rect 1941 10149 1943 10201
rect 1887 10147 1943 10149
rect 2207 10201 2263 10203
rect 2207 10149 2209 10201
rect 2209 10149 2261 10201
rect 2261 10149 2263 10201
rect 2207 10147 2263 10149
rect 2517 10201 2573 10203
rect 2517 10149 2519 10201
rect 2519 10149 2571 10201
rect 2571 10149 2573 10201
rect 2517 10147 2573 10149
rect 2837 10201 2893 10203
rect 2837 10149 2839 10201
rect 2839 10149 2891 10201
rect 2891 10149 2893 10201
rect 2837 10147 2893 10149
rect 3157 10201 3213 10203
rect 3157 10149 3159 10201
rect 3159 10149 3211 10201
rect 3211 10149 3213 10201
rect 3157 10147 3213 10149
rect 3467 10201 3523 10203
rect 3467 10149 3469 10201
rect 3469 10149 3521 10201
rect 3521 10149 3523 10201
rect 3467 10147 3523 10149
rect 3787 10201 3843 10203
rect 3787 10149 3789 10201
rect 3789 10149 3841 10201
rect 3841 10149 3843 10201
rect 3787 10147 3843 10149
rect 4097 10201 4153 10203
rect 4097 10149 4099 10201
rect 4099 10149 4151 10201
rect 4151 10149 4153 10201
rect 4097 10147 4153 10149
rect 4417 10201 4473 10203
rect 4417 10149 4419 10201
rect 4419 10149 4471 10201
rect 4471 10149 4473 10201
rect 4417 10147 4473 10149
rect 4737 10201 4793 10203
rect 4737 10149 4739 10201
rect 4739 10149 4791 10201
rect 4791 10149 4793 10201
rect 4737 10147 4793 10149
rect 5047 10201 5103 10203
rect 5047 10149 5049 10201
rect 5049 10149 5101 10201
rect 5101 10149 5103 10201
rect 5047 10147 5103 10149
rect 9587 10201 9643 10203
rect 9587 10149 9589 10201
rect 9589 10149 9641 10201
rect 9641 10149 9643 10201
rect 9587 10147 9643 10149
rect -5913 10091 -5857 10093
rect -5913 10039 -5911 10091
rect -5911 10039 -5859 10091
rect -5859 10039 -5857 10091
rect -5913 10037 -5857 10039
rect 9697 10091 9753 10093
rect 9697 10039 9699 10091
rect 9699 10039 9751 10091
rect 9751 10039 9753 10091
rect 9697 10037 9753 10039
rect -1113 9831 -1057 9833
rect -1113 9779 -1111 9831
rect -1111 9779 -1059 9831
rect -1059 9779 -1057 9831
rect -1113 9777 -1057 9779
rect -803 9831 -747 9833
rect -803 9779 -801 9831
rect -801 9779 -749 9831
rect -749 9779 -747 9831
rect -803 9777 -747 9779
rect -483 9831 -427 9833
rect -483 9779 -481 9831
rect -481 9779 -429 9831
rect -429 9779 -427 9831
rect -483 9777 -427 9779
rect -163 9831 -107 9833
rect -163 9779 -161 9831
rect -161 9779 -109 9831
rect -109 9779 -107 9831
rect -163 9777 -107 9779
rect 147 9831 203 9833
rect 147 9779 149 9831
rect 149 9779 201 9831
rect 201 9779 203 9831
rect 147 9777 203 9779
rect 467 9831 523 9833
rect 467 9779 469 9831
rect 469 9779 521 9831
rect 521 9779 523 9831
rect 467 9777 523 9779
rect 777 9831 833 9833
rect 777 9779 779 9831
rect 779 9779 831 9831
rect 831 9779 833 9831
rect 777 9777 833 9779
rect 1097 9831 1153 9833
rect 1097 9779 1099 9831
rect 1099 9779 1151 9831
rect 1151 9779 1153 9831
rect 1097 9777 1153 9779
rect 1417 9831 1473 9833
rect 1417 9779 1419 9831
rect 1419 9779 1471 9831
rect 1471 9779 1473 9831
rect 1417 9777 1473 9779
rect 1727 9831 1783 9833
rect 1727 9779 1729 9831
rect 1729 9779 1781 9831
rect 1781 9779 1783 9831
rect 1727 9777 1783 9779
rect 2047 9831 2103 9833
rect 2047 9779 2049 9831
rect 2049 9779 2101 9831
rect 2101 9779 2103 9831
rect 2047 9777 2103 9779
rect 2367 9831 2423 9833
rect 2367 9779 2369 9831
rect 2369 9779 2421 9831
rect 2421 9779 2423 9831
rect 2367 9777 2423 9779
rect 2677 9831 2733 9833
rect 2677 9779 2679 9831
rect 2679 9779 2731 9831
rect 2731 9779 2733 9831
rect 2677 9777 2733 9779
rect 2997 9831 3053 9833
rect 2997 9779 2999 9831
rect 2999 9779 3051 9831
rect 3051 9779 3053 9831
rect 2997 9777 3053 9779
rect 3307 9831 3363 9833
rect 3307 9779 3309 9831
rect 3309 9779 3361 9831
rect 3361 9779 3363 9831
rect 3307 9777 3363 9779
rect 3627 9831 3683 9833
rect 3627 9779 3629 9831
rect 3629 9779 3681 9831
rect 3681 9779 3683 9831
rect 3627 9777 3683 9779
rect 3947 9831 4003 9833
rect 3947 9779 3949 9831
rect 3949 9779 4001 9831
rect 4001 9779 4003 9831
rect 3947 9777 4003 9779
rect 4257 9831 4313 9833
rect 4257 9779 4259 9831
rect 4259 9779 4311 9831
rect 4311 9779 4313 9831
rect 4257 9777 4313 9779
rect 4577 9831 4633 9833
rect 4577 9779 4579 9831
rect 4579 9779 4631 9831
rect 4631 9779 4633 9831
rect 4577 9777 4633 9779
rect 4897 9831 4953 9833
rect 4897 9779 4899 9831
rect 4899 9779 4951 9831
rect 4951 9779 4953 9831
rect 4897 9777 4953 9779
rect -1113 9591 -1057 9593
rect -1113 9539 -1111 9591
rect -1111 9539 -1059 9591
rect -1059 9539 -1057 9591
rect -1113 9537 -1057 9539
rect -803 9591 -747 9593
rect -803 9539 -801 9591
rect -801 9539 -749 9591
rect -749 9539 -747 9591
rect -803 9537 -747 9539
rect -483 9591 -427 9593
rect -483 9539 -481 9591
rect -481 9539 -429 9591
rect -429 9539 -427 9591
rect -483 9537 -427 9539
rect -163 9591 -107 9593
rect -163 9539 -161 9591
rect -161 9539 -109 9591
rect -109 9539 -107 9591
rect -163 9537 -107 9539
rect 147 9591 203 9593
rect 147 9539 149 9591
rect 149 9539 201 9591
rect 201 9539 203 9591
rect 147 9537 203 9539
rect 467 9591 523 9593
rect 467 9539 469 9591
rect 469 9539 521 9591
rect 521 9539 523 9591
rect 467 9537 523 9539
rect 777 9591 833 9593
rect 777 9539 779 9591
rect 779 9539 831 9591
rect 831 9539 833 9591
rect 777 9537 833 9539
rect 1097 9591 1153 9593
rect 1097 9539 1099 9591
rect 1099 9539 1151 9591
rect 1151 9539 1153 9591
rect 1097 9537 1153 9539
rect 1417 9591 1473 9593
rect 1417 9539 1419 9591
rect 1419 9539 1471 9591
rect 1471 9539 1473 9591
rect 1417 9537 1473 9539
rect 1727 9591 1783 9593
rect 1727 9539 1729 9591
rect 1729 9539 1781 9591
rect 1781 9539 1783 9591
rect 1727 9537 1783 9539
rect 2047 9591 2103 9593
rect 2047 9539 2049 9591
rect 2049 9539 2101 9591
rect 2101 9539 2103 9591
rect 2047 9537 2103 9539
rect 2367 9591 2423 9593
rect 2367 9539 2369 9591
rect 2369 9539 2421 9591
rect 2421 9539 2423 9591
rect 2367 9537 2423 9539
rect 2677 9591 2733 9593
rect 2677 9539 2679 9591
rect 2679 9539 2731 9591
rect 2731 9539 2733 9591
rect 2677 9537 2733 9539
rect 2997 9591 3053 9593
rect 2997 9539 2999 9591
rect 2999 9539 3051 9591
rect 3051 9539 3053 9591
rect 2997 9537 3053 9539
rect 3307 9591 3363 9593
rect 3307 9539 3309 9591
rect 3309 9539 3361 9591
rect 3361 9539 3363 9591
rect 3307 9537 3363 9539
rect 3627 9591 3683 9593
rect 3627 9539 3629 9591
rect 3629 9539 3681 9591
rect 3681 9539 3683 9591
rect 3627 9537 3683 9539
rect 3947 9591 4003 9593
rect 3947 9539 3949 9591
rect 3949 9539 4001 9591
rect 4001 9539 4003 9591
rect 3947 9537 4003 9539
rect 4257 9591 4313 9593
rect 4257 9539 4259 9591
rect 4259 9539 4311 9591
rect 4311 9539 4313 9591
rect 4257 9537 4313 9539
rect 4577 9591 4633 9593
rect 4577 9539 4579 9591
rect 4579 9539 4631 9591
rect 4631 9539 4633 9591
rect 4577 9537 4633 9539
rect 4897 9591 4953 9593
rect 4897 9539 4899 9591
rect 4899 9539 4951 9591
rect 4951 9539 4953 9591
rect 4897 9537 4953 9539
rect -1113 9167 -1057 9223
rect -4018 8726 -3962 8728
rect -3938 8726 -3882 8728
rect -4018 8674 -3988 8726
rect -3988 8674 -3976 8726
rect -3976 8674 -3962 8726
rect -3938 8674 -3924 8726
rect -3924 8674 -3912 8726
rect -3912 8674 -3882 8726
rect -4018 8672 -3962 8674
rect -3938 8672 -3882 8674
rect -3598 8726 -3542 8728
rect -3518 8726 -3462 8728
rect -3598 8674 -3568 8726
rect -3568 8674 -3556 8726
rect -3556 8674 -3542 8726
rect -3518 8674 -3504 8726
rect -3504 8674 -3492 8726
rect -3492 8674 -3462 8726
rect -3598 8672 -3542 8674
rect -3518 8672 -3462 8674
rect 1297 9047 1513 9263
rect 2347 9047 2563 9263
rect 227 8771 283 8773
rect 227 8719 229 8771
rect 229 8719 281 8771
rect 281 8719 283 8771
rect 227 8717 283 8719
rect 547 8771 603 8773
rect 547 8719 549 8771
rect 549 8719 601 8771
rect 601 8719 603 8771
rect 547 8717 603 8719
rect 857 8771 913 8773
rect 857 8719 859 8771
rect 859 8719 911 8771
rect 911 8719 913 8771
rect 857 8717 913 8719
rect 1177 8771 1233 8773
rect 1177 8719 1179 8771
rect 1179 8719 1231 8771
rect 1231 8719 1233 8771
rect 1177 8717 1233 8719
rect 1497 8771 1553 8773
rect 1497 8719 1499 8771
rect 1499 8719 1551 8771
rect 1551 8719 1553 8771
rect 1497 8717 1553 8719
rect 1807 8771 1863 8773
rect 1807 8719 1809 8771
rect 1809 8719 1861 8771
rect 1861 8719 1863 8771
rect 1807 8717 1863 8719
rect 2127 8771 2183 8773
rect 2127 8719 2129 8771
rect 2129 8719 2181 8771
rect 2181 8719 2183 8771
rect 2127 8717 2183 8719
rect 2447 8771 2503 8773
rect 2447 8719 2449 8771
rect 2449 8719 2501 8771
rect 2501 8719 2503 8771
rect 2447 8717 2503 8719
rect 2757 8771 2813 8773
rect 2757 8719 2759 8771
rect 2759 8719 2811 8771
rect 2811 8719 2813 8771
rect 2757 8717 2813 8719
rect 3077 8771 3133 8773
rect 3077 8719 3079 8771
rect 3079 8719 3131 8771
rect 3131 8719 3133 8771
rect 3077 8717 3133 8719
rect 3387 8771 3443 8773
rect 3387 8719 3389 8771
rect 3389 8719 3441 8771
rect 3441 8719 3443 8771
rect 3387 8717 3443 8719
rect 227 8561 283 8563
rect 227 8509 229 8561
rect 229 8509 281 8561
rect 281 8509 283 8561
rect 227 8507 283 8509
rect 547 8561 603 8563
rect 547 8509 549 8561
rect 549 8509 601 8561
rect 601 8509 603 8561
rect 547 8507 603 8509
rect 857 8561 913 8563
rect 857 8509 859 8561
rect 859 8509 911 8561
rect 911 8509 913 8561
rect 857 8507 913 8509
rect 1177 8561 1233 8563
rect 1177 8509 1179 8561
rect 1179 8509 1231 8561
rect 1231 8509 1233 8561
rect 1177 8507 1233 8509
rect 1497 8561 1553 8563
rect 1497 8509 1499 8561
rect 1499 8509 1551 8561
rect 1551 8509 1553 8561
rect 1497 8507 1553 8509
rect 1807 8561 1863 8563
rect 1807 8509 1809 8561
rect 1809 8509 1861 8561
rect 1861 8509 1863 8561
rect 1807 8507 1863 8509
rect 2127 8561 2183 8563
rect 2127 8509 2129 8561
rect 2129 8509 2181 8561
rect 2181 8509 2183 8561
rect 2127 8507 2183 8509
rect 2447 8561 2503 8563
rect 2447 8509 2449 8561
rect 2449 8509 2501 8561
rect 2501 8509 2503 8561
rect 2447 8507 2503 8509
rect 2757 8561 2813 8563
rect 2757 8509 2759 8561
rect 2759 8509 2811 8561
rect 2811 8509 2813 8561
rect 2757 8507 2813 8509
rect 3077 8561 3133 8563
rect 3077 8509 3079 8561
rect 3079 8509 3131 8561
rect 3131 8509 3133 8561
rect 3077 8507 3133 8509
rect 3387 8561 3443 8563
rect 3387 8509 3389 8561
rect 3389 8509 3441 8561
rect 3441 8509 3443 8561
rect 3387 8507 3443 8509
rect -148 8062 -92 8118
rect 387 8131 443 8133
rect 387 8079 389 8131
rect 389 8079 441 8131
rect 441 8079 443 8131
rect 387 8077 443 8079
rect 707 8131 763 8133
rect 707 8079 709 8131
rect 709 8079 761 8131
rect 761 8079 763 8131
rect 707 8077 763 8079
rect 1017 8131 1073 8133
rect 1017 8079 1019 8131
rect 1019 8079 1071 8131
rect 1071 8079 1073 8131
rect 1017 8077 1073 8079
rect 1337 8131 1393 8133
rect 1337 8079 1339 8131
rect 1339 8079 1391 8131
rect 1391 8079 1393 8131
rect 1337 8077 1393 8079
rect 1657 8131 1713 8133
rect 1657 8079 1659 8131
rect 1659 8079 1711 8131
rect 1711 8079 1713 8131
rect 1657 8077 1713 8079
rect 1967 8131 2023 8133
rect 1967 8079 1969 8131
rect 1969 8079 2021 8131
rect 2021 8079 2023 8131
rect 1967 8077 2023 8079
rect 2287 8131 2343 8133
rect 2287 8079 2289 8131
rect 2289 8079 2341 8131
rect 2341 8079 2343 8131
rect 2287 8077 2343 8079
rect 2597 8131 2653 8133
rect 2597 8079 2599 8131
rect 2599 8079 2651 8131
rect 2651 8079 2653 8131
rect 2597 8077 2653 8079
rect 2917 8131 2973 8133
rect 2917 8079 2919 8131
rect 2919 8079 2971 8131
rect 2971 8079 2973 8131
rect 2917 8077 2973 8079
rect 3237 8131 3293 8133
rect 3237 8079 3239 8131
rect 3239 8079 3291 8131
rect 3291 8079 3293 8131
rect 3237 8077 3293 8079
rect 3547 8131 3603 8133
rect 3547 8079 3549 8131
rect 3549 8079 3601 8131
rect 3601 8079 3603 8131
rect 3547 8077 3603 8079
rect 3912 8062 3968 8118
rect -148 7882 -92 7938
rect 387 7921 443 7923
rect 387 7869 389 7921
rect 389 7869 441 7921
rect 441 7869 443 7921
rect 387 7867 443 7869
rect 707 7921 763 7923
rect 707 7869 709 7921
rect 709 7869 761 7921
rect 761 7869 763 7921
rect 707 7867 763 7869
rect 1017 7921 1073 7923
rect 1017 7869 1019 7921
rect 1019 7869 1071 7921
rect 1071 7869 1073 7921
rect 1017 7867 1073 7869
rect 1337 7921 1393 7923
rect 1337 7869 1339 7921
rect 1339 7869 1391 7921
rect 1391 7869 1393 7921
rect 1337 7867 1393 7869
rect 1657 7921 1713 7923
rect 1657 7869 1659 7921
rect 1659 7869 1711 7921
rect 1711 7869 1713 7921
rect 1657 7867 1713 7869
rect 1967 7921 2023 7923
rect 1967 7869 1969 7921
rect 1969 7869 2021 7921
rect 2021 7869 2023 7921
rect 1967 7867 2023 7869
rect 2287 7921 2343 7923
rect 2287 7869 2289 7921
rect 2289 7869 2341 7921
rect 2341 7869 2343 7921
rect 2287 7867 2343 7869
rect 2597 7921 2653 7923
rect 2597 7869 2599 7921
rect 2599 7869 2651 7921
rect 2651 7869 2653 7921
rect 2597 7867 2653 7869
rect 2917 7921 2973 7923
rect 2917 7869 2919 7921
rect 2919 7869 2971 7921
rect 2971 7869 2973 7921
rect 2917 7867 2973 7869
rect 3237 7921 3293 7923
rect 3237 7869 3239 7921
rect 3239 7869 3291 7921
rect 3291 7869 3293 7921
rect 3237 7867 3293 7869
rect 3547 7921 3603 7923
rect 3547 7869 3549 7921
rect 3549 7869 3601 7921
rect 3601 7869 3603 7921
rect 3547 7867 3603 7869
rect 3912 7882 3968 7938
rect 1062 7442 1278 7658
rect 2562 7442 2778 7658
rect 227 7221 283 7223
rect 227 7169 229 7221
rect 229 7169 281 7221
rect 281 7169 283 7221
rect 227 7167 283 7169
rect 547 7221 603 7223
rect 547 7169 549 7221
rect 549 7169 601 7221
rect 601 7169 603 7221
rect 547 7167 603 7169
rect 857 7221 913 7223
rect 857 7169 859 7221
rect 859 7169 911 7221
rect 911 7169 913 7221
rect 857 7167 913 7169
rect 1177 7221 1233 7223
rect 1177 7169 1179 7221
rect 1179 7169 1231 7221
rect 1231 7169 1233 7221
rect 1177 7167 1233 7169
rect 1497 7221 1553 7223
rect 1497 7169 1499 7221
rect 1499 7169 1551 7221
rect 1551 7169 1553 7221
rect 1497 7167 1553 7169
rect 1807 7221 1863 7223
rect 1807 7169 1809 7221
rect 1809 7169 1861 7221
rect 1861 7169 1863 7221
rect 1807 7167 1863 7169
rect 2127 7221 2183 7223
rect 2127 7169 2129 7221
rect 2129 7169 2181 7221
rect 2181 7169 2183 7221
rect 2127 7167 2183 7169
rect 2437 7221 2493 7223
rect 2437 7169 2439 7221
rect 2439 7169 2491 7221
rect 2491 7169 2493 7221
rect 2437 7167 2493 7169
rect 2757 7221 2813 7223
rect 2757 7169 2759 7221
rect 2759 7169 2811 7221
rect 2811 7169 2813 7221
rect 2757 7167 2813 7169
rect 3077 7221 3133 7223
rect 3077 7169 3079 7221
rect 3079 7169 3131 7221
rect 3131 7169 3133 7221
rect 3077 7167 3133 7169
rect 3387 7221 3443 7223
rect 3387 7169 3389 7221
rect 3389 7169 3441 7221
rect 3441 7169 3443 7221
rect 3387 7167 3443 7169
rect 227 7011 283 7013
rect 227 6959 229 7011
rect 229 6959 281 7011
rect 281 6959 283 7011
rect 227 6957 283 6959
rect 547 7011 603 7013
rect 547 6959 549 7011
rect 549 6959 601 7011
rect 601 6959 603 7011
rect 547 6957 603 6959
rect 857 7011 913 7013
rect 857 6959 859 7011
rect 859 6959 911 7011
rect 911 6959 913 7011
rect 857 6957 913 6959
rect 1177 7011 1233 7013
rect 1177 6959 1179 7011
rect 1179 6959 1231 7011
rect 1231 6959 1233 7011
rect 1177 6957 1233 6959
rect 1497 7011 1553 7013
rect 1497 6959 1499 7011
rect 1499 6959 1551 7011
rect 1551 6959 1553 7011
rect 1497 6957 1553 6959
rect 1807 7011 1863 7013
rect 1807 6959 1809 7011
rect 1809 6959 1861 7011
rect 1861 6959 1863 7011
rect 1807 6957 1863 6959
rect 2127 7011 2183 7013
rect 2127 6959 2129 7011
rect 2129 6959 2181 7011
rect 2181 6959 2183 7011
rect 2127 6957 2183 6959
rect 2437 7011 2493 7013
rect 2437 6959 2439 7011
rect 2439 6959 2491 7011
rect 2491 6959 2493 7011
rect 2437 6957 2493 6959
rect 2757 7011 2813 7013
rect 2757 6959 2759 7011
rect 2759 6959 2811 7011
rect 2811 6959 2813 7011
rect 2757 6957 2813 6959
rect 3077 7011 3133 7013
rect 3077 6959 3079 7011
rect 3079 6959 3131 7011
rect 3131 6959 3133 7011
rect 3077 6957 3133 6959
rect 3387 7011 3443 7013
rect 3387 6959 3389 7011
rect 3389 6959 3441 7011
rect 3441 6959 3443 7011
rect 3387 6957 3443 6959
rect 387 6591 443 6593
rect 387 6539 389 6591
rect 389 6539 441 6591
rect 441 6539 443 6591
rect 387 6537 443 6539
rect 707 6591 763 6593
rect 707 6539 709 6591
rect 709 6539 761 6591
rect 761 6539 763 6591
rect 707 6537 763 6539
rect 387 6381 443 6383
rect 387 6329 389 6381
rect 389 6329 441 6381
rect 441 6329 443 6381
rect 387 6327 443 6329
rect 1017 6591 1073 6593
rect 1017 6539 1019 6591
rect 1019 6539 1071 6591
rect 1071 6539 1073 6591
rect 1017 6537 1073 6539
rect 1337 6591 1393 6593
rect 1337 6539 1339 6591
rect 1339 6539 1391 6591
rect 1391 6539 1393 6591
rect 1337 6537 1393 6539
rect 1647 6591 1703 6593
rect 1647 6539 1649 6591
rect 1649 6539 1701 6591
rect 1701 6539 1703 6591
rect 1647 6537 1703 6539
rect 1967 6591 2023 6593
rect 1967 6539 1969 6591
rect 1969 6539 2021 6591
rect 2021 6539 2023 6591
rect 1967 6537 2023 6539
rect 2287 6591 2343 6593
rect 2287 6539 2289 6591
rect 2289 6539 2341 6591
rect 2341 6539 2343 6591
rect 2287 6537 2343 6539
rect 2597 6591 2653 6593
rect 2597 6539 2599 6591
rect 2599 6539 2651 6591
rect 2651 6539 2653 6591
rect 2597 6537 2653 6539
rect 2917 6591 2973 6593
rect 2917 6539 2919 6591
rect 2919 6539 2971 6591
rect 2971 6539 2973 6591
rect 2917 6537 2973 6539
rect 3227 6591 3283 6593
rect 3227 6539 3229 6591
rect 3229 6539 3281 6591
rect 3281 6539 3283 6591
rect 3227 6537 3283 6539
rect 707 6381 763 6383
rect 707 6329 709 6381
rect 709 6329 761 6381
rect 761 6329 763 6381
rect 707 6327 763 6329
rect -148 5572 -92 5628
rect -148 5352 -92 5408
rect 92 5012 148 5068
rect 92 4792 148 4848
rect 92 4052 148 4108
rect 92 3832 148 3888
rect -1113 2557 -1057 2613
rect -1113 2397 -1057 2453
rect 1017 6381 1073 6383
rect 1017 6329 1019 6381
rect 1019 6329 1071 6381
rect 1071 6329 1073 6381
rect 1017 6327 1073 6329
rect 1337 6381 1393 6383
rect 1337 6329 1339 6381
rect 1339 6329 1391 6381
rect 1391 6329 1393 6381
rect 1337 6327 1393 6329
rect 1647 6381 1703 6383
rect 1647 6329 1649 6381
rect 1649 6329 1701 6381
rect 1701 6329 1703 6381
rect 1647 6327 1703 6329
rect 1967 6381 2023 6383
rect 1967 6329 1969 6381
rect 1969 6329 2021 6381
rect 2021 6329 2023 6381
rect 1967 6327 2023 6329
rect 2287 6381 2343 6383
rect 2287 6329 2289 6381
rect 2289 6329 2341 6381
rect 2341 6329 2343 6381
rect 2287 6327 2343 6329
rect 2597 6381 2653 6383
rect 2597 6329 2599 6381
rect 2599 6329 2651 6381
rect 2651 6329 2653 6381
rect 2597 6327 2653 6329
rect 2917 6381 2973 6383
rect 2917 6329 2919 6381
rect 2919 6329 2971 6381
rect 2971 6329 2973 6381
rect 2917 6327 2973 6329
rect 3547 6591 3603 6593
rect 3547 6539 3549 6591
rect 3549 6539 3601 6591
rect 3601 6539 3603 6591
rect 3547 6537 3603 6539
rect 3227 6381 3283 6383
rect 3227 6329 3229 6381
rect 3229 6329 3281 6381
rect 3281 6329 3283 6381
rect 3227 6327 3283 6329
rect 1327 5661 1383 5663
rect 1327 5609 1329 5661
rect 1329 5609 1381 5661
rect 1381 5609 1383 5661
rect 1327 5607 1383 5609
rect 1647 5661 1703 5663
rect 1647 5609 1649 5661
rect 1649 5609 1701 5661
rect 1701 5609 1703 5661
rect 1647 5607 1703 5609
rect 1957 5661 2013 5663
rect 1957 5609 1959 5661
rect 1959 5609 2011 5661
rect 2011 5609 2013 5661
rect 1957 5607 2013 5609
rect 2277 5661 2333 5663
rect 2277 5609 2279 5661
rect 2279 5609 2331 5661
rect 2331 5609 2333 5661
rect 2277 5607 2333 5609
rect 1327 5371 1383 5373
rect 1327 5319 1329 5371
rect 1329 5319 1381 5371
rect 1381 5319 1383 5371
rect 1327 5317 1383 5319
rect 1647 5371 1703 5373
rect 1647 5319 1649 5371
rect 1649 5319 1701 5371
rect 1701 5319 1703 5371
rect 1647 5317 1703 5319
rect 1957 5371 2013 5373
rect 1957 5319 1959 5371
rect 1959 5319 2011 5371
rect 2011 5319 2013 5371
rect 1957 5317 2013 5319
rect 2277 5371 2333 5373
rect 2277 5319 2279 5371
rect 2279 5319 2331 5371
rect 2331 5319 2333 5371
rect 2277 5317 2333 5319
rect 1487 5101 1543 5103
rect 1487 5049 1489 5101
rect 1489 5049 1541 5101
rect 1541 5049 1543 5101
rect 1487 5047 1543 5049
rect 1797 5101 1853 5103
rect 1797 5049 1799 5101
rect 1799 5049 1851 5101
rect 1851 5049 1853 5101
rect 1797 5047 1853 5049
rect 2117 5101 2173 5103
rect 2117 5049 2119 5101
rect 2119 5049 2171 5101
rect 2171 5049 2173 5101
rect 2117 5047 2173 5049
rect 2437 5101 2493 5103
rect 2437 5049 2439 5101
rect 2439 5049 2491 5101
rect 2491 5049 2493 5101
rect 2437 5047 2493 5049
rect 1487 4811 1543 4813
rect 1487 4759 1489 4811
rect 1489 4759 1541 4811
rect 1541 4759 1543 4811
rect 1487 4757 1543 4759
rect 1797 4811 1853 4813
rect 1797 4759 1799 4811
rect 1799 4759 1851 4811
rect 1851 4759 1853 4811
rect 1797 4757 1853 4759
rect 2117 4811 2173 4813
rect 2117 4759 2119 4811
rect 2119 4759 2171 4811
rect 2171 4759 2173 4811
rect 2117 4757 2173 4759
rect 2437 4811 2493 4813
rect 2437 4759 2439 4811
rect 2439 4759 2491 4811
rect 2491 4759 2493 4811
rect 2437 4757 2493 4759
rect 1802 4342 2018 4558
rect 1327 4141 1383 4143
rect 1327 4089 1329 4141
rect 1329 4089 1381 4141
rect 1381 4089 1383 4141
rect 1327 4087 1383 4089
rect 1647 4141 1703 4143
rect 1647 4089 1649 4141
rect 1649 4089 1701 4141
rect 1701 4089 1703 4141
rect 1647 4087 1703 4089
rect 1957 4141 2013 4143
rect 1957 4089 1959 4141
rect 1959 4089 2011 4141
rect 2011 4089 2013 4141
rect 1957 4087 2013 4089
rect 2277 4141 2333 4143
rect 2277 4089 2279 4141
rect 2279 4089 2331 4141
rect 2331 4089 2333 4141
rect 2277 4087 2333 4089
rect 1327 3851 1383 3853
rect 1327 3799 1329 3851
rect 1329 3799 1381 3851
rect 1381 3799 1383 3851
rect 1327 3797 1383 3799
rect 1647 3851 1703 3853
rect 1647 3799 1649 3851
rect 1649 3799 1701 3851
rect 1701 3799 1703 3851
rect 1647 3797 1703 3799
rect 1957 3851 2013 3853
rect 1957 3799 1959 3851
rect 1959 3799 2011 3851
rect 2011 3799 2013 3851
rect 1957 3797 2013 3799
rect 2277 3851 2333 3853
rect 2277 3799 2279 3851
rect 2279 3799 2331 3851
rect 2331 3799 2333 3851
rect 2277 3797 2333 3799
rect 707 3507 763 3563
rect 1487 3581 1543 3583
rect 1487 3529 1489 3581
rect 1489 3529 1541 3581
rect 1541 3529 1543 3581
rect 1487 3527 1543 3529
rect 1797 3581 1853 3583
rect 1797 3529 1799 3581
rect 1799 3529 1851 3581
rect 1851 3529 1853 3581
rect 1797 3527 1853 3529
rect 2117 3581 2173 3583
rect 2117 3529 2119 3581
rect 2119 3529 2171 3581
rect 2171 3529 2173 3581
rect 2117 3527 2173 3529
rect 2437 3581 2493 3583
rect 2437 3529 2439 3581
rect 2439 3529 2491 3581
rect 2491 3529 2493 3581
rect 2437 3527 2493 3529
rect 3547 6381 3603 6383
rect 3547 6329 3549 6381
rect 3549 6329 3601 6381
rect 3601 6329 3603 6381
rect 3547 6327 3603 6329
rect 3912 5572 3968 5628
rect 3912 5352 3968 5408
rect 4897 9167 4953 9223
rect 707 3257 763 3313
rect 3227 3507 3283 3563
rect 1487 3291 1543 3293
rect 1487 3239 1489 3291
rect 1489 3239 1541 3291
rect 1541 3239 1543 3291
rect 1487 3237 1543 3239
rect 1797 3291 1853 3293
rect 1797 3239 1799 3291
rect 1799 3239 1851 3291
rect 1851 3239 1853 3291
rect 1797 3237 1853 3239
rect 2117 3291 2173 3293
rect 2117 3239 2119 3291
rect 2119 3239 2171 3291
rect 2171 3239 2173 3291
rect 2117 3237 2173 3239
rect 2437 3291 2493 3293
rect 2437 3239 2439 3291
rect 2439 3239 2491 3291
rect 2491 3239 2493 3291
rect 2437 3237 2493 3239
rect 3227 3257 3283 3313
rect 3672 5012 3728 5068
rect 3672 4792 3728 4848
rect 3672 4052 3728 4108
rect 3672 3832 3728 3888
rect 1802 2822 2018 3038
rect 337 2621 393 2623
rect 337 2569 339 2621
rect 339 2569 391 2621
rect 391 2569 393 2621
rect 337 2567 393 2569
rect 857 2621 913 2623
rect 857 2569 859 2621
rect 859 2569 911 2621
rect 911 2569 913 2621
rect 857 2567 913 2569
rect 1367 2621 1423 2623
rect 1367 2569 1369 2621
rect 1369 2569 1421 2621
rect 1421 2569 1423 2621
rect 1367 2567 1423 2569
rect 1887 2621 1943 2623
rect 1887 2569 1889 2621
rect 1889 2569 1941 2621
rect 1941 2569 1943 2621
rect 1887 2567 1943 2569
rect 2397 2621 2453 2623
rect 2397 2569 2399 2621
rect 2399 2569 2451 2621
rect 2451 2569 2453 2621
rect 2397 2567 2453 2569
rect 2917 2621 2973 2623
rect 2917 2569 2919 2621
rect 2919 2569 2971 2621
rect 2971 2569 2973 2621
rect 2917 2567 2973 2569
rect 3437 2621 3493 2623
rect 3437 2569 3439 2621
rect 3439 2569 3491 2621
rect 3491 2569 3493 2621
rect 3437 2567 3493 2569
rect 337 2441 393 2443
rect 337 2389 339 2441
rect 339 2389 391 2441
rect 391 2389 393 2441
rect 337 2387 393 2389
rect 857 2441 913 2443
rect 857 2389 859 2441
rect 859 2389 911 2441
rect 911 2389 913 2441
rect 857 2387 913 2389
rect 1367 2441 1423 2443
rect 1367 2389 1369 2441
rect 1369 2389 1421 2441
rect 1421 2389 1423 2441
rect 1367 2387 1423 2389
rect 1887 2441 1943 2443
rect 1887 2389 1889 2441
rect 1889 2389 1941 2441
rect 1941 2389 1943 2441
rect 1887 2387 1943 2389
rect 2397 2441 2453 2443
rect 2397 2389 2399 2441
rect 2399 2389 2451 2441
rect 2451 2389 2453 2441
rect 2397 2387 2453 2389
rect 2917 2441 2973 2443
rect 2917 2389 2919 2441
rect 2919 2389 2971 2441
rect 2971 2389 2973 2441
rect 2917 2387 2973 2389
rect 3437 2441 3493 2443
rect 3437 2389 3439 2441
rect 3439 2389 3491 2441
rect 3491 2389 3493 2441
rect 3437 2387 3493 2389
rect 597 1951 653 1953
rect 597 1899 599 1951
rect 599 1899 651 1951
rect 651 1899 653 1951
rect 597 1897 653 1899
rect 1107 1951 1163 1953
rect 1107 1899 1109 1951
rect 1109 1899 1161 1951
rect 1161 1899 1163 1951
rect 1107 1897 1163 1899
rect 1627 1951 1683 1953
rect 1627 1899 1629 1951
rect 1629 1899 1681 1951
rect 1681 1899 1683 1951
rect 1627 1897 1683 1899
rect 2147 1951 2203 1953
rect 2147 1899 2149 1951
rect 2149 1899 2201 1951
rect 2201 1899 2203 1951
rect 2147 1897 2203 1899
rect 2657 1951 2713 1953
rect 2657 1899 2659 1951
rect 2659 1899 2711 1951
rect 2711 1899 2713 1951
rect 2657 1897 2713 1899
rect 3177 1951 3233 1953
rect 3177 1899 3179 1951
rect 3179 1899 3231 1951
rect 3231 1899 3233 1951
rect 3177 1897 3233 1899
rect 597 1771 653 1773
rect 597 1719 599 1771
rect 599 1719 651 1771
rect 651 1719 653 1771
rect 597 1717 653 1719
rect 1107 1771 1163 1773
rect 1107 1719 1109 1771
rect 1109 1719 1161 1771
rect 1161 1719 1163 1771
rect 1107 1717 1163 1719
rect 1627 1771 1683 1773
rect 1627 1719 1629 1771
rect 1629 1719 1681 1771
rect 1681 1719 1683 1771
rect 1627 1717 1683 1719
rect 2147 1771 2203 1773
rect 2147 1719 2149 1771
rect 2149 1719 2201 1771
rect 2201 1719 2203 1771
rect 2147 1717 2203 1719
rect 2657 1771 2713 1773
rect 2657 1719 2659 1771
rect 2659 1719 2711 1771
rect 2711 1719 2713 1771
rect 2657 1717 2713 1719
rect 3177 1771 3233 1773
rect 3177 1719 3179 1771
rect 3179 1719 3231 1771
rect 3231 1719 3233 1771
rect 3177 1717 3233 1719
rect 1807 1307 2023 1523
rect 77 1101 133 1103
rect 77 1049 79 1101
rect 79 1049 131 1101
rect 131 1049 133 1101
rect 77 1047 133 1049
rect 597 1101 653 1103
rect 597 1049 599 1101
rect 599 1049 651 1101
rect 651 1049 653 1101
rect 597 1047 653 1049
rect 1107 1101 1163 1103
rect 1107 1049 1109 1101
rect 1109 1049 1161 1101
rect 1161 1049 1163 1101
rect 1107 1047 1163 1049
rect 1627 1101 1683 1103
rect 1627 1049 1629 1101
rect 1629 1049 1681 1101
rect 1681 1049 1683 1101
rect 1627 1047 1683 1049
rect 2137 1101 2193 1103
rect 2137 1049 2139 1101
rect 2139 1049 2191 1101
rect 2191 1049 2193 1101
rect 2137 1047 2193 1049
rect 2657 1101 2713 1103
rect 2657 1049 2659 1101
rect 2659 1049 2711 1101
rect 2711 1049 2713 1101
rect 2657 1047 2713 1049
rect 3177 1101 3233 1103
rect 3177 1049 3179 1101
rect 3179 1049 3231 1101
rect 3231 1049 3233 1101
rect 3177 1047 3233 1049
rect 3687 1101 3743 1103
rect 3687 1049 3689 1101
rect 3689 1049 3741 1101
rect 3741 1049 3743 1101
rect 3687 1047 3743 1049
rect 77 921 133 923
rect 77 869 79 921
rect 79 869 131 921
rect 131 869 133 921
rect 77 867 133 869
rect 597 921 653 923
rect 597 869 599 921
rect 599 869 651 921
rect 651 869 653 921
rect 597 867 653 869
rect 1107 921 1163 923
rect 1107 869 1109 921
rect 1109 869 1161 921
rect 1161 869 1163 921
rect 1107 867 1163 869
rect 1627 921 1683 923
rect 1627 869 1629 921
rect 1629 869 1681 921
rect 1681 869 1683 921
rect 1627 867 1683 869
rect 2137 921 2193 923
rect 2137 869 2139 921
rect 2139 869 2191 921
rect 2191 869 2193 921
rect 2137 867 2193 869
rect 2657 921 2713 923
rect 2657 869 2659 921
rect 2659 869 2711 921
rect 2711 869 2713 921
rect 2657 867 2713 869
rect 3177 921 3233 923
rect 3177 869 3179 921
rect 3179 869 3231 921
rect 3231 869 3233 921
rect 3177 867 3233 869
rect 3687 921 3743 923
rect 3687 869 3689 921
rect 3689 869 3741 921
rect 3741 869 3743 921
rect 3687 867 3743 869
rect 7232 8726 7288 8728
rect 7312 8726 7368 8728
rect 7232 8674 7262 8726
rect 7262 8674 7274 8726
rect 7274 8674 7288 8726
rect 7312 8674 7326 8726
rect 7326 8674 7338 8726
rect 7338 8674 7368 8726
rect 7232 8672 7288 8674
rect 7312 8672 7368 8674
rect 7652 8726 7708 8728
rect 7732 8726 7788 8728
rect 7652 8674 7682 8726
rect 7682 8674 7694 8726
rect 7694 8674 7708 8726
rect 7732 8674 7746 8726
rect 7746 8674 7758 8726
rect 7758 8674 7788 8726
rect 7652 8672 7708 8674
rect 7732 8672 7788 8674
rect 4897 2557 4953 2613
rect 4897 2397 4953 2453
rect 337 431 393 433
rect 337 379 339 431
rect 339 379 391 431
rect 391 379 393 431
rect 337 377 393 379
rect 847 431 903 433
rect 847 379 849 431
rect 849 379 901 431
rect 901 379 903 431
rect 847 377 903 379
rect 1367 431 1423 433
rect 1367 379 1369 431
rect 1369 379 1421 431
rect 1421 379 1423 431
rect 1367 377 1423 379
rect 1887 431 1943 433
rect 1887 379 1889 431
rect 1889 379 1941 431
rect 1941 379 1943 431
rect 1887 377 1943 379
rect 2397 431 2453 433
rect 2397 379 2399 431
rect 2399 379 2451 431
rect 2451 379 2453 431
rect 2397 377 2453 379
rect 2917 431 2973 433
rect 2917 379 2919 431
rect 2919 379 2971 431
rect 2971 379 2973 431
rect 2917 377 2973 379
rect 3427 431 3483 433
rect 3427 379 3429 431
rect 3429 379 3481 431
rect 3481 379 3483 431
rect 3427 377 3483 379
rect 337 251 393 253
rect 337 199 339 251
rect 339 199 391 251
rect 391 199 393 251
rect 337 197 393 199
rect 847 251 903 253
rect 847 199 849 251
rect 849 199 901 251
rect 901 199 903 251
rect 847 197 903 199
rect 1367 251 1423 253
rect 1367 199 1369 251
rect 1369 199 1421 251
rect 1421 199 1423 251
rect 1367 197 1423 199
rect 1887 251 1943 253
rect 1887 199 1889 251
rect 1889 199 1941 251
rect 1941 199 1943 251
rect 1887 197 1943 199
rect 2397 251 2453 253
rect 2397 199 2399 251
rect 2399 199 2451 251
rect 2451 199 2453 251
rect 2397 197 2453 199
rect 2917 251 2973 253
rect 2917 199 2919 251
rect 2919 199 2971 251
rect 2971 199 2973 251
rect 2917 197 2973 199
rect 3427 251 3483 253
rect 3427 199 3429 251
rect 3429 199 3481 251
rect 3481 199 3483 251
rect 3427 197 3483 199
rect 1807 -223 2023 -7
<< metal3 >>
rect 1260 10907 1550 10935
rect 1260 10683 1293 10907
rect 1517 10683 1550 10907
rect 1260 10655 1550 10683
rect 2310 10907 2600 10935
rect 2310 10683 2343 10907
rect 2567 10683 2600 10907
rect 2310 10655 2600 10683
rect -1280 10455 5110 10460
rect -1290 10443 5120 10455
rect -1290 10387 -1273 10443
rect -1217 10387 -953 10443
rect -897 10417 -643 10443
rect -897 10387 -887 10417
rect -1290 10375 -887 10387
rect -5940 10207 -5720 10230
rect -1280 10215 -887 10375
rect -5940 10143 -5807 10207
rect -5743 10143 -5720 10207
rect -5940 10097 -5720 10143
rect -1290 10203 -887 10215
rect -1290 10147 -1273 10203
rect -1217 10147 -953 10203
rect -897 10193 -887 10203
rect -663 10387 -643 10417
rect -587 10387 -323 10443
rect -267 10387 -13 10443
rect 43 10387 307 10443
rect 363 10387 627 10443
rect 683 10387 937 10443
rect 993 10407 1257 10443
rect 993 10387 1013 10407
rect -663 10203 1013 10387
rect -663 10193 -643 10203
rect -897 10147 -643 10193
rect -587 10147 -323 10203
rect -267 10147 -13 10203
rect 43 10147 307 10203
rect 363 10147 627 10203
rect 683 10147 937 10203
rect 993 10183 1013 10203
rect 1237 10387 1257 10407
rect 1313 10387 1577 10443
rect 1633 10387 1887 10443
rect 1943 10387 2207 10443
rect 2263 10387 2517 10443
rect 2573 10407 2837 10443
rect 2573 10387 2593 10407
rect 1237 10203 2593 10387
rect 1237 10183 1257 10203
rect 993 10147 1257 10183
rect 1313 10147 1577 10203
rect 1633 10147 1887 10203
rect 1943 10147 2207 10203
rect 2263 10147 2517 10203
rect 2573 10183 2593 10203
rect 2817 10387 2837 10407
rect 2893 10387 3157 10443
rect 3213 10387 3467 10443
rect 3523 10387 3787 10443
rect 3843 10387 4097 10443
rect 4153 10387 4417 10443
rect 4473 10407 4737 10443
rect 4473 10387 4493 10407
rect 2817 10203 4493 10387
rect 2817 10183 2837 10203
rect 2573 10147 2837 10183
rect 2893 10147 3157 10203
rect 3213 10147 3467 10203
rect 3523 10147 3787 10203
rect 3843 10147 4097 10203
rect 4153 10147 4417 10203
rect 4473 10183 4493 10203
rect 4717 10387 4737 10407
rect 4793 10387 5047 10443
rect 5103 10387 5120 10443
rect 4717 10375 5120 10387
rect 4717 10215 5110 10375
rect 4717 10203 5120 10215
rect 4717 10183 4737 10203
rect 4473 10147 4737 10183
rect 4793 10147 5047 10203
rect 5103 10147 5120 10203
rect -1290 10135 5120 10147
rect 9560 10207 9780 10230
rect 9560 10143 9583 10207
rect 9647 10143 9780 10207
rect -1280 10130 5110 10135
rect -5940 10033 -5917 10097
rect -5853 10033 -5720 10097
rect -5940 10010 -5720 10033
rect 9560 10097 9780 10143
rect 9560 10033 9693 10097
rect 9757 10033 9780 10097
rect 9560 10010 9780 10033
rect -1280 9833 5110 9850
rect -1280 9777 -1113 9833
rect -1057 9777 -803 9833
rect -747 9777 -483 9833
rect -427 9777 -163 9833
rect -107 9777 147 9833
rect 203 9777 467 9833
rect 523 9777 777 9833
rect 833 9777 1097 9833
rect 1153 9777 1417 9833
rect 1473 9777 1727 9833
rect 1783 9777 2047 9833
rect 2103 9777 2367 9833
rect 2423 9777 2677 9833
rect 2733 9777 2997 9833
rect 3053 9777 3307 9833
rect 3363 9777 3627 9833
rect 3683 9777 3947 9833
rect 4003 9777 4257 9833
rect 4313 9777 4577 9833
rect 4633 9777 4897 9833
rect 4953 9777 5110 9833
rect -1280 9593 5110 9777
rect -1280 9537 -1113 9593
rect -1057 9537 -803 9593
rect -747 9537 -483 9593
rect -427 9537 -163 9593
rect -107 9537 147 9593
rect 203 9537 467 9593
rect 523 9537 777 9593
rect 833 9537 1097 9593
rect 1153 9537 1417 9593
rect 1473 9537 1727 9593
rect 1783 9537 2047 9593
rect 2103 9537 2367 9593
rect 2423 9537 2677 9593
rect 2733 9537 2997 9593
rect 3053 9537 3307 9593
rect 3363 9537 3627 9593
rect 3683 9537 3947 9593
rect 4003 9537 4257 9593
rect 4313 9537 4577 9593
rect 4633 9537 4897 9593
rect 4953 9537 5110 9593
rect -1280 9520 5110 9537
rect -2050 9232 -1020 9270
rect -2050 9168 -2017 9232
rect -1953 9168 -1827 9232
rect -1763 9223 -1020 9232
rect -1763 9168 -1113 9223
rect -2050 9167 -1113 9168
rect -1057 9167 -1020 9223
rect -2050 9130 -1020 9167
rect 1260 9267 1550 9295
rect 1260 9043 1293 9267
rect 1517 9043 1550 9267
rect 1260 9015 1550 9043
rect 2310 9267 2600 9295
rect 2310 9043 2343 9267
rect 2567 9043 2600 9267
rect 4860 9232 5880 9270
rect 4860 9223 5593 9232
rect 4860 9167 4897 9223
rect 4953 9168 5593 9223
rect 5657 9168 5783 9232
rect 5847 9168 5880 9232
rect 4953 9167 5880 9168
rect 4860 9130 5880 9167
rect 2310 9015 2600 9043
rect 220 8785 3610 8790
rect 210 8773 3610 8785
rect -4050 8732 -3850 8755
rect -4050 8668 -4022 8732
rect -3958 8668 -3942 8732
rect -3878 8668 -3850 8732
rect -4050 8645 -3850 8668
rect -3630 8732 -3430 8755
rect -3630 8668 -3602 8732
rect -3538 8668 -3522 8732
rect -3458 8668 -3430 8732
rect 210 8717 227 8773
rect 283 8717 547 8773
rect 603 8752 857 8773
rect 603 8717 618 8752
rect 210 8705 618 8717
rect -3630 8645 -3430 8668
rect 220 8575 618 8705
rect 210 8563 618 8575
rect 210 8507 227 8563
rect 283 8507 547 8563
rect 603 8528 618 8563
rect 842 8717 857 8752
rect 913 8717 1177 8773
rect 1233 8717 1497 8773
rect 1553 8717 1807 8773
rect 1863 8752 2127 8773
rect 1863 8717 1888 8752
rect 842 8563 1888 8717
rect 842 8528 857 8563
rect 603 8507 857 8528
rect 913 8507 1177 8563
rect 1233 8507 1497 8563
rect 1553 8507 1807 8563
rect 1863 8528 1888 8563
rect 2112 8717 2127 8752
rect 2183 8717 2447 8773
rect 2503 8717 2757 8773
rect 2813 8717 3077 8773
rect 3133 8752 3387 8773
rect 3133 8717 3148 8752
rect 2112 8563 3148 8717
rect 2112 8528 2127 8563
rect 1863 8507 2127 8528
rect 2183 8507 2447 8563
rect 2503 8507 2757 8563
rect 2813 8507 3077 8563
rect 3133 8528 3148 8563
rect 3372 8717 3387 8752
rect 3443 8717 3610 8773
rect 3372 8563 3610 8717
rect 7200 8732 7400 8755
rect 7200 8668 7228 8732
rect 7292 8668 7308 8732
rect 7372 8668 7400 8732
rect 7200 8645 7400 8668
rect 7620 8732 7820 8755
rect 7620 8668 7648 8732
rect 7712 8668 7728 8732
rect 7792 8668 7820 8732
rect 7620 8645 7820 8668
rect 3372 8528 3387 8563
rect 3133 8507 3387 8528
rect 3443 8507 3610 8563
rect 210 8495 3610 8507
rect 220 8490 3610 8495
rect -200 8133 4020 8150
rect -200 8118 387 8133
rect -200 8062 -148 8118
rect -92 8077 387 8118
rect 443 8077 707 8133
rect 763 8077 1017 8133
rect 1073 8077 1337 8133
rect 1393 8077 1657 8133
rect 1713 8077 1967 8133
rect 2023 8077 2287 8133
rect 2343 8077 2597 8133
rect 2653 8077 2917 8133
rect 2973 8077 3237 8133
rect 3293 8077 3547 8133
rect 3603 8118 4020 8133
rect 3603 8077 3912 8118
rect -92 8062 3912 8077
rect 3968 8062 4020 8118
rect -200 7938 4020 8062
rect -200 7882 -148 7938
rect -92 7923 3912 7938
rect -92 7882 387 7923
rect -200 7867 387 7882
rect 443 7867 707 7923
rect 763 7867 1017 7923
rect 1073 7867 1337 7923
rect 1393 7867 1657 7923
rect 1713 7867 1967 7923
rect 2023 7867 2287 7923
rect 2343 7867 2597 7923
rect 2653 7867 2917 7923
rect 2973 7867 3237 7923
rect 3293 7867 3547 7923
rect 3603 7882 3912 7923
rect 3968 7882 4020 7938
rect 3603 7867 4020 7882
rect -200 7850 4020 7867
rect 1030 7662 1310 7685
rect 1030 7438 1058 7662
rect 1282 7438 1310 7662
rect 1030 7415 1310 7438
rect 2530 7662 2810 7685
rect 2530 7438 2558 7662
rect 2782 7438 2810 7662
rect 2530 7415 2810 7438
rect 220 7235 3610 7240
rect 210 7223 3610 7235
rect 210 7167 227 7223
rect 283 7167 547 7223
rect 603 7202 857 7223
rect 603 7167 618 7202
rect 210 7155 618 7167
rect 220 7025 618 7155
rect 210 7013 618 7025
rect 210 6957 227 7013
rect 283 6957 547 7013
rect 603 6978 618 7013
rect 842 7167 857 7202
rect 913 7167 1177 7223
rect 1233 7167 1497 7223
rect 1553 7167 1807 7223
rect 1863 7202 2127 7223
rect 1863 7167 1888 7202
rect 842 7013 1888 7167
rect 842 6978 857 7013
rect 603 6957 857 6978
rect 913 6957 1177 7013
rect 1233 6957 1497 7013
rect 1553 6957 1807 7013
rect 1863 6978 1888 7013
rect 2112 7167 2127 7202
rect 2183 7167 2437 7223
rect 2493 7167 2757 7223
rect 2813 7167 3077 7223
rect 3133 7202 3387 7223
rect 3133 7167 3148 7202
rect 2112 7013 3148 7167
rect 2112 6978 2127 7013
rect 1863 6957 2127 6978
rect 2183 6957 2437 7013
rect 2493 6957 2757 7013
rect 2813 6957 3077 7013
rect 3133 6978 3148 7013
rect 3372 7167 3387 7202
rect 3443 7167 3610 7223
rect 3372 7013 3610 7167
rect 3372 6978 3387 7013
rect 3133 6957 3387 6978
rect 3443 6957 3610 7013
rect 210 6945 3610 6957
rect 220 6940 3610 6945
rect 220 6605 3610 6610
rect 220 6593 3620 6605
rect 220 6537 387 6593
rect 443 6537 707 6593
rect 763 6537 1017 6593
rect 1073 6537 1337 6593
rect 1393 6537 1647 6593
rect 1703 6537 1967 6593
rect 2023 6537 2287 6593
rect 2343 6537 2597 6593
rect 2653 6537 2917 6593
rect 2973 6537 3227 6593
rect 3283 6537 3547 6593
rect 3603 6537 3620 6593
rect 220 6525 3620 6537
rect 220 6395 3610 6525
rect 220 6383 3620 6395
rect 220 6327 387 6383
rect 443 6327 707 6383
rect 763 6327 1017 6383
rect 1073 6327 1337 6383
rect 1393 6327 1647 6383
rect 1703 6327 1967 6383
rect 2023 6327 2287 6383
rect 2343 6327 2597 6383
rect 2653 6327 2917 6383
rect 2973 6327 3227 6383
rect 3283 6327 3547 6383
rect 3603 6327 3620 6383
rect 220 6315 3620 6327
rect 220 6310 3610 6315
rect -200 5663 4020 5680
rect -200 5628 1327 5663
rect -200 5572 -148 5628
rect -92 5607 1327 5628
rect 1383 5607 1647 5663
rect 1703 5607 1957 5663
rect 2013 5607 2277 5663
rect 2333 5628 4020 5663
rect 2333 5607 3912 5628
rect -92 5572 3912 5607
rect 3968 5572 4020 5628
rect -200 5408 4020 5572
rect -200 5352 -148 5408
rect -92 5373 3912 5408
rect -92 5352 1327 5373
rect -200 5317 1327 5352
rect 1383 5317 1647 5373
rect 1703 5317 1957 5373
rect 2013 5317 2277 5373
rect 2333 5352 3912 5373
rect 3968 5352 4020 5408
rect 2333 5317 4020 5352
rect -200 5300 4020 5317
rect 40 5103 3780 5120
rect 40 5068 1487 5103
rect 40 5012 92 5068
rect 148 5047 1487 5068
rect 1543 5047 1797 5103
rect 1853 5047 2117 5103
rect 2173 5047 2437 5103
rect 2493 5068 3780 5103
rect 2493 5047 3672 5068
rect 148 5012 3672 5047
rect 3728 5012 3780 5068
rect 40 4848 3780 5012
rect 40 4792 92 4848
rect 148 4813 3672 4848
rect 148 4792 1487 4813
rect 40 4757 1487 4792
rect 1543 4757 1797 4813
rect 1853 4757 2117 4813
rect 2173 4757 2437 4813
rect 2493 4792 3672 4813
rect 3728 4792 3780 4848
rect 2493 4757 3780 4792
rect 40 4740 3780 4757
rect 1770 4562 2050 4585
rect 1770 4338 1798 4562
rect 2022 4338 2050 4562
rect 1770 4315 2050 4338
rect 40 4143 3780 4160
rect 40 4108 1327 4143
rect 40 4052 92 4108
rect 148 4087 1327 4108
rect 1383 4087 1647 4143
rect 1703 4087 1957 4143
rect 2013 4087 2277 4143
rect 2333 4108 3780 4143
rect 2333 4087 3672 4108
rect 148 4052 3672 4087
rect 3728 4052 3780 4108
rect 40 3888 3780 4052
rect 40 3832 92 3888
rect 148 3853 3672 3888
rect 148 3832 1327 3853
rect 40 3797 1327 3832
rect 1383 3797 1647 3853
rect 1703 3797 1957 3853
rect 2013 3797 2277 3853
rect 2333 3832 3672 3853
rect 3728 3832 3780 3888
rect 2333 3797 3780 3832
rect 40 3780 3780 3797
rect 670 3583 3320 3600
rect 670 3563 1487 3583
rect 670 3507 707 3563
rect 763 3527 1487 3563
rect 1543 3527 1797 3583
rect 1853 3527 2117 3583
rect 2173 3527 2437 3583
rect 2493 3563 3320 3583
rect 2493 3527 3227 3563
rect 763 3507 3227 3527
rect 3283 3507 3320 3563
rect 670 3313 3320 3507
rect 670 3257 707 3313
rect 763 3293 3227 3313
rect 763 3257 1487 3293
rect 670 3237 1487 3257
rect 1543 3237 1797 3293
rect 1853 3237 2117 3293
rect 2173 3237 2437 3293
rect 2493 3257 3227 3293
rect 3283 3257 3320 3313
rect 2493 3237 3320 3257
rect 670 3220 3320 3237
rect 1770 3042 2050 3065
rect 1770 2818 1798 3042
rect 2022 2818 2050 3042
rect 1770 2795 2050 2818
rect -1150 2623 4990 2640
rect -1150 2613 337 2623
rect -1150 2557 -1113 2613
rect -1057 2567 337 2613
rect 393 2567 857 2623
rect 913 2567 1367 2623
rect 1423 2567 1887 2623
rect 1943 2567 2397 2623
rect 2453 2567 2917 2623
rect 2973 2567 3437 2623
rect 3493 2613 4990 2623
rect 3493 2567 4897 2613
rect -1057 2557 4897 2567
rect 4953 2557 4990 2613
rect -1150 2453 4990 2557
rect -1150 2397 -1113 2453
rect -1057 2443 4897 2453
rect -1057 2397 337 2443
rect -1150 2387 337 2397
rect 393 2387 857 2443
rect 913 2387 1367 2443
rect 1423 2387 1887 2443
rect 1943 2387 2397 2443
rect 2453 2387 2917 2443
rect 2973 2387 3437 2443
rect 3493 2397 4897 2443
rect 4953 2397 4990 2453
rect 3493 2387 4990 2397
rect -1150 2370 4990 2387
rect 330 1953 3500 1970
rect 330 1897 597 1953
rect 653 1947 1107 1953
rect 653 1897 773 1947
rect 330 1773 773 1897
rect 330 1717 597 1773
rect 653 1723 773 1773
rect 997 1897 1107 1947
rect 1163 1897 1627 1953
rect 1683 1897 2147 1953
rect 2203 1897 2657 1953
rect 2713 1947 3177 1953
rect 2713 1897 2833 1947
rect 997 1773 2833 1897
rect 997 1723 1107 1773
rect 653 1717 1107 1723
rect 1163 1717 1627 1773
rect 1683 1717 2147 1773
rect 2203 1717 2657 1773
rect 2713 1723 2833 1773
rect 3057 1897 3177 1947
rect 3233 1897 3500 1953
rect 3057 1773 3500 1897
rect 3057 1723 3177 1773
rect 2713 1717 3177 1723
rect 3233 1717 3500 1773
rect 330 1700 3500 1717
rect 1780 1527 2050 1545
rect 1780 1303 1803 1527
rect 2027 1303 2050 1527
rect 1780 1285 2050 1303
rect 70 1115 3750 1120
rect 60 1103 3760 1115
rect 60 1047 77 1103
rect 133 1047 597 1103
rect 653 1047 1107 1103
rect 1163 1047 1627 1103
rect 1683 1047 2137 1103
rect 2193 1047 2657 1103
rect 2713 1047 3177 1103
rect 3233 1047 3687 1103
rect 3743 1047 3760 1103
rect 60 1035 3760 1047
rect 70 935 3750 1035
rect 60 923 3760 935
rect 60 867 77 923
rect 133 867 597 923
rect 653 867 1107 923
rect 1163 867 1627 923
rect 1683 867 2137 923
rect 2193 867 2657 923
rect 2713 867 3177 923
rect 3233 867 3687 923
rect 3743 867 3760 923
rect 60 855 3760 867
rect 70 850 3750 855
rect 70 433 3750 450
rect 70 377 337 433
rect 393 427 847 433
rect 393 377 513 427
rect 70 253 513 377
rect 70 197 337 253
rect 393 203 513 253
rect 737 377 847 427
rect 903 377 1367 433
rect 1423 377 1887 433
rect 1943 377 2397 433
rect 2453 377 2917 433
rect 2973 427 3427 433
rect 2973 377 3093 427
rect 737 253 3093 377
rect 737 203 847 253
rect 393 197 847 203
rect 903 197 1367 253
rect 1423 197 1887 253
rect 1943 197 2397 253
rect 2453 197 2917 253
rect 2973 203 3093 253
rect 3317 377 3427 427
rect 3483 377 3750 433
rect 3317 253 3750 377
rect 3317 203 3427 253
rect 2973 197 3427 203
rect 3483 197 3750 253
rect 70 180 3750 197
rect 1780 -3 2050 15
rect 1780 -227 1803 -3
rect 2027 -227 2050 -3
rect 1780 -245 2050 -227
<< via3 >>
rect 1293 10903 1517 10907
rect 1293 10687 1297 10903
rect 1297 10687 1513 10903
rect 1513 10687 1517 10903
rect 1293 10683 1517 10687
rect 2343 10903 2567 10907
rect 2343 10687 2347 10903
rect 2347 10687 2563 10903
rect 2563 10687 2567 10903
rect 2343 10683 2567 10687
rect -5807 10203 -5743 10207
rect -5807 10147 -5803 10203
rect -5803 10147 -5747 10203
rect -5747 10147 -5743 10203
rect -5807 10143 -5743 10147
rect -887 10193 -663 10417
rect 1013 10183 1237 10407
rect 2593 10183 2817 10407
rect 4493 10183 4717 10407
rect 9583 10203 9647 10207
rect 9583 10147 9587 10203
rect 9587 10147 9643 10203
rect 9643 10147 9647 10203
rect 9583 10143 9647 10147
rect -5917 10093 -5853 10097
rect -5917 10037 -5913 10093
rect -5913 10037 -5857 10093
rect -5857 10037 -5853 10093
rect -5917 10033 -5853 10037
rect 9693 10093 9757 10097
rect 9693 10037 9697 10093
rect 9697 10037 9753 10093
rect 9753 10037 9757 10093
rect 9693 10033 9757 10037
rect -2017 9168 -1953 9232
rect -1827 9168 -1763 9232
rect 1293 9263 1517 9267
rect 1293 9047 1297 9263
rect 1297 9047 1513 9263
rect 1513 9047 1517 9263
rect 1293 9043 1517 9047
rect 2343 9263 2567 9267
rect 2343 9047 2347 9263
rect 2347 9047 2563 9263
rect 2563 9047 2567 9263
rect 2343 9043 2567 9047
rect 5593 9168 5657 9232
rect 5783 9168 5847 9232
rect -4022 8728 -3958 8732
rect -4022 8672 -4018 8728
rect -4018 8672 -3962 8728
rect -3962 8672 -3958 8728
rect -4022 8668 -3958 8672
rect -3942 8728 -3878 8732
rect -3942 8672 -3938 8728
rect -3938 8672 -3882 8728
rect -3882 8672 -3878 8728
rect -3942 8668 -3878 8672
rect -3602 8728 -3538 8732
rect -3602 8672 -3598 8728
rect -3598 8672 -3542 8728
rect -3542 8672 -3538 8728
rect -3602 8668 -3538 8672
rect -3522 8728 -3458 8732
rect -3522 8672 -3518 8728
rect -3518 8672 -3462 8728
rect -3462 8672 -3458 8728
rect -3522 8668 -3458 8672
rect 618 8528 842 8752
rect 1888 8528 2112 8752
rect 3148 8528 3372 8752
rect 7228 8728 7292 8732
rect 7228 8672 7232 8728
rect 7232 8672 7288 8728
rect 7288 8672 7292 8728
rect 7228 8668 7292 8672
rect 7308 8728 7372 8732
rect 7308 8672 7312 8728
rect 7312 8672 7368 8728
rect 7368 8672 7372 8728
rect 7308 8668 7372 8672
rect 7648 8728 7712 8732
rect 7648 8672 7652 8728
rect 7652 8672 7708 8728
rect 7708 8672 7712 8728
rect 7648 8668 7712 8672
rect 7728 8728 7792 8732
rect 7728 8672 7732 8728
rect 7732 8672 7788 8728
rect 7788 8672 7792 8728
rect 7728 8668 7792 8672
rect 1058 7658 1282 7662
rect 1058 7442 1062 7658
rect 1062 7442 1278 7658
rect 1278 7442 1282 7658
rect 1058 7438 1282 7442
rect 2558 7658 2782 7662
rect 2558 7442 2562 7658
rect 2562 7442 2778 7658
rect 2778 7442 2782 7658
rect 2558 7438 2782 7442
rect 618 6978 842 7202
rect 1888 6978 2112 7202
rect 3148 6978 3372 7202
rect 1798 4558 2022 4562
rect 1798 4342 1802 4558
rect 1802 4342 2018 4558
rect 2018 4342 2022 4558
rect 1798 4338 2022 4342
rect 1798 3038 2022 3042
rect 1798 2822 1802 3038
rect 1802 2822 2018 3038
rect 2018 2822 2022 3038
rect 1798 2818 2022 2822
rect 773 1723 997 1947
rect 2833 1723 3057 1947
rect 1803 1523 2027 1527
rect 1803 1307 1807 1523
rect 1807 1307 2023 1523
rect 2023 1307 2027 1523
rect 1803 1303 2027 1307
rect 513 203 737 427
rect 3093 203 3317 427
rect 1803 -7 2027 -3
rect 1803 -223 1807 -7
rect 1807 -223 2023 -7
rect 2023 -223 2027 -7
rect 1803 -227 2027 -223
<< metal4 >>
rect -5940 16310 9780 16550
rect -5940 10207 -5720 16310
rect -2350 14480 9150 14840
rect -5940 10143 -5807 10207
rect -5743 10143 -5720 10207
rect -5940 10097 -5720 10143
rect -5940 10033 -5917 10097
rect -5853 10033 -5720 10097
rect -5940 10010 -5720 10033
rect -2050 9232 -1730 14480
rect 1269 10913 1541 10931
rect 1269 10677 1287 10913
rect 1523 10677 1541 10913
rect 1269 10659 1541 10677
rect 2319 10913 2591 10931
rect 2319 10677 2337 10913
rect 2573 10677 2591 10913
rect 2319 10659 2591 10677
rect -901 10423 -649 10431
rect -901 10187 -893 10423
rect -657 10187 -649 10423
rect -901 10179 -649 10187
rect 999 10413 1251 10421
rect 999 10177 1007 10413
rect 1243 10177 1251 10413
rect 999 10169 1251 10177
rect 2579 10413 2831 10421
rect 2579 10177 2587 10413
rect 2823 10177 2831 10413
rect 2579 10169 2831 10177
rect 4479 10413 4731 10421
rect 4479 10177 4487 10413
rect 4723 10177 4731 10413
rect 4479 10169 4731 10177
rect -2050 9168 -2017 9232
rect -1953 9168 -1827 9232
rect -1763 9168 -1730 9232
rect -2050 9130 -1730 9168
rect 1269 9273 1541 9291
rect 1269 9037 1287 9273
rect 1523 9037 1541 9273
rect 1269 9019 1541 9037
rect 2319 9273 2591 9291
rect 2319 9037 2337 9273
rect 2573 9037 2591 9273
rect 5560 9232 5880 14480
rect 9560 10207 9780 16310
rect 9560 10143 9583 10207
rect 9647 10143 9780 10207
rect 9560 10097 9780 10143
rect 9560 10033 9693 10097
rect 9757 10033 9780 10097
rect 9560 10010 9780 10033
rect 5560 9168 5593 9232
rect 5657 9168 5783 9232
rect 5847 9168 5880 9232
rect 5560 9130 5880 9168
rect 2319 9019 2591 9037
rect -4070 8732 -3410 8780
rect -4070 8668 -4022 8732
rect -3958 8668 -3942 8732
rect -3878 8668 -3602 8732
rect -3538 8668 -3522 8732
rect -3458 8668 -3410 8732
rect -4070 1308 -3410 8668
rect 599 8758 861 8771
rect 599 8522 612 8758
rect 848 8522 861 8758
rect 599 8509 861 8522
rect 1869 8758 2131 8771
rect 1869 8522 1882 8758
rect 2118 8522 2131 8758
rect 1869 8509 2131 8522
rect 3129 8758 3391 8771
rect 3129 8522 3142 8758
rect 3378 8522 3391 8758
rect 3129 8509 3391 8522
rect 7180 8732 7840 8780
rect 7180 8668 7228 8732
rect 7292 8668 7308 8732
rect 7372 8668 7648 8732
rect 7712 8668 7728 8732
rect 7792 8668 7840 8732
rect 1039 7668 1301 7681
rect 1039 7432 1052 7668
rect 1288 7432 1301 7668
rect 1039 7419 1301 7432
rect 2539 7668 2801 7681
rect 2539 7432 2552 7668
rect 2788 7432 2801 7668
rect 2539 7419 2801 7432
rect 599 7208 861 7221
rect 599 6972 612 7208
rect 848 6972 861 7208
rect 599 6959 861 6972
rect 1869 7208 2131 7221
rect 1869 6972 1882 7208
rect 2118 6972 2131 7208
rect 1869 6959 2131 6972
rect 3129 7208 3391 7221
rect 3129 6972 3142 7208
rect 3378 6972 3391 7208
rect 3129 6959 3391 6972
rect 1779 4568 2041 4581
rect 1779 4332 1792 4568
rect 2028 4332 2041 4568
rect 1779 4319 2041 4332
rect 1779 3048 2041 3061
rect 1779 2812 1792 3048
rect 2028 2812 2041 3048
rect 1779 2799 2041 2812
rect 759 1953 1011 1961
rect 759 1717 767 1953
rect 1003 1717 1011 1953
rect 759 1709 1011 1717
rect 2819 1953 3071 1961
rect 2819 1717 2827 1953
rect 3063 1717 3071 1953
rect 2819 1709 3071 1717
rect -4070 1072 -4038 1308
rect -3802 1072 -3678 1308
rect -3442 1072 -3410 1308
rect 1789 1533 2041 1541
rect 1789 1297 1797 1533
rect 2033 1297 2041 1533
rect 1789 1289 2041 1297
rect 7180 1308 7840 8668
rect -4070 968 -3410 1072
rect -4070 732 -4038 968
rect -3802 732 -3678 968
rect -3442 732 -3410 968
rect -4070 700 -3410 732
rect 7180 1072 7212 1308
rect 7448 1072 7572 1308
rect 7808 1072 7840 1308
rect 7180 968 7840 1072
rect 7180 732 7212 968
rect 7448 732 7572 968
rect 7808 732 7840 968
rect 7180 700 7840 732
rect 499 433 751 441
rect 499 197 507 433
rect 743 197 751 433
rect 499 189 751 197
rect 3079 433 3331 441
rect 3079 197 3087 433
rect 3323 197 3331 433
rect 3079 189 3331 197
rect 1789 3 2041 11
rect 1789 -233 1797 3
rect 2033 -233 2041 3
rect 1789 -241 2041 -233
<< via4 >>
rect 1287 10907 1523 10913
rect 1287 10683 1293 10907
rect 1293 10683 1517 10907
rect 1517 10683 1523 10907
rect 1287 10677 1523 10683
rect 2337 10907 2573 10913
rect 2337 10683 2343 10907
rect 2343 10683 2567 10907
rect 2567 10683 2573 10907
rect 2337 10677 2573 10683
rect -893 10417 -657 10423
rect -893 10193 -887 10417
rect -887 10193 -663 10417
rect -663 10193 -657 10417
rect -893 10187 -657 10193
rect 1007 10407 1243 10413
rect 1007 10183 1013 10407
rect 1013 10183 1237 10407
rect 1237 10183 1243 10407
rect 1007 10177 1243 10183
rect 2587 10407 2823 10413
rect 2587 10183 2593 10407
rect 2593 10183 2817 10407
rect 2817 10183 2823 10407
rect 2587 10177 2823 10183
rect 4487 10407 4723 10413
rect 4487 10183 4493 10407
rect 4493 10183 4717 10407
rect 4717 10183 4723 10407
rect 4487 10177 4723 10183
rect 1287 9267 1523 9273
rect 1287 9043 1293 9267
rect 1293 9043 1517 9267
rect 1517 9043 1523 9267
rect 1287 9037 1523 9043
rect 2337 9267 2573 9273
rect 2337 9043 2343 9267
rect 2343 9043 2567 9267
rect 2567 9043 2573 9267
rect 2337 9037 2573 9043
rect 612 8752 848 8758
rect 612 8528 618 8752
rect 618 8528 842 8752
rect 842 8528 848 8752
rect 612 8522 848 8528
rect 1882 8752 2118 8758
rect 1882 8528 1888 8752
rect 1888 8528 2112 8752
rect 2112 8528 2118 8752
rect 1882 8522 2118 8528
rect 3142 8752 3378 8758
rect 3142 8528 3148 8752
rect 3148 8528 3372 8752
rect 3372 8528 3378 8752
rect 3142 8522 3378 8528
rect 1052 7662 1288 7668
rect 1052 7438 1058 7662
rect 1058 7438 1282 7662
rect 1282 7438 1288 7662
rect 1052 7432 1288 7438
rect 2552 7662 2788 7668
rect 2552 7438 2558 7662
rect 2558 7438 2782 7662
rect 2782 7438 2788 7662
rect 2552 7432 2788 7438
rect 612 7202 848 7208
rect 612 6978 618 7202
rect 618 6978 842 7202
rect 842 6978 848 7202
rect 612 6972 848 6978
rect 1882 7202 2118 7208
rect 1882 6978 1888 7202
rect 1888 6978 2112 7202
rect 2112 6978 2118 7202
rect 1882 6972 2118 6978
rect 3142 7202 3378 7208
rect 3142 6978 3148 7202
rect 3148 6978 3372 7202
rect 3372 6978 3378 7202
rect 3142 6972 3378 6978
rect 1792 4562 2028 4568
rect 1792 4338 1798 4562
rect 1798 4338 2022 4562
rect 2022 4338 2028 4562
rect 1792 4332 2028 4338
rect 1792 3042 2028 3048
rect 1792 2818 1798 3042
rect 1798 2818 2022 3042
rect 2022 2818 2028 3042
rect 1792 2812 2028 2818
rect 767 1947 1003 1953
rect 767 1723 773 1947
rect 773 1723 997 1947
rect 997 1723 1003 1947
rect 767 1717 1003 1723
rect 2827 1947 3063 1953
rect 2827 1723 2833 1947
rect 2833 1723 3057 1947
rect 3057 1723 3063 1947
rect 2827 1717 3063 1723
rect -4038 1072 -3802 1308
rect -3678 1072 -3442 1308
rect 1797 1527 2033 1533
rect 1797 1303 1803 1527
rect 1803 1303 2027 1527
rect 2027 1303 2033 1527
rect 1797 1297 2033 1303
rect -4038 732 -3802 968
rect -3678 732 -3442 968
rect 7212 1072 7448 1308
rect 7572 1072 7808 1308
rect 7212 732 7448 968
rect 7572 732 7808 968
rect 507 427 743 433
rect 507 203 513 427
rect 513 203 737 427
rect 737 203 743 427
rect 507 197 743 203
rect 3087 427 3323 433
rect 3087 203 3093 427
rect 3093 203 3317 427
rect 3317 203 3323 427
rect 3087 197 3323 203
rect 1797 -3 2033 3
rect 1797 -227 1803 -3
rect 1803 -227 2027 -3
rect 2027 -227 2033 -3
rect 1797 -233 2033 -227
<< metal5 >>
rect 1240 10913 2620 10980
rect 1240 10677 1287 10913
rect 1523 10677 2337 10913
rect 2573 10677 2620 10913
rect 1240 10460 2620 10677
rect -930 10423 4770 10460
rect -930 10187 -893 10423
rect -657 10413 4770 10423
rect -657 10187 1007 10413
rect -930 10177 1007 10187
rect 1243 10177 2587 10413
rect 2823 10177 4487 10413
rect 4723 10177 4770 10413
rect -930 10130 4770 10177
rect 1240 9273 2620 10130
rect 1240 9037 1287 9273
rect 1523 9037 2337 9273
rect 2573 9037 2620 9273
rect 1240 8800 2620 9037
rect 450 8758 3430 8800
rect 450 8522 612 8758
rect 848 8522 1882 8758
rect 2118 8522 3142 8758
rect 3378 8522 3430 8758
rect 450 8480 3430 8522
rect 1240 7710 2620 8480
rect 1010 7668 2830 7710
rect 1010 7432 1052 7668
rect 1288 7432 2552 7668
rect 2788 7432 2830 7668
rect 1010 7250 2830 7432
rect 560 7208 3430 7250
rect 560 6972 612 7208
rect 848 6972 1882 7208
rect 2118 6972 3142 7208
rect 3378 6972 3430 7208
rect 560 6930 3430 6972
rect 1690 4568 2130 4620
rect 1690 4332 1792 4568
rect 2028 4332 2130 4568
rect 1690 3048 2130 4332
rect 1690 2812 1792 3048
rect 2028 2812 2130 3048
rect 1690 2000 2130 2812
rect -920 1953 4720 2000
rect -920 1717 767 1953
rect 1003 1717 2827 1953
rect 3063 1717 4720 1953
rect -920 1533 4720 1717
rect -920 1340 1797 1533
rect -4070 1308 1797 1340
rect -4070 1072 -4038 1308
rect -3802 1072 -3678 1308
rect -3442 1297 1797 1308
rect 2033 1340 4720 1533
rect 2033 1308 7840 1340
rect 2033 1297 7212 1308
rect -3442 1072 7212 1297
rect 7448 1072 7572 1308
rect 7808 1072 7840 1308
rect -4070 968 7840 1072
rect -4070 732 -4038 968
rect -3802 732 -3678 968
rect -3442 732 7212 968
rect 7448 732 7572 968
rect 7808 732 7840 968
rect -4070 700 7840 732
rect -920 433 4720 700
rect -920 197 507 433
rect 743 197 3087 433
rect 3323 197 4720 433
rect -920 150 4720 197
rect 1700 3 2140 150
rect 1700 -233 1797 3
rect 2033 -233 2140 3
rect 1700 -310 2140 -233
use sky130_fd_pr__cap_mim_m3_1_95KK7Z  sky130_fd_pr__cap_mim_m3_1_95KK7Z_0
timestamp 1710000196
transform 0 -1 7610 1 0 14670
box -1750 -1700 1749 1700
use sky130_fd_pr__cap_mim_m3_1_95KK7Z  sky130_fd_pr__cap_mim_m3_1_95KK7Z_1
timestamp 1710000196
transform 0 -1 3810 1 0 14670
box -1750 -1700 1749 1700
use sky130_fd_pr__cap_mim_m3_1_95KK7Z  sky130_fd_pr__cap_mim_m3_1_95KK7Z_2
timestamp 1710000196
transform 0 -1 10 1 0 14670
box -1750 -1700 1749 1700
use sky130_fd_pr__cap_mim_m3_1_95KK7Z  sky130_fd_pr__cap_mim_m3_1_95KK7Z_3
timestamp 1710000196
transform 0 -1 -3790 1 0 14670
box -1750 -1700 1749 1700
use sky130_fd_pr__nfet_01v8_EJ3ASN  sky130_fd_pr__nfet_01v8_EJ3ASN_0
timestamp 1710000196
transform 1 0 1911 0 1 5211
box -710 -700 710 700
use sky130_fd_pr__nfet_01v8_EJ3ASN  sky130_fd_pr__nfet_01v8_EJ3ASN_1
timestamp 1710000196
transform 1 0 1911 0 1 3691
box -710 -700 710 700
use sky130_fd_pr__nfet_01v8_JEXVB9  sky130_fd_pr__nfet_01v8_JEXVB9_0
timestamp 1710000196
transform 1 0 1915 0 1 2170
box -1705 -700 1705 700
use sky130_fd_pr__nfet_01v8_JT3SH9  sky130_fd_pr__nfet_01v8_JT3SH9_0
timestamp 1710000196
transform 1 0 1913 0 1 650
box -1963 -700 1963 700
use sky130_fd_pr__pfet_01v8_9F67JW  sky130_fd_pr__pfet_01v8_9F67JW_0
timestamp 1710000196
transform 1 0 1917 0 1 9989
box -3327 -719 3327 719
use sky130_fd_pr__pfet_01v8_49C6SK  sky130_fd_pr__pfet_01v8_49C6SK_0
timestamp 1710000196
transform 1 0 1916 0 1 8319
box -1826 -719 1826 719
use sky130_fd_pr__pfet_01v8_GNAJ57  sky130_fd_pr__pfet_01v8_GNAJ57_0
timestamp 1710000196
transform 1 0 1916 0 1 6779
box -1826 -719 1826 719
use sky130_fd_pr__res_xhigh_po_5p73_F7BMVG  sky130_fd_pr__res_xhigh_po_5p73_F7BMVG_0
timestamp 1710000196
transform 0 1 -3615 -1 0 10846
box -729 -1588 729 1588
use sky130_fd_pr__res_xhigh_po_5p73_F7BMVG  sky130_fd_pr__res_xhigh_po_5p73_F7BMVG_1
timestamp 1710000196
transform 0 1 -3615 -1 0 9386
box -729 -1588 729 1588
use sky130_fd_pr__res_xhigh_po_5p73_F7BMVG  sky130_fd_pr__res_xhigh_po_5p73_F7BMVG_2
timestamp 1710000196
transform 0 1 7455 -1 0 9386
box -729 -1588 729 1588
use sky130_fd_pr__res_xhigh_po_5p73_F7BMVG  sky130_fd_pr__res_xhigh_po_5p73_F7BMVG_3
timestamp 1710000196
transform 0 1 7455 -1 0 10846
box -729 -1588 729 1588
<< end >>
