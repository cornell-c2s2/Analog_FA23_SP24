** sch_path: /foss/designs/Analog_FA23_SP24/flashADC/xschem/frontAnalog_v0p0p1.sch
.lib /foss/pdks/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.include /foss/pdks/sky130A/libs.ref/sky130_fd_sc_hd/spice/sky130_fd_sc_hd.spice

.subckt frontAnalog_v0p0p1 VDD GND VN VIN IB CLK Q
*.PININFO VDD:I GND:I VN:I VIN:I IB:I CLK:I Q:O
x63 net1 GND GND VDD VDD net4 sky130_fd_sc_hd__buf_1
x65 net2 GND GND VDD VDD net5 sky130_fd_sc_hd__buf_1
* noconn #net6
x1 VDD net4 net5 Q net6 GND RSfetsym
x2 net3 net1 net2 VN VIN IB CLK GND class_AB_v4_sym
.ends



.GLOBAL GND
.GLOBAL VDD
.end
