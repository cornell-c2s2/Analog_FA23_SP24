magic
tech sky130A
magscale 1 2
timestamp 1710000196
<< nwell >>
rect -1826 -719 1826 719
<< pmos >>
rect -1630 -500 -1530 500
rect -1472 -500 -1372 500
rect -1314 -500 -1214 500
rect -1156 -500 -1056 500
rect -998 -500 -898 500
rect -840 -500 -740 500
rect -682 -500 -582 500
rect -524 -500 -424 500
rect -366 -500 -266 500
rect -208 -500 -108 500
rect -50 -500 50 500
rect 108 -500 208 500
rect 266 -500 366 500
rect 424 -500 524 500
rect 582 -500 682 500
rect 740 -500 840 500
rect 898 -500 998 500
rect 1056 -500 1156 500
rect 1214 -500 1314 500
rect 1372 -500 1472 500
rect 1530 -500 1630 500
<< pdiff >>
rect -1688 459 -1630 500
rect -1688 425 -1676 459
rect -1642 425 -1630 459
rect -1688 391 -1630 425
rect -1688 357 -1676 391
rect -1642 357 -1630 391
rect -1688 323 -1630 357
rect -1688 289 -1676 323
rect -1642 289 -1630 323
rect -1688 255 -1630 289
rect -1688 221 -1676 255
rect -1642 221 -1630 255
rect -1688 187 -1630 221
rect -1688 153 -1676 187
rect -1642 153 -1630 187
rect -1688 119 -1630 153
rect -1688 85 -1676 119
rect -1642 85 -1630 119
rect -1688 51 -1630 85
rect -1688 17 -1676 51
rect -1642 17 -1630 51
rect -1688 -17 -1630 17
rect -1688 -51 -1676 -17
rect -1642 -51 -1630 -17
rect -1688 -85 -1630 -51
rect -1688 -119 -1676 -85
rect -1642 -119 -1630 -85
rect -1688 -153 -1630 -119
rect -1688 -187 -1676 -153
rect -1642 -187 -1630 -153
rect -1688 -221 -1630 -187
rect -1688 -255 -1676 -221
rect -1642 -255 -1630 -221
rect -1688 -289 -1630 -255
rect -1688 -323 -1676 -289
rect -1642 -323 -1630 -289
rect -1688 -357 -1630 -323
rect -1688 -391 -1676 -357
rect -1642 -391 -1630 -357
rect -1688 -425 -1630 -391
rect -1688 -459 -1676 -425
rect -1642 -459 -1630 -425
rect -1688 -500 -1630 -459
rect -1530 459 -1472 500
rect -1530 425 -1518 459
rect -1484 425 -1472 459
rect -1530 391 -1472 425
rect -1530 357 -1518 391
rect -1484 357 -1472 391
rect -1530 323 -1472 357
rect -1530 289 -1518 323
rect -1484 289 -1472 323
rect -1530 255 -1472 289
rect -1530 221 -1518 255
rect -1484 221 -1472 255
rect -1530 187 -1472 221
rect -1530 153 -1518 187
rect -1484 153 -1472 187
rect -1530 119 -1472 153
rect -1530 85 -1518 119
rect -1484 85 -1472 119
rect -1530 51 -1472 85
rect -1530 17 -1518 51
rect -1484 17 -1472 51
rect -1530 -17 -1472 17
rect -1530 -51 -1518 -17
rect -1484 -51 -1472 -17
rect -1530 -85 -1472 -51
rect -1530 -119 -1518 -85
rect -1484 -119 -1472 -85
rect -1530 -153 -1472 -119
rect -1530 -187 -1518 -153
rect -1484 -187 -1472 -153
rect -1530 -221 -1472 -187
rect -1530 -255 -1518 -221
rect -1484 -255 -1472 -221
rect -1530 -289 -1472 -255
rect -1530 -323 -1518 -289
rect -1484 -323 -1472 -289
rect -1530 -357 -1472 -323
rect -1530 -391 -1518 -357
rect -1484 -391 -1472 -357
rect -1530 -425 -1472 -391
rect -1530 -459 -1518 -425
rect -1484 -459 -1472 -425
rect -1530 -500 -1472 -459
rect -1372 459 -1314 500
rect -1372 425 -1360 459
rect -1326 425 -1314 459
rect -1372 391 -1314 425
rect -1372 357 -1360 391
rect -1326 357 -1314 391
rect -1372 323 -1314 357
rect -1372 289 -1360 323
rect -1326 289 -1314 323
rect -1372 255 -1314 289
rect -1372 221 -1360 255
rect -1326 221 -1314 255
rect -1372 187 -1314 221
rect -1372 153 -1360 187
rect -1326 153 -1314 187
rect -1372 119 -1314 153
rect -1372 85 -1360 119
rect -1326 85 -1314 119
rect -1372 51 -1314 85
rect -1372 17 -1360 51
rect -1326 17 -1314 51
rect -1372 -17 -1314 17
rect -1372 -51 -1360 -17
rect -1326 -51 -1314 -17
rect -1372 -85 -1314 -51
rect -1372 -119 -1360 -85
rect -1326 -119 -1314 -85
rect -1372 -153 -1314 -119
rect -1372 -187 -1360 -153
rect -1326 -187 -1314 -153
rect -1372 -221 -1314 -187
rect -1372 -255 -1360 -221
rect -1326 -255 -1314 -221
rect -1372 -289 -1314 -255
rect -1372 -323 -1360 -289
rect -1326 -323 -1314 -289
rect -1372 -357 -1314 -323
rect -1372 -391 -1360 -357
rect -1326 -391 -1314 -357
rect -1372 -425 -1314 -391
rect -1372 -459 -1360 -425
rect -1326 -459 -1314 -425
rect -1372 -500 -1314 -459
rect -1214 459 -1156 500
rect -1214 425 -1202 459
rect -1168 425 -1156 459
rect -1214 391 -1156 425
rect -1214 357 -1202 391
rect -1168 357 -1156 391
rect -1214 323 -1156 357
rect -1214 289 -1202 323
rect -1168 289 -1156 323
rect -1214 255 -1156 289
rect -1214 221 -1202 255
rect -1168 221 -1156 255
rect -1214 187 -1156 221
rect -1214 153 -1202 187
rect -1168 153 -1156 187
rect -1214 119 -1156 153
rect -1214 85 -1202 119
rect -1168 85 -1156 119
rect -1214 51 -1156 85
rect -1214 17 -1202 51
rect -1168 17 -1156 51
rect -1214 -17 -1156 17
rect -1214 -51 -1202 -17
rect -1168 -51 -1156 -17
rect -1214 -85 -1156 -51
rect -1214 -119 -1202 -85
rect -1168 -119 -1156 -85
rect -1214 -153 -1156 -119
rect -1214 -187 -1202 -153
rect -1168 -187 -1156 -153
rect -1214 -221 -1156 -187
rect -1214 -255 -1202 -221
rect -1168 -255 -1156 -221
rect -1214 -289 -1156 -255
rect -1214 -323 -1202 -289
rect -1168 -323 -1156 -289
rect -1214 -357 -1156 -323
rect -1214 -391 -1202 -357
rect -1168 -391 -1156 -357
rect -1214 -425 -1156 -391
rect -1214 -459 -1202 -425
rect -1168 -459 -1156 -425
rect -1214 -500 -1156 -459
rect -1056 459 -998 500
rect -1056 425 -1044 459
rect -1010 425 -998 459
rect -1056 391 -998 425
rect -1056 357 -1044 391
rect -1010 357 -998 391
rect -1056 323 -998 357
rect -1056 289 -1044 323
rect -1010 289 -998 323
rect -1056 255 -998 289
rect -1056 221 -1044 255
rect -1010 221 -998 255
rect -1056 187 -998 221
rect -1056 153 -1044 187
rect -1010 153 -998 187
rect -1056 119 -998 153
rect -1056 85 -1044 119
rect -1010 85 -998 119
rect -1056 51 -998 85
rect -1056 17 -1044 51
rect -1010 17 -998 51
rect -1056 -17 -998 17
rect -1056 -51 -1044 -17
rect -1010 -51 -998 -17
rect -1056 -85 -998 -51
rect -1056 -119 -1044 -85
rect -1010 -119 -998 -85
rect -1056 -153 -998 -119
rect -1056 -187 -1044 -153
rect -1010 -187 -998 -153
rect -1056 -221 -998 -187
rect -1056 -255 -1044 -221
rect -1010 -255 -998 -221
rect -1056 -289 -998 -255
rect -1056 -323 -1044 -289
rect -1010 -323 -998 -289
rect -1056 -357 -998 -323
rect -1056 -391 -1044 -357
rect -1010 -391 -998 -357
rect -1056 -425 -998 -391
rect -1056 -459 -1044 -425
rect -1010 -459 -998 -425
rect -1056 -500 -998 -459
rect -898 459 -840 500
rect -898 425 -886 459
rect -852 425 -840 459
rect -898 391 -840 425
rect -898 357 -886 391
rect -852 357 -840 391
rect -898 323 -840 357
rect -898 289 -886 323
rect -852 289 -840 323
rect -898 255 -840 289
rect -898 221 -886 255
rect -852 221 -840 255
rect -898 187 -840 221
rect -898 153 -886 187
rect -852 153 -840 187
rect -898 119 -840 153
rect -898 85 -886 119
rect -852 85 -840 119
rect -898 51 -840 85
rect -898 17 -886 51
rect -852 17 -840 51
rect -898 -17 -840 17
rect -898 -51 -886 -17
rect -852 -51 -840 -17
rect -898 -85 -840 -51
rect -898 -119 -886 -85
rect -852 -119 -840 -85
rect -898 -153 -840 -119
rect -898 -187 -886 -153
rect -852 -187 -840 -153
rect -898 -221 -840 -187
rect -898 -255 -886 -221
rect -852 -255 -840 -221
rect -898 -289 -840 -255
rect -898 -323 -886 -289
rect -852 -323 -840 -289
rect -898 -357 -840 -323
rect -898 -391 -886 -357
rect -852 -391 -840 -357
rect -898 -425 -840 -391
rect -898 -459 -886 -425
rect -852 -459 -840 -425
rect -898 -500 -840 -459
rect -740 459 -682 500
rect -740 425 -728 459
rect -694 425 -682 459
rect -740 391 -682 425
rect -740 357 -728 391
rect -694 357 -682 391
rect -740 323 -682 357
rect -740 289 -728 323
rect -694 289 -682 323
rect -740 255 -682 289
rect -740 221 -728 255
rect -694 221 -682 255
rect -740 187 -682 221
rect -740 153 -728 187
rect -694 153 -682 187
rect -740 119 -682 153
rect -740 85 -728 119
rect -694 85 -682 119
rect -740 51 -682 85
rect -740 17 -728 51
rect -694 17 -682 51
rect -740 -17 -682 17
rect -740 -51 -728 -17
rect -694 -51 -682 -17
rect -740 -85 -682 -51
rect -740 -119 -728 -85
rect -694 -119 -682 -85
rect -740 -153 -682 -119
rect -740 -187 -728 -153
rect -694 -187 -682 -153
rect -740 -221 -682 -187
rect -740 -255 -728 -221
rect -694 -255 -682 -221
rect -740 -289 -682 -255
rect -740 -323 -728 -289
rect -694 -323 -682 -289
rect -740 -357 -682 -323
rect -740 -391 -728 -357
rect -694 -391 -682 -357
rect -740 -425 -682 -391
rect -740 -459 -728 -425
rect -694 -459 -682 -425
rect -740 -500 -682 -459
rect -582 459 -524 500
rect -582 425 -570 459
rect -536 425 -524 459
rect -582 391 -524 425
rect -582 357 -570 391
rect -536 357 -524 391
rect -582 323 -524 357
rect -582 289 -570 323
rect -536 289 -524 323
rect -582 255 -524 289
rect -582 221 -570 255
rect -536 221 -524 255
rect -582 187 -524 221
rect -582 153 -570 187
rect -536 153 -524 187
rect -582 119 -524 153
rect -582 85 -570 119
rect -536 85 -524 119
rect -582 51 -524 85
rect -582 17 -570 51
rect -536 17 -524 51
rect -582 -17 -524 17
rect -582 -51 -570 -17
rect -536 -51 -524 -17
rect -582 -85 -524 -51
rect -582 -119 -570 -85
rect -536 -119 -524 -85
rect -582 -153 -524 -119
rect -582 -187 -570 -153
rect -536 -187 -524 -153
rect -582 -221 -524 -187
rect -582 -255 -570 -221
rect -536 -255 -524 -221
rect -582 -289 -524 -255
rect -582 -323 -570 -289
rect -536 -323 -524 -289
rect -582 -357 -524 -323
rect -582 -391 -570 -357
rect -536 -391 -524 -357
rect -582 -425 -524 -391
rect -582 -459 -570 -425
rect -536 -459 -524 -425
rect -582 -500 -524 -459
rect -424 459 -366 500
rect -424 425 -412 459
rect -378 425 -366 459
rect -424 391 -366 425
rect -424 357 -412 391
rect -378 357 -366 391
rect -424 323 -366 357
rect -424 289 -412 323
rect -378 289 -366 323
rect -424 255 -366 289
rect -424 221 -412 255
rect -378 221 -366 255
rect -424 187 -366 221
rect -424 153 -412 187
rect -378 153 -366 187
rect -424 119 -366 153
rect -424 85 -412 119
rect -378 85 -366 119
rect -424 51 -366 85
rect -424 17 -412 51
rect -378 17 -366 51
rect -424 -17 -366 17
rect -424 -51 -412 -17
rect -378 -51 -366 -17
rect -424 -85 -366 -51
rect -424 -119 -412 -85
rect -378 -119 -366 -85
rect -424 -153 -366 -119
rect -424 -187 -412 -153
rect -378 -187 -366 -153
rect -424 -221 -366 -187
rect -424 -255 -412 -221
rect -378 -255 -366 -221
rect -424 -289 -366 -255
rect -424 -323 -412 -289
rect -378 -323 -366 -289
rect -424 -357 -366 -323
rect -424 -391 -412 -357
rect -378 -391 -366 -357
rect -424 -425 -366 -391
rect -424 -459 -412 -425
rect -378 -459 -366 -425
rect -424 -500 -366 -459
rect -266 459 -208 500
rect -266 425 -254 459
rect -220 425 -208 459
rect -266 391 -208 425
rect -266 357 -254 391
rect -220 357 -208 391
rect -266 323 -208 357
rect -266 289 -254 323
rect -220 289 -208 323
rect -266 255 -208 289
rect -266 221 -254 255
rect -220 221 -208 255
rect -266 187 -208 221
rect -266 153 -254 187
rect -220 153 -208 187
rect -266 119 -208 153
rect -266 85 -254 119
rect -220 85 -208 119
rect -266 51 -208 85
rect -266 17 -254 51
rect -220 17 -208 51
rect -266 -17 -208 17
rect -266 -51 -254 -17
rect -220 -51 -208 -17
rect -266 -85 -208 -51
rect -266 -119 -254 -85
rect -220 -119 -208 -85
rect -266 -153 -208 -119
rect -266 -187 -254 -153
rect -220 -187 -208 -153
rect -266 -221 -208 -187
rect -266 -255 -254 -221
rect -220 -255 -208 -221
rect -266 -289 -208 -255
rect -266 -323 -254 -289
rect -220 -323 -208 -289
rect -266 -357 -208 -323
rect -266 -391 -254 -357
rect -220 -391 -208 -357
rect -266 -425 -208 -391
rect -266 -459 -254 -425
rect -220 -459 -208 -425
rect -266 -500 -208 -459
rect -108 459 -50 500
rect -108 425 -96 459
rect -62 425 -50 459
rect -108 391 -50 425
rect -108 357 -96 391
rect -62 357 -50 391
rect -108 323 -50 357
rect -108 289 -96 323
rect -62 289 -50 323
rect -108 255 -50 289
rect -108 221 -96 255
rect -62 221 -50 255
rect -108 187 -50 221
rect -108 153 -96 187
rect -62 153 -50 187
rect -108 119 -50 153
rect -108 85 -96 119
rect -62 85 -50 119
rect -108 51 -50 85
rect -108 17 -96 51
rect -62 17 -50 51
rect -108 -17 -50 17
rect -108 -51 -96 -17
rect -62 -51 -50 -17
rect -108 -85 -50 -51
rect -108 -119 -96 -85
rect -62 -119 -50 -85
rect -108 -153 -50 -119
rect -108 -187 -96 -153
rect -62 -187 -50 -153
rect -108 -221 -50 -187
rect -108 -255 -96 -221
rect -62 -255 -50 -221
rect -108 -289 -50 -255
rect -108 -323 -96 -289
rect -62 -323 -50 -289
rect -108 -357 -50 -323
rect -108 -391 -96 -357
rect -62 -391 -50 -357
rect -108 -425 -50 -391
rect -108 -459 -96 -425
rect -62 -459 -50 -425
rect -108 -500 -50 -459
rect 50 459 108 500
rect 50 425 62 459
rect 96 425 108 459
rect 50 391 108 425
rect 50 357 62 391
rect 96 357 108 391
rect 50 323 108 357
rect 50 289 62 323
rect 96 289 108 323
rect 50 255 108 289
rect 50 221 62 255
rect 96 221 108 255
rect 50 187 108 221
rect 50 153 62 187
rect 96 153 108 187
rect 50 119 108 153
rect 50 85 62 119
rect 96 85 108 119
rect 50 51 108 85
rect 50 17 62 51
rect 96 17 108 51
rect 50 -17 108 17
rect 50 -51 62 -17
rect 96 -51 108 -17
rect 50 -85 108 -51
rect 50 -119 62 -85
rect 96 -119 108 -85
rect 50 -153 108 -119
rect 50 -187 62 -153
rect 96 -187 108 -153
rect 50 -221 108 -187
rect 50 -255 62 -221
rect 96 -255 108 -221
rect 50 -289 108 -255
rect 50 -323 62 -289
rect 96 -323 108 -289
rect 50 -357 108 -323
rect 50 -391 62 -357
rect 96 -391 108 -357
rect 50 -425 108 -391
rect 50 -459 62 -425
rect 96 -459 108 -425
rect 50 -500 108 -459
rect 208 459 266 500
rect 208 425 220 459
rect 254 425 266 459
rect 208 391 266 425
rect 208 357 220 391
rect 254 357 266 391
rect 208 323 266 357
rect 208 289 220 323
rect 254 289 266 323
rect 208 255 266 289
rect 208 221 220 255
rect 254 221 266 255
rect 208 187 266 221
rect 208 153 220 187
rect 254 153 266 187
rect 208 119 266 153
rect 208 85 220 119
rect 254 85 266 119
rect 208 51 266 85
rect 208 17 220 51
rect 254 17 266 51
rect 208 -17 266 17
rect 208 -51 220 -17
rect 254 -51 266 -17
rect 208 -85 266 -51
rect 208 -119 220 -85
rect 254 -119 266 -85
rect 208 -153 266 -119
rect 208 -187 220 -153
rect 254 -187 266 -153
rect 208 -221 266 -187
rect 208 -255 220 -221
rect 254 -255 266 -221
rect 208 -289 266 -255
rect 208 -323 220 -289
rect 254 -323 266 -289
rect 208 -357 266 -323
rect 208 -391 220 -357
rect 254 -391 266 -357
rect 208 -425 266 -391
rect 208 -459 220 -425
rect 254 -459 266 -425
rect 208 -500 266 -459
rect 366 459 424 500
rect 366 425 378 459
rect 412 425 424 459
rect 366 391 424 425
rect 366 357 378 391
rect 412 357 424 391
rect 366 323 424 357
rect 366 289 378 323
rect 412 289 424 323
rect 366 255 424 289
rect 366 221 378 255
rect 412 221 424 255
rect 366 187 424 221
rect 366 153 378 187
rect 412 153 424 187
rect 366 119 424 153
rect 366 85 378 119
rect 412 85 424 119
rect 366 51 424 85
rect 366 17 378 51
rect 412 17 424 51
rect 366 -17 424 17
rect 366 -51 378 -17
rect 412 -51 424 -17
rect 366 -85 424 -51
rect 366 -119 378 -85
rect 412 -119 424 -85
rect 366 -153 424 -119
rect 366 -187 378 -153
rect 412 -187 424 -153
rect 366 -221 424 -187
rect 366 -255 378 -221
rect 412 -255 424 -221
rect 366 -289 424 -255
rect 366 -323 378 -289
rect 412 -323 424 -289
rect 366 -357 424 -323
rect 366 -391 378 -357
rect 412 -391 424 -357
rect 366 -425 424 -391
rect 366 -459 378 -425
rect 412 -459 424 -425
rect 366 -500 424 -459
rect 524 459 582 500
rect 524 425 536 459
rect 570 425 582 459
rect 524 391 582 425
rect 524 357 536 391
rect 570 357 582 391
rect 524 323 582 357
rect 524 289 536 323
rect 570 289 582 323
rect 524 255 582 289
rect 524 221 536 255
rect 570 221 582 255
rect 524 187 582 221
rect 524 153 536 187
rect 570 153 582 187
rect 524 119 582 153
rect 524 85 536 119
rect 570 85 582 119
rect 524 51 582 85
rect 524 17 536 51
rect 570 17 582 51
rect 524 -17 582 17
rect 524 -51 536 -17
rect 570 -51 582 -17
rect 524 -85 582 -51
rect 524 -119 536 -85
rect 570 -119 582 -85
rect 524 -153 582 -119
rect 524 -187 536 -153
rect 570 -187 582 -153
rect 524 -221 582 -187
rect 524 -255 536 -221
rect 570 -255 582 -221
rect 524 -289 582 -255
rect 524 -323 536 -289
rect 570 -323 582 -289
rect 524 -357 582 -323
rect 524 -391 536 -357
rect 570 -391 582 -357
rect 524 -425 582 -391
rect 524 -459 536 -425
rect 570 -459 582 -425
rect 524 -500 582 -459
rect 682 459 740 500
rect 682 425 694 459
rect 728 425 740 459
rect 682 391 740 425
rect 682 357 694 391
rect 728 357 740 391
rect 682 323 740 357
rect 682 289 694 323
rect 728 289 740 323
rect 682 255 740 289
rect 682 221 694 255
rect 728 221 740 255
rect 682 187 740 221
rect 682 153 694 187
rect 728 153 740 187
rect 682 119 740 153
rect 682 85 694 119
rect 728 85 740 119
rect 682 51 740 85
rect 682 17 694 51
rect 728 17 740 51
rect 682 -17 740 17
rect 682 -51 694 -17
rect 728 -51 740 -17
rect 682 -85 740 -51
rect 682 -119 694 -85
rect 728 -119 740 -85
rect 682 -153 740 -119
rect 682 -187 694 -153
rect 728 -187 740 -153
rect 682 -221 740 -187
rect 682 -255 694 -221
rect 728 -255 740 -221
rect 682 -289 740 -255
rect 682 -323 694 -289
rect 728 -323 740 -289
rect 682 -357 740 -323
rect 682 -391 694 -357
rect 728 -391 740 -357
rect 682 -425 740 -391
rect 682 -459 694 -425
rect 728 -459 740 -425
rect 682 -500 740 -459
rect 840 459 898 500
rect 840 425 852 459
rect 886 425 898 459
rect 840 391 898 425
rect 840 357 852 391
rect 886 357 898 391
rect 840 323 898 357
rect 840 289 852 323
rect 886 289 898 323
rect 840 255 898 289
rect 840 221 852 255
rect 886 221 898 255
rect 840 187 898 221
rect 840 153 852 187
rect 886 153 898 187
rect 840 119 898 153
rect 840 85 852 119
rect 886 85 898 119
rect 840 51 898 85
rect 840 17 852 51
rect 886 17 898 51
rect 840 -17 898 17
rect 840 -51 852 -17
rect 886 -51 898 -17
rect 840 -85 898 -51
rect 840 -119 852 -85
rect 886 -119 898 -85
rect 840 -153 898 -119
rect 840 -187 852 -153
rect 886 -187 898 -153
rect 840 -221 898 -187
rect 840 -255 852 -221
rect 886 -255 898 -221
rect 840 -289 898 -255
rect 840 -323 852 -289
rect 886 -323 898 -289
rect 840 -357 898 -323
rect 840 -391 852 -357
rect 886 -391 898 -357
rect 840 -425 898 -391
rect 840 -459 852 -425
rect 886 -459 898 -425
rect 840 -500 898 -459
rect 998 459 1056 500
rect 998 425 1010 459
rect 1044 425 1056 459
rect 998 391 1056 425
rect 998 357 1010 391
rect 1044 357 1056 391
rect 998 323 1056 357
rect 998 289 1010 323
rect 1044 289 1056 323
rect 998 255 1056 289
rect 998 221 1010 255
rect 1044 221 1056 255
rect 998 187 1056 221
rect 998 153 1010 187
rect 1044 153 1056 187
rect 998 119 1056 153
rect 998 85 1010 119
rect 1044 85 1056 119
rect 998 51 1056 85
rect 998 17 1010 51
rect 1044 17 1056 51
rect 998 -17 1056 17
rect 998 -51 1010 -17
rect 1044 -51 1056 -17
rect 998 -85 1056 -51
rect 998 -119 1010 -85
rect 1044 -119 1056 -85
rect 998 -153 1056 -119
rect 998 -187 1010 -153
rect 1044 -187 1056 -153
rect 998 -221 1056 -187
rect 998 -255 1010 -221
rect 1044 -255 1056 -221
rect 998 -289 1056 -255
rect 998 -323 1010 -289
rect 1044 -323 1056 -289
rect 998 -357 1056 -323
rect 998 -391 1010 -357
rect 1044 -391 1056 -357
rect 998 -425 1056 -391
rect 998 -459 1010 -425
rect 1044 -459 1056 -425
rect 998 -500 1056 -459
rect 1156 459 1214 500
rect 1156 425 1168 459
rect 1202 425 1214 459
rect 1156 391 1214 425
rect 1156 357 1168 391
rect 1202 357 1214 391
rect 1156 323 1214 357
rect 1156 289 1168 323
rect 1202 289 1214 323
rect 1156 255 1214 289
rect 1156 221 1168 255
rect 1202 221 1214 255
rect 1156 187 1214 221
rect 1156 153 1168 187
rect 1202 153 1214 187
rect 1156 119 1214 153
rect 1156 85 1168 119
rect 1202 85 1214 119
rect 1156 51 1214 85
rect 1156 17 1168 51
rect 1202 17 1214 51
rect 1156 -17 1214 17
rect 1156 -51 1168 -17
rect 1202 -51 1214 -17
rect 1156 -85 1214 -51
rect 1156 -119 1168 -85
rect 1202 -119 1214 -85
rect 1156 -153 1214 -119
rect 1156 -187 1168 -153
rect 1202 -187 1214 -153
rect 1156 -221 1214 -187
rect 1156 -255 1168 -221
rect 1202 -255 1214 -221
rect 1156 -289 1214 -255
rect 1156 -323 1168 -289
rect 1202 -323 1214 -289
rect 1156 -357 1214 -323
rect 1156 -391 1168 -357
rect 1202 -391 1214 -357
rect 1156 -425 1214 -391
rect 1156 -459 1168 -425
rect 1202 -459 1214 -425
rect 1156 -500 1214 -459
rect 1314 459 1372 500
rect 1314 425 1326 459
rect 1360 425 1372 459
rect 1314 391 1372 425
rect 1314 357 1326 391
rect 1360 357 1372 391
rect 1314 323 1372 357
rect 1314 289 1326 323
rect 1360 289 1372 323
rect 1314 255 1372 289
rect 1314 221 1326 255
rect 1360 221 1372 255
rect 1314 187 1372 221
rect 1314 153 1326 187
rect 1360 153 1372 187
rect 1314 119 1372 153
rect 1314 85 1326 119
rect 1360 85 1372 119
rect 1314 51 1372 85
rect 1314 17 1326 51
rect 1360 17 1372 51
rect 1314 -17 1372 17
rect 1314 -51 1326 -17
rect 1360 -51 1372 -17
rect 1314 -85 1372 -51
rect 1314 -119 1326 -85
rect 1360 -119 1372 -85
rect 1314 -153 1372 -119
rect 1314 -187 1326 -153
rect 1360 -187 1372 -153
rect 1314 -221 1372 -187
rect 1314 -255 1326 -221
rect 1360 -255 1372 -221
rect 1314 -289 1372 -255
rect 1314 -323 1326 -289
rect 1360 -323 1372 -289
rect 1314 -357 1372 -323
rect 1314 -391 1326 -357
rect 1360 -391 1372 -357
rect 1314 -425 1372 -391
rect 1314 -459 1326 -425
rect 1360 -459 1372 -425
rect 1314 -500 1372 -459
rect 1472 459 1530 500
rect 1472 425 1484 459
rect 1518 425 1530 459
rect 1472 391 1530 425
rect 1472 357 1484 391
rect 1518 357 1530 391
rect 1472 323 1530 357
rect 1472 289 1484 323
rect 1518 289 1530 323
rect 1472 255 1530 289
rect 1472 221 1484 255
rect 1518 221 1530 255
rect 1472 187 1530 221
rect 1472 153 1484 187
rect 1518 153 1530 187
rect 1472 119 1530 153
rect 1472 85 1484 119
rect 1518 85 1530 119
rect 1472 51 1530 85
rect 1472 17 1484 51
rect 1518 17 1530 51
rect 1472 -17 1530 17
rect 1472 -51 1484 -17
rect 1518 -51 1530 -17
rect 1472 -85 1530 -51
rect 1472 -119 1484 -85
rect 1518 -119 1530 -85
rect 1472 -153 1530 -119
rect 1472 -187 1484 -153
rect 1518 -187 1530 -153
rect 1472 -221 1530 -187
rect 1472 -255 1484 -221
rect 1518 -255 1530 -221
rect 1472 -289 1530 -255
rect 1472 -323 1484 -289
rect 1518 -323 1530 -289
rect 1472 -357 1530 -323
rect 1472 -391 1484 -357
rect 1518 -391 1530 -357
rect 1472 -425 1530 -391
rect 1472 -459 1484 -425
rect 1518 -459 1530 -425
rect 1472 -500 1530 -459
rect 1630 459 1688 500
rect 1630 425 1642 459
rect 1676 425 1688 459
rect 1630 391 1688 425
rect 1630 357 1642 391
rect 1676 357 1688 391
rect 1630 323 1688 357
rect 1630 289 1642 323
rect 1676 289 1688 323
rect 1630 255 1688 289
rect 1630 221 1642 255
rect 1676 221 1688 255
rect 1630 187 1688 221
rect 1630 153 1642 187
rect 1676 153 1688 187
rect 1630 119 1688 153
rect 1630 85 1642 119
rect 1676 85 1688 119
rect 1630 51 1688 85
rect 1630 17 1642 51
rect 1676 17 1688 51
rect 1630 -17 1688 17
rect 1630 -51 1642 -17
rect 1676 -51 1688 -17
rect 1630 -85 1688 -51
rect 1630 -119 1642 -85
rect 1676 -119 1688 -85
rect 1630 -153 1688 -119
rect 1630 -187 1642 -153
rect 1676 -187 1688 -153
rect 1630 -221 1688 -187
rect 1630 -255 1642 -221
rect 1676 -255 1688 -221
rect 1630 -289 1688 -255
rect 1630 -323 1642 -289
rect 1676 -323 1688 -289
rect 1630 -357 1688 -323
rect 1630 -391 1642 -357
rect 1676 -391 1688 -357
rect 1630 -425 1688 -391
rect 1630 -459 1642 -425
rect 1676 -459 1688 -425
rect 1630 -500 1688 -459
<< pdiffc >>
rect -1676 425 -1642 459
rect -1676 357 -1642 391
rect -1676 289 -1642 323
rect -1676 221 -1642 255
rect -1676 153 -1642 187
rect -1676 85 -1642 119
rect -1676 17 -1642 51
rect -1676 -51 -1642 -17
rect -1676 -119 -1642 -85
rect -1676 -187 -1642 -153
rect -1676 -255 -1642 -221
rect -1676 -323 -1642 -289
rect -1676 -391 -1642 -357
rect -1676 -459 -1642 -425
rect -1518 425 -1484 459
rect -1518 357 -1484 391
rect -1518 289 -1484 323
rect -1518 221 -1484 255
rect -1518 153 -1484 187
rect -1518 85 -1484 119
rect -1518 17 -1484 51
rect -1518 -51 -1484 -17
rect -1518 -119 -1484 -85
rect -1518 -187 -1484 -153
rect -1518 -255 -1484 -221
rect -1518 -323 -1484 -289
rect -1518 -391 -1484 -357
rect -1518 -459 -1484 -425
rect -1360 425 -1326 459
rect -1360 357 -1326 391
rect -1360 289 -1326 323
rect -1360 221 -1326 255
rect -1360 153 -1326 187
rect -1360 85 -1326 119
rect -1360 17 -1326 51
rect -1360 -51 -1326 -17
rect -1360 -119 -1326 -85
rect -1360 -187 -1326 -153
rect -1360 -255 -1326 -221
rect -1360 -323 -1326 -289
rect -1360 -391 -1326 -357
rect -1360 -459 -1326 -425
rect -1202 425 -1168 459
rect -1202 357 -1168 391
rect -1202 289 -1168 323
rect -1202 221 -1168 255
rect -1202 153 -1168 187
rect -1202 85 -1168 119
rect -1202 17 -1168 51
rect -1202 -51 -1168 -17
rect -1202 -119 -1168 -85
rect -1202 -187 -1168 -153
rect -1202 -255 -1168 -221
rect -1202 -323 -1168 -289
rect -1202 -391 -1168 -357
rect -1202 -459 -1168 -425
rect -1044 425 -1010 459
rect -1044 357 -1010 391
rect -1044 289 -1010 323
rect -1044 221 -1010 255
rect -1044 153 -1010 187
rect -1044 85 -1010 119
rect -1044 17 -1010 51
rect -1044 -51 -1010 -17
rect -1044 -119 -1010 -85
rect -1044 -187 -1010 -153
rect -1044 -255 -1010 -221
rect -1044 -323 -1010 -289
rect -1044 -391 -1010 -357
rect -1044 -459 -1010 -425
rect -886 425 -852 459
rect -886 357 -852 391
rect -886 289 -852 323
rect -886 221 -852 255
rect -886 153 -852 187
rect -886 85 -852 119
rect -886 17 -852 51
rect -886 -51 -852 -17
rect -886 -119 -852 -85
rect -886 -187 -852 -153
rect -886 -255 -852 -221
rect -886 -323 -852 -289
rect -886 -391 -852 -357
rect -886 -459 -852 -425
rect -728 425 -694 459
rect -728 357 -694 391
rect -728 289 -694 323
rect -728 221 -694 255
rect -728 153 -694 187
rect -728 85 -694 119
rect -728 17 -694 51
rect -728 -51 -694 -17
rect -728 -119 -694 -85
rect -728 -187 -694 -153
rect -728 -255 -694 -221
rect -728 -323 -694 -289
rect -728 -391 -694 -357
rect -728 -459 -694 -425
rect -570 425 -536 459
rect -570 357 -536 391
rect -570 289 -536 323
rect -570 221 -536 255
rect -570 153 -536 187
rect -570 85 -536 119
rect -570 17 -536 51
rect -570 -51 -536 -17
rect -570 -119 -536 -85
rect -570 -187 -536 -153
rect -570 -255 -536 -221
rect -570 -323 -536 -289
rect -570 -391 -536 -357
rect -570 -459 -536 -425
rect -412 425 -378 459
rect -412 357 -378 391
rect -412 289 -378 323
rect -412 221 -378 255
rect -412 153 -378 187
rect -412 85 -378 119
rect -412 17 -378 51
rect -412 -51 -378 -17
rect -412 -119 -378 -85
rect -412 -187 -378 -153
rect -412 -255 -378 -221
rect -412 -323 -378 -289
rect -412 -391 -378 -357
rect -412 -459 -378 -425
rect -254 425 -220 459
rect -254 357 -220 391
rect -254 289 -220 323
rect -254 221 -220 255
rect -254 153 -220 187
rect -254 85 -220 119
rect -254 17 -220 51
rect -254 -51 -220 -17
rect -254 -119 -220 -85
rect -254 -187 -220 -153
rect -254 -255 -220 -221
rect -254 -323 -220 -289
rect -254 -391 -220 -357
rect -254 -459 -220 -425
rect -96 425 -62 459
rect -96 357 -62 391
rect -96 289 -62 323
rect -96 221 -62 255
rect -96 153 -62 187
rect -96 85 -62 119
rect -96 17 -62 51
rect -96 -51 -62 -17
rect -96 -119 -62 -85
rect -96 -187 -62 -153
rect -96 -255 -62 -221
rect -96 -323 -62 -289
rect -96 -391 -62 -357
rect -96 -459 -62 -425
rect 62 425 96 459
rect 62 357 96 391
rect 62 289 96 323
rect 62 221 96 255
rect 62 153 96 187
rect 62 85 96 119
rect 62 17 96 51
rect 62 -51 96 -17
rect 62 -119 96 -85
rect 62 -187 96 -153
rect 62 -255 96 -221
rect 62 -323 96 -289
rect 62 -391 96 -357
rect 62 -459 96 -425
rect 220 425 254 459
rect 220 357 254 391
rect 220 289 254 323
rect 220 221 254 255
rect 220 153 254 187
rect 220 85 254 119
rect 220 17 254 51
rect 220 -51 254 -17
rect 220 -119 254 -85
rect 220 -187 254 -153
rect 220 -255 254 -221
rect 220 -323 254 -289
rect 220 -391 254 -357
rect 220 -459 254 -425
rect 378 425 412 459
rect 378 357 412 391
rect 378 289 412 323
rect 378 221 412 255
rect 378 153 412 187
rect 378 85 412 119
rect 378 17 412 51
rect 378 -51 412 -17
rect 378 -119 412 -85
rect 378 -187 412 -153
rect 378 -255 412 -221
rect 378 -323 412 -289
rect 378 -391 412 -357
rect 378 -459 412 -425
rect 536 425 570 459
rect 536 357 570 391
rect 536 289 570 323
rect 536 221 570 255
rect 536 153 570 187
rect 536 85 570 119
rect 536 17 570 51
rect 536 -51 570 -17
rect 536 -119 570 -85
rect 536 -187 570 -153
rect 536 -255 570 -221
rect 536 -323 570 -289
rect 536 -391 570 -357
rect 536 -459 570 -425
rect 694 425 728 459
rect 694 357 728 391
rect 694 289 728 323
rect 694 221 728 255
rect 694 153 728 187
rect 694 85 728 119
rect 694 17 728 51
rect 694 -51 728 -17
rect 694 -119 728 -85
rect 694 -187 728 -153
rect 694 -255 728 -221
rect 694 -323 728 -289
rect 694 -391 728 -357
rect 694 -459 728 -425
rect 852 425 886 459
rect 852 357 886 391
rect 852 289 886 323
rect 852 221 886 255
rect 852 153 886 187
rect 852 85 886 119
rect 852 17 886 51
rect 852 -51 886 -17
rect 852 -119 886 -85
rect 852 -187 886 -153
rect 852 -255 886 -221
rect 852 -323 886 -289
rect 852 -391 886 -357
rect 852 -459 886 -425
rect 1010 425 1044 459
rect 1010 357 1044 391
rect 1010 289 1044 323
rect 1010 221 1044 255
rect 1010 153 1044 187
rect 1010 85 1044 119
rect 1010 17 1044 51
rect 1010 -51 1044 -17
rect 1010 -119 1044 -85
rect 1010 -187 1044 -153
rect 1010 -255 1044 -221
rect 1010 -323 1044 -289
rect 1010 -391 1044 -357
rect 1010 -459 1044 -425
rect 1168 425 1202 459
rect 1168 357 1202 391
rect 1168 289 1202 323
rect 1168 221 1202 255
rect 1168 153 1202 187
rect 1168 85 1202 119
rect 1168 17 1202 51
rect 1168 -51 1202 -17
rect 1168 -119 1202 -85
rect 1168 -187 1202 -153
rect 1168 -255 1202 -221
rect 1168 -323 1202 -289
rect 1168 -391 1202 -357
rect 1168 -459 1202 -425
rect 1326 425 1360 459
rect 1326 357 1360 391
rect 1326 289 1360 323
rect 1326 221 1360 255
rect 1326 153 1360 187
rect 1326 85 1360 119
rect 1326 17 1360 51
rect 1326 -51 1360 -17
rect 1326 -119 1360 -85
rect 1326 -187 1360 -153
rect 1326 -255 1360 -221
rect 1326 -323 1360 -289
rect 1326 -391 1360 -357
rect 1326 -459 1360 -425
rect 1484 425 1518 459
rect 1484 357 1518 391
rect 1484 289 1518 323
rect 1484 221 1518 255
rect 1484 153 1518 187
rect 1484 85 1518 119
rect 1484 17 1518 51
rect 1484 -51 1518 -17
rect 1484 -119 1518 -85
rect 1484 -187 1518 -153
rect 1484 -255 1518 -221
rect 1484 -323 1518 -289
rect 1484 -391 1518 -357
rect 1484 -459 1518 -425
rect 1642 425 1676 459
rect 1642 357 1676 391
rect 1642 289 1676 323
rect 1642 221 1676 255
rect 1642 153 1676 187
rect 1642 85 1676 119
rect 1642 17 1676 51
rect 1642 -51 1676 -17
rect 1642 -119 1676 -85
rect 1642 -187 1676 -153
rect 1642 -255 1676 -221
rect 1642 -323 1676 -289
rect 1642 -391 1676 -357
rect 1642 -459 1676 -425
<< nsubdiff >>
rect -1790 649 -1683 683
rect -1649 649 -1615 683
rect -1581 649 -1547 683
rect -1513 649 -1479 683
rect -1445 649 -1411 683
rect -1377 649 -1343 683
rect -1309 649 -1275 683
rect -1241 649 -1207 683
rect -1173 649 -1139 683
rect -1105 649 -1071 683
rect -1037 649 -1003 683
rect -969 649 -935 683
rect -901 649 -867 683
rect -833 649 -799 683
rect -765 649 -731 683
rect -697 649 -663 683
rect -629 649 -595 683
rect -561 649 -527 683
rect -493 649 -459 683
rect -425 649 -391 683
rect -357 649 -323 683
rect -289 649 -255 683
rect -221 649 -187 683
rect -153 649 -119 683
rect -85 649 -51 683
rect -17 649 17 683
rect 51 649 85 683
rect 119 649 153 683
rect 187 649 221 683
rect 255 649 289 683
rect 323 649 357 683
rect 391 649 425 683
rect 459 649 493 683
rect 527 649 561 683
rect 595 649 629 683
rect 663 649 697 683
rect 731 649 765 683
rect 799 649 833 683
rect 867 649 901 683
rect 935 649 969 683
rect 1003 649 1037 683
rect 1071 649 1105 683
rect 1139 649 1173 683
rect 1207 649 1241 683
rect 1275 649 1309 683
rect 1343 649 1377 683
rect 1411 649 1445 683
rect 1479 649 1513 683
rect 1547 649 1581 683
rect 1615 649 1649 683
rect 1683 649 1790 683
rect -1790 561 -1756 649
rect -1790 493 -1756 527
rect 1756 561 1790 649
rect -1790 425 -1756 459
rect -1790 357 -1756 391
rect -1790 289 -1756 323
rect -1790 221 -1756 255
rect -1790 153 -1756 187
rect -1790 85 -1756 119
rect -1790 17 -1756 51
rect -1790 -51 -1756 -17
rect -1790 -119 -1756 -85
rect -1790 -187 -1756 -153
rect -1790 -255 -1756 -221
rect -1790 -323 -1756 -289
rect -1790 -391 -1756 -357
rect -1790 -459 -1756 -425
rect -1790 -527 -1756 -493
rect 1756 493 1790 527
rect 1756 425 1790 459
rect 1756 357 1790 391
rect 1756 289 1790 323
rect 1756 221 1790 255
rect 1756 153 1790 187
rect 1756 85 1790 119
rect 1756 17 1790 51
rect 1756 -51 1790 -17
rect 1756 -119 1790 -85
rect 1756 -187 1790 -153
rect 1756 -255 1790 -221
rect 1756 -323 1790 -289
rect 1756 -391 1790 -357
rect 1756 -459 1790 -425
rect -1790 -649 -1756 -561
rect 1756 -527 1790 -493
rect 1756 -649 1790 -561
rect -1790 -683 -1683 -649
rect -1649 -683 -1615 -649
rect -1581 -683 -1547 -649
rect -1513 -683 -1479 -649
rect -1445 -683 -1411 -649
rect -1377 -683 -1343 -649
rect -1309 -683 -1275 -649
rect -1241 -683 -1207 -649
rect -1173 -683 -1139 -649
rect -1105 -683 -1071 -649
rect -1037 -683 -1003 -649
rect -969 -683 -935 -649
rect -901 -683 -867 -649
rect -833 -683 -799 -649
rect -765 -683 -731 -649
rect -697 -683 -663 -649
rect -629 -683 -595 -649
rect -561 -683 -527 -649
rect -493 -683 -459 -649
rect -425 -683 -391 -649
rect -357 -683 -323 -649
rect -289 -683 -255 -649
rect -221 -683 -187 -649
rect -153 -683 -119 -649
rect -85 -683 -51 -649
rect -17 -683 17 -649
rect 51 -683 85 -649
rect 119 -683 153 -649
rect 187 -683 221 -649
rect 255 -683 289 -649
rect 323 -683 357 -649
rect 391 -683 425 -649
rect 459 -683 493 -649
rect 527 -683 561 -649
rect 595 -683 629 -649
rect 663 -683 697 -649
rect 731 -683 765 -649
rect 799 -683 833 -649
rect 867 -683 901 -649
rect 935 -683 969 -649
rect 1003 -683 1037 -649
rect 1071 -683 1105 -649
rect 1139 -683 1173 -649
rect 1207 -683 1241 -649
rect 1275 -683 1309 -649
rect 1343 -683 1377 -649
rect 1411 -683 1445 -649
rect 1479 -683 1513 -649
rect 1547 -683 1581 -649
rect 1615 -683 1649 -649
rect 1683 -683 1790 -649
<< nsubdiffcont >>
rect -1683 649 -1649 683
rect -1615 649 -1581 683
rect -1547 649 -1513 683
rect -1479 649 -1445 683
rect -1411 649 -1377 683
rect -1343 649 -1309 683
rect -1275 649 -1241 683
rect -1207 649 -1173 683
rect -1139 649 -1105 683
rect -1071 649 -1037 683
rect -1003 649 -969 683
rect -935 649 -901 683
rect -867 649 -833 683
rect -799 649 -765 683
rect -731 649 -697 683
rect -663 649 -629 683
rect -595 649 -561 683
rect -527 649 -493 683
rect -459 649 -425 683
rect -391 649 -357 683
rect -323 649 -289 683
rect -255 649 -221 683
rect -187 649 -153 683
rect -119 649 -85 683
rect -51 649 -17 683
rect 17 649 51 683
rect 85 649 119 683
rect 153 649 187 683
rect 221 649 255 683
rect 289 649 323 683
rect 357 649 391 683
rect 425 649 459 683
rect 493 649 527 683
rect 561 649 595 683
rect 629 649 663 683
rect 697 649 731 683
rect 765 649 799 683
rect 833 649 867 683
rect 901 649 935 683
rect 969 649 1003 683
rect 1037 649 1071 683
rect 1105 649 1139 683
rect 1173 649 1207 683
rect 1241 649 1275 683
rect 1309 649 1343 683
rect 1377 649 1411 683
rect 1445 649 1479 683
rect 1513 649 1547 683
rect 1581 649 1615 683
rect 1649 649 1683 683
rect -1790 527 -1756 561
rect 1756 527 1790 561
rect -1790 459 -1756 493
rect -1790 391 -1756 425
rect -1790 323 -1756 357
rect -1790 255 -1756 289
rect -1790 187 -1756 221
rect -1790 119 -1756 153
rect -1790 51 -1756 85
rect -1790 -17 -1756 17
rect -1790 -85 -1756 -51
rect -1790 -153 -1756 -119
rect -1790 -221 -1756 -187
rect -1790 -289 -1756 -255
rect -1790 -357 -1756 -323
rect -1790 -425 -1756 -391
rect -1790 -493 -1756 -459
rect 1756 459 1790 493
rect 1756 391 1790 425
rect 1756 323 1790 357
rect 1756 255 1790 289
rect 1756 187 1790 221
rect 1756 119 1790 153
rect 1756 51 1790 85
rect 1756 -17 1790 17
rect 1756 -85 1790 -51
rect 1756 -153 1790 -119
rect 1756 -221 1790 -187
rect 1756 -289 1790 -255
rect 1756 -357 1790 -323
rect 1756 -425 1790 -391
rect 1756 -493 1790 -459
rect -1790 -561 -1756 -527
rect 1756 -561 1790 -527
rect -1683 -683 -1649 -649
rect -1615 -683 -1581 -649
rect -1547 -683 -1513 -649
rect -1479 -683 -1445 -649
rect -1411 -683 -1377 -649
rect -1343 -683 -1309 -649
rect -1275 -683 -1241 -649
rect -1207 -683 -1173 -649
rect -1139 -683 -1105 -649
rect -1071 -683 -1037 -649
rect -1003 -683 -969 -649
rect -935 -683 -901 -649
rect -867 -683 -833 -649
rect -799 -683 -765 -649
rect -731 -683 -697 -649
rect -663 -683 -629 -649
rect -595 -683 -561 -649
rect -527 -683 -493 -649
rect -459 -683 -425 -649
rect -391 -683 -357 -649
rect -323 -683 -289 -649
rect -255 -683 -221 -649
rect -187 -683 -153 -649
rect -119 -683 -85 -649
rect -51 -683 -17 -649
rect 17 -683 51 -649
rect 85 -683 119 -649
rect 153 -683 187 -649
rect 221 -683 255 -649
rect 289 -683 323 -649
rect 357 -683 391 -649
rect 425 -683 459 -649
rect 493 -683 527 -649
rect 561 -683 595 -649
rect 629 -683 663 -649
rect 697 -683 731 -649
rect 765 -683 799 -649
rect 833 -683 867 -649
rect 901 -683 935 -649
rect 969 -683 1003 -649
rect 1037 -683 1071 -649
rect 1105 -683 1139 -649
rect 1173 -683 1207 -649
rect 1241 -683 1275 -649
rect 1309 -683 1343 -649
rect 1377 -683 1411 -649
rect 1445 -683 1479 -649
rect 1513 -683 1547 -649
rect 1581 -683 1615 -649
rect 1649 -683 1683 -649
<< poly >>
rect -1630 581 -1530 597
rect -1630 547 -1597 581
rect -1563 547 -1530 581
rect -1630 500 -1530 547
rect -1472 581 -1372 597
rect -1472 547 -1439 581
rect -1405 547 -1372 581
rect -1472 500 -1372 547
rect -1314 581 -1214 597
rect -1314 547 -1281 581
rect -1247 547 -1214 581
rect -1314 500 -1214 547
rect -1156 581 -1056 597
rect -1156 547 -1123 581
rect -1089 547 -1056 581
rect -1156 500 -1056 547
rect -998 581 -898 597
rect -998 547 -965 581
rect -931 547 -898 581
rect -998 500 -898 547
rect -840 581 -740 597
rect -840 547 -807 581
rect -773 547 -740 581
rect -840 500 -740 547
rect -682 581 -582 597
rect -682 547 -649 581
rect -615 547 -582 581
rect -682 500 -582 547
rect -524 581 -424 597
rect -524 547 -491 581
rect -457 547 -424 581
rect -524 500 -424 547
rect -366 581 -266 597
rect -366 547 -333 581
rect -299 547 -266 581
rect -366 500 -266 547
rect -208 581 -108 597
rect -208 547 -175 581
rect -141 547 -108 581
rect -208 500 -108 547
rect -50 581 50 597
rect -50 547 -17 581
rect 17 547 50 581
rect -50 500 50 547
rect 108 581 208 597
rect 108 547 141 581
rect 175 547 208 581
rect 108 500 208 547
rect 266 581 366 597
rect 266 547 299 581
rect 333 547 366 581
rect 266 500 366 547
rect 424 581 524 597
rect 424 547 457 581
rect 491 547 524 581
rect 424 500 524 547
rect 582 581 682 597
rect 582 547 615 581
rect 649 547 682 581
rect 582 500 682 547
rect 740 581 840 597
rect 740 547 773 581
rect 807 547 840 581
rect 740 500 840 547
rect 898 581 998 597
rect 898 547 931 581
rect 965 547 998 581
rect 898 500 998 547
rect 1056 581 1156 597
rect 1056 547 1089 581
rect 1123 547 1156 581
rect 1056 500 1156 547
rect 1214 581 1314 597
rect 1214 547 1247 581
rect 1281 547 1314 581
rect 1214 500 1314 547
rect 1372 581 1472 597
rect 1372 547 1405 581
rect 1439 547 1472 581
rect 1372 500 1472 547
rect 1530 581 1630 597
rect 1530 547 1563 581
rect 1597 547 1630 581
rect 1530 500 1630 547
rect -1630 -547 -1530 -500
rect -1630 -581 -1597 -547
rect -1563 -581 -1530 -547
rect -1630 -597 -1530 -581
rect -1472 -547 -1372 -500
rect -1472 -581 -1439 -547
rect -1405 -581 -1372 -547
rect -1472 -597 -1372 -581
rect -1314 -547 -1214 -500
rect -1314 -581 -1281 -547
rect -1247 -581 -1214 -547
rect -1314 -597 -1214 -581
rect -1156 -547 -1056 -500
rect -1156 -581 -1123 -547
rect -1089 -581 -1056 -547
rect -1156 -597 -1056 -581
rect -998 -547 -898 -500
rect -998 -581 -965 -547
rect -931 -581 -898 -547
rect -998 -597 -898 -581
rect -840 -547 -740 -500
rect -840 -581 -807 -547
rect -773 -581 -740 -547
rect -840 -597 -740 -581
rect -682 -547 -582 -500
rect -682 -581 -649 -547
rect -615 -581 -582 -547
rect -682 -597 -582 -581
rect -524 -547 -424 -500
rect -524 -581 -491 -547
rect -457 -581 -424 -547
rect -524 -597 -424 -581
rect -366 -547 -266 -500
rect -366 -581 -333 -547
rect -299 -581 -266 -547
rect -366 -597 -266 -581
rect -208 -547 -108 -500
rect -208 -581 -175 -547
rect -141 -581 -108 -547
rect -208 -597 -108 -581
rect -50 -547 50 -500
rect -50 -581 -17 -547
rect 17 -581 50 -547
rect -50 -597 50 -581
rect 108 -547 208 -500
rect 108 -581 141 -547
rect 175 -581 208 -547
rect 108 -597 208 -581
rect 266 -547 366 -500
rect 266 -581 299 -547
rect 333 -581 366 -547
rect 266 -597 366 -581
rect 424 -547 524 -500
rect 424 -581 457 -547
rect 491 -581 524 -547
rect 424 -597 524 -581
rect 582 -547 682 -500
rect 582 -581 615 -547
rect 649 -581 682 -547
rect 582 -597 682 -581
rect 740 -547 840 -500
rect 740 -581 773 -547
rect 807 -581 840 -547
rect 740 -597 840 -581
rect 898 -547 998 -500
rect 898 -581 931 -547
rect 965 -581 998 -547
rect 898 -597 998 -581
rect 1056 -547 1156 -500
rect 1056 -581 1089 -547
rect 1123 -581 1156 -547
rect 1056 -597 1156 -581
rect 1214 -547 1314 -500
rect 1214 -581 1247 -547
rect 1281 -581 1314 -547
rect 1214 -597 1314 -581
rect 1372 -547 1472 -500
rect 1372 -581 1405 -547
rect 1439 -581 1472 -547
rect 1372 -597 1472 -581
rect 1530 -547 1630 -500
rect 1530 -581 1563 -547
rect 1597 -581 1630 -547
rect 1530 -597 1630 -581
<< polycont >>
rect -1597 547 -1563 581
rect -1439 547 -1405 581
rect -1281 547 -1247 581
rect -1123 547 -1089 581
rect -965 547 -931 581
rect -807 547 -773 581
rect -649 547 -615 581
rect -491 547 -457 581
rect -333 547 -299 581
rect -175 547 -141 581
rect -17 547 17 581
rect 141 547 175 581
rect 299 547 333 581
rect 457 547 491 581
rect 615 547 649 581
rect 773 547 807 581
rect 931 547 965 581
rect 1089 547 1123 581
rect 1247 547 1281 581
rect 1405 547 1439 581
rect 1563 547 1597 581
rect -1597 -581 -1563 -547
rect -1439 -581 -1405 -547
rect -1281 -581 -1247 -547
rect -1123 -581 -1089 -547
rect -965 -581 -931 -547
rect -807 -581 -773 -547
rect -649 -581 -615 -547
rect -491 -581 -457 -547
rect -333 -581 -299 -547
rect -175 -581 -141 -547
rect -17 -581 17 -547
rect 141 -581 175 -547
rect 299 -581 333 -547
rect 457 -581 491 -547
rect 615 -581 649 -547
rect 773 -581 807 -547
rect 931 -581 965 -547
rect 1089 -581 1123 -547
rect 1247 -581 1281 -547
rect 1405 -581 1439 -547
rect 1563 -581 1597 -547
<< locali >>
rect -1790 649 -1683 683
rect -1649 649 -1615 683
rect -1581 649 -1547 683
rect -1513 649 -1479 683
rect -1445 649 -1411 683
rect -1377 649 -1343 683
rect -1309 649 -1275 683
rect -1241 649 -1207 683
rect -1173 649 -1139 683
rect -1105 649 -1071 683
rect -1037 649 -1003 683
rect -969 649 -935 683
rect -901 649 -867 683
rect -833 649 -799 683
rect -765 649 -731 683
rect -697 649 -663 683
rect -629 649 -595 683
rect -561 649 -527 683
rect -493 649 -459 683
rect -425 649 -391 683
rect -357 649 -323 683
rect -289 649 -255 683
rect -221 649 -187 683
rect -153 649 -119 683
rect -85 649 -51 683
rect -17 649 17 683
rect 51 649 85 683
rect 119 649 153 683
rect 187 649 221 683
rect 255 649 289 683
rect 323 649 357 683
rect 391 649 425 683
rect 459 649 493 683
rect 527 649 561 683
rect 595 649 629 683
rect 663 649 697 683
rect 731 649 765 683
rect 799 649 833 683
rect 867 649 901 683
rect 935 649 969 683
rect 1003 649 1037 683
rect 1071 649 1105 683
rect 1139 649 1173 683
rect 1207 649 1241 683
rect 1275 649 1309 683
rect 1343 649 1377 683
rect 1411 649 1445 683
rect 1479 649 1513 683
rect 1547 649 1581 683
rect 1615 649 1649 683
rect 1683 649 1790 683
rect -1790 561 -1756 649
rect -1630 547 -1597 581
rect -1563 547 -1530 581
rect -1472 547 -1439 581
rect -1405 547 -1372 581
rect -1314 547 -1281 581
rect -1247 547 -1214 581
rect -1156 547 -1123 581
rect -1089 547 -1056 581
rect -998 547 -965 581
rect -931 547 -898 581
rect -840 547 -807 581
rect -773 547 -740 581
rect -682 547 -649 581
rect -615 547 -582 581
rect -524 547 -491 581
rect -457 547 -424 581
rect -366 547 -333 581
rect -299 547 -266 581
rect -208 547 -175 581
rect -141 547 -108 581
rect -50 547 -17 581
rect 17 547 50 581
rect 108 547 141 581
rect 175 547 208 581
rect 266 547 299 581
rect 333 547 366 581
rect 424 547 457 581
rect 491 547 524 581
rect 582 547 615 581
rect 649 547 682 581
rect 740 547 773 581
rect 807 547 840 581
rect 898 547 931 581
rect 965 547 998 581
rect 1056 547 1089 581
rect 1123 547 1156 581
rect 1214 547 1247 581
rect 1281 547 1314 581
rect 1372 547 1405 581
rect 1439 547 1472 581
rect 1530 547 1563 581
rect 1597 547 1630 581
rect 1756 561 1790 649
rect -1790 493 -1756 527
rect -1790 425 -1756 459
rect -1790 357 -1756 391
rect -1790 289 -1756 323
rect -1790 221 -1756 255
rect -1790 153 -1756 187
rect -1790 85 -1756 119
rect -1790 17 -1756 51
rect -1790 -51 -1756 -17
rect -1790 -119 -1756 -85
rect -1790 -187 -1756 -153
rect -1790 -255 -1756 -221
rect -1790 -323 -1756 -289
rect -1790 -391 -1756 -357
rect -1790 -459 -1756 -425
rect -1790 -527 -1756 -493
rect -1676 485 -1642 504
rect -1676 413 -1642 425
rect -1676 341 -1642 357
rect -1676 269 -1642 289
rect -1676 197 -1642 221
rect -1676 125 -1642 153
rect -1676 53 -1642 85
rect -1676 -17 -1642 17
rect -1676 -85 -1642 -53
rect -1676 -153 -1642 -125
rect -1676 -221 -1642 -197
rect -1676 -289 -1642 -269
rect -1676 -357 -1642 -341
rect -1676 -425 -1642 -413
rect -1676 -504 -1642 -485
rect -1518 485 -1484 504
rect -1518 413 -1484 425
rect -1518 341 -1484 357
rect -1518 269 -1484 289
rect -1518 197 -1484 221
rect -1518 125 -1484 153
rect -1518 53 -1484 85
rect -1518 -17 -1484 17
rect -1518 -85 -1484 -53
rect -1518 -153 -1484 -125
rect -1518 -221 -1484 -197
rect -1518 -289 -1484 -269
rect -1518 -357 -1484 -341
rect -1518 -425 -1484 -413
rect -1518 -504 -1484 -485
rect -1360 485 -1326 504
rect -1360 413 -1326 425
rect -1360 341 -1326 357
rect -1360 269 -1326 289
rect -1360 197 -1326 221
rect -1360 125 -1326 153
rect -1360 53 -1326 85
rect -1360 -17 -1326 17
rect -1360 -85 -1326 -53
rect -1360 -153 -1326 -125
rect -1360 -221 -1326 -197
rect -1360 -289 -1326 -269
rect -1360 -357 -1326 -341
rect -1360 -425 -1326 -413
rect -1360 -504 -1326 -485
rect -1202 485 -1168 504
rect -1202 413 -1168 425
rect -1202 341 -1168 357
rect -1202 269 -1168 289
rect -1202 197 -1168 221
rect -1202 125 -1168 153
rect -1202 53 -1168 85
rect -1202 -17 -1168 17
rect -1202 -85 -1168 -53
rect -1202 -153 -1168 -125
rect -1202 -221 -1168 -197
rect -1202 -289 -1168 -269
rect -1202 -357 -1168 -341
rect -1202 -425 -1168 -413
rect -1202 -504 -1168 -485
rect -1044 485 -1010 504
rect -1044 413 -1010 425
rect -1044 341 -1010 357
rect -1044 269 -1010 289
rect -1044 197 -1010 221
rect -1044 125 -1010 153
rect -1044 53 -1010 85
rect -1044 -17 -1010 17
rect -1044 -85 -1010 -53
rect -1044 -153 -1010 -125
rect -1044 -221 -1010 -197
rect -1044 -289 -1010 -269
rect -1044 -357 -1010 -341
rect -1044 -425 -1010 -413
rect -1044 -504 -1010 -485
rect -886 485 -852 504
rect -886 413 -852 425
rect -886 341 -852 357
rect -886 269 -852 289
rect -886 197 -852 221
rect -886 125 -852 153
rect -886 53 -852 85
rect -886 -17 -852 17
rect -886 -85 -852 -53
rect -886 -153 -852 -125
rect -886 -221 -852 -197
rect -886 -289 -852 -269
rect -886 -357 -852 -341
rect -886 -425 -852 -413
rect -886 -504 -852 -485
rect -728 485 -694 504
rect -728 413 -694 425
rect -728 341 -694 357
rect -728 269 -694 289
rect -728 197 -694 221
rect -728 125 -694 153
rect -728 53 -694 85
rect -728 -17 -694 17
rect -728 -85 -694 -53
rect -728 -153 -694 -125
rect -728 -221 -694 -197
rect -728 -289 -694 -269
rect -728 -357 -694 -341
rect -728 -425 -694 -413
rect -728 -504 -694 -485
rect -570 485 -536 504
rect -570 413 -536 425
rect -570 341 -536 357
rect -570 269 -536 289
rect -570 197 -536 221
rect -570 125 -536 153
rect -570 53 -536 85
rect -570 -17 -536 17
rect -570 -85 -536 -53
rect -570 -153 -536 -125
rect -570 -221 -536 -197
rect -570 -289 -536 -269
rect -570 -357 -536 -341
rect -570 -425 -536 -413
rect -570 -504 -536 -485
rect -412 485 -378 504
rect -412 413 -378 425
rect -412 341 -378 357
rect -412 269 -378 289
rect -412 197 -378 221
rect -412 125 -378 153
rect -412 53 -378 85
rect -412 -17 -378 17
rect -412 -85 -378 -53
rect -412 -153 -378 -125
rect -412 -221 -378 -197
rect -412 -289 -378 -269
rect -412 -357 -378 -341
rect -412 -425 -378 -413
rect -412 -504 -378 -485
rect -254 485 -220 504
rect -254 413 -220 425
rect -254 341 -220 357
rect -254 269 -220 289
rect -254 197 -220 221
rect -254 125 -220 153
rect -254 53 -220 85
rect -254 -17 -220 17
rect -254 -85 -220 -53
rect -254 -153 -220 -125
rect -254 -221 -220 -197
rect -254 -289 -220 -269
rect -254 -357 -220 -341
rect -254 -425 -220 -413
rect -254 -504 -220 -485
rect -96 485 -62 504
rect -96 413 -62 425
rect -96 341 -62 357
rect -96 269 -62 289
rect -96 197 -62 221
rect -96 125 -62 153
rect -96 53 -62 85
rect -96 -17 -62 17
rect -96 -85 -62 -53
rect -96 -153 -62 -125
rect -96 -221 -62 -197
rect -96 -289 -62 -269
rect -96 -357 -62 -341
rect -96 -425 -62 -413
rect -96 -504 -62 -485
rect 62 485 96 504
rect 62 413 96 425
rect 62 341 96 357
rect 62 269 96 289
rect 62 197 96 221
rect 62 125 96 153
rect 62 53 96 85
rect 62 -17 96 17
rect 62 -85 96 -53
rect 62 -153 96 -125
rect 62 -221 96 -197
rect 62 -289 96 -269
rect 62 -357 96 -341
rect 62 -425 96 -413
rect 62 -504 96 -485
rect 220 485 254 504
rect 220 413 254 425
rect 220 341 254 357
rect 220 269 254 289
rect 220 197 254 221
rect 220 125 254 153
rect 220 53 254 85
rect 220 -17 254 17
rect 220 -85 254 -53
rect 220 -153 254 -125
rect 220 -221 254 -197
rect 220 -289 254 -269
rect 220 -357 254 -341
rect 220 -425 254 -413
rect 220 -504 254 -485
rect 378 485 412 504
rect 378 413 412 425
rect 378 341 412 357
rect 378 269 412 289
rect 378 197 412 221
rect 378 125 412 153
rect 378 53 412 85
rect 378 -17 412 17
rect 378 -85 412 -53
rect 378 -153 412 -125
rect 378 -221 412 -197
rect 378 -289 412 -269
rect 378 -357 412 -341
rect 378 -425 412 -413
rect 378 -504 412 -485
rect 536 485 570 504
rect 536 413 570 425
rect 536 341 570 357
rect 536 269 570 289
rect 536 197 570 221
rect 536 125 570 153
rect 536 53 570 85
rect 536 -17 570 17
rect 536 -85 570 -53
rect 536 -153 570 -125
rect 536 -221 570 -197
rect 536 -289 570 -269
rect 536 -357 570 -341
rect 536 -425 570 -413
rect 536 -504 570 -485
rect 694 485 728 504
rect 694 413 728 425
rect 694 341 728 357
rect 694 269 728 289
rect 694 197 728 221
rect 694 125 728 153
rect 694 53 728 85
rect 694 -17 728 17
rect 694 -85 728 -53
rect 694 -153 728 -125
rect 694 -221 728 -197
rect 694 -289 728 -269
rect 694 -357 728 -341
rect 694 -425 728 -413
rect 694 -504 728 -485
rect 852 485 886 504
rect 852 413 886 425
rect 852 341 886 357
rect 852 269 886 289
rect 852 197 886 221
rect 852 125 886 153
rect 852 53 886 85
rect 852 -17 886 17
rect 852 -85 886 -53
rect 852 -153 886 -125
rect 852 -221 886 -197
rect 852 -289 886 -269
rect 852 -357 886 -341
rect 852 -425 886 -413
rect 852 -504 886 -485
rect 1010 485 1044 504
rect 1010 413 1044 425
rect 1010 341 1044 357
rect 1010 269 1044 289
rect 1010 197 1044 221
rect 1010 125 1044 153
rect 1010 53 1044 85
rect 1010 -17 1044 17
rect 1010 -85 1044 -53
rect 1010 -153 1044 -125
rect 1010 -221 1044 -197
rect 1010 -289 1044 -269
rect 1010 -357 1044 -341
rect 1010 -425 1044 -413
rect 1010 -504 1044 -485
rect 1168 485 1202 504
rect 1168 413 1202 425
rect 1168 341 1202 357
rect 1168 269 1202 289
rect 1168 197 1202 221
rect 1168 125 1202 153
rect 1168 53 1202 85
rect 1168 -17 1202 17
rect 1168 -85 1202 -53
rect 1168 -153 1202 -125
rect 1168 -221 1202 -197
rect 1168 -289 1202 -269
rect 1168 -357 1202 -341
rect 1168 -425 1202 -413
rect 1168 -504 1202 -485
rect 1326 485 1360 504
rect 1326 413 1360 425
rect 1326 341 1360 357
rect 1326 269 1360 289
rect 1326 197 1360 221
rect 1326 125 1360 153
rect 1326 53 1360 85
rect 1326 -17 1360 17
rect 1326 -85 1360 -53
rect 1326 -153 1360 -125
rect 1326 -221 1360 -197
rect 1326 -289 1360 -269
rect 1326 -357 1360 -341
rect 1326 -425 1360 -413
rect 1326 -504 1360 -485
rect 1484 485 1518 504
rect 1484 413 1518 425
rect 1484 341 1518 357
rect 1484 269 1518 289
rect 1484 197 1518 221
rect 1484 125 1518 153
rect 1484 53 1518 85
rect 1484 -17 1518 17
rect 1484 -85 1518 -53
rect 1484 -153 1518 -125
rect 1484 -221 1518 -197
rect 1484 -289 1518 -269
rect 1484 -357 1518 -341
rect 1484 -425 1518 -413
rect 1484 -504 1518 -485
rect 1642 485 1676 504
rect 1642 413 1676 425
rect 1642 341 1676 357
rect 1642 269 1676 289
rect 1642 197 1676 221
rect 1642 125 1676 153
rect 1642 53 1676 85
rect 1642 -17 1676 17
rect 1642 -85 1676 -53
rect 1642 -153 1676 -125
rect 1642 -221 1676 -197
rect 1642 -289 1676 -269
rect 1642 -357 1676 -341
rect 1642 -425 1676 -413
rect 1642 -504 1676 -485
rect 1756 493 1790 527
rect 1756 425 1790 459
rect 1756 357 1790 391
rect 1756 289 1790 323
rect 1756 221 1790 255
rect 1756 153 1790 187
rect 1756 85 1790 119
rect 1756 17 1790 51
rect 1756 -51 1790 -17
rect 1756 -119 1790 -85
rect 1756 -187 1790 -153
rect 1756 -255 1790 -221
rect 1756 -323 1790 -289
rect 1756 -391 1790 -357
rect 1756 -459 1790 -425
rect 1756 -527 1790 -493
rect -1790 -649 -1756 -561
rect -1630 -581 -1597 -547
rect -1563 -581 -1530 -547
rect -1472 -581 -1439 -547
rect -1405 -581 -1372 -547
rect -1314 -581 -1281 -547
rect -1247 -581 -1214 -547
rect -1156 -581 -1123 -547
rect -1089 -581 -1056 -547
rect -998 -581 -965 -547
rect -931 -581 -898 -547
rect -840 -581 -807 -547
rect -773 -581 -740 -547
rect -682 -581 -649 -547
rect -615 -581 -582 -547
rect -524 -581 -491 -547
rect -457 -581 -424 -547
rect -366 -581 -333 -547
rect -299 -581 -266 -547
rect -208 -581 -175 -547
rect -141 -581 -108 -547
rect -50 -581 -17 -547
rect 17 -581 50 -547
rect 108 -581 141 -547
rect 175 -581 208 -547
rect 266 -581 299 -547
rect 333 -581 366 -547
rect 424 -581 457 -547
rect 491 -581 524 -547
rect 582 -581 615 -547
rect 649 -581 682 -547
rect 740 -581 773 -547
rect 807 -581 840 -547
rect 898 -581 931 -547
rect 965 -581 998 -547
rect 1056 -581 1089 -547
rect 1123 -581 1156 -547
rect 1214 -581 1247 -547
rect 1281 -581 1314 -547
rect 1372 -581 1405 -547
rect 1439 -581 1472 -547
rect 1530 -581 1563 -547
rect 1597 -581 1630 -547
rect 1756 -649 1790 -561
rect -1790 -683 -1683 -649
rect -1649 -683 -1615 -649
rect -1581 -683 -1547 -649
rect -1513 -683 -1479 -649
rect -1445 -683 -1411 -649
rect -1377 -683 -1343 -649
rect -1309 -683 -1275 -649
rect -1241 -683 -1207 -649
rect -1173 -683 -1139 -649
rect -1105 -683 -1071 -649
rect -1037 -683 -1003 -649
rect -969 -683 -935 -649
rect -901 -683 -867 -649
rect -833 -683 -799 -649
rect -765 -683 -731 -649
rect -697 -683 -663 -649
rect -629 -683 -595 -649
rect -561 -683 -527 -649
rect -493 -683 -459 -649
rect -425 -683 -391 -649
rect -357 -683 -323 -649
rect -289 -683 -255 -649
rect -221 -683 -187 -649
rect -153 -683 -119 -649
rect -85 -683 -51 -649
rect -17 -683 17 -649
rect 51 -683 85 -649
rect 119 -683 153 -649
rect 187 -683 221 -649
rect 255 -683 289 -649
rect 323 -683 357 -649
rect 391 -683 425 -649
rect 459 -683 493 -649
rect 527 -683 561 -649
rect 595 -683 629 -649
rect 663 -683 697 -649
rect 731 -683 765 -649
rect 799 -683 833 -649
rect 867 -683 901 -649
rect 935 -683 969 -649
rect 1003 -683 1037 -649
rect 1071 -683 1105 -649
rect 1139 -683 1173 -649
rect 1207 -683 1241 -649
rect 1275 -683 1309 -649
rect 1343 -683 1377 -649
rect 1411 -683 1445 -649
rect 1479 -683 1513 -649
rect 1547 -683 1581 -649
rect 1615 -683 1649 -649
rect 1683 -683 1790 -649
<< viali >>
rect -1597 547 -1563 581
rect -1439 547 -1405 581
rect -1281 547 -1247 581
rect -1123 547 -1089 581
rect -965 547 -931 581
rect -807 547 -773 581
rect -649 547 -615 581
rect -491 547 -457 581
rect -333 547 -299 581
rect -175 547 -141 581
rect -17 547 17 581
rect 141 547 175 581
rect 299 547 333 581
rect 457 547 491 581
rect 615 547 649 581
rect 773 547 807 581
rect 931 547 965 581
rect 1089 547 1123 581
rect 1247 547 1281 581
rect 1405 547 1439 581
rect 1563 547 1597 581
rect -1676 459 -1642 485
rect -1676 451 -1642 459
rect -1676 391 -1642 413
rect -1676 379 -1642 391
rect -1676 323 -1642 341
rect -1676 307 -1642 323
rect -1676 255 -1642 269
rect -1676 235 -1642 255
rect -1676 187 -1642 197
rect -1676 163 -1642 187
rect -1676 119 -1642 125
rect -1676 91 -1642 119
rect -1676 51 -1642 53
rect -1676 19 -1642 51
rect -1676 -51 -1642 -19
rect -1676 -53 -1642 -51
rect -1676 -119 -1642 -91
rect -1676 -125 -1642 -119
rect -1676 -187 -1642 -163
rect -1676 -197 -1642 -187
rect -1676 -255 -1642 -235
rect -1676 -269 -1642 -255
rect -1676 -323 -1642 -307
rect -1676 -341 -1642 -323
rect -1676 -391 -1642 -379
rect -1676 -413 -1642 -391
rect -1676 -459 -1642 -451
rect -1676 -485 -1642 -459
rect -1518 459 -1484 485
rect -1518 451 -1484 459
rect -1518 391 -1484 413
rect -1518 379 -1484 391
rect -1518 323 -1484 341
rect -1518 307 -1484 323
rect -1518 255 -1484 269
rect -1518 235 -1484 255
rect -1518 187 -1484 197
rect -1518 163 -1484 187
rect -1518 119 -1484 125
rect -1518 91 -1484 119
rect -1518 51 -1484 53
rect -1518 19 -1484 51
rect -1518 -51 -1484 -19
rect -1518 -53 -1484 -51
rect -1518 -119 -1484 -91
rect -1518 -125 -1484 -119
rect -1518 -187 -1484 -163
rect -1518 -197 -1484 -187
rect -1518 -255 -1484 -235
rect -1518 -269 -1484 -255
rect -1518 -323 -1484 -307
rect -1518 -341 -1484 -323
rect -1518 -391 -1484 -379
rect -1518 -413 -1484 -391
rect -1518 -459 -1484 -451
rect -1518 -485 -1484 -459
rect -1360 459 -1326 485
rect -1360 451 -1326 459
rect -1360 391 -1326 413
rect -1360 379 -1326 391
rect -1360 323 -1326 341
rect -1360 307 -1326 323
rect -1360 255 -1326 269
rect -1360 235 -1326 255
rect -1360 187 -1326 197
rect -1360 163 -1326 187
rect -1360 119 -1326 125
rect -1360 91 -1326 119
rect -1360 51 -1326 53
rect -1360 19 -1326 51
rect -1360 -51 -1326 -19
rect -1360 -53 -1326 -51
rect -1360 -119 -1326 -91
rect -1360 -125 -1326 -119
rect -1360 -187 -1326 -163
rect -1360 -197 -1326 -187
rect -1360 -255 -1326 -235
rect -1360 -269 -1326 -255
rect -1360 -323 -1326 -307
rect -1360 -341 -1326 -323
rect -1360 -391 -1326 -379
rect -1360 -413 -1326 -391
rect -1360 -459 -1326 -451
rect -1360 -485 -1326 -459
rect -1202 459 -1168 485
rect -1202 451 -1168 459
rect -1202 391 -1168 413
rect -1202 379 -1168 391
rect -1202 323 -1168 341
rect -1202 307 -1168 323
rect -1202 255 -1168 269
rect -1202 235 -1168 255
rect -1202 187 -1168 197
rect -1202 163 -1168 187
rect -1202 119 -1168 125
rect -1202 91 -1168 119
rect -1202 51 -1168 53
rect -1202 19 -1168 51
rect -1202 -51 -1168 -19
rect -1202 -53 -1168 -51
rect -1202 -119 -1168 -91
rect -1202 -125 -1168 -119
rect -1202 -187 -1168 -163
rect -1202 -197 -1168 -187
rect -1202 -255 -1168 -235
rect -1202 -269 -1168 -255
rect -1202 -323 -1168 -307
rect -1202 -341 -1168 -323
rect -1202 -391 -1168 -379
rect -1202 -413 -1168 -391
rect -1202 -459 -1168 -451
rect -1202 -485 -1168 -459
rect -1044 459 -1010 485
rect -1044 451 -1010 459
rect -1044 391 -1010 413
rect -1044 379 -1010 391
rect -1044 323 -1010 341
rect -1044 307 -1010 323
rect -1044 255 -1010 269
rect -1044 235 -1010 255
rect -1044 187 -1010 197
rect -1044 163 -1010 187
rect -1044 119 -1010 125
rect -1044 91 -1010 119
rect -1044 51 -1010 53
rect -1044 19 -1010 51
rect -1044 -51 -1010 -19
rect -1044 -53 -1010 -51
rect -1044 -119 -1010 -91
rect -1044 -125 -1010 -119
rect -1044 -187 -1010 -163
rect -1044 -197 -1010 -187
rect -1044 -255 -1010 -235
rect -1044 -269 -1010 -255
rect -1044 -323 -1010 -307
rect -1044 -341 -1010 -323
rect -1044 -391 -1010 -379
rect -1044 -413 -1010 -391
rect -1044 -459 -1010 -451
rect -1044 -485 -1010 -459
rect -886 459 -852 485
rect -886 451 -852 459
rect -886 391 -852 413
rect -886 379 -852 391
rect -886 323 -852 341
rect -886 307 -852 323
rect -886 255 -852 269
rect -886 235 -852 255
rect -886 187 -852 197
rect -886 163 -852 187
rect -886 119 -852 125
rect -886 91 -852 119
rect -886 51 -852 53
rect -886 19 -852 51
rect -886 -51 -852 -19
rect -886 -53 -852 -51
rect -886 -119 -852 -91
rect -886 -125 -852 -119
rect -886 -187 -852 -163
rect -886 -197 -852 -187
rect -886 -255 -852 -235
rect -886 -269 -852 -255
rect -886 -323 -852 -307
rect -886 -341 -852 -323
rect -886 -391 -852 -379
rect -886 -413 -852 -391
rect -886 -459 -852 -451
rect -886 -485 -852 -459
rect -728 459 -694 485
rect -728 451 -694 459
rect -728 391 -694 413
rect -728 379 -694 391
rect -728 323 -694 341
rect -728 307 -694 323
rect -728 255 -694 269
rect -728 235 -694 255
rect -728 187 -694 197
rect -728 163 -694 187
rect -728 119 -694 125
rect -728 91 -694 119
rect -728 51 -694 53
rect -728 19 -694 51
rect -728 -51 -694 -19
rect -728 -53 -694 -51
rect -728 -119 -694 -91
rect -728 -125 -694 -119
rect -728 -187 -694 -163
rect -728 -197 -694 -187
rect -728 -255 -694 -235
rect -728 -269 -694 -255
rect -728 -323 -694 -307
rect -728 -341 -694 -323
rect -728 -391 -694 -379
rect -728 -413 -694 -391
rect -728 -459 -694 -451
rect -728 -485 -694 -459
rect -570 459 -536 485
rect -570 451 -536 459
rect -570 391 -536 413
rect -570 379 -536 391
rect -570 323 -536 341
rect -570 307 -536 323
rect -570 255 -536 269
rect -570 235 -536 255
rect -570 187 -536 197
rect -570 163 -536 187
rect -570 119 -536 125
rect -570 91 -536 119
rect -570 51 -536 53
rect -570 19 -536 51
rect -570 -51 -536 -19
rect -570 -53 -536 -51
rect -570 -119 -536 -91
rect -570 -125 -536 -119
rect -570 -187 -536 -163
rect -570 -197 -536 -187
rect -570 -255 -536 -235
rect -570 -269 -536 -255
rect -570 -323 -536 -307
rect -570 -341 -536 -323
rect -570 -391 -536 -379
rect -570 -413 -536 -391
rect -570 -459 -536 -451
rect -570 -485 -536 -459
rect -412 459 -378 485
rect -412 451 -378 459
rect -412 391 -378 413
rect -412 379 -378 391
rect -412 323 -378 341
rect -412 307 -378 323
rect -412 255 -378 269
rect -412 235 -378 255
rect -412 187 -378 197
rect -412 163 -378 187
rect -412 119 -378 125
rect -412 91 -378 119
rect -412 51 -378 53
rect -412 19 -378 51
rect -412 -51 -378 -19
rect -412 -53 -378 -51
rect -412 -119 -378 -91
rect -412 -125 -378 -119
rect -412 -187 -378 -163
rect -412 -197 -378 -187
rect -412 -255 -378 -235
rect -412 -269 -378 -255
rect -412 -323 -378 -307
rect -412 -341 -378 -323
rect -412 -391 -378 -379
rect -412 -413 -378 -391
rect -412 -459 -378 -451
rect -412 -485 -378 -459
rect -254 459 -220 485
rect -254 451 -220 459
rect -254 391 -220 413
rect -254 379 -220 391
rect -254 323 -220 341
rect -254 307 -220 323
rect -254 255 -220 269
rect -254 235 -220 255
rect -254 187 -220 197
rect -254 163 -220 187
rect -254 119 -220 125
rect -254 91 -220 119
rect -254 51 -220 53
rect -254 19 -220 51
rect -254 -51 -220 -19
rect -254 -53 -220 -51
rect -254 -119 -220 -91
rect -254 -125 -220 -119
rect -254 -187 -220 -163
rect -254 -197 -220 -187
rect -254 -255 -220 -235
rect -254 -269 -220 -255
rect -254 -323 -220 -307
rect -254 -341 -220 -323
rect -254 -391 -220 -379
rect -254 -413 -220 -391
rect -254 -459 -220 -451
rect -254 -485 -220 -459
rect -96 459 -62 485
rect -96 451 -62 459
rect -96 391 -62 413
rect -96 379 -62 391
rect -96 323 -62 341
rect -96 307 -62 323
rect -96 255 -62 269
rect -96 235 -62 255
rect -96 187 -62 197
rect -96 163 -62 187
rect -96 119 -62 125
rect -96 91 -62 119
rect -96 51 -62 53
rect -96 19 -62 51
rect -96 -51 -62 -19
rect -96 -53 -62 -51
rect -96 -119 -62 -91
rect -96 -125 -62 -119
rect -96 -187 -62 -163
rect -96 -197 -62 -187
rect -96 -255 -62 -235
rect -96 -269 -62 -255
rect -96 -323 -62 -307
rect -96 -341 -62 -323
rect -96 -391 -62 -379
rect -96 -413 -62 -391
rect -96 -459 -62 -451
rect -96 -485 -62 -459
rect 62 459 96 485
rect 62 451 96 459
rect 62 391 96 413
rect 62 379 96 391
rect 62 323 96 341
rect 62 307 96 323
rect 62 255 96 269
rect 62 235 96 255
rect 62 187 96 197
rect 62 163 96 187
rect 62 119 96 125
rect 62 91 96 119
rect 62 51 96 53
rect 62 19 96 51
rect 62 -51 96 -19
rect 62 -53 96 -51
rect 62 -119 96 -91
rect 62 -125 96 -119
rect 62 -187 96 -163
rect 62 -197 96 -187
rect 62 -255 96 -235
rect 62 -269 96 -255
rect 62 -323 96 -307
rect 62 -341 96 -323
rect 62 -391 96 -379
rect 62 -413 96 -391
rect 62 -459 96 -451
rect 62 -485 96 -459
rect 220 459 254 485
rect 220 451 254 459
rect 220 391 254 413
rect 220 379 254 391
rect 220 323 254 341
rect 220 307 254 323
rect 220 255 254 269
rect 220 235 254 255
rect 220 187 254 197
rect 220 163 254 187
rect 220 119 254 125
rect 220 91 254 119
rect 220 51 254 53
rect 220 19 254 51
rect 220 -51 254 -19
rect 220 -53 254 -51
rect 220 -119 254 -91
rect 220 -125 254 -119
rect 220 -187 254 -163
rect 220 -197 254 -187
rect 220 -255 254 -235
rect 220 -269 254 -255
rect 220 -323 254 -307
rect 220 -341 254 -323
rect 220 -391 254 -379
rect 220 -413 254 -391
rect 220 -459 254 -451
rect 220 -485 254 -459
rect 378 459 412 485
rect 378 451 412 459
rect 378 391 412 413
rect 378 379 412 391
rect 378 323 412 341
rect 378 307 412 323
rect 378 255 412 269
rect 378 235 412 255
rect 378 187 412 197
rect 378 163 412 187
rect 378 119 412 125
rect 378 91 412 119
rect 378 51 412 53
rect 378 19 412 51
rect 378 -51 412 -19
rect 378 -53 412 -51
rect 378 -119 412 -91
rect 378 -125 412 -119
rect 378 -187 412 -163
rect 378 -197 412 -187
rect 378 -255 412 -235
rect 378 -269 412 -255
rect 378 -323 412 -307
rect 378 -341 412 -323
rect 378 -391 412 -379
rect 378 -413 412 -391
rect 378 -459 412 -451
rect 378 -485 412 -459
rect 536 459 570 485
rect 536 451 570 459
rect 536 391 570 413
rect 536 379 570 391
rect 536 323 570 341
rect 536 307 570 323
rect 536 255 570 269
rect 536 235 570 255
rect 536 187 570 197
rect 536 163 570 187
rect 536 119 570 125
rect 536 91 570 119
rect 536 51 570 53
rect 536 19 570 51
rect 536 -51 570 -19
rect 536 -53 570 -51
rect 536 -119 570 -91
rect 536 -125 570 -119
rect 536 -187 570 -163
rect 536 -197 570 -187
rect 536 -255 570 -235
rect 536 -269 570 -255
rect 536 -323 570 -307
rect 536 -341 570 -323
rect 536 -391 570 -379
rect 536 -413 570 -391
rect 536 -459 570 -451
rect 536 -485 570 -459
rect 694 459 728 485
rect 694 451 728 459
rect 694 391 728 413
rect 694 379 728 391
rect 694 323 728 341
rect 694 307 728 323
rect 694 255 728 269
rect 694 235 728 255
rect 694 187 728 197
rect 694 163 728 187
rect 694 119 728 125
rect 694 91 728 119
rect 694 51 728 53
rect 694 19 728 51
rect 694 -51 728 -19
rect 694 -53 728 -51
rect 694 -119 728 -91
rect 694 -125 728 -119
rect 694 -187 728 -163
rect 694 -197 728 -187
rect 694 -255 728 -235
rect 694 -269 728 -255
rect 694 -323 728 -307
rect 694 -341 728 -323
rect 694 -391 728 -379
rect 694 -413 728 -391
rect 694 -459 728 -451
rect 694 -485 728 -459
rect 852 459 886 485
rect 852 451 886 459
rect 852 391 886 413
rect 852 379 886 391
rect 852 323 886 341
rect 852 307 886 323
rect 852 255 886 269
rect 852 235 886 255
rect 852 187 886 197
rect 852 163 886 187
rect 852 119 886 125
rect 852 91 886 119
rect 852 51 886 53
rect 852 19 886 51
rect 852 -51 886 -19
rect 852 -53 886 -51
rect 852 -119 886 -91
rect 852 -125 886 -119
rect 852 -187 886 -163
rect 852 -197 886 -187
rect 852 -255 886 -235
rect 852 -269 886 -255
rect 852 -323 886 -307
rect 852 -341 886 -323
rect 852 -391 886 -379
rect 852 -413 886 -391
rect 852 -459 886 -451
rect 852 -485 886 -459
rect 1010 459 1044 485
rect 1010 451 1044 459
rect 1010 391 1044 413
rect 1010 379 1044 391
rect 1010 323 1044 341
rect 1010 307 1044 323
rect 1010 255 1044 269
rect 1010 235 1044 255
rect 1010 187 1044 197
rect 1010 163 1044 187
rect 1010 119 1044 125
rect 1010 91 1044 119
rect 1010 51 1044 53
rect 1010 19 1044 51
rect 1010 -51 1044 -19
rect 1010 -53 1044 -51
rect 1010 -119 1044 -91
rect 1010 -125 1044 -119
rect 1010 -187 1044 -163
rect 1010 -197 1044 -187
rect 1010 -255 1044 -235
rect 1010 -269 1044 -255
rect 1010 -323 1044 -307
rect 1010 -341 1044 -323
rect 1010 -391 1044 -379
rect 1010 -413 1044 -391
rect 1010 -459 1044 -451
rect 1010 -485 1044 -459
rect 1168 459 1202 485
rect 1168 451 1202 459
rect 1168 391 1202 413
rect 1168 379 1202 391
rect 1168 323 1202 341
rect 1168 307 1202 323
rect 1168 255 1202 269
rect 1168 235 1202 255
rect 1168 187 1202 197
rect 1168 163 1202 187
rect 1168 119 1202 125
rect 1168 91 1202 119
rect 1168 51 1202 53
rect 1168 19 1202 51
rect 1168 -51 1202 -19
rect 1168 -53 1202 -51
rect 1168 -119 1202 -91
rect 1168 -125 1202 -119
rect 1168 -187 1202 -163
rect 1168 -197 1202 -187
rect 1168 -255 1202 -235
rect 1168 -269 1202 -255
rect 1168 -323 1202 -307
rect 1168 -341 1202 -323
rect 1168 -391 1202 -379
rect 1168 -413 1202 -391
rect 1168 -459 1202 -451
rect 1168 -485 1202 -459
rect 1326 459 1360 485
rect 1326 451 1360 459
rect 1326 391 1360 413
rect 1326 379 1360 391
rect 1326 323 1360 341
rect 1326 307 1360 323
rect 1326 255 1360 269
rect 1326 235 1360 255
rect 1326 187 1360 197
rect 1326 163 1360 187
rect 1326 119 1360 125
rect 1326 91 1360 119
rect 1326 51 1360 53
rect 1326 19 1360 51
rect 1326 -51 1360 -19
rect 1326 -53 1360 -51
rect 1326 -119 1360 -91
rect 1326 -125 1360 -119
rect 1326 -187 1360 -163
rect 1326 -197 1360 -187
rect 1326 -255 1360 -235
rect 1326 -269 1360 -255
rect 1326 -323 1360 -307
rect 1326 -341 1360 -323
rect 1326 -391 1360 -379
rect 1326 -413 1360 -391
rect 1326 -459 1360 -451
rect 1326 -485 1360 -459
rect 1484 459 1518 485
rect 1484 451 1518 459
rect 1484 391 1518 413
rect 1484 379 1518 391
rect 1484 323 1518 341
rect 1484 307 1518 323
rect 1484 255 1518 269
rect 1484 235 1518 255
rect 1484 187 1518 197
rect 1484 163 1518 187
rect 1484 119 1518 125
rect 1484 91 1518 119
rect 1484 51 1518 53
rect 1484 19 1518 51
rect 1484 -51 1518 -19
rect 1484 -53 1518 -51
rect 1484 -119 1518 -91
rect 1484 -125 1518 -119
rect 1484 -187 1518 -163
rect 1484 -197 1518 -187
rect 1484 -255 1518 -235
rect 1484 -269 1518 -255
rect 1484 -323 1518 -307
rect 1484 -341 1518 -323
rect 1484 -391 1518 -379
rect 1484 -413 1518 -391
rect 1484 -459 1518 -451
rect 1484 -485 1518 -459
rect 1642 459 1676 485
rect 1642 451 1676 459
rect 1642 391 1676 413
rect 1642 379 1676 391
rect 1642 323 1676 341
rect 1642 307 1676 323
rect 1642 255 1676 269
rect 1642 235 1676 255
rect 1642 187 1676 197
rect 1642 163 1676 187
rect 1642 119 1676 125
rect 1642 91 1676 119
rect 1642 51 1676 53
rect 1642 19 1676 51
rect 1642 -51 1676 -19
rect 1642 -53 1676 -51
rect 1642 -119 1676 -91
rect 1642 -125 1676 -119
rect 1642 -187 1676 -163
rect 1642 -197 1676 -187
rect 1642 -255 1676 -235
rect 1642 -269 1676 -255
rect 1642 -323 1676 -307
rect 1642 -341 1676 -323
rect 1642 -391 1676 -379
rect 1642 -413 1676 -391
rect 1642 -459 1676 -451
rect 1642 -485 1676 -459
rect -1597 -581 -1563 -547
rect -1439 -581 -1405 -547
rect -1281 -581 -1247 -547
rect -1123 -581 -1089 -547
rect -965 -581 -931 -547
rect -807 -581 -773 -547
rect -649 -581 -615 -547
rect -491 -581 -457 -547
rect -333 -581 -299 -547
rect -175 -581 -141 -547
rect -17 -581 17 -547
rect 141 -581 175 -547
rect 299 -581 333 -547
rect 457 -581 491 -547
rect 615 -581 649 -547
rect 773 -581 807 -547
rect 931 -581 965 -547
rect 1089 -581 1123 -547
rect 1247 -581 1281 -547
rect 1405 -581 1439 -547
rect 1563 -581 1597 -547
<< metal1 >>
rect -1626 581 -1534 587
rect -1626 547 -1597 581
rect -1563 547 -1534 581
rect -1626 541 -1534 547
rect -1468 581 -1376 587
rect -1468 547 -1439 581
rect -1405 547 -1376 581
rect -1468 541 -1376 547
rect -1310 581 -1218 587
rect -1310 547 -1281 581
rect -1247 547 -1218 581
rect -1310 541 -1218 547
rect -1152 581 -1060 587
rect -1152 547 -1123 581
rect -1089 547 -1060 581
rect -1152 541 -1060 547
rect -994 581 -902 587
rect -994 547 -965 581
rect -931 547 -902 581
rect -994 541 -902 547
rect -836 581 -744 587
rect -836 547 -807 581
rect -773 547 -744 581
rect -836 541 -744 547
rect -678 581 -586 587
rect -678 547 -649 581
rect -615 547 -586 581
rect -678 541 -586 547
rect -520 581 -428 587
rect -520 547 -491 581
rect -457 547 -428 581
rect -520 541 -428 547
rect -362 581 -270 587
rect -362 547 -333 581
rect -299 547 -270 581
rect -362 541 -270 547
rect -204 581 -112 587
rect -204 547 -175 581
rect -141 547 -112 581
rect -204 541 -112 547
rect -46 581 46 587
rect -46 547 -17 581
rect 17 547 46 581
rect -46 541 46 547
rect 112 581 204 587
rect 112 547 141 581
rect 175 547 204 581
rect 112 541 204 547
rect 270 581 362 587
rect 270 547 299 581
rect 333 547 362 581
rect 270 541 362 547
rect 428 581 520 587
rect 428 547 457 581
rect 491 547 520 581
rect 428 541 520 547
rect 586 581 678 587
rect 586 547 615 581
rect 649 547 678 581
rect 586 541 678 547
rect 744 581 836 587
rect 744 547 773 581
rect 807 547 836 581
rect 744 541 836 547
rect 902 581 994 587
rect 902 547 931 581
rect 965 547 994 581
rect 902 541 994 547
rect 1060 581 1152 587
rect 1060 547 1089 581
rect 1123 547 1152 581
rect 1060 541 1152 547
rect 1218 581 1310 587
rect 1218 547 1247 581
rect 1281 547 1310 581
rect 1218 541 1310 547
rect 1376 581 1468 587
rect 1376 547 1405 581
rect 1439 547 1468 581
rect 1376 541 1468 547
rect 1534 581 1626 587
rect 1534 547 1563 581
rect 1597 547 1626 581
rect 1534 541 1626 547
rect -1682 485 -1636 500
rect -1682 451 -1676 485
rect -1642 451 -1636 485
rect -1682 413 -1636 451
rect -1682 379 -1676 413
rect -1642 379 -1636 413
rect -1682 341 -1636 379
rect -1682 307 -1676 341
rect -1642 307 -1636 341
rect -1682 269 -1636 307
rect -1682 235 -1676 269
rect -1642 235 -1636 269
rect -1682 197 -1636 235
rect -1682 163 -1676 197
rect -1642 163 -1636 197
rect -1682 125 -1636 163
rect -1682 91 -1676 125
rect -1642 91 -1636 125
rect -1682 53 -1636 91
rect -1682 19 -1676 53
rect -1642 19 -1636 53
rect -1682 -19 -1636 19
rect -1682 -53 -1676 -19
rect -1642 -53 -1636 -19
rect -1682 -91 -1636 -53
rect -1682 -125 -1676 -91
rect -1642 -125 -1636 -91
rect -1682 -163 -1636 -125
rect -1682 -197 -1676 -163
rect -1642 -197 -1636 -163
rect -1682 -235 -1636 -197
rect -1682 -269 -1676 -235
rect -1642 -269 -1636 -235
rect -1682 -307 -1636 -269
rect -1682 -341 -1676 -307
rect -1642 -341 -1636 -307
rect -1682 -379 -1636 -341
rect -1682 -413 -1676 -379
rect -1642 -413 -1636 -379
rect -1682 -451 -1636 -413
rect -1682 -485 -1676 -451
rect -1642 -485 -1636 -451
rect -1682 -500 -1636 -485
rect -1524 485 -1478 500
rect -1524 451 -1518 485
rect -1484 451 -1478 485
rect -1524 413 -1478 451
rect -1524 379 -1518 413
rect -1484 379 -1478 413
rect -1524 341 -1478 379
rect -1524 307 -1518 341
rect -1484 307 -1478 341
rect -1524 269 -1478 307
rect -1524 235 -1518 269
rect -1484 235 -1478 269
rect -1524 197 -1478 235
rect -1524 163 -1518 197
rect -1484 163 -1478 197
rect -1524 125 -1478 163
rect -1524 91 -1518 125
rect -1484 91 -1478 125
rect -1524 53 -1478 91
rect -1524 19 -1518 53
rect -1484 19 -1478 53
rect -1524 -19 -1478 19
rect -1524 -53 -1518 -19
rect -1484 -53 -1478 -19
rect -1524 -91 -1478 -53
rect -1524 -125 -1518 -91
rect -1484 -125 -1478 -91
rect -1524 -163 -1478 -125
rect -1524 -197 -1518 -163
rect -1484 -197 -1478 -163
rect -1524 -235 -1478 -197
rect -1524 -269 -1518 -235
rect -1484 -269 -1478 -235
rect -1524 -307 -1478 -269
rect -1524 -341 -1518 -307
rect -1484 -341 -1478 -307
rect -1524 -379 -1478 -341
rect -1524 -413 -1518 -379
rect -1484 -413 -1478 -379
rect -1524 -451 -1478 -413
rect -1524 -485 -1518 -451
rect -1484 -485 -1478 -451
rect -1524 -500 -1478 -485
rect -1366 485 -1320 500
rect -1366 451 -1360 485
rect -1326 451 -1320 485
rect -1366 413 -1320 451
rect -1366 379 -1360 413
rect -1326 379 -1320 413
rect -1366 341 -1320 379
rect -1366 307 -1360 341
rect -1326 307 -1320 341
rect -1366 269 -1320 307
rect -1366 235 -1360 269
rect -1326 235 -1320 269
rect -1366 197 -1320 235
rect -1366 163 -1360 197
rect -1326 163 -1320 197
rect -1366 125 -1320 163
rect -1366 91 -1360 125
rect -1326 91 -1320 125
rect -1366 53 -1320 91
rect -1366 19 -1360 53
rect -1326 19 -1320 53
rect -1366 -19 -1320 19
rect -1366 -53 -1360 -19
rect -1326 -53 -1320 -19
rect -1366 -91 -1320 -53
rect -1366 -125 -1360 -91
rect -1326 -125 -1320 -91
rect -1366 -163 -1320 -125
rect -1366 -197 -1360 -163
rect -1326 -197 -1320 -163
rect -1366 -235 -1320 -197
rect -1366 -269 -1360 -235
rect -1326 -269 -1320 -235
rect -1366 -307 -1320 -269
rect -1366 -341 -1360 -307
rect -1326 -341 -1320 -307
rect -1366 -379 -1320 -341
rect -1366 -413 -1360 -379
rect -1326 -413 -1320 -379
rect -1366 -451 -1320 -413
rect -1366 -485 -1360 -451
rect -1326 -485 -1320 -451
rect -1366 -500 -1320 -485
rect -1208 485 -1162 500
rect -1208 451 -1202 485
rect -1168 451 -1162 485
rect -1208 413 -1162 451
rect -1208 379 -1202 413
rect -1168 379 -1162 413
rect -1208 341 -1162 379
rect -1208 307 -1202 341
rect -1168 307 -1162 341
rect -1208 269 -1162 307
rect -1208 235 -1202 269
rect -1168 235 -1162 269
rect -1208 197 -1162 235
rect -1208 163 -1202 197
rect -1168 163 -1162 197
rect -1208 125 -1162 163
rect -1208 91 -1202 125
rect -1168 91 -1162 125
rect -1208 53 -1162 91
rect -1208 19 -1202 53
rect -1168 19 -1162 53
rect -1208 -19 -1162 19
rect -1208 -53 -1202 -19
rect -1168 -53 -1162 -19
rect -1208 -91 -1162 -53
rect -1208 -125 -1202 -91
rect -1168 -125 -1162 -91
rect -1208 -163 -1162 -125
rect -1208 -197 -1202 -163
rect -1168 -197 -1162 -163
rect -1208 -235 -1162 -197
rect -1208 -269 -1202 -235
rect -1168 -269 -1162 -235
rect -1208 -307 -1162 -269
rect -1208 -341 -1202 -307
rect -1168 -341 -1162 -307
rect -1208 -379 -1162 -341
rect -1208 -413 -1202 -379
rect -1168 -413 -1162 -379
rect -1208 -451 -1162 -413
rect -1208 -485 -1202 -451
rect -1168 -485 -1162 -451
rect -1208 -500 -1162 -485
rect -1050 485 -1004 500
rect -1050 451 -1044 485
rect -1010 451 -1004 485
rect -1050 413 -1004 451
rect -1050 379 -1044 413
rect -1010 379 -1004 413
rect -1050 341 -1004 379
rect -1050 307 -1044 341
rect -1010 307 -1004 341
rect -1050 269 -1004 307
rect -1050 235 -1044 269
rect -1010 235 -1004 269
rect -1050 197 -1004 235
rect -1050 163 -1044 197
rect -1010 163 -1004 197
rect -1050 125 -1004 163
rect -1050 91 -1044 125
rect -1010 91 -1004 125
rect -1050 53 -1004 91
rect -1050 19 -1044 53
rect -1010 19 -1004 53
rect -1050 -19 -1004 19
rect -1050 -53 -1044 -19
rect -1010 -53 -1004 -19
rect -1050 -91 -1004 -53
rect -1050 -125 -1044 -91
rect -1010 -125 -1004 -91
rect -1050 -163 -1004 -125
rect -1050 -197 -1044 -163
rect -1010 -197 -1004 -163
rect -1050 -235 -1004 -197
rect -1050 -269 -1044 -235
rect -1010 -269 -1004 -235
rect -1050 -307 -1004 -269
rect -1050 -341 -1044 -307
rect -1010 -341 -1004 -307
rect -1050 -379 -1004 -341
rect -1050 -413 -1044 -379
rect -1010 -413 -1004 -379
rect -1050 -451 -1004 -413
rect -1050 -485 -1044 -451
rect -1010 -485 -1004 -451
rect -1050 -500 -1004 -485
rect -892 485 -846 500
rect -892 451 -886 485
rect -852 451 -846 485
rect -892 413 -846 451
rect -892 379 -886 413
rect -852 379 -846 413
rect -892 341 -846 379
rect -892 307 -886 341
rect -852 307 -846 341
rect -892 269 -846 307
rect -892 235 -886 269
rect -852 235 -846 269
rect -892 197 -846 235
rect -892 163 -886 197
rect -852 163 -846 197
rect -892 125 -846 163
rect -892 91 -886 125
rect -852 91 -846 125
rect -892 53 -846 91
rect -892 19 -886 53
rect -852 19 -846 53
rect -892 -19 -846 19
rect -892 -53 -886 -19
rect -852 -53 -846 -19
rect -892 -91 -846 -53
rect -892 -125 -886 -91
rect -852 -125 -846 -91
rect -892 -163 -846 -125
rect -892 -197 -886 -163
rect -852 -197 -846 -163
rect -892 -235 -846 -197
rect -892 -269 -886 -235
rect -852 -269 -846 -235
rect -892 -307 -846 -269
rect -892 -341 -886 -307
rect -852 -341 -846 -307
rect -892 -379 -846 -341
rect -892 -413 -886 -379
rect -852 -413 -846 -379
rect -892 -451 -846 -413
rect -892 -485 -886 -451
rect -852 -485 -846 -451
rect -892 -500 -846 -485
rect -734 485 -688 500
rect -734 451 -728 485
rect -694 451 -688 485
rect -734 413 -688 451
rect -734 379 -728 413
rect -694 379 -688 413
rect -734 341 -688 379
rect -734 307 -728 341
rect -694 307 -688 341
rect -734 269 -688 307
rect -734 235 -728 269
rect -694 235 -688 269
rect -734 197 -688 235
rect -734 163 -728 197
rect -694 163 -688 197
rect -734 125 -688 163
rect -734 91 -728 125
rect -694 91 -688 125
rect -734 53 -688 91
rect -734 19 -728 53
rect -694 19 -688 53
rect -734 -19 -688 19
rect -734 -53 -728 -19
rect -694 -53 -688 -19
rect -734 -91 -688 -53
rect -734 -125 -728 -91
rect -694 -125 -688 -91
rect -734 -163 -688 -125
rect -734 -197 -728 -163
rect -694 -197 -688 -163
rect -734 -235 -688 -197
rect -734 -269 -728 -235
rect -694 -269 -688 -235
rect -734 -307 -688 -269
rect -734 -341 -728 -307
rect -694 -341 -688 -307
rect -734 -379 -688 -341
rect -734 -413 -728 -379
rect -694 -413 -688 -379
rect -734 -451 -688 -413
rect -734 -485 -728 -451
rect -694 -485 -688 -451
rect -734 -500 -688 -485
rect -576 485 -530 500
rect -576 451 -570 485
rect -536 451 -530 485
rect -576 413 -530 451
rect -576 379 -570 413
rect -536 379 -530 413
rect -576 341 -530 379
rect -576 307 -570 341
rect -536 307 -530 341
rect -576 269 -530 307
rect -576 235 -570 269
rect -536 235 -530 269
rect -576 197 -530 235
rect -576 163 -570 197
rect -536 163 -530 197
rect -576 125 -530 163
rect -576 91 -570 125
rect -536 91 -530 125
rect -576 53 -530 91
rect -576 19 -570 53
rect -536 19 -530 53
rect -576 -19 -530 19
rect -576 -53 -570 -19
rect -536 -53 -530 -19
rect -576 -91 -530 -53
rect -576 -125 -570 -91
rect -536 -125 -530 -91
rect -576 -163 -530 -125
rect -576 -197 -570 -163
rect -536 -197 -530 -163
rect -576 -235 -530 -197
rect -576 -269 -570 -235
rect -536 -269 -530 -235
rect -576 -307 -530 -269
rect -576 -341 -570 -307
rect -536 -341 -530 -307
rect -576 -379 -530 -341
rect -576 -413 -570 -379
rect -536 -413 -530 -379
rect -576 -451 -530 -413
rect -576 -485 -570 -451
rect -536 -485 -530 -451
rect -576 -500 -530 -485
rect -418 485 -372 500
rect -418 451 -412 485
rect -378 451 -372 485
rect -418 413 -372 451
rect -418 379 -412 413
rect -378 379 -372 413
rect -418 341 -372 379
rect -418 307 -412 341
rect -378 307 -372 341
rect -418 269 -372 307
rect -418 235 -412 269
rect -378 235 -372 269
rect -418 197 -372 235
rect -418 163 -412 197
rect -378 163 -372 197
rect -418 125 -372 163
rect -418 91 -412 125
rect -378 91 -372 125
rect -418 53 -372 91
rect -418 19 -412 53
rect -378 19 -372 53
rect -418 -19 -372 19
rect -418 -53 -412 -19
rect -378 -53 -372 -19
rect -418 -91 -372 -53
rect -418 -125 -412 -91
rect -378 -125 -372 -91
rect -418 -163 -372 -125
rect -418 -197 -412 -163
rect -378 -197 -372 -163
rect -418 -235 -372 -197
rect -418 -269 -412 -235
rect -378 -269 -372 -235
rect -418 -307 -372 -269
rect -418 -341 -412 -307
rect -378 -341 -372 -307
rect -418 -379 -372 -341
rect -418 -413 -412 -379
rect -378 -413 -372 -379
rect -418 -451 -372 -413
rect -418 -485 -412 -451
rect -378 -485 -372 -451
rect -418 -500 -372 -485
rect -260 485 -214 500
rect -260 451 -254 485
rect -220 451 -214 485
rect -260 413 -214 451
rect -260 379 -254 413
rect -220 379 -214 413
rect -260 341 -214 379
rect -260 307 -254 341
rect -220 307 -214 341
rect -260 269 -214 307
rect -260 235 -254 269
rect -220 235 -214 269
rect -260 197 -214 235
rect -260 163 -254 197
rect -220 163 -214 197
rect -260 125 -214 163
rect -260 91 -254 125
rect -220 91 -214 125
rect -260 53 -214 91
rect -260 19 -254 53
rect -220 19 -214 53
rect -260 -19 -214 19
rect -260 -53 -254 -19
rect -220 -53 -214 -19
rect -260 -91 -214 -53
rect -260 -125 -254 -91
rect -220 -125 -214 -91
rect -260 -163 -214 -125
rect -260 -197 -254 -163
rect -220 -197 -214 -163
rect -260 -235 -214 -197
rect -260 -269 -254 -235
rect -220 -269 -214 -235
rect -260 -307 -214 -269
rect -260 -341 -254 -307
rect -220 -341 -214 -307
rect -260 -379 -214 -341
rect -260 -413 -254 -379
rect -220 -413 -214 -379
rect -260 -451 -214 -413
rect -260 -485 -254 -451
rect -220 -485 -214 -451
rect -260 -500 -214 -485
rect -102 485 -56 500
rect -102 451 -96 485
rect -62 451 -56 485
rect -102 413 -56 451
rect -102 379 -96 413
rect -62 379 -56 413
rect -102 341 -56 379
rect -102 307 -96 341
rect -62 307 -56 341
rect -102 269 -56 307
rect -102 235 -96 269
rect -62 235 -56 269
rect -102 197 -56 235
rect -102 163 -96 197
rect -62 163 -56 197
rect -102 125 -56 163
rect -102 91 -96 125
rect -62 91 -56 125
rect -102 53 -56 91
rect -102 19 -96 53
rect -62 19 -56 53
rect -102 -19 -56 19
rect -102 -53 -96 -19
rect -62 -53 -56 -19
rect -102 -91 -56 -53
rect -102 -125 -96 -91
rect -62 -125 -56 -91
rect -102 -163 -56 -125
rect -102 -197 -96 -163
rect -62 -197 -56 -163
rect -102 -235 -56 -197
rect -102 -269 -96 -235
rect -62 -269 -56 -235
rect -102 -307 -56 -269
rect -102 -341 -96 -307
rect -62 -341 -56 -307
rect -102 -379 -56 -341
rect -102 -413 -96 -379
rect -62 -413 -56 -379
rect -102 -451 -56 -413
rect -102 -485 -96 -451
rect -62 -485 -56 -451
rect -102 -500 -56 -485
rect 56 485 102 500
rect 56 451 62 485
rect 96 451 102 485
rect 56 413 102 451
rect 56 379 62 413
rect 96 379 102 413
rect 56 341 102 379
rect 56 307 62 341
rect 96 307 102 341
rect 56 269 102 307
rect 56 235 62 269
rect 96 235 102 269
rect 56 197 102 235
rect 56 163 62 197
rect 96 163 102 197
rect 56 125 102 163
rect 56 91 62 125
rect 96 91 102 125
rect 56 53 102 91
rect 56 19 62 53
rect 96 19 102 53
rect 56 -19 102 19
rect 56 -53 62 -19
rect 96 -53 102 -19
rect 56 -91 102 -53
rect 56 -125 62 -91
rect 96 -125 102 -91
rect 56 -163 102 -125
rect 56 -197 62 -163
rect 96 -197 102 -163
rect 56 -235 102 -197
rect 56 -269 62 -235
rect 96 -269 102 -235
rect 56 -307 102 -269
rect 56 -341 62 -307
rect 96 -341 102 -307
rect 56 -379 102 -341
rect 56 -413 62 -379
rect 96 -413 102 -379
rect 56 -451 102 -413
rect 56 -485 62 -451
rect 96 -485 102 -451
rect 56 -500 102 -485
rect 214 485 260 500
rect 214 451 220 485
rect 254 451 260 485
rect 214 413 260 451
rect 214 379 220 413
rect 254 379 260 413
rect 214 341 260 379
rect 214 307 220 341
rect 254 307 260 341
rect 214 269 260 307
rect 214 235 220 269
rect 254 235 260 269
rect 214 197 260 235
rect 214 163 220 197
rect 254 163 260 197
rect 214 125 260 163
rect 214 91 220 125
rect 254 91 260 125
rect 214 53 260 91
rect 214 19 220 53
rect 254 19 260 53
rect 214 -19 260 19
rect 214 -53 220 -19
rect 254 -53 260 -19
rect 214 -91 260 -53
rect 214 -125 220 -91
rect 254 -125 260 -91
rect 214 -163 260 -125
rect 214 -197 220 -163
rect 254 -197 260 -163
rect 214 -235 260 -197
rect 214 -269 220 -235
rect 254 -269 260 -235
rect 214 -307 260 -269
rect 214 -341 220 -307
rect 254 -341 260 -307
rect 214 -379 260 -341
rect 214 -413 220 -379
rect 254 -413 260 -379
rect 214 -451 260 -413
rect 214 -485 220 -451
rect 254 -485 260 -451
rect 214 -500 260 -485
rect 372 485 418 500
rect 372 451 378 485
rect 412 451 418 485
rect 372 413 418 451
rect 372 379 378 413
rect 412 379 418 413
rect 372 341 418 379
rect 372 307 378 341
rect 412 307 418 341
rect 372 269 418 307
rect 372 235 378 269
rect 412 235 418 269
rect 372 197 418 235
rect 372 163 378 197
rect 412 163 418 197
rect 372 125 418 163
rect 372 91 378 125
rect 412 91 418 125
rect 372 53 418 91
rect 372 19 378 53
rect 412 19 418 53
rect 372 -19 418 19
rect 372 -53 378 -19
rect 412 -53 418 -19
rect 372 -91 418 -53
rect 372 -125 378 -91
rect 412 -125 418 -91
rect 372 -163 418 -125
rect 372 -197 378 -163
rect 412 -197 418 -163
rect 372 -235 418 -197
rect 372 -269 378 -235
rect 412 -269 418 -235
rect 372 -307 418 -269
rect 372 -341 378 -307
rect 412 -341 418 -307
rect 372 -379 418 -341
rect 372 -413 378 -379
rect 412 -413 418 -379
rect 372 -451 418 -413
rect 372 -485 378 -451
rect 412 -485 418 -451
rect 372 -500 418 -485
rect 530 485 576 500
rect 530 451 536 485
rect 570 451 576 485
rect 530 413 576 451
rect 530 379 536 413
rect 570 379 576 413
rect 530 341 576 379
rect 530 307 536 341
rect 570 307 576 341
rect 530 269 576 307
rect 530 235 536 269
rect 570 235 576 269
rect 530 197 576 235
rect 530 163 536 197
rect 570 163 576 197
rect 530 125 576 163
rect 530 91 536 125
rect 570 91 576 125
rect 530 53 576 91
rect 530 19 536 53
rect 570 19 576 53
rect 530 -19 576 19
rect 530 -53 536 -19
rect 570 -53 576 -19
rect 530 -91 576 -53
rect 530 -125 536 -91
rect 570 -125 576 -91
rect 530 -163 576 -125
rect 530 -197 536 -163
rect 570 -197 576 -163
rect 530 -235 576 -197
rect 530 -269 536 -235
rect 570 -269 576 -235
rect 530 -307 576 -269
rect 530 -341 536 -307
rect 570 -341 576 -307
rect 530 -379 576 -341
rect 530 -413 536 -379
rect 570 -413 576 -379
rect 530 -451 576 -413
rect 530 -485 536 -451
rect 570 -485 576 -451
rect 530 -500 576 -485
rect 688 485 734 500
rect 688 451 694 485
rect 728 451 734 485
rect 688 413 734 451
rect 688 379 694 413
rect 728 379 734 413
rect 688 341 734 379
rect 688 307 694 341
rect 728 307 734 341
rect 688 269 734 307
rect 688 235 694 269
rect 728 235 734 269
rect 688 197 734 235
rect 688 163 694 197
rect 728 163 734 197
rect 688 125 734 163
rect 688 91 694 125
rect 728 91 734 125
rect 688 53 734 91
rect 688 19 694 53
rect 728 19 734 53
rect 688 -19 734 19
rect 688 -53 694 -19
rect 728 -53 734 -19
rect 688 -91 734 -53
rect 688 -125 694 -91
rect 728 -125 734 -91
rect 688 -163 734 -125
rect 688 -197 694 -163
rect 728 -197 734 -163
rect 688 -235 734 -197
rect 688 -269 694 -235
rect 728 -269 734 -235
rect 688 -307 734 -269
rect 688 -341 694 -307
rect 728 -341 734 -307
rect 688 -379 734 -341
rect 688 -413 694 -379
rect 728 -413 734 -379
rect 688 -451 734 -413
rect 688 -485 694 -451
rect 728 -485 734 -451
rect 688 -500 734 -485
rect 846 485 892 500
rect 846 451 852 485
rect 886 451 892 485
rect 846 413 892 451
rect 846 379 852 413
rect 886 379 892 413
rect 846 341 892 379
rect 846 307 852 341
rect 886 307 892 341
rect 846 269 892 307
rect 846 235 852 269
rect 886 235 892 269
rect 846 197 892 235
rect 846 163 852 197
rect 886 163 892 197
rect 846 125 892 163
rect 846 91 852 125
rect 886 91 892 125
rect 846 53 892 91
rect 846 19 852 53
rect 886 19 892 53
rect 846 -19 892 19
rect 846 -53 852 -19
rect 886 -53 892 -19
rect 846 -91 892 -53
rect 846 -125 852 -91
rect 886 -125 892 -91
rect 846 -163 892 -125
rect 846 -197 852 -163
rect 886 -197 892 -163
rect 846 -235 892 -197
rect 846 -269 852 -235
rect 886 -269 892 -235
rect 846 -307 892 -269
rect 846 -341 852 -307
rect 886 -341 892 -307
rect 846 -379 892 -341
rect 846 -413 852 -379
rect 886 -413 892 -379
rect 846 -451 892 -413
rect 846 -485 852 -451
rect 886 -485 892 -451
rect 846 -500 892 -485
rect 1004 485 1050 500
rect 1004 451 1010 485
rect 1044 451 1050 485
rect 1004 413 1050 451
rect 1004 379 1010 413
rect 1044 379 1050 413
rect 1004 341 1050 379
rect 1004 307 1010 341
rect 1044 307 1050 341
rect 1004 269 1050 307
rect 1004 235 1010 269
rect 1044 235 1050 269
rect 1004 197 1050 235
rect 1004 163 1010 197
rect 1044 163 1050 197
rect 1004 125 1050 163
rect 1004 91 1010 125
rect 1044 91 1050 125
rect 1004 53 1050 91
rect 1004 19 1010 53
rect 1044 19 1050 53
rect 1004 -19 1050 19
rect 1004 -53 1010 -19
rect 1044 -53 1050 -19
rect 1004 -91 1050 -53
rect 1004 -125 1010 -91
rect 1044 -125 1050 -91
rect 1004 -163 1050 -125
rect 1004 -197 1010 -163
rect 1044 -197 1050 -163
rect 1004 -235 1050 -197
rect 1004 -269 1010 -235
rect 1044 -269 1050 -235
rect 1004 -307 1050 -269
rect 1004 -341 1010 -307
rect 1044 -341 1050 -307
rect 1004 -379 1050 -341
rect 1004 -413 1010 -379
rect 1044 -413 1050 -379
rect 1004 -451 1050 -413
rect 1004 -485 1010 -451
rect 1044 -485 1050 -451
rect 1004 -500 1050 -485
rect 1162 485 1208 500
rect 1162 451 1168 485
rect 1202 451 1208 485
rect 1162 413 1208 451
rect 1162 379 1168 413
rect 1202 379 1208 413
rect 1162 341 1208 379
rect 1162 307 1168 341
rect 1202 307 1208 341
rect 1162 269 1208 307
rect 1162 235 1168 269
rect 1202 235 1208 269
rect 1162 197 1208 235
rect 1162 163 1168 197
rect 1202 163 1208 197
rect 1162 125 1208 163
rect 1162 91 1168 125
rect 1202 91 1208 125
rect 1162 53 1208 91
rect 1162 19 1168 53
rect 1202 19 1208 53
rect 1162 -19 1208 19
rect 1162 -53 1168 -19
rect 1202 -53 1208 -19
rect 1162 -91 1208 -53
rect 1162 -125 1168 -91
rect 1202 -125 1208 -91
rect 1162 -163 1208 -125
rect 1162 -197 1168 -163
rect 1202 -197 1208 -163
rect 1162 -235 1208 -197
rect 1162 -269 1168 -235
rect 1202 -269 1208 -235
rect 1162 -307 1208 -269
rect 1162 -341 1168 -307
rect 1202 -341 1208 -307
rect 1162 -379 1208 -341
rect 1162 -413 1168 -379
rect 1202 -413 1208 -379
rect 1162 -451 1208 -413
rect 1162 -485 1168 -451
rect 1202 -485 1208 -451
rect 1162 -500 1208 -485
rect 1320 485 1366 500
rect 1320 451 1326 485
rect 1360 451 1366 485
rect 1320 413 1366 451
rect 1320 379 1326 413
rect 1360 379 1366 413
rect 1320 341 1366 379
rect 1320 307 1326 341
rect 1360 307 1366 341
rect 1320 269 1366 307
rect 1320 235 1326 269
rect 1360 235 1366 269
rect 1320 197 1366 235
rect 1320 163 1326 197
rect 1360 163 1366 197
rect 1320 125 1366 163
rect 1320 91 1326 125
rect 1360 91 1366 125
rect 1320 53 1366 91
rect 1320 19 1326 53
rect 1360 19 1366 53
rect 1320 -19 1366 19
rect 1320 -53 1326 -19
rect 1360 -53 1366 -19
rect 1320 -91 1366 -53
rect 1320 -125 1326 -91
rect 1360 -125 1366 -91
rect 1320 -163 1366 -125
rect 1320 -197 1326 -163
rect 1360 -197 1366 -163
rect 1320 -235 1366 -197
rect 1320 -269 1326 -235
rect 1360 -269 1366 -235
rect 1320 -307 1366 -269
rect 1320 -341 1326 -307
rect 1360 -341 1366 -307
rect 1320 -379 1366 -341
rect 1320 -413 1326 -379
rect 1360 -413 1366 -379
rect 1320 -451 1366 -413
rect 1320 -485 1326 -451
rect 1360 -485 1366 -451
rect 1320 -500 1366 -485
rect 1478 485 1524 500
rect 1478 451 1484 485
rect 1518 451 1524 485
rect 1478 413 1524 451
rect 1478 379 1484 413
rect 1518 379 1524 413
rect 1478 341 1524 379
rect 1478 307 1484 341
rect 1518 307 1524 341
rect 1478 269 1524 307
rect 1478 235 1484 269
rect 1518 235 1524 269
rect 1478 197 1524 235
rect 1478 163 1484 197
rect 1518 163 1524 197
rect 1478 125 1524 163
rect 1478 91 1484 125
rect 1518 91 1524 125
rect 1478 53 1524 91
rect 1478 19 1484 53
rect 1518 19 1524 53
rect 1478 -19 1524 19
rect 1478 -53 1484 -19
rect 1518 -53 1524 -19
rect 1478 -91 1524 -53
rect 1478 -125 1484 -91
rect 1518 -125 1524 -91
rect 1478 -163 1524 -125
rect 1478 -197 1484 -163
rect 1518 -197 1524 -163
rect 1478 -235 1524 -197
rect 1478 -269 1484 -235
rect 1518 -269 1524 -235
rect 1478 -307 1524 -269
rect 1478 -341 1484 -307
rect 1518 -341 1524 -307
rect 1478 -379 1524 -341
rect 1478 -413 1484 -379
rect 1518 -413 1524 -379
rect 1478 -451 1524 -413
rect 1478 -485 1484 -451
rect 1518 -485 1524 -451
rect 1478 -500 1524 -485
rect 1636 485 1682 500
rect 1636 451 1642 485
rect 1676 451 1682 485
rect 1636 413 1682 451
rect 1636 379 1642 413
rect 1676 379 1682 413
rect 1636 341 1682 379
rect 1636 307 1642 341
rect 1676 307 1682 341
rect 1636 269 1682 307
rect 1636 235 1642 269
rect 1676 235 1682 269
rect 1636 197 1682 235
rect 1636 163 1642 197
rect 1676 163 1682 197
rect 1636 125 1682 163
rect 1636 91 1642 125
rect 1676 91 1682 125
rect 1636 53 1682 91
rect 1636 19 1642 53
rect 1676 19 1682 53
rect 1636 -19 1682 19
rect 1636 -53 1642 -19
rect 1676 -53 1682 -19
rect 1636 -91 1682 -53
rect 1636 -125 1642 -91
rect 1676 -125 1682 -91
rect 1636 -163 1682 -125
rect 1636 -197 1642 -163
rect 1676 -197 1682 -163
rect 1636 -235 1682 -197
rect 1636 -269 1642 -235
rect 1676 -269 1682 -235
rect 1636 -307 1682 -269
rect 1636 -341 1642 -307
rect 1676 -341 1682 -307
rect 1636 -379 1682 -341
rect 1636 -413 1642 -379
rect 1676 -413 1682 -379
rect 1636 -451 1682 -413
rect 1636 -485 1642 -451
rect 1676 -485 1682 -451
rect 1636 -500 1682 -485
rect -1626 -547 -1534 -541
rect -1626 -581 -1597 -547
rect -1563 -581 -1534 -547
rect -1626 -587 -1534 -581
rect -1468 -547 -1376 -541
rect -1468 -581 -1439 -547
rect -1405 -581 -1376 -547
rect -1468 -587 -1376 -581
rect -1310 -547 -1218 -541
rect -1310 -581 -1281 -547
rect -1247 -581 -1218 -547
rect -1310 -587 -1218 -581
rect -1152 -547 -1060 -541
rect -1152 -581 -1123 -547
rect -1089 -581 -1060 -547
rect -1152 -587 -1060 -581
rect -994 -547 -902 -541
rect -994 -581 -965 -547
rect -931 -581 -902 -547
rect -994 -587 -902 -581
rect -836 -547 -744 -541
rect -836 -581 -807 -547
rect -773 -581 -744 -547
rect -836 -587 -744 -581
rect -678 -547 -586 -541
rect -678 -581 -649 -547
rect -615 -581 -586 -547
rect -678 -587 -586 -581
rect -520 -547 -428 -541
rect -520 -581 -491 -547
rect -457 -581 -428 -547
rect -520 -587 -428 -581
rect -362 -547 -270 -541
rect -362 -581 -333 -547
rect -299 -581 -270 -547
rect -362 -587 -270 -581
rect -204 -547 -112 -541
rect -204 -581 -175 -547
rect -141 -581 -112 -547
rect -204 -587 -112 -581
rect -46 -547 46 -541
rect -46 -581 -17 -547
rect 17 -581 46 -547
rect -46 -587 46 -581
rect 112 -547 204 -541
rect 112 -581 141 -547
rect 175 -581 204 -547
rect 112 -587 204 -581
rect 270 -547 362 -541
rect 270 -581 299 -547
rect 333 -581 362 -547
rect 270 -587 362 -581
rect 428 -547 520 -541
rect 428 -581 457 -547
rect 491 -581 520 -547
rect 428 -587 520 -581
rect 586 -547 678 -541
rect 586 -581 615 -547
rect 649 -581 678 -547
rect 586 -587 678 -581
rect 744 -547 836 -541
rect 744 -581 773 -547
rect 807 -581 836 -547
rect 744 -587 836 -581
rect 902 -547 994 -541
rect 902 -581 931 -547
rect 965 -581 994 -547
rect 902 -587 994 -581
rect 1060 -547 1152 -541
rect 1060 -581 1089 -547
rect 1123 -581 1152 -547
rect 1060 -587 1152 -581
rect 1218 -547 1310 -541
rect 1218 -581 1247 -547
rect 1281 -581 1310 -547
rect 1218 -587 1310 -581
rect 1376 -547 1468 -541
rect 1376 -581 1405 -547
rect 1439 -581 1468 -547
rect 1376 -587 1468 -581
rect 1534 -547 1626 -541
rect 1534 -581 1563 -547
rect 1597 -581 1626 -547
rect 1534 -587 1626 -581
<< properties >>
string FIXED_BBOX -1773 -666 1773 666
<< end >>
