magic
tech sky130A
magscale 1 2
timestamp 1716868724
<< xpolycontact >>
rect -573 6900 573 7332
rect -573 -7332 573 -6900
<< xpolyres >>
rect -573 -6900 573 6900
<< viali >>
rect -557 6918 557 7312
rect -557 -7313 557 -6919
<< metal1 >>
rect -569 7312 569 7320
rect -569 6918 -557 7312
rect 557 6918 569 7312
rect -569 6911 569 6918
rect -569 -6919 569 -6911
rect -569 -7313 -557 -6919
rect 557 -7313 569 -6919
rect -569 -7320 569 -7313
<< end >>
