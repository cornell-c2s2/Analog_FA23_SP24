magic
tech sky130A
magscale 1 2
timestamp 1713140669
<< pwell >>
rect -739 -7482 739 7482
<< psubdiff >>
rect -703 7412 -607 7446
rect 607 7412 703 7446
rect -703 7350 -669 7412
rect 669 7350 703 7412
rect -703 -7412 -669 -7350
rect 669 -7412 703 -7350
rect -703 -7446 -607 -7412
rect 607 -7446 703 -7412
<< psubdiffcont >>
rect -607 7412 607 7446
rect -703 -7350 -669 7350
rect 669 -7350 703 7350
rect -607 -7446 607 -7412
<< xpolycontact >>
rect -573 6884 573 7316
rect -573 -7316 573 -6884
<< xpolyres >>
rect -573 -6884 573 6884
<< locali >>
rect -703 7412 -607 7446
rect 607 7412 703 7446
rect -703 7350 -669 7412
rect 669 7350 703 7412
rect -703 -7412 -669 -7350
rect 669 -7412 703 -7350
rect -703 -7446 -607 -7412
rect 607 -7446 703 -7412
<< viali >>
rect -557 6901 557 7298
rect -557 -7298 557 -6901
<< metal1 >>
rect -569 7298 569 7304
rect -569 6901 -557 7298
rect 557 6901 569 7298
rect -569 6895 569 6901
rect -569 -6901 569 -6895
rect -569 -7298 -557 -6901
rect 557 -7298 569 -6901
rect -569 -7304 569 -7298
<< properties >>
string FIXED_BBOX -686 -7429 686 7429
string gencell sky130_fd_pr__res_xhigh_po_5p73
string library sky130
string parameters w 5.730 l 69.0 m 1 nx 1 wmin 5.730 lmin 0.50 rho 2000 val 24.149k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 5.730 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
