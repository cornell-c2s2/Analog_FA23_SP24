magic
tech sky130A
magscale 1 2
timestamp 1716869746
<< metal4 >>
rect -21094 38239 -14396 38280
rect -21094 32161 -14652 38239
rect -14416 32161 -14396 38239
rect -21094 32120 -14396 32161
rect -13996 38239 -7298 38280
rect -13996 32161 -7554 38239
rect -7318 32161 -7298 38239
rect -13996 32120 -7298 32161
rect -6898 38239 -200 38280
rect -6898 32161 -456 38239
rect -220 32161 -200 38239
rect -6898 32120 -200 32161
rect 200 38239 6898 38280
rect 200 32161 6642 38239
rect 6878 32161 6898 38239
rect 200 32120 6898 32161
rect 7298 38239 13996 38280
rect 7298 32161 13740 38239
rect 13976 32161 13996 38239
rect 7298 32120 13996 32161
rect 14396 38239 21094 38280
rect 14396 32161 20838 38239
rect 21074 32161 21094 38239
rect 14396 32120 21094 32161
rect -21094 31839 -14396 31880
rect -21094 25761 -14652 31839
rect -14416 25761 -14396 31839
rect -21094 25720 -14396 25761
rect -13996 31839 -7298 31880
rect -13996 25761 -7554 31839
rect -7318 25761 -7298 31839
rect -13996 25720 -7298 25761
rect -6898 31839 -200 31880
rect -6898 25761 -456 31839
rect -220 25761 -200 31839
rect -6898 25720 -200 25761
rect 200 31839 6898 31880
rect 200 25761 6642 31839
rect 6878 25761 6898 31839
rect 200 25720 6898 25761
rect 7298 31839 13996 31880
rect 7298 25761 13740 31839
rect 13976 25761 13996 31839
rect 7298 25720 13996 25761
rect 14396 31839 21094 31880
rect 14396 25761 20838 31839
rect 21074 25761 21094 31839
rect 14396 25720 21094 25761
rect -21094 25439 -14396 25480
rect -21094 19361 -14652 25439
rect -14416 19361 -14396 25439
rect -21094 19320 -14396 19361
rect -13996 25439 -7298 25480
rect -13996 19361 -7554 25439
rect -7318 19361 -7298 25439
rect -13996 19320 -7298 19361
rect -6898 25439 -200 25480
rect -6898 19361 -456 25439
rect -220 19361 -200 25439
rect -6898 19320 -200 19361
rect 200 25439 6898 25480
rect 200 19361 6642 25439
rect 6878 19361 6898 25439
rect 200 19320 6898 19361
rect 7298 25439 13996 25480
rect 7298 19361 13740 25439
rect 13976 19361 13996 25439
rect 7298 19320 13996 19361
rect 14396 25439 21094 25480
rect 14396 19361 20838 25439
rect 21074 19361 21094 25439
rect 14396 19320 21094 19361
rect -21094 19039 -14396 19080
rect -21094 12961 -14652 19039
rect -14416 12961 -14396 19039
rect -21094 12920 -14396 12961
rect -13996 19039 -7298 19080
rect -13996 12961 -7554 19039
rect -7318 12961 -7298 19039
rect -13996 12920 -7298 12961
rect -6898 19039 -200 19080
rect -6898 12961 -456 19039
rect -220 12961 -200 19039
rect -6898 12920 -200 12961
rect 200 19039 6898 19080
rect 200 12961 6642 19039
rect 6878 12961 6898 19039
rect 200 12920 6898 12961
rect 7298 19039 13996 19080
rect 7298 12961 13740 19039
rect 13976 12961 13996 19039
rect 7298 12920 13996 12961
rect 14396 19039 21094 19080
rect 14396 12961 20838 19039
rect 21074 12961 21094 19039
rect 14396 12920 21094 12961
rect -21094 12639 -14396 12680
rect -21094 6561 -14652 12639
rect -14416 6561 -14396 12639
rect -21094 6520 -14396 6561
rect -13996 12639 -7298 12680
rect -13996 6561 -7554 12639
rect -7318 6561 -7298 12639
rect -13996 6520 -7298 6561
rect -6898 12639 -200 12680
rect -6898 6561 -456 12639
rect -220 6561 -200 12639
rect -6898 6520 -200 6561
rect 200 12639 6898 12680
rect 200 6561 6642 12639
rect 6878 6561 6898 12639
rect 200 6520 6898 6561
rect 7298 12639 13996 12680
rect 7298 6561 13740 12639
rect 13976 6561 13996 12639
rect 7298 6520 13996 6561
rect 14396 12639 21094 12680
rect 14396 6561 20838 12639
rect 21074 6561 21094 12639
rect 14396 6520 21094 6561
rect -21094 6239 -14396 6280
rect -21094 161 -14652 6239
rect -14416 161 -14396 6239
rect -21094 120 -14396 161
rect -13996 6239 -7298 6280
rect -13996 161 -7554 6239
rect -7318 161 -7298 6239
rect -13996 120 -7298 161
rect -6898 6239 -200 6280
rect -6898 161 -456 6239
rect -220 161 -200 6239
rect -6898 120 -200 161
rect 200 6239 6898 6280
rect 200 161 6642 6239
rect 6878 161 6898 6239
rect 200 120 6898 161
rect 7298 6239 13996 6280
rect 7298 161 13740 6239
rect 13976 161 13996 6239
rect 7298 120 13996 161
rect 14396 6239 21094 6280
rect 14396 161 20838 6239
rect 21074 161 21094 6239
rect 14396 120 21094 161
rect -21094 -161 -14396 -120
rect -21094 -6239 -14652 -161
rect -14416 -6239 -14396 -161
rect -21094 -6280 -14396 -6239
rect -13996 -161 -7298 -120
rect -13996 -6239 -7554 -161
rect -7318 -6239 -7298 -161
rect -13996 -6280 -7298 -6239
rect -6898 -161 -200 -120
rect -6898 -6239 -456 -161
rect -220 -6239 -200 -161
rect -6898 -6280 -200 -6239
rect 200 -161 6898 -120
rect 200 -6239 6642 -161
rect 6878 -6239 6898 -161
rect 200 -6280 6898 -6239
rect 7298 -161 13996 -120
rect 7298 -6239 13740 -161
rect 13976 -6239 13996 -161
rect 7298 -6280 13996 -6239
rect 14396 -161 21094 -120
rect 14396 -6239 20838 -161
rect 21074 -6239 21094 -161
rect 14396 -6280 21094 -6239
rect -21094 -6561 -14396 -6520
rect -21094 -12639 -14652 -6561
rect -14416 -12639 -14396 -6561
rect -21094 -12680 -14396 -12639
rect -13996 -6561 -7298 -6520
rect -13996 -12639 -7554 -6561
rect -7318 -12639 -7298 -6561
rect -13996 -12680 -7298 -12639
rect -6898 -6561 -200 -6520
rect -6898 -12639 -456 -6561
rect -220 -12639 -200 -6561
rect -6898 -12680 -200 -12639
rect 200 -6561 6898 -6520
rect 200 -12639 6642 -6561
rect 6878 -12639 6898 -6561
rect 200 -12680 6898 -12639
rect 7298 -6561 13996 -6520
rect 7298 -12639 13740 -6561
rect 13976 -12639 13996 -6561
rect 7298 -12680 13996 -12639
rect 14396 -6561 21094 -6520
rect 14396 -12639 20838 -6561
rect 21074 -12639 21094 -6561
rect 14396 -12680 21094 -12639
rect -21094 -12961 -14396 -12920
rect -21094 -19039 -14652 -12961
rect -14416 -19039 -14396 -12961
rect -21094 -19080 -14396 -19039
rect -13996 -12961 -7298 -12920
rect -13996 -19039 -7554 -12961
rect -7318 -19039 -7298 -12961
rect -13996 -19080 -7298 -19039
rect -6898 -12961 -200 -12920
rect -6898 -19039 -456 -12961
rect -220 -19039 -200 -12961
rect -6898 -19080 -200 -19039
rect 200 -12961 6898 -12920
rect 200 -19039 6642 -12961
rect 6878 -19039 6898 -12961
rect 200 -19080 6898 -19039
rect 7298 -12961 13996 -12920
rect 7298 -19039 13740 -12961
rect 13976 -19039 13996 -12961
rect 7298 -19080 13996 -19039
rect 14396 -12961 21094 -12920
rect 14396 -19039 20838 -12961
rect 21074 -19039 21094 -12961
rect 14396 -19080 21094 -19039
rect -21094 -19361 -14396 -19320
rect -21094 -25439 -14652 -19361
rect -14416 -25439 -14396 -19361
rect -21094 -25480 -14396 -25439
rect -13996 -19361 -7298 -19320
rect -13996 -25439 -7554 -19361
rect -7318 -25439 -7298 -19361
rect -13996 -25480 -7298 -25439
rect -6898 -19361 -200 -19320
rect -6898 -25439 -456 -19361
rect -220 -25439 -200 -19361
rect -6898 -25480 -200 -25439
rect 200 -19361 6898 -19320
rect 200 -25439 6642 -19361
rect 6878 -25439 6898 -19361
rect 200 -25480 6898 -25439
rect 7298 -19361 13996 -19320
rect 7298 -25439 13740 -19361
rect 13976 -25439 13996 -19361
rect 7298 -25480 13996 -25439
rect 14396 -19361 21094 -19320
rect 14396 -25439 20838 -19361
rect 21074 -25439 21094 -19361
rect 14396 -25480 21094 -25439
rect -21094 -25761 -14396 -25720
rect -21094 -31839 -14652 -25761
rect -14416 -31839 -14396 -25761
rect -21094 -31880 -14396 -31839
rect -13996 -25761 -7298 -25720
rect -13996 -31839 -7554 -25761
rect -7318 -31839 -7298 -25761
rect -13996 -31880 -7298 -31839
rect -6898 -25761 -200 -25720
rect -6898 -31839 -456 -25761
rect -220 -31839 -200 -25761
rect -6898 -31880 -200 -31839
rect 200 -25761 6898 -25720
rect 200 -31839 6642 -25761
rect 6878 -31839 6898 -25761
rect 200 -31880 6898 -31839
rect 7298 -25761 13996 -25720
rect 7298 -31839 13740 -25761
rect 13976 -31839 13996 -25761
rect 7298 -31880 13996 -31839
rect 14396 -25761 21094 -25720
rect 14396 -31839 20838 -25761
rect 21074 -31839 21094 -25761
rect 14396 -31880 21094 -31839
rect -21094 -32161 -14396 -32120
rect -21094 -38239 -14652 -32161
rect -14416 -38239 -14396 -32161
rect -21094 -38280 -14396 -38239
rect -13996 -32161 -7298 -32120
rect -13996 -38239 -7554 -32161
rect -7318 -38239 -7298 -32161
rect -13996 -38280 -7298 -38239
rect -6898 -32161 -200 -32120
rect -6898 -38239 -456 -32161
rect -220 -38239 -200 -32161
rect -6898 -38280 -200 -38239
rect 200 -32161 6898 -32120
rect 200 -38239 6642 -32161
rect 6878 -38239 6898 -32161
rect 200 -38280 6898 -38239
rect 7298 -32161 13996 -32120
rect 7298 -38239 13740 -32161
rect 13976 -38239 13996 -32161
rect 7298 -38280 13996 -38239
rect 14396 -32161 21094 -32120
rect 14396 -38239 20838 -32161
rect 21074 -38239 21094 -32161
rect 14396 -38280 21094 -38239
<< via4 >>
rect -14652 32161 -14416 38239
rect -7554 32161 -7318 38239
rect -456 32161 -220 38239
rect 6642 32161 6878 38239
rect 13740 32161 13976 38239
rect 20838 32161 21074 38239
rect -14652 25761 -14416 31839
rect -7554 25761 -7318 31839
rect -456 25761 -220 31839
rect 6642 25761 6878 31839
rect 13740 25761 13976 31839
rect 20838 25761 21074 31839
rect -14652 19361 -14416 25439
rect -7554 19361 -7318 25439
rect -456 19361 -220 25439
rect 6642 19361 6878 25439
rect 13740 19361 13976 25439
rect 20838 19361 21074 25439
rect -14652 12961 -14416 19039
rect -7554 12961 -7318 19039
rect -456 12961 -220 19039
rect 6642 12961 6878 19039
rect 13740 12961 13976 19039
rect 20838 12961 21074 19039
rect -14652 6561 -14416 12639
rect -7554 6561 -7318 12639
rect -456 6561 -220 12639
rect 6642 6561 6878 12639
rect 13740 6561 13976 12639
rect 20838 6561 21074 12639
rect -14652 161 -14416 6239
rect -7554 161 -7318 6239
rect -456 161 -220 6239
rect 6642 161 6878 6239
rect 13740 161 13976 6239
rect 20838 161 21074 6239
rect -14652 -6239 -14416 -161
rect -7554 -6239 -7318 -161
rect -456 -6239 -220 -161
rect 6642 -6239 6878 -161
rect 13740 -6239 13976 -161
rect 20838 -6239 21074 -161
rect -14652 -12639 -14416 -6561
rect -7554 -12639 -7318 -6561
rect -456 -12639 -220 -6561
rect 6642 -12639 6878 -6561
rect 13740 -12639 13976 -6561
rect 20838 -12639 21074 -6561
rect -14652 -19039 -14416 -12961
rect -7554 -19039 -7318 -12961
rect -456 -19039 -220 -12961
rect 6642 -19039 6878 -12961
rect 13740 -19039 13976 -12961
rect 20838 -19039 21074 -12961
rect -14652 -25439 -14416 -19361
rect -7554 -25439 -7318 -19361
rect -456 -25439 -220 -19361
rect 6642 -25439 6878 -19361
rect 13740 -25439 13976 -19361
rect 20838 -25439 21074 -19361
rect -14652 -31839 -14416 -25761
rect -7554 -31839 -7318 -25761
rect -456 -31839 -220 -25761
rect 6642 -31839 6878 -25761
rect 13740 -31839 13976 -25761
rect 20838 -31839 21074 -25761
rect -14652 -38239 -14416 -32161
rect -7554 -38239 -7318 -32161
rect -456 -38239 -220 -32161
rect 6642 -38239 6878 -32161
rect 13740 -38239 13976 -32161
rect 20838 -38239 21074 -32161
<< mimcap2 >>
rect -21014 38160 -15014 38200
rect -21014 32240 -20974 38160
rect -15054 32240 -15014 38160
rect -21014 32200 -15014 32240
rect -13916 38160 -7916 38200
rect -13916 32240 -13876 38160
rect -7956 32240 -7916 38160
rect -13916 32200 -7916 32240
rect -6818 38160 -818 38200
rect -6818 32240 -6778 38160
rect -858 32240 -818 38160
rect -6818 32200 -818 32240
rect 280 38160 6280 38200
rect 280 32240 320 38160
rect 6240 32240 6280 38160
rect 280 32200 6280 32240
rect 7378 38160 13378 38200
rect 7378 32240 7418 38160
rect 13338 32240 13378 38160
rect 7378 32200 13378 32240
rect 14476 38160 20476 38200
rect 14476 32240 14516 38160
rect 20436 32240 20476 38160
rect 14476 32200 20476 32240
rect -21014 31760 -15014 31800
rect -21014 25840 -20974 31760
rect -15054 25840 -15014 31760
rect -21014 25800 -15014 25840
rect -13916 31760 -7916 31800
rect -13916 25840 -13876 31760
rect -7956 25840 -7916 31760
rect -13916 25800 -7916 25840
rect -6818 31760 -818 31800
rect -6818 25840 -6778 31760
rect -858 25840 -818 31760
rect -6818 25800 -818 25840
rect 280 31760 6280 31800
rect 280 25840 320 31760
rect 6240 25840 6280 31760
rect 280 25800 6280 25840
rect 7378 31760 13378 31800
rect 7378 25840 7418 31760
rect 13338 25840 13378 31760
rect 7378 25800 13378 25840
rect 14476 31760 20476 31800
rect 14476 25840 14516 31760
rect 20436 25840 20476 31760
rect 14476 25800 20476 25840
rect -21014 25360 -15014 25400
rect -21014 19440 -20974 25360
rect -15054 19440 -15014 25360
rect -21014 19400 -15014 19440
rect -13916 25360 -7916 25400
rect -13916 19440 -13876 25360
rect -7956 19440 -7916 25360
rect -13916 19400 -7916 19440
rect -6818 25360 -818 25400
rect -6818 19440 -6778 25360
rect -858 19440 -818 25360
rect -6818 19400 -818 19440
rect 280 25360 6280 25400
rect 280 19440 320 25360
rect 6240 19440 6280 25360
rect 280 19400 6280 19440
rect 7378 25360 13378 25400
rect 7378 19440 7418 25360
rect 13338 19440 13378 25360
rect 7378 19400 13378 19440
rect 14476 25360 20476 25400
rect 14476 19440 14516 25360
rect 20436 19440 20476 25360
rect 14476 19400 20476 19440
rect -21014 18960 -15014 19000
rect -21014 13040 -20974 18960
rect -15054 13040 -15014 18960
rect -21014 13000 -15014 13040
rect -13916 18960 -7916 19000
rect -13916 13040 -13876 18960
rect -7956 13040 -7916 18960
rect -13916 13000 -7916 13040
rect -6818 18960 -818 19000
rect -6818 13040 -6778 18960
rect -858 13040 -818 18960
rect -6818 13000 -818 13040
rect 280 18960 6280 19000
rect 280 13040 320 18960
rect 6240 13040 6280 18960
rect 280 13000 6280 13040
rect 7378 18960 13378 19000
rect 7378 13040 7418 18960
rect 13338 13040 13378 18960
rect 7378 13000 13378 13040
rect 14476 18960 20476 19000
rect 14476 13040 14516 18960
rect 20436 13040 20476 18960
rect 14476 13000 20476 13040
rect -21014 12560 -15014 12600
rect -21014 6640 -20974 12560
rect -15054 6640 -15014 12560
rect -21014 6600 -15014 6640
rect -13916 12560 -7916 12600
rect -13916 6640 -13876 12560
rect -7956 6640 -7916 12560
rect -13916 6600 -7916 6640
rect -6818 12560 -818 12600
rect -6818 6640 -6778 12560
rect -858 6640 -818 12560
rect -6818 6600 -818 6640
rect 280 12560 6280 12600
rect 280 6640 320 12560
rect 6240 6640 6280 12560
rect 280 6600 6280 6640
rect 7378 12560 13378 12600
rect 7378 6640 7418 12560
rect 13338 6640 13378 12560
rect 7378 6600 13378 6640
rect 14476 12560 20476 12600
rect 14476 6640 14516 12560
rect 20436 6640 20476 12560
rect 14476 6600 20476 6640
rect -21014 6160 -15014 6200
rect -21014 240 -20974 6160
rect -15054 240 -15014 6160
rect -21014 200 -15014 240
rect -13916 6160 -7916 6200
rect -13916 240 -13876 6160
rect -7956 240 -7916 6160
rect -13916 200 -7916 240
rect -6818 6160 -818 6200
rect -6818 240 -6778 6160
rect -858 240 -818 6160
rect -6818 200 -818 240
rect 280 6160 6280 6200
rect 280 240 320 6160
rect 6240 240 6280 6160
rect 280 200 6280 240
rect 7378 6160 13378 6200
rect 7378 240 7418 6160
rect 13338 240 13378 6160
rect 7378 200 13378 240
rect 14476 6160 20476 6200
rect 14476 240 14516 6160
rect 20436 240 20476 6160
rect 14476 200 20476 240
rect -21014 -240 -15014 -200
rect -21014 -6160 -20974 -240
rect -15054 -6160 -15014 -240
rect -21014 -6200 -15014 -6160
rect -13916 -240 -7916 -200
rect -13916 -6160 -13876 -240
rect -7956 -6160 -7916 -240
rect -13916 -6200 -7916 -6160
rect -6818 -240 -818 -200
rect -6818 -6160 -6778 -240
rect -858 -6160 -818 -240
rect -6818 -6200 -818 -6160
rect 280 -240 6280 -200
rect 280 -6160 320 -240
rect 6240 -6160 6280 -240
rect 280 -6200 6280 -6160
rect 7378 -240 13378 -200
rect 7378 -6160 7418 -240
rect 13338 -6160 13378 -240
rect 7378 -6200 13378 -6160
rect 14476 -240 20476 -200
rect 14476 -6160 14516 -240
rect 20436 -6160 20476 -240
rect 14476 -6200 20476 -6160
rect -21014 -6640 -15014 -6600
rect -21014 -12560 -20974 -6640
rect -15054 -12560 -15014 -6640
rect -21014 -12600 -15014 -12560
rect -13916 -6640 -7916 -6600
rect -13916 -12560 -13876 -6640
rect -7956 -12560 -7916 -6640
rect -13916 -12600 -7916 -12560
rect -6818 -6640 -818 -6600
rect -6818 -12560 -6778 -6640
rect -858 -12560 -818 -6640
rect -6818 -12600 -818 -12560
rect 280 -6640 6280 -6600
rect 280 -12560 320 -6640
rect 6240 -12560 6280 -6640
rect 280 -12600 6280 -12560
rect 7378 -6640 13378 -6600
rect 7378 -12560 7418 -6640
rect 13338 -12560 13378 -6640
rect 7378 -12600 13378 -12560
rect 14476 -6640 20476 -6600
rect 14476 -12560 14516 -6640
rect 20436 -12560 20476 -6640
rect 14476 -12600 20476 -12560
rect -21014 -13040 -15014 -13000
rect -21014 -18960 -20974 -13040
rect -15054 -18960 -15014 -13040
rect -21014 -19000 -15014 -18960
rect -13916 -13040 -7916 -13000
rect -13916 -18960 -13876 -13040
rect -7956 -18960 -7916 -13040
rect -13916 -19000 -7916 -18960
rect -6818 -13040 -818 -13000
rect -6818 -18960 -6778 -13040
rect -858 -18960 -818 -13040
rect -6818 -19000 -818 -18960
rect 280 -13040 6280 -13000
rect 280 -18960 320 -13040
rect 6240 -18960 6280 -13040
rect 280 -19000 6280 -18960
rect 7378 -13040 13378 -13000
rect 7378 -18960 7418 -13040
rect 13338 -18960 13378 -13040
rect 7378 -19000 13378 -18960
rect 14476 -13040 20476 -13000
rect 14476 -18960 14516 -13040
rect 20436 -18960 20476 -13040
rect 14476 -19000 20476 -18960
rect -21014 -19440 -15014 -19400
rect -21014 -25360 -20974 -19440
rect -15054 -25360 -15014 -19440
rect -21014 -25400 -15014 -25360
rect -13916 -19440 -7916 -19400
rect -13916 -25360 -13876 -19440
rect -7956 -25360 -7916 -19440
rect -13916 -25400 -7916 -25360
rect -6818 -19440 -818 -19400
rect -6818 -25360 -6778 -19440
rect -858 -25360 -818 -19440
rect -6818 -25400 -818 -25360
rect 280 -19440 6280 -19400
rect 280 -25360 320 -19440
rect 6240 -25360 6280 -19440
rect 280 -25400 6280 -25360
rect 7378 -19440 13378 -19400
rect 7378 -25360 7418 -19440
rect 13338 -25360 13378 -19440
rect 7378 -25400 13378 -25360
rect 14476 -19440 20476 -19400
rect 14476 -25360 14516 -19440
rect 20436 -25360 20476 -19440
rect 14476 -25400 20476 -25360
rect -21014 -25840 -15014 -25800
rect -21014 -31760 -20974 -25840
rect -15054 -31760 -15014 -25840
rect -21014 -31800 -15014 -31760
rect -13916 -25840 -7916 -25800
rect -13916 -31760 -13876 -25840
rect -7956 -31760 -7916 -25840
rect -13916 -31800 -7916 -31760
rect -6818 -25840 -818 -25800
rect -6818 -31760 -6778 -25840
rect -858 -31760 -818 -25840
rect -6818 -31800 -818 -31760
rect 280 -25840 6280 -25800
rect 280 -31760 320 -25840
rect 6240 -31760 6280 -25840
rect 280 -31800 6280 -31760
rect 7378 -25840 13378 -25800
rect 7378 -31760 7418 -25840
rect 13338 -31760 13378 -25840
rect 7378 -31800 13378 -31760
rect 14476 -25840 20476 -25800
rect 14476 -31760 14516 -25840
rect 20436 -31760 20476 -25840
rect 14476 -31800 20476 -31760
rect -21014 -32240 -15014 -32200
rect -21014 -38160 -20974 -32240
rect -15054 -38160 -15014 -32240
rect -21014 -38200 -15014 -38160
rect -13916 -32240 -7916 -32200
rect -13916 -38160 -13876 -32240
rect -7956 -38160 -7916 -32240
rect -13916 -38200 -7916 -38160
rect -6818 -32240 -818 -32200
rect -6818 -38160 -6778 -32240
rect -858 -38160 -818 -32240
rect -6818 -38200 -818 -38160
rect 280 -32240 6280 -32200
rect 280 -38160 320 -32240
rect 6240 -38160 6280 -32240
rect 280 -38200 6280 -38160
rect 7378 -32240 13378 -32200
rect 7378 -38160 7418 -32240
rect 13338 -38160 13378 -32240
rect 7378 -38200 13378 -38160
rect 14476 -32240 20476 -32200
rect 14476 -38160 14516 -32240
rect 20436 -38160 20476 -32240
rect 14476 -38200 20476 -38160
<< mimcap2contact >>
rect -20974 32240 -15054 38160
rect -13876 32240 -7956 38160
rect -6778 32240 -858 38160
rect 320 32240 6240 38160
rect 7418 32240 13338 38160
rect 14516 32240 20436 38160
rect -20974 25840 -15054 31760
rect -13876 25840 -7956 31760
rect -6778 25840 -858 31760
rect 320 25840 6240 31760
rect 7418 25840 13338 31760
rect 14516 25840 20436 31760
rect -20974 19440 -15054 25360
rect -13876 19440 -7956 25360
rect -6778 19440 -858 25360
rect 320 19440 6240 25360
rect 7418 19440 13338 25360
rect 14516 19440 20436 25360
rect -20974 13040 -15054 18960
rect -13876 13040 -7956 18960
rect -6778 13040 -858 18960
rect 320 13040 6240 18960
rect 7418 13040 13338 18960
rect 14516 13040 20436 18960
rect -20974 6640 -15054 12560
rect -13876 6640 -7956 12560
rect -6778 6640 -858 12560
rect 320 6640 6240 12560
rect 7418 6640 13338 12560
rect 14516 6640 20436 12560
rect -20974 240 -15054 6160
rect -13876 240 -7956 6160
rect -6778 240 -858 6160
rect 320 240 6240 6160
rect 7418 240 13338 6160
rect 14516 240 20436 6160
rect -20974 -6160 -15054 -240
rect -13876 -6160 -7956 -240
rect -6778 -6160 -858 -240
rect 320 -6160 6240 -240
rect 7418 -6160 13338 -240
rect 14516 -6160 20436 -240
rect -20974 -12560 -15054 -6640
rect -13876 -12560 -7956 -6640
rect -6778 -12560 -858 -6640
rect 320 -12560 6240 -6640
rect 7418 -12560 13338 -6640
rect 14516 -12560 20436 -6640
rect -20974 -18960 -15054 -13040
rect -13876 -18960 -7956 -13040
rect -6778 -18960 -858 -13040
rect 320 -18960 6240 -13040
rect 7418 -18960 13338 -13040
rect 14516 -18960 20436 -13040
rect -20974 -25360 -15054 -19440
rect -13876 -25360 -7956 -19440
rect -6778 -25360 -858 -19440
rect 320 -25360 6240 -19440
rect 7418 -25360 13338 -19440
rect 14516 -25360 20436 -19440
rect -20974 -31760 -15054 -25840
rect -13876 -31760 -7956 -25840
rect -6778 -31760 -858 -25840
rect 320 -31760 6240 -25840
rect 7418 -31760 13338 -25840
rect 14516 -31760 20436 -25840
rect -20974 -38160 -15054 -32240
rect -13876 -38160 -7956 -32240
rect -6778 -38160 -858 -32240
rect 320 -38160 6240 -32240
rect 7418 -38160 13338 -32240
rect 14516 -38160 20436 -32240
<< metal5 >>
rect -18174 38184 -17854 38400
rect -14694 38239 -14374 38400
rect -20998 38160 -15030 38184
rect -20998 32240 -20974 38160
rect -15054 32240 -15030 38160
rect -20998 32216 -15030 32240
rect -18174 31784 -17854 32216
rect -14694 32161 -14652 38239
rect -14416 32161 -14374 38239
rect -11076 38184 -10756 38400
rect -7596 38239 -7276 38400
rect -13900 38160 -7932 38184
rect -13900 32240 -13876 38160
rect -7956 32240 -7932 38160
rect -13900 32216 -7932 32240
rect -14694 31839 -14374 32161
rect -20998 31760 -15030 31784
rect -20998 25840 -20974 31760
rect -15054 25840 -15030 31760
rect -20998 25816 -15030 25840
rect -18174 25384 -17854 25816
rect -14694 25761 -14652 31839
rect -14416 25761 -14374 31839
rect -11076 31784 -10756 32216
rect -7596 32161 -7554 38239
rect -7318 32161 -7276 38239
rect -3978 38184 -3658 38400
rect -498 38239 -178 38400
rect -6802 38160 -834 38184
rect -6802 32240 -6778 38160
rect -858 32240 -834 38160
rect -6802 32216 -834 32240
rect -7596 31839 -7276 32161
rect -13900 31760 -7932 31784
rect -13900 25840 -13876 31760
rect -7956 25840 -7932 31760
rect -13900 25816 -7932 25840
rect -14694 25439 -14374 25761
rect -20998 25360 -15030 25384
rect -20998 19440 -20974 25360
rect -15054 19440 -15030 25360
rect -20998 19416 -15030 19440
rect -18174 18984 -17854 19416
rect -14694 19361 -14652 25439
rect -14416 19361 -14374 25439
rect -11076 25384 -10756 25816
rect -7596 25761 -7554 31839
rect -7318 25761 -7276 31839
rect -3978 31784 -3658 32216
rect -498 32161 -456 38239
rect -220 32161 -178 38239
rect 3120 38184 3440 38400
rect 6600 38239 6920 38400
rect 296 38160 6264 38184
rect 296 32240 320 38160
rect 6240 32240 6264 38160
rect 296 32216 6264 32240
rect -498 31839 -178 32161
rect -6802 31760 -834 31784
rect -6802 25840 -6778 31760
rect -858 25840 -834 31760
rect -6802 25816 -834 25840
rect -7596 25439 -7276 25761
rect -13900 25360 -7932 25384
rect -13900 19440 -13876 25360
rect -7956 19440 -7932 25360
rect -13900 19416 -7932 19440
rect -14694 19039 -14374 19361
rect -20998 18960 -15030 18984
rect -20998 13040 -20974 18960
rect -15054 13040 -15030 18960
rect -20998 13016 -15030 13040
rect -18174 12584 -17854 13016
rect -14694 12961 -14652 19039
rect -14416 12961 -14374 19039
rect -11076 18984 -10756 19416
rect -7596 19361 -7554 25439
rect -7318 19361 -7276 25439
rect -3978 25384 -3658 25816
rect -498 25761 -456 31839
rect -220 25761 -178 31839
rect 3120 31784 3440 32216
rect 6600 32161 6642 38239
rect 6878 32161 6920 38239
rect 10218 38184 10538 38400
rect 13698 38239 14018 38400
rect 7394 38160 13362 38184
rect 7394 32240 7418 38160
rect 13338 32240 13362 38160
rect 7394 32216 13362 32240
rect 6600 31839 6920 32161
rect 296 31760 6264 31784
rect 296 25840 320 31760
rect 6240 25840 6264 31760
rect 296 25816 6264 25840
rect -498 25439 -178 25761
rect -6802 25360 -834 25384
rect -6802 19440 -6778 25360
rect -858 19440 -834 25360
rect -6802 19416 -834 19440
rect -7596 19039 -7276 19361
rect -13900 18960 -7932 18984
rect -13900 13040 -13876 18960
rect -7956 13040 -7932 18960
rect -13900 13016 -7932 13040
rect -14694 12639 -14374 12961
rect -20998 12560 -15030 12584
rect -20998 6640 -20974 12560
rect -15054 6640 -15030 12560
rect -20998 6616 -15030 6640
rect -18174 6184 -17854 6616
rect -14694 6561 -14652 12639
rect -14416 6561 -14374 12639
rect -11076 12584 -10756 13016
rect -7596 12961 -7554 19039
rect -7318 12961 -7276 19039
rect -3978 18984 -3658 19416
rect -498 19361 -456 25439
rect -220 19361 -178 25439
rect 3120 25384 3440 25816
rect 6600 25761 6642 31839
rect 6878 25761 6920 31839
rect 10218 31784 10538 32216
rect 13698 32161 13740 38239
rect 13976 32161 14018 38239
rect 17316 38184 17636 38400
rect 20796 38239 21116 38400
rect 14492 38160 20460 38184
rect 14492 32240 14516 38160
rect 20436 32240 20460 38160
rect 14492 32216 20460 32240
rect 13698 31839 14018 32161
rect 7394 31760 13362 31784
rect 7394 25840 7418 31760
rect 13338 25840 13362 31760
rect 7394 25816 13362 25840
rect 6600 25439 6920 25761
rect 296 25360 6264 25384
rect 296 19440 320 25360
rect 6240 19440 6264 25360
rect 296 19416 6264 19440
rect -498 19039 -178 19361
rect -6802 18960 -834 18984
rect -6802 13040 -6778 18960
rect -858 13040 -834 18960
rect -6802 13016 -834 13040
rect -7596 12639 -7276 12961
rect -13900 12560 -7932 12584
rect -13900 6640 -13876 12560
rect -7956 6640 -7932 12560
rect -13900 6616 -7932 6640
rect -14694 6239 -14374 6561
rect -20998 6160 -15030 6184
rect -20998 240 -20974 6160
rect -15054 240 -15030 6160
rect -20998 216 -15030 240
rect -18174 -216 -17854 216
rect -14694 161 -14652 6239
rect -14416 161 -14374 6239
rect -11076 6184 -10756 6616
rect -7596 6561 -7554 12639
rect -7318 6561 -7276 12639
rect -3978 12584 -3658 13016
rect -498 12961 -456 19039
rect -220 12961 -178 19039
rect 3120 18984 3440 19416
rect 6600 19361 6642 25439
rect 6878 19361 6920 25439
rect 10218 25384 10538 25816
rect 13698 25761 13740 31839
rect 13976 25761 14018 31839
rect 17316 31784 17636 32216
rect 20796 32161 20838 38239
rect 21074 32161 21116 38239
rect 20796 31839 21116 32161
rect 14492 31760 20460 31784
rect 14492 25840 14516 31760
rect 20436 25840 20460 31760
rect 14492 25816 20460 25840
rect 13698 25439 14018 25761
rect 7394 25360 13362 25384
rect 7394 19440 7418 25360
rect 13338 19440 13362 25360
rect 7394 19416 13362 19440
rect 6600 19039 6920 19361
rect 296 18960 6264 18984
rect 296 13040 320 18960
rect 6240 13040 6264 18960
rect 296 13016 6264 13040
rect -498 12639 -178 12961
rect -6802 12560 -834 12584
rect -6802 6640 -6778 12560
rect -858 6640 -834 12560
rect -6802 6616 -834 6640
rect -7596 6239 -7276 6561
rect -13900 6160 -7932 6184
rect -13900 240 -13876 6160
rect -7956 240 -7932 6160
rect -13900 216 -7932 240
rect -14694 -161 -14374 161
rect -20998 -240 -15030 -216
rect -20998 -6160 -20974 -240
rect -15054 -6160 -15030 -240
rect -20998 -6184 -15030 -6160
rect -18174 -6616 -17854 -6184
rect -14694 -6239 -14652 -161
rect -14416 -6239 -14374 -161
rect -11076 -216 -10756 216
rect -7596 161 -7554 6239
rect -7318 161 -7276 6239
rect -3978 6184 -3658 6616
rect -498 6561 -456 12639
rect -220 6561 -178 12639
rect 3120 12584 3440 13016
rect 6600 12961 6642 19039
rect 6878 12961 6920 19039
rect 10218 18984 10538 19416
rect 13698 19361 13740 25439
rect 13976 19361 14018 25439
rect 17316 25384 17636 25816
rect 20796 25761 20838 31839
rect 21074 25761 21116 31839
rect 20796 25439 21116 25761
rect 14492 25360 20460 25384
rect 14492 19440 14516 25360
rect 20436 19440 20460 25360
rect 14492 19416 20460 19440
rect 13698 19039 14018 19361
rect 7394 18960 13362 18984
rect 7394 13040 7418 18960
rect 13338 13040 13362 18960
rect 7394 13016 13362 13040
rect 6600 12639 6920 12961
rect 296 12560 6264 12584
rect 296 6640 320 12560
rect 6240 6640 6264 12560
rect 296 6616 6264 6640
rect -498 6239 -178 6561
rect -6802 6160 -834 6184
rect -6802 240 -6778 6160
rect -858 240 -834 6160
rect -6802 216 -834 240
rect -7596 -161 -7276 161
rect -13900 -240 -7932 -216
rect -13900 -6160 -13876 -240
rect -7956 -6160 -7932 -240
rect -13900 -6184 -7932 -6160
rect -14694 -6561 -14374 -6239
rect -20998 -6640 -15030 -6616
rect -20998 -12560 -20974 -6640
rect -15054 -12560 -15030 -6640
rect -20998 -12584 -15030 -12560
rect -18174 -13016 -17854 -12584
rect -14694 -12639 -14652 -6561
rect -14416 -12639 -14374 -6561
rect -11076 -6616 -10756 -6184
rect -7596 -6239 -7554 -161
rect -7318 -6239 -7276 -161
rect -3978 -216 -3658 216
rect -498 161 -456 6239
rect -220 161 -178 6239
rect 3120 6184 3440 6616
rect 6600 6561 6642 12639
rect 6878 6561 6920 12639
rect 10218 12584 10538 13016
rect 13698 12961 13740 19039
rect 13976 12961 14018 19039
rect 17316 18984 17636 19416
rect 20796 19361 20838 25439
rect 21074 19361 21116 25439
rect 20796 19039 21116 19361
rect 14492 18960 20460 18984
rect 14492 13040 14516 18960
rect 20436 13040 20460 18960
rect 14492 13016 20460 13040
rect 13698 12639 14018 12961
rect 7394 12560 13362 12584
rect 7394 6640 7418 12560
rect 13338 6640 13362 12560
rect 7394 6616 13362 6640
rect 6600 6239 6920 6561
rect 296 6160 6264 6184
rect 296 240 320 6160
rect 6240 240 6264 6160
rect 296 216 6264 240
rect -498 -161 -178 161
rect -6802 -240 -834 -216
rect -6802 -6160 -6778 -240
rect -858 -6160 -834 -240
rect -6802 -6184 -834 -6160
rect -7596 -6561 -7276 -6239
rect -13900 -6640 -7932 -6616
rect -13900 -12560 -13876 -6640
rect -7956 -12560 -7932 -6640
rect -13900 -12584 -7932 -12560
rect -14694 -12961 -14374 -12639
rect -20998 -13040 -15030 -13016
rect -20998 -18960 -20974 -13040
rect -15054 -18960 -15030 -13040
rect -20998 -18984 -15030 -18960
rect -18174 -19416 -17854 -18984
rect -14694 -19039 -14652 -12961
rect -14416 -19039 -14374 -12961
rect -11076 -13016 -10756 -12584
rect -7596 -12639 -7554 -6561
rect -7318 -12639 -7276 -6561
rect -3978 -6616 -3658 -6184
rect -498 -6239 -456 -161
rect -220 -6239 -178 -161
rect 3120 -216 3440 216
rect 6600 161 6642 6239
rect 6878 161 6920 6239
rect 10218 6184 10538 6616
rect 13698 6561 13740 12639
rect 13976 6561 14018 12639
rect 17316 12584 17636 13016
rect 20796 12961 20838 19039
rect 21074 12961 21116 19039
rect 20796 12639 21116 12961
rect 14492 12560 20460 12584
rect 14492 6640 14516 12560
rect 20436 6640 20460 12560
rect 14492 6616 20460 6640
rect 13698 6239 14018 6561
rect 7394 6160 13362 6184
rect 7394 240 7418 6160
rect 13338 240 13362 6160
rect 7394 216 13362 240
rect 6600 -161 6920 161
rect 296 -240 6264 -216
rect 296 -6160 320 -240
rect 6240 -6160 6264 -240
rect 296 -6184 6264 -6160
rect -498 -6561 -178 -6239
rect -6802 -6640 -834 -6616
rect -6802 -12560 -6778 -6640
rect -858 -12560 -834 -6640
rect -6802 -12584 -834 -12560
rect -7596 -12961 -7276 -12639
rect -13900 -13040 -7932 -13016
rect -13900 -18960 -13876 -13040
rect -7956 -18960 -7932 -13040
rect -13900 -18984 -7932 -18960
rect -14694 -19361 -14374 -19039
rect -20998 -19440 -15030 -19416
rect -20998 -25360 -20974 -19440
rect -15054 -25360 -15030 -19440
rect -20998 -25384 -15030 -25360
rect -18174 -25816 -17854 -25384
rect -14694 -25439 -14652 -19361
rect -14416 -25439 -14374 -19361
rect -11076 -19416 -10756 -18984
rect -7596 -19039 -7554 -12961
rect -7318 -19039 -7276 -12961
rect -3978 -13016 -3658 -12584
rect -498 -12639 -456 -6561
rect -220 -12639 -178 -6561
rect 3120 -6616 3440 -6184
rect 6600 -6239 6642 -161
rect 6878 -6239 6920 -161
rect 10218 -216 10538 216
rect 13698 161 13740 6239
rect 13976 161 14018 6239
rect 17316 6184 17636 6616
rect 20796 6561 20838 12639
rect 21074 6561 21116 12639
rect 20796 6239 21116 6561
rect 14492 6160 20460 6184
rect 14492 240 14516 6160
rect 20436 240 20460 6160
rect 14492 216 20460 240
rect 13698 -161 14018 161
rect 7394 -240 13362 -216
rect 7394 -6160 7418 -240
rect 13338 -6160 13362 -240
rect 7394 -6184 13362 -6160
rect 6600 -6561 6920 -6239
rect 296 -6640 6264 -6616
rect 296 -12560 320 -6640
rect 6240 -12560 6264 -6640
rect 296 -12584 6264 -12560
rect -498 -12961 -178 -12639
rect -6802 -13040 -834 -13016
rect -6802 -18960 -6778 -13040
rect -858 -18960 -834 -13040
rect -6802 -18984 -834 -18960
rect -7596 -19361 -7276 -19039
rect -13900 -19440 -7932 -19416
rect -13900 -25360 -13876 -19440
rect -7956 -25360 -7932 -19440
rect -13900 -25384 -7932 -25360
rect -14694 -25761 -14374 -25439
rect -20998 -25840 -15030 -25816
rect -20998 -31760 -20974 -25840
rect -15054 -31760 -15030 -25840
rect -20998 -31784 -15030 -31760
rect -18174 -32216 -17854 -31784
rect -14694 -31839 -14652 -25761
rect -14416 -31839 -14374 -25761
rect -11076 -25816 -10756 -25384
rect -7596 -25439 -7554 -19361
rect -7318 -25439 -7276 -19361
rect -3978 -19416 -3658 -18984
rect -498 -19039 -456 -12961
rect -220 -19039 -178 -12961
rect 3120 -13016 3440 -12584
rect 6600 -12639 6642 -6561
rect 6878 -12639 6920 -6561
rect 10218 -6616 10538 -6184
rect 13698 -6239 13740 -161
rect 13976 -6239 14018 -161
rect 17316 -216 17636 216
rect 20796 161 20838 6239
rect 21074 161 21116 6239
rect 20796 -161 21116 161
rect 14492 -240 20460 -216
rect 14492 -6160 14516 -240
rect 20436 -6160 20460 -240
rect 14492 -6184 20460 -6160
rect 13698 -6561 14018 -6239
rect 7394 -6640 13362 -6616
rect 7394 -12560 7418 -6640
rect 13338 -12560 13362 -6640
rect 7394 -12584 13362 -12560
rect 6600 -12961 6920 -12639
rect 296 -13040 6264 -13016
rect 296 -18960 320 -13040
rect 6240 -18960 6264 -13040
rect 296 -18984 6264 -18960
rect -498 -19361 -178 -19039
rect -6802 -19440 -834 -19416
rect -6802 -25360 -6778 -19440
rect -858 -25360 -834 -19440
rect -6802 -25384 -834 -25360
rect -7596 -25761 -7276 -25439
rect -13900 -25840 -7932 -25816
rect -13900 -31760 -13876 -25840
rect -7956 -31760 -7932 -25840
rect -13900 -31784 -7932 -31760
rect -14694 -32161 -14374 -31839
rect -20998 -32240 -15030 -32216
rect -20998 -38160 -20974 -32240
rect -15054 -38160 -15030 -32240
rect -20998 -38184 -15030 -38160
rect -18174 -38400 -17854 -38184
rect -14694 -38239 -14652 -32161
rect -14416 -38239 -14374 -32161
rect -11076 -32216 -10756 -31784
rect -7596 -31839 -7554 -25761
rect -7318 -31839 -7276 -25761
rect -3978 -25816 -3658 -25384
rect -498 -25439 -456 -19361
rect -220 -25439 -178 -19361
rect 3120 -19416 3440 -18984
rect 6600 -19039 6642 -12961
rect 6878 -19039 6920 -12961
rect 10218 -13016 10538 -12584
rect 13698 -12639 13740 -6561
rect 13976 -12639 14018 -6561
rect 17316 -6616 17636 -6184
rect 20796 -6239 20838 -161
rect 21074 -6239 21116 -161
rect 20796 -6561 21116 -6239
rect 14492 -6640 20460 -6616
rect 14492 -12560 14516 -6640
rect 20436 -12560 20460 -6640
rect 14492 -12584 20460 -12560
rect 13698 -12961 14018 -12639
rect 7394 -13040 13362 -13016
rect 7394 -18960 7418 -13040
rect 13338 -18960 13362 -13040
rect 7394 -18984 13362 -18960
rect 6600 -19361 6920 -19039
rect 296 -19440 6264 -19416
rect 296 -25360 320 -19440
rect 6240 -25360 6264 -19440
rect 296 -25384 6264 -25360
rect -498 -25761 -178 -25439
rect -6802 -25840 -834 -25816
rect -6802 -31760 -6778 -25840
rect -858 -31760 -834 -25840
rect -6802 -31784 -834 -31760
rect -7596 -32161 -7276 -31839
rect -13900 -32240 -7932 -32216
rect -13900 -38160 -13876 -32240
rect -7956 -38160 -7932 -32240
rect -13900 -38184 -7932 -38160
rect -14694 -38400 -14374 -38239
rect -11076 -38400 -10756 -38184
rect -7596 -38239 -7554 -32161
rect -7318 -38239 -7276 -32161
rect -3978 -32216 -3658 -31784
rect -498 -31839 -456 -25761
rect -220 -31839 -178 -25761
rect 3120 -25816 3440 -25384
rect 6600 -25439 6642 -19361
rect 6878 -25439 6920 -19361
rect 10218 -19416 10538 -18984
rect 13698 -19039 13740 -12961
rect 13976 -19039 14018 -12961
rect 17316 -13016 17636 -12584
rect 20796 -12639 20838 -6561
rect 21074 -12639 21116 -6561
rect 20796 -12961 21116 -12639
rect 14492 -13040 20460 -13016
rect 14492 -18960 14516 -13040
rect 20436 -18960 20460 -13040
rect 14492 -18984 20460 -18960
rect 13698 -19361 14018 -19039
rect 7394 -19440 13362 -19416
rect 7394 -25360 7418 -19440
rect 13338 -25360 13362 -19440
rect 7394 -25384 13362 -25360
rect 6600 -25761 6920 -25439
rect 296 -25840 6264 -25816
rect 296 -31760 320 -25840
rect 6240 -31760 6264 -25840
rect 296 -31784 6264 -31760
rect -498 -32161 -178 -31839
rect -6802 -32240 -834 -32216
rect -6802 -38160 -6778 -32240
rect -858 -38160 -834 -32240
rect -6802 -38184 -834 -38160
rect -7596 -38400 -7276 -38239
rect -3978 -38400 -3658 -38184
rect -498 -38239 -456 -32161
rect -220 -38239 -178 -32161
rect 3120 -32216 3440 -31784
rect 6600 -31839 6642 -25761
rect 6878 -31839 6920 -25761
rect 10218 -25816 10538 -25384
rect 13698 -25439 13740 -19361
rect 13976 -25439 14018 -19361
rect 17316 -19416 17636 -18984
rect 20796 -19039 20838 -12961
rect 21074 -19039 21116 -12961
rect 20796 -19361 21116 -19039
rect 14492 -19440 20460 -19416
rect 14492 -25360 14516 -19440
rect 20436 -25360 20460 -19440
rect 14492 -25384 20460 -25360
rect 13698 -25761 14018 -25439
rect 7394 -25840 13362 -25816
rect 7394 -31760 7418 -25840
rect 13338 -31760 13362 -25840
rect 7394 -31784 13362 -31760
rect 6600 -32161 6920 -31839
rect 296 -32240 6264 -32216
rect 296 -38160 320 -32240
rect 6240 -38160 6264 -32240
rect 296 -38184 6264 -38160
rect -498 -38400 -178 -38239
rect 3120 -38400 3440 -38184
rect 6600 -38239 6642 -32161
rect 6878 -38239 6920 -32161
rect 10218 -32216 10538 -31784
rect 13698 -31839 13740 -25761
rect 13976 -31839 14018 -25761
rect 17316 -25816 17636 -25384
rect 20796 -25439 20838 -19361
rect 21074 -25439 21116 -19361
rect 20796 -25761 21116 -25439
rect 14492 -25840 20460 -25816
rect 14492 -31760 14516 -25840
rect 20436 -31760 20460 -25840
rect 14492 -31784 20460 -31760
rect 13698 -32161 14018 -31839
rect 7394 -32240 13362 -32216
rect 7394 -38160 7418 -32240
rect 13338 -38160 13362 -32240
rect 7394 -38184 13362 -38160
rect 6600 -38400 6920 -38239
rect 10218 -38400 10538 -38184
rect 13698 -38239 13740 -32161
rect 13976 -38239 14018 -32161
rect 17316 -32216 17636 -31784
rect 20796 -31839 20838 -25761
rect 21074 -31839 21116 -25761
rect 20796 -32161 21116 -31839
rect 14492 -32240 20460 -32216
rect 14492 -38160 14516 -32240
rect 20436 -38160 20460 -32240
rect 14492 -38184 20460 -38160
rect 13698 -38400 14018 -38239
rect 17316 -38400 17636 -38184
rect 20796 -38239 20838 -32161
rect 21074 -38239 21116 -32161
rect 20796 -38400 21116 -38239
<< properties >>
string FIXED_BBOX 14396 32120 20556 38280
string gencell sky130_fd_pr__cap_mim_m3_2
string library sky130
string parameters w 30 l 30 val 1.822k carea 2.00 cperi 0.19 nx 6 ny 12 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
