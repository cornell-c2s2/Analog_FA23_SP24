magic
tech sky130A
magscale 1 2
timestamp 1713027243
<< error_p >>
rect 6403 686267 6408 686273
rect 6409 686261 6415 686266
<< error_s >>
rect 6409 687586 6415 687591
rect 6403 687579 6408 687585
rect 57858 684084 57864 684090
rect 58852 684084 58858 684090
rect 57852 684078 57858 684084
rect 58858 684078 58864 684084
<< metal1 >>
rect 16988 698810 17948 698830
rect 16988 698690 17008 698810
rect 17128 698690 17208 698810
rect 17328 698690 17408 698810
rect 17528 698690 17608 698810
rect 17728 698690 17808 698810
rect 17928 698690 17948 698810
rect 16988 698670 17948 698690
rect 61024 694920 61924 694960
rect 61024 694740 61044 694920
rect 61224 694740 61384 694920
rect 61564 694740 61724 694920
rect 61904 694740 61924 694920
rect 61024 694700 61924 694740
rect 47100 690276 47400 690400
rect 47100 690224 47224 690276
rect 47276 690224 47400 690276
rect 47100 690010 47400 690224
rect 43870 689830 43950 690010
rect 45350 689990 47400 690010
rect 45350 689938 47224 689990
rect 47276 689938 47400 689990
rect 45350 689926 47400 689938
rect 45350 689874 47224 689926
rect 47276 689874 47400 689926
rect 45350 689862 47400 689874
rect 45350 689830 47224 689862
rect 47100 689810 47224 689830
rect 47276 689810 47400 689862
rect 18048 689650 18208 689690
rect 18048 689530 18068 689650
rect 18188 689530 18208 689650
rect 18048 689470 18208 689530
rect 18048 689350 18068 689470
rect 18188 689350 18208 689470
rect 47100 689576 47400 689810
rect 47100 689524 47224 689576
rect 47276 689524 47400 689576
rect 47100 689400 47400 689524
rect 18048 689290 18208 689350
rect 18048 689170 18068 689290
rect 18188 689170 18208 689290
rect 18048 689110 18208 689170
rect 18048 688990 18068 689110
rect 18188 688990 18208 689110
rect 18048 688930 18208 688990
rect 18048 688810 18068 688930
rect 18188 688810 18208 688930
rect 41900 688676 42200 688800
rect 41900 688624 42024 688676
rect 42076 688624 42200 688676
rect 6408 688530 7728 688610
rect 6408 688330 6508 688530
rect 6708 688330 6808 688530
rect 7008 688330 7108 688530
rect 7308 688330 7408 688530
rect 7608 688330 7728 688530
rect 6408 688230 7728 688330
rect 41900 688490 42200 688624
rect 41900 688438 42024 688490
rect 42076 688438 43870 688490
rect 41900 688426 43870 688438
rect 41900 688374 42024 688426
rect 42076 688374 43870 688426
rect 41900 688362 43870 688374
rect 41900 688310 42024 688362
rect 42076 688310 43870 688362
rect 41900 688176 42200 688310
rect 41900 688124 42024 688176
rect 42076 688124 42200 688176
rect 41900 688000 42200 688124
rect 60664 685660 60864 685700
rect 60664 685520 60704 685660
rect 60844 685520 60864 685660
rect 60664 685460 60864 685520
rect 60664 685320 60704 685460
rect 60844 685320 60864 685460
rect 60664 685280 60864 685320
rect 62024 685660 62224 685700
rect 62024 685520 62044 685660
rect 62184 685520 62224 685660
rect 62024 685460 62224 685520
rect 62024 685320 62044 685460
rect 62184 685320 62224 685460
rect 62024 685280 62224 685320
rect 71064 685660 71264 685700
rect 71064 685520 71104 685660
rect 71244 685520 71264 685660
rect 71064 685460 71264 685520
rect 71064 685320 71104 685460
rect 71244 685320 71264 685460
rect 71064 685280 71264 685320
rect 71204 684480 72484 684640
rect 40920 662800 48300 663400
<< via1 >>
rect 17008 698690 17128 698810
rect 17208 698690 17328 698810
rect 17408 698690 17528 698810
rect 17608 698690 17728 698810
rect 17808 698690 17928 698810
rect 61044 694740 61224 694920
rect 61384 694740 61564 694920
rect 61724 694740 61904 694920
rect 47224 690224 47276 690276
rect 47224 689938 47276 689990
rect 47224 689874 47276 689926
rect 47224 689810 47276 689862
rect 18068 689530 18188 689650
rect 18068 689350 18188 689470
rect 47224 689524 47276 689576
rect 18068 689170 18188 689290
rect 18068 688990 18188 689110
rect 18068 688810 18188 688930
rect 42024 688624 42076 688676
rect 6508 688330 6708 688530
rect 6808 688330 7008 688530
rect 7108 688330 7308 688530
rect 7408 688330 7608 688530
rect 42024 688438 42076 688490
rect 42024 688374 42076 688426
rect 42024 688310 42076 688362
rect 42024 688124 42076 688176
rect 60704 685520 60844 685660
rect 60704 685320 60844 685460
rect 62044 685520 62184 685660
rect 62044 685320 62184 685460
rect 71104 685520 71244 685660
rect 71104 685320 71244 685460
<< metal2 >>
rect 17008 698810 17128 698820
rect 17008 698680 17128 698690
rect 17208 698810 17328 698820
rect 17208 698680 17328 698690
rect 17408 698810 17528 698820
rect 17408 698680 17528 698690
rect 17608 698810 17728 698820
rect 17608 698680 17728 698690
rect 17808 698810 17928 698820
rect 17808 698680 17928 698690
rect 61044 694920 61224 694930
rect 61044 694730 61224 694740
rect 61384 694920 61564 694930
rect 61384 694730 61564 694740
rect 61724 694920 61904 694930
rect 61724 694730 61904 694740
rect 47200 690278 47300 690310
rect 47200 690222 47222 690278
rect 47278 690222 47300 690278
rect 47200 690190 47300 690222
rect 47200 689990 47300 690010
rect 47200 689968 47224 689990
rect 47276 689968 47300 689990
rect 47200 689912 47222 689968
rect 47278 689912 47300 689968
rect 47200 689888 47224 689912
rect 47276 689888 47300 689912
rect 47200 689832 47222 689888
rect 47278 689832 47300 689888
rect 47200 689810 47224 689832
rect 47276 689810 47300 689832
rect 47200 689790 47300 689810
rect 18068 689650 18188 689660
rect 18068 689520 18188 689530
rect 47200 689578 47300 689610
rect 47200 689522 47222 689578
rect 47278 689522 47300 689578
rect 47200 689490 47300 689522
rect 18068 689470 18188 689480
rect 18068 689340 18188 689350
rect 18068 689290 18188 689300
rect 18068 689160 18188 689170
rect 18068 689110 18188 689120
rect 18068 688980 18188 688990
rect 18068 688930 18188 688940
rect 18068 688800 18188 688810
rect 42000 688678 42100 688710
rect 42000 688622 42022 688678
rect 42078 688622 42100 688678
rect 42000 688590 42100 688622
rect 6508 688530 6708 688540
rect 6508 688320 6708 688330
rect 6808 688530 7008 688540
rect 6808 688320 7008 688330
rect 7108 688530 7308 688540
rect 7108 688320 7308 688330
rect 7408 688530 7608 688540
rect 7408 688320 7608 688330
rect 42000 688490 42100 688510
rect 42000 688468 42024 688490
rect 42076 688468 42100 688490
rect 42000 688412 42022 688468
rect 42078 688412 42100 688468
rect 42000 688388 42024 688412
rect 42076 688388 42100 688412
rect 42000 688332 42022 688388
rect 42078 688332 42100 688388
rect 42000 688310 42024 688332
rect 42076 688310 42100 688332
rect 42000 688290 42100 688310
rect 42000 688178 42100 688210
rect 42000 688122 42022 688178
rect 42078 688122 42100 688178
rect 42000 688090 42100 688122
rect 60704 685660 60844 685670
rect 60704 685510 60844 685520
rect 62044 685660 62184 685670
rect 62044 685510 62184 685520
rect 71104 685660 71244 685670
rect 71104 685510 71244 685520
rect 60704 685460 60844 685470
rect 60704 685310 60844 685320
rect 62044 685460 62184 685470
rect 62044 685310 62184 685320
rect 71104 685460 71244 685470
rect 71104 685310 71244 685320
rect 42240 683108 42640 684610
rect 42240 683052 42272 683108
rect 42328 683052 42412 683108
rect 42468 683052 42552 683108
rect 42608 683052 42640 683108
rect 42240 683020 42640 683052
rect 46640 683108 47040 684610
rect 46640 683052 46672 683108
rect 46728 683052 46812 683108
rect 46868 683052 46952 683108
rect 47008 683052 47040 683108
rect 46640 683020 47040 683052
<< via2 >>
rect 17008 698690 17128 698810
rect 17208 698690 17328 698810
rect 17408 698690 17528 698810
rect 17608 698690 17728 698810
rect 17808 698690 17928 698810
rect 61044 694740 61224 694920
rect 61384 694740 61564 694920
rect 61724 694740 61904 694920
rect 47222 690276 47278 690278
rect 47222 690224 47224 690276
rect 47224 690224 47276 690276
rect 47276 690224 47278 690276
rect 47222 690222 47278 690224
rect 47222 689938 47224 689968
rect 47224 689938 47276 689968
rect 47276 689938 47278 689968
rect 47222 689926 47278 689938
rect 47222 689912 47224 689926
rect 47224 689912 47276 689926
rect 47276 689912 47278 689926
rect 47222 689874 47224 689888
rect 47224 689874 47276 689888
rect 47276 689874 47278 689888
rect 47222 689862 47278 689874
rect 47222 689832 47224 689862
rect 47224 689832 47276 689862
rect 47276 689832 47278 689862
rect 18068 689530 18188 689650
rect 47222 689576 47278 689578
rect 47222 689524 47224 689576
rect 47224 689524 47276 689576
rect 47276 689524 47278 689576
rect 47222 689522 47278 689524
rect 18068 689350 18188 689470
rect 18068 689170 18188 689290
rect 18068 688990 18188 689110
rect 18068 688810 18188 688930
rect 42022 688676 42078 688678
rect 42022 688624 42024 688676
rect 42024 688624 42076 688676
rect 42076 688624 42078 688676
rect 42022 688622 42078 688624
rect 6508 688330 6708 688530
rect 6808 688330 7008 688530
rect 7108 688330 7308 688530
rect 7408 688330 7608 688530
rect 42022 688438 42024 688468
rect 42024 688438 42076 688468
rect 42076 688438 42078 688468
rect 42022 688426 42078 688438
rect 42022 688412 42024 688426
rect 42024 688412 42076 688426
rect 42076 688412 42078 688426
rect 42022 688374 42024 688388
rect 42024 688374 42076 688388
rect 42076 688374 42078 688388
rect 42022 688362 42078 688374
rect 42022 688332 42024 688362
rect 42024 688332 42076 688362
rect 42076 688332 42078 688362
rect 42022 688176 42078 688178
rect 42022 688124 42024 688176
rect 42024 688124 42076 688176
rect 42076 688124 42078 688176
rect 42022 688122 42078 688124
rect 60704 685520 60844 685660
rect 62044 685520 62184 685660
rect 71104 685520 71244 685660
rect 60704 685320 60844 685460
rect 62044 685320 62184 685460
rect 71104 685320 71244 685460
rect 42272 683052 42328 683108
rect 42412 683052 42468 683108
rect 42552 683052 42608 683108
rect 46672 683052 46728 683108
rect 46812 683052 46868 683108
rect 46952 683052 47008 683108
<< metal3 >>
rect 16998 698810 17138 698815
rect 16998 698690 17008 698810
rect 17128 698690 17138 698810
rect 16998 698685 17138 698690
rect 17198 698810 17338 698815
rect 17198 698690 17208 698810
rect 17328 698690 17338 698810
rect 17198 698685 17338 698690
rect 17398 698810 17538 698815
rect 17398 698690 17408 698810
rect 17528 698690 17538 698810
rect 17398 698685 17538 698690
rect 17598 698810 17738 698815
rect 17598 698690 17608 698810
rect 17728 698690 17738 698810
rect 17598 698685 17738 698690
rect 17798 698810 17938 698815
rect 17798 698690 17808 698810
rect 17928 698690 17938 698810
rect 17798 698685 17938 698690
rect 61034 694920 61234 694925
rect 6598 694630 6608 694830
rect 6808 694630 6818 694830
rect 7198 694630 7208 694830
rect 7408 694630 7418 694830
rect 16998 694630 17008 694830
rect 17208 694630 17218 694830
rect 17398 694630 17408 694830
rect 17608 694630 17618 694830
rect 17798 694630 17808 694830
rect 18008 694630 18018 694830
rect 61034 694740 61044 694920
rect 61224 694740 61234 694920
rect 61034 694735 61234 694740
rect 61374 694920 61574 694925
rect 61374 694740 61384 694920
rect 61564 694740 61574 694920
rect 61374 694735 61574 694740
rect 61714 694920 61914 694925
rect 61714 694740 61724 694920
rect 61904 694740 61914 694920
rect 61714 694735 61914 694740
rect 6598 694230 6608 694430
rect 6808 694230 6818 694430
rect 7198 694230 7208 694430
rect 7408 694230 7418 694430
rect 16998 694230 17008 694430
rect 17208 694230 17218 694430
rect 17398 694230 17408 694430
rect 17608 694230 17618 694430
rect 17798 694230 17808 694430
rect 18008 694230 18018 694430
rect 16998 693830 17008 694030
rect 17208 693830 17218 694030
rect 17398 693830 17408 694030
rect 17608 693830 17618 694030
rect 17798 693830 17808 694030
rect 18008 693830 18018 694030
rect 6598 693630 6608 693830
rect 6808 693630 6818 693830
rect 7198 693630 7208 693830
rect 7408 693630 7418 693830
rect 16998 693430 17008 693630
rect 17208 693430 17218 693630
rect 17398 693430 17408 693630
rect 17608 693430 17618 693630
rect 17798 693430 17808 693630
rect 18008 693430 18018 693630
rect 6598 693230 6608 693430
rect 6808 693230 6818 693430
rect 7198 693230 7208 693430
rect 7408 693230 7418 693430
rect 16908 693230 18008 693330
rect 16908 693030 17008 693230
rect 17208 693030 17408 693230
rect 17608 693030 17808 693230
rect 18008 693030 18018 693230
rect 46320 691800 56400 692040
rect 46320 691560 52800 691800
rect 46400 691400 52800 691560
rect 46600 691200 52800 691400
rect 53400 691200 54000 691800
rect 54600 691200 55200 691800
rect 55800 691200 56400 691800
rect 25008 690212 38420 691132
rect 39340 690212 39346 691132
rect 46600 691000 56400 691200
rect 71374 690660 71384 690860
rect 71584 690660 71594 690860
rect 71974 690660 71984 690860
rect 72184 690660 72194 690860
rect 47100 690278 58858 690400
rect 47100 690222 47222 690278
rect 47278 690222 58858 690278
rect 71374 690260 71384 690460
rect 71584 690260 71594 690460
rect 71974 690260 71984 690460
rect 72184 690260 72194 690460
rect 25008 689690 25928 690212
rect 47100 689968 58858 690222
rect 47100 689912 47222 689968
rect 47278 689912 58858 689968
rect 47100 689888 58858 689912
rect 47100 689832 47222 689888
rect 47278 689832 58858 689888
rect 71374 689860 71384 690060
rect 71584 689860 71594 690060
rect 71974 689860 71984 690060
rect 72184 689860 72194 690060
rect 18048 689650 27236 689690
rect 18048 689530 18068 689650
rect 18188 689530 27236 689650
rect 18048 689470 27236 689530
rect 18048 689350 18068 689470
rect 18188 689350 27236 689470
rect 47100 689578 58858 689832
rect 47100 689522 47222 689578
rect 47278 689522 58858 689578
rect 47100 689400 58858 689522
rect 71374 689460 71384 689660
rect 71584 689460 71594 689660
rect 71974 689460 71984 689660
rect 72184 689460 72194 689660
rect 18048 689290 27236 689350
rect 18048 689170 18068 689290
rect 18188 689170 27236 689290
rect 18048 689110 27236 689170
rect 18048 688990 18068 689110
rect 18188 688990 27236 689110
rect 18048 688930 27236 688990
rect 18048 688810 18068 688930
rect 18188 688810 27236 688930
rect 18048 688770 27236 688810
rect 6498 688530 6718 688535
rect 6498 688330 6508 688530
rect 6708 688330 6718 688530
rect 6498 688325 6718 688330
rect 6798 688530 7018 688535
rect 6798 688330 6808 688530
rect 7008 688330 7018 688530
rect 6798 688325 7018 688330
rect 7098 688530 7318 688535
rect 7098 688330 7108 688530
rect 7308 688330 7318 688530
rect 7098 688325 7318 688330
rect 7398 688530 7618 688535
rect 7398 688330 7408 688530
rect 7608 688330 7618 688530
rect 7398 688325 7618 688330
rect 19548 687586 20868 688770
rect 29800 688678 42200 688800
rect 29800 688622 42022 688678
rect 42078 688622 42200 688678
rect 29800 688582 42200 688622
rect 6408 687585 20868 687586
rect 6408 686267 6409 687585
rect 7727 686267 20868 687585
rect 27964 688468 42200 688582
rect 27964 688412 42022 688468
rect 42078 688412 42200 688468
rect 27964 688388 42200 688412
rect 27964 688332 42022 688388
rect 42078 688332 42200 688388
rect 27964 688178 42200 688332
rect 57858 688225 58858 689400
rect 71374 689060 71384 689260
rect 71584 689060 71594 689260
rect 71974 689060 71984 689260
rect 72184 689060 72194 689260
rect 27964 688122 42022 688178
rect 42078 688122 42200 688178
rect 27964 687800 42200 688122
rect 27964 687782 30846 687800
rect 27964 687364 28764 687782
rect 6408 686266 20868 686267
rect 26436 686564 28764 687364
rect 29800 687000 47800 687400
rect 57853 687227 57859 688225
rect 58857 687227 58863 688225
rect 26436 685430 27236 686564
rect 29800 686400 42900 687000
rect 9808 685330 27236 685430
rect 9808 685130 10008 685330
rect 10208 685130 10408 685330
rect 10608 685130 10808 685330
rect 11008 685130 11208 685330
rect 11408 685130 11608 685330
rect 11808 685130 12008 685330
rect 12208 685130 12408 685330
rect 12608 685130 12808 685330
rect 13008 685130 13208 685330
rect 13408 685130 13608 685330
rect 13808 685130 14008 685330
rect 14208 685130 14408 685330
rect 14608 685130 27236 685330
rect 50138 685700 50558 685706
rect 50558 685660 60864 685700
rect 50558 685520 60704 685660
rect 60844 685520 60864 685660
rect 50558 685460 60864 685520
rect 50558 685320 60704 685460
rect 60844 685320 60864 685460
rect 50558 685280 60864 685320
rect 62024 685660 71264 685700
rect 62024 685520 62044 685660
rect 62184 685520 71104 685660
rect 71244 685520 71264 685660
rect 62024 685460 71264 685520
rect 62024 685320 62044 685460
rect 62184 685320 71104 685460
rect 71244 685320 71264 685460
rect 62024 685280 71264 685320
rect 50138 685274 50558 685280
rect 9808 684930 27236 685130
rect 9808 684730 10008 684930
rect 10208 684730 10408 684930
rect 10608 684730 10808 684930
rect 11008 684730 11208 684930
rect 11408 684730 11608 684930
rect 11808 684730 12008 684930
rect 12208 684730 12408 684930
rect 12608 684730 12808 684930
rect 13008 684730 13208 684930
rect 13408 684730 13608 684930
rect 13808 684730 14008 684930
rect 14208 684730 14408 684930
rect 14608 684730 27236 684930
rect 9808 684630 27236 684730
rect 42240 683108 43910 683140
rect 42240 683052 42272 683108
rect 42328 683052 42412 683108
rect 42468 683052 42552 683108
rect 42608 683052 43910 683108
rect 42240 683020 43910 683052
rect 45360 683108 47040 683140
rect 45360 683052 46672 683108
rect 46728 683052 46812 683108
rect 46868 683052 46952 683108
rect 47008 683052 47040 683108
rect 45360 683020 47040 683052
rect 58858 683084 60120 683204
rect 57858 683060 60120 683084
rect 57858 682860 69184 683060
rect 57858 682660 64384 682860
rect 64584 682660 64784 682860
rect 64984 682660 65184 682860
rect 65384 682660 65584 682860
rect 65784 682660 65984 682860
rect 66184 682660 66384 682860
rect 66584 682660 66784 682860
rect 66984 682660 67184 682860
rect 67384 682660 67584 682860
rect 67784 682660 67984 682860
rect 68184 682660 68384 682860
rect 68584 682660 68784 682860
rect 68984 682660 69184 682860
rect 45400 682400 56400 682600
rect 45400 681800 52800 682400
rect 53400 681800 54000 682400
rect 54600 681800 55200 682400
rect 55800 681800 56400 682400
rect 57858 682460 69184 682660
rect 57858 682260 64384 682460
rect 64584 682260 64784 682460
rect 64984 682260 65184 682460
rect 65384 682260 65584 682460
rect 65784 682260 65984 682460
rect 66184 682260 66384 682460
rect 66584 682260 66784 682460
rect 66984 682260 67184 682460
rect 67384 682260 67584 682460
rect 67784 682260 67984 682460
rect 68184 682260 68384 682460
rect 68584 682260 68784 682460
rect 68984 682260 69184 682460
rect 57858 682204 69184 682260
rect 59250 682060 69184 682204
rect 45400 681600 56400 681800
<< via3 >>
rect 17008 698690 17128 698810
rect 17208 698690 17328 698810
rect 17408 698690 17528 698810
rect 17608 698690 17728 698810
rect 17808 698690 17928 698810
rect 6608 694630 6808 694830
rect 7208 694630 7408 694830
rect 17008 694630 17208 694830
rect 17408 694630 17608 694830
rect 17808 694630 18008 694830
rect 61044 694740 61224 694920
rect 61384 694740 61564 694920
rect 61724 694740 61904 694920
rect 6608 694230 6808 694430
rect 7208 694230 7408 694430
rect 17008 694230 17208 694430
rect 17408 694230 17608 694430
rect 17808 694230 18008 694430
rect 17008 693830 17208 694030
rect 17408 693830 17608 694030
rect 17808 693830 18008 694030
rect 6608 693630 6808 693830
rect 7208 693630 7408 693830
rect 17008 693430 17208 693630
rect 17408 693430 17608 693630
rect 17808 693430 18008 693630
rect 6608 693230 6808 693430
rect 7208 693230 7408 693430
rect 17008 693030 17208 693230
rect 17408 693030 17608 693230
rect 17808 693030 18008 693230
rect 52800 691200 53400 691800
rect 54000 691200 54600 691800
rect 55200 691200 55800 691800
rect 38420 690212 39340 691132
rect 71384 690660 71584 690860
rect 71984 690660 72184 690860
rect 71384 690260 71584 690460
rect 71984 690260 72184 690460
rect 71384 689860 71584 690060
rect 71984 689860 72184 690060
rect 71384 689460 71584 689660
rect 71984 689460 72184 689660
rect 6508 688330 6708 688530
rect 6808 688330 7008 688530
rect 7108 688330 7308 688530
rect 7408 688330 7608 688530
rect 6409 686267 7727 687585
rect 71384 689060 71584 689260
rect 71984 689060 72184 689260
rect 57859 687227 58857 688225
rect 10008 685130 10208 685330
rect 10408 685130 10608 685330
rect 10808 685130 11008 685330
rect 11208 685130 11408 685330
rect 11608 685130 11808 685330
rect 12008 685130 12208 685330
rect 12408 685130 12608 685330
rect 12808 685130 13008 685330
rect 13208 685130 13408 685330
rect 13608 685130 13808 685330
rect 14008 685130 14208 685330
rect 14408 685130 14608 685330
rect 50138 685280 50558 685700
rect 10008 684730 10208 684930
rect 10408 684730 10608 684930
rect 10808 684730 11008 684930
rect 11208 684730 11408 684930
rect 11608 684730 11808 684930
rect 12008 684730 12208 684930
rect 12408 684730 12608 684930
rect 12808 684730 13008 684930
rect 13208 684730 13408 684930
rect 13608 684730 13808 684930
rect 14008 684730 14208 684930
rect 14408 684730 14608 684930
rect 57858 683084 58858 684084
rect 64384 682660 64584 682860
rect 64784 682660 64984 682860
rect 65184 682660 65384 682860
rect 65584 682660 65784 682860
rect 65984 682660 66184 682860
rect 66384 682660 66584 682860
rect 66784 682660 66984 682860
rect 67184 682660 67384 682860
rect 67584 682660 67784 682860
rect 67984 682660 68184 682860
rect 68384 682660 68584 682860
rect 68784 682660 68984 682860
rect 52800 681800 53400 682400
rect 54000 681800 54600 682400
rect 55200 681800 55800 682400
rect 64384 682260 64584 682460
rect 64784 682260 64984 682460
rect 65184 682260 65384 682460
rect 65584 682260 65784 682460
rect 65984 682260 66184 682460
rect 66384 682260 66584 682460
rect 66784 682260 66984 682460
rect 67184 682260 67384 682460
rect 67584 682260 67784 682460
rect 67984 682260 68184 682460
rect 68384 682260 68584 682460
rect 68784 682260 68984 682460
<< metal4 >>
rect 9808 698810 17948 698930
rect 9808 698690 17008 698810
rect 17128 698690 17208 698810
rect 17328 698690 17408 698810
rect 17528 698690 17608 698810
rect 17728 698690 17808 698810
rect 17928 698690 17948 698810
rect 9808 698570 17948 698690
rect 9808 695030 14808 698570
rect 6408 694830 14808 695030
rect 6408 694630 6608 694830
rect 6808 694630 7208 694830
rect 7408 694630 14808 694830
rect 6408 694430 14808 694630
rect 6408 694230 6608 694430
rect 6808 694230 7208 694430
rect 7408 694230 14808 694430
rect 6408 693830 14808 694230
rect 6408 693630 6608 693830
rect 6808 693630 7208 693830
rect 7408 693630 14808 693830
rect 6408 693430 14808 693630
rect 6408 693230 6608 693430
rect 6808 693230 7208 693430
rect 7408 693230 14808 693430
rect 6408 693030 14808 693230
rect 6408 688530 7728 688610
rect 6408 688330 6508 688530
rect 6708 688330 6808 688530
rect 7008 688330 7108 688530
rect 7308 688330 7408 688530
rect 7608 688330 7728 688530
rect 6408 687585 7728 688330
rect 6408 686267 6409 687585
rect 7727 686267 7728 687585
rect 6408 684074 7728 686267
rect 9808 685330 14808 693030
rect 16808 694830 18208 695030
rect 16808 694630 17008 694830
rect 17208 694630 17408 694830
rect 17608 694630 17808 694830
rect 18008 694630 18208 694830
rect 61024 694920 69184 694960
rect 61024 694740 61044 694920
rect 61224 694740 61384 694920
rect 61564 694740 61724 694920
rect 61904 694740 69184 694920
rect 61024 694700 69184 694740
rect 16808 694430 18208 694630
rect 16808 694230 17008 694430
rect 17208 694230 17408 694430
rect 17608 694230 17808 694430
rect 18008 694230 18208 694430
rect 16808 694030 18208 694230
rect 16808 693830 17008 694030
rect 17208 693830 17408 694030
rect 17608 693830 17808 694030
rect 18008 693830 18208 694030
rect 16808 693630 18208 693830
rect 16808 693430 17008 693630
rect 17208 693430 17408 693630
rect 17608 693430 17808 693630
rect 18008 693430 18208 693630
rect 16808 693230 18208 693430
rect 16808 693030 17008 693230
rect 17208 693030 17408 693230
rect 17608 693030 17808 693230
rect 18008 693030 18208 693230
rect 16808 686728 18208 693030
rect 52400 691800 56400 692000
rect 52400 691200 52800 691800
rect 53400 691200 54000 691800
rect 54600 691200 55200 691800
rect 55800 691200 56400 691800
rect 38419 691132 39341 691133
rect 38419 690212 38420 691132
rect 39340 690212 39341 691132
rect 38419 690211 39341 690212
rect 52400 690594 56400 691200
rect 64184 691060 69184 694700
rect 59250 690594 61984 691060
rect 52400 688860 61984 690594
rect 64184 690860 72384 691060
rect 64184 690660 71384 690860
rect 71584 690660 71984 690860
rect 72184 690660 72384 690860
rect 64184 690460 72384 690660
rect 64184 690260 71384 690460
rect 71584 690260 71984 690460
rect 72184 690260 72384 690460
rect 64184 690060 72384 690260
rect 64184 689860 71384 690060
rect 71584 689860 71984 690060
rect 72184 689860 72384 690060
rect 64184 689660 72384 689860
rect 64184 689460 71384 689660
rect 71584 689460 71984 689660
rect 72184 689460 72384 689660
rect 64184 689260 72384 689460
rect 64184 689060 71384 689260
rect 71584 689060 71984 689260
rect 72184 689060 72384 689260
rect 64184 688860 72384 689060
rect 9808 685130 10008 685330
rect 10208 685130 10408 685330
rect 10608 685130 10808 685330
rect 11008 685130 11208 685330
rect 11408 685130 11608 685330
rect 11808 685130 12008 685330
rect 12208 685130 12408 685330
rect 12608 685130 12808 685330
rect 13008 685130 13208 685330
rect 13408 685130 13608 685330
rect 13808 685130 14008 685330
rect 14208 685130 14408 685330
rect 14608 685130 14808 685330
rect 9808 684930 14808 685130
rect 9808 684730 10008 684930
rect 10208 684730 10408 684930
rect 10608 684730 10808 684930
rect 11008 684730 11208 684930
rect 11408 684730 11608 684930
rect 11808 684730 12008 684930
rect 12208 684730 12408 684930
rect 12608 684730 12808 684930
rect 13008 684730 13208 684930
rect 13408 684730 13608 684930
rect 13808 684730 14008 684930
rect 14208 684730 14408 684930
rect 14608 684730 14808 684930
rect 16662 684928 20612 686728
rect 9808 684630 14808 684730
rect 16808 684074 18208 684928
rect 18812 658978 20612 684928
rect 38670 682003 39330 686050
rect 49920 685700 50580 686100
rect 49920 685280 50138 685700
rect 50558 685280 50580 685700
rect 35200 673800 40000 682003
rect 35200 673000 35600 673800
rect 36400 673000 37200 673800
rect 38000 673000 38800 673800
rect 39600 673000 40000 673800
rect 35200 670600 40000 673000
rect 49920 673968 50580 685280
rect 52400 682400 56400 688860
rect 57858 688225 58858 688226
rect 57858 687227 57859 688225
rect 58857 687227 58858 688225
rect 57858 684085 58858 687227
rect 57857 684084 58859 684085
rect 57857 683084 57858 684084
rect 58858 683084 58859 684084
rect 57857 683083 58859 683084
rect 52400 681800 52800 682400
rect 53400 681800 54000 682400
rect 54600 681800 55200 682400
rect 55800 681800 56400 682400
rect 64184 682860 69184 688860
rect 64184 682660 64384 682860
rect 64584 682660 64784 682860
rect 64984 682660 65184 682860
rect 65384 682660 65584 682860
rect 65784 682660 65984 682860
rect 66184 682660 66384 682860
rect 66584 682660 66784 682860
rect 66984 682660 67184 682860
rect 67384 682660 67584 682860
rect 67784 682660 67984 682860
rect 68184 682660 68384 682860
rect 68584 682660 68784 682860
rect 68984 682660 69184 682860
rect 64184 682460 69184 682660
rect 64184 682260 64384 682460
rect 64584 682260 64784 682460
rect 64984 682260 65184 682460
rect 65384 682260 65584 682460
rect 65784 682260 65984 682460
rect 66184 682260 66384 682460
rect 66584 682260 66784 682460
rect 66984 682260 67184 682460
rect 67384 682260 67584 682460
rect 67784 682260 67984 682460
rect 68184 682260 68384 682460
rect 68584 682260 68784 682460
rect 68984 682260 69184 682460
rect 64184 682060 69184 682260
rect 52400 680000 56400 681800
rect 49920 673732 50132 673968
rect 50368 673732 50580 673968
rect 49920 673568 50580 673732
rect 49920 673332 50132 673568
rect 50368 673332 50580 673568
rect 49920 673168 50580 673332
rect 49920 672932 50132 673168
rect 50368 672932 50580 673168
rect 49920 672700 50580 672932
rect 35200 669800 35600 670600
rect 36400 669800 37200 670600
rect 38000 669800 38800 670600
rect 39600 669800 40000 670600
rect 35200 667200 40000 669800
rect 35200 666400 35600 667200
rect 36400 666400 37200 667200
rect 38000 666400 38800 667200
rect 39600 666400 40000 667200
rect 35200 662800 40000 666400
rect 54448 658978 56248 680000
rect 18812 657178 56248 658978
<< via4 >>
rect 35600 673000 36400 673800
rect 37200 673000 38000 673800
rect 38800 673000 39600 673800
rect 50132 673732 50368 673968
rect 50132 673332 50368 673568
rect 50132 672932 50368 673168
rect 35600 669800 36400 670600
rect 37200 669800 38000 670600
rect 38800 669800 39600 670600
rect 35600 666400 36400 667200
rect 37200 666400 38000 667200
rect 38800 666400 39600 667200
<< metal5 >>
rect 35200 673968 51300 674200
rect 35200 673800 50132 673968
rect 35200 673000 35600 673800
rect 36400 673000 37200 673800
rect 38000 673000 38800 673800
rect 39600 673732 50132 673800
rect 50368 673732 51300 673968
rect 39600 673568 51300 673732
rect 39600 673332 50132 673568
rect 50368 673332 51300 673568
rect 39600 673168 51300 673332
rect 39600 673000 50132 673168
rect 35200 672932 50132 673000
rect 50368 672932 51300 673168
rect 35200 672700 51300 672932
rect 35200 670600 48300 670900
rect 35200 669800 35600 670600
rect 36400 669800 37200 670600
rect 38000 669800 38800 670600
rect 39600 669800 48300 670600
rect 35200 669500 48300 669800
rect 35200 667200 48300 667600
rect 35200 666400 35600 667200
rect 36400 666400 37200 667200
rect 38000 666400 38800 667200
rect 39600 666400 48300 667200
rect 35200 666200 48300 666400
use constant_gm_fingers#0  constant_gm_fingers#0_0
timestamp 1713027117
transform 1 0 43810 0 1 682900
box -2700 -20020 4420 1140
use diode_connected_nmos  diode_connected_nmos_0 /foss/designs/C2S2_Analog_TestChip/mag
timestamp 1683391037
transform 1 0 16868 0 1 688490
box -60 -60 1254 10360
use diode_connected_nmos  diode_connected_nmos_1
timestamp 1683391037
transform 1 0 6468 0 1 688490
box -60 -60 1254 10360
use diode_connected_nmos  diode_connected_nmos_3
timestamp 1683391037
transform 1 0 60844 0 1 684520
box -60 -60 1254 10360
use diode_connected_nmos  diode_connected_nmos_7
timestamp 1683391037
transform 1 0 71244 0 1 684520
box -60 -60 1254 10360
use OTA_fingers_031123_NON_FLAT#0  OTA_fingers_031123_NON_FLAT#0_0
timestamp 1713027127
transform 1 0 42740 0 1 684710
box -5940 -310 9780 16550
<< labels >>
rlabel metal3 56683 689400 57683 690400 1 VP
port 3 n
rlabel metal3 29800 686400 30800 687400 1 VOUT
port 6 n
rlabel metal3 29800 687800 30800 688800 1 VN
port 7 n
rlabel metal4 35200 662800 40000 665000 1 VSS
port 8 n
rlabel metal4 52400 680000 56400 684000 1 VDDA
port 5 n
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
