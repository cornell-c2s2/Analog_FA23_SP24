magic
tech sky130A
magscale 1 2
timestamp 1712004182
<< error_s >>
rect 4730 1360 4792 1366
rect 4730 1326 4742 1360
rect 4730 1320 4792 1326
rect 3521 605 3579 611
rect 3521 571 3533 605
rect 3521 565 3579 571
rect 4730 432 4792 438
rect 4730 398 4742 432
rect 4730 392 4792 398
rect 3521 295 3579 301
rect 3521 261 3533 295
rect 3521 255 3579 261
<< nwell >>
rect 1270 -630 1560 -620
rect 1258 -651 1560 -630
rect 1260 -1233 1560 -652
rect 1258 -1260 1560 -1233
rect 1880 -630 2170 -620
rect 1880 -1260 2182 -630
<< pwell >>
rect 1090 -620 2340 -480
rect 1090 -630 1270 -620
rect 1090 -1260 1258 -630
rect 1560 -1260 1880 -620
rect 2170 -630 2340 -620
rect 2182 -1260 2340 -630
rect 1090 -1320 2340 -1260
rect 1090 -1390 1260 -1320
rect 1740 -1330 1750 -1320
rect 2170 -1390 2340 -1320
rect 1090 -1426 1296 -1390
rect 2142 -1426 2340 -1390
<< psubdiff >>
rect 1150 -560 2290 -520
rect 1150 -1356 1190 -560
rect 1700 -660 1740 -560
rect 1150 -1360 1296 -1356
rect 1700 -1360 1740 -1100
rect 2250 -1356 2290 -560
rect 1150 -1380 1330 -1360
rect 1150 -1390 1296 -1380
rect 2142 -1390 2290 -1356
<< psubdiffcont >>
rect 1700 -1100 1740 -660
<< locali >>
rect 1150 -560 2290 -520
rect 1150 -1356 1190 -560
rect 1700 -660 1740 -560
rect 1150 -1360 1296 -1356
rect 1700 -1360 1740 -1100
rect 2250 -1356 2290 -560
rect 1150 -1380 1330 -1360
rect 1150 -1390 1296 -1380
rect 2142 -1390 2290 -1356
<< metal1 >>
rect -2090 590 -1890 790
rect -1360 530 -1160 730
rect -880 490 -680 690
rect -2190 140 -1990 340
rect -1640 150 -1440 350
rect -1310 -20 -1110 180
rect -670 -30 -470 170
rect 0 0 200 200
rect 760 -200 2660 -20
rect 760 -260 1560 -200
rect 1870 -260 2660 -200
rect 640 -380 650 -290
rect 730 -380 740 -290
rect 1600 -380 1670 -290
rect 1760 -380 1840 -290
rect 2700 -380 2710 -290
rect 2790 -380 2800 -290
rect 760 -450 1560 -410
rect 1880 -440 2670 -410
rect 1870 -450 2670 -440
rect 760 -480 1590 -450
rect 480 -630 1440 -540
rect 480 -680 1170 -630
rect 1160 -720 1170 -680
rect 1270 -720 1440 -630
rect 470 -830 480 -740
rect 580 -750 1060 -740
rect 1530 -750 1590 -480
rect 580 -820 880 -750
rect 580 -830 590 -820
rect 870 -830 880 -820
rect 1050 -830 1060 -750
rect 1510 -760 1590 -750
rect 870 -850 1060 -830
rect 880 -860 1060 -850
rect 1480 -810 1590 -760
rect 1840 -480 2670 -450
rect 1840 -750 1910 -480
rect 2160 -640 2170 -630
rect 2000 -720 2170 -640
rect 2270 -720 2280 -630
rect 1840 -760 1930 -750
rect 1840 -810 1960 -760
rect 880 -880 1020 -860
rect 600 -940 840 -880
rect 600 -1270 650 -940
rect 1480 -1060 1560 -810
rect 1870 -1060 1960 -810
rect 2600 -949 2840 -889
rect 1480 -1120 1570 -1060
rect 1650 -1120 1660 -1060
rect 1800 -1130 1960 -1060
rect 1160 -1260 1170 -1170
rect 1270 -1250 1440 -1170
rect 1270 -1260 1280 -1250
rect 350 -1340 650 -1270
rect 700 -1340 710 -1270
rect 800 -1340 810 -1270
rect 1800 -1300 1880 -1130
rect 2000 -1240 2170 -1170
rect 2160 -1260 2170 -1240
rect 2270 -1260 2280 -1170
rect 2790 -1279 2840 -949
rect 600 -1380 650 -1340
rect 1340 -1360 1880 -1300
rect 2020 -1340 2030 -1280
rect 2100 -1340 2110 -1280
rect 2040 -1350 2110 -1340
rect 2620 -1350 2630 -1280
rect 2730 -1350 2740 -1280
rect 2790 -1349 3090 -1279
rect 600 -1390 670 -1380
rect 430 -1510 470 -1410
rect 550 -1510 560 -1410
rect 430 -2170 550 -1510
rect 600 -2180 680 -1390
rect 790 -1750 860 -1390
rect 1340 -1530 1400 -1360
rect 1460 -1420 1580 -1410
rect 1460 -1490 1470 -1420
rect 1560 -1490 1580 -1420
rect 1860 -1420 1980 -1410
rect 1860 -1490 1880 -1420
rect 1960 -1490 1980 -1420
rect 1860 -1500 1980 -1490
rect 2040 -1530 2100 -1350
rect 2790 -1380 2840 -1349
rect 2750 -1390 2840 -1380
rect 1340 -1540 1410 -1530
rect 2030 -1540 2100 -1530
rect 1340 -1550 1440 -1540
rect 1360 -1750 1440 -1550
rect 790 -1940 1440 -1750
rect 790 -2170 860 -1940
rect 600 -2210 670 -2180
rect 600 -2220 640 -2210
rect 350 -2290 640 -2220
rect 710 -2240 850 -2230
rect 710 -2310 730 -2240
rect 830 -2310 850 -2240
rect 710 -2320 850 -2310
rect 1360 -2320 1440 -1940
rect 1590 -2320 1850 -1540
rect 2000 -1550 2100 -1540
rect 2000 -1750 2080 -1550
rect 2580 -1750 2650 -1400
rect 2000 -1940 2650 -1750
rect 2000 -2320 2080 -1940
rect 2580 -2180 2650 -1940
rect 2740 -1402 2840 -1390
rect 2740 -2178 2746 -1402
rect 2760 -2178 2840 -1402
rect 2740 -2190 2840 -2178
rect 2770 -2219 2840 -2190
rect 2800 -2229 2840 -2219
rect 2600 -2250 2740 -2240
rect 2600 -2310 2640 -2250
rect 2720 -2310 2740 -2250
rect 2800 -2299 3090 -2229
rect 2600 -2320 2740 -2310
rect 1660 -2340 1770 -2320
rect 1150 -2400 1160 -2340
rect 1270 -2360 1280 -2340
rect 1270 -2400 1580 -2360
rect 1150 -2420 1580 -2400
rect 1670 -2500 1760 -2340
rect 2160 -2360 2170 -2340
rect 1860 -2410 2170 -2360
rect 2280 -2410 2290 -2340
rect 1860 -2430 2290 -2410
rect 820 -2580 2620 -2500
rect 820 -2620 1600 -2580
rect 1840 -2620 2620 -2580
rect 1650 -2750 1790 -2630
<< via1 >>
rect 650 -380 730 -290
rect 1670 -380 1760 -290
rect 2710 -380 2790 -290
rect 1170 -720 1270 -630
rect 480 -830 580 -740
rect 880 -830 1050 -750
rect 2170 -720 2270 -630
rect 1570 -1120 1650 -1060
rect 1170 -1260 1270 -1170
rect 710 -1340 800 -1270
rect 2170 -1260 2270 -1170
rect 2030 -1340 2100 -1280
rect 2630 -1350 2730 -1280
rect 470 -1510 550 -1410
rect 1470 -1490 1560 -1420
rect 1880 -1490 1960 -1420
rect 730 -2310 830 -2240
rect 2640 -2310 2720 -2250
rect 1160 -2400 1270 -2340
rect 2170 -2410 2280 -2340
<< metal2 >>
rect 650 -290 780 -280
rect 730 -380 780 -290
rect 650 -410 780 -380
rect 1670 -290 1760 -280
rect 1670 -390 1760 -380
rect 2650 -290 2820 -280
rect 2650 -380 2710 -290
rect 2790 -380 2820 -290
rect 470 -740 580 -730
rect 470 -830 480 -740
rect 470 -1410 580 -830
rect 680 -1260 780 -410
rect 2650 -410 2820 -380
rect 1170 -630 1270 -620
rect 1160 -720 1170 -660
rect 880 -750 1050 -740
rect 880 -840 1050 -830
rect 1160 -1170 1270 -720
rect 2170 -630 2280 -620
rect 2270 -720 2280 -630
rect 1160 -1260 1170 -1170
rect 680 -1270 800 -1260
rect 680 -1340 710 -1270
rect 680 -1350 800 -1340
rect 470 -1520 550 -1510
rect 680 -2230 780 -1350
rect 1160 -1410 1270 -1260
rect 1570 -1060 1650 -1050
rect 1570 -1280 1650 -1120
rect 2170 -1170 2280 -720
rect 2270 -1260 2280 -1170
rect 2030 -1280 2100 -1270
rect 1570 -1340 2030 -1280
rect 2030 -1350 2100 -1340
rect 2170 -1410 2280 -1260
rect 2650 -1270 2750 -410
rect 2630 -1280 2750 -1270
rect 2730 -1350 2750 -1280
rect 2630 -1360 2750 -1350
rect 1160 -1420 1560 -1410
rect 1160 -1490 1470 -1420
rect 680 -2240 830 -2230
rect 680 -2310 730 -2240
rect 680 -2320 830 -2310
rect 1160 -2340 1270 -1490
rect 1470 -1500 1560 -1490
rect 1880 -1420 2280 -1410
rect 1960 -1490 2280 -1420
rect 1880 -1500 1960 -1490
rect 1160 -2410 1270 -2400
rect 2170 -2340 2280 -1490
rect 2640 -2250 2750 -1360
rect 2720 -2310 2750 -2250
rect 2640 -2320 2750 -2310
rect 2170 -2420 2280 -2410
<< via2 >>
rect 650 -380 730 -290
rect 1670 -380 1760 -290
rect 2710 -380 2790 -290
rect 880 -830 1050 -750
<< metal3 >>
rect 690 -285 2750 -280
rect 640 -290 2800 -285
rect 640 -380 650 -290
rect 730 -380 1670 -290
rect 1760 -380 2710 -290
rect 2790 -380 2800 -290
rect 640 -385 2800 -380
rect 690 -390 2750 -385
rect 870 -750 1060 -745
rect 870 -830 880 -750
rect 1050 -830 1060 -750
rect 870 -835 1060 -830
use sky130_fd_pr__cap_var_lvt_CYVAFU  XC1
timestamp 1711936448
transform 1 0 1409 0 1 -942
box -151 -318 151 318
use sky130_fd_pr__cap_var_lvt_CYVAFU  XC2
timestamp 1711936448
transform 1 0 2031 0 1 -942
box -151 -318 151 318
use sky130_fd_pr__nfet_01v8_lvt_648S5X  XM1
timestamp 1711936448
transform 1 0 3550 0 1 433
box -211 -310 211 310
use sky130_fd_pr__pfet_01v8_lvt_4QFHB3  XM2
timestamp 1712003522
transform 1 0 4761 0 1 879
box -231 -619 231 619
use sky130_fd_pr__nfet_01v8_lvt_AWHWK2  XM3
timestamp 1711942804
transform 0 1 2274 -1 0 -334
box -256 -610 256 610
use sky130_fd_pr__nfet_01v8_lvt_AWHWK2  XM4
timestamp 1711942804
transform 0 1 1160 -1 0 -334
box -256 -610 256 610
use sky130_fd_pr__pfet_01v8_lvt_4QFHB3  XM6
timestamp 1712003522
transform 1 0 3057 0 1 -1791
box -231 -619 231 619
use sky130_fd_pr__pfet_01v8_lvt_4QFHB3  XM7
timestamp 1712003522
transform 1 0 385 0 1 -1781
box -231 -619 231 619
use sky130_fd_pr__pfet_01v8_lvt_4QFHB3  XM9
timestamp 1712003522
transform -1 0 2701 0 -1 -1791
box -231 -619 231 619
use sky130_fd_pr__nfet_01v8_lvt_64Z3AY  XM10
timestamp 1712001983
transform 0 -1 941 1 0 -909
box -211 -279 211 279
use sky130_fd_pr__nfet_01v8_lvt_64Z3AY  XM11
timestamp 1712001983
transform 0 1 2499 -1 0 -919
box -211 -279 211 279
use sky130_fd_pr__nfet_01v8_lvt_AWHWK2  XM12
timestamp 1711942804
transform 1 0 550 0 1 1678
box -256 -610 256 610
use sky130_fd_pr__nfet_01v8_lvt_T2JW3B  XM13
timestamp 1711941703
transform 0 1 1719 -1 0 -2690
box -256 -1119 256 1119
use sky130_fd_pr__pfet_01v8_lvt_4QFHB3  XM14
timestamp 1712003522
transform -1 0 741 0 -1 -1781
box -231 -619 231 619
use sky130_fd_pr__nfet_01v8_lvt_AWHWK2  XM15
timestamp 1711942804
transform 1 0 1922 0 1 -1930
box -256 -610 256 610
use sky130_fd_pr__nfet_01v8_lvt_AWHWK2  XM17
timestamp 1711942804
transform 1 0 1516 0 1 -1930
box -256 -610 256 610
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 VDD
port 0 nsew
flabel metal1 -1310 -20 -1110 180 0 FreeSans 256 0 0 0 CLK
port 6 nsew
flabel metal1 -670 -30 -470 170 0 FreeSans 256 0 0 0 VIP
port 4 nsew
flabel metal1 -880 490 -680 690 0 FreeSans 256 0 0 0 IB
port 5 nsew
flabel metal1 -1360 530 -1160 730 0 FreeSans 256 0 0 0 VIN
port 3 nsew
flabel metal1 -1640 150 -1440 350 0 FreeSans 256 0 0 0 VON
port 2 nsew
flabel metal1 -2090 590 -1890 790 0 FreeSans 256 0 0 0 VOP
port 1 nsew
flabel metal1 -2190 140 -1990 340 0 FreeSans 256 0 0 0 VSS
port 7 nsew
<< end >>
