magic
tech sky130A
magscale 1 2
timestamp 1714802873
<< nwell >>
rect 5120 4210 5470 4700
rect 5120 2070 5480 2690
<< nsubdiff >>
rect 5190 4630 5420 4660
rect 5190 4560 5220 4630
rect 5380 4560 5420 4630
rect 5190 4530 5420 4560
rect 5220 2240 5380 2270
rect 5220 2140 5250 2240
rect 5350 2140 5380 2240
rect 5220 2110 5380 2140
<< nsubdiffcont >>
rect 5220 4560 5380 4630
rect 5250 2140 5350 2240
<< viali >>
rect 5190 4630 5420 4660
rect 5190 4560 5220 4630
rect 5220 4560 5380 4630
rect 5380 4560 5420 4630
rect 5190 4530 5420 4560
rect 5182 4136 5242 4186
rect 5390 4150 5430 4190
rect 5182 2686 5232 2736
rect 5390 2720 5440 2760
rect 5220 2240 5380 2270
rect 5220 2140 5250 2240
rect 5250 2140 5350 2240
rect 5350 2140 5380 2240
rect 5220 2110 5380 2140
<< metal1 >>
rect 3640 5290 3840 5490
rect 6870 5050 7050 5110
rect 1650 4790 1850 4990
rect 4210 4950 5430 5000
rect 4210 4700 4570 4950
rect 5080 4796 5430 4950
rect 5650 4850 7050 5050
rect 8020 4980 8220 5180
rect 5080 4700 5432 4796
rect 4210 4660 5432 4700
rect 4210 4580 5190 4660
rect 4792 4556 5190 4580
rect 5162 4530 5190 4556
rect 5420 4530 5432 4660
rect 5162 4436 5432 4530
rect 5650 4200 5770 4850
rect 5430 4196 5770 4200
rect 5042 4192 5252 4196
rect 5042 4186 5254 4192
rect 5042 4136 5182 4186
rect 5242 4136 5254 4186
rect 5378 4190 5770 4196
rect 5378 4150 5390 4190
rect 5430 4150 5770 4190
rect 5378 4144 5770 4150
rect 5430 4140 5770 4144
rect 5042 4130 5254 4136
rect 5042 4126 5252 4130
rect 5162 3966 5432 3976
rect 5162 3816 5432 3826
rect 5100 3340 5300 3540
rect 5162 3056 5432 3066
rect 1120 2780 1320 2980
rect 5162 2906 5432 2916
rect 5420 2766 5740 2780
rect 5378 2760 5740 2766
rect 5062 2746 5242 2756
rect 5022 2736 5242 2746
rect 5022 2686 5182 2736
rect 5232 2686 5242 2736
rect 5378 2720 5390 2760
rect 5440 2720 5740 2760
rect 5378 2714 5740 2720
rect 5420 2700 5740 2714
rect 5062 2676 5242 2686
rect 5176 2674 5238 2676
rect 5160 2350 5440 2410
rect 5130 2340 5440 2350
rect 4490 2326 5440 2340
rect 4462 2270 5440 2326
rect 4462 2250 5220 2270
rect 4370 2180 5220 2250
rect 4370 1830 4580 2180
rect 5110 2110 5220 2180
rect 5380 2110 5440 2270
rect 5110 1830 5440 2110
rect 4370 1630 5440 1830
rect 5620 1920 5740 2700
rect 5620 1720 6950 1920
rect 3770 1130 3970 1330
<< via1 >>
rect 4570 4700 5080 4950
rect 5162 3826 5432 3966
rect 5162 2916 5432 3056
rect 4580 1830 5110 2180
<< metal2 >>
rect 4570 4950 5080 4960
rect 4570 4690 5080 4700
rect 5152 3826 5162 3966
rect 5432 3826 5442 3966
rect 5152 2916 5162 3056
rect 5432 2916 5442 3056
rect 4580 2190 5110 2200
rect 4580 1810 5110 1820
<< via2 >>
rect 4570 4700 5080 4950
rect 5162 3826 5432 3966
rect 5162 2916 5432 3056
rect 4580 2180 5110 2190
rect 4580 1830 5110 2180
rect 4580 1820 5110 1830
<< metal3 >>
rect 4560 4950 5090 4955
rect 4560 4700 4570 4950
rect 5080 4700 5090 4950
rect 4560 4695 5090 4700
rect 5157 3966 5437 3976
rect 5157 3826 5162 3966
rect 5432 3826 5437 3966
rect 5157 3816 5437 3826
rect 5157 3056 5437 3066
rect 5157 2916 5162 3056
rect 5432 2916 5437 3056
rect 5157 2906 5437 2916
rect 9260 2790 9270 2980
rect 9480 2790 9490 2980
rect 4570 2190 5120 2195
rect 4570 1820 4580 2190
rect 5110 1820 5120 2190
rect 4570 1815 5120 1820
<< via3 >>
rect 4570 4700 5080 4950
rect 5162 3826 5432 3966
rect 5162 2916 5432 3056
rect 9270 2790 9480 2980
rect 4580 1820 5110 2190
<< metal4 >>
rect 4569 4950 5081 4951
rect 4569 4700 4570 4950
rect 5080 4700 5081 4950
rect 4569 4699 5081 4700
rect 4122 3966 5442 3976
rect 4122 3826 5162 3966
rect 5432 3826 5442 3966
rect 4122 3816 5442 3826
rect 4122 3056 5442 3066
rect 4122 2916 5162 3056
rect 5432 2916 5442 3056
rect 4122 2906 5442 2916
rect 9240 2980 9500 3000
rect 9240 2790 9270 2980
rect 9480 2790 9500 2980
rect 4579 2190 5111 2191
rect 4579 1840 4580 2190
rect 3170 1820 4580 1840
rect 5110 1840 5111 2190
rect 9240 1840 9500 2790
rect 5110 1820 9500 1840
rect 3170 1590 9500 1820
<< via4 >>
rect 4570 4700 5080 4950
rect 4580 1820 5110 2190
<< metal5 >>
rect 4540 4950 6960 5060
rect 4540 4700 4570 4950
rect 5080 4700 6960 4950
rect 4540 4650 6960 4700
rect 6460 4580 6960 4650
rect 4550 2190 6950 2450
rect 4550 1820 4580 2190
rect 5110 1820 6950 2190
rect 4550 1800 6950 1820
rect 4556 1796 5134 1800
use class_AB_v3_sym  class_AB_v3_sym_0 /foss/designs/Analog_FA23_SP24/ComparatorLayout/magic
timestamp 1713498221
transform 0 1 4324 -1 0 5162
box -330 -3260 4030 800
use RSfetsym  RSfetsym_0 /foss/designs/Analog_FA23_SP24/RSlatch/magic
timestamp 1714233353
transform 0 -1 6750 1 0 1970
box -350 -3040 3210 290
use sky130_fd_sc_hd__buf_1  x63 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 5160 0 -1 2948
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  x65
timestamp 1701704242
transform 1 0 5160 0 1 3924
box -38 -48 314 592
<< labels >>
flabel metal1 5160 4770 5360 4970 0 FreeSans 256 0 0 0 VDD
port 0 nsew
flabel metal1 1120 2780 1320 2980 0 FreeSans 256 0 0 0 GND
port 1 nsew
flabel metal1 1650 4790 1850 4990 0 FreeSans 256 0 0 0 IB
port 4 nsew
flabel metal1 3640 5290 3840 5490 0 FreeSans 256 0 0 0 VIN
port 3 nsew
flabel metal1 3770 1130 3970 1330 0 FreeSans 256 0 0 0 VN
port 2 nsew
flabel metal1 5100 3340 5300 3540 0 FreeSans 256 0 0 0 CLK
port 5 nsew
flabel metal1 8020 4980 8220 5180 0 FreeSans 256 0 0 0 Q
port 6 nsew
<< end >>
