magic
tech sky130A
magscale 1 2
timestamp 1709390584
<< error_p >>
rect 3875 12931 3910 12965
rect 48634 12931 48669 12965
rect 3876 12912 3910 12931
rect 48635 12912 48669 12931
rect 3895 11617 3910 12912
rect 3929 12878 3964 12912
rect 5262 12878 5297 12912
rect 3929 11617 3963 12878
rect 5263 12859 5297 12878
rect 6667 12859 6720 12860
rect 3929 11583 3944 11617
rect 5282 11564 5297 12859
rect 5316 12825 5351 12859
rect 6649 12825 6720 12859
rect 5316 11564 5350 12825
rect 6650 12824 6720 12825
rect 6667 12790 6738 12824
rect 10248 12790 10283 12824
rect 5316 11530 5331 11564
rect 6667 11511 6737 12790
rect 10249 12771 10283 12790
rect 6667 11475 6720 11511
rect 10268 11458 10283 12771
rect 10302 12737 10337 12771
rect 13847 12737 13882 12771
rect 10302 11458 10336 12737
rect 13848 12718 13882 12737
rect 10302 11424 10317 11458
rect 13867 11405 13882 12718
rect 13901 12684 13936 12718
rect 20448 12684 20483 12701
rect 13901 11405 13935 12684
rect 20449 12683 20483 12684
rect 20449 12647 20519 12683
rect 20466 12613 20537 12647
rect 13901 11371 13916 11405
rect 20466 11352 20536 12613
rect 48654 11617 48669 12912
rect 48688 12878 48723 12912
rect 50021 12878 50056 12912
rect 48688 11617 48722 12878
rect 50022 12859 50056 12878
rect 51426 12859 51479 12860
rect 48688 11583 48703 11617
rect 50041 11564 50056 12859
rect 50075 12825 50110 12859
rect 51408 12825 51479 12859
rect 50075 11564 50109 12825
rect 51409 12824 51479 12825
rect 51426 12790 51497 12824
rect 55007 12790 55042 12824
rect 50075 11530 50090 11564
rect 51426 11511 51496 12790
rect 55008 12771 55042 12790
rect 51426 11475 51479 11511
rect 55027 11458 55042 12771
rect 55061 12737 55096 12771
rect 58606 12737 58641 12771
rect 55061 11458 55095 12737
rect 58607 12718 58641 12737
rect 55061 11424 55076 11458
rect 58626 11405 58641 12718
rect 58660 12684 58695 12718
rect 65207 12684 65242 12701
rect 58660 11405 58694 12684
rect 65208 12683 65242 12684
rect 65208 12647 65278 12683
rect 65225 12613 65296 12647
rect 58660 11371 58675 11405
rect 65225 11352 65295 12613
rect 20466 11316 20519 11352
rect 65225 11316 65278 11352
rect 40905 10509 40940 10543
rect 85664 10509 85699 10543
rect 40906 10490 40940 10509
rect 85665 10490 85699 10509
rect 39947 10441 40005 10447
rect 40143 10441 40201 10447
rect 40339 10441 40397 10447
rect 40535 10441 40593 10447
rect 40731 10441 40789 10447
rect 39947 10407 39959 10441
rect 40143 10407 40155 10441
rect 40339 10407 40351 10441
rect 40535 10407 40547 10441
rect 40731 10407 40743 10441
rect 39947 10401 40005 10407
rect 40143 10401 40201 10407
rect 40339 10401 40397 10407
rect 40535 10401 40593 10407
rect 40731 10401 40789 10407
rect 28823 1915 28857 1933
rect 28823 1879 28893 1915
rect 28840 1845 28911 1879
rect 30651 1845 30686 1879
rect 28840 566 28910 1845
rect 30652 1826 30686 1845
rect 28840 530 28893 566
rect 30671 513 30686 1826
rect 30705 1792 30740 1826
rect 32480 1792 32515 1809
rect 30705 513 30739 1792
rect 32481 1791 32515 1792
rect 32481 1755 32551 1791
rect 32498 1721 32569 1755
rect 30705 479 30720 513
rect 32498 460 32568 1721
rect 34310 952 34344 1006
rect 32498 424 32551 460
rect 34329 407 34344 952
rect 34363 918 34398 952
rect 34363 407 34397 918
rect 34363 373 34378 407
rect 35642 354 35657 952
rect 35676 354 35710 1006
rect 35676 320 35691 354
rect 36239 301 36254 1149
rect 36273 301 36307 1203
rect 39849 331 39907 337
rect 40045 331 40103 337
rect 40241 331 40299 337
rect 40437 331 40495 337
rect 40633 331 40691 337
rect 36273 267 36288 301
rect 39849 297 39861 331
rect 40045 297 40057 331
rect 40241 297 40253 331
rect 40437 297 40449 331
rect 40633 297 40645 331
rect 39849 291 39907 297
rect 40045 291 40103 297
rect 40241 291 40299 297
rect 40437 291 40495 297
rect 40633 291 40691 297
rect 40925 195 40940 10490
rect 40959 10456 40994 10490
rect 42166 10456 42201 10490
rect 40959 195 40993 10456
rect 42167 10437 42201 10456
rect 84706 10441 84764 10447
rect 84902 10441 84960 10447
rect 85098 10441 85156 10447
rect 85294 10441 85352 10447
rect 85490 10441 85548 10447
rect 41208 10388 41266 10394
rect 41404 10388 41462 10394
rect 41600 10388 41658 10394
rect 41796 10388 41854 10394
rect 41992 10388 42050 10394
rect 41208 10354 41220 10388
rect 41404 10354 41416 10388
rect 41600 10354 41612 10388
rect 41796 10354 41808 10388
rect 41992 10354 42004 10388
rect 41208 10348 41266 10354
rect 41404 10348 41462 10354
rect 41600 10348 41658 10354
rect 41796 10348 41854 10354
rect 41992 10348 42050 10354
rect 41110 278 41168 284
rect 41306 278 41364 284
rect 41502 278 41560 284
rect 41698 278 41756 284
rect 41894 278 41952 284
rect 41110 244 41122 278
rect 41306 244 41318 278
rect 41502 244 41514 278
rect 41698 244 41710 278
rect 41894 244 41906 278
rect 41110 238 41168 244
rect 41306 238 41364 244
rect 41502 238 41560 244
rect 41698 238 41756 244
rect 41894 238 41952 244
rect 40959 161 40974 195
rect 42186 142 42201 10437
rect 42220 10403 42255 10437
rect 43427 10403 43462 10437
rect 42220 142 42254 10403
rect 43428 10384 43462 10403
rect 84706 10407 84718 10441
rect 84902 10407 84914 10441
rect 85098 10407 85110 10441
rect 85294 10407 85306 10441
rect 85490 10407 85502 10441
rect 84706 10401 84764 10407
rect 84902 10401 84960 10407
rect 85098 10401 85156 10407
rect 85294 10401 85352 10407
rect 85490 10401 85548 10407
rect 42469 10335 42527 10341
rect 42665 10335 42723 10341
rect 42861 10335 42919 10341
rect 43057 10335 43115 10341
rect 43253 10335 43311 10341
rect 42469 10301 42481 10335
rect 42665 10301 42677 10335
rect 42861 10301 42873 10335
rect 43057 10301 43069 10335
rect 43253 10301 43265 10335
rect 42469 10295 42527 10301
rect 42665 10295 42723 10301
rect 42861 10295 42919 10301
rect 43057 10295 43115 10301
rect 43253 10295 43311 10301
rect 42371 225 42429 231
rect 42567 225 42625 231
rect 42763 225 42821 231
rect 42959 225 43017 231
rect 43155 225 43213 231
rect 42371 191 42383 225
rect 42567 191 42579 225
rect 42763 191 42775 225
rect 42959 191 42971 225
rect 43155 191 43167 225
rect 42371 185 42429 191
rect 42567 185 42625 191
rect 42763 185 42821 191
rect 42959 185 43017 191
rect 43155 185 43213 191
rect 42220 108 42235 142
rect 43447 89 43462 10384
rect 43481 89 43499 10384
rect 73582 1915 73616 1933
rect 73582 1879 73652 1915
rect 73599 1845 73670 1879
rect 75410 1845 75445 1879
rect 73599 566 73669 1845
rect 75411 1826 75445 1845
rect 73599 530 73652 566
rect 75430 513 75445 1826
rect 75464 1792 75499 1826
rect 77239 1792 77274 1809
rect 75464 513 75498 1792
rect 77240 1791 77274 1792
rect 77240 1755 77310 1791
rect 77257 1721 77328 1755
rect 75464 479 75479 513
rect 77257 460 77327 1721
rect 79069 952 79103 1006
rect 77257 424 77310 460
rect 79088 407 79103 952
rect 79122 918 79157 952
rect 79122 407 79156 918
rect 79122 373 79137 407
rect 80401 354 80416 952
rect 80435 354 80469 1006
rect 80435 320 80450 354
rect 80998 301 81013 1149
rect 81032 301 81066 1203
rect 84608 331 84666 337
rect 84804 331 84862 337
rect 85000 331 85058 337
rect 85196 331 85254 337
rect 85392 331 85450 337
rect 81032 267 81047 301
rect 84608 297 84620 331
rect 84804 297 84816 331
rect 85000 297 85012 331
rect 85196 297 85208 331
rect 85392 297 85404 331
rect 84608 291 84666 297
rect 84804 291 84862 297
rect 85000 291 85058 297
rect 85196 291 85254 297
rect 85392 291 85450 297
rect 85684 195 85699 10490
rect 85718 10456 85753 10490
rect 86925 10456 86960 10490
rect 85718 195 85752 10456
rect 86926 10437 86960 10456
rect 85967 10388 86025 10394
rect 86163 10388 86221 10394
rect 86359 10388 86417 10394
rect 86555 10388 86613 10394
rect 86751 10388 86809 10394
rect 85967 10354 85979 10388
rect 86163 10354 86175 10388
rect 86359 10354 86371 10388
rect 86555 10354 86567 10388
rect 86751 10354 86763 10388
rect 85967 10348 86025 10354
rect 86163 10348 86221 10354
rect 86359 10348 86417 10354
rect 86555 10348 86613 10354
rect 86751 10348 86809 10354
rect 85869 278 85927 284
rect 86065 278 86123 284
rect 86261 278 86319 284
rect 86457 278 86515 284
rect 86653 278 86711 284
rect 85869 244 85881 278
rect 86065 244 86077 278
rect 86261 244 86273 278
rect 86457 244 86469 278
rect 86653 244 86665 278
rect 85869 238 85927 244
rect 86065 238 86123 244
rect 86261 238 86319 244
rect 86457 238 86515 244
rect 86653 238 86711 244
rect 85718 161 85733 195
rect 86945 142 86960 10437
rect 86979 10403 87014 10437
rect 88186 10403 88221 10437
rect 86979 142 87013 10403
rect 88187 10384 88221 10403
rect 87228 10335 87286 10341
rect 87424 10335 87482 10341
rect 87620 10335 87678 10341
rect 87816 10335 87874 10341
rect 88012 10335 88070 10341
rect 87228 10301 87240 10335
rect 87424 10301 87436 10335
rect 87620 10301 87632 10335
rect 87816 10301 87828 10335
rect 88012 10301 88024 10335
rect 87228 10295 87286 10301
rect 87424 10295 87482 10301
rect 87620 10295 87678 10301
rect 87816 10295 87874 10301
rect 88012 10295 88070 10301
rect 87130 225 87188 231
rect 87326 225 87384 231
rect 87522 225 87580 231
rect 87718 225 87776 231
rect 87914 225 87972 231
rect 87130 191 87142 225
rect 87326 191 87338 225
rect 87522 191 87534 225
rect 87718 191 87730 225
rect 87914 191 87926 225
rect 87130 185 87188 191
rect 87326 185 87384 191
rect 87522 185 87580 191
rect 87718 185 87776 191
rect 87914 185 87972 191
rect 86979 108 86994 142
rect 88206 89 88221 10384
rect 88240 10350 88275 10384
rect 88240 5245 88274 10350
rect 88489 10282 88547 10288
rect 88685 10282 88743 10288
rect 88881 10282 88939 10288
rect 89077 10282 89135 10288
rect 89273 10282 89331 10288
rect 88489 10248 88501 10282
rect 88685 10248 88697 10282
rect 88881 10248 88893 10282
rect 89077 10248 89089 10282
rect 89273 10248 89285 10282
rect 88489 10242 88547 10248
rect 88685 10242 88743 10248
rect 88881 10242 88939 10248
rect 89077 10242 89135 10248
rect 89273 10242 89331 10248
rect 88240 89 88258 5245
rect 99236 3915 99271 3932
rect 99237 3914 99271 3915
rect 99237 3878 99254 3914
rect 98409 3847 98449 3853
rect 98583 3847 98641 3853
rect 98775 3847 98833 3853
rect 98967 3847 99025 3853
rect 98583 3813 98595 3847
rect 98775 3813 98787 3847
rect 98967 3813 98979 3847
rect 98409 3807 98449 3813
rect 98583 3807 98641 3813
rect 98775 3807 98833 3813
rect 98967 3807 99025 3813
rect 98487 2719 98545 2725
rect 98679 2719 98737 2725
rect 98871 2719 98929 2725
rect 99063 2719 99121 2725
rect 98487 2685 98499 2719
rect 98679 2685 98691 2719
rect 98871 2685 98883 2719
rect 99063 2685 99075 2719
rect 98487 2679 98545 2685
rect 98679 2679 98737 2685
rect 98871 2679 98929 2685
rect 99063 2679 99121 2685
rect 100399 3878 100452 3879
rect 99307 3844 99325 3878
rect 100381 3844 100452 3878
rect 99307 2583 99324 3844
rect 100382 3843 100452 3844
rect 100399 3809 100470 3843
rect 102486 3809 102521 3826
rect 99536 3776 99594 3782
rect 99728 3776 99786 3782
rect 99920 3776 99978 3782
rect 100112 3776 100170 3782
rect 99536 3742 99548 3776
rect 99728 3742 99740 3776
rect 99920 3742 99932 3776
rect 100112 3742 100124 3776
rect 99536 3736 99594 3742
rect 99728 3736 99786 3742
rect 99920 3736 99978 3742
rect 100112 3736 100170 3742
rect 99440 2666 99498 2672
rect 99632 2666 99690 2672
rect 99824 2666 99882 2672
rect 100016 2666 100074 2672
rect 100208 2666 100266 2672
rect 99440 2632 99452 2666
rect 99632 2632 99644 2666
rect 99824 2632 99836 2666
rect 100016 2632 100028 2666
rect 100208 2632 100220 2666
rect 99440 2626 99498 2632
rect 99632 2626 99690 2632
rect 99824 2626 99882 2632
rect 100016 2626 100074 2632
rect 100208 2626 100266 2632
rect 100399 2530 100469 3809
rect 102487 3808 102521 3809
rect 102487 3772 102504 3808
rect 100681 3741 100739 3747
rect 100873 3741 100931 3747
rect 101065 3741 101123 3747
rect 101257 3741 101315 3747
rect 101449 3741 101507 3747
rect 101641 3741 101699 3747
rect 101833 3741 101891 3747
rect 102025 3741 102083 3747
rect 102217 3741 102275 3747
rect 100681 3707 100693 3741
rect 100873 3707 100885 3741
rect 101065 3707 101077 3741
rect 101257 3707 101269 3741
rect 101449 3707 101461 3741
rect 101641 3707 101653 3741
rect 101833 3707 101845 3741
rect 102025 3707 102037 3741
rect 102217 3707 102229 3741
rect 100681 3701 100739 3707
rect 100873 3701 100931 3707
rect 101065 3701 101123 3707
rect 101257 3701 101315 3707
rect 101449 3701 101507 3707
rect 101641 3701 101699 3707
rect 101833 3701 101891 3707
rect 102025 3701 102083 3707
rect 102217 3701 102275 3707
rect 100585 2613 100643 2619
rect 100777 2613 100835 2619
rect 100969 2613 101027 2619
rect 101161 2613 101219 2619
rect 101353 2613 101411 2619
rect 101545 2613 101603 2619
rect 101737 2613 101795 2619
rect 101929 2613 101987 2619
rect 102121 2613 102179 2619
rect 102313 2613 102371 2619
rect 100585 2579 100597 2613
rect 100777 2579 100789 2613
rect 100969 2579 100981 2613
rect 101161 2579 101173 2613
rect 101353 2579 101365 2613
rect 101545 2579 101557 2613
rect 101737 2579 101749 2613
rect 101929 2579 101941 2613
rect 102121 2579 102133 2613
rect 102313 2579 102325 2613
rect 100585 2573 100643 2579
rect 100777 2573 100835 2579
rect 100969 2573 101027 2579
rect 101161 2573 101219 2579
rect 101353 2573 101411 2579
rect 101545 2573 101603 2579
rect 101737 2573 101795 2579
rect 101929 2573 101987 2579
rect 102121 2573 102179 2579
rect 102313 2573 102371 2579
rect 100399 2494 100452 2530
rect 102557 3738 102575 3772
rect 102557 2477 102574 3738
rect 102786 3670 102844 3676
rect 102978 3670 103036 3676
rect 103170 3670 103228 3676
rect 103362 3670 103420 3676
rect 102786 3636 102798 3670
rect 102978 3636 102990 3670
rect 103170 3636 103182 3670
rect 103362 3636 103374 3670
rect 102786 3630 102844 3636
rect 102978 3630 103036 3636
rect 103170 3630 103228 3636
rect 103362 3630 103420 3636
rect 102690 2560 102748 2566
rect 102882 2560 102940 2566
rect 103074 2560 103132 2566
rect 103266 2560 103324 2566
rect 103458 2560 103516 2566
rect 102690 2526 102702 2560
rect 102882 2526 102894 2560
rect 103074 2526 103086 2560
rect 103266 2526 103278 2560
rect 103458 2526 103470 2560
rect 102690 2520 102748 2526
rect 102882 2520 102940 2526
rect 103074 2520 103132 2526
rect 103266 2520 103324 2526
rect 103458 2520 103516 2526
rect 43481 55 43496 89
rect 88240 55 88255 89
<< error_s >>
rect 114410 58341 114445 58375
rect 114411 58322 114445 58341
rect 43499 10350 43516 10384
rect 43499 89 43515 10350
rect 43730 10282 43788 10288
rect 43926 10282 43984 10288
rect 44122 10282 44180 10288
rect 44318 10282 44376 10288
rect 44514 10282 44572 10288
rect 43730 10248 43742 10282
rect 43926 10248 43938 10282
rect 44122 10248 44134 10282
rect 44318 10248 44330 10282
rect 44514 10248 44526 10282
rect 43730 10242 43788 10248
rect 43926 10242 43984 10248
rect 44122 10242 44180 10248
rect 44318 10242 44376 10248
rect 44514 10242 44572 10248
rect 43632 172 43690 178
rect 43828 172 43886 178
rect 44024 172 44082 178
rect 44220 172 44278 178
rect 44416 172 44474 178
rect 43632 138 43644 172
rect 43828 138 43840 172
rect 44024 138 44036 172
rect 44220 138 44232 172
rect 44416 138 44428 172
rect 43632 132 43690 138
rect 43828 132 43886 138
rect 44024 132 44082 138
rect 44220 132 44278 138
rect 44416 132 44474 138
rect 88258 89 88274 5245
rect 91605 3915 91640 3932
rect 91606 3914 91640 3915
rect 91606 3878 91676 3914
rect 92768 3878 92821 3879
rect 89800 3847 89858 3853
rect 89992 3847 90050 3853
rect 90184 3847 90242 3853
rect 90376 3847 90434 3853
rect 90568 3847 90626 3853
rect 90760 3847 90818 3853
rect 90952 3847 91010 3853
rect 91144 3847 91202 3853
rect 91336 3847 91394 3853
rect 89800 3813 89812 3847
rect 89992 3813 90004 3847
rect 90184 3813 90196 3847
rect 90376 3813 90388 3847
rect 90568 3813 90580 3847
rect 90760 3813 90772 3847
rect 90952 3813 90964 3847
rect 91144 3813 91156 3847
rect 91336 3813 91348 3847
rect 91623 3844 91694 3878
rect 92750 3844 92821 3878
rect 89800 3807 89858 3813
rect 89992 3807 90050 3813
rect 90184 3807 90242 3813
rect 90376 3807 90434 3813
rect 90568 3807 90626 3813
rect 90760 3807 90818 3813
rect 90952 3807 91010 3813
rect 91144 3807 91202 3813
rect 91336 3807 91394 3813
rect 89704 2719 89762 2725
rect 89896 2719 89954 2725
rect 90088 2719 90146 2725
rect 90280 2719 90338 2725
rect 90472 2719 90530 2725
rect 90664 2719 90722 2725
rect 90856 2719 90914 2725
rect 91048 2719 91106 2725
rect 91240 2719 91298 2725
rect 91432 2719 91490 2725
rect 89704 2685 89716 2719
rect 89896 2685 89908 2719
rect 90088 2685 90100 2719
rect 90280 2685 90292 2719
rect 90472 2685 90484 2719
rect 90664 2685 90676 2719
rect 90856 2685 90868 2719
rect 91048 2685 91060 2719
rect 91240 2685 91252 2719
rect 91432 2685 91444 2719
rect 89704 2679 89762 2685
rect 89896 2679 89954 2685
rect 90088 2679 90146 2685
rect 90280 2679 90338 2685
rect 90472 2679 90530 2685
rect 90664 2679 90722 2685
rect 90856 2679 90914 2685
rect 91048 2679 91106 2685
rect 91240 2679 91298 2685
rect 91432 2679 91490 2685
rect 91623 2583 91693 3844
rect 92751 3843 92821 3844
rect 97431 3847 97489 3853
rect 97623 3847 97681 3853
rect 97815 3847 97873 3853
rect 98007 3847 98065 3853
rect 98199 3847 98257 3853
rect 98391 3847 98409 3853
rect 92768 3809 92839 3843
rect 94855 3809 94890 3826
rect 91905 3776 91963 3782
rect 92097 3776 92155 3782
rect 92289 3776 92347 3782
rect 92481 3776 92539 3782
rect 91905 3742 91917 3776
rect 92097 3742 92109 3776
rect 92289 3742 92301 3776
rect 92481 3742 92493 3776
rect 91905 3736 91963 3742
rect 92097 3736 92155 3742
rect 92289 3736 92347 3742
rect 92481 3736 92539 3742
rect 91809 2666 91867 2672
rect 92001 2666 92059 2672
rect 92193 2666 92251 2672
rect 92385 2666 92443 2672
rect 92577 2666 92635 2672
rect 91809 2632 91821 2666
rect 92001 2632 92013 2666
rect 92193 2632 92205 2666
rect 92385 2632 92397 2666
rect 92577 2632 92589 2666
rect 91809 2626 91867 2632
rect 92001 2626 92059 2632
rect 92193 2626 92251 2632
rect 92385 2626 92443 2632
rect 92577 2626 92635 2632
rect 91623 2547 91676 2583
rect 92768 2530 92838 3809
rect 94856 3808 94890 3809
rect 97431 3813 97443 3847
rect 97623 3813 97635 3847
rect 97815 3813 97827 3847
rect 98007 3813 98019 3847
rect 98199 3813 98211 3847
rect 98391 3813 98403 3847
rect 94856 3772 94926 3808
rect 97431 3807 97489 3813
rect 97623 3807 97681 3813
rect 97815 3807 97873 3813
rect 98007 3807 98065 3813
rect 98199 3807 98257 3813
rect 98391 3807 98409 3813
rect 96018 3772 96071 3773
rect 93050 3741 93108 3747
rect 93242 3741 93300 3747
rect 93434 3741 93492 3747
rect 93626 3741 93684 3747
rect 93818 3741 93876 3747
rect 94010 3741 94068 3747
rect 94202 3741 94260 3747
rect 94394 3741 94452 3747
rect 94586 3741 94644 3747
rect 93050 3707 93062 3741
rect 93242 3707 93254 3741
rect 93434 3707 93446 3741
rect 93626 3707 93638 3741
rect 93818 3707 93830 3741
rect 94010 3707 94022 3741
rect 94202 3707 94214 3741
rect 94394 3707 94406 3741
rect 94586 3707 94598 3741
rect 94873 3738 94944 3772
rect 96000 3738 96071 3772
rect 93050 3701 93108 3707
rect 93242 3701 93300 3707
rect 93434 3701 93492 3707
rect 93626 3701 93684 3707
rect 93818 3701 93876 3707
rect 94010 3701 94068 3707
rect 94202 3701 94260 3707
rect 94394 3701 94452 3707
rect 94586 3701 94644 3707
rect 92954 2613 93012 2619
rect 93146 2613 93204 2619
rect 93338 2613 93396 2619
rect 93530 2613 93588 2619
rect 93722 2613 93780 2619
rect 93914 2613 93972 2619
rect 94106 2613 94164 2619
rect 94298 2613 94356 2619
rect 94490 2613 94548 2619
rect 94682 2613 94740 2619
rect 92954 2579 92966 2613
rect 93146 2579 93158 2613
rect 93338 2579 93350 2613
rect 93530 2579 93542 2613
rect 93722 2579 93734 2613
rect 93914 2579 93926 2613
rect 94106 2579 94118 2613
rect 94298 2579 94310 2613
rect 94490 2579 94502 2613
rect 94682 2579 94694 2613
rect 92954 2573 93012 2579
rect 93146 2573 93204 2579
rect 93338 2573 93396 2579
rect 93530 2573 93588 2579
rect 93722 2573 93780 2579
rect 93914 2573 93972 2579
rect 94106 2573 94164 2579
rect 94298 2573 94356 2579
rect 94490 2573 94548 2579
rect 94682 2573 94740 2579
rect 92768 2494 92821 2530
rect 94873 2477 94943 3738
rect 96001 3737 96071 3738
rect 96018 3703 96089 3737
rect 96539 3703 96574 3720
rect 95155 3670 95213 3676
rect 95347 3670 95405 3676
rect 95539 3670 95597 3676
rect 95731 3670 95789 3676
rect 95155 3636 95167 3670
rect 95347 3636 95359 3670
rect 95539 3636 95551 3670
rect 95731 3636 95743 3670
rect 95155 3630 95213 3636
rect 95347 3630 95405 3636
rect 95539 3630 95597 3636
rect 95731 3630 95789 3636
rect 95059 2560 95117 2566
rect 95251 2560 95309 2566
rect 95443 2560 95501 2566
rect 95635 2560 95693 2566
rect 95827 2560 95885 2566
rect 95059 2526 95071 2560
rect 95251 2526 95263 2560
rect 95443 2526 95455 2560
rect 95635 2526 95647 2560
rect 95827 2526 95839 2560
rect 95059 2520 95117 2526
rect 95251 2520 95309 2526
rect 95443 2520 95501 2526
rect 95635 2520 95693 2526
rect 95827 2520 95885 2526
rect 94873 2441 94926 2477
rect 96018 2424 96088 3703
rect 96540 3702 96574 3703
rect 96540 3666 96610 3702
rect 96557 3632 96628 3666
rect 96018 2388 96071 2424
rect 96557 2371 96627 3632
rect 97335 2719 97393 2725
rect 97527 2719 97585 2725
rect 97719 2719 97777 2725
rect 97911 2719 97969 2725
rect 98103 2719 98161 2725
rect 98295 2719 98353 2725
rect 97335 2685 97347 2719
rect 97527 2685 97539 2719
rect 97719 2685 97731 2719
rect 97911 2685 97923 2719
rect 98103 2685 98115 2719
rect 98295 2685 98307 2719
rect 97335 2679 97393 2685
rect 97527 2679 97585 2685
rect 97719 2679 97777 2685
rect 97911 2679 97969 2685
rect 98103 2679 98161 2685
rect 98295 2679 98353 2685
rect 103649 3772 103702 3773
rect 103631 3738 103702 3772
rect 103632 3737 103702 3738
rect 103649 3703 103720 3737
rect 104170 3703 104205 3720
rect 103649 2424 103719 3703
rect 104171 3702 104205 3703
rect 104171 3666 104241 3702
rect 104188 3632 104259 3666
rect 103649 2388 103702 2424
rect 104188 2371 104258 3632
rect 113039 2702 113052 2715
rect 108742 2621 108773 2653
rect 113003 2381 113056 2702
rect 96557 2335 96610 2371
rect 104188 2335 104241 2371
rect 113005 2103 113018 2137
rect 113039 2069 113052 2171
rect 88391 172 88449 178
rect 88587 172 88645 178
rect 88783 172 88841 178
rect 88979 172 89037 178
rect 89175 172 89233 178
rect 88391 138 88403 172
rect 88587 138 88599 172
rect 88783 138 88795 172
rect 88979 138 88991 172
rect 89175 138 89187 172
rect 88391 132 88449 138
rect 88587 132 88645 138
rect 88783 132 88841 138
rect 88979 132 89037 138
rect 89175 132 89233 138
rect 114430 -17 114445 58322
rect 114464 58288 114499 58322
rect 115835 58288 115870 58322
rect 114464 -17 114498 58288
rect 115836 58269 115870 58288
rect 114464 -51 114479 -17
rect 115855 -70 115870 58269
rect 115889 58235 115924 58269
rect 117260 58235 117295 58269
rect 115889 -70 115923 58235
rect 117261 58216 117295 58235
rect 115889 -104 115904 -70
rect 117280 -123 117295 58216
rect 117314 58182 117349 58216
rect 117314 -123 117348 58182
rect 117314 -157 117329 -123
<< error_ps >>
rect 99254 2547 99307 3914
rect 102504 2441 102557 3808
use C2S2_Amp_F_I  x1
timestamp 1709390584
transform 1 0 53 0 1 11034
box -53 -11034 44706 4392
use C2S2_Amp_F_I  x2
timestamp 1709390584
transform 1 0 44812 0 1 11034
box -53 -11034 44706 4392
use 1Bit_Clk_ADC  x3
timestamp 1709390584
transform 1 0 104818 0 1 2000
box -38 -2000 8238 1192
use 1Bit_DAC  x4
timestamp 1709390584
transform 1 0 97202 0 1 2000
box -53 -2000 7578 1985
use 1Bit_DAC_Inv  x5
timestamp 1709390584
transform 1 0 89571 0 1 2000
box -53 -2000 7578 1985
use sky130_fd_pr__res_xhigh_po_5p73_7B4CKM  XR1
timestamp 1709390584
transform 1 0 115167 0 1 29126
box -739 -29232 739 29232
use sky130_fd_pr__res_xhigh_po_5p73_7B4CKM  XR2
timestamp 1709390584
transform 1 0 116592 0 1 29073
box -739 -29232 739 29232
use sky130_fd_pr__res_xhigh_po_5p73_7B4CKM  XR3
timestamp 1709390584
transform 1 0 118017 0 1 29020
box -739 -29232 739 29232
use sky130_fd_pr__res_xhigh_po_5p73_7B4CKM  XR5
timestamp 1709390584
transform 1 0 113742 0 1 29179
box -739 -29232 739 29232
<< end >>
