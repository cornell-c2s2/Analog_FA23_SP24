magic
tech sky130A
magscale 1 2
timestamp 1717123183
<< nwell >>
rect 5120 4210 5470 4700
rect 5120 2070 5480 2690
<< pwell >>
rect 5150 3720 5440 4100
rect 5072 2770 5526 3212
<< psubdiff >>
rect 5150 3820 5440 3850
rect 5150 3750 5180 3820
rect 5410 3750 5440 3820
rect 5150 3720 5440 3750
rect 5120 3160 5480 3190
rect 5120 3080 5160 3160
rect 5440 3080 5480 3160
rect 5120 3050 5480 3080
<< nsubdiff >>
rect 5190 4630 5420 4660
rect 5190 4560 5220 4630
rect 5380 4560 5420 4630
rect 5190 4530 5420 4560
rect 5220 2240 5380 2270
rect 5220 2140 5250 2240
rect 5350 2140 5380 2240
rect 5220 2110 5380 2140
<< psubdiffcont >>
rect 5180 3750 5410 3820
rect 5160 3080 5440 3160
<< nsubdiffcont >>
rect 5220 4560 5380 4630
rect 5250 2140 5350 2240
<< viali >>
rect 5190 4630 5420 4660
rect 5190 4560 5220 4630
rect 5220 4560 5380 4630
rect 5380 4560 5420 4630
rect 5190 4530 5420 4560
rect 5182 4136 5242 4186
rect 5390 4150 5430 4190
rect 5150 3820 5440 3850
rect 5150 3750 5180 3820
rect 5180 3750 5410 3820
rect 5410 3750 5440 3820
rect 5150 3720 5440 3750
rect 5120 3160 5480 3190
rect 5120 3080 5160 3160
rect 5160 3080 5440 3160
rect 5440 3080 5480 3160
rect 5120 3050 5480 3080
rect 5182 2686 5232 2736
rect 5390 2720 5440 2760
rect 5220 2240 5380 2270
rect 5220 2140 5250 2240
rect 5250 2140 5350 2240
rect 5350 2140 5380 2240
rect 5220 2110 5380 2140
<< metal1 >>
rect 3640 5290 3840 5490
rect 6870 5050 7050 5110
rect 1650 4790 1850 4990
rect 4210 4950 5430 5000
rect 4210 4700 4570 4950
rect 5080 4796 5430 4950
rect 5650 4850 7050 5050
rect 5080 4700 5432 4796
rect 4210 4660 5432 4700
rect 4210 4580 5190 4660
rect 4792 4556 5190 4580
rect 5162 4530 5190 4556
rect 5420 4530 5432 4660
rect 5162 4436 5432 4530
rect 5650 4200 5770 4850
rect 5430 4196 5770 4200
rect 5042 4192 5252 4196
rect 5042 4186 5254 4192
rect 5042 4136 5182 4186
rect 5242 4136 5254 4186
rect 5378 4190 5770 4196
rect 5378 4150 5390 4190
rect 5430 4150 5770 4190
rect 5378 4144 5770 4150
rect 5430 4140 5770 4144
rect 5042 4130 5254 4136
rect 5042 4126 5252 4130
rect 5162 3966 5432 3976
rect 5130 3850 5162 3880
rect 5432 3850 5460 3880
rect 5130 3720 5150 3850
rect 5440 3720 5460 3850
rect 5130 3690 5460 3720
rect 5100 3340 5300 3540
rect 5100 3190 5510 3200
rect 5100 3050 5120 3190
rect 5480 3050 5510 3190
rect 5100 3030 5162 3050
rect 1120 2780 1320 2980
rect 5432 3030 5510 3050
rect 5162 2906 5432 2916
rect 5420 2766 5740 2780
rect 5378 2760 5740 2766
rect 5062 2746 5242 2756
rect 5022 2736 5242 2746
rect 5022 2686 5182 2736
rect 5232 2686 5242 2736
rect 5378 2720 5390 2760
rect 5440 2720 5740 2760
rect 5378 2714 5740 2720
rect 5420 2700 5740 2714
rect 5062 2676 5242 2686
rect 5176 2674 5238 2676
rect 5160 2350 5440 2410
rect 5130 2340 5440 2350
rect 4490 2326 5440 2340
rect 4462 2270 5440 2326
rect 4462 2262 5220 2270
rect 4462 2250 4718 2262
rect 4370 2044 4718 2250
rect 5062 2110 5220 2262
rect 5380 2110 5440 2270
rect 5062 2044 5440 2110
rect 4370 1630 5440 2044
rect 5620 1920 5740 2700
rect 5620 1720 6950 1920
rect 8020 1620 8220 1820
rect 3770 1130 3970 1330
<< via1 >>
rect 4570 4700 5080 4950
rect 5162 3850 5432 3966
rect 5162 3826 5432 3850
rect 5162 3050 5432 3056
rect 5162 2916 5432 3050
rect 4718 2044 5062 2262
<< metal2 >>
rect 4570 4950 5080 4960
rect 4570 4690 5080 4700
rect 5152 3826 5162 3966
rect 5432 3826 5442 3966
rect 5152 2916 5162 3056
rect 5432 2916 5442 3056
rect 4718 2262 5062 2272
rect 4718 2034 5062 2044
<< via2 >>
rect 4570 4700 5080 4950
rect 5162 3826 5432 3966
rect 5162 2916 5432 3056
rect 4718 2044 5062 2262
<< metal3 >>
rect 4560 4950 5090 4955
rect 4560 4700 4570 4950
rect 5080 4700 5090 4950
rect 4560 4695 5090 4700
rect 5157 3966 5437 3976
rect 5157 3826 5162 3966
rect 5432 3826 5437 3966
rect 5157 3816 5437 3826
rect 5157 3056 5437 3066
rect 5157 2916 5162 3056
rect 5432 2916 5437 3056
rect 5157 2906 5437 2916
rect 9260 2790 9490 2980
rect 4708 2262 5072 2267
rect 4708 2044 4718 2262
rect 5062 2044 5072 2262
rect 4708 2039 5072 2044
<< via3 >>
rect 4570 4700 5080 4950
rect 5162 3826 5432 3966
rect 5162 2916 5432 3056
rect 4718 2044 5062 2262
<< metal4 >>
rect 4569 4950 5081 4951
rect 4569 4700 4570 4950
rect 5080 4700 5081 4950
rect 4569 4699 5081 4700
rect 4122 3966 5442 3976
rect 4122 3826 5162 3966
rect 5432 3826 5442 3966
rect 4122 3816 5442 3826
rect 9250 3810 10170 4020
rect 4122 3056 5442 3066
rect 4122 2916 5162 3056
rect 5432 2916 5442 3056
rect 4122 2906 5442 2916
rect 9900 1840 10170 3810
rect 3170 1590 10170 1840
<< via4 >>
rect 4570 4700 5080 4950
rect 4692 2262 5090 2308
rect 4692 2044 4718 2262
rect 4718 2044 5062 2262
rect 5062 2044 5090 2262
rect 4692 2004 5090 2044
<< metal5 >>
rect 4540 4950 6960 5060
rect 4540 4700 4570 4950
rect 5080 4700 6960 4950
rect 4540 4650 6960 4700
rect 6460 4580 6960 4650
rect 4550 2308 6950 2450
rect 4550 2004 4692 2308
rect 5090 2004 6950 2308
rect 4550 1920 6950 2004
use class_AB_v3_sym  class_AB_v3_sym_0 /foss/designs/Analog_FA23_SP24/ComparatorLayout/magic
timestamp 1716869746
transform 0 1 4324 -1 0 5162
box -330 -3260 4030 800
use RSfetsym  RSfetsym_0 /foss/designs/Analog_FA23_SP24/RSlatch/magic
timestamp 1717123183
transform 0 -1 6750 -1 0 4830
box -350 -3040 3210 290
use sky130_fd_sc_hd__buf_1  x63 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1716869746
transform 1 0 5160 0 -1 2948
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  x65
timestamp 1716869746
transform 1 0 5160 0 1 3924
box -38 -48 314 592
<< labels >>
flabel metal1 5160 4770 5360 4970 0 FreeSans 256 0 0 0 VDD
port 0 nsew
flabel metal1 1120 2780 1320 2980 0 FreeSans 256 0 0 0 GND
port 1 nsew
flabel metal1 1650 4790 1850 4990 0 FreeSans 256 0 0 0 IB
port 4 nsew
flabel metal1 3640 5290 3840 5490 0 FreeSans 256 0 0 0 VIN
port 3 nsew
flabel metal1 3770 1130 3970 1330 0 FreeSans 256 0 0 0 VN
port 2 nsew
flabel metal1 5100 3340 5300 3540 0 FreeSans 256 0 0 0 CLK
port 5 nsew
flabel metal1 8020 1620 8220 1820 0 FreeSans 256 0 0 0 Q
port 6 nsew
<< end >>
