magic
tech sky130A
magscale 1 2
timestamp 1713626893
<< error_p >>
rect 3875 12931 3910 12965
rect 48634 12931 48669 12965
rect 3876 12912 3910 12931
rect 48635 12912 48669 12931
rect 3895 11617 3910 12912
rect 3929 12878 3964 12912
rect 5262 12878 5297 12912
rect 3929 11617 3963 12878
rect 5263 12859 5297 12878
rect 6667 12859 6720 12860
rect 3929 11583 3944 11617
rect 5282 11564 5297 12859
rect 5316 12825 5351 12859
rect 6649 12825 6720 12859
rect 5316 11564 5350 12825
rect 6650 12824 6720 12825
rect 6667 12790 6738 12824
rect 10248 12790 10283 12824
rect 5316 11530 5331 11564
rect 6667 11511 6737 12790
rect 10249 12771 10283 12790
rect 6667 11475 6720 11511
rect 10268 11458 10283 12771
rect 10302 12737 10337 12771
rect 13847 12737 13882 12771
rect 10302 11458 10336 12737
rect 13848 12718 13882 12737
rect 10302 11424 10317 11458
rect 13867 11405 13882 12718
rect 13901 12684 13936 12718
rect 20448 12684 20483 12701
rect 13901 11405 13935 12684
rect 20449 12683 20483 12684
rect 20449 12647 20519 12683
rect 20466 12613 20537 12647
rect 13901 11371 13916 11405
rect 20466 11352 20536 12613
rect 48654 11617 48669 12912
rect 48688 12878 48723 12912
rect 50021 12878 50056 12912
rect 48688 11617 48722 12878
rect 50022 12859 50056 12878
rect 51426 12859 51479 12860
rect 48688 11583 48703 11617
rect 50041 11564 50056 12859
rect 50075 12825 50110 12859
rect 51408 12825 51479 12859
rect 50075 11564 50109 12825
rect 51409 12824 51479 12825
rect 51426 12790 51497 12824
rect 55007 12790 55042 12824
rect 50075 11530 50090 11564
rect 51426 11511 51496 12790
rect 55008 12771 55042 12790
rect 51426 11475 51479 11511
rect 55027 11458 55042 12771
rect 55061 12737 55096 12771
rect 58606 12737 58641 12771
rect 55061 11458 55095 12737
rect 58607 12718 58641 12737
rect 55061 11424 55076 11458
rect 58626 11405 58641 12718
rect 58660 12684 58695 12718
rect 65207 12684 65242 12701
rect 58660 11405 58694 12684
rect 65208 12683 65242 12684
rect 65208 12647 65278 12683
rect 65225 12613 65296 12647
rect 58660 11371 58675 11405
rect 65225 11352 65295 12613
rect 20466 11316 20519 11352
rect 65225 11316 65278 11352
rect 40905 10509 40940 10543
rect 40906 10490 40940 10509
rect 39947 10441 40005 10447
rect 40143 10441 40201 10447
rect 40339 10441 40397 10447
rect 40535 10441 40593 10447
rect 40731 10441 40789 10447
rect 39947 10407 39959 10441
rect 40143 10407 40155 10441
rect 40339 10407 40351 10441
rect 40535 10407 40547 10441
rect 40731 10407 40743 10441
rect 39947 10401 40005 10407
rect 40143 10401 40201 10407
rect 40339 10401 40397 10407
rect 40535 10401 40593 10407
rect 40731 10401 40789 10407
rect 28823 1915 28857 1933
rect 28823 1879 28893 1915
rect 28840 1845 28911 1879
rect 30651 1845 30686 1879
rect 28840 566 28910 1845
rect 30652 1826 30686 1845
rect 28840 530 28893 566
rect 30671 513 30686 1826
rect 30705 1792 30740 1826
rect 32480 1792 32515 1809
rect 30705 513 30739 1792
rect 32481 1791 32515 1792
rect 32481 1755 32551 1791
rect 32498 1721 32569 1755
rect 30705 479 30720 513
rect 32498 460 32568 1721
rect 34310 952 34344 1006
rect 32498 424 32551 460
rect 34329 407 34344 952
rect 34363 918 34398 952
rect 34363 407 34397 918
rect 34363 373 34378 407
rect 35642 354 35657 952
rect 35676 354 35710 1006
rect 35676 320 35691 354
rect 36239 301 36254 1149
rect 36273 301 36307 1203
rect 39849 331 39907 337
rect 40045 331 40103 337
rect 40241 331 40299 337
rect 40437 331 40495 337
rect 40633 331 40691 337
rect 36273 267 36288 301
rect 39849 297 39861 331
rect 40045 297 40057 331
rect 40241 297 40253 331
rect 40437 297 40449 331
rect 40633 297 40645 331
rect 39849 291 39907 297
rect 40045 291 40103 297
rect 40241 291 40299 297
rect 40437 291 40495 297
rect 40633 291 40691 297
rect 40925 195 40940 10490
rect 40959 10456 40994 10490
rect 42166 10456 42201 10490
rect 40959 195 40993 10456
rect 42167 10437 42201 10456
rect 41208 10388 41266 10394
rect 41404 10388 41462 10394
rect 41600 10388 41658 10394
rect 41796 10388 41854 10394
rect 41992 10388 42050 10394
rect 41208 10354 41220 10388
rect 41404 10354 41416 10388
rect 41600 10354 41612 10388
rect 41796 10354 41808 10388
rect 41992 10354 42004 10388
rect 41208 10348 41266 10354
rect 41404 10348 41462 10354
rect 41600 10348 41658 10354
rect 41796 10348 41854 10354
rect 41992 10348 42050 10354
rect 41110 278 41168 284
rect 41306 278 41364 284
rect 41502 278 41560 284
rect 41698 278 41756 284
rect 41894 278 41952 284
rect 41110 244 41122 278
rect 41306 244 41318 278
rect 41502 244 41514 278
rect 41698 244 41710 278
rect 41894 244 41906 278
rect 41110 238 41168 244
rect 41306 238 41364 244
rect 41502 238 41560 244
rect 41698 238 41756 244
rect 41894 238 41952 244
rect 40959 161 40974 195
rect 42186 142 42201 10437
rect 42220 10403 42255 10437
rect 43427 10403 43462 10437
rect 42220 142 42254 10403
rect 43428 10384 43462 10403
rect 42469 10335 42527 10341
rect 42665 10335 42723 10341
rect 42861 10335 42919 10341
rect 43057 10335 43115 10341
rect 43253 10335 43311 10341
rect 42469 10301 42481 10335
rect 42665 10301 42677 10335
rect 42861 10301 42873 10335
rect 43057 10301 43069 10335
rect 43253 10301 43265 10335
rect 42469 10295 42527 10301
rect 42665 10295 42723 10301
rect 42861 10295 42919 10301
rect 43057 10295 43115 10301
rect 43253 10295 43311 10301
rect 42371 225 42429 231
rect 42567 225 42625 231
rect 42763 225 42821 231
rect 42959 225 43017 231
rect 43155 225 43213 231
rect 42371 191 42383 225
rect 42567 191 42579 225
rect 42763 191 42775 225
rect 42959 191 42971 225
rect 43155 191 43167 225
rect 42371 185 42429 191
rect 42567 185 42625 191
rect 42763 185 42821 191
rect 42959 185 43017 191
rect 43155 185 43213 191
rect 42220 108 42235 142
rect 43447 89 43462 10384
rect 43481 89 43499 10384
rect 73582 1915 73616 1933
rect 73582 1879 73652 1915
rect 73599 1845 73670 1879
rect 75410 1845 75445 1879
rect 73599 566 73669 1845
rect 75411 1826 75445 1845
rect 73599 530 73652 566
rect 75430 513 75445 1826
rect 75464 1792 75499 1826
rect 77239 1792 77274 1809
rect 75464 513 75498 1792
rect 77240 1791 77274 1792
rect 77240 1755 77310 1791
rect 77257 1721 77328 1755
rect 75464 479 75479 513
rect 77257 460 77327 1721
rect 79069 952 79103 1006
rect 77257 424 77310 460
rect 79088 407 79103 952
rect 79122 918 79157 952
rect 79122 407 79156 918
rect 79122 373 79137 407
rect 80401 354 80416 952
rect 80435 354 80469 1006
rect 80435 320 80450 354
rect 80998 301 81013 1149
rect 81032 301 81058 1203
rect 81032 267 81047 301
rect 43481 55 43496 89
<< error_s >>
rect 114410 58341 114445 58375
rect 114411 58322 114445 58341
rect 43499 10350 43516 10384
rect 43499 89 43515 10350
rect 43730 10282 43788 10288
rect 43926 10282 43984 10288
rect 44122 10282 44180 10288
rect 44318 10282 44376 10288
rect 44514 10282 44572 10288
rect 43730 10248 43742 10282
rect 43926 10248 43938 10282
rect 44122 10248 44134 10282
rect 44318 10248 44330 10282
rect 44514 10248 44526 10282
rect 43730 10242 43788 10248
rect 43926 10242 43984 10248
rect 44122 10242 44180 10248
rect 44318 10242 44376 10248
rect 44514 10242 44572 10248
rect 113039 2702 113052 2715
rect 113003 2381 113056 2702
rect 96355 2138 96397 2156
rect 96214 2083 96215 2100
rect 96227 2071 96397 2138
rect 113005 2103 113018 2137
rect 96219 2068 96397 2071
rect 113039 2069 113052 2171
rect 96227 1923 96397 2068
rect 96219 1919 96397 1923
rect 96214 1860 96397 1919
rect 96214 1752 96379 1860
rect 96219 1660 96379 1752
rect 96592 1728 96594 1732
rect 96564 1700 96566 1704
rect 96219 1652 96229 1660
rect 94159 1444 94193 1549
rect 94257 1444 94268 1455
rect 94280 1444 94291 1455
rect 94359 1444 94374 1459
rect 96226 1444 96241 1459
rect 93741 930 93807 958
rect 93837 930 93903 958
rect 93933 930 94016 958
rect 93688 915 93695 930
rect 93696 919 94016 930
rect 93696 878 93988 919
rect 93696 872 94002 878
rect 93696 850 94009 872
rect 93696 838 93996 850
rect 93997 838 94009 850
rect 93696 700 93988 838
rect 94244 770 94298 1444
rect 94359 1012 95435 1444
rect 94359 919 95390 1012
rect 94421 888 94451 919
rect 94517 893 94547 919
rect 94613 888 94643 919
rect 94709 893 94739 919
rect 94805 888 94835 919
rect 94901 893 94931 919
rect 94997 888 95027 919
rect 95093 893 95123 919
rect 95189 888 95219 919
rect 95285 893 95315 919
rect 95381 888 95390 919
rect 94403 822 94469 888
rect 94595 822 94661 888
rect 94787 822 94853 888
rect 94979 822 95045 888
rect 95171 822 95237 888
rect 95363 822 95390 888
rect 95794 919 96241 1444
rect 96309 1444 96320 1455
rect 96332 1444 96343 1455
rect 95794 888 95795 919
rect 95861 893 95891 919
rect 95957 888 95987 919
rect 96053 893 96083 919
rect 96149 888 96179 919
rect 95794 822 95813 888
rect 95939 822 96005 888
rect 96131 822 96197 888
rect 96309 770 96343 1444
rect 96564 982 96571 1700
rect 96592 1010 96599 1728
rect 98850 1444 98852 1478
rect 98862 1444 98886 1462
rect 100044 1460 100064 1478
rect 99267 1444 99282 1459
rect 98862 992 99282 1444
rect 98884 934 99282 992
rect 98869 919 99282 934
rect 99350 1444 99361 1455
rect 99373 1444 99384 1455
rect 98902 888 98932 919
rect 98998 893 99028 919
rect 99094 888 99124 919
rect 99190 893 99220 919
rect 98884 822 98950 888
rect 99076 822 99142 888
rect 99350 770 99384 1444
rect 94244 759 95401 770
rect 95783 759 96343 770
rect 98873 759 99384 770
rect 94244 747 95390 759
rect 95794 747 96343 759
rect 98884 747 99384 759
rect 94244 736 95401 747
rect 95783 736 96343 747
rect 98873 736 99384 747
rect 99738 1444 99749 1455
rect 99761 1444 99772 1455
rect 99738 770 99772 1444
rect 99840 1444 99855 1459
rect 100038 1444 100064 1460
rect 99840 1012 100064 1444
rect 99840 934 100030 1012
rect 100038 995 100064 1012
rect 100044 978 100064 995
rect 99840 931 100044 934
rect 99840 919 100045 931
rect 100368 930 100478 958
rect 100508 930 100574 958
rect 100604 930 100716 958
rect 100368 919 100716 930
rect 99902 888 99932 919
rect 99980 888 100030 919
rect 100094 888 100124 919
rect 99884 822 99950 888
rect 100076 822 100126 888
rect 99738 759 100041 770
rect 99738 747 100030 759
rect 99738 736 100041 747
rect 93734 668 93971 700
rect 93723 641 93971 668
rect 93771 600 93831 641
rect 93911 600 93971 641
rect 94244 634 94279 730
rect 100396 700 100688 919
rect 100402 652 100662 700
rect 94244 600 95383 634
rect 98873 623 99242 634
rect 98884 611 99242 623
rect 98873 600 99242 611
rect 100402 600 100462 652
rect 100602 600 100662 652
rect 100688 616 100716 634
rect 100688 600 100696 616
rect 93674 310 93691 510
rect 93702 338 93719 538
rect 93674 190 93701 310
rect 43632 172 43690 178
rect 43828 172 43886 178
rect 44024 172 44082 178
rect 44220 172 44278 178
rect 44416 172 44474 178
rect 43632 138 43644 172
rect 43828 138 43840 172
rect 44024 138 44036 172
rect 44220 138 44232 172
rect 44416 138 44428 172
rect 93702 162 93729 338
rect 43632 132 43690 138
rect 43828 132 43886 138
rect 44024 132 44082 138
rect 44220 132 44278 138
rect 44416 132 44474 138
rect 94244 -680 94291 600
rect 94421 460 94451 486
rect 94499 482 94565 548
rect 94517 460 94547 482
rect 94613 460 94643 486
rect 94691 482 94757 548
rect 94709 460 94739 482
rect 94805 460 94835 486
rect 94883 482 94949 548
rect 94901 460 94931 482
rect 94997 460 95027 486
rect 95075 482 95141 548
rect 95093 460 95123 482
rect 95189 460 95219 486
rect 94359 -540 95281 460
rect 94421 -562 94451 -540
rect 94403 -628 94469 -562
rect 94517 -566 94547 -540
rect 94613 -562 94643 -540
rect 94595 -628 94661 -562
rect 94709 -566 94739 -540
rect 94805 -562 94835 -540
rect 94787 -628 94853 -562
rect 94901 -566 94931 -540
rect 94997 -562 95027 -540
rect 94979 -628 95045 -562
rect 95093 -566 95123 -540
rect 95189 -562 95219 -540
rect 95171 -628 95237 -562
rect 95349 -680 95383 600
rect 98884 460 98918 600
rect 98952 460 98982 486
rect 99030 482 99096 548
rect 99048 460 99078 482
rect 98884 -540 99140 460
rect 98884 -680 98918 -540
rect 98952 -562 98982 -540
rect 98934 -628 99000 -562
rect 99048 -566 99078 -540
rect 99208 -680 99242 600
rect 114430 -17 114445 58322
rect 114464 58288 114499 58322
rect 115835 58288 115870 58322
rect 114464 -17 114498 58288
rect 115836 58269 115870 58288
rect 114464 -51 114479 -17
rect 115855 -70 115870 58269
rect 115889 58235 115924 58269
rect 117260 58235 117295 58269
rect 115889 -70 115923 58235
rect 117261 58216 117295 58235
rect 115889 -104 115904 -70
rect 117280 -123 117295 58216
rect 117314 58182 117349 58216
rect 117314 -123 117348 58182
rect 117314 -157 117329 -123
rect 94244 -714 95383 -680
rect 98873 -691 99242 -680
rect 98884 -703 99242 -691
rect 98873 -714 99242 -703
use C2S2_Amp_F_I  x1 ~/Analog_FA23_SP24/SP24_caravel_user_project_analog/mag
timestamp 1713626893
transform 1 0 53 0 1 11034
box 29796 662788 57684 701260
use C2S2_Amp_F_I  x2
timestamp 1713626893
transform 1 0 44812 0 1 11034
box 29796 662788 57684 701260
use 1Bit_Clk_ADC  x3 ~/Analog_FA23_SP24/SP24_caravel_user_project_analog/mag
timestamp 1713626893
transform 1 0 104818 0 1 2000
box -22500 -15300 5388 23160
use 1Bit_DAC  x4 ~/Analog_FA23_SP24/SP24_caravel_user_project_analog/mag
timestamp 1713148681
transform 1 0 97202 0 1 2000
box 1490 -2780 7005 210
use 1Bit_DAC_Inv  x5 ~/Analog_FA23_SP24/SP24_caravel_user_project_analog/mag
timestamp 1713148681
transform 1 0 89571 0 1 2000
box 1490 -2780 7005 210
use sky130_fd_pr__res_xhigh_po_5p73_7B4CKM  XR1
timestamp 1709390584
transform 1 0 115167 0 1 29126
box -739 -29232 739 29232
use sky130_fd_pr__res_xhigh_po_5p73_7B4CKM  XR2
timestamp 1709390584
transform 1 0 116592 0 1 29073
box -739 -29232 739 29232
use sky130_fd_pr__res_xhigh_po_5p73_7B4CKM  XR3
timestamp 1709390584
transform 1 0 118017 0 1 29020
box -739 -29232 739 29232
use sky130_fd_pr__res_xhigh_po_5p73_7B4CKM  XR5
timestamp 1709390584
transform 1 0 113742 0 1 29179
box -739 -29232 739 29232
<< end >>
