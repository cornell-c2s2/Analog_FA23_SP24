* NGSPICE file created from 16to4_PriorityEncoder_v0p0p1.ext - technology: sky130A

.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
X0 VGND A a_68_297# VNB sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 a_68_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X2 X a_68_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1 ps=0.985 w=0.65 l=0.15
X3 VPWR A a_150_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X4 X a_68_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.146 ps=1.34 w=1 l=0.15
X5 a_150_297# B a_68_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
X0 a_27_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 a_27_297# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X2 a_277_297# B a_205_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X3 VPWR A a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 X a_27_297# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.102 ps=0.99 w=0.65 l=0.15
X5 a_205_297# C a_109_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X6 X a_27_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.148 ps=1.34 w=1 l=0.15
X7 VGND C a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X8 a_109_297# D a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X9 VGND A a_27_297# VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__inv_1 A VGND VNB VPB VPWR Y
X0 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
X0 X a_29_53# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.148 ps=1.34 w=1 l=0.15
X1 a_111_297# C a_29_53# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X2 X a_29_53# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.102 ps=0.99 w=0.65 l=0.15
X3 a_183_297# B a_111_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X4 VPWR A a_183_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X5 a_29_53# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X6 VGND C a_29_53# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X7 VGND A a_29_53# VNB sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
X0 VPWR B a_59_75# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X1 X a_59_75# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.167 ps=1.39 w=1 l=0.15
X2 VGND B a_145_75# VNB sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X3 a_59_75# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X4 X a_59_75# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.112 ps=1.04 w=0.65 l=0.15
X5 a_145_75# A a_59_75# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1 VPWR C a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X2 a_181_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X3 VGND C a_181_47# VNB sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X4 a_27_47# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X5 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X6 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X7 a_109_47# A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
X0 a_27_47# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X1 a_197_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.312 ps=1.68 w=1 l=0.15
X3 a_303_47# C a_197_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X4 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.109 ps=1.36 w=0.42 l=0.15
X5 VPWR D a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.312 pd=1.68 as=0.0588 ps=0.7 w=0.42 l=0.15
X6 VGND D a_303_47# VNB sky130_fd_pr__nfet_01v8 ad=0.196 pd=1.33 as=0.0693 ps=0.75 w=0.42 l=0.15
X7 VPWR B a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X8 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.196 ps=1.33 w=0.65 l=0.15
X9 a_109_47# A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.109 ps=1.36 w=0.42 l=0.15
.ends

.subckt x8to3_Priority_Encoder_v0p2p0 I1 I0 I7 EO GS A2 EI A0 I5 I2 I3 I4 I6 x9/VPB
+ A1 x9/VNB
Xx1 I0 I1 I2 I3 x9/VNB x9/VNB x9/VPB x9/VPB x4/B sky130_fd_sc_hd__or4_1
Xx2 I4 I5 I6 I7 x9/VNB x9/VNB x9/VPB x9/VPB x4/C sky130_fd_sc_hd__or4_1
Xx3 I6 x9/VNB x9/VNB x9/VPB x9/VPB x3/Y sky130_fd_sc_hd__inv_1
Xx4 x9/Y x4/B x4/C x9/VNB x9/VNB x9/VPB x9/VPB EO sky130_fd_sc_hd__or3_1
Xx5 I5 x9/VNB x9/VNB x9/VPB x9/VPB x5/Y sky130_fd_sc_hd__inv_1
Xx6 I4 x9/VNB x9/VNB x9/VPB x9/VPB x6/Y sky130_fd_sc_hd__inv_1
Xx7 I2 x9/VNB x9/VNB x9/VPB x9/VPB x7/Y sky130_fd_sc_hd__inv_1
Xx8 EO EI x9/VNB x9/VNB x9/VPB x9/VPB GS sky130_fd_sc_hd__and2_1
Xx9 EI x9/VNB x9/VNB x9/VPB x9/VPB x9/Y sky130_fd_sc_hd__inv_1
Xx20 I5 x3/Y EI x9/VNB x9/VNB x9/VPB x9/VPB x22/D sky130_fd_sc_hd__and3_1
Xx10 EI I4 x9/VNB x9/VNB x9/VPB x9/VPB x14/A sky130_fd_sc_hd__and2_1
Xx21 EI x21/B x9/VNB x9/VNB x9/VPB x9/VPB x22/B sky130_fd_sc_hd__and2_1
Xx11 EI I5 x9/VNB x9/VNB x9/VPB x9/VPB x14/B sky130_fd_sc_hd__and2_1
Xx22 x22/A x22/B x22/C x22/D x9/VNB x9/VNB x9/VPB x9/VPB A0 sky130_fd_sc_hd__or4_1
Xx12 EI I6 x9/VNB x9/VNB x9/VPB x9/VPB x17/A sky130_fd_sc_hd__and2_1
Xx13 EI I7 x9/VNB x9/VNB x9/VPB x9/VPB x22/A sky130_fd_sc_hd__and2_1
Xx14 x14/A x14/B x17/A x22/A x9/VNB x9/VNB x9/VPB x9/VPB A2 sky130_fd_sc_hd__or4_1
Xx15 I2 x6/Y x5/Y EI x9/VNB x9/VNB x9/VPB x9/VPB x17/C sky130_fd_sc_hd__and4_1
Xx16 I3 x6/Y x5/Y EI x9/VNB x9/VNB x9/VPB x9/VPB x17/D sky130_fd_sc_hd__and4_1
Xx17 x17/A x22/A x17/C x17/D x9/VNB x9/VNB x9/VPB x9/VPB A1 sky130_fd_sc_hd__or4_1
Xx18 x6/Y I1 x7/Y x3/Y x9/VNB x9/VNB x9/VPB x9/VPB x21/B sky130_fd_sc_hd__and4_1
Xx19 EI I3 x6/Y x3/Y x9/VNB x9/VNB x9/VPB x9/VPB x22/C sky130_fd_sc_hd__and4_1
.ends

.subckt sky130_fd_sc_hd__inv_16 A VGND VNB VPB VPWR Y
X0 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X6 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X8 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X10 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X12 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X16 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X17 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X18 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X19 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X20 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X21 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X22 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X23 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X24 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X25 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X26 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X27 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X28 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X29 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X30 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X31 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
X0 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X5 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X6 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
.ends

.subckt x16to4_PriorityEncoder_v0p0p1 A3 EI I15 I14 I13 I12 I11 I10 A2 I9 I8 I7 I6
+ I5 I4 A1 I3 I2 I1 I0 A0
Xx1 x1/A x1/B x9/VNB x9/VNB x9/VPB x9/VPB x1/X sky130_fd_sc_hd__or2_1
Xx2 x2/A x2/B x9/VNB x9/VNB x9/VPB x9/VPB x2/X sky130_fd_sc_hd__or2_1
Xx3 I1 I0 I7 x3/EO x3/GS x3/A2 x7/Y x2/B I5 I2 I3 I4 I6 x9/VPB x1/B x9/VNB x8to3_Priority_Encoder_v0p2p0
Xx4 x9/A x9/VNB x9/VNB x9/VPB x9/VPB A3 sky130_fd_sc_hd__inv_16
Xx5 I9 I8 I15 x7/A x5/GS x5/A2 EI x2/A I13 I10 I11 I12 I14 x9/VPB x1/A x9/VNB x8to3_Priority_Encoder_v0p2p0
Xx6 x9/A x9/VNB x9/VNB x9/VPB x9/VPB A3 sky130_fd_sc_hd__inv_16
Xx7 x7/A x9/VNB x9/VNB x9/VPB x9/VPB x7/Y sky130_fd_sc_hd__inv_1
Xx8 x9/A x9/VNB x9/VNB x9/VPB x9/VPB A3 sky130_fd_sc_hd__inv_16
Xx9 x9/A x9/VNB x9/VNB x9/VPB x9/VPB A3 sky130_fd_sc_hd__inv_16
Xx41 x5/GS x9/VNB x9/VNB x9/VPB x9/VPB x42/A sky130_fd_sc_hd__inv_1
Xx42 x42/A x9/VNB x9/VNB x9/VPB x9/VPB x43/A sky130_fd_sc_hd__inv_4
Xx20 x2/X x9/VNB x9/VNB x9/VPB x9/VPB x21/A sky130_fd_sc_hd__inv_1
Xx43 x43/A x9/VNB x9/VNB x9/VPB x9/VPB x9/A sky130_fd_sc_hd__inv_16
Xx10 x36/Y x9/VNB x9/VNB x9/VPB x9/VPB A2 sky130_fd_sc_hd__inv_16
Xx21 x21/A x9/VNB x9/VNB x9/VPB x9/VPB x22/A sky130_fd_sc_hd__inv_4
Xx11 x5/A2 x3/A2 x9/VNB x9/VNB x9/VPB x9/VPB x34/A sky130_fd_sc_hd__or2_1
Xx22 x22/A x9/VNB x9/VNB x9/VPB x9/VPB x25/A sky130_fd_sc_hd__inv_16
Xx12 x36/Y x9/VNB x9/VNB x9/VPB x9/VPB A2 sky130_fd_sc_hd__inv_16
Xx34 x34/A x9/VNB x9/VNB x9/VPB x9/VPB x35/A sky130_fd_sc_hd__inv_1
Xx23 x25/A x9/VNB x9/VNB x9/VPB x9/VPB A0 sky130_fd_sc_hd__inv_16
Xx13 x36/Y x9/VNB x9/VNB x9/VPB x9/VPB A2 sky130_fd_sc_hd__inv_16
Xx35 x35/A x9/VNB x9/VNB x9/VPB x9/VPB x36/A sky130_fd_sc_hd__inv_4
Xx24 x25/A x9/VNB x9/VNB x9/VPB x9/VPB A0 sky130_fd_sc_hd__inv_16
Xx14 x36/Y x9/VNB x9/VNB x9/VPB x9/VPB A2 sky130_fd_sc_hd__inv_16
Xx36 x36/A x9/VNB x9/VNB x9/VPB x9/VPB x36/Y sky130_fd_sc_hd__inv_16
Xx25 x25/A x9/VNB x9/VNB x9/VPB x9/VPB A0 sky130_fd_sc_hd__inv_16
Xx15 x29/Y x9/VNB x9/VNB x9/VPB x9/VPB A1 sky130_fd_sc_hd__inv_16
Xx16 x29/Y x9/VNB x9/VNB x9/VPB x9/VPB A1 sky130_fd_sc_hd__inv_16
Xx27 x1/X x9/VNB x9/VNB x9/VPB x9/VPB x28/A sky130_fd_sc_hd__inv_1
Xx17 x29/Y x9/VNB x9/VNB x9/VPB x9/VPB A1 sky130_fd_sc_hd__inv_16
Xx28 x28/A x9/VNB x9/VNB x9/VPB x9/VPB x29/A sky130_fd_sc_hd__inv_4
Xx18 x29/Y x9/VNB x9/VNB x9/VPB x9/VPB A1 sky130_fd_sc_hd__inv_16
Xx29 x29/A x9/VNB x9/VNB x9/VPB x9/VPB x29/Y sky130_fd_sc_hd__inv_16
Xx19 x25/A x9/VNB x9/VNB x9/VPB x9/VPB A0 sky130_fd_sc_hd__inv_16
.ends

