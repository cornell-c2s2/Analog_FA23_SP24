magic
tech sky130A
timestamp 1717028336
<< metal1 >>
rect 25800 11100 25900 11200
rect 32700 11100 32900 11200
rect 52000 11100 52200 11200
rect 59000 11100 59100 11200
rect 62600 11100 62700 11200
rect 36100 11200 36200 11300
rect 46600 11200 46800 11300
rect 54000 11200 54100 11300
rect 64400 11200 64500 11300
rect 75000 11200 75100 11300
rect 27700 11300 27900 11500
rect 33000 11300 33100 11500
rect 57000 11300 57200 11500
rect 35900 11500 36100 11600
rect 40900 12000 41100 12200
rect 43800 12000 44000 12200
rect 23300 20200 23400 20400
rect 86800 23000 86900 23100
rect 86900 23100 87000 23300
rect 87200 23800 87300 24000
rect 46100 24500 46200 24700
rect 13600 25000 13700 25100
rect 47000 25100 47200 25200
rect 86900 25100 87000 25200
rect 47200 25200 47300 25400
rect 14000 25400 14100 25500
rect 47600 25500 47700 25600
rect 48100 26200 48300 26300
rect 48400 26600 48600 26800
rect 87200 29700 87300 29800
rect 86900 30400 87000 30500
rect 86800 30500 86900 30600
rect 13700 33600 13800 33700
rect 72900 34800 73000 35000
rect 48600 35000 48700 35100
rect 48300 35400 48400 35500
rect 73300 35400 73400 35500
rect 26900 35800 27000 35900
rect 73600 35800 73700 35900
rect 47600 36300 47700 36500
rect 47500 36500 47600 36600
rect 78000 38400 78100 38600
rect 86600 38700 86800 38800
rect 86800 38800 86900 39000
rect 86900 39000 87000 39100
rect 26600 43700 26800 43800
rect 13700 44100 13800 44300
rect 86900 44100 87000 44300
rect 72600 45600 72700 45800
rect 86900 46200 87000 46300
rect 71500 46300 71600 46500
rect 86800 46300 86900 46500
rect 71300 46500 71500 46600
rect 29500 46600 29700 46800
rect 70200 46800 70400 46900
rect 29800 48600 30000 48700
rect 87200 50100 87300 50200
rect 87200 50800 87300 50900
rect 87000 51100 87200 51200
rect 86900 51300 87000 51500
rect 26600 51600 26800 51800
rect 70600 57700 70800 57900
rect 72900 59000 73000 59100
rect 86800 59800 86900 60000
rect 13700 60000 13800 60100
rect 73600 60000 73700 60100
rect 52700 60400 52900 60500
rect 86900 61900 87000 62000
rect 14000 62200 14100 62300
rect 86600 65000 86800 65100
rect 86900 65200 87000 65400
rect 87200 65900 87300 66100
rect 14000 67500 14100 67600
rect 26600 67900 26800 68000
rect 72600 69800 72700 70000
rect 14100 70100 14300 70200
rect 71500 70500 71600 70600
rect 13600 70600 13700 70800
rect 29500 70800 29700 70900
rect 70200 70900 70400 71100
rect 86800 72600 86900 72700
rect 51600 84000 51800 84100
rect 70000 84000 70100 84100
rect 75200 84000 75400 84100
rect 35900 84100 36100 84300
rect 25500 84300 25600 84400
rect 33000 84300 33100 84400
rect 57000 84300 57200 84400
rect 27600 84400 27700 84500
rect 32900 84400 33000 84500
rect 48700 84400 48800 84500
rect 25800 84500 25900 84700
rect 38000 84500 38100 84700
rect 64300 84500 64400 84700
rect 67900 84500 68000 84700
<< metal2 >>
rect 27500 11100 27600 11200
rect 53700 11100 53800 11200
rect 67900 11100 68000 11200
rect 32900 11200 33000 11300
rect 41300 11200 41500 11300
rect 48700 11200 48800 11300
rect 51900 11200 52000 11300
rect 59300 11200 59400 11300
rect 22900 20500 23000 20600
rect 86800 25200 86900 25400
rect 48700 27300 48800 27500
rect 86800 28300 86900 28400
rect 86900 33700 87000 33800
rect 13700 35600 13800 35800
rect 13800 35800 14000 35900
rect 26600 36500 26800 36600
rect 26500 36800 26600 36900
rect 86600 44000 86800 44100
rect 27000 44700 27200 44800
rect 27500 45200 27600 45400
rect 28000 45800 28100 45900
rect 28300 46100 28400 46200
rect 14300 46500 14400 46600
rect 70900 46600 71100 46800
rect 86800 51500 86900 51600
rect 13800 54500 14000 54700
rect 13700 54700 13800 54800
rect 86600 56900 86800 57000
rect 51500 57700 51600 57900
rect 73700 60200 73800 60400
rect 13800 65100 14000 65200
rect 86800 65100 86900 65200
rect 27000 68800 27200 69000
rect 28000 70000 28100 70100
rect 28300 70200 28400 70400
rect 86800 70400 86900 70500
rect 77300 75400 77500 75500
rect 43700 83700 43800 83800
rect 62200 84000 62300 84100
rect 36200 84400 36300 84500
rect 62500 84400 62600 84500
rect 32700 84500 32900 84700
rect 52000 84500 52200 84700
rect 59000 84500 59100 84700
<< metal3 >>
rect 31100 11100 31200 11200
rect 43400 11200 43600 11300
rect 69700 11200 69800 11300
rect 62300 11300 62500 11500
rect 30600 11500 30800 11600
rect 54100 11500 54300 11600
rect 25400 11600 25500 11800
rect 23000 20400 23100 20500
rect 13600 23400 13700 23600
rect 45500 24400 45600 24500
rect 86900 28400 87000 28600
rect 44500 28700 44700 28800
rect 56100 28700 56200 28800
rect 13600 30100 13700 30200
rect 14100 30600 14300 30800
rect 86500 30600 86600 30800
rect 27500 35000 27600 35100
rect 47700 36200 47900 36300
rect 69500 37900 69700 38000
rect 26300 42300 26500 42500
rect 26800 44100 26900 44300
rect 27200 45000 27300 45100
rect 27600 45400 27700 45500
rect 27700 45500 27900 45600
rect 87000 45800 87200 45900
rect 13600 45900 13700 46100
rect 86900 49500 87000 49700
rect 27600 49800 27700 50000
rect 26500 51800 26600 51900
rect 56100 52900 56200 53000
rect 86900 54700 87000 54800
rect 87000 61600 87200 61800
rect 13800 62000 14000 62200
rect 69500 62000 69700 62200
rect 26300 66500 26500 66600
rect 26800 68300 26900 68400
rect 27200 69100 27300 69300
rect 27600 69500 27700 69700
rect 27700 69700 27900 69800
rect 86900 70500 87000 70600
rect 70900 70800 71100 70900
rect 86500 72700 86600 72900
rect 64700 84000 64800 84100
rect 36100 84300 36200 84400
rect 62300 84300 62500 84400
rect 31100 84500 31200 84700
rect 62600 84500 62700 84700
<< metal4 >>
rect 48400 11100 48600 11200
rect 57200 11200 57300 11300
rect 72900 11200 73000 11300
rect 77200 20200 77300 20400
rect 86800 33600 86900 33700
rect 52500 35900 52600 36100
rect 52600 36100 52700 36200
rect 73700 44100 73800 44300
rect 27300 45100 27500 45200
rect 72700 45500 72900 45600
rect 28100 45900 28300 46100
rect 28100 49400 28300 49500
rect 86600 51600 86800 51800
rect 52500 60100 52600 60200
rect 73700 68300 73800 68400
rect 73300 69100 73400 69300
rect 72700 69700 72900 69800
rect 28100 70100 28300 70200
rect 59400 84000 59500 84100
rect 27700 84300 27900 84400
rect 74800 84400 75000 84500
rect 53700 84500 53800 84700
rect -600 0 -500 100000
rect 100500 0 100600 100000
<< metal5 >>
rect 26100 10900 27300 11100
rect 31300 10900 32600 11100
rect 36600 10900 37700 11100
rect 41900 10900 43000 11100
rect 47200 10900 48300 11100
rect 52300 10900 53600 11100
rect 57700 10900 58700 11100
rect 63000 10900 64000 11100
rect 68100 10900 69300 11100
rect 73400 10900 74500 11100
rect 25900 11100 27500 11200
rect 31200 11100 32700 11200
rect 36300 11100 38000 11200
rect 41600 11100 43300 11200
rect 46900 11100 48400 11200
rect 52200 11100 53700 11200
rect 57500 11100 59000 11200
rect 62700 11100 64300 11200
rect 68000 11100 69500 11200
rect 73100 11100 74800 11200
rect 25600 11200 27700 11300
rect 30900 11200 32900 11300
rect 36200 11200 38300 11300
rect 41500 11200 43400 11300
rect 46800 11200 48700 11300
rect 52000 11200 54000 11300
rect 57300 11200 59300 11300
rect 62500 11200 64400 11300
rect 67700 11200 69700 11300
rect 73000 11200 75000 11300
rect 25500 11300 27700 11500
rect 30800 11300 33000 11500
rect 36100 11300 38300 11500
rect 41300 11300 43600 11500
rect 46600 11300 48800 11500
rect 51900 11300 54100 11500
rect 57200 11300 59400 11500
rect 62500 11300 64500 11500
rect 67600 11300 69800 11500
rect 72900 11300 75100 11500
rect 25500 11500 27900 11600
rect 30800 11500 33100 11600
rect 36100 11500 38400 11600
rect 41200 11500 43700 11600
rect 46500 11500 49000 11600
rect 51800 11500 54100 11600
rect 57000 11500 59400 11600
rect 62300 11500 64700 11600
rect 67600 11500 70000 11600
rect 72700 11500 75200 11600
rect 25500 11600 28000 11800
rect 30600 11600 33300 11800
rect 35900 11600 38600 11800
rect 41200 11600 43700 11800
rect 46300 11600 49000 11800
rect 51600 11600 54300 11800
rect 56900 11600 59500 11800
rect 62200 11600 64800 11800
rect 67500 11600 70100 11800
rect 72700 11600 75400 11800
rect 25400 11800 28100 11900
rect 30600 11800 33300 11900
rect 35900 11800 38600 11900
rect 41200 11800 43700 11900
rect 46300 11800 49000 11900
rect 51600 11800 54300 11900
rect 56900 11800 59700 11900
rect 62200 11800 64800 11900
rect 67300 11800 70100 11900
rect 72700 11800 75400 11900
rect 25400 11900 28100 12000
rect 30600 11900 33300 12000
rect 35900 11900 38600 12000
rect 41100 11900 43800 12000
rect 46300 11900 49000 12000
rect 51600 11900 54300 12000
rect 56900 11900 59700 12000
rect 62200 11900 64800 12000
rect 67300 11900 70100 12000
rect 72700 11900 75400 12000
rect 25400 12000 28100 12200
rect 30600 12000 33400 12200
rect 35900 12000 38600 12200
rect 41100 12000 43800 12200
rect 46300 12000 49100 12200
rect 51500 12000 54300 12200
rect 56900 12000 59700 12200
rect 62200 12000 65000 12200
rect 67300 12000 70100 12200
rect 72700 12000 75500 12200
rect 25400 12200 28100 12300
rect 30600 12200 33400 12300
rect 35900 12200 38600 12300
rect 40900 12200 44000 12300
rect 46300 12200 49100 12300
rect 51500 12200 54300 12300
rect 56900 12200 59700 12300
rect 62000 12200 65000 12300
rect 67300 12200 70100 12300
rect 72700 12200 75500 12300
rect 25400 12300 28100 12500
rect 30600 12300 33400 12500
rect 35900 12300 38700 12500
rect 40900 12300 44000 12500
rect 46300 12300 49100 12500
rect 51500 12300 54300 12500
rect 56900 12300 59700 12500
rect 62000 12300 65000 12500
rect 67300 12300 70100 12500
rect 72700 12300 75500 12500
rect 25400 12500 28100 12600
rect 30600 12500 33400 12600
rect 35900 12500 38700 12600
rect 40900 12500 44000 12600
rect 46200 12500 49100 12600
rect 51500 12500 54300 12600
rect 56900 12500 59700 12600
rect 62000 12500 65000 12600
rect 67300 12500 70100 12600
rect 72700 12500 75500 12600
rect 25400 12600 28100 12700
rect 30600 12600 33400 12700
rect 35900 12600 38700 12700
rect 40900 12600 44000 12700
rect 46200 12600 49100 12700
rect 51500 12600 54400 12700
rect 56900 12600 59700 12700
rect 62000 12600 65000 12700
rect 67300 12600 70200 12700
rect 72700 12600 75500 12700
rect 25400 12700 28100 12900
rect 30600 12700 33400 12900
rect 35900 12700 38700 12900
rect 40900 12700 44000 12900
rect 46200 12700 49100 12900
rect 51500 12700 54400 12900
rect 56900 12700 59700 12900
rect 62000 12700 65000 12900
rect 67300 12700 70200 12900
rect 72700 12700 75500 12900
rect 25400 12900 28100 13000
rect 30600 12900 33400 13000
rect 35900 12900 38700 13000
rect 40900 12900 44000 13000
rect 46200 12900 49100 13000
rect 51500 12900 54400 13000
rect 56900 12900 59700 13000
rect 62000 12900 65000 13000
rect 67300 12900 70200 13000
rect 72700 12900 75500 13000
rect 25400 13000 28100 13100
rect 30600 13000 33400 13100
rect 35900 13000 38700 13100
rect 40900 13000 44000 13100
rect 46200 13000 49100 13100
rect 51500 13000 54400 13100
rect 56900 13000 59700 13100
rect 62000 13000 65000 13100
rect 67300 13000 70200 13100
rect 72700 13000 75500 13100
rect 25400 13100 28100 13300
rect 30600 13100 33400 13300
rect 35900 13100 38700 13300
rect 40900 13100 44000 13300
rect 46200 13100 49100 13300
rect 51500 13100 54400 13300
rect 56900 13100 59700 13300
rect 62000 13100 65000 13300
rect 67300 13100 70200 13300
rect 72700 13100 75500 13300
rect 25400 13300 28100 13400
rect 30500 13300 33400 13400
rect 35900 13300 38700 13400
rect 40900 13300 44000 13400
rect 46200 13300 49100 13400
rect 51500 13300 54400 13400
rect 56800 13300 59700 13400
rect 62000 13300 65000 13400
rect 67300 13300 70200 13400
rect 72600 13300 75500 13400
rect 25400 13400 28100 13600
rect 30500 13400 33400 13600
rect 35900 13400 38700 13600
rect 40900 13400 44000 13600
rect 46200 13400 49100 13600
rect 51500 13400 54400 13600
rect 56800 13400 59700 13600
rect 62000 13400 65000 13600
rect 67300 13400 70200 13600
rect 72600 13400 75500 13600
rect 25400 13600 28100 13700
rect 30500 13600 33400 13700
rect 35900 13600 38700 13700
rect 40900 13600 44000 13700
rect 46200 13600 49100 13700
rect 51500 13600 54400 13700
rect 56800 13600 59700 13700
rect 62000 13600 65000 13700
rect 67300 13600 70200 13700
rect 72600 13600 75500 13700
rect 25400 13700 28100 13800
rect 30500 13700 33400 13800
rect 35900 13700 38700 13800
rect 40900 13700 44000 13800
rect 46200 13700 49100 13800
rect 51500 13700 54400 13800
rect 56800 13700 59700 13800
rect 62000 13700 65000 13800
rect 67300 13700 70200 13800
rect 72600 13700 75500 13800
rect 25400 13800 28100 14000
rect 30500 13800 33400 14000
rect 35900 13800 38700 14000
rect 40900 13800 44000 14000
rect 46200 13800 49100 14000
rect 51500 13800 54400 14000
rect 56800 13800 59700 14000
rect 62000 13800 65000 14000
rect 67300 13800 70200 14000
rect 72600 13800 75500 14000
rect 25400 14000 28100 14100
rect 30500 14000 33400 14100
rect 35900 14000 38700 14100
rect 40900 14000 44000 14100
rect 46200 14000 49100 14100
rect 51500 14000 54400 14100
rect 56800 14000 59700 14100
rect 62000 14000 65000 14100
rect 67300 14000 70200 14100
rect 72600 14000 75500 14100
rect 25400 14100 28100 14300
rect 30500 14100 33400 14300
rect 35900 14100 38700 14300
rect 40900 14100 44000 14300
rect 46200 14100 49100 14300
rect 51500 14100 54400 14300
rect 56800 14100 59700 14300
rect 62000 14100 65000 14300
rect 67300 14100 70200 14300
rect 72600 14100 75500 14300
rect 25400 14300 28100 14400
rect 30500 14300 33400 14400
rect 35900 14300 38700 14400
rect 40900 14300 44000 14400
rect 46200 14300 49100 14400
rect 51500 14300 54400 14400
rect 56800 14300 59700 14400
rect 62000 14300 65000 14400
rect 67300 14300 70200 14400
rect 72600 14300 75500 14400
rect 25400 14400 28100 14500
rect 30500 14400 33400 14500
rect 35900 14400 38700 14500
rect 40900 14400 44000 14500
rect 46200 14400 49100 14500
rect 51500 14400 54400 14500
rect 56800 14400 59700 14500
rect 62000 14400 65000 14500
rect 67300 14400 70200 14500
rect 72600 14400 75500 14500
rect 25400 14500 28100 14700
rect 30500 14500 33400 14700
rect 35900 14500 38700 14700
rect 40900 14500 44000 14700
rect 46200 14500 49100 14700
rect 51500 14500 54400 14700
rect 56800 14500 59700 14700
rect 62000 14500 65000 14700
rect 67300 14500 70200 14700
rect 72600 14500 75500 14700
rect 25400 14700 28100 14800
rect 30500 14700 33400 14800
rect 35900 14700 38700 14800
rect 40900 14700 44000 14800
rect 46200 14700 49100 14800
rect 51500 14700 54400 14800
rect 56800 14700 59700 14800
rect 62000 14700 65000 14800
rect 67300 14700 70200 14800
rect 72600 14700 75500 14800
rect 25400 14800 28100 15000
rect 30500 14800 33400 15000
rect 35900 14800 38700 15000
rect 40900 14800 44000 15000
rect 46200 14800 49100 15000
rect 51500 14800 54400 15000
rect 56800 14800 59700 15000
rect 62000 14800 65000 15000
rect 67300 14800 70200 15000
rect 72600 14800 75500 15000
rect 25400 15000 28100 15100
rect 30500 15000 33400 15100
rect 35900 15000 38700 15100
rect 40900 15000 44000 15100
rect 46200 15000 49100 15100
rect 51500 15000 54400 15100
rect 56800 15000 59700 15100
rect 62000 15000 65000 15100
rect 67300 15000 70200 15100
rect 72600 15000 75500 15100
rect 25400 15100 28100 15200
rect 30500 15100 33400 15200
rect 35900 15100 38700 15200
rect 40900 15100 44000 15200
rect 46200 15100 49100 15200
rect 51500 15100 54400 15200
rect 56800 15100 59700 15200
rect 62000 15100 65000 15200
rect 67300 15100 70200 15200
rect 72600 15100 75500 15200
rect 25400 15200 28100 15400
rect 30500 15200 33400 15400
rect 35900 15200 38700 15400
rect 40900 15200 44000 15400
rect 46200 15200 49100 15400
rect 51500 15200 54400 15400
rect 56800 15200 59700 15400
rect 62000 15200 65000 15400
rect 67300 15200 70200 15400
rect 72600 15200 75500 15400
rect 25400 15400 28100 15500
rect 30500 15400 33400 15500
rect 35900 15400 38700 15500
rect 40900 15400 44000 15500
rect 46200 15400 49100 15500
rect 51500 15400 54400 15500
rect 56800 15400 59700 15500
rect 62000 15400 65000 15500
rect 67300 15400 70200 15500
rect 72600 15400 75500 15500
rect 25400 15500 28100 15600
rect 30500 15500 33400 15600
rect 35900 15500 38700 15600
rect 40900 15500 44000 15600
rect 46200 15500 49100 15600
rect 51500 15500 54400 15600
rect 56800 15500 59700 15600
rect 62000 15500 65000 15600
rect 67300 15500 70200 15600
rect 72600 15500 75500 15600
rect 25400 15600 28100 15800
rect 30500 15600 33400 15800
rect 35900 15600 38700 15800
rect 40900 15600 44000 15800
rect 46200 15600 49100 15800
rect 51500 15600 54400 15800
rect 56800 15600 59700 15800
rect 62000 15600 65000 15800
rect 67300 15600 70200 15800
rect 72600 15600 75500 15800
rect 25400 15800 28100 15900
rect 30500 15800 33400 15900
rect 35900 15800 38700 15900
rect 40900 15800 44000 15900
rect 46200 15800 49100 15900
rect 51500 15800 54400 15900
rect 56800 15800 59700 15900
rect 62000 15800 65000 15900
rect 67300 15800 70200 15900
rect 72600 15800 75500 15900
rect 25400 15900 28100 16100
rect 30500 15900 33400 16100
rect 35900 15900 38700 16100
rect 40900 15900 44000 16100
rect 46200 15900 49100 16100
rect 51500 15900 54400 16100
rect 56800 15900 59700 16100
rect 62000 15900 65000 16100
rect 67300 15900 70200 16100
rect 72600 15900 75500 16100
rect 25400 16100 28100 16200
rect 30500 16100 33400 16200
rect 35900 16100 38700 16200
rect 40900 16100 44000 16200
rect 46200 16100 49100 16200
rect 51500 16100 54400 16200
rect 56800 16100 59700 16200
rect 62000 16100 65000 16200
rect 67300 16100 70200 16200
rect 72600 16100 75500 16200
rect 25200 16200 28100 16300
rect 30500 16200 33400 16300
rect 35900 16200 38700 16300
rect 40900 16200 44000 16300
rect 46200 16200 49100 16300
rect 51500 16200 54400 16300
rect 56800 16200 59700 16300
rect 62000 16200 65000 16300
rect 67300 16200 70200 16300
rect 72600 16200 75500 16300
rect 25200 16300 28100 16500
rect 30500 16300 33400 16500
rect 35900 16300 38700 16500
rect 40900 16300 44000 16500
rect 46200 16300 49100 16500
rect 51500 16300 54400 16500
rect 56800 16300 59700 16500
rect 62000 16300 65000 16500
rect 67300 16300 70200 16500
rect 72600 16300 75500 16500
rect 25200 16500 28100 16600
rect 30500 16500 33400 16600
rect 35900 16500 38700 16600
rect 40900 16500 44000 16600
rect 46200 16500 49100 16600
rect 51500 16500 54400 16600
rect 56800 16500 59700 16600
rect 62000 16500 65000 16600
rect 67300 16500 70200 16600
rect 72600 16500 75500 16600
rect 25200 16600 28100 16800
rect 30500 16600 33400 16800
rect 35900 16600 38700 16800
rect 40900 16600 44000 16800
rect 46200 16600 49100 16800
rect 51500 16600 54400 16800
rect 56800 16600 59700 16800
rect 62000 16600 65000 16800
rect 67300 16600 70200 16800
rect 72600 16600 75500 16800
rect 25200 16800 28100 16900
rect 30500 16800 33400 16900
rect 35900 16800 38700 16900
rect 40900 16800 44000 16900
rect 46200 16800 49100 16900
rect 51500 16800 54400 16900
rect 56800 16800 59700 16900
rect 62000 16800 65000 16900
rect 67300 16800 70200 16900
rect 72600 16800 75500 16900
rect 25200 16900 28100 17000
rect 30500 16900 33400 17000
rect 35900 16900 38700 17000
rect 40900 16900 44000 17000
rect 46200 16900 49100 17000
rect 51500 16900 54400 17000
rect 56800 16900 59700 17000
rect 62000 16900 65000 17000
rect 67300 16900 70200 17000
rect 72600 16900 75500 17000
rect 25200 17000 28100 17200
rect 30500 17000 33400 17200
rect 35900 17000 38700 17200
rect 40900 17000 44000 17200
rect 46200 17000 49100 17200
rect 51500 17000 54400 17200
rect 56800 17000 59700 17200
rect 62000 17000 65000 17200
rect 67300 17000 70200 17200
rect 72600 17000 75500 17200
rect 25200 17200 28100 17300
rect 30500 17200 33400 17300
rect 35900 17200 38700 17300
rect 40900 17200 44000 17300
rect 46200 17200 49100 17300
rect 51500 17200 54400 17300
rect 56800 17200 59700 17300
rect 62000 17200 65000 17300
rect 67300 17200 70200 17300
rect 72600 17200 75500 17300
rect 25200 17300 28100 17500
rect 30500 17300 33400 17500
rect 35900 17300 38700 17500
rect 40900 17300 44000 17500
rect 46200 17300 49100 17500
rect 51500 17300 54400 17500
rect 56800 17300 59700 17500
rect 62000 17300 65000 17500
rect 67300 17300 70200 17500
rect 72600 17300 75500 17500
rect 25200 17500 28100 17600
rect 30500 17500 33400 17600
rect 35900 17500 38700 17600
rect 40900 17500 44000 17600
rect 46200 17500 49100 17600
rect 51500 17500 54400 17600
rect 56800 17500 59700 17600
rect 62000 17500 65000 17600
rect 67300 17500 70200 17600
rect 72600 17500 75500 17600
rect 25200 17600 28100 17700
rect 30500 17600 33400 17700
rect 35900 17600 38700 17700
rect 40900 17600 44000 17700
rect 46200 17600 49100 17700
rect 51500 17600 54400 17700
rect 56800 17600 59700 17700
rect 62000 17600 65000 17700
rect 67300 17600 70200 17700
rect 72600 17600 75500 17700
rect 25200 17700 28100 17900
rect 30500 17700 33400 17900
rect 35900 17700 38700 17900
rect 40900 17700 44000 17900
rect 46200 17700 49100 17900
rect 51500 17700 54400 17900
rect 56800 17700 59700 17900
rect 62000 17700 65000 17900
rect 67300 17700 70200 17900
rect 72600 17700 75500 17900
rect 25200 17900 28100 18000
rect 30500 17900 33400 18000
rect 35900 17900 38700 18000
rect 40900 17900 44000 18000
rect 46200 17900 49100 18000
rect 51500 17900 54400 18000
rect 56800 17900 59700 18000
rect 62000 17900 65000 18000
rect 67300 17900 70200 18000
rect 72600 17900 75500 18000
rect 25200 18000 28100 18100
rect 30500 18000 33400 18100
rect 35900 18000 38700 18100
rect 40900 18000 44000 18100
rect 46200 18000 49100 18100
rect 51500 18000 54400 18100
rect 56800 18000 59700 18100
rect 62000 18000 65000 18100
rect 67300 18000 70200 18100
rect 72600 18000 75500 18100
rect 25200 18100 28100 18300
rect 30500 18100 33400 18300
rect 35900 18100 38700 18300
rect 40900 18100 44000 18300
rect 46200 18100 49100 18300
rect 51500 18100 54400 18300
rect 56800 18100 59700 18300
rect 62000 18100 65000 18300
rect 67300 18100 70200 18300
rect 72600 18100 75500 18300
rect 25200 18300 28100 18400
rect 30500 18300 33400 18400
rect 35900 18300 38700 18400
rect 40900 18300 44000 18400
rect 46200 18300 49100 18400
rect 51500 18300 54400 18400
rect 56800 18300 59700 18400
rect 62000 18300 65000 18400
rect 67300 18300 70200 18400
rect 72600 18300 75500 18400
rect 25200 18400 28100 18600
rect 30500 18400 33400 18600
rect 35900 18400 38700 18600
rect 40900 18400 44000 18600
rect 46200 18400 49100 18600
rect 51500 18400 54400 18600
rect 56800 18400 59700 18600
rect 62000 18400 65000 18600
rect 67300 18400 70200 18600
rect 72600 18400 75500 18600
rect 25200 18600 28100 18700
rect 30500 18600 33400 18700
rect 35900 18600 38700 18700
rect 40900 18600 44000 18700
rect 46200 18600 49100 18700
rect 51500 18600 54400 18700
rect 56800 18600 59700 18700
rect 62000 18600 65000 18700
rect 67300 18600 70200 18700
rect 72600 18600 75500 18700
rect 25200 18700 28100 18800
rect 30500 18700 33400 18800
rect 35900 18700 38700 18800
rect 40900 18700 44000 18800
rect 46200 18700 49100 18800
rect 51500 18700 54400 18800
rect 56800 18700 59700 18800
rect 62000 18700 65000 18800
rect 67300 18700 70200 18800
rect 72600 18700 75500 18800
rect 25200 18800 28100 19000
rect 30500 18800 33400 19000
rect 35900 18800 38700 19000
rect 40900 18800 44000 19000
rect 46200 18800 49100 19000
rect 51500 18800 54400 19000
rect 56800 18800 59700 19000
rect 62000 18800 65000 19000
rect 67300 18800 70200 19000
rect 72600 18800 75500 19000
rect 25200 19000 28100 19100
rect 30500 19000 33400 19100
rect 35900 19000 38700 19100
rect 40900 19000 44000 19100
rect 46200 19000 49100 19100
rect 51500 19000 54400 19100
rect 56800 19000 59700 19100
rect 62000 19000 65000 19100
rect 67300 19000 70200 19100
rect 72600 19000 75500 19100
rect 25200 19100 28100 19300
rect 30500 19100 33400 19300
rect 35900 19100 38700 19300
rect 40900 19100 44000 19300
rect 46200 19100 49100 19300
rect 51500 19100 54400 19300
rect 56800 19100 59700 19300
rect 62000 19100 65000 19300
rect 67300 19100 70200 19300
rect 72600 19100 75500 19300
rect 25200 19300 28100 19400
rect 30500 19300 33400 19400
rect 35900 19300 38700 19400
rect 40900 19300 44000 19400
rect 46200 19300 49100 19400
rect 51500 19300 54400 19400
rect 56800 19300 59700 19400
rect 62000 19300 65000 19400
rect 67300 19300 70200 19400
rect 72600 19300 75500 19400
rect 25200 19400 28100 19500
rect 30500 19400 33400 19500
rect 35900 19400 38700 19500
rect 40900 19400 44000 19500
rect 46200 19400 49100 19500
rect 51500 19400 54400 19500
rect 56800 19400 59700 19500
rect 62000 19400 65000 19500
rect 67300 19400 70200 19500
rect 72600 19400 75500 19500
rect 25200 19500 28100 19700
rect 30500 19500 33400 19700
rect 35900 19500 38700 19700
rect 40900 19500 44000 19700
rect 46200 19500 49100 19700
rect 51500 19500 54300 19700
rect 56800 19500 59700 19700
rect 62000 19500 65000 19700
rect 67300 19500 70200 19700
rect 72600 19500 75500 19700
rect 25200 19700 28100 19800
rect 30500 19700 33400 19800
rect 35900 19700 38700 19800
rect 40900 19700 44000 19800
rect 46200 19700 49100 19800
rect 51500 19700 54300 19800
rect 56800 19700 59700 19800
rect 62000 19700 65000 19800
rect 67300 19700 70100 19800
rect 72600 19700 75500 19800
rect 25200 19800 28100 20000
rect 30500 19800 33400 20000
rect 35900 19800 38700 20000
rect 40900 19800 44000 20000
rect 46200 19800 49100 20000
rect 51500 19800 54300 20000
rect 56800 19800 59700 20000
rect 62000 19800 65000 20000
rect 67300 19800 70100 20000
rect 72600 19800 75500 20000
rect 25200 20000 28100 20100
rect 30500 20000 33400 20100
rect 35900 20000 38700 20100
rect 40900 20000 44000 20100
rect 46200 20000 49100 20100
rect 51500 20000 54300 20100
rect 56800 20000 59700 20100
rect 62000 20000 65000 20100
rect 67300 20000 70100 20100
rect 72600 20000 75500 20100
rect 23800 20100 29300 20200
rect 29400 20100 34400 20200
rect 34700 20100 39700 20200
rect 40000 20100 45000 20200
rect 45200 20100 50200 20200
rect 50500 20100 55500 20200
rect 55800 20100 60600 20200
rect 61100 20100 65900 20200
rect 66200 20100 71200 20200
rect 71500 20100 76900 20200
rect 23400 20200 77200 20400
rect 23100 20400 77600 20500
rect 23000 20500 77700 20600
rect 22900 20600 77900 20800
rect 22700 20800 77900 20900
rect 22700 20900 78000 21100
rect 22700 21100 78000 21200
rect 22700 21200 78000 21300
rect 22600 21300 78100 21500
rect 22600 21500 78100 21600
rect 22600 21600 78100 21800
rect 22600 21800 78100 21900
rect 22600 21900 78100 22000
rect 22600 22000 78100 22200
rect 22600 22200 78100 22300
rect 22600 22300 78100 22500
rect 22600 22500 78100 22600
rect 22600 22600 78100 22700
rect 14300 22700 86500 22900
rect 14100 22900 86600 23000
rect 13800 23000 86800 23100
rect 13700 23100 86900 23300
rect 13700 23300 87000 23400
rect 13700 23400 87000 23600
rect 13600 23600 87200 23700
rect 13400 23700 87200 23800
rect 13400 23800 87200 24000
rect 13400 24000 87300 24100
rect 13400 24100 87300 24300
rect 13400 24300 34400 24400
rect 37600 24300 60900 24400
rect 64800 24300 87300 24400
rect 13400 24400 26500 24500
rect 45600 24400 51500 24500
rect 74100 24400 87300 24500
rect 13400 24500 26500 24700
rect 46200 24500 51500 24700
rect 74100 24500 87300 24700
rect 13600 24700 26500 24800
rect 46300 24700 51500 24800
rect 74100 24700 87200 24800
rect 13600 24800 26500 25000
rect 46600 24800 51500 25000
rect 74100 24800 87200 25000
rect 13700 25000 26500 25100
rect 46900 25000 51500 25100
rect 74100 25000 87000 25100
rect 13700 25100 26500 25200
rect 47200 25100 51500 25200
rect 74100 25100 86900 25200
rect 13800 25200 26500 25400
rect 47300 25200 51500 25400
rect 74100 25200 86800 25400
rect 14100 25400 26500 25500
rect 47500 25400 51500 25500
rect 74100 25400 86600 25500
rect 15800 25500 26500 25600
rect 47700 25500 51500 25600
rect 74100 25500 85100 25600
rect 22600 25600 26500 25800
rect 47700 25600 51500 25800
rect 74100 25600 78100 25800
rect 22600 25800 26500 25900
rect 47900 25800 51500 25900
rect 74100 25800 78100 25900
rect 22600 25900 26500 26100
rect 48000 25900 51500 26100
rect 74100 25900 78100 26100
rect 22600 26100 26500 26200
rect 48100 26100 51500 26200
rect 74100 26100 78100 26200
rect 22600 26200 26500 26300
rect 48300 26200 51500 26300
rect 74100 26200 78100 26300
rect 22600 26300 26500 26500
rect 48300 26300 51500 26500
rect 74100 26300 78100 26500
rect 22700 26500 26500 26600
rect 48400 26500 51500 26600
rect 74300 26500 78100 26600
rect 22700 26600 26500 26800
rect 48600 26600 51500 26800
rect 74100 26600 78100 26800
rect 22700 26800 26500 26900
rect 48600 26800 51500 26900
rect 74100 26800 78100 26900
rect 22700 26900 26500 27000
rect 48700 26900 51500 27000
rect 74100 26900 78100 27000
rect 22600 27000 26500 27200
rect 48700 27000 51500 27200
rect 74100 27000 78100 27200
rect 22600 27200 26500 27300
rect 48700 27200 51500 27300
rect 74100 27200 78100 27300
rect 22600 27300 26500 27500
rect 48800 27300 51500 27500
rect 74100 27300 78100 27500
rect 22600 27500 26500 27600
rect 48800 27500 51500 27600
rect 74100 27500 78100 27600
rect 22600 27600 26500 27700
rect 48800 27600 51500 27700
rect 74100 27600 78100 27700
rect 22600 27700 26500 27900
rect 48800 27700 51500 27900
rect 74100 27700 78000 27900
rect 22600 27900 26500 28000
rect 48800 27900 51500 28000
rect 74100 27900 78000 28000
rect 15800 28000 26300 28100
rect 49000 28000 51500 28100
rect 74100 28000 85100 28100
rect 14100 28100 26300 28300
rect 49000 28100 51500 28300
rect 74100 28100 86600 28300
rect 13800 28300 26300 28400
rect 49000 28300 51500 28400
rect 74100 28300 86800 28400
rect 13700 28400 26300 28600
rect 49000 28400 51500 28600
rect 74100 28400 86900 28600
rect 13700 28600 35200 28700
rect 49000 28600 51500 28700
rect 65600 28600 87000 28700
rect 13600 28700 44500 28800
rect 49000 28700 51500 28800
rect 56200 28700 87200 28800
rect 13600 28800 44700 29000
rect 49000 28800 51500 29000
rect 56100 28800 87200 29000
rect 13400 29000 44700 29100
rect 49000 29000 51500 29100
rect 56100 29000 87300 29100
rect 13400 29100 44700 29300
rect 49000 29100 51500 29300
rect 56100 29100 87300 29300
rect 13400 29300 44700 29400
rect 49000 29300 51500 29400
rect 56100 29300 87300 29400
rect 13400 29400 44800 29500
rect 49000 29400 51500 29500
rect 55900 29400 87300 29500
rect 13400 29500 44800 29700
rect 49000 29500 51500 29700
rect 55900 29500 87300 29700
rect 13400 29700 44800 29800
rect 49100 29700 51500 29800
rect 55900 29700 87200 29800
rect 13400 29800 44800 30000
rect 49100 29800 51500 30000
rect 55900 29800 87200 30000
rect 13600 30000 44800 30100
rect 49100 30000 51500 30100
rect 55900 30000 87200 30100
rect 13700 30100 44800 30200
rect 49100 30100 51500 30200
rect 55900 30100 87000 30200
rect 13700 30200 44800 30400
rect 49100 30200 51500 30400
rect 55900 30200 87000 30400
rect 13700 30400 44800 30500
rect 49100 30400 51500 30500
rect 55900 30400 86900 30500
rect 13800 30500 44800 30600
rect 49100 30500 51500 30600
rect 55900 30500 86800 30600
rect 14300 30600 44800 30800
rect 49100 30600 51500 30800
rect 55900 30600 86500 30800
rect 18700 30800 44800 30900
rect 49100 30800 51500 30900
rect 55900 30800 82200 30900
rect 22600 30900 44800 31100
rect 49100 30900 51500 31100
rect 55900 30900 78100 31100
rect 22600 31100 44800 31200
rect 49100 31100 51500 31200
rect 55900 31100 78100 31200
rect 22600 31200 44800 31300
rect 49100 31200 51500 31300
rect 55900 31200 78100 31300
rect 22600 31300 44800 31500
rect 49100 31300 51500 31500
rect 55900 31300 78100 31500
rect 22600 31500 44800 31600
rect 49100 31500 51500 31600
rect 55900 31500 78100 31600
rect 22600 31600 44800 31800
rect 49100 31600 51500 31800
rect 55900 31600 78100 31800
rect 22600 31800 44800 31900
rect 49100 31800 51500 31900
rect 55900 31800 78100 31900
rect 22700 31900 44800 32000
rect 49100 31900 51500 32000
rect 55900 31900 78100 32000
rect 22700 32000 44800 32200
rect 49100 32000 51500 32200
rect 55900 32000 78100 32200
rect 22700 32200 44800 32300
rect 49100 32200 51500 32300
rect 55900 32200 78100 32300
rect 22600 32300 44800 32500
rect 49100 32300 51500 32500
rect 55900 32300 78100 32500
rect 22600 32500 44800 32600
rect 49100 32500 51500 32600
rect 55900 32500 78100 32600
rect 22600 32600 44800 32700
rect 49000 32600 51500 32700
rect 55900 32600 78100 32700
rect 22600 32700 44800 32900
rect 49000 32700 51500 32900
rect 55900 32700 78100 32900
rect 22600 32900 44700 33000
rect 49000 32900 51500 33000
rect 56100 32900 78100 33000
rect 22600 33000 44700 33100
rect 49000 33000 51500 33100
rect 56100 33000 78000 33100
rect 22600 33100 44700 33300
rect 49000 33100 51500 33300
rect 56100 33100 78000 33300
rect 14700 33300 44700 33400
rect 49000 33300 51500 33400
rect 56100 33300 86100 33400
rect 14000 33400 42000 33600
rect 49000 33400 51500 33600
rect 58800 33400 86600 33600
rect 13800 33600 29800 33700
rect 49000 33600 51600 33700
rect 70800 33600 86800 33700
rect 13700 33700 29400 33800
rect 49000 33700 51600 33800
rect 71300 33700 86900 33800
rect 13600 33800 29100 34000
rect 49000 33800 51600 34000
rect 71500 33800 87000 34000
rect 13600 34000 28800 34100
rect 48800 34000 51800 34100
rect 71800 34000 87200 34100
rect 13600 34100 28600 34300
rect 48800 34100 51800 34300
rect 72000 34100 87200 34300
rect 13400 34300 28400 34400
rect 48800 34300 51800 34400
rect 72300 34300 87300 34400
rect 13400 34400 28100 34500
rect 48800 34400 51800 34500
rect 72500 34400 87300 34500
rect 13400 34500 28000 34700
rect 48800 34500 51800 34700
rect 72600 34500 87300 34700
rect 13400 34700 27900 34800
rect 48700 34700 51900 34800
rect 72900 34700 87300 34800
rect 13400 34800 27600 35000
rect 48700 34800 51900 35000
rect 73000 34800 87300 35000
rect 13400 35000 27500 35100
rect 48700 35000 51900 35100
rect 73000 35000 87200 35100
rect 13400 35100 27500 35200
rect 48600 35100 52000 35200
rect 73100 35100 87200 35200
rect 13600 35200 27300 35400
rect 48400 35200 52000 35400
rect 73300 35200 87200 35400
rect 13600 35400 27300 35500
rect 48400 35400 52200 35500
rect 73400 35400 87000 35500
rect 13700 35500 27200 35600
rect 48300 35500 52300 35600
rect 73400 35500 87000 35600
rect 13800 35600 27000 35800
rect 48300 35600 52300 35800
rect 73600 35600 86900 35800
rect 14000 35800 26900 35900
rect 48100 35800 52500 35900
rect 73700 35800 86800 35900
rect 14100 35900 26900 36100
rect 48000 35900 52500 36100
rect 73700 35900 86500 36100
rect 14800 36100 26800 36200
rect 47900 36100 52600 36200
rect 73800 36100 85900 36200
rect 22600 36200 26800 36300
rect 47900 36200 52900 36300
rect 73800 36200 78100 36300
rect 22600 36300 26800 36500
rect 47700 36300 52900 36500
rect 73800 36300 78100 36500
rect 22600 36500 26600 36600
rect 47600 36500 53000 36600
rect 73800 36500 78100 36600
rect 22600 36600 26600 36800
rect 47300 36600 53300 36800
rect 74000 36600 78100 36800
rect 22600 36800 26500 36900
rect 47200 36800 53400 36900
rect 74000 36800 78100 36900
rect 22600 36900 26500 37000
rect 47000 36900 53600 37000
rect 74000 36900 78100 37000
rect 22600 37000 26500 37200
rect 46800 37000 53800 37200
rect 74100 37000 78100 37200
rect 22700 37200 26500 37300
rect 46500 37200 54100 37300
rect 74100 37200 78100 37300
rect 22700 37300 26500 37500
rect 46300 37300 54300 37500
rect 74100 37300 78100 37500
rect 22700 37500 26500 37600
rect 45900 37500 54700 37600
rect 74100 37500 78100 37600
rect 22600 37600 26500 37700
rect 45200 37600 55400 37700
rect 74100 37600 78100 37700
rect 22600 37700 26500 37900
rect 38400 37700 62300 37900
rect 74100 37700 78100 37900
rect 22600 37900 26500 38000
rect 30900 37900 69500 38000
rect 74100 37900 78100 38000
rect 22600 38000 26500 38100
rect 30900 38000 69700 38100
rect 74100 38000 78100 38100
rect 22600 38100 26500 38300
rect 30900 38100 69700 38300
rect 74100 38100 78000 38300
rect 22600 38300 26500 38400
rect 30800 38300 69700 38400
rect 74100 38300 78000 38400
rect 22600 38400 26500 38600
rect 30800 38400 69700 38600
rect 74100 38400 78000 38600
rect 14100 38600 26500 38700
rect 30800 38600 69800 38700
rect 74100 38600 86500 38700
rect 14000 38700 26500 38800
rect 30800 38700 69800 38800
rect 74100 38700 86600 38800
rect 13800 38800 26500 39000
rect 30800 38800 69800 39000
rect 74100 38800 86800 39000
rect 13700 39000 26500 39100
rect 30800 39000 69800 39100
rect 74100 39000 86900 39100
rect 13600 39100 26500 39300
rect 30800 39100 69800 39300
rect 74100 39100 87000 39300
rect 13600 39300 26500 39400
rect 30800 39300 69800 39400
rect 74100 39300 87200 39400
rect 13600 39400 26500 39500
rect 30800 39400 69800 39500
rect 74100 39400 87200 39500
rect 13400 39500 26500 39700
rect 30800 39500 69800 39700
rect 74100 39500 87300 39700
rect 13400 39700 26500 39800
rect 30800 39700 69800 39800
rect 74100 39700 87300 39800
rect 13400 39800 26500 40000
rect 30800 39800 69800 40000
rect 74100 39800 87300 40000
rect 13400 40000 26500 40100
rect 30800 40000 69800 40100
rect 74300 40000 87300 40100
rect 13400 40100 26500 40200
rect 30800 40100 69800 40200
rect 74300 40100 87300 40200
rect 13400 40200 26500 40400
rect 30800 40200 69800 40400
rect 74100 40200 87300 40400
rect 13400 40400 26500 40500
rect 30800 40400 69800 40500
rect 74100 40400 87200 40500
rect 13600 40500 26500 40600
rect 30800 40500 69800 40600
rect 74100 40500 87200 40600
rect 13600 40600 26500 40800
rect 30800 40600 69800 40800
rect 74100 40600 87000 40800
rect 13700 40800 26500 40900
rect 30800 40800 69800 40900
rect 74100 40800 87000 40900
rect 13800 40900 26500 41100
rect 30800 40900 69800 41100
rect 74100 40900 86900 41100
rect 14000 41100 26500 41200
rect 30800 41100 69800 41200
rect 74100 41100 86800 41200
rect 14300 41200 26500 41300
rect 30800 41200 69800 41300
rect 74100 41200 86500 41300
rect 15900 41300 26500 41500
rect 30800 41300 69800 41500
rect 74100 41300 85000 41500
rect 22600 41500 26500 41600
rect 30800 41500 69800 41600
rect 74100 41500 78100 41600
rect 22600 41600 26500 41800
rect 30800 41600 69800 41800
rect 74100 41600 78100 41800
rect 22600 41800 26300 41900
rect 30800 41800 69800 41900
rect 74100 41800 78100 41900
rect 22600 41900 26300 42000
rect 30800 41900 69800 42000
rect 74100 41900 78100 42000
rect 22600 42000 26300 42200
rect 30800 42000 69700 42200
rect 74100 42000 78100 42200
rect 22600 42200 26300 42300
rect 30800 42200 69700 42300
rect 74100 42200 78100 42300
rect 22700 42300 26300 42500
rect 30900 42300 69700 42500
rect 74100 42300 78100 42500
rect 22700 42500 26500 42600
rect 30900 42500 69700 42600
rect 74100 42500 78100 42600
rect 22700 42600 26500 42700
rect 34300 42600 66500 42700
rect 74100 42600 78100 42700
rect 22700 42700 26500 42900
rect 49000 42700 51500 42900
rect 74100 42700 78100 42900
rect 22600 42900 26500 43000
rect 49000 42900 51500 43000
rect 74100 42900 78100 43000
rect 22600 43000 26500 43100
rect 49000 43000 51500 43100
rect 74100 43000 78100 43100
rect 22600 43100 26500 43300
rect 49000 43100 51500 43300
rect 74000 43100 78100 43300
rect 22600 43300 26500 43400
rect 49000 43300 51500 43400
rect 74000 43300 78100 43400
rect 22600 43400 26500 43600
rect 49000 43400 51500 43600
rect 74000 43400 78100 43600
rect 22600 43600 26600 43700
rect 49100 43600 51500 43700
rect 74000 43600 78000 43700
rect 22600 43700 26600 43800
rect 49100 43700 51500 43800
rect 73800 43700 78000 43800
rect 15600 43800 26800 44000
rect 49100 43800 51500 44000
rect 73800 43800 85100 44000
rect 14000 44000 26800 44100
rect 49100 44000 51500 44100
rect 73800 44000 86600 44100
rect 13800 44100 26800 44300
rect 49100 44100 51500 44300
rect 73800 44100 86900 44300
rect 13700 44300 26900 44400
rect 49100 44300 51500 44400
rect 73700 44300 87000 44400
rect 13600 44400 26900 44500
rect 49100 44400 51500 44500
rect 73700 44400 87000 44500
rect 13600 44500 27000 44700
rect 49100 44500 51500 44700
rect 73600 44500 87200 44700
rect 13400 44700 27000 44800
rect 49100 44700 51500 44800
rect 73400 44700 87200 44800
rect 13400 44800 27200 45000
rect 49100 44800 51500 45000
rect 73400 44800 87300 45000
rect 13400 45000 27200 45100
rect 49100 45000 51500 45100
rect 73300 45000 87300 45100
rect 13400 45100 27300 45200
rect 49100 45100 51500 45200
rect 73100 45100 87300 45200
rect 13400 45200 27500 45400
rect 49100 45200 51500 45400
rect 73000 45200 87300 45400
rect 13400 45400 27600 45500
rect 49100 45400 51500 45500
rect 72900 45400 87300 45500
rect 13400 45500 27700 45600
rect 49100 45500 51500 45600
rect 72900 45500 87300 45600
rect 13600 45600 27900 45800
rect 49100 45600 51500 45800
rect 72700 45600 87200 45800
rect 13600 45800 28000 45900
rect 49100 45800 51500 45900
rect 72500 45800 87000 45900
rect 13700 45900 28100 46100
rect 49100 45900 51500 46100
rect 72300 45900 87000 46100
rect 13700 46100 28300 46200
rect 49000 46100 51500 46200
rect 72200 46100 87000 46200
rect 13800 46200 28700 46300
rect 49000 46200 51500 46300
rect 71900 46200 86900 46300
rect 14000 46300 29000 46500
rect 49000 46300 51500 46500
rect 71600 46300 86800 46500
rect 14400 46500 29300 46600
rect 49000 46500 51500 46600
rect 71500 46500 86500 46600
rect 14500 46600 29500 46800
rect 49000 46600 51500 46800
rect 71100 46600 86300 46800
rect 22600 46800 30200 46900
rect 49000 46800 51500 46900
rect 70400 46800 78100 46900
rect 22600 46900 78100 47000
rect 22600 47000 78100 47200
rect 22600 47200 78100 47300
rect 22600 47300 78100 47500
rect 22600 47500 78100 47600
rect 22700 47600 78100 47700
rect 22700 47700 78100 47900
rect 22700 47900 78100 48000
rect 22700 48000 78100 48100
rect 22600 48100 78100 48300
rect 22600 48300 78100 48400
rect 22600 48400 78100 48600
rect 22600 48600 29800 48700
rect 49000 48600 51500 48700
rect 74100 48600 78100 48700
rect 22600 48700 29400 48800
rect 49000 48700 51500 48800
rect 74100 48700 78000 48800
rect 22600 48800 29100 49000
rect 49000 48800 51500 49000
rect 74100 48800 78000 49000
rect 14500 49000 28800 49100
rect 49000 49000 51500 49100
rect 74100 49000 86200 49100
rect 14100 49100 28600 49300
rect 49000 49100 51500 49300
rect 74100 49100 86600 49300
rect 14000 49300 28400 49400
rect 49000 49300 51500 49400
rect 74100 49300 86800 49400
rect 13800 49400 28100 49500
rect 49100 49400 51500 49500
rect 74100 49400 86900 49500
rect 13700 49500 28000 49700
rect 49100 49500 51500 49700
rect 74100 49500 86900 49700
rect 13600 49700 27900 49800
rect 49100 49700 51500 49800
rect 74100 49700 87000 49800
rect 13600 49800 27600 50000
rect 49100 49800 51500 50000
rect 74100 49800 87200 50000
rect 13400 50000 27600 50100
rect 49100 50000 51500 50100
rect 74100 50000 87200 50100
rect 13400 50100 27500 50200
rect 49100 50100 51500 50200
rect 74100 50100 87200 50200
rect 13400 50200 27300 50400
rect 49100 50200 51500 50400
rect 74100 50200 87300 50400
rect 13400 50400 27300 50500
rect 49100 50400 51500 50500
rect 74100 50400 87300 50500
rect 13400 50500 27200 50600
rect 49100 50500 51500 50600
rect 74100 50500 87300 50600
rect 13400 50600 27000 50800
rect 49100 50600 51500 50800
rect 74300 50600 87300 50800
rect 13400 50800 27000 50900
rect 49100 50800 51500 50900
rect 74100 50800 87200 50900
rect 13400 50900 26900 51100
rect 49100 50900 51500 51100
rect 74100 50900 87200 51100
rect 13600 51100 26800 51200
rect 49100 51100 51500 51200
rect 74100 51100 87000 51200
rect 13600 51200 26800 51300
rect 49100 51200 51500 51300
rect 74100 51200 87000 51300
rect 13700 51300 26800 51500
rect 49100 51300 51500 51500
rect 74100 51300 86900 51500
rect 13800 51500 26800 51600
rect 49100 51500 51500 51600
rect 74100 51500 86800 51600
rect 14000 51600 26600 51800
rect 49100 51600 51500 51800
rect 74100 51600 86600 51800
rect 14300 51800 26500 51900
rect 49100 51800 51500 51900
rect 74100 51800 86500 51900
rect 15000 51900 26500 52000
rect 49000 51900 51500 52000
rect 74100 51900 85800 52000
rect 22600 52000 26500 52200
rect 49000 52000 51500 52200
rect 74100 52000 78100 52200
rect 22600 52200 26500 52300
rect 49000 52200 51500 52300
rect 74100 52200 78100 52300
rect 22600 52300 26500 52500
rect 49000 52300 51500 52500
rect 74100 52300 78100 52500
rect 22600 52500 26500 52600
rect 49000 52500 51500 52600
rect 74100 52500 78100 52600
rect 22600 52600 26500 52700
rect 49000 52600 51500 52700
rect 74100 52600 78100 52700
rect 22600 52700 26500 52900
rect 40500 52700 51500 52900
rect 65600 52700 78100 52900
rect 22700 52900 26500 53000
rect 30900 52900 51500 53000
rect 56200 52900 78100 53000
rect 22700 53000 26500 53100
rect 30900 53000 51500 53100
rect 56100 53000 78100 53100
rect 22700 53100 26500 53300
rect 30900 53100 51500 53300
rect 56100 53100 78100 53300
rect 22600 53300 26500 53400
rect 30900 53300 51500 53400
rect 56100 53300 78100 53400
rect 22600 53400 26500 53600
rect 30800 53400 51500 53600
rect 56100 53400 78100 53600
rect 22600 53600 26500 53700
rect 30800 53600 51500 53700
rect 55900 53600 78100 53700
rect 22600 53700 26500 53800
rect 30800 53700 51500 53800
rect 55900 53700 78100 53800
rect 22600 53800 26500 54000
rect 30800 53800 51500 54000
rect 55900 53800 78100 54000
rect 22600 54000 26500 54100
rect 30800 54000 51500 54100
rect 55900 54000 78000 54100
rect 22600 54100 26500 54300
rect 30800 54100 51500 54300
rect 55900 54100 78000 54300
rect 14400 54300 26500 54400
rect 30800 54300 51500 54400
rect 55900 54300 86300 54400
rect 14300 54400 26500 54500
rect 30800 54400 51500 54500
rect 55900 54400 86500 54500
rect 14000 54500 26500 54700
rect 30800 54500 51500 54700
rect 55900 54500 86800 54700
rect 13800 54700 26500 54800
rect 30800 54700 51500 54800
rect 55900 54700 86900 54800
rect 13700 54800 26500 55000
rect 30800 54800 51500 55000
rect 55900 54800 87000 55000
rect 13600 55000 26500 55100
rect 30800 55000 51500 55100
rect 55900 55000 87000 55100
rect 13600 55100 26500 55200
rect 30800 55100 51500 55200
rect 55900 55100 87200 55200
rect 13400 55200 26500 55400
rect 30800 55200 51500 55400
rect 55900 55200 87200 55400
rect 13400 55400 26500 55500
rect 30800 55400 51500 55500
rect 55900 55400 87300 55500
rect 13400 55500 26500 55600
rect 30800 55500 51500 55600
rect 55900 55500 87300 55600
rect 13400 55600 26500 55800
rect 30800 55600 51500 55800
rect 55900 55600 87300 55800
rect 13400 55800 26500 55900
rect 30800 55800 51500 55900
rect 55900 55800 87300 55900
rect 13400 55900 26500 56100
rect 30800 55900 51500 56100
rect 55900 55900 87300 56100
rect 13400 56100 26500 56200
rect 30800 56100 51500 56200
rect 55900 56100 87300 56200
rect 13400 56200 26500 56300
rect 30800 56200 51500 56300
rect 55900 56200 87200 56300
rect 13600 56300 26500 56500
rect 30800 56300 51500 56500
rect 55900 56300 87200 56500
rect 13600 56500 26500 56600
rect 30800 56500 51500 56600
rect 55900 56500 87000 56600
rect 13700 56600 26500 56800
rect 30800 56600 51500 56800
rect 55900 56600 87000 56800
rect 13800 56800 26500 56900
rect 30800 56800 51500 56900
rect 55900 56800 86900 56900
rect 14000 56900 26500 57000
rect 30800 56900 51500 57000
rect 55900 56900 86600 57000
rect 18700 57000 26500 57200
rect 30800 57000 51500 57200
rect 56100 57000 82200 57200
rect 22600 57200 26500 57300
rect 30800 57200 51500 57300
rect 56100 57200 78100 57300
rect 22600 57300 26500 57500
rect 30800 57300 51500 57500
rect 56100 57300 78100 57500
rect 22600 57500 26500 57600
rect 30800 57500 51500 57600
rect 56100 57500 78100 57600
rect 22600 57600 26500 57700
rect 30800 57600 51500 57700
rect 58800 57600 78100 57700
rect 22600 57700 26500 57900
rect 30800 57700 51500 57900
rect 70800 57700 78100 57900
rect 22600 57900 26500 58000
rect 30800 57900 51600 58000
rect 71300 57900 78100 58000
rect 22700 58000 26500 58100
rect 30800 58000 51600 58100
rect 71500 58000 78100 58100
rect 22700 58100 26500 58300
rect 30800 58100 51600 58300
rect 71800 58100 78100 58300
rect 22700 58300 26500 58400
rect 30800 58300 51800 58400
rect 72000 58300 78100 58400
rect 22700 58400 26500 58600
rect 30800 58400 51800 58600
rect 72300 58400 78100 58600
rect 22600 58600 26500 58700
rect 30800 58600 51800 58700
rect 72500 58600 78100 58700
rect 22600 58700 26500 58800
rect 30800 58700 51800 58800
rect 72600 58700 78100 58800
rect 22600 58800 26500 59000
rect 30800 58800 51900 59000
rect 72900 58800 78100 59000
rect 22600 59000 26500 59100
rect 30800 59000 51900 59100
rect 73000 59000 78100 59100
rect 22600 59100 26500 59300
rect 30800 59100 51900 59300
rect 73000 59100 78100 59300
rect 22600 59300 26500 59400
rect 30800 59300 52000 59400
rect 73100 59300 78000 59400
rect 22600 59400 26500 59500
rect 30800 59400 52000 59500
rect 73300 59400 78000 59500
rect 14800 59500 26500 59700
rect 30800 59500 52200 59700
rect 73300 59500 85900 59700
rect 14100 59700 26500 59800
rect 30800 59700 52300 59800
rect 73400 59700 86600 59800
rect 13800 59800 26500 60000
rect 30800 59800 52300 60000
rect 73600 59800 86800 60000
rect 13800 60000 26500 60100
rect 30800 60000 52500 60100
rect 73700 60000 87000 60100
rect 13700 60100 26500 60200
rect 30800 60100 52500 60200
rect 73700 60100 87000 60200
rect 13600 60200 26500 60400
rect 30800 60200 52700 60400
rect 73800 60200 87200 60400
rect 13600 60400 26500 60500
rect 30800 60400 52700 60500
rect 73800 60400 87200 60500
rect 13400 60500 26500 60600
rect 30800 60500 52900 60600
rect 73800 60500 87200 60600
rect 13400 60600 26500 60800
rect 30800 60600 53000 60800
rect 73800 60600 87300 60800
rect 13400 60800 26500 60900
rect 30800 60800 53300 60900
rect 74000 60800 87300 60900
rect 13400 60900 26500 61100
rect 30800 60900 53400 61100
rect 74000 60900 87300 61100
rect 13400 61100 26500 61200
rect 30800 61100 53600 61200
rect 74000 61100 87300 61200
rect 13400 61200 26500 61300
rect 30800 61200 53800 61300
rect 74100 61200 87300 61300
rect 13400 61300 26500 61500
rect 30800 61300 54100 61500
rect 74100 61300 87300 61500
rect 13600 61500 26500 61600
rect 30800 61500 54300 61600
rect 74100 61500 87200 61600
rect 13600 61600 26500 61800
rect 30800 61600 54700 61800
rect 74100 61600 87000 61800
rect 13600 61800 26500 61900
rect 30800 61800 55400 61900
rect 74100 61800 87000 61900
rect 13700 61900 26500 62000
rect 30800 61900 62300 62000
rect 74100 61900 86900 62000
rect 14000 62000 26500 62200
rect 30800 62000 69500 62200
rect 74100 62000 86800 62200
rect 14100 62200 26500 62300
rect 30800 62200 69700 62300
rect 74100 62200 86600 62300
rect 22600 62300 26500 62500
rect 30800 62300 69700 62500
rect 74100 62300 78100 62500
rect 22600 62500 26500 62600
rect 30800 62500 69700 62600
rect 74100 62500 78100 62600
rect 22600 62600 26500 62700
rect 30800 62600 69700 62700
rect 74100 62600 78100 62700
rect 22600 62700 26500 62900
rect 30800 62700 69800 62900
rect 74100 62700 78100 62900
rect 22600 62900 26500 63000
rect 30800 62900 69800 63000
rect 74100 62900 78100 63000
rect 22600 63000 26500 63100
rect 30800 63000 69800 63100
rect 74100 63000 78100 63100
rect 22600 63100 26500 63300
rect 30800 63100 69800 63300
rect 74100 63100 78100 63300
rect 22600 63300 26500 63400
rect 30800 63300 69800 63400
rect 74100 63300 78100 63400
rect 22700 63400 26500 63600
rect 30800 63400 69800 63600
rect 74100 63400 78100 63600
rect 22700 63600 26500 63700
rect 30800 63600 69800 63700
rect 74100 63600 78100 63700
rect 22700 63700 26500 63800
rect 30800 63700 69800 63800
rect 74100 63700 78100 63800
rect 22600 63800 26500 64000
rect 30800 63800 69800 64000
rect 74100 63800 78100 64000
rect 22600 64000 26500 64100
rect 30800 64000 69800 64100
rect 74100 64000 78100 64100
rect 22600 64100 26500 64300
rect 30800 64100 69800 64300
rect 74300 64100 78100 64300
rect 22600 64300 26300 64400
rect 30800 64300 69800 64400
rect 74300 64300 78100 64400
rect 22600 64400 26300 64500
rect 30800 64400 69800 64500
rect 74100 64400 78100 64500
rect 22600 64500 26300 64700
rect 30800 64500 69800 64700
rect 74100 64500 78000 64700
rect 22600 64700 26300 64800
rect 30800 64700 69800 64800
rect 74100 64700 78000 64800
rect 14300 64800 26300 65000
rect 30800 64800 69800 65000
rect 74100 64800 86300 65000
rect 14100 65000 26300 65100
rect 30800 65000 69800 65100
rect 74100 65000 86600 65100
rect 14000 65100 26300 65200
rect 30800 65100 69800 65200
rect 74100 65100 86800 65200
rect 13800 65200 26300 65400
rect 30800 65200 69800 65400
rect 74100 65200 86900 65400
rect 13700 65400 26300 65500
rect 30800 65400 69800 65500
rect 74100 65400 87000 65500
rect 13600 65500 26300 65600
rect 30800 65500 69800 65600
rect 74100 65500 87000 65600
rect 13600 65600 26300 65800
rect 30800 65600 69800 65800
rect 74100 65600 87200 65800
rect 13400 65800 26300 65900
rect 30800 65800 69800 65900
rect 74100 65800 87200 65900
rect 13400 65900 26300 66100
rect 30800 65900 69800 66100
rect 74100 65900 87200 66100
rect 13400 66100 26300 66200
rect 30800 66100 69800 66200
rect 74100 66100 87300 66200
rect 13400 66200 26300 66300
rect 30900 66200 69700 66300
rect 74100 66200 87300 66300
rect 13400 66300 26300 66500
rect 30900 66300 69700 66500
rect 74100 66300 87300 66500
rect 13400 66500 26300 66600
rect 30900 66500 69700 66600
rect 74100 66500 87300 66600
rect 13400 66600 26500 66800
rect 30900 66600 69700 66800
rect 74100 66600 87300 66800
rect 13600 66800 26500 66900
rect 34300 66800 66500 66900
rect 74100 66800 87200 66900
rect 13600 66900 26500 67000
rect 49000 66900 51500 67000
rect 74100 66900 87200 67000
rect 13700 67000 26500 67200
rect 49000 67000 51500 67200
rect 74100 67000 87000 67200
rect 13700 67200 26500 67300
rect 49000 67200 51500 67300
rect 74100 67200 86900 67300
rect 13800 67300 26500 67500
rect 49000 67300 51500 67500
rect 74000 67300 86800 67500
rect 14100 67500 26500 67600
rect 49000 67500 51500 67600
rect 74000 67500 86600 67600
rect 15800 67600 26500 67700
rect 49000 67600 51500 67700
rect 74000 67600 85100 67700
rect 22600 67700 26600 67900
rect 49100 67700 51500 67900
rect 74000 67700 78100 67900
rect 22600 67900 26600 68000
rect 49100 67900 51500 68000
rect 73800 67900 78100 68000
rect 22600 68000 26800 68100
rect 49100 68000 51500 68100
rect 73800 68000 78100 68100
rect 22600 68100 26800 68300
rect 49100 68100 51500 68300
rect 73800 68100 78100 68300
rect 22600 68300 26800 68400
rect 49100 68300 51500 68400
rect 73800 68300 78100 68400
rect 22600 68400 26900 68600
rect 49100 68400 51500 68600
rect 73700 68400 78100 68600
rect 22700 68600 26900 68700
rect 49100 68600 51500 68700
rect 73700 68600 78100 68700
rect 22700 68700 27000 68800
rect 49100 68700 51500 68800
rect 73600 68700 78100 68800
rect 22700 68800 27000 69000
rect 49100 68800 51500 69000
rect 73400 68800 78100 69000
rect 22700 69000 27200 69100
rect 49100 69000 51500 69100
rect 73400 69000 78100 69100
rect 22600 69100 27200 69300
rect 49100 69100 51500 69300
rect 73400 69100 78100 69300
rect 22600 69300 27500 69400
rect 49100 69300 51500 69400
rect 73300 69300 78100 69400
rect 22600 69400 27600 69500
rect 49100 69400 51500 69500
rect 73000 69400 78100 69500
rect 22600 69500 27600 69700
rect 49100 69500 51500 69700
rect 72900 69500 78100 69700
rect 22600 69700 27700 69800
rect 49100 69700 51500 69800
rect 72900 69700 78100 69800
rect 22600 69800 27900 70000
rect 49100 69800 51500 70000
rect 72700 69800 78000 70000
rect 22600 70000 28000 70100
rect 49100 70000 51500 70100
rect 72500 70000 78000 70100
rect 14300 70100 28100 70200
rect 49100 70100 51500 70200
rect 72300 70100 86500 70200
rect 14100 70200 28300 70400
rect 49000 70200 51500 70400
rect 72200 70200 86600 70400
rect 13800 70400 28700 70500
rect 49000 70400 51500 70500
rect 71900 70400 86800 70500
rect 13700 70500 29000 70600
rect 49000 70500 51500 70600
rect 71600 70500 86900 70600
rect 13700 70600 29300 70800
rect 49000 70600 51500 70800
rect 71500 70600 87000 70800
rect 13600 70800 29500 70900
rect 49000 70800 51500 70900
rect 71100 70800 87000 70900
rect 13600 70900 30200 71100
rect 49000 70900 51500 71100
rect 70400 70900 87200 71100
rect 13400 71100 35000 71200
rect 44700 71100 56200 71200
rect 65900 71100 87200 71200
rect 13400 71200 87300 71300
rect 13400 71300 87300 71500
rect 13400 71500 87300 71600
rect 13400 71600 87300 71800
rect 13400 71800 87300 71900
rect 13400 71900 87300 72000
rect 13600 72000 87200 72200
rect 13600 72200 87200 72300
rect 13700 72300 87000 72500
rect 13700 72500 86900 72600
rect 13800 72600 86800 72700
rect 14100 72700 86500 72900
rect 18700 72900 82200 73000
rect 22600 73000 78100 73100
rect 22600 73100 78100 73300
rect 22600 73300 78100 73400
rect 22600 73400 78100 73600
rect 22600 73600 78100 73700
rect 22600 73700 78100 73800
rect 22600 73800 78100 74000
rect 22600 74000 78100 74100
rect 22600 74100 78000 74300
rect 22600 74300 78000 74400
rect 22700 74400 78000 74500
rect 22700 74500 78000 74700
rect 22700 74700 77900 74800
rect 22700 74800 77900 75000
rect 22900 75000 77900 75100
rect 23000 75100 77700 75200
rect 23100 75200 77600 75400
rect 23300 75400 77300 75500
rect 23800 75500 29300 75600
rect 29500 75500 34400 75600
rect 34800 75500 39700 75600
rect 40000 75500 45000 75600
rect 45200 75500 50100 75600
rect 50500 75500 55400 75600
rect 55600 75500 60600 75600
rect 61100 75500 65900 75600
rect 66300 75500 71200 75600
rect 71500 75500 76900 75600
rect 25200 75600 28100 75800
rect 30500 75600 33400 75800
rect 35900 75600 38700 75800
rect 40900 75600 44000 75800
rect 46200 75600 49100 75800
rect 51500 75600 54400 75800
rect 56800 75600 59700 75800
rect 62000 75600 65000 75800
rect 67300 75600 70200 75800
rect 72600 75600 75500 75800
rect 25200 75800 28100 75900
rect 30500 75800 33400 75900
rect 35900 75800 38700 75900
rect 40900 75800 44000 75900
rect 46200 75800 49100 75900
rect 51500 75800 54400 75900
rect 56800 75800 59700 75900
rect 62000 75800 65000 75900
rect 67300 75800 70200 75900
rect 72600 75800 75500 75900
rect 25200 75900 28100 76100
rect 30500 75900 33400 76100
rect 35900 75900 38700 76100
rect 40900 75900 44000 76100
rect 46200 75900 49100 76100
rect 51500 75900 54400 76100
rect 56800 75900 59700 76100
rect 62000 75900 65000 76100
rect 67300 75900 70200 76100
rect 72600 75900 75500 76100
rect 25200 76100 28100 76200
rect 30500 76100 33400 76200
rect 35900 76100 38700 76200
rect 40900 76100 44000 76200
rect 46200 76100 49100 76200
rect 51500 76100 54400 76200
rect 56800 76100 59700 76200
rect 62000 76100 65000 76200
rect 67300 76100 70200 76200
rect 72600 76100 75500 76200
rect 25200 76200 28100 76300
rect 30500 76200 33400 76300
rect 35900 76200 38700 76300
rect 40900 76200 44000 76300
rect 46200 76200 49100 76300
rect 51500 76200 54400 76300
rect 56800 76200 59700 76300
rect 62000 76200 65000 76300
rect 67300 76200 70200 76300
rect 72600 76200 75500 76300
rect 25200 76300 28100 76500
rect 30500 76300 33400 76500
rect 35900 76300 38700 76500
rect 40900 76300 44000 76500
rect 46200 76300 49100 76500
rect 51500 76300 54400 76500
rect 56800 76300 59700 76500
rect 62000 76300 65000 76500
rect 67300 76300 70200 76500
rect 72600 76300 75500 76500
rect 25200 76500 28100 76600
rect 30500 76500 33400 76600
rect 35900 76500 38700 76600
rect 40900 76500 44000 76600
rect 46200 76500 49100 76600
rect 51500 76500 54400 76600
rect 56800 76500 59700 76600
rect 62000 76500 65000 76600
rect 67300 76500 70200 76600
rect 72600 76500 75500 76600
rect 25200 76600 28100 76800
rect 30500 76600 33400 76800
rect 35900 76600 38700 76800
rect 40900 76600 44000 76800
rect 46200 76600 49100 76800
rect 51500 76600 54400 76800
rect 56800 76600 59700 76800
rect 62000 76600 65000 76800
rect 67300 76600 70200 76800
rect 72600 76600 75500 76800
rect 25200 76800 28100 76900
rect 30500 76800 33400 76900
rect 35900 76800 38700 76900
rect 40900 76800 44000 76900
rect 46200 76800 49100 76900
rect 51500 76800 54400 76900
rect 56800 76800 59700 76900
rect 62000 76800 65000 76900
rect 67300 76800 70200 76900
rect 72600 76800 75500 76900
rect 25200 76900 28100 77000
rect 30500 76900 33400 77000
rect 35900 76900 38700 77000
rect 40900 76900 44000 77000
rect 46200 76900 49100 77000
rect 51500 76900 54400 77000
rect 56800 76900 59700 77000
rect 62000 76900 65000 77000
rect 67300 76900 70200 77000
rect 72600 76900 75500 77000
rect 25200 77000 28100 77200
rect 30500 77000 33400 77200
rect 35900 77000 38700 77200
rect 40900 77000 44000 77200
rect 46200 77000 49100 77200
rect 51500 77000 54400 77200
rect 56800 77000 59700 77200
rect 62000 77000 65000 77200
rect 67300 77000 70200 77200
rect 72600 77000 75500 77200
rect 25200 77200 28100 77300
rect 30500 77200 33400 77300
rect 35900 77200 38700 77300
rect 40900 77200 44000 77300
rect 46200 77200 49100 77300
rect 51500 77200 54400 77300
rect 56800 77200 59700 77300
rect 62000 77200 65000 77300
rect 67300 77200 70200 77300
rect 72600 77200 75500 77300
rect 25200 77300 28100 77500
rect 30500 77300 33400 77500
rect 35900 77300 38700 77500
rect 40900 77300 44000 77500
rect 46200 77300 49100 77500
rect 51500 77300 54400 77500
rect 56800 77300 59700 77500
rect 62000 77300 65000 77500
rect 67300 77300 70200 77500
rect 72600 77300 75500 77500
rect 25200 77500 28100 77600
rect 30500 77500 33400 77600
rect 35900 77500 38700 77600
rect 40900 77500 44000 77600
rect 46200 77500 49100 77600
rect 51500 77500 54400 77600
rect 56800 77500 59700 77600
rect 62000 77500 65000 77600
rect 67300 77500 70200 77600
rect 72600 77500 75500 77600
rect 25200 77600 28100 77700
rect 30500 77600 33400 77700
rect 35900 77600 38700 77700
rect 40900 77600 44000 77700
rect 46200 77600 49100 77700
rect 51500 77600 54400 77700
rect 56800 77600 59700 77700
rect 62000 77600 65000 77700
rect 67300 77600 70200 77700
rect 72600 77600 75500 77700
rect 25200 77700 28100 77900
rect 30500 77700 33400 77900
rect 35900 77700 38700 77900
rect 40900 77700 44000 77900
rect 46200 77700 49100 77900
rect 51500 77700 54400 77900
rect 56800 77700 59700 77900
rect 62000 77700 65000 77900
rect 67300 77700 70200 77900
rect 72600 77700 75500 77900
rect 25200 77900 28100 78000
rect 30500 77900 33400 78000
rect 35900 77900 38700 78000
rect 40900 77900 44000 78000
rect 46200 77900 49100 78000
rect 51500 77900 54400 78000
rect 56800 77900 59700 78000
rect 62000 77900 65000 78000
rect 67300 77900 70200 78000
rect 72600 77900 75500 78000
rect 25200 78000 28100 78100
rect 30500 78000 33400 78100
rect 35900 78000 38700 78100
rect 40900 78000 44000 78100
rect 46200 78000 49100 78100
rect 51500 78000 54400 78100
rect 56800 78000 59700 78100
rect 62000 78000 65000 78100
rect 67300 78000 70200 78100
rect 72600 78000 75500 78100
rect 25200 78100 28100 78300
rect 30500 78100 33400 78300
rect 35900 78100 38700 78300
rect 40900 78100 44000 78300
rect 46200 78100 49100 78300
rect 51500 78100 54400 78300
rect 56800 78100 59700 78300
rect 62000 78100 65000 78300
rect 67300 78100 70200 78300
rect 72600 78100 75500 78300
rect 25200 78300 28100 78400
rect 30500 78300 33400 78400
rect 35900 78300 38700 78400
rect 40900 78300 44000 78400
rect 46200 78300 49100 78400
rect 51500 78300 54400 78400
rect 56800 78300 59700 78400
rect 62000 78300 65000 78400
rect 67300 78300 70200 78400
rect 72600 78300 75500 78400
rect 25200 78400 28100 78600
rect 30500 78400 33400 78600
rect 35900 78400 38700 78600
rect 40900 78400 44000 78600
rect 46200 78400 49100 78600
rect 51500 78400 54400 78600
rect 56800 78400 59700 78600
rect 62000 78400 65000 78600
rect 67300 78400 70200 78600
rect 72600 78400 75500 78600
rect 25200 78600 28100 78700
rect 30500 78600 33400 78700
rect 35900 78600 38700 78700
rect 40900 78600 44000 78700
rect 46200 78600 49100 78700
rect 51500 78600 54400 78700
rect 56800 78600 59700 78700
rect 62000 78600 65000 78700
rect 67300 78600 70200 78700
rect 72600 78600 75500 78700
rect 25200 78700 28100 78800
rect 30500 78700 33400 78800
rect 35900 78700 38700 78800
rect 40900 78700 44000 78800
rect 46200 78700 49100 78800
rect 51500 78700 54400 78800
rect 56800 78700 59700 78800
rect 62000 78700 65000 78800
rect 67300 78700 70200 78800
rect 72600 78700 75500 78800
rect 25200 78800 28100 79000
rect 30500 78800 33400 79000
rect 35900 78800 38700 79000
rect 40900 78800 44000 79000
rect 46200 78800 49100 79000
rect 51500 78800 54400 79000
rect 56800 78800 59700 79000
rect 62000 78800 65000 79000
rect 67300 78800 70200 79000
rect 72600 78800 75500 79000
rect 25200 79000 28100 79100
rect 30500 79000 33400 79100
rect 35900 79000 38700 79100
rect 40900 79000 44000 79100
rect 46200 79000 49100 79100
rect 51500 79000 54400 79100
rect 56800 79000 59700 79100
rect 62000 79000 65000 79100
rect 67300 79000 70200 79100
rect 72600 79000 75500 79100
rect 25200 79100 28100 79300
rect 30500 79100 33400 79300
rect 35900 79100 38700 79300
rect 40900 79100 44000 79300
rect 46200 79100 49100 79300
rect 51500 79100 54400 79300
rect 56800 79100 59700 79300
rect 62000 79100 65000 79300
rect 67300 79100 70200 79300
rect 72600 79100 75500 79300
rect 25200 79300 28100 79400
rect 30500 79300 33400 79400
rect 35900 79300 38700 79400
rect 40900 79300 44000 79400
rect 46200 79300 49100 79400
rect 51500 79300 54400 79400
rect 56800 79300 59700 79400
rect 62000 79300 65000 79400
rect 67300 79300 70200 79400
rect 72600 79300 75500 79400
rect 25400 79400 28100 79500
rect 30500 79400 33400 79500
rect 35900 79400 38700 79500
rect 40900 79400 44000 79500
rect 46200 79400 49100 79500
rect 51500 79400 54400 79500
rect 56800 79400 59700 79500
rect 62000 79400 65000 79500
rect 67300 79400 70200 79500
rect 72600 79400 75500 79500
rect 25400 79500 28100 79700
rect 30500 79500 33400 79700
rect 35900 79500 38700 79700
rect 40900 79500 44000 79700
rect 46200 79500 49100 79700
rect 51500 79500 54400 79700
rect 56800 79500 59700 79700
rect 62000 79500 65000 79700
rect 67300 79500 70200 79700
rect 72600 79500 75500 79700
rect 25400 79700 28100 79800
rect 30500 79700 33400 79800
rect 35900 79700 38700 79800
rect 40900 79700 44000 79800
rect 46200 79700 49100 79800
rect 51500 79700 54400 79800
rect 56800 79700 59700 79800
rect 62000 79700 65000 79800
rect 67300 79700 70200 79800
rect 72600 79700 75500 79800
rect 25400 79800 28100 80000
rect 30500 79800 33400 80000
rect 35900 79800 38700 80000
rect 40900 79800 44000 80000
rect 46200 79800 49100 80000
rect 51500 79800 54400 80000
rect 56800 79800 59700 80000
rect 62000 79800 65000 80000
rect 67300 79800 70200 80000
rect 72600 79800 75500 80000
rect 25400 80000 28100 80100
rect 30500 80000 33400 80100
rect 35900 80000 38700 80100
rect 40900 80000 44000 80100
rect 46200 80000 49100 80100
rect 51500 80000 54400 80100
rect 56800 80000 59700 80100
rect 62000 80000 65000 80100
rect 67300 80000 70200 80100
rect 72600 80000 75500 80100
rect 25400 80100 28100 80200
rect 30500 80100 33400 80200
rect 35900 80100 38700 80200
rect 40900 80100 44000 80200
rect 46200 80100 49100 80200
rect 51500 80100 54400 80200
rect 56800 80100 59700 80200
rect 62000 80100 65000 80200
rect 67300 80100 70200 80200
rect 72600 80100 75500 80200
rect 25400 80200 28100 80400
rect 30500 80200 33400 80400
rect 35900 80200 38700 80400
rect 40900 80200 44000 80400
rect 46200 80200 49100 80400
rect 51500 80200 54400 80400
rect 56800 80200 59700 80400
rect 62000 80200 65000 80400
rect 67300 80200 70200 80400
rect 72600 80200 75500 80400
rect 25400 80400 28100 80500
rect 30500 80400 33400 80500
rect 35900 80400 38700 80500
rect 40900 80400 44000 80500
rect 46200 80400 49100 80500
rect 51500 80400 54400 80500
rect 56800 80400 59700 80500
rect 62000 80400 65000 80500
rect 67300 80400 70200 80500
rect 72600 80400 75500 80500
rect 25400 80500 28100 80600
rect 30500 80500 33400 80600
rect 35900 80500 38700 80600
rect 40900 80500 44000 80600
rect 46200 80500 49100 80600
rect 51500 80500 54400 80600
rect 56800 80500 59700 80600
rect 62000 80500 65000 80600
rect 67300 80500 70200 80600
rect 72600 80500 75500 80600
rect 25400 80600 28100 80800
rect 30500 80600 33400 80800
rect 35900 80600 38700 80800
rect 40900 80600 44000 80800
rect 46200 80600 49100 80800
rect 51500 80600 54400 80800
rect 56800 80600 59700 80800
rect 62000 80600 65000 80800
rect 67300 80600 70200 80800
rect 72600 80600 75500 80800
rect 25400 80800 28100 80900
rect 30500 80800 33400 80900
rect 35900 80800 38700 80900
rect 40900 80800 44000 80900
rect 46200 80800 49100 80900
rect 51500 80800 54400 80900
rect 56800 80800 59700 80900
rect 62000 80800 65000 80900
rect 67300 80800 70200 80900
rect 72600 80800 75500 80900
rect 25400 80900 28100 81100
rect 30500 80900 33400 81100
rect 35900 80900 38700 81100
rect 40900 80900 44000 81100
rect 46200 80900 49100 81100
rect 51500 80900 54400 81100
rect 56800 80900 59700 81100
rect 62000 80900 65000 81100
rect 67300 80900 70200 81100
rect 72600 80900 75500 81100
rect 25400 81100 28100 81200
rect 30500 81100 33400 81200
rect 35900 81100 38700 81200
rect 40900 81100 44000 81200
rect 46200 81100 49100 81200
rect 51500 81100 54400 81200
rect 56800 81100 59700 81200
rect 62000 81100 65000 81200
rect 67300 81100 70200 81200
rect 72600 81100 75500 81200
rect 25400 81200 28100 81300
rect 30500 81200 33400 81300
rect 35900 81200 38700 81300
rect 40900 81200 44000 81300
rect 46200 81200 49100 81300
rect 51500 81200 54400 81300
rect 56800 81200 59700 81300
rect 62000 81200 65000 81300
rect 67300 81200 70200 81300
rect 72600 81200 75500 81300
rect 25400 81300 28100 81500
rect 30500 81300 33400 81500
rect 35900 81300 38700 81500
rect 40900 81300 44000 81500
rect 46200 81300 49100 81500
rect 51500 81300 54400 81500
rect 56800 81300 59700 81500
rect 62000 81300 65000 81500
rect 67300 81300 70200 81500
rect 72600 81300 75500 81500
rect 25400 81500 28100 81600
rect 30500 81500 33400 81600
rect 35900 81500 38700 81600
rect 40900 81500 44000 81600
rect 46200 81500 49100 81600
rect 51500 81500 54400 81600
rect 56800 81500 59700 81600
rect 62000 81500 65000 81600
rect 67300 81500 70200 81600
rect 72600 81500 75500 81600
rect 25400 81600 28100 81800
rect 30500 81600 33400 81800
rect 35900 81600 38700 81800
rect 40900 81600 44000 81800
rect 46200 81600 49100 81800
rect 51500 81600 54400 81800
rect 56800 81600 59700 81800
rect 62000 81600 65000 81800
rect 67300 81600 70200 81800
rect 72600 81600 75500 81800
rect 25400 81800 28100 81900
rect 30500 81800 33400 81900
rect 35900 81800 38700 81900
rect 40900 81800 44000 81900
rect 46200 81800 49100 81900
rect 51500 81800 54400 81900
rect 56800 81800 59700 81900
rect 62000 81800 65000 81900
rect 67300 81800 70200 81900
rect 72600 81800 75500 81900
rect 25400 81900 28100 82000
rect 30500 81900 33400 82000
rect 35900 81900 38700 82000
rect 40900 81900 44000 82000
rect 46200 81900 49100 82000
rect 51500 81900 54400 82000
rect 56800 81900 59700 82000
rect 62000 81900 65000 82000
rect 67300 81900 70200 82000
rect 72600 81900 75500 82000
rect 25400 82000 28100 82200
rect 30500 82000 33400 82200
rect 35900 82000 38700 82200
rect 40900 82000 44000 82200
rect 46200 82000 49100 82200
rect 51500 82000 54400 82200
rect 56800 82000 59700 82200
rect 62000 82000 65000 82200
rect 67300 82000 70200 82200
rect 72600 82000 75500 82200
rect 25400 82200 28100 82300
rect 30500 82200 33400 82300
rect 35900 82200 38700 82300
rect 40900 82200 44000 82300
rect 46200 82200 49100 82300
rect 51500 82200 54400 82300
rect 56800 82200 59700 82300
rect 62000 82200 65000 82300
rect 67300 82200 70200 82300
rect 72600 82200 75500 82300
rect 25400 82300 28100 82500
rect 30600 82300 33400 82500
rect 35900 82300 38700 82500
rect 40900 82300 44000 82500
rect 46200 82300 49100 82500
rect 51500 82300 54300 82500
rect 56900 82300 59700 82500
rect 62000 82300 65000 82500
rect 67300 82300 70100 82500
rect 72600 82300 75500 82500
rect 25400 82500 28100 82600
rect 30600 82500 33400 82600
rect 35900 82500 38700 82600
rect 40900 82500 44000 82600
rect 46200 82500 49100 82600
rect 51500 82500 54300 82600
rect 56900 82500 59700 82600
rect 62000 82500 65000 82600
rect 67300 82500 70100 82600
rect 72700 82500 75500 82600
rect 25400 82600 28100 82700
rect 30600 82600 33400 82700
rect 35900 82600 38700 82700
rect 40900 82600 44000 82700
rect 46200 82600 49100 82700
rect 51500 82600 54300 82700
rect 56900 82600 59700 82700
rect 62000 82600 65000 82700
rect 67300 82600 70100 82700
rect 72700 82600 75500 82700
rect 25400 82700 28100 82900
rect 30600 82700 33400 82900
rect 35900 82700 38700 82900
rect 40900 82700 44000 82900
rect 46200 82700 49100 82900
rect 51500 82700 54300 82900
rect 56900 82700 59700 82900
rect 62000 82700 65000 82900
rect 67300 82700 70100 82900
rect 72700 82700 75500 82900
rect 25400 82900 28100 83000
rect 30600 82900 33400 83000
rect 35900 82900 38700 83000
rect 40900 82900 44000 83000
rect 46200 82900 49100 83000
rect 51500 82900 54300 83000
rect 56900 82900 59700 83000
rect 62000 82900 65000 83000
rect 67300 82900 70100 83000
rect 72700 82900 75500 83000
rect 25400 83000 28100 83100
rect 30600 83000 33400 83100
rect 35900 83000 38700 83100
rect 40900 83000 44000 83100
rect 46200 83000 49100 83100
rect 51500 83000 54300 83100
rect 56900 83000 59700 83100
rect 62000 83000 65000 83100
rect 67300 83000 70100 83100
rect 72700 83000 75500 83100
rect 25400 83100 28100 83300
rect 30600 83100 33400 83300
rect 35900 83100 38600 83300
rect 40900 83100 44000 83300
rect 46300 83100 49100 83300
rect 51500 83100 54300 83300
rect 56900 83100 59700 83300
rect 62000 83100 65000 83300
rect 67300 83100 70100 83300
rect 72700 83100 75500 83300
rect 25400 83300 28100 83400
rect 30600 83300 33400 83400
rect 35900 83300 38600 83400
rect 40900 83300 44000 83400
rect 46300 83300 49100 83400
rect 51500 83300 54300 83400
rect 56900 83300 59700 83400
rect 62200 83300 64800 83400
rect 67300 83300 70100 83400
rect 72700 83300 75500 83400
rect 25400 83400 28100 83600
rect 30600 83400 33400 83600
rect 35900 83400 38600 83600
rect 40900 83400 44000 83600
rect 46300 83400 49000 83600
rect 51500 83400 54300 83600
rect 56900 83400 59700 83600
rect 62200 83400 64800 83600
rect 67300 83400 70100 83600
rect 72700 83400 75500 83600
rect 25400 83600 28100 83700
rect 30600 83600 33400 83700
rect 35900 83600 38600 83700
rect 41100 83600 43800 83700
rect 46300 83600 49000 83700
rect 51500 83600 54300 83700
rect 56900 83600 59700 83700
rect 62200 83600 64800 83700
rect 67300 83600 70100 83700
rect 72700 83600 75500 83700
rect 25400 83700 28100 83800
rect 30600 83700 33300 83800
rect 35900 83700 38600 83800
rect 41200 83700 43700 83800
rect 46300 83700 49000 83800
rect 51600 83700 54300 83800
rect 56900 83700 59700 83800
rect 62200 83700 64800 83800
rect 67300 83700 70100 83800
rect 72700 83700 75400 83800
rect 25400 83800 28100 84000
rect 30600 83800 33300 84000
rect 35900 83800 38600 84000
rect 41200 83800 43700 84000
rect 46300 83800 49000 84000
rect 51600 83800 54300 84000
rect 56900 83800 59500 84000
rect 62200 83800 64800 84000
rect 67500 83800 70100 84000
rect 72700 83800 75400 84000
rect 25500 84000 28000 84100
rect 30600 84000 33300 84100
rect 35900 84000 38400 84100
rect 41200 84000 43700 84100
rect 46500 84000 49000 84100
rect 51800 84000 54300 84100
rect 57000 84000 59400 84100
rect 62300 84000 64700 84100
rect 67500 84000 70000 84100
rect 72700 84000 75200 84100
rect 25500 84100 27900 84300
rect 30800 84100 33100 84300
rect 36100 84100 38400 84300
rect 41200 84100 43700 84300
rect 46500 84100 49000 84300
rect 51800 84100 54100 84300
rect 57000 84100 59400 84300
rect 62300 84100 64700 84300
rect 67600 84100 70000 84300
rect 72700 84100 75200 84300
rect 25600 84300 27700 84400
rect 30800 84300 33000 84400
rect 36200 84300 38300 84400
rect 41300 84300 43600 84400
rect 46600 84300 48800 84400
rect 51900 84300 54100 84400
rect 57200 84300 59400 84400
rect 62500 84300 64700 84400
rect 67600 84300 69800 84400
rect 72900 84300 75100 84400
rect 25800 84400 27600 84500
rect 30900 84400 32900 84500
rect 36300 84400 38100 84500
rect 41500 84400 43400 84500
rect 46800 84400 48700 84500
rect 52000 84400 54000 84500
rect 57300 84400 59300 84500
rect 62600 84400 64500 84500
rect 67700 84400 69700 84500
rect 73000 84400 74800 84500
rect 25900 84500 27500 84700
rect 31200 84500 32700 84700
rect 36300 84500 38000 84700
rect 41600 84500 43300 84700
rect 46900 84500 48600 84700
rect 52200 84500 53700 84700
rect 57500 84500 59000 84700
rect 62700 84500 64300 84700
rect 68000 84500 69500 84700
rect 73100 84500 74800 84700
rect 26100 84700 27200 84800
rect 31300 84700 32600 84800
rect 36600 84700 37700 84800
rect 41900 84700 43000 84800
rect 47200 84700 48300 84800
rect 52300 84700 53600 84800
rect 57700 84700 58700 84800
rect 63000 84700 64000 84800
rect 68100 84700 69300 84800
rect 73400 84700 74500 84800
<< labels >>
rlabel metal4 s 100500 0 100600 100000 6 vccd1
port 1 nsew power input
rlabel metal4 s -600 0 -500 100000 6 vssd1
port 2 nsew ground input
<< end >>
