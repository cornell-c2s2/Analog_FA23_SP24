magic
tech sky130A
magscale 1 2
timestamp 1709390584
<< pwell >>
rect -739 -1582 739 1582
<< psubdiff >>
rect -703 1512 -607 1546
rect 607 1512 703 1546
rect -703 1450 -669 1512
rect 669 1450 703 1512
rect -703 -1512 -669 -1450
rect 669 -1512 703 -1450
rect -703 -1546 -607 -1512
rect 607 -1546 703 -1512
<< psubdiffcont >>
rect -607 1512 607 1546
rect -703 -1450 -669 1450
rect 669 -1450 703 1450
rect -607 -1546 607 -1512
<< xpolycontact >>
rect -573 984 573 1416
rect -573 -1416 573 -984
<< xpolyres >>
rect -573 -984 573 984
<< locali >>
rect -703 1512 -607 1546
rect 607 1512 703 1546
rect -703 1450 -669 1512
rect 669 1450 703 1512
rect -703 -1512 -669 -1450
rect 669 -1512 703 -1450
rect -703 -1546 -607 -1512
rect 607 -1546 703 -1512
<< viali >>
rect -557 1001 557 1398
rect -557 -1398 557 -1001
<< metal1 >>
rect -569 1398 569 1404
rect -569 1001 -557 1398
rect 557 1001 569 1398
rect -569 995 569 1001
rect -569 -1001 569 -995
rect -569 -1398 -557 -1001
rect 557 -1398 569 -1001
rect -569 -1404 569 -1398
<< properties >>
string FIXED_BBOX -686 -1529 686 1529
string gencell sky130_fd_pr__res_xhigh_po_5p73
string library sky130
string parameters w 5.730 l 10.0 m 1 nx 1 wmin 5.730 lmin 0.50 rho 2000 val 3.556k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 5.730 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
