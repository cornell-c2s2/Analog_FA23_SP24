magic
tech sky130A
magscale 1 2
timestamp 1713142167
<< metal3 >>
rect -5508 6772 -1996 6800
rect -5508 3608 -2080 6772
rect -2016 3608 -1996 6772
rect -5508 3580 -1996 3608
rect -1756 6772 1756 6800
rect -1756 3608 1672 6772
rect 1736 3608 1756 6772
rect -1756 3580 1756 3608
rect 1996 6772 5508 6800
rect 1996 3608 5424 6772
rect 5488 3608 5508 6772
rect 1996 3580 5508 3608
rect -5508 3312 -1996 3340
rect -5508 148 -2080 3312
rect -2016 148 -1996 3312
rect -5508 120 -1996 148
rect -1756 3312 1756 3340
rect -1756 148 1672 3312
rect 1736 148 1756 3312
rect -1756 120 1756 148
rect 1996 3312 5508 3340
rect 1996 148 5424 3312
rect 5488 148 5508 3312
rect 1996 120 5508 148
rect -5508 -148 -1996 -120
rect -5508 -3312 -2080 -148
rect -2016 -3312 -1996 -148
rect -5508 -3340 -1996 -3312
rect -1756 -148 1756 -120
rect -1756 -3312 1672 -148
rect 1736 -3312 1756 -148
rect -1756 -3340 1756 -3312
rect 1996 -148 5508 -120
rect 1996 -3312 5424 -148
rect 5488 -3312 5508 -148
rect 1996 -3340 5508 -3312
rect -5508 -3608 -1996 -3580
rect -5508 -6772 -2080 -3608
rect -2016 -6772 -1996 -3608
rect -5508 -6800 -1996 -6772
rect -1756 -3608 1756 -3580
rect -1756 -6772 1672 -3608
rect 1736 -6772 1756 -3608
rect -1756 -6800 1756 -6772
rect 1996 -3608 5508 -3580
rect 1996 -6772 5424 -3608
rect 5488 -6772 5508 -3608
rect 1996 -6800 5508 -6772
<< via3 >>
rect -2080 3608 -2016 6772
rect 1672 3608 1736 6772
rect 5424 3608 5488 6772
rect -2080 148 -2016 3312
rect 1672 148 1736 3312
rect 5424 148 5488 3312
rect -2080 -3312 -2016 -148
rect 1672 -3312 1736 -148
rect 5424 -3312 5488 -148
rect -2080 -6772 -2016 -3608
rect 1672 -6772 1736 -3608
rect 5424 -6772 5488 -3608
<< mimcap >>
rect -5468 6720 -2328 6760
rect -5468 3660 -5428 6720
rect -2368 3660 -2328 6720
rect -5468 3620 -2328 3660
rect -1716 6720 1424 6760
rect -1716 3660 -1676 6720
rect 1384 3660 1424 6720
rect -1716 3620 1424 3660
rect 2036 6720 5176 6760
rect 2036 3660 2076 6720
rect 5136 3660 5176 6720
rect 2036 3620 5176 3660
rect -5468 3260 -2328 3300
rect -5468 200 -5428 3260
rect -2368 200 -2328 3260
rect -5468 160 -2328 200
rect -1716 3260 1424 3300
rect -1716 200 -1676 3260
rect 1384 200 1424 3260
rect -1716 160 1424 200
rect 2036 3260 5176 3300
rect 2036 200 2076 3260
rect 5136 200 5176 3260
rect 2036 160 5176 200
rect -5468 -200 -2328 -160
rect -5468 -3260 -5428 -200
rect -2368 -3260 -2328 -200
rect -5468 -3300 -2328 -3260
rect -1716 -200 1424 -160
rect -1716 -3260 -1676 -200
rect 1384 -3260 1424 -200
rect -1716 -3300 1424 -3260
rect 2036 -200 5176 -160
rect 2036 -3260 2076 -200
rect 5136 -3260 5176 -200
rect 2036 -3300 5176 -3260
rect -5468 -3660 -2328 -3620
rect -5468 -6720 -5428 -3660
rect -2368 -6720 -2328 -3660
rect -5468 -6760 -2328 -6720
rect -1716 -3660 1424 -3620
rect -1716 -6720 -1676 -3660
rect 1384 -6720 1424 -3660
rect -1716 -6760 1424 -6720
rect 2036 -3660 5176 -3620
rect 2036 -6720 2076 -3660
rect 5136 -6720 5176 -3660
rect 2036 -6760 5176 -6720
<< mimcapcontact >>
rect -5428 3660 -2368 6720
rect -1676 3660 1384 6720
rect 2076 3660 5136 6720
rect -5428 200 -2368 3260
rect -1676 200 1384 3260
rect 2076 200 5136 3260
rect -5428 -3260 -2368 -200
rect -1676 -3260 1384 -200
rect 2076 -3260 5136 -200
rect -5428 -6720 -2368 -3660
rect -1676 -6720 1384 -3660
rect 2076 -6720 5136 -3660
<< metal4 >>
rect -3950 6721 -3846 6920
rect -2100 6772 -1996 6920
rect -5429 6720 -2367 6721
rect -5429 3660 -5428 6720
rect -2368 3660 -2367 6720
rect -5429 3659 -2367 3660
rect -3950 3261 -3846 3659
rect -2100 3608 -2080 6772
rect -2016 3608 -1996 6772
rect -198 6721 -94 6920
rect 1652 6772 1756 6920
rect -1677 6720 1385 6721
rect -1677 3660 -1676 6720
rect 1384 3660 1385 6720
rect -1677 3659 1385 3660
rect -2100 3312 -1996 3608
rect -5429 3260 -2367 3261
rect -5429 200 -5428 3260
rect -2368 200 -2367 3260
rect -5429 199 -2367 200
rect -3950 -199 -3846 199
rect -2100 148 -2080 3312
rect -2016 148 -1996 3312
rect -198 3261 -94 3659
rect 1652 3608 1672 6772
rect 1736 3608 1756 6772
rect 3554 6721 3658 6920
rect 5404 6772 5508 6920
rect 2075 6720 5137 6721
rect 2075 3660 2076 6720
rect 5136 3660 5137 6720
rect 2075 3659 5137 3660
rect 1652 3312 1756 3608
rect -1677 3260 1385 3261
rect -1677 200 -1676 3260
rect 1384 200 1385 3260
rect -1677 199 1385 200
rect -2100 -148 -1996 148
rect -5429 -200 -2367 -199
rect -5429 -3260 -5428 -200
rect -2368 -3260 -2367 -200
rect -5429 -3261 -2367 -3260
rect -3950 -3659 -3846 -3261
rect -2100 -3312 -2080 -148
rect -2016 -3312 -1996 -148
rect -198 -199 -94 199
rect 1652 148 1672 3312
rect 1736 148 1756 3312
rect 3554 3261 3658 3659
rect 5404 3608 5424 6772
rect 5488 3608 5508 6772
rect 5404 3312 5508 3608
rect 2075 3260 5137 3261
rect 2075 200 2076 3260
rect 5136 200 5137 3260
rect 2075 199 5137 200
rect 1652 -148 1756 148
rect -1677 -200 1385 -199
rect -1677 -3260 -1676 -200
rect 1384 -3260 1385 -200
rect -1677 -3261 1385 -3260
rect -2100 -3608 -1996 -3312
rect -5429 -3660 -2367 -3659
rect -5429 -6720 -5428 -3660
rect -2368 -6720 -2367 -3660
rect -5429 -6721 -2367 -6720
rect -3950 -6920 -3846 -6721
rect -2100 -6772 -2080 -3608
rect -2016 -6772 -1996 -3608
rect -198 -3659 -94 -3261
rect 1652 -3312 1672 -148
rect 1736 -3312 1756 -148
rect 3554 -199 3658 199
rect 5404 148 5424 3312
rect 5488 148 5508 3312
rect 5404 -148 5508 148
rect 2075 -200 5137 -199
rect 2075 -3260 2076 -200
rect 5136 -3260 5137 -200
rect 2075 -3261 5137 -3260
rect 1652 -3608 1756 -3312
rect -1677 -3660 1385 -3659
rect -1677 -6720 -1676 -3660
rect 1384 -6720 1385 -3660
rect -1677 -6721 1385 -6720
rect -2100 -6920 -1996 -6772
rect -198 -6920 -94 -6721
rect 1652 -6772 1672 -3608
rect 1736 -6772 1756 -3608
rect 3554 -3659 3658 -3261
rect 5404 -3312 5424 -148
rect 5488 -3312 5508 -148
rect 5404 -3608 5508 -3312
rect 2075 -3660 5137 -3659
rect 2075 -6720 2076 -3660
rect 5136 -6720 5137 -3660
rect 2075 -6721 5137 -6720
rect 1652 -6920 1756 -6772
rect 3554 -6920 3658 -6721
rect 5404 -6772 5424 -3608
rect 5488 -6772 5508 -3608
rect 5404 -6920 5508 -6772
<< properties >>
string FIXED_BBOX 1996 3580 5216 6800
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 15.7 l 15.7 val 504.912 carea 2.00 cperi 0.19 nx 3 ny 4 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
