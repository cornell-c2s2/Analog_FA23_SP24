magic
tech sky130A
magscale 1 2
timestamp 1714790421
<< pwell >>
rect -5086 -13704 5086 13704
<< psubdiff >>
rect -5050 13634 -4954 13668
rect 4954 13634 5050 13668
rect -5050 13572 -5016 13634
rect 5016 13572 5050 13634
rect -5050 -13634 -5016 -13572
rect 5016 -13634 5050 -13572
rect -5050 -13668 -4954 -13634
rect 4954 -13668 5050 -13634
<< psubdiffcont >>
rect -4954 13634 4954 13668
rect -5050 -13572 -5016 13572
rect 5016 -13572 5050 13572
rect -4954 -13668 4954 -13634
<< xpolycontact >>
rect -4920 13106 -3774 13538
rect -4920 12132 -3774 12564
rect -3678 13106 -2532 13538
rect -3678 12132 -2532 12564
rect -2436 13106 -1290 13538
rect -2436 12132 -1290 12564
rect -1194 13106 -48 13538
rect -1194 12132 -48 12564
rect 48 13106 1194 13538
rect 48 12132 1194 12564
rect 1290 13106 2436 13538
rect 1290 12132 2436 12564
rect 2532 13106 3678 13538
rect 2532 12132 3678 12564
rect 3774 13106 4920 13538
rect 3774 12132 4920 12564
rect -4920 11596 -3774 12028
rect -4920 10622 -3774 11054
rect -3678 11596 -2532 12028
rect -3678 10622 -2532 11054
rect -2436 11596 -1290 12028
rect -2436 10622 -1290 11054
rect -1194 11596 -48 12028
rect -1194 10622 -48 11054
rect 48 11596 1194 12028
rect 48 10622 1194 11054
rect 1290 11596 2436 12028
rect 1290 10622 2436 11054
rect 2532 11596 3678 12028
rect 2532 10622 3678 11054
rect 3774 11596 4920 12028
rect 3774 10622 4920 11054
rect -4920 10086 -3774 10518
rect -4920 9112 -3774 9544
rect -3678 10086 -2532 10518
rect -3678 9112 -2532 9544
rect -2436 10086 -1290 10518
rect -2436 9112 -1290 9544
rect -1194 10086 -48 10518
rect -1194 9112 -48 9544
rect 48 10086 1194 10518
rect 48 9112 1194 9544
rect 1290 10086 2436 10518
rect 1290 9112 2436 9544
rect 2532 10086 3678 10518
rect 2532 9112 3678 9544
rect 3774 10086 4920 10518
rect 3774 9112 4920 9544
rect -4920 8576 -3774 9008
rect -4920 7602 -3774 8034
rect -3678 8576 -2532 9008
rect -3678 7602 -2532 8034
rect -2436 8576 -1290 9008
rect -2436 7602 -1290 8034
rect -1194 8576 -48 9008
rect -1194 7602 -48 8034
rect 48 8576 1194 9008
rect 48 7602 1194 8034
rect 1290 8576 2436 9008
rect 1290 7602 2436 8034
rect 2532 8576 3678 9008
rect 2532 7602 3678 8034
rect 3774 8576 4920 9008
rect 3774 7602 4920 8034
rect -4920 7066 -3774 7498
rect -4920 6092 -3774 6524
rect -3678 7066 -2532 7498
rect -3678 6092 -2532 6524
rect -2436 7066 -1290 7498
rect -2436 6092 -1290 6524
rect -1194 7066 -48 7498
rect -1194 6092 -48 6524
rect 48 7066 1194 7498
rect 48 6092 1194 6524
rect 1290 7066 2436 7498
rect 1290 6092 2436 6524
rect 2532 7066 3678 7498
rect 2532 6092 3678 6524
rect 3774 7066 4920 7498
rect 3774 6092 4920 6524
rect -4920 5556 -3774 5988
rect -4920 4582 -3774 5014
rect -3678 5556 -2532 5988
rect -3678 4582 -2532 5014
rect -2436 5556 -1290 5988
rect -2436 4582 -1290 5014
rect -1194 5556 -48 5988
rect -1194 4582 -48 5014
rect 48 5556 1194 5988
rect 48 4582 1194 5014
rect 1290 5556 2436 5988
rect 1290 4582 2436 5014
rect 2532 5556 3678 5988
rect 2532 4582 3678 5014
rect 3774 5556 4920 5988
rect 3774 4582 4920 5014
rect -4920 4046 -3774 4478
rect -4920 3072 -3774 3504
rect -3678 4046 -2532 4478
rect -3678 3072 -2532 3504
rect -2436 4046 -1290 4478
rect -2436 3072 -1290 3504
rect -1194 4046 -48 4478
rect -1194 3072 -48 3504
rect 48 4046 1194 4478
rect 48 3072 1194 3504
rect 1290 4046 2436 4478
rect 1290 3072 2436 3504
rect 2532 4046 3678 4478
rect 2532 3072 3678 3504
rect 3774 4046 4920 4478
rect 3774 3072 4920 3504
rect -4920 2536 -3774 2968
rect -4920 1562 -3774 1994
rect -3678 2536 -2532 2968
rect -3678 1562 -2532 1994
rect -2436 2536 -1290 2968
rect -2436 1562 -1290 1994
rect -1194 2536 -48 2968
rect -1194 1562 -48 1994
rect 48 2536 1194 2968
rect 48 1562 1194 1994
rect 1290 2536 2436 2968
rect 1290 1562 2436 1994
rect 2532 2536 3678 2968
rect 2532 1562 3678 1994
rect 3774 2536 4920 2968
rect 3774 1562 4920 1994
rect -4920 1026 -3774 1458
rect -4920 52 -3774 484
rect -3678 1026 -2532 1458
rect -3678 52 -2532 484
rect -2436 1026 -1290 1458
rect -2436 52 -1290 484
rect -1194 1026 -48 1458
rect -1194 52 -48 484
rect 48 1026 1194 1458
rect 48 52 1194 484
rect 1290 1026 2436 1458
rect 1290 52 2436 484
rect 2532 1026 3678 1458
rect 2532 52 3678 484
rect 3774 1026 4920 1458
rect 3774 52 4920 484
rect -4920 -484 -3774 -52
rect -4920 -1458 -3774 -1026
rect -3678 -484 -2532 -52
rect -3678 -1458 -2532 -1026
rect -2436 -484 -1290 -52
rect -2436 -1458 -1290 -1026
rect -1194 -484 -48 -52
rect -1194 -1458 -48 -1026
rect 48 -484 1194 -52
rect 48 -1458 1194 -1026
rect 1290 -484 2436 -52
rect 1290 -1458 2436 -1026
rect 2532 -484 3678 -52
rect 2532 -1458 3678 -1026
rect 3774 -484 4920 -52
rect 3774 -1458 4920 -1026
rect -4920 -1994 -3774 -1562
rect -4920 -2968 -3774 -2536
rect -3678 -1994 -2532 -1562
rect -3678 -2968 -2532 -2536
rect -2436 -1994 -1290 -1562
rect -2436 -2968 -1290 -2536
rect -1194 -1994 -48 -1562
rect -1194 -2968 -48 -2536
rect 48 -1994 1194 -1562
rect 48 -2968 1194 -2536
rect 1290 -1994 2436 -1562
rect 1290 -2968 2436 -2536
rect 2532 -1994 3678 -1562
rect 2532 -2968 3678 -2536
rect 3774 -1994 4920 -1562
rect 3774 -2968 4920 -2536
rect -4920 -3504 -3774 -3072
rect -4920 -4478 -3774 -4046
rect -3678 -3504 -2532 -3072
rect -3678 -4478 -2532 -4046
rect -2436 -3504 -1290 -3072
rect -2436 -4478 -1290 -4046
rect -1194 -3504 -48 -3072
rect -1194 -4478 -48 -4046
rect 48 -3504 1194 -3072
rect 48 -4478 1194 -4046
rect 1290 -3504 2436 -3072
rect 1290 -4478 2436 -4046
rect 2532 -3504 3678 -3072
rect 2532 -4478 3678 -4046
rect 3774 -3504 4920 -3072
rect 3774 -4478 4920 -4046
rect -4920 -5014 -3774 -4582
rect -4920 -5988 -3774 -5556
rect -3678 -5014 -2532 -4582
rect -3678 -5988 -2532 -5556
rect -2436 -5014 -1290 -4582
rect -2436 -5988 -1290 -5556
rect -1194 -5014 -48 -4582
rect -1194 -5988 -48 -5556
rect 48 -5014 1194 -4582
rect 48 -5988 1194 -5556
rect 1290 -5014 2436 -4582
rect 1290 -5988 2436 -5556
rect 2532 -5014 3678 -4582
rect 2532 -5988 3678 -5556
rect 3774 -5014 4920 -4582
rect 3774 -5988 4920 -5556
rect -4920 -6524 -3774 -6092
rect -4920 -7498 -3774 -7066
rect -3678 -6524 -2532 -6092
rect -3678 -7498 -2532 -7066
rect -2436 -6524 -1290 -6092
rect -2436 -7498 -1290 -7066
rect -1194 -6524 -48 -6092
rect -1194 -7498 -48 -7066
rect 48 -6524 1194 -6092
rect 48 -7498 1194 -7066
rect 1290 -6524 2436 -6092
rect 1290 -7498 2436 -7066
rect 2532 -6524 3678 -6092
rect 2532 -7498 3678 -7066
rect 3774 -6524 4920 -6092
rect 3774 -7498 4920 -7066
rect -4920 -8034 -3774 -7602
rect -4920 -9008 -3774 -8576
rect -3678 -8034 -2532 -7602
rect -3678 -9008 -2532 -8576
rect -2436 -8034 -1290 -7602
rect -2436 -9008 -1290 -8576
rect -1194 -8034 -48 -7602
rect -1194 -9008 -48 -8576
rect 48 -8034 1194 -7602
rect 48 -9008 1194 -8576
rect 1290 -8034 2436 -7602
rect 1290 -9008 2436 -8576
rect 2532 -8034 3678 -7602
rect 2532 -9008 3678 -8576
rect 3774 -8034 4920 -7602
rect 3774 -9008 4920 -8576
rect -4920 -9544 -3774 -9112
rect -4920 -10518 -3774 -10086
rect -3678 -9544 -2532 -9112
rect -3678 -10518 -2532 -10086
rect -2436 -9544 -1290 -9112
rect -2436 -10518 -1290 -10086
rect -1194 -9544 -48 -9112
rect -1194 -10518 -48 -10086
rect 48 -9544 1194 -9112
rect 48 -10518 1194 -10086
rect 1290 -9544 2436 -9112
rect 1290 -10518 2436 -10086
rect 2532 -9544 3678 -9112
rect 2532 -10518 3678 -10086
rect 3774 -9544 4920 -9112
rect 3774 -10518 4920 -10086
rect -4920 -11054 -3774 -10622
rect -4920 -12028 -3774 -11596
rect -3678 -11054 -2532 -10622
rect -3678 -12028 -2532 -11596
rect -2436 -11054 -1290 -10622
rect -2436 -12028 -1290 -11596
rect -1194 -11054 -48 -10622
rect -1194 -12028 -48 -11596
rect 48 -11054 1194 -10622
rect 48 -12028 1194 -11596
rect 1290 -11054 2436 -10622
rect 1290 -12028 2436 -11596
rect 2532 -11054 3678 -10622
rect 2532 -12028 3678 -11596
rect 3774 -11054 4920 -10622
rect 3774 -12028 4920 -11596
rect -4920 -12564 -3774 -12132
rect -4920 -13538 -3774 -13106
rect -3678 -12564 -2532 -12132
rect -3678 -13538 -2532 -13106
rect -2436 -12564 -1290 -12132
rect -2436 -13538 -1290 -13106
rect -1194 -12564 -48 -12132
rect -1194 -13538 -48 -13106
rect 48 -12564 1194 -12132
rect 48 -13538 1194 -13106
rect 1290 -12564 2436 -12132
rect 1290 -13538 2436 -13106
rect 2532 -12564 3678 -12132
rect 2532 -13538 3678 -13106
rect 3774 -12564 4920 -12132
rect 3774 -13538 4920 -13106
<< xpolyres >>
rect -4920 12564 -3774 13106
rect -3678 12564 -2532 13106
rect -2436 12564 -1290 13106
rect -1194 12564 -48 13106
rect 48 12564 1194 13106
rect 1290 12564 2436 13106
rect 2532 12564 3678 13106
rect 3774 12564 4920 13106
rect -4920 11054 -3774 11596
rect -3678 11054 -2532 11596
rect -2436 11054 -1290 11596
rect -1194 11054 -48 11596
rect 48 11054 1194 11596
rect 1290 11054 2436 11596
rect 2532 11054 3678 11596
rect 3774 11054 4920 11596
rect -4920 9544 -3774 10086
rect -3678 9544 -2532 10086
rect -2436 9544 -1290 10086
rect -1194 9544 -48 10086
rect 48 9544 1194 10086
rect 1290 9544 2436 10086
rect 2532 9544 3678 10086
rect 3774 9544 4920 10086
rect -4920 8034 -3774 8576
rect -3678 8034 -2532 8576
rect -2436 8034 -1290 8576
rect -1194 8034 -48 8576
rect 48 8034 1194 8576
rect 1290 8034 2436 8576
rect 2532 8034 3678 8576
rect 3774 8034 4920 8576
rect -4920 6524 -3774 7066
rect -3678 6524 -2532 7066
rect -2436 6524 -1290 7066
rect -1194 6524 -48 7066
rect 48 6524 1194 7066
rect 1290 6524 2436 7066
rect 2532 6524 3678 7066
rect 3774 6524 4920 7066
rect -4920 5014 -3774 5556
rect -3678 5014 -2532 5556
rect -2436 5014 -1290 5556
rect -1194 5014 -48 5556
rect 48 5014 1194 5556
rect 1290 5014 2436 5556
rect 2532 5014 3678 5556
rect 3774 5014 4920 5556
rect -4920 3504 -3774 4046
rect -3678 3504 -2532 4046
rect -2436 3504 -1290 4046
rect -1194 3504 -48 4046
rect 48 3504 1194 4046
rect 1290 3504 2436 4046
rect 2532 3504 3678 4046
rect 3774 3504 4920 4046
rect -4920 1994 -3774 2536
rect -3678 1994 -2532 2536
rect -2436 1994 -1290 2536
rect -1194 1994 -48 2536
rect 48 1994 1194 2536
rect 1290 1994 2436 2536
rect 2532 1994 3678 2536
rect 3774 1994 4920 2536
rect -4920 484 -3774 1026
rect -3678 484 -2532 1026
rect -2436 484 -1290 1026
rect -1194 484 -48 1026
rect 48 484 1194 1026
rect 1290 484 2436 1026
rect 2532 484 3678 1026
rect 3774 484 4920 1026
rect -4920 -1026 -3774 -484
rect -3678 -1026 -2532 -484
rect -2436 -1026 -1290 -484
rect -1194 -1026 -48 -484
rect 48 -1026 1194 -484
rect 1290 -1026 2436 -484
rect 2532 -1026 3678 -484
rect 3774 -1026 4920 -484
rect -4920 -2536 -3774 -1994
rect -3678 -2536 -2532 -1994
rect -2436 -2536 -1290 -1994
rect -1194 -2536 -48 -1994
rect 48 -2536 1194 -1994
rect 1290 -2536 2436 -1994
rect 2532 -2536 3678 -1994
rect 3774 -2536 4920 -1994
rect -4920 -4046 -3774 -3504
rect -3678 -4046 -2532 -3504
rect -2436 -4046 -1290 -3504
rect -1194 -4046 -48 -3504
rect 48 -4046 1194 -3504
rect 1290 -4046 2436 -3504
rect 2532 -4046 3678 -3504
rect 3774 -4046 4920 -3504
rect -4920 -5556 -3774 -5014
rect -3678 -5556 -2532 -5014
rect -2436 -5556 -1290 -5014
rect -1194 -5556 -48 -5014
rect 48 -5556 1194 -5014
rect 1290 -5556 2436 -5014
rect 2532 -5556 3678 -5014
rect 3774 -5556 4920 -5014
rect -4920 -7066 -3774 -6524
rect -3678 -7066 -2532 -6524
rect -2436 -7066 -1290 -6524
rect -1194 -7066 -48 -6524
rect 48 -7066 1194 -6524
rect 1290 -7066 2436 -6524
rect 2532 -7066 3678 -6524
rect 3774 -7066 4920 -6524
rect -4920 -8576 -3774 -8034
rect -3678 -8576 -2532 -8034
rect -2436 -8576 -1290 -8034
rect -1194 -8576 -48 -8034
rect 48 -8576 1194 -8034
rect 1290 -8576 2436 -8034
rect 2532 -8576 3678 -8034
rect 3774 -8576 4920 -8034
rect -4920 -10086 -3774 -9544
rect -3678 -10086 -2532 -9544
rect -2436 -10086 -1290 -9544
rect -1194 -10086 -48 -9544
rect 48 -10086 1194 -9544
rect 1290 -10086 2436 -9544
rect 2532 -10086 3678 -9544
rect 3774 -10086 4920 -9544
rect -4920 -11596 -3774 -11054
rect -3678 -11596 -2532 -11054
rect -2436 -11596 -1290 -11054
rect -1194 -11596 -48 -11054
rect 48 -11596 1194 -11054
rect 1290 -11596 2436 -11054
rect 2532 -11596 3678 -11054
rect 3774 -11596 4920 -11054
rect -4920 -13106 -3774 -12564
rect -3678 -13106 -2532 -12564
rect -2436 -13106 -1290 -12564
rect -1194 -13106 -48 -12564
rect 48 -13106 1194 -12564
rect 1290 -13106 2436 -12564
rect 2532 -13106 3678 -12564
rect 3774 -13106 4920 -12564
<< locali >>
rect -5050 13634 -4954 13668
rect 4954 13634 5050 13668
rect -5050 13572 -5016 13634
rect 5016 13572 5050 13634
rect -5050 -13634 -5016 -13572
rect 5016 -13634 5050 -13572
rect -5050 -13668 -4954 -13634
rect 4954 -13668 5050 -13634
<< viali >>
rect -4904 13123 -3790 13520
rect -3662 13123 -2548 13520
rect -2420 13123 -1306 13520
rect -1178 13123 -64 13520
rect 64 13123 1178 13520
rect 1306 13123 2420 13520
rect 2548 13123 3662 13520
rect 3790 13123 4904 13520
rect -4904 12150 -3790 12547
rect -3662 12150 -2548 12547
rect -2420 12150 -1306 12547
rect -1178 12150 -64 12547
rect 64 12150 1178 12547
rect 1306 12150 2420 12547
rect 2548 12150 3662 12547
rect 3790 12150 4904 12547
rect -4904 11613 -3790 12010
rect -3662 11613 -2548 12010
rect -2420 11613 -1306 12010
rect -1178 11613 -64 12010
rect 64 11613 1178 12010
rect 1306 11613 2420 12010
rect 2548 11613 3662 12010
rect 3790 11613 4904 12010
rect -4904 10640 -3790 11037
rect -3662 10640 -2548 11037
rect -2420 10640 -1306 11037
rect -1178 10640 -64 11037
rect 64 10640 1178 11037
rect 1306 10640 2420 11037
rect 2548 10640 3662 11037
rect 3790 10640 4904 11037
rect -4904 10103 -3790 10500
rect -3662 10103 -2548 10500
rect -2420 10103 -1306 10500
rect -1178 10103 -64 10500
rect 64 10103 1178 10500
rect 1306 10103 2420 10500
rect 2548 10103 3662 10500
rect 3790 10103 4904 10500
rect -4904 9130 -3790 9527
rect -3662 9130 -2548 9527
rect -2420 9130 -1306 9527
rect -1178 9130 -64 9527
rect 64 9130 1178 9527
rect 1306 9130 2420 9527
rect 2548 9130 3662 9527
rect 3790 9130 4904 9527
rect -4904 8593 -3790 8990
rect -3662 8593 -2548 8990
rect -2420 8593 -1306 8990
rect -1178 8593 -64 8990
rect 64 8593 1178 8990
rect 1306 8593 2420 8990
rect 2548 8593 3662 8990
rect 3790 8593 4904 8990
rect -4904 7620 -3790 8017
rect -3662 7620 -2548 8017
rect -2420 7620 -1306 8017
rect -1178 7620 -64 8017
rect 64 7620 1178 8017
rect 1306 7620 2420 8017
rect 2548 7620 3662 8017
rect 3790 7620 4904 8017
rect -4904 7083 -3790 7480
rect -3662 7083 -2548 7480
rect -2420 7083 -1306 7480
rect -1178 7083 -64 7480
rect 64 7083 1178 7480
rect 1306 7083 2420 7480
rect 2548 7083 3662 7480
rect 3790 7083 4904 7480
rect -4904 6110 -3790 6507
rect -3662 6110 -2548 6507
rect -2420 6110 -1306 6507
rect -1178 6110 -64 6507
rect 64 6110 1178 6507
rect 1306 6110 2420 6507
rect 2548 6110 3662 6507
rect 3790 6110 4904 6507
rect -4904 5573 -3790 5970
rect -3662 5573 -2548 5970
rect -2420 5573 -1306 5970
rect -1178 5573 -64 5970
rect 64 5573 1178 5970
rect 1306 5573 2420 5970
rect 2548 5573 3662 5970
rect 3790 5573 4904 5970
rect -4904 4600 -3790 4997
rect -3662 4600 -2548 4997
rect -2420 4600 -1306 4997
rect -1178 4600 -64 4997
rect 64 4600 1178 4997
rect 1306 4600 2420 4997
rect 2548 4600 3662 4997
rect 3790 4600 4904 4997
rect -4904 4063 -3790 4460
rect -3662 4063 -2548 4460
rect -2420 4063 -1306 4460
rect -1178 4063 -64 4460
rect 64 4063 1178 4460
rect 1306 4063 2420 4460
rect 2548 4063 3662 4460
rect 3790 4063 4904 4460
rect -4904 3090 -3790 3487
rect -3662 3090 -2548 3487
rect -2420 3090 -1306 3487
rect -1178 3090 -64 3487
rect 64 3090 1178 3487
rect 1306 3090 2420 3487
rect 2548 3090 3662 3487
rect 3790 3090 4904 3487
rect -4904 2553 -3790 2950
rect -3662 2553 -2548 2950
rect -2420 2553 -1306 2950
rect -1178 2553 -64 2950
rect 64 2553 1178 2950
rect 1306 2553 2420 2950
rect 2548 2553 3662 2950
rect 3790 2553 4904 2950
rect -4904 1580 -3790 1977
rect -3662 1580 -2548 1977
rect -2420 1580 -1306 1977
rect -1178 1580 -64 1977
rect 64 1580 1178 1977
rect 1306 1580 2420 1977
rect 2548 1580 3662 1977
rect 3790 1580 4904 1977
rect -4904 1043 -3790 1440
rect -3662 1043 -2548 1440
rect -2420 1043 -1306 1440
rect -1178 1043 -64 1440
rect 64 1043 1178 1440
rect 1306 1043 2420 1440
rect 2548 1043 3662 1440
rect 3790 1043 4904 1440
rect -4904 70 -3790 467
rect -3662 70 -2548 467
rect -2420 70 -1306 467
rect -1178 70 -64 467
rect 64 70 1178 467
rect 1306 70 2420 467
rect 2548 70 3662 467
rect 3790 70 4904 467
rect -4904 -467 -3790 -70
rect -3662 -467 -2548 -70
rect -2420 -467 -1306 -70
rect -1178 -467 -64 -70
rect 64 -467 1178 -70
rect 1306 -467 2420 -70
rect 2548 -467 3662 -70
rect 3790 -467 4904 -70
rect -4904 -1440 -3790 -1043
rect -3662 -1440 -2548 -1043
rect -2420 -1440 -1306 -1043
rect -1178 -1440 -64 -1043
rect 64 -1440 1178 -1043
rect 1306 -1440 2420 -1043
rect 2548 -1440 3662 -1043
rect 3790 -1440 4904 -1043
rect -4904 -1977 -3790 -1580
rect -3662 -1977 -2548 -1580
rect -2420 -1977 -1306 -1580
rect -1178 -1977 -64 -1580
rect 64 -1977 1178 -1580
rect 1306 -1977 2420 -1580
rect 2548 -1977 3662 -1580
rect 3790 -1977 4904 -1580
rect -4904 -2950 -3790 -2553
rect -3662 -2950 -2548 -2553
rect -2420 -2950 -1306 -2553
rect -1178 -2950 -64 -2553
rect 64 -2950 1178 -2553
rect 1306 -2950 2420 -2553
rect 2548 -2950 3662 -2553
rect 3790 -2950 4904 -2553
rect -4904 -3487 -3790 -3090
rect -3662 -3487 -2548 -3090
rect -2420 -3487 -1306 -3090
rect -1178 -3487 -64 -3090
rect 64 -3487 1178 -3090
rect 1306 -3487 2420 -3090
rect 2548 -3487 3662 -3090
rect 3790 -3487 4904 -3090
rect -4904 -4460 -3790 -4063
rect -3662 -4460 -2548 -4063
rect -2420 -4460 -1306 -4063
rect -1178 -4460 -64 -4063
rect 64 -4460 1178 -4063
rect 1306 -4460 2420 -4063
rect 2548 -4460 3662 -4063
rect 3790 -4460 4904 -4063
rect -4904 -4997 -3790 -4600
rect -3662 -4997 -2548 -4600
rect -2420 -4997 -1306 -4600
rect -1178 -4997 -64 -4600
rect 64 -4997 1178 -4600
rect 1306 -4997 2420 -4600
rect 2548 -4997 3662 -4600
rect 3790 -4997 4904 -4600
rect -4904 -5970 -3790 -5573
rect -3662 -5970 -2548 -5573
rect -2420 -5970 -1306 -5573
rect -1178 -5970 -64 -5573
rect 64 -5970 1178 -5573
rect 1306 -5970 2420 -5573
rect 2548 -5970 3662 -5573
rect 3790 -5970 4904 -5573
rect -4904 -6507 -3790 -6110
rect -3662 -6507 -2548 -6110
rect -2420 -6507 -1306 -6110
rect -1178 -6507 -64 -6110
rect 64 -6507 1178 -6110
rect 1306 -6507 2420 -6110
rect 2548 -6507 3662 -6110
rect 3790 -6507 4904 -6110
rect -4904 -7480 -3790 -7083
rect -3662 -7480 -2548 -7083
rect -2420 -7480 -1306 -7083
rect -1178 -7480 -64 -7083
rect 64 -7480 1178 -7083
rect 1306 -7480 2420 -7083
rect 2548 -7480 3662 -7083
rect 3790 -7480 4904 -7083
rect -4904 -8017 -3790 -7620
rect -3662 -8017 -2548 -7620
rect -2420 -8017 -1306 -7620
rect -1178 -8017 -64 -7620
rect 64 -8017 1178 -7620
rect 1306 -8017 2420 -7620
rect 2548 -8017 3662 -7620
rect 3790 -8017 4904 -7620
rect -4904 -8990 -3790 -8593
rect -3662 -8990 -2548 -8593
rect -2420 -8990 -1306 -8593
rect -1178 -8990 -64 -8593
rect 64 -8990 1178 -8593
rect 1306 -8990 2420 -8593
rect 2548 -8990 3662 -8593
rect 3790 -8990 4904 -8593
rect -4904 -9527 -3790 -9130
rect -3662 -9527 -2548 -9130
rect -2420 -9527 -1306 -9130
rect -1178 -9527 -64 -9130
rect 64 -9527 1178 -9130
rect 1306 -9527 2420 -9130
rect 2548 -9527 3662 -9130
rect 3790 -9527 4904 -9130
rect -4904 -10500 -3790 -10103
rect -3662 -10500 -2548 -10103
rect -2420 -10500 -1306 -10103
rect -1178 -10500 -64 -10103
rect 64 -10500 1178 -10103
rect 1306 -10500 2420 -10103
rect 2548 -10500 3662 -10103
rect 3790 -10500 4904 -10103
rect -4904 -11037 -3790 -10640
rect -3662 -11037 -2548 -10640
rect -2420 -11037 -1306 -10640
rect -1178 -11037 -64 -10640
rect 64 -11037 1178 -10640
rect 1306 -11037 2420 -10640
rect 2548 -11037 3662 -10640
rect 3790 -11037 4904 -10640
rect -4904 -12010 -3790 -11613
rect -3662 -12010 -2548 -11613
rect -2420 -12010 -1306 -11613
rect -1178 -12010 -64 -11613
rect 64 -12010 1178 -11613
rect 1306 -12010 2420 -11613
rect 2548 -12010 3662 -11613
rect 3790 -12010 4904 -11613
rect -4904 -12547 -3790 -12150
rect -3662 -12547 -2548 -12150
rect -2420 -12547 -1306 -12150
rect -1178 -12547 -64 -12150
rect 64 -12547 1178 -12150
rect 1306 -12547 2420 -12150
rect 2548 -12547 3662 -12150
rect 3790 -12547 4904 -12150
rect -4904 -13520 -3790 -13123
rect -3662 -13520 -2548 -13123
rect -2420 -13520 -1306 -13123
rect -1178 -13520 -64 -13123
rect 64 -13520 1178 -13123
rect 1306 -13520 2420 -13123
rect 2548 -13520 3662 -13123
rect 3790 -13520 4904 -13123
<< metal1 >>
rect -4916 13520 -3778 13526
rect -4916 13123 -4904 13520
rect -3790 13123 -3778 13520
rect -4916 13117 -3778 13123
rect -3674 13520 -2536 13526
rect -3674 13123 -3662 13520
rect -2548 13123 -2536 13520
rect -3674 13117 -2536 13123
rect -2432 13520 -1294 13526
rect -2432 13123 -2420 13520
rect -1306 13123 -1294 13520
rect -2432 13117 -1294 13123
rect -1190 13520 -52 13526
rect -1190 13123 -1178 13520
rect -64 13123 -52 13520
rect -1190 13117 -52 13123
rect 52 13520 1190 13526
rect 52 13123 64 13520
rect 1178 13123 1190 13520
rect 52 13117 1190 13123
rect 1294 13520 2432 13526
rect 1294 13123 1306 13520
rect 2420 13123 2432 13520
rect 1294 13117 2432 13123
rect 2536 13520 3674 13526
rect 2536 13123 2548 13520
rect 3662 13123 3674 13520
rect 2536 13117 3674 13123
rect 3778 13520 4916 13526
rect 3778 13123 3790 13520
rect 4904 13123 4916 13520
rect 3778 13117 4916 13123
rect -4916 12547 -3778 12553
rect -4916 12150 -4904 12547
rect -3790 12150 -3778 12547
rect -4916 12144 -3778 12150
rect -3674 12547 -2536 12553
rect -3674 12150 -3662 12547
rect -2548 12150 -2536 12547
rect -3674 12144 -2536 12150
rect -2432 12547 -1294 12553
rect -2432 12150 -2420 12547
rect -1306 12150 -1294 12547
rect -2432 12144 -1294 12150
rect -1190 12547 -52 12553
rect -1190 12150 -1178 12547
rect -64 12150 -52 12547
rect -1190 12144 -52 12150
rect 52 12547 1190 12553
rect 52 12150 64 12547
rect 1178 12150 1190 12547
rect 52 12144 1190 12150
rect 1294 12547 2432 12553
rect 1294 12150 1306 12547
rect 2420 12150 2432 12547
rect 1294 12144 2432 12150
rect 2536 12547 3674 12553
rect 2536 12150 2548 12547
rect 3662 12150 3674 12547
rect 2536 12144 3674 12150
rect 3778 12547 4916 12553
rect 3778 12150 3790 12547
rect 4904 12150 4916 12547
rect 3778 12144 4916 12150
rect -4916 12010 -3778 12016
rect -4916 11613 -4904 12010
rect -3790 11613 -3778 12010
rect -4916 11607 -3778 11613
rect -3674 12010 -2536 12016
rect -3674 11613 -3662 12010
rect -2548 11613 -2536 12010
rect -3674 11607 -2536 11613
rect -2432 12010 -1294 12016
rect -2432 11613 -2420 12010
rect -1306 11613 -1294 12010
rect -2432 11607 -1294 11613
rect -1190 12010 -52 12016
rect -1190 11613 -1178 12010
rect -64 11613 -52 12010
rect -1190 11607 -52 11613
rect 52 12010 1190 12016
rect 52 11613 64 12010
rect 1178 11613 1190 12010
rect 52 11607 1190 11613
rect 1294 12010 2432 12016
rect 1294 11613 1306 12010
rect 2420 11613 2432 12010
rect 1294 11607 2432 11613
rect 2536 12010 3674 12016
rect 2536 11613 2548 12010
rect 3662 11613 3674 12010
rect 2536 11607 3674 11613
rect 3778 12010 4916 12016
rect 3778 11613 3790 12010
rect 4904 11613 4916 12010
rect 3778 11607 4916 11613
rect -4916 11037 -3778 11043
rect -4916 10640 -4904 11037
rect -3790 10640 -3778 11037
rect -4916 10634 -3778 10640
rect -3674 11037 -2536 11043
rect -3674 10640 -3662 11037
rect -2548 10640 -2536 11037
rect -3674 10634 -2536 10640
rect -2432 11037 -1294 11043
rect -2432 10640 -2420 11037
rect -1306 10640 -1294 11037
rect -2432 10634 -1294 10640
rect -1190 11037 -52 11043
rect -1190 10640 -1178 11037
rect -64 10640 -52 11037
rect -1190 10634 -52 10640
rect 52 11037 1190 11043
rect 52 10640 64 11037
rect 1178 10640 1190 11037
rect 52 10634 1190 10640
rect 1294 11037 2432 11043
rect 1294 10640 1306 11037
rect 2420 10640 2432 11037
rect 1294 10634 2432 10640
rect 2536 11037 3674 11043
rect 2536 10640 2548 11037
rect 3662 10640 3674 11037
rect 2536 10634 3674 10640
rect 3778 11037 4916 11043
rect 3778 10640 3790 11037
rect 4904 10640 4916 11037
rect 3778 10634 4916 10640
rect -4916 10500 -3778 10506
rect -4916 10103 -4904 10500
rect -3790 10103 -3778 10500
rect -4916 10097 -3778 10103
rect -3674 10500 -2536 10506
rect -3674 10103 -3662 10500
rect -2548 10103 -2536 10500
rect -3674 10097 -2536 10103
rect -2432 10500 -1294 10506
rect -2432 10103 -2420 10500
rect -1306 10103 -1294 10500
rect -2432 10097 -1294 10103
rect -1190 10500 -52 10506
rect -1190 10103 -1178 10500
rect -64 10103 -52 10500
rect -1190 10097 -52 10103
rect 52 10500 1190 10506
rect 52 10103 64 10500
rect 1178 10103 1190 10500
rect 52 10097 1190 10103
rect 1294 10500 2432 10506
rect 1294 10103 1306 10500
rect 2420 10103 2432 10500
rect 1294 10097 2432 10103
rect 2536 10500 3674 10506
rect 2536 10103 2548 10500
rect 3662 10103 3674 10500
rect 2536 10097 3674 10103
rect 3778 10500 4916 10506
rect 3778 10103 3790 10500
rect 4904 10103 4916 10500
rect 3778 10097 4916 10103
rect -4916 9527 -3778 9533
rect -4916 9130 -4904 9527
rect -3790 9130 -3778 9527
rect -4916 9124 -3778 9130
rect -3674 9527 -2536 9533
rect -3674 9130 -3662 9527
rect -2548 9130 -2536 9527
rect -3674 9124 -2536 9130
rect -2432 9527 -1294 9533
rect -2432 9130 -2420 9527
rect -1306 9130 -1294 9527
rect -2432 9124 -1294 9130
rect -1190 9527 -52 9533
rect -1190 9130 -1178 9527
rect -64 9130 -52 9527
rect -1190 9124 -52 9130
rect 52 9527 1190 9533
rect 52 9130 64 9527
rect 1178 9130 1190 9527
rect 52 9124 1190 9130
rect 1294 9527 2432 9533
rect 1294 9130 1306 9527
rect 2420 9130 2432 9527
rect 1294 9124 2432 9130
rect 2536 9527 3674 9533
rect 2536 9130 2548 9527
rect 3662 9130 3674 9527
rect 2536 9124 3674 9130
rect 3778 9527 4916 9533
rect 3778 9130 3790 9527
rect 4904 9130 4916 9527
rect 3778 9124 4916 9130
rect -4916 8990 -3778 8996
rect -4916 8593 -4904 8990
rect -3790 8593 -3778 8990
rect -4916 8587 -3778 8593
rect -3674 8990 -2536 8996
rect -3674 8593 -3662 8990
rect -2548 8593 -2536 8990
rect -3674 8587 -2536 8593
rect -2432 8990 -1294 8996
rect -2432 8593 -2420 8990
rect -1306 8593 -1294 8990
rect -2432 8587 -1294 8593
rect -1190 8990 -52 8996
rect -1190 8593 -1178 8990
rect -64 8593 -52 8990
rect -1190 8587 -52 8593
rect 52 8990 1190 8996
rect 52 8593 64 8990
rect 1178 8593 1190 8990
rect 52 8587 1190 8593
rect 1294 8990 2432 8996
rect 1294 8593 1306 8990
rect 2420 8593 2432 8990
rect 1294 8587 2432 8593
rect 2536 8990 3674 8996
rect 2536 8593 2548 8990
rect 3662 8593 3674 8990
rect 2536 8587 3674 8593
rect 3778 8990 4916 8996
rect 3778 8593 3790 8990
rect 4904 8593 4916 8990
rect 3778 8587 4916 8593
rect -4916 8017 -3778 8023
rect -4916 7620 -4904 8017
rect -3790 7620 -3778 8017
rect -4916 7614 -3778 7620
rect -3674 8017 -2536 8023
rect -3674 7620 -3662 8017
rect -2548 7620 -2536 8017
rect -3674 7614 -2536 7620
rect -2432 8017 -1294 8023
rect -2432 7620 -2420 8017
rect -1306 7620 -1294 8017
rect -2432 7614 -1294 7620
rect -1190 8017 -52 8023
rect -1190 7620 -1178 8017
rect -64 7620 -52 8017
rect -1190 7614 -52 7620
rect 52 8017 1190 8023
rect 52 7620 64 8017
rect 1178 7620 1190 8017
rect 52 7614 1190 7620
rect 1294 8017 2432 8023
rect 1294 7620 1306 8017
rect 2420 7620 2432 8017
rect 1294 7614 2432 7620
rect 2536 8017 3674 8023
rect 2536 7620 2548 8017
rect 3662 7620 3674 8017
rect 2536 7614 3674 7620
rect 3778 8017 4916 8023
rect 3778 7620 3790 8017
rect 4904 7620 4916 8017
rect 3778 7614 4916 7620
rect -4916 7480 -3778 7486
rect -4916 7083 -4904 7480
rect -3790 7083 -3778 7480
rect -4916 7077 -3778 7083
rect -3674 7480 -2536 7486
rect -3674 7083 -3662 7480
rect -2548 7083 -2536 7480
rect -3674 7077 -2536 7083
rect -2432 7480 -1294 7486
rect -2432 7083 -2420 7480
rect -1306 7083 -1294 7480
rect -2432 7077 -1294 7083
rect -1190 7480 -52 7486
rect -1190 7083 -1178 7480
rect -64 7083 -52 7480
rect -1190 7077 -52 7083
rect 52 7480 1190 7486
rect 52 7083 64 7480
rect 1178 7083 1190 7480
rect 52 7077 1190 7083
rect 1294 7480 2432 7486
rect 1294 7083 1306 7480
rect 2420 7083 2432 7480
rect 1294 7077 2432 7083
rect 2536 7480 3674 7486
rect 2536 7083 2548 7480
rect 3662 7083 3674 7480
rect 2536 7077 3674 7083
rect 3778 7480 4916 7486
rect 3778 7083 3790 7480
rect 4904 7083 4916 7480
rect 3778 7077 4916 7083
rect -4916 6507 -3778 6513
rect -4916 6110 -4904 6507
rect -3790 6110 -3778 6507
rect -4916 6104 -3778 6110
rect -3674 6507 -2536 6513
rect -3674 6110 -3662 6507
rect -2548 6110 -2536 6507
rect -3674 6104 -2536 6110
rect -2432 6507 -1294 6513
rect -2432 6110 -2420 6507
rect -1306 6110 -1294 6507
rect -2432 6104 -1294 6110
rect -1190 6507 -52 6513
rect -1190 6110 -1178 6507
rect -64 6110 -52 6507
rect -1190 6104 -52 6110
rect 52 6507 1190 6513
rect 52 6110 64 6507
rect 1178 6110 1190 6507
rect 52 6104 1190 6110
rect 1294 6507 2432 6513
rect 1294 6110 1306 6507
rect 2420 6110 2432 6507
rect 1294 6104 2432 6110
rect 2536 6507 3674 6513
rect 2536 6110 2548 6507
rect 3662 6110 3674 6507
rect 2536 6104 3674 6110
rect 3778 6507 4916 6513
rect 3778 6110 3790 6507
rect 4904 6110 4916 6507
rect 3778 6104 4916 6110
rect -4916 5970 -3778 5976
rect -4916 5573 -4904 5970
rect -3790 5573 -3778 5970
rect -4916 5567 -3778 5573
rect -3674 5970 -2536 5976
rect -3674 5573 -3662 5970
rect -2548 5573 -2536 5970
rect -3674 5567 -2536 5573
rect -2432 5970 -1294 5976
rect -2432 5573 -2420 5970
rect -1306 5573 -1294 5970
rect -2432 5567 -1294 5573
rect -1190 5970 -52 5976
rect -1190 5573 -1178 5970
rect -64 5573 -52 5970
rect -1190 5567 -52 5573
rect 52 5970 1190 5976
rect 52 5573 64 5970
rect 1178 5573 1190 5970
rect 52 5567 1190 5573
rect 1294 5970 2432 5976
rect 1294 5573 1306 5970
rect 2420 5573 2432 5970
rect 1294 5567 2432 5573
rect 2536 5970 3674 5976
rect 2536 5573 2548 5970
rect 3662 5573 3674 5970
rect 2536 5567 3674 5573
rect 3778 5970 4916 5976
rect 3778 5573 3790 5970
rect 4904 5573 4916 5970
rect 3778 5567 4916 5573
rect -4916 4997 -3778 5003
rect -4916 4600 -4904 4997
rect -3790 4600 -3778 4997
rect -4916 4594 -3778 4600
rect -3674 4997 -2536 5003
rect -3674 4600 -3662 4997
rect -2548 4600 -2536 4997
rect -3674 4594 -2536 4600
rect -2432 4997 -1294 5003
rect -2432 4600 -2420 4997
rect -1306 4600 -1294 4997
rect -2432 4594 -1294 4600
rect -1190 4997 -52 5003
rect -1190 4600 -1178 4997
rect -64 4600 -52 4997
rect -1190 4594 -52 4600
rect 52 4997 1190 5003
rect 52 4600 64 4997
rect 1178 4600 1190 4997
rect 52 4594 1190 4600
rect 1294 4997 2432 5003
rect 1294 4600 1306 4997
rect 2420 4600 2432 4997
rect 1294 4594 2432 4600
rect 2536 4997 3674 5003
rect 2536 4600 2548 4997
rect 3662 4600 3674 4997
rect 2536 4594 3674 4600
rect 3778 4997 4916 5003
rect 3778 4600 3790 4997
rect 4904 4600 4916 4997
rect 3778 4594 4916 4600
rect -4916 4460 -3778 4466
rect -4916 4063 -4904 4460
rect -3790 4063 -3778 4460
rect -4916 4057 -3778 4063
rect -3674 4460 -2536 4466
rect -3674 4063 -3662 4460
rect -2548 4063 -2536 4460
rect -3674 4057 -2536 4063
rect -2432 4460 -1294 4466
rect -2432 4063 -2420 4460
rect -1306 4063 -1294 4460
rect -2432 4057 -1294 4063
rect -1190 4460 -52 4466
rect -1190 4063 -1178 4460
rect -64 4063 -52 4460
rect -1190 4057 -52 4063
rect 52 4460 1190 4466
rect 52 4063 64 4460
rect 1178 4063 1190 4460
rect 52 4057 1190 4063
rect 1294 4460 2432 4466
rect 1294 4063 1306 4460
rect 2420 4063 2432 4460
rect 1294 4057 2432 4063
rect 2536 4460 3674 4466
rect 2536 4063 2548 4460
rect 3662 4063 3674 4460
rect 2536 4057 3674 4063
rect 3778 4460 4916 4466
rect 3778 4063 3790 4460
rect 4904 4063 4916 4460
rect 3778 4057 4916 4063
rect -4916 3487 -3778 3493
rect -4916 3090 -4904 3487
rect -3790 3090 -3778 3487
rect -4916 3084 -3778 3090
rect -3674 3487 -2536 3493
rect -3674 3090 -3662 3487
rect -2548 3090 -2536 3487
rect -3674 3084 -2536 3090
rect -2432 3487 -1294 3493
rect -2432 3090 -2420 3487
rect -1306 3090 -1294 3487
rect -2432 3084 -1294 3090
rect -1190 3487 -52 3493
rect -1190 3090 -1178 3487
rect -64 3090 -52 3487
rect -1190 3084 -52 3090
rect 52 3487 1190 3493
rect 52 3090 64 3487
rect 1178 3090 1190 3487
rect 52 3084 1190 3090
rect 1294 3487 2432 3493
rect 1294 3090 1306 3487
rect 2420 3090 2432 3487
rect 1294 3084 2432 3090
rect 2536 3487 3674 3493
rect 2536 3090 2548 3487
rect 3662 3090 3674 3487
rect 2536 3084 3674 3090
rect 3778 3487 4916 3493
rect 3778 3090 3790 3487
rect 4904 3090 4916 3487
rect 3778 3084 4916 3090
rect -4916 2950 -3778 2956
rect -4916 2553 -4904 2950
rect -3790 2553 -3778 2950
rect -4916 2547 -3778 2553
rect -3674 2950 -2536 2956
rect -3674 2553 -3662 2950
rect -2548 2553 -2536 2950
rect -3674 2547 -2536 2553
rect -2432 2950 -1294 2956
rect -2432 2553 -2420 2950
rect -1306 2553 -1294 2950
rect -2432 2547 -1294 2553
rect -1190 2950 -52 2956
rect -1190 2553 -1178 2950
rect -64 2553 -52 2950
rect -1190 2547 -52 2553
rect 52 2950 1190 2956
rect 52 2553 64 2950
rect 1178 2553 1190 2950
rect 52 2547 1190 2553
rect 1294 2950 2432 2956
rect 1294 2553 1306 2950
rect 2420 2553 2432 2950
rect 1294 2547 2432 2553
rect 2536 2950 3674 2956
rect 2536 2553 2548 2950
rect 3662 2553 3674 2950
rect 2536 2547 3674 2553
rect 3778 2950 4916 2956
rect 3778 2553 3790 2950
rect 4904 2553 4916 2950
rect 3778 2547 4916 2553
rect -4916 1977 -3778 1983
rect -4916 1580 -4904 1977
rect -3790 1580 -3778 1977
rect -4916 1574 -3778 1580
rect -3674 1977 -2536 1983
rect -3674 1580 -3662 1977
rect -2548 1580 -2536 1977
rect -3674 1574 -2536 1580
rect -2432 1977 -1294 1983
rect -2432 1580 -2420 1977
rect -1306 1580 -1294 1977
rect -2432 1574 -1294 1580
rect -1190 1977 -52 1983
rect -1190 1580 -1178 1977
rect -64 1580 -52 1977
rect -1190 1574 -52 1580
rect 52 1977 1190 1983
rect 52 1580 64 1977
rect 1178 1580 1190 1977
rect 52 1574 1190 1580
rect 1294 1977 2432 1983
rect 1294 1580 1306 1977
rect 2420 1580 2432 1977
rect 1294 1574 2432 1580
rect 2536 1977 3674 1983
rect 2536 1580 2548 1977
rect 3662 1580 3674 1977
rect 2536 1574 3674 1580
rect 3778 1977 4916 1983
rect 3778 1580 3790 1977
rect 4904 1580 4916 1977
rect 3778 1574 4916 1580
rect -4916 1440 -3778 1446
rect -4916 1043 -4904 1440
rect -3790 1043 -3778 1440
rect -4916 1037 -3778 1043
rect -3674 1440 -2536 1446
rect -3674 1043 -3662 1440
rect -2548 1043 -2536 1440
rect -3674 1037 -2536 1043
rect -2432 1440 -1294 1446
rect -2432 1043 -2420 1440
rect -1306 1043 -1294 1440
rect -2432 1037 -1294 1043
rect -1190 1440 -52 1446
rect -1190 1043 -1178 1440
rect -64 1043 -52 1440
rect -1190 1037 -52 1043
rect 52 1440 1190 1446
rect 52 1043 64 1440
rect 1178 1043 1190 1440
rect 52 1037 1190 1043
rect 1294 1440 2432 1446
rect 1294 1043 1306 1440
rect 2420 1043 2432 1440
rect 1294 1037 2432 1043
rect 2536 1440 3674 1446
rect 2536 1043 2548 1440
rect 3662 1043 3674 1440
rect 2536 1037 3674 1043
rect 3778 1440 4916 1446
rect 3778 1043 3790 1440
rect 4904 1043 4916 1440
rect 3778 1037 4916 1043
rect -4916 467 -3778 473
rect -4916 70 -4904 467
rect -3790 70 -3778 467
rect -4916 64 -3778 70
rect -3674 467 -2536 473
rect -3674 70 -3662 467
rect -2548 70 -2536 467
rect -3674 64 -2536 70
rect -2432 467 -1294 473
rect -2432 70 -2420 467
rect -1306 70 -1294 467
rect -2432 64 -1294 70
rect -1190 467 -52 473
rect -1190 70 -1178 467
rect -64 70 -52 467
rect -1190 64 -52 70
rect 52 467 1190 473
rect 52 70 64 467
rect 1178 70 1190 467
rect 52 64 1190 70
rect 1294 467 2432 473
rect 1294 70 1306 467
rect 2420 70 2432 467
rect 1294 64 2432 70
rect 2536 467 3674 473
rect 2536 70 2548 467
rect 3662 70 3674 467
rect 2536 64 3674 70
rect 3778 467 4916 473
rect 3778 70 3790 467
rect 4904 70 4916 467
rect 3778 64 4916 70
rect -4916 -70 -3778 -64
rect -4916 -467 -4904 -70
rect -3790 -467 -3778 -70
rect -4916 -473 -3778 -467
rect -3674 -70 -2536 -64
rect -3674 -467 -3662 -70
rect -2548 -467 -2536 -70
rect -3674 -473 -2536 -467
rect -2432 -70 -1294 -64
rect -2432 -467 -2420 -70
rect -1306 -467 -1294 -70
rect -2432 -473 -1294 -467
rect -1190 -70 -52 -64
rect -1190 -467 -1178 -70
rect -64 -467 -52 -70
rect -1190 -473 -52 -467
rect 52 -70 1190 -64
rect 52 -467 64 -70
rect 1178 -467 1190 -70
rect 52 -473 1190 -467
rect 1294 -70 2432 -64
rect 1294 -467 1306 -70
rect 2420 -467 2432 -70
rect 1294 -473 2432 -467
rect 2536 -70 3674 -64
rect 2536 -467 2548 -70
rect 3662 -467 3674 -70
rect 2536 -473 3674 -467
rect 3778 -70 4916 -64
rect 3778 -467 3790 -70
rect 4904 -467 4916 -70
rect 3778 -473 4916 -467
rect -4916 -1043 -3778 -1037
rect -4916 -1440 -4904 -1043
rect -3790 -1440 -3778 -1043
rect -4916 -1446 -3778 -1440
rect -3674 -1043 -2536 -1037
rect -3674 -1440 -3662 -1043
rect -2548 -1440 -2536 -1043
rect -3674 -1446 -2536 -1440
rect -2432 -1043 -1294 -1037
rect -2432 -1440 -2420 -1043
rect -1306 -1440 -1294 -1043
rect -2432 -1446 -1294 -1440
rect -1190 -1043 -52 -1037
rect -1190 -1440 -1178 -1043
rect -64 -1440 -52 -1043
rect -1190 -1446 -52 -1440
rect 52 -1043 1190 -1037
rect 52 -1440 64 -1043
rect 1178 -1440 1190 -1043
rect 52 -1446 1190 -1440
rect 1294 -1043 2432 -1037
rect 1294 -1440 1306 -1043
rect 2420 -1440 2432 -1043
rect 1294 -1446 2432 -1440
rect 2536 -1043 3674 -1037
rect 2536 -1440 2548 -1043
rect 3662 -1440 3674 -1043
rect 2536 -1446 3674 -1440
rect 3778 -1043 4916 -1037
rect 3778 -1440 3790 -1043
rect 4904 -1440 4916 -1043
rect 3778 -1446 4916 -1440
rect -4916 -1580 -3778 -1574
rect -4916 -1977 -4904 -1580
rect -3790 -1977 -3778 -1580
rect -4916 -1983 -3778 -1977
rect -3674 -1580 -2536 -1574
rect -3674 -1977 -3662 -1580
rect -2548 -1977 -2536 -1580
rect -3674 -1983 -2536 -1977
rect -2432 -1580 -1294 -1574
rect -2432 -1977 -2420 -1580
rect -1306 -1977 -1294 -1580
rect -2432 -1983 -1294 -1977
rect -1190 -1580 -52 -1574
rect -1190 -1977 -1178 -1580
rect -64 -1977 -52 -1580
rect -1190 -1983 -52 -1977
rect 52 -1580 1190 -1574
rect 52 -1977 64 -1580
rect 1178 -1977 1190 -1580
rect 52 -1983 1190 -1977
rect 1294 -1580 2432 -1574
rect 1294 -1977 1306 -1580
rect 2420 -1977 2432 -1580
rect 1294 -1983 2432 -1977
rect 2536 -1580 3674 -1574
rect 2536 -1977 2548 -1580
rect 3662 -1977 3674 -1580
rect 2536 -1983 3674 -1977
rect 3778 -1580 4916 -1574
rect 3778 -1977 3790 -1580
rect 4904 -1977 4916 -1580
rect 3778 -1983 4916 -1977
rect -4916 -2553 -3778 -2547
rect -4916 -2950 -4904 -2553
rect -3790 -2950 -3778 -2553
rect -4916 -2956 -3778 -2950
rect -3674 -2553 -2536 -2547
rect -3674 -2950 -3662 -2553
rect -2548 -2950 -2536 -2553
rect -3674 -2956 -2536 -2950
rect -2432 -2553 -1294 -2547
rect -2432 -2950 -2420 -2553
rect -1306 -2950 -1294 -2553
rect -2432 -2956 -1294 -2950
rect -1190 -2553 -52 -2547
rect -1190 -2950 -1178 -2553
rect -64 -2950 -52 -2553
rect -1190 -2956 -52 -2950
rect 52 -2553 1190 -2547
rect 52 -2950 64 -2553
rect 1178 -2950 1190 -2553
rect 52 -2956 1190 -2950
rect 1294 -2553 2432 -2547
rect 1294 -2950 1306 -2553
rect 2420 -2950 2432 -2553
rect 1294 -2956 2432 -2950
rect 2536 -2553 3674 -2547
rect 2536 -2950 2548 -2553
rect 3662 -2950 3674 -2553
rect 2536 -2956 3674 -2950
rect 3778 -2553 4916 -2547
rect 3778 -2950 3790 -2553
rect 4904 -2950 4916 -2553
rect 3778 -2956 4916 -2950
rect -4916 -3090 -3778 -3084
rect -4916 -3487 -4904 -3090
rect -3790 -3487 -3778 -3090
rect -4916 -3493 -3778 -3487
rect -3674 -3090 -2536 -3084
rect -3674 -3487 -3662 -3090
rect -2548 -3487 -2536 -3090
rect -3674 -3493 -2536 -3487
rect -2432 -3090 -1294 -3084
rect -2432 -3487 -2420 -3090
rect -1306 -3487 -1294 -3090
rect -2432 -3493 -1294 -3487
rect -1190 -3090 -52 -3084
rect -1190 -3487 -1178 -3090
rect -64 -3487 -52 -3090
rect -1190 -3493 -52 -3487
rect 52 -3090 1190 -3084
rect 52 -3487 64 -3090
rect 1178 -3487 1190 -3090
rect 52 -3493 1190 -3487
rect 1294 -3090 2432 -3084
rect 1294 -3487 1306 -3090
rect 2420 -3487 2432 -3090
rect 1294 -3493 2432 -3487
rect 2536 -3090 3674 -3084
rect 2536 -3487 2548 -3090
rect 3662 -3487 3674 -3090
rect 2536 -3493 3674 -3487
rect 3778 -3090 4916 -3084
rect 3778 -3487 3790 -3090
rect 4904 -3487 4916 -3090
rect 3778 -3493 4916 -3487
rect -4916 -4063 -3778 -4057
rect -4916 -4460 -4904 -4063
rect -3790 -4460 -3778 -4063
rect -4916 -4466 -3778 -4460
rect -3674 -4063 -2536 -4057
rect -3674 -4460 -3662 -4063
rect -2548 -4460 -2536 -4063
rect -3674 -4466 -2536 -4460
rect -2432 -4063 -1294 -4057
rect -2432 -4460 -2420 -4063
rect -1306 -4460 -1294 -4063
rect -2432 -4466 -1294 -4460
rect -1190 -4063 -52 -4057
rect -1190 -4460 -1178 -4063
rect -64 -4460 -52 -4063
rect -1190 -4466 -52 -4460
rect 52 -4063 1190 -4057
rect 52 -4460 64 -4063
rect 1178 -4460 1190 -4063
rect 52 -4466 1190 -4460
rect 1294 -4063 2432 -4057
rect 1294 -4460 1306 -4063
rect 2420 -4460 2432 -4063
rect 1294 -4466 2432 -4460
rect 2536 -4063 3674 -4057
rect 2536 -4460 2548 -4063
rect 3662 -4460 3674 -4063
rect 2536 -4466 3674 -4460
rect 3778 -4063 4916 -4057
rect 3778 -4460 3790 -4063
rect 4904 -4460 4916 -4063
rect 3778 -4466 4916 -4460
rect -4916 -4600 -3778 -4594
rect -4916 -4997 -4904 -4600
rect -3790 -4997 -3778 -4600
rect -4916 -5003 -3778 -4997
rect -3674 -4600 -2536 -4594
rect -3674 -4997 -3662 -4600
rect -2548 -4997 -2536 -4600
rect -3674 -5003 -2536 -4997
rect -2432 -4600 -1294 -4594
rect -2432 -4997 -2420 -4600
rect -1306 -4997 -1294 -4600
rect -2432 -5003 -1294 -4997
rect -1190 -4600 -52 -4594
rect -1190 -4997 -1178 -4600
rect -64 -4997 -52 -4600
rect -1190 -5003 -52 -4997
rect 52 -4600 1190 -4594
rect 52 -4997 64 -4600
rect 1178 -4997 1190 -4600
rect 52 -5003 1190 -4997
rect 1294 -4600 2432 -4594
rect 1294 -4997 1306 -4600
rect 2420 -4997 2432 -4600
rect 1294 -5003 2432 -4997
rect 2536 -4600 3674 -4594
rect 2536 -4997 2548 -4600
rect 3662 -4997 3674 -4600
rect 2536 -5003 3674 -4997
rect 3778 -4600 4916 -4594
rect 3778 -4997 3790 -4600
rect 4904 -4997 4916 -4600
rect 3778 -5003 4916 -4997
rect -4916 -5573 -3778 -5567
rect -4916 -5970 -4904 -5573
rect -3790 -5970 -3778 -5573
rect -4916 -5976 -3778 -5970
rect -3674 -5573 -2536 -5567
rect -3674 -5970 -3662 -5573
rect -2548 -5970 -2536 -5573
rect -3674 -5976 -2536 -5970
rect -2432 -5573 -1294 -5567
rect -2432 -5970 -2420 -5573
rect -1306 -5970 -1294 -5573
rect -2432 -5976 -1294 -5970
rect -1190 -5573 -52 -5567
rect -1190 -5970 -1178 -5573
rect -64 -5970 -52 -5573
rect -1190 -5976 -52 -5970
rect 52 -5573 1190 -5567
rect 52 -5970 64 -5573
rect 1178 -5970 1190 -5573
rect 52 -5976 1190 -5970
rect 1294 -5573 2432 -5567
rect 1294 -5970 1306 -5573
rect 2420 -5970 2432 -5573
rect 1294 -5976 2432 -5970
rect 2536 -5573 3674 -5567
rect 2536 -5970 2548 -5573
rect 3662 -5970 3674 -5573
rect 2536 -5976 3674 -5970
rect 3778 -5573 4916 -5567
rect 3778 -5970 3790 -5573
rect 4904 -5970 4916 -5573
rect 3778 -5976 4916 -5970
rect -4916 -6110 -3778 -6104
rect -4916 -6507 -4904 -6110
rect -3790 -6507 -3778 -6110
rect -4916 -6513 -3778 -6507
rect -3674 -6110 -2536 -6104
rect -3674 -6507 -3662 -6110
rect -2548 -6507 -2536 -6110
rect -3674 -6513 -2536 -6507
rect -2432 -6110 -1294 -6104
rect -2432 -6507 -2420 -6110
rect -1306 -6507 -1294 -6110
rect -2432 -6513 -1294 -6507
rect -1190 -6110 -52 -6104
rect -1190 -6507 -1178 -6110
rect -64 -6507 -52 -6110
rect -1190 -6513 -52 -6507
rect 52 -6110 1190 -6104
rect 52 -6507 64 -6110
rect 1178 -6507 1190 -6110
rect 52 -6513 1190 -6507
rect 1294 -6110 2432 -6104
rect 1294 -6507 1306 -6110
rect 2420 -6507 2432 -6110
rect 1294 -6513 2432 -6507
rect 2536 -6110 3674 -6104
rect 2536 -6507 2548 -6110
rect 3662 -6507 3674 -6110
rect 2536 -6513 3674 -6507
rect 3778 -6110 4916 -6104
rect 3778 -6507 3790 -6110
rect 4904 -6507 4916 -6110
rect 3778 -6513 4916 -6507
rect -4916 -7083 -3778 -7077
rect -4916 -7480 -4904 -7083
rect -3790 -7480 -3778 -7083
rect -4916 -7486 -3778 -7480
rect -3674 -7083 -2536 -7077
rect -3674 -7480 -3662 -7083
rect -2548 -7480 -2536 -7083
rect -3674 -7486 -2536 -7480
rect -2432 -7083 -1294 -7077
rect -2432 -7480 -2420 -7083
rect -1306 -7480 -1294 -7083
rect -2432 -7486 -1294 -7480
rect -1190 -7083 -52 -7077
rect -1190 -7480 -1178 -7083
rect -64 -7480 -52 -7083
rect -1190 -7486 -52 -7480
rect 52 -7083 1190 -7077
rect 52 -7480 64 -7083
rect 1178 -7480 1190 -7083
rect 52 -7486 1190 -7480
rect 1294 -7083 2432 -7077
rect 1294 -7480 1306 -7083
rect 2420 -7480 2432 -7083
rect 1294 -7486 2432 -7480
rect 2536 -7083 3674 -7077
rect 2536 -7480 2548 -7083
rect 3662 -7480 3674 -7083
rect 2536 -7486 3674 -7480
rect 3778 -7083 4916 -7077
rect 3778 -7480 3790 -7083
rect 4904 -7480 4916 -7083
rect 3778 -7486 4916 -7480
rect -4916 -7620 -3778 -7614
rect -4916 -8017 -4904 -7620
rect -3790 -8017 -3778 -7620
rect -4916 -8023 -3778 -8017
rect -3674 -7620 -2536 -7614
rect -3674 -8017 -3662 -7620
rect -2548 -8017 -2536 -7620
rect -3674 -8023 -2536 -8017
rect -2432 -7620 -1294 -7614
rect -2432 -8017 -2420 -7620
rect -1306 -8017 -1294 -7620
rect -2432 -8023 -1294 -8017
rect -1190 -7620 -52 -7614
rect -1190 -8017 -1178 -7620
rect -64 -8017 -52 -7620
rect -1190 -8023 -52 -8017
rect 52 -7620 1190 -7614
rect 52 -8017 64 -7620
rect 1178 -8017 1190 -7620
rect 52 -8023 1190 -8017
rect 1294 -7620 2432 -7614
rect 1294 -8017 1306 -7620
rect 2420 -8017 2432 -7620
rect 1294 -8023 2432 -8017
rect 2536 -7620 3674 -7614
rect 2536 -8017 2548 -7620
rect 3662 -8017 3674 -7620
rect 2536 -8023 3674 -8017
rect 3778 -7620 4916 -7614
rect 3778 -8017 3790 -7620
rect 4904 -8017 4916 -7620
rect 3778 -8023 4916 -8017
rect -4916 -8593 -3778 -8587
rect -4916 -8990 -4904 -8593
rect -3790 -8990 -3778 -8593
rect -4916 -8996 -3778 -8990
rect -3674 -8593 -2536 -8587
rect -3674 -8990 -3662 -8593
rect -2548 -8990 -2536 -8593
rect -3674 -8996 -2536 -8990
rect -2432 -8593 -1294 -8587
rect -2432 -8990 -2420 -8593
rect -1306 -8990 -1294 -8593
rect -2432 -8996 -1294 -8990
rect -1190 -8593 -52 -8587
rect -1190 -8990 -1178 -8593
rect -64 -8990 -52 -8593
rect -1190 -8996 -52 -8990
rect 52 -8593 1190 -8587
rect 52 -8990 64 -8593
rect 1178 -8990 1190 -8593
rect 52 -8996 1190 -8990
rect 1294 -8593 2432 -8587
rect 1294 -8990 1306 -8593
rect 2420 -8990 2432 -8593
rect 1294 -8996 2432 -8990
rect 2536 -8593 3674 -8587
rect 2536 -8990 2548 -8593
rect 3662 -8990 3674 -8593
rect 2536 -8996 3674 -8990
rect 3778 -8593 4916 -8587
rect 3778 -8990 3790 -8593
rect 4904 -8990 4916 -8593
rect 3778 -8996 4916 -8990
rect -4916 -9130 -3778 -9124
rect -4916 -9527 -4904 -9130
rect -3790 -9527 -3778 -9130
rect -4916 -9533 -3778 -9527
rect -3674 -9130 -2536 -9124
rect -3674 -9527 -3662 -9130
rect -2548 -9527 -2536 -9130
rect -3674 -9533 -2536 -9527
rect -2432 -9130 -1294 -9124
rect -2432 -9527 -2420 -9130
rect -1306 -9527 -1294 -9130
rect -2432 -9533 -1294 -9527
rect -1190 -9130 -52 -9124
rect -1190 -9527 -1178 -9130
rect -64 -9527 -52 -9130
rect -1190 -9533 -52 -9527
rect 52 -9130 1190 -9124
rect 52 -9527 64 -9130
rect 1178 -9527 1190 -9130
rect 52 -9533 1190 -9527
rect 1294 -9130 2432 -9124
rect 1294 -9527 1306 -9130
rect 2420 -9527 2432 -9130
rect 1294 -9533 2432 -9527
rect 2536 -9130 3674 -9124
rect 2536 -9527 2548 -9130
rect 3662 -9527 3674 -9130
rect 2536 -9533 3674 -9527
rect 3778 -9130 4916 -9124
rect 3778 -9527 3790 -9130
rect 4904 -9527 4916 -9130
rect 3778 -9533 4916 -9527
rect -4916 -10103 -3778 -10097
rect -4916 -10500 -4904 -10103
rect -3790 -10500 -3778 -10103
rect -4916 -10506 -3778 -10500
rect -3674 -10103 -2536 -10097
rect -3674 -10500 -3662 -10103
rect -2548 -10500 -2536 -10103
rect -3674 -10506 -2536 -10500
rect -2432 -10103 -1294 -10097
rect -2432 -10500 -2420 -10103
rect -1306 -10500 -1294 -10103
rect -2432 -10506 -1294 -10500
rect -1190 -10103 -52 -10097
rect -1190 -10500 -1178 -10103
rect -64 -10500 -52 -10103
rect -1190 -10506 -52 -10500
rect 52 -10103 1190 -10097
rect 52 -10500 64 -10103
rect 1178 -10500 1190 -10103
rect 52 -10506 1190 -10500
rect 1294 -10103 2432 -10097
rect 1294 -10500 1306 -10103
rect 2420 -10500 2432 -10103
rect 1294 -10506 2432 -10500
rect 2536 -10103 3674 -10097
rect 2536 -10500 2548 -10103
rect 3662 -10500 3674 -10103
rect 2536 -10506 3674 -10500
rect 3778 -10103 4916 -10097
rect 3778 -10500 3790 -10103
rect 4904 -10500 4916 -10103
rect 3778 -10506 4916 -10500
rect -4916 -10640 -3778 -10634
rect -4916 -11037 -4904 -10640
rect -3790 -11037 -3778 -10640
rect -4916 -11043 -3778 -11037
rect -3674 -10640 -2536 -10634
rect -3674 -11037 -3662 -10640
rect -2548 -11037 -2536 -10640
rect -3674 -11043 -2536 -11037
rect -2432 -10640 -1294 -10634
rect -2432 -11037 -2420 -10640
rect -1306 -11037 -1294 -10640
rect -2432 -11043 -1294 -11037
rect -1190 -10640 -52 -10634
rect -1190 -11037 -1178 -10640
rect -64 -11037 -52 -10640
rect -1190 -11043 -52 -11037
rect 52 -10640 1190 -10634
rect 52 -11037 64 -10640
rect 1178 -11037 1190 -10640
rect 52 -11043 1190 -11037
rect 1294 -10640 2432 -10634
rect 1294 -11037 1306 -10640
rect 2420 -11037 2432 -10640
rect 1294 -11043 2432 -11037
rect 2536 -10640 3674 -10634
rect 2536 -11037 2548 -10640
rect 3662 -11037 3674 -10640
rect 2536 -11043 3674 -11037
rect 3778 -10640 4916 -10634
rect 3778 -11037 3790 -10640
rect 4904 -11037 4916 -10640
rect 3778 -11043 4916 -11037
rect -4916 -11613 -3778 -11607
rect -4916 -12010 -4904 -11613
rect -3790 -12010 -3778 -11613
rect -4916 -12016 -3778 -12010
rect -3674 -11613 -2536 -11607
rect -3674 -12010 -3662 -11613
rect -2548 -12010 -2536 -11613
rect -3674 -12016 -2536 -12010
rect -2432 -11613 -1294 -11607
rect -2432 -12010 -2420 -11613
rect -1306 -12010 -1294 -11613
rect -2432 -12016 -1294 -12010
rect -1190 -11613 -52 -11607
rect -1190 -12010 -1178 -11613
rect -64 -12010 -52 -11613
rect -1190 -12016 -52 -12010
rect 52 -11613 1190 -11607
rect 52 -12010 64 -11613
rect 1178 -12010 1190 -11613
rect 52 -12016 1190 -12010
rect 1294 -11613 2432 -11607
rect 1294 -12010 1306 -11613
rect 2420 -12010 2432 -11613
rect 1294 -12016 2432 -12010
rect 2536 -11613 3674 -11607
rect 2536 -12010 2548 -11613
rect 3662 -12010 3674 -11613
rect 2536 -12016 3674 -12010
rect 3778 -11613 4916 -11607
rect 3778 -12010 3790 -11613
rect 4904 -12010 4916 -11613
rect 3778 -12016 4916 -12010
rect -4916 -12150 -3778 -12144
rect -4916 -12547 -4904 -12150
rect -3790 -12547 -3778 -12150
rect -4916 -12553 -3778 -12547
rect -3674 -12150 -2536 -12144
rect -3674 -12547 -3662 -12150
rect -2548 -12547 -2536 -12150
rect -3674 -12553 -2536 -12547
rect -2432 -12150 -1294 -12144
rect -2432 -12547 -2420 -12150
rect -1306 -12547 -1294 -12150
rect -2432 -12553 -1294 -12547
rect -1190 -12150 -52 -12144
rect -1190 -12547 -1178 -12150
rect -64 -12547 -52 -12150
rect -1190 -12553 -52 -12547
rect 52 -12150 1190 -12144
rect 52 -12547 64 -12150
rect 1178 -12547 1190 -12150
rect 52 -12553 1190 -12547
rect 1294 -12150 2432 -12144
rect 1294 -12547 1306 -12150
rect 2420 -12547 2432 -12150
rect 1294 -12553 2432 -12547
rect 2536 -12150 3674 -12144
rect 2536 -12547 2548 -12150
rect 3662 -12547 3674 -12150
rect 2536 -12553 3674 -12547
rect 3778 -12150 4916 -12144
rect 3778 -12547 3790 -12150
rect 4904 -12547 4916 -12150
rect 3778 -12553 4916 -12547
rect -4916 -13123 -3778 -13117
rect -4916 -13520 -4904 -13123
rect -3790 -13520 -3778 -13123
rect -4916 -13526 -3778 -13520
rect -3674 -13123 -2536 -13117
rect -3674 -13520 -3662 -13123
rect -2548 -13520 -2536 -13123
rect -3674 -13526 -2536 -13520
rect -2432 -13123 -1294 -13117
rect -2432 -13520 -2420 -13123
rect -1306 -13520 -1294 -13123
rect -2432 -13526 -1294 -13520
rect -1190 -13123 -52 -13117
rect -1190 -13520 -1178 -13123
rect -64 -13520 -52 -13123
rect -1190 -13526 -52 -13520
rect 52 -13123 1190 -13117
rect 52 -13520 64 -13123
rect 1178 -13520 1190 -13123
rect 52 -13526 1190 -13520
rect 1294 -13123 2432 -13117
rect 1294 -13520 1306 -13123
rect 2420 -13520 2432 -13123
rect 1294 -13526 2432 -13520
rect 2536 -13123 3674 -13117
rect 2536 -13520 2548 -13123
rect 3662 -13520 3674 -13123
rect 2536 -13526 3674 -13520
rect 3778 -13123 4916 -13117
rect 3778 -13520 3790 -13123
rect 4904 -13520 4916 -13123
rect 3778 -13526 4916 -13520
<< properties >>
string FIXED_BBOX -5033 -13651 5033 13651
string gencell sky130_fd_pr__res_xhigh_po_5p73
string library sky130
string parameters w 5.73 l 2.865 m 18 nx 8 wmin 5.730 lmin 0.50 rho 2000 val 1.065k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 5.730 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
