magic
tech sky130A
magscale 1 2
timestamp 1714103463
<< locali >>
rect 6430 -1047 6432 -174
rect 6430 -1117 6431 -1047
<< viali >>
rect 2276 483 2326 4213
rect 2776 473 2826 4213
rect -2490 -80 6480 -20
rect 6430 -174 6480 -80
rect 6432 -1047 6480 -174
rect 6431 -1117 6480 -1047
rect 6430 -1152 6480 -1117
rect -2482 -1200 6480 -1152
rect -2482 -1212 6470 -1200
rect -2510 -1320 15790 -1260
rect -2510 -2640 -2440 -1320
rect 15700 -2640 15790 -1320
rect -2510 -2700 15794 -2640
rect -2510 -3990 -2440 -2700
rect 15700 -3990 15790 -2700
rect -2510 -4080 15800 -3990
<< metal1 >>
rect 2416 4620 2736 4693
rect 2416 4493 2460 4620
rect 2450 4490 2460 4493
rect 2690 4493 2736 4620
rect 2690 4490 2700 4493
rect 1956 4293 3146 4373
rect 1866 4227 1956 4243
rect 1864 473 1874 4227
rect 1948 473 1958 4227
rect 2166 4213 2446 4243
rect 2166 4133 2276 4213
rect 2326 4133 2446 4213
rect 2166 623 2256 4133
rect 2346 623 2446 4133
rect 2166 483 2276 623
rect 2326 483 2446 623
rect 1866 443 1956 473
rect 2166 453 2446 483
rect 2626 403 2716 4293
rect 2776 4225 2926 4243
rect 2770 4213 2926 4225
rect 2770 473 2776 4213
rect 2826 4133 2926 4213
rect 2886 623 2926 4133
rect 2826 473 2926 623
rect 2770 461 2926 473
rect 3130 470 3140 4230
rect 3210 470 3220 4230
rect 5800 670 6610 720
rect 5790 470 5800 670
rect 6260 470 6610 670
rect 2776 443 2926 461
rect 5800 460 6610 470
rect 1956 400 3146 403
rect 1450 330 2140 400
rect 2980 330 3146 400
rect 1450 323 3146 330
rect 1450 320 2050 323
rect 1450 180 1510 320
rect 1350 140 1510 180
rect 1450 80 1510 140
rect 1320 20 1330 80
rect 1410 20 1420 80
rect 6424 -14 6486 -8
rect -2502 -20 6492 -14
rect -2502 -80 -2490 -20
rect -2502 -86 6430 -80
rect -2450 -130 6100 -120
rect -2520 -180 6100 -130
rect -2520 -1050 -2450 -180
rect 1880 -210 1950 -180
rect -2413 -1004 -2403 -227
rect -2344 -1004 -2334 -227
rect -2210 -1005 -2200 -228
rect -2141 -1005 -2131 -228
rect -2007 -1004 -1997 -227
rect -1938 -1004 -1928 -227
rect -1804 -1005 -1794 -228
rect -1735 -1005 -1725 -228
rect -1601 -1004 -1591 -227
rect -1532 -1004 -1522 -227
rect -1398 -1005 -1388 -228
rect -1329 -1005 -1319 -228
rect -1195 -1004 -1185 -227
rect -1126 -1004 -1116 -227
rect -992 -1005 -982 -228
rect -923 -1005 -913 -228
rect -789 -1004 -779 -227
rect -720 -1004 -710 -227
rect -586 -1005 -576 -228
rect -517 -1005 -507 -228
rect -383 -1004 -373 -227
rect -314 -1004 -304 -227
rect -180 -1005 -170 -228
rect -111 -1005 -101 -228
rect 23 -1004 33 -227
rect 92 -1004 102 -227
rect 226 -1005 236 -228
rect 295 -1005 305 -228
rect 429 -1004 439 -227
rect 498 -1004 508 -227
rect 632 -1005 642 -228
rect 701 -1005 711 -228
rect 835 -1004 845 -227
rect 904 -1004 914 -227
rect 1038 -1005 1048 -228
rect 1107 -1005 1117 -228
rect 1241 -1004 1251 -227
rect 1310 -1004 1320 -227
rect 1444 -1005 1454 -228
rect 1513 -1005 1523 -228
rect 1647 -250 1726 -227
rect 1860 -228 1950 -210
rect 1640 -940 1650 -250
rect 1710 -940 1726 -250
rect 1647 -1004 1726 -940
rect 1850 -249 1950 -228
rect 1850 -939 1871 -249
rect 1931 -939 1950 -249
rect 1850 -1005 1950 -939
rect 2053 -1004 2063 -227
rect 2122 -1004 2132 -227
rect 2256 -1005 2266 -228
rect 2325 -1005 2335 -228
rect 2459 -1004 2469 -227
rect 2528 -1004 2538 -227
rect 2662 -1005 2672 -228
rect 2731 -1005 2741 -228
rect 2865 -1004 2875 -227
rect 2934 -1004 2944 -227
rect 3068 -1005 3078 -228
rect 3137 -1005 3147 -228
rect 3271 -1004 3281 -227
rect 3340 -1004 3350 -227
rect 3474 -1005 3484 -228
rect 3543 -1005 3553 -228
rect 3677 -1004 3687 -227
rect 3746 -1004 3756 -227
rect 3880 -1005 3890 -228
rect 3949 -1005 3959 -228
rect 4083 -1004 4093 -227
rect 4152 -1004 4162 -227
rect 4286 -1005 4296 -228
rect 4355 -1005 4365 -228
rect 4489 -1004 4499 -227
rect 4558 -1004 4568 -227
rect 4692 -1005 4702 -228
rect 4761 -1005 4771 -228
rect 4895 -1004 4905 -227
rect 4964 -1004 4974 -227
rect 5098 -1005 5108 -228
rect 5167 -1005 5177 -228
rect 5301 -1004 5311 -227
rect 5370 -1004 5380 -227
rect 5504 -1005 5514 -228
rect 5573 -1005 5583 -228
rect 5707 -1004 5717 -227
rect 5776 -1004 5786 -227
rect 5910 -1005 5920 -228
rect 5979 -1005 5989 -228
rect 1860 -1020 1950 -1005
rect 1880 -1050 1950 -1020
rect -2520 -1051 5910 -1050
rect 6030 -1051 6100 -180
rect -2520 -1110 6100 -1051
rect 6150 -190 6160 -120
rect 6280 -174 6320 -120
rect 6424 -174 6430 -86
rect 6480 -86 6492 -20
rect 6480 -160 6486 -86
rect 6280 -180 6316 -174
rect 6280 -190 6290 -180
rect 6150 -1050 6210 -190
rect 6424 -234 6432 -174
rect 6329 -266 6364 -234
rect 6423 -266 6432 -234
rect 6329 -934 6432 -266
rect 6329 -1002 6364 -934
rect 6329 -1004 6359 -1002
rect 6423 -1047 6432 -934
rect 6150 -1080 6240 -1050
rect 6423 -1117 6431 -1047
rect 6423 -1146 6430 -1117
rect -2494 -1152 6430 -1146
rect -2494 -1212 -2482 -1152
rect 6480 -1200 15800 -160
rect 6470 -1212 15800 -1200
rect -2494 -1218 1640 -1212
rect -2490 -1248 1640 -1218
rect -2516 -1260 1640 -1248
rect 1740 -1260 15800 -1212
rect -2516 -3984 -2510 -1260
rect -2440 -1326 15700 -1320
rect -2440 -2634 -2434 -1326
rect -2360 -2540 -2350 -1430
rect -1940 -2540 -1930 -1430
rect 15230 -2634 15700 -1326
rect -2440 -2640 15700 -2634
rect 15790 -1326 15800 -1260
rect 15790 -2634 15796 -1326
rect 15790 -2640 15806 -2634
rect 15794 -2700 15806 -2640
rect -2522 -4080 -2510 -3984
rect -2440 -2706 15700 -2700
rect -2440 -3984 -2434 -2706
rect -2360 -3920 -2350 -2810
rect -1940 -3920 -1930 -2810
rect 15230 -3984 15700 -2706
rect -2440 -3990 15700 -3984
rect 15790 -2706 15806 -2700
rect 15790 -3984 15796 -2706
rect 15790 -3990 15812 -3984
rect 15800 -4080 15812 -3990
rect -2522 -4086 15812 -4080
<< via1 >>
rect 2460 4490 2690 4620
rect 1874 473 1948 4227
rect 2256 623 2276 4133
rect 2276 623 2326 4133
rect 2326 623 2346 4133
rect 2796 623 2826 4133
rect 2826 623 2886 4133
rect 3140 470 3210 4230
rect 5800 470 6260 670
rect 2140 330 2980 400
rect 1330 20 1410 80
rect -2403 -1004 -2344 -227
rect -2200 -1005 -2141 -228
rect -1997 -1004 -1938 -227
rect -1794 -1005 -1735 -228
rect -1591 -1004 -1532 -227
rect -1388 -1005 -1329 -228
rect -1185 -1004 -1126 -227
rect -982 -1005 -923 -228
rect -779 -1004 -720 -227
rect -576 -1005 -517 -228
rect -373 -1004 -314 -227
rect -170 -1005 -111 -228
rect 33 -1004 92 -227
rect 236 -1005 295 -228
rect 439 -1004 498 -227
rect 642 -1005 701 -228
rect 845 -1004 904 -227
rect 1048 -1005 1107 -228
rect 1251 -1004 1310 -227
rect 1454 -1005 1513 -228
rect 1650 -940 1710 -250
rect 1871 -939 1931 -249
rect 2063 -1004 2122 -227
rect 2266 -1005 2325 -228
rect 2469 -1004 2528 -227
rect 2672 -1005 2731 -228
rect 2875 -1004 2934 -227
rect 3078 -1005 3137 -228
rect 3281 -1004 3340 -227
rect 3484 -1005 3543 -228
rect 3687 -1004 3746 -227
rect 3890 -1005 3949 -228
rect 4093 -1004 4152 -227
rect 4296 -1005 4355 -228
rect 4499 -1004 4558 -227
rect 4702 -1005 4761 -228
rect 4905 -1004 4964 -227
rect 5108 -1005 5167 -228
rect 5311 -1004 5370 -227
rect 5514 -1005 5573 -228
rect 5717 -1004 5776 -227
rect 5920 -1005 5979 -228
rect 6160 -190 6280 -120
rect 1640 -1212 1740 -1210
rect 1640 -1260 1740 -1212
rect 1640 -1290 1740 -1260
rect -2350 -2540 -1940 -1430
rect -2350 -3920 -1940 -2810
<< metal2 >>
rect 2226 4620 2926 4633
rect 2226 4490 2460 4620
rect 2690 4490 2926 4620
rect 2226 4423 2926 4490
rect 1874 4227 1948 4237
rect 2226 4133 2376 4423
rect 2226 4073 2256 4133
rect 2346 4073 2376 4133
rect 2786 4133 2926 4423
rect 2786 4073 2796 4133
rect 2256 613 2346 623
rect 2886 4073 2926 4133
rect 3140 4230 3210 4240
rect 2796 613 2886 623
rect 1874 463 1948 473
rect 3210 670 6280 680
rect 3210 470 5800 670
rect 6260 470 6280 670
rect 3140 460 6280 470
rect 2140 400 2980 410
rect 1870 100 1950 110
rect 1320 20 1330 80
rect 1410 20 1870 80
rect 1330 10 1870 20
rect 1870 0 1950 10
rect 2140 -80 2980 330
rect -2200 -120 5980 -80
rect 6160 -120 6280 460
rect -2200 -160 5979 -120
rect -2403 -227 -2344 -217
rect -2403 -1005 -2344 -1004
rect -2404 -1014 -2344 -1005
rect -2200 -228 -2141 -160
rect -1997 -227 -1938 -217
rect -1997 -1005 -1938 -1004
rect -2404 -1060 -2345 -1014
rect -2200 -1015 -2141 -1005
rect -1998 -1014 -1938 -1005
rect -1794 -228 -1735 -160
rect -1591 -227 -1532 -217
rect -1591 -1005 -1532 -1004
rect -1998 -1060 -1939 -1014
rect -1794 -1015 -1735 -1005
rect -1592 -1014 -1532 -1005
rect -1388 -228 -1329 -160
rect -1185 -227 -1126 -217
rect -1185 -1005 -1126 -1004
rect -1592 -1060 -1533 -1014
rect -1388 -1015 -1329 -1005
rect -1186 -1014 -1126 -1005
rect -982 -228 -923 -160
rect -779 -227 -720 -217
rect -779 -1005 -720 -1004
rect -1186 -1060 -1127 -1014
rect -982 -1015 -923 -1005
rect -780 -1014 -720 -1005
rect -576 -228 -517 -160
rect -373 -227 -314 -217
rect -373 -1005 -314 -1004
rect -780 -1060 -721 -1014
rect -576 -1015 -517 -1005
rect -374 -1014 -314 -1005
rect -170 -228 -111 -160
rect 33 -227 92 -217
rect 33 -1005 92 -1004
rect -374 -1060 -315 -1014
rect -170 -1015 -111 -1005
rect 32 -1014 92 -1005
rect 236 -228 295 -160
rect 439 -227 498 -217
rect 439 -1005 498 -1004
rect 32 -1060 91 -1014
rect 236 -1015 295 -1005
rect 438 -1014 498 -1005
rect 642 -228 701 -160
rect 845 -227 904 -217
rect 845 -1005 904 -1004
rect 438 -1060 497 -1014
rect 642 -1015 701 -1005
rect 844 -1014 904 -1005
rect 1048 -228 1107 -160
rect 1251 -227 1310 -217
rect 1251 -1005 1310 -1004
rect 844 -1060 903 -1014
rect 1048 -1015 1107 -1005
rect 1250 -1014 1310 -1005
rect 1454 -228 1513 -160
rect 2063 -227 2122 -217
rect 1650 -250 1710 -240
rect 1650 -950 1710 -940
rect 1871 -249 1931 -239
rect 1871 -949 1931 -939
rect 2063 -1005 2122 -1004
rect 1250 -1060 1309 -1014
rect 1454 -1015 1513 -1005
rect 2062 -1014 2122 -1005
rect 2266 -228 2325 -160
rect 2469 -227 2528 -217
rect 2469 -1005 2528 -1004
rect 2062 -1060 2121 -1014
rect 2266 -1015 2325 -1005
rect 2468 -1014 2528 -1005
rect 2672 -228 2731 -160
rect 2875 -227 2934 -217
rect 2875 -1005 2934 -1004
rect 2468 -1060 2527 -1014
rect 2672 -1015 2731 -1005
rect 2874 -1014 2934 -1005
rect 3078 -228 3137 -160
rect 3281 -227 3340 -217
rect 3281 -1005 3340 -1004
rect 2874 -1060 2933 -1014
rect 3078 -1015 3137 -1005
rect 3280 -1014 3340 -1005
rect 3484 -228 3543 -160
rect 3687 -227 3746 -217
rect 3687 -1005 3746 -1004
rect 3280 -1060 3339 -1014
rect 3484 -1015 3543 -1005
rect 3686 -1014 3746 -1005
rect 3890 -228 3949 -160
rect 4093 -227 4152 -217
rect 4093 -1005 4152 -1004
rect 3686 -1060 3745 -1014
rect 3890 -1015 3949 -1005
rect 4092 -1014 4152 -1005
rect 4296 -228 4355 -160
rect 4499 -227 4558 -217
rect 4499 -1005 4558 -1004
rect 4092 -1060 4151 -1014
rect 4296 -1015 4355 -1005
rect 4498 -1014 4558 -1005
rect 4702 -228 4761 -160
rect 4905 -227 4964 -217
rect 4905 -1005 4964 -1004
rect 4498 -1060 4557 -1014
rect 4702 -1015 4761 -1005
rect 4904 -1014 4964 -1005
rect 5108 -228 5167 -160
rect 5311 -227 5370 -217
rect 5311 -1005 5370 -1004
rect 4904 -1060 4963 -1014
rect 5108 -1015 5167 -1005
rect 5310 -1014 5370 -1005
rect 5514 -228 5573 -160
rect 5717 -227 5776 -217
rect 5717 -1005 5776 -1004
rect 5310 -1060 5369 -1014
rect 5514 -1015 5573 -1005
rect 5716 -1014 5776 -1005
rect 5920 -228 5979 -160
rect 6160 -200 6280 -190
rect 5716 -1060 5775 -1014
rect 5920 -1015 5979 -1005
rect -2404 -1112 5775 -1060
rect -2404 -1152 5776 -1112
rect -2404 -1153 -1930 -1152
rect -1592 -1153 -1533 -1152
rect -1186 -1153 -1127 -1152
rect -780 -1153 -721 -1152
rect -374 -1153 -315 -1152
rect 32 -1153 91 -1152
rect 438 -1153 497 -1152
rect 844 -1153 903 -1152
rect 1250 -1153 1309 -1152
rect 1656 -1153 1715 -1152
rect 2062 -1153 2121 -1152
rect 2468 -1153 2527 -1152
rect 2874 -1153 2933 -1152
rect 3280 -1153 3339 -1152
rect 3686 -1153 3745 -1152
rect 4092 -1153 4151 -1152
rect 4498 -1153 4557 -1152
rect 4904 -1153 4963 -1152
rect 5310 -1153 5369 -1152
rect 5716 -1153 5775 -1152
rect -2400 -1210 -1930 -1153
rect -2340 -1420 -1930 -1210
rect 1640 -1210 1740 -1200
rect 1640 -1300 1740 -1290
rect -2350 -1430 -1930 -1420
rect -1940 -2540 -1930 -1430
rect -2350 -2550 -1930 -2540
rect -2340 -2800 -1930 -2550
rect -2350 -2810 -1930 -2800
rect -1940 -3920 -1930 -2810
rect -2350 -3930 -1940 -3920
<< via2 >>
rect 1874 473 1948 4227
rect 1870 10 1950 100
rect 1650 -940 1710 -250
rect 1871 -939 1931 -249
rect 1640 -1290 1740 -1210
<< metal3 >>
rect 1864 4227 1958 4232
rect 1864 473 1874 4227
rect 1948 473 1958 4227
rect 1864 468 1958 473
rect 1871 105 1947 468
rect 1860 100 1960 105
rect 1860 10 1870 100
rect 1950 10 1960 100
rect 1860 5 1960 10
rect 1871 -130 1947 5
rect 1870 -244 1950 -130
rect 1640 -250 1720 -245
rect 1640 -940 1650 -250
rect 1710 -940 1720 -250
rect 1640 -945 1720 -940
rect 1861 -249 1950 -244
rect 1861 -939 1871 -249
rect 1931 -300 1950 -249
rect 1931 -939 1947 -300
rect 1861 -944 1941 -939
rect 1640 -1205 1710 -945
rect 1630 -1210 1750 -1205
rect 1630 -1290 1640 -1210
rect 1740 -1290 1750 -1210
rect 1630 -1295 1750 -1290
use sky130_fd_pr__nfet_01v8_BKH6ZK  sky130_fd_pr__nfet_01v8_BKH6ZK_0
timestamp 1714085375
transform 1 0 1382 0 1 -616
box -256 -610 256 610
use sky130_fd_pr__nfet_01v8_BKH6ZK  sky130_fd_pr__nfet_01v8_BKH6ZK_1
timestamp 1714085375
transform 1 0 2194 0 1 -616
box -256 -610 256 610
use sky130_fd_pr__nfet_01v8_BKH6ZK  sky130_fd_pr__nfet_01v8_BKH6ZK_2
timestamp 1714085375
transform 1 0 976 0 1 -616
box -256 -610 256 610
use sky130_fd_pr__nfet_01v8_BKH6ZK  sky130_fd_pr__nfet_01v8_BKH6ZK_3
timestamp 1714085375
transform 1 0 2600 0 1 -616
box -256 -610 256 610
use sky130_fd_pr__nfet_01v8_BKH6ZK  sky130_fd_pr__nfet_01v8_BKH6ZK_4
timestamp 1714085375
transform 1 0 3006 0 1 -616
box -256 -610 256 610
use sky130_fd_pr__nfet_01v8_BKH6ZK  sky130_fd_pr__nfet_01v8_BKH6ZK_5
timestamp 1714085375
transform 1 0 3412 0 1 -616
box -256 -610 256 610
use sky130_fd_pr__nfet_01v8_BKH6ZK  sky130_fd_pr__nfet_01v8_BKH6ZK_6
timestamp 1714085375
transform 1 0 3818 0 1 -616
box -256 -610 256 610
use sky130_fd_pr__nfet_01v8_BKH6ZK  sky130_fd_pr__nfet_01v8_BKH6ZK_7
timestamp 1714085375
transform 1 0 -2272 0 1 -616
box -256 -610 256 610
use sky130_fd_pr__nfet_01v8_BKH6ZK  sky130_fd_pr__nfet_01v8_BKH6ZK_8
timestamp 1714085375
transform 1 0 5442 0 1 -616
box -256 -610 256 610
use sky130_fd_pr__nfet_01v8_BKH6ZK  sky130_fd_pr__nfet_01v8_BKH6ZK_9
timestamp 1714085375
transform 1 0 5036 0 1 -616
box -256 -610 256 610
use sky130_fd_pr__nfet_01v8_BKH6ZK  sky130_fd_pr__nfet_01v8_BKH6ZK_10
timestamp 1714085375
transform 1 0 4630 0 1 -616
box -256 -610 256 610
use sky130_fd_pr__nfet_01v8_BKH6ZK  sky130_fd_pr__nfet_01v8_BKH6ZK_11
timestamp 1714085375
transform 1 0 5848 0 1 -616
box -256 -610 256 610
use sky130_fd_pr__nfet_01v8_BKH6ZK  sky130_fd_pr__nfet_01v8_BKH6ZK_12
timestamp 1714085375
transform 1 0 4224 0 1 -616
box -256 -610 256 610
use sky130_fd_pr__nfet_01v8_BKH6ZK  sky130_fd_pr__nfet_01v8_BKH6ZK_13
timestamp 1714085375
transform 1 0 570 0 1 -616
box -256 -610 256 610
use sky130_fd_pr__nfet_01v8_BKH6ZK  sky130_fd_pr__nfet_01v8_BKH6ZK_14
timestamp 1714085375
transform 1 0 164 0 1 -616
box -256 -610 256 610
use sky130_fd_pr__nfet_01v8_BKH6ZK  sky130_fd_pr__nfet_01v8_BKH6ZK_15
timestamp 1714085375
transform 1 0 -242 0 1 -616
box -256 -610 256 610
use sky130_fd_pr__nfet_01v8_BKH6ZK  sky130_fd_pr__nfet_01v8_BKH6ZK_16
timestamp 1714085375
transform 1 0 -648 0 1 -616
box -256 -610 256 610
use sky130_fd_pr__nfet_01v8_BKH6ZK  sky130_fd_pr__nfet_01v8_BKH6ZK_17
timestamp 1714085375
transform 1 0 -1054 0 1 -616
box -256 -610 256 610
use sky130_fd_pr__nfet_01v8_BKH6ZK  sky130_fd_pr__nfet_01v8_BKH6ZK_18
timestamp 1714085375
transform 1 0 -1460 0 1 -616
box -256 -610 256 610
use sky130_fd_pr__nfet_01v8_BKH6ZK  sky130_fd_pr__nfet_01v8_BKH6ZK_19
timestamp 1714085375
transform 1 0 -1866 0 1 -616
box -256 -610 256 610
use sky130_fd_pr__pfet_01v8_lvt_GUHUBJ  XM1
timestamp 1713931681
transform 1 0 2062 0 1 2346
box -296 -2119 296 2119
use sky130_fd_pr__pfet_01v8_lvt_GUHUBJ  XM2
timestamp 1713931681
transform 1 0 2548 0 1 2346
box -296 -2119 296 2119
use sky130_fd_pr__pfet_01v8_lvt_GUHUBJ  XM3
timestamp 1713931681
transform 1 0 3034 0 1 2346
box -296 -2119 296 2119
use sky130_fd_pr__nfet_01v8_lvt_AWHWK2  XM4
timestamp 1714103463
transform 1 0 1788 0 1 -616
box -256 -610 256 610
use sky130_fd_pr__nfet_01v8_lvt_B7MEP5  XM6
timestamp 1714102074
transform 0 1 1411 -1 0 111
box -211 -221 211 221
use sky130_fd_pr__nfet_01v8_lvt_AWHWK2  XM7
timestamp 1714103463
transform 1 0 6254 0 1 -616
box -256 -610 256 610
use sky130_fd_pr__res_xhigh_po_5p73_GWLG8Y  XR1
timestamp 1713929811
transform 0 1 6646 -1 0 -3359
box -739 -9176 739 9176
use sky130_fd_pr__res_xhigh_po_5p73_GWLG8Y  XR2
timestamp 1713929811
transform 0 1 6646 -1 0 -1987
box -739 -9176 739 9176
<< labels >>
flabel metal1 2466 4493 2666 4693 0 FreeSans 256 0 0 0 VDD
port 0 nsew
flabel metal1 6380 510 6580 710 0 FreeSans 256 0 0 0 VOUT
port 1 nsew
flabel metal1 9480 -990 9680 -790 0 FreeSans 256 0 0 0 VSS
port 2 nsew
<< end >>
