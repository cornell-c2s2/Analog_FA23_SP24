magic
tech sky130A
magscale 1 2
timestamp 1711862879
<< error_s >>
rect 4056 4299 4118 4305
rect 4056 4265 4068 4299
rect 4056 4259 4118 4265
rect 2492 3766 2554 3772
rect 2492 3732 2504 3766
rect 2492 3726 2554 3732
rect 4056 3371 4118 3377
rect 4056 3337 4068 3371
rect 4056 3331 4118 3337
rect 2492 2838 2554 2844
rect 2492 2804 2504 2838
rect 2492 2798 2554 2804
rect 3970 1230 4032 1236
rect 3970 1196 3982 1230
rect 3970 1190 4032 1196
rect 5246 1079 5281 1113
rect 5247 1060 5281 1079
rect 5055 1011 5117 1017
rect 5055 977 5067 1011
rect 5055 971 5117 977
rect 2952 779 2987 813
rect 2953 760 2987 779
rect 2783 711 2841 717
rect 2783 677 2795 711
rect 2783 671 2841 677
rect 2783 401 2841 407
rect 2783 367 2795 401
rect 2783 361 2841 367
rect 2972 265 2987 760
rect 3006 726 3041 760
rect 3321 726 3356 760
rect 3006 265 3040 726
rect 3322 707 3356 726
rect 3152 658 3210 664
rect 3152 624 3164 658
rect 3152 618 3210 624
rect 3152 348 3210 354
rect 3152 314 3164 348
rect 3152 308 3210 314
rect 3006 231 3021 265
rect 3341 212 3356 707
rect 3375 673 3410 707
rect 3375 212 3409 673
rect 3521 605 3579 611
rect 3521 571 3533 605
rect 3521 565 3579 571
rect 3970 302 4032 308
rect 3521 295 3579 301
rect 3521 261 3533 295
rect 3970 268 3982 302
rect 3970 262 4032 268
rect 3521 255 3579 261
rect 3375 178 3390 212
rect 5055 83 5117 89
rect 5055 49 5067 83
rect 5055 43 5117 49
rect 5266 -53 5281 1060
rect 5300 1026 5335 1060
rect 5655 1026 5690 1043
rect 5300 -53 5334 1026
rect 5656 1025 5690 1026
rect 5656 989 5726 1025
rect 5464 958 5526 964
rect 5464 924 5476 958
rect 5673 955 5744 989
rect 6114 955 6149 989
rect 5464 918 5526 924
rect 5464 30 5526 36
rect 5464 -4 5476 30
rect 5464 -10 5526 -4
rect 5300 -87 5315 -53
rect 5673 -106 5743 955
rect 6115 936 6149 955
rect 5673 -142 5726 -106
rect 6134 -159 6149 936
rect 6168 902 6203 936
rect 6168 -159 6202 902
rect 6168 -193 6183 -159
<< viali >>
rect 1000 -1680 2690 -1630
<< metal1 >>
rect 1520 460 1530 540
rect 1590 460 1750 540
rect 1990 460 2150 540
rect 2210 460 2220 540
rect 0 0 200 200
rect 1640 40 1774 420
rect 1970 40 2104 420
rect 1520 -80 1530 0
rect 1590 -80 1750 0
rect 1990 -80 2150 0
rect 2210 -80 2220 0
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
rect 1510 -1080 1520 -300
rect 1590 -1080 1600 -300
rect 1740 -1080 2000 -310
rect 2140 -1080 2150 -300
rect 2220 -1080 2230 -300
rect 1770 -1100 1970 -1080
rect 1800 -1290 1940 -1100
rect 1780 -1310 1960 -1290
rect 960 -1340 2770 -1310
rect 960 -1380 1760 -1340
rect 1970 -1380 2770 -1340
rect 0 -1600 200 -1400
rect 1800 -1510 1940 -1400
rect 970 -1570 1770 -1530
rect 1970 -1570 2770 -1530
rect 970 -1590 2770 -1570
rect 980 -1630 2760 -1590
rect 980 -1680 1000 -1630
rect 2690 -1640 2760 -1630
rect 2690 -1680 2770 -1640
rect 980 -1700 2770 -1680
rect 0 -2000 200 -1800
rect 0 -2400 200 -2200
rect 0 -2800 200 -2600
<< via1 >>
rect 1530 460 1590 540
rect 2150 460 2210 540
rect 1530 -80 1590 0
rect 2150 -80 2210 0
rect 1520 -1080 1590 -300
rect 2150 -1080 2220 -300
<< metal2 >>
rect 1520 540 1590 550
rect 1520 460 1530 540
rect 1520 0 1590 460
rect 1520 -80 1530 0
rect 1520 -300 1590 -80
rect 1520 -1090 1590 -1080
rect 2150 540 2220 550
rect 2210 460 2220 540
rect 2150 0 2220 460
rect 2210 -80 2220 0
rect 2150 -300 2220 -80
rect 2150 -1090 2220 -1080
use sky130_fd_pr__nfet_01v8_lvt_648S5X  XM1
timestamp 1711862879
transform 1 0 3550 0 1 433
box -211 -310 211 310
use sky130_fd_pr__pfet_01v8_lvt_4QFHB3  XM2
timestamp 1711862879
transform 1 0 4001 0 1 749
box -231 -619 231 619
use sky130_fd_pr__nfet_01v8_lvt_AWHWK2  XM3
timestamp 1711824350
transform 1 0 5929 0 1 415
box -256 -610 256 610
use sky130_fd_pr__nfet_01v8_lvt_AWHWK2  XM4
timestamp 1711824350
transform 1 0 6388 0 1 362
box -256 -610 256 610
use sky130_fd_pr__nfet_01v8_lvt_ATY4A8  XM5
timestamp 1711844308
transform 1 0 1711 0 1 230
box -211 -410 211 410
use sky130_fd_pr__pfet_01v8_lvt_4QFHB3  XM6
timestamp 1711862879
transform 1 0 4087 0 1 3818
box -231 -619 231 619
use sky130_fd_pr__pfet_01v8_lvt_4QFHB3  XM7
timestamp 1711862879
transform 1 0 2523 0 1 3285
box -231 -619 231 619
use sky130_fd_pr__nfet_01v8_lvt_LGA5SN  XM8
timestamp 1711825685
transform 1 0 2031 0 1 230
box -211 -410 211 410
use sky130_fd_pr__pfet_01v8_lvt_4QFHB3  XM9
timestamp 1711862879
transform 1 0 5086 0 1 530
box -231 -619 231 619
use sky130_fd_pr__nfet_01v8_lvt_648S5X  XM10
timestamp 1711862879
transform 1 0 2812 0 1 539
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_lvt_648S5X  XM11
timestamp 1711862879
transform 1 0 3181 0 1 486
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_lvt_AWHWK2  XM12
timestamp 1711824350
transform 1 0 662 0 1 1104
box -256 -610 256 610
use sky130_fd_pr__nfet_01v8_lvt_T2JW3B  XM13
timestamp 1711824350
transform 0 1 1869 -1 0 -1454
box -256 -1119 256 1119
use sky130_fd_pr__pfet_01v8_lvt_4QFHB3  XM14
timestamp 1711862879
transform 1 0 5495 0 1 477
box -231 -619 231 619
use sky130_fd_pr__nfet_01v8_lvt_UGLW3B  XM15
timestamp 1711825065
transform 1 0 2077 0 1 -689
box -256 -610 256 610
use sky130_fd_pr__nfet_01v8_lvt_AWHWK2  XM17
timestamp 1711824350
transform 1 0 1666 0 1 -690
box -256 -610 256 610
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 VDD
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 IB
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 VSS
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 VIP
port 3 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 256 0 0 0 VIN
port 4 nsew
flabel metal1 0 -2000 200 -1800 0 FreeSans 256 0 0 0 VON
port 5 nsew
flabel metal1 0 -2400 200 -2200 0 FreeSans 256 0 0 0 VOP
port 6 nsew
flabel metal1 0 -2800 200 -2600 0 FreeSans 256 0 0 0 CLK
port 7 nsew
<< end >>
