magic
tech sky130A
magscale 1 2
timestamp 1683376989
<< nwell >>
rect 41330 690750 47990 695500
rect 538289 685502 550909 690942
rect 43710 681100 45600 684040
rect 540434 680239 548644 681480
rect 540794 680238 548412 680239
<< pwell >>
rect 37527 693357 40723 696295
rect 48597 693357 51793 696295
rect 43931 689211 45371 690631
rect 43931 687691 45371 689111
rect 42940 686170 46370 687590
rect 42680 684650 46626 686070
rect 534556 685189 537752 688137
rect 540249 684722 548977 685214
rect 551616 685189 554812 688137
rect 540249 684222 548977 684714
rect 540809 683622 548319 684214
rect 540809 683002 548319 683594
rect 540249 682402 548977 682994
rect 540249 681802 548977 682394
rect 44310 680000 44960 680920
rect 43950 679250 45316 679920
rect 543564 679448 545638 680040
rect 43695 677750 45577 679170
rect 543784 678923 545422 679415
rect 540849 678298 548359 678890
rect 41150 662800 48180 677610
rect 541314 677290 547888 678108
rect 541314 671978 547894 677290
rect 541314 664522 547884 671978
rect 541312 663278 547884 664522
<< nmos >>
rect 44127 689421 44227 690421
rect 44285 689421 44385 690421
rect 44443 689421 44543 690421
rect 44601 689421 44701 690421
rect 44759 689421 44859 690421
rect 44917 689421 45017 690421
rect 45075 689421 45175 690421
rect 44127 687901 44227 688901
rect 44285 687901 44385 688901
rect 44443 687901 44543 688901
rect 44601 687901 44701 688901
rect 44759 687901 44859 688901
rect 44917 687901 45017 688901
rect 45075 687901 45175 688901
rect 43136 686380 43336 687380
rect 43394 686380 43594 687380
rect 43652 686380 43852 687380
rect 43910 686380 44110 687380
rect 44168 686380 44368 687380
rect 44426 686380 44626 687380
rect 44684 686380 44884 687380
rect 44942 686380 45142 687380
rect 45200 686380 45400 687380
rect 45458 686380 45658 687380
rect 45716 686380 45916 687380
rect 45974 686380 46174 687380
rect 42876 684860 43076 685860
rect 43134 684860 43334 685860
rect 43392 684860 43592 685860
rect 43650 684860 43850 685860
rect 43908 684860 44108 685860
rect 44166 684860 44366 685860
rect 44424 684860 44624 685860
rect 44682 684860 44882 685860
rect 44940 684860 45140 685860
rect 45198 684860 45398 685860
rect 45456 684860 45656 685860
rect 45714 684860 45914 685860
rect 45972 684860 46172 685860
rect 46230 684860 46430 685860
rect 540459 684918 541459 685018
rect 541677 684918 542677 685018
rect 542895 684918 543895 685018
rect 544113 684918 545113 685018
rect 545331 684918 546331 685018
rect 546549 684918 547549 685018
rect 547767 684918 548767 685018
rect 540459 684418 541459 684518
rect 541677 684418 542677 684518
rect 542895 684418 543895 684518
rect 544113 684418 545113 684518
rect 545331 684418 546331 684518
rect 546549 684418 547549 684518
rect 547767 684418 548767 684518
rect 541019 683818 542019 684018
rect 542237 683818 543237 684018
rect 543455 683818 544455 684018
rect 544673 683818 545673 684018
rect 545891 683818 546891 684018
rect 547109 683818 548109 684018
rect 541019 683198 542019 683398
rect 542237 683198 543237 683398
rect 543455 683198 544455 683398
rect 544673 683198 545673 683398
rect 545891 683198 546891 683398
rect 547109 683198 548109 683398
rect 540459 682598 541459 682798
rect 541677 682598 542677 682798
rect 542895 682598 543895 682798
rect 544113 682598 545113 682798
rect 545331 682598 546331 682798
rect 546549 682598 547549 682798
rect 547767 682598 548767 682798
rect 540459 681998 541459 682198
rect 541677 681998 542677 682198
rect 542895 681998 543895 682198
rect 544113 681998 545113 682198
rect 545331 681998 546331 682198
rect 546549 681998 547549 682198
rect 547767 681998 548767 682198
rect 44506 680210 44606 680710
rect 44664 680210 44764 680710
rect 44146 679460 44346 679710
rect 44404 679460 44604 679710
rect 44662 679460 44862 679710
rect 44920 679460 45120 679710
rect 543774 679644 544024 679844
rect 544242 679644 544492 679844
rect 544710 679644 544960 679844
rect 545178 679644 545428 679844
rect 43891 677960 44091 678960
rect 44149 677960 44349 678960
rect 44407 677960 44607 678960
rect 44665 677960 44865 678960
rect 44923 677960 45123 678960
rect 45181 677960 45381 678960
rect 543994 679119 544494 679219
rect 544712 679119 545212 679219
rect 541059 678494 542059 678694
rect 542277 678494 543277 678694
rect 543495 678494 544495 678694
rect 544713 678494 545713 678694
rect 545931 678494 546931 678694
rect 547149 678494 548149 678694
<< pmos >>
rect 41526 694199 41626 695199
rect 41684 694199 41784 695199
rect 41842 694199 41942 695199
rect 42000 694199 42100 695199
rect 42158 694199 42258 695199
rect 42316 694199 42416 695199
rect 42474 694199 42574 695199
rect 42632 694199 42732 695199
rect 42790 694199 42890 695199
rect 42948 694199 43048 695199
rect 43106 694199 43206 695199
rect 43264 694199 43364 695199
rect 43422 694199 43522 695199
rect 43580 694199 43680 695199
rect 43738 694199 43838 695199
rect 43896 694199 43996 695199
rect 44054 694199 44154 695199
rect 44212 694199 44312 695199
rect 44370 694199 44470 695199
rect 44528 694199 44628 695199
rect 44686 694199 44786 695199
rect 44844 694199 44944 695199
rect 45002 694199 45102 695199
rect 45160 694199 45260 695199
rect 45318 694199 45418 695199
rect 45476 694199 45576 695199
rect 45634 694199 45734 695199
rect 45792 694199 45892 695199
rect 45950 694199 46050 695199
rect 46108 694199 46208 695199
rect 46266 694199 46366 695199
rect 46424 694199 46524 695199
rect 46582 694199 46682 695199
rect 46740 694199 46840 695199
rect 46898 694199 46998 695199
rect 47056 694199 47156 695199
rect 47214 694199 47314 695199
rect 47372 694199 47472 695199
rect 47530 694199 47630 695199
rect 47688 694199 47788 695199
rect 43026 692529 43126 693529
rect 43184 692529 43284 693529
rect 43342 692529 43442 693529
rect 43500 692529 43600 693529
rect 43658 692529 43758 693529
rect 43816 692529 43916 693529
rect 43974 692529 44074 693529
rect 44132 692529 44232 693529
rect 44290 692529 44390 693529
rect 44448 692529 44548 693529
rect 44606 692529 44706 693529
rect 44764 692529 44864 693529
rect 44922 692529 45022 693529
rect 45080 692529 45180 693529
rect 45238 692529 45338 693529
rect 45396 692529 45496 693529
rect 45554 692529 45654 693529
rect 45712 692529 45812 693529
rect 45870 692529 45970 693529
rect 46028 692529 46128 693529
rect 46186 692529 46286 693529
rect 43026 690989 43126 691989
rect 43184 690989 43284 691989
rect 43342 690989 43442 691989
rect 43500 690989 43600 691989
rect 43658 690989 43758 691989
rect 43816 690989 43916 691989
rect 43974 690989 44074 691989
rect 44132 690989 44232 691989
rect 44290 690989 44390 691989
rect 44448 690989 44548 691989
rect 44606 690989 44706 691989
rect 44764 690989 44864 691989
rect 44922 690989 45022 691989
rect 45080 690989 45180 691989
rect 45238 690989 45338 691989
rect 45396 690989 45496 691989
rect 45554 690989 45654 691989
rect 45712 690989 45812 691989
rect 45870 690989 45970 691989
rect 46028 690989 46128 691989
rect 46186 690989 46286 691989
rect 540368 690638 541368 690738
rect 541604 690638 542604 690738
rect 542840 690638 543840 690738
rect 544076 690638 545076 690738
rect 545312 690638 546312 690738
rect 546548 690638 547548 690738
rect 547784 690638 548784 690738
rect 540368 690098 541368 690198
rect 541604 690098 542604 690198
rect 542840 690098 543840 690198
rect 544076 690098 545076 690198
rect 545312 690098 546312 690198
rect 546548 690098 547548 690198
rect 547784 690098 548784 690198
rect 540368 689558 541368 689658
rect 541604 689558 542604 689658
rect 542840 689558 543840 689658
rect 544076 689558 545076 689658
rect 545312 689558 546312 689658
rect 546548 689558 547548 689658
rect 547784 689558 548784 689658
rect 540368 689018 541368 689118
rect 541604 689018 542604 689118
rect 542840 689018 543840 689118
rect 544076 689018 545076 689118
rect 545312 689018 546312 689118
rect 546548 689018 547548 689118
rect 547784 689018 548784 689118
rect 540368 688438 541368 688538
rect 541604 688438 542604 688538
rect 542840 688438 543840 688538
rect 544076 688438 545076 688538
rect 545312 688438 546312 688538
rect 546548 688438 547548 688538
rect 547784 688438 548784 688538
rect 540368 687858 541368 687958
rect 541604 687858 542604 687958
rect 542840 687858 543840 687958
rect 544076 687858 545076 687958
rect 545312 687858 546312 687958
rect 546548 687858 547548 687958
rect 547784 687858 548784 687958
rect 538528 687318 539528 687418
rect 539764 687318 540764 687418
rect 541000 687318 542000 687418
rect 542236 687318 543236 687418
rect 543472 687318 544472 687418
rect 544708 687318 545708 687418
rect 545944 687318 546944 687418
rect 547180 687318 548180 687418
rect 548416 687318 549416 687418
rect 549652 687318 550652 687418
rect 538528 686778 539528 686878
rect 539764 686778 540764 686878
rect 541000 686778 542000 686878
rect 542236 686778 543236 686878
rect 543472 686778 544472 686878
rect 544708 686778 545708 686878
rect 545944 686778 546944 686878
rect 547180 686778 548180 686878
rect 548416 686778 549416 686878
rect 549652 686778 550652 686878
rect 538528 686238 539528 686338
rect 539764 686238 540764 686338
rect 541000 686238 542000 686338
rect 542236 686238 543236 686338
rect 543472 686238 544472 686338
rect 544708 686238 545708 686338
rect 545944 686238 546944 686338
rect 547180 686238 548180 686338
rect 548416 686238 549416 686338
rect 549652 686238 550652 686338
rect 538528 685698 539528 685798
rect 539764 685698 540764 685798
rect 541000 685698 542000 685798
rect 542236 685698 543236 685798
rect 543472 685698 544472 685798
rect 544708 685698 545708 685798
rect 545944 685698 546944 685798
rect 547180 685698 548180 685798
rect 548416 685698 549416 685798
rect 549652 685698 550652 685798
rect 43906 682819 44106 683819
rect 44164 682819 44364 683819
rect 44422 682819 44622 683819
rect 44680 682819 44880 683819
rect 44938 682819 45138 683819
rect 45196 682819 45396 683819
rect 43906 681319 44106 682319
rect 44164 681319 44364 682319
rect 44422 681319 44622 682319
rect 44680 681319 44880 682319
rect 44938 681319 45138 682319
rect 45196 681319 45396 682319
rect 541013 681024 542013 681224
rect 542249 681024 543249 681224
rect 543485 681024 544485 681224
rect 544721 681024 545721 681224
rect 545957 681024 546957 681224
rect 547193 681024 548193 681224
rect 541013 680434 542013 680634
rect 542249 680434 543249 680634
rect 543485 680434 544485 680634
rect 544721 680434 545721 680634
rect 545957 680434 546957 680634
rect 547193 680434 548193 680634
<< ndiff >>
rect 44069 690409 44127 690421
rect 44069 689433 44081 690409
rect 44115 689433 44127 690409
rect 44069 689421 44127 689433
rect 44227 690409 44285 690421
rect 44227 689433 44239 690409
rect 44273 689433 44285 690409
rect 44227 689421 44285 689433
rect 44385 690409 44443 690421
rect 44385 689433 44397 690409
rect 44431 689433 44443 690409
rect 44385 689421 44443 689433
rect 44543 690409 44601 690421
rect 44543 689433 44555 690409
rect 44589 689433 44601 690409
rect 44543 689421 44601 689433
rect 44701 690409 44759 690421
rect 44701 689433 44713 690409
rect 44747 689433 44759 690409
rect 44701 689421 44759 689433
rect 44859 690409 44917 690421
rect 44859 689433 44871 690409
rect 44905 689433 44917 690409
rect 44859 689421 44917 689433
rect 45017 690409 45075 690421
rect 45017 689433 45029 690409
rect 45063 689433 45075 690409
rect 45017 689421 45075 689433
rect 45175 690409 45233 690421
rect 45175 689433 45187 690409
rect 45221 689433 45233 690409
rect 45175 689421 45233 689433
rect 44069 688889 44127 688901
rect 44069 687913 44081 688889
rect 44115 687913 44127 688889
rect 44069 687901 44127 687913
rect 44227 688889 44285 688901
rect 44227 687913 44239 688889
rect 44273 687913 44285 688889
rect 44227 687901 44285 687913
rect 44385 688889 44443 688901
rect 44385 687913 44397 688889
rect 44431 687913 44443 688889
rect 44385 687901 44443 687913
rect 44543 688889 44601 688901
rect 44543 687913 44555 688889
rect 44589 687913 44601 688889
rect 44543 687901 44601 687913
rect 44701 688889 44759 688901
rect 44701 687913 44713 688889
rect 44747 687913 44759 688889
rect 44701 687901 44759 687913
rect 44859 688889 44917 688901
rect 44859 687913 44871 688889
rect 44905 687913 44917 688889
rect 44859 687901 44917 687913
rect 45017 688889 45075 688901
rect 45017 687913 45029 688889
rect 45063 687913 45075 688889
rect 45017 687901 45075 687913
rect 45175 688889 45233 688901
rect 45175 687913 45187 688889
rect 45221 687913 45233 688889
rect 45175 687901 45233 687913
rect 43078 687368 43136 687380
rect 43078 686392 43090 687368
rect 43124 686392 43136 687368
rect 43078 686380 43136 686392
rect 43336 687368 43394 687380
rect 43336 686392 43348 687368
rect 43382 686392 43394 687368
rect 43336 686380 43394 686392
rect 43594 687368 43652 687380
rect 43594 686392 43606 687368
rect 43640 686392 43652 687368
rect 43594 686380 43652 686392
rect 43852 687368 43910 687380
rect 43852 686392 43864 687368
rect 43898 686392 43910 687368
rect 43852 686380 43910 686392
rect 44110 687368 44168 687380
rect 44110 686392 44122 687368
rect 44156 686392 44168 687368
rect 44110 686380 44168 686392
rect 44368 687368 44426 687380
rect 44368 686392 44380 687368
rect 44414 686392 44426 687368
rect 44368 686380 44426 686392
rect 44626 687368 44684 687380
rect 44626 686392 44638 687368
rect 44672 686392 44684 687368
rect 44626 686380 44684 686392
rect 44884 687368 44942 687380
rect 44884 686392 44896 687368
rect 44930 686392 44942 687368
rect 44884 686380 44942 686392
rect 45142 687368 45200 687380
rect 45142 686392 45154 687368
rect 45188 686392 45200 687368
rect 45142 686380 45200 686392
rect 45400 687368 45458 687380
rect 45400 686392 45412 687368
rect 45446 686392 45458 687368
rect 45400 686380 45458 686392
rect 45658 687368 45716 687380
rect 45658 686392 45670 687368
rect 45704 686392 45716 687368
rect 45658 686380 45716 686392
rect 45916 687368 45974 687380
rect 45916 686392 45928 687368
rect 45962 686392 45974 687368
rect 45916 686380 45974 686392
rect 46174 687368 46232 687380
rect 46174 686392 46186 687368
rect 46220 686392 46232 687368
rect 46174 686380 46232 686392
rect 42818 685848 42876 685860
rect 42818 684872 42830 685848
rect 42864 684872 42876 685848
rect 42818 684860 42876 684872
rect 43076 685848 43134 685860
rect 43076 684872 43088 685848
rect 43122 684872 43134 685848
rect 43076 684860 43134 684872
rect 43334 685848 43392 685860
rect 43334 684872 43346 685848
rect 43380 684872 43392 685848
rect 43334 684860 43392 684872
rect 43592 685848 43650 685860
rect 43592 684872 43604 685848
rect 43638 684872 43650 685848
rect 43592 684860 43650 684872
rect 43850 685848 43908 685860
rect 43850 684872 43862 685848
rect 43896 684872 43908 685848
rect 43850 684860 43908 684872
rect 44108 685848 44166 685860
rect 44108 684872 44120 685848
rect 44154 684872 44166 685848
rect 44108 684860 44166 684872
rect 44366 685848 44424 685860
rect 44366 684872 44378 685848
rect 44412 684872 44424 685848
rect 44366 684860 44424 684872
rect 44624 685848 44682 685860
rect 44624 684872 44636 685848
rect 44670 684872 44682 685848
rect 44624 684860 44682 684872
rect 44882 685848 44940 685860
rect 44882 684872 44894 685848
rect 44928 684872 44940 685848
rect 44882 684860 44940 684872
rect 45140 685848 45198 685860
rect 45140 684872 45152 685848
rect 45186 684872 45198 685848
rect 45140 684860 45198 684872
rect 45398 685848 45456 685860
rect 45398 684872 45410 685848
rect 45444 684872 45456 685848
rect 45398 684860 45456 684872
rect 45656 685848 45714 685860
rect 45656 684872 45668 685848
rect 45702 684872 45714 685848
rect 45656 684860 45714 684872
rect 45914 685848 45972 685860
rect 45914 684872 45926 685848
rect 45960 684872 45972 685848
rect 45914 684860 45972 684872
rect 46172 685848 46230 685860
rect 46172 684872 46184 685848
rect 46218 684872 46230 685848
rect 46172 684860 46230 684872
rect 46430 685848 46488 685860
rect 46430 684872 46442 685848
rect 46476 684872 46488 685848
rect 46430 684860 46488 684872
rect 540459 685064 541459 685076
rect 540459 685030 540471 685064
rect 541447 685030 541459 685064
rect 540459 685018 541459 685030
rect 541677 685064 542677 685076
rect 541677 685030 541689 685064
rect 542665 685030 542677 685064
rect 541677 685018 542677 685030
rect 542895 685064 543895 685076
rect 542895 685030 542907 685064
rect 543883 685030 543895 685064
rect 542895 685018 543895 685030
rect 544113 685064 545113 685076
rect 544113 685030 544125 685064
rect 545101 685030 545113 685064
rect 544113 685018 545113 685030
rect 545331 685064 546331 685076
rect 545331 685030 545343 685064
rect 546319 685030 546331 685064
rect 545331 685018 546331 685030
rect 546549 685064 547549 685076
rect 546549 685030 546561 685064
rect 547537 685030 547549 685064
rect 546549 685018 547549 685030
rect 547767 685064 548767 685076
rect 547767 685030 547779 685064
rect 548755 685030 548767 685064
rect 547767 685018 548767 685030
rect 540459 684906 541459 684918
rect 540459 684872 540471 684906
rect 541447 684872 541459 684906
rect 540459 684860 541459 684872
rect 541677 684906 542677 684918
rect 541677 684872 541689 684906
rect 542665 684872 542677 684906
rect 541677 684860 542677 684872
rect 542895 684906 543895 684918
rect 542895 684872 542907 684906
rect 543883 684872 543895 684906
rect 542895 684860 543895 684872
rect 544113 684906 545113 684918
rect 544113 684872 544125 684906
rect 545101 684872 545113 684906
rect 544113 684860 545113 684872
rect 545331 684906 546331 684918
rect 545331 684872 545343 684906
rect 546319 684872 546331 684906
rect 545331 684860 546331 684872
rect 546549 684906 547549 684918
rect 546549 684872 546561 684906
rect 547537 684872 547549 684906
rect 546549 684860 547549 684872
rect 547767 684906 548767 684918
rect 547767 684872 547779 684906
rect 548755 684872 548767 684906
rect 547767 684860 548767 684872
rect 540459 684564 541459 684576
rect 540459 684530 540471 684564
rect 541447 684530 541459 684564
rect 540459 684518 541459 684530
rect 541677 684564 542677 684576
rect 541677 684530 541689 684564
rect 542665 684530 542677 684564
rect 541677 684518 542677 684530
rect 542895 684564 543895 684576
rect 542895 684530 542907 684564
rect 543883 684530 543895 684564
rect 542895 684518 543895 684530
rect 544113 684564 545113 684576
rect 544113 684530 544125 684564
rect 545101 684530 545113 684564
rect 544113 684518 545113 684530
rect 545331 684564 546331 684576
rect 545331 684530 545343 684564
rect 546319 684530 546331 684564
rect 545331 684518 546331 684530
rect 546549 684564 547549 684576
rect 546549 684530 546561 684564
rect 547537 684530 547549 684564
rect 546549 684518 547549 684530
rect 547767 684564 548767 684576
rect 547767 684530 547779 684564
rect 548755 684530 548767 684564
rect 547767 684518 548767 684530
rect 540459 684406 541459 684418
rect 540459 684372 540471 684406
rect 541447 684372 541459 684406
rect 540459 684360 541459 684372
rect 541677 684406 542677 684418
rect 541677 684372 541689 684406
rect 542665 684372 542677 684406
rect 541677 684360 542677 684372
rect 542895 684406 543895 684418
rect 542895 684372 542907 684406
rect 543883 684372 543895 684406
rect 542895 684360 543895 684372
rect 544113 684406 545113 684418
rect 544113 684372 544125 684406
rect 545101 684372 545113 684406
rect 544113 684360 545113 684372
rect 545331 684406 546331 684418
rect 545331 684372 545343 684406
rect 546319 684372 546331 684406
rect 545331 684360 546331 684372
rect 546549 684406 547549 684418
rect 546549 684372 546561 684406
rect 547537 684372 547549 684406
rect 546549 684360 547549 684372
rect 547767 684406 548767 684418
rect 547767 684372 547779 684406
rect 548755 684372 548767 684406
rect 547767 684360 548767 684372
rect 541019 684064 542019 684076
rect 541019 684030 541031 684064
rect 542007 684030 542019 684064
rect 541019 684018 542019 684030
rect 542237 684064 543237 684076
rect 542237 684030 542249 684064
rect 543225 684030 543237 684064
rect 542237 684018 543237 684030
rect 543455 684064 544455 684076
rect 543455 684030 543467 684064
rect 544443 684030 544455 684064
rect 543455 684018 544455 684030
rect 544673 684064 545673 684076
rect 544673 684030 544685 684064
rect 545661 684030 545673 684064
rect 544673 684018 545673 684030
rect 545891 684064 546891 684076
rect 545891 684030 545903 684064
rect 546879 684030 546891 684064
rect 545891 684018 546891 684030
rect 547109 684064 548109 684076
rect 547109 684030 547121 684064
rect 548097 684030 548109 684064
rect 547109 684018 548109 684030
rect 541019 683806 542019 683818
rect 541019 683772 541031 683806
rect 542007 683772 542019 683806
rect 541019 683760 542019 683772
rect 542237 683806 543237 683818
rect 542237 683772 542249 683806
rect 543225 683772 543237 683806
rect 542237 683760 543237 683772
rect 543455 683806 544455 683818
rect 543455 683772 543467 683806
rect 544443 683772 544455 683806
rect 543455 683760 544455 683772
rect 544673 683806 545673 683818
rect 544673 683772 544685 683806
rect 545661 683772 545673 683806
rect 544673 683760 545673 683772
rect 545891 683806 546891 683818
rect 545891 683772 545903 683806
rect 546879 683772 546891 683806
rect 545891 683760 546891 683772
rect 547109 683806 548109 683818
rect 547109 683772 547121 683806
rect 548097 683772 548109 683806
rect 547109 683760 548109 683772
rect 541019 683444 542019 683456
rect 541019 683410 541031 683444
rect 542007 683410 542019 683444
rect 541019 683398 542019 683410
rect 542237 683444 543237 683456
rect 542237 683410 542249 683444
rect 543225 683410 543237 683444
rect 542237 683398 543237 683410
rect 543455 683444 544455 683456
rect 543455 683410 543467 683444
rect 544443 683410 544455 683444
rect 543455 683398 544455 683410
rect 544673 683444 545673 683456
rect 544673 683410 544685 683444
rect 545661 683410 545673 683444
rect 544673 683398 545673 683410
rect 545891 683444 546891 683456
rect 545891 683410 545903 683444
rect 546879 683410 546891 683444
rect 545891 683398 546891 683410
rect 547109 683444 548109 683456
rect 547109 683410 547121 683444
rect 548097 683410 548109 683444
rect 547109 683398 548109 683410
rect 541019 683186 542019 683198
rect 541019 683152 541031 683186
rect 542007 683152 542019 683186
rect 541019 683140 542019 683152
rect 542237 683186 543237 683198
rect 542237 683152 542249 683186
rect 543225 683152 543237 683186
rect 542237 683140 543237 683152
rect 543455 683186 544455 683198
rect 543455 683152 543467 683186
rect 544443 683152 544455 683186
rect 543455 683140 544455 683152
rect 544673 683186 545673 683198
rect 544673 683152 544685 683186
rect 545661 683152 545673 683186
rect 544673 683140 545673 683152
rect 545891 683186 546891 683198
rect 545891 683152 545903 683186
rect 546879 683152 546891 683186
rect 545891 683140 546891 683152
rect 547109 683186 548109 683198
rect 547109 683152 547121 683186
rect 548097 683152 548109 683186
rect 547109 683140 548109 683152
rect 540459 682844 541459 682856
rect 540459 682810 540471 682844
rect 541447 682810 541459 682844
rect 540459 682798 541459 682810
rect 541677 682844 542677 682856
rect 541677 682810 541689 682844
rect 542665 682810 542677 682844
rect 541677 682798 542677 682810
rect 542895 682844 543895 682856
rect 542895 682810 542907 682844
rect 543883 682810 543895 682844
rect 542895 682798 543895 682810
rect 544113 682844 545113 682856
rect 544113 682810 544125 682844
rect 545101 682810 545113 682844
rect 544113 682798 545113 682810
rect 545331 682844 546331 682856
rect 545331 682810 545343 682844
rect 546319 682810 546331 682844
rect 545331 682798 546331 682810
rect 546549 682844 547549 682856
rect 546549 682810 546561 682844
rect 547537 682810 547549 682844
rect 546549 682798 547549 682810
rect 547767 682844 548767 682856
rect 547767 682810 547779 682844
rect 548755 682810 548767 682844
rect 547767 682798 548767 682810
rect 540459 682586 541459 682598
rect 540459 682552 540471 682586
rect 541447 682552 541459 682586
rect 540459 682540 541459 682552
rect 541677 682586 542677 682598
rect 541677 682552 541689 682586
rect 542665 682552 542677 682586
rect 541677 682540 542677 682552
rect 542895 682586 543895 682598
rect 542895 682552 542907 682586
rect 543883 682552 543895 682586
rect 542895 682540 543895 682552
rect 544113 682586 545113 682598
rect 544113 682552 544125 682586
rect 545101 682552 545113 682586
rect 544113 682540 545113 682552
rect 545331 682586 546331 682598
rect 545331 682552 545343 682586
rect 546319 682552 546331 682586
rect 545331 682540 546331 682552
rect 546549 682586 547549 682598
rect 546549 682552 546561 682586
rect 547537 682552 547549 682586
rect 546549 682540 547549 682552
rect 547767 682586 548767 682598
rect 547767 682552 547779 682586
rect 548755 682552 548767 682586
rect 547767 682540 548767 682552
rect 540459 682244 541459 682256
rect 540459 682210 540471 682244
rect 541447 682210 541459 682244
rect 540459 682198 541459 682210
rect 541677 682244 542677 682256
rect 541677 682210 541689 682244
rect 542665 682210 542677 682244
rect 541677 682198 542677 682210
rect 542895 682244 543895 682256
rect 542895 682210 542907 682244
rect 543883 682210 543895 682244
rect 542895 682198 543895 682210
rect 544113 682244 545113 682256
rect 544113 682210 544125 682244
rect 545101 682210 545113 682244
rect 544113 682198 545113 682210
rect 545331 682244 546331 682256
rect 545331 682210 545343 682244
rect 546319 682210 546331 682244
rect 545331 682198 546331 682210
rect 546549 682244 547549 682256
rect 546549 682210 546561 682244
rect 547537 682210 547549 682244
rect 546549 682198 547549 682210
rect 547767 682244 548767 682256
rect 547767 682210 547779 682244
rect 548755 682210 548767 682244
rect 547767 682198 548767 682210
rect 540459 681986 541459 681998
rect 540459 681952 540471 681986
rect 541447 681952 541459 681986
rect 540459 681940 541459 681952
rect 541677 681986 542677 681998
rect 541677 681952 541689 681986
rect 542665 681952 542677 681986
rect 541677 681940 542677 681952
rect 542895 681986 543895 681998
rect 542895 681952 542907 681986
rect 543883 681952 543895 681986
rect 542895 681940 543895 681952
rect 544113 681986 545113 681998
rect 544113 681952 544125 681986
rect 545101 681952 545113 681986
rect 544113 681940 545113 681952
rect 545331 681986 546331 681998
rect 545331 681952 545343 681986
rect 546319 681952 546331 681986
rect 545331 681940 546331 681952
rect 546549 681986 547549 681998
rect 546549 681952 546561 681986
rect 547537 681952 547549 681986
rect 546549 681940 547549 681952
rect 547767 681986 548767 681998
rect 547767 681952 547779 681986
rect 548755 681952 548767 681986
rect 547767 681940 548767 681952
rect 44448 680698 44506 680710
rect 44448 680222 44460 680698
rect 44494 680222 44506 680698
rect 44448 680210 44506 680222
rect 44606 680698 44664 680710
rect 44606 680222 44618 680698
rect 44652 680222 44664 680698
rect 44606 680210 44664 680222
rect 44764 680698 44822 680710
rect 44764 680222 44776 680698
rect 44810 680222 44822 680698
rect 44764 680210 44822 680222
rect 44088 679698 44146 679710
rect 44088 679472 44100 679698
rect 44134 679472 44146 679698
rect 44088 679460 44146 679472
rect 44346 679698 44404 679710
rect 44346 679472 44358 679698
rect 44392 679472 44404 679698
rect 44346 679460 44404 679472
rect 44604 679698 44662 679710
rect 44604 679472 44616 679698
rect 44650 679472 44662 679698
rect 44604 679460 44662 679472
rect 44862 679698 44920 679710
rect 44862 679472 44874 679698
rect 44908 679472 44920 679698
rect 44862 679460 44920 679472
rect 45120 679698 45178 679710
rect 45120 679472 45132 679698
rect 45166 679472 45178 679698
rect 45120 679460 45178 679472
rect 543774 679890 544024 679902
rect 543774 679856 543786 679890
rect 544012 679856 544024 679890
rect 543774 679844 544024 679856
rect 544242 679890 544492 679902
rect 544242 679856 544254 679890
rect 544480 679856 544492 679890
rect 544242 679844 544492 679856
rect 544710 679890 544960 679902
rect 544710 679856 544722 679890
rect 544948 679856 544960 679890
rect 544710 679844 544960 679856
rect 545178 679890 545428 679902
rect 545178 679856 545190 679890
rect 545416 679856 545428 679890
rect 545178 679844 545428 679856
rect 543774 679632 544024 679644
rect 543774 679598 543786 679632
rect 544012 679598 544024 679632
rect 543774 679586 544024 679598
rect 544242 679632 544492 679644
rect 544242 679598 544254 679632
rect 544480 679598 544492 679632
rect 544242 679586 544492 679598
rect 544710 679632 544960 679644
rect 544710 679598 544722 679632
rect 544948 679598 544960 679632
rect 544710 679586 544960 679598
rect 545178 679632 545428 679644
rect 545178 679598 545190 679632
rect 545416 679598 545428 679632
rect 545178 679586 545428 679598
rect 43833 678948 43891 678960
rect 43833 677972 43845 678948
rect 43879 677972 43891 678948
rect 43833 677960 43891 677972
rect 44091 678948 44149 678960
rect 44091 677972 44103 678948
rect 44137 677972 44149 678948
rect 44091 677960 44149 677972
rect 44349 678948 44407 678960
rect 44349 677972 44361 678948
rect 44395 677972 44407 678948
rect 44349 677960 44407 677972
rect 44607 678948 44665 678960
rect 44607 677972 44619 678948
rect 44653 677972 44665 678948
rect 44607 677960 44665 677972
rect 44865 678948 44923 678960
rect 44865 677972 44877 678948
rect 44911 677972 44923 678948
rect 44865 677960 44923 677972
rect 45123 678948 45181 678960
rect 45123 677972 45135 678948
rect 45169 677972 45181 678948
rect 45123 677960 45181 677972
rect 45381 678948 45439 678960
rect 45381 677972 45393 678948
rect 45427 677972 45439 678948
rect 45381 677960 45439 677972
rect 543994 679265 544494 679277
rect 543994 679231 544006 679265
rect 544482 679231 544494 679265
rect 543994 679219 544494 679231
rect 544712 679265 545212 679277
rect 544712 679231 544724 679265
rect 545200 679231 545212 679265
rect 544712 679219 545212 679231
rect 543994 679107 544494 679119
rect 543994 679073 544006 679107
rect 544482 679073 544494 679107
rect 543994 679061 544494 679073
rect 544712 679107 545212 679119
rect 544712 679073 544724 679107
rect 545200 679073 545212 679107
rect 544712 679061 545212 679073
rect 541059 678740 542059 678752
rect 541059 678706 541071 678740
rect 542047 678706 542059 678740
rect 541059 678694 542059 678706
rect 542277 678740 543277 678752
rect 542277 678706 542289 678740
rect 543265 678706 543277 678740
rect 542277 678694 543277 678706
rect 543495 678740 544495 678752
rect 543495 678706 543507 678740
rect 544483 678706 544495 678740
rect 543495 678694 544495 678706
rect 544713 678740 545713 678752
rect 544713 678706 544725 678740
rect 545701 678706 545713 678740
rect 544713 678694 545713 678706
rect 545931 678740 546931 678752
rect 545931 678706 545943 678740
rect 546919 678706 546931 678740
rect 545931 678694 546931 678706
rect 547149 678740 548149 678752
rect 547149 678706 547161 678740
rect 548137 678706 548149 678740
rect 547149 678694 548149 678706
rect 541059 678482 542059 678494
rect 541059 678448 541071 678482
rect 542047 678448 542059 678482
rect 541059 678436 542059 678448
rect 542277 678482 543277 678494
rect 542277 678448 542289 678482
rect 543265 678448 543277 678482
rect 542277 678436 543277 678448
rect 543495 678482 544495 678494
rect 543495 678448 543507 678482
rect 544483 678448 544495 678482
rect 543495 678436 544495 678448
rect 544713 678482 545713 678494
rect 544713 678448 544725 678482
rect 545701 678448 545713 678482
rect 544713 678436 545713 678448
rect 545931 678482 546931 678494
rect 545931 678448 545943 678482
rect 546919 678448 546931 678482
rect 545931 678436 546931 678448
rect 547149 678482 548149 678494
rect 547149 678448 547161 678482
rect 548137 678448 548149 678482
rect 547149 678436 548149 678448
<< pdiff >>
rect 41468 695187 41526 695199
rect 41468 694211 41480 695187
rect 41514 694211 41526 695187
rect 41468 694199 41526 694211
rect 41626 695187 41684 695199
rect 41626 694211 41638 695187
rect 41672 694211 41684 695187
rect 41626 694199 41684 694211
rect 41784 695187 41842 695199
rect 41784 694211 41796 695187
rect 41830 694211 41842 695187
rect 41784 694199 41842 694211
rect 41942 695187 42000 695199
rect 41942 694211 41954 695187
rect 41988 694211 42000 695187
rect 41942 694199 42000 694211
rect 42100 695187 42158 695199
rect 42100 694211 42112 695187
rect 42146 694211 42158 695187
rect 42100 694199 42158 694211
rect 42258 695187 42316 695199
rect 42258 694211 42270 695187
rect 42304 694211 42316 695187
rect 42258 694199 42316 694211
rect 42416 695187 42474 695199
rect 42416 694211 42428 695187
rect 42462 694211 42474 695187
rect 42416 694199 42474 694211
rect 42574 695187 42632 695199
rect 42574 694211 42586 695187
rect 42620 694211 42632 695187
rect 42574 694199 42632 694211
rect 42732 695187 42790 695199
rect 42732 694211 42744 695187
rect 42778 694211 42790 695187
rect 42732 694199 42790 694211
rect 42890 695187 42948 695199
rect 42890 694211 42902 695187
rect 42936 694211 42948 695187
rect 42890 694199 42948 694211
rect 43048 695187 43106 695199
rect 43048 694211 43060 695187
rect 43094 694211 43106 695187
rect 43048 694199 43106 694211
rect 43206 695187 43264 695199
rect 43206 694211 43218 695187
rect 43252 694211 43264 695187
rect 43206 694199 43264 694211
rect 43364 695187 43422 695199
rect 43364 694211 43376 695187
rect 43410 694211 43422 695187
rect 43364 694199 43422 694211
rect 43522 695187 43580 695199
rect 43522 694211 43534 695187
rect 43568 694211 43580 695187
rect 43522 694199 43580 694211
rect 43680 695187 43738 695199
rect 43680 694211 43692 695187
rect 43726 694211 43738 695187
rect 43680 694199 43738 694211
rect 43838 695187 43896 695199
rect 43838 694211 43850 695187
rect 43884 694211 43896 695187
rect 43838 694199 43896 694211
rect 43996 695187 44054 695199
rect 43996 694211 44008 695187
rect 44042 694211 44054 695187
rect 43996 694199 44054 694211
rect 44154 695187 44212 695199
rect 44154 694211 44166 695187
rect 44200 694211 44212 695187
rect 44154 694199 44212 694211
rect 44312 695187 44370 695199
rect 44312 694211 44324 695187
rect 44358 694211 44370 695187
rect 44312 694199 44370 694211
rect 44470 695187 44528 695199
rect 44470 694211 44482 695187
rect 44516 694211 44528 695187
rect 44470 694199 44528 694211
rect 44628 695187 44686 695199
rect 44628 694211 44640 695187
rect 44674 694211 44686 695187
rect 44628 694199 44686 694211
rect 44786 695187 44844 695199
rect 44786 694211 44798 695187
rect 44832 694211 44844 695187
rect 44786 694199 44844 694211
rect 44944 695187 45002 695199
rect 44944 694211 44956 695187
rect 44990 694211 45002 695187
rect 44944 694199 45002 694211
rect 45102 695187 45160 695199
rect 45102 694211 45114 695187
rect 45148 694211 45160 695187
rect 45102 694199 45160 694211
rect 45260 695187 45318 695199
rect 45260 694211 45272 695187
rect 45306 694211 45318 695187
rect 45260 694199 45318 694211
rect 45418 695187 45476 695199
rect 45418 694211 45430 695187
rect 45464 694211 45476 695187
rect 45418 694199 45476 694211
rect 45576 695187 45634 695199
rect 45576 694211 45588 695187
rect 45622 694211 45634 695187
rect 45576 694199 45634 694211
rect 45734 695187 45792 695199
rect 45734 694211 45746 695187
rect 45780 694211 45792 695187
rect 45734 694199 45792 694211
rect 45892 695187 45950 695199
rect 45892 694211 45904 695187
rect 45938 694211 45950 695187
rect 45892 694199 45950 694211
rect 46050 695187 46108 695199
rect 46050 694211 46062 695187
rect 46096 694211 46108 695187
rect 46050 694199 46108 694211
rect 46208 695187 46266 695199
rect 46208 694211 46220 695187
rect 46254 694211 46266 695187
rect 46208 694199 46266 694211
rect 46366 695187 46424 695199
rect 46366 694211 46378 695187
rect 46412 694211 46424 695187
rect 46366 694199 46424 694211
rect 46524 695187 46582 695199
rect 46524 694211 46536 695187
rect 46570 694211 46582 695187
rect 46524 694199 46582 694211
rect 46682 695187 46740 695199
rect 46682 694211 46694 695187
rect 46728 694211 46740 695187
rect 46682 694199 46740 694211
rect 46840 695187 46898 695199
rect 46840 694211 46852 695187
rect 46886 694211 46898 695187
rect 46840 694199 46898 694211
rect 46998 695187 47056 695199
rect 46998 694211 47010 695187
rect 47044 694211 47056 695187
rect 46998 694199 47056 694211
rect 47156 695187 47214 695199
rect 47156 694211 47168 695187
rect 47202 694211 47214 695187
rect 47156 694199 47214 694211
rect 47314 695187 47372 695199
rect 47314 694211 47326 695187
rect 47360 694211 47372 695187
rect 47314 694199 47372 694211
rect 47472 695187 47530 695199
rect 47472 694211 47484 695187
rect 47518 694211 47530 695187
rect 47472 694199 47530 694211
rect 47630 695187 47688 695199
rect 47630 694211 47642 695187
rect 47676 694211 47688 695187
rect 47630 694199 47688 694211
rect 47788 695187 47846 695199
rect 47788 694211 47800 695187
rect 47834 694211 47846 695187
rect 47788 694199 47846 694211
rect 42968 693517 43026 693529
rect 42968 692541 42980 693517
rect 43014 692541 43026 693517
rect 42968 692529 43026 692541
rect 43126 693517 43184 693529
rect 43126 692541 43138 693517
rect 43172 692541 43184 693517
rect 43126 692529 43184 692541
rect 43284 693517 43342 693529
rect 43284 692541 43296 693517
rect 43330 692541 43342 693517
rect 43284 692529 43342 692541
rect 43442 693517 43500 693529
rect 43442 692541 43454 693517
rect 43488 692541 43500 693517
rect 43442 692529 43500 692541
rect 43600 693517 43658 693529
rect 43600 692541 43612 693517
rect 43646 692541 43658 693517
rect 43600 692529 43658 692541
rect 43758 693517 43816 693529
rect 43758 692541 43770 693517
rect 43804 692541 43816 693517
rect 43758 692529 43816 692541
rect 43916 693517 43974 693529
rect 43916 692541 43928 693517
rect 43962 692541 43974 693517
rect 43916 692529 43974 692541
rect 44074 693517 44132 693529
rect 44074 692541 44086 693517
rect 44120 692541 44132 693517
rect 44074 692529 44132 692541
rect 44232 693517 44290 693529
rect 44232 692541 44244 693517
rect 44278 692541 44290 693517
rect 44232 692529 44290 692541
rect 44390 693517 44448 693529
rect 44390 692541 44402 693517
rect 44436 692541 44448 693517
rect 44390 692529 44448 692541
rect 44548 693517 44606 693529
rect 44548 692541 44560 693517
rect 44594 692541 44606 693517
rect 44548 692529 44606 692541
rect 44706 693517 44764 693529
rect 44706 692541 44718 693517
rect 44752 692541 44764 693517
rect 44706 692529 44764 692541
rect 44864 693517 44922 693529
rect 44864 692541 44876 693517
rect 44910 692541 44922 693517
rect 44864 692529 44922 692541
rect 45022 693517 45080 693529
rect 45022 692541 45034 693517
rect 45068 692541 45080 693517
rect 45022 692529 45080 692541
rect 45180 693517 45238 693529
rect 45180 692541 45192 693517
rect 45226 692541 45238 693517
rect 45180 692529 45238 692541
rect 45338 693517 45396 693529
rect 45338 692541 45350 693517
rect 45384 692541 45396 693517
rect 45338 692529 45396 692541
rect 45496 693517 45554 693529
rect 45496 692541 45508 693517
rect 45542 692541 45554 693517
rect 45496 692529 45554 692541
rect 45654 693517 45712 693529
rect 45654 692541 45666 693517
rect 45700 692541 45712 693517
rect 45654 692529 45712 692541
rect 45812 693517 45870 693529
rect 45812 692541 45824 693517
rect 45858 692541 45870 693517
rect 45812 692529 45870 692541
rect 45970 693517 46028 693529
rect 45970 692541 45982 693517
rect 46016 692541 46028 693517
rect 45970 692529 46028 692541
rect 46128 693517 46186 693529
rect 46128 692541 46140 693517
rect 46174 692541 46186 693517
rect 46128 692529 46186 692541
rect 46286 693517 46344 693529
rect 46286 692541 46298 693517
rect 46332 692541 46344 693517
rect 46286 692529 46344 692541
rect 42968 691977 43026 691989
rect 42968 691001 42980 691977
rect 43014 691001 43026 691977
rect 42968 690989 43026 691001
rect 43126 691977 43184 691989
rect 43126 691001 43138 691977
rect 43172 691001 43184 691977
rect 43126 690989 43184 691001
rect 43284 691977 43342 691989
rect 43284 691001 43296 691977
rect 43330 691001 43342 691977
rect 43284 690989 43342 691001
rect 43442 691977 43500 691989
rect 43442 691001 43454 691977
rect 43488 691001 43500 691977
rect 43442 690989 43500 691001
rect 43600 691977 43658 691989
rect 43600 691001 43612 691977
rect 43646 691001 43658 691977
rect 43600 690989 43658 691001
rect 43758 691977 43816 691989
rect 43758 691001 43770 691977
rect 43804 691001 43816 691977
rect 43758 690989 43816 691001
rect 43916 691977 43974 691989
rect 43916 691001 43928 691977
rect 43962 691001 43974 691977
rect 43916 690989 43974 691001
rect 44074 691977 44132 691989
rect 44074 691001 44086 691977
rect 44120 691001 44132 691977
rect 44074 690989 44132 691001
rect 44232 691977 44290 691989
rect 44232 691001 44244 691977
rect 44278 691001 44290 691977
rect 44232 690989 44290 691001
rect 44390 691977 44448 691989
rect 44390 691001 44402 691977
rect 44436 691001 44448 691977
rect 44390 690989 44448 691001
rect 44548 691977 44606 691989
rect 44548 691001 44560 691977
rect 44594 691001 44606 691977
rect 44548 690989 44606 691001
rect 44706 691977 44764 691989
rect 44706 691001 44718 691977
rect 44752 691001 44764 691977
rect 44706 690989 44764 691001
rect 44864 691977 44922 691989
rect 44864 691001 44876 691977
rect 44910 691001 44922 691977
rect 44864 690989 44922 691001
rect 45022 691977 45080 691989
rect 45022 691001 45034 691977
rect 45068 691001 45080 691977
rect 45022 690989 45080 691001
rect 45180 691977 45238 691989
rect 45180 691001 45192 691977
rect 45226 691001 45238 691977
rect 45180 690989 45238 691001
rect 45338 691977 45396 691989
rect 45338 691001 45350 691977
rect 45384 691001 45396 691977
rect 45338 690989 45396 691001
rect 45496 691977 45554 691989
rect 45496 691001 45508 691977
rect 45542 691001 45554 691977
rect 45496 690989 45554 691001
rect 45654 691977 45712 691989
rect 45654 691001 45666 691977
rect 45700 691001 45712 691977
rect 45654 690989 45712 691001
rect 45812 691977 45870 691989
rect 45812 691001 45824 691977
rect 45858 691001 45870 691977
rect 45812 690989 45870 691001
rect 45970 691977 46028 691989
rect 45970 691001 45982 691977
rect 46016 691001 46028 691977
rect 45970 690989 46028 691001
rect 46128 691977 46186 691989
rect 46128 691001 46140 691977
rect 46174 691001 46186 691977
rect 46128 690989 46186 691001
rect 46286 691977 46344 691989
rect 46286 691001 46298 691977
rect 46332 691001 46344 691977
rect 46286 690989 46344 691001
rect 540368 690784 541368 690796
rect 540368 690750 540380 690784
rect 541356 690750 541368 690784
rect 540368 690738 541368 690750
rect 541604 690784 542604 690796
rect 541604 690750 541616 690784
rect 542592 690750 542604 690784
rect 541604 690738 542604 690750
rect 542840 690784 543840 690796
rect 542840 690750 542852 690784
rect 543828 690750 543840 690784
rect 542840 690738 543840 690750
rect 544076 690784 545076 690796
rect 544076 690750 544088 690784
rect 545064 690750 545076 690784
rect 544076 690738 545076 690750
rect 545312 690784 546312 690796
rect 545312 690750 545324 690784
rect 546300 690750 546312 690784
rect 545312 690738 546312 690750
rect 546548 690784 547548 690796
rect 546548 690750 546560 690784
rect 547536 690750 547548 690784
rect 546548 690738 547548 690750
rect 547784 690784 548784 690796
rect 547784 690750 547796 690784
rect 548772 690750 548784 690784
rect 547784 690738 548784 690750
rect 540368 690626 541368 690638
rect 540368 690592 540380 690626
rect 541356 690592 541368 690626
rect 540368 690580 541368 690592
rect 541604 690626 542604 690638
rect 541604 690592 541616 690626
rect 542592 690592 542604 690626
rect 541604 690580 542604 690592
rect 542840 690626 543840 690638
rect 542840 690592 542852 690626
rect 543828 690592 543840 690626
rect 542840 690580 543840 690592
rect 544076 690626 545076 690638
rect 544076 690592 544088 690626
rect 545064 690592 545076 690626
rect 544076 690580 545076 690592
rect 545312 690626 546312 690638
rect 545312 690592 545324 690626
rect 546300 690592 546312 690626
rect 545312 690580 546312 690592
rect 546548 690626 547548 690638
rect 546548 690592 546560 690626
rect 547536 690592 547548 690626
rect 546548 690580 547548 690592
rect 547784 690626 548784 690638
rect 547784 690592 547796 690626
rect 548772 690592 548784 690626
rect 547784 690580 548784 690592
rect 540368 690244 541368 690256
rect 540368 690210 540380 690244
rect 541356 690210 541368 690244
rect 540368 690198 541368 690210
rect 541604 690244 542604 690256
rect 541604 690210 541616 690244
rect 542592 690210 542604 690244
rect 541604 690198 542604 690210
rect 542840 690244 543840 690256
rect 542840 690210 542852 690244
rect 543828 690210 543840 690244
rect 542840 690198 543840 690210
rect 544076 690244 545076 690256
rect 544076 690210 544088 690244
rect 545064 690210 545076 690244
rect 544076 690198 545076 690210
rect 545312 690244 546312 690256
rect 545312 690210 545324 690244
rect 546300 690210 546312 690244
rect 545312 690198 546312 690210
rect 546548 690244 547548 690256
rect 546548 690210 546560 690244
rect 547536 690210 547548 690244
rect 546548 690198 547548 690210
rect 547784 690244 548784 690256
rect 547784 690210 547796 690244
rect 548772 690210 548784 690244
rect 547784 690198 548784 690210
rect 540368 690086 541368 690098
rect 540368 690052 540380 690086
rect 541356 690052 541368 690086
rect 540368 690040 541368 690052
rect 541604 690086 542604 690098
rect 541604 690052 541616 690086
rect 542592 690052 542604 690086
rect 541604 690040 542604 690052
rect 542840 690086 543840 690098
rect 542840 690052 542852 690086
rect 543828 690052 543840 690086
rect 542840 690040 543840 690052
rect 544076 690086 545076 690098
rect 544076 690052 544088 690086
rect 545064 690052 545076 690086
rect 544076 690040 545076 690052
rect 545312 690086 546312 690098
rect 545312 690052 545324 690086
rect 546300 690052 546312 690086
rect 545312 690040 546312 690052
rect 546548 690086 547548 690098
rect 546548 690052 546560 690086
rect 547536 690052 547548 690086
rect 546548 690040 547548 690052
rect 547784 690086 548784 690098
rect 547784 690052 547796 690086
rect 548772 690052 548784 690086
rect 547784 690040 548784 690052
rect 540368 689704 541368 689716
rect 540368 689670 540380 689704
rect 541356 689670 541368 689704
rect 540368 689658 541368 689670
rect 541604 689704 542604 689716
rect 541604 689670 541616 689704
rect 542592 689670 542604 689704
rect 541604 689658 542604 689670
rect 542840 689704 543840 689716
rect 542840 689670 542852 689704
rect 543828 689670 543840 689704
rect 542840 689658 543840 689670
rect 544076 689704 545076 689716
rect 544076 689670 544088 689704
rect 545064 689670 545076 689704
rect 544076 689658 545076 689670
rect 545312 689704 546312 689716
rect 545312 689670 545324 689704
rect 546300 689670 546312 689704
rect 545312 689658 546312 689670
rect 546548 689704 547548 689716
rect 546548 689670 546560 689704
rect 547536 689670 547548 689704
rect 546548 689658 547548 689670
rect 547784 689704 548784 689716
rect 547784 689670 547796 689704
rect 548772 689670 548784 689704
rect 547784 689658 548784 689670
rect 540368 689546 541368 689558
rect 540368 689512 540380 689546
rect 541356 689512 541368 689546
rect 540368 689500 541368 689512
rect 541604 689546 542604 689558
rect 541604 689512 541616 689546
rect 542592 689512 542604 689546
rect 541604 689500 542604 689512
rect 542840 689546 543840 689558
rect 542840 689512 542852 689546
rect 543828 689512 543840 689546
rect 542840 689500 543840 689512
rect 544076 689546 545076 689558
rect 544076 689512 544088 689546
rect 545064 689512 545076 689546
rect 544076 689500 545076 689512
rect 545312 689546 546312 689558
rect 545312 689512 545324 689546
rect 546300 689512 546312 689546
rect 545312 689500 546312 689512
rect 546548 689546 547548 689558
rect 546548 689512 546560 689546
rect 547536 689512 547548 689546
rect 546548 689500 547548 689512
rect 547784 689546 548784 689558
rect 547784 689512 547796 689546
rect 548772 689512 548784 689546
rect 547784 689500 548784 689512
rect 540368 689164 541368 689176
rect 540368 689130 540380 689164
rect 541356 689130 541368 689164
rect 540368 689118 541368 689130
rect 541604 689164 542604 689176
rect 541604 689130 541616 689164
rect 542592 689130 542604 689164
rect 541604 689118 542604 689130
rect 542840 689164 543840 689176
rect 542840 689130 542852 689164
rect 543828 689130 543840 689164
rect 542840 689118 543840 689130
rect 544076 689164 545076 689176
rect 544076 689130 544088 689164
rect 545064 689130 545076 689164
rect 544076 689118 545076 689130
rect 545312 689164 546312 689176
rect 545312 689130 545324 689164
rect 546300 689130 546312 689164
rect 545312 689118 546312 689130
rect 546548 689164 547548 689176
rect 546548 689130 546560 689164
rect 547536 689130 547548 689164
rect 546548 689118 547548 689130
rect 547784 689164 548784 689176
rect 547784 689130 547796 689164
rect 548772 689130 548784 689164
rect 547784 689118 548784 689130
rect 540368 689006 541368 689018
rect 540368 688972 540380 689006
rect 541356 688972 541368 689006
rect 540368 688960 541368 688972
rect 541604 689006 542604 689018
rect 541604 688972 541616 689006
rect 542592 688972 542604 689006
rect 541604 688960 542604 688972
rect 542840 689006 543840 689018
rect 542840 688972 542852 689006
rect 543828 688972 543840 689006
rect 542840 688960 543840 688972
rect 544076 689006 545076 689018
rect 544076 688972 544088 689006
rect 545064 688972 545076 689006
rect 544076 688960 545076 688972
rect 545312 689006 546312 689018
rect 545312 688972 545324 689006
rect 546300 688972 546312 689006
rect 545312 688960 546312 688972
rect 546548 689006 547548 689018
rect 546548 688972 546560 689006
rect 547536 688972 547548 689006
rect 546548 688960 547548 688972
rect 547784 689006 548784 689018
rect 547784 688972 547796 689006
rect 548772 688972 548784 689006
rect 547784 688960 548784 688972
rect 540368 688584 541368 688596
rect 540368 688550 540380 688584
rect 541356 688550 541368 688584
rect 540368 688538 541368 688550
rect 541604 688584 542604 688596
rect 541604 688550 541616 688584
rect 542592 688550 542604 688584
rect 541604 688538 542604 688550
rect 542840 688584 543840 688596
rect 542840 688550 542852 688584
rect 543828 688550 543840 688584
rect 542840 688538 543840 688550
rect 544076 688584 545076 688596
rect 544076 688550 544088 688584
rect 545064 688550 545076 688584
rect 544076 688538 545076 688550
rect 545312 688584 546312 688596
rect 545312 688550 545324 688584
rect 546300 688550 546312 688584
rect 545312 688538 546312 688550
rect 546548 688584 547548 688596
rect 546548 688550 546560 688584
rect 547536 688550 547548 688584
rect 546548 688538 547548 688550
rect 547784 688584 548784 688596
rect 547784 688550 547796 688584
rect 548772 688550 548784 688584
rect 547784 688538 548784 688550
rect 540368 688426 541368 688438
rect 540368 688392 540380 688426
rect 541356 688392 541368 688426
rect 540368 688380 541368 688392
rect 541604 688426 542604 688438
rect 541604 688392 541616 688426
rect 542592 688392 542604 688426
rect 541604 688380 542604 688392
rect 542840 688426 543840 688438
rect 542840 688392 542852 688426
rect 543828 688392 543840 688426
rect 542840 688380 543840 688392
rect 544076 688426 545076 688438
rect 544076 688392 544088 688426
rect 545064 688392 545076 688426
rect 544076 688380 545076 688392
rect 545312 688426 546312 688438
rect 545312 688392 545324 688426
rect 546300 688392 546312 688426
rect 545312 688380 546312 688392
rect 546548 688426 547548 688438
rect 546548 688392 546560 688426
rect 547536 688392 547548 688426
rect 546548 688380 547548 688392
rect 547784 688426 548784 688438
rect 547784 688392 547796 688426
rect 548772 688392 548784 688426
rect 547784 688380 548784 688392
rect 540368 688004 541368 688016
rect 540368 687970 540380 688004
rect 541356 687970 541368 688004
rect 540368 687958 541368 687970
rect 541604 688004 542604 688016
rect 541604 687970 541616 688004
rect 542592 687970 542604 688004
rect 541604 687958 542604 687970
rect 542840 688004 543840 688016
rect 542840 687970 542852 688004
rect 543828 687970 543840 688004
rect 542840 687958 543840 687970
rect 544076 688004 545076 688016
rect 544076 687970 544088 688004
rect 545064 687970 545076 688004
rect 544076 687958 545076 687970
rect 545312 688004 546312 688016
rect 545312 687970 545324 688004
rect 546300 687970 546312 688004
rect 545312 687958 546312 687970
rect 546548 688004 547548 688016
rect 546548 687970 546560 688004
rect 547536 687970 547548 688004
rect 546548 687958 547548 687970
rect 547784 688004 548784 688016
rect 547784 687970 547796 688004
rect 548772 687970 548784 688004
rect 547784 687958 548784 687970
rect 540368 687846 541368 687858
rect 540368 687812 540380 687846
rect 541356 687812 541368 687846
rect 540368 687800 541368 687812
rect 541604 687846 542604 687858
rect 541604 687812 541616 687846
rect 542592 687812 542604 687846
rect 541604 687800 542604 687812
rect 542840 687846 543840 687858
rect 542840 687812 542852 687846
rect 543828 687812 543840 687846
rect 542840 687800 543840 687812
rect 544076 687846 545076 687858
rect 544076 687812 544088 687846
rect 545064 687812 545076 687846
rect 544076 687800 545076 687812
rect 545312 687846 546312 687858
rect 545312 687812 545324 687846
rect 546300 687812 546312 687846
rect 545312 687800 546312 687812
rect 546548 687846 547548 687858
rect 546548 687812 546560 687846
rect 547536 687812 547548 687846
rect 546548 687800 547548 687812
rect 547784 687846 548784 687858
rect 547784 687812 547796 687846
rect 548772 687812 548784 687846
rect 547784 687800 548784 687812
rect 538528 687464 539528 687476
rect 538528 687430 538540 687464
rect 539516 687430 539528 687464
rect 538528 687418 539528 687430
rect 539764 687464 540764 687476
rect 539764 687430 539776 687464
rect 540752 687430 540764 687464
rect 539764 687418 540764 687430
rect 541000 687464 542000 687476
rect 541000 687430 541012 687464
rect 541988 687430 542000 687464
rect 541000 687418 542000 687430
rect 542236 687464 543236 687476
rect 542236 687430 542248 687464
rect 543224 687430 543236 687464
rect 542236 687418 543236 687430
rect 543472 687464 544472 687476
rect 543472 687430 543484 687464
rect 544460 687430 544472 687464
rect 543472 687418 544472 687430
rect 544708 687464 545708 687476
rect 544708 687430 544720 687464
rect 545696 687430 545708 687464
rect 544708 687418 545708 687430
rect 545944 687464 546944 687476
rect 545944 687430 545956 687464
rect 546932 687430 546944 687464
rect 545944 687418 546944 687430
rect 547180 687464 548180 687476
rect 547180 687430 547192 687464
rect 548168 687430 548180 687464
rect 547180 687418 548180 687430
rect 548416 687464 549416 687476
rect 548416 687430 548428 687464
rect 549404 687430 549416 687464
rect 548416 687418 549416 687430
rect 549652 687464 550652 687476
rect 549652 687430 549664 687464
rect 550640 687430 550652 687464
rect 549652 687418 550652 687430
rect 538528 687306 539528 687318
rect 538528 687272 538540 687306
rect 539516 687272 539528 687306
rect 538528 687260 539528 687272
rect 539764 687306 540764 687318
rect 539764 687272 539776 687306
rect 540752 687272 540764 687306
rect 539764 687260 540764 687272
rect 541000 687306 542000 687318
rect 541000 687272 541012 687306
rect 541988 687272 542000 687306
rect 541000 687260 542000 687272
rect 542236 687306 543236 687318
rect 542236 687272 542248 687306
rect 543224 687272 543236 687306
rect 542236 687260 543236 687272
rect 543472 687306 544472 687318
rect 543472 687272 543484 687306
rect 544460 687272 544472 687306
rect 543472 687260 544472 687272
rect 544708 687306 545708 687318
rect 544708 687272 544720 687306
rect 545696 687272 545708 687306
rect 544708 687260 545708 687272
rect 545944 687306 546944 687318
rect 545944 687272 545956 687306
rect 546932 687272 546944 687306
rect 545944 687260 546944 687272
rect 547180 687306 548180 687318
rect 547180 687272 547192 687306
rect 548168 687272 548180 687306
rect 547180 687260 548180 687272
rect 548416 687306 549416 687318
rect 548416 687272 548428 687306
rect 549404 687272 549416 687306
rect 548416 687260 549416 687272
rect 549652 687306 550652 687318
rect 549652 687272 549664 687306
rect 550640 687272 550652 687306
rect 549652 687260 550652 687272
rect 538528 686924 539528 686936
rect 538528 686890 538540 686924
rect 539516 686890 539528 686924
rect 538528 686878 539528 686890
rect 539764 686924 540764 686936
rect 539764 686890 539776 686924
rect 540752 686890 540764 686924
rect 539764 686878 540764 686890
rect 541000 686924 542000 686936
rect 541000 686890 541012 686924
rect 541988 686890 542000 686924
rect 541000 686878 542000 686890
rect 542236 686924 543236 686936
rect 542236 686890 542248 686924
rect 543224 686890 543236 686924
rect 542236 686878 543236 686890
rect 543472 686924 544472 686936
rect 543472 686890 543484 686924
rect 544460 686890 544472 686924
rect 543472 686878 544472 686890
rect 544708 686924 545708 686936
rect 544708 686890 544720 686924
rect 545696 686890 545708 686924
rect 544708 686878 545708 686890
rect 545944 686924 546944 686936
rect 545944 686890 545956 686924
rect 546932 686890 546944 686924
rect 545944 686878 546944 686890
rect 547180 686924 548180 686936
rect 547180 686890 547192 686924
rect 548168 686890 548180 686924
rect 547180 686878 548180 686890
rect 548416 686924 549416 686936
rect 548416 686890 548428 686924
rect 549404 686890 549416 686924
rect 548416 686878 549416 686890
rect 549652 686924 550652 686936
rect 549652 686890 549664 686924
rect 550640 686890 550652 686924
rect 549652 686878 550652 686890
rect 538528 686766 539528 686778
rect 538528 686732 538540 686766
rect 539516 686732 539528 686766
rect 538528 686720 539528 686732
rect 539764 686766 540764 686778
rect 539764 686732 539776 686766
rect 540752 686732 540764 686766
rect 539764 686720 540764 686732
rect 541000 686766 542000 686778
rect 541000 686732 541012 686766
rect 541988 686732 542000 686766
rect 541000 686720 542000 686732
rect 542236 686766 543236 686778
rect 542236 686732 542248 686766
rect 543224 686732 543236 686766
rect 542236 686720 543236 686732
rect 543472 686766 544472 686778
rect 543472 686732 543484 686766
rect 544460 686732 544472 686766
rect 543472 686720 544472 686732
rect 544708 686766 545708 686778
rect 544708 686732 544720 686766
rect 545696 686732 545708 686766
rect 544708 686720 545708 686732
rect 545944 686766 546944 686778
rect 545944 686732 545956 686766
rect 546932 686732 546944 686766
rect 545944 686720 546944 686732
rect 547180 686766 548180 686778
rect 547180 686732 547192 686766
rect 548168 686732 548180 686766
rect 547180 686720 548180 686732
rect 548416 686766 549416 686778
rect 548416 686732 548428 686766
rect 549404 686732 549416 686766
rect 548416 686720 549416 686732
rect 549652 686766 550652 686778
rect 549652 686732 549664 686766
rect 550640 686732 550652 686766
rect 549652 686720 550652 686732
rect 538528 686384 539528 686396
rect 538528 686350 538540 686384
rect 539516 686350 539528 686384
rect 538528 686338 539528 686350
rect 539764 686384 540764 686396
rect 539764 686350 539776 686384
rect 540752 686350 540764 686384
rect 539764 686338 540764 686350
rect 541000 686384 542000 686396
rect 541000 686350 541012 686384
rect 541988 686350 542000 686384
rect 541000 686338 542000 686350
rect 542236 686384 543236 686396
rect 542236 686350 542248 686384
rect 543224 686350 543236 686384
rect 542236 686338 543236 686350
rect 543472 686384 544472 686396
rect 543472 686350 543484 686384
rect 544460 686350 544472 686384
rect 543472 686338 544472 686350
rect 544708 686384 545708 686396
rect 544708 686350 544720 686384
rect 545696 686350 545708 686384
rect 544708 686338 545708 686350
rect 545944 686384 546944 686396
rect 545944 686350 545956 686384
rect 546932 686350 546944 686384
rect 545944 686338 546944 686350
rect 547180 686384 548180 686396
rect 547180 686350 547192 686384
rect 548168 686350 548180 686384
rect 547180 686338 548180 686350
rect 548416 686384 549416 686396
rect 548416 686350 548428 686384
rect 549404 686350 549416 686384
rect 548416 686338 549416 686350
rect 549652 686384 550652 686396
rect 549652 686350 549664 686384
rect 550640 686350 550652 686384
rect 549652 686338 550652 686350
rect 538528 686226 539528 686238
rect 538528 686192 538540 686226
rect 539516 686192 539528 686226
rect 538528 686180 539528 686192
rect 539764 686226 540764 686238
rect 539764 686192 539776 686226
rect 540752 686192 540764 686226
rect 539764 686180 540764 686192
rect 541000 686226 542000 686238
rect 541000 686192 541012 686226
rect 541988 686192 542000 686226
rect 541000 686180 542000 686192
rect 542236 686226 543236 686238
rect 542236 686192 542248 686226
rect 543224 686192 543236 686226
rect 542236 686180 543236 686192
rect 543472 686226 544472 686238
rect 543472 686192 543484 686226
rect 544460 686192 544472 686226
rect 543472 686180 544472 686192
rect 544708 686226 545708 686238
rect 544708 686192 544720 686226
rect 545696 686192 545708 686226
rect 544708 686180 545708 686192
rect 545944 686226 546944 686238
rect 545944 686192 545956 686226
rect 546932 686192 546944 686226
rect 545944 686180 546944 686192
rect 547180 686226 548180 686238
rect 547180 686192 547192 686226
rect 548168 686192 548180 686226
rect 547180 686180 548180 686192
rect 548416 686226 549416 686238
rect 548416 686192 548428 686226
rect 549404 686192 549416 686226
rect 548416 686180 549416 686192
rect 549652 686226 550652 686238
rect 549652 686192 549664 686226
rect 550640 686192 550652 686226
rect 549652 686180 550652 686192
rect 538528 685844 539528 685856
rect 538528 685810 538540 685844
rect 539516 685810 539528 685844
rect 538528 685798 539528 685810
rect 539764 685844 540764 685856
rect 539764 685810 539776 685844
rect 540752 685810 540764 685844
rect 539764 685798 540764 685810
rect 541000 685844 542000 685856
rect 541000 685810 541012 685844
rect 541988 685810 542000 685844
rect 541000 685798 542000 685810
rect 542236 685844 543236 685856
rect 542236 685810 542248 685844
rect 543224 685810 543236 685844
rect 542236 685798 543236 685810
rect 543472 685844 544472 685856
rect 543472 685810 543484 685844
rect 544460 685810 544472 685844
rect 543472 685798 544472 685810
rect 544708 685844 545708 685856
rect 544708 685810 544720 685844
rect 545696 685810 545708 685844
rect 544708 685798 545708 685810
rect 545944 685844 546944 685856
rect 545944 685810 545956 685844
rect 546932 685810 546944 685844
rect 545944 685798 546944 685810
rect 547180 685844 548180 685856
rect 547180 685810 547192 685844
rect 548168 685810 548180 685844
rect 547180 685798 548180 685810
rect 548416 685844 549416 685856
rect 548416 685810 548428 685844
rect 549404 685810 549416 685844
rect 548416 685798 549416 685810
rect 549652 685844 550652 685856
rect 549652 685810 549664 685844
rect 550640 685810 550652 685844
rect 549652 685798 550652 685810
rect 538528 685686 539528 685698
rect 538528 685652 538540 685686
rect 539516 685652 539528 685686
rect 538528 685640 539528 685652
rect 539764 685686 540764 685698
rect 539764 685652 539776 685686
rect 540752 685652 540764 685686
rect 539764 685640 540764 685652
rect 541000 685686 542000 685698
rect 541000 685652 541012 685686
rect 541988 685652 542000 685686
rect 541000 685640 542000 685652
rect 542236 685686 543236 685698
rect 542236 685652 542248 685686
rect 543224 685652 543236 685686
rect 542236 685640 543236 685652
rect 543472 685686 544472 685698
rect 543472 685652 543484 685686
rect 544460 685652 544472 685686
rect 543472 685640 544472 685652
rect 544708 685686 545708 685698
rect 544708 685652 544720 685686
rect 545696 685652 545708 685686
rect 544708 685640 545708 685652
rect 545944 685686 546944 685698
rect 545944 685652 545956 685686
rect 546932 685652 546944 685686
rect 545944 685640 546944 685652
rect 547180 685686 548180 685698
rect 547180 685652 547192 685686
rect 548168 685652 548180 685686
rect 547180 685640 548180 685652
rect 548416 685686 549416 685698
rect 548416 685652 548428 685686
rect 549404 685652 549416 685686
rect 548416 685640 549416 685652
rect 549652 685686 550652 685698
rect 549652 685652 549664 685686
rect 550640 685652 550652 685686
rect 549652 685640 550652 685652
rect 43848 683807 43906 683819
rect 43848 682831 43860 683807
rect 43894 682831 43906 683807
rect 43848 682819 43906 682831
rect 44106 683807 44164 683819
rect 44106 682831 44118 683807
rect 44152 682831 44164 683807
rect 44106 682819 44164 682831
rect 44364 683807 44422 683819
rect 44364 682831 44376 683807
rect 44410 682831 44422 683807
rect 44364 682819 44422 682831
rect 44622 683807 44680 683819
rect 44622 682831 44634 683807
rect 44668 682831 44680 683807
rect 44622 682819 44680 682831
rect 44880 683807 44938 683819
rect 44880 682831 44892 683807
rect 44926 682831 44938 683807
rect 44880 682819 44938 682831
rect 45138 683807 45196 683819
rect 45138 682831 45150 683807
rect 45184 682831 45196 683807
rect 45138 682819 45196 682831
rect 45396 683807 45454 683819
rect 45396 682831 45408 683807
rect 45442 682831 45454 683807
rect 45396 682819 45454 682831
rect 43848 682307 43906 682319
rect 43848 681331 43860 682307
rect 43894 681331 43906 682307
rect 43848 681319 43906 681331
rect 44106 682307 44164 682319
rect 44106 681331 44118 682307
rect 44152 681331 44164 682307
rect 44106 681319 44164 681331
rect 44364 682307 44422 682319
rect 44364 681331 44376 682307
rect 44410 681331 44422 682307
rect 44364 681319 44422 681331
rect 44622 682307 44680 682319
rect 44622 681331 44634 682307
rect 44668 681331 44680 682307
rect 44622 681319 44680 681331
rect 44880 682307 44938 682319
rect 44880 681331 44892 682307
rect 44926 681331 44938 682307
rect 44880 681319 44938 681331
rect 45138 682307 45196 682319
rect 45138 681331 45150 682307
rect 45184 681331 45196 682307
rect 45138 681319 45196 681331
rect 45396 682307 45454 682319
rect 45396 681331 45408 682307
rect 45442 681331 45454 682307
rect 45396 681319 45454 681331
rect 541013 681270 542013 681282
rect 541013 681236 541025 681270
rect 542001 681236 542013 681270
rect 541013 681224 542013 681236
rect 542249 681270 543249 681282
rect 542249 681236 542261 681270
rect 543237 681236 543249 681270
rect 542249 681224 543249 681236
rect 543485 681270 544485 681282
rect 543485 681236 543497 681270
rect 544473 681236 544485 681270
rect 543485 681224 544485 681236
rect 544721 681270 545721 681282
rect 544721 681236 544733 681270
rect 545709 681236 545721 681270
rect 544721 681224 545721 681236
rect 545957 681270 546957 681282
rect 545957 681236 545969 681270
rect 546945 681236 546957 681270
rect 545957 681224 546957 681236
rect 547193 681270 548193 681282
rect 547193 681236 547205 681270
rect 548181 681236 548193 681270
rect 547193 681224 548193 681236
rect 541013 681012 542013 681024
rect 541013 680978 541025 681012
rect 542001 680978 542013 681012
rect 541013 680966 542013 680978
rect 542249 681012 543249 681024
rect 542249 680978 542261 681012
rect 543237 680978 543249 681012
rect 542249 680966 543249 680978
rect 543485 681012 544485 681024
rect 543485 680978 543497 681012
rect 544473 680978 544485 681012
rect 543485 680966 544485 680978
rect 544721 681012 545721 681024
rect 544721 680978 544733 681012
rect 545709 680978 545721 681012
rect 544721 680966 545721 680978
rect 545957 681012 546957 681024
rect 545957 680978 545969 681012
rect 546945 680978 546957 681012
rect 545957 680966 546957 680978
rect 547193 681012 548193 681024
rect 547193 680978 547205 681012
rect 548181 680978 548193 681012
rect 547193 680966 548193 680978
rect 541013 680680 542013 680692
rect 541013 680646 541025 680680
rect 542001 680646 542013 680680
rect 541013 680634 542013 680646
rect 542249 680680 543249 680692
rect 542249 680646 542261 680680
rect 543237 680646 543249 680680
rect 542249 680634 543249 680646
rect 543485 680680 544485 680692
rect 543485 680646 543497 680680
rect 544473 680646 544485 680680
rect 543485 680634 544485 680646
rect 544721 680680 545721 680692
rect 544721 680646 544733 680680
rect 545709 680646 545721 680680
rect 544721 680634 545721 680646
rect 545957 680680 546957 680692
rect 545957 680646 545969 680680
rect 546945 680646 546957 680680
rect 545957 680634 546957 680646
rect 547193 680680 548193 680692
rect 547193 680646 547205 680680
rect 548181 680646 548193 680680
rect 547193 680634 548193 680646
rect 541013 680422 542013 680434
rect 541013 680388 541025 680422
rect 542001 680388 542013 680422
rect 541013 680376 542013 680388
rect 542249 680422 543249 680434
rect 542249 680388 542261 680422
rect 543237 680388 543249 680422
rect 542249 680376 543249 680388
rect 543485 680422 544485 680434
rect 543485 680388 543497 680422
rect 544473 680388 544485 680422
rect 543485 680376 544485 680388
rect 544721 680422 545721 680434
rect 544721 680388 544733 680422
rect 545709 680388 545721 680422
rect 544721 680376 545721 680388
rect 545957 680422 546957 680434
rect 545957 680388 545969 680422
rect 546945 680388 546957 680422
rect 545957 680376 546957 680388
rect 547193 680422 548193 680434
rect 547193 680388 547205 680422
rect 548181 680388 548193 680422
rect 547193 680376 548193 680388
<< ndiffc >>
rect 44081 689433 44115 690409
rect 44239 689433 44273 690409
rect 44397 689433 44431 690409
rect 44555 689433 44589 690409
rect 44713 689433 44747 690409
rect 44871 689433 44905 690409
rect 45029 689433 45063 690409
rect 45187 689433 45221 690409
rect 44081 687913 44115 688889
rect 44239 687913 44273 688889
rect 44397 687913 44431 688889
rect 44555 687913 44589 688889
rect 44713 687913 44747 688889
rect 44871 687913 44905 688889
rect 45029 687913 45063 688889
rect 45187 687913 45221 688889
rect 43090 686392 43124 687368
rect 43348 686392 43382 687368
rect 43606 686392 43640 687368
rect 43864 686392 43898 687368
rect 44122 686392 44156 687368
rect 44380 686392 44414 687368
rect 44638 686392 44672 687368
rect 44896 686392 44930 687368
rect 45154 686392 45188 687368
rect 45412 686392 45446 687368
rect 45670 686392 45704 687368
rect 45928 686392 45962 687368
rect 46186 686392 46220 687368
rect 42830 684872 42864 685848
rect 43088 684872 43122 685848
rect 43346 684872 43380 685848
rect 43604 684872 43638 685848
rect 43862 684872 43896 685848
rect 44120 684872 44154 685848
rect 44378 684872 44412 685848
rect 44636 684872 44670 685848
rect 44894 684872 44928 685848
rect 45152 684872 45186 685848
rect 45410 684872 45444 685848
rect 45668 684872 45702 685848
rect 45926 684872 45960 685848
rect 46184 684872 46218 685848
rect 46442 684872 46476 685848
rect 540471 685030 541447 685064
rect 541689 685030 542665 685064
rect 542907 685030 543883 685064
rect 544125 685030 545101 685064
rect 545343 685030 546319 685064
rect 546561 685030 547537 685064
rect 547779 685030 548755 685064
rect 540471 684872 541447 684906
rect 541689 684872 542665 684906
rect 542907 684872 543883 684906
rect 544125 684872 545101 684906
rect 545343 684872 546319 684906
rect 546561 684872 547537 684906
rect 547779 684872 548755 684906
rect 540471 684530 541447 684564
rect 541689 684530 542665 684564
rect 542907 684530 543883 684564
rect 544125 684530 545101 684564
rect 545343 684530 546319 684564
rect 546561 684530 547537 684564
rect 547779 684530 548755 684564
rect 540471 684372 541447 684406
rect 541689 684372 542665 684406
rect 542907 684372 543883 684406
rect 544125 684372 545101 684406
rect 545343 684372 546319 684406
rect 546561 684372 547537 684406
rect 547779 684372 548755 684406
rect 541031 684030 542007 684064
rect 542249 684030 543225 684064
rect 543467 684030 544443 684064
rect 544685 684030 545661 684064
rect 545903 684030 546879 684064
rect 547121 684030 548097 684064
rect 541031 683772 542007 683806
rect 542249 683772 543225 683806
rect 543467 683772 544443 683806
rect 544685 683772 545661 683806
rect 545903 683772 546879 683806
rect 547121 683772 548097 683806
rect 541031 683410 542007 683444
rect 542249 683410 543225 683444
rect 543467 683410 544443 683444
rect 544685 683410 545661 683444
rect 545903 683410 546879 683444
rect 547121 683410 548097 683444
rect 541031 683152 542007 683186
rect 542249 683152 543225 683186
rect 543467 683152 544443 683186
rect 544685 683152 545661 683186
rect 545903 683152 546879 683186
rect 547121 683152 548097 683186
rect 540471 682810 541447 682844
rect 541689 682810 542665 682844
rect 542907 682810 543883 682844
rect 544125 682810 545101 682844
rect 545343 682810 546319 682844
rect 546561 682810 547537 682844
rect 547779 682810 548755 682844
rect 540471 682552 541447 682586
rect 541689 682552 542665 682586
rect 542907 682552 543883 682586
rect 544125 682552 545101 682586
rect 545343 682552 546319 682586
rect 546561 682552 547537 682586
rect 547779 682552 548755 682586
rect 540471 682210 541447 682244
rect 541689 682210 542665 682244
rect 542907 682210 543883 682244
rect 544125 682210 545101 682244
rect 545343 682210 546319 682244
rect 546561 682210 547537 682244
rect 547779 682210 548755 682244
rect 540471 681952 541447 681986
rect 541689 681952 542665 681986
rect 542907 681952 543883 681986
rect 544125 681952 545101 681986
rect 545343 681952 546319 681986
rect 546561 681952 547537 681986
rect 547779 681952 548755 681986
rect 44460 680222 44494 680698
rect 44618 680222 44652 680698
rect 44776 680222 44810 680698
rect 44100 679472 44134 679698
rect 44358 679472 44392 679698
rect 44616 679472 44650 679698
rect 44874 679472 44908 679698
rect 45132 679472 45166 679698
rect 543786 679856 544012 679890
rect 544254 679856 544480 679890
rect 544722 679856 544948 679890
rect 545190 679856 545416 679890
rect 543786 679598 544012 679632
rect 544254 679598 544480 679632
rect 544722 679598 544948 679632
rect 545190 679598 545416 679632
rect 43845 677972 43879 678948
rect 44103 677972 44137 678948
rect 44361 677972 44395 678948
rect 44619 677972 44653 678948
rect 44877 677972 44911 678948
rect 45135 677972 45169 678948
rect 45393 677972 45427 678948
rect 544006 679231 544482 679265
rect 544724 679231 545200 679265
rect 544006 679073 544482 679107
rect 544724 679073 545200 679107
rect 541071 678706 542047 678740
rect 542289 678706 543265 678740
rect 543507 678706 544483 678740
rect 544725 678706 545701 678740
rect 545943 678706 546919 678740
rect 547161 678706 548137 678740
rect 541071 678448 542047 678482
rect 542289 678448 543265 678482
rect 543507 678448 544483 678482
rect 544725 678448 545701 678482
rect 545943 678448 546919 678482
rect 547161 678448 548137 678482
<< pdiffc >>
rect 41480 694211 41514 695187
rect 41638 694211 41672 695187
rect 41796 694211 41830 695187
rect 41954 694211 41988 695187
rect 42112 694211 42146 695187
rect 42270 694211 42304 695187
rect 42428 694211 42462 695187
rect 42586 694211 42620 695187
rect 42744 694211 42778 695187
rect 42902 694211 42936 695187
rect 43060 694211 43094 695187
rect 43218 694211 43252 695187
rect 43376 694211 43410 695187
rect 43534 694211 43568 695187
rect 43692 694211 43726 695187
rect 43850 694211 43884 695187
rect 44008 694211 44042 695187
rect 44166 694211 44200 695187
rect 44324 694211 44358 695187
rect 44482 694211 44516 695187
rect 44640 694211 44674 695187
rect 44798 694211 44832 695187
rect 44956 694211 44990 695187
rect 45114 694211 45148 695187
rect 45272 694211 45306 695187
rect 45430 694211 45464 695187
rect 45588 694211 45622 695187
rect 45746 694211 45780 695187
rect 45904 694211 45938 695187
rect 46062 694211 46096 695187
rect 46220 694211 46254 695187
rect 46378 694211 46412 695187
rect 46536 694211 46570 695187
rect 46694 694211 46728 695187
rect 46852 694211 46886 695187
rect 47010 694211 47044 695187
rect 47168 694211 47202 695187
rect 47326 694211 47360 695187
rect 47484 694211 47518 695187
rect 47642 694211 47676 695187
rect 47800 694211 47834 695187
rect 42980 692541 43014 693517
rect 43138 692541 43172 693517
rect 43296 692541 43330 693517
rect 43454 692541 43488 693517
rect 43612 692541 43646 693517
rect 43770 692541 43804 693517
rect 43928 692541 43962 693517
rect 44086 692541 44120 693517
rect 44244 692541 44278 693517
rect 44402 692541 44436 693517
rect 44560 692541 44594 693517
rect 44718 692541 44752 693517
rect 44876 692541 44910 693517
rect 45034 692541 45068 693517
rect 45192 692541 45226 693517
rect 45350 692541 45384 693517
rect 45508 692541 45542 693517
rect 45666 692541 45700 693517
rect 45824 692541 45858 693517
rect 45982 692541 46016 693517
rect 46140 692541 46174 693517
rect 46298 692541 46332 693517
rect 42980 691001 43014 691977
rect 43138 691001 43172 691977
rect 43296 691001 43330 691977
rect 43454 691001 43488 691977
rect 43612 691001 43646 691977
rect 43770 691001 43804 691977
rect 43928 691001 43962 691977
rect 44086 691001 44120 691977
rect 44244 691001 44278 691977
rect 44402 691001 44436 691977
rect 44560 691001 44594 691977
rect 44718 691001 44752 691977
rect 44876 691001 44910 691977
rect 45034 691001 45068 691977
rect 45192 691001 45226 691977
rect 45350 691001 45384 691977
rect 45508 691001 45542 691977
rect 45666 691001 45700 691977
rect 45824 691001 45858 691977
rect 45982 691001 46016 691977
rect 46140 691001 46174 691977
rect 46298 691001 46332 691977
rect 540380 690750 541356 690784
rect 541616 690750 542592 690784
rect 542852 690750 543828 690784
rect 544088 690750 545064 690784
rect 545324 690750 546300 690784
rect 546560 690750 547536 690784
rect 547796 690750 548772 690784
rect 540380 690592 541356 690626
rect 541616 690592 542592 690626
rect 542852 690592 543828 690626
rect 544088 690592 545064 690626
rect 545324 690592 546300 690626
rect 546560 690592 547536 690626
rect 547796 690592 548772 690626
rect 540380 690210 541356 690244
rect 541616 690210 542592 690244
rect 542852 690210 543828 690244
rect 544088 690210 545064 690244
rect 545324 690210 546300 690244
rect 546560 690210 547536 690244
rect 547796 690210 548772 690244
rect 540380 690052 541356 690086
rect 541616 690052 542592 690086
rect 542852 690052 543828 690086
rect 544088 690052 545064 690086
rect 545324 690052 546300 690086
rect 546560 690052 547536 690086
rect 547796 690052 548772 690086
rect 540380 689670 541356 689704
rect 541616 689670 542592 689704
rect 542852 689670 543828 689704
rect 544088 689670 545064 689704
rect 545324 689670 546300 689704
rect 546560 689670 547536 689704
rect 547796 689670 548772 689704
rect 540380 689512 541356 689546
rect 541616 689512 542592 689546
rect 542852 689512 543828 689546
rect 544088 689512 545064 689546
rect 545324 689512 546300 689546
rect 546560 689512 547536 689546
rect 547796 689512 548772 689546
rect 540380 689130 541356 689164
rect 541616 689130 542592 689164
rect 542852 689130 543828 689164
rect 544088 689130 545064 689164
rect 545324 689130 546300 689164
rect 546560 689130 547536 689164
rect 547796 689130 548772 689164
rect 540380 688972 541356 689006
rect 541616 688972 542592 689006
rect 542852 688972 543828 689006
rect 544088 688972 545064 689006
rect 545324 688972 546300 689006
rect 546560 688972 547536 689006
rect 547796 688972 548772 689006
rect 540380 688550 541356 688584
rect 541616 688550 542592 688584
rect 542852 688550 543828 688584
rect 544088 688550 545064 688584
rect 545324 688550 546300 688584
rect 546560 688550 547536 688584
rect 547796 688550 548772 688584
rect 540380 688392 541356 688426
rect 541616 688392 542592 688426
rect 542852 688392 543828 688426
rect 544088 688392 545064 688426
rect 545324 688392 546300 688426
rect 546560 688392 547536 688426
rect 547796 688392 548772 688426
rect 540380 687970 541356 688004
rect 541616 687970 542592 688004
rect 542852 687970 543828 688004
rect 544088 687970 545064 688004
rect 545324 687970 546300 688004
rect 546560 687970 547536 688004
rect 547796 687970 548772 688004
rect 540380 687812 541356 687846
rect 541616 687812 542592 687846
rect 542852 687812 543828 687846
rect 544088 687812 545064 687846
rect 545324 687812 546300 687846
rect 546560 687812 547536 687846
rect 547796 687812 548772 687846
rect 538540 687430 539516 687464
rect 539776 687430 540752 687464
rect 541012 687430 541988 687464
rect 542248 687430 543224 687464
rect 543484 687430 544460 687464
rect 544720 687430 545696 687464
rect 545956 687430 546932 687464
rect 547192 687430 548168 687464
rect 548428 687430 549404 687464
rect 549664 687430 550640 687464
rect 538540 687272 539516 687306
rect 539776 687272 540752 687306
rect 541012 687272 541988 687306
rect 542248 687272 543224 687306
rect 543484 687272 544460 687306
rect 544720 687272 545696 687306
rect 545956 687272 546932 687306
rect 547192 687272 548168 687306
rect 548428 687272 549404 687306
rect 549664 687272 550640 687306
rect 538540 686890 539516 686924
rect 539776 686890 540752 686924
rect 541012 686890 541988 686924
rect 542248 686890 543224 686924
rect 543484 686890 544460 686924
rect 544720 686890 545696 686924
rect 545956 686890 546932 686924
rect 547192 686890 548168 686924
rect 548428 686890 549404 686924
rect 549664 686890 550640 686924
rect 538540 686732 539516 686766
rect 539776 686732 540752 686766
rect 541012 686732 541988 686766
rect 542248 686732 543224 686766
rect 543484 686732 544460 686766
rect 544720 686732 545696 686766
rect 545956 686732 546932 686766
rect 547192 686732 548168 686766
rect 548428 686732 549404 686766
rect 549664 686732 550640 686766
rect 538540 686350 539516 686384
rect 539776 686350 540752 686384
rect 541012 686350 541988 686384
rect 542248 686350 543224 686384
rect 543484 686350 544460 686384
rect 544720 686350 545696 686384
rect 545956 686350 546932 686384
rect 547192 686350 548168 686384
rect 548428 686350 549404 686384
rect 549664 686350 550640 686384
rect 538540 686192 539516 686226
rect 539776 686192 540752 686226
rect 541012 686192 541988 686226
rect 542248 686192 543224 686226
rect 543484 686192 544460 686226
rect 544720 686192 545696 686226
rect 545956 686192 546932 686226
rect 547192 686192 548168 686226
rect 548428 686192 549404 686226
rect 549664 686192 550640 686226
rect 538540 685810 539516 685844
rect 539776 685810 540752 685844
rect 541012 685810 541988 685844
rect 542248 685810 543224 685844
rect 543484 685810 544460 685844
rect 544720 685810 545696 685844
rect 545956 685810 546932 685844
rect 547192 685810 548168 685844
rect 548428 685810 549404 685844
rect 549664 685810 550640 685844
rect 538540 685652 539516 685686
rect 539776 685652 540752 685686
rect 541012 685652 541988 685686
rect 542248 685652 543224 685686
rect 543484 685652 544460 685686
rect 544720 685652 545696 685686
rect 545956 685652 546932 685686
rect 547192 685652 548168 685686
rect 548428 685652 549404 685686
rect 549664 685652 550640 685686
rect 43860 682831 43894 683807
rect 44118 682831 44152 683807
rect 44376 682831 44410 683807
rect 44634 682831 44668 683807
rect 44892 682831 44926 683807
rect 45150 682831 45184 683807
rect 45408 682831 45442 683807
rect 43860 681331 43894 682307
rect 44118 681331 44152 682307
rect 44376 681331 44410 682307
rect 44634 681331 44668 682307
rect 44892 681331 44926 682307
rect 45150 681331 45184 682307
rect 45408 681331 45442 682307
rect 541025 681236 542001 681270
rect 542261 681236 543237 681270
rect 543497 681236 544473 681270
rect 544733 681236 545709 681270
rect 545969 681236 546945 681270
rect 547205 681236 548181 681270
rect 541025 680978 542001 681012
rect 542261 680978 543237 681012
rect 543497 680978 544473 681012
rect 544733 680978 545709 681012
rect 545969 680978 546945 681012
rect 547205 680978 548181 681012
rect 541025 680646 542001 680680
rect 542261 680646 543237 680680
rect 543497 680646 544473 680680
rect 544733 680646 545709 680680
rect 545969 680646 546945 680680
rect 547205 680646 548181 680680
rect 541025 680388 542001 680422
rect 542261 680388 543237 680422
rect 543497 680388 544473 680422
rect 544733 680388 545709 680422
rect 545969 680388 546945 680422
rect 547205 680388 548181 680422
<< psubdiff >>
rect 37563 696225 37659 696259
rect 40591 696225 40687 696259
rect 37563 696163 37597 696225
rect 40653 696163 40687 696225
rect 37563 694887 37597 694949
rect 48633 696225 48729 696259
rect 51661 696225 51757 696259
rect 48633 696163 48667 696225
rect 40653 694887 40687 694949
rect 37563 694853 37659 694887
rect 40591 694853 40687 694887
rect 37563 694765 37659 694799
rect 40591 694765 40687 694799
rect 37563 694703 37597 694765
rect 40653 694703 40687 694765
rect 37563 693427 37597 693489
rect 51723 696163 51757 696225
rect 48633 694887 48667 694949
rect 51723 694887 51757 694949
rect 48633 694853 48729 694887
rect 51661 694853 51757 694887
rect 48633 694765 48729 694799
rect 51661 694765 51757 694799
rect 48633 694703 48667 694765
rect 40653 693427 40687 693489
rect 37563 693393 37659 693427
rect 40591 693393 40687 693427
rect 51723 694703 51757 694765
rect 48633 693427 48667 693489
rect 51723 693427 51757 693489
rect 48633 693393 48729 693427
rect 51661 693393 51757 693427
rect 43967 690561 44063 690595
rect 45239 690561 45335 690595
rect 43967 690499 44001 690561
rect 45301 690499 45335 690561
rect 43967 689281 44001 689343
rect 45301 689281 45335 689343
rect 43967 689247 44063 689281
rect 45239 689247 45335 689281
rect 43967 689041 44063 689075
rect 45239 689041 45335 689075
rect 43967 688979 44001 689041
rect 45301 688979 45335 689041
rect 43967 687761 44001 687823
rect 45301 687761 45335 687823
rect 43967 687727 44063 687761
rect 45239 687727 45335 687761
rect 534592 688067 534688 688101
rect 537620 688067 537716 688101
rect 534592 688005 534626 688067
rect 42976 687520 43072 687554
rect 46238 687520 46334 687554
rect 42976 687458 43010 687520
rect 46300 687458 46334 687520
rect 42976 686240 43010 686302
rect 537682 688005 537716 688067
rect 534592 686729 534626 686791
rect 551652 688067 551748 688101
rect 554680 688067 554776 688101
rect 551652 688005 551686 688067
rect 537682 686729 537716 686791
rect 534592 686695 534688 686729
rect 537620 686695 537716 686729
rect 554742 688005 554776 688067
rect 551652 686729 551686 686791
rect 554742 686729 554776 686791
rect 551652 686695 551748 686729
rect 554680 686695 554776 686729
rect 46300 686240 46334 686302
rect 42976 686206 43072 686240
rect 46238 686206 46334 686240
rect 534592 686597 534688 686631
rect 537620 686597 537716 686631
rect 534592 686535 534626 686597
rect 42716 686000 42812 686034
rect 46494 686000 46590 686034
rect 42716 685938 42750 686000
rect 46556 685938 46590 686000
rect 42716 684720 42750 684782
rect 537682 686535 537716 686597
rect 534592 685259 534626 685321
rect 551652 686597 551748 686631
rect 554680 686597 554776 686631
rect 551652 686535 551686 686597
rect 537682 685259 537716 685321
rect 534592 685225 534688 685259
rect 537620 685225 537716 685259
rect 554742 686535 554776 686597
rect 551652 685259 551686 685321
rect 554742 685259 554776 685321
rect 551652 685225 551748 685259
rect 554680 685225 554776 685259
rect 46556 684720 46590 684782
rect 540285 685144 540381 685178
rect 548845 685144 548941 685178
rect 540285 685082 540319 685144
rect 548907 685082 548941 685144
rect 540285 684792 540319 684854
rect 548907 684792 548941 684854
rect 540285 684758 540381 684792
rect 548845 684758 548941 684792
rect 42716 684686 42812 684720
rect 46494 684686 46590 684720
rect 540285 684644 540381 684678
rect 548845 684644 548941 684678
rect 540285 684582 540319 684644
rect 548907 684582 548941 684644
rect 540285 684292 540319 684354
rect 548907 684292 548941 684354
rect 540285 684258 540381 684292
rect 548845 684258 548941 684292
rect 540845 684144 540941 684178
rect 548187 684144 548283 684178
rect 540845 684082 540879 684144
rect 548249 684082 548283 684144
rect 540845 683692 540879 683754
rect 548249 683692 548283 683754
rect 540845 683658 540941 683692
rect 548187 683658 548283 683692
rect 540845 683524 540941 683558
rect 548187 683524 548283 683558
rect 540845 683462 540879 683524
rect 548249 683462 548283 683524
rect 540845 683072 540879 683134
rect 548249 683072 548283 683134
rect 540845 683038 540941 683072
rect 548187 683038 548283 683072
rect 540285 682924 540381 682958
rect 548845 682924 548941 682958
rect 540285 682862 540319 682924
rect 548907 682862 548941 682924
rect 540285 682472 540319 682534
rect 548907 682472 548941 682534
rect 540285 682438 540381 682472
rect 548845 682438 548941 682472
rect 540285 682324 540381 682358
rect 548845 682324 548941 682358
rect 540285 682262 540319 682324
rect 548907 682262 548941 682324
rect 540285 681872 540319 681934
rect 548907 681872 548941 681934
rect 540285 681838 540381 681872
rect 548845 681838 548941 681872
rect 44346 680850 44442 680884
rect 44828 680850 44924 680884
rect 44346 680788 44380 680850
rect 44890 680788 44924 680850
rect 44346 680070 44380 680132
rect 44890 680070 44924 680132
rect 44346 680036 44442 680070
rect 44828 680036 44924 680070
rect 543600 679970 543696 680004
rect 545506 679970 545602 680004
rect 543600 679908 543634 679970
rect 43986 679850 44082 679884
rect 45184 679850 45280 679884
rect 43986 679788 44020 679850
rect 45246 679788 45280 679850
rect 43986 679320 44020 679382
rect 545568 679908 545602 679970
rect 543600 679518 543634 679580
rect 545568 679518 545602 679580
rect 543600 679484 543696 679518
rect 545506 679484 545602 679518
rect 45246 679320 45280 679382
rect 43986 679286 44082 679320
rect 45184 679286 45280 679320
rect 543820 679345 543916 679379
rect 545290 679345 545386 679379
rect 543820 679283 543854 679345
rect 43731 679100 43827 679134
rect 45445 679100 45541 679134
rect 43731 679038 43765 679100
rect 45507 679038 45541 679100
rect 43731 677820 43765 677882
rect 545352 679283 545386 679345
rect 543820 678993 543854 679055
rect 545352 678993 545386 679055
rect 543820 678959 543916 678993
rect 545290 678959 545386 678993
rect 540885 678820 540981 678854
rect 548227 678820 548323 678854
rect 540885 678758 540919 678820
rect 548289 678758 548323 678820
rect 540885 678368 540919 678430
rect 548289 678368 548323 678430
rect 540885 678334 540981 678368
rect 548227 678334 548323 678368
rect 45507 677820 45541 677882
rect 43731 677786 43827 677820
rect 45445 677786 45541 677820
rect 41200 676980 41440 677004
rect 41200 676716 41440 676740
rect 41200 675260 41440 675284
rect 41200 674996 41440 675020
rect 41200 673540 41440 673564
rect 41200 673276 41440 673300
rect 41200 672060 41440 672084
rect 41200 671796 41440 671820
rect 41200 670340 41440 670364
rect 41200 670076 41440 670100
rect 41200 668740 41440 668764
rect 41200 668476 41440 668500
rect 41200 667020 41440 667044
rect 41200 666756 41440 666780
rect 41200 665420 41440 665444
rect 41200 665156 41440 665180
rect 41200 663700 41440 663724
rect 41200 663436 41440 663460
rect 541364 677058 541484 677082
rect 47900 676980 48140 677004
rect 541364 676914 541484 676938
rect 47900 676716 48140 676740
rect 47900 675260 48140 675284
rect 47900 674996 48140 675020
rect 541364 674058 541484 674082
rect 541364 673914 541484 673938
rect 47900 673540 48140 673564
rect 47900 673276 48140 673300
rect 47900 672060 48140 672084
rect 47900 671796 48140 671820
rect 541364 671058 541484 671082
rect 541364 670914 541484 670938
rect 47900 670340 48140 670364
rect 47900 670076 48140 670100
rect 47900 668740 48140 668764
rect 47900 668476 48140 668500
rect 541364 668058 541484 668082
rect 541364 667914 541484 667938
rect 47900 667020 48140 667044
rect 47900 666756 48140 666780
rect 47900 665420 48140 665444
rect 47900 665156 48140 665180
rect 541364 665058 541484 665082
rect 541364 664914 541484 664938
rect 47900 663700 48140 663724
rect 47900 663436 48140 663460
rect 547734 677058 547854 677082
rect 547734 676914 547854 676938
rect 547734 674058 547854 674082
rect 547734 673914 547854 673938
rect 547734 671058 547854 671082
rect 547734 670914 547854 670938
rect 547734 668058 547854 668082
rect 547734 667914 547854 667938
rect 547734 665058 547854 665082
rect 547734 664914 547854 664938
<< nsubdiff >>
rect 41366 695348 41462 695382
rect 47852 695348 47948 695382
rect 41366 695286 41400 695348
rect 47914 695286 47948 695348
rect 41366 694050 41400 694112
rect 47914 694050 47948 694112
rect 41366 694016 41462 694050
rect 47852 694016 47948 694050
rect 42866 693678 42962 693712
rect 46350 693678 46446 693712
rect 42866 693616 42900 693678
rect 46412 693616 46446 693678
rect 42866 692380 42900 692442
rect 46412 692380 46446 692442
rect 42866 692346 42962 692380
rect 46350 692346 46446 692380
rect 42866 692138 42962 692172
rect 46350 692138 46446 692172
rect 42866 692076 42900 692138
rect 46412 692076 46446 692138
rect 42866 690840 42900 690902
rect 46412 690840 46446 690902
rect 42866 690806 42962 690840
rect 46350 690806 46446 690840
rect 540185 690864 540281 690898
rect 548871 690864 548967 690898
rect 540185 690802 540219 690864
rect 548933 690802 548967 690864
rect 540185 690512 540219 690574
rect 548933 690512 548967 690574
rect 540185 690478 540281 690512
rect 548871 690478 548967 690512
rect 540185 690324 540281 690358
rect 548871 690324 548967 690358
rect 540185 690262 540219 690324
rect 548933 690262 548967 690324
rect 540185 689972 540219 690034
rect 548933 689972 548967 690034
rect 540185 689938 540281 689972
rect 548871 689938 548967 689972
rect 540185 689784 540281 689818
rect 548871 689784 548967 689818
rect 540185 689722 540219 689784
rect 548933 689722 548967 689784
rect 540185 689432 540219 689494
rect 548933 689432 548967 689494
rect 540185 689398 540281 689432
rect 548871 689398 548967 689432
rect 540185 689244 540281 689278
rect 548871 689244 548967 689278
rect 540185 689182 540219 689244
rect 548933 689182 548967 689244
rect 540185 688892 540219 688954
rect 548933 688892 548967 688954
rect 540185 688858 540281 688892
rect 548871 688858 548967 688892
rect 540185 688664 540281 688698
rect 548871 688664 548967 688698
rect 540185 688602 540219 688664
rect 548933 688602 548967 688664
rect 540185 688312 540219 688374
rect 548933 688312 548967 688374
rect 540185 688278 540281 688312
rect 548871 688278 548967 688312
rect 540185 688084 540281 688118
rect 548871 688084 548967 688118
rect 540185 688022 540219 688084
rect 548933 688022 548967 688084
rect 540185 687732 540219 687794
rect 548933 687732 548967 687794
rect 540185 687698 540281 687732
rect 548871 687698 548967 687732
rect 538345 687544 538441 687578
rect 550739 687544 550835 687578
rect 538345 687482 538379 687544
rect 550801 687482 550835 687544
rect 538345 687192 538379 687254
rect 550801 687192 550835 687254
rect 538345 687158 538441 687192
rect 550739 687158 550835 687192
rect 538345 687004 538441 687038
rect 550739 687004 550835 687038
rect 538345 686942 538379 687004
rect 550801 686942 550835 687004
rect 538345 686652 538379 686714
rect 550801 686652 550835 686714
rect 538345 686618 538441 686652
rect 550739 686618 550835 686652
rect 538345 686464 538441 686498
rect 550739 686464 550835 686498
rect 538345 686402 538379 686464
rect 550801 686402 550835 686464
rect 538345 686112 538379 686174
rect 550801 686112 550835 686174
rect 538345 686078 538441 686112
rect 550739 686078 550835 686112
rect 538345 685924 538441 685958
rect 550739 685924 550835 685958
rect 538345 685862 538379 685924
rect 550801 685862 550835 685924
rect 538345 685572 538379 685634
rect 550801 685572 550835 685634
rect 538345 685538 538441 685572
rect 550739 685538 550835 685572
rect 43746 683968 43842 684002
rect 45460 683968 45556 684002
rect 43746 683906 43780 683968
rect 45522 683906 45556 683968
rect 43746 682670 43780 682732
rect 45522 682670 45556 682732
rect 43746 682636 43842 682670
rect 45460 682636 45556 682670
rect 43746 682468 43842 682502
rect 45460 682468 45556 682502
rect 43746 682406 43780 682468
rect 45522 682406 45556 682468
rect 43746 681170 43780 681232
rect 45522 681170 45556 681232
rect 43746 681136 43842 681170
rect 45460 681136 45556 681170
rect 540830 681350 540926 681384
rect 548280 681350 548376 681384
rect 540830 681288 540864 681350
rect 548342 681288 548376 681350
rect 540830 680898 540864 680960
rect 548342 680898 548376 680960
rect 540830 680864 540926 680898
rect 548280 680864 548376 680898
rect 540830 680760 540926 680794
rect 548280 680760 548376 680794
rect 540830 680698 540864 680760
rect 548342 680698 548376 680760
rect 540830 680308 540864 680370
rect 548342 680308 548376 680370
rect 540830 680274 540926 680308
rect 548280 680274 548376 680308
<< psubdiffcont >>
rect 37659 696225 40591 696259
rect 37563 694949 37597 696163
rect 40653 694949 40687 696163
rect 48729 696225 51661 696259
rect 37659 694853 40591 694887
rect 37659 694765 40591 694799
rect 37563 693489 37597 694703
rect 40653 693489 40687 694703
rect 48633 694949 48667 696163
rect 51723 694949 51757 696163
rect 48729 694853 51661 694887
rect 48729 694765 51661 694799
rect 37659 693393 40591 693427
rect 48633 693489 48667 694703
rect 51723 693489 51757 694703
rect 48729 693393 51661 693427
rect 44063 690561 45239 690595
rect 43967 689343 44001 690499
rect 45301 689343 45335 690499
rect 44063 689247 45239 689281
rect 44063 689041 45239 689075
rect 43967 687823 44001 688979
rect 45301 687823 45335 688979
rect 44063 687727 45239 687761
rect 534688 688067 537620 688101
rect 43072 687520 46238 687554
rect 42976 686302 43010 687458
rect 46300 686302 46334 687458
rect 534592 686791 534626 688005
rect 537682 686791 537716 688005
rect 551748 688067 554680 688101
rect 534688 686695 537620 686729
rect 551652 686791 551686 688005
rect 554742 686791 554776 688005
rect 551748 686695 554680 686729
rect 43072 686206 46238 686240
rect 534688 686597 537620 686631
rect 42812 686000 46494 686034
rect 42716 684782 42750 685938
rect 46556 684782 46590 685938
rect 534592 685321 534626 686535
rect 537682 685321 537716 686535
rect 551748 686597 554680 686631
rect 534688 685225 537620 685259
rect 551652 685321 551686 686535
rect 554742 685321 554776 686535
rect 551748 685225 554680 685259
rect 540381 685144 548845 685178
rect 540285 684854 540319 685082
rect 548907 684854 548941 685082
rect 540381 684758 548845 684792
rect 42812 684686 46494 684720
rect 540381 684644 548845 684678
rect 540285 684354 540319 684582
rect 548907 684354 548941 684582
rect 540381 684258 548845 684292
rect 540941 684144 548187 684178
rect 540845 683754 540879 684082
rect 548249 683754 548283 684082
rect 540941 683658 548187 683692
rect 540941 683524 548187 683558
rect 540845 683134 540879 683462
rect 548249 683134 548283 683462
rect 540941 683038 548187 683072
rect 540381 682924 548845 682958
rect 540285 682534 540319 682862
rect 548907 682534 548941 682862
rect 540381 682438 548845 682472
rect 540381 682324 548845 682358
rect 540285 681934 540319 682262
rect 548907 681934 548941 682262
rect 540381 681838 548845 681872
rect 44442 680850 44828 680884
rect 44346 680132 44380 680788
rect 44890 680132 44924 680788
rect 44442 680036 44828 680070
rect 543696 679970 545506 680004
rect 44082 679850 45184 679884
rect 43986 679382 44020 679788
rect 45246 679382 45280 679788
rect 543600 679580 543634 679908
rect 545568 679580 545602 679908
rect 543696 679484 545506 679518
rect 44082 679286 45184 679320
rect 543916 679345 545290 679379
rect 43827 679100 45445 679134
rect 43731 677882 43765 679038
rect 45507 677882 45541 679038
rect 543820 679055 543854 679283
rect 545352 679055 545386 679283
rect 543916 678959 545290 678993
rect 540981 678820 548227 678854
rect 540885 678430 540919 678758
rect 548289 678430 548323 678758
rect 540981 678334 548227 678368
rect 43827 677786 45445 677820
rect 41200 676740 41440 676980
rect 41200 675020 41440 675260
rect 41200 673300 41440 673540
rect 41200 671820 41440 672060
rect 41200 670100 41440 670340
rect 41200 668500 41440 668740
rect 41200 666780 41440 667020
rect 41200 665180 41440 665420
rect 41200 663460 41440 663700
rect 47900 676740 48140 676980
rect 541364 676938 541484 677058
rect 47900 675020 48140 675260
rect 541364 673938 541484 674058
rect 47900 673300 48140 673540
rect 47900 671820 48140 672060
rect 541364 670938 541484 671058
rect 47900 670100 48140 670340
rect 47900 668500 48140 668740
rect 541364 667938 541484 668058
rect 47900 666780 48140 667020
rect 47900 665180 48140 665420
rect 541364 664938 541484 665058
rect 47900 663460 48140 663700
rect 547734 676938 547854 677058
rect 547734 673938 547854 674058
rect 547734 670938 547854 671058
rect 547734 667938 547854 668058
rect 547734 664938 547854 665058
<< nsubdiffcont >>
rect 41462 695348 47852 695382
rect 41366 694112 41400 695286
rect 47914 694112 47948 695286
rect 41462 694016 47852 694050
rect 42962 693678 46350 693712
rect 42866 692442 42900 693616
rect 46412 692442 46446 693616
rect 42962 692346 46350 692380
rect 42962 692138 46350 692172
rect 42866 690902 42900 692076
rect 46412 690902 46446 692076
rect 42962 690806 46350 690840
rect 540281 690864 548871 690898
rect 540185 690574 540219 690802
rect 548933 690574 548967 690802
rect 540281 690478 548871 690512
rect 540281 690324 548871 690358
rect 540185 690034 540219 690262
rect 548933 690034 548967 690262
rect 540281 689938 548871 689972
rect 540281 689784 548871 689818
rect 540185 689494 540219 689722
rect 548933 689494 548967 689722
rect 540281 689398 548871 689432
rect 540281 689244 548871 689278
rect 540185 688954 540219 689182
rect 548933 688954 548967 689182
rect 540281 688858 548871 688892
rect 540281 688664 548871 688698
rect 540185 688374 540219 688602
rect 548933 688374 548967 688602
rect 540281 688278 548871 688312
rect 540281 688084 548871 688118
rect 540185 687794 540219 688022
rect 548933 687794 548967 688022
rect 540281 687698 548871 687732
rect 538441 687544 550739 687578
rect 538345 687254 538379 687482
rect 550801 687254 550835 687482
rect 538441 687158 550739 687192
rect 538441 687004 550739 687038
rect 538345 686714 538379 686942
rect 550801 686714 550835 686942
rect 538441 686618 550739 686652
rect 538441 686464 550739 686498
rect 538345 686174 538379 686402
rect 550801 686174 550835 686402
rect 538441 686078 550739 686112
rect 538441 685924 550739 685958
rect 538345 685634 538379 685862
rect 550801 685634 550835 685862
rect 538441 685538 550739 685572
rect 43842 683968 45460 684002
rect 43746 682732 43780 683906
rect 45522 682732 45556 683906
rect 43842 682636 45460 682670
rect 43842 682468 45460 682502
rect 43746 681232 43780 682406
rect 45522 681232 45556 682406
rect 43842 681136 45460 681170
rect 540926 681350 548280 681384
rect 540830 680960 540864 681288
rect 548342 680960 548376 681288
rect 540926 680864 548280 680898
rect 540926 680760 548280 680794
rect 540830 680370 540864 680698
rect 548342 680370 548376 680698
rect 540926 680274 548280 680308
<< poly >>
rect 41526 695280 41626 695296
rect 41526 695246 41542 695280
rect 41610 695246 41626 695280
rect 41526 695199 41626 695246
rect 41684 695280 41784 695296
rect 41684 695246 41700 695280
rect 41768 695246 41784 695280
rect 41684 695199 41784 695246
rect 41842 695280 41942 695296
rect 41842 695246 41858 695280
rect 41926 695246 41942 695280
rect 41842 695199 41942 695246
rect 42000 695280 42100 695296
rect 42000 695246 42016 695280
rect 42084 695246 42100 695280
rect 42000 695199 42100 695246
rect 42158 695280 42258 695296
rect 42158 695246 42174 695280
rect 42242 695246 42258 695280
rect 42158 695199 42258 695246
rect 42316 695280 42416 695296
rect 42316 695246 42332 695280
rect 42400 695246 42416 695280
rect 42316 695199 42416 695246
rect 42474 695280 42574 695296
rect 42474 695246 42490 695280
rect 42558 695246 42574 695280
rect 42474 695199 42574 695246
rect 42632 695280 42732 695296
rect 42632 695246 42648 695280
rect 42716 695246 42732 695280
rect 42632 695199 42732 695246
rect 42790 695280 42890 695296
rect 42790 695246 42806 695280
rect 42874 695246 42890 695280
rect 42790 695199 42890 695246
rect 42948 695280 43048 695296
rect 42948 695246 42964 695280
rect 43032 695246 43048 695280
rect 42948 695199 43048 695246
rect 43106 695280 43206 695296
rect 43106 695246 43122 695280
rect 43190 695246 43206 695280
rect 43106 695199 43206 695246
rect 43264 695280 43364 695296
rect 43264 695246 43280 695280
rect 43348 695246 43364 695280
rect 43264 695199 43364 695246
rect 43422 695280 43522 695296
rect 43422 695246 43438 695280
rect 43506 695246 43522 695280
rect 43422 695199 43522 695246
rect 43580 695280 43680 695296
rect 43580 695246 43596 695280
rect 43664 695246 43680 695280
rect 43580 695199 43680 695246
rect 43738 695280 43838 695296
rect 43738 695246 43754 695280
rect 43822 695246 43838 695280
rect 43738 695199 43838 695246
rect 43896 695280 43996 695296
rect 43896 695246 43912 695280
rect 43980 695246 43996 695280
rect 43896 695199 43996 695246
rect 44054 695280 44154 695296
rect 44054 695246 44070 695280
rect 44138 695246 44154 695280
rect 44054 695199 44154 695246
rect 44212 695280 44312 695296
rect 44212 695246 44228 695280
rect 44296 695246 44312 695280
rect 44212 695199 44312 695246
rect 44370 695280 44470 695296
rect 44370 695246 44386 695280
rect 44454 695246 44470 695280
rect 44370 695199 44470 695246
rect 44528 695280 44628 695296
rect 44528 695246 44544 695280
rect 44612 695246 44628 695280
rect 44528 695199 44628 695246
rect 44686 695280 44786 695296
rect 44686 695246 44702 695280
rect 44770 695246 44786 695280
rect 44686 695199 44786 695246
rect 44844 695280 44944 695296
rect 44844 695246 44860 695280
rect 44928 695246 44944 695280
rect 44844 695199 44944 695246
rect 45002 695280 45102 695296
rect 45002 695246 45018 695280
rect 45086 695246 45102 695280
rect 45002 695199 45102 695246
rect 45160 695280 45260 695296
rect 45160 695246 45176 695280
rect 45244 695246 45260 695280
rect 45160 695199 45260 695246
rect 45318 695280 45418 695296
rect 45318 695246 45334 695280
rect 45402 695246 45418 695280
rect 45318 695199 45418 695246
rect 45476 695280 45576 695296
rect 45476 695246 45492 695280
rect 45560 695246 45576 695280
rect 45476 695199 45576 695246
rect 45634 695280 45734 695296
rect 45634 695246 45650 695280
rect 45718 695246 45734 695280
rect 45634 695199 45734 695246
rect 45792 695280 45892 695296
rect 45792 695246 45808 695280
rect 45876 695246 45892 695280
rect 45792 695199 45892 695246
rect 45950 695280 46050 695296
rect 45950 695246 45966 695280
rect 46034 695246 46050 695280
rect 45950 695199 46050 695246
rect 46108 695280 46208 695296
rect 46108 695246 46124 695280
rect 46192 695246 46208 695280
rect 46108 695199 46208 695246
rect 46266 695280 46366 695296
rect 46266 695246 46282 695280
rect 46350 695246 46366 695280
rect 46266 695199 46366 695246
rect 46424 695280 46524 695296
rect 46424 695246 46440 695280
rect 46508 695246 46524 695280
rect 46424 695199 46524 695246
rect 46582 695280 46682 695296
rect 46582 695246 46598 695280
rect 46666 695246 46682 695280
rect 46582 695199 46682 695246
rect 46740 695280 46840 695296
rect 46740 695246 46756 695280
rect 46824 695246 46840 695280
rect 46740 695199 46840 695246
rect 46898 695280 46998 695296
rect 46898 695246 46914 695280
rect 46982 695246 46998 695280
rect 46898 695199 46998 695246
rect 47056 695280 47156 695296
rect 47056 695246 47072 695280
rect 47140 695246 47156 695280
rect 47056 695199 47156 695246
rect 47214 695280 47314 695296
rect 47214 695246 47230 695280
rect 47298 695246 47314 695280
rect 47214 695199 47314 695246
rect 47372 695280 47472 695296
rect 47372 695246 47388 695280
rect 47456 695246 47472 695280
rect 47372 695199 47472 695246
rect 47530 695280 47630 695296
rect 47530 695246 47546 695280
rect 47614 695246 47630 695280
rect 47530 695199 47630 695246
rect 47688 695280 47788 695296
rect 47688 695246 47704 695280
rect 47772 695246 47788 695280
rect 47688 695199 47788 695246
rect 41526 694152 41626 694199
rect 41526 694118 41542 694152
rect 41610 694118 41626 694152
rect 41526 694102 41626 694118
rect 41684 694152 41784 694199
rect 41684 694118 41700 694152
rect 41768 694118 41784 694152
rect 41684 694102 41784 694118
rect 41842 694152 41942 694199
rect 41842 694118 41858 694152
rect 41926 694118 41942 694152
rect 41842 694102 41942 694118
rect 42000 694152 42100 694199
rect 42000 694118 42016 694152
rect 42084 694118 42100 694152
rect 42000 694102 42100 694118
rect 42158 694152 42258 694199
rect 42158 694118 42174 694152
rect 42242 694118 42258 694152
rect 42158 694102 42258 694118
rect 42316 694152 42416 694199
rect 42316 694118 42332 694152
rect 42400 694118 42416 694152
rect 42316 694102 42416 694118
rect 42474 694152 42574 694199
rect 42474 694118 42490 694152
rect 42558 694118 42574 694152
rect 42474 694102 42574 694118
rect 42632 694152 42732 694199
rect 42632 694118 42648 694152
rect 42716 694118 42732 694152
rect 42632 694102 42732 694118
rect 42790 694152 42890 694199
rect 42790 694118 42806 694152
rect 42874 694118 42890 694152
rect 42790 694102 42890 694118
rect 42948 694152 43048 694199
rect 42948 694118 42964 694152
rect 43032 694118 43048 694152
rect 42948 694102 43048 694118
rect 43106 694152 43206 694199
rect 43106 694118 43122 694152
rect 43190 694118 43206 694152
rect 43106 694102 43206 694118
rect 43264 694152 43364 694199
rect 43264 694118 43280 694152
rect 43348 694118 43364 694152
rect 43264 694102 43364 694118
rect 43422 694152 43522 694199
rect 43422 694118 43438 694152
rect 43506 694118 43522 694152
rect 43422 694102 43522 694118
rect 43580 694152 43680 694199
rect 43580 694118 43596 694152
rect 43664 694118 43680 694152
rect 43580 694102 43680 694118
rect 43738 694152 43838 694199
rect 43738 694118 43754 694152
rect 43822 694118 43838 694152
rect 43738 694102 43838 694118
rect 43896 694152 43996 694199
rect 43896 694118 43912 694152
rect 43980 694118 43996 694152
rect 43896 694102 43996 694118
rect 44054 694152 44154 694199
rect 44054 694118 44070 694152
rect 44138 694118 44154 694152
rect 44054 694102 44154 694118
rect 44212 694152 44312 694199
rect 44212 694118 44228 694152
rect 44296 694118 44312 694152
rect 44212 694102 44312 694118
rect 44370 694152 44470 694199
rect 44370 694118 44386 694152
rect 44454 694118 44470 694152
rect 44370 694102 44470 694118
rect 44528 694152 44628 694199
rect 44528 694118 44544 694152
rect 44612 694118 44628 694152
rect 44528 694102 44628 694118
rect 44686 694152 44786 694199
rect 44686 694118 44702 694152
rect 44770 694118 44786 694152
rect 44686 694102 44786 694118
rect 44844 694152 44944 694199
rect 44844 694118 44860 694152
rect 44928 694118 44944 694152
rect 44844 694102 44944 694118
rect 45002 694152 45102 694199
rect 45002 694118 45018 694152
rect 45086 694118 45102 694152
rect 45002 694102 45102 694118
rect 45160 694152 45260 694199
rect 45160 694118 45176 694152
rect 45244 694118 45260 694152
rect 45160 694102 45260 694118
rect 45318 694152 45418 694199
rect 45318 694118 45334 694152
rect 45402 694118 45418 694152
rect 45318 694102 45418 694118
rect 45476 694152 45576 694199
rect 45476 694118 45492 694152
rect 45560 694118 45576 694152
rect 45476 694102 45576 694118
rect 45634 694152 45734 694199
rect 45634 694118 45650 694152
rect 45718 694118 45734 694152
rect 45634 694102 45734 694118
rect 45792 694152 45892 694199
rect 45792 694118 45808 694152
rect 45876 694118 45892 694152
rect 45792 694102 45892 694118
rect 45950 694152 46050 694199
rect 45950 694118 45966 694152
rect 46034 694118 46050 694152
rect 45950 694102 46050 694118
rect 46108 694152 46208 694199
rect 46108 694118 46124 694152
rect 46192 694118 46208 694152
rect 46108 694102 46208 694118
rect 46266 694152 46366 694199
rect 46266 694118 46282 694152
rect 46350 694118 46366 694152
rect 46266 694102 46366 694118
rect 46424 694152 46524 694199
rect 46424 694118 46440 694152
rect 46508 694118 46524 694152
rect 46424 694102 46524 694118
rect 46582 694152 46682 694199
rect 46582 694118 46598 694152
rect 46666 694118 46682 694152
rect 46582 694102 46682 694118
rect 46740 694152 46840 694199
rect 46740 694118 46756 694152
rect 46824 694118 46840 694152
rect 46740 694102 46840 694118
rect 46898 694152 46998 694199
rect 46898 694118 46914 694152
rect 46982 694118 46998 694152
rect 46898 694102 46998 694118
rect 47056 694152 47156 694199
rect 47056 694118 47072 694152
rect 47140 694118 47156 694152
rect 47056 694102 47156 694118
rect 47214 694152 47314 694199
rect 47214 694118 47230 694152
rect 47298 694118 47314 694152
rect 47214 694102 47314 694118
rect 47372 694152 47472 694199
rect 47372 694118 47388 694152
rect 47456 694118 47472 694152
rect 47372 694102 47472 694118
rect 47530 694152 47630 694199
rect 47530 694118 47546 694152
rect 47614 694118 47630 694152
rect 47530 694102 47630 694118
rect 47688 694152 47788 694199
rect 47688 694118 47704 694152
rect 47772 694118 47788 694152
rect 47688 694102 47788 694118
rect 43026 693610 43126 693626
rect 43026 693576 43042 693610
rect 43110 693576 43126 693610
rect 43026 693529 43126 693576
rect 43184 693610 43284 693626
rect 43184 693576 43200 693610
rect 43268 693576 43284 693610
rect 43184 693529 43284 693576
rect 43342 693610 43442 693626
rect 43342 693576 43358 693610
rect 43426 693576 43442 693610
rect 43342 693529 43442 693576
rect 43500 693610 43600 693626
rect 43500 693576 43516 693610
rect 43584 693576 43600 693610
rect 43500 693529 43600 693576
rect 43658 693610 43758 693626
rect 43658 693576 43674 693610
rect 43742 693576 43758 693610
rect 43658 693529 43758 693576
rect 43816 693610 43916 693626
rect 43816 693576 43832 693610
rect 43900 693576 43916 693610
rect 43816 693529 43916 693576
rect 43974 693610 44074 693626
rect 43974 693576 43990 693610
rect 44058 693576 44074 693610
rect 43974 693529 44074 693576
rect 44132 693610 44232 693626
rect 44132 693576 44148 693610
rect 44216 693576 44232 693610
rect 44132 693529 44232 693576
rect 44290 693610 44390 693626
rect 44290 693576 44306 693610
rect 44374 693576 44390 693610
rect 44290 693529 44390 693576
rect 44448 693610 44548 693626
rect 44448 693576 44464 693610
rect 44532 693576 44548 693610
rect 44448 693529 44548 693576
rect 44606 693610 44706 693626
rect 44606 693576 44622 693610
rect 44690 693576 44706 693610
rect 44606 693529 44706 693576
rect 44764 693610 44864 693626
rect 44764 693576 44780 693610
rect 44848 693576 44864 693610
rect 44764 693529 44864 693576
rect 44922 693610 45022 693626
rect 44922 693576 44938 693610
rect 45006 693576 45022 693610
rect 44922 693529 45022 693576
rect 45080 693610 45180 693626
rect 45080 693576 45096 693610
rect 45164 693576 45180 693610
rect 45080 693529 45180 693576
rect 45238 693610 45338 693626
rect 45238 693576 45254 693610
rect 45322 693576 45338 693610
rect 45238 693529 45338 693576
rect 45396 693610 45496 693626
rect 45396 693576 45412 693610
rect 45480 693576 45496 693610
rect 45396 693529 45496 693576
rect 45554 693610 45654 693626
rect 45554 693576 45570 693610
rect 45638 693576 45654 693610
rect 45554 693529 45654 693576
rect 45712 693610 45812 693626
rect 45712 693576 45728 693610
rect 45796 693576 45812 693610
rect 45712 693529 45812 693576
rect 45870 693610 45970 693626
rect 45870 693576 45886 693610
rect 45954 693576 45970 693610
rect 45870 693529 45970 693576
rect 46028 693610 46128 693626
rect 46028 693576 46044 693610
rect 46112 693576 46128 693610
rect 46028 693529 46128 693576
rect 46186 693610 46286 693626
rect 46186 693576 46202 693610
rect 46270 693576 46286 693610
rect 46186 693529 46286 693576
rect 43026 692482 43126 692529
rect 43026 692448 43042 692482
rect 43110 692448 43126 692482
rect 43026 692432 43126 692448
rect 43184 692482 43284 692529
rect 43184 692448 43200 692482
rect 43268 692448 43284 692482
rect 43184 692432 43284 692448
rect 43342 692482 43442 692529
rect 43342 692448 43358 692482
rect 43426 692448 43442 692482
rect 43342 692432 43442 692448
rect 43500 692482 43600 692529
rect 43500 692448 43516 692482
rect 43584 692448 43600 692482
rect 43500 692432 43600 692448
rect 43658 692482 43758 692529
rect 43658 692448 43674 692482
rect 43742 692448 43758 692482
rect 43658 692432 43758 692448
rect 43816 692482 43916 692529
rect 43816 692448 43832 692482
rect 43900 692448 43916 692482
rect 43816 692432 43916 692448
rect 43974 692482 44074 692529
rect 43974 692448 43990 692482
rect 44058 692448 44074 692482
rect 43974 692432 44074 692448
rect 44132 692482 44232 692529
rect 44132 692448 44148 692482
rect 44216 692448 44232 692482
rect 44132 692432 44232 692448
rect 44290 692482 44390 692529
rect 44290 692448 44306 692482
rect 44374 692448 44390 692482
rect 44290 692432 44390 692448
rect 44448 692482 44548 692529
rect 44448 692448 44464 692482
rect 44532 692448 44548 692482
rect 44448 692432 44548 692448
rect 44606 692482 44706 692529
rect 44606 692448 44622 692482
rect 44690 692448 44706 692482
rect 44606 692432 44706 692448
rect 44764 692482 44864 692529
rect 44764 692448 44780 692482
rect 44848 692448 44864 692482
rect 44764 692432 44864 692448
rect 44922 692482 45022 692529
rect 44922 692448 44938 692482
rect 45006 692448 45022 692482
rect 44922 692432 45022 692448
rect 45080 692482 45180 692529
rect 45080 692448 45096 692482
rect 45164 692448 45180 692482
rect 45080 692432 45180 692448
rect 45238 692482 45338 692529
rect 45238 692448 45254 692482
rect 45322 692448 45338 692482
rect 45238 692432 45338 692448
rect 45396 692482 45496 692529
rect 45396 692448 45412 692482
rect 45480 692448 45496 692482
rect 45396 692432 45496 692448
rect 45554 692482 45654 692529
rect 45554 692448 45570 692482
rect 45638 692448 45654 692482
rect 45554 692432 45654 692448
rect 45712 692482 45812 692529
rect 45712 692448 45728 692482
rect 45796 692448 45812 692482
rect 45712 692432 45812 692448
rect 45870 692482 45970 692529
rect 45870 692448 45886 692482
rect 45954 692448 45970 692482
rect 45870 692432 45970 692448
rect 46028 692482 46128 692529
rect 46028 692448 46044 692482
rect 46112 692448 46128 692482
rect 46028 692432 46128 692448
rect 46186 692482 46286 692529
rect 46186 692448 46202 692482
rect 46270 692448 46286 692482
rect 46186 692432 46286 692448
rect 43026 692070 43126 692086
rect 43026 692036 43042 692070
rect 43110 692036 43126 692070
rect 43026 691989 43126 692036
rect 43184 692070 43284 692086
rect 43184 692036 43200 692070
rect 43268 692036 43284 692070
rect 43184 691989 43284 692036
rect 43342 692070 43442 692086
rect 43342 692036 43358 692070
rect 43426 692036 43442 692070
rect 43342 691989 43442 692036
rect 43500 692070 43600 692086
rect 43500 692036 43516 692070
rect 43584 692036 43600 692070
rect 43500 691989 43600 692036
rect 43658 692070 43758 692086
rect 43658 692036 43674 692070
rect 43742 692036 43758 692070
rect 43658 691989 43758 692036
rect 43816 692070 43916 692086
rect 43816 692036 43832 692070
rect 43900 692036 43916 692070
rect 43816 691989 43916 692036
rect 43974 692070 44074 692086
rect 43974 692036 43990 692070
rect 44058 692036 44074 692070
rect 43974 691989 44074 692036
rect 44132 692070 44232 692086
rect 44132 692036 44148 692070
rect 44216 692036 44232 692070
rect 44132 691989 44232 692036
rect 44290 692070 44390 692086
rect 44290 692036 44306 692070
rect 44374 692036 44390 692070
rect 44290 691989 44390 692036
rect 44448 692070 44548 692086
rect 44448 692036 44464 692070
rect 44532 692036 44548 692070
rect 44448 691989 44548 692036
rect 44606 692070 44706 692086
rect 44606 692036 44622 692070
rect 44690 692036 44706 692070
rect 44606 691989 44706 692036
rect 44764 692070 44864 692086
rect 44764 692036 44780 692070
rect 44848 692036 44864 692070
rect 44764 691989 44864 692036
rect 44922 692070 45022 692086
rect 44922 692036 44938 692070
rect 45006 692036 45022 692070
rect 44922 691989 45022 692036
rect 45080 692070 45180 692086
rect 45080 692036 45096 692070
rect 45164 692036 45180 692070
rect 45080 691989 45180 692036
rect 45238 692070 45338 692086
rect 45238 692036 45254 692070
rect 45322 692036 45338 692070
rect 45238 691989 45338 692036
rect 45396 692070 45496 692086
rect 45396 692036 45412 692070
rect 45480 692036 45496 692070
rect 45396 691989 45496 692036
rect 45554 692070 45654 692086
rect 45554 692036 45570 692070
rect 45638 692036 45654 692070
rect 45554 691989 45654 692036
rect 45712 692070 45812 692086
rect 45712 692036 45728 692070
rect 45796 692036 45812 692070
rect 45712 691989 45812 692036
rect 45870 692070 45970 692086
rect 45870 692036 45886 692070
rect 45954 692036 45970 692070
rect 45870 691989 45970 692036
rect 46028 692070 46128 692086
rect 46028 692036 46044 692070
rect 46112 692036 46128 692070
rect 46028 691989 46128 692036
rect 46186 692070 46286 692086
rect 46186 692036 46202 692070
rect 46270 692036 46286 692070
rect 46186 691989 46286 692036
rect 43026 690942 43126 690989
rect 43026 690908 43042 690942
rect 43110 690908 43126 690942
rect 43026 690892 43126 690908
rect 43184 690942 43284 690989
rect 43184 690908 43200 690942
rect 43268 690908 43284 690942
rect 43184 690892 43284 690908
rect 43342 690942 43442 690989
rect 43342 690908 43358 690942
rect 43426 690908 43442 690942
rect 43342 690892 43442 690908
rect 43500 690942 43600 690989
rect 43500 690908 43516 690942
rect 43584 690908 43600 690942
rect 43500 690892 43600 690908
rect 43658 690942 43758 690989
rect 43658 690908 43674 690942
rect 43742 690908 43758 690942
rect 43658 690892 43758 690908
rect 43816 690942 43916 690989
rect 43816 690908 43832 690942
rect 43900 690908 43916 690942
rect 43816 690892 43916 690908
rect 43974 690942 44074 690989
rect 43974 690908 43990 690942
rect 44058 690908 44074 690942
rect 43974 690892 44074 690908
rect 44132 690942 44232 690989
rect 44132 690908 44148 690942
rect 44216 690908 44232 690942
rect 44132 690892 44232 690908
rect 44290 690942 44390 690989
rect 44290 690908 44306 690942
rect 44374 690908 44390 690942
rect 44290 690892 44390 690908
rect 44448 690942 44548 690989
rect 44448 690908 44464 690942
rect 44532 690908 44548 690942
rect 44448 690892 44548 690908
rect 44606 690942 44706 690989
rect 44606 690908 44622 690942
rect 44690 690908 44706 690942
rect 44606 690892 44706 690908
rect 44764 690942 44864 690989
rect 44764 690908 44780 690942
rect 44848 690908 44864 690942
rect 44764 690892 44864 690908
rect 44922 690942 45022 690989
rect 44922 690908 44938 690942
rect 45006 690908 45022 690942
rect 44922 690892 45022 690908
rect 45080 690942 45180 690989
rect 45080 690908 45096 690942
rect 45164 690908 45180 690942
rect 45080 690892 45180 690908
rect 45238 690942 45338 690989
rect 45238 690908 45254 690942
rect 45322 690908 45338 690942
rect 45238 690892 45338 690908
rect 45396 690942 45496 690989
rect 45396 690908 45412 690942
rect 45480 690908 45496 690942
rect 45396 690892 45496 690908
rect 45554 690942 45654 690989
rect 45554 690908 45570 690942
rect 45638 690908 45654 690942
rect 45554 690892 45654 690908
rect 45712 690942 45812 690989
rect 45712 690908 45728 690942
rect 45796 690908 45812 690942
rect 45712 690892 45812 690908
rect 45870 690942 45970 690989
rect 45870 690908 45886 690942
rect 45954 690908 45970 690942
rect 45870 690892 45970 690908
rect 46028 690942 46128 690989
rect 46028 690908 46044 690942
rect 46112 690908 46128 690942
rect 46028 690892 46128 690908
rect 46186 690942 46286 690989
rect 46186 690908 46202 690942
rect 46270 690908 46286 690942
rect 46186 690892 46286 690908
rect 44127 690493 44227 690509
rect 44127 690459 44143 690493
rect 44211 690459 44227 690493
rect 44127 690421 44227 690459
rect 44285 690493 44385 690509
rect 44285 690459 44301 690493
rect 44369 690459 44385 690493
rect 44285 690421 44385 690459
rect 44443 690493 44543 690509
rect 44443 690459 44459 690493
rect 44527 690459 44543 690493
rect 44443 690421 44543 690459
rect 44601 690493 44701 690509
rect 44601 690459 44617 690493
rect 44685 690459 44701 690493
rect 44601 690421 44701 690459
rect 44759 690493 44859 690509
rect 44759 690459 44775 690493
rect 44843 690459 44859 690493
rect 44759 690421 44859 690459
rect 44917 690493 45017 690509
rect 44917 690459 44933 690493
rect 45001 690459 45017 690493
rect 44917 690421 45017 690459
rect 45075 690493 45175 690509
rect 45075 690459 45091 690493
rect 45159 690459 45175 690493
rect 45075 690421 45175 690459
rect 44127 689383 44227 689421
rect 44127 689349 44143 689383
rect 44211 689349 44227 689383
rect 44127 689333 44227 689349
rect 44285 689383 44385 689421
rect 44285 689349 44301 689383
rect 44369 689349 44385 689383
rect 44285 689333 44385 689349
rect 44443 689383 44543 689421
rect 44443 689349 44459 689383
rect 44527 689349 44543 689383
rect 44443 689333 44543 689349
rect 44601 689383 44701 689421
rect 44601 689349 44617 689383
rect 44685 689349 44701 689383
rect 44601 689333 44701 689349
rect 44759 689383 44859 689421
rect 44759 689349 44775 689383
rect 44843 689349 44859 689383
rect 44759 689333 44859 689349
rect 44917 689383 45017 689421
rect 44917 689349 44933 689383
rect 45001 689349 45017 689383
rect 44917 689333 45017 689349
rect 45075 689383 45175 689421
rect 45075 689349 45091 689383
rect 45159 689349 45175 689383
rect 45075 689333 45175 689349
rect 540271 690722 540368 690738
rect 540271 690654 540287 690722
rect 540321 690654 540368 690722
rect 540271 690638 540368 690654
rect 541368 690722 541465 690738
rect 541368 690654 541415 690722
rect 541449 690654 541465 690722
rect 541368 690638 541465 690654
rect 541507 690722 541604 690738
rect 541507 690654 541523 690722
rect 541557 690654 541604 690722
rect 541507 690638 541604 690654
rect 542604 690722 542701 690738
rect 542604 690654 542651 690722
rect 542685 690654 542701 690722
rect 542604 690638 542701 690654
rect 542743 690722 542840 690738
rect 542743 690654 542759 690722
rect 542793 690654 542840 690722
rect 542743 690638 542840 690654
rect 543840 690722 543937 690738
rect 543840 690654 543887 690722
rect 543921 690654 543937 690722
rect 543840 690638 543937 690654
rect 543979 690722 544076 690738
rect 543979 690654 543995 690722
rect 544029 690654 544076 690722
rect 543979 690638 544076 690654
rect 545076 690722 545173 690738
rect 545076 690654 545123 690722
rect 545157 690654 545173 690722
rect 545076 690638 545173 690654
rect 545215 690722 545312 690738
rect 545215 690654 545231 690722
rect 545265 690654 545312 690722
rect 545215 690638 545312 690654
rect 546312 690722 546409 690738
rect 546312 690654 546359 690722
rect 546393 690654 546409 690722
rect 546312 690638 546409 690654
rect 546451 690722 546548 690738
rect 546451 690654 546467 690722
rect 546501 690654 546548 690722
rect 546451 690638 546548 690654
rect 547548 690722 547645 690738
rect 547548 690654 547595 690722
rect 547629 690654 547645 690722
rect 547548 690638 547645 690654
rect 547687 690722 547784 690738
rect 547687 690654 547703 690722
rect 547737 690654 547784 690722
rect 547687 690638 547784 690654
rect 548784 690722 548881 690738
rect 548784 690654 548831 690722
rect 548865 690654 548881 690722
rect 548784 690638 548881 690654
rect 540271 690182 540368 690198
rect 540271 690114 540287 690182
rect 540321 690114 540368 690182
rect 540271 690098 540368 690114
rect 541368 690182 541465 690198
rect 541368 690114 541415 690182
rect 541449 690114 541465 690182
rect 541368 690098 541465 690114
rect 541507 690182 541604 690198
rect 541507 690114 541523 690182
rect 541557 690114 541604 690182
rect 541507 690098 541604 690114
rect 542604 690182 542701 690198
rect 542604 690114 542651 690182
rect 542685 690114 542701 690182
rect 542604 690098 542701 690114
rect 542743 690182 542840 690198
rect 542743 690114 542759 690182
rect 542793 690114 542840 690182
rect 542743 690098 542840 690114
rect 543840 690182 543937 690198
rect 543840 690114 543887 690182
rect 543921 690114 543937 690182
rect 543840 690098 543937 690114
rect 543979 690182 544076 690198
rect 543979 690114 543995 690182
rect 544029 690114 544076 690182
rect 543979 690098 544076 690114
rect 545076 690182 545173 690198
rect 545076 690114 545123 690182
rect 545157 690114 545173 690182
rect 545076 690098 545173 690114
rect 545215 690182 545312 690198
rect 545215 690114 545231 690182
rect 545265 690114 545312 690182
rect 545215 690098 545312 690114
rect 546312 690182 546409 690198
rect 546312 690114 546359 690182
rect 546393 690114 546409 690182
rect 546312 690098 546409 690114
rect 546451 690182 546548 690198
rect 546451 690114 546467 690182
rect 546501 690114 546548 690182
rect 546451 690098 546548 690114
rect 547548 690182 547645 690198
rect 547548 690114 547595 690182
rect 547629 690114 547645 690182
rect 547548 690098 547645 690114
rect 547687 690182 547784 690198
rect 547687 690114 547703 690182
rect 547737 690114 547784 690182
rect 547687 690098 547784 690114
rect 548784 690182 548881 690198
rect 548784 690114 548831 690182
rect 548865 690114 548881 690182
rect 548784 690098 548881 690114
rect 540271 689642 540368 689658
rect 540271 689574 540287 689642
rect 540321 689574 540368 689642
rect 540271 689558 540368 689574
rect 541368 689642 541465 689658
rect 541368 689574 541415 689642
rect 541449 689574 541465 689642
rect 541368 689558 541465 689574
rect 541507 689642 541604 689658
rect 541507 689574 541523 689642
rect 541557 689574 541604 689642
rect 541507 689558 541604 689574
rect 542604 689642 542701 689658
rect 542604 689574 542651 689642
rect 542685 689574 542701 689642
rect 542604 689558 542701 689574
rect 542743 689642 542840 689658
rect 542743 689574 542759 689642
rect 542793 689574 542840 689642
rect 542743 689558 542840 689574
rect 543840 689642 543937 689658
rect 543840 689574 543887 689642
rect 543921 689574 543937 689642
rect 543840 689558 543937 689574
rect 543979 689642 544076 689658
rect 543979 689574 543995 689642
rect 544029 689574 544076 689642
rect 543979 689558 544076 689574
rect 545076 689642 545173 689658
rect 545076 689574 545123 689642
rect 545157 689574 545173 689642
rect 545076 689558 545173 689574
rect 545215 689642 545312 689658
rect 545215 689574 545231 689642
rect 545265 689574 545312 689642
rect 545215 689558 545312 689574
rect 546312 689642 546409 689658
rect 546312 689574 546359 689642
rect 546393 689574 546409 689642
rect 546312 689558 546409 689574
rect 546451 689642 546548 689658
rect 546451 689574 546467 689642
rect 546501 689574 546548 689642
rect 546451 689558 546548 689574
rect 547548 689642 547645 689658
rect 547548 689574 547595 689642
rect 547629 689574 547645 689642
rect 547548 689558 547645 689574
rect 547687 689642 547784 689658
rect 547687 689574 547703 689642
rect 547737 689574 547784 689642
rect 547687 689558 547784 689574
rect 548784 689642 548881 689658
rect 548784 689574 548831 689642
rect 548865 689574 548881 689642
rect 548784 689558 548881 689574
rect 44127 688973 44227 688989
rect 44127 688939 44143 688973
rect 44211 688939 44227 688973
rect 44127 688901 44227 688939
rect 44285 688973 44385 688989
rect 44285 688939 44301 688973
rect 44369 688939 44385 688973
rect 44285 688901 44385 688939
rect 44443 688973 44543 688989
rect 44443 688939 44459 688973
rect 44527 688939 44543 688973
rect 44443 688901 44543 688939
rect 44601 688973 44701 688989
rect 44601 688939 44617 688973
rect 44685 688939 44701 688973
rect 44601 688901 44701 688939
rect 44759 688973 44859 688989
rect 44759 688939 44775 688973
rect 44843 688939 44859 688973
rect 44759 688901 44859 688939
rect 44917 688973 45017 688989
rect 44917 688939 44933 688973
rect 45001 688939 45017 688973
rect 44917 688901 45017 688939
rect 45075 688973 45175 688989
rect 45075 688939 45091 688973
rect 45159 688939 45175 688973
rect 45075 688901 45175 688939
rect 44127 687863 44227 687901
rect 44127 687829 44143 687863
rect 44211 687829 44227 687863
rect 44127 687813 44227 687829
rect 44285 687863 44385 687901
rect 44285 687829 44301 687863
rect 44369 687829 44385 687863
rect 44285 687813 44385 687829
rect 44443 687863 44543 687901
rect 44443 687829 44459 687863
rect 44527 687829 44543 687863
rect 44443 687813 44543 687829
rect 44601 687863 44701 687901
rect 44601 687829 44617 687863
rect 44685 687829 44701 687863
rect 44601 687813 44701 687829
rect 44759 687863 44859 687901
rect 44759 687829 44775 687863
rect 44843 687829 44859 687863
rect 44759 687813 44859 687829
rect 44917 687863 45017 687901
rect 44917 687829 44933 687863
rect 45001 687829 45017 687863
rect 44917 687813 45017 687829
rect 45075 687863 45175 687901
rect 45075 687829 45091 687863
rect 45159 687829 45175 687863
rect 45075 687813 45175 687829
rect 540271 689102 540368 689118
rect 540271 689034 540287 689102
rect 540321 689034 540368 689102
rect 540271 689018 540368 689034
rect 541368 689102 541465 689118
rect 541368 689034 541415 689102
rect 541449 689034 541465 689102
rect 541368 689018 541465 689034
rect 541507 689102 541604 689118
rect 541507 689034 541523 689102
rect 541557 689034 541604 689102
rect 541507 689018 541604 689034
rect 542604 689102 542701 689118
rect 542604 689034 542651 689102
rect 542685 689034 542701 689102
rect 542604 689018 542701 689034
rect 542743 689102 542840 689118
rect 542743 689034 542759 689102
rect 542793 689034 542840 689102
rect 542743 689018 542840 689034
rect 543840 689102 543937 689118
rect 543840 689034 543887 689102
rect 543921 689034 543937 689102
rect 543840 689018 543937 689034
rect 543979 689102 544076 689118
rect 543979 689034 543995 689102
rect 544029 689034 544076 689102
rect 543979 689018 544076 689034
rect 545076 689102 545173 689118
rect 545076 689034 545123 689102
rect 545157 689034 545173 689102
rect 545076 689018 545173 689034
rect 545215 689102 545312 689118
rect 545215 689034 545231 689102
rect 545265 689034 545312 689102
rect 545215 689018 545312 689034
rect 546312 689102 546409 689118
rect 546312 689034 546359 689102
rect 546393 689034 546409 689102
rect 546312 689018 546409 689034
rect 546451 689102 546548 689118
rect 546451 689034 546467 689102
rect 546501 689034 546548 689102
rect 546451 689018 546548 689034
rect 547548 689102 547645 689118
rect 547548 689034 547595 689102
rect 547629 689034 547645 689102
rect 547548 689018 547645 689034
rect 547687 689102 547784 689118
rect 547687 689034 547703 689102
rect 547737 689034 547784 689102
rect 547687 689018 547784 689034
rect 548784 689102 548881 689118
rect 548784 689034 548831 689102
rect 548865 689034 548881 689102
rect 548784 689018 548881 689034
rect 540271 688522 540368 688538
rect 540271 688454 540287 688522
rect 540321 688454 540368 688522
rect 540271 688438 540368 688454
rect 541368 688522 541465 688538
rect 541368 688454 541415 688522
rect 541449 688454 541465 688522
rect 541368 688438 541465 688454
rect 541507 688522 541604 688538
rect 541507 688454 541523 688522
rect 541557 688454 541604 688522
rect 541507 688438 541604 688454
rect 542604 688522 542701 688538
rect 542604 688454 542651 688522
rect 542685 688454 542701 688522
rect 542604 688438 542701 688454
rect 542743 688522 542840 688538
rect 542743 688454 542759 688522
rect 542793 688454 542840 688522
rect 542743 688438 542840 688454
rect 543840 688522 543937 688538
rect 543840 688454 543887 688522
rect 543921 688454 543937 688522
rect 543840 688438 543937 688454
rect 543979 688522 544076 688538
rect 543979 688454 543995 688522
rect 544029 688454 544076 688522
rect 543979 688438 544076 688454
rect 545076 688522 545173 688538
rect 545076 688454 545123 688522
rect 545157 688454 545173 688522
rect 545076 688438 545173 688454
rect 545215 688522 545312 688538
rect 545215 688454 545231 688522
rect 545265 688454 545312 688522
rect 545215 688438 545312 688454
rect 546312 688522 546409 688538
rect 546312 688454 546359 688522
rect 546393 688454 546409 688522
rect 546312 688438 546409 688454
rect 546451 688522 546548 688538
rect 546451 688454 546467 688522
rect 546501 688454 546548 688522
rect 546451 688438 546548 688454
rect 547548 688522 547645 688538
rect 547548 688454 547595 688522
rect 547629 688454 547645 688522
rect 547548 688438 547645 688454
rect 547687 688522 547784 688538
rect 547687 688454 547703 688522
rect 547737 688454 547784 688522
rect 547687 688438 547784 688454
rect 548784 688522 548881 688538
rect 548784 688454 548831 688522
rect 548865 688454 548881 688522
rect 548784 688438 548881 688454
rect 43136 687452 43336 687468
rect 43136 687418 43152 687452
rect 43320 687418 43336 687452
rect 43136 687380 43336 687418
rect 43394 687452 43594 687468
rect 43394 687418 43410 687452
rect 43578 687418 43594 687452
rect 43394 687380 43594 687418
rect 43652 687452 43852 687468
rect 43652 687418 43668 687452
rect 43836 687418 43852 687452
rect 43652 687380 43852 687418
rect 43910 687452 44110 687468
rect 43910 687418 43926 687452
rect 44094 687418 44110 687452
rect 43910 687380 44110 687418
rect 44168 687452 44368 687468
rect 44168 687418 44184 687452
rect 44352 687418 44368 687452
rect 44168 687380 44368 687418
rect 44426 687452 44626 687468
rect 44426 687418 44442 687452
rect 44610 687418 44626 687452
rect 44426 687380 44626 687418
rect 44684 687452 44884 687468
rect 44684 687418 44700 687452
rect 44868 687418 44884 687452
rect 44684 687380 44884 687418
rect 44942 687452 45142 687468
rect 44942 687418 44958 687452
rect 45126 687418 45142 687452
rect 44942 687380 45142 687418
rect 45200 687452 45400 687468
rect 45200 687418 45216 687452
rect 45384 687418 45400 687452
rect 45200 687380 45400 687418
rect 45458 687452 45658 687468
rect 45458 687418 45474 687452
rect 45642 687418 45658 687452
rect 45458 687380 45658 687418
rect 45716 687452 45916 687468
rect 45716 687418 45732 687452
rect 45900 687418 45916 687452
rect 45716 687380 45916 687418
rect 45974 687452 46174 687468
rect 45974 687418 45990 687452
rect 46158 687418 46174 687452
rect 45974 687380 46174 687418
rect 43136 686342 43336 686380
rect 43136 686308 43152 686342
rect 43320 686308 43336 686342
rect 43136 686292 43336 686308
rect 43394 686342 43594 686380
rect 43394 686308 43410 686342
rect 43578 686308 43594 686342
rect 43394 686292 43594 686308
rect 43652 686342 43852 686380
rect 43652 686308 43668 686342
rect 43836 686308 43852 686342
rect 43652 686292 43852 686308
rect 43910 686342 44110 686380
rect 43910 686308 43926 686342
rect 44094 686308 44110 686342
rect 43910 686292 44110 686308
rect 44168 686342 44368 686380
rect 44168 686308 44184 686342
rect 44352 686308 44368 686342
rect 44168 686292 44368 686308
rect 44426 686342 44626 686380
rect 44426 686308 44442 686342
rect 44610 686308 44626 686342
rect 44426 686292 44626 686308
rect 44684 686342 44884 686380
rect 44684 686308 44700 686342
rect 44868 686308 44884 686342
rect 44684 686292 44884 686308
rect 44942 686342 45142 686380
rect 44942 686308 44958 686342
rect 45126 686308 45142 686342
rect 44942 686292 45142 686308
rect 45200 686342 45400 686380
rect 45200 686308 45216 686342
rect 45384 686308 45400 686342
rect 45200 686292 45400 686308
rect 45458 686342 45658 686380
rect 45458 686308 45474 686342
rect 45642 686308 45658 686342
rect 45458 686292 45658 686308
rect 45716 686342 45916 686380
rect 45716 686308 45732 686342
rect 45900 686308 45916 686342
rect 45716 686292 45916 686308
rect 45974 686342 46174 686380
rect 45974 686308 45990 686342
rect 46158 686308 46174 686342
rect 45974 686292 46174 686308
rect 540271 687942 540368 687958
rect 540271 687874 540287 687942
rect 540321 687874 540368 687942
rect 540271 687858 540368 687874
rect 541368 687942 541465 687958
rect 541368 687874 541415 687942
rect 541449 687874 541465 687942
rect 541368 687858 541465 687874
rect 541507 687942 541604 687958
rect 541507 687874 541523 687942
rect 541557 687874 541604 687942
rect 541507 687858 541604 687874
rect 542604 687942 542701 687958
rect 542604 687874 542651 687942
rect 542685 687874 542701 687942
rect 542604 687858 542701 687874
rect 542743 687942 542840 687958
rect 542743 687874 542759 687942
rect 542793 687874 542840 687942
rect 542743 687858 542840 687874
rect 543840 687942 543937 687958
rect 543840 687874 543887 687942
rect 543921 687874 543937 687942
rect 543840 687858 543937 687874
rect 543979 687942 544076 687958
rect 543979 687874 543995 687942
rect 544029 687874 544076 687942
rect 543979 687858 544076 687874
rect 545076 687942 545173 687958
rect 545076 687874 545123 687942
rect 545157 687874 545173 687942
rect 545076 687858 545173 687874
rect 545215 687942 545312 687958
rect 545215 687874 545231 687942
rect 545265 687874 545312 687942
rect 545215 687858 545312 687874
rect 546312 687942 546409 687958
rect 546312 687874 546359 687942
rect 546393 687874 546409 687942
rect 546312 687858 546409 687874
rect 546451 687942 546548 687958
rect 546451 687874 546467 687942
rect 546501 687874 546548 687942
rect 546451 687858 546548 687874
rect 547548 687942 547645 687958
rect 547548 687874 547595 687942
rect 547629 687874 547645 687942
rect 547548 687858 547645 687874
rect 547687 687942 547784 687958
rect 547687 687874 547703 687942
rect 547737 687874 547784 687942
rect 547687 687858 547784 687874
rect 548784 687942 548881 687958
rect 548784 687874 548831 687942
rect 548865 687874 548881 687942
rect 548784 687858 548881 687874
rect 538431 687402 538528 687418
rect 538431 687334 538447 687402
rect 538481 687334 538528 687402
rect 538431 687318 538528 687334
rect 539528 687402 539625 687418
rect 539528 687334 539575 687402
rect 539609 687334 539625 687402
rect 539528 687318 539625 687334
rect 539667 687402 539764 687418
rect 539667 687334 539683 687402
rect 539717 687334 539764 687402
rect 539667 687318 539764 687334
rect 540764 687402 540861 687418
rect 540764 687334 540811 687402
rect 540845 687334 540861 687402
rect 540764 687318 540861 687334
rect 540903 687402 541000 687418
rect 540903 687334 540919 687402
rect 540953 687334 541000 687402
rect 540903 687318 541000 687334
rect 542000 687402 542097 687418
rect 542000 687334 542047 687402
rect 542081 687334 542097 687402
rect 542000 687318 542097 687334
rect 542139 687402 542236 687418
rect 542139 687334 542155 687402
rect 542189 687334 542236 687402
rect 542139 687318 542236 687334
rect 543236 687402 543333 687418
rect 543236 687334 543283 687402
rect 543317 687334 543333 687402
rect 543236 687318 543333 687334
rect 543375 687402 543472 687418
rect 543375 687334 543391 687402
rect 543425 687334 543472 687402
rect 543375 687318 543472 687334
rect 544472 687402 544569 687418
rect 544472 687334 544519 687402
rect 544553 687334 544569 687402
rect 544472 687318 544569 687334
rect 544611 687402 544708 687418
rect 544611 687334 544627 687402
rect 544661 687334 544708 687402
rect 544611 687318 544708 687334
rect 545708 687402 545805 687418
rect 545708 687334 545755 687402
rect 545789 687334 545805 687402
rect 545708 687318 545805 687334
rect 545847 687402 545944 687418
rect 545847 687334 545863 687402
rect 545897 687334 545944 687402
rect 545847 687318 545944 687334
rect 546944 687402 547041 687418
rect 546944 687334 546991 687402
rect 547025 687334 547041 687402
rect 546944 687318 547041 687334
rect 547083 687402 547180 687418
rect 547083 687334 547099 687402
rect 547133 687334 547180 687402
rect 547083 687318 547180 687334
rect 548180 687402 548277 687418
rect 548180 687334 548227 687402
rect 548261 687334 548277 687402
rect 548180 687318 548277 687334
rect 548319 687402 548416 687418
rect 548319 687334 548335 687402
rect 548369 687334 548416 687402
rect 548319 687318 548416 687334
rect 549416 687402 549513 687418
rect 549416 687334 549463 687402
rect 549497 687334 549513 687402
rect 549416 687318 549513 687334
rect 549555 687402 549652 687418
rect 549555 687334 549571 687402
rect 549605 687334 549652 687402
rect 549555 687318 549652 687334
rect 550652 687402 550749 687418
rect 550652 687334 550699 687402
rect 550733 687334 550749 687402
rect 550652 687318 550749 687334
rect 538431 686862 538528 686878
rect 538431 686794 538447 686862
rect 538481 686794 538528 686862
rect 538431 686778 538528 686794
rect 539528 686862 539625 686878
rect 539528 686794 539575 686862
rect 539609 686794 539625 686862
rect 539528 686778 539625 686794
rect 539667 686862 539764 686878
rect 539667 686794 539683 686862
rect 539717 686794 539764 686862
rect 539667 686778 539764 686794
rect 540764 686862 540861 686878
rect 540764 686794 540811 686862
rect 540845 686794 540861 686862
rect 540764 686778 540861 686794
rect 540903 686862 541000 686878
rect 540903 686794 540919 686862
rect 540953 686794 541000 686862
rect 540903 686778 541000 686794
rect 542000 686862 542097 686878
rect 542000 686794 542047 686862
rect 542081 686794 542097 686862
rect 542000 686778 542097 686794
rect 542139 686862 542236 686878
rect 542139 686794 542155 686862
rect 542189 686794 542236 686862
rect 542139 686778 542236 686794
rect 543236 686862 543333 686878
rect 543236 686794 543283 686862
rect 543317 686794 543333 686862
rect 543236 686778 543333 686794
rect 543375 686862 543472 686878
rect 543375 686794 543391 686862
rect 543425 686794 543472 686862
rect 543375 686778 543472 686794
rect 544472 686862 544569 686878
rect 544472 686794 544519 686862
rect 544553 686794 544569 686862
rect 544472 686778 544569 686794
rect 544611 686862 544708 686878
rect 544611 686794 544627 686862
rect 544661 686794 544708 686862
rect 544611 686778 544708 686794
rect 545708 686862 545805 686878
rect 545708 686794 545755 686862
rect 545789 686794 545805 686862
rect 545708 686778 545805 686794
rect 545847 686862 545944 686878
rect 545847 686794 545863 686862
rect 545897 686794 545944 686862
rect 545847 686778 545944 686794
rect 546944 686862 547041 686878
rect 546944 686794 546991 686862
rect 547025 686794 547041 686862
rect 546944 686778 547041 686794
rect 547083 686862 547180 686878
rect 547083 686794 547099 686862
rect 547133 686794 547180 686862
rect 547083 686778 547180 686794
rect 548180 686862 548277 686878
rect 548180 686794 548227 686862
rect 548261 686794 548277 686862
rect 548180 686778 548277 686794
rect 548319 686862 548416 686878
rect 548319 686794 548335 686862
rect 548369 686794 548416 686862
rect 548319 686778 548416 686794
rect 549416 686862 549513 686878
rect 549416 686794 549463 686862
rect 549497 686794 549513 686862
rect 549416 686778 549513 686794
rect 549555 686862 549652 686878
rect 549555 686794 549571 686862
rect 549605 686794 549652 686862
rect 549555 686778 549652 686794
rect 550652 686862 550749 686878
rect 550652 686794 550699 686862
rect 550733 686794 550749 686862
rect 550652 686778 550749 686794
rect 42876 685932 43076 685948
rect 42876 685898 42892 685932
rect 43060 685898 43076 685932
rect 42876 685860 43076 685898
rect 43134 685932 43334 685948
rect 43134 685898 43150 685932
rect 43318 685898 43334 685932
rect 43134 685860 43334 685898
rect 43392 685932 43592 685948
rect 43392 685898 43408 685932
rect 43576 685898 43592 685932
rect 43392 685860 43592 685898
rect 43650 685932 43850 685948
rect 43650 685898 43666 685932
rect 43834 685898 43850 685932
rect 43650 685860 43850 685898
rect 43908 685932 44108 685948
rect 43908 685898 43924 685932
rect 44092 685898 44108 685932
rect 43908 685860 44108 685898
rect 44166 685932 44366 685948
rect 44166 685898 44182 685932
rect 44350 685898 44366 685932
rect 44166 685860 44366 685898
rect 44424 685932 44624 685948
rect 44424 685898 44440 685932
rect 44608 685898 44624 685932
rect 44424 685860 44624 685898
rect 44682 685932 44882 685948
rect 44682 685898 44698 685932
rect 44866 685898 44882 685932
rect 44682 685860 44882 685898
rect 44940 685932 45140 685948
rect 44940 685898 44956 685932
rect 45124 685898 45140 685932
rect 44940 685860 45140 685898
rect 45198 685932 45398 685948
rect 45198 685898 45214 685932
rect 45382 685898 45398 685932
rect 45198 685860 45398 685898
rect 45456 685932 45656 685948
rect 45456 685898 45472 685932
rect 45640 685898 45656 685932
rect 45456 685860 45656 685898
rect 45714 685932 45914 685948
rect 45714 685898 45730 685932
rect 45898 685898 45914 685932
rect 45714 685860 45914 685898
rect 45972 685932 46172 685948
rect 45972 685898 45988 685932
rect 46156 685898 46172 685932
rect 45972 685860 46172 685898
rect 46230 685932 46430 685948
rect 46230 685898 46246 685932
rect 46414 685898 46430 685932
rect 46230 685860 46430 685898
rect 42876 684822 43076 684860
rect 42876 684788 42892 684822
rect 43060 684788 43076 684822
rect 42876 684772 43076 684788
rect 43134 684822 43334 684860
rect 43134 684788 43150 684822
rect 43318 684788 43334 684822
rect 43134 684772 43334 684788
rect 43392 684822 43592 684860
rect 43392 684788 43408 684822
rect 43576 684788 43592 684822
rect 43392 684772 43592 684788
rect 43650 684822 43850 684860
rect 43650 684788 43666 684822
rect 43834 684788 43850 684822
rect 43650 684772 43850 684788
rect 43908 684822 44108 684860
rect 43908 684788 43924 684822
rect 44092 684788 44108 684822
rect 43908 684772 44108 684788
rect 44166 684822 44366 684860
rect 44166 684788 44182 684822
rect 44350 684788 44366 684822
rect 44166 684772 44366 684788
rect 44424 684822 44624 684860
rect 44424 684788 44440 684822
rect 44608 684788 44624 684822
rect 44424 684772 44624 684788
rect 44682 684822 44882 684860
rect 44682 684788 44698 684822
rect 44866 684788 44882 684822
rect 44682 684772 44882 684788
rect 44940 684822 45140 684860
rect 44940 684788 44956 684822
rect 45124 684788 45140 684822
rect 44940 684772 45140 684788
rect 45198 684822 45398 684860
rect 45198 684788 45214 684822
rect 45382 684788 45398 684822
rect 45198 684772 45398 684788
rect 45456 684822 45656 684860
rect 45456 684788 45472 684822
rect 45640 684788 45656 684822
rect 45456 684772 45656 684788
rect 45714 684822 45914 684860
rect 45714 684788 45730 684822
rect 45898 684788 45914 684822
rect 45714 684772 45914 684788
rect 45972 684822 46172 684860
rect 45972 684788 45988 684822
rect 46156 684788 46172 684822
rect 45972 684772 46172 684788
rect 46230 684822 46430 684860
rect 46230 684788 46246 684822
rect 46414 684788 46430 684822
rect 46230 684772 46430 684788
rect 538431 686322 538528 686338
rect 538431 686254 538447 686322
rect 538481 686254 538528 686322
rect 538431 686238 538528 686254
rect 539528 686322 539625 686338
rect 539528 686254 539575 686322
rect 539609 686254 539625 686322
rect 539528 686238 539625 686254
rect 539667 686322 539764 686338
rect 539667 686254 539683 686322
rect 539717 686254 539764 686322
rect 539667 686238 539764 686254
rect 540764 686322 540861 686338
rect 540764 686254 540811 686322
rect 540845 686254 540861 686322
rect 540764 686238 540861 686254
rect 540903 686322 541000 686338
rect 540903 686254 540919 686322
rect 540953 686254 541000 686322
rect 540903 686238 541000 686254
rect 542000 686322 542097 686338
rect 542000 686254 542047 686322
rect 542081 686254 542097 686322
rect 542000 686238 542097 686254
rect 542139 686322 542236 686338
rect 542139 686254 542155 686322
rect 542189 686254 542236 686322
rect 542139 686238 542236 686254
rect 543236 686322 543333 686338
rect 543236 686254 543283 686322
rect 543317 686254 543333 686322
rect 543236 686238 543333 686254
rect 543375 686322 543472 686338
rect 543375 686254 543391 686322
rect 543425 686254 543472 686322
rect 543375 686238 543472 686254
rect 544472 686322 544569 686338
rect 544472 686254 544519 686322
rect 544553 686254 544569 686322
rect 544472 686238 544569 686254
rect 544611 686322 544708 686338
rect 544611 686254 544627 686322
rect 544661 686254 544708 686322
rect 544611 686238 544708 686254
rect 545708 686322 545805 686338
rect 545708 686254 545755 686322
rect 545789 686254 545805 686322
rect 545708 686238 545805 686254
rect 545847 686322 545944 686338
rect 545847 686254 545863 686322
rect 545897 686254 545944 686322
rect 545847 686238 545944 686254
rect 546944 686322 547041 686338
rect 546944 686254 546991 686322
rect 547025 686254 547041 686322
rect 546944 686238 547041 686254
rect 547083 686322 547180 686338
rect 547083 686254 547099 686322
rect 547133 686254 547180 686322
rect 547083 686238 547180 686254
rect 548180 686322 548277 686338
rect 548180 686254 548227 686322
rect 548261 686254 548277 686322
rect 548180 686238 548277 686254
rect 548319 686322 548416 686338
rect 548319 686254 548335 686322
rect 548369 686254 548416 686322
rect 548319 686238 548416 686254
rect 549416 686322 549513 686338
rect 549416 686254 549463 686322
rect 549497 686254 549513 686322
rect 549416 686238 549513 686254
rect 549555 686322 549652 686338
rect 549555 686254 549571 686322
rect 549605 686254 549652 686322
rect 549555 686238 549652 686254
rect 550652 686322 550749 686338
rect 550652 686254 550699 686322
rect 550733 686254 550749 686322
rect 550652 686238 550749 686254
rect 538431 685782 538528 685798
rect 538431 685714 538447 685782
rect 538481 685714 538528 685782
rect 538431 685698 538528 685714
rect 539528 685782 539625 685798
rect 539528 685714 539575 685782
rect 539609 685714 539625 685782
rect 539528 685698 539625 685714
rect 539667 685782 539764 685798
rect 539667 685714 539683 685782
rect 539717 685714 539764 685782
rect 539667 685698 539764 685714
rect 540764 685782 540861 685798
rect 540764 685714 540811 685782
rect 540845 685714 540861 685782
rect 540764 685698 540861 685714
rect 540903 685782 541000 685798
rect 540903 685714 540919 685782
rect 540953 685714 541000 685782
rect 540903 685698 541000 685714
rect 542000 685782 542097 685798
rect 542000 685714 542047 685782
rect 542081 685714 542097 685782
rect 542000 685698 542097 685714
rect 542139 685782 542236 685798
rect 542139 685714 542155 685782
rect 542189 685714 542236 685782
rect 542139 685698 542236 685714
rect 543236 685782 543333 685798
rect 543236 685714 543283 685782
rect 543317 685714 543333 685782
rect 543236 685698 543333 685714
rect 543375 685782 543472 685798
rect 543375 685714 543391 685782
rect 543425 685714 543472 685782
rect 543375 685698 543472 685714
rect 544472 685782 544569 685798
rect 544472 685714 544519 685782
rect 544553 685714 544569 685782
rect 544472 685698 544569 685714
rect 544611 685782 544708 685798
rect 544611 685714 544627 685782
rect 544661 685714 544708 685782
rect 544611 685698 544708 685714
rect 545708 685782 545805 685798
rect 545708 685714 545755 685782
rect 545789 685714 545805 685782
rect 545708 685698 545805 685714
rect 545847 685782 545944 685798
rect 545847 685714 545863 685782
rect 545897 685714 545944 685782
rect 545847 685698 545944 685714
rect 546944 685782 547041 685798
rect 546944 685714 546991 685782
rect 547025 685714 547041 685782
rect 546944 685698 547041 685714
rect 547083 685782 547180 685798
rect 547083 685714 547099 685782
rect 547133 685714 547180 685782
rect 547083 685698 547180 685714
rect 548180 685782 548277 685798
rect 548180 685714 548227 685782
rect 548261 685714 548277 685782
rect 548180 685698 548277 685714
rect 548319 685782 548416 685798
rect 548319 685714 548335 685782
rect 548369 685714 548416 685782
rect 548319 685698 548416 685714
rect 549416 685782 549513 685798
rect 549416 685714 549463 685782
rect 549497 685714 549513 685782
rect 549416 685698 549513 685714
rect 549555 685782 549652 685798
rect 549555 685714 549571 685782
rect 549605 685714 549652 685782
rect 549555 685698 549652 685714
rect 550652 685782 550749 685798
rect 550652 685714 550699 685782
rect 550733 685714 550749 685782
rect 550652 685698 550749 685714
rect 540371 685002 540459 685018
rect 540371 684934 540387 685002
rect 540421 684934 540459 685002
rect 540371 684918 540459 684934
rect 541459 685002 541547 685018
rect 541459 684934 541497 685002
rect 541531 684934 541547 685002
rect 541459 684918 541547 684934
rect 541589 685002 541677 685018
rect 541589 684934 541605 685002
rect 541639 684934 541677 685002
rect 541589 684918 541677 684934
rect 542677 685002 542765 685018
rect 542677 684934 542715 685002
rect 542749 684934 542765 685002
rect 542677 684918 542765 684934
rect 542807 685002 542895 685018
rect 542807 684934 542823 685002
rect 542857 684934 542895 685002
rect 542807 684918 542895 684934
rect 543895 685002 543983 685018
rect 543895 684934 543933 685002
rect 543967 684934 543983 685002
rect 543895 684918 543983 684934
rect 544025 685002 544113 685018
rect 544025 684934 544041 685002
rect 544075 684934 544113 685002
rect 544025 684918 544113 684934
rect 545113 685002 545201 685018
rect 545113 684934 545151 685002
rect 545185 684934 545201 685002
rect 545113 684918 545201 684934
rect 545243 685002 545331 685018
rect 545243 684934 545259 685002
rect 545293 684934 545331 685002
rect 545243 684918 545331 684934
rect 546331 685002 546419 685018
rect 546331 684934 546369 685002
rect 546403 684934 546419 685002
rect 546331 684918 546419 684934
rect 546461 685002 546549 685018
rect 546461 684934 546477 685002
rect 546511 684934 546549 685002
rect 546461 684918 546549 684934
rect 547549 685002 547637 685018
rect 547549 684934 547587 685002
rect 547621 684934 547637 685002
rect 547549 684918 547637 684934
rect 547679 685002 547767 685018
rect 547679 684934 547695 685002
rect 547729 684934 547767 685002
rect 547679 684918 547767 684934
rect 548767 685002 548855 685018
rect 548767 684934 548805 685002
rect 548839 684934 548855 685002
rect 548767 684918 548855 684934
rect 540371 684502 540459 684518
rect 540371 684434 540387 684502
rect 540421 684434 540459 684502
rect 540371 684418 540459 684434
rect 541459 684502 541547 684518
rect 541459 684434 541497 684502
rect 541531 684434 541547 684502
rect 541459 684418 541547 684434
rect 541589 684502 541677 684518
rect 541589 684434 541605 684502
rect 541639 684434 541677 684502
rect 541589 684418 541677 684434
rect 542677 684502 542765 684518
rect 542677 684434 542715 684502
rect 542749 684434 542765 684502
rect 542677 684418 542765 684434
rect 542807 684502 542895 684518
rect 542807 684434 542823 684502
rect 542857 684434 542895 684502
rect 542807 684418 542895 684434
rect 543895 684502 543983 684518
rect 543895 684434 543933 684502
rect 543967 684434 543983 684502
rect 543895 684418 543983 684434
rect 544025 684502 544113 684518
rect 544025 684434 544041 684502
rect 544075 684434 544113 684502
rect 544025 684418 544113 684434
rect 545113 684502 545201 684518
rect 545113 684434 545151 684502
rect 545185 684434 545201 684502
rect 545113 684418 545201 684434
rect 545243 684502 545331 684518
rect 545243 684434 545259 684502
rect 545293 684434 545331 684502
rect 545243 684418 545331 684434
rect 546331 684502 546419 684518
rect 546331 684434 546369 684502
rect 546403 684434 546419 684502
rect 546331 684418 546419 684434
rect 546461 684502 546549 684518
rect 546461 684434 546477 684502
rect 546511 684434 546549 684502
rect 546461 684418 546549 684434
rect 547549 684502 547637 684518
rect 547549 684434 547587 684502
rect 547621 684434 547637 684502
rect 547549 684418 547637 684434
rect 547679 684502 547767 684518
rect 547679 684434 547695 684502
rect 547729 684434 547767 684502
rect 547679 684418 547767 684434
rect 548767 684502 548855 684518
rect 548767 684434 548805 684502
rect 548839 684434 548855 684502
rect 548767 684418 548855 684434
rect 43906 683900 44106 683916
rect 43906 683866 43922 683900
rect 44090 683866 44106 683900
rect 43906 683819 44106 683866
rect 44164 683900 44364 683916
rect 44164 683866 44180 683900
rect 44348 683866 44364 683900
rect 44164 683819 44364 683866
rect 44422 683900 44622 683916
rect 44422 683866 44438 683900
rect 44606 683866 44622 683900
rect 44422 683819 44622 683866
rect 44680 683900 44880 683916
rect 44680 683866 44696 683900
rect 44864 683866 44880 683900
rect 44680 683819 44880 683866
rect 44938 683900 45138 683916
rect 44938 683866 44954 683900
rect 45122 683866 45138 683900
rect 44938 683819 45138 683866
rect 45196 683900 45396 683916
rect 45196 683866 45212 683900
rect 45380 683866 45396 683900
rect 45196 683819 45396 683866
rect 43906 682772 44106 682819
rect 43906 682738 43922 682772
rect 44090 682738 44106 682772
rect 43906 682722 44106 682738
rect 44164 682772 44364 682819
rect 44164 682738 44180 682772
rect 44348 682738 44364 682772
rect 44164 682722 44364 682738
rect 44422 682772 44622 682819
rect 44422 682738 44438 682772
rect 44606 682738 44622 682772
rect 44422 682722 44622 682738
rect 44680 682772 44880 682819
rect 44680 682738 44696 682772
rect 44864 682738 44880 682772
rect 44680 682722 44880 682738
rect 44938 682772 45138 682819
rect 44938 682738 44954 682772
rect 45122 682738 45138 682772
rect 44938 682722 45138 682738
rect 45196 682772 45396 682819
rect 45196 682738 45212 682772
rect 45380 682738 45396 682772
rect 45196 682722 45396 682738
rect 540931 684002 541019 684018
rect 540931 683834 540947 684002
rect 540981 683834 541019 684002
rect 540931 683818 541019 683834
rect 542019 684002 542107 684018
rect 542019 683834 542057 684002
rect 542091 683834 542107 684002
rect 542019 683818 542107 683834
rect 542149 684002 542237 684018
rect 542149 683834 542165 684002
rect 542199 683834 542237 684002
rect 542149 683818 542237 683834
rect 543237 684002 543325 684018
rect 543237 683834 543275 684002
rect 543309 683834 543325 684002
rect 543237 683818 543325 683834
rect 543367 684002 543455 684018
rect 543367 683834 543383 684002
rect 543417 683834 543455 684002
rect 543367 683818 543455 683834
rect 544455 684002 544543 684018
rect 544455 683834 544493 684002
rect 544527 683834 544543 684002
rect 544455 683818 544543 683834
rect 544585 684002 544673 684018
rect 544585 683834 544601 684002
rect 544635 683834 544673 684002
rect 544585 683818 544673 683834
rect 545673 684002 545761 684018
rect 545673 683834 545711 684002
rect 545745 683834 545761 684002
rect 545673 683818 545761 683834
rect 545803 684002 545891 684018
rect 545803 683834 545819 684002
rect 545853 683834 545891 684002
rect 545803 683818 545891 683834
rect 546891 684002 546979 684018
rect 546891 683834 546929 684002
rect 546963 683834 546979 684002
rect 546891 683818 546979 683834
rect 547021 684002 547109 684018
rect 547021 683834 547037 684002
rect 547071 683834 547109 684002
rect 547021 683818 547109 683834
rect 548109 684002 548197 684018
rect 548109 683834 548147 684002
rect 548181 683834 548197 684002
rect 548109 683818 548197 683834
rect 540931 683382 541019 683398
rect 540931 683214 540947 683382
rect 540981 683214 541019 683382
rect 540931 683198 541019 683214
rect 542019 683382 542107 683398
rect 542019 683214 542057 683382
rect 542091 683214 542107 683382
rect 542019 683198 542107 683214
rect 542149 683382 542237 683398
rect 542149 683214 542165 683382
rect 542199 683214 542237 683382
rect 542149 683198 542237 683214
rect 543237 683382 543325 683398
rect 543237 683214 543275 683382
rect 543309 683214 543325 683382
rect 543237 683198 543325 683214
rect 543367 683382 543455 683398
rect 543367 683214 543383 683382
rect 543417 683214 543455 683382
rect 543367 683198 543455 683214
rect 544455 683382 544543 683398
rect 544455 683214 544493 683382
rect 544527 683214 544543 683382
rect 544455 683198 544543 683214
rect 544585 683382 544673 683398
rect 544585 683214 544601 683382
rect 544635 683214 544673 683382
rect 544585 683198 544673 683214
rect 545673 683382 545761 683398
rect 545673 683214 545711 683382
rect 545745 683214 545761 683382
rect 545673 683198 545761 683214
rect 545803 683382 545891 683398
rect 545803 683214 545819 683382
rect 545853 683214 545891 683382
rect 545803 683198 545891 683214
rect 546891 683382 546979 683398
rect 546891 683214 546929 683382
rect 546963 683214 546979 683382
rect 546891 683198 546979 683214
rect 547021 683382 547109 683398
rect 547021 683214 547037 683382
rect 547071 683214 547109 683382
rect 547021 683198 547109 683214
rect 548109 683382 548197 683398
rect 548109 683214 548147 683382
rect 548181 683214 548197 683382
rect 548109 683198 548197 683214
rect 540371 682782 540459 682798
rect 540371 682614 540387 682782
rect 540421 682614 540459 682782
rect 540371 682598 540459 682614
rect 541459 682782 541547 682798
rect 541459 682614 541497 682782
rect 541531 682614 541547 682782
rect 541459 682598 541547 682614
rect 541589 682782 541677 682798
rect 541589 682614 541605 682782
rect 541639 682614 541677 682782
rect 541589 682598 541677 682614
rect 542677 682782 542765 682798
rect 542677 682614 542715 682782
rect 542749 682614 542765 682782
rect 542677 682598 542765 682614
rect 542807 682782 542895 682798
rect 542807 682614 542823 682782
rect 542857 682614 542895 682782
rect 542807 682598 542895 682614
rect 543895 682782 543983 682798
rect 543895 682614 543933 682782
rect 543967 682614 543983 682782
rect 543895 682598 543983 682614
rect 544025 682782 544113 682798
rect 544025 682614 544041 682782
rect 544075 682614 544113 682782
rect 544025 682598 544113 682614
rect 545113 682782 545201 682798
rect 545113 682614 545151 682782
rect 545185 682614 545201 682782
rect 545113 682598 545201 682614
rect 545243 682782 545331 682798
rect 545243 682614 545259 682782
rect 545293 682614 545331 682782
rect 545243 682598 545331 682614
rect 546331 682782 546419 682798
rect 546331 682614 546369 682782
rect 546403 682614 546419 682782
rect 546331 682598 546419 682614
rect 546461 682782 546549 682798
rect 546461 682614 546477 682782
rect 546511 682614 546549 682782
rect 546461 682598 546549 682614
rect 547549 682782 547637 682798
rect 547549 682614 547587 682782
rect 547621 682614 547637 682782
rect 547549 682598 547637 682614
rect 547679 682782 547767 682798
rect 547679 682614 547695 682782
rect 547729 682614 547767 682782
rect 547679 682598 547767 682614
rect 548767 682782 548855 682798
rect 548767 682614 548805 682782
rect 548839 682614 548855 682782
rect 548767 682598 548855 682614
rect 43906 682400 44106 682416
rect 43906 682366 43922 682400
rect 44090 682366 44106 682400
rect 43906 682319 44106 682366
rect 44164 682400 44364 682416
rect 44164 682366 44180 682400
rect 44348 682366 44364 682400
rect 44164 682319 44364 682366
rect 44422 682400 44622 682416
rect 44422 682366 44438 682400
rect 44606 682366 44622 682400
rect 44422 682319 44622 682366
rect 44680 682400 44880 682416
rect 44680 682366 44696 682400
rect 44864 682366 44880 682400
rect 44680 682319 44880 682366
rect 44938 682400 45138 682416
rect 44938 682366 44954 682400
rect 45122 682366 45138 682400
rect 44938 682319 45138 682366
rect 45196 682400 45396 682416
rect 45196 682366 45212 682400
rect 45380 682366 45396 682400
rect 45196 682319 45396 682366
rect 43906 681272 44106 681319
rect 43906 681238 43922 681272
rect 44090 681238 44106 681272
rect 43906 681222 44106 681238
rect 44164 681272 44364 681319
rect 44164 681238 44180 681272
rect 44348 681238 44364 681272
rect 44164 681222 44364 681238
rect 44422 681272 44622 681319
rect 44422 681238 44438 681272
rect 44606 681238 44622 681272
rect 44422 681222 44622 681238
rect 44680 681272 44880 681319
rect 44680 681238 44696 681272
rect 44864 681238 44880 681272
rect 44680 681222 44880 681238
rect 44938 681272 45138 681319
rect 44938 681238 44954 681272
rect 45122 681238 45138 681272
rect 44938 681222 45138 681238
rect 45196 681272 45396 681319
rect 45196 681238 45212 681272
rect 45380 681238 45396 681272
rect 45196 681222 45396 681238
rect 540371 682182 540459 682198
rect 540371 682014 540387 682182
rect 540421 682014 540459 682182
rect 540371 681998 540459 682014
rect 541459 682182 541547 682198
rect 541459 682014 541497 682182
rect 541531 682014 541547 682182
rect 541459 681998 541547 682014
rect 541589 682182 541677 682198
rect 541589 682014 541605 682182
rect 541639 682014 541677 682182
rect 541589 681998 541677 682014
rect 542677 682182 542765 682198
rect 542677 682014 542715 682182
rect 542749 682014 542765 682182
rect 542677 681998 542765 682014
rect 542807 682182 542895 682198
rect 542807 682014 542823 682182
rect 542857 682014 542895 682182
rect 542807 681998 542895 682014
rect 543895 682182 543983 682198
rect 543895 682014 543933 682182
rect 543967 682014 543983 682182
rect 543895 681998 543983 682014
rect 544025 682182 544113 682198
rect 544025 682014 544041 682182
rect 544075 682014 544113 682182
rect 544025 681998 544113 682014
rect 545113 682182 545201 682198
rect 545113 682014 545151 682182
rect 545185 682014 545201 682182
rect 545113 681998 545201 682014
rect 545243 682182 545331 682198
rect 545243 682014 545259 682182
rect 545293 682014 545331 682182
rect 545243 681998 545331 682014
rect 546331 682182 546419 682198
rect 546331 682014 546369 682182
rect 546403 682014 546419 682182
rect 546331 681998 546419 682014
rect 546461 682182 546549 682198
rect 546461 682014 546477 682182
rect 546511 682014 546549 682182
rect 546461 681998 546549 682014
rect 547549 682182 547637 682198
rect 547549 682014 547587 682182
rect 547621 682014 547637 682182
rect 547549 681998 547637 682014
rect 547679 682182 547767 682198
rect 547679 682014 547695 682182
rect 547729 682014 547767 682182
rect 547679 681998 547767 682014
rect 548767 682182 548855 682198
rect 548767 682014 548805 682182
rect 548839 682014 548855 682182
rect 548767 681998 548855 682014
rect 540916 681208 541013 681224
rect 540916 681040 540932 681208
rect 540966 681040 541013 681208
rect 540916 681024 541013 681040
rect 542013 681208 542110 681224
rect 542013 681040 542060 681208
rect 542094 681040 542110 681208
rect 542013 681024 542110 681040
rect 542152 681208 542249 681224
rect 542152 681040 542168 681208
rect 542202 681040 542249 681208
rect 542152 681024 542249 681040
rect 543249 681208 543346 681224
rect 543249 681040 543296 681208
rect 543330 681040 543346 681208
rect 543249 681024 543346 681040
rect 543388 681208 543485 681224
rect 543388 681040 543404 681208
rect 543438 681040 543485 681208
rect 543388 681024 543485 681040
rect 544485 681208 544582 681224
rect 544485 681040 544532 681208
rect 544566 681040 544582 681208
rect 544485 681024 544582 681040
rect 544624 681208 544721 681224
rect 544624 681040 544640 681208
rect 544674 681040 544721 681208
rect 544624 681024 544721 681040
rect 545721 681208 545818 681224
rect 545721 681040 545768 681208
rect 545802 681040 545818 681208
rect 545721 681024 545818 681040
rect 545860 681208 545957 681224
rect 545860 681040 545876 681208
rect 545910 681040 545957 681208
rect 545860 681024 545957 681040
rect 546957 681208 547054 681224
rect 546957 681040 547004 681208
rect 547038 681040 547054 681208
rect 546957 681024 547054 681040
rect 547096 681208 547193 681224
rect 547096 681040 547112 681208
rect 547146 681040 547193 681208
rect 547096 681024 547193 681040
rect 548193 681208 548290 681224
rect 548193 681040 548240 681208
rect 548274 681040 548290 681208
rect 548193 681024 548290 681040
rect 44506 680782 44606 680798
rect 44506 680748 44522 680782
rect 44590 680748 44606 680782
rect 44506 680710 44606 680748
rect 44664 680782 44764 680798
rect 44664 680748 44680 680782
rect 44748 680748 44764 680782
rect 44664 680710 44764 680748
rect 44506 680172 44606 680210
rect 44506 680138 44522 680172
rect 44590 680138 44606 680172
rect 44506 680122 44606 680138
rect 44664 680172 44764 680210
rect 44664 680138 44680 680172
rect 44748 680138 44764 680172
rect 44664 680122 44764 680138
rect 540916 680618 541013 680634
rect 540916 680450 540932 680618
rect 540966 680450 541013 680618
rect 540916 680434 541013 680450
rect 542013 680618 542110 680634
rect 542013 680450 542060 680618
rect 542094 680450 542110 680618
rect 542013 680434 542110 680450
rect 542152 680618 542249 680634
rect 542152 680450 542168 680618
rect 542202 680450 542249 680618
rect 542152 680434 542249 680450
rect 543249 680618 543346 680634
rect 543249 680450 543296 680618
rect 543330 680450 543346 680618
rect 543249 680434 543346 680450
rect 543388 680618 543485 680634
rect 543388 680450 543404 680618
rect 543438 680450 543485 680618
rect 543388 680434 543485 680450
rect 544485 680618 544582 680634
rect 544485 680450 544532 680618
rect 544566 680450 544582 680618
rect 544485 680434 544582 680450
rect 544624 680618 544721 680634
rect 544624 680450 544640 680618
rect 544674 680450 544721 680618
rect 544624 680434 544721 680450
rect 545721 680618 545818 680634
rect 545721 680450 545768 680618
rect 545802 680450 545818 680618
rect 545721 680434 545818 680450
rect 545860 680618 545957 680634
rect 545860 680450 545876 680618
rect 545910 680450 545957 680618
rect 545860 680434 545957 680450
rect 546957 680618 547054 680634
rect 546957 680450 547004 680618
rect 547038 680450 547054 680618
rect 546957 680434 547054 680450
rect 547096 680618 547193 680634
rect 547096 680450 547112 680618
rect 547146 680450 547193 680618
rect 547096 680434 547193 680450
rect 548193 680618 548290 680634
rect 548193 680450 548240 680618
rect 548274 680450 548290 680618
rect 548193 680434 548290 680450
rect 44146 679782 44346 679798
rect 44146 679748 44162 679782
rect 44330 679748 44346 679782
rect 44146 679710 44346 679748
rect 44404 679782 44604 679798
rect 44404 679748 44420 679782
rect 44588 679748 44604 679782
rect 44404 679710 44604 679748
rect 44662 679782 44862 679798
rect 44662 679748 44678 679782
rect 44846 679748 44862 679782
rect 44662 679710 44862 679748
rect 44920 679782 45120 679798
rect 44920 679748 44936 679782
rect 45104 679748 45120 679782
rect 44920 679710 45120 679748
rect 44146 679422 44346 679460
rect 44146 679388 44162 679422
rect 44330 679388 44346 679422
rect 44146 679372 44346 679388
rect 44404 679422 44604 679460
rect 44404 679388 44420 679422
rect 44588 679388 44604 679422
rect 44404 679372 44604 679388
rect 44662 679422 44862 679460
rect 44662 679388 44678 679422
rect 44846 679388 44862 679422
rect 44662 679372 44862 679388
rect 44920 679422 45120 679460
rect 44920 679388 44936 679422
rect 45104 679388 45120 679422
rect 44920 679372 45120 679388
rect 543686 679828 543774 679844
rect 543686 679660 543702 679828
rect 543736 679660 543774 679828
rect 543686 679644 543774 679660
rect 544024 679828 544112 679844
rect 544024 679660 544062 679828
rect 544096 679660 544112 679828
rect 544024 679644 544112 679660
rect 544154 679828 544242 679844
rect 544154 679660 544170 679828
rect 544204 679660 544242 679828
rect 544154 679644 544242 679660
rect 544492 679828 544580 679844
rect 544492 679660 544530 679828
rect 544564 679660 544580 679828
rect 544492 679644 544580 679660
rect 544622 679828 544710 679844
rect 544622 679660 544638 679828
rect 544672 679660 544710 679828
rect 544622 679644 544710 679660
rect 544960 679828 545048 679844
rect 544960 679660 544998 679828
rect 545032 679660 545048 679828
rect 544960 679644 545048 679660
rect 545090 679828 545178 679844
rect 545090 679660 545106 679828
rect 545140 679660 545178 679828
rect 545090 679644 545178 679660
rect 545428 679828 545516 679844
rect 545428 679660 545466 679828
rect 545500 679660 545516 679828
rect 545428 679644 545516 679660
rect 43891 679032 44091 679048
rect 43891 678998 43907 679032
rect 44075 678998 44091 679032
rect 43891 678960 44091 678998
rect 44149 679032 44349 679048
rect 44149 678998 44165 679032
rect 44333 678998 44349 679032
rect 44149 678960 44349 678998
rect 44407 679032 44607 679048
rect 44407 678998 44423 679032
rect 44591 678998 44607 679032
rect 44407 678960 44607 678998
rect 44665 679032 44865 679048
rect 44665 678998 44681 679032
rect 44849 678998 44865 679032
rect 44665 678960 44865 678998
rect 44923 679032 45123 679048
rect 44923 678998 44939 679032
rect 45107 678998 45123 679032
rect 44923 678960 45123 678998
rect 45181 679032 45381 679048
rect 45181 678998 45197 679032
rect 45365 678998 45381 679032
rect 45181 678960 45381 678998
rect 43891 677922 44091 677960
rect 43891 677888 43907 677922
rect 44075 677888 44091 677922
rect 43891 677872 44091 677888
rect 44149 677922 44349 677960
rect 44149 677888 44165 677922
rect 44333 677888 44349 677922
rect 44149 677872 44349 677888
rect 44407 677922 44607 677960
rect 44407 677888 44423 677922
rect 44591 677888 44607 677922
rect 44407 677872 44607 677888
rect 44665 677922 44865 677960
rect 44665 677888 44681 677922
rect 44849 677888 44865 677922
rect 44665 677872 44865 677888
rect 44923 677922 45123 677960
rect 44923 677888 44939 677922
rect 45107 677888 45123 677922
rect 44923 677872 45123 677888
rect 45181 677922 45381 677960
rect 45181 677888 45197 677922
rect 45365 677888 45381 677922
rect 45181 677872 45381 677888
rect 543906 679203 543994 679219
rect 543906 679135 543922 679203
rect 543956 679135 543994 679203
rect 543906 679119 543994 679135
rect 544494 679203 544582 679219
rect 544494 679135 544532 679203
rect 544566 679135 544582 679203
rect 544494 679119 544582 679135
rect 544624 679203 544712 679219
rect 544624 679135 544640 679203
rect 544674 679135 544712 679203
rect 544624 679119 544712 679135
rect 545212 679203 545300 679219
rect 545212 679135 545250 679203
rect 545284 679135 545300 679203
rect 545212 679119 545300 679135
rect 540971 678678 541059 678694
rect 540971 678510 540987 678678
rect 541021 678510 541059 678678
rect 540971 678494 541059 678510
rect 542059 678678 542147 678694
rect 542059 678510 542097 678678
rect 542131 678510 542147 678678
rect 542059 678494 542147 678510
rect 542189 678678 542277 678694
rect 542189 678510 542205 678678
rect 542239 678510 542277 678678
rect 542189 678494 542277 678510
rect 543277 678678 543365 678694
rect 543277 678510 543315 678678
rect 543349 678510 543365 678678
rect 543277 678494 543365 678510
rect 543407 678678 543495 678694
rect 543407 678510 543423 678678
rect 543457 678510 543495 678678
rect 543407 678494 543495 678510
rect 544495 678678 544583 678694
rect 544495 678510 544533 678678
rect 544567 678510 544583 678678
rect 544495 678494 544583 678510
rect 544625 678678 544713 678694
rect 544625 678510 544641 678678
rect 544675 678510 544713 678678
rect 544625 678494 544713 678510
rect 545713 678678 545801 678694
rect 545713 678510 545751 678678
rect 545785 678510 545801 678678
rect 545713 678494 545801 678510
rect 545843 678678 545931 678694
rect 545843 678510 545859 678678
rect 545893 678510 545931 678678
rect 545843 678494 545931 678510
rect 546931 678678 547019 678694
rect 546931 678510 546969 678678
rect 547003 678510 547019 678678
rect 546931 678494 547019 678510
rect 547061 678678 547149 678694
rect 547061 678510 547077 678678
rect 547111 678510 547149 678678
rect 547061 678494 547149 678510
rect 548149 678678 548237 678694
rect 548149 678510 548187 678678
rect 548221 678510 548237 678678
rect 548149 678494 548237 678510
<< polycont >>
rect 41542 695246 41610 695280
rect 41700 695246 41768 695280
rect 41858 695246 41926 695280
rect 42016 695246 42084 695280
rect 42174 695246 42242 695280
rect 42332 695246 42400 695280
rect 42490 695246 42558 695280
rect 42648 695246 42716 695280
rect 42806 695246 42874 695280
rect 42964 695246 43032 695280
rect 43122 695246 43190 695280
rect 43280 695246 43348 695280
rect 43438 695246 43506 695280
rect 43596 695246 43664 695280
rect 43754 695246 43822 695280
rect 43912 695246 43980 695280
rect 44070 695246 44138 695280
rect 44228 695246 44296 695280
rect 44386 695246 44454 695280
rect 44544 695246 44612 695280
rect 44702 695246 44770 695280
rect 44860 695246 44928 695280
rect 45018 695246 45086 695280
rect 45176 695246 45244 695280
rect 45334 695246 45402 695280
rect 45492 695246 45560 695280
rect 45650 695246 45718 695280
rect 45808 695246 45876 695280
rect 45966 695246 46034 695280
rect 46124 695246 46192 695280
rect 46282 695246 46350 695280
rect 46440 695246 46508 695280
rect 46598 695246 46666 695280
rect 46756 695246 46824 695280
rect 46914 695246 46982 695280
rect 47072 695246 47140 695280
rect 47230 695246 47298 695280
rect 47388 695246 47456 695280
rect 47546 695246 47614 695280
rect 47704 695246 47772 695280
rect 41542 694118 41610 694152
rect 41700 694118 41768 694152
rect 41858 694118 41926 694152
rect 42016 694118 42084 694152
rect 42174 694118 42242 694152
rect 42332 694118 42400 694152
rect 42490 694118 42558 694152
rect 42648 694118 42716 694152
rect 42806 694118 42874 694152
rect 42964 694118 43032 694152
rect 43122 694118 43190 694152
rect 43280 694118 43348 694152
rect 43438 694118 43506 694152
rect 43596 694118 43664 694152
rect 43754 694118 43822 694152
rect 43912 694118 43980 694152
rect 44070 694118 44138 694152
rect 44228 694118 44296 694152
rect 44386 694118 44454 694152
rect 44544 694118 44612 694152
rect 44702 694118 44770 694152
rect 44860 694118 44928 694152
rect 45018 694118 45086 694152
rect 45176 694118 45244 694152
rect 45334 694118 45402 694152
rect 45492 694118 45560 694152
rect 45650 694118 45718 694152
rect 45808 694118 45876 694152
rect 45966 694118 46034 694152
rect 46124 694118 46192 694152
rect 46282 694118 46350 694152
rect 46440 694118 46508 694152
rect 46598 694118 46666 694152
rect 46756 694118 46824 694152
rect 46914 694118 46982 694152
rect 47072 694118 47140 694152
rect 47230 694118 47298 694152
rect 47388 694118 47456 694152
rect 47546 694118 47614 694152
rect 47704 694118 47772 694152
rect 43042 693576 43110 693610
rect 43200 693576 43268 693610
rect 43358 693576 43426 693610
rect 43516 693576 43584 693610
rect 43674 693576 43742 693610
rect 43832 693576 43900 693610
rect 43990 693576 44058 693610
rect 44148 693576 44216 693610
rect 44306 693576 44374 693610
rect 44464 693576 44532 693610
rect 44622 693576 44690 693610
rect 44780 693576 44848 693610
rect 44938 693576 45006 693610
rect 45096 693576 45164 693610
rect 45254 693576 45322 693610
rect 45412 693576 45480 693610
rect 45570 693576 45638 693610
rect 45728 693576 45796 693610
rect 45886 693576 45954 693610
rect 46044 693576 46112 693610
rect 46202 693576 46270 693610
rect 43042 692448 43110 692482
rect 43200 692448 43268 692482
rect 43358 692448 43426 692482
rect 43516 692448 43584 692482
rect 43674 692448 43742 692482
rect 43832 692448 43900 692482
rect 43990 692448 44058 692482
rect 44148 692448 44216 692482
rect 44306 692448 44374 692482
rect 44464 692448 44532 692482
rect 44622 692448 44690 692482
rect 44780 692448 44848 692482
rect 44938 692448 45006 692482
rect 45096 692448 45164 692482
rect 45254 692448 45322 692482
rect 45412 692448 45480 692482
rect 45570 692448 45638 692482
rect 45728 692448 45796 692482
rect 45886 692448 45954 692482
rect 46044 692448 46112 692482
rect 46202 692448 46270 692482
rect 43042 692036 43110 692070
rect 43200 692036 43268 692070
rect 43358 692036 43426 692070
rect 43516 692036 43584 692070
rect 43674 692036 43742 692070
rect 43832 692036 43900 692070
rect 43990 692036 44058 692070
rect 44148 692036 44216 692070
rect 44306 692036 44374 692070
rect 44464 692036 44532 692070
rect 44622 692036 44690 692070
rect 44780 692036 44848 692070
rect 44938 692036 45006 692070
rect 45096 692036 45164 692070
rect 45254 692036 45322 692070
rect 45412 692036 45480 692070
rect 45570 692036 45638 692070
rect 45728 692036 45796 692070
rect 45886 692036 45954 692070
rect 46044 692036 46112 692070
rect 46202 692036 46270 692070
rect 43042 690908 43110 690942
rect 43200 690908 43268 690942
rect 43358 690908 43426 690942
rect 43516 690908 43584 690942
rect 43674 690908 43742 690942
rect 43832 690908 43900 690942
rect 43990 690908 44058 690942
rect 44148 690908 44216 690942
rect 44306 690908 44374 690942
rect 44464 690908 44532 690942
rect 44622 690908 44690 690942
rect 44780 690908 44848 690942
rect 44938 690908 45006 690942
rect 45096 690908 45164 690942
rect 45254 690908 45322 690942
rect 45412 690908 45480 690942
rect 45570 690908 45638 690942
rect 45728 690908 45796 690942
rect 45886 690908 45954 690942
rect 46044 690908 46112 690942
rect 46202 690908 46270 690942
rect 44143 690459 44211 690493
rect 44301 690459 44369 690493
rect 44459 690459 44527 690493
rect 44617 690459 44685 690493
rect 44775 690459 44843 690493
rect 44933 690459 45001 690493
rect 45091 690459 45159 690493
rect 44143 689349 44211 689383
rect 44301 689349 44369 689383
rect 44459 689349 44527 689383
rect 44617 689349 44685 689383
rect 44775 689349 44843 689383
rect 44933 689349 45001 689383
rect 45091 689349 45159 689383
rect 540287 690654 540321 690722
rect 541415 690654 541449 690722
rect 541523 690654 541557 690722
rect 542651 690654 542685 690722
rect 542759 690654 542793 690722
rect 543887 690654 543921 690722
rect 543995 690654 544029 690722
rect 545123 690654 545157 690722
rect 545231 690654 545265 690722
rect 546359 690654 546393 690722
rect 546467 690654 546501 690722
rect 547595 690654 547629 690722
rect 547703 690654 547737 690722
rect 548831 690654 548865 690722
rect 540287 690114 540321 690182
rect 541415 690114 541449 690182
rect 541523 690114 541557 690182
rect 542651 690114 542685 690182
rect 542759 690114 542793 690182
rect 543887 690114 543921 690182
rect 543995 690114 544029 690182
rect 545123 690114 545157 690182
rect 545231 690114 545265 690182
rect 546359 690114 546393 690182
rect 546467 690114 546501 690182
rect 547595 690114 547629 690182
rect 547703 690114 547737 690182
rect 548831 690114 548865 690182
rect 540287 689574 540321 689642
rect 541415 689574 541449 689642
rect 541523 689574 541557 689642
rect 542651 689574 542685 689642
rect 542759 689574 542793 689642
rect 543887 689574 543921 689642
rect 543995 689574 544029 689642
rect 545123 689574 545157 689642
rect 545231 689574 545265 689642
rect 546359 689574 546393 689642
rect 546467 689574 546501 689642
rect 547595 689574 547629 689642
rect 547703 689574 547737 689642
rect 548831 689574 548865 689642
rect 44143 688939 44211 688973
rect 44301 688939 44369 688973
rect 44459 688939 44527 688973
rect 44617 688939 44685 688973
rect 44775 688939 44843 688973
rect 44933 688939 45001 688973
rect 45091 688939 45159 688973
rect 44143 687829 44211 687863
rect 44301 687829 44369 687863
rect 44459 687829 44527 687863
rect 44617 687829 44685 687863
rect 44775 687829 44843 687863
rect 44933 687829 45001 687863
rect 45091 687829 45159 687863
rect 540287 689034 540321 689102
rect 541415 689034 541449 689102
rect 541523 689034 541557 689102
rect 542651 689034 542685 689102
rect 542759 689034 542793 689102
rect 543887 689034 543921 689102
rect 543995 689034 544029 689102
rect 545123 689034 545157 689102
rect 545231 689034 545265 689102
rect 546359 689034 546393 689102
rect 546467 689034 546501 689102
rect 547595 689034 547629 689102
rect 547703 689034 547737 689102
rect 548831 689034 548865 689102
rect 540287 688454 540321 688522
rect 541415 688454 541449 688522
rect 541523 688454 541557 688522
rect 542651 688454 542685 688522
rect 542759 688454 542793 688522
rect 543887 688454 543921 688522
rect 543995 688454 544029 688522
rect 545123 688454 545157 688522
rect 545231 688454 545265 688522
rect 546359 688454 546393 688522
rect 546467 688454 546501 688522
rect 547595 688454 547629 688522
rect 547703 688454 547737 688522
rect 548831 688454 548865 688522
rect 43152 687418 43320 687452
rect 43410 687418 43578 687452
rect 43668 687418 43836 687452
rect 43926 687418 44094 687452
rect 44184 687418 44352 687452
rect 44442 687418 44610 687452
rect 44700 687418 44868 687452
rect 44958 687418 45126 687452
rect 45216 687418 45384 687452
rect 45474 687418 45642 687452
rect 45732 687418 45900 687452
rect 45990 687418 46158 687452
rect 43152 686308 43320 686342
rect 43410 686308 43578 686342
rect 43668 686308 43836 686342
rect 43926 686308 44094 686342
rect 44184 686308 44352 686342
rect 44442 686308 44610 686342
rect 44700 686308 44868 686342
rect 44958 686308 45126 686342
rect 45216 686308 45384 686342
rect 45474 686308 45642 686342
rect 45732 686308 45900 686342
rect 45990 686308 46158 686342
rect 540287 687874 540321 687942
rect 541415 687874 541449 687942
rect 541523 687874 541557 687942
rect 542651 687874 542685 687942
rect 542759 687874 542793 687942
rect 543887 687874 543921 687942
rect 543995 687874 544029 687942
rect 545123 687874 545157 687942
rect 545231 687874 545265 687942
rect 546359 687874 546393 687942
rect 546467 687874 546501 687942
rect 547595 687874 547629 687942
rect 547703 687874 547737 687942
rect 548831 687874 548865 687942
rect 538447 687334 538481 687402
rect 539575 687334 539609 687402
rect 539683 687334 539717 687402
rect 540811 687334 540845 687402
rect 540919 687334 540953 687402
rect 542047 687334 542081 687402
rect 542155 687334 542189 687402
rect 543283 687334 543317 687402
rect 543391 687334 543425 687402
rect 544519 687334 544553 687402
rect 544627 687334 544661 687402
rect 545755 687334 545789 687402
rect 545863 687334 545897 687402
rect 546991 687334 547025 687402
rect 547099 687334 547133 687402
rect 548227 687334 548261 687402
rect 548335 687334 548369 687402
rect 549463 687334 549497 687402
rect 549571 687334 549605 687402
rect 550699 687334 550733 687402
rect 538447 686794 538481 686862
rect 539575 686794 539609 686862
rect 539683 686794 539717 686862
rect 540811 686794 540845 686862
rect 540919 686794 540953 686862
rect 542047 686794 542081 686862
rect 542155 686794 542189 686862
rect 543283 686794 543317 686862
rect 543391 686794 543425 686862
rect 544519 686794 544553 686862
rect 544627 686794 544661 686862
rect 545755 686794 545789 686862
rect 545863 686794 545897 686862
rect 546991 686794 547025 686862
rect 547099 686794 547133 686862
rect 548227 686794 548261 686862
rect 548335 686794 548369 686862
rect 549463 686794 549497 686862
rect 549571 686794 549605 686862
rect 550699 686794 550733 686862
rect 42892 685898 43060 685932
rect 43150 685898 43318 685932
rect 43408 685898 43576 685932
rect 43666 685898 43834 685932
rect 43924 685898 44092 685932
rect 44182 685898 44350 685932
rect 44440 685898 44608 685932
rect 44698 685898 44866 685932
rect 44956 685898 45124 685932
rect 45214 685898 45382 685932
rect 45472 685898 45640 685932
rect 45730 685898 45898 685932
rect 45988 685898 46156 685932
rect 46246 685898 46414 685932
rect 42892 684788 43060 684822
rect 43150 684788 43318 684822
rect 43408 684788 43576 684822
rect 43666 684788 43834 684822
rect 43924 684788 44092 684822
rect 44182 684788 44350 684822
rect 44440 684788 44608 684822
rect 44698 684788 44866 684822
rect 44956 684788 45124 684822
rect 45214 684788 45382 684822
rect 45472 684788 45640 684822
rect 45730 684788 45898 684822
rect 45988 684788 46156 684822
rect 46246 684788 46414 684822
rect 538447 686254 538481 686322
rect 539575 686254 539609 686322
rect 539683 686254 539717 686322
rect 540811 686254 540845 686322
rect 540919 686254 540953 686322
rect 542047 686254 542081 686322
rect 542155 686254 542189 686322
rect 543283 686254 543317 686322
rect 543391 686254 543425 686322
rect 544519 686254 544553 686322
rect 544627 686254 544661 686322
rect 545755 686254 545789 686322
rect 545863 686254 545897 686322
rect 546991 686254 547025 686322
rect 547099 686254 547133 686322
rect 548227 686254 548261 686322
rect 548335 686254 548369 686322
rect 549463 686254 549497 686322
rect 549571 686254 549605 686322
rect 550699 686254 550733 686322
rect 538447 685714 538481 685782
rect 539575 685714 539609 685782
rect 539683 685714 539717 685782
rect 540811 685714 540845 685782
rect 540919 685714 540953 685782
rect 542047 685714 542081 685782
rect 542155 685714 542189 685782
rect 543283 685714 543317 685782
rect 543391 685714 543425 685782
rect 544519 685714 544553 685782
rect 544627 685714 544661 685782
rect 545755 685714 545789 685782
rect 545863 685714 545897 685782
rect 546991 685714 547025 685782
rect 547099 685714 547133 685782
rect 548227 685714 548261 685782
rect 548335 685714 548369 685782
rect 549463 685714 549497 685782
rect 549571 685714 549605 685782
rect 550699 685714 550733 685782
rect 540387 684934 540421 685002
rect 541497 684934 541531 685002
rect 541605 684934 541639 685002
rect 542715 684934 542749 685002
rect 542823 684934 542857 685002
rect 543933 684934 543967 685002
rect 544041 684934 544075 685002
rect 545151 684934 545185 685002
rect 545259 684934 545293 685002
rect 546369 684934 546403 685002
rect 546477 684934 546511 685002
rect 547587 684934 547621 685002
rect 547695 684934 547729 685002
rect 548805 684934 548839 685002
rect 540387 684434 540421 684502
rect 541497 684434 541531 684502
rect 541605 684434 541639 684502
rect 542715 684434 542749 684502
rect 542823 684434 542857 684502
rect 543933 684434 543967 684502
rect 544041 684434 544075 684502
rect 545151 684434 545185 684502
rect 545259 684434 545293 684502
rect 546369 684434 546403 684502
rect 546477 684434 546511 684502
rect 547587 684434 547621 684502
rect 547695 684434 547729 684502
rect 548805 684434 548839 684502
rect 43922 683866 44090 683900
rect 44180 683866 44348 683900
rect 44438 683866 44606 683900
rect 44696 683866 44864 683900
rect 44954 683866 45122 683900
rect 45212 683866 45380 683900
rect 43922 682738 44090 682772
rect 44180 682738 44348 682772
rect 44438 682738 44606 682772
rect 44696 682738 44864 682772
rect 44954 682738 45122 682772
rect 45212 682738 45380 682772
rect 540947 683834 540981 684002
rect 542057 683834 542091 684002
rect 542165 683834 542199 684002
rect 543275 683834 543309 684002
rect 543383 683834 543417 684002
rect 544493 683834 544527 684002
rect 544601 683834 544635 684002
rect 545711 683834 545745 684002
rect 545819 683834 545853 684002
rect 546929 683834 546963 684002
rect 547037 683834 547071 684002
rect 548147 683834 548181 684002
rect 540947 683214 540981 683382
rect 542057 683214 542091 683382
rect 542165 683214 542199 683382
rect 543275 683214 543309 683382
rect 543383 683214 543417 683382
rect 544493 683214 544527 683382
rect 544601 683214 544635 683382
rect 545711 683214 545745 683382
rect 545819 683214 545853 683382
rect 546929 683214 546963 683382
rect 547037 683214 547071 683382
rect 548147 683214 548181 683382
rect 540387 682614 540421 682782
rect 541497 682614 541531 682782
rect 541605 682614 541639 682782
rect 542715 682614 542749 682782
rect 542823 682614 542857 682782
rect 543933 682614 543967 682782
rect 544041 682614 544075 682782
rect 545151 682614 545185 682782
rect 545259 682614 545293 682782
rect 546369 682614 546403 682782
rect 546477 682614 546511 682782
rect 547587 682614 547621 682782
rect 547695 682614 547729 682782
rect 548805 682614 548839 682782
rect 43922 682366 44090 682400
rect 44180 682366 44348 682400
rect 44438 682366 44606 682400
rect 44696 682366 44864 682400
rect 44954 682366 45122 682400
rect 45212 682366 45380 682400
rect 43922 681238 44090 681272
rect 44180 681238 44348 681272
rect 44438 681238 44606 681272
rect 44696 681238 44864 681272
rect 44954 681238 45122 681272
rect 45212 681238 45380 681272
rect 540387 682014 540421 682182
rect 541497 682014 541531 682182
rect 541605 682014 541639 682182
rect 542715 682014 542749 682182
rect 542823 682014 542857 682182
rect 543933 682014 543967 682182
rect 544041 682014 544075 682182
rect 545151 682014 545185 682182
rect 545259 682014 545293 682182
rect 546369 682014 546403 682182
rect 546477 682014 546511 682182
rect 547587 682014 547621 682182
rect 547695 682014 547729 682182
rect 548805 682014 548839 682182
rect 540932 681040 540966 681208
rect 542060 681040 542094 681208
rect 542168 681040 542202 681208
rect 543296 681040 543330 681208
rect 543404 681040 543438 681208
rect 544532 681040 544566 681208
rect 544640 681040 544674 681208
rect 545768 681040 545802 681208
rect 545876 681040 545910 681208
rect 547004 681040 547038 681208
rect 547112 681040 547146 681208
rect 548240 681040 548274 681208
rect 44522 680748 44590 680782
rect 44680 680748 44748 680782
rect 44522 680138 44590 680172
rect 44680 680138 44748 680172
rect 540932 680450 540966 680618
rect 542060 680450 542094 680618
rect 542168 680450 542202 680618
rect 543296 680450 543330 680618
rect 543404 680450 543438 680618
rect 544532 680450 544566 680618
rect 544640 680450 544674 680618
rect 545768 680450 545802 680618
rect 545876 680450 545910 680618
rect 547004 680450 547038 680618
rect 547112 680450 547146 680618
rect 548240 680450 548274 680618
rect 44162 679748 44330 679782
rect 44420 679748 44588 679782
rect 44678 679748 44846 679782
rect 44936 679748 45104 679782
rect 44162 679388 44330 679422
rect 44420 679388 44588 679422
rect 44678 679388 44846 679422
rect 44936 679388 45104 679422
rect 543702 679660 543736 679828
rect 544062 679660 544096 679828
rect 544170 679660 544204 679828
rect 544530 679660 544564 679828
rect 544638 679660 544672 679828
rect 544998 679660 545032 679828
rect 545106 679660 545140 679828
rect 545466 679660 545500 679828
rect 43907 678998 44075 679032
rect 44165 678998 44333 679032
rect 44423 678998 44591 679032
rect 44681 678998 44849 679032
rect 44939 678998 45107 679032
rect 45197 678998 45365 679032
rect 43907 677888 44075 677922
rect 44165 677888 44333 677922
rect 44423 677888 44591 677922
rect 44681 677888 44849 677922
rect 44939 677888 45107 677922
rect 45197 677888 45365 677922
rect 543922 679135 543956 679203
rect 544532 679135 544566 679203
rect 544640 679135 544674 679203
rect 545250 679135 545284 679203
rect 540987 678510 541021 678678
rect 542097 678510 542131 678678
rect 542205 678510 542239 678678
rect 543315 678510 543349 678678
rect 543423 678510 543457 678678
rect 544533 678510 544567 678678
rect 544641 678510 544675 678678
rect 545751 678510 545785 678678
rect 545859 678510 545893 678678
rect 546969 678510 547003 678678
rect 547077 678510 547111 678678
rect 548187 678510 548221 678678
<< xpolycontact >>
rect 37693 694983 38125 696129
rect 40125 694983 40557 696129
rect 37693 693523 38125 694669
rect 40125 693523 40557 694669
rect 48763 694983 49195 696129
rect 51195 694983 51627 696129
rect 48763 693523 49195 694669
rect 51195 693523 51627 694669
rect 534722 686825 535154 687971
rect 537154 686825 537586 687971
rect 551782 686825 552214 687971
rect 554214 686825 554646 687971
rect 534722 685355 535154 686501
rect 537154 685355 537586 686501
rect 551782 685355 552214 686501
rect 554214 685355 554646 686501
rect 541761 677570 542907 678002
rect 41722 677112 42868 677544
rect 41722 662880 42868 663312
rect 43272 677112 44418 677544
rect 43272 662880 44418 663312
rect 44812 677112 45958 677544
rect 44812 662880 45958 663312
rect 46362 677112 47508 677544
rect 541761 663338 542907 663770
rect 543281 677570 544427 678002
rect 543281 663338 544427 663770
rect 544791 677576 545937 678008
rect 544791 663344 545937 663776
rect 546301 677576 547447 678008
rect 546301 663344 547447 663776
rect 46362 662880 47508 663312
<< xpolyres >>
rect 38125 694983 40125 696129
rect 38125 693523 40125 694669
rect 49195 694983 51195 696129
rect 49195 693523 51195 694669
rect 535154 686825 537154 687971
rect 552214 686825 554214 687971
rect 535154 685355 537154 686501
rect 552214 685355 554214 686501
rect 41722 663312 42868 677112
rect 43272 663312 44418 677112
rect 44812 663312 45958 677112
rect 46362 663312 47508 677112
rect 541761 663770 542907 677570
rect 543281 663770 544427 677570
rect 544791 663776 545937 677576
rect 546301 663776 547447 677576
<< locali >>
rect 37563 696225 37659 696259
rect 40591 696225 40687 696259
rect 37563 696163 37597 696225
rect 40653 696163 40687 696225
rect 37563 694887 37597 694949
rect 48633 696225 48729 696259
rect 51661 696225 51757 696259
rect 48633 696163 48667 696225
rect 38670 694887 39330 694890
rect 40653 694887 40687 694949
rect 37563 694853 37659 694887
rect 40591 694853 40687 694887
rect 41366 695348 41462 695382
rect 47852 695348 47948 695382
rect 41366 695286 41400 695348
rect 38670 694799 39330 694853
rect 37563 694765 37659 694799
rect 40591 694765 40687 694799
rect 37563 694703 37597 694765
rect 40653 694703 40687 694765
rect 37563 693427 37597 693489
rect 47914 695286 47948 695348
rect 41526 695246 41542 695280
rect 41610 695246 41626 695280
rect 41684 695246 41700 695280
rect 41768 695246 41784 695280
rect 41842 695246 41858 695280
rect 41926 695246 41942 695280
rect 42000 695246 42016 695280
rect 42084 695246 42100 695280
rect 42158 695246 42174 695280
rect 42242 695246 42258 695280
rect 42316 695246 42332 695280
rect 42400 695246 42416 695280
rect 42474 695246 42490 695280
rect 42558 695246 42574 695280
rect 42632 695246 42648 695280
rect 42716 695246 42732 695280
rect 42790 695246 42806 695280
rect 42874 695246 42890 695280
rect 42948 695246 42964 695280
rect 43032 695246 43048 695280
rect 43106 695246 43122 695280
rect 43190 695246 43206 695280
rect 43264 695246 43280 695280
rect 43348 695246 43364 695280
rect 43422 695246 43438 695280
rect 43506 695246 43522 695280
rect 43580 695246 43596 695280
rect 43664 695246 43680 695280
rect 43738 695246 43754 695280
rect 43822 695246 43838 695280
rect 43896 695246 43912 695280
rect 43980 695246 43996 695280
rect 44054 695246 44070 695280
rect 44138 695246 44154 695280
rect 44212 695246 44228 695280
rect 44296 695246 44312 695280
rect 44370 695246 44386 695280
rect 44454 695246 44470 695280
rect 44528 695246 44544 695280
rect 44612 695246 44628 695280
rect 44686 695246 44702 695280
rect 44770 695246 44786 695280
rect 44844 695246 44860 695280
rect 44928 695246 44944 695280
rect 45002 695246 45018 695280
rect 45086 695246 45102 695280
rect 45160 695246 45176 695280
rect 45244 695246 45260 695280
rect 45318 695246 45334 695280
rect 45402 695246 45418 695280
rect 45476 695246 45492 695280
rect 45560 695246 45576 695280
rect 45634 695246 45650 695280
rect 45718 695246 45734 695280
rect 45792 695246 45808 695280
rect 45876 695246 45892 695280
rect 45950 695246 45966 695280
rect 46034 695246 46050 695280
rect 46108 695246 46124 695280
rect 46192 695246 46208 695280
rect 46266 695246 46282 695280
rect 46350 695246 46366 695280
rect 46424 695246 46440 695280
rect 46508 695246 46524 695280
rect 46582 695246 46598 695280
rect 46666 695246 46682 695280
rect 46740 695246 46756 695280
rect 46824 695246 46840 695280
rect 46898 695246 46914 695280
rect 46982 695246 46998 695280
rect 47056 695246 47072 695280
rect 47140 695246 47156 695280
rect 47214 695246 47230 695280
rect 47298 695246 47314 695280
rect 47372 695246 47388 695280
rect 47456 695246 47472 695280
rect 47530 695246 47546 695280
rect 47614 695246 47630 695280
rect 47688 695246 47704 695280
rect 47772 695246 47788 695280
rect 41480 695187 41514 695203
rect 41480 694195 41514 694211
rect 41638 695187 41672 695203
rect 41638 694195 41672 694211
rect 41796 695187 41830 695203
rect 41796 694195 41830 694211
rect 41954 695187 41988 695203
rect 41954 694195 41988 694211
rect 42112 695187 42146 695203
rect 42112 694195 42146 694211
rect 42270 695187 42304 695203
rect 42270 694195 42304 694211
rect 42428 695187 42462 695203
rect 42428 694195 42462 694211
rect 42586 695187 42620 695203
rect 42586 694195 42620 694211
rect 42744 695187 42778 695203
rect 42744 694195 42778 694211
rect 42902 695187 42936 695203
rect 42902 694195 42936 694211
rect 43060 695187 43094 695203
rect 43060 694195 43094 694211
rect 43218 695187 43252 695203
rect 43218 694195 43252 694211
rect 43376 695187 43410 695203
rect 43376 694195 43410 694211
rect 43534 695187 43568 695203
rect 43534 694195 43568 694211
rect 43692 695187 43726 695203
rect 43692 694195 43726 694211
rect 43850 695187 43884 695203
rect 43850 694195 43884 694211
rect 44008 695187 44042 695203
rect 44008 694195 44042 694211
rect 44166 695187 44200 695203
rect 44166 694195 44200 694211
rect 44324 695187 44358 695203
rect 44324 694195 44358 694211
rect 44482 695187 44516 695203
rect 44482 694195 44516 694211
rect 44640 695187 44674 695203
rect 44640 694195 44674 694211
rect 44798 695187 44832 695203
rect 44798 694195 44832 694211
rect 44956 695187 44990 695203
rect 44956 694195 44990 694211
rect 45114 695187 45148 695203
rect 45114 694195 45148 694211
rect 45272 695187 45306 695203
rect 45272 694195 45306 694211
rect 45430 695187 45464 695203
rect 45430 694195 45464 694211
rect 45588 695187 45622 695203
rect 45588 694195 45622 694211
rect 45746 695187 45780 695203
rect 45746 694195 45780 694211
rect 45904 695187 45938 695203
rect 45904 694195 45938 694211
rect 46062 695187 46096 695203
rect 46062 694195 46096 694211
rect 46220 695187 46254 695203
rect 46220 694195 46254 694211
rect 46378 695187 46412 695203
rect 46378 694195 46412 694211
rect 46536 695187 46570 695203
rect 46536 694195 46570 694211
rect 46694 695187 46728 695203
rect 46694 694195 46728 694211
rect 46852 695187 46886 695203
rect 46852 694195 46886 694211
rect 47010 695187 47044 695203
rect 47010 694195 47044 694211
rect 47168 695187 47202 695203
rect 47168 694195 47202 694211
rect 47326 695187 47360 695203
rect 47326 694195 47360 694211
rect 47484 695187 47518 695203
rect 47484 694195 47518 694211
rect 47642 695187 47676 695203
rect 47642 694195 47676 694211
rect 47800 695187 47834 695203
rect 47800 694195 47834 694211
rect 41526 694118 41542 694152
rect 41610 694118 41626 694152
rect 41684 694118 41700 694152
rect 41768 694118 41784 694152
rect 41842 694118 41858 694152
rect 41926 694118 41942 694152
rect 42000 694118 42016 694152
rect 42084 694118 42100 694152
rect 42158 694118 42174 694152
rect 42242 694118 42258 694152
rect 42316 694118 42332 694152
rect 42400 694118 42416 694152
rect 42474 694118 42490 694152
rect 42558 694118 42574 694152
rect 42632 694118 42648 694152
rect 42716 694118 42732 694152
rect 42790 694118 42806 694152
rect 42874 694118 42890 694152
rect 42948 694118 42964 694152
rect 43032 694118 43048 694152
rect 43106 694118 43122 694152
rect 43190 694118 43206 694152
rect 43264 694118 43280 694152
rect 43348 694118 43364 694152
rect 43422 694118 43438 694152
rect 43506 694118 43522 694152
rect 43580 694118 43596 694152
rect 43664 694118 43680 694152
rect 43738 694118 43754 694152
rect 43822 694118 43838 694152
rect 43896 694118 43912 694152
rect 43980 694118 43996 694152
rect 44054 694118 44070 694152
rect 44138 694118 44154 694152
rect 44212 694118 44228 694152
rect 44296 694118 44312 694152
rect 44370 694118 44386 694152
rect 44454 694118 44470 694152
rect 44528 694118 44544 694152
rect 44612 694118 44628 694152
rect 44686 694118 44702 694152
rect 44770 694118 44786 694152
rect 44844 694118 44860 694152
rect 44928 694118 44944 694152
rect 45002 694118 45018 694152
rect 45086 694118 45102 694152
rect 45160 694118 45176 694152
rect 45244 694118 45260 694152
rect 45318 694118 45334 694152
rect 45402 694118 45418 694152
rect 45476 694118 45492 694152
rect 45560 694118 45576 694152
rect 45634 694118 45650 694152
rect 45718 694118 45734 694152
rect 45792 694118 45808 694152
rect 45876 694118 45892 694152
rect 45950 694118 45966 694152
rect 46034 694118 46050 694152
rect 46108 694118 46124 694152
rect 46192 694118 46208 694152
rect 46266 694118 46282 694152
rect 46350 694118 46366 694152
rect 46424 694118 46440 694152
rect 46508 694118 46524 694152
rect 46582 694118 46598 694152
rect 46666 694118 46682 694152
rect 46740 694118 46756 694152
rect 46824 694118 46840 694152
rect 46898 694118 46914 694152
rect 46982 694118 46998 694152
rect 47056 694118 47072 694152
rect 47140 694118 47156 694152
rect 47214 694118 47230 694152
rect 47298 694118 47314 694152
rect 47372 694118 47388 694152
rect 47456 694118 47472 694152
rect 47530 694118 47546 694152
rect 47614 694118 47630 694152
rect 47688 694118 47704 694152
rect 47772 694118 47788 694152
rect 41366 694050 41400 694112
rect 51723 696163 51757 696225
rect 48633 694887 48667 694949
rect 49920 694887 50580 694890
rect 51723 694887 51757 694949
rect 48633 694853 48729 694887
rect 51661 694853 51757 694887
rect 49920 694799 50580 694853
rect 47914 694050 47948 694112
rect 41366 694016 41462 694050
rect 47852 694016 47948 694050
rect 48633 694765 48729 694799
rect 51661 694765 51757 694799
rect 48633 694703 48667 694765
rect 40653 693427 40687 693489
rect 37563 693393 37659 693427
rect 40591 693393 40687 693427
rect 42866 693678 42962 693712
rect 46350 693678 46446 693712
rect 42866 693616 42900 693678
rect 46412 693616 46446 693678
rect 43026 693576 43042 693610
rect 43110 693576 43126 693610
rect 43184 693576 43200 693610
rect 43268 693576 43284 693610
rect 43342 693576 43358 693610
rect 43426 693576 43442 693610
rect 43500 693576 43516 693610
rect 43584 693576 43600 693610
rect 43658 693576 43674 693610
rect 43742 693576 43758 693610
rect 43816 693576 43832 693610
rect 43900 693576 43916 693610
rect 43974 693576 43990 693610
rect 44058 693576 44074 693610
rect 44132 693576 44148 693610
rect 44216 693576 44232 693610
rect 44290 693576 44306 693610
rect 44374 693576 44390 693610
rect 44448 693576 44464 693610
rect 44532 693576 44548 693610
rect 44606 693576 44622 693610
rect 44690 693576 44706 693610
rect 44764 693576 44780 693610
rect 44848 693576 44864 693610
rect 44922 693576 44938 693610
rect 45006 693576 45022 693610
rect 45080 693576 45096 693610
rect 45164 693576 45180 693610
rect 45238 693576 45254 693610
rect 45322 693576 45338 693610
rect 45396 693576 45412 693610
rect 45480 693576 45496 693610
rect 45554 693576 45570 693610
rect 45638 693576 45654 693610
rect 45712 693576 45728 693610
rect 45796 693576 45812 693610
rect 45870 693576 45886 693610
rect 45954 693576 45970 693610
rect 46028 693576 46044 693610
rect 46112 693576 46128 693610
rect 46186 693576 46202 693610
rect 46270 693576 46286 693610
rect 42980 693517 43014 693533
rect 42980 692525 43014 692541
rect 43138 693517 43172 693533
rect 43138 692525 43172 692541
rect 43296 693517 43330 693533
rect 43296 692525 43330 692541
rect 43454 693517 43488 693533
rect 43454 692525 43488 692541
rect 43612 693517 43646 693533
rect 43612 692525 43646 692541
rect 43770 693517 43804 693533
rect 43770 692525 43804 692541
rect 43928 693517 43962 693533
rect 43928 692525 43962 692541
rect 44086 693517 44120 693533
rect 44086 692525 44120 692541
rect 44244 693517 44278 693533
rect 44244 692525 44278 692541
rect 44402 693517 44436 693533
rect 44402 692525 44436 692541
rect 44560 693517 44594 693533
rect 44560 692525 44594 692541
rect 44718 693517 44752 693533
rect 44718 692525 44752 692541
rect 44876 693517 44910 693533
rect 44876 692525 44910 692541
rect 45034 693517 45068 693533
rect 45034 692525 45068 692541
rect 45192 693517 45226 693533
rect 45192 692525 45226 692541
rect 45350 693517 45384 693533
rect 45350 692525 45384 692541
rect 45508 693517 45542 693533
rect 45508 692525 45542 692541
rect 45666 693517 45700 693533
rect 45666 692525 45700 692541
rect 45824 693517 45858 693533
rect 45824 692525 45858 692541
rect 45982 693517 46016 693533
rect 45982 692525 46016 692541
rect 46140 693517 46174 693533
rect 46140 692525 46174 692541
rect 46298 693517 46332 693533
rect 46298 692525 46332 692541
rect 43026 692448 43042 692482
rect 43110 692448 43126 692482
rect 43184 692448 43200 692482
rect 43268 692448 43284 692482
rect 43342 692448 43358 692482
rect 43426 692448 43442 692482
rect 43500 692448 43516 692482
rect 43584 692448 43600 692482
rect 43658 692448 43674 692482
rect 43742 692448 43758 692482
rect 43816 692448 43832 692482
rect 43900 692448 43916 692482
rect 43974 692448 43990 692482
rect 44058 692448 44074 692482
rect 44132 692448 44148 692482
rect 44216 692448 44232 692482
rect 44290 692448 44306 692482
rect 44374 692448 44390 692482
rect 44448 692448 44464 692482
rect 44532 692448 44548 692482
rect 44606 692448 44622 692482
rect 44690 692448 44706 692482
rect 44764 692448 44780 692482
rect 44848 692448 44864 692482
rect 44922 692448 44938 692482
rect 45006 692448 45022 692482
rect 45080 692448 45096 692482
rect 45164 692448 45180 692482
rect 45238 692448 45254 692482
rect 45322 692448 45338 692482
rect 45396 692448 45412 692482
rect 45480 692448 45496 692482
rect 45554 692448 45570 692482
rect 45638 692448 45654 692482
rect 45712 692448 45728 692482
rect 45796 692448 45812 692482
rect 45870 692448 45886 692482
rect 45954 692448 45970 692482
rect 46028 692448 46044 692482
rect 46112 692448 46128 692482
rect 46186 692448 46202 692482
rect 46270 692448 46286 692482
rect 42866 692380 42900 692442
rect 51723 694703 51757 694765
rect 48633 693427 48667 693489
rect 51723 693427 51757 693489
rect 48633 693393 48729 693427
rect 51661 693393 51757 693427
rect 46412 692380 46446 692442
rect 42866 692346 42962 692380
rect 46350 692346 46446 692380
rect 42866 692138 42962 692172
rect 46350 692138 46446 692172
rect 42866 692076 42900 692138
rect 46412 692076 46446 692138
rect 43026 692036 43042 692070
rect 43110 692036 43126 692070
rect 43184 692036 43200 692070
rect 43268 692036 43284 692070
rect 43342 692036 43358 692070
rect 43426 692036 43442 692070
rect 43500 692036 43516 692070
rect 43584 692036 43600 692070
rect 43658 692036 43674 692070
rect 43742 692036 43758 692070
rect 43816 692036 43832 692070
rect 43900 692036 43916 692070
rect 43974 692036 43990 692070
rect 44058 692036 44074 692070
rect 44132 692036 44148 692070
rect 44216 692036 44232 692070
rect 44290 692036 44306 692070
rect 44374 692036 44390 692070
rect 44448 692036 44464 692070
rect 44532 692036 44548 692070
rect 44606 692036 44622 692070
rect 44690 692036 44706 692070
rect 44764 692036 44780 692070
rect 44848 692036 44864 692070
rect 44922 692036 44938 692070
rect 45006 692036 45022 692070
rect 45080 692036 45096 692070
rect 45164 692036 45180 692070
rect 45238 692036 45254 692070
rect 45322 692036 45338 692070
rect 45396 692036 45412 692070
rect 45480 692036 45496 692070
rect 45554 692036 45570 692070
rect 45638 692036 45654 692070
rect 45712 692036 45728 692070
rect 45796 692036 45812 692070
rect 45870 692036 45886 692070
rect 45954 692036 45970 692070
rect 46028 692036 46044 692070
rect 46112 692036 46128 692070
rect 46186 692036 46202 692070
rect 46270 692036 46286 692070
rect 42980 691977 43014 691993
rect 42980 690985 43014 691001
rect 43138 691977 43172 691993
rect 43138 690985 43172 691001
rect 43296 691977 43330 691993
rect 43296 690985 43330 691001
rect 43454 691977 43488 691993
rect 43454 690985 43488 691001
rect 43612 691977 43646 691993
rect 43612 690985 43646 691001
rect 43770 691977 43804 691993
rect 43770 690985 43804 691001
rect 43928 691977 43962 691993
rect 43928 690985 43962 691001
rect 44086 691977 44120 691993
rect 44086 690985 44120 691001
rect 44244 691977 44278 691993
rect 44244 690985 44278 691001
rect 44402 691977 44436 691993
rect 44402 690985 44436 691001
rect 44560 691977 44594 691993
rect 44560 690985 44594 691001
rect 44718 691977 44752 691993
rect 44718 690985 44752 691001
rect 44876 691977 44910 691993
rect 44876 690985 44910 691001
rect 45034 691977 45068 691993
rect 45034 690985 45068 691001
rect 45192 691977 45226 691993
rect 45192 690985 45226 691001
rect 45350 691977 45384 691993
rect 45350 690985 45384 691001
rect 45508 691977 45542 691993
rect 45508 690985 45542 691001
rect 45666 691977 45700 691993
rect 45666 690985 45700 691001
rect 45824 691977 45858 691993
rect 45824 690985 45858 691001
rect 45982 691977 46016 691993
rect 45982 690985 46016 691001
rect 46140 691977 46174 691993
rect 46140 690985 46174 691001
rect 46298 691977 46332 691993
rect 46298 690985 46332 691001
rect 43026 690908 43042 690942
rect 43110 690908 43126 690942
rect 43184 690908 43200 690942
rect 43268 690908 43284 690942
rect 43342 690908 43358 690942
rect 43426 690908 43442 690942
rect 43500 690908 43516 690942
rect 43584 690908 43600 690942
rect 43658 690908 43674 690942
rect 43742 690908 43758 690942
rect 43816 690908 43832 690942
rect 43900 690908 43916 690942
rect 43974 690908 43990 690942
rect 44058 690908 44074 690942
rect 44132 690908 44148 690942
rect 44216 690908 44232 690942
rect 44290 690908 44306 690942
rect 44374 690908 44390 690942
rect 44448 690908 44464 690942
rect 44532 690908 44548 690942
rect 44606 690908 44622 690942
rect 44690 690908 44706 690942
rect 44764 690908 44780 690942
rect 44848 690908 44864 690942
rect 44922 690908 44938 690942
rect 45006 690908 45022 690942
rect 45080 690908 45096 690942
rect 45164 690908 45180 690942
rect 45238 690908 45254 690942
rect 45322 690908 45338 690942
rect 45396 690908 45412 690942
rect 45480 690908 45496 690942
rect 45554 690908 45570 690942
rect 45638 690908 45654 690942
rect 45712 690908 45728 690942
rect 45796 690908 45812 690942
rect 45870 690908 45886 690942
rect 45954 690908 45970 690942
rect 46028 690908 46044 690942
rect 46112 690908 46128 690942
rect 46186 690908 46202 690942
rect 46270 690908 46286 690942
rect 42866 690840 42900 690902
rect 46412 690840 46446 690902
rect 42866 690806 42962 690840
rect 46350 690806 46446 690840
rect 540185 690864 540281 690898
rect 548871 690864 548967 690898
rect 540185 690802 540219 690864
rect 43967 690561 44063 690595
rect 45239 690561 45335 690595
rect 43967 690499 44001 690561
rect 45301 690499 45335 690561
rect 44127 690459 44143 690493
rect 44211 690459 44227 690493
rect 44285 690459 44301 690493
rect 44369 690459 44385 690493
rect 44443 690459 44459 690493
rect 44527 690459 44543 690493
rect 44601 690459 44617 690493
rect 44685 690459 44701 690493
rect 44759 690459 44775 690493
rect 44843 690459 44859 690493
rect 44917 690459 44933 690493
rect 45001 690459 45017 690493
rect 45075 690459 45091 690493
rect 45159 690459 45175 690493
rect 44081 690409 44115 690425
rect 44081 689417 44115 689433
rect 44239 690409 44273 690425
rect 44239 689417 44273 689433
rect 44397 690409 44431 690425
rect 44397 689417 44431 689433
rect 44555 690409 44589 690425
rect 44555 689417 44589 689433
rect 44713 690409 44747 690425
rect 44713 689417 44747 689433
rect 44871 690409 44905 690425
rect 44871 689417 44905 689433
rect 45029 690409 45063 690425
rect 45029 689417 45063 689433
rect 45187 690409 45221 690425
rect 45187 689417 45221 689433
rect 44127 689349 44143 689383
rect 44211 689349 44227 689383
rect 44285 689349 44301 689383
rect 44369 689349 44385 689383
rect 44443 689349 44459 689383
rect 44527 689349 44543 689383
rect 44601 689349 44617 689383
rect 44685 689349 44701 689383
rect 44759 689349 44775 689383
rect 44843 689349 44859 689383
rect 44917 689349 44933 689383
rect 45001 689349 45017 689383
rect 45075 689349 45091 689383
rect 45159 689349 45175 689383
rect 43967 689281 44001 689343
rect 548933 690802 548967 690864
rect 540364 690750 540380 690784
rect 541356 690750 541372 690784
rect 541600 690750 541616 690784
rect 542592 690750 542608 690784
rect 542836 690750 542852 690784
rect 543828 690750 543844 690784
rect 544072 690750 544088 690784
rect 545064 690750 545080 690784
rect 545308 690750 545324 690784
rect 546300 690750 546316 690784
rect 546544 690750 546560 690784
rect 547536 690750 547552 690784
rect 547780 690750 547796 690784
rect 548772 690750 548788 690784
rect 540287 690722 540321 690738
rect 540287 690638 540321 690654
rect 541415 690722 541449 690738
rect 541415 690638 541449 690654
rect 541523 690722 541557 690738
rect 541523 690638 541557 690654
rect 542651 690722 542685 690738
rect 542651 690638 542685 690654
rect 542759 690722 542793 690738
rect 542759 690638 542793 690654
rect 543887 690722 543921 690738
rect 543887 690638 543921 690654
rect 543995 690722 544029 690738
rect 543995 690638 544029 690654
rect 545123 690722 545157 690738
rect 545123 690638 545157 690654
rect 545231 690722 545265 690738
rect 545231 690638 545265 690654
rect 546359 690722 546393 690738
rect 546359 690638 546393 690654
rect 546467 690722 546501 690738
rect 546467 690638 546501 690654
rect 547595 690722 547629 690738
rect 547595 690638 547629 690654
rect 547703 690722 547737 690738
rect 547703 690638 547737 690654
rect 548831 690722 548865 690738
rect 548831 690638 548865 690654
rect 540364 690592 540380 690626
rect 541356 690592 541372 690626
rect 541600 690592 541616 690626
rect 542592 690592 542608 690626
rect 542836 690592 542852 690626
rect 543828 690592 543844 690626
rect 544072 690592 544088 690626
rect 545064 690592 545080 690626
rect 545308 690592 545324 690626
rect 546300 690592 546316 690626
rect 546544 690592 546560 690626
rect 547536 690592 547552 690626
rect 547780 690592 547796 690626
rect 548772 690592 548788 690626
rect 540185 690512 540219 690574
rect 548933 690512 548967 690574
rect 540185 690478 540281 690512
rect 548871 690478 548967 690512
rect 540185 690324 540281 690358
rect 548871 690324 548967 690358
rect 540185 690262 540219 690324
rect 548933 690262 548967 690324
rect 540364 690210 540380 690244
rect 541356 690210 541372 690244
rect 541600 690210 541616 690244
rect 542592 690210 542608 690244
rect 542836 690210 542852 690244
rect 543828 690210 543844 690244
rect 544072 690210 544088 690244
rect 545064 690210 545080 690244
rect 545308 690210 545324 690244
rect 546300 690210 546316 690244
rect 546544 690210 546560 690244
rect 547536 690210 547552 690244
rect 547780 690210 547796 690244
rect 548772 690210 548788 690244
rect 540287 690182 540321 690198
rect 540287 690098 540321 690114
rect 541415 690182 541449 690198
rect 541415 690098 541449 690114
rect 541523 690182 541557 690198
rect 541523 690098 541557 690114
rect 542651 690182 542685 690198
rect 542651 690098 542685 690114
rect 542759 690182 542793 690198
rect 542759 690098 542793 690114
rect 543887 690182 543921 690198
rect 543887 690098 543921 690114
rect 543995 690182 544029 690198
rect 543995 690098 544029 690114
rect 545123 690182 545157 690198
rect 545123 690098 545157 690114
rect 545231 690182 545265 690198
rect 545231 690098 545265 690114
rect 546359 690182 546393 690198
rect 546359 690098 546393 690114
rect 546467 690182 546501 690198
rect 546467 690098 546501 690114
rect 547595 690182 547629 690198
rect 547595 690098 547629 690114
rect 547703 690182 547737 690198
rect 547703 690098 547737 690114
rect 548831 690182 548865 690198
rect 548831 690098 548865 690114
rect 540364 690052 540380 690086
rect 541356 690052 541372 690086
rect 541600 690052 541616 690086
rect 542592 690052 542608 690086
rect 542836 690052 542852 690086
rect 543828 690052 543844 690086
rect 544072 690052 544088 690086
rect 545064 690052 545080 690086
rect 545308 690052 545324 690086
rect 546300 690052 546316 690086
rect 546544 690052 546560 690086
rect 547536 690052 547552 690086
rect 547780 690052 547796 690086
rect 548772 690052 548788 690086
rect 540185 689972 540219 690034
rect 548933 689972 548967 690034
rect 540185 689938 540281 689972
rect 548871 689938 548967 689972
rect 541969 689912 542229 689938
rect 541969 689842 541979 689912
rect 542069 689842 542119 689912
rect 542209 689842 542229 689912
rect 541969 689818 542229 689842
rect 544439 689922 544729 689938
rect 544439 689912 544619 689922
rect 544439 689842 544459 689912
rect 544549 689852 544619 689912
rect 544709 689852 544729 689922
rect 544549 689842 544729 689852
rect 544439 689818 544729 689842
rect 546899 689922 547189 689938
rect 546899 689852 546919 689922
rect 546999 689852 547089 689922
rect 547169 689852 547189 689922
rect 546899 689818 547189 689852
rect 540185 689784 540281 689818
rect 548871 689784 548967 689818
rect 540185 689722 540219 689784
rect 548933 689722 548967 689784
rect 540364 689670 540380 689704
rect 541356 689670 541372 689704
rect 541600 689670 541616 689704
rect 542592 689670 542608 689704
rect 542836 689670 542852 689704
rect 543828 689670 543844 689704
rect 544072 689670 544088 689704
rect 545064 689670 545080 689704
rect 545308 689670 545324 689704
rect 546300 689670 546316 689704
rect 546544 689670 546560 689704
rect 547536 689670 547552 689704
rect 547780 689670 547796 689704
rect 548772 689670 548788 689704
rect 540287 689642 540321 689658
rect 540287 689558 540321 689574
rect 541415 689642 541449 689658
rect 541415 689558 541449 689574
rect 541523 689642 541557 689658
rect 541523 689558 541557 689574
rect 542651 689642 542685 689658
rect 542651 689558 542685 689574
rect 542759 689642 542793 689658
rect 542759 689558 542793 689574
rect 543887 689642 543921 689658
rect 543887 689558 543921 689574
rect 543995 689642 544029 689658
rect 543995 689558 544029 689574
rect 545123 689642 545157 689658
rect 545123 689558 545157 689574
rect 545231 689642 545265 689658
rect 545231 689558 545265 689574
rect 546359 689642 546393 689658
rect 546359 689558 546393 689574
rect 546467 689642 546501 689658
rect 546467 689558 546501 689574
rect 547595 689642 547629 689658
rect 547595 689558 547629 689574
rect 547703 689642 547737 689658
rect 547703 689558 547737 689574
rect 548831 689642 548865 689658
rect 548831 689558 548865 689574
rect 540364 689512 540380 689546
rect 541356 689512 541372 689546
rect 541600 689512 541616 689546
rect 542592 689512 542608 689546
rect 542836 689512 542852 689546
rect 543828 689512 543844 689546
rect 544072 689512 544088 689546
rect 545064 689512 545080 689546
rect 545308 689512 545324 689546
rect 546300 689512 546316 689546
rect 546544 689512 546560 689546
rect 547536 689512 547552 689546
rect 547780 689512 547796 689546
rect 548772 689512 548788 689546
rect 540185 689432 540219 689494
rect 548933 689432 548967 689494
rect 540185 689398 540281 689432
rect 548871 689398 548967 689432
rect 45301 689281 45335 689343
rect 43967 689247 44063 689281
rect 45239 689247 45335 689281
rect 541959 689382 542249 689398
rect 541959 689302 541979 689382
rect 542059 689302 542149 689382
rect 542229 689302 542249 689382
rect 541959 689278 542249 689302
rect 544439 689382 544729 689398
rect 544439 689302 544459 689382
rect 544539 689302 544629 689382
rect 544709 689302 544729 689382
rect 544439 689278 544729 689302
rect 546899 689382 547189 689398
rect 546899 689302 546919 689382
rect 546999 689302 547089 689382
rect 547169 689302 547189 689382
rect 546899 689278 547189 689302
rect 540185 689244 540281 689278
rect 548871 689244 548967 689278
rect 540185 689182 540219 689244
rect 43967 689041 44063 689075
rect 45239 689041 45335 689075
rect 43967 688979 44001 689041
rect 45301 688979 45335 689041
rect 44127 688939 44143 688973
rect 44211 688939 44227 688973
rect 44285 688939 44301 688973
rect 44369 688939 44385 688973
rect 44443 688939 44459 688973
rect 44527 688939 44543 688973
rect 44601 688939 44617 688973
rect 44685 688939 44701 688973
rect 44759 688939 44775 688973
rect 44843 688939 44859 688973
rect 44917 688939 44933 688973
rect 45001 688939 45017 688973
rect 45075 688939 45091 688973
rect 45159 688939 45175 688973
rect 44081 688889 44115 688905
rect 44081 687897 44115 687913
rect 44239 688889 44273 688905
rect 44239 687897 44273 687913
rect 44397 688889 44431 688905
rect 44397 687897 44431 687913
rect 44555 688889 44589 688905
rect 44555 687897 44589 687913
rect 44713 688889 44747 688905
rect 44713 687897 44747 687913
rect 44871 688889 44905 688905
rect 44871 687897 44905 687913
rect 45029 688889 45063 688905
rect 45029 687897 45063 687913
rect 45187 688889 45221 688905
rect 45187 687897 45221 687913
rect 44127 687829 44143 687863
rect 44211 687829 44227 687863
rect 44285 687829 44301 687863
rect 44369 687829 44385 687863
rect 44443 687829 44459 687863
rect 44527 687829 44543 687863
rect 44601 687829 44617 687863
rect 44685 687829 44701 687863
rect 44759 687829 44775 687863
rect 44843 687829 44859 687863
rect 44917 687829 44933 687863
rect 45001 687829 45017 687863
rect 45075 687829 45091 687863
rect 45159 687829 45175 687863
rect 43967 687761 44001 687823
rect 548933 689182 548967 689244
rect 540364 689130 540380 689164
rect 541356 689130 541372 689164
rect 541600 689130 541616 689164
rect 542592 689130 542608 689164
rect 542836 689130 542852 689164
rect 543828 689130 543844 689164
rect 544072 689130 544088 689164
rect 545064 689130 545080 689164
rect 545308 689130 545324 689164
rect 546300 689130 546316 689164
rect 546544 689130 546560 689164
rect 547536 689130 547552 689164
rect 547780 689130 547796 689164
rect 548772 689130 548788 689164
rect 540287 689102 540321 689118
rect 540287 689018 540321 689034
rect 541415 689102 541449 689118
rect 541415 689018 541449 689034
rect 541523 689102 541557 689118
rect 541523 689018 541557 689034
rect 542651 689102 542685 689118
rect 542651 689018 542685 689034
rect 542759 689102 542793 689118
rect 542759 689018 542793 689034
rect 543887 689102 543921 689118
rect 543887 689018 543921 689034
rect 543995 689102 544029 689118
rect 543995 689018 544029 689034
rect 545123 689102 545157 689118
rect 545123 689018 545157 689034
rect 545231 689102 545265 689118
rect 545231 689018 545265 689034
rect 546359 689102 546393 689118
rect 546359 689018 546393 689034
rect 546467 689102 546501 689118
rect 546467 689018 546501 689034
rect 547595 689102 547629 689118
rect 547595 689018 547629 689034
rect 547703 689102 547737 689118
rect 547703 689018 547737 689034
rect 548831 689102 548865 689118
rect 548831 689018 548865 689034
rect 540364 688972 540380 689006
rect 541356 688972 541372 689006
rect 541600 688972 541616 689006
rect 542592 688972 542608 689006
rect 542836 688972 542852 689006
rect 543828 688972 543844 689006
rect 544072 688972 544088 689006
rect 545064 688972 545080 689006
rect 545308 688972 545324 689006
rect 546300 688972 546316 689006
rect 546544 688972 546560 689006
rect 547536 688972 547552 689006
rect 547780 688972 547796 689006
rect 548772 688972 548788 689006
rect 540185 688892 540219 688954
rect 548933 688892 548967 688954
rect 540185 688858 540281 688892
rect 548871 688858 548967 688892
rect 540185 688664 540281 688698
rect 548871 688664 548967 688698
rect 540185 688602 540219 688664
rect 548933 688602 548967 688664
rect 540364 688550 540380 688584
rect 541356 688550 541372 688584
rect 541600 688550 541616 688584
rect 542592 688550 542608 688584
rect 542836 688550 542852 688584
rect 543828 688550 543844 688584
rect 544072 688550 544088 688584
rect 545064 688550 545080 688584
rect 545308 688550 545324 688584
rect 546300 688550 546316 688584
rect 546544 688550 546560 688584
rect 547536 688550 547552 688584
rect 547780 688550 547796 688584
rect 548772 688550 548788 688584
rect 540287 688522 540321 688538
rect 540287 688438 540321 688454
rect 541415 688522 541449 688538
rect 541415 688438 541449 688454
rect 541523 688522 541557 688538
rect 541523 688438 541557 688454
rect 542651 688522 542685 688538
rect 542651 688438 542685 688454
rect 542759 688522 542793 688538
rect 542759 688438 542793 688454
rect 543887 688522 543921 688538
rect 543887 688438 543921 688454
rect 543995 688522 544029 688538
rect 543995 688438 544029 688454
rect 545123 688522 545157 688538
rect 545123 688438 545157 688454
rect 545231 688522 545265 688538
rect 545231 688438 545265 688454
rect 546359 688522 546393 688538
rect 546359 688438 546393 688454
rect 546467 688522 546501 688538
rect 546467 688438 546501 688454
rect 547595 688522 547629 688538
rect 547595 688438 547629 688454
rect 547703 688522 547737 688538
rect 547703 688438 547737 688454
rect 548831 688522 548865 688538
rect 548831 688438 548865 688454
rect 540364 688392 540380 688426
rect 541356 688392 541372 688426
rect 541600 688392 541616 688426
rect 542592 688392 542608 688426
rect 542836 688392 542852 688426
rect 543828 688392 543844 688426
rect 544072 688392 544088 688426
rect 545064 688392 545080 688426
rect 545308 688392 545324 688426
rect 546300 688392 546316 688426
rect 546544 688392 546560 688426
rect 547536 688392 547552 688426
rect 547780 688392 547796 688426
rect 548772 688392 548788 688426
rect 540185 688312 540219 688374
rect 548933 688312 548967 688374
rect 540185 688278 540281 688312
rect 548871 688278 548967 688312
rect 541959 688222 542249 688278
rect 541959 688142 541979 688222
rect 542069 688142 542139 688222
rect 542229 688142 542249 688222
rect 541959 688118 542249 688142
rect 544439 688212 544729 688278
rect 544439 688142 544459 688212
rect 544539 688142 544629 688212
rect 544709 688142 544729 688212
rect 544439 688118 544729 688142
rect 546899 688212 547189 688278
rect 546899 688142 546919 688212
rect 546999 688142 547089 688212
rect 547169 688142 547189 688212
rect 546899 688118 547189 688142
rect 45301 687761 45335 687823
rect 43967 687727 44063 687761
rect 45239 687727 45335 687761
rect 534592 688067 534688 688101
rect 537620 688067 537716 688101
rect 534592 688005 534626 688067
rect 42976 687520 43072 687554
rect 46238 687520 46334 687554
rect 42976 687458 43010 687520
rect 46300 687458 46334 687520
rect 43136 687418 43152 687452
rect 43320 687418 43336 687452
rect 43394 687418 43410 687452
rect 43578 687418 43594 687452
rect 43652 687418 43668 687452
rect 43836 687418 43852 687452
rect 43910 687418 43926 687452
rect 44094 687418 44110 687452
rect 44168 687418 44184 687452
rect 44352 687418 44368 687452
rect 44426 687418 44442 687452
rect 44610 687418 44626 687452
rect 44684 687418 44700 687452
rect 44868 687418 44884 687452
rect 44942 687418 44958 687452
rect 45126 687418 45142 687452
rect 45200 687418 45216 687452
rect 45384 687418 45400 687452
rect 45458 687418 45474 687452
rect 45642 687418 45658 687452
rect 45716 687418 45732 687452
rect 45900 687418 45916 687452
rect 45974 687418 45990 687452
rect 46158 687418 46174 687452
rect 43090 687368 43124 687384
rect 43090 686376 43124 686392
rect 43348 687368 43382 687384
rect 43348 686376 43382 686392
rect 43606 687368 43640 687384
rect 43606 686376 43640 686392
rect 43864 687368 43898 687384
rect 43864 686376 43898 686392
rect 44122 687368 44156 687384
rect 44122 686376 44156 686392
rect 44380 687368 44414 687384
rect 44380 686376 44414 686392
rect 44638 687368 44672 687384
rect 44638 686376 44672 686392
rect 44896 687368 44930 687384
rect 44896 686376 44930 686392
rect 45154 687368 45188 687384
rect 45154 686376 45188 686392
rect 45412 687368 45446 687384
rect 45412 686376 45446 686392
rect 45670 687368 45704 687384
rect 45670 686376 45704 686392
rect 45928 687368 45962 687384
rect 45928 686376 45962 686392
rect 46186 687368 46220 687384
rect 46186 686376 46220 686392
rect 43136 686308 43152 686342
rect 43320 686308 43336 686342
rect 43394 686308 43410 686342
rect 43578 686308 43594 686342
rect 43652 686308 43668 686342
rect 43836 686308 43852 686342
rect 43910 686308 43926 686342
rect 44094 686308 44110 686342
rect 44168 686308 44184 686342
rect 44352 686308 44368 686342
rect 44426 686308 44442 686342
rect 44610 686308 44626 686342
rect 44684 686308 44700 686342
rect 44868 686308 44884 686342
rect 44942 686308 44958 686342
rect 45126 686308 45142 686342
rect 45200 686308 45216 686342
rect 45384 686308 45400 686342
rect 45458 686308 45474 686342
rect 45642 686308 45658 686342
rect 45716 686308 45732 686342
rect 45900 686308 45916 686342
rect 45974 686308 45990 686342
rect 46158 686308 46174 686342
rect 42976 686240 43010 686302
rect 537682 688005 537716 688067
rect 534592 686729 534626 686791
rect 540185 688084 540281 688118
rect 548871 688084 548967 688118
rect 540185 688022 540219 688084
rect 548933 688022 548967 688084
rect 540364 687970 540380 688004
rect 541356 687970 541372 688004
rect 541600 687970 541616 688004
rect 542592 687970 542608 688004
rect 542836 687970 542852 688004
rect 543828 687970 543844 688004
rect 544072 687970 544088 688004
rect 545064 687970 545080 688004
rect 545308 687970 545324 688004
rect 546300 687970 546316 688004
rect 546544 687970 546560 688004
rect 547536 687970 547552 688004
rect 547780 687970 547796 688004
rect 548772 687970 548788 688004
rect 540287 687942 540321 687958
rect 540287 687858 540321 687874
rect 541415 687942 541449 687958
rect 541415 687858 541449 687874
rect 541523 687942 541557 687958
rect 541523 687858 541557 687874
rect 542651 687942 542685 687958
rect 542651 687858 542685 687874
rect 542759 687942 542793 687958
rect 542759 687858 542793 687874
rect 543887 687942 543921 687958
rect 543887 687858 543921 687874
rect 543995 687942 544029 687958
rect 543995 687858 544029 687874
rect 545123 687942 545157 687958
rect 545123 687858 545157 687874
rect 545231 687942 545265 687958
rect 545231 687858 545265 687874
rect 546359 687942 546393 687958
rect 546359 687858 546393 687874
rect 546467 687942 546501 687958
rect 546467 687858 546501 687874
rect 547595 687942 547629 687958
rect 547595 687858 547629 687874
rect 547703 687942 547737 687958
rect 547703 687858 547737 687874
rect 548831 687942 548865 687958
rect 548831 687858 548865 687874
rect 540364 687812 540380 687846
rect 541356 687812 541372 687846
rect 541600 687812 541616 687846
rect 542592 687812 542608 687846
rect 542836 687812 542852 687846
rect 543828 687812 543844 687846
rect 544072 687812 544088 687846
rect 545064 687812 545080 687846
rect 545308 687812 545324 687846
rect 546300 687812 546316 687846
rect 546544 687812 546560 687846
rect 547536 687812 547552 687846
rect 547780 687812 547796 687846
rect 548772 687812 548788 687846
rect 540185 687732 540219 687794
rect 548933 687732 548967 687794
rect 540185 687698 540281 687732
rect 548871 687698 548967 687732
rect 551652 688067 551748 688101
rect 554680 688067 554776 688101
rect 551652 688005 551686 688067
rect 538345 687544 538441 687578
rect 550739 687544 550835 687578
rect 538345 687482 538379 687544
rect 550801 687482 550835 687544
rect 538524 687430 538540 687464
rect 539516 687430 539532 687464
rect 539760 687430 539776 687464
rect 540752 687430 540768 687464
rect 540996 687430 541012 687464
rect 541988 687430 542004 687464
rect 542232 687430 542248 687464
rect 543224 687430 543240 687464
rect 543468 687430 543484 687464
rect 544460 687430 544476 687464
rect 544704 687430 544720 687464
rect 545696 687430 545712 687464
rect 545940 687430 545956 687464
rect 546932 687430 546948 687464
rect 547176 687430 547192 687464
rect 548168 687430 548184 687464
rect 548412 687430 548428 687464
rect 549404 687430 549420 687464
rect 549648 687430 549664 687464
rect 550640 687430 550656 687464
rect 538447 687402 538481 687418
rect 538447 687318 538481 687334
rect 539575 687402 539609 687418
rect 539575 687318 539609 687334
rect 539683 687402 539717 687418
rect 539683 687318 539717 687334
rect 540811 687402 540845 687418
rect 540811 687318 540845 687334
rect 540919 687402 540953 687418
rect 540919 687318 540953 687334
rect 542047 687402 542081 687418
rect 542047 687318 542081 687334
rect 542155 687402 542189 687418
rect 542155 687318 542189 687334
rect 543283 687402 543317 687418
rect 543283 687318 543317 687334
rect 543391 687402 543425 687418
rect 543391 687318 543425 687334
rect 544519 687402 544553 687418
rect 544519 687318 544553 687334
rect 544627 687402 544661 687418
rect 544627 687318 544661 687334
rect 545755 687402 545789 687418
rect 545755 687318 545789 687334
rect 545863 687402 545897 687418
rect 545863 687318 545897 687334
rect 546991 687402 547025 687418
rect 546991 687318 547025 687334
rect 547099 687402 547133 687418
rect 547099 687318 547133 687334
rect 548227 687402 548261 687418
rect 548227 687318 548261 687334
rect 548335 687402 548369 687418
rect 548335 687318 548369 687334
rect 549463 687402 549497 687418
rect 549463 687318 549497 687334
rect 549571 687402 549605 687418
rect 549571 687318 549605 687334
rect 550699 687402 550733 687418
rect 550699 687318 550733 687334
rect 538524 687272 538540 687306
rect 539516 687272 539532 687306
rect 539760 687272 539776 687306
rect 540752 687272 540768 687306
rect 540996 687272 541012 687306
rect 541988 687272 542004 687306
rect 542232 687272 542248 687306
rect 543224 687272 543240 687306
rect 543468 687272 543484 687306
rect 544460 687272 544476 687306
rect 544704 687272 544720 687306
rect 545696 687272 545712 687306
rect 545940 687272 545956 687306
rect 546932 687272 546948 687306
rect 547176 687272 547192 687306
rect 548168 687272 548184 687306
rect 548412 687272 548428 687306
rect 549404 687272 549420 687306
rect 549648 687272 549664 687306
rect 550640 687272 550656 687306
rect 538345 687192 538379 687254
rect 550801 687192 550835 687254
rect 538345 687158 538441 687192
rect 550739 687158 550835 687192
rect 540099 687142 540409 687158
rect 540099 687062 540119 687142
rect 540209 687062 540299 687142
rect 540389 687062 540409 687142
rect 540099 687038 540409 687062
rect 542629 687142 542919 687158
rect 542629 687062 542649 687142
rect 542739 687062 542809 687142
rect 542899 687062 542919 687142
rect 542629 687038 542919 687062
rect 545099 687142 545389 687158
rect 545099 687062 545119 687142
rect 545209 687062 545279 687142
rect 545369 687062 545389 687142
rect 545099 687038 545389 687062
rect 547549 687142 547839 687158
rect 547549 687062 547569 687142
rect 547659 687062 547729 687142
rect 547819 687062 547839 687142
rect 547549 687038 547839 687062
rect 550049 687142 550339 687158
rect 550049 687062 550069 687142
rect 550159 687062 550229 687142
rect 550319 687062 550339 687142
rect 550049 687038 550339 687062
rect 535779 686729 535869 686742
rect 537682 686729 537716 686791
rect 534592 686695 534688 686729
rect 537620 686695 537716 686729
rect 538345 687004 538441 687038
rect 550739 687004 550835 687038
rect 538345 686942 538379 687004
rect 550801 686942 550835 687004
rect 538524 686890 538540 686924
rect 539516 686890 539532 686924
rect 539760 686890 539776 686924
rect 540752 686890 540768 686924
rect 540996 686890 541012 686924
rect 541988 686890 542004 686924
rect 542232 686890 542248 686924
rect 543224 686890 543240 686924
rect 543468 686890 543484 686924
rect 544460 686890 544476 686924
rect 544704 686890 544720 686924
rect 545696 686890 545712 686924
rect 545940 686890 545956 686924
rect 546932 686890 546948 686924
rect 547176 686890 547192 686924
rect 548168 686890 548184 686924
rect 548412 686890 548428 686924
rect 549404 686890 549420 686924
rect 549648 686890 549664 686924
rect 550640 686890 550656 686924
rect 538447 686862 538481 686878
rect 538447 686778 538481 686794
rect 539575 686862 539609 686878
rect 539575 686778 539609 686794
rect 539683 686862 539717 686878
rect 539683 686778 539717 686794
rect 540811 686862 540845 686878
rect 540811 686778 540845 686794
rect 540919 686862 540953 686878
rect 540919 686778 540953 686794
rect 542047 686862 542081 686878
rect 542047 686778 542081 686794
rect 542155 686862 542189 686878
rect 542155 686778 542189 686794
rect 543283 686862 543317 686878
rect 543283 686778 543317 686794
rect 543391 686862 543425 686878
rect 543391 686778 543425 686794
rect 544519 686862 544553 686878
rect 544519 686778 544553 686794
rect 544627 686862 544661 686878
rect 544627 686778 544661 686794
rect 545755 686862 545789 686878
rect 545755 686778 545789 686794
rect 545863 686862 545897 686878
rect 545863 686778 545897 686794
rect 546991 686862 547025 686878
rect 546991 686778 547025 686794
rect 547099 686862 547133 686878
rect 547099 686778 547133 686794
rect 548227 686862 548261 686878
rect 548227 686778 548261 686794
rect 548335 686862 548369 686878
rect 548335 686778 548369 686794
rect 549463 686862 549497 686878
rect 549463 686778 549497 686794
rect 549571 686862 549605 686878
rect 549571 686778 549605 686794
rect 550699 686862 550733 686878
rect 550699 686778 550733 686794
rect 538524 686732 538540 686766
rect 539516 686732 539532 686766
rect 539760 686732 539776 686766
rect 540752 686732 540768 686766
rect 540996 686732 541012 686766
rect 541988 686732 542004 686766
rect 542232 686732 542248 686766
rect 543224 686732 543240 686766
rect 543468 686732 543484 686766
rect 544460 686732 544476 686766
rect 544704 686732 544720 686766
rect 545696 686732 545712 686766
rect 545940 686732 545956 686766
rect 546932 686732 546948 686766
rect 547176 686732 547192 686766
rect 548168 686732 548184 686766
rect 548412 686732 548428 686766
rect 549404 686732 549420 686766
rect 549648 686732 549664 686766
rect 550640 686732 550656 686766
rect 535779 686631 535869 686695
rect 538345 686652 538379 686714
rect 550801 686652 550835 686714
rect 554742 688005 554776 688067
rect 551652 686729 551686 686791
rect 554742 686729 554776 686791
rect 551652 686695 551748 686729
rect 554680 686695 554776 686729
rect 46300 686240 46334 686302
rect 42976 686206 43072 686240
rect 46238 686206 46334 686240
rect 534592 686597 534688 686631
rect 537620 686597 537716 686631
rect 538345 686618 538441 686652
rect 550739 686618 550835 686652
rect 553029 686631 553169 686695
rect 534592 686535 534626 686597
rect 42716 686000 42812 686034
rect 46494 686000 46590 686034
rect 42716 685938 42750 686000
rect 46556 685938 46590 686000
rect 42876 685898 42892 685932
rect 43060 685898 43076 685932
rect 43134 685898 43150 685932
rect 43318 685898 43334 685932
rect 43392 685898 43408 685932
rect 43576 685898 43592 685932
rect 43650 685898 43666 685932
rect 43834 685898 43850 685932
rect 43908 685898 43924 685932
rect 44092 685898 44108 685932
rect 44166 685898 44182 685932
rect 44350 685898 44366 685932
rect 44424 685898 44440 685932
rect 44608 685898 44624 685932
rect 44682 685898 44698 685932
rect 44866 685898 44882 685932
rect 44940 685898 44956 685932
rect 45124 685898 45140 685932
rect 45198 685898 45214 685932
rect 45382 685898 45398 685932
rect 45456 685898 45472 685932
rect 45640 685898 45656 685932
rect 45714 685898 45730 685932
rect 45898 685898 45914 685932
rect 45972 685898 45988 685932
rect 46156 685898 46172 685932
rect 46230 685898 46246 685932
rect 46414 685898 46430 685932
rect 42830 685848 42864 685864
rect 42830 684856 42864 684872
rect 43088 685848 43122 685864
rect 43088 684856 43122 684872
rect 43346 685848 43380 685864
rect 43346 684856 43380 684872
rect 43604 685848 43638 685864
rect 43604 684856 43638 684872
rect 43862 685848 43896 685864
rect 43862 684856 43896 684872
rect 44120 685848 44154 685864
rect 44120 684856 44154 684872
rect 44378 685848 44412 685864
rect 44378 684856 44412 684872
rect 44636 685848 44670 685864
rect 44636 684856 44670 684872
rect 44894 685848 44928 685864
rect 44894 684856 44928 684872
rect 45152 685848 45186 685864
rect 45152 684856 45186 684872
rect 45410 685848 45444 685864
rect 45410 684856 45444 684872
rect 45668 685848 45702 685864
rect 45668 684856 45702 684872
rect 45926 685848 45960 685864
rect 45926 684856 45960 684872
rect 46184 685848 46218 685864
rect 46184 684856 46218 684872
rect 46442 685848 46476 685864
rect 46442 684856 46476 684872
rect 42876 684788 42892 684822
rect 43060 684788 43076 684822
rect 43134 684788 43150 684822
rect 43318 684788 43334 684822
rect 43392 684788 43408 684822
rect 43576 684788 43592 684822
rect 43650 684788 43666 684822
rect 43834 684788 43850 684822
rect 43908 684788 43924 684822
rect 44092 684788 44108 684822
rect 44166 684788 44182 684822
rect 44350 684788 44366 684822
rect 44424 684788 44440 684822
rect 44608 684788 44624 684822
rect 44682 684788 44698 684822
rect 44866 684788 44882 684822
rect 44940 684788 44956 684822
rect 45124 684788 45140 684822
rect 45198 684788 45214 684822
rect 45382 684788 45398 684822
rect 45456 684788 45472 684822
rect 45640 684788 45656 684822
rect 45714 684788 45730 684822
rect 45898 684788 45914 684822
rect 45972 684788 45988 684822
rect 46156 684788 46172 684822
rect 46230 684788 46246 684822
rect 46414 684788 46430 684822
rect 42716 684720 42750 684782
rect 537682 686535 537716 686597
rect 534592 685259 534626 685321
rect 551652 686597 551748 686631
rect 554680 686597 554776 686631
rect 551652 686535 551686 686597
rect 538345 686464 538441 686498
rect 550739 686464 550835 686498
rect 538345 686402 538379 686464
rect 550801 686402 550835 686464
rect 538524 686350 538540 686384
rect 539516 686350 539532 686384
rect 539760 686350 539776 686384
rect 540752 686350 540768 686384
rect 540996 686350 541012 686384
rect 541988 686350 542004 686384
rect 542232 686350 542248 686384
rect 543224 686350 543240 686384
rect 543468 686350 543484 686384
rect 544460 686350 544476 686384
rect 544704 686350 544720 686384
rect 545696 686350 545712 686384
rect 545940 686350 545956 686384
rect 546932 686350 546948 686384
rect 547176 686350 547192 686384
rect 548168 686350 548184 686384
rect 548412 686350 548428 686384
rect 549404 686350 549420 686384
rect 549648 686350 549664 686384
rect 550640 686350 550656 686384
rect 538447 686322 538481 686338
rect 538447 686238 538481 686254
rect 539575 686322 539609 686338
rect 539575 686238 539609 686254
rect 539683 686322 539717 686338
rect 539683 686238 539717 686254
rect 540811 686322 540845 686338
rect 540811 686238 540845 686254
rect 540919 686322 540953 686338
rect 540919 686238 540953 686254
rect 542047 686322 542081 686338
rect 542047 686238 542081 686254
rect 542155 686322 542189 686338
rect 542155 686238 542189 686254
rect 543283 686322 543317 686338
rect 543283 686238 543317 686254
rect 543391 686322 543425 686338
rect 543391 686238 543425 686254
rect 544519 686322 544553 686338
rect 544519 686238 544553 686254
rect 544627 686322 544661 686338
rect 544627 686238 544661 686254
rect 545755 686322 545789 686338
rect 545755 686238 545789 686254
rect 545863 686322 545897 686338
rect 545863 686238 545897 686254
rect 546991 686322 547025 686338
rect 546991 686238 547025 686254
rect 547099 686322 547133 686338
rect 547099 686238 547133 686254
rect 548227 686322 548261 686338
rect 548227 686238 548261 686254
rect 548335 686322 548369 686338
rect 548335 686238 548369 686254
rect 549463 686322 549497 686338
rect 549463 686238 549497 686254
rect 549571 686322 549605 686338
rect 549571 686238 549605 686254
rect 550699 686322 550733 686338
rect 550699 686238 550733 686254
rect 538524 686192 538540 686226
rect 539516 686192 539532 686226
rect 539760 686192 539776 686226
rect 540752 686192 540768 686226
rect 540996 686192 541012 686226
rect 541988 686192 542004 686226
rect 542232 686192 542248 686226
rect 543224 686192 543240 686226
rect 543468 686192 543484 686226
rect 544460 686192 544476 686226
rect 544704 686192 544720 686226
rect 545696 686192 545712 686226
rect 545940 686192 545956 686226
rect 546932 686192 546948 686226
rect 547176 686192 547192 686226
rect 548168 686192 548184 686226
rect 548412 686192 548428 686226
rect 549404 686192 549420 686226
rect 549648 686192 549664 686226
rect 550640 686192 550656 686226
rect 538345 686112 538379 686174
rect 550801 686112 550835 686174
rect 538345 686078 538441 686112
rect 550739 686078 550835 686112
rect 540099 686072 540409 686078
rect 540099 686062 540299 686072
rect 540099 685982 540119 686062
rect 540209 685992 540299 686062
rect 540389 685992 540409 686072
rect 540209 685982 540409 685992
rect 540099 685958 540409 685982
rect 542629 686062 542919 686078
rect 542629 685982 542649 686062
rect 542739 685982 542809 686062
rect 542899 685982 542919 686062
rect 542629 685958 542919 685982
rect 545099 686062 545389 686078
rect 545099 685982 545119 686062
rect 545209 685982 545279 686062
rect 545369 685982 545389 686062
rect 545099 685958 545389 685982
rect 547549 686062 547839 686078
rect 547549 685982 547569 686062
rect 547659 685982 547729 686062
rect 547819 685982 547839 686062
rect 547549 685958 547839 685982
rect 550049 686062 550339 686078
rect 550049 685982 550069 686062
rect 550159 685982 550229 686062
rect 550319 685982 550339 686062
rect 550049 685958 550339 685982
rect 538345 685924 538441 685958
rect 550739 685924 550835 685958
rect 538345 685862 538379 685924
rect 550801 685862 550835 685924
rect 538524 685810 538540 685844
rect 539516 685810 539532 685844
rect 539760 685810 539776 685844
rect 540752 685810 540768 685844
rect 540996 685810 541012 685844
rect 541988 685810 542004 685844
rect 542232 685810 542248 685844
rect 543224 685810 543240 685844
rect 543468 685810 543484 685844
rect 544460 685810 544476 685844
rect 544704 685810 544720 685844
rect 545696 685810 545712 685844
rect 545940 685810 545956 685844
rect 546932 685810 546948 685844
rect 547176 685810 547192 685844
rect 548168 685810 548184 685844
rect 548412 685810 548428 685844
rect 549404 685810 549420 685844
rect 549648 685810 549664 685844
rect 550640 685810 550656 685844
rect 538447 685782 538481 685798
rect 538447 685698 538481 685714
rect 539575 685782 539609 685798
rect 539575 685698 539609 685714
rect 539683 685782 539717 685798
rect 539683 685698 539717 685714
rect 540811 685782 540845 685798
rect 540811 685698 540845 685714
rect 540919 685782 540953 685798
rect 540919 685698 540953 685714
rect 542047 685782 542081 685798
rect 542047 685698 542081 685714
rect 542155 685782 542189 685798
rect 542155 685698 542189 685714
rect 543283 685782 543317 685798
rect 543283 685698 543317 685714
rect 543391 685782 543425 685798
rect 543391 685698 543425 685714
rect 544519 685782 544553 685798
rect 544519 685698 544553 685714
rect 544627 685782 544661 685798
rect 544627 685698 544661 685714
rect 545755 685782 545789 685798
rect 545755 685698 545789 685714
rect 545863 685782 545897 685798
rect 545863 685698 545897 685714
rect 546991 685782 547025 685798
rect 546991 685698 547025 685714
rect 547099 685782 547133 685798
rect 547099 685698 547133 685714
rect 548227 685782 548261 685798
rect 548227 685698 548261 685714
rect 548335 685782 548369 685798
rect 548335 685698 548369 685714
rect 549463 685782 549497 685798
rect 549463 685698 549497 685714
rect 549571 685782 549605 685798
rect 549571 685698 549605 685714
rect 550699 685782 550733 685798
rect 550699 685698 550733 685714
rect 538524 685652 538540 685686
rect 539516 685652 539532 685686
rect 539760 685652 539776 685686
rect 540752 685652 540768 685686
rect 540996 685652 541012 685686
rect 541988 685652 542004 685686
rect 542232 685652 542248 685686
rect 543224 685652 543240 685686
rect 543468 685652 543484 685686
rect 544460 685652 544476 685686
rect 544704 685652 544720 685686
rect 545696 685652 545712 685686
rect 545940 685652 545956 685686
rect 546932 685652 546948 685686
rect 547176 685652 547192 685686
rect 548168 685652 548184 685686
rect 548412 685652 548428 685686
rect 549404 685652 549420 685686
rect 549648 685652 549664 685686
rect 550640 685652 550656 685686
rect 538345 685572 538379 685634
rect 550801 685572 550835 685634
rect 538345 685538 538441 685572
rect 550739 685538 550835 685572
rect 537682 685259 537716 685321
rect 534592 685225 534688 685259
rect 537620 685225 537716 685259
rect 554742 686535 554776 686597
rect 551652 685259 551686 685321
rect 554742 685259 554776 685321
rect 551652 685225 551748 685259
rect 554680 685225 554776 685259
rect 540285 685144 540381 685178
rect 548845 685144 548941 685178
rect 46556 684720 46590 684782
rect 540285 685082 540319 685144
rect 548907 685082 548941 685144
rect 540455 685030 540471 685064
rect 541447 685030 541463 685064
rect 541673 685030 541689 685064
rect 542665 685030 542681 685064
rect 542891 685030 542907 685064
rect 543883 685030 543899 685064
rect 544109 685030 544125 685064
rect 545101 685030 545117 685064
rect 545327 685030 545343 685064
rect 546319 685030 546335 685064
rect 546545 685030 546561 685064
rect 547537 685030 547553 685064
rect 547763 685030 547779 685064
rect 548755 685030 548771 685064
rect 540387 685002 540421 685018
rect 540387 684918 540421 684934
rect 541497 685002 541531 685018
rect 541497 684918 541531 684934
rect 541605 685002 541639 685018
rect 541605 684918 541639 684934
rect 542715 685002 542749 685018
rect 542715 684918 542749 684934
rect 542823 685002 542857 685018
rect 542823 684918 542857 684934
rect 543933 685002 543967 685018
rect 543933 684918 543967 684934
rect 544041 685002 544075 685018
rect 544041 684918 544075 684934
rect 545151 685002 545185 685018
rect 545151 684918 545185 684934
rect 545259 685002 545293 685018
rect 545259 684918 545293 684934
rect 546369 685002 546403 685018
rect 546369 684918 546403 684934
rect 546477 685002 546511 685018
rect 546477 684918 546511 684934
rect 547587 685002 547621 685018
rect 547587 684918 547621 684934
rect 547695 685002 547729 685018
rect 547695 684918 547729 684934
rect 548805 685002 548839 685018
rect 548805 684918 548839 684934
rect 540455 684872 540471 684906
rect 541447 684872 541463 684906
rect 541673 684872 541689 684906
rect 542665 684872 542681 684906
rect 542891 684872 542907 684906
rect 543883 684872 543899 684906
rect 544109 684872 544125 684906
rect 545101 684872 545117 684906
rect 545327 684872 545343 684906
rect 546319 684872 546335 684906
rect 546545 684872 546561 684906
rect 547537 684872 547553 684906
rect 547763 684872 547779 684906
rect 548755 684872 548771 684906
rect 540285 684792 540319 684854
rect 548907 684792 548941 684854
rect 540285 684758 540381 684792
rect 548845 684758 548941 684792
rect 42716 684686 42812 684720
rect 46494 684686 46590 684720
rect 540285 684644 540381 684678
rect 548845 684644 548941 684678
rect 540285 684582 540319 684644
rect 548907 684582 548941 684644
rect 540455 684530 540471 684564
rect 541447 684530 541463 684564
rect 541673 684530 541689 684564
rect 542665 684530 542681 684564
rect 542891 684530 542907 684564
rect 543883 684530 543899 684564
rect 544109 684530 544125 684564
rect 545101 684530 545117 684564
rect 545327 684530 545343 684564
rect 546319 684530 546335 684564
rect 546545 684530 546561 684564
rect 547537 684530 547553 684564
rect 547763 684530 547779 684564
rect 548755 684530 548771 684564
rect 540387 684502 540421 684518
rect 540387 684418 540421 684434
rect 541497 684502 541531 684518
rect 541497 684418 541531 684434
rect 541605 684502 541639 684518
rect 541605 684418 541639 684434
rect 542715 684502 542749 684518
rect 542715 684418 542749 684434
rect 542823 684502 542857 684518
rect 542823 684418 542857 684434
rect 543933 684502 543967 684518
rect 543933 684418 543967 684434
rect 544041 684502 544075 684518
rect 544041 684418 544075 684434
rect 545151 684502 545185 684518
rect 545151 684418 545185 684434
rect 545259 684502 545293 684518
rect 545259 684418 545293 684434
rect 546369 684502 546403 684518
rect 546369 684418 546403 684434
rect 546477 684502 546511 684518
rect 546477 684418 546511 684434
rect 547587 684502 547621 684518
rect 547587 684418 547621 684434
rect 547695 684502 547729 684518
rect 547695 684418 547729 684434
rect 548805 684502 548839 684518
rect 548805 684418 548839 684434
rect 540455 684372 540471 684406
rect 541447 684372 541463 684406
rect 541673 684372 541689 684406
rect 542665 684372 542681 684406
rect 542891 684372 542907 684406
rect 543883 684372 543899 684406
rect 544109 684372 544125 684406
rect 545101 684372 545117 684406
rect 545327 684372 545343 684406
rect 546319 684372 546335 684406
rect 546545 684372 546561 684406
rect 547537 684372 547553 684406
rect 547763 684372 547779 684406
rect 548755 684372 548771 684406
rect 540285 684292 540319 684354
rect 548907 684292 548941 684354
rect 540285 684258 540381 684292
rect 548845 684258 548941 684292
rect 540845 684144 540941 684178
rect 548187 684144 548283 684178
rect 540845 684082 540879 684144
rect 43746 683968 43842 684002
rect 45460 683968 45556 684002
rect 43746 683906 43780 683968
rect 45522 683906 45556 683968
rect 43906 683866 43922 683900
rect 44090 683866 44106 683900
rect 44164 683866 44180 683900
rect 44348 683866 44364 683900
rect 44422 683866 44438 683900
rect 44606 683866 44622 683900
rect 44680 683866 44696 683900
rect 44864 683866 44880 683900
rect 44938 683866 44954 683900
rect 45122 683866 45138 683900
rect 45196 683866 45212 683900
rect 45380 683866 45396 683900
rect 43860 683807 43894 683823
rect 43860 682815 43894 682831
rect 44118 683807 44152 683823
rect 44118 682815 44152 682831
rect 44376 683807 44410 683823
rect 44376 682815 44410 682831
rect 44634 683807 44668 683823
rect 44634 682815 44668 682831
rect 44892 683807 44926 683823
rect 44892 682815 44926 682831
rect 45150 683807 45184 683823
rect 45150 682815 45184 682831
rect 45408 683807 45442 683823
rect 548249 684082 548283 684144
rect 541015 684030 541031 684064
rect 542007 684030 542023 684064
rect 542233 684030 542249 684064
rect 543225 684030 543241 684064
rect 543451 684030 543467 684064
rect 544443 684030 544459 684064
rect 544669 684030 544685 684064
rect 545661 684030 545677 684064
rect 545887 684030 545903 684064
rect 546879 684030 546895 684064
rect 547105 684030 547121 684064
rect 548097 684030 548113 684064
rect 540947 684002 540981 684018
rect 540947 683818 540981 683834
rect 542057 684002 542091 684018
rect 542057 683818 542091 683834
rect 542165 684002 542199 684018
rect 542165 683818 542199 683834
rect 543275 684002 543309 684018
rect 543275 683818 543309 683834
rect 543383 684002 543417 684018
rect 543383 683818 543417 683834
rect 544493 684002 544527 684018
rect 544493 683818 544527 683834
rect 544601 684002 544635 684018
rect 544601 683818 544635 683834
rect 545711 684002 545745 684018
rect 545711 683818 545745 683834
rect 545819 684002 545853 684018
rect 545819 683818 545853 683834
rect 546929 684002 546963 684018
rect 546929 683818 546963 683834
rect 547037 684002 547071 684018
rect 547037 683818 547071 683834
rect 548147 684002 548181 684018
rect 548147 683818 548181 683834
rect 541015 683772 541031 683806
rect 542007 683772 542023 683806
rect 542233 683772 542249 683806
rect 543225 683772 543241 683806
rect 543451 683772 543467 683806
rect 544443 683772 544459 683806
rect 544669 683772 544685 683806
rect 545661 683772 545677 683806
rect 545887 683772 545903 683806
rect 546879 683772 546895 683806
rect 547105 683772 547121 683806
rect 548097 683772 548113 683806
rect 540845 683692 540879 683754
rect 548249 683692 548283 683754
rect 540845 683658 540941 683692
rect 548187 683658 548283 683692
rect 541539 683652 541709 683658
rect 541539 683562 541569 683652
rect 541679 683562 541709 683652
rect 541539 683558 541709 683562
rect 546449 683652 546619 683658
rect 546449 683562 546479 683652
rect 546589 683562 546619 683652
rect 546449 683558 546619 683562
rect 540845 683524 540941 683558
rect 548187 683524 548283 683558
rect 540845 683462 540879 683524
rect 45408 682815 45442 682831
rect 43906 682738 43922 682772
rect 44090 682738 44106 682772
rect 44164 682738 44180 682772
rect 44348 682738 44364 682772
rect 44422 682738 44438 682772
rect 44606 682738 44622 682772
rect 44680 682738 44696 682772
rect 44864 682738 44880 682772
rect 44938 682738 44954 682772
rect 45122 682738 45138 682772
rect 45196 682738 45212 682772
rect 45380 682738 45396 682772
rect 43746 682670 43780 682732
rect 548249 683462 548283 683524
rect 541015 683410 541031 683444
rect 542007 683410 542023 683444
rect 542233 683410 542249 683444
rect 543225 683410 543241 683444
rect 543451 683410 543467 683444
rect 544443 683410 544459 683444
rect 544669 683410 544685 683444
rect 545661 683410 545677 683444
rect 545887 683410 545903 683444
rect 546879 683410 546895 683444
rect 547105 683410 547121 683444
rect 548097 683410 548113 683444
rect 540947 683382 540981 683398
rect 540947 683198 540981 683214
rect 542057 683382 542091 683398
rect 542057 683198 542091 683214
rect 542165 683382 542199 683398
rect 542165 683198 542199 683214
rect 543275 683382 543309 683398
rect 543275 683198 543309 683214
rect 543383 683382 543417 683398
rect 543383 683198 543417 683214
rect 544493 683382 544527 683398
rect 544493 683198 544527 683214
rect 544601 683382 544635 683398
rect 544601 683198 544635 683214
rect 545711 683382 545745 683398
rect 545711 683198 545745 683214
rect 545819 683382 545853 683398
rect 545819 683198 545853 683214
rect 546929 683382 546963 683398
rect 546929 683198 546963 683214
rect 547037 683382 547071 683398
rect 547037 683198 547071 683214
rect 548147 683382 548181 683398
rect 548147 683198 548181 683214
rect 541015 683152 541031 683186
rect 542007 683152 542023 683186
rect 542233 683152 542249 683186
rect 543225 683152 543241 683186
rect 543451 683152 543467 683186
rect 544443 683152 544459 683186
rect 544669 683152 544685 683186
rect 545661 683152 545677 683186
rect 545887 683152 545903 683186
rect 546879 683152 546895 683186
rect 547105 683152 547121 683186
rect 548097 683152 548113 683186
rect 540845 683072 540879 683134
rect 548249 683072 548283 683134
rect 540845 683038 540941 683072
rect 548187 683038 548283 683072
rect 45522 682670 45556 682732
rect 43746 682636 43842 682670
rect 45460 682636 45556 682670
rect 540285 682924 540381 682958
rect 548845 682924 548941 682958
rect 540285 682862 540319 682924
rect 548907 682862 548941 682924
rect 540455 682810 540471 682844
rect 541447 682810 541463 682844
rect 541673 682810 541689 682844
rect 542665 682810 542681 682844
rect 542891 682810 542907 682844
rect 543883 682810 543899 682844
rect 544109 682810 544125 682844
rect 545101 682810 545117 682844
rect 545327 682810 545343 682844
rect 546319 682810 546335 682844
rect 546545 682810 546561 682844
rect 547537 682810 547553 682844
rect 547763 682810 547779 682844
rect 548755 682810 548771 682844
rect 540387 682782 540421 682798
rect 540387 682598 540421 682614
rect 541497 682782 541531 682798
rect 541497 682598 541531 682614
rect 541605 682782 541639 682798
rect 541605 682598 541639 682614
rect 542715 682782 542749 682798
rect 542715 682598 542749 682614
rect 542823 682782 542857 682798
rect 542823 682598 542857 682614
rect 543933 682782 543967 682798
rect 543933 682598 543967 682614
rect 544041 682782 544075 682798
rect 544041 682598 544075 682614
rect 545151 682782 545185 682798
rect 545151 682598 545185 682614
rect 545259 682782 545293 682798
rect 545259 682598 545293 682614
rect 546369 682782 546403 682798
rect 546369 682598 546403 682614
rect 546477 682782 546511 682798
rect 546477 682598 546511 682614
rect 547587 682782 547621 682798
rect 547587 682598 547621 682614
rect 547695 682782 547729 682798
rect 547695 682598 547729 682614
rect 548805 682782 548839 682798
rect 548805 682598 548839 682614
rect 540455 682552 540471 682586
rect 541447 682552 541463 682586
rect 541673 682552 541689 682586
rect 542665 682552 542681 682586
rect 542891 682552 542907 682586
rect 543883 682552 543899 682586
rect 544109 682552 544125 682586
rect 545101 682552 545117 682586
rect 545327 682552 545343 682586
rect 546319 682552 546335 682586
rect 546545 682552 546561 682586
rect 547537 682552 547553 682586
rect 547763 682552 547779 682586
rect 548755 682552 548771 682586
rect 43746 682468 43842 682502
rect 45460 682468 45556 682502
rect 43746 682406 43780 682468
rect 45522 682406 45556 682468
rect 540285 682472 540319 682534
rect 548907 682472 548941 682534
rect 540285 682438 540381 682472
rect 548845 682438 548941 682472
rect 43906 682366 43922 682400
rect 44090 682366 44106 682400
rect 44164 682366 44180 682400
rect 44348 682366 44364 682400
rect 44422 682366 44438 682400
rect 44606 682366 44622 682400
rect 44680 682366 44696 682400
rect 44864 682366 44880 682400
rect 44938 682366 44954 682400
rect 45122 682366 45138 682400
rect 45196 682366 45212 682400
rect 45380 682366 45396 682400
rect 43860 682307 43894 682323
rect 43860 681315 43894 681331
rect 44118 682307 44152 682323
rect 44118 681315 44152 681331
rect 44376 682307 44410 682323
rect 44376 681315 44410 681331
rect 44634 682307 44668 682323
rect 44634 681315 44668 681331
rect 44892 682307 44926 682323
rect 44892 681315 44926 681331
rect 45150 682307 45184 682323
rect 45150 681315 45184 681331
rect 45408 682307 45442 682323
rect 540285 682324 540381 682358
rect 548845 682324 548941 682358
rect 540285 682262 540319 682324
rect 548907 682262 548941 682324
rect 540455 682210 540471 682244
rect 541447 682210 541463 682244
rect 541673 682210 541689 682244
rect 542665 682210 542681 682244
rect 542891 682210 542907 682244
rect 543883 682210 543899 682244
rect 544109 682210 544125 682244
rect 545101 682210 545117 682244
rect 545327 682210 545343 682244
rect 546319 682210 546335 682244
rect 546545 682210 546561 682244
rect 547537 682210 547553 682244
rect 547763 682210 547779 682244
rect 548755 682210 548771 682244
rect 540387 682182 540421 682198
rect 540387 681998 540421 682014
rect 541497 682182 541531 682198
rect 541497 681998 541531 682014
rect 541605 682182 541639 682198
rect 541605 681998 541639 682014
rect 542715 682182 542749 682198
rect 542715 681998 542749 682014
rect 542823 682182 542857 682198
rect 542823 681998 542857 682014
rect 543933 682182 543967 682198
rect 543933 681998 543967 682014
rect 544041 682182 544075 682198
rect 544041 681998 544075 682014
rect 545151 682182 545185 682198
rect 545151 681998 545185 682014
rect 545259 682182 545293 682198
rect 545259 681998 545293 682014
rect 546369 682182 546403 682198
rect 546369 681998 546403 682014
rect 546477 682182 546511 682198
rect 546477 681998 546511 682014
rect 547587 682182 547621 682198
rect 547587 681998 547621 682014
rect 547695 682182 547729 682198
rect 547695 681998 547729 682014
rect 548805 682182 548839 682198
rect 548805 681998 548839 682014
rect 540455 681952 540471 681986
rect 541447 681952 541463 681986
rect 541673 681952 541689 681986
rect 542665 681952 542681 681986
rect 542891 681952 542907 681986
rect 543883 681952 543899 681986
rect 544109 681952 544125 681986
rect 545101 681952 545117 681986
rect 545327 681952 545343 681986
rect 546319 681952 546335 681986
rect 546545 681952 546561 681986
rect 547537 681952 547553 681986
rect 547763 681952 547779 681986
rect 548755 681952 548771 681986
rect 540285 681872 540319 681934
rect 548907 681872 548941 681934
rect 540285 681838 540381 681872
rect 548845 681838 548941 681872
rect 45408 681315 45442 681331
rect 43906 681238 43922 681272
rect 44090 681238 44106 681272
rect 44164 681238 44180 681272
rect 44348 681238 44364 681272
rect 44606 681238 44622 681272
rect 44680 681238 44696 681272
rect 44864 681238 44880 681272
rect 44938 681238 44954 681272
rect 45122 681238 45138 681272
rect 45196 681238 45212 681272
rect 45380 681238 45396 681272
rect 43746 681170 43780 681232
rect 45522 681170 45556 681232
rect 43746 681136 43842 681170
rect 45460 681136 45556 681170
rect 540830 681350 540926 681384
rect 548280 681350 548376 681384
rect 540830 681288 540864 681350
rect 548342 681288 548376 681350
rect 541009 681236 541025 681270
rect 542001 681236 542017 681270
rect 542245 681236 542261 681270
rect 543237 681236 543253 681270
rect 543481 681236 543497 681270
rect 544473 681236 544489 681270
rect 544717 681236 544733 681270
rect 545709 681236 545725 681270
rect 545953 681236 545969 681270
rect 546945 681236 546961 681270
rect 547189 681236 547205 681270
rect 548181 681236 548197 681270
rect 540932 681208 540966 681224
rect 540932 681024 540966 681040
rect 542060 681208 542094 681224
rect 542060 681024 542094 681040
rect 542168 681208 542202 681224
rect 542168 681024 542202 681040
rect 543296 681208 543330 681224
rect 543296 681024 543330 681040
rect 543404 681208 543438 681224
rect 543404 681024 543438 681040
rect 544532 681208 544566 681224
rect 544532 681024 544566 681040
rect 544640 681208 544674 681224
rect 544640 681024 544674 681040
rect 545768 681208 545802 681224
rect 545768 681024 545802 681040
rect 545876 681208 545910 681224
rect 545876 681024 545910 681040
rect 547004 681208 547038 681224
rect 547004 681024 547038 681040
rect 547112 681208 547146 681224
rect 547112 681024 547146 681040
rect 548240 681208 548274 681224
rect 548240 681024 548274 681040
rect 541009 680978 541025 681012
rect 542001 680978 542017 681012
rect 542245 680978 542261 681012
rect 543237 680978 543253 681012
rect 543481 680978 543497 681012
rect 544473 680978 544489 681012
rect 544717 680978 544733 681012
rect 545709 680978 545725 681012
rect 545953 680978 545969 681012
rect 546945 680978 546961 681012
rect 547189 680978 547205 681012
rect 548181 680978 548197 681012
rect 540830 680898 540864 680960
rect 548342 680898 548376 680960
rect 44346 680850 44442 680884
rect 44828 680850 44924 680884
rect 540830 680864 540926 680898
rect 548280 680864 548376 680898
rect 44346 680788 44380 680850
rect 44890 680788 44924 680850
rect 44506 680748 44522 680782
rect 44590 680748 44606 680782
rect 44664 680748 44680 680782
rect 44748 680748 44764 680782
rect 44460 680698 44494 680714
rect 44460 680206 44494 680222
rect 44618 680698 44652 680714
rect 44618 680206 44652 680222
rect 44776 680698 44810 680714
rect 44776 680206 44810 680222
rect 540830 680760 540926 680794
rect 548280 680760 548376 680794
rect 540830 680698 540864 680760
rect 548342 680698 548376 680760
rect 541009 680646 541025 680680
rect 542001 680646 542017 680680
rect 542245 680646 542261 680680
rect 543237 680646 543253 680680
rect 543481 680646 543497 680680
rect 544473 680646 544489 680680
rect 544717 680646 544733 680680
rect 545709 680646 545725 680680
rect 545953 680646 545969 680680
rect 546945 680646 546961 680680
rect 547189 680646 547205 680680
rect 548181 680646 548197 680680
rect 540932 680618 540966 680634
rect 540932 680434 540966 680450
rect 542060 680618 542094 680634
rect 542060 680434 542094 680450
rect 542168 680618 542202 680634
rect 542168 680434 542202 680450
rect 543296 680618 543330 680634
rect 543296 680434 543330 680450
rect 543404 680618 543438 680634
rect 543404 680434 543438 680450
rect 544532 680618 544566 680634
rect 544532 680434 544566 680450
rect 544640 680618 544674 680634
rect 544640 680434 544674 680450
rect 545768 680618 545802 680634
rect 545768 680434 545802 680450
rect 545876 680618 545910 680634
rect 545876 680434 545910 680450
rect 547004 680618 547038 680634
rect 547004 680434 547038 680450
rect 547112 680618 547146 680634
rect 547112 680434 547146 680450
rect 548240 680618 548274 680634
rect 548240 680434 548274 680450
rect 541009 680388 541025 680422
rect 542001 680388 542017 680422
rect 542245 680388 542261 680422
rect 543237 680388 543253 680422
rect 543481 680388 543497 680422
rect 544473 680388 544489 680422
rect 544717 680388 544733 680422
rect 545709 680388 545725 680422
rect 545953 680388 545969 680422
rect 546945 680388 546961 680422
rect 547189 680388 547205 680422
rect 548181 680388 548197 680422
rect 44506 680138 44522 680172
rect 44590 680138 44606 680172
rect 44664 680138 44680 680172
rect 44748 680138 44764 680172
rect 44346 680070 44380 680132
rect 540830 680308 540864 680370
rect 548342 680308 548376 680370
rect 540830 680274 540926 680308
rect 548280 680274 548376 680308
rect 44890 680070 44924 680132
rect 44346 680036 44442 680070
rect 44828 680036 44924 680070
rect 543600 679970 543696 680004
rect 545506 679970 545602 680004
rect 543600 679908 543634 679970
rect 43986 679850 44082 679884
rect 45184 679850 45280 679884
rect 43986 679788 44020 679850
rect 45246 679788 45280 679850
rect 44146 679748 44162 679782
rect 44330 679748 44346 679782
rect 44404 679748 44420 679782
rect 44588 679748 44604 679782
rect 44662 679748 44678 679782
rect 44846 679748 44862 679782
rect 44920 679748 44936 679782
rect 45104 679748 45120 679782
rect 44100 679698 44134 679714
rect 44100 679456 44134 679472
rect 44358 679698 44392 679714
rect 44358 679456 44392 679472
rect 44616 679698 44650 679714
rect 44616 679456 44650 679472
rect 44874 679698 44908 679714
rect 44874 679456 44908 679472
rect 45132 679698 45166 679714
rect 545568 679908 545602 679970
rect 543770 679856 543786 679890
rect 544012 679856 544028 679890
rect 544238 679856 544254 679890
rect 544480 679856 544496 679890
rect 544706 679856 544722 679890
rect 544948 679856 544964 679890
rect 545174 679856 545190 679890
rect 545416 679856 545432 679890
rect 543702 679828 543736 679844
rect 543702 679644 543736 679660
rect 544062 679828 544096 679844
rect 544062 679644 544096 679660
rect 544170 679828 544204 679844
rect 544170 679644 544204 679660
rect 544530 679828 544564 679844
rect 544530 679644 544564 679660
rect 544638 679828 544672 679844
rect 544638 679644 544672 679660
rect 544998 679828 545032 679844
rect 544998 679644 545032 679660
rect 545106 679828 545140 679844
rect 545106 679644 545140 679660
rect 545466 679828 545500 679844
rect 545466 679644 545500 679660
rect 543770 679598 543786 679632
rect 544012 679598 544028 679632
rect 544238 679598 544254 679632
rect 544480 679598 544496 679632
rect 544706 679598 544722 679632
rect 544948 679598 544964 679632
rect 545174 679598 545190 679632
rect 545416 679598 545432 679632
rect 45132 679456 45166 679472
rect 44146 679388 44162 679422
rect 44330 679388 44346 679422
rect 44404 679388 44420 679422
rect 44588 679388 44604 679422
rect 44662 679388 44678 679422
rect 44846 679388 44862 679422
rect 44920 679388 44936 679422
rect 45104 679388 45120 679422
rect 43986 679320 44020 679382
rect 543600 679518 543634 679580
rect 545568 679518 545602 679580
rect 543600 679484 543696 679518
rect 545506 679484 545602 679518
rect 45246 679320 45280 679382
rect 43986 679286 44082 679320
rect 45184 679286 45280 679320
rect 543820 679345 543916 679368
rect 545290 679345 545386 679368
rect 543820 679283 543854 679345
rect 43731 679100 43827 679134
rect 45445 679100 45541 679134
rect 43731 679038 43765 679100
rect 45507 679038 45541 679100
rect 43891 678998 43907 679032
rect 44075 678998 44091 679032
rect 44149 678998 44165 679032
rect 44333 678998 44349 679032
rect 44407 678998 44423 679032
rect 44591 678998 44607 679032
rect 44665 678998 44681 679032
rect 44849 678998 44865 679032
rect 44923 678998 44939 679032
rect 45107 678998 45123 679032
rect 45181 678998 45197 679032
rect 45365 678998 45381 679032
rect 43845 678948 43879 678964
rect 43845 677956 43879 677972
rect 44103 678948 44137 678964
rect 44103 677956 44137 677972
rect 44361 678948 44395 678964
rect 44361 677956 44395 677972
rect 44619 678948 44653 678964
rect 44619 677956 44653 677972
rect 44877 678948 44911 678964
rect 44877 677956 44911 677972
rect 45135 678948 45169 678964
rect 45135 677956 45169 677972
rect 45393 678948 45427 678964
rect 45393 677956 45427 677972
rect 43891 677888 43907 677922
rect 44075 677888 44091 677922
rect 44149 677888 44165 677922
rect 44333 677888 44349 677922
rect 44407 677888 44423 677922
rect 44591 677888 44607 677922
rect 44665 677888 44681 677922
rect 44849 677888 44865 677922
rect 44923 677888 44939 677922
rect 45107 677888 45123 677922
rect 45181 677888 45197 677922
rect 45365 677888 45381 677922
rect 43731 677820 43765 677882
rect 545352 679283 545386 679345
rect 543990 679231 544006 679265
rect 544482 679231 544498 679265
rect 544708 679231 544724 679265
rect 545200 679231 545216 679265
rect 543922 679203 543956 679219
rect 543922 679119 543956 679135
rect 544532 679203 544566 679219
rect 544532 679119 544566 679135
rect 544640 679203 544674 679219
rect 544640 679119 544674 679135
rect 545250 679203 545284 679219
rect 545250 679119 545284 679135
rect 543990 679073 544006 679107
rect 544482 679073 544498 679107
rect 544708 679073 544724 679107
rect 545200 679073 545216 679107
rect 543820 678993 543854 679055
rect 545352 678993 545386 679055
rect 543820 678959 543916 678993
rect 545290 678959 545386 678993
rect 540885 678820 540981 678854
rect 548227 678820 548323 678854
rect 540885 678758 540919 678820
rect 548289 678758 548323 678820
rect 541055 678706 541071 678740
rect 542047 678706 542063 678740
rect 542273 678706 542289 678740
rect 543265 678706 543281 678740
rect 543491 678706 543507 678740
rect 544483 678706 544499 678740
rect 544709 678706 544725 678740
rect 545701 678706 545717 678740
rect 545927 678706 545943 678740
rect 546919 678706 546935 678740
rect 547145 678706 547161 678740
rect 548137 678706 548153 678740
rect 540987 678678 541021 678694
rect 540987 678494 541021 678510
rect 542097 678678 542131 678694
rect 542097 678494 542131 678510
rect 542205 678678 542239 678694
rect 542205 678494 542239 678510
rect 543315 678678 543349 678694
rect 543315 678494 543349 678510
rect 543423 678678 543457 678694
rect 543423 678494 543457 678510
rect 544533 678678 544567 678694
rect 544533 678494 544567 678510
rect 544641 678678 544675 678694
rect 544641 678494 544675 678510
rect 545751 678678 545785 678694
rect 545751 678494 545785 678510
rect 545859 678678 545893 678694
rect 545859 678494 545893 678510
rect 546969 678678 547003 678694
rect 546969 678494 547003 678510
rect 547077 678678 547111 678694
rect 547077 678494 547111 678510
rect 548187 678678 548221 678694
rect 548187 678494 548221 678510
rect 541055 678448 541071 678482
rect 542047 678448 542063 678482
rect 542273 678448 542289 678482
rect 543265 678448 543281 678482
rect 543491 678448 543507 678482
rect 544483 678448 544499 678482
rect 544709 678448 544725 678482
rect 545701 678448 545717 678482
rect 545927 678448 545943 678482
rect 546919 678448 546935 678482
rect 547145 678448 547161 678482
rect 548137 678448 548153 678482
rect 540885 678368 540919 678430
rect 548289 678368 548323 678430
rect 540885 678334 540981 678368
rect 548227 678334 548323 678368
rect 45507 677820 45541 677882
rect 43731 677786 43827 677820
rect 45445 677786 45541 677820
rect 541364 677058 541484 677074
rect 41200 676980 41440 676996
rect 41200 676724 41440 676740
rect 47900 676980 48140 676996
rect 541364 676922 541484 676938
rect 547734 677058 547854 677074
rect 547734 676922 547854 676938
rect 47900 676724 48140 676740
rect 41200 675260 41440 675276
rect 41200 675004 41440 675020
rect 47900 675260 48140 675276
rect 47900 675004 48140 675020
rect 541364 674058 541484 674074
rect 541364 673922 541484 673938
rect 547734 674058 547854 674074
rect 547734 673922 547854 673938
rect 41200 673540 41440 673556
rect 41200 673284 41440 673300
rect 47900 673540 48140 673556
rect 47900 673284 48140 673300
rect 41200 672060 41440 672076
rect 41200 671804 41440 671820
rect 47900 672060 48140 672076
rect 47900 671804 48140 671820
rect 541364 671058 541484 671074
rect 541364 670922 541484 670938
rect 547734 671058 547854 671074
rect 547734 670922 547854 670938
rect 41200 670340 41440 670356
rect 41200 670084 41440 670100
rect 47900 670340 48140 670356
rect 47900 670084 48140 670100
rect 41200 668740 41440 668756
rect 41200 668484 41440 668500
rect 47900 668740 48140 668756
rect 47900 668484 48140 668500
rect 541364 668058 541484 668074
rect 541364 667922 541484 667938
rect 547734 668058 547854 668074
rect 547734 667922 547854 667938
rect 41200 667020 41440 667036
rect 41200 666764 41440 666780
rect 47900 667020 48140 667036
rect 47900 666764 48140 666780
rect 41200 665420 41440 665436
rect 41200 665164 41440 665180
rect 47900 665420 48140 665436
rect 47900 665164 48140 665180
rect 541364 665058 541484 665074
rect 541364 664922 541484 664938
rect 547734 665058 547854 665074
rect 547734 664922 547854 664938
rect 41200 663700 41440 663716
rect 41200 663444 41440 663460
rect 47900 663700 48140 663716
rect 47900 663444 48140 663460
<< viali >>
rect 37711 694999 38108 696113
rect 40142 694999 40539 696113
rect 43029 695348 46285 695382
rect 37711 693539 38108 694653
rect 40142 693539 40539 694653
rect 41542 695246 41610 695280
rect 41700 695246 41768 695280
rect 41858 695246 41926 695280
rect 42016 695246 42084 695280
rect 42174 695246 42242 695280
rect 42332 695246 42400 695280
rect 42490 695246 42558 695280
rect 42648 695246 42716 695280
rect 42806 695246 42874 695280
rect 42964 695246 43032 695280
rect 43122 695246 43190 695280
rect 43280 695246 43348 695280
rect 43438 695246 43506 695280
rect 43596 695246 43664 695280
rect 43754 695246 43822 695280
rect 43912 695246 43980 695280
rect 44070 695246 44138 695280
rect 44228 695246 44296 695280
rect 44386 695246 44454 695280
rect 44544 695246 44612 695280
rect 44702 695246 44770 695280
rect 44860 695246 44928 695280
rect 45018 695246 45086 695280
rect 45176 695246 45244 695280
rect 45334 695246 45402 695280
rect 45492 695246 45560 695280
rect 45650 695246 45718 695280
rect 45808 695246 45876 695280
rect 45966 695246 46034 695280
rect 46124 695246 46192 695280
rect 46282 695246 46350 695280
rect 46440 695246 46508 695280
rect 46598 695246 46666 695280
rect 46756 695246 46824 695280
rect 46914 695246 46982 695280
rect 47072 695246 47140 695280
rect 47230 695246 47298 695280
rect 47388 695246 47456 695280
rect 47546 695246 47614 695280
rect 47704 695246 47772 695280
rect 41480 694211 41514 695187
rect 41638 694211 41672 695187
rect 41796 694211 41830 695187
rect 41954 694211 41988 695187
rect 42112 694211 42146 695187
rect 42270 694211 42304 695187
rect 42428 694211 42462 695187
rect 42586 694211 42620 695187
rect 42744 694211 42778 695187
rect 42902 694211 42936 695187
rect 43060 694211 43094 695187
rect 43218 694211 43252 695187
rect 43376 694211 43410 695187
rect 43534 694211 43568 695187
rect 43692 694211 43726 695187
rect 43850 694211 43884 695187
rect 44008 694211 44042 695187
rect 44166 694211 44200 695187
rect 44324 694211 44358 695187
rect 44482 694211 44516 695187
rect 44640 694211 44674 695187
rect 44798 694211 44832 695187
rect 44956 694211 44990 695187
rect 45114 694211 45148 695187
rect 45272 694211 45306 695187
rect 45430 694211 45464 695187
rect 45588 694211 45622 695187
rect 45746 694211 45780 695187
rect 45904 694211 45938 695187
rect 46062 694211 46096 695187
rect 46220 694211 46254 695187
rect 46378 694211 46412 695187
rect 46536 694211 46570 695187
rect 46694 694211 46728 695187
rect 46852 694211 46886 695187
rect 47010 694211 47044 695187
rect 47168 694211 47202 695187
rect 47326 694211 47360 695187
rect 47484 694211 47518 695187
rect 47642 694211 47676 695187
rect 47800 694211 47834 695187
rect 41542 694118 41610 694152
rect 41700 694118 41768 694152
rect 41858 694118 41926 694152
rect 42016 694118 42084 694152
rect 42174 694118 42242 694152
rect 42332 694118 42400 694152
rect 42490 694118 42558 694152
rect 42648 694118 42716 694152
rect 42806 694118 42874 694152
rect 42964 694118 43032 694152
rect 43122 694118 43190 694152
rect 43280 694118 43348 694152
rect 43438 694118 43506 694152
rect 43596 694118 43664 694152
rect 43754 694118 43822 694152
rect 43912 694118 43980 694152
rect 44070 694118 44138 694152
rect 44228 694118 44296 694152
rect 44386 694118 44454 694152
rect 44544 694118 44612 694152
rect 44702 694118 44770 694152
rect 44860 694118 44928 694152
rect 45018 694118 45086 694152
rect 45176 694118 45244 694152
rect 45334 694118 45402 694152
rect 45492 694118 45560 694152
rect 45650 694118 45718 694152
rect 45808 694118 45876 694152
rect 45966 694118 46034 694152
rect 46124 694118 46192 694152
rect 46282 694118 46350 694152
rect 46440 694118 46508 694152
rect 46598 694118 46666 694152
rect 46756 694118 46824 694152
rect 46914 694118 46982 694152
rect 47072 694118 47140 694152
rect 47230 694118 47298 694152
rect 47388 694118 47456 694152
rect 47546 694118 47614 694152
rect 47704 694118 47772 694152
rect 48781 694999 49178 696113
rect 51212 694999 51609 696113
rect 43029 694016 46285 694050
rect 38700 693427 38880 693460
rect 39120 693427 39300 693460
rect 38700 693393 38880 693427
rect 39120 693393 39300 693427
rect 43778 693678 45534 693712
rect 38700 693360 38880 693393
rect 39120 693360 39300 693393
rect 43042 693576 43110 693610
rect 43200 693576 43268 693610
rect 43358 693576 43426 693610
rect 43516 693576 43584 693610
rect 43674 693576 43742 693610
rect 43832 693576 43900 693610
rect 43990 693576 44058 693610
rect 44148 693576 44216 693610
rect 44306 693576 44374 693610
rect 44464 693576 44532 693610
rect 44622 693576 44690 693610
rect 44780 693576 44848 693610
rect 44938 693576 45006 693610
rect 45096 693576 45164 693610
rect 45254 693576 45322 693610
rect 45412 693576 45480 693610
rect 45570 693576 45638 693610
rect 45728 693576 45796 693610
rect 45886 693576 45954 693610
rect 46044 693576 46112 693610
rect 46202 693576 46270 693610
rect 42980 692541 43014 693517
rect 43138 692541 43172 693517
rect 43296 692541 43330 693517
rect 43454 692541 43488 693517
rect 43612 692541 43646 693517
rect 43770 692541 43804 693517
rect 43928 692541 43962 693517
rect 44086 692541 44120 693517
rect 44244 692541 44278 693517
rect 44402 692541 44436 693517
rect 44560 692541 44594 693517
rect 44718 692541 44752 693517
rect 44876 692541 44910 693517
rect 45034 692541 45068 693517
rect 45192 692541 45226 693517
rect 45350 692541 45384 693517
rect 45508 692541 45542 693517
rect 45666 692541 45700 693517
rect 45824 692541 45858 693517
rect 45982 692541 46016 693517
rect 46140 692541 46174 693517
rect 46298 692541 46332 693517
rect 43042 692448 43110 692482
rect 43200 692448 43268 692482
rect 43358 692448 43426 692482
rect 43516 692448 43584 692482
rect 43674 692448 43742 692482
rect 43832 692448 43900 692482
rect 43990 692448 44058 692482
rect 44148 692448 44216 692482
rect 44306 692448 44374 692482
rect 44464 692448 44532 692482
rect 44622 692448 44690 692482
rect 44780 692448 44848 692482
rect 44938 692448 45006 692482
rect 45096 692448 45164 692482
rect 45254 692448 45322 692482
rect 45412 692448 45480 692482
rect 45570 692448 45638 692482
rect 45728 692448 45796 692482
rect 45886 692448 45954 692482
rect 46044 692448 46112 692482
rect 46202 692448 46270 692482
rect 48781 693539 49178 694653
rect 51212 693539 51609 694653
rect 49950 693427 50130 693460
rect 50370 693427 50550 693460
rect 49950 693393 50130 693427
rect 50370 693393 50550 693427
rect 49950 693360 50130 693393
rect 50370 693360 50550 693393
rect 43640 692346 44210 692380
rect 45110 692346 45680 692380
rect 43640 692172 44210 692346
rect 45110 692172 45680 692346
rect 43640 692140 44210 692172
rect 45110 692140 45680 692172
rect 43042 692036 43110 692070
rect 43200 692036 43268 692070
rect 43358 692036 43426 692070
rect 43516 692036 43584 692070
rect 43674 692036 43742 692070
rect 43832 692036 43900 692070
rect 43990 692036 44058 692070
rect 44148 692036 44216 692070
rect 44306 692036 44374 692070
rect 44464 692036 44532 692070
rect 44622 692036 44690 692070
rect 44780 692036 44848 692070
rect 44938 692036 45006 692070
rect 45096 692036 45164 692070
rect 45254 692036 45322 692070
rect 45412 692036 45480 692070
rect 45570 692036 45638 692070
rect 45728 692036 45796 692070
rect 45886 692036 45954 692070
rect 46044 692036 46112 692070
rect 46202 692036 46270 692070
rect 42980 691001 43014 691977
rect 43138 691001 43172 691977
rect 43296 691001 43330 691977
rect 43454 691001 43488 691977
rect 43612 691001 43646 691977
rect 43770 691001 43804 691977
rect 43928 691001 43962 691977
rect 44086 691001 44120 691977
rect 44244 691001 44278 691977
rect 44402 691001 44436 691977
rect 44560 691001 44594 691977
rect 44718 691001 44752 691977
rect 44876 691001 44910 691977
rect 45034 691001 45068 691977
rect 45192 691001 45226 691977
rect 45350 691001 45384 691977
rect 45508 691001 45542 691977
rect 45666 691001 45700 691977
rect 45824 691001 45858 691977
rect 45982 691001 46016 691977
rect 46140 691001 46174 691977
rect 46298 691001 46332 691977
rect 43042 690908 43110 690942
rect 43200 690908 43268 690942
rect 43358 690908 43426 690942
rect 43516 690908 43584 690942
rect 43674 690908 43742 690942
rect 43832 690908 43900 690942
rect 43990 690908 44058 690942
rect 44148 690908 44216 690942
rect 44306 690908 44374 690942
rect 44464 690908 44532 690942
rect 44622 690908 44690 690942
rect 44780 690908 44848 690942
rect 44938 690908 45006 690942
rect 45096 690908 45164 690942
rect 45254 690908 45322 690942
rect 45412 690908 45480 690942
rect 45570 690908 45638 690942
rect 45728 690908 45796 690942
rect 45886 690908 45954 690942
rect 46044 690908 46112 690942
rect 46202 690908 46270 690942
rect 541969 690898 542059 690962
rect 542139 690898 542229 690962
rect 544459 690898 544549 690962
rect 544629 690898 544719 690962
rect 546919 690898 546999 690972
rect 547089 690898 547169 690972
rect 541969 690892 542059 690898
rect 542139 690892 542229 690898
rect 544459 690892 544549 690898
rect 544629 690892 544719 690898
rect 546919 690892 546999 690898
rect 547089 690892 547169 690898
rect 44326 690561 44976 690595
rect 44143 690459 44211 690493
rect 44301 690459 44369 690493
rect 44459 690459 44527 690493
rect 44617 690459 44685 690493
rect 44775 690459 44843 690493
rect 44933 690459 45001 690493
rect 45091 690459 45159 690493
rect 44081 689433 44115 690409
rect 44239 689433 44273 690409
rect 44397 689433 44431 690409
rect 44555 689433 44589 690409
rect 44713 689433 44747 690409
rect 44871 689433 44905 690409
rect 45029 689433 45063 690409
rect 45187 689433 45221 690409
rect 44143 689349 44211 689383
rect 44301 689349 44369 689383
rect 44459 689349 44527 689383
rect 44617 689349 44685 689383
rect 44775 689349 44843 689383
rect 44933 689349 45001 689383
rect 45091 689349 45159 689383
rect 540380 690750 541356 690784
rect 541616 690750 542592 690784
rect 542852 690750 543828 690784
rect 544088 690750 545064 690784
rect 545324 690750 546300 690784
rect 546560 690750 547536 690784
rect 547796 690750 548772 690784
rect 540287 690654 540321 690722
rect 541415 690654 541449 690722
rect 541523 690654 541557 690722
rect 542651 690654 542685 690722
rect 542759 690654 542793 690722
rect 543887 690654 543921 690722
rect 543995 690654 544029 690722
rect 545123 690654 545157 690722
rect 545231 690654 545265 690722
rect 546359 690654 546393 690722
rect 546467 690654 546501 690722
rect 547595 690654 547629 690722
rect 547703 690654 547737 690722
rect 548831 690654 548865 690722
rect 540380 690592 541356 690626
rect 541616 690592 542592 690626
rect 542852 690592 543828 690626
rect 544088 690592 545064 690626
rect 545324 690592 546300 690626
rect 546560 690592 547536 690626
rect 547796 690592 548772 690626
rect 540380 690210 541356 690244
rect 541616 690210 542592 690244
rect 542852 690210 543828 690244
rect 544088 690210 545064 690244
rect 545324 690210 546300 690244
rect 546560 690210 547536 690244
rect 547796 690210 548772 690244
rect 540287 690114 540321 690182
rect 541415 690114 541449 690182
rect 541523 690114 541557 690182
rect 542651 690114 542685 690182
rect 542759 690114 542793 690182
rect 543887 690114 543921 690182
rect 543995 690114 544029 690182
rect 545123 690114 545157 690182
rect 545231 690114 545265 690182
rect 546359 690114 546393 690182
rect 546467 690114 546501 690182
rect 547595 690114 547629 690182
rect 547703 690114 547737 690182
rect 548831 690114 548865 690182
rect 540380 690052 541356 690086
rect 541616 690052 542592 690086
rect 542852 690052 543828 690086
rect 544088 690052 545064 690086
rect 545324 690052 546300 690086
rect 546560 690052 547536 690086
rect 547796 690052 548772 690086
rect 541979 689842 542069 689912
rect 542119 689842 542209 689912
rect 544459 689842 544549 689912
rect 544619 689852 544709 689922
rect 546919 689852 546999 689922
rect 547089 689852 547169 689922
rect 540380 689670 541356 689704
rect 541616 689670 542592 689704
rect 542852 689670 543828 689704
rect 544088 689670 545064 689704
rect 545324 689670 546300 689704
rect 546560 689670 547536 689704
rect 547796 689670 548772 689704
rect 540287 689574 540321 689642
rect 541415 689574 541449 689642
rect 541523 689574 541557 689642
rect 542651 689574 542685 689642
rect 542759 689574 542793 689642
rect 543887 689574 543921 689642
rect 543995 689574 544029 689642
rect 545123 689574 545157 689642
rect 545231 689574 545265 689642
rect 546359 689574 546393 689642
rect 546467 689574 546501 689642
rect 547595 689574 547629 689642
rect 547703 689574 547737 689642
rect 548831 689574 548865 689642
rect 540380 689512 541356 689546
rect 541616 689512 542592 689546
rect 542852 689512 543828 689546
rect 544088 689512 545064 689546
rect 545324 689512 546300 689546
rect 546560 689512 547536 689546
rect 547796 689512 548772 689546
rect 44326 689247 44976 689281
rect 541979 689302 542059 689382
rect 542149 689302 542229 689382
rect 544459 689302 544539 689382
rect 544629 689302 544709 689382
rect 546919 689302 546999 689382
rect 547089 689302 547169 689382
rect 44326 689041 44976 689075
rect 44143 688939 44211 688973
rect 44301 688939 44369 688973
rect 44459 688939 44527 688973
rect 44617 688939 44685 688973
rect 44775 688939 44843 688973
rect 44933 688939 45001 688973
rect 45091 688939 45159 688973
rect 44081 687913 44115 688889
rect 44239 687913 44273 688889
rect 44397 687913 44431 688889
rect 44555 687913 44589 688889
rect 44713 687913 44747 688889
rect 44871 687913 44905 688889
rect 45029 687913 45063 688889
rect 45187 687913 45221 688889
rect 44143 687829 44211 687863
rect 44301 687829 44369 687863
rect 44459 687829 44527 687863
rect 44617 687829 44685 687863
rect 44775 687829 44843 687863
rect 44933 687829 45001 687863
rect 45091 687829 45159 687863
rect 540380 689130 541356 689164
rect 541616 689130 542592 689164
rect 542852 689130 543828 689164
rect 544088 689130 545064 689164
rect 545324 689130 546300 689164
rect 546560 689130 547536 689164
rect 547796 689130 548772 689164
rect 540287 689034 540321 689102
rect 541415 689034 541449 689102
rect 541523 689034 541557 689102
rect 542651 689034 542685 689102
rect 542759 689034 542793 689102
rect 543887 689034 543921 689102
rect 543995 689034 544029 689102
rect 545123 689034 545157 689102
rect 545231 689034 545265 689102
rect 546359 689034 546393 689102
rect 546467 689034 546501 689102
rect 547595 689034 547629 689102
rect 547703 689034 547737 689102
rect 548831 689034 548865 689102
rect 540380 688972 541356 689006
rect 541616 688972 542592 689006
rect 542852 688972 543828 689006
rect 544088 688972 545064 689006
rect 545324 688972 546300 689006
rect 546560 688972 547536 689006
rect 547796 688972 548772 689006
rect 540380 688550 541356 688584
rect 541616 688550 542592 688584
rect 542852 688550 543828 688584
rect 544088 688550 545064 688584
rect 545324 688550 546300 688584
rect 546560 688550 547536 688584
rect 547796 688550 548772 688584
rect 540287 688454 540321 688522
rect 541415 688454 541449 688522
rect 541523 688454 541557 688522
rect 542651 688454 542685 688522
rect 542759 688454 542793 688522
rect 543887 688454 543921 688522
rect 543995 688454 544029 688522
rect 545123 688454 545157 688522
rect 545231 688454 545265 688522
rect 546359 688454 546393 688522
rect 546467 688454 546501 688522
rect 547595 688454 547629 688522
rect 547703 688454 547737 688522
rect 548831 688454 548865 688522
rect 540380 688392 541356 688426
rect 541616 688392 542592 688426
rect 542852 688392 543828 688426
rect 544088 688392 545064 688426
rect 545324 688392 546300 688426
rect 546560 688392 547536 688426
rect 547796 688392 548772 688426
rect 541979 688142 542069 688222
rect 542139 688142 542229 688222
rect 544459 688142 544539 688212
rect 544629 688142 544709 688212
rect 546919 688142 546999 688212
rect 547089 688142 547169 688212
rect 44326 687727 44976 687761
rect 43833 687520 45477 687554
rect 43152 687418 43320 687452
rect 43410 687418 43578 687452
rect 43668 687418 43836 687452
rect 43926 687418 44094 687452
rect 44184 687418 44352 687452
rect 44442 687418 44610 687452
rect 44700 687418 44868 687452
rect 44958 687418 45126 687452
rect 45216 687418 45384 687452
rect 45474 687418 45642 687452
rect 45732 687418 45900 687452
rect 45990 687418 46158 687452
rect 43090 686392 43124 687368
rect 43348 686392 43382 687368
rect 43606 686392 43640 687368
rect 43864 686392 43898 687368
rect 44122 686392 44156 687368
rect 44380 686392 44414 687368
rect 44638 686392 44672 687368
rect 44896 686392 44930 687368
rect 45154 686392 45188 687368
rect 45412 686392 45446 687368
rect 45670 686392 45704 687368
rect 45928 686392 45962 687368
rect 46186 686392 46220 687368
rect 43152 686308 43320 686342
rect 43410 686308 43578 686342
rect 43668 686308 43836 686342
rect 43926 686308 44094 686342
rect 44184 686308 44352 686342
rect 44442 686308 44610 686342
rect 44700 686308 44868 686342
rect 44958 686308 45126 686342
rect 45216 686308 45384 686342
rect 45474 686308 45642 686342
rect 45732 686308 45900 686342
rect 45990 686308 46158 686342
rect 534740 686841 535137 687955
rect 537171 686841 537568 687955
rect 540380 687970 541356 688004
rect 541616 687970 542592 688004
rect 542852 687970 543828 688004
rect 544088 687970 545064 688004
rect 545324 687970 546300 688004
rect 546560 687970 547536 688004
rect 547796 687970 548772 688004
rect 540287 687874 540321 687942
rect 541415 687874 541449 687942
rect 541523 687874 541557 687942
rect 542651 687874 542685 687942
rect 542759 687874 542793 687942
rect 543887 687874 543921 687942
rect 543995 687874 544029 687942
rect 545123 687874 545157 687942
rect 545231 687874 545265 687942
rect 546359 687874 546393 687942
rect 546467 687874 546501 687942
rect 547595 687874 547629 687942
rect 547703 687874 547737 687942
rect 548831 687874 548865 687942
rect 540380 687812 541356 687846
rect 541616 687812 542592 687846
rect 542852 687812 543828 687846
rect 544088 687812 545064 687846
rect 545324 687812 546300 687846
rect 546560 687812 547536 687846
rect 547796 687812 548772 687846
rect 538540 687430 539516 687464
rect 539776 687430 540752 687464
rect 541012 687430 541988 687464
rect 542248 687430 543224 687464
rect 543484 687430 544460 687464
rect 544720 687430 545696 687464
rect 545956 687430 546932 687464
rect 547192 687430 548168 687464
rect 548428 687430 549404 687464
rect 549664 687430 550640 687464
rect 538447 687334 538481 687402
rect 539575 687334 539609 687402
rect 539683 687334 539717 687402
rect 540811 687334 540845 687402
rect 540919 687334 540953 687402
rect 542047 687334 542081 687402
rect 542155 687334 542189 687402
rect 543283 687334 543317 687402
rect 543391 687334 543425 687402
rect 544519 687334 544553 687402
rect 544627 687334 544661 687402
rect 545755 687334 545789 687402
rect 545863 687334 545897 687402
rect 546991 687334 547025 687402
rect 547099 687334 547133 687402
rect 548227 687334 548261 687402
rect 548335 687334 548369 687402
rect 549463 687334 549497 687402
rect 549571 687334 549605 687402
rect 550699 687334 550733 687402
rect 538540 687272 539516 687306
rect 539776 687272 540752 687306
rect 541012 687272 541988 687306
rect 542248 687272 543224 687306
rect 543484 687272 544460 687306
rect 544720 687272 545696 687306
rect 545956 687272 546932 687306
rect 547192 687272 548168 687306
rect 548428 687272 549404 687306
rect 549664 687272 550640 687306
rect 540119 687062 540209 687142
rect 540299 687062 540389 687142
rect 542649 687062 542739 687142
rect 542809 687062 542899 687142
rect 545119 687062 545209 687142
rect 545279 687062 545369 687142
rect 547569 687062 547659 687142
rect 547729 687062 547819 687142
rect 550069 687062 550159 687142
rect 550229 687062 550319 687142
rect 538540 686890 539516 686924
rect 539776 686890 540752 686924
rect 541012 686890 541988 686924
rect 542248 686890 543224 686924
rect 543484 686890 544460 686924
rect 544720 686890 545696 686924
rect 545956 686890 546932 686924
rect 547192 686890 548168 686924
rect 548428 686890 549404 686924
rect 549664 686890 550640 686924
rect 538447 686794 538481 686862
rect 539575 686794 539609 686862
rect 539683 686794 539717 686862
rect 540811 686794 540845 686862
rect 540919 686794 540953 686862
rect 542047 686794 542081 686862
rect 542155 686794 542189 686862
rect 543283 686794 543317 686862
rect 543391 686794 543425 686862
rect 544519 686794 544553 686862
rect 544627 686794 544661 686862
rect 545755 686794 545789 686862
rect 545863 686794 545897 686862
rect 546991 686794 547025 686862
rect 547099 686794 547133 686862
rect 548227 686794 548261 686862
rect 548335 686794 548369 686862
rect 549463 686794 549497 686862
rect 549571 686794 549605 686862
rect 550699 686794 550733 686862
rect 538540 686732 539516 686766
rect 539776 686732 540752 686766
rect 541012 686732 541988 686766
rect 542248 686732 543224 686766
rect 543484 686732 544460 686766
rect 544720 686732 545696 686766
rect 545956 686732 546932 686766
rect 547192 686732 548168 686766
rect 548428 686732 549404 686766
rect 549664 686732 550640 686766
rect 551800 686841 552197 687955
rect 554231 686841 554628 687955
rect 43833 686206 45477 686240
rect 43702 686000 45604 686034
rect 42892 685898 43060 685932
rect 43150 685898 43318 685932
rect 43408 685898 43576 685932
rect 43666 685898 43834 685932
rect 43924 685898 44092 685932
rect 44182 685898 44350 685932
rect 44440 685898 44608 685932
rect 44698 685898 44866 685932
rect 44956 685898 45124 685932
rect 45214 685898 45382 685932
rect 45472 685898 45640 685932
rect 45730 685898 45898 685932
rect 45988 685898 46156 685932
rect 46246 685898 46414 685932
rect 42830 684872 42864 685848
rect 43088 684872 43122 685848
rect 43346 684872 43380 685848
rect 43604 684872 43638 685848
rect 43862 684872 43896 685848
rect 44120 684872 44154 685848
rect 44378 684872 44412 685848
rect 44636 684872 44670 685848
rect 44894 684872 44928 685848
rect 45152 684872 45186 685848
rect 45410 684872 45444 685848
rect 45668 684872 45702 685848
rect 45926 684872 45960 685848
rect 46184 684872 46218 685848
rect 46442 684872 46476 685848
rect 42892 684788 43060 684822
rect 43150 684788 43318 684822
rect 43408 684788 43576 684822
rect 43666 684788 43834 684822
rect 43924 684788 44092 684822
rect 44182 684788 44350 684822
rect 44440 684788 44608 684822
rect 44698 684788 44866 684822
rect 44956 684788 45124 684822
rect 45214 684788 45382 684822
rect 45472 684788 45640 684822
rect 45730 684788 45898 684822
rect 45988 684788 46156 684822
rect 46246 684788 46414 684822
rect 534740 685371 535137 686485
rect 537171 685371 537568 686485
rect 538540 686350 539516 686384
rect 539776 686350 540752 686384
rect 541012 686350 541988 686384
rect 542248 686350 543224 686384
rect 543484 686350 544460 686384
rect 544720 686350 545696 686384
rect 545956 686350 546932 686384
rect 547192 686350 548168 686384
rect 548428 686350 549404 686384
rect 549664 686350 550640 686384
rect 538447 686254 538481 686322
rect 539575 686254 539609 686322
rect 539683 686254 539717 686322
rect 540811 686254 540845 686322
rect 540919 686254 540953 686322
rect 542047 686254 542081 686322
rect 542155 686254 542189 686322
rect 543283 686254 543317 686322
rect 543391 686254 543425 686322
rect 544519 686254 544553 686322
rect 544627 686254 544661 686322
rect 545755 686254 545789 686322
rect 545863 686254 545897 686322
rect 546991 686254 547025 686322
rect 547099 686254 547133 686322
rect 548227 686254 548261 686322
rect 548335 686254 548369 686322
rect 549463 686254 549497 686322
rect 549571 686254 549605 686322
rect 550699 686254 550733 686322
rect 538540 686192 539516 686226
rect 539776 686192 540752 686226
rect 541012 686192 541988 686226
rect 542248 686192 543224 686226
rect 543484 686192 544460 686226
rect 544720 686192 545696 686226
rect 545956 686192 546932 686226
rect 547192 686192 548168 686226
rect 548428 686192 549404 686226
rect 549664 686192 550640 686226
rect 540119 685982 540209 686062
rect 540299 685992 540389 686072
rect 542649 685982 542739 686062
rect 542809 685982 542899 686062
rect 545119 685982 545209 686062
rect 545279 685982 545369 686062
rect 547569 685982 547659 686062
rect 547729 685982 547819 686062
rect 550069 685982 550159 686062
rect 550229 685982 550319 686062
rect 538540 685810 539516 685844
rect 539776 685810 540752 685844
rect 541012 685810 541988 685844
rect 542248 685810 543224 685844
rect 543484 685810 544460 685844
rect 544720 685810 545696 685844
rect 545956 685810 546932 685844
rect 547192 685810 548168 685844
rect 548428 685810 549404 685844
rect 549664 685810 550640 685844
rect 538447 685714 538481 685782
rect 539575 685714 539609 685782
rect 539683 685714 539717 685782
rect 540811 685714 540845 685782
rect 540919 685714 540953 685782
rect 542047 685714 542081 685782
rect 542155 685714 542189 685782
rect 543283 685714 543317 685782
rect 543391 685714 543425 685782
rect 544519 685714 544553 685782
rect 544627 685714 544661 685782
rect 545755 685714 545789 685782
rect 545863 685714 545897 685782
rect 546991 685714 547025 685782
rect 547099 685714 547133 685782
rect 548227 685714 548261 685782
rect 548335 685714 548369 685782
rect 549463 685714 549497 685782
rect 549571 685714 549605 685782
rect 550699 685714 550733 685782
rect 538540 685652 539516 685686
rect 539776 685652 540752 685686
rect 541012 685652 541988 685686
rect 542248 685652 543224 685686
rect 543484 685652 544460 685686
rect 544720 685652 545696 685686
rect 545956 685652 546932 685686
rect 547192 685652 548168 685686
rect 548428 685652 549404 685686
rect 549664 685652 550640 685686
rect 535759 685225 535849 685252
rect 535969 685225 536059 685252
rect 551800 685371 552197 686485
rect 554231 685371 554628 686485
rect 553069 685225 553139 685242
rect 553229 685225 553299 685242
rect 535759 685122 535849 685225
rect 535969 685122 536059 685225
rect 553069 685152 553139 685225
rect 553229 685152 553299 685225
rect 540471 685030 541447 685064
rect 541689 685030 542665 685064
rect 542907 685030 543883 685064
rect 544125 685030 545101 685064
rect 545343 685030 546319 685064
rect 546561 685030 547537 685064
rect 547779 685030 548755 685064
rect 540387 684934 540421 685002
rect 541497 684934 541531 685002
rect 541605 684934 541639 685002
rect 542715 684934 542749 685002
rect 542823 684934 542857 685002
rect 543933 684934 543967 685002
rect 544041 684934 544075 685002
rect 545151 684934 545185 685002
rect 545259 684934 545293 685002
rect 546369 684934 546403 685002
rect 546477 684934 546511 685002
rect 547587 684934 547621 685002
rect 547695 684934 547729 685002
rect 548805 684934 548839 685002
rect 540471 684872 541447 684906
rect 541689 684872 542665 684906
rect 542907 684872 543883 684906
rect 544125 684872 545101 684906
rect 545343 684872 546319 684906
rect 546561 684872 547537 684906
rect 547779 684872 548755 684906
rect 542279 684758 542389 684772
rect 543139 684758 543249 684772
rect 544349 684758 544459 684772
rect 545199 684758 545309 684772
rect 546769 684758 546879 684772
rect 547649 684758 547759 684772
rect 43702 684686 45604 684720
rect 542279 684678 542389 684758
rect 543139 684678 543249 684758
rect 544349 684678 544459 684758
rect 545199 684678 545309 684758
rect 546769 684678 546879 684758
rect 547649 684678 547759 684758
rect 542279 684662 542389 684678
rect 543139 684662 543249 684678
rect 544349 684662 544459 684678
rect 545199 684662 545309 684678
rect 546769 684662 546879 684678
rect 547649 684662 547759 684678
rect 540471 684530 541447 684564
rect 541689 684530 542665 684564
rect 542907 684530 543883 684564
rect 544125 684530 545101 684564
rect 545343 684530 546319 684564
rect 546561 684530 547537 684564
rect 547779 684530 548755 684564
rect 540387 684434 540421 684502
rect 541497 684434 541531 684502
rect 541605 684434 541639 684502
rect 542715 684434 542749 684502
rect 542823 684434 542857 684502
rect 543933 684434 543967 684502
rect 544041 684434 544075 684502
rect 545151 684434 545185 684502
rect 545259 684434 545293 684502
rect 546369 684434 546403 684502
rect 546477 684434 546511 684502
rect 547587 684434 547621 684502
rect 547695 684434 547729 684502
rect 548805 684434 548839 684502
rect 540471 684372 541447 684406
rect 541689 684372 542665 684406
rect 542907 684372 543883 684406
rect 544125 684372 545101 684406
rect 545343 684372 546319 684406
rect 546561 684372 547537 684406
rect 547779 684372 548755 684406
rect 43922 683866 44090 683900
rect 44180 683866 44348 683900
rect 44438 683866 44606 683900
rect 44696 683866 44864 683900
rect 44954 683866 45122 683900
rect 45212 683866 45380 683900
rect 43740 683200 43746 683430
rect 43746 683200 43780 683430
rect 43860 682831 43894 683807
rect 44118 682831 44152 683807
rect 44376 682831 44410 683807
rect 44634 682831 44668 683807
rect 44892 682831 44926 683807
rect 45150 682831 45184 683807
rect 45408 682831 45442 683807
rect 541031 684030 542007 684064
rect 542249 684030 543225 684064
rect 543467 684030 544443 684064
rect 544685 684030 545661 684064
rect 545903 684030 546879 684064
rect 547121 684030 548097 684064
rect 540947 683834 540981 684002
rect 542057 683834 542091 684002
rect 542165 683834 542199 684002
rect 543275 683834 543309 684002
rect 543383 683834 543417 684002
rect 544493 683834 544527 684002
rect 544601 683834 544635 684002
rect 545711 683834 545745 684002
rect 545819 683834 545853 684002
rect 546929 683834 546963 684002
rect 547037 683834 547071 684002
rect 548147 683834 548181 684002
rect 541031 683772 542007 683806
rect 542249 683772 543225 683806
rect 543467 683772 544443 683806
rect 544685 683772 545661 683806
rect 545903 683772 546879 683806
rect 547121 683772 548097 683806
rect 541569 683562 541679 683652
rect 546479 683562 546589 683652
rect 45520 683200 45522 683430
rect 45522 683200 45556 683430
rect 45556 683200 45560 683430
rect 43922 682738 44090 682772
rect 44180 682738 44348 682772
rect 44438 682738 44606 682772
rect 44696 682738 44864 682772
rect 44954 682738 45122 682772
rect 45212 682738 45380 682772
rect 541031 683410 542007 683444
rect 542249 683410 543225 683444
rect 543467 683410 544443 683444
rect 544685 683410 545661 683444
rect 545903 683410 546879 683444
rect 547121 683410 548097 683444
rect 540947 683214 540981 683382
rect 542057 683214 542091 683382
rect 542165 683214 542199 683382
rect 543275 683214 543309 683382
rect 543383 683214 543417 683382
rect 544493 683214 544527 683382
rect 544601 683214 544635 683382
rect 545711 683214 545745 683382
rect 545819 683214 545853 683382
rect 546929 683214 546963 683382
rect 547037 683214 547071 683382
rect 548147 683214 548181 683382
rect 541031 683152 542007 683186
rect 542249 683152 543225 683186
rect 543467 683152 544443 683186
rect 544685 683152 545661 683186
rect 545903 683152 546879 683186
rect 547121 683152 548097 683186
rect 540471 682810 541447 682844
rect 541689 682810 542665 682844
rect 542907 682810 543883 682844
rect 544125 682810 545101 682844
rect 545343 682810 546319 682844
rect 546561 682810 547537 682844
rect 547779 682810 548755 682844
rect 540387 682614 540421 682782
rect 541497 682614 541531 682782
rect 541605 682614 541639 682782
rect 542715 682614 542749 682782
rect 542823 682614 542857 682782
rect 543933 682614 543967 682782
rect 544041 682614 544075 682782
rect 545151 682614 545185 682782
rect 545259 682614 545293 682782
rect 546369 682614 546403 682782
rect 546477 682614 546511 682782
rect 547587 682614 547621 682782
rect 547695 682614 547729 682782
rect 548805 682614 548839 682782
rect 540471 682552 541447 682586
rect 541689 682552 542665 682586
rect 542907 682552 543883 682586
rect 544125 682552 545101 682586
rect 545343 682552 546319 682586
rect 546561 682552 547537 682586
rect 547779 682552 548755 682586
rect 541509 682438 541629 682452
rect 542729 682438 542849 682452
rect 543939 682438 544059 682452
rect 545159 682438 545279 682452
rect 546389 682438 546509 682442
rect 547599 682438 547719 682452
rect 43922 682366 44090 682400
rect 44180 682366 44348 682400
rect 44438 682366 44606 682400
rect 44696 682366 44864 682400
rect 44954 682366 45122 682400
rect 45212 682366 45380 682400
rect 43740 681690 43746 681920
rect 43746 681690 43780 681920
rect 43860 681331 43894 682307
rect 44118 681331 44152 682307
rect 44376 681331 44410 682307
rect 44634 681331 44668 682307
rect 44892 681331 44926 682307
rect 45150 681331 45184 682307
rect 45408 681331 45442 682307
rect 541509 682358 541629 682438
rect 542729 682358 542849 682438
rect 543939 682358 544059 682438
rect 545159 682358 545279 682438
rect 546389 682358 546509 682438
rect 547599 682358 547719 682438
rect 541509 682352 541629 682358
rect 542729 682352 542849 682358
rect 543939 682352 544059 682358
rect 545159 682352 545279 682358
rect 546389 682342 546509 682358
rect 547599 682352 547719 682358
rect 540471 682210 541447 682244
rect 541689 682210 542665 682244
rect 542907 682210 543883 682244
rect 544125 682210 545101 682244
rect 545343 682210 546319 682244
rect 546561 682210 547537 682244
rect 547779 682210 548755 682244
rect 540387 682014 540421 682182
rect 541497 682014 541531 682182
rect 541605 682014 541639 682182
rect 542715 682014 542749 682182
rect 542823 682014 542857 682182
rect 543933 682014 543967 682182
rect 544041 682014 544075 682182
rect 545151 682014 545185 682182
rect 545259 682014 545293 682182
rect 546369 682014 546403 682182
rect 546477 682014 546511 682182
rect 547587 682014 547621 682182
rect 547695 682014 547729 682182
rect 548805 682014 548839 682182
rect 540471 681952 541447 681986
rect 541689 681952 542665 681986
rect 542907 681952 543883 681986
rect 544125 681952 545101 681986
rect 545343 681952 546319 681986
rect 546561 681952 547537 681986
rect 547779 681952 548755 681986
rect 45520 681690 45522 681920
rect 45522 681690 45556 681920
rect 45556 681690 45560 681920
rect 44420 681272 44582 681274
rect 43922 681238 44090 681272
rect 44180 681238 44348 681272
rect 44420 681238 44438 681272
rect 44438 681238 44606 681272
rect 44696 681238 44864 681272
rect 44954 681238 45122 681272
rect 45212 681238 45380 681272
rect 44420 681234 44582 681238
rect 541384 681384 541544 681478
rect 542444 681384 542604 681478
rect 543904 681384 544064 681478
rect 545124 681384 545284 681478
rect 546604 681384 546764 681478
rect 547604 681384 547764 681478
rect 541384 681350 541544 681384
rect 542444 681350 542604 681384
rect 543904 681350 544064 681384
rect 545124 681350 545284 681384
rect 546604 681350 546764 681384
rect 547604 681350 547764 681384
rect 541384 681318 541544 681350
rect 542444 681318 542604 681350
rect 543904 681318 544064 681350
rect 545124 681318 545284 681350
rect 546604 681318 546764 681350
rect 547604 681318 547764 681350
rect 541025 681236 542001 681270
rect 542261 681236 543237 681270
rect 543497 681236 544473 681270
rect 544733 681236 545709 681270
rect 545969 681236 546945 681270
rect 547205 681236 548181 681270
rect 540932 681040 540966 681208
rect 542060 681040 542094 681208
rect 542168 681040 542202 681208
rect 543296 681040 543330 681208
rect 543404 681040 543438 681208
rect 544532 681040 544566 681208
rect 544640 681040 544674 681208
rect 545768 681040 545802 681208
rect 545876 681040 545910 681208
rect 547004 681040 547038 681208
rect 547112 681040 547146 681208
rect 548240 681040 548274 681208
rect 541025 680978 542001 681012
rect 542261 680978 543237 681012
rect 543497 680978 544473 681012
rect 544733 680978 545709 681012
rect 545969 680978 546945 681012
rect 547205 680978 548181 681012
rect 541384 680864 541544 680898
rect 542444 680864 542604 680898
rect 543904 680864 544064 680898
rect 545124 680864 545284 680898
rect 546604 680864 546764 680898
rect 547604 680864 547764 680898
rect 541384 680794 541544 680864
rect 542444 680794 542604 680864
rect 543904 680794 544064 680864
rect 545124 680794 545284 680864
rect 546604 680794 546764 680864
rect 547604 680794 547764 680864
rect 44522 680748 44590 680782
rect 44680 680748 44748 680782
rect 44340 680350 44346 680580
rect 44346 680350 44380 680580
rect 44460 680222 44494 680698
rect 44618 680222 44652 680698
rect 44776 680222 44810 680698
rect 541384 680760 541544 680794
rect 542444 680760 542604 680794
rect 543904 680760 544064 680794
rect 545124 680760 545284 680794
rect 546604 680760 546764 680794
rect 547604 680760 547764 680794
rect 541384 680738 541544 680760
rect 542444 680738 542604 680760
rect 543904 680738 544064 680760
rect 545124 680738 545284 680760
rect 546604 680738 546764 680760
rect 547604 680738 547764 680760
rect 44890 680350 44924 680580
rect 44924 680350 44930 680580
rect 541025 680646 542001 680680
rect 542261 680646 543237 680680
rect 543497 680646 544473 680680
rect 544733 680646 545709 680680
rect 545969 680646 546945 680680
rect 547205 680646 548181 680680
rect 540932 680450 540966 680618
rect 542060 680450 542094 680618
rect 542168 680450 542202 680618
rect 543296 680450 543330 680618
rect 543404 680450 543438 680618
rect 544532 680450 544566 680618
rect 544640 680450 544674 680618
rect 545768 680450 545802 680618
rect 545876 680450 545910 680618
rect 547004 680450 547038 680618
rect 547112 680450 547146 680618
rect 548240 680450 548274 680618
rect 541025 680388 542001 680422
rect 542261 680388 543237 680422
rect 543497 680388 544473 680422
rect 544733 680388 545709 680422
rect 545969 680388 546945 680422
rect 547205 680388 548181 680422
rect 44522 680138 44590 680172
rect 44680 680138 44748 680172
rect 44162 679748 44330 679782
rect 44420 679748 44588 679782
rect 44678 679748 44846 679782
rect 44936 679748 45104 679782
rect 43960 679540 43986 679630
rect 43986 679540 44020 679630
rect 44020 679540 44050 679630
rect 44100 679472 44134 679698
rect 44358 679472 44392 679698
rect 44616 679472 44650 679698
rect 44874 679472 44908 679698
rect 45132 679472 45166 679698
rect 45220 679550 45246 679630
rect 45246 679550 45280 679630
rect 45280 679550 45300 679630
rect 543786 679856 544012 679890
rect 544254 679856 544480 679890
rect 544722 679856 544948 679890
rect 545190 679856 545416 679890
rect 543702 679660 543736 679828
rect 544062 679660 544096 679828
rect 544170 679660 544204 679828
rect 544530 679660 544564 679828
rect 544638 679660 544672 679828
rect 544998 679660 545032 679828
rect 545106 679660 545140 679828
rect 545466 679660 545500 679828
rect 543786 679598 544012 679632
rect 544254 679598 544480 679632
rect 544722 679598 544948 679632
rect 545190 679598 545416 679632
rect 44162 679388 44330 679422
rect 44420 679388 44588 679422
rect 44678 679388 44846 679422
rect 44936 679388 45104 679422
rect 543764 679484 543984 679518
rect 544284 679484 544504 679518
rect 544704 679484 544924 679518
rect 545254 679484 545474 679518
rect 543764 679379 543984 679484
rect 544284 679379 544504 679484
rect 544704 679379 544924 679484
rect 545254 679379 545474 679484
rect 543764 679368 543916 679379
rect 543916 679368 543984 679379
rect 544284 679368 544504 679379
rect 544704 679368 544924 679379
rect 545254 679368 545290 679379
rect 545290 679368 545474 679379
rect 44500 679286 44740 679320
rect 44500 679280 44740 679286
rect 44500 679134 44740 679140
rect 44500 679100 44740 679134
rect 43907 678998 44075 679032
rect 44165 678998 44333 679032
rect 44423 678998 44591 679032
rect 44681 678998 44849 679032
rect 44939 678998 45107 679032
rect 45197 678998 45365 679032
rect 43845 677972 43879 678948
rect 44103 677972 44137 678948
rect 44361 677972 44395 678948
rect 44619 677972 44653 678948
rect 44877 677972 44911 678948
rect 45135 677972 45169 678948
rect 45393 677972 45427 678948
rect 43907 677888 44075 677922
rect 44165 677888 44333 677922
rect 44423 677888 44591 677922
rect 44681 677888 44849 677922
rect 44939 677888 45107 677922
rect 45197 677888 45365 677922
rect 544006 679231 544482 679265
rect 544724 679231 545200 679265
rect 543922 679135 543956 679203
rect 544532 679135 544566 679203
rect 544640 679135 544674 679203
rect 545250 679135 545284 679203
rect 544006 679073 544482 679107
rect 544724 679073 545200 679107
rect 541404 678854 541584 678958
rect 542544 678854 542724 678958
rect 543524 678854 543704 678968
rect 544294 678959 544474 678968
rect 544734 678959 544914 678968
rect 544294 678854 544474 678959
rect 544734 678854 544914 678959
rect 545454 678854 545634 678958
rect 546524 678854 546704 678968
rect 547524 678854 547704 678968
rect 541404 678828 541584 678854
rect 542544 678828 542724 678854
rect 543524 678838 543704 678854
rect 544294 678838 544474 678854
rect 544734 678838 544914 678854
rect 545454 678828 545634 678854
rect 546524 678838 546704 678854
rect 547524 678838 547704 678854
rect 541071 678706 542047 678740
rect 542289 678706 543265 678740
rect 543507 678706 544483 678740
rect 544725 678706 545701 678740
rect 545943 678706 546919 678740
rect 547161 678706 548137 678740
rect 540987 678510 541021 678678
rect 542097 678510 542131 678678
rect 542205 678510 542239 678678
rect 543315 678510 543349 678678
rect 543423 678510 543457 678678
rect 544533 678510 544567 678678
rect 544641 678510 544675 678678
rect 545751 678510 545785 678678
rect 545859 678510 545893 678678
rect 546969 678510 547003 678678
rect 547077 678510 547111 678678
rect 548187 678510 548221 678678
rect 541071 678448 542047 678482
rect 542289 678448 543265 678482
rect 543507 678448 544483 678482
rect 544725 678448 545701 678482
rect 545943 678448 546919 678482
rect 547161 678448 548137 678482
rect 44500 677786 44740 677820
rect 44500 677780 44740 677786
rect 541777 677587 542891 677984
rect 543297 677587 544411 677984
rect 544807 677593 545921 677990
rect 546317 677593 547431 677990
rect 41738 677129 42852 677526
rect 43288 677129 44402 677526
rect 44828 677129 45942 677526
rect 46378 677129 47492 677526
rect 41200 676740 41440 676980
rect 47900 676740 48140 676980
rect 541364 676938 541484 677058
rect 547734 676938 547854 677058
rect 41200 675020 41440 675260
rect 47900 675020 48140 675260
rect 541364 673938 541484 674058
rect 547734 673938 547854 674058
rect 41200 673300 41440 673540
rect 47900 673300 48140 673540
rect 41200 671820 41440 672060
rect 47900 671820 48140 672060
rect 541364 670938 541484 671058
rect 547734 670938 547854 671058
rect 41200 670100 41440 670340
rect 47900 670100 48140 670340
rect 41200 668500 41440 668740
rect 47900 668500 48140 668740
rect 541364 667938 541484 668058
rect 547734 667938 547854 668058
rect 41200 666780 41440 667020
rect 47900 666780 48140 667020
rect 41200 665180 41440 665420
rect 47900 665180 48140 665420
rect 541364 664938 541484 665058
rect 547734 664938 547854 665058
rect 41200 663460 41440 663700
rect 47900 663460 48140 663700
rect 541777 663356 542891 663753
rect 543297 663356 544411 663753
rect 544807 663362 545921 663759
rect 546317 663362 547431 663759
rect 41738 662898 42852 663295
rect 43288 662898 44402 663295
rect 44828 662898 45942 663295
rect 46378 662898 47492 663295
<< metal1 >>
rect 37690 696113 38130 696130
rect 37690 694999 37711 696113
rect 38108 694999 38130 696113
rect 37690 694940 38130 694999
rect 36800 694920 38130 694940
rect 36800 694850 36930 694920
rect 37000 694850 38130 694920
rect 36800 694810 38130 694850
rect 36800 694740 36820 694810
rect 36890 694740 38130 694810
rect 36800 694720 38130 694740
rect 37690 694653 38130 694720
rect 37690 693539 37711 694653
rect 38108 693539 38130 694653
rect 37690 693520 38130 693539
rect 40120 696113 40560 696140
rect 40120 694999 40142 696113
rect 40539 694999 40560 696113
rect 48760 696113 49190 696130
rect 43980 695640 45360 695690
rect 43980 695388 44010 695640
rect 43017 695382 44010 695388
rect 44280 695382 45060 695640
rect 45330 695388 45360 695640
rect 45330 695382 46297 695388
rect 43017 695348 43029 695382
rect 46285 695348 46297 695382
rect 43017 695342 46297 695348
rect 40120 694860 40560 694999
rect 41330 695280 47990 695290
rect 41330 695246 41542 695280
rect 41610 695246 41700 695280
rect 41768 695246 41858 695280
rect 41926 695246 42016 695280
rect 42084 695246 42174 695280
rect 42242 695246 42332 695280
rect 42400 695246 42490 695280
rect 42558 695246 42648 695280
rect 42716 695246 42806 695280
rect 42874 695246 42964 695280
rect 43032 695246 43122 695280
rect 43190 695246 43280 695280
rect 43348 695246 43438 695280
rect 43506 695246 43596 695280
rect 43664 695246 43754 695280
rect 43822 695246 43912 695280
rect 43980 695246 44070 695280
rect 44138 695246 44228 695280
rect 44296 695246 44386 695280
rect 44454 695246 44544 695280
rect 44612 695246 44702 695280
rect 44770 695246 44860 695280
rect 44928 695246 45018 695280
rect 45086 695246 45176 695280
rect 45244 695246 45334 695280
rect 45402 695246 45492 695280
rect 45560 695246 45650 695280
rect 45718 695246 45808 695280
rect 45876 695246 45966 695280
rect 46034 695246 46124 695280
rect 46192 695246 46282 695280
rect 46350 695246 46440 695280
rect 46508 695246 46598 695280
rect 46666 695246 46756 695280
rect 46824 695246 46914 695280
rect 46982 695246 47072 695280
rect 47140 695246 47230 695280
rect 47298 695246 47388 695280
rect 47456 695246 47546 695280
rect 47614 695246 47704 695280
rect 47772 695246 47990 695280
rect 41330 695240 47990 695246
rect 41330 694860 41410 695240
rect 41474 695187 41520 695199
rect 41474 695160 41480 695187
rect 41514 695160 41520 695187
rect 41632 695187 41678 695199
rect 41450 695090 41460 695160
rect 41530 695090 41540 695160
rect 41474 694920 41480 695090
rect 41514 694920 41520 695090
rect 40120 694653 41410 694860
rect 41450 694850 41460 694920
rect 41530 694850 41540 694920
rect 40120 693539 40142 694653
rect 40539 694570 41410 694653
rect 40539 693539 40560 694570
rect 41330 694160 41410 694570
rect 41474 694211 41480 694850
rect 41514 694211 41520 694850
rect 41632 694550 41638 695187
rect 41672 694550 41678 695187
rect 41790 695187 41836 695199
rect 41790 695160 41796 695187
rect 41830 695160 41836 695187
rect 41948 695187 41994 695199
rect 41770 695090 41780 695160
rect 41850 695090 41860 695160
rect 41790 694920 41796 695090
rect 41830 694920 41836 695090
rect 41770 694850 41780 694920
rect 41850 694850 41860 694920
rect 41610 694480 41620 694550
rect 41690 694480 41700 694550
rect 41632 694310 41638 694480
rect 41672 694310 41678 694480
rect 41610 694240 41620 694310
rect 41690 694240 41700 694310
rect 41474 694199 41520 694211
rect 41632 694211 41638 694240
rect 41672 694211 41678 694240
rect 41632 694199 41678 694211
rect 41790 694211 41796 694850
rect 41830 694211 41836 694850
rect 41948 694550 41954 695187
rect 41988 694550 41994 695187
rect 42106 695187 42152 695199
rect 42106 695160 42112 695187
rect 42146 695160 42152 695187
rect 42264 695187 42310 695199
rect 42080 695090 42090 695160
rect 42160 695090 42170 695160
rect 42106 694920 42112 695090
rect 42146 694920 42152 695090
rect 42080 694850 42090 694920
rect 42160 694850 42170 694920
rect 41920 694480 41930 694550
rect 42000 694480 42010 694550
rect 41948 694310 41954 694480
rect 41988 694310 41994 694480
rect 41920 694240 41930 694310
rect 42000 694240 42010 694310
rect 41790 694199 41836 694211
rect 41948 694211 41954 694240
rect 41988 694211 41994 694240
rect 41948 694199 41994 694211
rect 42106 694211 42112 694850
rect 42146 694211 42152 694850
rect 42264 694550 42270 695187
rect 42304 694550 42310 695187
rect 42422 695187 42468 695199
rect 42422 695160 42428 695187
rect 42462 695160 42468 695187
rect 42580 695187 42626 695199
rect 42400 695090 42410 695160
rect 42480 695090 42490 695160
rect 42422 694920 42428 695090
rect 42462 694920 42468 695090
rect 42400 694850 42410 694920
rect 42480 694850 42490 694920
rect 42240 694480 42250 694550
rect 42320 694480 42330 694550
rect 42264 694310 42270 694480
rect 42304 694310 42310 694480
rect 42240 694240 42250 694310
rect 42320 694240 42330 694310
rect 42106 694199 42152 694211
rect 42264 694211 42270 694240
rect 42304 694211 42310 694240
rect 42264 694199 42310 694211
rect 42422 694211 42428 694850
rect 42462 694211 42468 694850
rect 42580 694550 42586 695187
rect 42620 694550 42626 695187
rect 42738 695187 42784 695199
rect 42738 695160 42744 695187
rect 42778 695160 42784 695187
rect 42896 695187 42942 695199
rect 42710 695090 42720 695160
rect 42790 695090 42800 695160
rect 42738 694920 42744 695090
rect 42778 694920 42784 695090
rect 42710 694850 42720 694920
rect 42790 694850 42800 694920
rect 42560 694480 42570 694550
rect 42640 694480 42650 694550
rect 42580 694310 42586 694480
rect 42620 694310 42626 694480
rect 42560 694240 42570 694310
rect 42640 694240 42650 694310
rect 42422 694199 42468 694211
rect 42580 694211 42586 694240
rect 42620 694211 42626 694240
rect 42580 694199 42626 694211
rect 42738 694211 42744 694850
rect 42778 694211 42784 694850
rect 42896 694550 42902 695187
rect 42936 694550 42942 695187
rect 43054 695187 43100 695199
rect 43054 695160 43060 695187
rect 43094 695160 43100 695187
rect 43212 695187 43258 695199
rect 43030 695090 43040 695160
rect 43110 695090 43120 695160
rect 43054 694920 43060 695090
rect 43094 694920 43100 695090
rect 43030 694850 43040 694920
rect 43110 694850 43120 694920
rect 42870 694480 42880 694550
rect 42950 694480 42960 694550
rect 42896 694310 42902 694480
rect 42936 694310 42942 694480
rect 42870 694240 42880 694310
rect 42950 694240 42960 694310
rect 42738 694199 42784 694211
rect 42896 694211 42902 694240
rect 42936 694211 42942 694240
rect 42896 694199 42942 694211
rect 43054 694211 43060 694850
rect 43094 694211 43100 694850
rect 43212 694550 43218 695187
rect 43252 694550 43258 695187
rect 43370 695187 43416 695199
rect 43370 695160 43376 695187
rect 43410 695160 43416 695187
rect 43528 695187 43574 695199
rect 43350 695090 43360 695160
rect 43430 695090 43440 695160
rect 43370 694920 43376 695090
rect 43410 694920 43416 695090
rect 43350 694850 43360 694920
rect 43430 694850 43440 694920
rect 43190 694480 43200 694550
rect 43270 694480 43280 694550
rect 43212 694310 43218 694480
rect 43252 694310 43258 694480
rect 43190 694240 43200 694310
rect 43270 694240 43280 694310
rect 43054 694199 43100 694211
rect 43212 694211 43218 694240
rect 43252 694211 43258 694240
rect 43212 694199 43258 694211
rect 43370 694211 43376 694850
rect 43410 694211 43416 694850
rect 43528 694550 43534 695187
rect 43568 694550 43574 695187
rect 43686 695187 43732 695199
rect 43686 695160 43692 695187
rect 43726 695160 43732 695187
rect 43844 695187 43890 695199
rect 43660 695090 43670 695160
rect 43740 695090 43750 695160
rect 43686 694920 43692 695090
rect 43726 694920 43732 695090
rect 43660 694850 43670 694920
rect 43740 694850 43750 694920
rect 43500 694480 43510 694550
rect 43580 694480 43590 694550
rect 43528 694310 43534 694480
rect 43568 694310 43574 694480
rect 43500 694240 43510 694310
rect 43580 694240 43590 694310
rect 43370 694199 43416 694211
rect 43528 694211 43534 694240
rect 43568 694211 43574 694240
rect 43528 694199 43574 694211
rect 43686 694211 43692 694850
rect 43726 694211 43732 694850
rect 43844 694550 43850 695187
rect 43884 694550 43890 695187
rect 44002 695187 44048 695199
rect 44002 695160 44008 695187
rect 44042 695160 44048 695187
rect 44160 695187 44206 695199
rect 43980 695090 43990 695160
rect 44060 695090 44070 695160
rect 44002 694920 44008 695090
rect 44042 694920 44048 695090
rect 43980 694850 43990 694920
rect 44060 694850 44070 694920
rect 43820 694480 43830 694550
rect 43900 694480 43910 694550
rect 43844 694310 43850 694480
rect 43884 694310 43890 694480
rect 43820 694240 43830 694310
rect 43900 694240 43910 694310
rect 43686 694199 43732 694211
rect 43844 694211 43850 694240
rect 43884 694211 43890 694240
rect 43844 694199 43890 694211
rect 44002 694211 44008 694850
rect 44042 694211 44048 694850
rect 44160 694550 44166 695187
rect 44200 694550 44206 695187
rect 44318 695187 44364 695199
rect 44318 695160 44324 695187
rect 44358 695160 44364 695187
rect 44476 695187 44522 695199
rect 44300 695090 44310 695160
rect 44380 695090 44390 695160
rect 44318 694920 44324 695090
rect 44358 694920 44364 695090
rect 44300 694850 44310 694920
rect 44380 694850 44390 694920
rect 44140 694480 44150 694550
rect 44220 694480 44230 694550
rect 44160 694310 44166 694480
rect 44200 694310 44206 694480
rect 44140 694240 44150 694310
rect 44220 694240 44230 694310
rect 44002 694199 44048 694211
rect 44160 694211 44166 694240
rect 44200 694211 44206 694240
rect 44160 694199 44206 694211
rect 44318 694211 44324 694850
rect 44358 694211 44364 694850
rect 44476 694550 44482 695187
rect 44516 694550 44522 695187
rect 44634 695187 44680 695199
rect 44634 695160 44640 695187
rect 44674 695160 44680 695187
rect 44792 695187 44838 695199
rect 44610 695090 44620 695160
rect 44690 695090 44700 695160
rect 44634 694920 44640 695090
rect 44674 694920 44680 695090
rect 44610 694850 44620 694920
rect 44690 694850 44700 694920
rect 44450 694480 44460 694550
rect 44530 694480 44540 694550
rect 44476 694310 44482 694480
rect 44516 694310 44522 694480
rect 44450 694240 44460 694310
rect 44530 694240 44540 694310
rect 44318 694199 44364 694211
rect 44476 694211 44482 694240
rect 44516 694211 44522 694240
rect 44476 694199 44522 694211
rect 44634 694211 44640 694850
rect 44674 694211 44680 694850
rect 44792 694550 44798 695187
rect 44832 694550 44838 695187
rect 44950 695187 44996 695199
rect 44950 695160 44956 695187
rect 44990 695160 44996 695187
rect 45108 695187 45154 695199
rect 44930 695090 44940 695160
rect 45010 695090 45020 695160
rect 44950 694920 44956 695090
rect 44990 694920 44996 695090
rect 44930 694850 44940 694920
rect 45010 694850 45020 694920
rect 44770 694480 44780 694550
rect 44850 694480 44860 694550
rect 44792 694310 44798 694480
rect 44832 694310 44838 694480
rect 44770 694240 44780 694310
rect 44850 694240 44860 694310
rect 44634 694199 44680 694211
rect 44792 694211 44798 694240
rect 44832 694211 44838 694240
rect 44792 694199 44838 694211
rect 44950 694211 44956 694850
rect 44990 694211 44996 694850
rect 45108 694550 45114 695187
rect 45148 694550 45154 695187
rect 45266 695187 45312 695199
rect 45266 695160 45272 695187
rect 45306 695160 45312 695187
rect 45424 695187 45470 695199
rect 45240 695090 45250 695160
rect 45320 695090 45330 695160
rect 45266 694920 45272 695090
rect 45306 694920 45312 695090
rect 45240 694850 45250 694920
rect 45320 694850 45330 694920
rect 45090 694480 45100 694550
rect 45170 694480 45180 694550
rect 45108 694310 45114 694480
rect 45148 694310 45154 694480
rect 45090 694240 45100 694310
rect 45170 694240 45180 694310
rect 44950 694199 44996 694211
rect 45108 694211 45114 694240
rect 45148 694211 45154 694240
rect 45108 694199 45154 694211
rect 45266 694211 45272 694850
rect 45306 694211 45312 694850
rect 45424 694550 45430 695187
rect 45464 694550 45470 695187
rect 45582 695187 45628 695199
rect 45582 695160 45588 695187
rect 45622 695160 45628 695187
rect 45740 695187 45786 695199
rect 45560 695090 45570 695160
rect 45640 695090 45650 695160
rect 45582 694920 45588 695090
rect 45622 694920 45628 695090
rect 45560 694850 45570 694920
rect 45640 694850 45650 694920
rect 45400 694480 45410 694550
rect 45480 694480 45490 694550
rect 45424 694310 45430 694480
rect 45464 694310 45470 694480
rect 45400 694240 45410 694310
rect 45480 694240 45490 694310
rect 45266 694199 45312 694211
rect 45424 694211 45430 694240
rect 45464 694211 45470 694240
rect 45424 694199 45470 694211
rect 45582 694211 45588 694850
rect 45622 694211 45628 694850
rect 45740 694550 45746 695187
rect 45780 694550 45786 695187
rect 45898 695187 45944 695199
rect 45898 695160 45904 695187
rect 45938 695160 45944 695187
rect 46056 695187 46102 695199
rect 45880 695090 45890 695160
rect 45960 695090 45970 695160
rect 45898 694920 45904 695090
rect 45938 694920 45944 695090
rect 45880 694850 45890 694920
rect 45960 694850 45970 694920
rect 45720 694480 45730 694550
rect 45800 694480 45810 694550
rect 45740 694310 45746 694480
rect 45780 694310 45786 694480
rect 45720 694240 45730 694310
rect 45800 694240 45810 694310
rect 45582 694199 45628 694211
rect 45740 694211 45746 694240
rect 45780 694211 45786 694240
rect 45740 694199 45786 694211
rect 45898 694211 45904 694850
rect 45938 694211 45944 694850
rect 46056 694550 46062 695187
rect 46096 694550 46102 695187
rect 46214 695187 46260 695199
rect 46214 695160 46220 695187
rect 46254 695160 46260 695187
rect 46372 695187 46418 695199
rect 46190 695090 46200 695160
rect 46270 695090 46280 695160
rect 46214 694920 46220 695090
rect 46254 694920 46260 695090
rect 46190 694850 46200 694920
rect 46270 694850 46280 694920
rect 46030 694480 46040 694550
rect 46110 694480 46120 694550
rect 46056 694310 46062 694480
rect 46096 694310 46102 694480
rect 46030 694240 46040 694310
rect 46110 694240 46120 694310
rect 45898 694199 45944 694211
rect 46056 694211 46062 694240
rect 46096 694211 46102 694240
rect 46056 694199 46102 694211
rect 46214 694211 46220 694850
rect 46254 694211 46260 694850
rect 46372 694550 46378 695187
rect 46412 694550 46418 695187
rect 46530 695187 46576 695199
rect 46530 695160 46536 695187
rect 46570 695160 46576 695187
rect 46688 695187 46734 695199
rect 46510 695090 46520 695160
rect 46590 695090 46600 695160
rect 46530 694920 46536 695090
rect 46570 694920 46576 695090
rect 46510 694850 46520 694920
rect 46590 694850 46600 694920
rect 46350 694480 46360 694550
rect 46430 694480 46440 694550
rect 46372 694310 46378 694480
rect 46412 694310 46418 694480
rect 46350 694240 46360 694310
rect 46430 694240 46440 694310
rect 46214 694199 46260 694211
rect 46372 694211 46378 694240
rect 46412 694211 46418 694240
rect 46372 694199 46418 694211
rect 46530 694211 46536 694850
rect 46570 694211 46576 694850
rect 46688 694550 46694 695187
rect 46728 694550 46734 695187
rect 46846 695187 46892 695199
rect 46846 695160 46852 695187
rect 46886 695160 46892 695187
rect 47004 695187 47050 695199
rect 46820 695090 46830 695160
rect 46900 695090 46910 695160
rect 46846 694920 46852 695090
rect 46886 694920 46892 695090
rect 46820 694850 46830 694920
rect 46900 694850 46910 694920
rect 46670 694480 46680 694550
rect 46750 694480 46760 694550
rect 46688 694310 46694 694480
rect 46728 694310 46734 694480
rect 46670 694240 46680 694310
rect 46750 694240 46760 694310
rect 46530 694199 46576 694211
rect 46688 694211 46694 694240
rect 46728 694211 46734 694240
rect 46688 694199 46734 694211
rect 46846 694211 46852 694850
rect 46886 694211 46892 694850
rect 47004 694550 47010 695187
rect 47044 694550 47050 695187
rect 47162 695187 47208 695199
rect 47162 695160 47168 695187
rect 47202 695160 47208 695187
rect 47320 695187 47366 695199
rect 47140 695090 47150 695160
rect 47220 695090 47230 695160
rect 47162 694920 47168 695090
rect 47202 694920 47208 695090
rect 47140 694850 47150 694920
rect 47220 694850 47230 694920
rect 46980 694480 46990 694550
rect 47060 694480 47070 694550
rect 47004 694310 47010 694480
rect 47044 694310 47050 694480
rect 46980 694240 46990 694310
rect 47060 694240 47070 694310
rect 46846 694199 46892 694211
rect 47004 694211 47010 694240
rect 47044 694211 47050 694240
rect 47004 694199 47050 694211
rect 47162 694211 47168 694850
rect 47202 694211 47208 694850
rect 47320 694550 47326 695187
rect 47360 694550 47366 695187
rect 47478 695187 47524 695199
rect 47478 695160 47484 695187
rect 47518 695160 47524 695187
rect 47636 695187 47682 695199
rect 47460 695090 47470 695160
rect 47540 695090 47550 695160
rect 47478 694920 47484 695090
rect 47518 694920 47524 695090
rect 47460 694850 47470 694920
rect 47540 694850 47550 694920
rect 47300 694480 47310 694550
rect 47380 694480 47390 694550
rect 47320 694310 47326 694480
rect 47360 694310 47366 694480
rect 47300 694240 47310 694310
rect 47380 694240 47390 694310
rect 47162 694199 47208 694211
rect 47320 694211 47326 694240
rect 47360 694211 47366 694240
rect 47320 694199 47366 694211
rect 47478 694211 47484 694850
rect 47518 694211 47524 694850
rect 47636 694550 47642 695187
rect 47676 694550 47682 695187
rect 47794 695187 47840 695199
rect 47794 695160 47800 695187
rect 47834 695160 47840 695187
rect 47770 695090 47780 695160
rect 47850 695090 47860 695160
rect 47794 694920 47800 695090
rect 47834 694920 47840 695090
rect 47770 694850 47780 694920
rect 47850 694850 47860 694920
rect 47910 694860 47990 695240
rect 48760 694999 48781 696113
rect 49178 694999 49190 696113
rect 48760 694860 49190 694999
rect 47620 694480 47630 694550
rect 47700 694480 47710 694550
rect 47636 694310 47642 694480
rect 47676 694310 47682 694480
rect 47620 694240 47630 694310
rect 47700 694240 47710 694310
rect 47478 694199 47524 694211
rect 47636 694211 47642 694240
rect 47676 694211 47682 694240
rect 47636 694199 47682 694211
rect 47794 694211 47800 694850
rect 47834 694211 47840 694850
rect 47794 694199 47840 694211
rect 47910 694653 49190 694860
rect 47910 694570 48781 694653
rect 47910 694160 47990 694570
rect 41330 694152 47990 694160
rect 41330 694118 41542 694152
rect 41610 694118 41700 694152
rect 41768 694118 41858 694152
rect 41926 694118 42016 694152
rect 42084 694118 42174 694152
rect 42242 694118 42332 694152
rect 42400 694118 42490 694152
rect 42558 694140 42648 694152
rect 42558 694118 42580 694140
rect 42716 694118 42806 694152
rect 42874 694118 42964 694152
rect 43032 694118 43122 694152
rect 43190 694118 43280 694152
rect 43348 694118 43438 694152
rect 43506 694118 43596 694152
rect 43664 694118 43754 694152
rect 43822 694118 43912 694152
rect 43980 694118 44070 694152
rect 44138 694118 44228 694152
rect 44296 694118 44386 694152
rect 44454 694118 44544 694152
rect 44612 694118 44702 694152
rect 44770 694118 44860 694152
rect 44928 694118 45018 694152
rect 45086 694118 45176 694152
rect 45244 694118 45334 694152
rect 45402 694118 45492 694152
rect 45560 694118 45650 694152
rect 45718 694118 45808 694152
rect 45876 694118 45966 694152
rect 46034 694118 46124 694152
rect 46192 694118 46282 694152
rect 46350 694118 46440 694152
rect 46508 694118 46598 694152
rect 46666 694140 46756 694152
rect 46720 694118 46756 694140
rect 46824 694118 46914 694152
rect 46982 694118 47072 694152
rect 47140 694118 47230 694152
rect 47298 694118 47388 694152
rect 47456 694118 47546 694152
rect 47614 694118 47704 694152
rect 47772 694118 47990 694152
rect 41330 694110 42580 694118
rect 42540 694060 42580 694110
rect 42660 694110 46640 694118
rect 42660 694060 42700 694110
rect 46600 694060 46640 694110
rect 46720 694110 47990 694118
rect 46720 694060 46760 694110
rect 42540 694050 42700 694060
rect 43760 694056 45550 694060
rect 43017 694050 46297 694056
rect 46600 694050 46760 694060
rect 43017 694016 43029 694050
rect 46285 694016 46297 694050
rect 43017 694010 46297 694016
rect 43760 694000 45550 694010
rect 43760 693730 44010 694000
rect 44280 693730 45060 694000
rect 45330 693730 45550 694000
rect 43760 693712 45550 693730
rect 43760 693678 43778 693712
rect 45534 693678 45550 693712
rect 43760 693670 45550 693678
rect 40120 693520 40560 693539
rect 42830 693610 46480 693620
rect 42830 693576 43042 693610
rect 43110 693576 43200 693610
rect 43268 693576 43358 693610
rect 43426 693576 43516 693610
rect 43584 693576 43674 693610
rect 43742 693576 43832 693610
rect 43900 693576 43990 693610
rect 44058 693576 44148 693610
rect 44216 693576 44306 693610
rect 44374 693576 44464 693610
rect 44532 693576 44622 693610
rect 44690 693576 44780 693610
rect 44848 693576 44938 693610
rect 45006 693576 45096 693610
rect 45164 693576 45254 693610
rect 45322 693576 45412 693610
rect 45480 693576 45570 693610
rect 45638 693576 45728 693610
rect 45796 693576 45886 693610
rect 45954 693576 46044 693610
rect 46112 693576 46202 693610
rect 46270 693576 46480 693610
rect 42830 693570 46480 693576
rect 38688 693460 38892 693466
rect 38688 693360 38700 693460
rect 38880 693360 38892 693460
rect 38688 693354 38892 693360
rect 39108 693460 39312 693466
rect 39108 693360 39120 693460
rect 39300 693360 39312 693460
rect 39108 693354 39312 693360
rect 42830 692490 42910 693570
rect 42974 693517 43020 693529
rect 42974 693490 42980 693517
rect 43014 693490 43020 693517
rect 43132 693517 43178 693529
rect 42950 693420 42960 693490
rect 43030 693420 43040 693490
rect 42974 693280 42980 693420
rect 43014 693280 43020 693420
rect 42950 693210 42960 693280
rect 43030 693210 43040 693280
rect 42974 692541 42980 693210
rect 43014 692541 43020 693210
rect 43132 692850 43138 693517
rect 43172 692850 43178 693517
rect 43290 693517 43336 693529
rect 43290 693490 43296 693517
rect 43330 693490 43336 693517
rect 43448 693517 43494 693529
rect 43270 693420 43280 693490
rect 43350 693420 43360 693490
rect 43290 693280 43296 693420
rect 43330 693280 43336 693420
rect 43270 693210 43280 693280
rect 43350 693210 43360 693280
rect 43110 692780 43120 692850
rect 43190 692780 43200 692850
rect 43132 692640 43138 692780
rect 43172 692640 43178 692780
rect 43110 692570 43120 692640
rect 43190 692570 43200 692640
rect 42974 692529 43020 692541
rect 43132 692541 43138 692570
rect 43172 692541 43178 692570
rect 43132 692529 43178 692541
rect 43290 692541 43296 693210
rect 43330 692541 43336 693210
rect 43448 692850 43454 693517
rect 43488 692850 43494 693517
rect 43606 693517 43652 693529
rect 43606 693490 43612 693517
rect 43646 693490 43652 693517
rect 43764 693517 43810 693529
rect 43580 693420 43590 693490
rect 43660 693420 43670 693490
rect 43606 693280 43612 693420
rect 43646 693280 43652 693420
rect 43580 693210 43590 693280
rect 43660 693210 43670 693280
rect 43430 692780 43440 692850
rect 43510 692780 43520 692850
rect 43448 692640 43454 692780
rect 43488 692640 43494 692780
rect 43430 692570 43440 692640
rect 43510 692570 43520 692640
rect 43290 692529 43336 692541
rect 43448 692541 43454 692570
rect 43488 692541 43494 692570
rect 43448 692529 43494 692541
rect 43606 692541 43612 693210
rect 43646 692541 43652 693210
rect 43764 692850 43770 693517
rect 43804 692850 43810 693517
rect 43922 693517 43968 693529
rect 43922 693490 43928 693517
rect 43962 693490 43968 693517
rect 44080 693517 44126 693529
rect 43900 693420 43910 693490
rect 43980 693420 43990 693490
rect 43922 693280 43928 693420
rect 43962 693280 43968 693420
rect 43900 693210 43910 693280
rect 43980 693210 43990 693280
rect 43740 692780 43750 692850
rect 43820 692780 43830 692850
rect 43764 692640 43770 692780
rect 43804 692640 43810 692780
rect 43740 692570 43750 692640
rect 43820 692570 43830 692640
rect 43606 692529 43652 692541
rect 43764 692541 43770 692570
rect 43804 692541 43810 692570
rect 43764 692529 43810 692541
rect 43922 692541 43928 693210
rect 43962 692541 43968 693210
rect 44080 692850 44086 693517
rect 44120 692850 44126 693517
rect 44238 693517 44284 693529
rect 44238 693490 44244 693517
rect 44278 693490 44284 693517
rect 44396 693517 44442 693529
rect 44220 693420 44230 693490
rect 44300 693420 44310 693490
rect 44238 693280 44244 693420
rect 44278 693280 44284 693420
rect 44220 693210 44230 693280
rect 44300 693210 44310 693280
rect 44060 692780 44070 692850
rect 44140 692780 44150 692850
rect 44080 692640 44086 692780
rect 44120 692640 44126 692780
rect 44060 692570 44070 692640
rect 44140 692570 44150 692640
rect 43922 692529 43968 692541
rect 44080 692541 44086 692570
rect 44120 692541 44126 692570
rect 44080 692529 44126 692541
rect 44238 692541 44244 693210
rect 44278 692541 44284 693210
rect 44396 692850 44402 693517
rect 44436 692850 44442 693517
rect 44554 693517 44600 693529
rect 44554 693490 44560 693517
rect 44594 693490 44600 693517
rect 44712 693517 44758 693529
rect 44530 693420 44540 693490
rect 44610 693420 44620 693490
rect 44554 693280 44560 693420
rect 44594 693280 44600 693420
rect 44530 693210 44540 693280
rect 44610 693210 44620 693280
rect 44380 692780 44390 692850
rect 44460 692780 44470 692850
rect 44396 692640 44402 692780
rect 44436 692640 44442 692780
rect 44380 692570 44390 692640
rect 44460 692570 44470 692640
rect 44238 692529 44284 692541
rect 44396 692541 44402 692570
rect 44436 692541 44442 692570
rect 44396 692529 44442 692541
rect 44554 692541 44560 693210
rect 44594 692541 44600 693210
rect 44712 692850 44718 693517
rect 44752 692850 44758 693517
rect 44870 693517 44916 693529
rect 44870 693490 44876 693517
rect 44910 693490 44916 693517
rect 45028 693517 45074 693529
rect 44850 693420 44860 693490
rect 44930 693420 44940 693490
rect 44870 693280 44876 693420
rect 44910 693280 44916 693420
rect 44850 693210 44860 693280
rect 44930 693210 44940 693280
rect 44690 692780 44700 692850
rect 44770 692780 44780 692850
rect 44712 692640 44718 692780
rect 44752 692640 44758 692780
rect 44690 692570 44700 692640
rect 44770 692570 44780 692640
rect 44554 692529 44600 692541
rect 44712 692541 44718 692570
rect 44752 692541 44758 692570
rect 44712 692529 44758 692541
rect 44870 692541 44876 693210
rect 44910 692541 44916 693210
rect 45028 692850 45034 693517
rect 45068 692850 45074 693517
rect 45186 693517 45232 693529
rect 45186 693490 45192 693517
rect 45226 693490 45232 693517
rect 45344 693517 45390 693529
rect 45170 693420 45180 693490
rect 45250 693420 45260 693490
rect 45186 693280 45192 693420
rect 45226 693280 45232 693420
rect 45170 693210 45180 693280
rect 45250 693210 45260 693280
rect 45010 692780 45020 692850
rect 45090 692780 45100 692850
rect 45028 692640 45034 692780
rect 45068 692640 45074 692780
rect 45010 692570 45020 692640
rect 45090 692570 45100 692640
rect 44870 692529 44916 692541
rect 45028 692541 45034 692570
rect 45068 692541 45074 692570
rect 45028 692529 45074 692541
rect 45186 692541 45192 693210
rect 45226 692541 45232 693210
rect 45344 692850 45350 693517
rect 45384 692850 45390 693517
rect 45502 693517 45548 693529
rect 45502 693490 45508 693517
rect 45542 693490 45548 693517
rect 45660 693517 45706 693529
rect 45480 693420 45490 693490
rect 45560 693420 45570 693490
rect 45502 693280 45508 693420
rect 45542 693280 45548 693420
rect 45480 693210 45490 693280
rect 45560 693210 45570 693280
rect 45320 692780 45330 692850
rect 45400 692780 45410 692850
rect 45344 692640 45350 692780
rect 45384 692640 45390 692780
rect 45320 692570 45330 692640
rect 45400 692570 45410 692640
rect 45186 692529 45232 692541
rect 45344 692541 45350 692570
rect 45384 692541 45390 692570
rect 45344 692529 45390 692541
rect 45502 692541 45508 693210
rect 45542 692541 45548 693210
rect 45660 692850 45666 693517
rect 45700 692850 45706 693517
rect 45818 693517 45864 693529
rect 45818 693490 45824 693517
rect 45858 693490 45864 693517
rect 45976 693517 46022 693529
rect 45800 693420 45810 693490
rect 45880 693420 45890 693490
rect 45818 693280 45824 693420
rect 45858 693280 45864 693420
rect 45800 693210 45810 693280
rect 45880 693210 45890 693280
rect 45640 692780 45650 692850
rect 45720 692780 45730 692850
rect 45660 692640 45666 692780
rect 45700 692640 45706 692780
rect 45640 692570 45650 692640
rect 45720 692570 45730 692640
rect 45502 692529 45548 692541
rect 45660 692541 45666 692570
rect 45700 692541 45706 692570
rect 45660 692529 45706 692541
rect 45818 692541 45824 693210
rect 45858 692541 45864 693210
rect 45976 692850 45982 693517
rect 46016 692850 46022 693517
rect 46134 693517 46180 693529
rect 46134 693490 46140 693517
rect 46174 693490 46180 693517
rect 46292 693517 46338 693529
rect 46110 693420 46120 693490
rect 46190 693420 46200 693490
rect 46134 693280 46140 693420
rect 46174 693280 46180 693420
rect 46110 693210 46120 693280
rect 46190 693210 46200 693280
rect 45960 692780 45970 692850
rect 46040 692780 46050 692850
rect 45976 692640 45982 692780
rect 46016 692640 46022 692780
rect 45960 692570 45970 692640
rect 46040 692570 46050 692640
rect 45818 692529 45864 692541
rect 45976 692541 45982 692570
rect 46016 692541 46022 692570
rect 45976 692529 46022 692541
rect 46134 692541 46140 693210
rect 46174 692541 46180 693210
rect 46292 692850 46298 693517
rect 46332 692850 46338 693517
rect 46270 692780 46280 692850
rect 46350 692780 46360 692850
rect 46292 692640 46298 692780
rect 46332 692640 46338 692780
rect 46270 692570 46280 692640
rect 46350 692570 46360 692640
rect 46134 692529 46180 692541
rect 46292 692541 46298 692570
rect 46332 692541 46338 692570
rect 46292 692529 46338 692541
rect 46400 692490 46480 693570
rect 48760 693539 48781 694570
rect 49178 693539 49190 694653
rect 48760 693520 49190 693539
rect 51190 696113 51630 696130
rect 51190 694999 51212 696113
rect 51609 694999 51630 696113
rect 51190 694940 51630 694999
rect 51190 694920 52520 694940
rect 51190 694850 52320 694920
rect 52390 694850 52520 694920
rect 51190 694810 52520 694850
rect 51190 694740 52430 694810
rect 52500 694740 52520 694810
rect 51190 694720 52520 694740
rect 51190 694653 51630 694720
rect 51190 693539 51212 694653
rect 51609 693539 51630 694653
rect 51190 693520 51630 693539
rect 49938 693460 50142 693466
rect 49938 693360 49950 693460
rect 50130 693360 50142 693460
rect 49938 693354 50142 693360
rect 50358 693460 50562 693466
rect 50358 693360 50370 693460
rect 50550 693360 50562 693460
rect 50358 693354 50562 693360
rect 42830 692482 46480 692490
rect 42830 692448 43042 692482
rect 43110 692448 43200 692482
rect 43268 692448 43358 692482
rect 43426 692448 43516 692482
rect 43584 692448 43674 692482
rect 43742 692448 43832 692482
rect 43900 692448 43990 692482
rect 44058 692448 44148 692482
rect 44216 692448 44306 692482
rect 44374 692448 44464 692482
rect 44532 692448 44622 692482
rect 44690 692448 44780 692482
rect 44848 692448 44938 692482
rect 45006 692448 45096 692482
rect 45164 692448 45254 692482
rect 45322 692448 45412 692482
rect 45480 692448 45570 692482
rect 45638 692448 45728 692482
rect 45796 692448 45886 692482
rect 45954 692448 46044 692482
rect 46112 692448 46202 692482
rect 46270 692448 46480 692482
rect 42830 692440 46480 692448
rect 43020 692080 43290 692440
rect 43770 692386 43780 692390
rect 43628 692380 43780 692386
rect 44040 692386 44050 692390
rect 44040 692380 44222 692386
rect 43628 692140 43640 692380
rect 44210 692140 44222 692380
rect 43628 692134 43780 692140
rect 43770 692130 43780 692134
rect 44040 692134 44222 692140
rect 44040 692130 44050 692134
rect 44520 692080 44790 692440
rect 45270 692386 45280 692390
rect 45098 692380 45280 692386
rect 45540 692386 45550 692390
rect 45540 692380 45692 692386
rect 45098 692140 45110 692380
rect 45680 692140 45692 692380
rect 45098 692134 45280 692140
rect 45270 692130 45280 692134
rect 45540 692134 45692 692140
rect 45540 692130 45550 692134
rect 46020 692080 46290 692440
rect 43020 692070 46290 692080
rect 43020 692036 43042 692070
rect 43110 692036 43200 692070
rect 43268 692036 43358 692070
rect 43426 692036 43516 692070
rect 43584 692036 43674 692070
rect 43742 692036 43832 692070
rect 43900 692036 43990 692070
rect 44058 692036 44148 692070
rect 44216 692036 44306 692070
rect 44374 692036 44464 692070
rect 44532 692036 44622 692070
rect 44690 692036 44780 692070
rect 44848 692036 44938 692070
rect 45006 692036 45096 692070
rect 45164 692036 45254 692070
rect 45322 692036 45412 692070
rect 45480 692036 45570 692070
rect 45638 692036 45728 692070
rect 45796 692036 45886 692070
rect 45954 692036 46044 692070
rect 46112 692036 46202 692070
rect 46270 692036 46290 692070
rect 43020 692030 46290 692036
rect 42974 691977 43020 691989
rect 42974 691940 42980 691977
rect 43014 691940 43020 691977
rect 43132 691977 43178 691989
rect 42950 691870 42960 691940
rect 43030 691870 43040 691940
rect 42974 691730 42980 691870
rect 43014 691730 43020 691870
rect 42950 691660 42960 691730
rect 43030 691660 43040 691730
rect 42974 691001 42980 691660
rect 43014 691001 43020 691660
rect 43132 691310 43138 691977
rect 43172 691310 43178 691977
rect 43290 691977 43336 691989
rect 43290 691940 43296 691977
rect 43330 691940 43336 691977
rect 43440 691977 43500 692030
rect 43270 691870 43280 691940
rect 43350 691870 43360 691940
rect 43290 691730 43296 691870
rect 43330 691730 43336 691870
rect 43270 691660 43280 691730
rect 43350 691660 43360 691730
rect 43110 691240 43120 691310
rect 43190 691240 43200 691310
rect 43132 691100 43138 691240
rect 43172 691100 43178 691240
rect 43110 691030 43120 691100
rect 43190 691030 43200 691100
rect 42974 690989 43020 691001
rect 43132 691001 43138 691030
rect 43172 691001 43178 691030
rect 43132 690989 43178 691001
rect 43290 691001 43296 691660
rect 43330 691001 43336 691660
rect 43440 691310 43454 691977
rect 43488 691310 43500 691977
rect 43606 691977 43652 691989
rect 43606 691940 43612 691977
rect 43646 691940 43652 691977
rect 43760 691977 43820 692030
rect 43580 691870 43590 691940
rect 43660 691870 43670 691940
rect 43606 691730 43612 691870
rect 43646 691730 43652 691870
rect 43580 691660 43590 691730
rect 43660 691660 43670 691730
rect 43430 691240 43440 691310
rect 43510 691240 43520 691310
rect 43440 691100 43454 691240
rect 43488 691100 43500 691240
rect 43430 691030 43440 691100
rect 43510 691030 43520 691100
rect 43290 690989 43336 691001
rect 43440 691001 43454 691030
rect 43488 691001 43500 691030
rect 43440 690950 43500 691001
rect 43606 691001 43612 691660
rect 43646 691001 43652 691660
rect 43760 691310 43770 691977
rect 43804 691310 43820 691977
rect 43922 691977 43968 691989
rect 43922 691940 43928 691977
rect 43962 691940 43968 691977
rect 44080 691977 44126 691989
rect 43900 691870 43910 691940
rect 43980 691870 43990 691940
rect 43922 691730 43928 691870
rect 43962 691730 43968 691870
rect 43900 691660 43910 691730
rect 43980 691660 43990 691730
rect 43740 691240 43750 691310
rect 43820 691240 43830 691310
rect 43760 691100 43770 691240
rect 43804 691100 43820 691240
rect 43740 691030 43750 691100
rect 43820 691030 43830 691100
rect 43606 690989 43652 691001
rect 43760 691001 43770 691030
rect 43804 691001 43820 691030
rect 43760 690950 43820 691001
rect 43922 691001 43928 691660
rect 43962 691001 43968 691660
rect 44080 691310 44086 691977
rect 44120 691310 44126 691977
rect 44238 691977 44284 691989
rect 44238 691940 44244 691977
rect 44278 691940 44284 691977
rect 44396 691977 44442 691989
rect 44220 691870 44230 691940
rect 44300 691870 44310 691940
rect 44238 691730 44244 691870
rect 44278 691730 44284 691870
rect 44220 691660 44230 691730
rect 44300 691660 44310 691730
rect 44060 691240 44070 691310
rect 44140 691240 44150 691310
rect 44080 691100 44086 691240
rect 44120 691100 44126 691240
rect 44060 691030 44070 691100
rect 44140 691030 44150 691100
rect 43922 690989 43968 691001
rect 44080 691001 44086 691030
rect 44120 691001 44126 691030
rect 44080 690989 44126 691001
rect 44238 691001 44244 691660
rect 44278 691001 44284 691660
rect 44396 691310 44402 691977
rect 44436 691310 44442 691977
rect 44554 691977 44600 691989
rect 44554 691940 44560 691977
rect 44594 691940 44600 691977
rect 44712 691977 44758 691989
rect 44530 691870 44540 691940
rect 44610 691870 44620 691940
rect 44554 691730 44560 691870
rect 44594 691730 44600 691870
rect 44530 691660 44540 691730
rect 44610 691660 44620 691730
rect 44370 691240 44380 691310
rect 44450 691240 44460 691310
rect 44396 691100 44402 691240
rect 44436 691100 44442 691240
rect 44370 691030 44380 691100
rect 44450 691030 44460 691100
rect 44238 690989 44284 691001
rect 44396 691001 44402 691030
rect 44436 691001 44442 691030
rect 44396 690989 44442 691001
rect 44554 691001 44560 691660
rect 44594 691001 44600 691660
rect 44712 691310 44718 691977
rect 44752 691310 44758 691977
rect 44870 691977 44916 691989
rect 44870 691940 44876 691977
rect 44910 691940 44916 691977
rect 45028 691977 45074 691989
rect 44850 691870 44860 691940
rect 44930 691870 44940 691940
rect 44870 691730 44876 691870
rect 44910 691730 44916 691870
rect 44850 691660 44860 691730
rect 44930 691660 44940 691730
rect 44690 691240 44700 691310
rect 44770 691240 44780 691310
rect 44712 691100 44718 691240
rect 44752 691100 44758 691240
rect 44690 691030 44700 691100
rect 44770 691030 44780 691100
rect 44554 690989 44600 691001
rect 44712 691001 44718 691030
rect 44752 691001 44758 691030
rect 44712 690989 44758 691001
rect 44870 691001 44876 691660
rect 44910 691001 44916 691660
rect 45028 691310 45034 691977
rect 45068 691310 45074 691977
rect 45186 691977 45232 691989
rect 45186 691940 45192 691977
rect 45226 691940 45232 691977
rect 45344 691977 45390 691989
rect 45160 691870 45170 691940
rect 45240 691870 45250 691940
rect 45186 691730 45192 691870
rect 45226 691730 45232 691870
rect 45160 691660 45170 691730
rect 45240 691660 45250 691730
rect 45010 691240 45020 691310
rect 45090 691240 45100 691310
rect 45028 691100 45034 691240
rect 45068 691100 45074 691240
rect 45010 691030 45020 691100
rect 45090 691030 45100 691100
rect 44870 690989 44916 691001
rect 45028 691001 45034 691030
rect 45068 691001 45074 691030
rect 45028 690989 45074 691001
rect 45186 691001 45192 691660
rect 45226 691001 45232 691660
rect 45344 691310 45350 691977
rect 45384 691310 45390 691977
rect 45502 691977 45548 691989
rect 45502 691940 45508 691977
rect 45542 691940 45548 691977
rect 45650 691977 45710 692030
rect 45480 691870 45490 691940
rect 45560 691870 45570 691940
rect 45502 691730 45508 691870
rect 45542 691730 45548 691870
rect 45480 691660 45490 691730
rect 45560 691660 45570 691730
rect 45320 691240 45330 691310
rect 45400 691240 45410 691310
rect 45344 691100 45350 691240
rect 45384 691100 45390 691240
rect 45320 691030 45330 691100
rect 45400 691030 45410 691100
rect 45186 690989 45232 691001
rect 45344 691001 45350 691030
rect 45384 691001 45390 691030
rect 45344 690989 45390 691001
rect 45502 691001 45508 691660
rect 45542 691001 45548 691660
rect 45650 691310 45666 691977
rect 45700 691310 45710 691977
rect 45818 691977 45864 691989
rect 45818 691940 45824 691977
rect 45858 691940 45864 691977
rect 45970 691977 46030 692030
rect 45800 691870 45810 691940
rect 45880 691870 45890 691940
rect 45818 691730 45824 691870
rect 45858 691730 45864 691870
rect 45800 691660 45810 691730
rect 45880 691660 45890 691730
rect 45640 691240 45650 691310
rect 45720 691240 45730 691310
rect 45650 691100 45666 691240
rect 45700 691100 45710 691240
rect 45640 691030 45650 691100
rect 45720 691030 45730 691100
rect 45502 690989 45548 691001
rect 45650 691001 45666 691030
rect 45700 691001 45710 691030
rect 45650 690950 45710 691001
rect 45818 691001 45824 691660
rect 45858 691001 45864 691660
rect 45970 691310 45982 691977
rect 46016 691310 46030 691977
rect 46134 691977 46180 691989
rect 46134 691940 46140 691977
rect 46174 691940 46180 691977
rect 46292 691977 46338 691989
rect 46110 691870 46120 691940
rect 46190 691870 46200 691940
rect 46134 691730 46140 691870
rect 46174 691730 46180 691870
rect 46110 691660 46120 691730
rect 46190 691660 46200 691730
rect 45950 691240 45960 691310
rect 46030 691240 46040 691310
rect 45970 691100 45982 691240
rect 46016 691100 46030 691240
rect 45950 691030 45960 691100
rect 46030 691030 46040 691100
rect 45818 690989 45864 691001
rect 45970 691001 45982 691030
rect 46016 691001 46030 691030
rect 45970 690950 46030 691001
rect 46134 691001 46140 691660
rect 46174 691001 46180 691660
rect 46292 691310 46298 691977
rect 46332 691310 46338 691977
rect 46270 691240 46280 691310
rect 46350 691240 46360 691310
rect 46292 691100 46298 691240
rect 46332 691100 46338 691240
rect 566260 691100 571840 691320
rect 46270 691030 46280 691100
rect 46350 691030 46360 691100
rect 46134 690989 46180 691001
rect 46292 691001 46298 691030
rect 46332 691001 46338 691030
rect 46292 690989 46338 691001
rect 546907 690972 547011 690978
rect 541957 690962 542071 690968
rect 43020 690942 46290 690950
rect 43020 690908 43042 690942
rect 43110 690908 43200 690942
rect 43268 690908 43358 690942
rect 43426 690908 43516 690942
rect 43584 690908 43674 690942
rect 43742 690908 43832 690942
rect 43900 690908 43990 690942
rect 44058 690908 44148 690942
rect 44216 690908 44306 690942
rect 44374 690908 44464 690942
rect 44532 690908 44622 690942
rect 44690 690908 44780 690942
rect 44848 690908 44938 690942
rect 45006 690908 45096 690942
rect 45164 690908 45254 690942
rect 45322 690908 45412 690942
rect 45480 690908 45570 690942
rect 45638 690908 45728 690942
rect 45796 690908 45886 690942
rect 45954 690908 46044 690942
rect 46112 690908 46202 690942
rect 46270 690908 46290 690942
rect 43020 690900 46290 690908
rect 541957 690892 541969 690962
rect 542059 690892 542071 690962
rect 541957 690886 542071 690892
rect 542127 690962 542241 690968
rect 542127 690892 542139 690962
rect 542229 690892 542241 690962
rect 542127 690886 542241 690892
rect 544447 690962 544561 690968
rect 544447 690892 544459 690962
rect 544549 690892 544561 690962
rect 544447 690886 544561 690892
rect 544617 690962 544731 690968
rect 544617 690892 544629 690962
rect 544719 690892 544731 690962
rect 544617 690886 544731 690892
rect 546907 690892 546919 690972
rect 546999 690892 547011 690972
rect 546907 690886 547011 690892
rect 547077 690972 547181 690978
rect 547077 690892 547089 690972
rect 547169 690892 547181 690972
rect 547077 690886 547181 690892
rect 566260 690900 566300 691100
rect 566500 690900 566700 691100
rect 566900 690900 567100 691100
rect 567300 690900 567500 691100
rect 567700 690900 567900 691100
rect 568100 690900 568300 691100
rect 568500 690900 568700 691100
rect 568900 690900 569100 691100
rect 569300 690900 569500 691100
rect 569700 690900 569900 691100
rect 570100 690900 570300 691100
rect 570500 690900 570700 691100
rect 570900 690900 571100 691100
rect 571300 690900 571500 691100
rect 571700 690900 571840 691100
rect 541959 690802 541969 690852
rect 540359 690784 541969 690802
rect 542049 690802 542059 690852
rect 542129 690802 542139 690852
rect 542049 690784 542139 690802
rect 542219 690802 542229 690852
rect 544449 690802 544459 690852
rect 542219 690784 544459 690802
rect 544539 690802 544549 690852
rect 544619 690802 544629 690852
rect 544539 690784 544629 690802
rect 544709 690802 544719 690852
rect 546909 690802 546919 690842
rect 544709 690784 546919 690802
rect 546999 690802 547009 690842
rect 547079 690802 547089 690842
rect 546999 690784 547089 690802
rect 547169 690802 547179 690842
rect 547169 690784 548799 690802
rect 540359 690762 540380 690784
rect 540368 690750 540380 690762
rect 541356 690762 541616 690784
rect 541356 690750 541368 690762
rect 540368 690744 541368 690750
rect 541604 690750 541616 690762
rect 542592 690762 542852 690784
rect 542592 690750 542604 690762
rect 541604 690744 542604 690750
rect 542840 690750 542852 690762
rect 543828 690762 544088 690784
rect 543828 690750 543840 690762
rect 542840 690744 543840 690750
rect 544076 690750 544088 690762
rect 545064 690762 545324 690784
rect 545064 690750 545076 690762
rect 544076 690744 545076 690750
rect 545312 690750 545324 690762
rect 546300 690762 546560 690784
rect 547536 690762 547796 690784
rect 546300 690750 546312 690762
rect 545312 690744 546312 690750
rect 546548 690750 546560 690762
rect 547536 690750 547548 690762
rect 546548 690744 547548 690750
rect 547784 690750 547796 690762
rect 548772 690762 548799 690784
rect 548772 690750 548784 690762
rect 547784 690744 548784 690750
rect 540281 690722 540327 690734
rect 540281 690672 540287 690722
rect 540269 690654 540287 690672
rect 540321 690712 540327 690722
rect 541409 690722 541455 690734
rect 541517 690722 541563 690734
rect 541409 690712 541415 690722
rect 540321 690682 541415 690712
rect 540321 690654 541089 690682
rect 540269 690626 541089 690654
rect 541169 690626 541239 690682
rect 541319 690654 541415 690682
rect 541557 690712 541563 690722
rect 542645 690722 542691 690734
rect 542753 690722 542799 690734
rect 543881 690722 543927 690734
rect 543989 690722 544035 690734
rect 542645 690712 542651 690722
rect 541557 690654 542651 690712
rect 542793 690712 542799 690722
rect 543879 690712 543887 690722
rect 542793 690682 543887 690712
rect 542793 690654 543579 690682
rect 541319 690652 541419 690654
rect 541549 690652 542659 690654
rect 542789 690652 543579 690654
rect 541319 690626 543579 690652
rect 543659 690626 543729 690682
rect 543809 690654 543887 690682
rect 544029 690712 544035 690722
rect 545117 690722 545163 690734
rect 545225 690722 545271 690734
rect 545117 690712 545123 690722
rect 544029 690654 545123 690712
rect 545265 690712 545271 690722
rect 546353 690722 546399 690734
rect 546461 690722 546507 690734
rect 547589 690722 547635 690734
rect 547697 690722 547743 690734
rect 546353 690712 546359 690722
rect 545265 690682 546359 690712
rect 545265 690654 546059 690682
rect 543809 690652 543889 690654
rect 544019 690652 545129 690654
rect 545259 690652 546059 690654
rect 543809 690626 546059 690652
rect 546139 690626 546209 690682
rect 546289 690654 546359 690682
rect 546501 690712 546509 690722
rect 547589 690712 547595 690722
rect 546501 690654 547595 690712
rect 547737 690712 547743 690722
rect 548825 690722 548871 690734
rect 548825 690712 548831 690722
rect 547737 690654 548831 690712
rect 548865 690672 548871 690722
rect 566260 690700 571840 690900
rect 548865 690654 548879 690672
rect 546289 690652 546369 690654
rect 546499 690652 547599 690654
rect 547729 690652 548879 690654
rect 546289 690626 548879 690652
rect 44314 690595 44988 690601
rect 44314 690561 44326 690595
rect 44976 690561 44988 690595
rect 540269 690592 540380 690626
rect 541356 690592 541616 690626
rect 542592 690592 542852 690626
rect 543828 690592 544088 690626
rect 545064 690592 545324 690626
rect 546300 690592 546560 690626
rect 547536 690592 547796 690626
rect 548772 690592 548879 690626
rect 540269 690572 540699 690592
rect 44314 690555 44988 690561
rect 540689 690532 540699 690572
rect 540779 690572 540869 690592
rect 540779 690532 540789 690572
rect 540859 690532 540869 690572
rect 540949 690572 543219 690592
rect 540949 690532 540959 690572
rect 543209 690532 543219 690572
rect 543299 690572 543389 690592
rect 543299 690532 543309 690572
rect 543379 690532 543389 690572
rect 543469 690572 545709 690592
rect 543469 690532 543479 690572
rect 545699 690532 545709 690572
rect 545789 690572 545879 690592
rect 545789 690532 545799 690572
rect 545869 690532 545879 690572
rect 545959 690572 548159 690592
rect 545959 690532 545969 690572
rect 548149 690532 548159 690572
rect 548239 690572 548329 690592
rect 548239 690532 548249 690572
rect 548319 690532 548329 690572
rect 548409 690572 548879 690592
rect 548409 690532 548419 690572
rect 566260 690500 566300 690700
rect 566500 690500 566700 690700
rect 566900 690500 567100 690700
rect 567300 690500 567500 690700
rect 567700 690500 567900 690700
rect 568100 690500 568300 690700
rect 568500 690500 568700 690700
rect 568900 690500 569100 690700
rect 569300 690500 569500 690700
rect 569700 690500 569900 690700
rect 570100 690500 570300 690700
rect 570500 690500 570700 690700
rect 570900 690500 571100 690700
rect 571300 690500 571500 690700
rect 571700 690500 571840 690700
rect 43870 690493 45430 690500
rect 43870 690459 44143 690493
rect 44211 690459 44301 690493
rect 44369 690459 44459 690493
rect 44527 690459 44617 690493
rect 44685 690459 44775 690493
rect 44843 690459 44933 690493
rect 45001 690459 45091 690493
rect 45159 690459 45430 690493
rect 43870 690450 45430 690459
rect 43870 689390 43950 690450
rect 44075 690409 44121 690421
rect 44075 690380 44081 690409
rect 44115 690380 44121 690409
rect 44233 690409 44279 690421
rect 44050 690310 44060 690380
rect 44130 690310 44140 690380
rect 44075 690090 44081 690310
rect 44115 690090 44121 690310
rect 44050 690020 44060 690090
rect 44130 690020 44140 690090
rect 44075 689433 44081 690020
rect 44115 689433 44121 690020
rect 44233 689820 44239 690409
rect 44273 689820 44279 690409
rect 44391 690409 44437 690421
rect 44391 690380 44397 690409
rect 44431 690380 44437 690409
rect 44549 690409 44595 690421
rect 44370 690310 44380 690380
rect 44450 690310 44460 690380
rect 44391 690090 44397 690310
rect 44431 690090 44437 690310
rect 44370 690020 44380 690090
rect 44450 690020 44460 690090
rect 44210 689750 44220 689820
rect 44290 689750 44300 689820
rect 44233 689530 44239 689750
rect 44273 689530 44279 689750
rect 44210 689460 44220 689530
rect 44290 689460 44300 689530
rect 44075 689421 44121 689433
rect 44233 689433 44239 689460
rect 44273 689433 44279 689460
rect 44233 689421 44279 689433
rect 44391 689433 44397 690020
rect 44431 689433 44437 690020
rect 44549 689820 44555 690409
rect 44589 689820 44595 690409
rect 44707 690409 44753 690421
rect 44707 690380 44713 690409
rect 44747 690380 44753 690409
rect 44865 690409 44911 690421
rect 44680 690310 44690 690380
rect 44760 690310 44770 690380
rect 44707 690090 44713 690310
rect 44747 690090 44753 690310
rect 44680 690020 44690 690090
rect 44760 690020 44770 690090
rect 44520 689750 44530 689820
rect 44600 689750 44610 689820
rect 44549 689530 44555 689750
rect 44589 689530 44595 689750
rect 44520 689460 44530 689530
rect 44600 689460 44610 689530
rect 44391 689421 44437 689433
rect 44549 689433 44555 689460
rect 44589 689433 44595 689460
rect 44549 689421 44595 689433
rect 44707 689433 44713 690020
rect 44747 689433 44753 690020
rect 44865 689820 44871 690409
rect 44905 689820 44911 690409
rect 45023 690409 45069 690421
rect 45023 690380 45029 690409
rect 45063 690380 45069 690409
rect 45181 690409 45227 690421
rect 45000 690310 45010 690380
rect 45080 690310 45090 690380
rect 45023 690090 45029 690310
rect 45063 690090 45069 690310
rect 45000 690020 45010 690090
rect 45080 690020 45090 690090
rect 44840 689750 44850 689820
rect 44920 689750 44930 689820
rect 44865 689530 44871 689750
rect 44905 689530 44911 689750
rect 44840 689460 44850 689530
rect 44920 689460 44930 689530
rect 44707 689421 44753 689433
rect 44865 689433 44871 689460
rect 44905 689433 44911 689460
rect 44865 689421 44911 689433
rect 45023 689433 45029 690020
rect 45063 689433 45069 690020
rect 45181 689820 45187 690409
rect 45221 689820 45227 690409
rect 45350 690010 45430 690450
rect 47100 690300 47400 690400
rect 47100 690200 47200 690300
rect 47300 690200 47400 690300
rect 541959 690262 541969 690312
rect 540359 690244 541969 690262
rect 542049 690262 542059 690312
rect 542129 690262 542139 690312
rect 542049 690244 542139 690262
rect 542219 690262 542229 690312
rect 544449 690262 544459 690312
rect 542219 690244 544459 690262
rect 544539 690262 544549 690312
rect 544619 690262 544629 690312
rect 544539 690244 544629 690262
rect 544709 690262 544719 690312
rect 546909 690262 546919 690302
rect 544709 690244 546919 690262
rect 546999 690262 547009 690302
rect 547079 690262 547089 690302
rect 546999 690244 547089 690262
rect 547169 690262 547179 690302
rect 566260 690300 571840 690500
rect 547169 690244 548799 690262
rect 540359 690222 540380 690244
rect 540368 690210 540380 690222
rect 541356 690222 541616 690244
rect 541356 690210 541368 690222
rect 540368 690204 541368 690210
rect 541604 690210 541616 690222
rect 542592 690222 542852 690244
rect 542592 690210 542604 690222
rect 541604 690204 542604 690210
rect 542840 690210 542852 690222
rect 543828 690222 544088 690244
rect 543828 690210 543840 690222
rect 542840 690204 543840 690210
rect 544076 690210 544088 690222
rect 545064 690222 545324 690244
rect 545064 690210 545076 690222
rect 544076 690204 545076 690210
rect 545312 690210 545324 690222
rect 546300 690222 546560 690244
rect 547536 690222 547796 690244
rect 546300 690210 546312 690222
rect 545312 690204 546312 690210
rect 546548 690210 546560 690222
rect 547536 690210 547548 690222
rect 546548 690204 547548 690210
rect 547784 690210 547796 690222
rect 548772 690222 548799 690244
rect 548772 690210 548784 690222
rect 547784 690204 548784 690210
rect 47100 690010 47400 690200
rect 540281 690182 540327 690194
rect 540281 690132 540287 690182
rect 540279 690114 540287 690132
rect 540321 690172 540327 690182
rect 541409 690182 541455 690194
rect 541517 690182 541563 690194
rect 541409 690172 541415 690182
rect 540321 690142 541415 690172
rect 540321 690114 541089 690142
rect 540279 690086 541089 690114
rect 541169 690086 541239 690142
rect 541319 690114 541415 690142
rect 541557 690172 541563 690182
rect 542645 690182 542691 690194
rect 542753 690182 542799 690194
rect 543881 690182 543927 690194
rect 543989 690182 544035 690194
rect 542645 690172 542651 690182
rect 541557 690114 542651 690172
rect 542793 690172 542799 690182
rect 543879 690172 543887 690182
rect 542793 690142 543887 690172
rect 542793 690114 543579 690142
rect 541319 690112 541419 690114
rect 541549 690112 542659 690114
rect 542789 690112 543579 690114
rect 541319 690086 543579 690112
rect 543659 690086 543729 690142
rect 543809 690114 543887 690142
rect 544029 690172 544035 690182
rect 545117 690182 545163 690194
rect 545225 690182 545271 690194
rect 545117 690172 545123 690182
rect 544029 690114 545123 690172
rect 545265 690172 545271 690182
rect 546353 690182 546399 690194
rect 546461 690182 546507 690194
rect 547589 690182 547635 690194
rect 547697 690182 547743 690194
rect 546353 690172 546359 690182
rect 545265 690142 546359 690172
rect 545265 690114 546059 690142
rect 543809 690112 543889 690114
rect 544019 690112 545129 690114
rect 545259 690112 546059 690114
rect 543809 690086 546059 690112
rect 546139 690086 546209 690142
rect 546289 690114 546359 690142
rect 546501 690172 546509 690182
rect 547589 690172 547595 690182
rect 546501 690114 547595 690172
rect 547737 690172 547743 690182
rect 548825 690182 548871 690194
rect 548825 690172 548831 690182
rect 547737 690114 548831 690172
rect 548865 690114 548871 690182
rect 546289 690112 546369 690114
rect 546499 690112 547599 690114
rect 547729 690112 548871 690114
rect 546289 690102 548871 690112
rect 546289 690086 548859 690102
rect 540279 690052 540380 690086
rect 541356 690052 541616 690086
rect 542592 690052 542852 690086
rect 543828 690052 544088 690086
rect 545064 690052 545324 690086
rect 546300 690052 546560 690086
rect 547536 690052 547796 690086
rect 548772 690052 548859 690086
rect 540279 690032 540699 690052
rect 45350 690000 47400 690010
rect 45350 689830 47200 690000
rect 45160 689750 45170 689820
rect 45240 689750 45250 689820
rect 45181 689530 45187 689750
rect 45221 689530 45227 689750
rect 45160 689460 45170 689530
rect 45240 689460 45250 689530
rect 45023 689421 45069 689433
rect 45181 689433 45187 689460
rect 45221 689433 45227 689460
rect 45181 689421 45227 689433
rect 45350 689390 45430 689830
rect 47100 689800 47200 689830
rect 47300 689800 47400 690000
rect 540689 689992 540699 690032
rect 540779 690032 540869 690052
rect 540779 689992 540789 690032
rect 540859 689992 540869 690032
rect 540949 690032 543219 690052
rect 540949 689992 540959 690032
rect 543209 689992 543219 690032
rect 543299 690032 543389 690052
rect 543299 689992 543309 690032
rect 543379 689992 543389 690032
rect 543469 690032 545709 690052
rect 543469 689992 543479 690032
rect 545699 689992 545709 690032
rect 545789 690032 545879 690052
rect 545789 689992 545799 690032
rect 545869 689992 545879 690032
rect 545959 690032 548159 690052
rect 545959 689992 545969 690032
rect 548149 689982 548159 690032
rect 548239 690032 548329 690052
rect 548239 689982 548249 690032
rect 548319 689982 548329 690032
rect 548409 690032 548859 690052
rect 566260 690100 566300 690300
rect 566500 690100 566700 690300
rect 566900 690100 567100 690300
rect 567300 690100 567500 690300
rect 567700 690100 567900 690300
rect 568100 690100 568300 690300
rect 568500 690100 568700 690300
rect 568900 690100 569100 690300
rect 569300 690100 569500 690300
rect 569700 690100 569900 690300
rect 570100 690100 570300 690300
rect 570500 690100 570700 690300
rect 570900 690100 571100 690300
rect 571300 690100 571500 690300
rect 571700 690100 571840 690300
rect 548409 689982 548419 690032
rect 541969 689918 542229 689952
rect 544607 689922 544721 689928
rect 541967 689912 542229 689918
rect 541967 689842 541979 689912
rect 542069 689842 542119 689912
rect 542209 689842 542229 689912
rect 541967 689836 542229 689842
rect 544447 689912 544561 689918
rect 544447 689842 544459 689912
rect 544549 689842 544561 689912
rect 544607 689852 544619 689922
rect 544709 689852 544721 689922
rect 544607 689846 544721 689852
rect 546907 689922 547011 689928
rect 546907 689852 546919 689922
rect 546999 689852 547011 689922
rect 546907 689846 547011 689852
rect 547077 689922 547181 689928
rect 547077 689852 547089 689922
rect 547169 689852 547181 689922
rect 547077 689846 547181 689852
rect 566260 689900 571840 690100
rect 544447 689836 544561 689842
rect 541969 689802 542229 689836
rect 47100 689600 47400 689800
rect 541959 689722 541969 689772
rect 540359 689704 541969 689722
rect 542049 689722 542059 689772
rect 542129 689722 542139 689772
rect 542049 689704 542139 689722
rect 542219 689722 542229 689772
rect 544449 689722 544459 689782
rect 542219 689704 544459 689722
rect 544539 689722 544549 689782
rect 544619 689722 544629 689782
rect 544539 689704 544629 689722
rect 544709 689722 544719 689782
rect 546909 689722 546919 689762
rect 544709 689704 546919 689722
rect 546999 689722 547009 689762
rect 547079 689722 547089 689762
rect 546999 689704 547089 689722
rect 547169 689722 547179 689762
rect 547169 689704 548799 689722
rect 540359 689682 540380 689704
rect 540368 689670 540380 689682
rect 541356 689682 541616 689704
rect 541356 689670 541368 689682
rect 540368 689664 541368 689670
rect 541604 689670 541616 689682
rect 542592 689682 542852 689704
rect 542592 689670 542604 689682
rect 541604 689664 542604 689670
rect 542840 689670 542852 689682
rect 543828 689682 544088 689704
rect 543828 689670 543840 689682
rect 542840 689664 543840 689670
rect 544076 689670 544088 689682
rect 545064 689682 545324 689704
rect 545064 689670 545076 689682
rect 544076 689664 545076 689670
rect 545312 689670 545324 689682
rect 546300 689682 546560 689704
rect 547536 689682 547796 689704
rect 546300 689670 546312 689682
rect 545312 689664 546312 689670
rect 546548 689670 546560 689682
rect 547536 689670 547548 689682
rect 546548 689664 547548 689670
rect 547784 689670 547796 689682
rect 548772 689682 548799 689704
rect 566260 689700 566300 689900
rect 566500 689700 566700 689900
rect 566900 689700 567100 689900
rect 567300 689700 567500 689900
rect 567700 689700 567900 689900
rect 568100 689700 568300 689900
rect 568500 689700 568700 689900
rect 568900 689700 569100 689900
rect 569300 689700 569500 689900
rect 569700 689700 569900 689900
rect 570100 689700 570300 689900
rect 570500 689700 570700 689900
rect 570900 689700 571100 689900
rect 571300 689700 571500 689900
rect 571700 689700 571840 689900
rect 548772 689670 548784 689682
rect 547784 689664 548784 689670
rect 47100 689500 47200 689600
rect 47300 689500 47400 689600
rect 540281 689642 540327 689654
rect 540281 689574 540287 689642
rect 540321 689632 540327 689642
rect 541409 689642 541455 689654
rect 541517 689642 541563 689654
rect 541409 689632 541415 689642
rect 540321 689602 541415 689632
rect 540321 689574 541089 689602
rect 540281 689562 541089 689574
rect 47100 689400 47400 689500
rect 540289 689546 541089 689562
rect 541169 689546 541239 689602
rect 541319 689574 541415 689602
rect 541557 689632 541563 689642
rect 542645 689642 542691 689654
rect 542753 689642 542799 689654
rect 543881 689642 543927 689654
rect 543989 689642 544035 689654
rect 542645 689632 542651 689642
rect 541557 689574 542651 689632
rect 542793 689632 542799 689642
rect 543879 689632 543887 689642
rect 542793 689602 543887 689632
rect 542793 689574 543579 689602
rect 541319 689572 541419 689574
rect 541549 689572 542659 689574
rect 542789 689572 543579 689574
rect 541319 689546 543579 689572
rect 543659 689546 543729 689602
rect 543809 689574 543887 689602
rect 544029 689632 544035 689642
rect 545117 689642 545163 689654
rect 545225 689642 545271 689654
rect 545117 689632 545123 689642
rect 544029 689574 545123 689632
rect 545265 689632 545271 689642
rect 546353 689642 546399 689654
rect 546461 689642 546507 689654
rect 547589 689642 547635 689654
rect 547697 689642 547743 689654
rect 546353 689632 546359 689642
rect 545265 689602 546359 689632
rect 545265 689574 546069 689602
rect 543809 689572 543889 689574
rect 544019 689572 545129 689574
rect 545259 689572 546069 689574
rect 543809 689546 546069 689572
rect 546149 689546 546209 689602
rect 546289 689574 546359 689602
rect 546501 689632 546509 689642
rect 547589 689632 547595 689642
rect 546501 689574 547595 689632
rect 547737 689632 547743 689642
rect 548825 689642 548871 689654
rect 548825 689632 548831 689642
rect 547737 689574 548831 689632
rect 548865 689574 548871 689642
rect 546289 689572 546369 689574
rect 546499 689572 547599 689574
rect 547729 689572 548871 689574
rect 546289 689562 548871 689572
rect 546289 689546 548869 689562
rect 540289 689512 540380 689546
rect 541356 689512 541616 689546
rect 542592 689512 542852 689546
rect 543828 689512 544088 689546
rect 545064 689512 545324 689546
rect 546300 689512 546560 689546
rect 547536 689512 547796 689546
rect 548772 689512 548869 689546
rect 540289 689492 540699 689512
rect 540689 689452 540699 689492
rect 540779 689492 540869 689512
rect 540779 689452 540789 689492
rect 540859 689452 540869 689492
rect 540949 689492 543219 689512
rect 540949 689452 540959 689492
rect 543209 689452 543219 689492
rect 543299 689492 543389 689512
rect 543299 689452 543309 689492
rect 543379 689452 543389 689492
rect 543469 689492 545709 689512
rect 543469 689452 543479 689492
rect 545699 689442 545709 689492
rect 545789 689492 545879 689512
rect 545789 689442 545799 689492
rect 545869 689442 545879 689492
rect 545959 689492 548159 689512
rect 545959 689442 545969 689492
rect 548149 689452 548159 689492
rect 548239 689492 548329 689512
rect 548239 689452 548249 689492
rect 548319 689452 548329 689492
rect 548409 689492 548869 689512
rect 566260 689520 571840 689700
rect 566260 689500 571820 689520
rect 548409 689452 548419 689492
rect 43870 689383 45430 689390
rect 43870 689349 44143 689383
rect 44211 689349 44301 689383
rect 44369 689349 44459 689383
rect 44527 689349 44617 689383
rect 44685 689349 44775 689383
rect 44843 689349 44933 689383
rect 45001 689349 45091 689383
rect 45159 689349 45430 689383
rect 43870 689340 45430 689349
rect 541967 689382 542071 689388
rect 541967 689302 541979 689382
rect 542059 689302 542071 689382
rect 541967 689296 542071 689302
rect 542137 689382 542241 689388
rect 542137 689302 542149 689382
rect 542229 689302 542241 689382
rect 542137 689296 542241 689302
rect 544447 689382 544551 689388
rect 544447 689302 544459 689382
rect 544539 689302 544551 689382
rect 544447 689296 544551 689302
rect 544617 689382 544721 689388
rect 544617 689302 544629 689382
rect 544709 689302 544721 689382
rect 544617 689296 544721 689302
rect 546907 689382 547011 689388
rect 546907 689302 546919 689382
rect 546999 689302 547011 689382
rect 546907 689296 547011 689302
rect 547077 689382 547181 689388
rect 547077 689302 547089 689382
rect 547169 689302 547181 689382
rect 547077 689296 547181 689302
rect 566260 689300 566300 689500
rect 566500 689300 566700 689500
rect 566900 689300 567100 689500
rect 567300 689300 567500 689500
rect 567700 689300 567900 689500
rect 568100 689300 568300 689500
rect 568500 689300 568700 689500
rect 568900 689300 569100 689500
rect 569300 689300 569500 689500
rect 569700 689300 569900 689500
rect 570100 689300 570300 689500
rect 570500 689300 570700 689500
rect 570900 689300 571100 689500
rect 571300 689300 571500 689500
rect 571700 689300 571820 689500
rect 44510 689287 44520 689290
rect 44314 689281 44520 689287
rect 44780 689287 44790 689290
rect 44780 689281 44988 689287
rect 44314 689247 44326 689281
rect 44976 689247 44988 689281
rect 44314 689241 44520 689247
rect 44510 689081 44520 689241
rect 44314 689075 44520 689081
rect 44780 689241 44988 689247
rect 44780 689081 44790 689241
rect 541969 689192 541979 689252
rect 540369 689172 541979 689192
rect 542059 689192 542069 689252
rect 542139 689192 542149 689252
rect 542059 689172 542149 689192
rect 542229 689192 542239 689252
rect 544449 689192 544459 689262
rect 542229 689182 544459 689192
rect 544539 689192 544549 689262
rect 544619 689192 544629 689262
rect 544539 689182 544629 689192
rect 544709 689192 544719 689262
rect 546909 689192 546919 689252
rect 544709 689182 546919 689192
rect 542229 689172 546919 689182
rect 546999 689192 547009 689252
rect 547079 689192 547089 689252
rect 546999 689172 547089 689192
rect 547169 689192 547179 689252
rect 547169 689172 548809 689192
rect 540369 689170 548809 689172
rect 540368 689164 548809 689170
rect 540368 689130 540380 689164
rect 541356 689152 541616 689164
rect 541356 689130 541368 689152
rect 540368 689124 541368 689130
rect 541604 689130 541616 689152
rect 542592 689152 542852 689164
rect 542592 689130 542604 689152
rect 541604 689124 542604 689130
rect 542840 689130 542852 689152
rect 543828 689152 544088 689164
rect 543828 689130 543840 689152
rect 542840 689124 543840 689130
rect 544076 689130 544088 689152
rect 545064 689152 545324 689164
rect 545064 689130 545076 689152
rect 544076 689124 545076 689130
rect 545312 689130 545324 689152
rect 546300 689152 546560 689164
rect 546300 689130 546312 689152
rect 545312 689124 546312 689130
rect 546548 689130 546560 689152
rect 547536 689152 547796 689164
rect 547536 689130 547548 689152
rect 546548 689124 547548 689130
rect 547784 689130 547796 689152
rect 548772 689152 548809 689164
rect 548772 689130 548784 689152
rect 547784 689124 548784 689130
rect 540281 689102 540327 689114
rect 44780 689075 44988 689081
rect 44314 689041 44326 689075
rect 44976 689041 44988 689075
rect 44314 689035 44520 689041
rect 44510 689030 44520 689035
rect 44780 689035 44988 689041
rect 44780 689030 44790 689035
rect 540281 689034 540287 689102
rect 540321 689092 540327 689102
rect 541409 689102 541455 689114
rect 541517 689102 541563 689114
rect 541409 689092 541415 689102
rect 540321 689042 541415 689092
rect 540321 689034 540327 689042
rect 540281 689022 540327 689034
rect 541409 689034 541415 689042
rect 541557 689092 541563 689102
rect 542645 689102 542691 689114
rect 542753 689102 542799 689114
rect 543881 689102 543927 689114
rect 543989 689102 544035 689114
rect 542645 689092 542651 689102
rect 541557 689042 542651 689092
rect 541557 689034 541563 689042
rect 541409 689032 541419 689034
rect 541549 689032 541563 689034
rect 541409 689022 541455 689032
rect 541517 689022 541563 689032
rect 542645 689034 542651 689042
rect 542793 689092 542799 689102
rect 543879 689092 543887 689102
rect 542793 689042 543887 689092
rect 542793 689034 542799 689042
rect 542645 689032 542659 689034
rect 542789 689032 542799 689034
rect 543879 689034 543887 689042
rect 544029 689092 544035 689102
rect 545117 689102 545163 689114
rect 545225 689102 545271 689114
rect 546353 689102 546399 689114
rect 546461 689102 546507 689114
rect 545117 689092 545123 689102
rect 544029 689042 545123 689092
rect 544029 689034 544035 689042
rect 543879 689032 543889 689034
rect 544019 689032 544035 689034
rect 542645 689022 542691 689032
rect 542753 689022 542799 689032
rect 543881 689022 543927 689032
rect 543989 689022 544035 689032
rect 545117 689034 545123 689042
rect 545265 689092 545271 689102
rect 546349 689092 546359 689102
rect 545265 689042 546359 689092
rect 545265 689034 545271 689042
rect 545117 689032 545129 689034
rect 545259 689032 545271 689034
rect 546349 689032 546359 689042
rect 546501 689092 546507 689102
rect 547589 689102 547635 689114
rect 547697 689102 547743 689114
rect 547589 689092 547595 689102
rect 546501 689042 547595 689092
rect 546501 689034 546507 689042
rect 546489 689032 546507 689034
rect 545117 689022 545163 689032
rect 545225 689022 545271 689032
rect 546353 689022 546399 689032
rect 546461 689022 546507 689032
rect 547589 689034 547595 689042
rect 547737 689092 547743 689102
rect 548825 689102 548871 689114
rect 548825 689092 548831 689102
rect 547737 689042 548831 689092
rect 547737 689034 547743 689042
rect 547589 689032 547599 689034
rect 547729 689032 547743 689034
rect 547589 689022 547635 689032
rect 547697 689022 547743 689032
rect 548825 689034 548831 689042
rect 548865 689034 548871 689102
rect 548825 689022 548871 689034
rect 540368 689006 541368 689012
rect 540368 688992 540380 689006
rect 541356 688992 541368 689006
rect 541604 689006 542604 689012
rect 541604 688992 541616 689006
rect 43870 688973 45430 688980
rect 43870 688939 44143 688973
rect 44211 688939 44301 688973
rect 44369 688939 44459 688973
rect 44527 688939 44617 688973
rect 44685 688939 44775 688973
rect 44843 688939 44933 688973
rect 45001 688939 45091 688973
rect 45159 688939 45430 688973
rect 540359 688972 540380 688992
rect 541356 688972 541616 688992
rect 542592 688992 542604 689006
rect 542840 689006 543840 689012
rect 542840 688992 542852 689006
rect 543828 688992 543840 689006
rect 544076 689006 545076 689012
rect 544076 688992 544088 689006
rect 542592 688972 542852 688992
rect 543828 688972 544088 688992
rect 545064 688992 545076 689006
rect 545312 689006 546312 689012
rect 545312 688992 545324 689006
rect 546300 688992 546312 689006
rect 546548 689006 547548 689012
rect 546548 688992 546560 689006
rect 547536 688992 547548 689006
rect 547784 689006 548784 689012
rect 547784 688992 547796 689006
rect 548772 688992 548784 689006
rect 545064 688972 545324 688992
rect 546300 688972 546560 688992
rect 547536 688972 547796 688992
rect 548772 688972 548799 688992
rect 540359 688952 540699 688972
rect 43870 688930 45430 688939
rect 41900 688700 42200 688800
rect 41900 688600 42000 688700
rect 42100 688600 42200 688700
rect 41900 688500 42200 688600
rect 41900 688300 42000 688500
rect 42100 688490 42200 688500
rect 43870 688490 43950 688930
rect 44075 688889 44121 688901
rect 44075 688860 44081 688889
rect 44115 688860 44121 688889
rect 44233 688889 44279 688901
rect 44050 688790 44060 688860
rect 44130 688790 44140 688860
rect 44075 688570 44081 688790
rect 44115 688570 44121 688790
rect 44050 688500 44060 688570
rect 44130 688500 44140 688570
rect 42100 688310 43950 688490
rect 42100 688300 42200 688310
rect 41900 688200 42200 688300
rect 41900 688100 42000 688200
rect 42100 688100 42200 688200
rect 41900 688000 42200 688100
rect 43870 687870 43950 688310
rect 44075 687913 44081 688500
rect 44115 687913 44121 688500
rect 44233 688300 44239 688889
rect 44273 688300 44279 688889
rect 44391 688889 44437 688901
rect 44391 688860 44397 688889
rect 44431 688860 44437 688889
rect 44549 688889 44595 688901
rect 44370 688790 44380 688860
rect 44450 688790 44460 688860
rect 44391 688570 44397 688790
rect 44431 688570 44437 688790
rect 44370 688500 44380 688570
rect 44450 688500 44460 688570
rect 44210 688230 44220 688300
rect 44290 688230 44300 688300
rect 44233 688010 44239 688230
rect 44273 688010 44279 688230
rect 44210 687940 44220 688010
rect 44290 687940 44300 688010
rect 44075 687901 44121 687913
rect 44233 687913 44239 687940
rect 44273 687913 44279 687940
rect 44233 687901 44279 687913
rect 44391 687913 44397 688500
rect 44431 687913 44437 688500
rect 44549 688300 44555 688889
rect 44589 688300 44595 688889
rect 44707 688889 44753 688901
rect 44707 688860 44713 688889
rect 44747 688860 44753 688889
rect 44865 688889 44911 688901
rect 44680 688790 44690 688860
rect 44760 688790 44770 688860
rect 44707 688570 44713 688790
rect 44747 688570 44753 688790
rect 44680 688500 44690 688570
rect 44760 688500 44770 688570
rect 44520 688230 44530 688300
rect 44600 688230 44610 688300
rect 44549 688010 44555 688230
rect 44589 688010 44595 688230
rect 44520 687940 44530 688010
rect 44600 687940 44610 688010
rect 44391 687901 44437 687913
rect 44549 687913 44555 687940
rect 44589 687913 44595 687940
rect 44549 687901 44595 687913
rect 44707 687913 44713 688500
rect 44747 687913 44753 688500
rect 44865 688300 44871 688889
rect 44905 688300 44911 688889
rect 45023 688889 45069 688901
rect 45023 688860 45029 688889
rect 45063 688860 45069 688889
rect 45181 688889 45227 688901
rect 45000 688790 45010 688860
rect 45080 688790 45090 688860
rect 45023 688570 45029 688790
rect 45063 688570 45069 688790
rect 45000 688500 45010 688570
rect 45080 688500 45090 688570
rect 44840 688230 44850 688300
rect 44920 688230 44930 688300
rect 44865 688010 44871 688230
rect 44905 688010 44911 688230
rect 44840 687940 44850 688010
rect 44920 687940 44930 688010
rect 44707 687901 44753 687913
rect 44865 687913 44871 687940
rect 44905 687913 44911 687940
rect 44865 687901 44911 687913
rect 45023 687913 45029 688500
rect 45063 687913 45069 688500
rect 45181 688300 45187 688889
rect 45221 688300 45227 688889
rect 45160 688230 45170 688300
rect 45240 688230 45250 688300
rect 45181 688010 45187 688230
rect 45221 688010 45227 688230
rect 45160 687940 45170 688010
rect 45240 687940 45250 688010
rect 45023 687901 45069 687913
rect 45181 687913 45187 687940
rect 45221 687913 45227 687940
rect 45181 687901 45227 687913
rect 45350 687870 45430 688930
rect 540689 688912 540699 688952
rect 540779 688952 540869 688972
rect 540779 688912 540789 688952
rect 540859 688912 540869 688952
rect 540949 688952 542379 688972
rect 540949 688912 540959 688952
rect 542359 688922 542379 688952
rect 542459 688922 542489 688972
rect 542569 688952 543209 688972
rect 542569 688922 542589 688952
rect 542359 688892 542589 688922
rect 543199 688912 543209 688952
rect 543289 688952 543379 688972
rect 543289 688912 543299 688952
rect 543369 688912 543379 688952
rect 543459 688952 544789 688972
rect 543459 688912 543469 688952
rect 544769 688922 544789 688952
rect 544869 688922 544899 688972
rect 544979 688952 545699 688972
rect 544979 688922 544999 688952
rect 544769 688912 544999 688922
rect 545689 688912 545699 688952
rect 545779 688952 545869 688972
rect 545779 688912 545789 688952
rect 545859 688912 545869 688952
rect 545949 688952 547249 688972
rect 545949 688912 545959 688952
rect 547229 688912 547249 688952
rect 547329 688912 547359 688972
rect 547439 688952 548189 688972
rect 547439 688912 547459 688952
rect 548179 688912 548189 688952
rect 548269 688952 548359 688972
rect 548269 688912 548279 688952
rect 548349 688912 548359 688952
rect 548439 688952 548799 688972
rect 548439 688912 548449 688952
rect 547229 688892 547459 688912
rect 541969 688612 541979 688672
rect 540359 688592 541979 688612
rect 542059 688612 542069 688672
rect 542139 688612 542149 688672
rect 542059 688592 542149 688612
rect 542229 688612 542239 688672
rect 544449 688612 544459 688682
rect 542229 688602 544459 688612
rect 544539 688612 544549 688682
rect 544619 688612 544629 688682
rect 544539 688602 544629 688612
rect 544709 688612 544719 688682
rect 546909 688612 546919 688672
rect 544709 688602 546919 688612
rect 542229 688592 546919 688602
rect 546999 688612 547009 688672
rect 547079 688612 547089 688672
rect 546999 688592 547089 688612
rect 547169 688612 547179 688672
rect 547169 688592 548799 688612
rect 540359 688584 548799 688592
rect 540359 688572 540380 688584
rect 540368 688550 540380 688572
rect 541356 688572 541616 688584
rect 541356 688550 541368 688572
rect 540368 688544 541368 688550
rect 541604 688550 541616 688572
rect 542592 688572 542852 688584
rect 542592 688550 542604 688572
rect 541604 688544 542604 688550
rect 542840 688550 542852 688572
rect 543828 688572 544088 688584
rect 543828 688550 543840 688572
rect 542840 688544 543840 688550
rect 544076 688550 544088 688572
rect 545064 688572 545324 688584
rect 545064 688550 545076 688572
rect 544076 688544 545076 688550
rect 545312 688550 545324 688572
rect 546300 688572 546560 688584
rect 546300 688550 546312 688572
rect 545312 688544 546312 688550
rect 546548 688550 546560 688572
rect 547536 688572 547796 688584
rect 547536 688550 547548 688572
rect 546548 688544 547548 688550
rect 547784 688550 547796 688572
rect 548772 688572 548799 688584
rect 548772 688550 548784 688572
rect 547784 688544 548784 688550
rect 540281 688522 540327 688534
rect 540281 688454 540287 688522
rect 540321 688512 540327 688522
rect 541409 688522 541455 688534
rect 541517 688522 541563 688534
rect 541409 688512 541415 688522
rect 540321 688462 541415 688512
rect 540321 688454 540327 688462
rect 540281 688442 540327 688454
rect 541409 688454 541415 688462
rect 541557 688512 541563 688522
rect 542645 688522 542691 688534
rect 542753 688522 542799 688534
rect 542645 688512 542651 688522
rect 541557 688462 542651 688512
rect 541557 688454 541563 688462
rect 541409 688452 541419 688454
rect 541549 688452 541563 688454
rect 541409 688442 541455 688452
rect 541517 688442 541563 688452
rect 542645 688454 542651 688462
rect 542793 688512 542799 688522
rect 543881 688522 543927 688534
rect 543989 688522 544035 688534
rect 545117 688522 545163 688534
rect 545225 688522 545271 688534
rect 546353 688522 546399 688534
rect 546461 688522 546507 688534
rect 543881 688512 543887 688522
rect 542793 688462 543887 688512
rect 542793 688454 542799 688462
rect 542645 688452 542659 688454
rect 542789 688452 542799 688454
rect 542645 688442 542691 688452
rect 542753 688442 542799 688452
rect 543881 688454 543887 688462
rect 544029 688512 544039 688522
rect 545117 688512 545123 688522
rect 544029 688462 545123 688512
rect 543881 688452 543899 688454
rect 544029 688452 544039 688462
rect 545117 688454 545123 688462
rect 545265 688512 545271 688522
rect 546349 688512 546359 688522
rect 545265 688462 546359 688512
rect 545265 688454 545271 688462
rect 545117 688452 545129 688454
rect 545259 688452 545271 688454
rect 546349 688452 546359 688462
rect 546501 688512 546507 688522
rect 547589 688522 547635 688534
rect 547697 688522 547743 688534
rect 547589 688512 547595 688522
rect 546501 688462 547595 688512
rect 546501 688454 546507 688462
rect 546489 688452 546507 688454
rect 543881 688442 543927 688452
rect 543989 688442 544035 688452
rect 545117 688442 545163 688452
rect 545225 688442 545271 688452
rect 546353 688442 546399 688452
rect 546461 688442 546507 688452
rect 547589 688454 547595 688462
rect 547737 688512 547743 688522
rect 548825 688522 548871 688534
rect 548825 688512 548831 688522
rect 547737 688462 548831 688512
rect 547737 688454 547743 688462
rect 547589 688452 547599 688454
rect 547729 688452 547743 688454
rect 547589 688442 547635 688452
rect 547697 688442 547743 688452
rect 548825 688454 548831 688462
rect 548865 688454 548871 688522
rect 548825 688442 548871 688454
rect 540368 688426 541368 688432
rect 540368 688412 540380 688426
rect 541356 688412 541368 688426
rect 541604 688426 542604 688432
rect 541604 688412 541616 688426
rect 540359 688392 540380 688412
rect 541356 688392 541616 688412
rect 542592 688412 542604 688426
rect 542840 688426 543840 688432
rect 542840 688412 542852 688426
rect 543828 688412 543840 688426
rect 544076 688426 545076 688432
rect 544076 688412 544088 688426
rect 545064 688412 545076 688426
rect 545312 688426 546312 688432
rect 545312 688412 545324 688426
rect 542592 688392 542852 688412
rect 543828 688392 544088 688412
rect 545064 688392 545324 688412
rect 546300 688412 546312 688426
rect 546548 688426 547548 688432
rect 546548 688412 546560 688426
rect 547536 688412 547548 688426
rect 547784 688426 548784 688432
rect 547784 688412 547796 688426
rect 548772 688412 548784 688426
rect 546300 688392 546560 688412
rect 547536 688392 547796 688412
rect 548772 688392 548799 688412
rect 540359 688372 540699 688392
rect 540689 688332 540699 688372
rect 540779 688372 540869 688392
rect 540779 688332 540789 688372
rect 540859 688332 540869 688372
rect 540949 688372 542379 688392
rect 540949 688332 540959 688372
rect 542359 688312 542379 688372
rect 542459 688312 542489 688392
rect 542569 688372 543209 688392
rect 542569 688312 542589 688372
rect 543199 688332 543209 688372
rect 543289 688372 543379 688392
rect 543289 688332 543299 688372
rect 543369 688332 543379 688372
rect 543459 688372 544789 688392
rect 543459 688332 543469 688372
rect 544769 688332 544789 688372
rect 544869 688332 544899 688392
rect 544979 688372 545699 688392
rect 544979 688332 544999 688372
rect 544769 688312 544999 688332
rect 545689 688322 545699 688372
rect 545779 688372 545869 688392
rect 545779 688322 545789 688372
rect 545859 688322 545869 688372
rect 545949 688372 547249 688392
rect 545949 688322 545959 688372
rect 547229 688332 547249 688372
rect 547329 688332 547359 688392
rect 547439 688372 548189 688392
rect 547439 688332 547459 688372
rect 548179 688332 548189 688372
rect 548269 688372 548359 688392
rect 548269 688332 548279 688372
rect 548349 688332 548359 688372
rect 548439 688372 548799 688392
rect 548439 688332 548449 688372
rect 547229 688312 547459 688332
rect 542359 688302 542589 688312
rect 554109 688302 554539 688422
rect 43870 687863 45430 687870
rect 43870 687829 44143 687863
rect 44211 687829 44301 687863
rect 44369 687829 44459 687863
rect 44527 687829 44617 687863
rect 44685 687829 44775 687863
rect 44843 687829 44933 687863
rect 45001 687829 45091 687863
rect 45159 687829 45430 687863
rect 43870 687820 45430 687829
rect 534609 688132 535039 688252
rect 541967 688222 542081 688228
rect 541967 688142 541979 688222
rect 542069 688142 542081 688222
rect 541967 688136 542081 688142
rect 542127 688222 542241 688228
rect 542127 688142 542139 688222
rect 542229 688142 542241 688222
rect 542127 688136 542241 688142
rect 544447 688212 544551 688218
rect 544447 688142 544459 688212
rect 544539 688142 544551 688212
rect 544447 688136 544551 688142
rect 544617 688212 544721 688218
rect 544617 688142 544629 688212
rect 544709 688142 544721 688212
rect 544617 688136 544721 688142
rect 546907 688212 547011 688218
rect 546907 688142 546919 688212
rect 546999 688142 547011 688212
rect 546907 688136 547011 688142
rect 547077 688212 547181 688218
rect 547077 688142 547089 688212
rect 547169 688142 547181 688212
rect 547077 688136 547181 688142
rect 554109 688162 554129 688302
rect 554259 688162 554389 688302
rect 554519 688162 554539 688302
rect 534609 687992 534629 688132
rect 534759 687992 534879 688132
rect 535009 687992 535039 688132
rect 541969 688032 541979 688092
rect 540359 688012 541979 688032
rect 542059 688032 542069 688092
rect 542139 688032 542149 688092
rect 542059 688012 542149 688032
rect 542229 688032 542239 688092
rect 544449 688032 544459 688102
rect 542229 688022 544459 688032
rect 544539 688032 544549 688102
rect 544619 688032 544629 688102
rect 544539 688022 544629 688032
rect 544709 688032 544719 688102
rect 546909 688032 546919 688092
rect 544709 688022 546919 688032
rect 542229 688012 546919 688022
rect 546999 688032 547009 688092
rect 547079 688032 547089 688092
rect 546999 688012 547089 688032
rect 547169 688032 547179 688092
rect 547169 688012 548799 688032
rect 540359 688004 548799 688012
rect 540359 687992 540380 688004
rect 534609 687967 535039 687992
rect 540368 687970 540380 687992
rect 541356 687992 541616 688004
rect 541356 687970 541368 687992
rect 534609 687955 535143 687967
rect 44510 687767 44520 687770
rect 44314 687761 44520 687767
rect 44780 687767 44790 687770
rect 44780 687761 44988 687767
rect 44314 687727 44326 687761
rect 44976 687727 44988 687761
rect 44314 687721 44520 687727
rect 44510 687560 44520 687721
rect 43821 687554 44520 687560
rect 44780 687721 44988 687727
rect 44780 687560 44790 687721
rect 44780 687554 45489 687560
rect 43821 687520 43833 687554
rect 45477 687520 45489 687554
rect 43821 687514 44520 687520
rect 44510 687510 44520 687514
rect 44780 687514 45489 687520
rect 44780 687510 44790 687514
rect 42250 687460 42260 687490
rect 42240 687410 42260 687460
rect 42250 687380 42260 687410
rect 42370 687460 42380 687490
rect 42500 687460 42510 687490
rect 42370 687410 42510 687460
rect 42370 687380 42380 687410
rect 42500 687380 42510 687410
rect 42620 687460 42630 687490
rect 46650 687460 46660 687490
rect 42620 687452 46660 687460
rect 42620 687418 43152 687452
rect 43320 687418 43410 687452
rect 43578 687418 43668 687452
rect 43836 687418 43926 687452
rect 44094 687418 44184 687452
rect 44352 687418 44442 687452
rect 44610 687418 44700 687452
rect 44868 687418 44958 687452
rect 45126 687418 45216 687452
rect 45384 687418 45474 687452
rect 45642 687418 45732 687452
rect 45900 687418 45990 687452
rect 46158 687418 46660 687452
rect 42620 687410 46660 687418
rect 42620 687380 42630 687410
rect 46650 687380 46660 687410
rect 46770 687460 46780 687490
rect 46900 687460 46910 687490
rect 46770 687410 46910 687460
rect 46770 687380 46780 687410
rect 46900 687380 46910 687410
rect 47020 687460 47030 687490
rect 47020 687410 47040 687460
rect 47020 687380 47030 687410
rect 43084 687368 43130 687380
rect 43084 687340 43090 687368
rect 43124 687340 43130 687368
rect 43342 687368 43388 687380
rect 43060 687270 43070 687340
rect 43140 687270 43150 687340
rect 43084 687160 43090 687270
rect 43124 687160 43130 687270
rect 43060 687090 43070 687160
rect 43140 687090 43150 687160
rect 43084 686392 43090 687090
rect 43124 686392 43130 687090
rect 43342 686670 43348 687368
rect 43382 686670 43388 687368
rect 43600 687368 43646 687380
rect 43600 687340 43606 687368
rect 43640 687340 43646 687368
rect 43858 687368 43904 687380
rect 43580 687270 43590 687340
rect 43660 687270 43670 687340
rect 43600 687160 43606 687270
rect 43640 687160 43646 687270
rect 43580 687090 43590 687160
rect 43660 687090 43670 687160
rect 43320 686600 43330 686670
rect 43400 686600 43410 686670
rect 43342 686490 43348 686600
rect 43382 686490 43388 686600
rect 43320 686420 43330 686490
rect 43400 686420 43410 686490
rect 43084 686380 43130 686392
rect 43342 686392 43348 686420
rect 43382 686392 43388 686420
rect 43342 686380 43388 686392
rect 43600 686392 43606 687090
rect 43640 686392 43646 687090
rect 43858 686670 43864 687368
rect 43898 686670 43904 687368
rect 44116 687368 44162 687380
rect 44116 687340 44122 687368
rect 44156 687340 44162 687368
rect 44374 687368 44420 687380
rect 44090 687270 44100 687340
rect 44170 687270 44180 687340
rect 44116 687160 44122 687270
rect 44156 687160 44162 687270
rect 44090 687090 44100 687160
rect 44170 687090 44180 687160
rect 43830 686600 43840 686670
rect 43910 686600 43920 686670
rect 43858 686490 43864 686600
rect 43898 686490 43904 686600
rect 43830 686420 43840 686490
rect 43910 686420 43920 686490
rect 43600 686380 43646 686392
rect 43858 686392 43864 686420
rect 43898 686392 43904 686420
rect 43858 686380 43904 686392
rect 44116 686392 44122 687090
rect 44156 686392 44162 687090
rect 44374 686670 44380 687368
rect 44414 686670 44420 687368
rect 44632 687368 44678 687380
rect 44632 687340 44638 687368
rect 44672 687340 44678 687368
rect 44890 687368 44936 687380
rect 44610 687270 44620 687340
rect 44690 687270 44700 687340
rect 44632 687160 44638 687270
rect 44672 687160 44678 687270
rect 44610 687090 44620 687160
rect 44690 687090 44700 687160
rect 44350 686600 44360 686670
rect 44430 686600 44440 686670
rect 44374 686490 44380 686600
rect 44414 686490 44420 686600
rect 44350 686420 44360 686490
rect 44430 686420 44440 686490
rect 44116 686380 44162 686392
rect 44374 686392 44380 686420
rect 44414 686392 44420 686420
rect 44374 686380 44420 686392
rect 44632 686392 44638 687090
rect 44672 686392 44678 687090
rect 44890 686670 44896 687368
rect 44930 686670 44936 687368
rect 45148 687368 45194 687380
rect 45148 687340 45154 687368
rect 45188 687340 45194 687368
rect 45406 687368 45452 687380
rect 45120 687270 45130 687340
rect 45200 687270 45210 687340
rect 45148 687160 45154 687270
rect 45188 687160 45194 687270
rect 45120 687090 45130 687160
rect 45200 687090 45210 687160
rect 44870 686600 44880 686670
rect 44950 686600 44960 686670
rect 44890 686490 44896 686600
rect 44930 686490 44936 686600
rect 44870 686420 44880 686490
rect 44950 686420 44960 686490
rect 44632 686380 44678 686392
rect 44890 686392 44896 686420
rect 44930 686392 44936 686420
rect 44890 686380 44936 686392
rect 45148 686392 45154 687090
rect 45188 686392 45194 687090
rect 45406 686670 45412 687368
rect 45446 686670 45452 687368
rect 45664 687368 45710 687380
rect 45664 687340 45670 687368
rect 45704 687340 45710 687368
rect 45922 687368 45968 687380
rect 45640 687270 45650 687340
rect 45720 687270 45730 687340
rect 45664 687160 45670 687270
rect 45704 687160 45710 687270
rect 45640 687090 45650 687160
rect 45720 687090 45730 687160
rect 45380 686600 45390 686670
rect 45460 686600 45470 686670
rect 45406 686490 45412 686600
rect 45446 686490 45452 686600
rect 45380 686420 45390 686490
rect 45460 686420 45470 686490
rect 45148 686380 45194 686392
rect 45406 686392 45412 686420
rect 45446 686392 45452 686420
rect 45406 686380 45452 686392
rect 45664 686392 45670 687090
rect 45704 686392 45710 687090
rect 45922 686670 45928 687368
rect 45962 686670 45968 687368
rect 46180 687368 46226 687380
rect 46180 687340 46186 687368
rect 46220 687340 46226 687368
rect 46160 687270 46170 687340
rect 46240 687270 46250 687340
rect 46180 687160 46186 687270
rect 46220 687160 46226 687270
rect 46160 687090 46170 687160
rect 46240 687090 46250 687160
rect 45900 686600 45910 686670
rect 45980 686600 45990 686670
rect 45922 686490 45928 686600
rect 45962 686490 45968 686600
rect 45900 686420 45910 686490
rect 45980 686420 45990 686490
rect 45664 686380 45710 686392
rect 45922 686392 45928 686420
rect 45962 686392 45968 686420
rect 45922 686380 45968 686392
rect 46180 686392 46186 687090
rect 46220 686392 46226 687090
rect 46180 686380 46226 686392
rect 534609 686841 534740 687955
rect 535137 686841 535143 687955
rect 537165 687955 537574 687967
rect 540368 687964 541368 687970
rect 541604 687970 541616 687992
rect 542592 687992 542852 688004
rect 542592 687970 542604 687992
rect 541604 687964 542604 687970
rect 542840 687970 542852 687992
rect 543828 687992 544088 688004
rect 543828 687970 543840 687992
rect 542840 687964 543840 687970
rect 544076 687970 544088 687992
rect 545064 687992 545324 688004
rect 545064 687970 545076 687992
rect 544076 687964 545076 687970
rect 545312 687970 545324 687992
rect 546300 687992 546560 688004
rect 546300 687970 546312 687992
rect 545312 687964 546312 687970
rect 546548 687970 546560 687992
rect 547536 687992 547796 688004
rect 547536 687970 547548 687992
rect 546548 687964 547548 687970
rect 547784 687970 547796 687992
rect 548772 687992 548799 688004
rect 548772 687970 548784 687992
rect 547784 687964 548784 687970
rect 554109 687967 554539 688162
rect 537165 687862 537171 687955
rect 534609 686829 535143 686841
rect 537039 686841 537171 687862
rect 537568 687422 537574 687955
rect 551794 687955 552203 687967
rect 540281 687942 540327 687954
rect 540281 687874 540287 687942
rect 540321 687932 540327 687942
rect 541409 687942 541455 687954
rect 541517 687942 541563 687954
rect 541409 687932 541415 687942
rect 540321 687882 541415 687932
rect 540321 687874 540327 687882
rect 540281 687862 540327 687874
rect 541409 687874 541415 687882
rect 541557 687932 541563 687942
rect 542645 687942 542691 687954
rect 542753 687942 542799 687954
rect 543881 687942 543927 687954
rect 543989 687942 544035 687954
rect 542645 687932 542651 687942
rect 541557 687882 542651 687932
rect 541557 687874 541563 687882
rect 541409 687872 541419 687874
rect 541549 687872 541563 687874
rect 541409 687862 541455 687872
rect 541517 687862 541563 687872
rect 542645 687874 542651 687882
rect 542793 687932 542799 687942
rect 543879 687932 543887 687942
rect 542793 687882 543887 687932
rect 542793 687874 542799 687882
rect 542645 687872 542659 687874
rect 542789 687872 542799 687874
rect 543879 687874 543887 687882
rect 544029 687932 544035 687942
rect 545117 687942 545163 687954
rect 545225 687942 545271 687954
rect 546353 687942 546399 687954
rect 546461 687942 546507 687954
rect 545117 687932 545123 687942
rect 544029 687882 545123 687932
rect 544029 687874 544035 687882
rect 543879 687872 543889 687874
rect 544019 687872 544035 687874
rect 542645 687862 542691 687872
rect 542753 687862 542799 687872
rect 543881 687862 543927 687872
rect 543989 687862 544035 687872
rect 545117 687874 545123 687882
rect 545265 687932 545271 687942
rect 546349 687932 546359 687942
rect 545265 687882 546359 687932
rect 545265 687874 545271 687882
rect 545117 687872 545129 687874
rect 545259 687872 545271 687874
rect 546349 687872 546359 687882
rect 546501 687932 546507 687942
rect 547589 687942 547635 687954
rect 547697 687942 547743 687954
rect 547589 687932 547595 687942
rect 546501 687882 547595 687932
rect 546501 687874 546507 687882
rect 546489 687872 546507 687874
rect 545117 687862 545163 687872
rect 545225 687862 545271 687872
rect 546353 687862 546399 687872
rect 546461 687862 546507 687872
rect 547589 687874 547595 687882
rect 547737 687932 547743 687942
rect 548825 687942 548871 687954
rect 548825 687932 548831 687942
rect 547737 687882 548831 687932
rect 547737 687874 547743 687882
rect 547589 687872 547599 687874
rect 547729 687872 547743 687874
rect 547589 687862 547635 687872
rect 547697 687862 547743 687872
rect 548825 687874 548831 687882
rect 548865 687874 548871 687942
rect 548825 687862 548871 687874
rect 551794 687862 551800 687955
rect 540368 687846 541368 687852
rect 540368 687822 540380 687846
rect 540359 687812 540380 687822
rect 541356 687822 541368 687846
rect 541604 687846 542604 687852
rect 541604 687822 541616 687846
rect 541356 687812 541616 687822
rect 542592 687822 542604 687846
rect 542840 687846 543840 687852
rect 542840 687822 542852 687846
rect 542592 687812 542852 687822
rect 543828 687822 543840 687846
rect 544076 687846 545076 687852
rect 544076 687822 544088 687846
rect 543828 687812 544088 687822
rect 545064 687822 545076 687846
rect 545312 687846 546312 687852
rect 545312 687822 545324 687846
rect 545064 687812 545324 687822
rect 546300 687822 546312 687846
rect 546548 687846 547548 687852
rect 546548 687822 546560 687846
rect 546300 687812 546560 687822
rect 547536 687822 547548 687846
rect 547784 687846 548784 687852
rect 547784 687822 547796 687846
rect 547536 687812 547796 687822
rect 548772 687822 548784 687846
rect 548772 687812 548799 687822
rect 540359 687802 542380 687812
rect 540359 687782 540679 687802
rect 540669 687722 540679 687782
rect 540759 687782 540889 687802
rect 540759 687722 540769 687782
rect 540879 687722 540889 687782
rect 540969 687782 542380 687802
rect 540969 687722 540979 687782
rect 542359 687750 542380 687782
rect 542460 687750 542500 687812
rect 542580 687782 543209 687812
rect 542580 687750 542590 687782
rect 543199 687752 543209 687782
rect 543289 687782 543379 687812
rect 543289 687752 543299 687782
rect 543369 687752 543379 687782
rect 543459 687782 544789 687812
rect 543459 687752 543469 687782
rect 544769 687752 544789 687782
rect 544869 687752 544899 687812
rect 544979 687782 545699 687812
rect 544979 687752 544999 687782
rect 545689 687752 545699 687782
rect 545779 687782 545869 687812
rect 545779 687752 545789 687782
rect 545859 687752 545869 687782
rect 545949 687782 547249 687812
rect 545949 687752 545959 687782
rect 547229 687752 547249 687782
rect 547329 687752 547359 687812
rect 547439 687782 548189 687812
rect 547439 687752 547459 687782
rect 548179 687752 548189 687782
rect 548269 687782 548359 687812
rect 548269 687752 548279 687782
rect 548349 687752 548359 687782
rect 548439 687782 548799 687812
rect 548439 687752 548449 687782
rect 542359 687732 542589 687750
rect 544769 687732 544999 687752
rect 547229 687732 547459 687752
rect 540089 687492 540099 687562
rect 538519 687482 540099 687492
rect 540179 687492 540189 687562
rect 540319 687492 540329 687562
rect 540179 687482 540329 687492
rect 540409 687492 540419 687562
rect 542639 687492 542649 687552
rect 540409 687482 542649 687492
rect 538519 687472 542649 687482
rect 542729 687492 542739 687552
rect 542809 687492 542819 687552
rect 542729 687472 542819 687492
rect 542899 687492 542909 687552
rect 545099 687492 545109 687552
rect 542899 687472 545109 687492
rect 545189 687492 545199 687552
rect 545289 687492 545299 687552
rect 545189 687472 545299 687492
rect 545379 687492 545389 687552
rect 547549 687492 547559 687552
rect 545379 687472 547559 687492
rect 547639 687492 547649 687552
rect 547739 687492 547749 687552
rect 547639 687472 547749 687492
rect 547829 687492 547839 687552
rect 550059 687492 550069 687552
rect 547829 687472 550069 687492
rect 550149 687492 550159 687552
rect 550229 687492 550239 687552
rect 550149 687472 550239 687492
rect 550319 687492 550329 687552
rect 550319 687472 550669 687492
rect 538519 687464 550669 687472
rect 538519 687442 538540 687464
rect 538528 687430 538540 687442
rect 539516 687442 539776 687464
rect 539516 687430 539528 687442
rect 538528 687424 539528 687430
rect 539764 687430 539776 687442
rect 540752 687442 541012 687464
rect 540752 687430 540764 687442
rect 539764 687424 540764 687430
rect 541000 687430 541012 687442
rect 541988 687442 542248 687464
rect 541988 687430 542000 687442
rect 541000 687424 542000 687430
rect 542236 687430 542248 687442
rect 543224 687442 543484 687464
rect 543224 687430 543236 687442
rect 542236 687424 543236 687430
rect 543472 687430 543484 687442
rect 544460 687442 544720 687464
rect 544460 687430 544472 687442
rect 543472 687424 544472 687430
rect 544708 687430 544720 687442
rect 545696 687442 545956 687464
rect 545696 687430 545708 687442
rect 544708 687424 545708 687430
rect 545944 687430 545956 687442
rect 546932 687442 547192 687464
rect 546932 687430 546944 687442
rect 545944 687424 546944 687430
rect 547180 687430 547192 687442
rect 548168 687442 548428 687464
rect 548168 687430 548180 687442
rect 547180 687424 548180 687430
rect 548416 687430 548428 687442
rect 549404 687442 549664 687464
rect 549404 687430 549416 687442
rect 548416 687424 549416 687430
rect 549652 687430 549664 687442
rect 550640 687442 550669 687464
rect 550640 687430 550652 687442
rect 549652 687424 550652 687430
rect 551669 687422 551800 687862
rect 537568 687414 538479 687422
rect 550699 687414 551800 687422
rect 537568 687402 538487 687414
rect 537568 687334 538447 687402
rect 538481 687392 538487 687402
rect 539569 687402 539615 687414
rect 539677 687402 539723 687414
rect 539569 687392 539575 687402
rect 538481 687352 539575 687392
rect 538481 687334 538487 687352
rect 537568 687322 538487 687334
rect 539569 687334 539575 687352
rect 539717 687392 539723 687402
rect 540805 687402 540851 687414
rect 540913 687402 540959 687414
rect 542041 687402 542087 687414
rect 542149 687402 542195 687414
rect 540805 687392 540811 687402
rect 539717 687352 540811 687392
rect 539717 687334 539723 687352
rect 539569 687332 539579 687334
rect 539709 687332 539723 687334
rect 539569 687322 539615 687332
rect 539677 687322 539723 687332
rect 540805 687334 540811 687352
rect 540953 687392 540959 687402
rect 542039 687392 542047 687402
rect 540953 687352 542047 687392
rect 540953 687334 540959 687352
rect 540805 687332 540819 687334
rect 540949 687332 540959 687334
rect 542039 687334 542047 687352
rect 542189 687392 542195 687402
rect 543277 687402 543323 687414
rect 543385 687402 543431 687414
rect 543277 687392 543283 687402
rect 542189 687352 543283 687392
rect 542189 687334 542195 687352
rect 542039 687332 542049 687334
rect 542179 687332 542195 687334
rect 540805 687322 540851 687332
rect 540913 687322 540959 687332
rect 542041 687322 542087 687332
rect 542149 687322 542195 687332
rect 543277 687334 543283 687352
rect 543425 687392 543431 687402
rect 544513 687402 544559 687414
rect 544621 687402 544667 687414
rect 545749 687402 545795 687414
rect 545857 687402 545903 687414
rect 544513 687392 544519 687402
rect 543425 687352 544519 687392
rect 543425 687334 543431 687352
rect 543277 687332 543289 687334
rect 543419 687332 543431 687334
rect 543277 687322 543323 687332
rect 543385 687322 543431 687332
rect 544513 687334 544519 687352
rect 544661 687392 544669 687402
rect 545749 687392 545755 687402
rect 544661 687352 545755 687392
rect 544661 687334 544669 687352
rect 544513 687332 544529 687334
rect 544659 687332 544669 687334
rect 545749 687334 545755 687352
rect 545897 687392 545903 687402
rect 546985 687402 547031 687414
rect 547093 687402 547139 687414
rect 548221 687402 548267 687414
rect 548329 687402 548375 687414
rect 546985 687392 546991 687402
rect 545897 687352 546991 687392
rect 545897 687334 545903 687352
rect 545749 687332 545759 687334
rect 545889 687332 545903 687334
rect 544513 687322 544559 687332
rect 544621 687322 544667 687332
rect 545749 687322 545795 687332
rect 545857 687322 545903 687332
rect 546985 687334 546991 687352
rect 547133 687392 547139 687402
rect 548219 687392 548227 687402
rect 547133 687352 548227 687392
rect 547133 687334 547139 687352
rect 546985 687332 546999 687334
rect 547129 687332 547139 687334
rect 548219 687334 548227 687352
rect 548369 687392 548375 687402
rect 549457 687402 549503 687414
rect 549565 687402 549611 687414
rect 549457 687392 549463 687402
rect 548369 687352 549463 687392
rect 548369 687334 548375 687352
rect 548219 687332 548229 687334
rect 548359 687332 548375 687334
rect 546985 687322 547031 687332
rect 547093 687322 547139 687332
rect 548221 687322 548267 687332
rect 548329 687322 548375 687332
rect 549457 687334 549463 687352
rect 549605 687392 549611 687402
rect 550693 687402 551800 687414
rect 550693 687392 550699 687402
rect 549605 687352 550699 687392
rect 549605 687334 549611 687352
rect 549457 687332 549469 687334
rect 549599 687332 549611 687334
rect 549457 687322 549503 687332
rect 549565 687322 549611 687332
rect 550693 687334 550699 687352
rect 550733 687334 551800 687402
rect 550693 687322 551800 687334
rect 537568 686882 537574 687322
rect 538528 687306 539528 687312
rect 538528 687292 538540 687306
rect 538519 687272 538540 687292
rect 539516 687292 539528 687306
rect 539764 687306 540764 687312
rect 539764 687292 539776 687306
rect 539516 687272 539776 687292
rect 540752 687292 540764 687306
rect 541000 687306 542000 687312
rect 541000 687292 541012 687306
rect 540752 687272 541012 687292
rect 541988 687292 542000 687306
rect 542236 687306 543236 687312
rect 542236 687292 542248 687306
rect 541988 687272 542248 687292
rect 543224 687292 543236 687306
rect 543472 687306 544472 687312
rect 543472 687292 543484 687306
rect 543224 687272 543484 687292
rect 544460 687292 544472 687306
rect 544708 687306 545708 687312
rect 544708 687292 544720 687306
rect 544460 687272 544720 687292
rect 545696 687292 545708 687306
rect 545944 687306 546944 687312
rect 545944 687292 545956 687306
rect 545696 687272 545956 687292
rect 546932 687292 546944 687306
rect 547180 687306 548180 687312
rect 547180 687292 547192 687306
rect 546932 687272 547192 687292
rect 548168 687292 548180 687306
rect 548416 687306 549416 687312
rect 548416 687292 548428 687306
rect 548168 687272 548428 687292
rect 549404 687292 549416 687306
rect 549652 687306 550652 687312
rect 549652 687292 549664 687306
rect 549404 687272 549664 687292
rect 550640 687292 550652 687306
rect 550640 687272 550669 687292
rect 538519 687242 538849 687272
rect 538839 687202 538849 687242
rect 538929 687242 539059 687272
rect 538929 687202 538939 687242
rect 539049 687202 539059 687242
rect 539139 687242 541329 687272
rect 539139 687202 539149 687242
rect 541319 687202 541329 687242
rect 541409 687242 541549 687272
rect 541409 687202 541419 687242
rect 541539 687202 541549 687242
rect 541629 687242 543859 687272
rect 541629 687202 541639 687242
rect 543849 687202 543859 687242
rect 543939 687242 544039 687272
rect 543939 687202 543949 687242
rect 544029 687202 544039 687242
rect 544119 687242 546319 687272
rect 544119 687202 544129 687242
rect 546309 687192 546319 687242
rect 546399 687242 546499 687272
rect 546399 687192 546409 687242
rect 546489 687192 546499 687242
rect 546579 687242 548799 687272
rect 546579 687192 546589 687242
rect 548789 687192 548799 687242
rect 548879 687242 548969 687272
rect 548879 687192 548889 687242
rect 548959 687192 548969 687242
rect 549049 687242 550669 687272
rect 549049 687192 549059 687242
rect 540107 687142 540221 687148
rect 540107 687062 540119 687142
rect 540209 687062 540221 687142
rect 540107 687056 540221 687062
rect 540287 687142 540401 687148
rect 540287 687062 540299 687142
rect 540389 687062 540401 687142
rect 540287 687056 540401 687062
rect 542637 687142 542751 687148
rect 542637 687062 542649 687142
rect 542739 687062 542751 687142
rect 542637 687056 542751 687062
rect 542797 687142 542911 687148
rect 542797 687062 542809 687142
rect 542899 687062 542911 687142
rect 542797 687056 542911 687062
rect 545107 687142 545221 687148
rect 545107 687062 545119 687142
rect 545209 687062 545221 687142
rect 545107 687056 545221 687062
rect 545267 687142 545381 687148
rect 545267 687062 545279 687142
rect 545369 687062 545381 687142
rect 545267 687056 545381 687062
rect 547557 687142 547671 687148
rect 547557 687062 547569 687142
rect 547659 687062 547671 687142
rect 547557 687056 547671 687062
rect 547717 687142 547831 687148
rect 547717 687062 547729 687142
rect 547819 687062 547831 687142
rect 547717 687056 547831 687062
rect 550057 687142 550171 687148
rect 550057 687062 550069 687142
rect 550159 687062 550171 687142
rect 550057 687056 550171 687062
rect 550217 687142 550331 687148
rect 550217 687062 550229 687142
rect 550319 687062 550331 687142
rect 550217 687056 550331 687062
rect 540089 686962 540099 687022
rect 538519 686942 540099 686962
rect 540179 686962 540189 687022
rect 540319 686962 540329 687022
rect 540179 686942 540329 686962
rect 540409 686962 540419 687022
rect 542639 686962 542649 687012
rect 540409 686942 542649 686962
rect 538519 686932 542649 686942
rect 542729 686962 542739 687012
rect 542809 686962 542819 687022
rect 542729 686942 542819 686962
rect 542899 686962 542909 687022
rect 545099 686962 545109 687022
rect 542899 686942 545109 686962
rect 545189 686962 545199 687022
rect 545289 686962 545299 687022
rect 545189 686942 545299 686962
rect 545379 686962 545389 687022
rect 547549 686962 547559 687012
rect 545379 686942 547559 686962
rect 542729 686932 547559 686942
rect 547639 686962 547649 687012
rect 547739 686962 547749 687012
rect 547639 686932 547749 686962
rect 547829 686962 547839 687012
rect 550059 686962 550069 687012
rect 547829 686932 550069 686962
rect 550149 686962 550159 687012
rect 550229 686962 550239 687012
rect 550149 686932 550239 686962
rect 550319 686962 550329 687012
rect 550319 686932 550669 686962
rect 538519 686924 550669 686932
rect 538519 686912 538540 686924
rect 538528 686890 538540 686912
rect 539516 686912 539776 686924
rect 539516 686890 539528 686912
rect 538528 686884 539528 686890
rect 539764 686890 539776 686912
rect 540752 686912 541012 686924
rect 540752 686890 540764 686912
rect 539764 686884 540764 686890
rect 541000 686890 541012 686912
rect 541988 686912 542248 686924
rect 541988 686890 542000 686912
rect 541000 686884 542000 686890
rect 542236 686890 542248 686912
rect 543224 686912 543484 686924
rect 543224 686890 543236 686912
rect 542236 686884 543236 686890
rect 543472 686890 543484 686912
rect 544460 686912 544720 686924
rect 544460 686890 544472 686912
rect 543472 686884 544472 686890
rect 544708 686890 544720 686912
rect 545696 686912 545956 686924
rect 545696 686890 545708 686912
rect 544708 686884 545708 686890
rect 545944 686890 545956 686912
rect 546932 686912 547192 686924
rect 546932 686890 546944 686912
rect 545944 686884 546944 686890
rect 547180 686890 547192 686912
rect 548168 686912 548428 686924
rect 548168 686890 548180 686912
rect 547180 686884 548180 686890
rect 548416 686890 548428 686912
rect 549404 686912 549664 686924
rect 549404 686890 549416 686912
rect 548416 686884 549416 686890
rect 549652 686890 549664 686912
rect 550640 686912 550669 686924
rect 550640 686890 550652 686912
rect 549652 686884 550652 686890
rect 537568 686874 538479 686882
rect 537568 686862 538487 686874
rect 537568 686841 538447 686862
rect 534609 686497 535039 686829
rect 537039 686794 538447 686841
rect 538481 686852 538487 686862
rect 539569 686872 539615 686874
rect 539677 686872 539723 686874
rect 539569 686862 539579 686872
rect 539709 686862 539723 686872
rect 539569 686852 539575 686862
rect 538481 686812 539575 686852
rect 538481 686794 538487 686812
rect 537039 686782 538487 686794
rect 539569 686794 539575 686812
rect 539717 686852 539723 686862
rect 540805 686862 540851 686874
rect 540913 686862 540959 686874
rect 542041 686862 542087 686874
rect 542149 686862 542195 686874
rect 540805 686852 540811 686862
rect 539717 686812 540811 686852
rect 539609 686794 539615 686802
rect 539569 686782 539615 686794
rect 539677 686794 539683 686802
rect 539717 686794 539723 686812
rect 539677 686782 539723 686794
rect 540805 686794 540811 686812
rect 540953 686852 540959 686862
rect 542039 686852 542047 686862
rect 540953 686812 542047 686852
rect 540953 686794 540959 686812
rect 540805 686792 540819 686794
rect 540949 686792 540959 686794
rect 542039 686794 542047 686812
rect 542189 686852 542195 686862
rect 543277 686862 543323 686874
rect 543385 686862 543431 686874
rect 543277 686852 543283 686862
rect 542189 686812 543283 686852
rect 542189 686794 542195 686812
rect 542039 686792 542049 686794
rect 542179 686792 542195 686794
rect 540805 686782 540851 686792
rect 540913 686782 540959 686792
rect 542041 686782 542087 686792
rect 542149 686782 542195 686792
rect 543277 686794 543283 686812
rect 543425 686852 543431 686862
rect 544513 686862 544559 686874
rect 544621 686862 544667 686874
rect 545749 686862 545795 686874
rect 545857 686862 545903 686874
rect 544513 686852 544519 686862
rect 543425 686812 544519 686852
rect 543425 686794 543431 686812
rect 543277 686792 543289 686794
rect 543419 686792 543431 686794
rect 543277 686782 543323 686792
rect 543385 686782 543431 686792
rect 544513 686794 544519 686812
rect 544661 686852 544669 686862
rect 545749 686852 545755 686862
rect 544661 686812 545755 686852
rect 544661 686794 544669 686812
rect 544513 686792 544529 686794
rect 544659 686792 544669 686794
rect 545749 686794 545755 686812
rect 545897 686852 545903 686862
rect 546985 686862 547031 686874
rect 547093 686862 547139 686874
rect 548221 686862 548267 686874
rect 548329 686862 548375 686874
rect 546985 686852 546991 686862
rect 545897 686812 546991 686852
rect 545897 686794 545903 686812
rect 545749 686792 545759 686794
rect 545889 686792 545903 686794
rect 544513 686782 544559 686792
rect 544621 686782 544667 686792
rect 545749 686782 545795 686792
rect 545857 686782 545903 686792
rect 546985 686794 546991 686812
rect 547133 686852 547139 686862
rect 548219 686852 548227 686862
rect 547133 686812 548227 686852
rect 547133 686794 547139 686812
rect 546985 686792 546999 686794
rect 547129 686792 547139 686794
rect 548219 686794 548227 686812
rect 548369 686852 548375 686862
rect 549457 686862 549503 686874
rect 549565 686862 549611 686874
rect 549457 686852 549463 686862
rect 548369 686812 549463 686852
rect 548369 686794 548375 686812
rect 548219 686792 548229 686794
rect 548359 686792 548375 686794
rect 546985 686782 547031 686792
rect 547093 686782 547139 686792
rect 548221 686782 548267 686792
rect 548329 686782 548375 686792
rect 549457 686794 549463 686812
rect 549605 686852 549611 686862
rect 550693 686872 550739 686874
rect 551669 686872 551800 687322
rect 550693 686862 551800 686872
rect 550693 686852 550699 686862
rect 549605 686812 550699 686852
rect 549605 686794 549611 686812
rect 549457 686792 549469 686794
rect 549599 686792 549611 686794
rect 549457 686782 549503 686792
rect 549565 686782 549611 686792
rect 550693 686794 550699 686812
rect 550733 686841 551800 686862
rect 552197 686841 552203 687955
rect 550733 686829 552203 686841
rect 554109 687955 554634 687967
rect 554109 686841 554231 687955
rect 554628 686841 554634 687955
rect 554109 686829 554634 686841
rect 550733 686794 552099 686829
rect 550693 686782 552099 686794
rect 537039 686772 538479 686782
rect 550699 686772 552099 686782
rect 537039 686497 537469 686772
rect 538528 686766 539528 686772
rect 538528 686752 538540 686766
rect 538519 686732 538540 686752
rect 539516 686752 539528 686766
rect 539764 686766 540764 686772
rect 539764 686752 539776 686766
rect 539516 686732 539776 686752
rect 540752 686752 540764 686766
rect 541000 686766 542000 686772
rect 541000 686752 541012 686766
rect 540752 686732 541012 686752
rect 541988 686752 542000 686766
rect 542236 686766 543236 686772
rect 542236 686752 542248 686766
rect 541988 686732 542248 686752
rect 543224 686752 543236 686766
rect 543472 686766 544472 686772
rect 543472 686752 543484 686766
rect 543224 686732 543484 686752
rect 544460 686752 544472 686766
rect 544708 686766 545708 686772
rect 544708 686752 544720 686766
rect 544460 686732 544720 686752
rect 545696 686752 545708 686766
rect 545944 686766 546944 686772
rect 545944 686752 545956 686766
rect 545696 686732 545956 686752
rect 546932 686752 546944 686766
rect 547180 686766 548180 686772
rect 547180 686752 547192 686766
rect 546932 686732 547192 686752
rect 548168 686752 548180 686766
rect 548416 686766 549416 686772
rect 548416 686752 548428 686766
rect 548168 686732 548428 686752
rect 549404 686752 549416 686766
rect 549652 686766 550652 686772
rect 549652 686752 549664 686766
rect 549404 686732 549664 686752
rect 550640 686752 550652 686766
rect 550640 686732 550669 686752
rect 538519 686702 538849 686732
rect 538839 686662 538849 686702
rect 538929 686702 539059 686732
rect 538929 686662 538939 686702
rect 539049 686662 539059 686702
rect 539139 686702 541329 686732
rect 539139 686662 539149 686702
rect 541319 686662 541329 686702
rect 541409 686702 541549 686732
rect 541409 686662 541419 686702
rect 541539 686662 541549 686702
rect 541629 686702 543859 686732
rect 541629 686662 541639 686702
rect 543849 686662 543859 686702
rect 543939 686702 544049 686732
rect 543939 686662 543949 686702
rect 544039 686662 544049 686702
rect 544129 686702 546319 686732
rect 544129 686662 544139 686702
rect 546309 686652 546319 686702
rect 546399 686702 546499 686732
rect 546399 686652 546409 686702
rect 546489 686652 546499 686702
rect 546579 686702 548799 686732
rect 546579 686652 546589 686702
rect 548789 686652 548799 686702
rect 548879 686702 548969 686732
rect 548879 686652 548889 686702
rect 548959 686652 548969 686702
rect 549049 686702 550669 686732
rect 549049 686652 549059 686702
rect 551669 686497 552099 686772
rect 554109 686497 554539 686829
rect 534609 686485 535143 686497
rect 42250 686350 42260 686380
rect 42240 686300 42260 686350
rect 42250 686270 42260 686300
rect 42370 686350 42380 686380
rect 42500 686350 42510 686380
rect 42370 686300 42510 686350
rect 42370 686270 42380 686300
rect 42500 686270 42510 686300
rect 42620 686350 42630 686380
rect 46650 686350 46660 686380
rect 42620 686342 46660 686350
rect 42620 686308 43152 686342
rect 43320 686308 43410 686342
rect 43578 686308 43668 686342
rect 43836 686308 43926 686342
rect 44094 686308 44184 686342
rect 44352 686308 44442 686342
rect 44610 686308 44700 686342
rect 44868 686308 44958 686342
rect 45126 686308 45216 686342
rect 45384 686308 45474 686342
rect 45642 686308 45732 686342
rect 45900 686308 45990 686342
rect 46158 686308 46660 686342
rect 42620 686300 46660 686308
rect 42620 686270 42630 686300
rect 46650 686270 46660 686300
rect 46770 686350 46780 686380
rect 46900 686350 46910 686380
rect 46770 686300 46910 686350
rect 46770 686270 46780 686300
rect 46900 686270 46910 686300
rect 47020 686350 47030 686380
rect 47020 686300 47040 686350
rect 47020 686270 47030 686300
rect 44520 686246 44530 686250
rect 43821 686240 44530 686246
rect 44780 686246 44790 686250
rect 44780 686240 45489 686246
rect 43821 686206 43833 686240
rect 45477 686206 45489 686240
rect 43821 686200 44530 686206
rect 44520 686040 44530 686200
rect 43690 686034 44530 686040
rect 44780 686200 45489 686206
rect 44780 686040 44790 686200
rect 44780 686034 45616 686040
rect 43690 686000 43702 686034
rect 45604 686000 45616 686034
rect 43690 685994 45616 686000
rect 44520 685990 44790 685994
rect 42250 685940 42260 685970
rect 42240 685890 42260 685940
rect 42250 685860 42260 685890
rect 42370 685940 42380 685970
rect 42500 685940 42510 685970
rect 42370 685890 42510 685940
rect 42370 685860 42380 685890
rect 42500 685860 42510 685890
rect 42620 685940 42630 685970
rect 46650 685940 46660 685970
rect 42620 685932 46660 685940
rect 42620 685898 42892 685932
rect 43060 685898 43150 685932
rect 43318 685898 43408 685932
rect 43576 685898 43666 685932
rect 43834 685898 43924 685932
rect 44092 685898 44182 685932
rect 44350 685898 44440 685932
rect 44608 685898 44698 685932
rect 44866 685898 44956 685932
rect 45124 685898 45214 685932
rect 45382 685898 45472 685932
rect 45640 685898 45730 685932
rect 45898 685898 45988 685932
rect 46156 685898 46246 685932
rect 46414 685898 46660 685932
rect 42620 685890 46660 685898
rect 42620 685860 42630 685890
rect 46650 685860 46660 685890
rect 46770 685940 46780 685970
rect 46900 685940 46910 685970
rect 46770 685890 46910 685940
rect 46770 685860 46780 685890
rect 46900 685860 46910 685890
rect 47020 685940 47030 685970
rect 47020 685890 47040 685940
rect 47020 685860 47030 685890
rect 42824 685848 42870 685860
rect 42824 685820 42830 685848
rect 42864 685820 42870 685848
rect 43082 685848 43128 685860
rect 42800 685750 42810 685820
rect 42880 685750 42890 685820
rect 42824 685640 42830 685750
rect 42864 685640 42870 685750
rect 42800 685570 42810 685640
rect 42880 685570 42890 685640
rect 42824 684872 42830 685570
rect 42864 684872 42870 685570
rect 43082 685150 43088 685848
rect 43122 685150 43128 685848
rect 43340 685848 43386 685860
rect 43340 685820 43346 685848
rect 43380 685820 43386 685848
rect 43598 685848 43644 685860
rect 43320 685750 43330 685820
rect 43400 685750 43410 685820
rect 43340 685640 43346 685750
rect 43380 685640 43386 685750
rect 43320 685570 43330 685640
rect 43400 685570 43410 685640
rect 43060 685080 43070 685150
rect 43140 685080 43150 685150
rect 43082 684970 43088 685080
rect 43122 684970 43128 685080
rect 43060 684900 43070 684970
rect 43140 684900 43150 684970
rect 42824 684860 42870 684872
rect 43082 684872 43088 684900
rect 43122 684872 43128 684900
rect 43082 684860 43128 684872
rect 43340 684872 43346 685570
rect 43380 684872 43386 685570
rect 43598 685150 43604 685848
rect 43638 685150 43644 685848
rect 43856 685848 43902 685860
rect 43856 685820 43862 685848
rect 43896 685820 43902 685848
rect 44114 685848 44160 685860
rect 43830 685750 43840 685820
rect 43910 685750 43920 685820
rect 43856 685640 43862 685750
rect 43896 685640 43902 685750
rect 43830 685570 43840 685640
rect 43910 685570 43920 685640
rect 43570 685080 43580 685150
rect 43650 685080 43660 685150
rect 43598 684970 43604 685080
rect 43638 684970 43644 685080
rect 43570 684900 43580 684970
rect 43650 684900 43660 684970
rect 43340 684860 43386 684872
rect 43598 684872 43604 684900
rect 43638 684872 43644 684900
rect 43598 684860 43644 684872
rect 43856 684872 43862 685570
rect 43896 684872 43902 685570
rect 44114 685150 44120 685848
rect 44154 685150 44160 685848
rect 44372 685848 44418 685860
rect 44372 685820 44378 685848
rect 44412 685820 44418 685848
rect 44630 685848 44676 685860
rect 44350 685750 44360 685820
rect 44430 685750 44440 685820
rect 44372 685640 44378 685750
rect 44412 685640 44418 685750
rect 44350 685570 44360 685640
rect 44430 685570 44440 685640
rect 44090 685080 44100 685150
rect 44170 685080 44180 685150
rect 44114 684970 44120 685080
rect 44154 684970 44160 685080
rect 44090 684900 44100 684970
rect 44170 684900 44180 684970
rect 43856 684860 43902 684872
rect 44114 684872 44120 684900
rect 44154 684872 44160 684900
rect 44114 684860 44160 684872
rect 44372 684872 44378 685570
rect 44412 684872 44418 685570
rect 44630 685150 44636 685848
rect 44670 685150 44676 685848
rect 44888 685848 44934 685860
rect 44888 685820 44894 685848
rect 44928 685820 44934 685848
rect 45146 685848 45192 685860
rect 44860 685750 44870 685820
rect 44940 685750 44950 685820
rect 44888 685640 44894 685750
rect 44928 685640 44934 685750
rect 44860 685570 44870 685640
rect 44940 685570 44950 685640
rect 44610 685080 44620 685150
rect 44690 685080 44700 685150
rect 44630 684970 44636 685080
rect 44670 684970 44676 685080
rect 44610 684900 44620 684970
rect 44690 684900 44700 684970
rect 44372 684860 44418 684872
rect 44630 684872 44636 684900
rect 44670 684872 44676 684900
rect 44630 684860 44676 684872
rect 44888 684872 44894 685570
rect 44928 684872 44934 685570
rect 45146 685150 45152 685848
rect 45186 685150 45192 685848
rect 45404 685848 45450 685860
rect 45404 685820 45410 685848
rect 45444 685820 45450 685848
rect 45662 685848 45708 685860
rect 45380 685750 45390 685820
rect 45460 685750 45470 685820
rect 45404 685640 45410 685750
rect 45444 685640 45450 685750
rect 45380 685570 45390 685640
rect 45460 685570 45470 685640
rect 45120 685080 45130 685150
rect 45200 685080 45210 685150
rect 45146 684970 45152 685080
rect 45186 684970 45192 685080
rect 45120 684900 45130 684970
rect 45200 684900 45210 684970
rect 44888 684860 44934 684872
rect 45146 684872 45152 684900
rect 45186 684872 45192 684900
rect 45146 684860 45192 684872
rect 45404 684872 45410 685570
rect 45444 684872 45450 685570
rect 45662 685150 45668 685848
rect 45702 685150 45708 685848
rect 45920 685848 45966 685860
rect 45920 685820 45926 685848
rect 45960 685820 45966 685848
rect 46178 685848 46224 685860
rect 45900 685750 45910 685820
rect 45980 685750 45990 685820
rect 45920 685640 45926 685750
rect 45960 685640 45966 685750
rect 45900 685570 45910 685640
rect 45980 685570 45990 685640
rect 45640 685080 45650 685150
rect 45720 685080 45730 685150
rect 45662 684970 45668 685080
rect 45702 684970 45708 685080
rect 45640 684900 45650 684970
rect 45720 684900 45730 684970
rect 45404 684860 45450 684872
rect 45662 684872 45668 684900
rect 45702 684872 45708 684900
rect 45662 684860 45708 684872
rect 45920 684872 45926 685570
rect 45960 684872 45966 685570
rect 46178 685150 46184 685848
rect 46218 685150 46224 685848
rect 46436 685848 46482 685860
rect 46436 685820 46442 685848
rect 46476 685820 46482 685848
rect 46410 685750 46420 685820
rect 46490 685750 46500 685820
rect 46436 685640 46442 685750
rect 46476 685640 46482 685750
rect 46410 685570 46420 685640
rect 46490 685570 46500 685640
rect 46150 685080 46160 685150
rect 46230 685080 46240 685150
rect 46178 684970 46184 685080
rect 46218 684970 46224 685080
rect 46150 684900 46160 684970
rect 46230 684900 46240 684970
rect 45920 684860 45966 684872
rect 46178 684872 46184 684900
rect 46218 684872 46224 684900
rect 46178 684860 46224 684872
rect 46436 684872 46442 685570
rect 46476 684872 46482 685570
rect 534609 685392 534740 686485
rect 534734 685371 534740 685392
rect 535137 685371 535143 686485
rect 537039 686485 537574 686497
rect 537039 685382 537171 686485
rect 534734 685359 535143 685371
rect 537165 685371 537171 685382
rect 537568 686342 537574 686485
rect 551669 686485 552203 686497
rect 540089 686422 540099 686482
rect 538519 686402 540099 686422
rect 540179 686422 540189 686482
rect 540319 686422 540329 686482
rect 540179 686402 540329 686422
rect 540409 686422 540419 686482
rect 542629 686422 542639 686472
rect 540409 686402 542639 686422
rect 538519 686392 542639 686402
rect 542719 686422 542729 686472
rect 542799 686422 542809 686472
rect 542719 686392 542809 686422
rect 542889 686422 542899 686472
rect 545099 686422 545109 686472
rect 542889 686392 545109 686422
rect 545189 686422 545199 686472
rect 545279 686422 545289 686472
rect 545189 686392 545289 686422
rect 545369 686422 545379 686472
rect 547549 686422 547559 686472
rect 545369 686392 547559 686422
rect 547639 686422 547649 686472
rect 547739 686422 547749 686472
rect 547639 686392 547749 686422
rect 547829 686422 547839 686472
rect 550059 686422 550069 686472
rect 547829 686392 550069 686422
rect 550149 686422 550159 686472
rect 550229 686422 550239 686472
rect 550149 686392 550239 686422
rect 550319 686422 550329 686472
rect 550319 686392 550669 686422
rect 538519 686384 550669 686392
rect 538519 686372 538540 686384
rect 538528 686350 538540 686372
rect 539516 686372 539776 686384
rect 539516 686350 539528 686372
rect 538528 686344 539528 686350
rect 539764 686350 539776 686372
rect 540752 686372 541012 686384
rect 540752 686350 540764 686372
rect 539764 686344 540764 686350
rect 541000 686350 541012 686372
rect 541988 686372 542248 686384
rect 541988 686350 542000 686372
rect 541000 686344 542000 686350
rect 542236 686350 542248 686372
rect 543224 686372 543484 686384
rect 543224 686350 543236 686372
rect 542236 686344 543236 686350
rect 543472 686350 543484 686372
rect 544460 686372 544720 686384
rect 544460 686350 544472 686372
rect 543472 686344 544472 686350
rect 544708 686350 544720 686372
rect 545696 686372 545956 686384
rect 545696 686350 545708 686372
rect 544708 686344 545708 686350
rect 545944 686350 545956 686372
rect 546932 686372 547192 686384
rect 546932 686350 546944 686372
rect 545944 686344 546944 686350
rect 547180 686350 547192 686372
rect 548168 686372 548428 686384
rect 548168 686350 548180 686372
rect 547180 686344 548180 686350
rect 548416 686350 548428 686372
rect 549404 686372 549664 686384
rect 549404 686350 549416 686372
rect 548416 686344 549416 686350
rect 549652 686350 549664 686372
rect 550640 686372 550669 686384
rect 550640 686350 550652 686372
rect 549652 686344 550652 686350
rect 551669 686342 551800 686485
rect 537568 686322 538499 686342
rect 550699 686334 551800 686342
rect 537568 686254 538447 686322
rect 538481 686312 538499 686322
rect 539569 686322 539615 686334
rect 539677 686322 539723 686334
rect 539569 686312 539575 686322
rect 538481 686272 539575 686312
rect 538481 686254 538499 686272
rect 537568 686232 538499 686254
rect 539569 686254 539575 686272
rect 539717 686312 539723 686322
rect 540805 686322 540851 686334
rect 540913 686322 540959 686334
rect 542041 686322 542087 686334
rect 542149 686322 542195 686334
rect 540805 686312 540811 686322
rect 539717 686272 540811 686312
rect 539717 686254 539723 686272
rect 539569 686252 539579 686254
rect 539709 686252 539723 686254
rect 539569 686242 539615 686252
rect 539677 686242 539723 686252
rect 540805 686254 540811 686272
rect 540953 686312 540959 686322
rect 542039 686312 542047 686322
rect 540953 686272 542047 686312
rect 540953 686254 540959 686272
rect 540805 686252 540819 686254
rect 540949 686252 540959 686254
rect 542039 686254 542047 686272
rect 542189 686312 542195 686322
rect 543277 686322 543323 686334
rect 543385 686322 543431 686334
rect 543277 686312 543283 686322
rect 542189 686272 543283 686312
rect 542189 686254 542195 686272
rect 542039 686252 542049 686254
rect 542179 686252 542195 686254
rect 540805 686242 540851 686252
rect 540913 686242 540959 686252
rect 542041 686242 542087 686252
rect 542149 686242 542195 686252
rect 543277 686254 543283 686272
rect 543425 686312 543431 686322
rect 544513 686322 544559 686334
rect 544621 686322 544667 686334
rect 545749 686322 545795 686334
rect 545857 686322 545903 686334
rect 544513 686312 544519 686322
rect 543425 686272 544519 686312
rect 543425 686254 543431 686272
rect 543277 686252 543289 686254
rect 543419 686252 543431 686254
rect 543277 686242 543323 686252
rect 543385 686242 543431 686252
rect 544513 686254 544519 686272
rect 544661 686312 544669 686322
rect 545749 686312 545755 686322
rect 544661 686272 545755 686312
rect 544661 686254 544669 686272
rect 544513 686252 544529 686254
rect 544659 686252 544669 686254
rect 545749 686254 545755 686272
rect 545897 686312 545903 686322
rect 546985 686322 547031 686334
rect 547093 686322 547139 686334
rect 548221 686322 548267 686334
rect 548329 686322 548375 686334
rect 546985 686312 546991 686322
rect 545897 686272 546991 686312
rect 545897 686254 545903 686272
rect 545749 686252 545759 686254
rect 545889 686252 545903 686254
rect 544513 686242 544559 686252
rect 544621 686242 544667 686252
rect 545749 686242 545795 686252
rect 545857 686242 545903 686252
rect 546985 686254 546991 686272
rect 547133 686312 547139 686322
rect 548219 686312 548227 686322
rect 547133 686272 548227 686312
rect 547133 686254 547139 686272
rect 546985 686252 546999 686254
rect 547129 686252 547139 686254
rect 548219 686254 548227 686272
rect 548369 686312 548375 686322
rect 549457 686322 549503 686334
rect 549565 686322 549611 686334
rect 549457 686312 549463 686322
rect 548369 686272 549463 686312
rect 548369 686254 548375 686272
rect 548219 686252 548229 686254
rect 548359 686252 548375 686254
rect 546985 686242 547031 686252
rect 547093 686242 547139 686252
rect 548221 686242 548267 686252
rect 548329 686242 548375 686252
rect 549457 686254 549463 686272
rect 549605 686312 549611 686322
rect 550693 686322 551800 686334
rect 550693 686312 550699 686322
rect 549605 686272 550699 686312
rect 549605 686254 549611 686272
rect 549457 686252 549469 686254
rect 549599 686252 549611 686254
rect 549457 686242 549503 686252
rect 549565 686242 549611 686252
rect 550693 686254 550699 686272
rect 550733 686254 551800 686322
rect 550693 686242 551800 686254
rect 537568 685802 537574 686232
rect 538528 686226 539528 686232
rect 538528 686212 538540 686226
rect 538519 686192 538540 686212
rect 539516 686212 539528 686226
rect 539764 686226 540764 686232
rect 539764 686212 539776 686226
rect 539516 686192 539776 686212
rect 540752 686212 540764 686226
rect 541000 686226 542000 686232
rect 541000 686212 541012 686226
rect 540752 686192 541012 686212
rect 541988 686212 542000 686226
rect 542236 686226 543236 686232
rect 542236 686212 542248 686226
rect 541988 686192 542248 686212
rect 543224 686212 543236 686226
rect 543472 686226 544472 686232
rect 543472 686212 543484 686226
rect 543224 686192 543484 686212
rect 544460 686212 544472 686226
rect 544708 686226 545708 686232
rect 544708 686212 544720 686226
rect 544460 686192 544720 686212
rect 545696 686212 545708 686226
rect 545944 686226 546944 686232
rect 545944 686212 545956 686226
rect 545696 686192 545956 686212
rect 546932 686212 546944 686226
rect 547180 686226 548180 686232
rect 547180 686212 547192 686226
rect 546932 686192 547192 686212
rect 548168 686212 548180 686226
rect 548416 686226 549416 686232
rect 548416 686212 548428 686226
rect 548168 686192 548428 686212
rect 549404 686212 549416 686226
rect 549652 686226 550652 686232
rect 549652 686212 549664 686226
rect 549404 686192 549664 686212
rect 550640 686212 550652 686226
rect 550640 686192 550669 686212
rect 538519 686162 538849 686192
rect 538839 686122 538849 686162
rect 538929 686162 539059 686192
rect 538929 686122 538939 686162
rect 539049 686122 539059 686162
rect 539139 686162 541319 686192
rect 539139 686122 539149 686162
rect 541309 686122 541319 686162
rect 541399 686162 541559 686192
rect 541399 686122 541409 686162
rect 541549 686122 541559 686162
rect 541639 686162 543859 686192
rect 541639 686122 541649 686162
rect 543849 686122 543859 686162
rect 543939 686162 544039 686192
rect 543939 686122 543949 686162
rect 544029 686122 544039 686162
rect 544119 686162 546329 686192
rect 544119 686122 544129 686162
rect 546319 686112 546329 686162
rect 546409 686162 546499 686192
rect 546409 686112 546419 686162
rect 546489 686112 546499 686162
rect 546579 686162 548799 686192
rect 546579 686112 546589 686162
rect 548789 686112 548799 686162
rect 548879 686162 548969 686192
rect 548879 686112 548889 686162
rect 548959 686112 548969 686162
rect 549049 686162 550669 686192
rect 549049 686112 549059 686162
rect 540287 686072 540401 686078
rect 540107 686062 540221 686068
rect 540107 685982 540119 686062
rect 540209 685982 540221 686062
rect 540287 685992 540299 686072
rect 540389 685992 540401 686072
rect 540287 685986 540401 685992
rect 542637 686062 542751 686068
rect 540107 685976 540221 685982
rect 542637 685982 542649 686062
rect 542739 685982 542751 686062
rect 542637 685976 542751 685982
rect 542797 686062 542911 686068
rect 542797 685982 542809 686062
rect 542899 685982 542911 686062
rect 542797 685976 542911 685982
rect 545107 686062 545221 686068
rect 545107 685982 545119 686062
rect 545209 685982 545221 686062
rect 545107 685976 545221 685982
rect 545267 686062 545381 686068
rect 545267 685982 545279 686062
rect 545369 685982 545381 686062
rect 545267 685976 545381 685982
rect 547557 686062 547671 686068
rect 547557 685982 547569 686062
rect 547659 685982 547671 686062
rect 547557 685976 547671 685982
rect 547717 686062 547831 686068
rect 547717 685982 547729 686062
rect 547819 685982 547831 686062
rect 547717 685976 547831 685982
rect 550057 686062 550171 686068
rect 550057 685982 550069 686062
rect 550159 685982 550171 686062
rect 550057 685976 550171 685982
rect 550217 686062 550331 686068
rect 550217 685982 550229 686062
rect 550319 685982 550331 686062
rect 550217 685976 550331 685982
rect 540089 685882 540099 685932
rect 538519 685852 540099 685882
rect 540179 685882 540189 685932
rect 540319 685882 540329 685932
rect 540179 685852 540329 685882
rect 540409 685882 540419 685932
rect 542619 685882 542629 685942
rect 540409 685862 542629 685882
rect 542709 685882 542719 685942
rect 542809 685882 542819 685942
rect 542709 685862 542819 685882
rect 542899 685882 542909 685942
rect 545099 685882 545109 685932
rect 542899 685862 545109 685882
rect 540409 685852 545109 685862
rect 545189 685882 545199 685932
rect 545289 685882 545299 685932
rect 545189 685852 545299 685882
rect 545379 685882 545389 685932
rect 547549 685882 547559 685932
rect 545379 685852 547559 685882
rect 547639 685882 547649 685932
rect 547739 685882 547749 685932
rect 547639 685852 547749 685882
rect 547829 685882 547839 685932
rect 550059 685882 550069 685922
rect 547829 685852 550069 685882
rect 538519 685844 550069 685852
rect 550149 685882 550159 685922
rect 550229 685882 550239 685922
rect 550149 685844 550239 685882
rect 550319 685882 550329 685922
rect 550319 685844 550669 685882
rect 538519 685832 538540 685844
rect 538528 685810 538540 685832
rect 539516 685832 539776 685844
rect 539516 685810 539528 685832
rect 538528 685804 539528 685810
rect 539764 685810 539776 685832
rect 540752 685832 541012 685844
rect 540752 685810 540764 685832
rect 539764 685804 540764 685810
rect 541000 685810 541012 685832
rect 541988 685832 542248 685844
rect 541988 685810 542000 685832
rect 541000 685804 542000 685810
rect 542236 685810 542248 685832
rect 543224 685832 543484 685844
rect 543224 685810 543236 685832
rect 542236 685804 543236 685810
rect 543472 685810 543484 685832
rect 544460 685832 544720 685844
rect 544460 685810 544472 685832
rect 543472 685804 544472 685810
rect 544708 685810 544720 685832
rect 545696 685832 545956 685844
rect 545696 685810 545708 685832
rect 544708 685804 545708 685810
rect 545944 685810 545956 685832
rect 546932 685832 547192 685844
rect 546932 685810 546944 685832
rect 545944 685804 546944 685810
rect 547180 685810 547192 685832
rect 548168 685832 548428 685844
rect 548168 685810 548180 685832
rect 547180 685804 548180 685810
rect 548416 685810 548428 685832
rect 549404 685832 549664 685844
rect 549404 685810 549416 685832
rect 548416 685804 549416 685810
rect 549652 685810 549664 685832
rect 550640 685832 550669 685844
rect 550640 685810 550652 685832
rect 549652 685804 550652 685810
rect 551669 685802 551800 686242
rect 537568 685782 538489 685802
rect 550699 685794 551800 685802
rect 537568 685714 538447 685782
rect 538481 685772 538489 685782
rect 539569 685782 539615 685794
rect 539677 685782 539723 685794
rect 539569 685772 539575 685782
rect 538481 685732 539575 685772
rect 538481 685714 538489 685732
rect 537568 685692 538489 685714
rect 539569 685714 539575 685732
rect 539717 685772 539723 685782
rect 540805 685782 540851 685794
rect 540913 685782 540959 685794
rect 542041 685782 542087 685794
rect 542149 685782 542195 685794
rect 540805 685772 540811 685782
rect 539717 685732 540811 685772
rect 539717 685714 539723 685732
rect 539569 685712 539579 685714
rect 539709 685712 539723 685714
rect 539569 685702 539615 685712
rect 539677 685702 539723 685712
rect 540805 685714 540811 685732
rect 540953 685772 540959 685782
rect 542039 685772 542047 685782
rect 540953 685732 542047 685772
rect 540953 685714 540959 685732
rect 540805 685712 540819 685714
rect 540949 685712 540959 685714
rect 542039 685714 542047 685732
rect 542189 685772 542195 685782
rect 543277 685782 543323 685794
rect 543385 685782 543431 685794
rect 543277 685772 543283 685782
rect 542189 685732 543283 685772
rect 542189 685714 542195 685732
rect 542039 685712 542049 685714
rect 542179 685712 542195 685714
rect 540805 685702 540851 685712
rect 540913 685702 540959 685712
rect 542041 685702 542087 685712
rect 542149 685702 542195 685712
rect 543277 685714 543283 685732
rect 543425 685772 543431 685782
rect 544513 685782 544559 685794
rect 544621 685782 544667 685794
rect 545749 685782 545795 685794
rect 545857 685782 545903 685794
rect 544513 685772 544519 685782
rect 543425 685732 544519 685772
rect 543425 685714 543431 685732
rect 543277 685712 543289 685714
rect 543419 685712 543431 685714
rect 543277 685702 543323 685712
rect 543385 685702 543431 685712
rect 544513 685714 544519 685732
rect 544661 685772 544669 685782
rect 545749 685772 545755 685782
rect 544661 685732 545755 685772
rect 544661 685714 544669 685732
rect 544513 685712 544529 685714
rect 544659 685712 544669 685714
rect 545749 685714 545755 685732
rect 545897 685772 545903 685782
rect 546985 685782 547031 685794
rect 547093 685782 547139 685794
rect 548221 685782 548267 685794
rect 548329 685782 548375 685794
rect 546985 685772 546991 685782
rect 545897 685732 546991 685772
rect 545897 685714 545903 685732
rect 545749 685712 545759 685714
rect 545889 685712 545903 685714
rect 544513 685702 544559 685712
rect 544621 685702 544667 685712
rect 545749 685702 545795 685712
rect 545857 685702 545903 685712
rect 546985 685714 546991 685732
rect 547133 685772 547139 685782
rect 548219 685772 548227 685782
rect 547133 685732 548227 685772
rect 547133 685714 547139 685732
rect 546985 685712 546999 685714
rect 547129 685712 547139 685714
rect 548219 685714 548227 685732
rect 548369 685772 548375 685782
rect 549457 685782 549503 685794
rect 549565 685782 549611 685794
rect 549457 685772 549463 685782
rect 548369 685732 549463 685772
rect 548369 685714 548375 685732
rect 548219 685712 548229 685714
rect 548359 685712 548375 685714
rect 546985 685702 547031 685712
rect 547093 685702 547139 685712
rect 548221 685702 548267 685712
rect 548329 685702 548375 685712
rect 549457 685714 549463 685732
rect 549605 685772 549611 685782
rect 550693 685782 551800 685794
rect 550693 685772 550699 685782
rect 549605 685732 550699 685772
rect 549605 685714 549611 685732
rect 549457 685712 549469 685714
rect 549599 685712 549611 685714
rect 549457 685702 549503 685712
rect 549565 685702 549611 685712
rect 550693 685714 550699 685732
rect 550733 685714 551800 685782
rect 550693 685702 551800 685714
rect 537568 685371 537574 685692
rect 538528 685686 539528 685692
rect 538528 685672 538540 685686
rect 538519 685652 538540 685672
rect 539516 685672 539528 685686
rect 539764 685686 540764 685692
rect 539764 685672 539776 685686
rect 539516 685652 539776 685672
rect 540752 685672 540764 685686
rect 541000 685686 542000 685692
rect 541000 685672 541012 685686
rect 540752 685652 541012 685672
rect 541988 685672 542000 685686
rect 542236 685686 543236 685692
rect 542236 685672 542248 685686
rect 541988 685652 542248 685672
rect 543224 685672 543236 685686
rect 543472 685686 544472 685692
rect 543472 685672 543484 685686
rect 543224 685652 543484 685672
rect 544460 685672 544472 685686
rect 544708 685686 545708 685692
rect 544708 685672 544720 685686
rect 544460 685652 544720 685672
rect 545696 685672 545708 685686
rect 545944 685686 546944 685692
rect 545944 685672 545956 685686
rect 545696 685652 545956 685672
rect 546932 685672 546944 685686
rect 547180 685686 548180 685692
rect 547180 685672 547192 685686
rect 546932 685652 547192 685672
rect 548168 685672 548180 685686
rect 548416 685686 549416 685692
rect 548416 685672 548428 685686
rect 548168 685652 548428 685672
rect 549404 685672 549416 685686
rect 549652 685686 550652 685692
rect 549652 685672 549664 685686
rect 549404 685652 549664 685672
rect 550640 685672 550652 685686
rect 550640 685652 550669 685672
rect 538519 685622 538849 685652
rect 538839 685582 538849 685622
rect 538929 685622 539059 685652
rect 538929 685582 538939 685622
rect 539049 685582 539059 685622
rect 539139 685622 541319 685652
rect 539139 685582 539149 685622
rect 541309 685572 541319 685622
rect 541399 685622 541559 685652
rect 541399 685572 541409 685622
rect 541549 685572 541559 685622
rect 541639 685622 543859 685652
rect 541639 685572 541649 685622
rect 543849 685582 543859 685622
rect 543939 685622 544049 685652
rect 543939 685582 543949 685622
rect 544039 685582 544049 685622
rect 544129 685622 546319 685652
rect 544129 685582 544139 685622
rect 546309 685572 546319 685622
rect 546399 685622 546509 685652
rect 546399 685572 546409 685622
rect 546499 685572 546509 685622
rect 546589 685642 550669 685652
rect 546589 685622 548799 685642
rect 546589 685572 546599 685622
rect 548789 685562 548799 685622
rect 548879 685622 548969 685642
rect 548879 685562 548889 685622
rect 548959 685562 548969 685622
rect 549049 685622 550669 685642
rect 549049 685562 549059 685622
rect 551669 685382 551800 685702
rect 537165 685359 537574 685371
rect 551794 685371 551800 685382
rect 552197 685371 552203 686485
rect 551794 685359 552203 685371
rect 554109 686485 554634 686497
rect 554109 685371 554231 686485
rect 554628 685371 554634 686485
rect 554109 685362 554634 685371
rect 554225 685359 554634 685362
rect 535753 685252 535855 685264
rect 535963 685252 536065 685264
rect 535749 685122 535759 685252
rect 535849 685122 535859 685252
rect 535959 685122 535969 685252
rect 536059 685122 536069 685252
rect 553063 685242 553145 685254
rect 553223 685242 553305 685254
rect 553059 685152 553069 685242
rect 553139 685152 553149 685242
rect 553219 685152 553229 685242
rect 553299 685152 553309 685242
rect 542359 685132 542589 685142
rect 535753 685110 535855 685122
rect 535963 685110 536065 685122
rect 540809 685082 540819 685132
rect 540449 685064 540819 685082
rect 540949 685082 540959 685132
rect 542129 685122 542229 685132
rect 542039 685082 542049 685122
rect 540949 685064 542049 685082
rect 542179 685082 542229 685122
rect 542359 685082 542379 685132
rect 542179 685064 542379 685082
rect 542459 685064 542489 685132
rect 542569 685082 542589 685132
rect 544549 685122 544649 685152
rect 544769 685132 544999 685152
rect 547229 685142 547459 685152
rect 543279 685082 543289 685122
rect 542569 685064 543289 685082
rect 543419 685082 543429 685122
rect 544519 685082 544529 685122
rect 543419 685064 544529 685082
rect 544659 685082 544669 685122
rect 544769 685082 544789 685132
rect 544659 685064 544789 685082
rect 544869 685064 544899 685132
rect 544979 685082 544999 685132
rect 545749 685082 545759 685122
rect 544979 685064 545759 685082
rect 545889 685082 545899 685122
rect 546979 685082 546999 685142
rect 545889 685072 546999 685082
rect 547129 685082 547139 685142
rect 547229 685082 547249 685142
rect 547129 685072 547249 685082
rect 545889 685064 547249 685072
rect 547329 685064 547359 685142
rect 547439 685082 547459 685142
rect 553063 685140 553145 685152
rect 553223 685140 553305 685152
rect 548219 685082 548229 685122
rect 547439 685064 548229 685082
rect 548359 685082 548369 685122
rect 548359 685064 548779 685082
rect 566260 685080 571820 689300
rect 540449 685042 540471 685064
rect 540459 685030 540471 685042
rect 541447 685042 541689 685064
rect 541447 685030 541459 685042
rect 540459 685024 541459 685030
rect 541677 685030 541689 685042
rect 542665 685042 542907 685064
rect 542665 685030 542677 685042
rect 541677 685024 542677 685030
rect 542895 685030 542907 685042
rect 543883 685042 544125 685064
rect 543883 685030 543895 685042
rect 542895 685024 543895 685030
rect 544113 685030 544125 685042
rect 545101 685042 545343 685064
rect 545101 685030 545113 685042
rect 544113 685024 545113 685030
rect 545331 685030 545343 685042
rect 546319 685042 546561 685064
rect 546319 685030 546331 685042
rect 545331 685024 546331 685030
rect 546549 685030 546561 685042
rect 547537 685042 547779 685064
rect 547537 685030 547549 685042
rect 546549 685024 547549 685030
rect 547767 685030 547779 685042
rect 548755 685042 548779 685064
rect 548755 685030 548767 685042
rect 547767 685024 548767 685030
rect 548820 685014 571820 685080
rect 540381 685002 540427 685014
rect 540381 684992 540387 685002
rect 540379 684952 540387 684992
rect 540381 684934 540387 684952
rect 540421 684992 540427 685002
rect 541491 685002 541537 685014
rect 541491 684992 541497 685002
rect 540421 684952 541497 684992
rect 540421 684934 540427 684952
rect 540381 684922 540427 684934
rect 541491 684934 541497 684952
rect 541531 684992 541537 685002
rect 541599 685002 541645 685014
rect 541599 684992 541605 685002
rect 541531 684952 541605 684992
rect 541531 684934 541537 684952
rect 541491 684922 541537 684934
rect 541599 684934 541605 684952
rect 541639 684992 541645 685002
rect 542709 685002 542755 685014
rect 542817 685002 542863 685014
rect 542709 684992 542715 685002
rect 541639 684952 542715 684992
rect 541639 684934 541645 684952
rect 541599 684922 541645 684934
rect 542709 684934 542715 684952
rect 542749 684934 542823 685002
rect 542857 684992 542863 685002
rect 543927 685002 543973 685014
rect 544035 685002 544081 685014
rect 543927 684992 543933 685002
rect 542857 684952 543933 684992
rect 542857 684934 542863 684952
rect 542709 684932 542863 684934
rect 542709 684922 542755 684932
rect 542817 684922 542863 684932
rect 543927 684934 543933 684952
rect 543967 684934 544041 685002
rect 544075 684992 544081 685002
rect 545145 685002 545191 685014
rect 545253 685002 545299 685014
rect 545145 684992 545151 685002
rect 544075 684952 545151 684992
rect 544075 684934 544081 684952
rect 543927 684932 544081 684934
rect 543927 684922 543973 684932
rect 544035 684922 544081 684932
rect 545145 684934 545151 684952
rect 545185 684934 545259 685002
rect 545293 684992 545299 685002
rect 546363 685002 546409 685014
rect 546471 685002 546517 685014
rect 547581 685002 547627 685014
rect 547689 685002 547735 685014
rect 546363 684992 546369 685002
rect 545293 684952 546369 684992
rect 545293 684934 545299 684952
rect 545145 684932 545299 684934
rect 545145 684922 545191 684932
rect 545253 684922 545299 684932
rect 546363 684934 546369 684952
rect 546403 684934 546477 685002
rect 546511 684992 546519 685002
rect 547579 684992 547587 685002
rect 546511 684952 547587 684992
rect 546511 684934 546519 684952
rect 546363 684932 546519 684934
rect 547579 684934 547587 684952
rect 547621 684934 547695 685002
rect 547729 684992 547735 685002
rect 548799 685002 571820 685014
rect 548799 684992 548805 685002
rect 547729 684952 548805 684992
rect 547729 684934 547735 684952
rect 547579 684932 547735 684934
rect 546363 684922 546409 684932
rect 546471 684922 546517 684932
rect 547581 684922 547627 684932
rect 547689 684922 547735 684932
rect 548799 684934 548805 684952
rect 548839 684934 571820 685002
rect 548799 684922 571820 684934
rect 540459 684906 541459 684912
rect 540459 684892 540471 684906
rect 46436 684860 46482 684872
rect 540449 684872 540471 684892
rect 541447 684892 541459 684906
rect 541677 684906 542677 684912
rect 541677 684892 541689 684906
rect 541447 684872 541689 684892
rect 542665 684892 542677 684906
rect 542895 684906 543895 684912
rect 542895 684892 542907 684906
rect 542665 684872 542907 684892
rect 543883 684892 543895 684906
rect 544113 684906 545113 684912
rect 544113 684892 544125 684906
rect 543883 684872 544125 684892
rect 545101 684892 545113 684906
rect 545331 684906 546331 684912
rect 545331 684892 545343 684906
rect 545101 684872 545343 684892
rect 546319 684892 546331 684906
rect 546549 684906 547549 684912
rect 546549 684892 546561 684906
rect 546319 684872 546561 684892
rect 547537 684892 547549 684906
rect 547767 684906 548767 684912
rect 547767 684892 547779 684906
rect 547537 684872 547779 684892
rect 548755 684892 548767 684906
rect 548755 684872 548779 684892
rect 540449 684862 545769 684872
rect 42250 684830 42260 684860
rect 42240 684780 42260 684830
rect 42250 684750 42260 684780
rect 42370 684830 42380 684860
rect 42500 684830 42510 684860
rect 42370 684780 42510 684830
rect 42370 684750 42380 684780
rect 42500 684750 42510 684780
rect 42620 684830 42630 684860
rect 46650 684830 46660 684860
rect 42620 684822 46660 684830
rect 42620 684788 42892 684822
rect 43060 684788 43150 684822
rect 43318 684788 43408 684822
rect 43576 684788 43666 684822
rect 43834 684788 43924 684822
rect 44092 684788 44182 684822
rect 44350 684788 44440 684822
rect 44608 684788 44698 684822
rect 44866 684788 44956 684822
rect 45124 684788 45214 684822
rect 45382 684788 45472 684822
rect 45640 684788 45730 684822
rect 45898 684788 45988 684822
rect 46156 684788 46246 684822
rect 46414 684788 46660 684822
rect 42620 684780 46660 684788
rect 42620 684750 42630 684780
rect 46650 684750 46660 684780
rect 46770 684830 46780 684860
rect 46900 684830 46910 684860
rect 46770 684780 46910 684830
rect 46770 684750 46780 684780
rect 46900 684750 46910 684780
rect 47020 684830 47030 684860
rect 540449 684852 540759 684862
rect 47020 684780 47040 684830
rect 540749 684782 540759 684852
rect 540849 684782 540899 684862
rect 540989 684852 545769 684862
rect 540989 684782 540999 684852
rect 543339 684802 543439 684852
rect 545759 684802 545769 684852
rect 545859 684802 545909 684872
rect 545999 684852 548779 684872
rect 548820 684860 571820 684922
rect 545999 684802 546009 684852
rect 47020 684750 47030 684780
rect 43690 684720 45616 684726
rect 43690 684686 43702 684720
rect 45604 684686 45616 684720
rect 43690 684680 44530 684686
rect 44520 684470 44530 684680
rect 44780 684680 45616 684686
rect 44780 684470 44790 684680
rect 540759 684632 540989 684782
rect 542267 684772 542401 684778
rect 542267 684662 542279 684772
rect 542389 684662 542401 684772
rect 542267 684656 542401 684662
rect 543127 684772 543261 684778
rect 543127 684662 543139 684772
rect 543249 684662 543261 684772
rect 543127 684656 543261 684662
rect 544337 684772 544471 684778
rect 544337 684662 544349 684772
rect 544459 684662 544471 684772
rect 544337 684656 544471 684662
rect 545187 684772 545321 684778
rect 545187 684662 545199 684772
rect 545309 684662 545321 684772
rect 545187 684656 545321 684662
rect 540749 684582 540759 684632
rect 540449 684564 540759 684582
rect 540849 684564 540899 684632
rect 540989 684582 540999 684632
rect 542129 684582 542229 684632
rect 544549 684582 544649 684652
rect 545769 684622 545999 684802
rect 548219 684792 548319 684852
rect 546757 684772 546891 684778
rect 546757 684662 546769 684772
rect 546879 684662 546891 684772
rect 546757 684656 546891 684662
rect 547637 684772 547771 684778
rect 547637 684662 547649 684772
rect 547759 684662 547771 684772
rect 547637 684656 547771 684662
rect 545759 684582 545769 684622
rect 540989 684564 545769 684582
rect 545859 684564 545909 684622
rect 545999 684582 546009 684622
rect 546979 684582 547079 684642
rect 545999 684564 548779 684582
rect 540449 684542 540471 684564
rect 540459 684530 540471 684542
rect 541447 684542 541689 684564
rect 541447 684530 541459 684542
rect 540459 684524 541459 684530
rect 541677 684530 541689 684542
rect 542665 684542 542907 684564
rect 542665 684530 542677 684542
rect 541677 684524 542677 684530
rect 542895 684530 542907 684542
rect 543883 684542 544125 684564
rect 543883 684530 543895 684542
rect 542895 684524 543895 684530
rect 544113 684530 544125 684542
rect 545101 684542 545343 684564
rect 546319 684542 546561 684564
rect 545101 684530 545113 684542
rect 544113 684524 545113 684530
rect 545331 684530 545343 684542
rect 546319 684530 546331 684542
rect 545331 684524 546331 684530
rect 546549 684530 546561 684542
rect 547537 684542 547779 684564
rect 547537 684530 547549 684542
rect 546549 684524 547549 684530
rect 547767 684530 547779 684542
rect 548755 684542 548779 684564
rect 548755 684530 548767 684542
rect 547767 684524 548767 684530
rect 548820 684514 554960 684580
rect 540381 684502 540427 684514
rect 540381 684434 540387 684502
rect 540421 684492 540427 684502
rect 541491 684502 541537 684514
rect 541491 684492 541497 684502
rect 540421 684452 541497 684492
rect 540421 684434 540427 684452
rect 540381 684422 540427 684434
rect 541491 684434 541497 684452
rect 541531 684492 541537 684502
rect 541599 684502 541645 684514
rect 541599 684492 541605 684502
rect 541531 684452 541605 684492
rect 541531 684434 541537 684452
rect 541491 684422 541537 684434
rect 541599 684434 541605 684452
rect 541639 684492 541645 684502
rect 542709 684502 542755 684514
rect 542817 684502 542863 684514
rect 542709 684492 542715 684502
rect 541639 684452 542715 684492
rect 541639 684434 541645 684452
rect 541599 684422 541645 684434
rect 542709 684434 542715 684452
rect 542749 684434 542823 684502
rect 542857 684492 542863 684502
rect 543927 684502 543973 684514
rect 544035 684502 544081 684514
rect 543927 684492 543933 684502
rect 542857 684452 543933 684492
rect 542857 684434 542863 684452
rect 542709 684432 542863 684434
rect 542709 684422 542755 684432
rect 542817 684422 542863 684432
rect 543927 684434 543933 684452
rect 543967 684434 544041 684502
rect 544075 684492 544081 684502
rect 545145 684502 545191 684514
rect 545253 684502 545299 684514
rect 545145 684492 545151 684502
rect 544075 684452 545151 684492
rect 544075 684434 544081 684452
rect 543927 684432 544081 684434
rect 543927 684422 543973 684432
rect 544035 684422 544081 684432
rect 545145 684434 545151 684452
rect 545185 684434 545259 684502
rect 545293 684492 545299 684502
rect 546363 684502 546409 684514
rect 546471 684502 546517 684514
rect 547581 684502 547627 684514
rect 547689 684502 547735 684514
rect 546363 684492 546369 684502
rect 545293 684452 546369 684492
rect 545293 684434 545299 684452
rect 545145 684432 545299 684434
rect 545145 684422 545191 684432
rect 545253 684422 545299 684432
rect 546363 684434 546369 684452
rect 546403 684434 546477 684502
rect 546511 684492 546519 684502
rect 547579 684492 547587 684502
rect 546511 684452 547587 684492
rect 546511 684434 546519 684452
rect 546363 684432 546519 684434
rect 547579 684434 547587 684452
rect 547621 684434 547695 684502
rect 547729 684492 547735 684502
rect 548799 684502 554960 684514
rect 548799 684492 548805 684502
rect 547729 684452 548805 684492
rect 547729 684434 547735 684452
rect 547579 684432 547735 684434
rect 546363 684422 546409 684432
rect 546471 684422 546517 684432
rect 547581 684422 547627 684432
rect 547689 684422 547735 684432
rect 548799 684434 548805 684452
rect 548839 684434 554960 684502
rect 548799 684422 554960 684434
rect 540459 684406 541459 684412
rect 540459 684392 540471 684406
rect 540449 684372 540471 684392
rect 541447 684392 541459 684406
rect 541677 684406 542677 684412
rect 541677 684392 541689 684406
rect 541447 684372 541689 684392
rect 542665 684392 542677 684406
rect 542895 684406 543895 684412
rect 542895 684392 542907 684406
rect 543883 684392 543895 684406
rect 544113 684406 545113 684412
rect 544113 684392 544125 684406
rect 542665 684372 542907 684392
rect 543883 684372 544125 684392
rect 545101 684392 545113 684406
rect 545331 684406 546331 684412
rect 545331 684392 545343 684406
rect 546319 684392 546331 684406
rect 546549 684406 547549 684412
rect 546549 684392 546561 684406
rect 545101 684372 545343 684392
rect 546319 684372 546561 684392
rect 547537 684392 547549 684406
rect 547767 684406 548767 684412
rect 547767 684392 547779 684406
rect 547537 684372 547779 684392
rect 548755 684392 548767 684406
rect 548755 684372 548779 684392
rect 540449 684352 541089 684372
rect 540889 684302 540989 684352
rect 541079 684292 541089 684352
rect 541169 684352 541239 684372
rect 541169 684292 541179 684352
rect 541229 684292 541239 684352
rect 541319 684352 543579 684372
rect 541319 684292 541329 684352
rect 542039 684332 542189 684352
rect 543279 684322 543439 684352
rect 543339 684302 543439 684322
rect 543569 684312 543579 684352
rect 543659 684352 543729 684372
rect 543659 684312 543669 684352
rect 543719 684312 543729 684352
rect 543809 684352 546059 684372
rect 543809 684312 543819 684352
rect 544519 684322 544669 684352
rect 545779 684292 545879 684352
rect 546049 684312 546059 684352
rect 546139 684352 546199 684372
rect 546139 684312 546149 684352
rect 546189 684312 546199 684352
rect 546279 684352 548779 684372
rect 548820 684360 554960 684422
rect 546279 684312 546289 684352
rect 546989 684322 547139 684352
rect 548219 684322 548369 684352
rect 548219 684292 548319 684322
rect 541449 684142 541759 684172
rect 541329 684082 541539 684142
rect 541009 684064 541539 684082
rect 541619 684064 541649 684142
rect 541729 684082 541759 684142
rect 546389 684132 546609 684142
rect 543939 684082 543949 684112
rect 541729 684064 543949 684082
rect 544029 684082 544039 684112
rect 546389 684082 546399 684132
rect 544029 684064 546399 684082
rect 546479 684064 546519 684132
rect 546599 684082 546609 684132
rect 547589 684082 547599 684122
rect 546599 684064 547599 684082
rect 547679 684082 547689 684122
rect 547679 684064 548129 684082
rect 541009 684042 541031 684064
rect 541019 684030 541031 684042
rect 542007 684042 542249 684064
rect 542007 684030 542019 684042
rect 541019 684024 542019 684030
rect 542237 684030 542249 684042
rect 543225 684042 543467 684064
rect 543225 684030 543237 684042
rect 542237 684024 543237 684030
rect 543455 684030 543467 684042
rect 544443 684042 544685 684064
rect 544443 684030 544455 684042
rect 543455 684024 544455 684030
rect 544673 684030 544685 684042
rect 545661 684042 545903 684064
rect 545661 684030 545673 684042
rect 544673 684024 545673 684030
rect 545891 684030 545903 684042
rect 546879 684042 547121 684064
rect 548097 684042 548129 684064
rect 546879 684030 546891 684042
rect 545891 684024 546891 684030
rect 547109 684030 547121 684042
rect 548097 684030 548109 684042
rect 547109 684024 548109 684030
rect 540941 684002 540987 684014
rect 540941 683982 540947 684002
rect 43600 683900 45700 683910
rect 43600 683866 43922 683900
rect 44090 683866 44180 683900
rect 44348 683866 44438 683900
rect 44606 683866 44696 683900
rect 44864 683866 44954 683900
rect 45122 683866 45212 683900
rect 45380 683866 45700 683900
rect 43600 683860 45700 683866
rect 540929 683862 540947 683982
rect 43600 682780 43670 683860
rect 43854 683807 43900 683819
rect 43854 683600 43860 683807
rect 43894 683600 43900 683807
rect 44112 683807 44158 683819
rect 43830 683520 43840 683600
rect 43920 683520 43930 683600
rect 43854 683450 43860 683520
rect 43730 683430 43860 683450
rect 43730 683200 43740 683430
rect 43780 683200 43860 683430
rect 43730 683180 43860 683200
rect 43854 682831 43860 683180
rect 43894 682831 43900 683520
rect 44112 683120 44118 683807
rect 44152 683120 44158 683807
rect 44370 683807 44416 683819
rect 44370 683600 44376 683807
rect 44410 683600 44416 683807
rect 44628 683807 44674 683819
rect 44340 683520 44350 683600
rect 44430 683520 44440 683600
rect 44080 683040 44090 683120
rect 44170 683040 44180 683120
rect 43854 682819 43900 682831
rect 44112 682831 44118 683040
rect 44152 682831 44158 683040
rect 44112 682819 44158 682831
rect 44370 682831 44376 683520
rect 44410 682831 44416 683520
rect 44628 683120 44634 683807
rect 44668 683120 44674 683807
rect 44886 683807 44932 683819
rect 44886 683600 44892 683807
rect 44926 683600 44932 683807
rect 45144 683807 45190 683819
rect 44860 683520 44870 683600
rect 44950 683520 44960 683600
rect 44600 683040 44610 683120
rect 44690 683040 44700 683120
rect 44370 682819 44416 682831
rect 44628 682831 44634 683040
rect 44668 682831 44674 683040
rect 44628 682819 44674 682831
rect 44886 682831 44892 683520
rect 44926 682831 44932 683520
rect 45144 683120 45150 683807
rect 45184 683120 45190 683807
rect 45402 683807 45448 683819
rect 45402 683600 45408 683807
rect 45442 683600 45448 683807
rect 45380 683520 45390 683600
rect 45470 683520 45480 683600
rect 45402 683450 45408 683520
rect 45400 683180 45408 683450
rect 45120 683040 45130 683120
rect 45210 683040 45220 683120
rect 44886 682819 44932 682831
rect 45144 682831 45150 683040
rect 45184 682831 45190 683040
rect 45144 682819 45190 682831
rect 45402 682831 45408 683180
rect 45442 683450 45448 683520
rect 45442 683430 45570 683450
rect 45442 683200 45520 683430
rect 45560 683200 45570 683430
rect 45442 683180 45570 683200
rect 45442 682831 45448 683180
rect 45402 682819 45448 682831
rect 45630 682780 45700 683860
rect 540941 683834 540947 683862
rect 540981 683982 540987 684002
rect 542051 684002 542097 684014
rect 542051 683982 542057 684002
rect 540981 683862 542057 683982
rect 540981 683834 540987 683862
rect 540941 683822 540987 683834
rect 542051 683834 542057 683862
rect 542091 683982 542097 684002
rect 542159 684002 542205 684014
rect 542159 683982 542165 684002
rect 542091 683862 542165 683982
rect 542091 683834 542097 683862
rect 542051 683822 542097 683834
rect 542159 683834 542165 683862
rect 542199 683982 542205 684002
rect 543269 684002 543315 684014
rect 543269 683982 543275 684002
rect 542199 683962 543275 683982
rect 542199 683882 542719 683962
rect 542799 683882 543275 683962
rect 542199 683862 543275 683882
rect 542199 683834 542205 683862
rect 542159 683822 542205 683834
rect 543269 683834 543275 683862
rect 543309 683982 543315 684002
rect 543377 684002 543423 684014
rect 543377 683982 543383 684002
rect 543309 683862 543383 683982
rect 543309 683834 543315 683862
rect 543269 683822 543315 683834
rect 543377 683834 543383 683862
rect 543417 683982 543423 684002
rect 544487 684002 544533 684014
rect 544487 683982 544493 684002
rect 543417 683862 544493 683982
rect 543417 683834 543423 683862
rect 543377 683822 543423 683834
rect 544487 683834 544493 683862
rect 544527 683982 544533 684002
rect 544595 684002 544641 684014
rect 544595 683982 544601 684002
rect 544527 683862 544601 683982
rect 544527 683834 544533 683862
rect 544487 683822 544533 683834
rect 544595 683834 544601 683862
rect 544635 683982 544641 684002
rect 545705 684002 545751 684014
rect 545705 683982 545711 684002
rect 544635 683962 545711 683982
rect 544635 683882 545129 683962
rect 545209 683882 545711 683962
rect 544635 683862 545711 683882
rect 544635 683834 544641 683862
rect 544595 683822 544641 683834
rect 545705 683834 545711 683862
rect 545745 683982 545751 684002
rect 545813 684002 545859 684014
rect 545813 683982 545819 684002
rect 545745 683862 545819 683982
rect 545745 683834 545751 683862
rect 545705 683822 545751 683834
rect 545813 683834 545819 683862
rect 545853 683982 545859 684002
rect 546923 684002 546969 684014
rect 546923 683982 546929 684002
rect 545853 683862 546929 683982
rect 545853 683834 545859 683862
rect 545813 683822 545859 683834
rect 546923 683834 546929 683862
rect 546963 683982 546969 684002
rect 547031 684002 547077 684014
rect 547031 683982 547037 684002
rect 546963 683862 547037 683982
rect 546963 683834 546969 683862
rect 546923 683822 546969 683834
rect 547031 683834 547037 683862
rect 547071 683982 547077 684002
rect 548141 684002 548187 684014
rect 548141 683982 548147 684002
rect 547071 683862 548147 683982
rect 547071 683834 547077 683862
rect 547031 683822 547077 683834
rect 548141 683834 548147 683862
rect 548181 683834 548187 684002
rect 548141 683822 548187 683834
rect 541019 683806 542019 683812
rect 541019 683782 541031 683806
rect 542007 683782 542019 683806
rect 542237 683806 543237 683812
rect 542237 683782 542249 683806
rect 541009 683772 541031 683782
rect 542007 683772 542249 683782
rect 543225 683782 543237 683806
rect 543455 683806 544455 683812
rect 543455 683782 543467 683806
rect 543225 683772 543467 683782
rect 544443 683782 544455 683806
rect 544673 683806 545673 683812
rect 544673 683782 544685 683806
rect 544443 683772 544685 683782
rect 545661 683782 545673 683806
rect 545891 683806 546891 683812
rect 545891 683782 545903 683806
rect 546879 683782 546891 683806
rect 547109 683806 548109 683812
rect 547109 683782 547121 683806
rect 545661 683772 545903 683782
rect 546879 683772 547121 683782
rect 548097 683782 548109 683806
rect 548097 683772 548129 683782
rect 541009 683742 541459 683772
rect 541449 683702 541459 683742
rect 541539 683742 546349 683772
rect 541539 683702 541549 683742
rect 546339 683702 546349 683742
rect 546429 683742 548129 683772
rect 546429 683702 546439 683742
rect 541557 683652 541691 683658
rect 541557 683562 541569 683652
rect 541679 683562 541691 683652
rect 541557 683556 541691 683562
rect 546467 683652 546601 683658
rect 546467 683562 546479 683652
rect 546589 683562 546601 683652
rect 546467 683556 546601 683562
rect 543939 683462 543949 683492
rect 541009 683444 543949 683462
rect 544029 683462 544039 683492
rect 547589 683462 547599 683502
rect 544029 683444 547599 683462
rect 547679 683462 547689 683502
rect 547679 683444 548129 683462
rect 541009 683422 541031 683444
rect 541019 683410 541031 683422
rect 542007 683422 542249 683444
rect 542007 683410 542019 683422
rect 541019 683404 542019 683410
rect 542237 683410 542249 683422
rect 543225 683422 543467 683444
rect 543225 683410 543237 683422
rect 542237 683404 543237 683410
rect 543455 683410 543467 683422
rect 544443 683422 544685 683444
rect 544443 683410 544455 683422
rect 543455 683404 544455 683410
rect 544673 683410 544685 683422
rect 545661 683422 545903 683444
rect 545661 683410 545673 683422
rect 544673 683404 545673 683410
rect 545891 683410 545903 683422
rect 546879 683422 547121 683444
rect 548097 683422 548129 683444
rect 546879 683410 546891 683422
rect 545891 683404 546891 683410
rect 547109 683410 547121 683422
rect 548097 683410 548109 683422
rect 547109 683404 548109 683410
rect 540941 683382 540987 683394
rect 540941 683352 540947 683382
rect 540909 683252 540947 683352
rect 540941 683214 540947 683252
rect 540981 683362 540987 683382
rect 542051 683382 542097 683394
rect 542051 683362 542057 683382
rect 540981 683242 542057 683362
rect 540981 683214 540987 683242
rect 540941 683202 540987 683214
rect 542051 683214 542057 683242
rect 542091 683362 542097 683382
rect 542159 683382 542205 683394
rect 542159 683362 542165 683382
rect 542091 683342 542165 683362
rect 542199 683362 542205 683382
rect 543269 683382 543315 683394
rect 543269 683362 543275 683382
rect 542199 683342 543275 683362
rect 542091 683262 542109 683342
rect 542199 683262 542229 683342
rect 542319 683262 542719 683342
rect 542799 683262 543275 683342
rect 542091 683242 542165 683262
rect 542091 683214 542097 683242
rect 542051 683202 542097 683214
rect 542159 683214 542165 683242
rect 542199 683242 543275 683262
rect 542199 683214 542205 683242
rect 542159 683202 542205 683214
rect 543269 683214 543275 683242
rect 543309 683362 543315 683382
rect 543377 683382 543423 683394
rect 543377 683362 543383 683382
rect 543309 683242 543383 683362
rect 543309 683214 543315 683242
rect 543269 683202 543315 683214
rect 543377 683214 543383 683242
rect 543417 683362 543423 683382
rect 544487 683382 544533 683394
rect 544487 683362 544493 683382
rect 543417 683242 544493 683362
rect 543417 683214 543423 683242
rect 543377 683202 543423 683214
rect 544487 683214 544493 683242
rect 544527 683362 544533 683382
rect 544595 683382 544641 683394
rect 544595 683362 544601 683382
rect 544527 683342 544601 683362
rect 544635 683362 544641 683382
rect 545705 683382 545751 683394
rect 545705 683362 545711 683382
rect 544635 683342 545711 683362
rect 544527 683262 544559 683342
rect 544649 683262 544679 683342
rect 544769 683262 545129 683342
rect 545209 683262 545711 683342
rect 544527 683242 544601 683262
rect 544527 683214 544533 683242
rect 544487 683202 544533 683214
rect 544595 683214 544601 683242
rect 544635 683242 545711 683262
rect 544635 683214 544641 683242
rect 544595 683202 544641 683214
rect 545705 683214 545711 683242
rect 545745 683362 545751 683382
rect 545813 683382 545859 683394
rect 545813 683362 545819 683382
rect 545745 683242 545819 683362
rect 545745 683214 545751 683242
rect 545705 683202 545751 683214
rect 545813 683214 545819 683242
rect 545853 683362 545859 683382
rect 546923 683382 546969 683394
rect 546923 683362 546929 683382
rect 545853 683242 546929 683362
rect 545853 683214 545859 683242
rect 545813 683202 545859 683214
rect 546923 683214 546929 683242
rect 546963 683362 546969 683382
rect 547031 683382 547077 683394
rect 547031 683362 547037 683382
rect 546963 683342 547037 683362
rect 547071 683362 547077 683382
rect 548141 683382 548187 683394
rect 548141 683362 548147 683382
rect 547071 683342 548147 683362
rect 546963 683262 546989 683342
rect 547079 683262 547109 683342
rect 547199 683262 548147 683342
rect 546963 683242 547037 683262
rect 546963 683214 546969 683242
rect 546923 683202 546969 683214
rect 547031 683214 547037 683242
rect 547071 683242 548147 683262
rect 547071 683214 547077 683242
rect 547031 683202 547077 683214
rect 548141 683214 548147 683242
rect 548181 683362 548187 683382
rect 548181 683242 548189 683362
rect 548181 683214 548187 683242
rect 548141 683202 548187 683214
rect 541019 683186 542019 683192
rect 541019 683162 541031 683186
rect 542007 683162 542019 683186
rect 542237 683186 543237 683192
rect 542237 683162 542249 683186
rect 541009 683152 541031 683162
rect 542007 683152 542249 683162
rect 543225 683162 543237 683186
rect 543455 683186 544455 683192
rect 543455 683162 543467 683186
rect 543225 683152 543467 683162
rect 544443 683162 544455 683186
rect 544673 683186 545673 683192
rect 544673 683162 544685 683186
rect 544443 683152 544685 683162
rect 545661 683162 545673 683186
rect 545891 683186 546891 683192
rect 545891 683162 545903 683186
rect 546879 683162 546891 683186
rect 547109 683186 548109 683192
rect 547109 683162 547121 683186
rect 545661 683152 545903 683162
rect 546879 683152 547121 683162
rect 548097 683162 548109 683186
rect 548097 683152 548129 683162
rect 541009 683122 541459 683152
rect 541449 683082 541459 683122
rect 541539 683122 546349 683152
rect 541539 683082 541549 683122
rect 546339 683082 546349 683122
rect 546429 683122 548129 683152
rect 546429 683082 546439 683122
rect 543329 682882 543339 682912
rect 540449 682844 543339 682882
rect 543429 682882 543439 682912
rect 548209 682882 548219 682932
rect 543429 682852 548219 682882
rect 548309 682882 548319 682932
rect 548309 682852 548769 682882
rect 543429 682844 548769 682852
rect 540449 682842 540471 682844
rect 540459 682810 540471 682842
rect 541447 682842 541689 682844
rect 541447 682810 541459 682842
rect 540459 682804 541459 682810
rect 541677 682810 541689 682842
rect 542665 682842 542907 682844
rect 542665 682810 542677 682842
rect 541677 682804 542677 682810
rect 542895 682810 542907 682842
rect 543883 682842 544125 682844
rect 543883 682810 543895 682842
rect 542895 682804 543895 682810
rect 544113 682810 544125 682842
rect 545101 682842 545343 682844
rect 545101 682810 545113 682842
rect 544113 682804 545113 682810
rect 545331 682810 545343 682842
rect 546319 682842 546561 682844
rect 546319 682810 546331 682842
rect 545331 682804 546331 682810
rect 546549 682810 546561 682842
rect 547537 682842 547779 682844
rect 547537 682810 547549 682842
rect 546549 682804 547549 682810
rect 547767 682810 547779 682842
rect 548755 682842 548769 682844
rect 548755 682810 548767 682842
rect 547767 682804 548767 682810
rect 43600 682772 45700 682780
rect 43600 682770 43922 682772
rect 43600 682730 43920 682770
rect 44090 682738 44180 682772
rect 44348 682738 44438 682772
rect 44606 682770 44696 682772
rect 44606 682738 44620 682770
rect 43910 682700 43920 682730
rect 43990 682730 44620 682738
rect 43990 682700 44000 682730
rect 44610 682700 44620 682730
rect 44690 682738 44696 682770
rect 44864 682738 44954 682772
rect 45122 682738 45212 682772
rect 44690 682730 45310 682738
rect 44690 682700 44700 682730
rect 45300 682700 45310 682730
rect 45380 682730 45700 682772
rect 540381 682782 540427 682794
rect 540381 682762 540387 682782
rect 45380 682700 45390 682730
rect 540369 682642 540387 682762
rect 540381 682614 540387 682642
rect 540421 682762 540427 682782
rect 541491 682782 541537 682794
rect 541491 682762 541497 682782
rect 540421 682642 541497 682762
rect 540421 682614 540427 682642
rect 540381 682602 540427 682614
rect 541491 682614 541497 682642
rect 541531 682762 541537 682782
rect 541599 682782 541645 682794
rect 541599 682762 541605 682782
rect 541531 682642 541605 682762
rect 541531 682614 541537 682642
rect 541491 682602 541537 682614
rect 541599 682614 541605 682642
rect 541639 682762 541645 682782
rect 542709 682782 542755 682794
rect 542709 682762 542715 682782
rect 541639 682742 542715 682762
rect 541639 682662 542109 682742
rect 542199 682662 542229 682742
rect 542319 682662 542715 682742
rect 541639 682642 542715 682662
rect 541639 682614 541645 682642
rect 541599 682602 541645 682614
rect 542709 682614 542715 682642
rect 542749 682762 542755 682782
rect 542817 682782 542863 682794
rect 542817 682762 542823 682782
rect 542749 682642 542823 682762
rect 542749 682614 542755 682642
rect 542709 682602 542755 682614
rect 542817 682614 542823 682642
rect 542857 682762 542863 682782
rect 543927 682782 543973 682794
rect 543927 682762 543933 682782
rect 542857 682642 543933 682762
rect 542857 682614 542863 682642
rect 542817 682602 542863 682614
rect 543927 682614 543933 682642
rect 543967 682762 543973 682782
rect 544035 682782 544081 682794
rect 544035 682762 544041 682782
rect 543967 682642 544041 682762
rect 543967 682614 543973 682642
rect 543927 682602 543973 682614
rect 544035 682614 544041 682642
rect 544075 682762 544081 682782
rect 545145 682782 545191 682794
rect 545145 682762 545151 682782
rect 544075 682742 545151 682762
rect 544075 682662 544559 682742
rect 544649 682662 544679 682742
rect 544769 682662 545151 682742
rect 544075 682642 545151 682662
rect 544075 682614 544081 682642
rect 544035 682602 544081 682614
rect 545145 682614 545151 682642
rect 545185 682762 545191 682782
rect 545253 682782 545299 682794
rect 545253 682762 545259 682782
rect 545185 682642 545259 682762
rect 545185 682614 545191 682642
rect 545145 682602 545191 682614
rect 545253 682614 545259 682642
rect 545293 682762 545299 682782
rect 546363 682782 546409 682794
rect 546363 682762 546369 682782
rect 545293 682642 546369 682762
rect 545293 682614 545299 682642
rect 545253 682602 545299 682614
rect 546363 682614 546369 682642
rect 546403 682762 546409 682782
rect 546471 682782 546517 682794
rect 546471 682762 546477 682782
rect 546403 682642 546477 682762
rect 546403 682614 546409 682642
rect 546363 682602 546409 682614
rect 546471 682614 546477 682642
rect 546511 682762 546517 682782
rect 547581 682782 547627 682794
rect 547581 682762 547587 682782
rect 546511 682742 547587 682762
rect 546511 682662 546989 682742
rect 547079 682662 547109 682742
rect 547199 682662 547587 682742
rect 546511 682642 547587 682662
rect 546511 682614 546517 682642
rect 546471 682602 546517 682614
rect 547581 682614 547587 682642
rect 547621 682762 547627 682782
rect 547689 682782 547735 682794
rect 547689 682762 547695 682782
rect 547621 682642 547695 682762
rect 547621 682614 547627 682642
rect 547581 682602 547627 682614
rect 547689 682614 547695 682642
rect 547729 682762 547735 682782
rect 548799 682782 548845 682794
rect 548799 682762 548805 682782
rect 547729 682642 548805 682762
rect 547729 682614 547735 682642
rect 547689 682602 547735 682614
rect 548799 682614 548805 682642
rect 548839 682762 548845 682782
rect 548839 682642 548849 682762
rect 548839 682614 548845 682642
rect 548799 682602 548845 682614
rect 540459 682586 541459 682592
rect 540459 682562 540471 682586
rect 540449 682552 540471 682562
rect 541447 682562 541459 682586
rect 541677 682586 542677 682592
rect 541677 682562 541689 682586
rect 541447 682552 541689 682562
rect 542665 682562 542677 682586
rect 542895 682586 543895 682592
rect 542895 682562 542907 682586
rect 542665 682552 542907 682562
rect 543883 682562 543895 682586
rect 544113 682586 545113 682592
rect 544113 682562 544125 682586
rect 543883 682552 544125 682562
rect 545101 682562 545113 682586
rect 545331 682586 546331 682592
rect 545331 682562 545343 682586
rect 545101 682552 545343 682562
rect 546319 682562 546331 682586
rect 546549 682586 547549 682592
rect 546549 682562 546561 682586
rect 546319 682552 546561 682562
rect 547537 682562 547549 682586
rect 547767 682586 548767 682592
rect 547767 682562 547779 682586
rect 547537 682552 547779 682562
rect 548755 682562 548767 682586
rect 548755 682552 548769 682562
rect 540449 682522 540759 682552
rect 540749 682502 540759 682522
rect 540849 682522 540899 682552
rect 540849 682502 540859 682522
rect 540889 682502 540899 682522
rect 540989 682522 545769 682552
rect 540989 682502 540999 682522
rect 545759 682502 545769 682522
rect 545859 682522 545909 682552
rect 545859 682502 545869 682522
rect 545899 682502 545909 682522
rect 545999 682522 548769 682552
rect 545999 682502 546009 682522
rect 541489 682452 541649 682462
rect 43910 682410 43920 682440
rect 43900 682370 43920 682410
rect 43990 682410 44000 682440
rect 44610 682410 44620 682440
rect 43990 682400 44620 682410
rect 43900 682366 43922 682370
rect 44090 682366 44180 682400
rect 44348 682366 44438 682400
rect 44606 682370 44620 682400
rect 44690 682410 44700 682440
rect 45300 682410 45310 682440
rect 44690 682400 45310 682410
rect 45380 682410 45390 682440
rect 44690 682370 44696 682400
rect 44606 682366 44696 682370
rect 44864 682366 44954 682400
rect 45122 682366 45212 682400
rect 45380 682366 45400 682410
rect 43900 682360 45400 682366
rect 43854 682307 43900 682319
rect 43854 682140 43860 682307
rect 43894 682140 43900 682307
rect 44110 682307 44160 682360
rect 44630 682319 44680 682360
rect 44110 682200 44118 682307
rect 43830 682060 43840 682140
rect 43920 682060 43930 682140
rect 43570 681920 43790 681940
rect 43570 681840 43630 681920
rect 43710 681840 43740 681920
rect 43570 681780 43740 681840
rect 43570 681700 43630 681780
rect 43710 681700 43740 681780
rect 43570 681690 43740 681700
rect 43780 681690 43790 681920
rect 43570 681680 43790 681690
rect 43734 681678 43786 681680
rect 43854 681331 43860 682060
rect 43894 681331 43900 682060
rect 44112 681440 44118 682200
rect 43854 681319 43900 681331
rect 44110 681331 44118 681440
rect 44152 682200 44160 682307
rect 44370 682307 44416 682319
rect 44152 681440 44158 682200
rect 44370 682140 44376 682307
rect 44410 682140 44416 682307
rect 44628 682307 44680 682319
rect 44340 682060 44350 682140
rect 44430 682060 44440 682140
rect 44152 681331 44160 681440
rect 44110 681280 44160 681331
rect 44370 681331 44376 682060
rect 44410 681331 44416 682060
rect 44370 681319 44416 681331
rect 44628 681331 44634 682307
rect 44668 682200 44680 682307
rect 44886 682307 44932 682319
rect 44668 681450 44674 682200
rect 44886 682140 44892 682307
rect 44926 682140 44932 682307
rect 45140 682307 45190 682360
rect 541489 682352 541509 682452
rect 541629 682352 541649 682452
rect 45140 682200 45150 682307
rect 44860 682060 44870 682140
rect 44950 682060 44960 682140
rect 44668 681331 44680 681450
rect 44628 681319 44680 681331
rect 44886 681331 44892 682060
rect 44926 681331 44932 682060
rect 45144 681440 45150 682200
rect 44886 681319 44932 681331
rect 45140 681331 45150 681440
rect 45184 681331 45190 682307
rect 45402 682307 45448 682319
rect 45402 682140 45408 682307
rect 45442 682140 45448 682307
rect 541489 682282 541649 682352
rect 542709 682452 542869 682462
rect 542709 682352 542729 682452
rect 542849 682352 542869 682452
rect 542709 682282 542869 682352
rect 543919 682452 544079 682462
rect 545147 682452 545291 682458
rect 547587 682452 547731 682458
rect 543919 682352 543939 682452
rect 544059 682352 544079 682452
rect 543329 682282 543339 682312
rect 540449 682244 543339 682282
rect 543429 682282 543439 682312
rect 543919 682282 544079 682352
rect 545139 682352 545159 682452
rect 545279 682352 545299 682452
rect 546377 682442 546521 682448
rect 545139 682282 545299 682352
rect 546369 682342 546389 682442
rect 546509 682342 546529 682442
rect 546369 682282 546529 682342
rect 547579 682352 547599 682452
rect 547719 682352 547739 682452
rect 547579 682282 547739 682352
rect 548209 682282 548219 682332
rect 543429 682252 548219 682282
rect 548309 682282 548319 682332
rect 554420 682300 554960 684360
rect 548309 682252 548769 682282
rect 543429 682244 548769 682252
rect 540449 682242 540471 682244
rect 540459 682210 540471 682242
rect 541447 682242 541689 682244
rect 541447 682210 541459 682242
rect 540459 682204 541459 682210
rect 541677 682210 541689 682242
rect 542665 682242 542907 682244
rect 542665 682210 542677 682242
rect 541677 682204 542677 682210
rect 542895 682210 542907 682242
rect 543883 682242 544125 682244
rect 543883 682210 543895 682242
rect 542895 682204 543895 682210
rect 544113 682210 544125 682242
rect 545101 682242 545343 682244
rect 545101 682210 545113 682242
rect 544113 682204 545113 682210
rect 545331 682210 545343 682242
rect 546319 682242 546561 682244
rect 546319 682210 546331 682242
rect 545331 682204 546331 682210
rect 546549 682210 546561 682242
rect 547537 682242 547779 682244
rect 547537 682210 547549 682242
rect 546549 682204 547549 682210
rect 547767 682210 547779 682242
rect 548755 682242 548769 682244
rect 548755 682210 548767 682242
rect 547767 682204 548767 682210
rect 554420 682200 563740 682300
rect 540381 682182 540427 682194
rect 45380 682060 45390 682140
rect 45470 682060 45480 682140
rect 44630 681280 44680 681319
rect 45140 681280 45190 681331
rect 45402 681331 45408 682060
rect 45442 681331 45448 682060
rect 540381 682014 540387 682182
rect 540421 682162 540427 682182
rect 541491 682182 541537 682194
rect 541491 682162 541497 682182
rect 540421 682042 541497 682162
rect 540421 682014 540427 682042
rect 540381 682002 540427 682014
rect 541491 682014 541497 682042
rect 541531 682162 541537 682182
rect 541599 682182 541645 682194
rect 541599 682162 541605 682182
rect 541531 682042 541605 682162
rect 541531 682014 541537 682042
rect 541491 682002 541537 682014
rect 541599 682014 541605 682042
rect 541639 682162 541645 682182
rect 542709 682182 542755 682194
rect 542709 682162 542715 682182
rect 541639 682142 542715 682162
rect 541639 682062 542109 682142
rect 542199 682062 542229 682142
rect 542319 682062 542715 682142
rect 541639 682042 542715 682062
rect 541639 682014 541645 682042
rect 541599 682002 541645 682014
rect 542709 682014 542715 682042
rect 542749 682162 542755 682182
rect 542817 682182 542863 682194
rect 542817 682162 542823 682182
rect 542749 682042 542823 682162
rect 542749 682014 542755 682042
rect 542709 682002 542755 682014
rect 542817 682014 542823 682042
rect 542857 682162 542863 682182
rect 543927 682182 543973 682194
rect 543927 682162 543933 682182
rect 542857 682042 543933 682162
rect 542857 682014 542863 682042
rect 542817 682002 542863 682014
rect 543927 682014 543933 682042
rect 543967 682162 543973 682182
rect 544035 682182 544081 682194
rect 544035 682162 544041 682182
rect 543967 682042 544041 682162
rect 543967 682014 543973 682042
rect 543927 682002 543973 682014
rect 544035 682014 544041 682042
rect 544075 682162 544081 682182
rect 545145 682182 545191 682194
rect 545145 682162 545151 682182
rect 544075 682146 545151 682162
rect 544075 682056 544420 682146
rect 544508 682142 545151 682146
rect 544508 682062 544559 682142
rect 544649 682062 544679 682142
rect 544769 682062 545151 682142
rect 544508 682056 545151 682062
rect 544075 682042 545151 682056
rect 544075 682014 544081 682042
rect 544035 682002 544081 682014
rect 545145 682014 545151 682042
rect 545185 682162 545191 682182
rect 545253 682182 545299 682194
rect 545253 682162 545259 682182
rect 545185 682042 545259 682162
rect 545185 682014 545191 682042
rect 545145 682002 545191 682014
rect 545253 682014 545259 682042
rect 545293 682162 545299 682182
rect 546363 682182 546409 682194
rect 546363 682162 546369 682182
rect 545293 682042 546369 682162
rect 545293 682014 545299 682042
rect 545253 682002 545299 682014
rect 546363 682014 546369 682042
rect 546403 682162 546409 682182
rect 546471 682182 546517 682194
rect 546471 682162 546477 682182
rect 546403 682042 546477 682162
rect 546403 682014 546409 682042
rect 546363 682002 546409 682014
rect 546471 682014 546477 682042
rect 546511 682162 546517 682182
rect 547581 682182 547627 682194
rect 547581 682162 547587 682182
rect 546511 682142 547587 682162
rect 546511 682062 546989 682142
rect 547079 682062 547109 682142
rect 547199 682062 547587 682142
rect 546511 682042 547587 682062
rect 546511 682014 546517 682042
rect 546471 682002 546517 682014
rect 547581 682014 547587 682042
rect 547621 682162 547627 682182
rect 547689 682182 547735 682194
rect 547689 682162 547695 682182
rect 547621 682042 547695 682162
rect 547621 682014 547627 682042
rect 547581 682002 547627 682014
rect 547689 682014 547695 682042
rect 547729 682162 547735 682182
rect 548799 682182 548845 682194
rect 548799 682162 548805 682182
rect 547729 682042 548805 682162
rect 547729 682014 547735 682042
rect 547689 682002 547735 682014
rect 548799 682014 548805 682042
rect 548839 682162 548845 682182
rect 548839 682042 548849 682162
rect 548839 682014 548845 682042
rect 548799 682002 548845 682014
rect 554420 682000 561700 682200
rect 561900 682000 562100 682200
rect 562300 682000 562500 682200
rect 562700 682000 562900 682200
rect 563100 682000 563300 682200
rect 563500 682000 563740 682200
rect 540459 681986 541459 681992
rect 540459 681962 540471 681986
rect 541447 681962 541459 681986
rect 541677 681986 542677 681992
rect 541677 681962 541689 681986
rect 540449 681952 540471 681962
rect 541447 681952 541689 681962
rect 542665 681962 542677 681986
rect 542895 681986 543895 681992
rect 542895 681962 542907 681986
rect 542665 681952 542907 681962
rect 543883 681962 543895 681986
rect 544113 681986 545113 681992
rect 544113 681962 544125 681986
rect 543883 681952 544125 681962
rect 545101 681962 545113 681986
rect 545331 681986 546331 681992
rect 545331 681962 545343 681986
rect 545101 681952 545343 681962
rect 546319 681962 546331 681986
rect 546549 681986 547549 681992
rect 546549 681962 546561 681986
rect 546319 681952 546561 681962
rect 547537 681962 547549 681986
rect 547767 681986 548767 681992
rect 547767 681962 547779 681986
rect 547537 681952 547779 681962
rect 548755 681962 548767 681986
rect 548755 681952 548769 681962
rect 45510 681920 45730 681940
rect 540449 681922 540759 681952
rect 45510 681690 45520 681920
rect 45560 681840 45590 681920
rect 45670 681840 45730 681920
rect 540749 681882 540759 681922
rect 540849 681922 540899 681952
rect 540849 681882 540859 681922
rect 540889 681882 540899 681922
rect 540989 681922 545769 681952
rect 540989 681882 540999 681922
rect 545759 681902 545769 681922
rect 545859 681922 545909 681952
rect 545859 681902 545869 681922
rect 545899 681902 545909 681922
rect 545999 681922 548769 681952
rect 545999 681902 546009 681922
rect 45560 681780 45730 681840
rect 45560 681700 45590 681780
rect 45670 681700 45730 681780
rect 45560 681690 45730 681700
rect 45510 681680 45730 681690
rect 554420 681800 563740 682000
rect 45514 681678 45566 681680
rect 554420 681600 561700 681800
rect 561900 681600 562100 681800
rect 562300 681600 562500 681800
rect 562700 681600 562900 681800
rect 563100 681600 563300 681800
rect 563500 681600 563740 681800
rect 541372 681478 541556 681484
rect 542432 681478 542616 681484
rect 543892 681478 544076 681484
rect 545112 681478 545296 681484
rect 546592 681478 546776 681484
rect 547592 681478 547776 681484
rect 45402 681319 45448 681331
rect 541004 681318 541384 681478
rect 541544 681318 542444 681478
rect 542604 681318 543904 681478
rect 544064 681318 545124 681478
rect 545284 681318 546604 681478
rect 546764 681318 547604 681478
rect 547764 681318 548204 681478
rect 43790 681274 45480 681280
rect 43790 681272 44420 681274
rect 44582 681272 45480 681274
rect 43790 681270 43922 681272
rect 43790 681170 43810 681270
rect 43910 681238 43922 681270
rect 44090 681238 44180 681272
rect 44348 681238 44420 681272
rect 44606 681270 44696 681272
rect 44670 681238 44696 681270
rect 44864 681238 44954 681272
rect 45122 681238 45212 681272
rect 45380 681270 45480 681272
rect 43910 681234 44420 681238
rect 44582 681234 44600 681238
rect 43910 681230 44600 681234
rect 43910 681170 43930 681230
rect 44408 681228 44600 681230
rect 44590 681200 44600 681228
rect 44670 681230 45360 681238
rect 44670 681200 44680 681230
rect 43790 681160 43930 681170
rect 45340 681170 45360 681230
rect 45460 681170 45480 681270
rect 541004 681270 548204 681318
rect 541004 681236 541025 681270
rect 542001 681258 542261 681270
rect 542001 681236 542024 681258
rect 45340 681160 45480 681170
rect 540926 681208 540972 681220
rect 541004 681218 542024 681236
rect 542244 681236 542261 681258
rect 543237 681258 543497 681270
rect 543237 681236 543249 681258
rect 542244 681230 543249 681236
rect 543484 681236 543497 681258
rect 544473 681258 544733 681270
rect 544473 681236 544485 681258
rect 543484 681230 544485 681236
rect 544721 681236 544733 681258
rect 545709 681258 545969 681270
rect 545709 681236 545724 681258
rect 544721 681230 545724 681236
rect 540926 681040 540932 681208
rect 540966 681168 540972 681208
rect 542054 681208 542100 681220
rect 542054 681168 542060 681208
rect 540966 681040 542060 681168
rect 542094 681168 542100 681208
rect 542162 681208 542208 681220
rect 542244 681218 543244 681230
rect 542162 681168 542168 681208
rect 542094 681040 542168 681168
rect 542202 681168 542208 681208
rect 543290 681208 543336 681220
rect 543290 681168 543296 681208
rect 542202 681158 543296 681168
rect 542202 681088 542884 681158
rect 542954 681088 543104 681158
rect 543174 681088 543296 681158
rect 542202 681040 543296 681088
rect 543330 681168 543336 681208
rect 543398 681208 543444 681220
rect 543484 681218 544484 681230
rect 543398 681168 543404 681208
rect 543330 681040 543404 681168
rect 543438 681168 543444 681208
rect 544526 681208 544572 681220
rect 544526 681168 544532 681208
rect 543438 681040 544532 681168
rect 544566 681168 544572 681208
rect 544634 681208 544680 681220
rect 544724 681218 545724 681230
rect 545944 681236 545969 681258
rect 546945 681258 547205 681270
rect 546945 681236 546964 681258
rect 544634 681168 544640 681208
rect 544566 681040 544640 681168
rect 544674 681168 544680 681208
rect 545762 681208 545808 681220
rect 545762 681168 545768 681208
rect 544674 681040 545768 681168
rect 545802 681168 545808 681208
rect 545870 681208 545916 681220
rect 545944 681218 546964 681236
rect 547184 681236 547205 681258
rect 548181 681236 548204 681270
rect 545870 681168 545876 681208
rect 545802 681040 545876 681168
rect 545910 681168 545916 681208
rect 546998 681208 547044 681220
rect 546998 681168 547004 681208
rect 545910 681158 547004 681168
rect 545910 681088 546064 681158
rect 546134 681088 546304 681158
rect 546374 681088 547004 681158
rect 545910 681040 547004 681088
rect 547038 681168 547044 681208
rect 547106 681208 547152 681220
rect 547184 681218 548204 681236
rect 554420 681400 563740 681600
rect 547106 681168 547112 681208
rect 547038 681040 547112 681168
rect 547146 681168 547152 681208
rect 548234 681208 548280 681220
rect 548234 681168 548240 681208
rect 547146 681040 548240 681168
rect 548274 681040 548280 681208
rect 540926 681028 548280 681040
rect 554420 681200 561700 681400
rect 561900 681200 562100 681400
rect 562300 681200 562500 681400
rect 562700 681200 562900 681400
rect 563100 681200 563300 681400
rect 563500 681200 563740 681400
rect 540926 681012 548274 681028
rect 540926 680978 541025 681012
rect 542001 680978 542261 681012
rect 543237 680978 543497 681012
rect 544473 680978 544733 681012
rect 545709 680978 545969 681012
rect 546945 680978 547205 681012
rect 548181 680978 548274 681012
rect 540926 680956 548274 680978
rect 554420 681000 563740 681200
rect 541372 680898 541556 680904
rect 542432 680898 542616 680904
rect 543892 680898 544076 680904
rect 545112 680898 545296 680904
rect 546592 680898 546776 680904
rect 547592 680898 547776 680904
rect 44590 680790 44600 680830
rect 44450 680782 44600 680790
rect 44450 680748 44522 680782
rect 44590 680760 44600 680782
rect 44670 680790 44680 680830
rect 44670 680782 44820 680790
rect 44670 680760 44680 680782
rect 44590 680748 44680 680760
rect 44748 680748 44820 680782
rect 44450 680740 44820 680748
rect 44450 680698 44500 680740
rect 44334 680580 44386 680592
rect 44334 680520 44340 680580
rect 44380 680520 44386 680580
rect 44450 680550 44460 680698
rect 44260 680400 44270 680520
rect 44390 680400 44400 680520
rect 44334 680350 44340 680400
rect 44380 680350 44386 680400
rect 44334 680338 44386 680350
rect 44454 680222 44460 680550
rect 44494 680222 44500 680698
rect 44612 680698 44658 680710
rect 44612 680360 44618 680698
rect 44652 680360 44658 680698
rect 44770 680698 44820 680740
rect 44590 680290 44600 680360
rect 44670 680290 44680 680360
rect 44454 680220 44500 680222
rect 44450 680180 44500 680220
rect 44612 680222 44618 680290
rect 44652 680222 44658 680290
rect 44612 680210 44658 680222
rect 44770 680222 44776 680698
rect 44810 680550 44820 680698
rect 541004 680738 541384 680898
rect 541544 680738 542444 680898
rect 542604 680738 543904 680898
rect 544064 680738 545124 680898
rect 545284 680738 546604 680898
rect 546764 680738 547604 680898
rect 547764 680738 548204 680898
rect 541004 680680 548204 680738
rect 541004 680658 541025 680680
rect 541013 680646 541025 680658
rect 542001 680668 542261 680680
rect 542001 680646 542013 680668
rect 541013 680640 542013 680646
rect 542249 680646 542261 680668
rect 543237 680668 543497 680680
rect 543237 680646 543249 680668
rect 542249 680640 543249 680646
rect 543485 680646 543497 680668
rect 544473 680668 544733 680680
rect 544473 680646 544485 680668
rect 543485 680640 544485 680646
rect 544721 680646 544733 680668
rect 545709 680668 545969 680680
rect 545709 680646 545721 680668
rect 544721 680640 545721 680646
rect 545957 680646 545969 680668
rect 546945 680668 547205 680680
rect 546945 680646 546957 680668
rect 545957 680640 546957 680646
rect 547193 680646 547205 680668
rect 548181 680658 548204 680680
rect 554420 680800 561700 681000
rect 561900 680800 562100 681000
rect 562300 680800 562500 681000
rect 562700 680800 562900 681000
rect 563100 680800 563300 681000
rect 563500 680800 563740 681000
rect 548181 680646 548193 680658
rect 547193 680640 548193 680646
rect 540926 680618 540972 680630
rect 44884 680580 44936 680592
rect 44810 680222 44816 680550
rect 44884 680530 44890 680580
rect 44930 680530 44936 680580
rect 540926 680578 540932 680618
rect 44880 680410 44890 680530
rect 45010 680410 45020 680530
rect 540924 680488 540932 680578
rect 540926 680450 540932 680488
rect 540966 680578 540972 680618
rect 542054 680618 542100 680630
rect 542054 680578 542060 680618
rect 540966 680488 542060 680578
rect 540966 680450 540972 680488
rect 540926 680438 540972 680450
rect 542054 680450 542060 680488
rect 542094 680578 542100 680618
rect 542162 680618 542208 680630
rect 542162 680578 542168 680618
rect 542094 680488 542168 680578
rect 542094 680450 542100 680488
rect 542054 680438 542100 680450
rect 542162 680450 542168 680488
rect 542202 680578 542208 680618
rect 543290 680618 543336 680630
rect 543290 680578 543296 680618
rect 542202 680568 543296 680578
rect 542202 680498 542884 680568
rect 542954 680498 543104 680568
rect 543174 680498 543296 680568
rect 542202 680488 543296 680498
rect 542202 680450 542208 680488
rect 542162 680438 542208 680450
rect 543290 680450 543296 680488
rect 543330 680578 543336 680618
rect 543398 680618 543444 680630
rect 543398 680578 543404 680618
rect 543330 680488 543404 680578
rect 543330 680450 543336 680488
rect 543290 680438 543336 680450
rect 543398 680450 543404 680488
rect 543438 680578 543444 680618
rect 544526 680618 544572 680630
rect 544526 680578 544532 680618
rect 543438 680488 544532 680578
rect 543438 680450 543444 680488
rect 543398 680438 543444 680450
rect 544526 680450 544532 680488
rect 544566 680578 544572 680618
rect 544634 680618 544680 680630
rect 544634 680578 544640 680618
rect 544566 680488 544640 680578
rect 544566 680450 544572 680488
rect 544526 680438 544572 680450
rect 544634 680450 544640 680488
rect 544674 680578 544680 680618
rect 545762 680618 545808 680630
rect 545762 680578 545768 680618
rect 544674 680488 545768 680578
rect 544674 680450 544680 680488
rect 544634 680438 544680 680450
rect 545762 680450 545768 680488
rect 545802 680578 545808 680618
rect 545870 680618 545916 680630
rect 545870 680578 545876 680618
rect 545802 680488 545876 680578
rect 545802 680450 545808 680488
rect 545762 680438 545808 680450
rect 545870 680450 545876 680488
rect 545910 680578 545916 680618
rect 546998 680618 547044 680630
rect 546998 680578 547004 680618
rect 545910 680568 547004 680578
rect 545910 680498 546064 680568
rect 546134 680498 546304 680568
rect 546374 680498 547004 680568
rect 545910 680488 547004 680498
rect 545910 680450 545916 680488
rect 545870 680438 545916 680450
rect 546998 680450 547004 680488
rect 547038 680578 547044 680618
rect 547106 680618 547152 680630
rect 547106 680578 547112 680618
rect 547038 680488 547112 680578
rect 547038 680450 547044 680488
rect 546998 680438 547044 680450
rect 547106 680450 547112 680488
rect 547146 680578 547152 680618
rect 548234 680618 548280 680630
rect 548234 680578 548240 680618
rect 547146 680488 548240 680578
rect 547146 680450 547152 680488
rect 547106 680438 547152 680450
rect 548234 680450 548240 680488
rect 548274 680450 548280 680618
rect 548234 680438 548280 680450
rect 554420 680600 563740 680800
rect 541004 680422 542013 680428
rect 44884 680350 44890 680410
rect 44930 680350 44936 680410
rect 44884 680338 44936 680350
rect 541004 680388 541025 680422
rect 542001 680408 542013 680422
rect 542249 680422 543249 680428
rect 542249 680408 542261 680422
rect 542001 680388 542261 680408
rect 543237 680408 543249 680422
rect 543485 680422 544485 680428
rect 543485 680408 543497 680422
rect 544473 680408 544485 680422
rect 544721 680422 545721 680428
rect 544721 680408 544733 680422
rect 545709 680408 545721 680422
rect 545957 680422 546957 680428
rect 545957 680408 545969 680422
rect 543237 680388 543497 680408
rect 544473 680388 544733 680408
rect 545709 680388 545969 680408
rect 546945 680408 546957 680422
rect 547193 680422 548198 680428
rect 547193 680408 547205 680422
rect 546945 680388 547205 680408
rect 548181 680388 548198 680422
rect 541004 680338 544044 680388
rect 544114 680338 544154 680388
rect 544224 680338 544984 680388
rect 545054 680338 545094 680388
rect 545164 680338 548198 680388
rect 541004 680328 548198 680338
rect 554420 680400 561700 680600
rect 561900 680400 562100 680600
rect 562300 680400 562500 680600
rect 562700 680400 562900 680600
rect 563100 680400 563300 680600
rect 563500 680400 563740 680600
rect 44770 680220 44816 680222
rect 44770 680180 44820 680220
rect 44450 680172 44820 680180
rect 44450 680138 44522 680172
rect 44590 680138 44680 680172
rect 44748 680138 44820 680172
rect 44450 680130 44820 680138
rect 554420 680200 563740 680400
rect 554420 680000 561700 680200
rect 561900 680000 562100 680200
rect 562300 680000 562500 680200
rect 562700 680000 562900 680200
rect 563100 680000 563300 680200
rect 563500 680000 563740 680200
rect 544400 679918 544410 679926
rect 543684 679890 544410 679918
rect 544470 679890 544510 679926
rect 543684 679856 543786 679890
rect 544012 679856 544254 679890
rect 544480 679866 544510 679890
rect 544570 679866 544610 679926
rect 544670 679866 544710 679926
rect 544770 679918 544780 679926
rect 544770 679890 545504 679918
rect 544480 679856 544722 679866
rect 544948 679856 545190 679890
rect 545416 679856 545504 679890
rect 543684 679848 545504 679856
rect 543684 679838 544984 679848
rect 44080 679750 44090 679830
rect 44170 679790 44180 679830
rect 44590 679790 44600 679830
rect 44170 679782 44600 679790
rect 44080 679748 44162 679750
rect 44330 679748 44420 679782
rect 44588 679760 44600 679782
rect 44670 679790 44680 679830
rect 45120 679790 45130 679830
rect 44670 679782 45130 679790
rect 44670 679760 44678 679782
rect 44588 679748 44678 679760
rect 44846 679748 44936 679782
rect 45104 679750 45130 679782
rect 45210 679750 45220 679830
rect 543684 679828 544044 679838
rect 543684 679768 543702 679828
rect 45104 679748 45220 679750
rect 44080 679740 45220 679748
rect 44094 679698 44140 679710
rect 44350 679700 44400 679740
rect 44870 679710 44920 679740
rect 44094 679640 44100 679698
rect 43940 679630 44100 679640
rect 44134 679640 44140 679698
rect 44352 679698 44398 679700
rect 44134 679630 44170 679640
rect 43940 679540 43960 679630
rect 44050 679540 44070 679630
rect 44160 679540 44170 679630
rect 43940 679530 44100 679540
rect 44094 679472 44100 679530
rect 44134 679530 44170 679540
rect 44134 679472 44140 679530
rect 44094 679460 44140 679472
rect 44352 679472 44358 679698
rect 44392 679472 44398 679698
rect 44610 679698 44656 679710
rect 44610 679630 44616 679698
rect 44650 679630 44656 679698
rect 44868 679698 44914 679710
rect 44580 679540 44590 679630
rect 44680 679540 44690 679630
rect 44352 679470 44398 679472
rect 44610 679472 44616 679540
rect 44650 679472 44656 679540
rect 44350 679430 44400 679470
rect 44610 679460 44656 679472
rect 44868 679472 44874 679698
rect 44908 679472 44914 679698
rect 45126 679698 45172 679710
rect 45126 679630 45132 679698
rect 45166 679640 45172 679698
rect 543696 679660 543702 679768
rect 543736 679768 544044 679828
rect 544114 679768 544154 679838
rect 544224 679828 544984 679838
rect 544224 679768 544530 679828
rect 543736 679688 544062 679768
rect 543736 679660 543742 679688
rect 543696 679648 543742 679660
rect 544054 679660 544062 679688
rect 544096 679660 544170 679768
rect 544204 679688 544530 679768
rect 544204 679660 544214 679688
rect 544054 679648 544214 679660
rect 544524 679660 544530 679688
rect 544564 679660 544638 679828
rect 544672 679778 544984 679828
rect 545054 679778 545094 679848
rect 545164 679840 545504 679848
rect 545164 679828 545506 679840
rect 545164 679778 545466 679828
rect 544672 679688 544998 679778
rect 544672 679660 544679 679688
rect 544524 679648 544679 679660
rect 544992 679660 544998 679688
rect 545032 679660 545106 679778
rect 545140 679688 545466 679778
rect 545140 679660 545149 679688
rect 544992 679648 545149 679660
rect 545460 679660 545466 679688
rect 545500 679660 545506 679828
rect 545460 679648 545506 679660
rect 554420 679800 563740 680000
rect 45166 679630 45320 679640
rect 45090 679540 45100 679630
rect 45190 679550 45220 679630
rect 45300 679550 45320 679630
rect 543774 679632 544024 679638
rect 543774 679618 543786 679632
rect 45190 679540 45320 679550
rect 543764 679598 543786 679618
rect 544012 679618 544024 679632
rect 544242 679632 544492 679638
rect 544242 679618 544254 679632
rect 544012 679598 544254 679618
rect 544480 679618 544492 679632
rect 544710 679632 544960 679638
rect 544710 679618 544722 679632
rect 544480 679598 544722 679618
rect 544948 679618 544960 679632
rect 545178 679632 545428 679638
rect 545178 679618 545190 679632
rect 544948 679598 545190 679618
rect 545416 679618 545428 679632
rect 545416 679598 545434 679618
rect 543764 679578 545434 679598
rect 554420 679600 561700 679800
rect 561900 679600 562100 679800
rect 562300 679600 562500 679800
rect 562700 679600 562900 679800
rect 563100 679600 563300 679800
rect 563500 679600 563740 679800
rect 44868 679470 44914 679472
rect 45126 679472 45132 679540
rect 45166 679472 45172 679540
rect 543764 679524 545474 679578
rect 44868 679460 44920 679470
rect 45126 679460 45172 679472
rect 543752 679518 545486 679524
rect 44870 679430 44920 679460
rect 44140 679422 45120 679430
rect 44140 679388 44162 679422
rect 44330 679388 44420 679422
rect 44588 679388 44678 679422
rect 44846 679388 44936 679422
rect 45104 679388 45120 679422
rect 44140 679380 44220 679388
rect 44210 679360 44220 679380
rect 44280 679380 44990 679388
rect 44280 679360 44290 679380
rect 44980 679360 44990 679380
rect 45050 679380 45120 679388
rect 45050 679360 45060 679380
rect 543752 679368 543764 679518
rect 543984 679508 544284 679518
rect 543984 679368 543996 679508
rect 543752 679362 543996 679368
rect 544272 679368 544284 679508
rect 544504 679508 544704 679518
rect 544504 679368 544516 679508
rect 544272 679362 544516 679368
rect 544692 679368 544704 679508
rect 544924 679508 545254 679518
rect 544924 679368 544936 679508
rect 544692 679362 544936 679368
rect 545242 679368 545254 679508
rect 545474 679368 545486 679518
rect 545242 679362 545486 679368
rect 554420 679400 563740 679600
rect 44480 679320 44760 679330
rect 546044 679328 546394 679348
rect 44480 679280 44500 679320
rect 44740 679280 44760 679320
rect 44480 679250 44760 679280
rect 44480 679160 44580 679250
rect 44670 679160 44760 679250
rect 44480 679140 44760 679160
rect 44480 679100 44500 679140
rect 44740 679100 44760 679140
rect 542864 679308 546064 679328
rect 542864 679238 542884 679308
rect 542954 679238 543094 679308
rect 543164 679265 546064 679308
rect 543164 679238 544006 679265
rect 542864 679231 544006 679238
rect 544482 679231 544724 679265
rect 545200 679258 546064 679265
rect 546134 679258 546304 679328
rect 546374 679258 546394 679328
rect 545200 679238 546394 679258
rect 545200 679231 546064 679238
rect 542864 679218 546064 679231
rect 542864 679148 542884 679218
rect 542954 679148 543094 679218
rect 543164 679203 546064 679218
rect 543164 679148 543922 679203
rect 542864 679118 543194 679148
rect 543916 679135 543922 679148
rect 543956 679148 544532 679203
rect 543956 679135 543962 679148
rect 543916 679123 543962 679135
rect 544526 679135 544532 679148
rect 544566 679148 544640 679203
rect 544566 679135 544572 679148
rect 544526 679123 544572 679135
rect 544634 679135 544640 679148
rect 544674 679148 545250 679203
rect 544674 679135 544680 679148
rect 544634 679123 544680 679135
rect 545244 679135 545250 679148
rect 545284 679168 546064 679203
rect 546134 679168 546304 679238
rect 546374 679168 546394 679238
rect 545284 679148 546394 679168
rect 554420 679200 561700 679400
rect 561900 679200 562100 679400
rect 562300 679200 562500 679400
rect 562700 679200 562900 679400
rect 563100 679200 563300 679400
rect 563500 679200 563740 679400
rect 545284 679135 545290 679148
rect 545244 679123 545290 679135
rect 44480 679090 44760 679100
rect 543994 679107 544494 679113
rect 543994 679093 544006 679107
rect 543989 679078 544006 679093
rect 544482 679093 544494 679107
rect 544712 679107 545212 679113
rect 544712 679093 544724 679107
rect 543984 679073 544006 679078
rect 544482 679073 544724 679093
rect 545200 679093 545212 679107
rect 545200 679078 545224 679093
rect 545200 679073 545234 679078
rect 44210 679040 44220 679060
rect 43720 679032 44220 679040
rect 44280 679040 44290 679060
rect 44980 679040 44990 679060
rect 44280 679032 44990 679040
rect 45050 679040 45060 679060
rect 45050 679032 45550 679040
rect 43720 678998 43907 679032
rect 44075 678998 44165 679032
rect 44333 678998 44423 679032
rect 44591 678998 44681 679032
rect 44849 678998 44939 679032
rect 45107 678998 45197 679032
rect 45365 678998 45550 679032
rect 543984 679018 544044 679073
rect 544114 679018 544154 679073
rect 544224 679018 544984 679073
rect 545054 679018 545094 679073
rect 545164 679018 545234 679073
rect 543984 679008 545234 679018
rect 43720 678990 45550 678998
rect 43720 677930 43780 678990
rect 43839 678948 43885 678960
rect 43839 678690 43845 678948
rect 43879 678690 43885 678948
rect 44097 678948 44143 678960
rect 43820 678630 43830 678690
rect 43890 678630 43900 678690
rect 43839 677972 43845 678630
rect 43879 677972 43885 678630
rect 44097 678280 44103 678948
rect 44137 678280 44143 678948
rect 44355 678948 44401 678960
rect 44355 678690 44361 678948
rect 44395 678690 44401 678948
rect 44613 678948 44659 678960
rect 44340 678630 44350 678690
rect 44410 678630 44420 678690
rect 44080 678220 44090 678280
rect 44150 678220 44160 678280
rect 43839 677960 43885 677972
rect 44097 677972 44103 678220
rect 44137 677972 44143 678220
rect 44097 677960 44143 677972
rect 44355 677972 44361 678630
rect 44395 677972 44401 678630
rect 44613 678280 44619 678948
rect 44653 678280 44659 678948
rect 44871 678948 44917 678960
rect 44871 678720 44877 678948
rect 44911 678720 44917 678948
rect 45129 678948 45175 678960
rect 44820 678610 44830 678720
rect 44960 678610 44970 678720
rect 44600 678220 44610 678280
rect 44670 678220 44680 678280
rect 44355 677960 44401 677972
rect 44613 677972 44619 678220
rect 44653 677972 44659 678220
rect 44613 677960 44659 677972
rect 44871 677972 44877 678610
rect 44911 677972 44917 678610
rect 45129 678280 45135 678948
rect 45169 678280 45175 678948
rect 45387 678948 45433 678960
rect 45387 678690 45393 678948
rect 45427 678690 45433 678948
rect 45370 678630 45380 678690
rect 45440 678630 45450 678690
rect 45110 678220 45120 678280
rect 45180 678220 45190 678280
rect 44871 677960 44917 677972
rect 45129 677972 45135 678220
rect 45169 677972 45175 678220
rect 45129 677960 45175 677972
rect 45387 677972 45393 678630
rect 45427 677972 45433 678630
rect 45387 677960 45433 677972
rect 45490 677930 45550 678990
rect 554420 679000 563740 679200
rect 543512 678968 543716 678974
rect 541392 678958 541596 678964
rect 541392 678828 541404 678958
rect 541584 678828 541596 678958
rect 541392 678822 541596 678828
rect 542532 678958 542736 678964
rect 542532 678828 542544 678958
rect 542724 678828 542736 678958
rect 543512 678838 543524 678968
rect 543704 678838 543716 678968
rect 543512 678832 543716 678838
rect 544282 678968 544486 678974
rect 544282 678838 544294 678968
rect 544474 678838 544486 678968
rect 544282 678832 544486 678838
rect 544722 678968 544926 678974
rect 544722 678838 544734 678968
rect 544914 678838 544926 678968
rect 546512 678968 546716 678974
rect 544722 678832 544926 678838
rect 545442 678958 545646 678964
rect 542532 678822 542736 678828
rect 545442 678828 545454 678958
rect 545634 678828 545646 678958
rect 546512 678838 546524 678968
rect 546704 678838 546716 678968
rect 546512 678832 546716 678838
rect 547512 678968 547716 678974
rect 547512 678838 547524 678968
rect 547704 678838 547716 678968
rect 547512 678832 547716 678838
rect 545442 678822 545646 678828
rect 554420 678800 561700 679000
rect 561900 678800 562100 679000
rect 562300 678800 562500 679000
rect 562700 678800 562900 679000
rect 563100 678800 563300 679000
rect 563500 678800 563740 679000
rect 541054 678788 548144 678793
rect 541054 678740 542884 678788
rect 542954 678740 543104 678788
rect 543174 678740 546064 678788
rect 546134 678740 546304 678788
rect 546374 678746 548144 678788
rect 546374 678740 548149 678746
rect 541054 678718 541071 678740
rect 541059 678706 541071 678718
rect 542047 678718 542289 678740
rect 543265 678718 543507 678740
rect 542047 678706 542059 678718
rect 541059 678700 542059 678706
rect 542277 678706 542289 678718
rect 543265 678706 543277 678718
rect 542277 678700 543277 678706
rect 543495 678706 543507 678718
rect 544483 678718 544725 678740
rect 544483 678706 544495 678718
rect 543495 678700 544495 678706
rect 544713 678706 544725 678718
rect 545701 678718 545943 678740
rect 546919 678718 547161 678740
rect 545701 678706 545713 678718
rect 544713 678700 545713 678706
rect 545931 678706 545943 678718
rect 546919 678706 546931 678718
rect 545931 678700 546931 678706
rect 547149 678706 547161 678718
rect 548137 678706 548149 678740
rect 547149 678700 548149 678706
rect 540981 678678 541027 678690
rect 540981 678510 540987 678678
rect 541021 678643 541027 678678
rect 542091 678678 542137 678690
rect 542091 678643 542097 678678
rect 541021 678558 542097 678643
rect 541021 678510 541027 678558
rect 540981 678498 541027 678510
rect 542091 678510 542097 678558
rect 542131 678643 542137 678678
rect 542199 678678 542245 678690
rect 542199 678643 542205 678678
rect 542131 678558 542205 678643
rect 542131 678510 542137 678558
rect 542091 678498 542137 678510
rect 542199 678510 542205 678558
rect 542239 678643 542245 678678
rect 543309 678678 543355 678690
rect 543309 678643 543315 678678
rect 542239 678558 543315 678643
rect 542239 678510 542245 678558
rect 542199 678498 542245 678510
rect 543309 678510 543315 678558
rect 543349 678643 543355 678678
rect 543417 678678 543463 678690
rect 543417 678643 543423 678678
rect 543349 678558 543423 678643
rect 543349 678510 543355 678558
rect 543309 678498 543355 678510
rect 543417 678510 543423 678558
rect 543457 678643 543463 678678
rect 544527 678678 544573 678690
rect 544527 678643 544533 678678
rect 543457 678638 544533 678643
rect 543457 678568 544044 678638
rect 544114 678568 544154 678638
rect 544224 678568 544533 678638
rect 543457 678558 544533 678568
rect 543457 678510 543463 678558
rect 543417 678498 543463 678510
rect 544527 678510 544533 678558
rect 544567 678643 544573 678678
rect 544635 678678 544681 678690
rect 544635 678643 544641 678678
rect 544567 678558 544641 678643
rect 544567 678510 544573 678558
rect 544527 678498 544573 678510
rect 544635 678510 544641 678558
rect 544675 678643 544681 678678
rect 545745 678678 545791 678690
rect 545745 678643 545751 678678
rect 544675 678638 545751 678643
rect 544675 678568 544984 678638
rect 545054 678568 545094 678638
rect 545164 678568 545751 678638
rect 544675 678558 545751 678568
rect 544675 678510 544681 678558
rect 544635 678498 544681 678510
rect 545745 678510 545751 678558
rect 545785 678643 545791 678678
rect 545853 678678 545899 678690
rect 545853 678643 545859 678678
rect 545785 678558 545859 678643
rect 545785 678510 545791 678558
rect 545745 678498 545791 678510
rect 545853 678510 545859 678558
rect 545893 678643 545899 678678
rect 546963 678678 547009 678690
rect 546963 678643 546969 678678
rect 545893 678558 546969 678643
rect 545893 678510 545899 678558
rect 545853 678498 545899 678510
rect 546963 678510 546969 678558
rect 547003 678643 547009 678678
rect 547071 678678 547117 678690
rect 547071 678643 547077 678678
rect 547003 678558 547077 678643
rect 547003 678510 547009 678558
rect 546963 678498 547009 678510
rect 547071 678510 547077 678558
rect 547111 678643 547117 678678
rect 548181 678678 548227 678690
rect 548181 678643 548187 678678
rect 547111 678558 548187 678643
rect 547111 678510 547117 678558
rect 547071 678498 547117 678510
rect 548181 678510 548187 678558
rect 548221 678510 548227 678678
rect 548181 678498 548227 678510
rect 554420 678600 563740 678800
rect 541059 678482 542059 678488
rect 541059 678468 541071 678482
rect 541054 678448 541071 678468
rect 542047 678468 542059 678482
rect 542277 678482 543277 678488
rect 542277 678468 542289 678482
rect 542047 678448 542289 678468
rect 543265 678468 543277 678482
rect 543495 678482 544495 678488
rect 543495 678468 543507 678482
rect 543265 678448 543507 678468
rect 544483 678468 544495 678482
rect 544713 678482 545713 678488
rect 544713 678468 544725 678482
rect 544483 678448 544725 678468
rect 545701 678468 545713 678482
rect 545931 678482 546931 678488
rect 545931 678468 545943 678482
rect 545701 678448 545943 678468
rect 546919 678468 546931 678482
rect 547149 678482 548149 678488
rect 547149 678468 547161 678482
rect 546919 678448 547161 678468
rect 548137 678448 548149 678482
rect 541054 678442 548149 678448
rect 541054 678393 548144 678442
rect 554420 678400 561700 678600
rect 561900 678400 562100 678600
rect 562300 678400 562500 678600
rect 562700 678400 562900 678600
rect 563100 678400 563300 678600
rect 563500 678400 563740 678600
rect 542404 678098 542804 678393
rect 543804 678098 544204 678393
rect 545104 678098 545504 678393
rect 546394 678098 546804 678393
rect 554420 678340 563740 678400
rect 43720 677922 45550 677930
rect 43720 677888 43907 677922
rect 44075 677888 44165 677922
rect 44333 677888 44423 677922
rect 44591 677888 44681 677922
rect 44849 677888 44939 677922
rect 45107 677888 45197 677922
rect 45365 677888 45550 677922
rect 43720 677880 45550 677888
rect 541604 677990 547604 678098
rect 541604 677984 544807 677990
rect 44480 677820 44760 677830
rect 44480 677780 44500 677820
rect 44740 677780 44760 677820
rect 44480 677720 44580 677780
rect 44670 677720 44760 677780
rect 44480 677710 44760 677720
rect 541604 677587 541777 677984
rect 542891 677587 543297 677984
rect 544411 677593 544807 677984
rect 545921 677593 546317 677990
rect 547431 677593 547604 677990
rect 544411 677587 547604 677593
rect 42590 677532 46960 677550
rect 41726 677530 47504 677532
rect 41726 677526 44090 677530
rect 44150 677526 45120 677530
rect 45180 677526 47504 677530
rect 41726 677129 41738 677526
rect 42852 677129 43288 677526
rect 44402 677129 44828 677526
rect 45942 677129 46378 677526
rect 47492 677129 47504 677526
rect 541604 677498 547604 677587
rect 41726 677123 47504 677129
rect 42590 677110 46960 677123
rect 541352 677058 541496 677064
rect 41188 676980 41452 676986
rect 41188 676740 41200 676980
rect 41440 676740 41452 676980
rect 41188 676734 41452 676740
rect 47888 676980 48152 676986
rect 47888 676740 47900 676980
rect 48140 676740 48152 676980
rect 541352 676938 541364 677058
rect 541484 676938 541496 677058
rect 541352 676932 541496 676938
rect 547722 677058 547866 677064
rect 547722 676938 547734 677058
rect 547854 676938 547866 677058
rect 547722 676932 547866 676938
rect 47888 676734 48152 676740
rect 41188 675260 41452 675266
rect 41188 675020 41200 675260
rect 41440 675020 41452 675260
rect 41188 675014 41452 675020
rect 47888 675260 48152 675266
rect 47888 675020 47900 675260
rect 48140 675020 48152 675260
rect 47888 675014 48152 675020
rect 541352 674058 541496 674064
rect 541352 673938 541364 674058
rect 541484 673938 541496 674058
rect 541352 673932 541496 673938
rect 547722 674058 547866 674064
rect 547722 673938 547734 674058
rect 547854 673938 547866 674058
rect 547722 673932 547866 673938
rect 41188 673540 41452 673546
rect 41188 673300 41200 673540
rect 41440 673300 41452 673540
rect 41188 673294 41452 673300
rect 47888 673540 48152 673546
rect 47888 673300 47900 673540
rect 48140 673300 48152 673540
rect 47888 673294 48152 673300
rect 41188 672060 41452 672066
rect 41188 671820 41200 672060
rect 41440 671820 41452 672060
rect 41188 671814 41452 671820
rect 47888 672060 48152 672066
rect 47888 671820 47900 672060
rect 48140 671820 48152 672060
rect 47888 671814 48152 671820
rect 541352 671058 541496 671064
rect 541352 670938 541364 671058
rect 541484 670938 541496 671058
rect 541352 670932 541496 670938
rect 547722 671058 547866 671064
rect 547722 670938 547734 671058
rect 547854 670938 547866 671058
rect 547722 670932 547866 670938
rect 41188 670340 41452 670346
rect 41188 670100 41200 670340
rect 41440 670100 41452 670340
rect 41188 670094 41452 670100
rect 47888 670340 48152 670346
rect 47888 670100 47900 670340
rect 48140 670100 48152 670340
rect 47888 670094 48152 670100
rect 41188 668740 41452 668746
rect 41188 668500 41200 668740
rect 41440 668500 41452 668740
rect 41188 668494 41452 668500
rect 47888 668740 48152 668746
rect 47888 668500 47900 668740
rect 48140 668500 48152 668740
rect 47888 668494 48152 668500
rect 541352 668058 541496 668064
rect 541352 667938 541364 668058
rect 541484 667938 541496 668058
rect 541352 667932 541496 667938
rect 547722 668058 547866 668064
rect 547722 667938 547734 668058
rect 547854 667938 547866 668058
rect 547722 667932 547866 667938
rect 41188 667020 41452 667026
rect 41188 666780 41200 667020
rect 41440 666780 41452 667020
rect 41188 666774 41452 666780
rect 47888 667020 48152 667026
rect 47888 666780 47900 667020
rect 48140 666780 48152 667020
rect 47888 666774 48152 666780
rect 41188 665420 41452 665426
rect 41188 665180 41200 665420
rect 41440 665180 41452 665420
rect 41188 665174 41452 665180
rect 47888 665420 48152 665426
rect 47888 665180 47900 665420
rect 48140 665180 48152 665420
rect 47888 665174 48152 665180
rect 541352 665058 541496 665064
rect 541352 664938 541364 665058
rect 541484 664938 541496 665058
rect 541352 664932 541496 664938
rect 547722 665058 547866 665064
rect 547722 664938 547734 665058
rect 547854 664938 547866 665058
rect 547722 664932 547866 664938
rect 541604 663759 547604 663798
rect 541604 663753 544807 663759
rect 541604 663728 541777 663753
rect 542891 663728 543297 663753
rect 544411 663728 544807 663753
rect 545921 663738 546317 663759
rect 547431 663738 547604 663759
rect 545921 663728 546294 663738
rect 41188 663700 41452 663706
rect 41188 663460 41200 663700
rect 41440 663460 41452 663700
rect 41188 663454 41452 663460
rect 47888 663700 48152 663706
rect 47888 663460 47900 663700
rect 48140 663460 48152 663700
rect 47888 663454 48152 663460
rect 32600 663300 48300 663400
rect 32600 663000 32800 663300
rect 33100 663000 33300 663300
rect 33600 663000 33800 663300
rect 34100 663000 34300 663300
rect 34600 663000 34800 663300
rect 35100 663000 35300 663300
rect 35600 663000 35800 663300
rect 36100 663000 36300 663300
rect 36600 663000 36800 663300
rect 37100 663000 37300 663300
rect 37600 663000 37800 663300
rect 38100 663000 38300 663300
rect 38600 663000 38800 663300
rect 39100 663000 39300 663300
rect 39600 663000 39800 663300
rect 40100 663000 40300 663300
rect 40600 663295 48300 663300
rect 541604 663318 541744 663728
rect 542914 663318 543254 663728
rect 544424 663318 544774 663728
rect 545944 663328 546294 663728
rect 547464 663328 547604 663738
rect 545944 663318 547604 663328
rect 541604 663298 547604 663318
rect 40600 663220 41738 663295
rect 40600 663000 41200 663220
rect 32600 662980 41200 663000
rect 41440 662980 41738 663220
rect 32600 662898 41738 662980
rect 42852 662898 43288 663295
rect 44402 662898 44828 663295
rect 45942 662898 46378 663295
rect 47492 663220 48300 663295
rect 47492 662980 47900 663220
rect 48140 662980 48300 663220
rect 47492 662898 48300 662980
rect 32600 662800 48300 662898
<< via1 >>
rect 36930 694850 37000 694920
rect 36820 694740 36890 694810
rect 44010 695382 44280 695640
rect 45060 695382 45330 695640
rect 44010 695370 44280 695382
rect 45060 695370 45330 695382
rect 41460 695090 41480 695160
rect 41480 695090 41514 695160
rect 41514 695090 41530 695160
rect 41460 694850 41480 694920
rect 41480 694850 41514 694920
rect 41514 694850 41530 694920
rect 41780 695090 41796 695160
rect 41796 695090 41830 695160
rect 41830 695090 41850 695160
rect 41780 694850 41796 694920
rect 41796 694850 41830 694920
rect 41830 694850 41850 694920
rect 41620 694480 41638 694550
rect 41638 694480 41672 694550
rect 41672 694480 41690 694550
rect 41620 694240 41638 694310
rect 41638 694240 41672 694310
rect 41672 694240 41690 694310
rect 42090 695090 42112 695160
rect 42112 695090 42146 695160
rect 42146 695090 42160 695160
rect 42090 694850 42112 694920
rect 42112 694850 42146 694920
rect 42146 694850 42160 694920
rect 41930 694480 41954 694550
rect 41954 694480 41988 694550
rect 41988 694480 42000 694550
rect 41930 694240 41954 694310
rect 41954 694240 41988 694310
rect 41988 694240 42000 694310
rect 42410 695090 42428 695160
rect 42428 695090 42462 695160
rect 42462 695090 42480 695160
rect 42410 694850 42428 694920
rect 42428 694850 42462 694920
rect 42462 694850 42480 694920
rect 42250 694480 42270 694550
rect 42270 694480 42304 694550
rect 42304 694480 42320 694550
rect 42250 694240 42270 694310
rect 42270 694240 42304 694310
rect 42304 694240 42320 694310
rect 42720 695090 42744 695160
rect 42744 695090 42778 695160
rect 42778 695090 42790 695160
rect 42720 694850 42744 694920
rect 42744 694850 42778 694920
rect 42778 694850 42790 694920
rect 42570 694480 42586 694550
rect 42586 694480 42620 694550
rect 42620 694480 42640 694550
rect 42570 694240 42586 694310
rect 42586 694240 42620 694310
rect 42620 694240 42640 694310
rect 43040 695090 43060 695160
rect 43060 695090 43094 695160
rect 43094 695090 43110 695160
rect 43040 694850 43060 694920
rect 43060 694850 43094 694920
rect 43094 694850 43110 694920
rect 42880 694480 42902 694550
rect 42902 694480 42936 694550
rect 42936 694480 42950 694550
rect 42880 694240 42902 694310
rect 42902 694240 42936 694310
rect 42936 694240 42950 694310
rect 43360 695090 43376 695160
rect 43376 695090 43410 695160
rect 43410 695090 43430 695160
rect 43360 694850 43376 694920
rect 43376 694850 43410 694920
rect 43410 694850 43430 694920
rect 43200 694480 43218 694550
rect 43218 694480 43252 694550
rect 43252 694480 43270 694550
rect 43200 694240 43218 694310
rect 43218 694240 43252 694310
rect 43252 694240 43270 694310
rect 43670 695090 43692 695160
rect 43692 695090 43726 695160
rect 43726 695090 43740 695160
rect 43670 694850 43692 694920
rect 43692 694850 43726 694920
rect 43726 694850 43740 694920
rect 43510 694480 43534 694550
rect 43534 694480 43568 694550
rect 43568 694480 43580 694550
rect 43510 694240 43534 694310
rect 43534 694240 43568 694310
rect 43568 694240 43580 694310
rect 43990 695090 44008 695160
rect 44008 695090 44042 695160
rect 44042 695090 44060 695160
rect 43990 694850 44008 694920
rect 44008 694850 44042 694920
rect 44042 694850 44060 694920
rect 43830 694480 43850 694550
rect 43850 694480 43884 694550
rect 43884 694480 43900 694550
rect 43830 694240 43850 694310
rect 43850 694240 43884 694310
rect 43884 694240 43900 694310
rect 44310 695090 44324 695160
rect 44324 695090 44358 695160
rect 44358 695090 44380 695160
rect 44310 694850 44324 694920
rect 44324 694850 44358 694920
rect 44358 694850 44380 694920
rect 44150 694480 44166 694550
rect 44166 694480 44200 694550
rect 44200 694480 44220 694550
rect 44150 694240 44166 694310
rect 44166 694240 44200 694310
rect 44200 694240 44220 694310
rect 44620 695090 44640 695160
rect 44640 695090 44674 695160
rect 44674 695090 44690 695160
rect 44620 694850 44640 694920
rect 44640 694850 44674 694920
rect 44674 694850 44690 694920
rect 44460 694480 44482 694550
rect 44482 694480 44516 694550
rect 44516 694480 44530 694550
rect 44460 694240 44482 694310
rect 44482 694240 44516 694310
rect 44516 694240 44530 694310
rect 44940 695090 44956 695160
rect 44956 695090 44990 695160
rect 44990 695090 45010 695160
rect 44940 694850 44956 694920
rect 44956 694850 44990 694920
rect 44990 694850 45010 694920
rect 44780 694480 44798 694550
rect 44798 694480 44832 694550
rect 44832 694480 44850 694550
rect 44780 694240 44798 694310
rect 44798 694240 44832 694310
rect 44832 694240 44850 694310
rect 45250 695090 45272 695160
rect 45272 695090 45306 695160
rect 45306 695090 45320 695160
rect 45250 694850 45272 694920
rect 45272 694850 45306 694920
rect 45306 694850 45320 694920
rect 45100 694480 45114 694550
rect 45114 694480 45148 694550
rect 45148 694480 45170 694550
rect 45100 694240 45114 694310
rect 45114 694240 45148 694310
rect 45148 694240 45170 694310
rect 45570 695090 45588 695160
rect 45588 695090 45622 695160
rect 45622 695090 45640 695160
rect 45570 694850 45588 694920
rect 45588 694850 45622 694920
rect 45622 694850 45640 694920
rect 45410 694480 45430 694550
rect 45430 694480 45464 694550
rect 45464 694480 45480 694550
rect 45410 694240 45430 694310
rect 45430 694240 45464 694310
rect 45464 694240 45480 694310
rect 45890 695090 45904 695160
rect 45904 695090 45938 695160
rect 45938 695090 45960 695160
rect 45890 694850 45904 694920
rect 45904 694850 45938 694920
rect 45938 694850 45960 694920
rect 45730 694480 45746 694550
rect 45746 694480 45780 694550
rect 45780 694480 45800 694550
rect 45730 694240 45746 694310
rect 45746 694240 45780 694310
rect 45780 694240 45800 694310
rect 46200 695090 46220 695160
rect 46220 695090 46254 695160
rect 46254 695090 46270 695160
rect 46200 694850 46220 694920
rect 46220 694850 46254 694920
rect 46254 694850 46270 694920
rect 46040 694480 46062 694550
rect 46062 694480 46096 694550
rect 46096 694480 46110 694550
rect 46040 694240 46062 694310
rect 46062 694240 46096 694310
rect 46096 694240 46110 694310
rect 46520 695090 46536 695160
rect 46536 695090 46570 695160
rect 46570 695090 46590 695160
rect 46520 694850 46536 694920
rect 46536 694850 46570 694920
rect 46570 694850 46590 694920
rect 46360 694480 46378 694550
rect 46378 694480 46412 694550
rect 46412 694480 46430 694550
rect 46360 694240 46378 694310
rect 46378 694240 46412 694310
rect 46412 694240 46430 694310
rect 46830 695090 46852 695160
rect 46852 695090 46886 695160
rect 46886 695090 46900 695160
rect 46830 694850 46852 694920
rect 46852 694850 46886 694920
rect 46886 694850 46900 694920
rect 46680 694480 46694 694550
rect 46694 694480 46728 694550
rect 46728 694480 46750 694550
rect 46680 694240 46694 694310
rect 46694 694240 46728 694310
rect 46728 694240 46750 694310
rect 47150 695090 47168 695160
rect 47168 695090 47202 695160
rect 47202 695090 47220 695160
rect 47150 694850 47168 694920
rect 47168 694850 47202 694920
rect 47202 694850 47220 694920
rect 46990 694480 47010 694550
rect 47010 694480 47044 694550
rect 47044 694480 47060 694550
rect 46990 694240 47010 694310
rect 47010 694240 47044 694310
rect 47044 694240 47060 694310
rect 47470 695090 47484 695160
rect 47484 695090 47518 695160
rect 47518 695090 47540 695160
rect 47470 694850 47484 694920
rect 47484 694850 47518 694920
rect 47518 694850 47540 694920
rect 47310 694480 47326 694550
rect 47326 694480 47360 694550
rect 47360 694480 47380 694550
rect 47310 694240 47326 694310
rect 47326 694240 47360 694310
rect 47360 694240 47380 694310
rect 47780 695090 47800 695160
rect 47800 695090 47834 695160
rect 47834 695090 47850 695160
rect 47780 694850 47800 694920
rect 47800 694850 47834 694920
rect 47834 694850 47850 694920
rect 47630 694480 47642 694550
rect 47642 694480 47676 694550
rect 47676 694480 47700 694550
rect 47630 694240 47642 694310
rect 47642 694240 47676 694310
rect 47676 694240 47700 694310
rect 42580 694118 42648 694140
rect 42648 694118 42660 694140
rect 46640 694118 46666 694140
rect 46666 694118 46720 694140
rect 42580 694060 42660 694118
rect 46640 694060 46720 694118
rect 44010 693730 44280 694000
rect 45060 693730 45330 694000
rect 38700 693360 38880 693460
rect 39120 693360 39300 693460
rect 42960 693420 42980 693490
rect 42980 693420 43014 693490
rect 43014 693420 43030 693490
rect 42960 693210 42980 693280
rect 42980 693210 43014 693280
rect 43014 693210 43030 693280
rect 43280 693420 43296 693490
rect 43296 693420 43330 693490
rect 43330 693420 43350 693490
rect 43280 693210 43296 693280
rect 43296 693210 43330 693280
rect 43330 693210 43350 693280
rect 43120 692780 43138 692850
rect 43138 692780 43172 692850
rect 43172 692780 43190 692850
rect 43120 692570 43138 692640
rect 43138 692570 43172 692640
rect 43172 692570 43190 692640
rect 43590 693420 43612 693490
rect 43612 693420 43646 693490
rect 43646 693420 43660 693490
rect 43590 693210 43612 693280
rect 43612 693210 43646 693280
rect 43646 693210 43660 693280
rect 43440 692780 43454 692850
rect 43454 692780 43488 692850
rect 43488 692780 43510 692850
rect 43440 692570 43454 692640
rect 43454 692570 43488 692640
rect 43488 692570 43510 692640
rect 43910 693420 43928 693490
rect 43928 693420 43962 693490
rect 43962 693420 43980 693490
rect 43910 693210 43928 693280
rect 43928 693210 43962 693280
rect 43962 693210 43980 693280
rect 43750 692780 43770 692850
rect 43770 692780 43804 692850
rect 43804 692780 43820 692850
rect 43750 692570 43770 692640
rect 43770 692570 43804 692640
rect 43804 692570 43820 692640
rect 44230 693420 44244 693490
rect 44244 693420 44278 693490
rect 44278 693420 44300 693490
rect 44230 693210 44244 693280
rect 44244 693210 44278 693280
rect 44278 693210 44300 693280
rect 44070 692780 44086 692850
rect 44086 692780 44120 692850
rect 44120 692780 44140 692850
rect 44070 692570 44086 692640
rect 44086 692570 44120 692640
rect 44120 692570 44140 692640
rect 44540 693420 44560 693490
rect 44560 693420 44594 693490
rect 44594 693420 44610 693490
rect 44540 693210 44560 693280
rect 44560 693210 44594 693280
rect 44594 693210 44610 693280
rect 44390 692780 44402 692850
rect 44402 692780 44436 692850
rect 44436 692780 44460 692850
rect 44390 692570 44402 692640
rect 44402 692570 44436 692640
rect 44436 692570 44460 692640
rect 44860 693420 44876 693490
rect 44876 693420 44910 693490
rect 44910 693420 44930 693490
rect 44860 693210 44876 693280
rect 44876 693210 44910 693280
rect 44910 693210 44930 693280
rect 44700 692780 44718 692850
rect 44718 692780 44752 692850
rect 44752 692780 44770 692850
rect 44700 692570 44718 692640
rect 44718 692570 44752 692640
rect 44752 692570 44770 692640
rect 45180 693420 45192 693490
rect 45192 693420 45226 693490
rect 45226 693420 45250 693490
rect 45180 693210 45192 693280
rect 45192 693210 45226 693280
rect 45226 693210 45250 693280
rect 45020 692780 45034 692850
rect 45034 692780 45068 692850
rect 45068 692780 45090 692850
rect 45020 692570 45034 692640
rect 45034 692570 45068 692640
rect 45068 692570 45090 692640
rect 45490 693420 45508 693490
rect 45508 693420 45542 693490
rect 45542 693420 45560 693490
rect 45490 693210 45508 693280
rect 45508 693210 45542 693280
rect 45542 693210 45560 693280
rect 45330 692780 45350 692850
rect 45350 692780 45384 692850
rect 45384 692780 45400 692850
rect 45330 692570 45350 692640
rect 45350 692570 45384 692640
rect 45384 692570 45400 692640
rect 45810 693420 45824 693490
rect 45824 693420 45858 693490
rect 45858 693420 45880 693490
rect 45810 693210 45824 693280
rect 45824 693210 45858 693280
rect 45858 693210 45880 693280
rect 45650 692780 45666 692850
rect 45666 692780 45700 692850
rect 45700 692780 45720 692850
rect 45650 692570 45666 692640
rect 45666 692570 45700 692640
rect 45700 692570 45720 692640
rect 46120 693420 46140 693490
rect 46140 693420 46174 693490
rect 46174 693420 46190 693490
rect 46120 693210 46140 693280
rect 46140 693210 46174 693280
rect 46174 693210 46190 693280
rect 45970 692780 45982 692850
rect 45982 692780 46016 692850
rect 46016 692780 46040 692850
rect 45970 692570 45982 692640
rect 45982 692570 46016 692640
rect 46016 692570 46040 692640
rect 46280 692780 46298 692850
rect 46298 692780 46332 692850
rect 46332 692780 46350 692850
rect 46280 692570 46298 692640
rect 46298 692570 46332 692640
rect 46332 692570 46350 692640
rect 52320 694850 52390 694920
rect 52430 694740 52500 694810
rect 49950 693360 50130 693460
rect 50370 693360 50550 693460
rect 43780 692380 44040 692390
rect 43780 692140 44040 692380
rect 43780 692130 44040 692140
rect 45280 692380 45540 692390
rect 45280 692140 45540 692380
rect 45280 692130 45540 692140
rect 42960 691870 42980 691940
rect 42980 691870 43014 691940
rect 43014 691870 43030 691940
rect 42960 691660 42980 691730
rect 42980 691660 43014 691730
rect 43014 691660 43030 691730
rect 43280 691870 43296 691940
rect 43296 691870 43330 691940
rect 43330 691870 43350 691940
rect 43280 691660 43296 691730
rect 43296 691660 43330 691730
rect 43330 691660 43350 691730
rect 43120 691240 43138 691310
rect 43138 691240 43172 691310
rect 43172 691240 43190 691310
rect 43120 691030 43138 691100
rect 43138 691030 43172 691100
rect 43172 691030 43190 691100
rect 43590 691870 43612 691940
rect 43612 691870 43646 691940
rect 43646 691870 43660 691940
rect 43590 691660 43612 691730
rect 43612 691660 43646 691730
rect 43646 691660 43660 691730
rect 43440 691240 43454 691310
rect 43454 691240 43488 691310
rect 43488 691240 43510 691310
rect 43440 691030 43454 691100
rect 43454 691030 43488 691100
rect 43488 691030 43510 691100
rect 43910 691870 43928 691940
rect 43928 691870 43962 691940
rect 43962 691870 43980 691940
rect 43910 691660 43928 691730
rect 43928 691660 43962 691730
rect 43962 691660 43980 691730
rect 43750 691240 43770 691310
rect 43770 691240 43804 691310
rect 43804 691240 43820 691310
rect 43750 691030 43770 691100
rect 43770 691030 43804 691100
rect 43804 691030 43820 691100
rect 44230 691870 44244 691940
rect 44244 691870 44278 691940
rect 44278 691870 44300 691940
rect 44230 691660 44244 691730
rect 44244 691660 44278 691730
rect 44278 691660 44300 691730
rect 44070 691240 44086 691310
rect 44086 691240 44120 691310
rect 44120 691240 44140 691310
rect 44070 691030 44086 691100
rect 44086 691030 44120 691100
rect 44120 691030 44140 691100
rect 44540 691870 44560 691940
rect 44560 691870 44594 691940
rect 44594 691870 44610 691940
rect 44540 691660 44560 691730
rect 44560 691660 44594 691730
rect 44594 691660 44610 691730
rect 44380 691240 44402 691310
rect 44402 691240 44436 691310
rect 44436 691240 44450 691310
rect 44380 691030 44402 691100
rect 44402 691030 44436 691100
rect 44436 691030 44450 691100
rect 44860 691870 44876 691940
rect 44876 691870 44910 691940
rect 44910 691870 44930 691940
rect 44860 691660 44876 691730
rect 44876 691660 44910 691730
rect 44910 691660 44930 691730
rect 44700 691240 44718 691310
rect 44718 691240 44752 691310
rect 44752 691240 44770 691310
rect 44700 691030 44718 691100
rect 44718 691030 44752 691100
rect 44752 691030 44770 691100
rect 45170 691870 45192 691940
rect 45192 691870 45226 691940
rect 45226 691870 45240 691940
rect 45170 691660 45192 691730
rect 45192 691660 45226 691730
rect 45226 691660 45240 691730
rect 45020 691240 45034 691310
rect 45034 691240 45068 691310
rect 45068 691240 45090 691310
rect 45020 691030 45034 691100
rect 45034 691030 45068 691100
rect 45068 691030 45090 691100
rect 45490 691870 45508 691940
rect 45508 691870 45542 691940
rect 45542 691870 45560 691940
rect 45490 691660 45508 691730
rect 45508 691660 45542 691730
rect 45542 691660 45560 691730
rect 45330 691240 45350 691310
rect 45350 691240 45384 691310
rect 45384 691240 45400 691310
rect 45330 691030 45350 691100
rect 45350 691030 45384 691100
rect 45384 691030 45400 691100
rect 45810 691870 45824 691940
rect 45824 691870 45858 691940
rect 45858 691870 45880 691940
rect 45810 691660 45824 691730
rect 45824 691660 45858 691730
rect 45858 691660 45880 691730
rect 45650 691240 45666 691310
rect 45666 691240 45700 691310
rect 45700 691240 45720 691310
rect 45650 691030 45666 691100
rect 45666 691030 45700 691100
rect 45700 691030 45720 691100
rect 46120 691870 46140 691940
rect 46140 691870 46174 691940
rect 46174 691870 46190 691940
rect 46120 691660 46140 691730
rect 46140 691660 46174 691730
rect 46174 691660 46190 691730
rect 45960 691240 45982 691310
rect 45982 691240 46016 691310
rect 46016 691240 46030 691310
rect 45960 691030 45982 691100
rect 45982 691030 46016 691100
rect 46016 691030 46030 691100
rect 46280 691240 46298 691310
rect 46298 691240 46332 691310
rect 46332 691240 46350 691310
rect 46280 691030 46298 691100
rect 46298 691030 46332 691100
rect 46332 691030 46350 691100
rect 541969 690892 542059 690962
rect 542139 690892 542229 690962
rect 544459 690892 544549 690962
rect 544629 690892 544719 690962
rect 546919 690892 546999 690972
rect 547089 690892 547169 690972
rect 566300 690900 566500 691100
rect 566700 690900 566900 691100
rect 567100 690900 567300 691100
rect 567500 690900 567700 691100
rect 567900 690900 568100 691100
rect 568300 690900 568500 691100
rect 568700 690900 568900 691100
rect 569100 690900 569300 691100
rect 569500 690900 569700 691100
rect 569900 690900 570100 691100
rect 570300 690900 570500 691100
rect 570700 690900 570900 691100
rect 571100 690900 571300 691100
rect 571500 690900 571700 691100
rect 541969 690784 542049 690852
rect 542139 690784 542219 690852
rect 544459 690784 544539 690852
rect 544629 690784 544709 690852
rect 546919 690784 546999 690842
rect 547089 690784 547169 690842
rect 541969 690772 542049 690784
rect 542139 690772 542219 690784
rect 544459 690772 544539 690784
rect 544629 690772 544709 690784
rect 546919 690762 546999 690784
rect 547089 690762 547169 690784
rect 541089 690626 541169 690682
rect 541239 690626 541319 690682
rect 541419 690654 541449 690722
rect 541449 690654 541523 690722
rect 541523 690654 541549 690722
rect 542659 690654 542685 690722
rect 542685 690654 542759 690722
rect 542759 690654 542789 690722
rect 541419 690652 541549 690654
rect 542659 690652 542789 690654
rect 543579 690626 543659 690682
rect 543729 690626 543809 690682
rect 543889 690654 543921 690722
rect 543921 690654 543995 690722
rect 543995 690654 544019 690722
rect 545129 690654 545157 690722
rect 545157 690654 545231 690722
rect 545231 690654 545259 690722
rect 543889 690652 544019 690654
rect 545129 690652 545259 690654
rect 546059 690626 546139 690682
rect 546209 690626 546289 690682
rect 546369 690654 546393 690722
rect 546393 690654 546467 690722
rect 546467 690654 546499 690722
rect 547599 690654 547629 690722
rect 547629 690654 547703 690722
rect 547703 690654 547729 690722
rect 546369 690652 546499 690654
rect 547599 690652 547729 690654
rect 540699 690592 540779 690612
rect 540869 690592 540949 690612
rect 541089 690602 541169 690626
rect 541239 690602 541319 690626
rect 543219 690592 543299 690612
rect 543389 690592 543469 690612
rect 543579 690602 543659 690626
rect 543729 690602 543809 690626
rect 545709 690592 545789 690612
rect 545879 690592 545959 690612
rect 546059 690602 546139 690626
rect 546209 690602 546289 690626
rect 548159 690592 548239 690612
rect 548329 690592 548409 690612
rect 540699 690532 540779 690592
rect 540869 690532 540949 690592
rect 543219 690532 543299 690592
rect 543389 690532 543469 690592
rect 545709 690532 545789 690592
rect 545879 690532 545959 690592
rect 548159 690532 548239 690592
rect 548329 690532 548409 690592
rect 566300 690500 566500 690700
rect 566700 690500 566900 690700
rect 567100 690500 567300 690700
rect 567500 690500 567700 690700
rect 567900 690500 568100 690700
rect 568300 690500 568500 690700
rect 568700 690500 568900 690700
rect 569100 690500 569300 690700
rect 569500 690500 569700 690700
rect 569900 690500 570100 690700
rect 570300 690500 570500 690700
rect 570700 690500 570900 690700
rect 571100 690500 571300 690700
rect 571500 690500 571700 690700
rect 44060 690310 44081 690380
rect 44081 690310 44115 690380
rect 44115 690310 44130 690380
rect 44060 690020 44081 690090
rect 44081 690020 44115 690090
rect 44115 690020 44130 690090
rect 44380 690310 44397 690380
rect 44397 690310 44431 690380
rect 44431 690310 44450 690380
rect 44380 690020 44397 690090
rect 44397 690020 44431 690090
rect 44431 690020 44450 690090
rect 44220 689750 44239 689820
rect 44239 689750 44273 689820
rect 44273 689750 44290 689820
rect 44220 689460 44239 689530
rect 44239 689460 44273 689530
rect 44273 689460 44290 689530
rect 44690 690310 44713 690380
rect 44713 690310 44747 690380
rect 44747 690310 44760 690380
rect 44690 690020 44713 690090
rect 44713 690020 44747 690090
rect 44747 690020 44760 690090
rect 44530 689750 44555 689820
rect 44555 689750 44589 689820
rect 44589 689750 44600 689820
rect 44530 689460 44555 689530
rect 44555 689460 44589 689530
rect 44589 689460 44600 689530
rect 45010 690310 45029 690380
rect 45029 690310 45063 690380
rect 45063 690310 45080 690380
rect 45010 690020 45029 690090
rect 45029 690020 45063 690090
rect 45063 690020 45080 690090
rect 44850 689750 44871 689820
rect 44871 689750 44905 689820
rect 44905 689750 44920 689820
rect 44850 689460 44871 689530
rect 44871 689460 44905 689530
rect 44905 689460 44920 689530
rect 47200 690200 47300 690300
rect 541969 690244 542049 690312
rect 542139 690244 542219 690312
rect 544459 690244 544539 690312
rect 544629 690244 544709 690312
rect 546919 690244 546999 690302
rect 547089 690244 547169 690302
rect 541969 690232 542049 690244
rect 542139 690232 542219 690244
rect 544459 690232 544539 690244
rect 544629 690232 544709 690244
rect 546919 690222 546999 690244
rect 547089 690222 547169 690244
rect 541089 690086 541169 690142
rect 541239 690086 541319 690142
rect 541419 690114 541449 690182
rect 541449 690114 541523 690182
rect 541523 690114 541549 690182
rect 542659 690114 542685 690182
rect 542685 690114 542759 690182
rect 542759 690114 542789 690182
rect 541419 690112 541549 690114
rect 542659 690112 542789 690114
rect 543579 690086 543659 690142
rect 543729 690086 543809 690142
rect 543889 690114 543921 690182
rect 543921 690114 543995 690182
rect 543995 690114 544019 690182
rect 545129 690114 545157 690182
rect 545157 690114 545231 690182
rect 545231 690114 545259 690182
rect 543889 690112 544019 690114
rect 545129 690112 545259 690114
rect 546059 690086 546139 690142
rect 546209 690086 546289 690142
rect 546369 690114 546393 690182
rect 546393 690114 546467 690182
rect 546467 690114 546499 690182
rect 547599 690114 547629 690182
rect 547629 690114 547703 690182
rect 547703 690114 547729 690182
rect 546369 690112 546499 690114
rect 547599 690112 547729 690114
rect 540699 690052 540779 690072
rect 540869 690052 540949 690072
rect 541089 690062 541169 690086
rect 541239 690062 541319 690086
rect 543219 690052 543299 690072
rect 543389 690052 543469 690072
rect 543579 690062 543659 690086
rect 543729 690062 543809 690086
rect 545709 690052 545789 690072
rect 545879 690052 545959 690072
rect 546059 690062 546139 690086
rect 546209 690062 546289 690086
rect 548159 690052 548239 690062
rect 548329 690052 548409 690062
rect 45170 689750 45187 689820
rect 45187 689750 45221 689820
rect 45221 689750 45240 689820
rect 45170 689460 45187 689530
rect 45187 689460 45221 689530
rect 45221 689460 45240 689530
rect 47200 689800 47300 690000
rect 540699 689992 540779 690052
rect 540869 689992 540949 690052
rect 543219 689992 543299 690052
rect 543389 689992 543469 690052
rect 545709 689992 545789 690052
rect 545879 689992 545959 690052
rect 548159 689982 548239 690052
rect 548329 689982 548409 690052
rect 566300 690100 566500 690300
rect 566700 690100 566900 690300
rect 567100 690100 567300 690300
rect 567500 690100 567700 690300
rect 567900 690100 568100 690300
rect 568300 690100 568500 690300
rect 568700 690100 568900 690300
rect 569100 690100 569300 690300
rect 569500 690100 569700 690300
rect 569900 690100 570100 690300
rect 570300 690100 570500 690300
rect 570700 690100 570900 690300
rect 571100 690100 571300 690300
rect 571500 690100 571700 690300
rect 541979 689842 542069 689912
rect 542119 689842 542209 689912
rect 544459 689842 544549 689912
rect 544619 689852 544709 689922
rect 546919 689852 546999 689922
rect 547089 689852 547169 689922
rect 541969 689704 542049 689772
rect 542139 689704 542219 689772
rect 544459 689704 544539 689782
rect 544629 689704 544709 689782
rect 546919 689704 546999 689762
rect 547089 689704 547169 689762
rect 541969 689692 542049 689704
rect 542139 689692 542219 689704
rect 544459 689702 544539 689704
rect 544629 689702 544709 689704
rect 546919 689682 546999 689704
rect 547089 689682 547169 689704
rect 566300 689700 566500 689900
rect 566700 689700 566900 689900
rect 567100 689700 567300 689900
rect 567500 689700 567700 689900
rect 567900 689700 568100 689900
rect 568300 689700 568500 689900
rect 568700 689700 568900 689900
rect 569100 689700 569300 689900
rect 569500 689700 569700 689900
rect 569900 689700 570100 689900
rect 570300 689700 570500 689900
rect 570700 689700 570900 689900
rect 571100 689700 571300 689900
rect 571500 689700 571700 689900
rect 47200 689500 47300 689600
rect 541089 689546 541169 689602
rect 541239 689546 541319 689602
rect 541419 689574 541449 689642
rect 541449 689574 541523 689642
rect 541523 689574 541549 689642
rect 542659 689574 542685 689642
rect 542685 689574 542759 689642
rect 542759 689574 542789 689642
rect 541419 689572 541549 689574
rect 542659 689572 542789 689574
rect 543579 689546 543659 689602
rect 543729 689546 543809 689602
rect 543889 689574 543921 689642
rect 543921 689574 543995 689642
rect 543995 689574 544019 689642
rect 545129 689574 545157 689642
rect 545157 689574 545231 689642
rect 545231 689574 545259 689642
rect 543889 689572 544019 689574
rect 545129 689572 545259 689574
rect 546069 689546 546149 689602
rect 546209 689546 546289 689602
rect 546369 689574 546393 689642
rect 546393 689574 546467 689642
rect 546467 689574 546499 689642
rect 547599 689574 547629 689642
rect 547629 689574 547703 689642
rect 547703 689574 547729 689642
rect 546369 689572 546499 689574
rect 547599 689572 547729 689574
rect 540699 689512 540779 689532
rect 540869 689512 540949 689532
rect 541089 689522 541169 689546
rect 541239 689522 541319 689546
rect 543219 689512 543299 689532
rect 543389 689512 543469 689532
rect 543579 689522 543659 689546
rect 543729 689522 543809 689546
rect 546069 689522 546149 689546
rect 546209 689522 546289 689546
rect 545709 689512 545789 689522
rect 545879 689512 545959 689522
rect 548159 689512 548239 689532
rect 548329 689512 548409 689532
rect 540699 689452 540779 689512
rect 540869 689452 540949 689512
rect 543219 689452 543299 689512
rect 543389 689452 543469 689512
rect 545709 689442 545789 689512
rect 545879 689442 545959 689512
rect 548159 689452 548239 689512
rect 548329 689452 548409 689512
rect 541979 689302 542059 689382
rect 542149 689302 542229 689382
rect 544459 689302 544539 689382
rect 544629 689302 544709 689382
rect 546919 689302 546999 689382
rect 547089 689302 547169 689382
rect 566300 689300 566500 689500
rect 566700 689300 566900 689500
rect 567100 689300 567300 689500
rect 567500 689300 567700 689500
rect 567900 689300 568100 689500
rect 568300 689300 568500 689500
rect 568700 689300 568900 689500
rect 569100 689300 569300 689500
rect 569500 689300 569700 689500
rect 569900 689300 570100 689500
rect 570300 689300 570500 689500
rect 570700 689300 570900 689500
rect 571100 689300 571300 689500
rect 571500 689300 571700 689500
rect 44520 689281 44780 689290
rect 44520 689247 44780 689281
rect 44520 689075 44780 689247
rect 541979 689172 542059 689252
rect 542149 689172 542229 689252
rect 544459 689182 544539 689262
rect 544629 689182 544709 689262
rect 546919 689172 546999 689252
rect 547089 689172 547169 689252
rect 44520 689041 44780 689075
rect 44520 689030 44780 689041
rect 541419 689034 541449 689102
rect 541449 689034 541523 689102
rect 541523 689034 541549 689102
rect 541419 689032 541549 689034
rect 542659 689034 542685 689102
rect 542685 689034 542759 689102
rect 542759 689034 542789 689102
rect 542659 689032 542789 689034
rect 543889 689034 543921 689102
rect 543921 689034 543995 689102
rect 543995 689034 544019 689102
rect 543889 689032 544019 689034
rect 545129 689034 545157 689102
rect 545157 689034 545231 689102
rect 545231 689034 545259 689102
rect 545129 689032 545259 689034
rect 546359 689034 546393 689102
rect 546393 689034 546467 689102
rect 546467 689034 546489 689102
rect 546359 689032 546489 689034
rect 547599 689034 547629 689102
rect 547629 689034 547703 689102
rect 547703 689034 547729 689102
rect 547599 689032 547729 689034
rect 540699 688972 540779 688992
rect 540869 688972 540949 688992
rect 542379 688972 542459 689002
rect 542489 688972 542569 689002
rect 543209 688972 543289 688992
rect 543379 688972 543459 688992
rect 544789 688972 544869 689002
rect 544899 688972 544979 689002
rect 545699 688972 545779 688992
rect 545869 688972 545949 688992
rect 547249 688972 547329 688992
rect 547359 688972 547439 688992
rect 548189 688972 548269 688992
rect 548359 688972 548439 688992
rect 42000 688600 42100 688700
rect 42000 688300 42100 688500
rect 44060 688790 44081 688860
rect 44081 688790 44115 688860
rect 44115 688790 44130 688860
rect 44060 688500 44081 688570
rect 44081 688500 44115 688570
rect 44115 688500 44130 688570
rect 42000 688100 42100 688200
rect 44380 688790 44397 688860
rect 44397 688790 44431 688860
rect 44431 688790 44450 688860
rect 44380 688500 44397 688570
rect 44397 688500 44431 688570
rect 44431 688500 44450 688570
rect 44220 688230 44239 688300
rect 44239 688230 44273 688300
rect 44273 688230 44290 688300
rect 44220 687940 44239 688010
rect 44239 687940 44273 688010
rect 44273 687940 44290 688010
rect 44690 688790 44713 688860
rect 44713 688790 44747 688860
rect 44747 688790 44760 688860
rect 44690 688500 44713 688570
rect 44713 688500 44747 688570
rect 44747 688500 44760 688570
rect 44530 688230 44555 688300
rect 44555 688230 44589 688300
rect 44589 688230 44600 688300
rect 44530 687940 44555 688010
rect 44555 687940 44589 688010
rect 44589 687940 44600 688010
rect 45010 688790 45029 688860
rect 45029 688790 45063 688860
rect 45063 688790 45080 688860
rect 45010 688500 45029 688570
rect 45029 688500 45063 688570
rect 45063 688500 45080 688570
rect 44850 688230 44871 688300
rect 44871 688230 44905 688300
rect 44905 688230 44920 688300
rect 44850 687940 44871 688010
rect 44871 687940 44905 688010
rect 44905 687940 44920 688010
rect 45170 688230 45187 688300
rect 45187 688230 45221 688300
rect 45221 688230 45240 688300
rect 45170 687940 45187 688010
rect 45187 687940 45221 688010
rect 45221 687940 45240 688010
rect 540699 688912 540779 688972
rect 540869 688912 540949 688972
rect 542379 688922 542459 688972
rect 542489 688922 542569 688972
rect 543209 688912 543289 688972
rect 543379 688912 543459 688972
rect 544789 688922 544869 688972
rect 544899 688922 544979 688972
rect 545699 688912 545779 688972
rect 545869 688912 545949 688972
rect 547249 688912 547329 688972
rect 547359 688912 547439 688972
rect 548189 688912 548269 688972
rect 548359 688912 548439 688972
rect 541979 688592 542059 688672
rect 542149 688592 542229 688672
rect 544459 688602 544539 688682
rect 544629 688602 544709 688682
rect 546919 688592 546999 688672
rect 547089 688592 547169 688672
rect 541419 688454 541449 688522
rect 541449 688454 541523 688522
rect 541523 688454 541549 688522
rect 541419 688452 541549 688454
rect 542659 688454 542685 688522
rect 542685 688454 542759 688522
rect 542759 688454 542789 688522
rect 542659 688452 542789 688454
rect 543899 688454 543921 688522
rect 543921 688454 543995 688522
rect 543995 688454 544029 688522
rect 543899 688452 544029 688454
rect 545129 688454 545157 688522
rect 545157 688454 545231 688522
rect 545231 688454 545259 688522
rect 545129 688452 545259 688454
rect 546359 688454 546393 688522
rect 546393 688454 546467 688522
rect 546467 688454 546489 688522
rect 546359 688452 546489 688454
rect 547599 688454 547629 688522
rect 547629 688454 547703 688522
rect 547703 688454 547729 688522
rect 547599 688452 547729 688454
rect 540699 688392 540779 688412
rect 540869 688392 540949 688412
rect 543209 688392 543289 688412
rect 543379 688392 543459 688412
rect 544789 688392 544869 688412
rect 544899 688392 544979 688412
rect 545699 688392 545779 688402
rect 545869 688392 545949 688402
rect 547249 688392 547329 688412
rect 547359 688392 547439 688412
rect 548189 688392 548269 688412
rect 548359 688392 548439 688412
rect 540699 688332 540779 688392
rect 540869 688332 540949 688392
rect 542379 688312 542459 688392
rect 542489 688312 542569 688392
rect 543209 688332 543289 688392
rect 543379 688332 543459 688392
rect 544789 688332 544869 688392
rect 544899 688332 544979 688392
rect 545699 688322 545779 688392
rect 545869 688322 545949 688392
rect 547249 688332 547329 688392
rect 547359 688332 547439 688392
rect 548189 688332 548269 688392
rect 548359 688332 548439 688392
rect 541979 688142 542069 688222
rect 542139 688142 542229 688222
rect 544459 688142 544539 688212
rect 544629 688142 544709 688212
rect 546919 688142 546999 688212
rect 547089 688142 547169 688212
rect 554129 688162 554259 688302
rect 554389 688162 554519 688302
rect 534629 687992 534759 688132
rect 534879 687992 535009 688132
rect 541979 688012 542059 688092
rect 542149 688012 542229 688092
rect 544459 688022 544539 688102
rect 544629 688022 544709 688102
rect 546919 688012 546999 688092
rect 547089 688012 547169 688092
rect 44520 687761 44780 687770
rect 44520 687727 44780 687761
rect 44520 687554 44780 687727
rect 44520 687520 44780 687554
rect 44520 687510 44780 687520
rect 42260 687380 42370 687490
rect 42510 687380 42620 687490
rect 46660 687380 46770 687490
rect 46910 687380 47020 687490
rect 43070 687270 43090 687340
rect 43090 687270 43124 687340
rect 43124 687270 43140 687340
rect 43070 687090 43090 687160
rect 43090 687090 43124 687160
rect 43124 687090 43140 687160
rect 43590 687270 43606 687340
rect 43606 687270 43640 687340
rect 43640 687270 43660 687340
rect 43590 687090 43606 687160
rect 43606 687090 43640 687160
rect 43640 687090 43660 687160
rect 43330 686600 43348 686670
rect 43348 686600 43382 686670
rect 43382 686600 43400 686670
rect 43330 686420 43348 686490
rect 43348 686420 43382 686490
rect 43382 686420 43400 686490
rect 44100 687270 44122 687340
rect 44122 687270 44156 687340
rect 44156 687270 44170 687340
rect 44100 687090 44122 687160
rect 44122 687090 44156 687160
rect 44156 687090 44170 687160
rect 43840 686600 43864 686670
rect 43864 686600 43898 686670
rect 43898 686600 43910 686670
rect 43840 686420 43864 686490
rect 43864 686420 43898 686490
rect 43898 686420 43910 686490
rect 44620 687270 44638 687340
rect 44638 687270 44672 687340
rect 44672 687270 44690 687340
rect 44620 687090 44638 687160
rect 44638 687090 44672 687160
rect 44672 687090 44690 687160
rect 44360 686600 44380 686670
rect 44380 686600 44414 686670
rect 44414 686600 44430 686670
rect 44360 686420 44380 686490
rect 44380 686420 44414 686490
rect 44414 686420 44430 686490
rect 45130 687270 45154 687340
rect 45154 687270 45188 687340
rect 45188 687270 45200 687340
rect 45130 687090 45154 687160
rect 45154 687090 45188 687160
rect 45188 687090 45200 687160
rect 44880 686600 44896 686670
rect 44896 686600 44930 686670
rect 44930 686600 44950 686670
rect 44880 686420 44896 686490
rect 44896 686420 44930 686490
rect 44930 686420 44950 686490
rect 45650 687270 45670 687340
rect 45670 687270 45704 687340
rect 45704 687270 45720 687340
rect 45650 687090 45670 687160
rect 45670 687090 45704 687160
rect 45704 687090 45720 687160
rect 45390 686600 45412 686670
rect 45412 686600 45446 686670
rect 45446 686600 45460 686670
rect 45390 686420 45412 686490
rect 45412 686420 45446 686490
rect 45446 686420 45460 686490
rect 46170 687270 46186 687340
rect 46186 687270 46220 687340
rect 46220 687270 46240 687340
rect 46170 687090 46186 687160
rect 46186 687090 46220 687160
rect 46220 687090 46240 687160
rect 45910 686600 45928 686670
rect 45928 686600 45962 686670
rect 45962 686600 45980 686670
rect 45910 686420 45928 686490
rect 45928 686420 45962 686490
rect 45962 686420 45980 686490
rect 541419 687874 541449 687942
rect 541449 687874 541523 687942
rect 541523 687874 541549 687942
rect 541419 687872 541549 687874
rect 542659 687874 542685 687942
rect 542685 687874 542759 687942
rect 542759 687874 542789 687942
rect 542659 687872 542789 687874
rect 543889 687874 543921 687942
rect 543921 687874 543995 687942
rect 543995 687874 544019 687942
rect 543889 687872 544019 687874
rect 545129 687874 545157 687942
rect 545157 687874 545231 687942
rect 545231 687874 545259 687942
rect 545129 687872 545259 687874
rect 546359 687874 546393 687942
rect 546393 687874 546467 687942
rect 546467 687874 546489 687942
rect 546359 687872 546489 687874
rect 547599 687874 547629 687942
rect 547629 687874 547703 687942
rect 547703 687874 547729 687942
rect 547599 687872 547729 687874
rect 542380 687812 542460 687830
rect 542500 687812 542580 687830
rect 543209 687812 543289 687832
rect 543379 687812 543459 687832
rect 544789 687812 544869 687832
rect 544899 687812 544979 687832
rect 545699 687812 545779 687832
rect 545869 687812 545949 687832
rect 547249 687812 547329 687832
rect 547359 687812 547439 687832
rect 548189 687812 548269 687832
rect 548359 687812 548439 687832
rect 540679 687722 540759 687802
rect 540889 687722 540969 687802
rect 542380 687750 542460 687812
rect 542500 687750 542580 687812
rect 543209 687752 543289 687812
rect 543379 687752 543459 687812
rect 544789 687752 544869 687812
rect 544899 687752 544979 687812
rect 545699 687752 545779 687812
rect 545869 687752 545949 687812
rect 547249 687752 547329 687812
rect 547359 687752 547439 687812
rect 548189 687752 548269 687812
rect 548359 687752 548439 687812
rect 540099 687482 540179 687562
rect 540329 687482 540409 687562
rect 542649 687472 542729 687552
rect 542819 687472 542899 687552
rect 545109 687472 545189 687552
rect 545299 687472 545379 687552
rect 547559 687472 547639 687552
rect 547749 687472 547829 687552
rect 550069 687472 550149 687552
rect 550239 687472 550319 687552
rect 539579 687334 539609 687402
rect 539609 687334 539683 687402
rect 539683 687334 539709 687402
rect 539579 687332 539709 687334
rect 540819 687334 540845 687402
rect 540845 687334 540919 687402
rect 540919 687334 540949 687402
rect 540819 687332 540949 687334
rect 542049 687334 542081 687402
rect 542081 687334 542155 687402
rect 542155 687334 542179 687402
rect 542049 687332 542179 687334
rect 543289 687334 543317 687402
rect 543317 687334 543391 687402
rect 543391 687334 543419 687402
rect 543289 687332 543419 687334
rect 544529 687334 544553 687402
rect 544553 687334 544627 687402
rect 544627 687334 544659 687402
rect 544529 687332 544659 687334
rect 545759 687334 545789 687402
rect 545789 687334 545863 687402
rect 545863 687334 545889 687402
rect 545759 687332 545889 687334
rect 546999 687334 547025 687402
rect 547025 687334 547099 687402
rect 547099 687334 547129 687402
rect 546999 687332 547129 687334
rect 548229 687334 548261 687402
rect 548261 687334 548335 687402
rect 548335 687334 548359 687402
rect 548229 687332 548359 687334
rect 549469 687334 549497 687402
rect 549497 687334 549571 687402
rect 549571 687334 549599 687402
rect 549469 687332 549599 687334
rect 538849 687272 538929 687282
rect 539059 687272 539139 687282
rect 541329 687272 541409 687282
rect 541549 687272 541629 687282
rect 543859 687272 543939 687282
rect 544039 687272 544119 687282
rect 538849 687202 538929 687272
rect 539059 687202 539139 687272
rect 541329 687202 541409 687272
rect 541549 687202 541629 687272
rect 543859 687202 543939 687272
rect 544039 687202 544119 687272
rect 546319 687192 546399 687272
rect 546499 687192 546579 687272
rect 548799 687192 548879 687272
rect 548969 687192 549049 687272
rect 540119 687062 540209 687142
rect 540299 687062 540389 687142
rect 542649 687062 542739 687142
rect 542809 687062 542899 687142
rect 545119 687062 545209 687142
rect 545279 687062 545369 687142
rect 547569 687062 547659 687142
rect 547729 687062 547819 687142
rect 550069 687062 550159 687142
rect 550229 687062 550319 687142
rect 540099 686942 540179 687022
rect 540329 686942 540409 687022
rect 542649 686932 542729 687012
rect 542819 686942 542899 687022
rect 545109 686942 545189 687022
rect 545299 686942 545379 687022
rect 547559 686932 547639 687012
rect 547749 686932 547829 687012
rect 550069 686932 550149 687012
rect 550239 686932 550319 687012
rect 539579 686862 539709 686872
rect 539579 686802 539609 686862
rect 539609 686802 539683 686862
rect 539683 686802 539709 686862
rect 540819 686794 540845 686862
rect 540845 686794 540919 686862
rect 540919 686794 540949 686862
rect 540819 686792 540949 686794
rect 542049 686794 542081 686862
rect 542081 686794 542155 686862
rect 542155 686794 542179 686862
rect 542049 686792 542179 686794
rect 543289 686794 543317 686862
rect 543317 686794 543391 686862
rect 543391 686794 543419 686862
rect 543289 686792 543419 686794
rect 544529 686794 544553 686862
rect 544553 686794 544627 686862
rect 544627 686794 544659 686862
rect 544529 686792 544659 686794
rect 545759 686794 545789 686862
rect 545789 686794 545863 686862
rect 545863 686794 545889 686862
rect 545759 686792 545889 686794
rect 546999 686794 547025 686862
rect 547025 686794 547099 686862
rect 547099 686794 547129 686862
rect 546999 686792 547129 686794
rect 548229 686794 548261 686862
rect 548261 686794 548335 686862
rect 548335 686794 548359 686862
rect 548229 686792 548359 686794
rect 549469 686794 549497 686862
rect 549497 686794 549571 686862
rect 549571 686794 549599 686862
rect 549469 686792 549599 686794
rect 538849 686732 538929 686742
rect 539059 686732 539139 686742
rect 541329 686732 541409 686742
rect 541549 686732 541629 686742
rect 543859 686732 543939 686742
rect 544049 686732 544129 686742
rect 538849 686662 538929 686732
rect 539059 686662 539139 686732
rect 541329 686662 541409 686732
rect 541549 686662 541629 686732
rect 543859 686662 543939 686732
rect 544049 686662 544129 686732
rect 546319 686652 546399 686732
rect 546499 686652 546579 686732
rect 548799 686652 548879 686732
rect 548969 686652 549049 686732
rect 42260 686270 42370 686380
rect 42510 686270 42620 686380
rect 46660 686270 46770 686380
rect 46910 686270 47020 686380
rect 44530 686240 44780 686250
rect 44530 686206 44780 686240
rect 44530 686034 44780 686206
rect 44530 686000 44780 686034
rect 42260 685860 42370 685970
rect 42510 685860 42620 685970
rect 46660 685860 46770 685970
rect 46910 685860 47020 685970
rect 42810 685750 42830 685820
rect 42830 685750 42864 685820
rect 42864 685750 42880 685820
rect 42810 685570 42830 685640
rect 42830 685570 42864 685640
rect 42864 685570 42880 685640
rect 43330 685750 43346 685820
rect 43346 685750 43380 685820
rect 43380 685750 43400 685820
rect 43330 685570 43346 685640
rect 43346 685570 43380 685640
rect 43380 685570 43400 685640
rect 43070 685080 43088 685150
rect 43088 685080 43122 685150
rect 43122 685080 43140 685150
rect 43070 684900 43088 684970
rect 43088 684900 43122 684970
rect 43122 684900 43140 684970
rect 43840 685750 43862 685820
rect 43862 685750 43896 685820
rect 43896 685750 43910 685820
rect 43840 685570 43862 685640
rect 43862 685570 43896 685640
rect 43896 685570 43910 685640
rect 43580 685080 43604 685150
rect 43604 685080 43638 685150
rect 43638 685080 43650 685150
rect 43580 684900 43604 684970
rect 43604 684900 43638 684970
rect 43638 684900 43650 684970
rect 44360 685750 44378 685820
rect 44378 685750 44412 685820
rect 44412 685750 44430 685820
rect 44360 685570 44378 685640
rect 44378 685570 44412 685640
rect 44412 685570 44430 685640
rect 44100 685080 44120 685150
rect 44120 685080 44154 685150
rect 44154 685080 44170 685150
rect 44100 684900 44120 684970
rect 44120 684900 44154 684970
rect 44154 684900 44170 684970
rect 44870 685750 44894 685820
rect 44894 685750 44928 685820
rect 44928 685750 44940 685820
rect 44870 685570 44894 685640
rect 44894 685570 44928 685640
rect 44928 685570 44940 685640
rect 44620 685080 44636 685150
rect 44636 685080 44670 685150
rect 44670 685080 44690 685150
rect 44620 684900 44636 684970
rect 44636 684900 44670 684970
rect 44670 684900 44690 684970
rect 45390 685750 45410 685820
rect 45410 685750 45444 685820
rect 45444 685750 45460 685820
rect 45390 685570 45410 685640
rect 45410 685570 45444 685640
rect 45444 685570 45460 685640
rect 45130 685080 45152 685150
rect 45152 685080 45186 685150
rect 45186 685080 45200 685150
rect 45130 684900 45152 684970
rect 45152 684900 45186 684970
rect 45186 684900 45200 684970
rect 45910 685750 45926 685820
rect 45926 685750 45960 685820
rect 45960 685750 45980 685820
rect 45910 685570 45926 685640
rect 45926 685570 45960 685640
rect 45960 685570 45980 685640
rect 45650 685080 45668 685150
rect 45668 685080 45702 685150
rect 45702 685080 45720 685150
rect 45650 684900 45668 684970
rect 45668 684900 45702 684970
rect 45702 684900 45720 684970
rect 46420 685750 46442 685820
rect 46442 685750 46476 685820
rect 46476 685750 46490 685820
rect 46420 685570 46442 685640
rect 46442 685570 46476 685640
rect 46476 685570 46490 685640
rect 46160 685080 46184 685150
rect 46184 685080 46218 685150
rect 46218 685080 46230 685150
rect 46160 684900 46184 684970
rect 46184 684900 46218 684970
rect 46218 684900 46230 684970
rect 540099 686402 540179 686482
rect 540329 686402 540409 686482
rect 542639 686392 542719 686472
rect 542809 686392 542889 686472
rect 545109 686392 545189 686472
rect 545289 686392 545369 686472
rect 547559 686392 547639 686472
rect 547749 686392 547829 686472
rect 550069 686392 550149 686472
rect 550239 686392 550319 686472
rect 539579 686254 539609 686322
rect 539609 686254 539683 686322
rect 539683 686254 539709 686322
rect 539579 686252 539709 686254
rect 540819 686254 540845 686322
rect 540845 686254 540919 686322
rect 540919 686254 540949 686322
rect 540819 686252 540949 686254
rect 542049 686254 542081 686322
rect 542081 686254 542155 686322
rect 542155 686254 542179 686322
rect 542049 686252 542179 686254
rect 543289 686254 543317 686322
rect 543317 686254 543391 686322
rect 543391 686254 543419 686322
rect 543289 686252 543419 686254
rect 544529 686254 544553 686322
rect 544553 686254 544627 686322
rect 544627 686254 544659 686322
rect 544529 686252 544659 686254
rect 545759 686254 545789 686322
rect 545789 686254 545863 686322
rect 545863 686254 545889 686322
rect 545759 686252 545889 686254
rect 546999 686254 547025 686322
rect 547025 686254 547099 686322
rect 547099 686254 547129 686322
rect 546999 686252 547129 686254
rect 548229 686254 548261 686322
rect 548261 686254 548335 686322
rect 548335 686254 548359 686322
rect 548229 686252 548359 686254
rect 549469 686254 549497 686322
rect 549497 686254 549571 686322
rect 549571 686254 549599 686322
rect 549469 686252 549599 686254
rect 538849 686192 538929 686202
rect 539059 686192 539139 686202
rect 541319 686192 541399 686202
rect 541559 686192 541639 686202
rect 543859 686192 543939 686202
rect 544039 686192 544119 686202
rect 538849 686122 538929 686192
rect 539059 686122 539139 686192
rect 541319 686122 541399 686192
rect 541559 686122 541639 686192
rect 543859 686122 543939 686192
rect 544039 686122 544119 686192
rect 546329 686112 546409 686192
rect 546499 686112 546579 686192
rect 548799 686112 548879 686192
rect 548969 686112 549049 686192
rect 540119 685982 540209 686062
rect 540299 685992 540389 686072
rect 542649 685982 542739 686062
rect 542809 685982 542899 686062
rect 545119 685982 545209 686062
rect 545279 685982 545369 686062
rect 547569 685982 547659 686062
rect 547729 685982 547819 686062
rect 550069 685982 550159 686062
rect 550229 685982 550319 686062
rect 540099 685852 540179 685932
rect 540329 685852 540409 685932
rect 542629 685862 542709 685942
rect 542819 685862 542899 685942
rect 545109 685852 545189 685932
rect 545299 685852 545379 685932
rect 547559 685852 547639 685932
rect 547749 685852 547829 685932
rect 550069 685844 550149 685922
rect 550239 685844 550319 685922
rect 550069 685842 550149 685844
rect 550239 685842 550319 685844
rect 539579 685714 539609 685782
rect 539609 685714 539683 685782
rect 539683 685714 539709 685782
rect 539579 685712 539709 685714
rect 540819 685714 540845 685782
rect 540845 685714 540919 685782
rect 540919 685714 540949 685782
rect 540819 685712 540949 685714
rect 542049 685714 542081 685782
rect 542081 685714 542155 685782
rect 542155 685714 542179 685782
rect 542049 685712 542179 685714
rect 543289 685714 543317 685782
rect 543317 685714 543391 685782
rect 543391 685714 543419 685782
rect 543289 685712 543419 685714
rect 544529 685714 544553 685782
rect 544553 685714 544627 685782
rect 544627 685714 544659 685782
rect 544529 685712 544659 685714
rect 545759 685714 545789 685782
rect 545789 685714 545863 685782
rect 545863 685714 545889 685782
rect 545759 685712 545889 685714
rect 546999 685714 547025 685782
rect 547025 685714 547099 685782
rect 547099 685714 547129 685782
rect 546999 685712 547129 685714
rect 548229 685714 548261 685782
rect 548261 685714 548335 685782
rect 548335 685714 548359 685782
rect 548229 685712 548359 685714
rect 549469 685714 549497 685782
rect 549497 685714 549571 685782
rect 549571 685714 549599 685782
rect 549469 685712 549599 685714
rect 538849 685652 538929 685662
rect 539059 685652 539139 685662
rect 543859 685652 543939 685662
rect 544049 685652 544129 685662
rect 538849 685582 538929 685652
rect 539059 685582 539139 685652
rect 541319 685572 541399 685652
rect 541559 685572 541639 685652
rect 543859 685582 543939 685652
rect 544049 685582 544129 685652
rect 546319 685572 546399 685652
rect 546509 685572 546589 685652
rect 548799 685562 548879 685642
rect 548969 685562 549049 685642
rect 535759 685122 535849 685252
rect 535969 685122 536059 685252
rect 553069 685152 553139 685242
rect 553229 685152 553299 685242
rect 540819 685064 540949 685132
rect 542049 685064 542179 685122
rect 542379 685064 542459 685132
rect 542489 685064 542569 685132
rect 543289 685064 543419 685122
rect 544529 685064 544659 685122
rect 544789 685064 544869 685132
rect 544899 685064 544979 685132
rect 545759 685064 545889 685122
rect 546999 685072 547129 685142
rect 547249 685064 547329 685142
rect 547359 685064 547439 685142
rect 548229 685064 548359 685122
rect 540819 685062 540949 685064
rect 542049 685052 542179 685064
rect 542379 685052 542459 685064
rect 542489 685052 542569 685064
rect 543289 685052 543419 685064
rect 544529 685052 544659 685064
rect 544789 685052 544869 685064
rect 544899 685052 544979 685064
rect 545759 685052 545889 685064
rect 547249 685062 547329 685064
rect 547359 685062 547439 685064
rect 548229 685052 548359 685064
rect 545769 684872 545859 684882
rect 545909 684872 545999 684882
rect 42260 684750 42370 684860
rect 42510 684750 42620 684860
rect 46660 684750 46770 684860
rect 46910 684750 47020 684860
rect 540759 684782 540849 684862
rect 540899 684782 540989 684862
rect 545769 684802 545859 684872
rect 545909 684802 545999 684872
rect 44530 684686 44780 684720
rect 44530 684470 44780 684686
rect 542279 684662 542389 684772
rect 543139 684662 543249 684772
rect 544349 684662 544459 684772
rect 545199 684662 545309 684772
rect 540759 684564 540849 684632
rect 540899 684564 540989 684632
rect 546769 684662 546879 684772
rect 547649 684662 547759 684772
rect 545769 684564 545859 684622
rect 545909 684564 545999 684622
rect 540759 684552 540849 684564
rect 540899 684552 540989 684564
rect 545769 684542 545859 684564
rect 545909 684542 545999 684564
rect 543579 684372 543659 684392
rect 543729 684372 543809 684392
rect 546059 684372 546139 684392
rect 546199 684372 546279 684392
rect 541089 684292 541169 684372
rect 541239 684292 541319 684372
rect 543579 684312 543659 684372
rect 543729 684312 543809 684372
rect 546059 684312 546139 684372
rect 546199 684312 546279 684372
rect 541539 684064 541619 684142
rect 541649 684064 541729 684142
rect 543949 684064 544029 684112
rect 546399 684064 546479 684132
rect 546519 684064 546599 684132
rect 547599 684064 547679 684122
rect 541539 684062 541619 684064
rect 541649 684062 541729 684064
rect 543949 684032 544029 684064
rect 546399 684052 546479 684064
rect 546519 684052 546599 684064
rect 547599 684042 547679 684064
rect 43840 683520 43860 683600
rect 43860 683520 43894 683600
rect 43894 683520 43920 683600
rect 44350 683520 44376 683600
rect 44376 683520 44410 683600
rect 44410 683520 44430 683600
rect 44090 683040 44118 683120
rect 44118 683040 44152 683120
rect 44152 683040 44170 683120
rect 44870 683520 44892 683600
rect 44892 683520 44926 683600
rect 44926 683520 44950 683600
rect 44610 683040 44634 683120
rect 44634 683040 44668 683120
rect 44668 683040 44690 683120
rect 45390 683520 45408 683600
rect 45408 683520 45442 683600
rect 45442 683520 45470 683600
rect 45130 683040 45150 683120
rect 45150 683040 45184 683120
rect 45184 683040 45210 683120
rect 542719 683882 542799 683962
rect 545129 683882 545209 683962
rect 541459 683772 541539 683782
rect 546349 683772 546429 683782
rect 541459 683702 541539 683772
rect 546349 683702 546429 683772
rect 541569 683562 541679 683652
rect 546479 683562 546589 683652
rect 543949 683444 544029 683492
rect 547599 683444 547679 683502
rect 543949 683412 544029 683444
rect 547599 683422 547679 683444
rect 542109 683262 542165 683342
rect 542165 683262 542199 683342
rect 542229 683262 542319 683342
rect 542719 683262 542799 683342
rect 544559 683262 544601 683342
rect 544601 683262 544635 683342
rect 544635 683262 544649 683342
rect 544679 683262 544769 683342
rect 545129 683262 545209 683342
rect 546989 683262 547037 683342
rect 547037 683262 547071 683342
rect 547071 683262 547079 683342
rect 547109 683262 547199 683342
rect 541459 683152 541539 683162
rect 546349 683152 546429 683162
rect 541459 683082 541539 683152
rect 546349 683082 546429 683152
rect 543339 682844 543429 682912
rect 548219 682852 548309 682932
rect 543339 682832 543429 682844
rect 43920 682738 43922 682770
rect 43922 682738 43990 682770
rect 43920 682700 43990 682738
rect 44620 682700 44690 682770
rect 45310 682738 45380 682770
rect 45310 682700 45380 682738
rect 542109 682662 542199 682742
rect 542229 682662 542319 682742
rect 544559 682662 544649 682742
rect 544679 682662 544769 682742
rect 546989 682662 547079 682742
rect 547109 682662 547199 682742
rect 540759 682552 540849 682582
rect 540899 682552 540989 682582
rect 545769 682552 545859 682582
rect 545909 682552 545999 682582
rect 540759 682502 540849 682552
rect 540899 682502 540989 682552
rect 545769 682502 545859 682552
rect 545909 682502 545999 682552
rect 43920 682400 43990 682440
rect 43920 682370 43922 682400
rect 43922 682370 43990 682400
rect 44620 682370 44690 682440
rect 45310 682400 45380 682440
rect 45310 682370 45380 682400
rect 43840 682060 43860 682140
rect 43860 682060 43894 682140
rect 43894 682060 43920 682140
rect 43630 681840 43710 681920
rect 43630 681700 43710 681780
rect 44350 682060 44376 682140
rect 44376 682060 44410 682140
rect 44410 682060 44430 682140
rect 541509 682352 541629 682452
rect 44870 682060 44892 682140
rect 44892 682060 44926 682140
rect 44926 682060 44950 682140
rect 542729 682352 542849 682452
rect 543939 682352 544059 682452
rect 543339 682244 543429 682312
rect 545159 682352 545279 682452
rect 546389 682342 546509 682442
rect 547599 682352 547719 682452
rect 548219 682252 548309 682332
rect 543339 682232 543429 682244
rect 45390 682060 45408 682140
rect 45408 682060 45442 682140
rect 45442 682060 45470 682140
rect 542109 682062 542199 682142
rect 542229 682062 542319 682142
rect 544420 682056 544508 682146
rect 544559 682062 544649 682142
rect 544679 682062 544769 682142
rect 546989 682062 547079 682142
rect 547109 682062 547199 682142
rect 561700 682000 561900 682200
rect 562100 682000 562300 682200
rect 562500 682000 562700 682200
rect 562900 682000 563100 682200
rect 563300 682000 563500 682200
rect 540759 681952 540849 681962
rect 540899 681952 540989 681962
rect 545769 681952 545859 681982
rect 545909 681952 545999 681982
rect 45590 681840 45670 681920
rect 540759 681882 540849 681952
rect 540899 681882 540989 681952
rect 545769 681902 545859 681952
rect 545909 681902 545999 681952
rect 45590 681700 45670 681780
rect 561700 681600 561900 681800
rect 562100 681600 562300 681800
rect 562500 681600 562700 681800
rect 562900 681600 563100 681800
rect 563300 681600 563500 681800
rect 541384 681318 541544 681478
rect 542444 681318 542604 681478
rect 543904 681318 544064 681478
rect 545124 681318 545284 681478
rect 546604 681318 546764 681478
rect 547604 681318 547764 681478
rect 43810 681170 43910 681270
rect 44600 681238 44606 681270
rect 44606 681238 44670 681270
rect 45360 681238 45380 681270
rect 45380 681238 45460 681270
rect 44600 681200 44670 681238
rect 45360 681170 45460 681238
rect 542884 681088 542954 681158
rect 543104 681088 543174 681158
rect 546064 681088 546134 681158
rect 546304 681088 546374 681158
rect 561700 681200 561900 681400
rect 562100 681200 562300 681400
rect 562500 681200 562700 681400
rect 562900 681200 563100 681400
rect 563300 681200 563500 681400
rect 44600 680760 44670 680830
rect 44270 680400 44340 680520
rect 44340 680400 44380 680520
rect 44380 680400 44390 680520
rect 44600 680290 44618 680360
rect 44618 680290 44652 680360
rect 44652 680290 44670 680360
rect 541384 680738 541544 680898
rect 542444 680738 542604 680898
rect 543904 680738 544064 680898
rect 545124 680738 545284 680898
rect 546604 680738 546764 680898
rect 547604 680738 547764 680898
rect 561700 680800 561900 681000
rect 562100 680800 562300 681000
rect 562500 680800 562700 681000
rect 562900 680800 563100 681000
rect 563300 680800 563500 681000
rect 44890 680410 44930 680530
rect 44930 680410 45010 680530
rect 542884 680498 542954 680568
rect 543104 680498 543174 680568
rect 546064 680498 546134 680568
rect 546304 680498 546374 680568
rect 544044 680388 544114 680408
rect 544154 680388 544224 680408
rect 544984 680388 545054 680408
rect 545094 680388 545164 680408
rect 544044 680338 544114 680388
rect 544154 680338 544224 680388
rect 544984 680338 545054 680388
rect 545094 680338 545164 680388
rect 561700 680400 561900 680600
rect 562100 680400 562300 680600
rect 562500 680400 562700 680600
rect 562900 680400 563100 680600
rect 563300 680400 563500 680600
rect 561700 680000 561900 680200
rect 562100 680000 562300 680200
rect 562500 680000 562700 680200
rect 562900 680000 563100 680200
rect 563300 680000 563500 680200
rect 544410 679890 544470 679926
rect 544410 679866 544470 679890
rect 544510 679866 544570 679926
rect 544610 679866 544670 679926
rect 544710 679890 544770 679926
rect 544710 679866 544722 679890
rect 544722 679866 544770 679890
rect 44090 679782 44170 679830
rect 44090 679750 44162 679782
rect 44162 679750 44170 679782
rect 44600 679760 44670 679830
rect 45130 679750 45210 679830
rect 544044 679828 544114 679838
rect 44070 679540 44100 679630
rect 44100 679540 44134 679630
rect 44134 679540 44160 679630
rect 44590 679540 44616 679630
rect 44616 679540 44650 679630
rect 44650 679540 44680 679630
rect 544044 679768 544062 679828
rect 544062 679768 544096 679828
rect 544096 679768 544114 679828
rect 544154 679828 544224 679838
rect 544984 679828 545054 679848
rect 544154 679768 544170 679828
rect 544170 679768 544204 679828
rect 544204 679768 544224 679828
rect 544984 679778 544998 679828
rect 544998 679778 545032 679828
rect 545032 679778 545054 679828
rect 545094 679828 545164 679848
rect 545094 679778 545106 679828
rect 545106 679778 545140 679828
rect 545140 679778 545164 679828
rect 45100 679540 45132 679630
rect 45132 679540 45166 679630
rect 45166 679540 45190 679630
rect 561700 679600 561900 679800
rect 562100 679600 562300 679800
rect 562500 679600 562700 679800
rect 562900 679600 563100 679800
rect 563300 679600 563500 679800
rect 44220 679388 44280 679420
rect 44990 679388 45050 679420
rect 44220 679360 44280 679388
rect 44990 679360 45050 679388
rect 543764 679368 543984 679518
rect 544284 679368 544504 679518
rect 544704 679368 544924 679518
rect 545254 679368 545474 679518
rect 44580 679160 44670 679250
rect 542884 679238 542954 679308
rect 543094 679238 543164 679308
rect 546064 679258 546134 679328
rect 546304 679258 546374 679328
rect 542884 679148 542954 679218
rect 543094 679148 543164 679218
rect 546064 679168 546134 679238
rect 546304 679168 546374 679238
rect 561700 679200 561900 679400
rect 562100 679200 562300 679400
rect 562500 679200 562700 679400
rect 562900 679200 563100 679400
rect 563300 679200 563500 679400
rect 544044 679073 544114 679088
rect 544154 679073 544224 679088
rect 544984 679073 545054 679088
rect 545094 679073 545164 679088
rect 44220 679032 44280 679060
rect 44990 679032 45050 679060
rect 44220 679000 44280 679032
rect 44990 679000 45050 679032
rect 544044 679018 544114 679073
rect 544154 679018 544224 679073
rect 544984 679018 545054 679073
rect 545094 679018 545164 679073
rect 43830 678630 43845 678690
rect 43845 678630 43879 678690
rect 43879 678630 43890 678690
rect 44350 678630 44361 678690
rect 44361 678630 44395 678690
rect 44395 678630 44410 678690
rect 44090 678220 44103 678280
rect 44103 678220 44137 678280
rect 44137 678220 44150 678280
rect 44830 678610 44877 678720
rect 44877 678610 44911 678720
rect 44911 678610 44960 678720
rect 44610 678220 44619 678280
rect 44619 678220 44653 678280
rect 44653 678220 44670 678280
rect 45380 678630 45393 678690
rect 45393 678630 45427 678690
rect 45427 678630 45440 678690
rect 45120 678220 45135 678280
rect 45135 678220 45169 678280
rect 45169 678220 45180 678280
rect 541404 678828 541584 678958
rect 542544 678828 542724 678958
rect 543524 678838 543704 678968
rect 544294 678838 544474 678968
rect 544734 678838 544914 678968
rect 545454 678828 545634 678958
rect 546524 678838 546704 678968
rect 547524 678838 547704 678968
rect 561700 678800 561900 679000
rect 562100 678800 562300 679000
rect 562500 678800 562700 679000
rect 562900 678800 563100 679000
rect 563300 678800 563500 679000
rect 542884 678740 542954 678788
rect 543104 678740 543174 678788
rect 546064 678740 546134 678788
rect 546304 678740 546374 678788
rect 542884 678718 542954 678740
rect 543104 678718 543174 678740
rect 546064 678718 546134 678740
rect 546304 678718 546374 678740
rect 544044 678568 544114 678638
rect 544154 678568 544224 678638
rect 544984 678568 545054 678638
rect 545094 678568 545164 678638
rect 561700 678400 561900 678600
rect 562100 678400 562300 678600
rect 562500 678400 562700 678600
rect 562900 678400 563100 678600
rect 563300 678400 563500 678600
rect 44580 677780 44670 677810
rect 44580 677720 44670 677780
rect 44090 677526 44150 677530
rect 45120 677526 45180 677530
rect 44090 677470 44150 677526
rect 44090 677300 44150 677360
rect 44090 677130 44150 677190
rect 45120 677470 45180 677526
rect 45120 677300 45180 677360
rect 45120 677130 45180 677190
rect 41200 676740 41440 676980
rect 47900 676740 48140 676980
rect 541364 676938 541484 677058
rect 547734 676938 547854 677058
rect 41200 675020 41440 675260
rect 47900 675020 48140 675260
rect 541364 673938 541484 674058
rect 547734 673938 547854 674058
rect 41200 673300 41440 673540
rect 47900 673300 48140 673540
rect 41200 671820 41440 672060
rect 47900 671820 48140 672060
rect 541364 670938 541484 671058
rect 547734 670938 547854 671058
rect 41200 670100 41440 670340
rect 47900 670100 48140 670340
rect 41200 668500 41440 668740
rect 47900 668500 48140 668740
rect 541364 667938 541484 668058
rect 547734 667938 547854 668058
rect 41200 666780 41440 667020
rect 47900 666780 48140 667020
rect 41200 665180 41440 665420
rect 47900 665180 48140 665420
rect 541364 664938 541484 665058
rect 547734 664938 547854 665058
rect 41200 663460 41440 663700
rect 47900 663460 48140 663700
rect 32800 663000 33100 663300
rect 33300 663000 33600 663300
rect 33800 663000 34100 663300
rect 34300 663000 34600 663300
rect 34800 663000 35100 663300
rect 35300 663000 35600 663300
rect 35800 663000 36100 663300
rect 36300 663000 36600 663300
rect 36800 663000 37100 663300
rect 37300 663000 37600 663300
rect 37800 663000 38100 663300
rect 38300 663000 38600 663300
rect 38800 663000 39100 663300
rect 39300 663000 39600 663300
rect 39800 663000 40100 663300
rect 40300 663000 40600 663300
rect 541744 663356 541777 663728
rect 541777 663356 542891 663728
rect 542891 663356 542914 663728
rect 541744 663318 542914 663356
rect 543254 663356 543297 663728
rect 543297 663356 544411 663728
rect 544411 663356 544424 663728
rect 543254 663318 544424 663356
rect 544774 663362 544807 663728
rect 544807 663362 545921 663728
rect 545921 663362 545944 663728
rect 544774 663318 545944 663362
rect 546294 663362 546317 663738
rect 546317 663362 547431 663738
rect 547431 663362 547464 663738
rect 546294 663328 547464 663362
rect 41200 662980 41440 663220
rect 47900 662980 48140 663220
<< metal2 >>
rect 44010 695640 44280 695650
rect 44010 695360 44280 695370
rect 45060 695640 45330 695650
rect 45060 695360 45330 695370
rect 41460 695160 41530 695170
rect 41460 695080 41530 695090
rect 41780 695160 41850 695170
rect 41780 695080 41850 695090
rect 42090 695160 42160 695170
rect 42090 695080 42160 695090
rect 42410 695160 42480 695170
rect 42410 695080 42480 695090
rect 42720 695160 42790 695170
rect 42720 695080 42790 695090
rect 43040 695160 43110 695170
rect 43040 695080 43110 695090
rect 43360 695160 43430 695170
rect 43360 695080 43430 695090
rect 43670 695160 43740 695170
rect 43670 695080 43740 695090
rect 43990 695160 44060 695170
rect 43990 695080 44060 695090
rect 44310 695160 44380 695170
rect 44310 695080 44380 695090
rect 44620 695160 44690 695170
rect 44620 695080 44690 695090
rect 44940 695160 45010 695170
rect 44940 695080 45010 695090
rect 45250 695160 45320 695170
rect 45250 695080 45320 695090
rect 45570 695160 45640 695170
rect 45570 695080 45640 695090
rect 45890 695160 45960 695170
rect 45890 695080 45960 695090
rect 46200 695160 46270 695170
rect 46200 695080 46270 695090
rect 46520 695160 46590 695170
rect 46520 695080 46590 695090
rect 46830 695160 46900 695170
rect 46830 695080 46900 695090
rect 47150 695160 47220 695170
rect 47150 695080 47220 695090
rect 47470 695160 47540 695170
rect 47470 695080 47540 695090
rect 47780 695160 47850 695170
rect 47780 695080 47850 695090
rect 36800 694920 37020 694940
rect 36800 694850 36930 694920
rect 37000 694850 37020 694920
rect 36800 694810 37020 694850
rect 41460 694920 41530 694930
rect 41460 694840 41530 694850
rect 41780 694920 41850 694930
rect 41780 694840 41850 694850
rect 42090 694920 42160 694930
rect 42090 694840 42160 694850
rect 42410 694920 42480 694930
rect 42410 694840 42480 694850
rect 42720 694920 42790 694930
rect 42720 694840 42790 694850
rect 43040 694920 43110 694930
rect 43040 694840 43110 694850
rect 43360 694920 43430 694930
rect 43360 694840 43430 694850
rect 43670 694920 43740 694930
rect 43670 694840 43740 694850
rect 43990 694920 44060 694930
rect 43990 694840 44060 694850
rect 44310 694920 44380 694930
rect 44310 694840 44380 694850
rect 44620 694920 44690 694930
rect 44620 694840 44690 694850
rect 44940 694920 45010 694930
rect 44940 694840 45010 694850
rect 45250 694920 45320 694930
rect 45250 694840 45320 694850
rect 45570 694920 45640 694930
rect 45570 694840 45640 694850
rect 45890 694920 45960 694930
rect 45890 694840 45960 694850
rect 46200 694920 46270 694930
rect 46200 694840 46270 694850
rect 46520 694920 46590 694930
rect 46520 694840 46590 694850
rect 46830 694920 46900 694930
rect 46830 694840 46900 694850
rect 47150 694920 47220 694930
rect 47150 694840 47220 694850
rect 47470 694920 47540 694930
rect 47470 694840 47540 694850
rect 47780 694920 47850 694930
rect 47780 694840 47850 694850
rect 52300 694920 52520 694940
rect 52300 694850 52320 694920
rect 52390 694850 52520 694920
rect 36800 694740 36820 694810
rect 36890 694740 37020 694810
rect 36800 694720 37020 694740
rect 52300 694810 52520 694850
rect 52300 694740 52430 694810
rect 52500 694740 52520 694810
rect 52300 694720 52520 694740
rect 41590 694550 41720 694560
rect 41590 694480 41620 694550
rect 41690 694480 41720 694550
rect 41590 694310 41720 694480
rect 41930 694550 42000 694560
rect 41930 694470 42000 694480
rect 42250 694550 42320 694560
rect 42250 694470 42320 694480
rect 42570 694550 42640 694560
rect 42570 694470 42640 694480
rect 42880 694550 42950 694560
rect 42880 694470 42950 694480
rect 43200 694550 43270 694560
rect 43200 694470 43270 694480
rect 43510 694550 43580 694560
rect 43510 694470 43580 694480
rect 43830 694550 43900 694560
rect 43830 694470 43900 694480
rect 44150 694550 44220 694560
rect 44150 694470 44220 694480
rect 44460 694550 44530 694560
rect 44460 694470 44530 694480
rect 44780 694550 44850 694560
rect 44780 694470 44850 694480
rect 45100 694550 45170 694560
rect 45100 694470 45170 694480
rect 45410 694550 45480 694560
rect 45410 694470 45480 694480
rect 45730 694550 45800 694560
rect 45730 694470 45800 694480
rect 46040 694550 46110 694560
rect 46040 694470 46110 694480
rect 46360 694550 46430 694560
rect 46360 694470 46430 694480
rect 46680 694550 46750 694560
rect 46680 694470 46750 694480
rect 46990 694550 47060 694560
rect 46990 694470 47060 694480
rect 47310 694550 47380 694560
rect 47310 694470 47380 694480
rect 47600 694550 47730 694560
rect 47600 694480 47630 694550
rect 47700 694480 47730 694550
rect 41590 694240 41620 694310
rect 41690 694240 41720 694310
rect 41590 693940 41720 694240
rect 41930 694310 42000 694320
rect 41930 694230 42000 694240
rect 42250 694310 42320 694320
rect 42250 694230 42320 694240
rect 42570 694310 42640 694320
rect 42570 694230 42640 694240
rect 42880 694310 42950 694320
rect 42880 694230 42950 694240
rect 43200 694310 43270 694320
rect 43200 694230 43270 694240
rect 43510 694310 43580 694320
rect 43510 694230 43580 694240
rect 43830 694310 43900 694320
rect 43830 694230 43900 694240
rect 44150 694310 44220 694320
rect 44150 694230 44220 694240
rect 44460 694310 44530 694320
rect 44460 694230 44530 694240
rect 44780 694310 44850 694320
rect 44780 694230 44850 694240
rect 45100 694310 45170 694320
rect 45100 694230 45170 694240
rect 45410 694310 45480 694320
rect 45410 694230 45480 694240
rect 45730 694310 45800 694320
rect 45730 694230 45800 694240
rect 46040 694310 46110 694320
rect 46040 694230 46110 694240
rect 46360 694310 46430 694320
rect 46360 694230 46430 694240
rect 46680 694310 46750 694320
rect 46680 694230 46750 694240
rect 46990 694310 47060 694320
rect 46990 694230 47060 694240
rect 47310 694310 47380 694320
rect 47310 694230 47380 694240
rect 47600 694310 47730 694480
rect 47600 694240 47630 694310
rect 47700 694240 47730 694310
rect 41590 693870 41620 693940
rect 41690 693870 41720 693940
rect 38700 693460 38880 693470
rect 38700 693350 38880 693360
rect 39120 693460 39300 693470
rect 39120 693350 39300 693360
rect 41590 687330 41720 693870
rect 42540 694140 42700 694160
rect 42540 694060 42580 694140
rect 42660 694060 42700 694140
rect 42540 692840 42700 694060
rect 46600 694140 46760 694160
rect 46600 694060 46640 694140
rect 46720 694060 46760 694140
rect 44010 694000 44280 694010
rect 44010 693720 44280 693730
rect 45060 694000 45330 694010
rect 45060 693720 45330 693730
rect 42960 693490 43030 693500
rect 42960 693410 43030 693420
rect 43280 693490 43350 693500
rect 43280 693410 43350 693420
rect 43590 693490 43660 693500
rect 43590 693410 43660 693420
rect 43910 693490 43980 693500
rect 43910 693410 43980 693420
rect 44230 693490 44300 693500
rect 44230 693410 44300 693420
rect 44540 693490 44610 693500
rect 44540 693410 44610 693420
rect 44860 693490 44930 693500
rect 44860 693410 44930 693420
rect 45180 693490 45250 693500
rect 45180 693410 45250 693420
rect 45490 693490 45560 693500
rect 45490 693410 45560 693420
rect 45810 693490 45880 693500
rect 45810 693410 45880 693420
rect 46120 693490 46190 693500
rect 46120 693410 46190 693420
rect 42960 693280 43030 693290
rect 42960 693200 43030 693210
rect 43280 693280 43350 693290
rect 43280 693200 43350 693210
rect 43590 693280 43660 693290
rect 43590 693200 43660 693210
rect 43910 693280 43980 693290
rect 43910 693200 43980 693210
rect 44230 693280 44300 693290
rect 44230 693200 44300 693210
rect 44540 693280 44610 693290
rect 44540 693200 44610 693210
rect 44860 693280 44930 693290
rect 44860 693200 44930 693210
rect 45180 693280 45250 693290
rect 45180 693200 45250 693210
rect 45490 693280 45560 693290
rect 45490 693200 45560 693210
rect 45810 693280 45880 693290
rect 45810 693200 45880 693210
rect 46120 693280 46190 693290
rect 46120 693200 46190 693210
rect 42540 692760 42580 692840
rect 42660 692760 42700 692840
rect 43120 692850 43190 692860
rect 43120 692770 43190 692780
rect 43440 692850 43510 692860
rect 43440 692770 43510 692780
rect 43750 692850 43820 692860
rect 43750 692770 43820 692780
rect 44070 692850 44140 692860
rect 44070 692770 44140 692780
rect 44390 692850 44460 692860
rect 44390 692770 44460 692780
rect 44700 692850 44770 692860
rect 44700 692770 44770 692780
rect 45020 692850 45090 692860
rect 45020 692770 45090 692780
rect 45330 692850 45400 692860
rect 45330 692770 45400 692780
rect 45650 692850 45720 692860
rect 45650 692770 45720 692780
rect 45970 692850 46040 692860
rect 45970 692770 46040 692780
rect 46280 692850 46350 692860
rect 46280 692770 46350 692780
rect 46600 692840 46760 694060
rect 42540 692660 42700 692760
rect 42540 692580 42580 692660
rect 42660 692580 42700 692660
rect 46600 692760 46640 692840
rect 46720 692760 46760 692840
rect 46600 692660 46760 692760
rect 42540 690370 42700 692580
rect 43120 692640 43190 692650
rect 43120 692560 43190 692570
rect 43440 692640 43510 692650
rect 43440 692560 43510 692570
rect 43750 692640 43820 692650
rect 43750 692560 43820 692570
rect 44070 692640 44140 692650
rect 44070 692560 44140 692570
rect 44390 692640 44460 692650
rect 44390 692560 44460 692570
rect 44700 692640 44770 692650
rect 44700 692560 44770 692570
rect 45020 692640 45090 692650
rect 45020 692560 45090 692570
rect 45330 692640 45400 692650
rect 45330 692560 45400 692570
rect 45650 692640 45720 692650
rect 45650 692560 45720 692570
rect 45970 692640 46040 692650
rect 45970 692560 46040 692570
rect 46280 692640 46350 692650
rect 46280 692560 46350 692570
rect 46600 692580 46640 692660
rect 46720 692580 46760 692660
rect 43780 692390 44040 692400
rect 43780 692120 44040 692130
rect 45280 692390 45540 692400
rect 45280 692120 45540 692130
rect 42960 691940 43030 691950
rect 42960 691860 43030 691870
rect 43280 691940 43350 691950
rect 43280 691860 43350 691870
rect 43590 691940 43660 691950
rect 43590 691860 43660 691870
rect 43910 691940 43980 691950
rect 43910 691860 43980 691870
rect 44230 691940 44300 691950
rect 44230 691860 44300 691870
rect 44540 691940 44610 691950
rect 44540 691860 44610 691870
rect 44860 691940 44930 691950
rect 44860 691860 44930 691870
rect 45170 691940 45240 691950
rect 45170 691860 45240 691870
rect 45490 691940 45560 691950
rect 45490 691860 45560 691870
rect 45810 691940 45880 691950
rect 45810 691860 45880 691870
rect 46120 691940 46190 691950
rect 46120 691860 46190 691870
rect 42960 691730 43030 691740
rect 42960 691650 43030 691660
rect 43280 691730 43350 691740
rect 43280 691650 43350 691660
rect 43590 691730 43660 691740
rect 43590 691650 43660 691660
rect 43910 691730 43980 691740
rect 43910 691650 43980 691660
rect 44230 691730 44300 691740
rect 44230 691650 44300 691660
rect 44540 691730 44610 691740
rect 44540 691650 44610 691660
rect 44860 691730 44930 691740
rect 44860 691650 44930 691660
rect 45170 691730 45240 691740
rect 45170 691650 45240 691660
rect 45490 691730 45560 691740
rect 45490 691650 45560 691660
rect 45810 691730 45880 691740
rect 45810 691650 45880 691660
rect 46120 691730 46190 691740
rect 46120 691650 46190 691660
rect 43120 691310 43190 691320
rect 43120 691230 43190 691240
rect 43410 691310 43540 691320
rect 43410 691240 43440 691310
rect 43510 691240 43540 691310
rect 43120 691100 43190 691110
rect 43120 691020 43190 691030
rect 43410 691100 43540 691240
rect 43750 691310 43820 691320
rect 43750 691230 43820 691240
rect 44070 691310 44140 691320
rect 44070 691230 44140 691240
rect 44380 691310 44450 691320
rect 44380 691230 44450 691240
rect 44700 691310 44770 691320
rect 44700 691230 44770 691240
rect 45020 691310 45090 691320
rect 45020 691230 45090 691240
rect 45330 691310 45400 691320
rect 45330 691230 45400 691240
rect 45650 691310 45720 691320
rect 45650 691230 45720 691240
rect 45930 691310 46060 691320
rect 45930 691240 45960 691310
rect 46030 691240 46060 691310
rect 43410 691030 43440 691100
rect 43510 691030 43540 691100
rect 42540 690250 42560 690370
rect 42680 690250 42700 690370
rect 42540 690150 42700 690250
rect 42540 690030 42560 690150
rect 42680 690030 42700 690150
rect 42540 690010 42700 690030
rect 42780 689810 42940 689830
rect 42780 689690 42800 689810
rect 42920 689690 42940 689810
rect 42780 689590 42940 689690
rect 42780 689470 42800 689590
rect 42920 689470 42940 689590
rect 42780 688850 42940 689470
rect 42780 688730 42800 688850
rect 42920 688730 42940 688850
rect 42000 688700 42100 688710
rect 42000 688590 42100 688600
rect 42780 688630 42940 688730
rect 42780 688510 42800 688630
rect 42920 688510 42940 688630
rect 42000 688500 42100 688510
rect 42000 688290 42100 688300
rect 42000 688200 42100 688210
rect 42000 688090 42100 688100
rect 41590 687260 41620 687330
rect 41690 687260 41720 687330
rect 41590 687170 41720 687260
rect 41590 687100 41620 687170
rect 41690 687100 41720 687170
rect 41590 687080 41720 687100
rect 42240 687490 42640 687610
rect 42240 687380 42260 687490
rect 42370 687380 42510 687490
rect 42620 687380 42640 687490
rect 42240 686380 42640 687380
rect 42240 686270 42260 686380
rect 42370 686270 42510 686380
rect 42620 686270 42640 686380
rect 42240 685970 42640 686270
rect 42240 685860 42260 685970
rect 42370 685860 42510 685970
rect 42620 685860 42640 685970
rect 42240 684860 42640 685860
rect 42780 685820 42940 688510
rect 43410 688280 43540 691030
rect 43750 691100 43820 691110
rect 43750 691020 43820 691030
rect 44070 691100 44140 691110
rect 44070 691020 44140 691030
rect 44380 691100 44450 691110
rect 44380 691020 44450 691030
rect 44700 691100 44770 691110
rect 44700 691020 44770 691030
rect 45020 691100 45090 691110
rect 45020 691020 45090 691030
rect 45330 691100 45400 691110
rect 45330 691020 45400 691030
rect 45650 691100 45720 691110
rect 45650 691020 45720 691030
rect 45930 691100 46060 691240
rect 46280 691310 46350 691320
rect 46280 691230 46350 691240
rect 45930 691030 45960 691100
rect 46030 691030 46060 691100
rect 44060 690380 44130 690390
rect 44060 690300 44130 690310
rect 44380 690380 44450 690390
rect 44380 690300 44450 690310
rect 44690 690380 44760 690390
rect 44690 690300 44760 690310
rect 45010 690380 45080 690390
rect 45010 690300 45080 690310
rect 44060 690090 44130 690100
rect 44060 690010 44130 690020
rect 44380 690090 44450 690100
rect 44380 690010 44450 690020
rect 44690 690090 44760 690100
rect 44690 690010 44760 690020
rect 45010 690090 45080 690100
rect 45010 690010 45080 690020
rect 44220 689820 44290 689830
rect 44220 689740 44290 689750
rect 44530 689820 44600 689830
rect 44530 689740 44600 689750
rect 44850 689820 44920 689830
rect 44850 689740 44920 689750
rect 45170 689820 45240 689830
rect 45170 689740 45240 689750
rect 44220 689530 44290 689540
rect 44220 689450 44290 689460
rect 44530 689530 44600 689540
rect 44530 689450 44600 689460
rect 44850 689530 44920 689540
rect 44850 689450 44920 689460
rect 45170 689530 45240 689540
rect 45170 689450 45240 689460
rect 44520 689290 44780 689300
rect 44520 689020 44780 689030
rect 44060 688860 44130 688870
rect 44060 688780 44130 688790
rect 44380 688860 44450 688870
rect 44380 688780 44450 688790
rect 44690 688860 44760 688870
rect 44690 688780 44760 688790
rect 45010 688860 45080 688870
rect 45010 688780 45080 688790
rect 44060 688570 44130 688580
rect 44060 688490 44130 688500
rect 44380 688570 44450 688580
rect 44380 688490 44450 688500
rect 44690 688570 44760 688580
rect 44690 688490 44760 688500
rect 45010 688570 45080 688580
rect 45010 688490 45080 688500
rect 43410 688210 43440 688280
rect 43510 688210 43540 688280
rect 44220 688300 44290 688310
rect 44220 688220 44290 688230
rect 44530 688300 44600 688310
rect 44530 688220 44600 688230
rect 44850 688300 44920 688310
rect 44850 688220 44920 688230
rect 45170 688300 45240 688310
rect 45170 688220 45240 688230
rect 45930 688280 46060 691030
rect 46280 691100 46350 691110
rect 46280 691020 46350 691030
rect 46600 690370 46760 692580
rect 46600 690250 46620 690370
rect 46740 690250 46760 690370
rect 47600 693940 47730 694240
rect 47600 693870 47630 693940
rect 47700 693870 47730 693940
rect 46600 690150 46760 690250
rect 47200 690300 47300 690310
rect 47200 690190 47300 690200
rect 46600 690030 46620 690150
rect 46740 690030 46760 690150
rect 46600 690010 46760 690030
rect 47200 690000 47300 690010
rect 43410 688030 43540 688210
rect 43410 687960 43440 688030
rect 43510 687960 43540 688030
rect 45930 688210 45960 688280
rect 46030 688210 46060 688280
rect 45930 688030 46060 688210
rect 43410 687930 43540 687960
rect 44220 688010 44290 688020
rect 44220 687930 44290 687940
rect 44530 688010 44600 688020
rect 44530 687930 44600 687940
rect 44850 688010 44920 688020
rect 44850 687930 44920 687940
rect 45170 688010 45240 688020
rect 45170 687930 45240 687940
rect 45930 687960 45960 688030
rect 46030 687960 46060 688030
rect 45930 687930 46060 687960
rect 46360 689810 46520 689830
rect 46360 689690 46380 689810
rect 46500 689690 46520 689810
rect 47200 689790 47300 689800
rect 46360 689590 46520 689690
rect 46360 689470 46380 689590
rect 46500 689470 46520 689590
rect 47200 689600 47300 689610
rect 47200 689490 47300 689500
rect 46360 688850 46520 689470
rect 46360 688730 46380 688850
rect 46500 688730 46520 688850
rect 46360 688630 46520 688730
rect 46360 688510 46380 688630
rect 46500 688510 46520 688630
rect 44520 687770 44780 687780
rect 44520 687500 44780 687510
rect 43070 687340 43140 687350
rect 43070 687260 43140 687270
rect 43590 687340 43660 687350
rect 43590 687260 43660 687270
rect 44100 687340 44170 687350
rect 44100 687260 44170 687270
rect 44620 687340 44690 687350
rect 44620 687260 44690 687270
rect 45130 687340 45200 687350
rect 45130 687260 45200 687270
rect 45650 687340 45720 687350
rect 45650 687260 45720 687270
rect 46170 687340 46240 687350
rect 46170 687260 46240 687270
rect 43070 687160 43140 687170
rect 43070 687080 43140 687090
rect 43590 687160 43660 687170
rect 43590 687080 43660 687090
rect 44100 687160 44170 687170
rect 44100 687080 44170 687090
rect 44620 687160 44690 687170
rect 44620 687080 44690 687090
rect 45130 687160 45200 687170
rect 45130 687080 45200 687090
rect 45650 687160 45720 687170
rect 45650 687080 45720 687090
rect 46170 687160 46240 687170
rect 46170 687080 46240 687090
rect 43330 686670 43400 686680
rect 43330 686590 43400 686600
rect 43840 686670 43910 686680
rect 43840 686590 43910 686600
rect 44360 686670 44430 686680
rect 44360 686590 44430 686600
rect 44880 686670 44950 686680
rect 44880 686590 44950 686600
rect 45390 686670 45460 686680
rect 45390 686590 45460 686600
rect 45910 686670 45980 686680
rect 45910 686590 45980 686600
rect 43330 686490 43400 686500
rect 43330 686410 43400 686420
rect 43840 686490 43910 686500
rect 43840 686410 43910 686420
rect 44360 686490 44430 686500
rect 44360 686410 44430 686420
rect 44880 686490 44950 686500
rect 44880 686410 44950 686420
rect 45390 686490 45460 686500
rect 45390 686410 45460 686420
rect 45910 686490 45980 686500
rect 45910 686410 45980 686420
rect 44530 686250 44780 686260
rect 44530 685990 44780 686000
rect 42780 685750 42810 685820
rect 42880 685750 42940 685820
rect 42780 685640 42940 685750
rect 43330 685820 43400 685830
rect 43330 685740 43400 685750
rect 43840 685820 43910 685830
rect 43840 685740 43910 685750
rect 44360 685820 44430 685830
rect 44360 685740 44430 685750
rect 44870 685820 44940 685830
rect 44870 685740 44940 685750
rect 45390 685820 45460 685830
rect 45390 685740 45460 685750
rect 45910 685820 45980 685830
rect 45910 685740 45980 685750
rect 46360 685820 46520 688510
rect 46360 685750 46420 685820
rect 46490 685750 46520 685820
rect 42780 685570 42810 685640
rect 42880 685570 42940 685640
rect 42780 685560 42940 685570
rect 43330 685640 43400 685650
rect 43330 685560 43400 685570
rect 43840 685640 43910 685650
rect 43840 685560 43910 685570
rect 44360 685640 44430 685650
rect 44360 685560 44430 685570
rect 44870 685640 44940 685650
rect 44870 685560 44940 685570
rect 45390 685640 45460 685650
rect 45390 685560 45460 685570
rect 45910 685640 45980 685650
rect 45910 685560 45980 685570
rect 46360 685640 46520 685750
rect 46360 685570 46420 685640
rect 46490 685570 46520 685640
rect 46360 685560 46520 685570
rect 46640 687490 47040 687610
rect 46640 687380 46660 687490
rect 46770 687380 46910 687490
rect 47020 687380 47040 687490
rect 46640 686380 47040 687380
rect 47600 687330 47730 693870
rect 49950 693460 50130 693470
rect 49950 693350 50130 693360
rect 50370 693460 50550 693470
rect 50370 693350 50550 693360
rect 541949 690962 542239 690982
rect 541949 690892 541969 690962
rect 542059 690892 542139 690962
rect 542229 690892 542239 690962
rect 541949 690852 542239 690892
rect 541949 690772 541969 690852
rect 542049 690772 542139 690852
rect 542219 690772 542239 690852
rect 544439 690962 544729 690982
rect 544439 690892 544459 690962
rect 544549 690892 544629 690962
rect 544719 690892 544729 690962
rect 544439 690852 544729 690892
rect 540679 690612 540969 690732
rect 541409 690722 541559 690772
rect 540679 690532 540699 690612
rect 540779 690532 540869 690612
rect 540949 690532 540969 690612
rect 541089 690682 541169 690692
rect 541089 690592 541169 690602
rect 541239 690682 541319 690692
rect 541239 690592 541319 690602
rect 541409 690652 541419 690722
rect 541549 690652 541559 690722
rect 540679 690072 540969 690532
rect 541409 690182 541559 690652
rect 540679 689992 540699 690072
rect 540779 689992 540869 690072
rect 540949 689992 540969 690072
rect 541089 690142 541169 690152
rect 541089 690052 541169 690062
rect 541239 690142 541319 690152
rect 541239 690052 541319 690062
rect 541409 690112 541419 690182
rect 541549 690112 541559 690182
rect 540679 689532 540969 689992
rect 541409 689642 541559 690112
rect 541949 690312 542239 690772
rect 541949 690232 541969 690312
rect 542049 690232 542139 690312
rect 542219 690232 542239 690312
rect 541949 689912 542239 690232
rect 541949 689842 541979 689912
rect 542069 689842 542119 689912
rect 542209 689842 542239 689912
rect 541949 689772 542239 689842
rect 541949 689692 541969 689772
rect 542049 689692 542139 689772
rect 542219 689692 542239 689772
rect 541949 689682 542239 689692
rect 542649 690722 542799 690782
rect 542649 690652 542659 690722
rect 542789 690652 542799 690722
rect 542649 690182 542799 690652
rect 542649 690112 542659 690182
rect 542789 690112 542799 690182
rect 540679 689452 540699 689532
rect 540779 689452 540869 689532
rect 540949 689452 540969 689532
rect 541089 689602 541169 689612
rect 541089 689512 541169 689522
rect 541239 689602 541319 689612
rect 541239 689512 541319 689522
rect 541409 689572 541419 689642
rect 541549 689572 541559 689642
rect 540679 689432 540969 689452
rect 541409 689102 541559 689572
rect 542649 689642 542799 690112
rect 542649 689572 542659 689642
rect 542789 689572 542799 689642
rect 541979 689382 542059 689392
rect 541979 689292 542059 689302
rect 542149 689382 542229 689392
rect 542149 689292 542229 689302
rect 541409 689032 541419 689102
rect 541549 689032 541559 689102
rect 540679 688992 540969 689022
rect 540679 688912 540699 688992
rect 540779 688912 540869 688992
rect 540949 688912 540969 688992
rect 540679 688412 540969 688912
rect 540679 688332 540699 688412
rect 540779 688332 540869 688412
rect 540949 688332 540969 688412
rect 534629 688132 534759 688142
rect 534629 687982 534759 687992
rect 534879 688132 535009 688142
rect 534879 687982 535009 687992
rect 540679 687802 540969 688332
rect 541409 688522 541559 689032
rect 541409 688452 541419 688522
rect 541549 688452 541559 688522
rect 541409 687942 541559 688452
rect 541959 689252 542249 689292
rect 541959 689172 541979 689252
rect 542059 689172 542149 689252
rect 542229 689172 542249 689252
rect 541959 688672 542249 689172
rect 542649 689102 542799 689572
rect 543199 690612 543489 690812
rect 544439 690772 544459 690852
rect 544539 690772 544629 690852
rect 544709 690772 544729 690852
rect 546899 690972 547189 691012
rect 546899 690892 546919 690972
rect 546999 690892 547089 690972
rect 547169 690892 547189 690972
rect 566290 690900 566300 691100
rect 566500 690900 566510 691100
rect 566690 690900 566700 691100
rect 566900 690900 566910 691100
rect 567090 690900 567100 691100
rect 567300 690900 567310 691100
rect 567490 690900 567500 691100
rect 567700 690900 567710 691100
rect 567890 690900 567900 691100
rect 568100 690900 568110 691100
rect 568290 690900 568300 691100
rect 568500 690900 568510 691100
rect 568690 690900 568700 691100
rect 568900 690900 568910 691100
rect 569090 690900 569100 691100
rect 569300 690900 569310 691100
rect 569490 690900 569500 691100
rect 569700 690900 569710 691100
rect 569890 690900 569900 691100
rect 570100 690900 570110 691100
rect 570290 690900 570300 691100
rect 570500 690900 570510 691100
rect 570690 690900 570700 691100
rect 570900 690900 570910 691100
rect 571090 690900 571100 691100
rect 571300 690900 571310 691100
rect 571490 690900 571500 691100
rect 571700 690900 571710 691100
rect 546899 690842 547189 690892
rect 543879 690722 544029 690772
rect 543199 690532 543219 690612
rect 543299 690532 543389 690612
rect 543469 690532 543489 690612
rect 543579 690682 543659 690692
rect 543579 690592 543659 690602
rect 543729 690682 543809 690692
rect 543729 690592 543809 690602
rect 543879 690652 543889 690722
rect 544019 690652 544029 690722
rect 543199 690072 543489 690532
rect 543879 690182 544029 690652
rect 543199 689992 543219 690072
rect 543299 689992 543389 690072
rect 543469 689992 543489 690072
rect 543579 690142 543659 690152
rect 543579 690052 543659 690062
rect 543729 690142 543809 690152
rect 543729 690052 543809 690062
rect 543879 690112 543889 690182
rect 544019 690112 544029 690182
rect 543199 689532 543489 689992
rect 543879 689642 544029 690112
rect 544439 690312 544729 690772
rect 544439 690232 544459 690312
rect 544539 690232 544629 690312
rect 544709 690232 544729 690312
rect 544439 689922 544729 690232
rect 544439 689912 544619 689922
rect 544439 689842 544459 689912
rect 544549 689852 544619 689912
rect 544709 689852 544729 689922
rect 544549 689842 544729 689852
rect 544439 689782 544729 689842
rect 544439 689702 544459 689782
rect 544539 689702 544629 689782
rect 544709 689702 544729 689782
rect 544439 689682 544729 689702
rect 545119 690722 545269 690772
rect 545119 690652 545129 690722
rect 545259 690652 545269 690722
rect 545119 690182 545269 690652
rect 545119 690112 545129 690182
rect 545259 690112 545269 690182
rect 543199 689452 543219 689532
rect 543299 689452 543389 689532
rect 543469 689452 543489 689532
rect 543579 689602 543659 689612
rect 543579 689512 543659 689522
rect 543729 689602 543809 689612
rect 543729 689512 543809 689522
rect 543879 689572 543889 689642
rect 544019 689572 544029 689642
rect 543199 689422 543489 689452
rect 542649 689032 542659 689102
rect 542789 689032 542799 689102
rect 543879 689102 544029 689572
rect 545119 689642 545269 690112
rect 545119 689572 545129 689642
rect 545259 689572 545269 689642
rect 544459 689382 544539 689392
rect 544629 689382 544709 689392
rect 542379 689002 542459 689012
rect 542379 688912 542459 688922
rect 542489 689002 542569 689012
rect 542489 688912 542569 688922
rect 541959 688592 541979 688672
rect 542059 688592 542149 688672
rect 542229 688592 542249 688672
rect 541959 688222 542249 688592
rect 542649 688522 542799 689032
rect 542649 688452 542659 688522
rect 542789 688452 542799 688522
rect 542379 688392 542459 688402
rect 542379 688302 542459 688312
rect 542489 688392 542569 688402
rect 542489 688302 542569 688312
rect 541959 688142 541979 688222
rect 542069 688142 542139 688222
rect 542229 688142 542249 688222
rect 541959 688092 542249 688142
rect 541959 688012 541979 688092
rect 542059 688012 542149 688092
rect 542229 688012 542249 688092
rect 541959 687992 542249 688012
rect 541409 687872 541419 687942
rect 541549 687872 541559 687942
rect 542649 687942 542799 688452
rect 541409 687832 541559 687872
rect 47600 687260 47630 687330
rect 47700 687260 47730 687330
rect 47600 687170 47730 687260
rect 47600 687100 47630 687170
rect 47700 687100 47730 687170
rect 47600 687080 47730 687100
rect 538849 687652 539139 687732
rect 540759 687722 540889 687802
rect 542350 687830 542600 687880
rect 542350 687750 542380 687830
rect 542460 687750 542500 687830
rect 542580 687750 542600 687830
rect 542649 687872 542659 687942
rect 542789 687872 542799 687942
rect 542649 687792 542799 687872
rect 543181 688992 543513 689042
rect 543181 688912 543209 688992
rect 543289 688912 543379 688992
rect 543459 688912 543513 688992
rect 543181 688412 543513 688912
rect 543181 688332 543209 688412
rect 543289 688332 543379 688412
rect 543459 688332 543513 688412
rect 543181 687832 543513 688332
rect 543879 689032 543889 689102
rect 544019 689032 544029 689102
rect 543879 688522 544029 689032
rect 543879 688452 543899 688522
rect 543879 687942 544029 688452
rect 544439 689262 544729 689302
rect 544439 689182 544459 689262
rect 544539 689182 544629 689262
rect 544709 689182 544729 689262
rect 544439 688682 544729 689182
rect 545119 689102 545269 689572
rect 545689 690612 545979 690812
rect 546899 690762 546919 690842
rect 546999 690762 547089 690842
rect 547169 690762 547189 690842
rect 546359 690722 546509 690762
rect 545689 690532 545709 690612
rect 545789 690532 545879 690612
rect 545959 690532 545979 690612
rect 546059 690682 546139 690692
rect 546059 690592 546139 690602
rect 546209 690682 546289 690692
rect 546209 690592 546289 690602
rect 546359 690652 546369 690722
rect 546499 690652 546509 690722
rect 545689 690072 545979 690532
rect 546359 690432 546509 690652
rect 546349 690182 546509 690432
rect 545689 689992 545709 690072
rect 545789 689992 545879 690072
rect 545959 689992 545979 690072
rect 546059 690142 546139 690152
rect 546059 690052 546139 690062
rect 546209 690142 546289 690152
rect 546209 690052 546289 690062
rect 546349 690112 546369 690182
rect 546499 690112 546509 690182
rect 545689 689522 545979 689992
rect 546349 689642 546509 690112
rect 545689 689442 545709 689522
rect 545789 689442 545879 689522
rect 545959 689442 545979 689522
rect 546069 689602 546149 689612
rect 546069 689512 546149 689522
rect 546209 689602 546289 689612
rect 546209 689512 546289 689522
rect 546349 689572 546369 689642
rect 546499 689572 546509 689642
rect 546349 689532 546509 689572
rect 546899 690302 547189 690762
rect 546899 690222 546919 690302
rect 546999 690222 547089 690302
rect 547169 690222 547189 690302
rect 546899 689922 547189 690222
rect 546899 689852 546919 689922
rect 546999 689852 547089 689922
rect 547169 689852 547189 689922
rect 546899 689762 547189 689852
rect 546899 689682 546919 689762
rect 546999 689682 547089 689762
rect 547169 689682 547189 689762
rect 545689 689422 545979 689442
rect 545119 689032 545129 689102
rect 545259 689032 545269 689102
rect 546349 689102 546499 689532
rect 546899 689432 547189 689682
rect 547589 690722 547739 690752
rect 547589 690652 547599 690722
rect 547729 690652 547739 690722
rect 547589 690182 547739 690652
rect 547589 690112 547599 690182
rect 547729 690112 547739 690182
rect 547589 689642 547739 690112
rect 547589 689572 547599 689642
rect 547729 689572 547739 689642
rect 546919 689382 546999 689392
rect 547089 689382 547169 689392
rect 546349 689032 546359 689102
rect 546489 689032 546499 689102
rect 544789 689002 544869 689012
rect 544789 688912 544869 688922
rect 544899 689002 544979 689012
rect 544899 688912 544979 688922
rect 544439 688602 544459 688682
rect 544539 688602 544629 688682
rect 544709 688602 544729 688682
rect 544439 688212 544729 688602
rect 545119 688522 545269 689032
rect 545119 688452 545129 688522
rect 545259 688452 545269 688522
rect 544789 688412 544869 688422
rect 544789 688322 544869 688332
rect 544899 688412 544979 688422
rect 544899 688322 544979 688332
rect 544439 688142 544459 688212
rect 544539 688142 544629 688212
rect 544709 688142 544729 688212
rect 544439 688102 544729 688142
rect 544439 688022 544459 688102
rect 544539 688022 544629 688102
rect 544709 688022 544729 688102
rect 544439 688002 544729 688022
rect 543879 687872 543889 687942
rect 544019 687872 544029 687942
rect 543879 687842 544029 687872
rect 545119 687942 545269 688452
rect 545119 687872 545129 687942
rect 545259 687872 545269 687942
rect 545119 687842 545269 687872
rect 545679 688992 545969 689032
rect 545679 688912 545699 688992
rect 545779 688912 545869 688992
rect 545949 688912 545969 688992
rect 545679 688402 545969 688912
rect 545679 688322 545699 688402
rect 545779 688322 545869 688402
rect 545949 688322 545969 688402
rect 542350 687730 542600 687750
rect 543181 687752 543209 687832
rect 543289 687752 543379 687832
rect 543459 687752 543513 687832
rect 540679 687712 540759 687722
rect 540889 687712 540969 687722
rect 543181 687694 543513 687752
rect 544789 687832 544869 687842
rect 544789 687742 544869 687752
rect 544899 687832 544979 687842
rect 544899 687742 544979 687752
rect 545679 687832 545969 688322
rect 546349 688522 546499 689032
rect 546349 688452 546359 688522
rect 546489 688452 546499 688522
rect 546349 687942 546499 688452
rect 546899 689252 547189 689302
rect 546899 689172 546919 689252
rect 546999 689172 547089 689252
rect 547169 689172 547189 689252
rect 546899 688672 547189 689172
rect 547589 689102 547739 689572
rect 548139 690612 548429 690882
rect 548139 690532 548159 690612
rect 548239 690532 548329 690612
rect 548409 690532 548429 690612
rect 548139 690062 548429 690532
rect 566290 690500 566300 690700
rect 566500 690500 566510 690700
rect 566690 690500 566700 690700
rect 566900 690500 566910 690700
rect 567090 690500 567100 690700
rect 567300 690500 567310 690700
rect 567490 690500 567500 690700
rect 567700 690500 567710 690700
rect 567890 690500 567900 690700
rect 568100 690500 568110 690700
rect 568290 690500 568300 690700
rect 568500 690500 568510 690700
rect 568690 690500 568700 690700
rect 568900 690500 568910 690700
rect 569090 690500 569100 690700
rect 569300 690500 569310 690700
rect 569490 690500 569500 690700
rect 569700 690500 569710 690700
rect 569890 690500 569900 690700
rect 570100 690500 570110 690700
rect 570290 690500 570300 690700
rect 570500 690500 570510 690700
rect 570690 690500 570700 690700
rect 570900 690500 570910 690700
rect 571090 690500 571100 690700
rect 571300 690500 571310 690700
rect 571490 690500 571500 690700
rect 571700 690500 571710 690700
rect 566290 690100 566300 690300
rect 566500 690100 566510 690300
rect 566690 690100 566700 690300
rect 566900 690100 566910 690300
rect 567090 690100 567100 690300
rect 567300 690100 567310 690300
rect 567490 690100 567500 690300
rect 567700 690100 567710 690300
rect 567890 690100 567900 690300
rect 568100 690100 568110 690300
rect 568290 690100 568300 690300
rect 568500 690100 568510 690300
rect 568690 690100 568700 690300
rect 568900 690100 568910 690300
rect 569090 690100 569100 690300
rect 569300 690100 569310 690300
rect 569490 690100 569500 690300
rect 569700 690100 569710 690300
rect 569890 690100 569900 690300
rect 570100 690100 570110 690300
rect 570290 690100 570300 690300
rect 570500 690100 570510 690300
rect 570690 690100 570700 690300
rect 570900 690100 570910 690300
rect 571090 690100 571100 690300
rect 571300 690100 571310 690300
rect 571490 690100 571500 690300
rect 571700 690100 571710 690300
rect 548139 689982 548159 690062
rect 548239 689982 548329 690062
rect 548409 689982 548429 690062
rect 548139 689532 548429 689982
rect 566290 689700 566300 689900
rect 566500 689700 566510 689900
rect 566690 689700 566700 689900
rect 566900 689700 566910 689900
rect 567090 689700 567100 689900
rect 567300 689700 567310 689900
rect 567490 689700 567500 689900
rect 567700 689700 567710 689900
rect 567890 689700 567900 689900
rect 568100 689700 568110 689900
rect 568290 689700 568300 689900
rect 568500 689700 568510 689900
rect 568690 689700 568700 689900
rect 568900 689700 568910 689900
rect 569090 689700 569100 689900
rect 569300 689700 569310 689900
rect 569490 689700 569500 689900
rect 569700 689700 569710 689900
rect 569890 689700 569900 689900
rect 570100 689700 570110 689900
rect 570290 689700 570300 689900
rect 570500 689700 570510 689900
rect 570690 689700 570700 689900
rect 570900 689700 570910 689900
rect 571090 689700 571100 689900
rect 571300 689700 571310 689900
rect 571490 689700 571500 689900
rect 571700 689700 571710 689900
rect 548139 689452 548159 689532
rect 548239 689452 548329 689532
rect 548409 689452 548429 689532
rect 548139 689442 548429 689452
rect 566290 689300 566300 689500
rect 566500 689300 566510 689500
rect 566690 689300 566700 689500
rect 566900 689300 566910 689500
rect 567090 689300 567100 689500
rect 567300 689300 567310 689500
rect 567490 689300 567500 689500
rect 567700 689300 567710 689500
rect 567890 689300 567900 689500
rect 568100 689300 568110 689500
rect 568290 689300 568300 689500
rect 568500 689300 568510 689500
rect 568690 689300 568700 689500
rect 568900 689300 568910 689500
rect 569090 689300 569100 689500
rect 569300 689300 569310 689500
rect 569490 689300 569500 689500
rect 569700 689300 569710 689500
rect 569890 689300 569900 689500
rect 570100 689300 570110 689500
rect 570290 689300 570300 689500
rect 570500 689300 570510 689500
rect 570690 689300 570700 689500
rect 570900 689300 570910 689500
rect 571090 689300 571100 689500
rect 571300 689300 571310 689500
rect 571490 689300 571500 689500
rect 571700 689300 571710 689500
rect 547589 689032 547599 689102
rect 547729 689032 547739 689102
rect 547249 688992 547329 689002
rect 547249 688902 547329 688912
rect 547359 688992 547439 689002
rect 547359 688902 547439 688912
rect 546899 688592 546919 688672
rect 546999 688592 547089 688672
rect 547169 688592 547189 688672
rect 546899 688212 547189 688592
rect 547589 688522 547739 689032
rect 547589 688452 547599 688522
rect 547729 688452 547739 688522
rect 547249 688412 547329 688422
rect 547249 688322 547329 688332
rect 547359 688412 547439 688422
rect 547359 688322 547439 688332
rect 546899 688142 546919 688212
rect 546999 688142 547089 688212
rect 547169 688142 547189 688212
rect 546899 688092 547189 688142
rect 546899 688012 546919 688092
rect 546999 688012 547089 688092
rect 547169 688012 547189 688092
rect 546899 688002 547189 688012
rect 546349 687872 546359 687942
rect 546489 687872 546499 687942
rect 546349 687832 546499 687872
rect 547589 687942 547739 688452
rect 547589 687872 547599 687942
rect 547729 687872 547739 687942
rect 547589 687842 547739 687872
rect 548169 688992 548459 689082
rect 548169 688912 548189 688992
rect 548269 688912 548359 688992
rect 548439 688912 548459 688992
rect 548169 688412 548459 688912
rect 548169 688332 548189 688412
rect 548269 688332 548359 688412
rect 548439 688332 548459 688412
rect 547249 687832 547329 687842
rect 545679 687752 545699 687832
rect 545779 687752 545869 687832
rect 545949 687752 545969 687832
rect 545679 687732 545969 687752
rect 547249 687742 547329 687752
rect 547359 687832 547439 687842
rect 547359 687742 547439 687752
rect 548169 687832 548459 688332
rect 554129 688302 554259 688312
rect 554129 688152 554259 688162
rect 554389 688302 554519 688312
rect 554389 688152 554519 688162
rect 548169 687752 548189 687832
rect 548269 687752 548359 687832
rect 548439 687752 548459 687832
rect 548169 687732 548459 687752
rect 538849 687542 538869 687652
rect 538959 687542 539029 687652
rect 539119 687542 539139 687652
rect 548779 687602 549069 687642
rect 538849 687282 539139 687542
rect 540099 687562 540409 687582
rect 540179 687482 540329 687562
rect 538929 687202 539059 687282
rect 46640 686270 46660 686380
rect 46770 686270 46910 686380
rect 47020 686270 47040 686380
rect 46640 685970 47040 686270
rect 46640 685860 46660 685970
rect 46770 685860 46910 685970
rect 47020 685860 47040 685970
rect 43070 685150 43140 685160
rect 43070 685070 43140 685080
rect 43580 685150 43650 685160
rect 43580 685070 43650 685080
rect 44100 685150 44170 685160
rect 44100 685070 44170 685080
rect 44620 685150 44690 685160
rect 44620 685070 44690 685080
rect 45130 685150 45200 685160
rect 45130 685070 45200 685080
rect 45650 685150 45720 685160
rect 45650 685070 45720 685080
rect 46160 685150 46230 685160
rect 46160 685070 46230 685080
rect 43070 684970 43140 684980
rect 43070 684890 43140 684900
rect 43580 684970 43650 684980
rect 43580 684890 43650 684900
rect 44100 684970 44170 684980
rect 44100 684890 44170 684900
rect 44620 684970 44690 684980
rect 44620 684890 44690 684900
rect 45130 684970 45200 684980
rect 45130 684890 45200 684900
rect 45650 684970 45720 684980
rect 45650 684890 45720 684900
rect 46160 684970 46230 684980
rect 46160 684890 46230 684900
rect 42240 684750 42260 684860
rect 42370 684750 42510 684860
rect 42620 684750 42640 684860
rect 42240 683120 42640 684750
rect 46640 684860 47040 685860
rect 538849 686742 539139 687202
rect 538929 686662 539059 686742
rect 538849 686202 539139 686662
rect 538929 686122 539059 686202
rect 538849 685662 539139 686122
rect 539569 687402 539719 687432
rect 539569 687332 539579 687402
rect 539709 687332 539719 687402
rect 539569 686872 539719 687332
rect 539569 686802 539579 686872
rect 539709 686802 539719 686872
rect 539569 686322 539719 686802
rect 539569 686252 539579 686322
rect 539709 686252 539719 686322
rect 539569 685782 539719 686252
rect 540099 687142 540409 687482
rect 542629 687552 542919 687582
rect 542629 687472 542649 687552
rect 542729 687472 542819 687552
rect 542899 687472 542919 687552
rect 540099 687062 540119 687142
rect 540209 687062 540299 687142
rect 540389 687062 540409 687142
rect 540099 687022 540409 687062
rect 540179 686942 540329 687022
rect 540099 686482 540409 686942
rect 540179 686402 540329 686482
rect 540099 686072 540409 686402
rect 540099 686062 540299 686072
rect 540099 685982 540119 686062
rect 540209 685992 540299 686062
rect 540389 685992 540409 686072
rect 540209 685982 540409 685992
rect 540099 685932 540409 685982
rect 540179 685852 540329 685932
rect 540099 685842 540409 685852
rect 540809 687402 540959 687442
rect 540809 687332 540819 687402
rect 540949 687332 540959 687402
rect 540809 686862 540959 687332
rect 542039 687402 542189 687432
rect 542039 687332 542049 687402
rect 542179 687332 542189 687402
rect 540809 686792 540819 686862
rect 540949 686792 540959 686862
rect 540809 686322 540959 686792
rect 540809 686252 540819 686322
rect 540949 686252 540959 686322
rect 539569 685712 539579 685782
rect 539709 685712 539719 685782
rect 539569 685672 539719 685712
rect 540809 685782 540959 686252
rect 540809 685712 540819 685782
rect 540949 685712 540959 685782
rect 538929 685582 539059 685662
rect 538849 685572 539139 685582
rect 535759 685252 535849 685262
rect 535759 685112 535849 685122
rect 535969 685252 536059 685262
rect 535969 685112 536059 685122
rect 540809 685132 540959 685712
rect 541319 687282 541639 687312
rect 541319 687202 541329 687282
rect 541409 687202 541549 687282
rect 541629 687202 541639 687282
rect 541319 686742 541639 687202
rect 541319 686662 541329 686742
rect 541409 686662 541549 686742
rect 541629 686662 541639 686742
rect 541319 686202 541639 686662
rect 541399 686122 541559 686202
rect 541319 685732 541639 686122
rect 542039 686862 542189 687332
rect 542039 686792 542049 686862
rect 542179 686792 542189 686862
rect 542039 686322 542189 686792
rect 542039 686252 542049 686322
rect 542179 686252 542189 686322
rect 542039 685782 542189 686252
rect 542629 687142 542919 687472
rect 545099 687552 545389 687592
rect 545099 687472 545109 687552
rect 545189 687472 545299 687552
rect 545379 687472 545389 687552
rect 542629 687062 542649 687142
rect 542739 687062 542809 687142
rect 542899 687062 542919 687142
rect 542629 687022 542919 687062
rect 542629 687012 542819 687022
rect 542629 686932 542649 687012
rect 542729 686942 542819 687012
rect 542899 686942 542919 687022
rect 542729 686932 542919 686942
rect 542629 686472 542919 686932
rect 542629 686392 542639 686472
rect 542719 686392 542809 686472
rect 542889 686392 542919 686472
rect 542629 686062 542919 686392
rect 542629 685982 542649 686062
rect 542739 685982 542809 686062
rect 542899 685982 542919 686062
rect 542629 685942 542919 685982
rect 542709 685862 542819 685942
rect 542899 685862 542919 685942
rect 542629 685832 542919 685862
rect 543279 687402 543429 687432
rect 543279 687332 543289 687402
rect 543419 687332 543429 687402
rect 544519 687402 544669 687422
rect 543279 686862 543429 687332
rect 543279 686792 543289 686862
rect 543419 686792 543429 686862
rect 543279 686322 543429 686792
rect 543279 686252 543289 686322
rect 543419 686252 543429 686322
rect 541319 685652 541729 685732
rect 541399 685572 541559 685652
rect 541639 685572 541729 685652
rect 541319 685472 541729 685572
rect 540809 685062 540819 685132
rect 540949 685062 540959 685132
rect 540809 685052 540959 685062
rect 46640 684750 46660 684860
rect 46770 684750 46910 684860
rect 47020 684750 47040 684860
rect 44530 684720 44780 684730
rect 44530 684460 44780 684470
rect 43840 683600 43920 683610
rect 43840 683510 43920 683520
rect 44350 683600 44430 683610
rect 44350 683510 44430 683520
rect 44870 683600 44950 683610
rect 44870 683510 44950 683520
rect 45390 683600 45470 683610
rect 45390 683510 45470 683520
rect 42240 683040 42260 683120
rect 42340 683040 42400 683120
rect 42480 683040 42540 683120
rect 42620 683040 42640 683120
rect 42240 683020 42640 683040
rect 44080 683120 44180 683130
rect 44080 683040 44090 683120
rect 44170 683040 44180 683120
rect 43900 682770 44010 682780
rect 43900 682700 43920 682770
rect 43990 682700 44010 682770
rect 43900 682440 44010 682700
rect 43900 682370 43920 682440
rect 43990 682370 44010 682440
rect 43900 682360 44010 682370
rect 43840 682140 43920 682150
rect 43840 682050 43920 682060
rect 43630 681920 43710 681930
rect 43630 681830 43710 681840
rect 43630 681780 43710 681790
rect 43630 681690 43710 681700
rect 43790 681270 43930 681280
rect 43790 681170 43810 681270
rect 43910 681170 43930 681270
rect 43790 678690 43930 681170
rect 44080 679830 44180 683040
rect 44610 683120 44690 683130
rect 44610 683030 44690 683040
rect 45120 683120 45220 683130
rect 45120 683040 45130 683120
rect 45210 683040 45220 683120
rect 44600 682770 44710 682780
rect 44600 682700 44620 682770
rect 44690 682700 44710 682770
rect 44600 682440 44710 682700
rect 44600 682370 44620 682440
rect 44690 682370 44710 682440
rect 44600 682360 44710 682370
rect 44350 682140 44430 682150
rect 44350 682050 44430 682060
rect 44870 682140 44950 682150
rect 44870 682050 44950 682060
rect 44590 681270 44680 681280
rect 44590 681200 44600 681270
rect 44670 681200 44680 681270
rect 44590 680830 44680 681200
rect 44590 680760 44600 680830
rect 44670 680760 44680 680830
rect 44590 680750 44680 680760
rect 44890 680530 45010 680540
rect 44270 680520 44390 680530
rect 44890 680400 45010 680410
rect 44270 680390 44390 680400
rect 44080 679750 44090 679830
rect 44170 679750 44180 679830
rect 44590 680360 44680 680370
rect 44590 680290 44600 680360
rect 44670 680290 44680 680360
rect 44590 679830 44680 680290
rect 44590 679790 44600 679830
rect 44670 679790 44680 679830
rect 45120 679830 45220 683040
rect 46640 683120 47040 684750
rect 46640 683040 46660 683120
rect 46740 683040 46800 683120
rect 46880 683040 46940 683120
rect 47020 683040 47040 683120
rect 46640 683020 47040 683040
rect 540759 684862 540849 684872
rect 540899 684862 540989 684872
rect 540849 684782 540899 684852
rect 540759 684632 540989 684782
rect 540849 684552 540899 684632
rect 45290 682770 45400 682780
rect 45290 682700 45310 682770
rect 45380 682700 45400 682770
rect 45290 682440 45400 682700
rect 45290 682370 45310 682440
rect 45380 682370 45400 682440
rect 45290 682360 45400 682370
rect 540759 682582 540989 684552
rect 541069 684372 541339 684382
rect 541069 684292 541089 684372
rect 541169 684292 541239 684372
rect 541319 684292 541339 684372
rect 541089 684282 541169 684292
rect 541239 684282 541319 684292
rect 541539 684172 541729 685472
rect 542039 685712 542049 685782
rect 542179 685712 542189 685782
rect 542039 685122 542189 685712
rect 543279 685782 543429 686252
rect 543279 685712 543289 685782
rect 543419 685712 543429 685782
rect 542039 685052 542049 685122
rect 542179 685052 542189 685122
rect 542039 685002 542189 685052
rect 542379 685132 542459 685142
rect 542379 685042 542459 685052
rect 542489 685132 542569 685142
rect 542489 685042 542569 685052
rect 543279 685122 543429 685712
rect 543279 685052 543289 685122
rect 543419 685052 543429 685122
rect 543279 684962 543429 685052
rect 543849 687282 544139 687372
rect 543849 687202 543859 687282
rect 543939 687202 544039 687282
rect 544119 687202 544139 687282
rect 543849 686742 544139 687202
rect 543849 686662 543859 686742
rect 543939 686662 544049 686742
rect 544129 686662 544139 686742
rect 543849 686202 544139 686662
rect 543849 686122 543859 686202
rect 543939 686122 544039 686202
rect 544119 686122 544139 686202
rect 543849 685662 544139 686122
rect 543849 685582 543859 685662
rect 543939 685582 544049 685662
rect 544129 685582 544139 685662
rect 542279 684772 542389 684782
rect 542279 684652 542389 684662
rect 543139 684772 543249 684782
rect 543139 684652 543249 684662
rect 543579 684392 543659 684402
rect 543579 684302 543659 684312
rect 543729 684392 543809 684402
rect 543729 684302 543809 684312
rect 541449 684142 541759 684172
rect 541449 684062 541539 684142
rect 541619 684062 541649 684142
rect 541729 684062 541759 684142
rect 543849 684112 544139 685582
rect 544519 687332 544529 687402
rect 544659 687332 544669 687402
rect 544519 686862 544669 687332
rect 544519 686792 544529 686862
rect 544659 686792 544669 686862
rect 544519 686322 544669 686792
rect 544519 686252 544529 686322
rect 544659 686252 544669 686322
rect 544519 685782 544669 686252
rect 545099 687142 545389 687472
rect 547549 687552 547839 687582
rect 547549 687472 547559 687552
rect 547639 687472 547749 687552
rect 547829 687472 547839 687552
rect 545099 687062 545119 687142
rect 545209 687062 545279 687142
rect 545369 687062 545389 687142
rect 545099 687022 545389 687062
rect 545099 686942 545109 687022
rect 545189 686942 545299 687022
rect 545379 686942 545389 687022
rect 545099 686472 545389 686942
rect 545099 686392 545109 686472
rect 545189 686392 545289 686472
rect 545369 686392 545389 686472
rect 545099 686062 545389 686392
rect 545099 685982 545119 686062
rect 545209 685982 545279 686062
rect 545369 685982 545389 686062
rect 545099 685932 545389 685982
rect 545099 685852 545109 685932
rect 545189 685852 545299 685932
rect 545379 685852 545389 685932
rect 545099 685842 545389 685852
rect 545749 687402 545899 687432
rect 545749 687332 545759 687402
rect 545889 687332 545899 687402
rect 546989 687402 547139 687452
rect 545749 686862 545899 687332
rect 545749 686792 545759 686862
rect 545889 686792 545899 686862
rect 545749 686322 545899 686792
rect 545749 686252 545759 686322
rect 545889 686252 545899 686322
rect 544519 685712 544529 685782
rect 544659 685712 544669 685782
rect 544519 685122 544669 685712
rect 545749 685782 545899 686252
rect 545749 685712 545759 685782
rect 545889 685712 545899 685782
rect 544519 685052 544529 685122
rect 544659 685052 544669 685122
rect 544519 684982 544669 685052
rect 544789 685132 544869 685142
rect 544789 685042 544869 685052
rect 544899 685132 544979 685142
rect 544899 685042 544979 685052
rect 545749 685122 545899 685712
rect 546309 687272 546599 687372
rect 546309 687192 546319 687272
rect 546399 687192 546499 687272
rect 546579 687192 546599 687272
rect 546309 686732 546599 687192
rect 546309 686652 546319 686732
rect 546399 686652 546499 686732
rect 546579 686652 546599 686732
rect 546309 686192 546599 686652
rect 546309 686112 546329 686192
rect 546409 686112 546499 686192
rect 546579 686112 546599 686192
rect 546309 685752 546599 686112
rect 546989 687332 546999 687402
rect 547129 687332 547139 687402
rect 546989 686862 547139 687332
rect 546989 686792 546999 686862
rect 547129 686792 547139 686862
rect 546989 686322 547139 686792
rect 546989 686252 546999 686322
rect 547129 686252 547139 686322
rect 546989 685782 547139 686252
rect 546309 685652 546609 685752
rect 546309 685572 546319 685652
rect 546399 685572 546509 685652
rect 546589 685572 546609 685652
rect 546309 685552 546609 685572
rect 545749 685052 545759 685122
rect 545889 685052 545899 685122
rect 545749 685042 545899 685052
rect 545769 684882 545859 684892
rect 545909 684882 545999 684892
rect 545859 684802 545909 684882
rect 544349 684772 544459 684782
rect 544349 684652 544459 684662
rect 545199 684772 545309 684782
rect 545199 684652 545309 684662
rect 543849 684062 543949 684112
rect 541449 684042 541759 684062
rect 544029 684062 544139 684112
rect 545769 684622 545999 684802
rect 545859 684542 545909 684622
rect 542719 683962 542799 683992
rect 541459 683782 541539 683812
rect 541459 683692 541539 683702
rect 541459 683652 541719 683692
rect 541459 683562 541569 683652
rect 541679 683562 541719 683652
rect 541459 683522 541719 683562
rect 541459 683162 541539 683522
rect 541459 683072 541539 683082
rect 542109 683342 542319 683362
rect 542199 683262 542229 683342
rect 540849 682502 540899 682582
rect 45390 682140 45470 682150
rect 45390 682050 45470 682060
rect 540759 681962 540989 682502
rect 542109 682742 542319 683262
rect 542719 683342 542799 683882
rect 543949 683492 544029 684032
rect 543949 683402 544029 683412
rect 545129 683962 545209 683992
rect 542719 683252 542799 683262
rect 544559 683342 544769 683362
rect 544649 683262 544679 683342
rect 542199 682662 542229 682742
rect 541509 682452 541629 682462
rect 541509 682342 541629 682352
rect 542109 682142 542319 682662
rect 543339 682912 543429 682942
rect 542729 682452 542849 682462
rect 542729 682342 542849 682352
rect 543339 682312 543429 682832
rect 544559 682742 544769 683262
rect 545129 683342 545209 683882
rect 545129 683252 545209 683262
rect 544649 682662 544679 682742
rect 543939 682452 544059 682462
rect 543939 682342 544059 682352
rect 543339 682222 543429 682232
rect 544559 682196 544769 682662
rect 545769 682582 545999 684542
rect 546059 684392 546139 684402
rect 546059 684302 546139 684312
rect 546199 684392 546279 684402
rect 546199 684302 546279 684312
rect 546389 684132 546609 685552
rect 546989 685712 546999 685782
rect 547129 685712 547139 685782
rect 546989 685142 547139 685712
rect 547549 687142 547839 687472
rect 548779 687522 548799 687602
rect 548879 687522 548969 687602
rect 549049 687522 549069 687602
rect 547549 687062 547569 687142
rect 547659 687062 547729 687142
rect 547819 687062 547839 687142
rect 547549 687012 547839 687062
rect 547549 686932 547559 687012
rect 547639 686932 547749 687012
rect 547829 686932 547839 687012
rect 547549 686472 547839 686932
rect 547549 686392 547559 686472
rect 547639 686392 547749 686472
rect 547829 686392 547839 686472
rect 547549 686062 547839 686392
rect 547549 685982 547569 686062
rect 547659 685982 547729 686062
rect 547819 685982 547839 686062
rect 547549 685932 547839 685982
rect 547549 685852 547559 685932
rect 547639 685852 547749 685932
rect 547829 685852 547839 685932
rect 547549 685602 547839 685852
rect 548219 687402 548369 687442
rect 548219 687332 548229 687402
rect 548359 687332 548369 687402
rect 548219 686862 548369 687332
rect 548219 686792 548229 686862
rect 548359 686792 548369 686862
rect 548219 686322 548369 686792
rect 548219 686252 548229 686322
rect 548359 686252 548369 686322
rect 548219 685782 548369 686252
rect 548219 685712 548229 685782
rect 548359 685712 548369 685782
rect 546989 685072 546999 685142
rect 547129 685072 547139 685142
rect 546989 685012 547139 685072
rect 547249 685142 547329 685152
rect 547249 685052 547329 685062
rect 547359 685142 547439 685152
rect 547359 685052 547439 685062
rect 548219 685122 548369 685712
rect 548779 687272 549069 687522
rect 550049 687552 550339 687572
rect 550049 687472 550069 687552
rect 550149 687472 550239 687552
rect 550319 687472 550339 687552
rect 548779 687192 548799 687272
rect 548879 687192 548969 687272
rect 549049 687192 549069 687272
rect 548779 686732 549069 687192
rect 548779 686652 548799 686732
rect 548879 686652 548969 686732
rect 549049 686652 549069 686732
rect 548779 686192 549069 686652
rect 548779 686112 548799 686192
rect 548879 686112 548969 686192
rect 549049 686112 549069 686192
rect 548779 685642 549069 686112
rect 549459 687402 549609 687442
rect 549459 687332 549469 687402
rect 549599 687332 549609 687402
rect 549459 686862 549609 687332
rect 549459 686792 549469 686862
rect 549599 686792 549609 686862
rect 549459 686322 549609 686792
rect 549459 686252 549469 686322
rect 549599 686252 549609 686322
rect 549459 685782 549609 686252
rect 550049 687142 550339 687472
rect 550049 687062 550069 687142
rect 550159 687062 550229 687142
rect 550319 687062 550339 687142
rect 550049 687012 550339 687062
rect 550049 686932 550069 687012
rect 550149 686932 550239 687012
rect 550319 686932 550339 687012
rect 550049 686472 550339 686932
rect 550049 686392 550069 686472
rect 550149 686392 550239 686472
rect 550319 686392 550339 686472
rect 550049 686062 550339 686392
rect 550049 685982 550069 686062
rect 550159 685982 550229 686062
rect 550319 685982 550339 686062
rect 550049 685922 550339 685982
rect 550049 685842 550069 685922
rect 550149 685842 550239 685922
rect 550319 685842 550339 685922
rect 550049 685822 550339 685842
rect 549459 685712 549469 685782
rect 549599 685712 549609 685782
rect 549459 685682 549609 685712
rect 548779 685562 548799 685642
rect 548879 685562 548969 685642
rect 549049 685562 549069 685642
rect 548779 685552 549069 685562
rect 553069 685242 553139 685252
rect 553069 685142 553139 685152
rect 553229 685242 553299 685252
rect 553229 685142 553299 685152
rect 548219 685052 548229 685122
rect 548359 685052 548369 685122
rect 548219 685012 548369 685052
rect 546769 684772 546879 684782
rect 546769 684652 546879 684662
rect 547649 684772 547759 684782
rect 547649 684652 547759 684662
rect 546389 684052 546399 684132
rect 546479 684052 546519 684132
rect 546599 684052 546609 684132
rect 547549 684122 547839 684132
rect 547549 684082 547599 684122
rect 546389 684042 546609 684052
rect 547679 684082 547839 684122
rect 546349 683782 546429 683812
rect 546349 683692 546429 683702
rect 546349 683652 546619 683692
rect 546349 683562 546479 683652
rect 546589 683562 546619 683652
rect 546349 683522 546619 683562
rect 546349 683162 546429 683522
rect 547599 683502 547679 684042
rect 547599 683412 547679 683422
rect 546349 683072 546429 683082
rect 546989 683342 547199 683362
rect 547079 683262 547109 683342
rect 545859 682502 545909 682582
rect 545159 682452 545279 682462
rect 545159 682342 545279 682352
rect 542199 682062 542229 682142
rect 542109 682052 542319 682062
rect 544390 682146 544790 682196
rect 544390 682056 544420 682146
rect 544508 682142 544790 682146
rect 544508 682062 544559 682142
rect 544649 682062 544679 682142
rect 544769 682062 544790 682142
rect 544508 682056 544790 682062
rect 45590 681920 45670 681930
rect 540849 681882 540899 681962
rect 540759 681872 540989 681882
rect 45590 681830 45670 681840
rect 45590 681780 45670 681790
rect 45590 681690 45670 681700
rect 541384 681478 541544 681488
rect 541384 681308 541544 681318
rect 542444 681478 542604 681488
rect 542444 681308 542604 681318
rect 543904 681478 544064 681488
rect 543904 681308 544064 681318
rect 44600 679750 44670 679760
rect 45120 679750 45130 679830
rect 45210 679750 45220 679830
rect 44080 679740 44180 679750
rect 45120 679740 45220 679750
rect 45340 681270 45480 681280
rect 45340 681170 45360 681270
rect 45460 681170 45480 681270
rect 44070 679630 44160 679640
rect 44070 679530 44160 679540
rect 44590 679630 44680 679640
rect 44590 679530 44680 679540
rect 45100 679630 45190 679640
rect 45100 679530 45190 679540
rect 44210 679420 44290 679430
rect 44210 679360 44220 679420
rect 44280 679360 44290 679420
rect 44210 679060 44290 679360
rect 44980 679420 45060 679430
rect 44980 679360 44990 679420
rect 45050 679360 45060 679420
rect 44580 679250 44670 679260
rect 44580 679150 44670 679160
rect 44210 679000 44220 679060
rect 44280 679000 44290 679060
rect 44210 678990 44290 679000
rect 44980 679060 45060 679360
rect 44980 679000 44990 679060
rect 45050 679000 45060 679060
rect 44980 678990 45060 679000
rect 44830 678720 44960 678730
rect 43790 678630 43830 678690
rect 43890 678630 43930 678690
rect 43790 678620 43930 678630
rect 44350 678690 44410 678700
rect 44350 678620 44410 678630
rect 45340 678690 45480 681170
rect 542864 681088 542884 681158
rect 542954 681088 543104 681158
rect 543174 681088 543194 681158
rect 541384 680898 541544 680908
rect 541384 680728 541544 680738
rect 542444 680898 542604 680908
rect 542444 680728 542604 680738
rect 542864 680568 543194 681088
rect 543904 680898 544064 680908
rect 543904 680728 544064 680738
rect 542864 680498 542884 680568
rect 542954 680498 543104 680568
rect 543174 680498 543194 680568
rect 542864 679308 543194 680498
rect 544024 680408 544244 680418
rect 544024 680338 544044 680408
rect 544114 680338 544154 680408
rect 544224 680338 544244 680408
rect 544024 679838 544244 680338
rect 544390 679926 544790 682056
rect 545769 681982 545999 682502
rect 546989 682742 547199 683262
rect 547079 682662 547109 682742
rect 546389 682442 546509 682452
rect 546389 682332 546509 682342
rect 546989 682142 547199 682662
rect 548219 682932 548309 682962
rect 547599 682452 547719 682462
rect 547599 682342 547719 682352
rect 548219 682332 548309 682852
rect 548219 682242 548309 682252
rect 547079 682062 547109 682142
rect 546989 682052 547199 682062
rect 561700 682200 561900 682210
rect 561700 681990 561900 682000
rect 562100 682200 562300 682210
rect 562100 681990 562300 682000
rect 562500 682200 562700 682210
rect 562500 681990 562700 682000
rect 562900 682200 563100 682210
rect 562900 681990 563100 682000
rect 563300 682200 563500 682210
rect 563300 681990 563500 682000
rect 545859 681902 545909 681982
rect 545769 681892 545999 681902
rect 561700 681800 561900 681810
rect 561700 681590 561900 681600
rect 562100 681800 562300 681810
rect 562100 681590 562300 681600
rect 562500 681800 562700 681810
rect 562500 681590 562700 681600
rect 562900 681800 563100 681810
rect 562900 681590 563100 681600
rect 563300 681800 563500 681810
rect 563300 681590 563500 681600
rect 545124 681478 545284 681488
rect 545124 681308 545284 681318
rect 546604 681478 546764 681488
rect 546604 681308 546764 681318
rect 547604 681478 547764 681488
rect 547604 681308 547764 681318
rect 561700 681400 561900 681410
rect 561700 681190 561900 681200
rect 562100 681400 562300 681410
rect 562100 681190 562300 681200
rect 562500 681400 562700 681410
rect 562500 681190 562700 681200
rect 562900 681400 563100 681410
rect 562900 681190 563100 681200
rect 563300 681400 563500 681410
rect 563300 681190 563500 681200
rect 546044 681158 546394 681168
rect 546044 681088 546064 681158
rect 546134 681088 546304 681158
rect 546374 681088 546394 681158
rect 545124 680898 545284 680908
rect 545124 680728 545284 680738
rect 546044 680568 546394 681088
rect 561700 681000 561900 681010
rect 546604 680898 546764 680908
rect 546604 680728 546764 680738
rect 547604 680898 547764 680908
rect 561700 680790 561900 680800
rect 562100 681000 562300 681010
rect 562100 680790 562300 680800
rect 562500 681000 562700 681010
rect 562500 680790 562700 680800
rect 562900 681000 563100 681010
rect 562900 680790 563100 680800
rect 563300 681000 563500 681010
rect 563300 680790 563500 680800
rect 547604 680728 547764 680738
rect 546044 680498 546064 680568
rect 546134 680498 546304 680568
rect 546374 680498 546394 680568
rect 544390 679866 544410 679926
rect 544470 679866 544510 679926
rect 544570 679866 544610 679926
rect 544670 679866 544710 679926
rect 544770 679866 544790 679926
rect 544390 679846 544790 679866
rect 544964 680408 545184 680428
rect 544964 680338 544984 680408
rect 545054 680338 545094 680408
rect 545164 680338 545184 680408
rect 544964 679848 545184 680338
rect 544024 679768 544044 679838
rect 544114 679768 544154 679838
rect 544224 679768 544244 679838
rect 543764 679518 543984 679528
rect 543764 679358 543984 679368
rect 542864 679238 542884 679308
rect 542954 679238 543094 679308
rect 543164 679238 543194 679308
rect 542864 679218 543194 679238
rect 542864 679148 542884 679218
rect 542954 679148 543094 679218
rect 543164 679148 543194 679218
rect 541404 678958 541584 678968
rect 541404 678818 541584 678828
rect 542544 678958 542724 678968
rect 542544 678818 542724 678828
rect 542864 678788 543194 679148
rect 544024 679088 544244 679768
rect 544964 679778 544984 679848
rect 545054 679778 545094 679848
rect 545164 679778 545184 679848
rect 544284 679518 544504 679528
rect 544284 679358 544504 679368
rect 544704 679518 544924 679528
rect 544704 679358 544924 679368
rect 544024 679018 544044 679088
rect 544114 679018 544154 679088
rect 544224 679018 544244 679088
rect 543524 678968 543704 678978
rect 543524 678828 543704 678838
rect 542864 678718 542884 678788
rect 542954 678718 543104 678788
rect 543174 678718 543194 678788
rect 542864 678708 543194 678718
rect 45340 678630 45380 678690
rect 45440 678630 45480 678690
rect 45340 678620 45480 678630
rect 544024 678638 544244 679018
rect 544964 679088 545184 679778
rect 545254 679518 545474 679528
rect 545254 679358 545474 679368
rect 544964 679018 544984 679088
rect 545054 679018 545094 679088
rect 545164 679018 545184 679088
rect 544294 678968 544474 678978
rect 544294 678828 544474 678838
rect 544734 678968 544914 678978
rect 544734 678828 544914 678838
rect 44830 678600 44960 678610
rect 544024 678568 544044 678638
rect 544114 678568 544154 678638
rect 544224 678568 544244 678638
rect 544024 678498 544244 678568
rect 544964 678638 545184 679018
rect 546044 679328 546394 680498
rect 561700 680600 561900 680610
rect 561700 680390 561900 680400
rect 562100 680600 562300 680610
rect 562100 680390 562300 680400
rect 562500 680600 562700 680610
rect 562500 680390 562700 680400
rect 562900 680600 563100 680610
rect 562900 680390 563100 680400
rect 563300 680600 563500 680610
rect 563300 680390 563500 680400
rect 561700 680200 561900 680210
rect 561700 679990 561900 680000
rect 562100 680200 562300 680210
rect 562100 679990 562300 680000
rect 562500 680200 562700 680210
rect 562500 679990 562700 680000
rect 562900 680200 563100 680210
rect 562900 679990 563100 680000
rect 563300 680200 563500 680210
rect 563300 679990 563500 680000
rect 561700 679800 561900 679810
rect 561700 679590 561900 679600
rect 562100 679800 562300 679810
rect 562100 679590 562300 679600
rect 562500 679800 562700 679810
rect 562500 679590 562700 679600
rect 562900 679800 563100 679810
rect 562900 679590 563100 679600
rect 563300 679800 563500 679810
rect 563300 679590 563500 679600
rect 546044 679258 546064 679328
rect 546134 679258 546304 679328
rect 546374 679258 546394 679328
rect 546044 679238 546394 679258
rect 546044 679168 546064 679238
rect 546134 679168 546304 679238
rect 546374 679168 546394 679238
rect 561700 679400 561900 679410
rect 561700 679190 561900 679200
rect 562100 679400 562300 679410
rect 562100 679190 562300 679200
rect 562500 679400 562700 679410
rect 562500 679190 562700 679200
rect 562900 679400 563100 679410
rect 562900 679190 563100 679200
rect 563300 679400 563500 679410
rect 563300 679190 563500 679200
rect 545454 678958 545634 678968
rect 545454 678818 545634 678828
rect 546044 678788 546394 679168
rect 561700 679000 561900 679010
rect 546524 678968 546704 678978
rect 546524 678828 546704 678838
rect 547524 678968 547704 678978
rect 547524 678828 547704 678838
rect 561700 678790 561900 678800
rect 562100 679000 562300 679010
rect 562100 678790 562300 678800
rect 562500 679000 562700 679010
rect 562500 678790 562700 678800
rect 562900 679000 563100 679010
rect 562900 678790 563100 678800
rect 563300 679000 563500 679010
rect 563300 678790 563500 678800
rect 546044 678718 546064 678788
rect 546134 678718 546304 678788
rect 546374 678718 546394 678788
rect 546044 678688 546394 678718
rect 544964 678568 544984 678638
rect 545054 678568 545094 678638
rect 545164 678568 545184 678638
rect 544964 678508 545184 678568
rect 561700 678600 561900 678610
rect 561700 678390 561900 678400
rect 562100 678600 562300 678610
rect 562100 678390 562300 678400
rect 562500 678600 562700 678610
rect 562500 678390 562700 678400
rect 562900 678600 563100 678610
rect 562900 678390 563100 678400
rect 563300 678600 563500 678610
rect 563300 678390 563500 678400
rect 44070 678280 44170 678290
rect 44070 678220 44090 678280
rect 44150 678220 44170 678280
rect 44070 677530 44170 678220
rect 44610 678280 44670 678290
rect 44610 678210 44670 678220
rect 45100 678280 45200 678290
rect 45100 678220 45120 678280
rect 45180 678220 45200 678280
rect 44580 677810 44670 677820
rect 44580 677710 44670 677720
rect 44070 677470 44090 677530
rect 44150 677470 44170 677530
rect 44070 677360 44170 677470
rect 44070 677300 44090 677360
rect 44150 677300 44170 677360
rect 44070 677190 44170 677300
rect 44070 677130 44090 677190
rect 44150 677130 44170 677190
rect 44070 677110 44170 677130
rect 45100 677530 45200 678220
rect 45100 677470 45120 677530
rect 45180 677470 45200 677530
rect 45100 677360 45200 677470
rect 45100 677300 45120 677360
rect 45180 677300 45200 677360
rect 45100 677190 45200 677300
rect 45100 677130 45120 677190
rect 45180 677130 45200 677190
rect 45100 677110 45200 677130
rect 541364 677058 541484 677068
rect 41180 676980 41460 677020
rect 41180 676740 41200 676980
rect 41440 676740 41460 676980
rect 41180 675260 41460 676740
rect 41180 675020 41200 675260
rect 41440 675020 41460 675260
rect 41180 673540 41460 675020
rect 41180 673300 41200 673540
rect 41440 673300 41460 673540
rect 41180 672060 41460 673300
rect 41180 671820 41200 672060
rect 41440 671820 41460 672060
rect 41180 670340 41460 671820
rect 41180 670100 41200 670340
rect 41440 670100 41460 670340
rect 41180 668740 41460 670100
rect 41180 668500 41200 668740
rect 41440 668500 41460 668740
rect 41180 667020 41460 668500
rect 41180 666780 41200 667020
rect 41440 666780 41460 667020
rect 41180 665420 41460 666780
rect 41180 665180 41200 665420
rect 41440 665180 41460 665420
rect 41180 663700 41460 665180
rect 41180 663460 41200 663700
rect 41440 663460 41460 663700
rect 32800 663300 33100 663310
rect 32800 662990 33100 663000
rect 33300 663300 33600 663310
rect 33300 662990 33600 663000
rect 33800 663300 34100 663310
rect 33800 662990 34100 663000
rect 34300 663300 34600 663310
rect 34300 662990 34600 663000
rect 34800 663300 35100 663310
rect 34800 662990 35100 663000
rect 35300 663300 35600 663310
rect 35300 662990 35600 663000
rect 35800 663300 36100 663310
rect 35800 662990 36100 663000
rect 36300 663300 36600 663310
rect 36300 662990 36600 663000
rect 36800 663300 37100 663310
rect 36800 662990 37100 663000
rect 37300 663300 37600 663310
rect 37300 662990 37600 663000
rect 37800 663300 38100 663310
rect 37800 662990 38100 663000
rect 38300 663300 38600 663310
rect 38300 662990 38600 663000
rect 38800 663300 39100 663310
rect 38800 662990 39100 663000
rect 39300 663300 39600 663310
rect 39300 662990 39600 663000
rect 39800 663300 40100 663310
rect 39800 662990 40100 663000
rect 40300 663300 40600 663310
rect 40300 662990 40600 663000
rect 41180 663220 41460 663460
rect 41180 662980 41200 663220
rect 41440 662980 41460 663220
rect 41180 662880 41460 662980
rect 47880 676980 48160 677020
rect 47880 676740 47900 676980
rect 48140 676740 48160 676980
rect 541364 676928 541484 676938
rect 547734 677058 547854 677068
rect 547734 676928 547854 676938
rect 47880 675260 48160 676740
rect 47880 675020 47900 675260
rect 48140 675020 48160 675260
rect 47880 673540 48160 675020
rect 541364 674058 541484 674068
rect 541364 673928 541484 673938
rect 547734 674058 547854 674068
rect 547734 673928 547854 673938
rect 47880 673300 47900 673540
rect 48140 673300 48160 673540
rect 47880 672060 48160 673300
rect 47880 671820 47900 672060
rect 48140 671820 48160 672060
rect 47880 670340 48160 671820
rect 541364 671058 541484 671068
rect 541364 670928 541484 670938
rect 547734 671058 547854 671068
rect 547734 670928 547854 670938
rect 47880 670100 47900 670340
rect 48140 670100 48160 670340
rect 47880 668740 48160 670100
rect 47880 668500 47900 668740
rect 48140 668500 48160 668740
rect 47880 667020 48160 668500
rect 541364 668058 541484 668068
rect 541364 667928 541484 667938
rect 547734 668058 547854 668068
rect 547734 667928 547854 667938
rect 47880 666780 47900 667020
rect 48140 666780 48160 667020
rect 47880 665420 48160 666780
rect 47880 665180 47900 665420
rect 48140 665180 48160 665420
rect 47880 663700 48160 665180
rect 541364 665058 541484 665068
rect 541364 664928 541484 664938
rect 547734 665058 547854 665068
rect 547734 664928 547854 664938
rect 546294 663738 547464 663748
rect 47880 663460 47900 663700
rect 48140 663460 48160 663700
rect 47880 663220 48160 663460
rect 541744 663728 542914 663738
rect 541744 663308 542914 663318
rect 543254 663728 544424 663738
rect 543254 663308 544424 663318
rect 544774 663728 545944 663738
rect 546294 663318 547464 663328
rect 544774 663308 545944 663318
rect 47880 662980 47900 663220
rect 48140 662980 48160 663220
rect 47880 662880 48160 662980
<< via2 >>
rect 44010 695370 44280 695640
rect 45060 695370 45330 695640
rect 41460 695090 41530 695160
rect 41780 695090 41850 695160
rect 42090 695090 42160 695160
rect 42410 695090 42480 695160
rect 42720 695090 42790 695160
rect 43040 695090 43110 695160
rect 43360 695090 43430 695160
rect 43670 695090 43740 695160
rect 43990 695090 44060 695160
rect 44310 695090 44380 695160
rect 44620 695090 44690 695160
rect 44940 695090 45010 695160
rect 45250 695090 45320 695160
rect 45570 695090 45640 695160
rect 45890 695090 45960 695160
rect 46200 695090 46270 695160
rect 46520 695090 46590 695160
rect 46830 695090 46900 695160
rect 47150 695090 47220 695160
rect 47470 695090 47540 695160
rect 47780 695090 47850 695160
rect 36930 694850 37000 694920
rect 41460 694850 41530 694920
rect 41780 694850 41850 694920
rect 42090 694850 42160 694920
rect 42410 694850 42480 694920
rect 42720 694850 42790 694920
rect 43040 694850 43110 694920
rect 43360 694850 43430 694920
rect 43670 694850 43740 694920
rect 43990 694850 44060 694920
rect 44310 694850 44380 694920
rect 44620 694850 44690 694920
rect 44940 694850 45010 694920
rect 45250 694850 45320 694920
rect 45570 694850 45640 694920
rect 45890 694850 45960 694920
rect 46200 694850 46270 694920
rect 46520 694850 46590 694920
rect 46830 694850 46900 694920
rect 47150 694850 47220 694920
rect 47470 694850 47540 694920
rect 47780 694850 47850 694920
rect 52320 694850 52390 694920
rect 36820 694740 36890 694810
rect 52430 694740 52500 694810
rect 41620 694480 41690 694550
rect 41930 694480 42000 694550
rect 42250 694480 42320 694550
rect 42570 694480 42640 694550
rect 42880 694480 42950 694550
rect 43200 694480 43270 694550
rect 43510 694480 43580 694550
rect 43830 694480 43900 694550
rect 44150 694480 44220 694550
rect 44460 694480 44530 694550
rect 44780 694480 44850 694550
rect 45100 694480 45170 694550
rect 45410 694480 45480 694550
rect 45730 694480 45800 694550
rect 46040 694480 46110 694550
rect 46360 694480 46430 694550
rect 46680 694480 46750 694550
rect 46990 694480 47060 694550
rect 47310 694480 47380 694550
rect 47630 694480 47700 694550
rect 41620 694240 41690 694310
rect 41930 694240 42000 694310
rect 42250 694240 42320 694310
rect 42570 694240 42640 694310
rect 42880 694240 42950 694310
rect 43200 694240 43270 694310
rect 43510 694240 43580 694310
rect 43830 694240 43900 694310
rect 44150 694240 44220 694310
rect 44460 694240 44530 694310
rect 44780 694240 44850 694310
rect 45100 694240 45170 694310
rect 45410 694240 45480 694310
rect 45730 694240 45800 694310
rect 46040 694240 46110 694310
rect 46360 694240 46430 694310
rect 46680 694240 46750 694310
rect 46990 694240 47060 694310
rect 47310 694240 47380 694310
rect 47630 694240 47700 694310
rect 41620 693870 41690 693940
rect 38700 693360 38880 693460
rect 39120 693360 39300 693460
rect 44010 693730 44280 694000
rect 45060 693730 45330 694000
rect 42960 693420 43030 693490
rect 43280 693420 43350 693490
rect 43590 693420 43660 693490
rect 43910 693420 43980 693490
rect 44230 693420 44300 693490
rect 44540 693420 44610 693490
rect 44860 693420 44930 693490
rect 45180 693420 45250 693490
rect 45490 693420 45560 693490
rect 45810 693420 45880 693490
rect 46120 693420 46190 693490
rect 42960 693210 43030 693280
rect 43280 693210 43350 693280
rect 43590 693210 43660 693280
rect 43910 693210 43980 693280
rect 44230 693210 44300 693280
rect 44540 693210 44610 693280
rect 44860 693210 44930 693280
rect 45180 693210 45250 693280
rect 45490 693210 45560 693280
rect 45810 693210 45880 693280
rect 46120 693210 46190 693280
rect 42580 692760 42660 692840
rect 43120 692780 43190 692850
rect 43440 692780 43510 692850
rect 43750 692780 43820 692850
rect 44070 692780 44140 692850
rect 44390 692780 44460 692850
rect 44700 692780 44770 692850
rect 45020 692780 45090 692850
rect 45330 692780 45400 692850
rect 45650 692780 45720 692850
rect 45970 692780 46040 692850
rect 46280 692780 46350 692850
rect 42580 692580 42660 692660
rect 46640 692760 46720 692840
rect 43120 692570 43190 692640
rect 43440 692570 43510 692640
rect 43750 692570 43820 692640
rect 44070 692570 44140 692640
rect 44390 692570 44460 692640
rect 44700 692570 44770 692640
rect 45020 692570 45090 692640
rect 45330 692570 45400 692640
rect 45650 692570 45720 692640
rect 45970 692570 46040 692640
rect 46280 692570 46350 692640
rect 46640 692580 46720 692660
rect 43780 692130 44040 692390
rect 45280 692130 45540 692390
rect 42960 691870 43030 691940
rect 43280 691870 43350 691940
rect 43590 691870 43660 691940
rect 43910 691870 43980 691940
rect 44230 691870 44300 691940
rect 44540 691870 44610 691940
rect 44860 691870 44930 691940
rect 45170 691870 45240 691940
rect 45490 691870 45560 691940
rect 45810 691870 45880 691940
rect 46120 691870 46190 691940
rect 42960 691660 43030 691730
rect 43280 691660 43350 691730
rect 43590 691660 43660 691730
rect 43910 691660 43980 691730
rect 44230 691660 44300 691730
rect 44540 691660 44610 691730
rect 44860 691660 44930 691730
rect 45170 691660 45240 691730
rect 45490 691660 45560 691730
rect 45810 691660 45880 691730
rect 46120 691660 46190 691730
rect 43120 691240 43190 691310
rect 43440 691240 43510 691310
rect 43120 691030 43190 691100
rect 43750 691240 43820 691310
rect 44070 691240 44140 691310
rect 44380 691240 44450 691310
rect 44700 691240 44770 691310
rect 45020 691240 45090 691310
rect 45330 691240 45400 691310
rect 45650 691240 45720 691310
rect 45960 691240 46030 691310
rect 43440 691030 43510 691100
rect 42560 690250 42680 690370
rect 42560 690030 42680 690150
rect 42800 689690 42920 689810
rect 42800 689470 42920 689590
rect 42800 688730 42920 688850
rect 42000 688600 42100 688700
rect 42800 688510 42920 688630
rect 42000 688300 42100 688500
rect 42000 688100 42100 688200
rect 41620 687260 41690 687330
rect 41620 687100 41690 687170
rect 43750 691030 43820 691100
rect 44070 691030 44140 691100
rect 44380 691030 44450 691100
rect 44700 691030 44770 691100
rect 45020 691030 45090 691100
rect 45330 691030 45400 691100
rect 45650 691030 45720 691100
rect 46280 691240 46350 691310
rect 45960 691030 46030 691100
rect 44060 690310 44130 690380
rect 44380 690310 44450 690380
rect 44690 690310 44760 690380
rect 45010 690310 45080 690380
rect 44060 690020 44130 690090
rect 44380 690020 44450 690090
rect 44690 690020 44760 690090
rect 45010 690020 45080 690090
rect 44220 689750 44290 689820
rect 44530 689750 44600 689820
rect 44850 689750 44920 689820
rect 45170 689750 45240 689820
rect 44220 689460 44290 689530
rect 44530 689460 44600 689530
rect 44850 689460 44920 689530
rect 45170 689460 45240 689530
rect 44520 689030 44780 689290
rect 44060 688790 44130 688860
rect 44380 688790 44450 688860
rect 44690 688790 44760 688860
rect 45010 688790 45080 688860
rect 44060 688500 44130 688570
rect 44380 688500 44450 688570
rect 44690 688500 44760 688570
rect 45010 688500 45080 688570
rect 43440 688210 43510 688280
rect 44220 688230 44290 688300
rect 44530 688230 44600 688300
rect 44850 688230 44920 688300
rect 45170 688230 45240 688300
rect 46280 691030 46350 691100
rect 46620 690250 46740 690370
rect 47630 693870 47700 693940
rect 47200 690200 47300 690300
rect 46620 690030 46740 690150
rect 43440 687960 43510 688030
rect 45960 688210 46030 688280
rect 44220 687940 44290 688010
rect 44530 687940 44600 688010
rect 44850 687940 44920 688010
rect 45170 687940 45240 688010
rect 45960 687960 46030 688030
rect 46380 689690 46500 689810
rect 47200 689800 47300 690000
rect 46380 689470 46500 689590
rect 47200 689500 47300 689600
rect 46380 688730 46500 688850
rect 46380 688510 46500 688630
rect 44520 687510 44780 687770
rect 43070 687270 43140 687340
rect 43590 687270 43660 687340
rect 44100 687270 44170 687340
rect 44620 687270 44690 687340
rect 45130 687270 45200 687340
rect 45650 687270 45720 687340
rect 46170 687270 46240 687340
rect 43070 687090 43140 687160
rect 43590 687090 43660 687160
rect 44100 687090 44170 687160
rect 44620 687090 44690 687160
rect 45130 687090 45200 687160
rect 45650 687090 45720 687160
rect 46170 687090 46240 687160
rect 43330 686600 43400 686670
rect 43840 686600 43910 686670
rect 44360 686600 44430 686670
rect 44880 686600 44950 686670
rect 45390 686600 45460 686670
rect 45910 686600 45980 686670
rect 43330 686420 43400 686490
rect 43840 686420 43910 686490
rect 44360 686420 44430 686490
rect 44880 686420 44950 686490
rect 45390 686420 45460 686490
rect 45910 686420 45980 686490
rect 44530 686000 44780 686250
rect 42810 685750 42880 685820
rect 43330 685750 43400 685820
rect 43840 685750 43910 685820
rect 44360 685750 44430 685820
rect 44870 685750 44940 685820
rect 45390 685750 45460 685820
rect 45910 685750 45980 685820
rect 46420 685750 46490 685820
rect 42810 685570 42880 685640
rect 43330 685570 43400 685640
rect 43840 685570 43910 685640
rect 44360 685570 44430 685640
rect 44870 685570 44940 685640
rect 45390 685570 45460 685640
rect 45910 685570 45980 685640
rect 46420 685570 46490 685640
rect 49950 693360 50130 693460
rect 50370 693360 50550 693460
rect 541969 690892 542059 690962
rect 542139 690892 542229 690962
rect 544459 690892 544549 690962
rect 544629 690892 544719 690962
rect 541089 690602 541169 690682
rect 541239 690602 541319 690682
rect 541089 690062 541169 690142
rect 541239 690062 541319 690142
rect 541979 689842 542069 689912
rect 542119 689842 542209 689912
rect 541089 689522 541169 689602
rect 541239 689522 541319 689602
rect 541979 689302 542059 689382
rect 542149 689302 542229 689382
rect 534629 687992 534759 688132
rect 534879 687992 535009 688132
rect 546919 690892 546999 690972
rect 547089 690892 547169 690972
rect 566300 690900 566500 691100
rect 566700 690900 566900 691100
rect 567100 690900 567300 691100
rect 567500 690900 567700 691100
rect 567900 690900 568100 691100
rect 568300 690900 568500 691100
rect 568700 690900 568900 691100
rect 569100 690900 569300 691100
rect 569500 690900 569700 691100
rect 569900 690900 570100 691100
rect 570300 690900 570500 691100
rect 570700 690900 570900 691100
rect 571100 690900 571300 691100
rect 571500 690900 571700 691100
rect 543579 690602 543659 690682
rect 543729 690602 543809 690682
rect 543579 690062 543659 690142
rect 543729 690062 543809 690142
rect 544459 689842 544549 689912
rect 544619 689852 544709 689922
rect 543579 689522 543659 689602
rect 543729 689522 543809 689602
rect 544459 689302 544539 689382
rect 544629 689302 544709 689382
rect 542379 688922 542459 689002
rect 542489 688922 542569 689002
rect 542379 688312 542459 688392
rect 542489 688312 542569 688392
rect 541979 688142 542069 688222
rect 542139 688142 542229 688222
rect 47630 687260 47700 687330
rect 47630 687100 47700 687170
rect 542380 687750 542460 687830
rect 542500 687750 542580 687830
rect 546059 690602 546139 690682
rect 546209 690602 546289 690682
rect 546059 690062 546139 690142
rect 546209 690062 546289 690142
rect 546069 689522 546149 689602
rect 546209 689522 546289 689602
rect 546919 689852 546999 689922
rect 547089 689852 547169 689922
rect 546919 689302 546999 689382
rect 547089 689302 547169 689382
rect 544789 688922 544869 689002
rect 544899 688922 544979 689002
rect 544789 688332 544869 688412
rect 544899 688332 544979 688412
rect 544459 688142 544539 688212
rect 544629 688142 544709 688212
rect 544789 687752 544869 687832
rect 544899 687752 544979 687832
rect 566300 690500 566500 690700
rect 566700 690500 566900 690700
rect 567100 690500 567300 690700
rect 567500 690500 567700 690700
rect 567900 690500 568100 690700
rect 568300 690500 568500 690700
rect 568700 690500 568900 690700
rect 569100 690500 569300 690700
rect 569500 690500 569700 690700
rect 569900 690500 570100 690700
rect 570300 690500 570500 690700
rect 570700 690500 570900 690700
rect 571100 690500 571300 690700
rect 571500 690500 571700 690700
rect 566300 690100 566500 690300
rect 566700 690100 566900 690300
rect 567100 690100 567300 690300
rect 567500 690100 567700 690300
rect 567900 690100 568100 690300
rect 568300 690100 568500 690300
rect 568700 690100 568900 690300
rect 569100 690100 569300 690300
rect 569500 690100 569700 690300
rect 569900 690100 570100 690300
rect 570300 690100 570500 690300
rect 570700 690100 570900 690300
rect 571100 690100 571300 690300
rect 571500 690100 571700 690300
rect 566300 689700 566500 689900
rect 566700 689700 566900 689900
rect 567100 689700 567300 689900
rect 567500 689700 567700 689900
rect 567900 689700 568100 689900
rect 568300 689700 568500 689900
rect 568700 689700 568900 689900
rect 569100 689700 569300 689900
rect 569500 689700 569700 689900
rect 569900 689700 570100 689900
rect 570300 689700 570500 689900
rect 570700 689700 570900 689900
rect 571100 689700 571300 689900
rect 571500 689700 571700 689900
rect 566300 689300 566500 689500
rect 566700 689300 566900 689500
rect 567100 689300 567300 689500
rect 567500 689300 567700 689500
rect 567900 689300 568100 689500
rect 568300 689300 568500 689500
rect 568700 689300 568900 689500
rect 569100 689300 569300 689500
rect 569500 689300 569700 689500
rect 569900 689300 570100 689500
rect 570300 689300 570500 689500
rect 570700 689300 570900 689500
rect 571100 689300 571300 689500
rect 571500 689300 571700 689500
rect 547249 688912 547329 688992
rect 547359 688912 547439 688992
rect 547249 688332 547329 688412
rect 547359 688332 547439 688412
rect 546919 688142 546999 688212
rect 547089 688142 547169 688212
rect 547249 687752 547329 687832
rect 547359 687752 547439 687832
rect 554129 688162 554259 688302
rect 554389 688162 554519 688302
rect 538869 687542 538959 687652
rect 539029 687542 539119 687652
rect 43070 685080 43140 685150
rect 43580 685080 43650 685150
rect 44100 685080 44170 685150
rect 44620 685080 44690 685150
rect 45130 685080 45200 685150
rect 45650 685080 45720 685150
rect 46160 685080 46230 685150
rect 43070 684900 43140 684970
rect 43580 684900 43650 684970
rect 44100 684900 44170 684970
rect 44620 684900 44690 684970
rect 45130 684900 45200 684970
rect 45650 684900 45720 684970
rect 46160 684900 46230 684970
rect 540119 687062 540209 687142
rect 540299 687062 540389 687142
rect 540119 685982 540209 686062
rect 540299 685992 540389 686072
rect 535759 685122 535849 685252
rect 535969 685122 536059 685252
rect 542649 687062 542739 687142
rect 542809 687062 542899 687142
rect 542649 685982 542739 686062
rect 542809 685982 542899 686062
rect 44530 684470 44780 684720
rect 43840 683520 43920 683600
rect 44350 683520 44430 683600
rect 44870 683520 44950 683600
rect 45390 683520 45470 683600
rect 42260 683040 42340 683120
rect 42400 683040 42480 683120
rect 42540 683040 42620 683120
rect 44090 683040 44170 683120
rect 43840 682060 43920 682140
rect 43630 681840 43710 681920
rect 43630 681700 43710 681780
rect 44610 683040 44690 683120
rect 45130 683040 45210 683120
rect 44350 682060 44430 682140
rect 44870 682060 44950 682140
rect 44270 680400 44390 680520
rect 44890 680410 45010 680530
rect 46660 683040 46740 683120
rect 46800 683040 46880 683120
rect 46940 683040 47020 683120
rect 541089 684292 541169 684372
rect 541239 684292 541319 684372
rect 542379 685052 542459 685132
rect 542489 685052 542569 685132
rect 542279 684662 542389 684772
rect 543139 684662 543249 684772
rect 543579 684312 543659 684392
rect 543729 684312 543809 684392
rect 545119 687062 545209 687142
rect 545279 687062 545369 687142
rect 545119 685982 545209 686062
rect 545279 685982 545369 686062
rect 544789 685052 544869 685132
rect 544899 685052 544979 685132
rect 544349 684662 544459 684772
rect 545199 684662 545309 684772
rect 541569 683562 541679 683652
rect 45390 682060 45470 682140
rect 541509 682352 541629 682452
rect 542729 682352 542849 682452
rect 543939 682352 544059 682452
rect 546059 684312 546139 684392
rect 546199 684312 546279 684392
rect 548799 687522 548879 687602
rect 548969 687522 549049 687602
rect 547569 687062 547659 687142
rect 547729 687062 547819 687142
rect 547569 685982 547659 686062
rect 547729 685982 547819 686062
rect 547249 685062 547329 685142
rect 547359 685062 547439 685142
rect 550069 687062 550159 687142
rect 550229 687062 550319 687142
rect 550069 685982 550159 686062
rect 550229 685982 550319 686062
rect 553069 685152 553139 685242
rect 553229 685152 553299 685242
rect 546769 684662 546879 684772
rect 547649 684662 547759 684772
rect 546479 683562 546589 683652
rect 545159 682352 545279 682452
rect 45590 681840 45670 681920
rect 45590 681700 45670 681780
rect 541384 681318 541544 681478
rect 542444 681318 542604 681478
rect 543904 681318 544064 681478
rect 44070 679540 44160 679630
rect 44590 679540 44680 679630
rect 45100 679540 45190 679630
rect 44580 679160 44670 679250
rect 43830 678630 43890 678690
rect 44350 678630 44410 678690
rect 44830 678610 44960 678720
rect 541384 680738 541544 680898
rect 542444 680738 542604 680898
rect 543904 680738 544064 680898
rect 547599 682352 547719 682452
rect 561700 682000 561900 682200
rect 562100 682000 562300 682200
rect 562500 682000 562700 682200
rect 562900 682000 563100 682200
rect 563300 682000 563500 682200
rect 561700 681600 561900 681800
rect 562100 681600 562300 681800
rect 562500 681600 562700 681800
rect 562900 681600 563100 681800
rect 563300 681600 563500 681800
rect 545124 681318 545284 681478
rect 546604 681318 546764 681478
rect 547604 681318 547764 681478
rect 561700 681200 561900 681400
rect 562100 681200 562300 681400
rect 562500 681200 562700 681400
rect 562900 681200 563100 681400
rect 563300 681200 563500 681400
rect 545124 680738 545284 680898
rect 546604 680738 546764 680898
rect 547604 680738 547764 680898
rect 561700 680800 561900 681000
rect 562100 680800 562300 681000
rect 562500 680800 562700 681000
rect 562900 680800 563100 681000
rect 563300 680800 563500 681000
rect 543764 679368 543984 679518
rect 541404 678828 541584 678958
rect 542544 678828 542724 678958
rect 544284 679368 544504 679518
rect 544704 679368 544924 679518
rect 543524 678838 543704 678968
rect 45380 678630 45440 678690
rect 545254 679368 545474 679518
rect 544294 678838 544474 678968
rect 544734 678838 544914 678968
rect 561700 680400 561900 680600
rect 562100 680400 562300 680600
rect 562500 680400 562700 680600
rect 562900 680400 563100 680600
rect 563300 680400 563500 680600
rect 561700 680000 561900 680200
rect 562100 680000 562300 680200
rect 562500 680000 562700 680200
rect 562900 680000 563100 680200
rect 563300 680000 563500 680200
rect 561700 679600 561900 679800
rect 562100 679600 562300 679800
rect 562500 679600 562700 679800
rect 562900 679600 563100 679800
rect 563300 679600 563500 679800
rect 561700 679200 561900 679400
rect 562100 679200 562300 679400
rect 562500 679200 562700 679400
rect 562900 679200 563100 679400
rect 563300 679200 563500 679400
rect 545454 678828 545634 678958
rect 546524 678838 546704 678968
rect 547524 678838 547704 678968
rect 561700 678800 561900 679000
rect 562100 678800 562300 679000
rect 562500 678800 562700 679000
rect 562900 678800 563100 679000
rect 563300 678800 563500 679000
rect 561700 678400 561900 678600
rect 562100 678400 562300 678600
rect 562500 678400 562700 678600
rect 562900 678400 563100 678600
rect 563300 678400 563500 678600
rect 44090 678220 44150 678280
rect 44610 678220 44670 678280
rect 45120 678220 45180 678280
rect 44580 677720 44670 677810
rect 41200 676740 41440 676980
rect 41200 675020 41440 675260
rect 41200 673300 41440 673540
rect 41200 671820 41440 672060
rect 41200 670100 41440 670340
rect 41200 668500 41440 668740
rect 41200 666780 41440 667020
rect 41200 665180 41440 665420
rect 41200 663460 41440 663700
rect 32800 663000 33100 663300
rect 33300 663000 33600 663300
rect 33800 663000 34100 663300
rect 34300 663000 34600 663300
rect 34800 663000 35100 663300
rect 35300 663000 35600 663300
rect 35800 663000 36100 663300
rect 36300 663000 36600 663300
rect 36800 663000 37100 663300
rect 37300 663000 37600 663300
rect 37800 663000 38100 663300
rect 38300 663000 38600 663300
rect 38800 663000 39100 663300
rect 39300 663000 39600 663300
rect 39800 663000 40100 663300
rect 40300 663000 40600 663300
rect 47900 676740 48140 676980
rect 541364 676938 541484 677058
rect 547734 676938 547854 677058
rect 47900 675020 48140 675260
rect 541364 673938 541484 674058
rect 547734 673938 547854 674058
rect 47900 673300 48140 673540
rect 47900 671820 48140 672060
rect 541364 670938 541484 671058
rect 547734 670938 547854 671058
rect 47900 670100 48140 670340
rect 47900 668500 48140 668740
rect 541364 667938 541484 668058
rect 547734 667938 547854 668058
rect 47900 666780 48140 667020
rect 47900 665180 48140 665420
rect 541364 664938 541484 665058
rect 547734 664938 547854 665058
rect 47900 663460 48140 663700
rect 541744 663318 542914 663728
rect 543254 663318 544424 663728
rect 544774 663318 545944 663728
rect 546294 663328 547464 663738
<< metal3 >>
rect 16194 702300 21194 704800
rect 68194 702300 73194 704800
rect 465394 703700 470394 704800
rect 16200 702200 21200 702300
rect 16200 702000 16400 702200
rect 16600 702000 16800 702200
rect 17000 702000 17200 702200
rect 17400 702000 17600 702200
rect 17800 702000 18000 702200
rect 18200 702000 18400 702200
rect 18600 702000 18800 702200
rect 19000 702000 19200 702200
rect 19400 702000 19600 702200
rect 19800 702000 20000 702200
rect 20200 702000 20400 702200
rect 20600 702000 20800 702200
rect 21000 702000 21200 702200
rect 16200 701800 21200 702000
rect 16200 701600 16400 701800
rect 16600 701600 16800 701800
rect 17000 701600 17200 701800
rect 17400 701600 17600 701800
rect 17800 701600 18000 701800
rect 18200 701600 18400 701800
rect 18600 701600 18800 701800
rect 19000 701600 19200 701800
rect 19400 701600 19600 701800
rect 19800 701600 20000 701800
rect 20200 701600 20400 701800
rect 20600 701600 20800 701800
rect 21000 701600 21200 701800
rect 16200 701400 21200 701600
rect 16200 701200 16400 701400
rect 16600 701200 16800 701400
rect 17000 701200 17200 701400
rect 17400 701200 17600 701400
rect 17800 701200 18000 701400
rect 18200 701200 18400 701400
rect 18600 701200 18800 701400
rect 19000 701200 19200 701400
rect 19400 701200 19600 701400
rect 19800 701200 20000 701400
rect 20200 701200 20400 701400
rect 20600 701200 20800 701400
rect 21000 701200 21200 701400
rect 16200 701000 21200 701200
rect 68200 702200 73200 702300
rect 68200 702000 68400 702200
rect 68600 702000 68800 702200
rect 69000 702000 69200 702200
rect 69400 702000 69600 702200
rect 69800 702000 70000 702200
rect 70200 702000 70400 702200
rect 70600 702000 70800 702200
rect 71000 702000 71200 702200
rect 71400 702000 71600 702200
rect 71800 702000 72000 702200
rect 72200 702000 72400 702200
rect 72600 702000 72800 702200
rect 73000 702000 73200 702200
rect 68200 701800 73200 702000
rect 68200 701600 68400 701800
rect 68600 701600 68800 701800
rect 69000 701600 69200 701800
rect 69400 701600 69600 701800
rect 69800 701600 70000 701800
rect 70200 701600 70400 701800
rect 70600 701600 70800 701800
rect 71000 701600 71200 701800
rect 71400 701600 71600 701800
rect 71800 701600 72000 701800
rect 72200 701600 72400 701800
rect 72600 701600 72800 701800
rect 73000 701600 73200 701800
rect 68200 701400 73200 701600
rect 68200 701200 68400 701400
rect 68600 701200 68800 701400
rect 69000 701200 69200 701400
rect 69400 701200 69600 701400
rect 69800 701200 70000 701400
rect 70200 701200 70400 701400
rect 70600 701200 70800 701400
rect 71000 701200 71200 701400
rect 71400 701200 71600 701400
rect 71800 701200 72000 701400
rect 72200 701200 72400 701400
rect 72600 701200 72800 701400
rect 73000 701200 73200 701400
rect 16200 700800 16400 701000
rect 16600 700800 16800 701000
rect 17000 700800 17200 701000
rect 17400 700800 17600 701000
rect 17800 700800 18000 701000
rect 18200 700800 18400 701000
rect 18600 700800 18800 701000
rect 19000 700800 19200 701000
rect 19400 700800 19600 701000
rect 19800 700800 20000 701000
rect 20200 700800 20400 701000
rect 20600 700800 20800 701000
rect 21000 700800 21200 701000
rect 16200 700600 21200 700800
rect 16200 700400 16400 700600
rect 16600 700400 16800 700600
rect 17000 700400 17200 700600
rect 17400 700400 17600 700600
rect 17800 700400 18000 700600
rect 18200 700400 18400 700600
rect 18600 700400 18800 700600
rect 19000 700400 19200 700600
rect 19400 700400 19600 700600
rect 19800 700400 20000 700600
rect 20200 700400 20400 700600
rect 20600 700400 20800 700600
rect 21000 700400 21200 700600
rect 16200 700200 21200 700400
rect 16200 700000 16400 700200
rect 16600 700000 16800 700200
rect 17000 700000 17200 700200
rect 17400 700000 17600 700200
rect 17800 700000 18000 700200
rect 18200 700000 18400 700200
rect 18600 700000 18800 700200
rect 19000 700000 19200 700200
rect 19400 700000 19600 700200
rect 19800 700000 20000 700200
rect 20200 700000 20400 700200
rect 20600 700000 20800 700200
rect 21000 700000 21200 700200
rect 16200 699800 21200 700000
rect 37250 701109 40650 701129
rect 37250 701045 37278 701109
rect 40622 701045 40650 701109
rect 37250 697630 40650 701045
rect 41050 701109 44450 701129
rect 41050 701045 41078 701109
rect 44422 701045 44450 701109
rect 41050 697630 44450 701045
rect 44850 701109 48250 701129
rect 44850 701045 44878 701109
rect 48222 701045 48250 701109
rect 44850 697630 48250 701045
rect 48650 701109 52050 701129
rect 48650 701045 48678 701109
rect 52022 701045 52050 701109
rect 48650 697630 52050 701045
rect 68200 701000 73200 701200
rect 68200 700800 68400 701000
rect 68600 700800 68800 701000
rect 69000 700800 69200 701000
rect 69400 700800 69600 701000
rect 69800 700800 70000 701000
rect 70200 700800 70400 701000
rect 70600 700800 70800 701000
rect 71000 700800 71200 701000
rect 71400 700800 71600 701000
rect 71800 700800 72000 701000
rect 72200 700800 72400 701000
rect 72600 700800 72800 701000
rect 73000 700800 73200 701000
rect 68200 700600 73200 700800
rect 68200 700400 68400 700600
rect 68600 700400 68800 700600
rect 69000 700400 69200 700600
rect 69400 700400 69600 700600
rect 69800 700400 70000 700600
rect 70200 700400 70400 700600
rect 70600 700400 70800 700600
rect 71000 700400 71200 700600
rect 71400 700400 71600 700600
rect 71800 700400 72000 700600
rect 72200 700400 72400 700600
rect 72600 700400 72800 700600
rect 73000 700400 73200 700600
rect 68200 700200 73200 700400
rect 68200 700000 68400 700200
rect 68600 700000 68800 700200
rect 69000 700000 69200 700200
rect 69400 700000 69600 700200
rect 69800 700000 70000 700200
rect 70200 700000 70400 700200
rect 70600 700000 70800 700200
rect 71000 700000 71200 700200
rect 71400 700000 71600 700200
rect 71800 700000 72000 700200
rect 72200 700000 72400 700200
rect 72600 700000 72800 700200
rect 73000 700000 73200 700200
rect 68200 699800 73200 700000
rect 44000 695640 44290 695645
rect 44000 695370 44010 695640
rect 44280 695370 44290 695640
rect 44000 695365 44290 695370
rect 45050 695640 45340 695645
rect 45050 695370 45060 695640
rect 45330 695370 45340 695640
rect 45050 695365 45340 695370
rect 41460 695165 47850 695170
rect 41450 695160 47860 695165
rect 41450 695090 41460 695160
rect 41530 695090 41780 695160
rect 41850 695140 42090 695160
rect 42160 695090 42410 695160
rect 42480 695090 42720 695160
rect 42790 695090 43040 695160
rect 43110 695090 43360 695160
rect 43430 695090 43670 695160
rect 43740 695130 43990 695160
rect 41450 695085 41840 695090
rect 36800 694920 37020 694940
rect 41460 694925 41840 695085
rect 36800 694850 36930 694920
rect 37000 694850 37020 694920
rect 36800 694810 37020 694850
rect 41450 694920 41840 694925
rect 42090 694920 43740 695090
rect 41450 694850 41460 694920
rect 41530 694850 41780 694920
rect 41850 694850 42090 694890
rect 42160 694850 42410 694920
rect 42480 694850 42720 694920
rect 42790 694850 43040 694920
rect 43110 694850 43360 694920
rect 43430 694850 43670 694920
rect 44060 695090 44310 695160
rect 44380 695090 44620 695160
rect 44690 695090 44940 695160
rect 45010 695090 45250 695160
rect 45320 695130 45570 695160
rect 43990 694920 45320 695090
rect 43740 694850 43990 694880
rect 44060 694850 44310 694920
rect 44380 694850 44620 694920
rect 44690 694850 44940 694920
rect 45010 694850 45250 694920
rect 45640 695090 45890 695160
rect 45960 695090 46200 695160
rect 46270 695090 46520 695160
rect 46590 695090 46830 695160
rect 46900 695090 47150 695160
rect 47220 695130 47470 695160
rect 45570 694920 47220 695090
rect 45320 694850 45570 694880
rect 45640 694850 45890 694920
rect 45960 694850 46200 694920
rect 46270 694850 46520 694920
rect 46590 694850 46830 694920
rect 46900 694850 47150 694920
rect 47540 695090 47780 695160
rect 47850 695090 47860 695160
rect 47470 695085 47860 695090
rect 47470 694925 47850 695085
rect 47470 694920 47860 694925
rect 47220 694850 47470 694880
rect 47540 694850 47780 694920
rect 47850 694850 47860 694920
rect 41450 694845 47860 694850
rect 52300 694920 52520 694940
rect 52300 694850 52320 694920
rect 52390 694850 52520 694920
rect 41460 694840 47850 694845
rect 36800 694740 36820 694810
rect 36890 694740 37020 694810
rect 36800 694720 37020 694740
rect 52300 694810 52520 694850
rect 52300 694740 52430 694810
rect 52500 694740 52520 694810
rect 52300 694720 52520 694740
rect 41460 694550 47850 694560
rect 41460 694480 41620 694550
rect 41690 694480 41930 694550
rect 42000 694480 42250 694550
rect 42320 694480 42570 694550
rect 42640 694480 42880 694550
rect 42950 694480 43200 694550
rect 43270 694480 43510 694550
rect 43580 694480 43830 694550
rect 43900 694480 44150 694550
rect 44220 694480 44460 694550
rect 44530 694480 44780 694550
rect 44850 694480 45100 694550
rect 45170 694480 45410 694550
rect 45480 694480 45730 694550
rect 45800 694480 46040 694550
rect 46110 694480 46360 694550
rect 46430 694480 46680 694550
rect 46750 694480 46990 694550
rect 47060 694480 47310 694550
rect 47380 694480 47630 694550
rect 47700 694480 47850 694550
rect 41460 694310 47850 694480
rect 41460 694240 41620 694310
rect 41690 694240 41930 694310
rect 42000 694240 42250 694310
rect 42320 694240 42570 694310
rect 42640 694240 42880 694310
rect 42950 694240 43200 694310
rect 43270 694240 43510 694310
rect 43580 694240 43830 694310
rect 43900 694240 44150 694310
rect 44220 694240 44460 694310
rect 44530 694240 44780 694310
rect 44850 694240 45100 694310
rect 45170 694240 45410 694310
rect 45480 694240 45730 694310
rect 45800 694240 46040 694310
rect 46110 694240 46360 694310
rect 46430 694240 46680 694310
rect 46750 694240 46990 694310
rect 47060 694240 47310 694310
rect 47380 694240 47630 694310
rect 47700 694240 47850 694310
rect 41460 694230 47850 694240
rect 44000 694000 44290 694005
rect 40690 693960 41720 693980
rect 40690 693860 40710 693960
rect 40800 693860 40900 693960
rect 40990 693940 41720 693960
rect 40990 693870 41620 693940
rect 41690 693870 41720 693940
rect 40990 693860 41720 693870
rect 40690 693840 41720 693860
rect 44000 693730 44010 694000
rect 44280 693730 44290 694000
rect 44000 693725 44290 693730
rect 45050 694000 45340 694005
rect 45050 693730 45060 694000
rect 45330 693730 45340 694000
rect 47600 693960 48620 693980
rect 47600 693940 48320 693960
rect 47600 693870 47630 693940
rect 47700 693870 48320 693940
rect 47600 693860 48320 693870
rect 48410 693860 48510 693960
rect 48600 693860 48620 693960
rect 47600 693840 48620 693860
rect 45050 693725 45340 693730
rect 42960 693495 46350 693500
rect 42950 693490 46350 693495
rect 38690 693460 38890 693465
rect 38690 693360 38700 693460
rect 38880 693360 38890 693460
rect 38690 693355 38890 693360
rect 39110 693460 39310 693465
rect 39110 693360 39120 693460
rect 39300 693360 39310 693460
rect 42950 693420 42960 693490
rect 43030 693420 43280 693490
rect 43350 693480 43590 693490
rect 43660 693420 43910 693490
rect 43980 693420 44230 693490
rect 44300 693420 44540 693490
rect 44610 693480 44860 693490
rect 44930 693420 45180 693490
rect 45250 693420 45490 693490
rect 45560 693420 45810 693490
rect 45880 693480 46120 693490
rect 46190 693420 46350 693490
rect 42950 693415 43340 693420
rect 39110 693355 39310 693360
rect 42960 693285 43340 693415
rect 42950 693280 43340 693285
rect 43600 693280 44610 693420
rect 44870 693280 45870 693420
rect 46130 693280 46350 693420
rect 49940 693460 50140 693465
rect 49940 693360 49950 693460
rect 50130 693360 50140 693460
rect 49940 693355 50140 693360
rect 50360 693460 50560 693465
rect 50360 693360 50370 693460
rect 50550 693360 50560 693460
rect 50360 693355 50560 693360
rect 42950 693210 42960 693280
rect 43030 693210 43280 693280
rect 43350 693210 43590 693220
rect 43660 693210 43910 693280
rect 43980 693210 44230 693280
rect 44300 693210 44540 693280
rect 44610 693210 44860 693220
rect 44930 693210 45180 693280
rect 45250 693210 45490 693280
rect 45560 693210 45810 693280
rect 45880 693210 46120 693220
rect 46190 693210 46350 693280
rect 42950 693205 46350 693210
rect 42960 693200 46350 693205
rect 42540 692850 46760 692860
rect 42540 692840 43120 692850
rect 42540 692760 42580 692840
rect 42660 692780 43120 692840
rect 43190 692780 43440 692850
rect 43510 692780 43750 692850
rect 43820 692780 44070 692850
rect 44140 692780 44390 692850
rect 44460 692780 44700 692850
rect 44770 692780 45020 692850
rect 45090 692780 45330 692850
rect 45400 692780 45650 692850
rect 45720 692780 45970 692850
rect 46040 692780 46280 692850
rect 46350 692840 46760 692850
rect 46350 692780 46640 692840
rect 42660 692760 46640 692780
rect 46720 692760 46760 692840
rect 42540 692660 46760 692760
rect 42540 692580 42580 692660
rect 42660 692640 46640 692660
rect 42660 692580 43120 692640
rect 42540 692570 43120 692580
rect 43190 692570 43440 692640
rect 43510 692570 43750 692640
rect 43820 692570 44070 692640
rect 44140 692570 44390 692640
rect 44460 692570 44700 692640
rect 44770 692570 45020 692640
rect 45090 692570 45330 692640
rect 45400 692570 45650 692640
rect 45720 692570 45970 692640
rect 46040 692570 46280 692640
rect 46350 692580 46640 692640
rect 46720 692580 46760 692660
rect 46350 692570 46760 692580
rect 42540 692560 46760 692570
rect 43770 692390 44050 692395
rect 43770 692130 43780 692390
rect 44040 692130 44050 692390
rect 43770 692125 44050 692130
rect 45270 692390 45550 692395
rect 45270 692130 45280 692390
rect 45540 692130 45550 692390
rect 45270 692125 45550 692130
rect 46320 691950 62200 692040
rect 42960 691945 62200 691950
rect 42950 691940 62200 691945
rect 42950 691870 42960 691940
rect 43030 691870 43280 691940
rect 43350 691930 43590 691940
rect 43660 691870 43910 691940
rect 43980 691870 44230 691940
rect 44300 691870 44540 691940
rect 44610 691930 44860 691940
rect 44930 691870 45170 691940
rect 45240 691870 45490 691940
rect 45560 691870 45810 691940
rect 45880 691930 46120 691940
rect 46190 691900 62200 691940
rect 46190 691870 58000 691900
rect 42950 691865 43340 691870
rect 42960 691735 43340 691865
rect 42950 691730 43340 691735
rect 43600 691730 44610 691870
rect 44870 691730 45870 691870
rect 46130 691730 58000 691870
rect 42950 691660 42960 691730
rect 43030 691660 43280 691730
rect 43350 691660 43590 691670
rect 43660 691660 43910 691730
rect 43980 691660 44230 691730
rect 44300 691660 44540 691730
rect 44610 691660 44860 691670
rect 44930 691660 45170 691730
rect 45240 691660 45490 691730
rect 45560 691660 45810 691730
rect 46190 691700 58000 691730
rect 58200 691700 58400 691900
rect 58600 691700 58800 691900
rect 59000 691700 59200 691900
rect 59400 691700 59600 691900
rect 59800 691700 60000 691900
rect 60200 691700 60400 691900
rect 60600 691700 60800 691900
rect 61000 691700 61200 691900
rect 61400 691700 61600 691900
rect 61800 691700 62200 691900
rect 45880 691660 46120 691670
rect 46190 691660 62200 691700
rect 42950 691655 62200 691660
rect 42960 691650 62200 691655
rect 46320 691560 62200 691650
rect 42960 691315 46350 691320
rect 42960 691310 46360 691315
rect 42960 691240 43120 691310
rect 43190 691240 43440 691310
rect 43510 691240 43750 691310
rect 43820 691240 44070 691310
rect 44140 691240 44380 691310
rect 44450 691240 44700 691310
rect 44770 691240 45020 691310
rect 45090 691240 45330 691310
rect 45400 691240 45650 691310
rect 45720 691240 45960 691310
rect 46030 691240 46280 691310
rect 46350 691240 46360 691310
rect 42960 691235 46360 691240
rect 42960 691105 46350 691235
rect 42960 691100 46360 691105
rect 42960 691030 43120 691100
rect 43190 691030 43440 691100
rect 43510 691030 43750 691100
rect 43820 691030 44070 691100
rect 44140 691030 44380 691100
rect 44450 691030 44700 691100
rect 44770 691030 45020 691100
rect 45090 691030 45330 691100
rect 45400 691030 45650 691100
rect 45720 691030 45960 691100
rect 46030 691030 46280 691100
rect 46350 691030 46360 691100
rect 42960 691025 46360 691030
rect 42960 691020 46350 691025
rect 465100 690500 470600 703700
rect 566594 703100 571594 704800
rect 534609 694992 535049 695042
rect 534609 694862 534639 694992
rect 534739 694862 534899 694992
rect 534999 694862 535049 694992
rect 554109 694992 554539 695052
rect 465100 690400 534200 690500
rect 42540 690380 46760 690390
rect 42540 690370 44060 690380
rect 42540 690250 42560 690370
rect 42680 690310 44060 690370
rect 44130 690310 44380 690380
rect 44450 690310 44690 690380
rect 44760 690310 45010 690380
rect 45080 690370 46760 690380
rect 45080 690310 46620 690370
rect 42680 690250 46620 690310
rect 46740 690250 46760 690370
rect 42540 690150 46760 690250
rect 42540 690030 42560 690150
rect 42680 690090 46620 690150
rect 42680 690030 44060 690090
rect 42540 690020 44060 690030
rect 44130 690020 44380 690090
rect 44450 690020 44690 690090
rect 44760 690020 45010 690090
rect 45080 690030 46620 690090
rect 46740 690030 46760 690150
rect 45080 690020 46760 690030
rect 42540 690010 46760 690020
rect 47100 690300 73200 690400
rect 47100 690200 47200 690300
rect 47300 690200 73200 690300
rect 47100 690000 68400 690200
rect 68600 690000 68800 690200
rect 69000 690000 69200 690200
rect 69400 690000 69600 690200
rect 69800 690000 70000 690200
rect 70200 690000 70400 690200
rect 70600 690000 70800 690200
rect 71000 690000 71200 690200
rect 71400 690000 71600 690200
rect 71800 690000 72000 690200
rect 72200 690000 72400 690200
rect 72600 690000 72800 690200
rect 73000 690000 73200 690200
rect 42780 689820 46520 689830
rect 42780 689810 44220 689820
rect 42780 689690 42800 689810
rect 42920 689750 44220 689810
rect 44290 689750 44530 689820
rect 44600 689750 44850 689820
rect 44920 689750 45170 689820
rect 45240 689810 46520 689820
rect 45240 689750 46380 689810
rect 42920 689690 46380 689750
rect 46500 689690 46520 689810
rect 42780 689590 46520 689690
rect 42780 689470 42800 689590
rect 42920 689530 46380 689590
rect 42920 689470 44220 689530
rect 42780 689460 44220 689470
rect 44290 689460 44530 689530
rect 44600 689460 44850 689530
rect 44920 689460 45170 689530
rect 45240 689470 46380 689530
rect 46500 689470 46520 689590
rect 45240 689460 46520 689470
rect 42780 689450 46520 689460
rect 47100 689800 47200 690000
rect 47300 689800 73200 690000
rect 47100 689600 68400 689800
rect 68600 689600 68800 689800
rect 69000 689600 69200 689800
rect 69400 689600 69600 689800
rect 69800 689600 70000 689800
rect 70200 689600 70400 689800
rect 70600 689600 70800 689800
rect 71000 689600 71200 689800
rect 71400 689600 71600 689800
rect 71800 689600 72000 689800
rect 72200 689600 72400 689800
rect 72600 689600 72800 689800
rect 73000 689600 73200 689800
rect 47100 689500 47200 689600
rect 47300 689500 73200 689600
rect 47100 689400 73200 689500
rect 465100 690200 532300 690400
rect 532500 690200 532700 690400
rect 532900 690200 533100 690400
rect 533300 690200 533500 690400
rect 533700 690200 533900 690400
rect 534100 690200 534200 690400
rect 465100 690100 534200 690200
rect 465100 689900 532300 690100
rect 532500 689900 532700 690100
rect 532900 689900 533100 690100
rect 533300 689900 533500 690100
rect 533700 689900 533900 690100
rect 534100 689900 534200 690100
rect 465100 689700 534200 689900
rect 465100 689500 532300 689700
rect 532500 689500 532700 689700
rect 532900 689500 533100 689700
rect 533300 689500 533500 689700
rect 533700 689500 533900 689700
rect 534100 689500 534200 689700
rect 465100 689300 534200 689500
rect 44510 689290 44790 689295
rect 44510 689030 44520 689290
rect 44780 689030 44790 689290
rect 44510 689025 44790 689030
rect 465100 689100 532300 689300
rect 532500 689100 532700 689300
rect 532900 689100 533100 689300
rect 533300 689100 533500 689300
rect 533700 689100 533900 689300
rect 534100 689100 534200 689300
rect 465100 688900 534200 689100
rect 42780 688860 46520 688870
rect 42780 688850 44060 688860
rect 16200 688700 42200 688800
rect 16200 688500 16400 688700
rect 16600 688500 16800 688700
rect 17000 688500 17200 688700
rect 17400 688500 17600 688700
rect 17800 688500 18000 688700
rect 18200 688500 18400 688700
rect 18600 688500 18800 688700
rect 19000 688500 19200 688700
rect 19400 688500 19600 688700
rect 19800 688500 20000 688700
rect 20200 688500 20400 688700
rect 20600 688500 20800 688700
rect 21000 688600 42000 688700
rect 42100 688600 42200 688700
rect 21000 688500 42200 688600
rect 16200 688300 42000 688500
rect 42100 688300 42200 688500
rect 42780 688730 42800 688850
rect 42920 688790 44060 688850
rect 44130 688790 44380 688860
rect 44450 688790 44690 688860
rect 44760 688790 45010 688860
rect 45080 688850 46520 688860
rect 45080 688790 46380 688850
rect 42920 688730 46380 688790
rect 46500 688730 46520 688850
rect 42780 688630 46520 688730
rect 42780 688510 42800 688630
rect 42920 688570 46380 688630
rect 42920 688510 44060 688570
rect 42780 688500 44060 688510
rect 44130 688500 44380 688570
rect 44450 688500 44690 688570
rect 44760 688500 45010 688570
rect 45080 688510 46380 688570
rect 46500 688510 46520 688630
rect 465100 688700 532300 688900
rect 532500 688700 532700 688900
rect 532900 688700 533100 688900
rect 533300 688700 533500 688900
rect 533700 688700 533900 688900
rect 534100 688700 534200 688900
rect 465100 688600 534200 688700
rect 45080 688500 46520 688510
rect 42780 688490 46520 688500
rect 16200 688100 16400 688300
rect 16600 688100 16800 688300
rect 17000 688100 17200 688300
rect 17400 688100 17600 688300
rect 17800 688100 18000 688300
rect 18200 688100 18400 688300
rect 18600 688100 18800 688300
rect 19000 688100 19200 688300
rect 19400 688100 19600 688300
rect 19800 688100 20000 688300
rect 20200 688100 20400 688300
rect 20600 688100 20800 688300
rect 21000 688200 42200 688300
rect 21000 688100 42000 688200
rect 42100 688100 42200 688200
rect 16200 688000 42200 688100
rect 43410 688300 46060 688310
rect 43410 688280 44220 688300
rect 43410 688210 43440 688280
rect 43510 688230 44220 688280
rect 44290 688230 44530 688300
rect 44600 688230 44850 688300
rect 44920 688230 45170 688300
rect 45240 688280 46060 688300
rect 45240 688230 45960 688280
rect 43510 688210 45960 688230
rect 46030 688210 46060 688280
rect 43410 688030 46060 688210
rect 43410 687960 43440 688030
rect 43510 688010 45960 688030
rect 43510 687960 44220 688010
rect 43410 687940 44220 687960
rect 44290 687940 44530 688010
rect 44600 687940 44850 688010
rect 44920 687940 45170 688010
rect 45240 687960 45960 688010
rect 46030 687960 46060 688030
rect 534609 688132 535049 694862
rect 537169 694921 540569 694941
rect 537169 694857 537197 694921
rect 540541 694857 540569 694921
rect 537169 691442 540569 694857
rect 540969 694921 544369 694941
rect 540969 694857 540997 694921
rect 544341 694857 544369 694921
rect 540969 691442 544369 694857
rect 544769 694921 548169 694941
rect 544769 694857 544797 694921
rect 548141 694857 548169 694921
rect 544769 691442 548169 694857
rect 548569 694921 551969 694941
rect 548569 694857 548597 694921
rect 551941 694857 551969 694921
rect 548569 691442 551969 694857
rect 554109 694862 554129 694992
rect 554239 694862 554389 694992
rect 554499 694862 554539 694992
rect 539919 690972 551499 691212
rect 539919 690962 546919 690972
rect 539919 690892 541969 690962
rect 542059 690892 542139 690962
rect 542229 690892 544459 690962
rect 544549 690892 544629 690962
rect 544719 690892 546919 690962
rect 546999 690892 547089 690972
rect 547169 690892 551499 690972
rect 539919 690852 551499 690892
rect 541069 690682 541339 690702
rect 541069 690602 541089 690682
rect 541169 690602 541239 690682
rect 541319 690602 541339 690682
rect 541069 690582 541339 690602
rect 543559 690682 543829 690692
rect 543559 690602 543579 690682
rect 543659 690602 543729 690682
rect 543809 690602 543829 690682
rect 543559 690582 543829 690602
rect 546039 690682 546309 690702
rect 546039 690602 546059 690682
rect 546139 690602 546209 690682
rect 546289 690602 546309 690682
rect 546039 690582 546309 690602
rect 541069 690142 541339 690162
rect 541069 690062 541089 690142
rect 541169 690062 541239 690142
rect 541319 690062 541339 690142
rect 541069 690042 541339 690062
rect 543559 690142 543829 690152
rect 543559 690062 543579 690142
rect 543659 690062 543729 690142
rect 543809 690062 543829 690142
rect 543559 690042 543829 690062
rect 546039 690142 546309 690162
rect 546039 690062 546059 690142
rect 546139 690062 546209 690142
rect 546289 690062 546309 690142
rect 546039 690042 546309 690062
rect 551089 689982 551499 690852
rect 539679 689922 551499 689982
rect 539679 689912 544619 689922
rect 539679 689842 541979 689912
rect 542069 689842 542119 689912
rect 542209 689842 544459 689912
rect 544549 689852 544619 689912
rect 544709 689852 546919 689922
rect 546999 689852 547089 689922
rect 547169 689852 551499 689922
rect 544549 689842 551499 689852
rect 539679 689752 551499 689842
rect 541069 689602 541339 689632
rect 541069 689522 541089 689602
rect 541169 689522 541239 689602
rect 541319 689522 541339 689602
rect 541069 689502 541339 689522
rect 543559 689602 543829 689612
rect 543559 689522 543579 689602
rect 543659 689522 543729 689602
rect 543809 689522 543829 689602
rect 543559 689502 543829 689522
rect 546039 689602 546309 689632
rect 546039 689522 546069 689602
rect 546149 689522 546209 689602
rect 546289 689522 546309 689602
rect 546039 689502 546309 689522
rect 551089 689392 551499 689752
rect 540069 689382 551499 689392
rect 540069 689302 541979 689382
rect 542059 689302 542149 689382
rect 542229 689302 544459 689382
rect 544539 689302 544629 689382
rect 544709 689302 546919 689382
rect 546999 689302 547089 689382
rect 547169 689302 551499 689382
rect 540069 689172 551499 689302
rect 542359 689002 542589 689022
rect 542359 688922 542379 689002
rect 542459 688922 542489 689002
rect 542569 688922 542589 689002
rect 542359 688892 542589 688922
rect 544769 689002 544999 689022
rect 544769 688922 544789 689002
rect 544869 688922 544899 689002
rect 544979 688922 544999 689002
rect 544769 688912 544999 688922
rect 547229 688992 547459 689002
rect 547229 688912 547249 688992
rect 547329 688912 547359 688992
rect 547439 688912 547459 688992
rect 547229 688892 547459 688912
rect 544769 688412 544999 688422
rect 542359 688392 542589 688402
rect 542359 688312 542379 688392
rect 542459 688312 542489 688392
rect 542569 688312 542589 688392
rect 544769 688332 544789 688412
rect 544869 688332 544899 688412
rect 544979 688332 544999 688412
rect 544769 688312 544999 688332
rect 547229 688412 547459 688422
rect 547229 688332 547249 688412
rect 547329 688332 547359 688412
rect 547439 688332 547459 688412
rect 547229 688312 547459 688332
rect 542359 688302 542589 688312
rect 551089 688232 551499 689172
rect 534609 687992 534629 688132
rect 534759 687992 534879 688132
rect 535009 687992 535049 688132
rect 539989 688222 551499 688232
rect 539989 688142 541979 688222
rect 542069 688142 542139 688222
rect 542229 688212 551499 688222
rect 542229 688142 544459 688212
rect 544539 688142 544629 688212
rect 544709 688142 546919 688212
rect 546999 688142 547089 688212
rect 547169 688142 551499 688212
rect 554109 688302 554539 694862
rect 566260 691320 571820 703100
rect 566260 691100 571840 691320
rect 566260 690900 566300 691100
rect 566500 690900 566700 691100
rect 566900 690900 567100 691100
rect 567300 690900 567500 691100
rect 567700 690900 567900 691100
rect 568100 690900 568300 691100
rect 568500 690900 568700 691100
rect 568900 690900 569100 691100
rect 569300 690900 569500 691100
rect 569700 690900 569900 691100
rect 570100 690900 570300 691100
rect 570500 690900 570700 691100
rect 570900 690900 571100 691100
rect 571300 690900 571500 691100
rect 571700 690900 571840 691100
rect 566260 690700 571840 690900
rect 566260 690500 566300 690700
rect 566500 690500 566700 690700
rect 566900 690500 567100 690700
rect 567300 690500 567500 690700
rect 567700 690500 567900 690700
rect 568100 690500 568300 690700
rect 568500 690500 568700 690700
rect 568900 690500 569100 690700
rect 569300 690500 569500 690700
rect 569700 690500 569900 690700
rect 570100 690500 570300 690700
rect 570500 690500 570700 690700
rect 570900 690500 571100 690700
rect 571300 690500 571500 690700
rect 571700 690500 571840 690700
rect 566260 690300 571840 690500
rect 566260 690100 566300 690300
rect 566500 690100 566700 690300
rect 566900 690100 567100 690300
rect 567300 690100 567500 690300
rect 567700 690100 567900 690300
rect 568100 690100 568300 690300
rect 568500 690100 568700 690300
rect 568900 690100 569100 690300
rect 569300 690100 569500 690300
rect 569700 690100 569900 690300
rect 570100 690100 570300 690300
rect 570500 690100 570700 690300
rect 570900 690100 571100 690300
rect 571300 690100 571500 690300
rect 571700 690100 571840 690300
rect 566260 689900 571840 690100
rect 566260 689700 566300 689900
rect 566500 689700 566700 689900
rect 566900 689700 567100 689900
rect 567300 689700 567500 689900
rect 567700 689700 567900 689900
rect 568100 689700 568300 689900
rect 568500 689700 568700 689900
rect 568900 689700 569100 689900
rect 569300 689700 569500 689900
rect 569700 689700 569900 689900
rect 570100 689700 570300 689900
rect 570500 689700 570700 689900
rect 570900 689700 571100 689900
rect 571300 689700 571500 689900
rect 571700 689700 571840 689900
rect 566260 689520 571840 689700
rect 566260 689500 571820 689520
rect 566260 689300 566300 689500
rect 566500 689300 566700 689500
rect 566900 689300 567100 689500
rect 567300 689300 567500 689500
rect 567700 689300 567900 689500
rect 568100 689300 568300 689500
rect 568500 689300 568700 689500
rect 568900 689300 569100 689500
rect 569300 689300 569500 689500
rect 569700 689300 569900 689500
rect 570100 689300 570300 689500
rect 570500 689300 570700 689500
rect 570900 689300 571100 689500
rect 571300 689300 571500 689500
rect 571700 689300 571820 689500
rect 566260 689200 571820 689300
rect 554109 688162 554129 688302
rect 554259 688162 554389 688302
rect 554519 688162 554539 688302
rect 554109 688152 554539 688162
rect 539989 688052 551499 688142
rect 534609 687972 535049 687992
rect 45240 687940 46060 687960
rect 43410 687930 46060 687940
rect 542350 687830 542600 687880
rect 44510 687770 44790 687775
rect 44510 687510 44520 687770
rect 44780 687510 44790 687770
rect 542350 687750 542380 687830
rect 542460 687750 542500 687830
rect 542580 687750 542600 687830
rect 542350 687730 542600 687750
rect 544769 687832 544999 687842
rect 544769 687752 544789 687832
rect 544869 687752 544899 687832
rect 544979 687752 544999 687832
rect 544769 687732 544999 687752
rect 547229 687832 547459 687842
rect 547229 687752 547249 687832
rect 547329 687752 547359 687832
rect 547439 687752 547459 687832
rect 547229 687732 547459 687752
rect 538849 687652 539139 687672
rect 538849 687542 538869 687652
rect 538959 687542 539029 687652
rect 539119 687542 539139 687652
rect 538849 687532 539139 687542
rect 548779 687602 549071 687612
rect 548779 687522 548799 687602
rect 548879 687522 548969 687602
rect 549049 687522 549071 687602
rect 548779 687514 549071 687522
rect 44510 687505 44790 687510
rect 36600 687340 47800 687400
rect 36600 687330 43070 687340
rect 36600 687300 41620 687330
rect 36600 687100 36800 687300
rect 37000 687100 37200 687300
rect 37400 687100 37600 687300
rect 37800 687100 38000 687300
rect 38200 687260 41620 687300
rect 41690 687270 43070 687330
rect 43140 687270 43590 687340
rect 43660 687270 44100 687340
rect 44170 687270 44620 687340
rect 44690 687270 45130 687340
rect 45200 687270 45650 687340
rect 45720 687270 46170 687340
rect 46240 687330 47800 687340
rect 46240 687270 47630 687330
rect 41690 687260 47630 687270
rect 47700 687260 47800 687330
rect 551089 687322 551499 688052
rect 38200 687170 47800 687260
rect 38200 687100 41620 687170
rect 41690 687160 47630 687170
rect 41690 687100 43070 687160
rect 36600 687090 43070 687100
rect 43140 687090 43590 687160
rect 43660 687090 44100 687160
rect 44170 687090 44620 687160
rect 44690 687090 45130 687160
rect 45200 687090 45650 687160
rect 45720 687090 46170 687160
rect 46240 687100 47630 687160
rect 47700 687100 47800 687170
rect 46240 687090 47800 687100
rect 36600 687000 47800 687090
rect 537839 687300 551499 687322
rect 537839 687200 551200 687300
rect 537839 687142 549900 687200
rect 550100 687142 550200 687200
rect 537839 687062 540119 687142
rect 540209 687062 540299 687142
rect 540389 687062 542649 687142
rect 542739 687062 542809 687142
rect 542899 687062 545119 687142
rect 545209 687062 545279 687142
rect 545369 687062 547569 687142
rect 547659 687062 547729 687142
rect 547819 687062 549900 687142
rect 550159 687062 550200 687142
rect 537839 687000 549900 687062
rect 550100 687000 550200 687062
rect 550400 687000 550500 687200
rect 550700 687000 550800 687200
rect 551000 687100 551200 687200
rect 551400 687100 551499 687300
rect 551000 687000 551499 687100
rect 537839 686962 551200 687000
rect 551089 686800 551200 686962
rect 551400 686800 551499 687000
rect 551089 686700 551499 686800
rect 43070 686670 46240 686680
rect 43070 686600 43330 686670
rect 43400 686600 43500 686670
rect 43070 686490 43500 686600
rect 43070 686420 43330 686490
rect 43400 686420 43500 686490
rect 43750 686600 43840 686670
rect 43910 686600 44360 686670
rect 44430 686600 44880 686670
rect 44950 686600 45390 686670
rect 45460 686600 45560 686670
rect 43750 686490 45560 686600
rect 43750 686420 43840 686490
rect 43910 686420 44360 686490
rect 44430 686420 44880 686490
rect 44950 686420 45390 686490
rect 45460 686420 45560 686490
rect 45810 686600 45910 686670
rect 45980 686600 46240 686670
rect 45810 686490 46240 686600
rect 45810 686420 45910 686490
rect 45980 686420 46240 686490
rect 43070 686410 46240 686420
rect 551089 686500 551200 686700
rect 551400 686500 551499 686700
rect 551089 686400 551499 686500
rect 44520 686250 44790 686255
rect 44520 686000 44530 686250
rect 44780 686000 44790 686250
rect 551089 686200 551200 686400
rect 551400 686200 551499 686400
rect 551089 686192 551499 686200
rect 44520 685995 44790 686000
rect 538209 686100 551499 686192
rect 538209 686072 549800 686100
rect 538209 686062 540299 686072
rect 538209 685982 540119 686062
rect 540209 685992 540299 686062
rect 540389 686062 549800 686072
rect 540389 685992 542649 686062
rect 540209 685982 542649 685992
rect 542739 685982 542809 686062
rect 542899 685982 545119 686062
rect 545209 685982 545279 686062
rect 545369 685982 547569 686062
rect 547659 685982 547729 686062
rect 547819 685982 549800 686062
rect 538209 685900 549800 685982
rect 550000 686062 550100 686100
rect 550300 686062 550400 686100
rect 550000 685982 550069 686062
rect 550319 685982 550400 686062
rect 550000 685900 550100 685982
rect 550300 685900 550400 685982
rect 550600 685900 550800 686100
rect 551000 685900 551499 686100
rect 538209 685852 551499 685900
rect 42810 685825 46490 685830
rect 42800 685820 46500 685825
rect 42800 685750 42810 685820
rect 42880 685750 43330 685820
rect 43400 685750 43840 685820
rect 43910 685750 44360 685820
rect 44430 685750 44870 685820
rect 44940 685750 45390 685820
rect 45460 685750 45910 685820
rect 45980 685750 46420 685820
rect 46490 685750 46500 685820
rect 42800 685745 46500 685750
rect 42810 685645 46490 685745
rect 42800 685640 46500 685645
rect 42800 685570 42810 685640
rect 42880 685570 43330 685640
rect 43400 685570 43840 685640
rect 43910 685570 44360 685640
rect 44430 685570 44870 685640
rect 44940 685570 45390 685640
rect 45460 685570 45910 685640
rect 45980 685570 46420 685640
rect 46490 685570 46500 685640
rect 42800 685565 46500 685570
rect 42810 685560 46490 685565
rect 0 685300 38400 685400
rect 0 685242 36800 685300
rect -800 685100 36800 685242
rect 37000 685100 37200 685300
rect 37400 685100 37600 685300
rect 37800 685100 38000 685300
rect 38200 685100 38400 685300
rect 535739 685252 536089 685262
rect -800 684900 38400 685100
rect -800 684700 36800 684900
rect 37000 684700 37200 684900
rect 37400 684700 37600 684900
rect 37800 684700 38000 684900
rect 38200 684700 38400 684900
rect 42810 685150 46490 685160
rect 42810 685080 43070 685150
rect 43140 685080 43240 685150
rect 42810 684970 43240 685080
rect 42810 684900 43070 684970
rect 43140 684900 43240 684970
rect 43490 685080 43580 685150
rect 43650 685080 44100 685150
rect 44170 685080 44620 685150
rect 44690 685080 45130 685150
rect 45200 685080 45650 685150
rect 45720 685080 45820 685150
rect 43490 684970 45820 685080
rect 43490 684900 43580 684970
rect 43650 684900 44100 684970
rect 44170 684900 44620 684970
rect 44690 684900 45130 684970
rect 45200 684900 45650 684970
rect 45720 684900 45820 684970
rect 46070 685080 46160 685150
rect 46230 685080 46490 685150
rect 46070 684970 46490 685080
rect 46070 684900 46160 684970
rect 46230 684900 46490 684970
rect 535739 685122 535759 685252
rect 535849 685122 535969 685252
rect 536059 685122 536089 685252
rect 553059 685242 553319 685252
rect 553059 685152 553069 685242
rect 553139 685152 553229 685242
rect 553299 685152 553319 685242
rect 535739 684940 536089 685122
rect 542359 685132 542589 685142
rect 542359 685052 542379 685132
rect 542459 685052 542489 685132
rect 542569 685052 542589 685132
rect 542359 685042 542589 685052
rect 544769 685132 544999 685152
rect 544769 685052 544789 685132
rect 544869 685052 544899 685132
rect 544979 685052 544999 685132
rect 547229 685142 547459 685152
rect 547229 685062 547249 685142
rect 547329 685062 547359 685142
rect 547439 685062 547459 685142
rect 547229 685052 547459 685062
rect 544769 685042 544999 685052
rect 42810 684890 46490 684900
rect 515500 684912 540560 684940
rect 553059 684912 553319 685152
rect 515500 684800 554449 684912
rect -800 684500 38400 684700
rect -800 684300 36800 684500
rect 37000 684300 37200 684500
rect 37400 684300 37600 684500
rect 37800 684300 38000 684500
rect 38200 684300 38400 684500
rect 44520 684720 44790 684725
rect 44520 684470 44530 684720
rect 44780 684470 44790 684720
rect 44520 684465 44790 684470
rect 515500 684600 515700 684800
rect 515900 684600 516100 684800
rect 516300 684600 516500 684800
rect 516700 684600 516900 684800
rect 517100 684600 517300 684800
rect 517500 684600 517700 684800
rect 517900 684600 518100 684800
rect 518300 684600 518500 684800
rect 518700 684600 518900 684800
rect 519100 684600 519300 684800
rect 519500 684600 519700 684800
rect 519900 684600 520100 684800
rect 520300 684600 520500 684800
rect 520700 684772 554449 684800
rect 520700 684662 542279 684772
rect 542389 684662 543139 684772
rect 543249 684662 544349 684772
rect 544459 684662 545199 684772
rect 545309 684662 546769 684772
rect 546879 684662 547649 684772
rect 547759 684662 554449 684772
rect 520700 684600 554449 684662
rect 515500 684552 554449 684600
rect -800 684100 38400 684300
rect -800 683900 36800 684100
rect 37000 683900 37200 684100
rect 37400 683900 37600 684100
rect 37800 683900 38000 684100
rect 38200 683900 38400 684100
rect -800 683700 38400 683900
rect -800 683500 36800 683700
rect 37000 683500 37200 683700
rect 37400 683500 37600 683700
rect 37800 683500 38000 683700
rect 38200 683500 38400 683700
rect 515500 684400 540560 684552
rect 549399 684542 554449 684552
rect 515500 684200 515700 684400
rect 515900 684200 516100 684400
rect 516300 684200 516500 684400
rect 516700 684200 516900 684400
rect 517100 684200 517300 684400
rect 517500 684200 517700 684400
rect 517900 684200 518100 684400
rect 518300 684200 518500 684400
rect 518700 684200 518900 684400
rect 519100 684200 519300 684400
rect 519500 684200 519700 684400
rect 519900 684200 520100 684400
rect 520300 684200 520500 684400
rect 520700 684200 540560 684400
rect 543559 684392 543829 684402
rect 541069 684372 541339 684392
rect 541069 684292 541089 684372
rect 541169 684292 541239 684372
rect 541319 684292 541339 684372
rect 543559 684312 543579 684392
rect 543659 684312 543729 684392
rect 543809 684312 543829 684392
rect 543559 684292 543829 684312
rect 546039 684392 546309 684402
rect 546039 684312 546059 684392
rect 546139 684312 546199 684392
rect 546279 684312 546309 684392
rect 546039 684292 546309 684312
rect 541069 684262 541339 684292
rect 515500 684000 540560 684200
rect 515500 683800 515700 684000
rect 515900 683800 516100 684000
rect 516300 683800 516500 684000
rect 516700 683800 516900 684000
rect 517100 683800 517300 684000
rect 517500 683800 517700 684000
rect 517900 683800 518100 684000
rect 518300 683800 518500 684000
rect 518700 683800 518900 684000
rect 519100 683800 519300 684000
rect 519500 683800 519700 684000
rect 519900 683800 520100 684000
rect 520300 683800 520500 684000
rect 520700 683852 540560 684000
rect 549469 683852 549689 684542
rect 520700 683800 549689 683852
rect 515500 683652 549689 683800
rect 43800 683500 43810 683620
rect 43930 683600 45480 683620
rect 43930 683520 44350 683600
rect 44430 683520 44870 683600
rect 44950 683520 45390 683600
rect 45470 683520 45480 683600
rect 43930 683500 45480 683520
rect 515500 683600 541569 683652
rect -800 683300 38400 683500
rect -800 683100 36800 683300
rect 37000 683100 37200 683300
rect 37400 683100 37600 683300
rect 37800 683100 38000 683300
rect 38200 683100 38400 683300
rect 515500 683400 515700 683600
rect 515900 683400 516100 683600
rect 516300 683400 516500 683600
rect 516700 683400 516900 683600
rect 517100 683400 517300 683600
rect 517500 683400 517700 683600
rect 517900 683400 518100 683600
rect 518300 683400 518500 683600
rect 518700 683400 518900 683600
rect 519100 683400 519300 683600
rect 519500 683400 519700 683600
rect 519900 683400 520100 683600
rect 520300 683400 520500 683600
rect 520700 683562 541569 683600
rect 541679 683562 546479 683652
rect 546589 683562 549689 683652
rect 520700 683400 549689 683562
rect 515500 683392 549689 683400
rect 515500 683200 540560 683392
rect -800 682900 38400 683100
rect 42240 683120 47040 683140
rect 42240 683040 42260 683120
rect 42340 683040 42400 683120
rect 42480 683040 42540 683120
rect 42620 683040 44090 683120
rect 44170 683040 44610 683120
rect 44690 683040 45130 683120
rect 45210 683040 46660 683120
rect 46740 683040 46800 683120
rect 46880 683040 46940 683120
rect 47020 683040 47040 683120
rect 42240 683020 47040 683040
rect -800 682700 36800 682900
rect 37000 682700 37200 682900
rect 37400 682700 37600 682900
rect 37800 682700 38000 682900
rect 38200 682700 38400 682900
rect -800 682500 38400 682700
rect -800 682300 36800 682500
rect 37000 682300 37200 682500
rect 37400 682300 37600 682500
rect 37800 682300 38000 682500
rect 38200 682300 38400 682500
rect 515500 683000 515700 683200
rect 515900 683000 516100 683200
rect 516300 683000 516500 683200
rect 516700 683000 516900 683200
rect 517100 683000 517300 683200
rect 517500 683000 517700 683200
rect 517900 683000 518100 683200
rect 518300 683000 518500 683200
rect 518700 683000 518900 683200
rect 519100 683000 519300 683200
rect 519500 683000 519700 683200
rect 519900 683000 520100 683200
rect 520300 683000 520500 683200
rect 520700 683000 540560 683200
rect 515500 682800 540560 683000
rect 515500 682600 515700 682800
rect 515900 682600 516100 682800
rect 516300 682600 516500 682800
rect 516700 682600 516900 682800
rect 517100 682600 517300 682800
rect 517500 682600 517700 682800
rect 517900 682600 518100 682800
rect 518300 682600 518500 682800
rect 518700 682600 518900 682800
rect 519100 682600 519300 682800
rect 519500 682600 519700 682800
rect 519900 682600 520100 682800
rect 520300 682600 520500 682800
rect 520700 682672 540560 682800
rect 549469 682672 549689 683392
rect 520700 682600 549689 682672
rect 515500 682460 549689 682600
rect 515500 682400 515600 682460
rect 539629 682452 549689 682460
rect 539629 682352 541509 682452
rect 541629 682352 542729 682452
rect 542849 682352 543939 682452
rect 544059 682352 545159 682452
rect 545279 682442 547599 682452
rect 545279 682352 546389 682442
rect 539629 682342 546389 682352
rect 546509 682352 547599 682442
rect 547719 682352 549689 682452
rect 546509 682342 549689 682352
rect -800 682100 38400 682300
rect 45440 682200 62200 682320
rect 539629 682212 549689 682342
rect 561620 682984 582320 683140
rect 45440 682160 58000 682200
rect -800 681900 36800 682100
rect 37000 681900 37200 682100
rect 37400 681900 37600 682100
rect 37800 681900 38000 682100
rect 38200 681900 38400 682100
rect 43570 682140 58000 682160
rect 43570 682060 43630 682140
rect 43710 682060 43840 682140
rect 43920 682060 44350 682140
rect 44430 682060 44870 682140
rect 44950 682060 45390 682140
rect 45470 682060 45590 682140
rect 45670 682060 58000 682140
rect 43570 682040 58000 682060
rect 45440 682000 58000 682040
rect 58200 682000 58400 682200
rect 58600 682000 58800 682200
rect 59000 682000 59200 682200
rect 59400 682000 59600 682200
rect 59800 682000 60000 682200
rect 60200 682000 60400 682200
rect 60600 682000 60800 682200
rect 61000 682000 61200 682200
rect 61400 682000 61600 682200
rect 61800 682000 62200 682200
rect -800 681700 38400 681900
rect -800 681500 36800 681700
rect 37000 681500 37200 681700
rect 37400 681500 37600 681700
rect 37800 681500 38000 681700
rect 38200 681500 38400 681700
rect 43610 681920 43730 681940
rect 43610 681840 43630 681920
rect 43710 681840 43730 681920
rect 45440 681920 62200 682000
rect 561620 682200 584800 682984
rect 561620 682000 561700 682200
rect 561900 682000 562100 682200
rect 562300 682000 562500 682200
rect 562700 682000 562900 682200
rect 563100 682000 563300 682200
rect 563500 682000 584800 682200
rect 45440 681860 45590 681920
rect 43610 681780 43730 681840
rect 43610 681700 43630 681780
rect 43710 681700 43730 681780
rect 43610 681680 43730 681700
rect 45570 681840 45590 681860
rect 45670 681860 62200 681920
rect 45670 681840 45690 681860
rect 45570 681780 45690 681840
rect 45570 681700 45590 681780
rect 45670 681700 45690 681780
rect 45570 681680 45690 681700
rect -800 681300 38400 681500
rect -800 681100 36800 681300
rect 37000 681100 37200 681300
rect 37400 681100 37600 681300
rect 37800 681100 38000 681300
rect 38200 681100 38400 681300
rect -800 680900 38400 681100
rect -800 680700 36800 680900
rect 37000 680700 37200 680900
rect 37400 680700 37600 680900
rect 37800 680700 38000 680900
rect 38200 680700 38400 680900
rect 541344 681500 547804 681938
rect 561620 681800 584800 682000
rect 561620 681600 561700 681800
rect 561900 681600 562100 681800
rect 562300 681600 562500 681800
rect 562700 681600 562900 681800
rect 563100 681600 563300 681800
rect 563500 681600 584800 681800
rect 541344 681478 553100 681500
rect 541344 681318 541384 681478
rect 541544 681318 542444 681478
rect 542604 681318 543904 681478
rect 544064 681318 545124 681478
rect 545284 681318 546604 681478
rect 546764 681318 547604 681478
rect 547764 681400 553100 681478
rect 547764 681318 549800 681400
rect 541344 681200 549800 681318
rect 550000 681200 550200 681400
rect 550400 681200 550600 681400
rect 550800 681200 551000 681400
rect 551200 681200 551400 681400
rect 551600 681200 551800 681400
rect 552000 681200 552200 681400
rect 552400 681200 552600 681400
rect 552800 681200 553100 681400
rect 541344 681000 553100 681200
rect 541344 680898 549800 681000
rect 541344 680738 541384 680898
rect 541544 680738 542444 680898
rect 542604 680738 543904 680898
rect 544064 680738 545124 680898
rect 545284 680738 546604 680898
rect 546764 680738 547604 680898
rect 547764 680800 549800 680898
rect 550000 680800 550200 681000
rect 550400 680800 550600 681000
rect 550800 680800 551000 681000
rect 551200 680800 551400 681000
rect 551600 680800 551800 681000
rect 552000 680800 552200 681000
rect 552400 680800 552600 681000
rect 552800 680800 553100 681000
rect 547764 680738 553100 680800
rect 541344 680718 553100 680738
rect 547600 680700 553100 680718
rect 561620 681400 584800 681600
rect 561620 681200 561700 681400
rect 561900 681200 562100 681400
rect 562300 681200 562500 681400
rect 562700 681200 562900 681400
rect 563100 681200 563300 681400
rect 563500 681200 584800 681400
rect 561620 681000 584800 681200
rect 561620 680800 561700 681000
rect 561900 680800 562100 681000
rect 562300 680800 562500 681000
rect 562700 680800 562900 681000
rect 563100 680800 563300 681000
rect 563500 680800 584800 681000
rect -800 680500 38400 680700
rect 561620 680600 584800 680800
rect 44880 680530 45020 680535
rect -800 680300 36800 680500
rect 37000 680300 37200 680500
rect 37400 680300 37600 680500
rect 37800 680300 38000 680500
rect 38200 680300 38400 680500
rect 44260 680520 44400 680525
rect 44260 680400 44270 680520
rect 44390 680400 44400 680520
rect 44880 680410 44890 680530
rect 45010 680410 45020 680530
rect 44880 680405 45020 680410
rect 44260 680395 44400 680400
rect 561620 680400 561700 680600
rect 561900 680400 562100 680600
rect 562300 680400 562500 680600
rect 562700 680400 562900 680600
rect 563100 680400 563300 680600
rect 563500 680400 584800 680600
rect -800 680242 38400 680300
rect 0 680200 38400 680242
rect 561620 680200 584800 680400
rect 561620 680000 561700 680200
rect 561900 680000 562100 680200
rect 562300 680000 562500 680200
rect 562700 680000 562900 680200
rect 563100 680000 563300 680200
rect 563500 680000 584800 680200
rect 561620 679800 584800 680000
rect 44050 679630 45210 679650
rect 44050 679540 44070 679630
rect 44160 679540 44590 679630
rect 44680 679540 45100 679630
rect 45190 679540 45210 679630
rect 561620 679600 561700 679800
rect 561900 679600 562100 679800
rect 562300 679600 562500 679800
rect 562700 679600 562900 679800
rect 563100 679600 563300 679800
rect 563500 679600 584800 679800
rect 44050 679520 45210 679540
rect 511150 679558 541760 679560
rect 511150 679518 547914 679558
rect 511150 679368 543764 679518
rect 543984 679368 544284 679518
rect 544504 679368 544704 679518
rect 544924 679368 545254 679518
rect 545474 679368 547914 679518
rect 44570 679250 44680 679255
rect 44570 679160 44580 679250
rect 44670 679160 44680 679250
rect 44570 679155 44680 679160
rect 511150 679200 547914 679368
rect 511150 679000 515900 679200
rect 516100 679000 516300 679200
rect 516500 679000 516700 679200
rect 516900 679000 517100 679200
rect 517300 679000 517500 679200
rect 517700 679000 517900 679200
rect 518100 679000 518300 679200
rect 518500 679000 518700 679200
rect 518900 679000 519100 679200
rect 519300 679000 519500 679200
rect 519700 679000 519900 679200
rect 520100 679000 520300 679200
rect 520500 679000 520700 679200
rect 520900 679000 547914 679200
rect 511150 678968 547914 679000
rect 511150 678958 543524 678968
rect 511150 678828 541404 678958
rect 541584 678828 542544 678958
rect 542724 678838 543524 678958
rect 543704 678838 544294 678968
rect 544474 678838 544734 678968
rect 544914 678958 546524 678968
rect 544914 678838 545454 678958
rect 542724 678828 545454 678838
rect 545634 678838 546524 678958
rect 546704 678838 547524 678968
rect 547704 678838 547914 678968
rect 545634 678828 547914 678838
rect 511150 678800 547914 678828
rect 44820 678720 44970 678725
rect 44820 678700 44830 678720
rect 43820 678690 44830 678700
rect 43820 678630 43830 678690
rect 43890 678630 44350 678690
rect 44410 678630 44830 678690
rect 43820 678620 44830 678630
rect 44820 678610 44830 678620
rect 44960 678700 44970 678720
rect 44960 678690 45450 678700
rect 44960 678630 45380 678690
rect 45440 678630 45450 678690
rect 44960 678620 45450 678630
rect 44960 678610 44970 678620
rect 44820 678605 44970 678610
rect 511150 678600 515900 678800
rect 516100 678600 516300 678800
rect 516500 678600 516700 678800
rect 516900 678600 517100 678800
rect 517300 678600 517500 678800
rect 517700 678600 517900 678800
rect 518100 678600 518300 678800
rect 518500 678600 518700 678800
rect 518900 678600 519100 678800
rect 519300 678600 519500 678800
rect 519700 678600 519900 678800
rect 520100 678600 520300 678800
rect 520500 678600 520700 678800
rect 520900 678798 547914 678800
rect 520900 678600 541760 678798
rect 511150 678400 541760 678600
rect 43840 678280 45430 678290
rect 43840 678220 44090 678280
rect 44150 678220 44610 678280
rect 44670 678220 45120 678280
rect 45180 678220 45430 678280
rect 43840 678210 45430 678220
rect 511150 678200 515900 678400
rect 516100 678200 516300 678400
rect 516500 678200 516700 678400
rect 516900 678200 517100 678400
rect 517300 678200 517500 678400
rect 517700 678200 517900 678400
rect 518100 678200 518300 678400
rect 518500 678200 518700 678400
rect 518900 678200 519100 678400
rect 519300 678200 519500 678400
rect 519700 678200 519900 678400
rect 520100 678200 520300 678400
rect 520500 678200 520700 678400
rect 520900 678200 541760 678400
rect 511150 678000 541760 678200
rect 44570 677810 44680 677815
rect 44570 677720 44580 677810
rect 44670 677720 44680 677810
rect 44570 677715 44680 677720
rect 511150 677800 515900 678000
rect 516100 677800 516300 678000
rect 516500 677800 516700 678000
rect 516900 677800 517100 678000
rect 517300 677800 517500 678000
rect 517700 677800 517900 678000
rect 518100 677800 518300 678000
rect 518500 677800 518700 678000
rect 518900 677800 519100 678000
rect 519300 677800 519500 678000
rect 519700 677800 519900 678000
rect 520100 677800 520300 678000
rect 520500 677800 520700 678000
rect 520900 677800 541760 678000
rect 511150 677600 541760 677800
rect 511150 677400 515900 677600
rect 516100 677400 516300 677600
rect 516500 677400 516700 677600
rect 516900 677400 517100 677600
rect 517300 677400 517500 677600
rect 517700 677400 517900 677600
rect 518100 677400 518300 677600
rect 518500 677400 518700 677600
rect 518900 677400 519100 677600
rect 519300 677400 519500 677600
rect 519700 677400 519900 677600
rect 520100 677400 520300 677600
rect 520500 677400 520700 677600
rect 520900 677400 541760 677600
rect 511150 677200 541760 677400
rect 511150 677000 515900 677200
rect 516100 677000 516300 677200
rect 516500 677000 516700 677200
rect 516900 677000 517100 677200
rect 517300 677000 517500 677200
rect 517700 677000 517900 677200
rect 518100 677000 518300 677200
rect 518500 677000 518700 677200
rect 518900 677000 519100 677200
rect 519300 677000 519500 677200
rect 519700 677000 519900 677200
rect 520100 677000 520300 677200
rect 520500 677000 520700 677200
rect 520900 677058 541760 677200
rect 520900 677000 541364 677058
rect 41190 676980 41450 676985
rect 41190 676740 41200 676980
rect 41440 676740 41450 676980
rect 41190 676735 41450 676740
rect 47890 676980 48150 676985
rect 47890 676740 47900 676980
rect 48140 676740 48150 676980
rect 47890 676735 48150 676740
rect 511150 676938 541364 677000
rect 541484 676938 541760 677058
rect 511150 676800 541760 676938
rect 511150 676600 515900 676800
rect 516100 676600 516300 676800
rect 516500 676600 516700 676800
rect 516900 676600 517100 676800
rect 517300 676600 517500 676800
rect 517700 676600 517900 676800
rect 518100 676600 518300 676800
rect 518500 676600 518700 676800
rect 518900 676600 519100 676800
rect 519300 676600 519500 676800
rect 519700 676600 519900 676800
rect 520100 676600 520300 676800
rect 520500 676600 520700 676800
rect 520900 676600 541760 676800
rect 511150 676460 541760 676600
rect 547594 677058 547914 678798
rect 561620 679400 584800 679600
rect 561620 679200 561700 679400
rect 561900 679200 562100 679400
rect 562300 679200 562500 679400
rect 562700 679200 562900 679400
rect 563100 679200 563300 679400
rect 563500 679200 584800 679400
rect 561620 679000 584800 679200
rect 561620 678800 561700 679000
rect 561900 678800 562100 679000
rect 562300 678800 562500 679000
rect 562700 678800 562900 679000
rect 563100 678800 563300 679000
rect 563500 678800 584800 679000
rect 561620 678600 584800 678800
rect 561620 678400 561700 678600
rect 561900 678400 562100 678600
rect 562300 678400 562500 678600
rect 562700 678400 562900 678600
rect 563100 678400 563300 678600
rect 563500 678400 584800 678600
rect 561620 677984 584800 678400
rect 561620 677940 582320 677984
rect 547594 676938 547734 677058
rect 547854 676938 547914 677058
rect 41190 675260 41450 675265
rect 41190 675020 41200 675260
rect 41440 675020 41450 675260
rect 41190 675015 41450 675020
rect 47890 675260 48150 675265
rect 47890 675020 47900 675260
rect 48140 675020 48150 675260
rect 47890 675015 48150 675020
rect 41190 673540 41450 673545
rect 41190 673300 41200 673540
rect 41440 673300 41450 673540
rect 41190 673295 41450 673300
rect 47890 673540 48150 673545
rect 47890 673300 47900 673540
rect 48140 673300 48150 673540
rect 47890 673295 48150 673300
rect 41190 672060 41450 672065
rect 41190 671820 41200 672060
rect 41440 671820 41450 672060
rect 41190 671815 41450 671820
rect 47890 672060 48150 672065
rect 47890 671820 47900 672060
rect 48140 671820 48150 672060
rect 47890 671815 48150 671820
rect 41190 670340 41450 670345
rect 41190 670100 41200 670340
rect 41440 670100 41450 670340
rect 41190 670095 41450 670100
rect 47890 670340 48150 670345
rect 47890 670100 47900 670340
rect 48140 670100 48150 670340
rect 47890 670095 48150 670100
rect 41190 668740 41450 668745
rect 41190 668500 41200 668740
rect 41440 668500 41450 668740
rect 41190 668495 41450 668500
rect 47890 668740 48150 668745
rect 47890 668500 47900 668740
rect 48140 668500 48150 668740
rect 47890 668495 48150 668500
rect 41190 667020 41450 667025
rect 41190 666780 41200 667020
rect 41440 666780 41450 667020
rect 41190 666775 41450 666780
rect 47890 667020 48150 667025
rect 47890 666780 47900 667020
rect 48140 666780 48150 667020
rect 47890 666775 48150 666780
rect 41190 665420 41450 665425
rect 41190 665180 41200 665420
rect 41440 665180 41450 665420
rect 41190 665175 41450 665180
rect 47890 665420 48150 665425
rect 47890 665180 47900 665420
rect 48140 665180 48150 665420
rect 47890 665175 48150 665180
rect 41190 663700 41450 663705
rect 41190 663460 41200 663700
rect 41440 663460 41450 663700
rect 41190 663455 41450 663460
rect 47890 663700 48150 663705
rect 47890 663460 47900 663700
rect 48140 663460 48150 663700
rect 47890 663455 48150 663460
rect 32790 663300 33110 663305
rect 32790 663000 32800 663300
rect 33100 663000 33110 663300
rect 32790 662995 33110 663000
rect 33290 663300 33610 663305
rect 33290 663000 33300 663300
rect 33600 663000 33610 663300
rect 33290 662995 33610 663000
rect 33790 663300 34110 663305
rect 33790 663000 33800 663300
rect 34100 663000 34110 663300
rect 33790 662995 34110 663000
rect 34290 663300 34610 663305
rect 34290 663000 34300 663300
rect 34600 663000 34610 663300
rect 34290 662995 34610 663000
rect 34790 663300 35110 663305
rect 34790 663000 34800 663300
rect 35100 663000 35110 663300
rect 34790 662995 35110 663000
rect 35290 663300 35610 663305
rect 35290 663000 35300 663300
rect 35600 663000 35610 663300
rect 35290 662995 35610 663000
rect 35790 663300 36110 663305
rect 35790 663000 35800 663300
rect 36100 663000 36110 663300
rect 35790 662995 36110 663000
rect 36290 663300 36610 663305
rect 36290 663000 36300 663300
rect 36600 663000 36610 663300
rect 36290 662995 36610 663000
rect 36790 663300 37110 663305
rect 36790 663000 36800 663300
rect 37100 663000 37110 663300
rect 36790 662995 37110 663000
rect 37290 663300 37610 663305
rect 37290 663000 37300 663300
rect 37600 663000 37610 663300
rect 37290 662995 37610 663000
rect 37790 663300 38110 663305
rect 37790 663000 37800 663300
rect 38100 663000 38110 663300
rect 37790 662995 38110 663000
rect 38290 663300 38610 663305
rect 38290 663000 38300 663300
rect 38600 663000 38610 663300
rect 38290 662995 38610 663000
rect 38790 663300 39110 663305
rect 38790 663000 38800 663300
rect 39100 663000 39110 663300
rect 38790 662995 39110 663000
rect 39290 663300 39610 663305
rect 39290 663000 39300 663300
rect 39600 663000 39610 663300
rect 39290 662995 39610 663000
rect 39790 663300 40110 663305
rect 39790 663000 39800 663300
rect 40100 663000 40110 663300
rect 39790 662995 40110 663000
rect 40290 663300 40610 663305
rect 40290 663000 40300 663300
rect 40600 663000 40610 663300
rect 40290 662995 40610 663000
rect 0 648642 4000 648800
rect -800 648600 4000 648642
rect -800 648300 2500 648600
rect 2800 648300 3000 648600
rect 3300 648300 3500 648600
rect 3800 648300 4000 648600
rect -800 648100 4000 648300
rect -800 647800 2500 648100
rect 2800 647800 3000 648100
rect 3300 647800 3500 648100
rect 3800 647800 4000 648100
rect -800 647600 4000 647800
rect -800 647300 2500 647600
rect 2800 647300 3000 647600
rect 3300 647300 3500 647600
rect 3800 647300 4000 647600
rect -800 647100 4000 647300
rect -800 646800 2500 647100
rect 2800 646800 3000 647100
rect 3300 646800 3500 647100
rect 3800 646800 4000 647100
rect -800 646600 4000 646800
rect -800 646300 2500 646600
rect 2800 646300 3000 646600
rect 3300 646300 3500 646600
rect 3800 646300 4000 646600
rect -800 646100 4000 646300
rect -800 645800 2500 646100
rect 2800 645800 3000 646100
rect 3300 645800 3500 646100
rect 3800 645800 4000 646100
rect -800 645600 4000 645800
rect -800 645300 2500 645600
rect 2800 645300 3000 645600
rect 3300 645300 3500 645600
rect 3800 645300 4000 645600
rect -800 645100 4000 645300
rect -800 644800 2500 645100
rect 2800 644800 3000 645100
rect 3300 644800 3500 645100
rect 3800 644800 4000 645100
rect -800 644600 4000 644800
rect -800 644300 2500 644600
rect 2800 644300 3000 644600
rect 3300 644300 3500 644600
rect 3800 644300 4000 644600
rect -800 644100 4000 644300
rect -800 643842 2500 644100
rect 0 643800 2500 643842
rect 2800 643800 3000 644100
rect 3300 643800 3500 644100
rect 3800 643800 4000 644100
rect 0 643600 4000 643800
rect 0 643300 2500 643600
rect 2800 643300 3000 643600
rect 3300 643300 3500 643600
rect 3800 643300 4000 643600
rect 0 643100 4000 643300
rect 0 642800 2500 643100
rect 2800 642800 3000 643100
rect 3300 642800 3500 643100
rect 3800 642800 4000 643100
rect 0 642600 4000 642800
rect 0 642300 2500 642600
rect 2800 642300 3000 642600
rect 3300 642300 3500 642600
rect 3800 642300 4000 642600
rect 0 642100 4000 642300
rect 0 641800 2500 642100
rect 2800 641800 3000 642100
rect 3300 641800 3500 642100
rect 3800 641800 4000 642100
rect 0 641600 4000 641800
rect 0 641300 2500 641600
rect 2800 641300 3000 641600
rect 3300 641300 3500 641600
rect 3800 641300 4000 641600
rect 0 641100 4000 641300
rect 0 640800 2500 641100
rect 2800 640800 3000 641100
rect 3300 640800 3500 641100
rect 3800 640800 4000 641100
rect 0 640600 4000 640800
rect 0 640300 2500 640600
rect 2800 640300 3000 640600
rect 3300 640300 3500 640600
rect 3800 640300 4000 640600
rect 0 640100 4000 640300
rect 0 639800 2500 640100
rect 2800 639800 3000 640100
rect 3300 639800 3500 640100
rect 3800 639800 4000 640100
rect 0 639600 4000 639800
rect 0 639300 2500 639600
rect 2800 639300 3000 639600
rect 3300 639300 3500 639600
rect 3800 639300 4000 639600
rect 0 639100 4000 639300
rect 0 638800 2500 639100
rect 2800 638800 3000 639100
rect 3300 638800 3500 639100
rect 3800 638800 4000 639100
rect 0 638642 4000 638800
rect -800 638600 4000 638642
rect -800 638300 2500 638600
rect 2800 638300 3000 638600
rect 3300 638300 3500 638600
rect 3800 638300 4000 638600
rect -800 638100 4000 638300
rect -800 637800 2500 638100
rect 2800 637800 3000 638100
rect 3300 637800 3500 638100
rect 3800 637800 4000 638100
rect -800 637600 4000 637800
rect -800 637300 2500 637600
rect 2800 637300 3000 637600
rect 3300 637300 3500 637600
rect 3800 637300 4000 637600
rect -800 637100 4000 637300
rect -800 636800 2500 637100
rect 2800 636800 3000 637100
rect 3300 636800 3500 637100
rect 3800 636800 4000 637100
rect -800 636600 4000 636800
rect -800 636300 2500 636600
rect 2800 636300 3000 636600
rect 3300 636300 3500 636600
rect 3800 636300 4000 636600
rect -800 636100 4000 636300
rect -800 635800 2500 636100
rect 2800 635800 3000 636100
rect 3300 635800 3500 636100
rect 3800 635800 4000 636100
rect -800 635600 4000 635800
rect -800 635300 2500 635600
rect 2800 635300 3000 635600
rect 3300 635300 3500 635600
rect 3800 635300 4000 635600
rect -800 635100 4000 635300
rect -800 634800 2500 635100
rect 2800 634800 3000 635100
rect 3300 634800 3500 635100
rect 3800 634800 4000 635100
rect -800 634600 4000 634800
rect -800 634300 2500 634600
rect 2800 634300 3000 634600
rect 3300 634300 3500 634600
rect 3800 634300 4000 634600
rect -800 633842 4000 634300
rect 0 633800 4000 633842
rect 511150 572960 521284 676460
rect 541294 674058 541614 676460
rect 541294 673938 541364 674058
rect 541484 673938 541614 674058
rect 541294 671058 541614 673938
rect 541294 670938 541364 671058
rect 541484 670938 541614 671058
rect 541294 668058 541614 670938
rect 541294 667938 541364 668058
rect 541484 667938 541614 668058
rect 541294 665058 541614 667938
rect 541294 664938 541364 665058
rect 541484 664938 541614 665058
rect 541294 663758 541614 664938
rect 547594 674058 547914 676938
rect 547594 673938 547734 674058
rect 547854 673938 547914 674058
rect 547594 671058 547914 673938
rect 547594 670938 547734 671058
rect 547854 670938 547914 671058
rect 547594 668058 547914 670938
rect 547594 667938 547734 668058
rect 547854 667938 547914 668058
rect 547594 665058 547914 667938
rect 547594 664938 547734 665058
rect 547854 664938 547914 665058
rect 547594 663758 547914 664938
rect 541294 663738 547914 663758
rect 541294 663728 546294 663738
rect 541294 663318 541744 663728
rect 542914 663318 543254 663728
rect 544424 663318 544774 663728
rect 545944 663328 546294 663728
rect 547464 663328 547914 663738
rect 545944 663318 547914 663328
rect 541294 663278 547914 663318
rect 549700 644600 584000 644700
rect 549700 644400 550000 644600
rect 550200 644400 550400 644600
rect 550600 644400 550800 644600
rect 551000 644400 551200 644600
rect 551400 644400 551600 644600
rect 551800 644400 552000 644600
rect 552200 644400 552400 644600
rect 552600 644400 552800 644600
rect 553000 644584 584000 644600
rect 553000 644400 584800 644584
rect 549700 644200 584800 644400
rect 549700 644000 550000 644200
rect 550200 644000 550400 644200
rect 550600 644000 550800 644200
rect 551000 644000 551200 644200
rect 551400 644000 551600 644200
rect 551800 644000 552000 644200
rect 552200 644000 552400 644200
rect 552600 644000 552800 644200
rect 553000 644000 584800 644200
rect 549700 643800 584800 644000
rect 549700 643600 550000 643800
rect 550200 643600 550400 643800
rect 550600 643600 550800 643800
rect 551000 643600 551200 643800
rect 551400 643600 551600 643800
rect 551800 643600 552000 643800
rect 552200 643600 552400 643800
rect 552600 643600 552800 643800
rect 553000 643600 584800 643800
rect 549700 643400 584800 643600
rect 549700 643200 550000 643400
rect 550200 643200 550400 643400
rect 550600 643200 550800 643400
rect 551000 643200 551200 643400
rect 551400 643200 551600 643400
rect 551800 643200 552000 643400
rect 552200 643200 552400 643400
rect 552600 643200 552800 643400
rect 553000 643200 584800 643400
rect 549700 643000 584800 643200
rect 549700 642800 550000 643000
rect 550200 642800 550400 643000
rect 550600 642800 550800 643000
rect 551000 642800 551200 643000
rect 551400 642800 551600 643000
rect 551800 642800 552000 643000
rect 552200 642800 552400 643000
rect 552600 642800 552800 643000
rect 553000 642800 584800 643000
rect 549700 642600 584800 642800
rect 549700 642400 550000 642600
rect 550200 642400 550400 642600
rect 550600 642400 550800 642600
rect 551000 642400 551200 642600
rect 551400 642400 551600 642600
rect 551800 642400 552000 642600
rect 552200 642400 552400 642600
rect 552600 642400 552800 642600
rect 553000 642400 584800 642600
rect 549700 642200 584800 642400
rect 549700 642000 550000 642200
rect 550200 642000 550400 642200
rect 550600 642000 550800 642200
rect 551000 642000 551200 642200
rect 551400 642000 551600 642200
rect 551800 642000 552000 642200
rect 552200 642000 552400 642200
rect 552600 642000 552800 642200
rect 553000 642000 584800 642200
rect 549700 641800 584800 642000
rect 549700 641600 550000 641800
rect 550200 641600 550400 641800
rect 550600 641600 550800 641800
rect 551000 641600 551200 641800
rect 551400 641600 551600 641800
rect 551800 641600 552000 641800
rect 552200 641600 552400 641800
rect 552600 641600 552800 641800
rect 553000 641600 584800 641800
rect 549700 641400 584800 641600
rect 549700 641200 550000 641400
rect 550200 641200 550400 641400
rect 550600 641200 550800 641400
rect 551000 641200 551200 641400
rect 551400 641200 551600 641400
rect 551800 641200 552000 641400
rect 552200 641200 552400 641400
rect 552600 641200 552800 641400
rect 553000 641200 584800 641400
rect 549700 641000 584800 641200
rect 549700 640800 550000 641000
rect 550200 640800 550400 641000
rect 550600 640800 550800 641000
rect 551000 640800 551200 641000
rect 551400 640800 551600 641000
rect 551800 640800 552000 641000
rect 552200 640800 552400 641000
rect 552600 640800 552800 641000
rect 553000 640800 584800 641000
rect 549700 640600 584800 640800
rect 549700 640400 550000 640600
rect 550200 640400 550400 640600
rect 550600 640400 550800 640600
rect 551000 640400 551200 640600
rect 551400 640400 551600 640600
rect 551800 640400 552000 640600
rect 552200 640400 552400 640600
rect 552600 640400 552800 640600
rect 553000 640400 584800 640600
rect 549700 640200 584800 640400
rect 549700 640000 550000 640200
rect 550200 640000 550400 640200
rect 550600 640000 550800 640200
rect 551000 640000 551200 640200
rect 551400 640000 551600 640200
rect 551800 640000 552000 640200
rect 552200 640000 552400 640200
rect 552600 640000 552800 640200
rect 553000 640000 584800 640200
rect 549700 639800 584800 640000
rect 549700 639600 550000 639800
rect 550200 639600 550400 639800
rect 550600 639600 550800 639800
rect 551000 639600 551200 639800
rect 551400 639600 551600 639800
rect 551800 639600 552000 639800
rect 552200 639600 552400 639800
rect 552600 639600 552800 639800
rect 553000 639784 584800 639800
rect 553000 639600 582600 639784
rect 549700 639400 582600 639600
rect 549700 639200 550000 639400
rect 550200 639200 550400 639400
rect 550600 639200 550800 639400
rect 551000 639200 551200 639400
rect 551400 639200 551600 639400
rect 551800 639200 552000 639400
rect 552200 639200 552400 639400
rect 552600 639200 552800 639400
rect 553000 639200 582600 639400
rect 549700 639000 582600 639200
rect 549700 638800 550000 639000
rect 550200 638800 550400 639000
rect 550600 638800 550800 639000
rect 551000 638800 551200 639000
rect 551400 638800 551600 639000
rect 551800 638800 552000 639000
rect 552200 638800 552400 639000
rect 552600 638800 552800 639000
rect 553000 638800 582600 639000
rect 549700 638600 582600 638800
rect 549700 638400 550000 638600
rect 550200 638400 550400 638600
rect 550600 638400 550800 638600
rect 551000 638400 551200 638600
rect 551400 638400 551600 638600
rect 551800 638400 552000 638600
rect 552200 638400 552400 638600
rect 552600 638400 552800 638600
rect 553000 638400 582600 638600
rect 549700 638200 582600 638400
rect 549700 638000 550000 638200
rect 550200 638000 550400 638200
rect 550600 638000 550800 638200
rect 551000 638000 551200 638200
rect 551400 638000 551600 638200
rect 551800 638000 552000 638200
rect 552200 638000 552400 638200
rect 552600 638000 552800 638200
rect 553000 638000 582600 638200
rect 549700 637800 582600 638000
rect 549700 637600 550000 637800
rect 550200 637600 550400 637800
rect 550600 637600 550800 637800
rect 551000 637600 551200 637800
rect 551400 637600 551600 637800
rect 551800 637600 552000 637800
rect 552200 637600 552400 637800
rect 552600 637600 552800 637800
rect 553000 637600 582600 637800
rect 549700 637400 582600 637600
rect 549700 637200 550000 637400
rect 550200 637200 550400 637400
rect 550600 637200 550800 637400
rect 551000 637200 551200 637400
rect 551400 637200 551600 637400
rect 551800 637200 552000 637400
rect 552200 637200 552400 637400
rect 552600 637200 552800 637400
rect 553000 637200 582600 637400
rect 549700 637000 582600 637200
rect 549700 636800 550000 637000
rect 550200 636800 550400 637000
rect 550600 636800 550800 637000
rect 551000 636800 551200 637000
rect 551400 636800 551600 637000
rect 551800 636800 552000 637000
rect 552200 636800 552400 637000
rect 552600 636800 552800 637000
rect 553000 636800 582600 637000
rect 549700 636600 582600 636800
rect 549700 636400 550000 636600
rect 550200 636400 550400 636600
rect 550600 636400 550800 636600
rect 551000 636400 551200 636600
rect 551400 636400 551600 636600
rect 551800 636400 552000 636600
rect 552200 636400 552400 636600
rect 552600 636400 552800 636600
rect 553000 636400 582600 636600
rect 549700 636200 582600 636400
rect 549700 636000 550000 636200
rect 550200 636000 550400 636200
rect 550600 636000 550800 636200
rect 551000 636000 551200 636200
rect 551400 636000 551600 636200
rect 551800 636000 552000 636200
rect 552200 636000 552400 636200
rect 552600 636000 552800 636200
rect 553000 636000 582600 636200
rect 549700 635800 582600 636000
rect 549700 635600 550000 635800
rect 550200 635600 550400 635800
rect 550600 635600 550800 635800
rect 551000 635600 551200 635800
rect 551400 635600 551600 635800
rect 551800 635600 552000 635800
rect 552200 635600 552400 635800
rect 552600 635600 552800 635800
rect 553000 635600 582600 635800
rect 549700 635400 582600 635600
rect 549700 635200 550000 635400
rect 550200 635200 550400 635400
rect 550600 635200 550800 635400
rect 551000 635200 551200 635400
rect 551400 635200 551600 635400
rect 551800 635200 552000 635400
rect 552200 635200 552400 635400
rect 552600 635200 552800 635400
rect 553000 635200 582600 635400
rect 549700 635000 582600 635200
rect 549700 634800 550000 635000
rect 550200 634800 550400 635000
rect 550600 634800 550800 635000
rect 551000 634800 551200 635000
rect 551400 634800 551600 635000
rect 551800 634800 552000 635000
rect 552200 634800 552400 635000
rect 552600 634800 552800 635000
rect 553000 634800 582600 635000
rect 549700 634600 582600 634800
rect 549700 634400 550000 634600
rect 550200 634400 550400 634600
rect 550600 634400 550800 634600
rect 551000 634400 551200 634600
rect 551400 634400 551600 634600
rect 551800 634400 552000 634600
rect 552200 634400 552400 634600
rect 552600 634400 552800 634600
rect 553000 634584 582600 634600
rect 553000 634400 584800 634584
rect 549700 634200 584800 634400
rect 549700 634000 550000 634200
rect 550200 634000 550400 634200
rect 550600 634000 550800 634200
rect 551000 634000 551200 634200
rect 551400 634000 551600 634200
rect 551800 634000 552000 634200
rect 552200 634000 552400 634200
rect 552600 634000 552800 634200
rect 553000 634000 584800 634200
rect 549700 633800 584800 634000
rect 549700 633600 550000 633800
rect 550200 633600 550400 633800
rect 550600 633600 550800 633800
rect 551000 633600 551200 633800
rect 551400 633600 551600 633800
rect 551800 633600 552000 633800
rect 552200 633600 552400 633800
rect 552600 633600 552800 633800
rect 553000 633600 584800 633800
rect 549700 633400 584800 633600
rect 549700 633200 550000 633400
rect 550200 633200 550400 633400
rect 550600 633200 550800 633400
rect 551000 633200 551200 633400
rect 551400 633200 551600 633400
rect 551800 633200 552000 633400
rect 552200 633200 552400 633400
rect 552600 633200 552800 633400
rect 553000 633200 584800 633400
rect 549700 633000 584800 633200
rect 549700 632800 550000 633000
rect 550200 632800 550400 633000
rect 550600 632800 550800 633000
rect 551000 632800 551200 633000
rect 551400 632800 551600 633000
rect 551800 632800 552000 633000
rect 552200 632800 552400 633000
rect 552600 632800 552800 633000
rect 553000 632800 584800 633000
rect 549700 632600 584800 632800
rect 549700 632400 550000 632600
rect 550200 632400 550400 632600
rect 550600 632400 550800 632600
rect 551000 632400 551200 632600
rect 551400 632400 551600 632600
rect 551800 632400 552000 632600
rect 552200 632400 552400 632600
rect 552600 632400 552800 632600
rect 553000 632400 584800 632600
rect 549700 632200 584800 632400
rect 549700 632000 550000 632200
rect 550200 632000 550400 632200
rect 550600 632000 550800 632200
rect 551000 632000 551200 632200
rect 551400 632000 551600 632200
rect 551800 632000 552000 632200
rect 552200 632000 552400 632200
rect 552600 632000 552800 632200
rect 553000 632000 584800 632200
rect 549700 631800 584800 632000
rect 549700 631600 550000 631800
rect 550200 631600 550400 631800
rect 550600 631600 550800 631800
rect 551000 631600 551200 631800
rect 551400 631600 551600 631800
rect 551800 631600 552000 631800
rect 552200 631600 552400 631800
rect 552600 631600 552800 631800
rect 553000 631600 584800 631800
rect 549700 631400 584800 631600
rect 549700 631200 550000 631400
rect 550200 631200 550400 631400
rect 550600 631200 550800 631400
rect 551000 631200 551200 631400
rect 551400 631200 551600 631400
rect 551800 631200 552000 631400
rect 552200 631200 552400 631400
rect 552600 631200 552800 631400
rect 553000 631200 584800 631400
rect 549700 631000 584800 631200
rect 549700 630800 550000 631000
rect 550200 630800 550400 631000
rect 550600 630800 550800 631000
rect 551000 630800 551200 631000
rect 551400 630800 551600 631000
rect 551800 630800 552000 631000
rect 552200 630800 552400 631000
rect 552600 630800 552800 631000
rect 553000 630800 584800 631000
rect 549700 630700 584800 630800
rect 549700 630500 550000 630700
rect 550200 630500 550400 630700
rect 550600 630500 550800 630700
rect 551000 630500 551200 630700
rect 551400 630500 551600 630700
rect 551800 630500 552000 630700
rect 552200 630500 552400 630700
rect 552600 630500 552800 630700
rect 553000 630500 584800 630700
rect 549700 630400 584800 630500
rect 549700 630200 550000 630400
rect 550200 630200 550400 630400
rect 550600 630200 550800 630400
rect 551000 630200 551200 630400
rect 551400 630200 551600 630400
rect 551800 630200 552000 630400
rect 552200 630200 552400 630400
rect 552600 630200 552800 630400
rect 553000 630200 584800 630400
rect 549700 630000 584800 630200
rect 549700 629800 550000 630000
rect 550200 629800 550400 630000
rect 550600 629800 550800 630000
rect 551000 629800 551200 630000
rect 551400 629800 551600 630000
rect 551800 629800 552000 630000
rect 552200 629800 552400 630000
rect 552600 629800 552800 630000
rect 553000 629800 584800 630000
rect 549700 629784 584800 629800
rect 549700 629700 582600 629784
rect 549700 629660 580096 629700
rect 568260 629656 580096 629660
rect 0 564242 40800 564300
rect -800 564100 40800 564242
rect -800 563900 32800 564100
rect 33000 563900 33200 564100
rect 33400 563900 33600 564100
rect 33800 563900 34000 564100
rect 34200 563900 34400 564100
rect 34600 563900 34800 564100
rect 35000 563900 35200 564100
rect 35400 563900 35600 564100
rect 35800 563900 36000 564100
rect 36200 563900 36400 564100
rect 36600 563900 36800 564100
rect 37000 563900 37200 564100
rect 37400 563900 37600 564100
rect 37800 563900 38000 564100
rect 38200 563900 38400 564100
rect 38600 563900 38800 564100
rect 39000 563900 39200 564100
rect 39400 563900 39600 564100
rect 39800 563900 40000 564100
rect 40200 563900 40400 564100
rect 40600 563900 40800 564100
rect -800 563700 40800 563900
rect -800 563500 32800 563700
rect 33000 563500 33200 563700
rect 33400 563500 33600 563700
rect 33800 563500 34000 563700
rect 34200 563500 34400 563700
rect 34600 563500 34800 563700
rect 35000 563500 35200 563700
rect 35400 563500 35600 563700
rect 35800 563500 36000 563700
rect 36200 563500 36400 563700
rect 36600 563500 36800 563700
rect 37000 563500 37200 563700
rect 37400 563500 37600 563700
rect 37800 563500 38000 563700
rect 38200 563500 38400 563700
rect 38600 563500 38800 563700
rect 39000 563500 39200 563700
rect 39400 563500 39600 563700
rect 39800 563500 40000 563700
rect 40200 563500 40400 563700
rect 40600 563500 40800 563700
rect -800 563300 40800 563500
rect -800 563100 32800 563300
rect 33000 563100 33200 563300
rect 33400 563100 33600 563300
rect 33800 563100 34000 563300
rect 34200 563100 34400 563300
rect 34600 563100 34800 563300
rect 35000 563100 35200 563300
rect 35400 563100 35600 563300
rect 35800 563100 36000 563300
rect 36200 563100 36400 563300
rect 36600 563100 36800 563300
rect 37000 563100 37200 563300
rect 37400 563100 37600 563300
rect 37800 563100 38000 563300
rect 38200 563100 38400 563300
rect 38600 563100 38800 563300
rect 39000 563100 39200 563300
rect 39400 563100 39600 563300
rect 39800 563100 40000 563300
rect 40200 563100 40400 563300
rect 40600 563124 40800 563300
rect 511150 563124 521280 572960
rect 40600 563100 521280 563124
rect -800 562900 521280 563100
rect -800 562700 32800 562900
rect 33000 562700 33200 562900
rect 33400 562700 33600 562900
rect 33800 562700 34000 562900
rect 34200 562700 34400 562900
rect 34600 562700 34800 562900
rect 35000 562700 35200 562900
rect 35400 562700 35600 562900
rect 35800 562700 36000 562900
rect 36200 562700 36400 562900
rect 36600 562700 36800 562900
rect 37000 562700 37200 562900
rect 37400 562700 37600 562900
rect 37800 562700 38000 562900
rect 38200 562700 38400 562900
rect 38600 562700 38800 562900
rect 39000 562700 39200 562900
rect 39400 562700 39600 562900
rect 39800 562700 40000 562900
rect 40200 562700 40400 562900
rect 40600 562700 521280 562900
rect -800 562500 521280 562700
rect -800 562300 32800 562500
rect 33000 562300 33200 562500
rect 33400 562300 33600 562500
rect 33800 562300 34000 562500
rect 34200 562300 34400 562500
rect 34600 562300 34800 562500
rect 35000 562300 35200 562500
rect 35400 562300 35600 562500
rect 35800 562300 36000 562500
rect 36200 562300 36400 562500
rect 36600 562300 36800 562500
rect 37000 562300 37200 562500
rect 37400 562300 37600 562500
rect 37800 562300 38000 562500
rect 38200 562300 38400 562500
rect 38600 562300 38800 562500
rect 39000 562300 39200 562500
rect 39400 562300 39600 562500
rect 39800 562300 40000 562500
rect 40200 562300 40400 562500
rect 40600 562300 521280 562500
rect -800 562100 521280 562300
rect -800 561900 32800 562100
rect 33000 561900 33200 562100
rect 33400 561900 33600 562100
rect 33800 561900 34000 562100
rect 34200 561900 34400 562100
rect 34600 561900 34800 562100
rect 35000 561900 35200 562100
rect 35400 561900 35600 562100
rect 35800 561900 36000 562100
rect 36200 561900 36400 562100
rect 36600 561900 36800 562100
rect 37000 561900 37200 562100
rect 37400 561900 37600 562100
rect 37800 561900 38000 562100
rect 38200 561900 38400 562100
rect 38600 561900 38800 562100
rect 39000 561900 39200 562100
rect 39400 561900 39600 562100
rect 39800 561900 40000 562100
rect 40200 561900 40400 562100
rect 40600 561900 521280 562100
rect -800 561700 521280 561900
rect -800 561500 32800 561700
rect 33000 561500 33200 561700
rect 33400 561500 33600 561700
rect 33800 561500 34000 561700
rect 34200 561500 34400 561700
rect 34600 561500 34800 561700
rect 35000 561500 35200 561700
rect 35400 561500 35600 561700
rect 35800 561500 36000 561700
rect 36200 561500 36400 561700
rect 36600 561500 36800 561700
rect 37000 561500 37200 561700
rect 37400 561500 37600 561700
rect 37800 561500 38000 561700
rect 38200 561500 38400 561700
rect 38600 561500 38800 561700
rect 39000 561500 39200 561700
rect 39400 561500 39600 561700
rect 39800 561500 40000 561700
rect 40200 561500 40400 561700
rect 40600 561500 521280 561700
rect -800 561300 521280 561500
rect -800 561100 32800 561300
rect 33000 561100 33200 561300
rect 33400 561100 33600 561300
rect 33800 561100 34000 561300
rect 34200 561100 34400 561300
rect 34600 561100 34800 561300
rect 35000 561100 35200 561300
rect 35400 561100 35600 561300
rect 35800 561100 36000 561300
rect 36200 561100 36400 561300
rect 36600 561100 36800 561300
rect 37000 561100 37200 561300
rect 37400 561100 37600 561300
rect 37800 561100 38000 561300
rect 38200 561100 38400 561300
rect 38600 561100 38800 561300
rect 39000 561100 39200 561300
rect 39400 561100 39600 561300
rect 39800 561100 40000 561300
rect 40200 561100 40400 561300
rect 40600 561100 521280 561300
rect -800 560900 521280 561100
rect -800 560700 32800 560900
rect 33000 560700 33200 560900
rect 33400 560700 33600 560900
rect 33800 560700 34000 560900
rect 34200 560700 34400 560900
rect 34600 560700 34800 560900
rect 35000 560700 35200 560900
rect 35400 560700 35600 560900
rect 35800 560700 36000 560900
rect 36200 560700 36400 560900
rect 36600 560700 36800 560900
rect 37000 560700 37200 560900
rect 37400 560700 37600 560900
rect 37800 560700 38000 560900
rect 38200 560700 38400 560900
rect 38600 560700 38800 560900
rect 39000 560700 39200 560900
rect 39400 560700 39600 560900
rect 39800 560700 40000 560900
rect 40200 560700 40400 560900
rect 40600 560700 521280 560900
rect -800 560500 521280 560700
rect -800 560300 32800 560500
rect 33000 560300 33200 560500
rect 33400 560300 33600 560500
rect 33800 560300 34000 560500
rect 34200 560300 34400 560500
rect 34600 560300 34800 560500
rect 35000 560300 35200 560500
rect 35400 560300 35600 560500
rect 35800 560300 36000 560500
rect 36200 560300 36400 560500
rect 36600 560300 36800 560500
rect 37000 560300 37200 560500
rect 37400 560300 37600 560500
rect 37800 560300 38000 560500
rect 38200 560300 38400 560500
rect 38600 560300 38800 560500
rect 39000 560300 39200 560500
rect 39400 560300 39600 560500
rect 39800 560300 40000 560500
rect 40200 560300 40400 560500
rect 40600 560300 521280 560500
rect -800 560100 521280 560300
rect -800 559900 32800 560100
rect 33000 559900 33200 560100
rect 33400 559900 33600 560100
rect 33800 559900 34000 560100
rect 34200 559900 34400 560100
rect 34600 559900 34800 560100
rect 35000 559900 35200 560100
rect 35400 559900 35600 560100
rect 35800 559900 36000 560100
rect 36200 559900 36400 560100
rect 36600 559900 36800 560100
rect 37000 559900 37200 560100
rect 37400 559900 37600 560100
rect 37800 559900 38000 560100
rect 38200 559900 38400 560100
rect 38600 559900 38800 560100
rect 39000 559900 39200 560100
rect 39400 559900 39600 560100
rect 39800 559900 40000 560100
rect 40200 559900 40400 560100
rect 40600 559900 521280 560100
rect -800 559700 521280 559900
rect -800 559500 32800 559700
rect 33000 559500 33200 559700
rect 33400 559500 33600 559700
rect 33800 559500 34000 559700
rect 34200 559500 34400 559700
rect 34600 559500 34800 559700
rect 35000 559500 35200 559700
rect 35400 559500 35600 559700
rect 35800 559500 36000 559700
rect 36200 559500 36400 559700
rect 36600 559500 36800 559700
rect 37000 559500 37200 559700
rect 37400 559500 37600 559700
rect 37800 559500 38000 559700
rect 38200 559500 38400 559700
rect 38600 559500 38800 559700
rect 39000 559500 39200 559700
rect 39400 559500 39600 559700
rect 39800 559500 40000 559700
rect 40200 559500 40400 559700
rect 40600 559500 521280 559700
rect -800 559442 521280 559500
rect 0 559300 521280 559442
rect 0 559100 32800 559300
rect 33000 559100 33200 559300
rect 33400 559100 33600 559300
rect 33800 559100 34000 559300
rect 34200 559100 34400 559300
rect 34600 559100 34800 559300
rect 35000 559100 35200 559300
rect 35400 559100 35600 559300
rect 35800 559100 36000 559300
rect 36200 559100 36400 559300
rect 36600 559100 36800 559300
rect 37000 559100 37200 559300
rect 37400 559100 37600 559300
rect 37800 559100 38000 559300
rect 38200 559100 38400 559300
rect 38600 559100 38800 559300
rect 39000 559100 39200 559300
rect 39400 559100 39600 559300
rect 39800 559100 40000 559300
rect 40200 559100 40400 559300
rect 40600 559100 521280 559300
rect 0 558900 521280 559100
rect 0 558700 32800 558900
rect 33000 558700 33200 558900
rect 33400 558700 33600 558900
rect 33800 558700 34000 558900
rect 34200 558700 34400 558900
rect 34600 558700 34800 558900
rect 35000 558700 35200 558900
rect 35400 558700 35600 558900
rect 35800 558700 36000 558900
rect 36200 558700 36400 558900
rect 36600 558700 36800 558900
rect 37000 558700 37200 558900
rect 37400 558700 37600 558900
rect 37800 558700 38000 558900
rect 38200 558700 38400 558900
rect 38600 558700 38800 558900
rect 39000 558700 39200 558900
rect 39400 558700 39600 558900
rect 39800 558700 40000 558900
rect 40200 558700 40400 558900
rect 40600 558700 521280 558900
rect 0 558500 521280 558700
rect 0 558300 32800 558500
rect 33000 558300 33200 558500
rect 33400 558300 33600 558500
rect 33800 558300 34000 558500
rect 34200 558300 34400 558500
rect 34600 558300 34800 558500
rect 35000 558300 35200 558500
rect 35400 558300 35600 558500
rect 35800 558300 36000 558500
rect 36200 558300 36400 558500
rect 36600 558300 36800 558500
rect 37000 558300 37200 558500
rect 37400 558300 37600 558500
rect 37800 558300 38000 558500
rect 38200 558300 38400 558500
rect 38600 558300 38800 558500
rect 39000 558300 39200 558500
rect 39400 558300 39600 558500
rect 39800 558300 40000 558500
rect 40200 558300 40400 558500
rect 40600 558300 521280 558500
rect 0 558100 521280 558300
rect 0 557900 32800 558100
rect 33000 557900 33200 558100
rect 33400 557900 33600 558100
rect 33800 557900 34000 558100
rect 34200 557900 34400 558100
rect 34600 557900 34800 558100
rect 35000 557900 35200 558100
rect 35400 557900 35600 558100
rect 35800 557900 36000 558100
rect 36200 557900 36400 558100
rect 36600 557900 36800 558100
rect 37000 557900 37200 558100
rect 37400 557900 37600 558100
rect 37800 557900 38000 558100
rect 38200 557900 38400 558100
rect 38600 557900 38800 558100
rect 39000 557900 39200 558100
rect 39400 557900 39600 558100
rect 39800 557900 40000 558100
rect 40200 557900 40400 558100
rect 40600 557900 521280 558100
rect 0 557700 521280 557900
rect 0 557500 32800 557700
rect 33000 557500 33200 557700
rect 33400 557500 33600 557700
rect 33800 557500 34000 557700
rect 34200 557500 34400 557700
rect 34600 557500 34800 557700
rect 35000 557500 35200 557700
rect 35400 557500 35600 557700
rect 35800 557500 36000 557700
rect 36200 557500 36400 557700
rect 36600 557500 36800 557700
rect 37000 557500 37200 557700
rect 37400 557500 37600 557700
rect 37800 557500 38000 557700
rect 38200 557500 38400 557700
rect 38600 557500 38800 557700
rect 39000 557500 39200 557700
rect 39400 557500 39600 557700
rect 39800 557500 40000 557700
rect 40200 557500 40400 557700
rect 40600 557500 521280 557700
rect 0 557300 521280 557500
rect 0 557100 32800 557300
rect 33000 557100 33200 557300
rect 33400 557100 33600 557300
rect 33800 557100 34000 557300
rect 34200 557100 34400 557300
rect 34600 557100 34800 557300
rect 35000 557100 35200 557300
rect 35400 557100 35600 557300
rect 35800 557100 36000 557300
rect 36200 557100 36400 557300
rect 36600 557100 36800 557300
rect 37000 557100 37200 557300
rect 37400 557100 37600 557300
rect 37800 557100 38000 557300
rect 38200 557100 38400 557300
rect 38600 557100 38800 557300
rect 39000 557100 39200 557300
rect 39400 557100 39600 557300
rect 39800 557100 40000 557300
rect 40200 557100 40400 557300
rect 40600 557100 521280 557300
rect 0 556900 521280 557100
rect 0 556700 32800 556900
rect 33000 556700 33200 556900
rect 33400 556700 33600 556900
rect 33800 556700 34000 556900
rect 34200 556700 34400 556900
rect 34600 556700 34800 556900
rect 35000 556700 35200 556900
rect 35400 556700 35600 556900
rect 35800 556700 36000 556900
rect 36200 556700 36400 556900
rect 36600 556700 36800 556900
rect 37000 556700 37200 556900
rect 37400 556700 37600 556900
rect 37800 556700 38000 556900
rect 38200 556700 38400 556900
rect 38600 556700 38800 556900
rect 39000 556700 39200 556900
rect 39400 556700 39600 556900
rect 39800 556700 40000 556900
rect 40200 556700 40400 556900
rect 40600 556700 521280 556900
rect 0 556500 521280 556700
rect 0 556300 32800 556500
rect 33000 556300 33200 556500
rect 33400 556300 33600 556500
rect 33800 556300 34000 556500
rect 34200 556300 34400 556500
rect 34600 556300 34800 556500
rect 35000 556300 35200 556500
rect 35400 556300 35600 556500
rect 35800 556300 36000 556500
rect 36200 556300 36400 556500
rect 36600 556300 36800 556500
rect 37000 556300 37200 556500
rect 37400 556300 37600 556500
rect 37800 556300 38000 556500
rect 38200 556300 38400 556500
rect 38600 556300 38800 556500
rect 39000 556300 39200 556500
rect 39400 556300 39600 556500
rect 39800 556300 40000 556500
rect 40200 556300 40400 556500
rect 40600 556300 521280 556500
rect 0 556100 521280 556300
rect 0 555900 32800 556100
rect 33000 555900 33200 556100
rect 33400 555900 33600 556100
rect 33800 555900 34000 556100
rect 34200 555900 34400 556100
rect 34600 555900 34800 556100
rect 35000 555900 35200 556100
rect 35400 555900 35600 556100
rect 35800 555900 36000 556100
rect 36200 555900 36400 556100
rect 36600 555900 36800 556100
rect 37000 555900 37200 556100
rect 37400 555900 37600 556100
rect 37800 555900 38000 556100
rect 38200 555900 38400 556100
rect 38600 555900 38800 556100
rect 39000 555900 39200 556100
rect 39400 555900 39600 556100
rect 39800 555900 40000 556100
rect 40200 555900 40400 556100
rect 40600 555900 521280 556100
rect 0 555700 521280 555900
rect 0 555500 32800 555700
rect 33000 555500 33200 555700
rect 33400 555500 33600 555700
rect 33800 555500 34000 555700
rect 34200 555500 34400 555700
rect 34600 555500 34800 555700
rect 35000 555500 35200 555700
rect 35400 555500 35600 555700
rect 35800 555500 36000 555700
rect 36200 555500 36400 555700
rect 36600 555500 36800 555700
rect 37000 555500 37200 555700
rect 37400 555500 37600 555700
rect 37800 555500 38000 555700
rect 38200 555500 38400 555700
rect 38600 555500 38800 555700
rect 39000 555500 39200 555700
rect 39400 555500 39600 555700
rect 39800 555500 40000 555700
rect 40200 555500 40400 555700
rect 40600 555500 521280 555700
rect 0 555300 521280 555500
rect 0 555100 32800 555300
rect 33000 555100 33200 555300
rect 33400 555100 33600 555300
rect 33800 555100 34000 555300
rect 34200 555100 34400 555300
rect 34600 555100 34800 555300
rect 35000 555100 35200 555300
rect 35400 555100 35600 555300
rect 35800 555100 36000 555300
rect 36200 555100 36400 555300
rect 36600 555100 36800 555300
rect 37000 555100 37200 555300
rect 37400 555100 37600 555300
rect 37800 555100 38000 555300
rect 38200 555100 38400 555300
rect 38600 555100 38800 555300
rect 39000 555100 39200 555300
rect 39400 555100 39600 555300
rect 39800 555100 40000 555300
rect 40200 555100 40400 555300
rect 40600 555100 521280 555300
rect 0 554900 521280 555100
rect 0 554700 32800 554900
rect 33000 554700 33200 554900
rect 33400 554700 33600 554900
rect 33800 554700 34000 554900
rect 34200 554700 34400 554900
rect 34600 554700 34800 554900
rect 35000 554700 35200 554900
rect 35400 554700 35600 554900
rect 35800 554700 36000 554900
rect 36200 554700 36400 554900
rect 36600 554700 36800 554900
rect 37000 554700 37200 554900
rect 37400 554700 37600 554900
rect 37800 554700 38000 554900
rect 38200 554700 38400 554900
rect 38600 554700 38800 554900
rect 39000 554700 39200 554900
rect 39400 554700 39600 554900
rect 39800 554700 40000 554900
rect 40200 554700 40400 554900
rect 40600 554700 521280 554900
rect 0 554500 521280 554700
rect 0 554300 32800 554500
rect 33000 554300 33200 554500
rect 33400 554300 33600 554500
rect 33800 554300 34000 554500
rect 34200 554300 34400 554500
rect 34600 554300 34800 554500
rect 35000 554300 35200 554500
rect 35400 554300 35600 554500
rect 35800 554300 36000 554500
rect 36200 554300 36400 554500
rect 36600 554300 36800 554500
rect 37000 554300 37200 554500
rect 37400 554300 37600 554500
rect 37800 554300 38000 554500
rect 38200 554300 38400 554500
rect 38600 554300 38800 554500
rect 39000 554300 39200 554500
rect 39400 554300 39600 554500
rect 39800 554300 40000 554500
rect 40200 554300 40400 554500
rect 40600 554300 521280 554500
rect 0 554242 521280 554300
rect -800 554100 521280 554242
rect -800 553900 32800 554100
rect 33000 553900 33200 554100
rect 33400 553900 33600 554100
rect 33800 553900 34000 554100
rect 34200 553900 34400 554100
rect 34600 553900 34800 554100
rect 35000 553900 35200 554100
rect 35400 553900 35600 554100
rect 35800 553900 36000 554100
rect 36200 553900 36400 554100
rect 36600 553900 36800 554100
rect 37000 553900 37200 554100
rect 37400 553900 37600 554100
rect 37800 553900 38000 554100
rect 38200 553900 38400 554100
rect 38600 553900 38800 554100
rect 39000 553900 39200 554100
rect 39400 553900 39600 554100
rect 39800 553900 40000 554100
rect 40200 553900 40400 554100
rect 40600 553900 521280 554100
rect -800 553700 521280 553900
rect -800 553500 32800 553700
rect 33000 553500 33200 553700
rect 33400 553500 33600 553700
rect 33800 553500 34000 553700
rect 34200 553500 34400 553700
rect 34600 553500 34800 553700
rect 35000 553500 35200 553700
rect 35400 553500 35600 553700
rect 35800 553500 36000 553700
rect 36200 553500 36400 553700
rect 36600 553500 36800 553700
rect 37000 553500 37200 553700
rect 37400 553500 37600 553700
rect 37800 553500 38000 553700
rect 38200 553500 38400 553700
rect 38600 553500 38800 553700
rect 39000 553500 39200 553700
rect 39400 553500 39600 553700
rect 39800 553500 40000 553700
rect 40200 553500 40400 553700
rect 40600 553500 521280 553700
rect -800 553300 521280 553500
rect -800 553100 32800 553300
rect 33000 553100 33200 553300
rect 33400 553100 33600 553300
rect 33800 553100 34000 553300
rect 34200 553100 34400 553300
rect 34600 553100 34800 553300
rect 35000 553100 35200 553300
rect 35400 553100 35600 553300
rect 35800 553100 36000 553300
rect 36200 553100 36400 553300
rect 36600 553100 36800 553300
rect 37000 553100 37200 553300
rect 37400 553100 37600 553300
rect 37800 553100 38000 553300
rect 38200 553100 38400 553300
rect 38600 553100 38800 553300
rect 39000 553100 39200 553300
rect 39400 553100 39600 553300
rect 39800 553100 40000 553300
rect 40200 553100 40400 553300
rect 40600 553100 521280 553300
rect -800 552900 521280 553100
rect -800 552700 32800 552900
rect 33000 552700 33200 552900
rect 33400 552700 33600 552900
rect 33800 552700 34000 552900
rect 34200 552700 34400 552900
rect 34600 552700 34800 552900
rect 35000 552700 35200 552900
rect 35400 552700 35600 552900
rect 35800 552700 36000 552900
rect 36200 552700 36400 552900
rect 36600 552700 36800 552900
rect 37000 552700 37200 552900
rect 37400 552700 37600 552900
rect 37800 552700 38000 552900
rect 38200 552700 38400 552900
rect 38600 552700 38800 552900
rect 39000 552700 39200 552900
rect 39400 552700 39600 552900
rect 39800 552700 40000 552900
rect 40200 552700 40400 552900
rect 40600 552700 521280 552900
rect -800 552500 521280 552700
rect -800 552300 32800 552500
rect 33000 552300 33200 552500
rect 33400 552300 33600 552500
rect 33800 552300 34000 552500
rect 34200 552300 34400 552500
rect 34600 552300 34800 552500
rect 35000 552300 35200 552500
rect 35400 552300 35600 552500
rect 35800 552300 36000 552500
rect 36200 552300 36400 552500
rect 36600 552300 36800 552500
rect 37000 552300 37200 552500
rect 37400 552300 37600 552500
rect 37800 552300 38000 552500
rect 38200 552300 38400 552500
rect 38600 552300 38800 552500
rect 39000 552300 39200 552500
rect 39400 552300 39600 552500
rect 39800 552300 40000 552500
rect 40200 552300 40400 552500
rect 40600 552300 521280 552500
rect -800 552100 521280 552300
rect -800 551900 32800 552100
rect 33000 551900 33200 552100
rect 33400 551900 33600 552100
rect 33800 551900 34000 552100
rect 34200 551900 34400 552100
rect 34600 551900 34800 552100
rect 35000 551900 35200 552100
rect 35400 551900 35600 552100
rect 35800 551900 36000 552100
rect 36200 551900 36400 552100
rect 36600 551900 36800 552100
rect 37000 551900 37200 552100
rect 37400 551900 37600 552100
rect 37800 551900 38000 552100
rect 38200 551900 38400 552100
rect 38600 551900 38800 552100
rect 39000 551900 39200 552100
rect 39400 551900 39600 552100
rect 39800 551900 40000 552100
rect 40200 551900 40400 552100
rect 40600 551900 521280 552100
rect -800 551700 521280 551900
rect -800 551500 32800 551700
rect 33000 551500 33200 551700
rect 33400 551500 33600 551700
rect 33800 551500 34000 551700
rect 34200 551500 34400 551700
rect 34600 551500 34800 551700
rect 35000 551500 35200 551700
rect 35400 551500 35600 551700
rect 35800 551500 36000 551700
rect 36200 551500 36400 551700
rect 36600 551500 36800 551700
rect 37000 551500 37200 551700
rect 37400 551500 37600 551700
rect 37800 551500 38000 551700
rect 38200 551500 38400 551700
rect 38600 551500 38800 551700
rect 39000 551500 39200 551700
rect 39400 551500 39600 551700
rect 39800 551500 40000 551700
rect 40200 551500 40400 551700
rect 40600 551500 521280 551700
rect -800 551300 521280 551500
rect -800 551100 32800 551300
rect 33000 551100 33200 551300
rect 33400 551100 33600 551300
rect 33800 551100 34000 551300
rect 34200 551100 34400 551300
rect 34600 551100 34800 551300
rect 35000 551100 35200 551300
rect 35400 551100 35600 551300
rect 35800 551100 36000 551300
rect 36200 551100 36400 551300
rect 36600 551100 36800 551300
rect 37000 551100 37200 551300
rect 37400 551100 37600 551300
rect 37800 551100 38000 551300
rect 38200 551100 38400 551300
rect 38600 551100 38800 551300
rect 39000 551100 39200 551300
rect 39400 551100 39600 551300
rect 39800 551100 40000 551300
rect 40200 551100 40400 551300
rect 40600 551100 521280 551300
rect -800 550900 521280 551100
rect -800 550700 32800 550900
rect 33000 550700 33200 550900
rect 33400 550700 33600 550900
rect 33800 550700 34000 550900
rect 34200 550700 34400 550900
rect 34600 550700 34800 550900
rect 35000 550700 35200 550900
rect 35400 550700 35600 550900
rect 35800 550700 36000 550900
rect 36200 550700 36400 550900
rect 36600 550700 36800 550900
rect 37000 550700 37200 550900
rect 37400 550700 37600 550900
rect 37800 550700 38000 550900
rect 38200 550700 38400 550900
rect 38600 550700 38800 550900
rect 39000 550700 39200 550900
rect 39400 550700 39600 550900
rect 39800 550700 40000 550900
rect 40200 550700 40400 550900
rect 40600 550700 521280 550900
rect -800 550500 521280 550700
rect -800 550300 32800 550500
rect 33000 550300 33200 550500
rect 33400 550300 33600 550500
rect 33800 550300 34000 550500
rect 34200 550300 34400 550500
rect 34600 550300 34800 550500
rect 35000 550300 35200 550500
rect 35400 550300 35600 550500
rect 35800 550300 36000 550500
rect 36200 550300 36400 550500
rect 36600 550300 36800 550500
rect 37000 550300 37200 550500
rect 37400 550300 37600 550500
rect 37800 550300 38000 550500
rect 38200 550300 38400 550500
rect 38600 550300 38800 550500
rect 39000 550300 39200 550500
rect 39400 550300 39600 550500
rect 39800 550300 40000 550500
rect 40200 550300 40400 550500
rect 40600 550300 521280 550500
rect -800 550100 521280 550300
rect -800 549900 32800 550100
rect 33000 549900 33200 550100
rect 33400 549900 33600 550100
rect 33800 549900 34000 550100
rect 34200 549900 34400 550100
rect 34600 549900 34800 550100
rect 35000 549900 35200 550100
rect 35400 549900 35600 550100
rect 35800 549900 36000 550100
rect 36200 549900 36400 550100
rect 36600 549900 36800 550100
rect 37000 549900 37200 550100
rect 37400 549900 37600 550100
rect 37800 549900 38000 550100
rect 38200 549900 38400 550100
rect 38600 549900 38800 550100
rect 39000 549900 39200 550100
rect 39400 549900 39600 550100
rect 39800 549900 40000 550100
rect 40200 549900 40400 550100
rect 40600 549900 521280 550100
rect -800 549700 521280 549900
rect -800 549500 32800 549700
rect 33000 549500 33200 549700
rect 33400 549500 33600 549700
rect 33800 549500 34000 549700
rect 34200 549500 34400 549700
rect 34600 549500 34800 549700
rect 35000 549500 35200 549700
rect 35400 549500 35600 549700
rect 35800 549500 36000 549700
rect 36200 549500 36400 549700
rect 36600 549500 36800 549700
rect 37000 549500 37200 549700
rect 37400 549500 37600 549700
rect 37800 549500 38000 549700
rect 38200 549500 38400 549700
rect 38600 549500 38800 549700
rect 39000 549500 39200 549700
rect 39400 549500 39600 549700
rect 39800 549500 40000 549700
rect 40200 549500 40400 549700
rect 40600 549500 521280 549700
rect -800 549442 521280 549500
rect 0 549400 521280 549442
rect 29612 548300 521280 549400
<< via3 >>
rect 16400 702000 16600 702200
rect 16800 702000 17000 702200
rect 17200 702000 17400 702200
rect 17600 702000 17800 702200
rect 18000 702000 18200 702200
rect 18400 702000 18600 702200
rect 18800 702000 19000 702200
rect 19200 702000 19400 702200
rect 19600 702000 19800 702200
rect 20000 702000 20200 702200
rect 20400 702000 20600 702200
rect 20800 702000 21000 702200
rect 16400 701600 16600 701800
rect 16800 701600 17000 701800
rect 17200 701600 17400 701800
rect 17600 701600 17800 701800
rect 18000 701600 18200 701800
rect 18400 701600 18600 701800
rect 18800 701600 19000 701800
rect 19200 701600 19400 701800
rect 19600 701600 19800 701800
rect 20000 701600 20200 701800
rect 20400 701600 20600 701800
rect 20800 701600 21000 701800
rect 16400 701200 16600 701400
rect 16800 701200 17000 701400
rect 17200 701200 17400 701400
rect 17600 701200 17800 701400
rect 18000 701200 18200 701400
rect 18400 701200 18600 701400
rect 18800 701200 19000 701400
rect 19200 701200 19400 701400
rect 19600 701200 19800 701400
rect 20000 701200 20200 701400
rect 20400 701200 20600 701400
rect 20800 701200 21000 701400
rect 68400 702000 68600 702200
rect 68800 702000 69000 702200
rect 69200 702000 69400 702200
rect 69600 702000 69800 702200
rect 70000 702000 70200 702200
rect 70400 702000 70600 702200
rect 70800 702000 71000 702200
rect 71200 702000 71400 702200
rect 71600 702000 71800 702200
rect 72000 702000 72200 702200
rect 72400 702000 72600 702200
rect 72800 702000 73000 702200
rect 68400 701600 68600 701800
rect 68800 701600 69000 701800
rect 69200 701600 69400 701800
rect 69600 701600 69800 701800
rect 70000 701600 70200 701800
rect 70400 701600 70600 701800
rect 70800 701600 71000 701800
rect 71200 701600 71400 701800
rect 71600 701600 71800 701800
rect 72000 701600 72200 701800
rect 72400 701600 72600 701800
rect 72800 701600 73000 701800
rect 68400 701200 68600 701400
rect 68800 701200 69000 701400
rect 69200 701200 69400 701400
rect 69600 701200 69800 701400
rect 70000 701200 70200 701400
rect 70400 701200 70600 701400
rect 70800 701200 71000 701400
rect 71200 701200 71400 701400
rect 71600 701200 71800 701400
rect 72000 701200 72200 701400
rect 72400 701200 72600 701400
rect 72800 701200 73000 701400
rect 16400 700800 16600 701000
rect 16800 700800 17000 701000
rect 17200 700800 17400 701000
rect 17600 700800 17800 701000
rect 18000 700800 18200 701000
rect 18400 700800 18600 701000
rect 18800 700800 19000 701000
rect 19200 700800 19400 701000
rect 19600 700800 19800 701000
rect 20000 700800 20200 701000
rect 20400 700800 20600 701000
rect 20800 700800 21000 701000
rect 16400 700400 16600 700600
rect 16800 700400 17000 700600
rect 17200 700400 17400 700600
rect 17600 700400 17800 700600
rect 18000 700400 18200 700600
rect 18400 700400 18600 700600
rect 18800 700400 19000 700600
rect 19200 700400 19400 700600
rect 19600 700400 19800 700600
rect 20000 700400 20200 700600
rect 20400 700400 20600 700600
rect 20800 700400 21000 700600
rect 16400 700000 16600 700200
rect 16800 700000 17000 700200
rect 17200 700000 17400 700200
rect 17600 700000 17800 700200
rect 18000 700000 18200 700200
rect 18400 700000 18600 700200
rect 18800 700000 19000 700200
rect 19200 700000 19400 700200
rect 19600 700000 19800 700200
rect 20000 700000 20200 700200
rect 20400 700000 20600 700200
rect 20800 700000 21000 700200
rect 37278 701045 40622 701109
rect 41078 701045 44422 701109
rect 44878 701045 48222 701109
rect 48678 701045 52022 701109
rect 68400 700800 68600 701000
rect 68800 700800 69000 701000
rect 69200 700800 69400 701000
rect 69600 700800 69800 701000
rect 70000 700800 70200 701000
rect 70400 700800 70600 701000
rect 70800 700800 71000 701000
rect 71200 700800 71400 701000
rect 71600 700800 71800 701000
rect 72000 700800 72200 701000
rect 72400 700800 72600 701000
rect 72800 700800 73000 701000
rect 68400 700400 68600 700600
rect 68800 700400 69000 700600
rect 69200 700400 69400 700600
rect 69600 700400 69800 700600
rect 70000 700400 70200 700600
rect 70400 700400 70600 700600
rect 70800 700400 71000 700600
rect 71200 700400 71400 700600
rect 71600 700400 71800 700600
rect 72000 700400 72200 700600
rect 72400 700400 72600 700600
rect 72800 700400 73000 700600
rect 68400 700000 68600 700200
rect 68800 700000 69000 700200
rect 69200 700000 69400 700200
rect 69600 700000 69800 700200
rect 70000 700000 70200 700200
rect 70400 700000 70600 700200
rect 70800 700000 71000 700200
rect 71200 700000 71400 700200
rect 71600 700000 71800 700200
rect 72000 700000 72200 700200
rect 72400 700000 72600 700200
rect 72800 700000 73000 700200
rect 44010 695370 44280 695640
rect 45060 695370 45330 695640
rect 41840 695090 41850 695140
rect 41850 695090 42090 695140
rect 36930 694850 37000 694920
rect 41840 694920 42090 695090
rect 41840 694890 41850 694920
rect 41850 694890 42090 694920
rect 43740 694880 43990 695130
rect 45320 694880 45570 695130
rect 47220 694880 47470 695130
rect 52320 694850 52390 694920
rect 36820 694740 36890 694810
rect 52430 694740 52500 694810
rect 40710 693860 40800 693960
rect 40900 693860 40990 693960
rect 44010 693730 44280 694000
rect 45060 693730 45330 694000
rect 48320 693860 48410 693960
rect 48510 693860 48600 693960
rect 38700 693360 38880 693460
rect 39120 693360 39300 693460
rect 43340 693420 43350 693480
rect 43350 693420 43590 693480
rect 43590 693420 43600 693480
rect 44610 693420 44860 693480
rect 44860 693420 44870 693480
rect 45870 693420 45880 693480
rect 45880 693420 46120 693480
rect 46120 693420 46130 693480
rect 43340 693280 43600 693420
rect 44610 693280 44870 693420
rect 45870 693280 46130 693420
rect 49950 693360 50130 693460
rect 50370 693360 50550 693460
rect 43340 693220 43350 693280
rect 43350 693220 43590 693280
rect 43590 693220 43600 693280
rect 44610 693220 44860 693280
rect 44860 693220 44870 693280
rect 45870 693220 45880 693280
rect 45880 693220 46120 693280
rect 46120 693220 46130 693280
rect 43780 692130 44040 692390
rect 45280 692130 45540 692390
rect 43340 691870 43350 691930
rect 43350 691870 43590 691930
rect 43590 691870 43600 691930
rect 44610 691870 44860 691930
rect 44860 691870 44870 691930
rect 45870 691870 45880 691930
rect 45880 691870 46120 691930
rect 46120 691870 46130 691930
rect 43340 691730 43600 691870
rect 44610 691730 44870 691870
rect 45870 691730 46130 691870
rect 43340 691670 43350 691730
rect 43350 691670 43590 691730
rect 43590 691670 43600 691730
rect 44610 691670 44860 691730
rect 44860 691670 44870 691730
rect 45870 691670 45880 691730
rect 45880 691670 46120 691730
rect 46120 691670 46130 691730
rect 58000 691700 58200 691900
rect 58400 691700 58600 691900
rect 58800 691700 59000 691900
rect 59200 691700 59400 691900
rect 59600 691700 59800 691900
rect 60000 691700 60200 691900
rect 60400 691700 60600 691900
rect 60800 691700 61000 691900
rect 61200 691700 61400 691900
rect 61600 691700 61800 691900
rect 534639 694862 534739 694992
rect 534899 694862 534999 694992
rect 68400 690000 68600 690200
rect 68800 690000 69000 690200
rect 69200 690000 69400 690200
rect 69600 690000 69800 690200
rect 70000 690000 70200 690200
rect 70400 690000 70600 690200
rect 70800 690000 71000 690200
rect 71200 690000 71400 690200
rect 71600 690000 71800 690200
rect 72000 690000 72200 690200
rect 72400 690000 72600 690200
rect 72800 690000 73000 690200
rect 68400 689600 68600 689800
rect 68800 689600 69000 689800
rect 69200 689600 69400 689800
rect 69600 689600 69800 689800
rect 70000 689600 70200 689800
rect 70400 689600 70600 689800
rect 70800 689600 71000 689800
rect 71200 689600 71400 689800
rect 71600 689600 71800 689800
rect 72000 689600 72200 689800
rect 72400 689600 72600 689800
rect 72800 689600 73000 689800
rect 532300 690200 532500 690400
rect 532700 690200 532900 690400
rect 533100 690200 533300 690400
rect 533500 690200 533700 690400
rect 533900 690200 534100 690400
rect 532300 689900 532500 690100
rect 532700 689900 532900 690100
rect 533100 689900 533300 690100
rect 533500 689900 533700 690100
rect 533900 689900 534100 690100
rect 532300 689500 532500 689700
rect 532700 689500 532900 689700
rect 533100 689500 533300 689700
rect 533500 689500 533700 689700
rect 533900 689500 534100 689700
rect 44520 689030 44780 689290
rect 532300 689100 532500 689300
rect 532700 689100 532900 689300
rect 533100 689100 533300 689300
rect 533500 689100 533700 689300
rect 533900 689100 534100 689300
rect 16400 688500 16600 688700
rect 16800 688500 17000 688700
rect 17200 688500 17400 688700
rect 17600 688500 17800 688700
rect 18000 688500 18200 688700
rect 18400 688500 18600 688700
rect 18800 688500 19000 688700
rect 19200 688500 19400 688700
rect 19600 688500 19800 688700
rect 20000 688500 20200 688700
rect 20400 688500 20600 688700
rect 20800 688500 21000 688700
rect 532300 688700 532500 688900
rect 532700 688700 532900 688900
rect 533100 688700 533300 688900
rect 533500 688700 533700 688900
rect 533900 688700 534100 688900
rect 16400 688100 16600 688300
rect 16800 688100 17000 688300
rect 17200 688100 17400 688300
rect 17600 688100 17800 688300
rect 18000 688100 18200 688300
rect 18400 688100 18600 688300
rect 18800 688100 19000 688300
rect 19200 688100 19400 688300
rect 19600 688100 19800 688300
rect 20000 688100 20200 688300
rect 20400 688100 20600 688300
rect 20800 688100 21000 688300
rect 537197 694857 540541 694921
rect 540997 694857 544341 694921
rect 544797 694857 548141 694921
rect 548597 694857 551941 694921
rect 554129 694862 554239 694992
rect 554389 694862 554499 694992
rect 541089 690602 541169 690682
rect 541239 690602 541319 690682
rect 543579 690602 543659 690682
rect 543729 690602 543809 690682
rect 546059 690602 546139 690682
rect 546209 690602 546289 690682
rect 541089 690062 541169 690142
rect 541239 690062 541319 690142
rect 543579 690062 543659 690142
rect 543729 690062 543809 690142
rect 546059 690062 546139 690142
rect 546209 690062 546289 690142
rect 541089 689522 541169 689602
rect 541239 689522 541319 689602
rect 543579 689522 543659 689602
rect 543729 689522 543809 689602
rect 546069 689522 546149 689602
rect 546209 689522 546289 689602
rect 542379 688922 542459 689002
rect 542489 688922 542569 689002
rect 544789 688922 544869 689002
rect 544899 688922 544979 689002
rect 547249 688912 547329 688992
rect 547359 688912 547439 688992
rect 542379 688312 542459 688392
rect 542489 688312 542569 688392
rect 544789 688332 544869 688412
rect 544899 688332 544979 688412
rect 547249 688332 547329 688412
rect 547359 688332 547439 688412
rect 44520 687510 44780 687770
rect 542380 687750 542460 687830
rect 542500 687750 542580 687830
rect 544789 687752 544869 687832
rect 544899 687752 544979 687832
rect 547249 687752 547329 687832
rect 547359 687752 547439 687832
rect 538869 687542 538959 687652
rect 539029 687542 539119 687652
rect 548799 687522 548879 687602
rect 548969 687522 549049 687602
rect 36800 687100 37000 687300
rect 37200 687100 37400 687300
rect 37600 687100 37800 687300
rect 38000 687100 38200 687300
rect 549900 687142 550100 687200
rect 550200 687142 550400 687200
rect 549900 687062 550069 687142
rect 550069 687062 550100 687142
rect 550200 687062 550229 687142
rect 550229 687062 550319 687142
rect 550319 687062 550400 687142
rect 549900 687000 550100 687062
rect 550200 687000 550400 687062
rect 550500 687000 550700 687200
rect 550800 687000 551000 687200
rect 551200 687100 551400 687300
rect 551200 686800 551400 687000
rect 43500 686420 43750 686670
rect 45560 686420 45810 686670
rect 551200 686500 551400 686700
rect 44530 686000 44780 686250
rect 551200 686200 551400 686400
rect 549800 685900 550000 686100
rect 550100 686062 550300 686100
rect 550100 685982 550159 686062
rect 550159 685982 550229 686062
rect 550229 685982 550300 686062
rect 550100 685900 550300 685982
rect 550400 685900 550600 686100
rect 550800 685900 551000 686100
rect 36800 685100 37000 685300
rect 37200 685100 37400 685300
rect 37600 685100 37800 685300
rect 38000 685100 38200 685300
rect 36800 684700 37000 684900
rect 37200 684700 37400 684900
rect 37600 684700 37800 684900
rect 38000 684700 38200 684900
rect 43240 684900 43490 685150
rect 45820 684900 46070 685150
rect 542379 685052 542459 685132
rect 542489 685052 542569 685132
rect 544789 685052 544869 685132
rect 544899 685052 544979 685132
rect 547249 685062 547329 685142
rect 547359 685062 547439 685142
rect 36800 684300 37000 684500
rect 37200 684300 37400 684500
rect 37600 684300 37800 684500
rect 38000 684300 38200 684500
rect 44530 684470 44780 684720
rect 515700 684600 515900 684800
rect 516100 684600 516300 684800
rect 516500 684600 516700 684800
rect 516900 684600 517100 684800
rect 517300 684600 517500 684800
rect 517700 684600 517900 684800
rect 518100 684600 518300 684800
rect 518500 684600 518700 684800
rect 518900 684600 519100 684800
rect 519300 684600 519500 684800
rect 519700 684600 519900 684800
rect 520100 684600 520300 684800
rect 520500 684600 520700 684800
rect 36800 683900 37000 684100
rect 37200 683900 37400 684100
rect 37600 683900 37800 684100
rect 38000 683900 38200 684100
rect 36800 683500 37000 683700
rect 37200 683500 37400 683700
rect 37600 683500 37800 683700
rect 38000 683500 38200 683700
rect 515700 684200 515900 684400
rect 516100 684200 516300 684400
rect 516500 684200 516700 684400
rect 516900 684200 517100 684400
rect 517300 684200 517500 684400
rect 517700 684200 517900 684400
rect 518100 684200 518300 684400
rect 518500 684200 518700 684400
rect 518900 684200 519100 684400
rect 519300 684200 519500 684400
rect 519700 684200 519900 684400
rect 520100 684200 520300 684400
rect 520500 684200 520700 684400
rect 541089 684292 541169 684372
rect 541239 684292 541319 684372
rect 543579 684312 543659 684392
rect 543729 684312 543809 684392
rect 546059 684312 546139 684392
rect 546199 684312 546279 684392
rect 515700 683800 515900 684000
rect 516100 683800 516300 684000
rect 516500 683800 516700 684000
rect 516900 683800 517100 684000
rect 517300 683800 517500 684000
rect 517700 683800 517900 684000
rect 518100 683800 518300 684000
rect 518500 683800 518700 684000
rect 518900 683800 519100 684000
rect 519300 683800 519500 684000
rect 519700 683800 519900 684000
rect 520100 683800 520300 684000
rect 520500 683800 520700 684000
rect 43810 683600 43930 683620
rect 43810 683520 43840 683600
rect 43840 683520 43920 683600
rect 43920 683520 43930 683600
rect 44350 683520 44430 683600
rect 44870 683520 44950 683600
rect 45390 683520 45470 683600
rect 43810 683500 43930 683520
rect 36800 683100 37000 683300
rect 37200 683100 37400 683300
rect 37600 683100 37800 683300
rect 38000 683100 38200 683300
rect 515700 683400 515900 683600
rect 516100 683400 516300 683600
rect 516500 683400 516700 683600
rect 516900 683400 517100 683600
rect 517300 683400 517500 683600
rect 517700 683400 517900 683600
rect 518100 683400 518300 683600
rect 518500 683400 518700 683600
rect 518900 683400 519100 683600
rect 519300 683400 519500 683600
rect 519700 683400 519900 683600
rect 520100 683400 520300 683600
rect 520500 683400 520700 683600
rect 36800 682700 37000 682900
rect 37200 682700 37400 682900
rect 37600 682700 37800 682900
rect 38000 682700 38200 682900
rect 36800 682300 37000 682500
rect 37200 682300 37400 682500
rect 37600 682300 37800 682500
rect 38000 682300 38200 682500
rect 515700 683000 515900 683200
rect 516100 683000 516300 683200
rect 516500 683000 516700 683200
rect 516900 683000 517100 683200
rect 517300 683000 517500 683200
rect 517700 683000 517900 683200
rect 518100 683000 518300 683200
rect 518500 683000 518700 683200
rect 518900 683000 519100 683200
rect 519300 683000 519500 683200
rect 519700 683000 519900 683200
rect 520100 683000 520300 683200
rect 520500 683000 520700 683200
rect 515700 682600 515900 682800
rect 516100 682600 516300 682800
rect 516500 682600 516700 682800
rect 516900 682600 517100 682800
rect 517300 682600 517500 682800
rect 517700 682600 517900 682800
rect 518100 682600 518300 682800
rect 518500 682600 518700 682800
rect 518900 682600 519100 682800
rect 519300 682600 519500 682800
rect 519700 682600 519900 682800
rect 520100 682600 520300 682800
rect 520500 682600 520700 682800
rect 546389 682342 546509 682442
rect 36800 681900 37000 682100
rect 37200 681900 37400 682100
rect 37600 681900 37800 682100
rect 38000 681900 38200 682100
rect 43630 682060 43710 682140
rect 45590 682060 45670 682140
rect 58000 682000 58200 682200
rect 58400 682000 58600 682200
rect 58800 682000 59000 682200
rect 59200 682000 59400 682200
rect 59600 682000 59800 682200
rect 60000 682000 60200 682200
rect 60400 682000 60600 682200
rect 60800 682000 61000 682200
rect 61200 682000 61400 682200
rect 61600 682000 61800 682200
rect 36800 681500 37000 681700
rect 37200 681500 37400 681700
rect 37600 681500 37800 681700
rect 38000 681500 38200 681700
rect 43630 681840 43710 681920
rect 43630 681700 43710 681780
rect 45590 681840 45670 681920
rect 45590 681700 45670 681780
rect 36800 681100 37000 681300
rect 37200 681100 37400 681300
rect 37600 681100 37800 681300
rect 38000 681100 38200 681300
rect 36800 680700 37000 680900
rect 37200 680700 37400 680900
rect 37600 680700 37800 680900
rect 38000 680700 38200 680900
rect 549800 681200 550000 681400
rect 550200 681200 550400 681400
rect 550600 681200 550800 681400
rect 551000 681200 551200 681400
rect 551400 681200 551600 681400
rect 551800 681200 552000 681400
rect 552200 681200 552400 681400
rect 552600 681200 552800 681400
rect 549800 680800 550000 681000
rect 550200 680800 550400 681000
rect 550600 680800 550800 681000
rect 551000 680800 551200 681000
rect 551400 680800 551600 681000
rect 551800 680800 552000 681000
rect 552200 680800 552400 681000
rect 552600 680800 552800 681000
rect 36800 680300 37000 680500
rect 37200 680300 37400 680500
rect 37600 680300 37800 680500
rect 38000 680300 38200 680500
rect 44270 680400 44390 680520
rect 44890 680410 45010 680530
rect 44590 679540 44680 679630
rect 44580 679160 44670 679250
rect 515900 679000 516100 679200
rect 516300 679000 516500 679200
rect 516700 679000 516900 679200
rect 517100 679000 517300 679200
rect 517500 679000 517700 679200
rect 517900 679000 518100 679200
rect 518300 679000 518500 679200
rect 518700 679000 518900 679200
rect 519100 679000 519300 679200
rect 519500 679000 519700 679200
rect 519900 679000 520100 679200
rect 520300 679000 520500 679200
rect 520700 679000 520900 679200
rect 515900 678600 516100 678800
rect 516300 678600 516500 678800
rect 516700 678600 516900 678800
rect 517100 678600 517300 678800
rect 517500 678600 517700 678800
rect 517900 678600 518100 678800
rect 518300 678600 518500 678800
rect 518700 678600 518900 678800
rect 519100 678600 519300 678800
rect 519500 678600 519700 678800
rect 519900 678600 520100 678800
rect 520300 678600 520500 678800
rect 520700 678600 520900 678800
rect 515900 678200 516100 678400
rect 516300 678200 516500 678400
rect 516700 678200 516900 678400
rect 517100 678200 517300 678400
rect 517500 678200 517700 678400
rect 517900 678200 518100 678400
rect 518300 678200 518500 678400
rect 518700 678200 518900 678400
rect 519100 678200 519300 678400
rect 519500 678200 519700 678400
rect 519900 678200 520100 678400
rect 520300 678200 520500 678400
rect 520700 678200 520900 678400
rect 44580 677720 44670 677810
rect 515900 677800 516100 678000
rect 516300 677800 516500 678000
rect 516700 677800 516900 678000
rect 517100 677800 517300 678000
rect 517500 677800 517700 678000
rect 517900 677800 518100 678000
rect 518300 677800 518500 678000
rect 518700 677800 518900 678000
rect 519100 677800 519300 678000
rect 519500 677800 519700 678000
rect 519900 677800 520100 678000
rect 520300 677800 520500 678000
rect 520700 677800 520900 678000
rect 515900 677400 516100 677600
rect 516300 677400 516500 677600
rect 516700 677400 516900 677600
rect 517100 677400 517300 677600
rect 517500 677400 517700 677600
rect 517900 677400 518100 677600
rect 518300 677400 518500 677600
rect 518700 677400 518900 677600
rect 519100 677400 519300 677600
rect 519500 677400 519700 677600
rect 519900 677400 520100 677600
rect 520300 677400 520500 677600
rect 520700 677400 520900 677600
rect 515900 677000 516100 677200
rect 516300 677000 516500 677200
rect 516700 677000 516900 677200
rect 517100 677000 517300 677200
rect 517500 677000 517700 677200
rect 517900 677000 518100 677200
rect 518300 677000 518500 677200
rect 518700 677000 518900 677200
rect 519100 677000 519300 677200
rect 519500 677000 519700 677200
rect 519900 677000 520100 677200
rect 520300 677000 520500 677200
rect 520700 677000 520900 677200
rect 515900 676600 516100 676800
rect 516300 676600 516500 676800
rect 516700 676600 516900 676800
rect 517100 676600 517300 676800
rect 517500 676600 517700 676800
rect 517900 676600 518100 676800
rect 518300 676600 518500 676800
rect 518700 676600 518900 676800
rect 519100 676600 519300 676800
rect 519500 676600 519700 676800
rect 519900 676600 520100 676800
rect 520300 676600 520500 676800
rect 520700 676600 520900 676800
rect 41200 673300 41440 673540
rect 47900 673300 48140 673540
rect 41200 670100 41440 670340
rect 47900 670100 48140 670340
rect 41200 666780 41440 667020
rect 47900 666780 48140 667020
rect 32800 663000 33100 663300
rect 33300 663000 33600 663300
rect 33800 663000 34100 663300
rect 34300 663000 34600 663300
rect 34800 663000 35100 663300
rect 35300 663000 35600 663300
rect 35800 663000 36100 663300
rect 36300 663000 36600 663300
rect 36800 663000 37100 663300
rect 37300 663000 37600 663300
rect 37800 663000 38100 663300
rect 38300 663000 38600 663300
rect 38800 663000 39100 663300
rect 39300 663000 39600 663300
rect 39800 663000 40100 663300
rect 40300 663000 40600 663300
rect 2500 648300 2800 648600
rect 3000 648300 3300 648600
rect 3500 648300 3800 648600
rect 2500 647800 2800 648100
rect 3000 647800 3300 648100
rect 3500 647800 3800 648100
rect 2500 647300 2800 647600
rect 3000 647300 3300 647600
rect 3500 647300 3800 647600
rect 2500 646800 2800 647100
rect 3000 646800 3300 647100
rect 3500 646800 3800 647100
rect 2500 646300 2800 646600
rect 3000 646300 3300 646600
rect 3500 646300 3800 646600
rect 2500 645800 2800 646100
rect 3000 645800 3300 646100
rect 3500 645800 3800 646100
rect 2500 645300 2800 645600
rect 3000 645300 3300 645600
rect 3500 645300 3800 645600
rect 2500 644800 2800 645100
rect 3000 644800 3300 645100
rect 3500 644800 3800 645100
rect 2500 644300 2800 644600
rect 3000 644300 3300 644600
rect 3500 644300 3800 644600
rect 2500 643800 2800 644100
rect 3000 643800 3300 644100
rect 3500 643800 3800 644100
rect 2500 643300 2800 643600
rect 3000 643300 3300 643600
rect 3500 643300 3800 643600
rect 2500 642800 2800 643100
rect 3000 642800 3300 643100
rect 3500 642800 3800 643100
rect 2500 642300 2800 642600
rect 3000 642300 3300 642600
rect 3500 642300 3800 642600
rect 2500 641800 2800 642100
rect 3000 641800 3300 642100
rect 3500 641800 3800 642100
rect 2500 641300 2800 641600
rect 3000 641300 3300 641600
rect 3500 641300 3800 641600
rect 2500 640800 2800 641100
rect 3000 640800 3300 641100
rect 3500 640800 3800 641100
rect 2500 640300 2800 640600
rect 3000 640300 3300 640600
rect 3500 640300 3800 640600
rect 2500 639800 2800 640100
rect 3000 639800 3300 640100
rect 3500 639800 3800 640100
rect 2500 639300 2800 639600
rect 3000 639300 3300 639600
rect 3500 639300 3800 639600
rect 2500 638800 2800 639100
rect 3000 638800 3300 639100
rect 3500 638800 3800 639100
rect 2500 638300 2800 638600
rect 3000 638300 3300 638600
rect 3500 638300 3800 638600
rect 2500 637800 2800 638100
rect 3000 637800 3300 638100
rect 3500 637800 3800 638100
rect 2500 637300 2800 637600
rect 3000 637300 3300 637600
rect 3500 637300 3800 637600
rect 2500 636800 2800 637100
rect 3000 636800 3300 637100
rect 3500 636800 3800 637100
rect 2500 636300 2800 636600
rect 3000 636300 3300 636600
rect 3500 636300 3800 636600
rect 2500 635800 2800 636100
rect 3000 635800 3300 636100
rect 3500 635800 3800 636100
rect 2500 635300 2800 635600
rect 3000 635300 3300 635600
rect 3500 635300 3800 635600
rect 2500 634800 2800 635100
rect 3000 634800 3300 635100
rect 3500 634800 3800 635100
rect 2500 634300 2800 634600
rect 3000 634300 3300 634600
rect 3500 634300 3800 634600
rect 550000 644400 550200 644600
rect 550400 644400 550600 644600
rect 550800 644400 551000 644600
rect 551200 644400 551400 644600
rect 551600 644400 551800 644600
rect 552000 644400 552200 644600
rect 552400 644400 552600 644600
rect 552800 644400 553000 644600
rect 550000 644000 550200 644200
rect 550400 644000 550600 644200
rect 550800 644000 551000 644200
rect 551200 644000 551400 644200
rect 551600 644000 551800 644200
rect 552000 644000 552200 644200
rect 552400 644000 552600 644200
rect 552800 644000 553000 644200
rect 550000 643600 550200 643800
rect 550400 643600 550600 643800
rect 550800 643600 551000 643800
rect 551200 643600 551400 643800
rect 551600 643600 551800 643800
rect 552000 643600 552200 643800
rect 552400 643600 552600 643800
rect 552800 643600 553000 643800
rect 550000 643200 550200 643400
rect 550400 643200 550600 643400
rect 550800 643200 551000 643400
rect 551200 643200 551400 643400
rect 551600 643200 551800 643400
rect 552000 643200 552200 643400
rect 552400 643200 552600 643400
rect 552800 643200 553000 643400
rect 550000 642800 550200 643000
rect 550400 642800 550600 643000
rect 550800 642800 551000 643000
rect 551200 642800 551400 643000
rect 551600 642800 551800 643000
rect 552000 642800 552200 643000
rect 552400 642800 552600 643000
rect 552800 642800 553000 643000
rect 550000 642400 550200 642600
rect 550400 642400 550600 642600
rect 550800 642400 551000 642600
rect 551200 642400 551400 642600
rect 551600 642400 551800 642600
rect 552000 642400 552200 642600
rect 552400 642400 552600 642600
rect 552800 642400 553000 642600
rect 550000 642000 550200 642200
rect 550400 642000 550600 642200
rect 550800 642000 551000 642200
rect 551200 642000 551400 642200
rect 551600 642000 551800 642200
rect 552000 642000 552200 642200
rect 552400 642000 552600 642200
rect 552800 642000 553000 642200
rect 550000 641600 550200 641800
rect 550400 641600 550600 641800
rect 550800 641600 551000 641800
rect 551200 641600 551400 641800
rect 551600 641600 551800 641800
rect 552000 641600 552200 641800
rect 552400 641600 552600 641800
rect 552800 641600 553000 641800
rect 550000 641200 550200 641400
rect 550400 641200 550600 641400
rect 550800 641200 551000 641400
rect 551200 641200 551400 641400
rect 551600 641200 551800 641400
rect 552000 641200 552200 641400
rect 552400 641200 552600 641400
rect 552800 641200 553000 641400
rect 550000 640800 550200 641000
rect 550400 640800 550600 641000
rect 550800 640800 551000 641000
rect 551200 640800 551400 641000
rect 551600 640800 551800 641000
rect 552000 640800 552200 641000
rect 552400 640800 552600 641000
rect 552800 640800 553000 641000
rect 550000 640400 550200 640600
rect 550400 640400 550600 640600
rect 550800 640400 551000 640600
rect 551200 640400 551400 640600
rect 551600 640400 551800 640600
rect 552000 640400 552200 640600
rect 552400 640400 552600 640600
rect 552800 640400 553000 640600
rect 550000 640000 550200 640200
rect 550400 640000 550600 640200
rect 550800 640000 551000 640200
rect 551200 640000 551400 640200
rect 551600 640000 551800 640200
rect 552000 640000 552200 640200
rect 552400 640000 552600 640200
rect 552800 640000 553000 640200
rect 550000 639600 550200 639800
rect 550400 639600 550600 639800
rect 550800 639600 551000 639800
rect 551200 639600 551400 639800
rect 551600 639600 551800 639800
rect 552000 639600 552200 639800
rect 552400 639600 552600 639800
rect 552800 639600 553000 639800
rect 550000 639200 550200 639400
rect 550400 639200 550600 639400
rect 550800 639200 551000 639400
rect 551200 639200 551400 639400
rect 551600 639200 551800 639400
rect 552000 639200 552200 639400
rect 552400 639200 552600 639400
rect 552800 639200 553000 639400
rect 550000 638800 550200 639000
rect 550400 638800 550600 639000
rect 550800 638800 551000 639000
rect 551200 638800 551400 639000
rect 551600 638800 551800 639000
rect 552000 638800 552200 639000
rect 552400 638800 552600 639000
rect 552800 638800 553000 639000
rect 550000 638400 550200 638600
rect 550400 638400 550600 638600
rect 550800 638400 551000 638600
rect 551200 638400 551400 638600
rect 551600 638400 551800 638600
rect 552000 638400 552200 638600
rect 552400 638400 552600 638600
rect 552800 638400 553000 638600
rect 550000 638000 550200 638200
rect 550400 638000 550600 638200
rect 550800 638000 551000 638200
rect 551200 638000 551400 638200
rect 551600 638000 551800 638200
rect 552000 638000 552200 638200
rect 552400 638000 552600 638200
rect 552800 638000 553000 638200
rect 550000 637600 550200 637800
rect 550400 637600 550600 637800
rect 550800 637600 551000 637800
rect 551200 637600 551400 637800
rect 551600 637600 551800 637800
rect 552000 637600 552200 637800
rect 552400 637600 552600 637800
rect 552800 637600 553000 637800
rect 550000 637200 550200 637400
rect 550400 637200 550600 637400
rect 550800 637200 551000 637400
rect 551200 637200 551400 637400
rect 551600 637200 551800 637400
rect 552000 637200 552200 637400
rect 552400 637200 552600 637400
rect 552800 637200 553000 637400
rect 550000 636800 550200 637000
rect 550400 636800 550600 637000
rect 550800 636800 551000 637000
rect 551200 636800 551400 637000
rect 551600 636800 551800 637000
rect 552000 636800 552200 637000
rect 552400 636800 552600 637000
rect 552800 636800 553000 637000
rect 550000 636400 550200 636600
rect 550400 636400 550600 636600
rect 550800 636400 551000 636600
rect 551200 636400 551400 636600
rect 551600 636400 551800 636600
rect 552000 636400 552200 636600
rect 552400 636400 552600 636600
rect 552800 636400 553000 636600
rect 550000 636000 550200 636200
rect 550400 636000 550600 636200
rect 550800 636000 551000 636200
rect 551200 636000 551400 636200
rect 551600 636000 551800 636200
rect 552000 636000 552200 636200
rect 552400 636000 552600 636200
rect 552800 636000 553000 636200
rect 550000 635600 550200 635800
rect 550400 635600 550600 635800
rect 550800 635600 551000 635800
rect 551200 635600 551400 635800
rect 551600 635600 551800 635800
rect 552000 635600 552200 635800
rect 552400 635600 552600 635800
rect 552800 635600 553000 635800
rect 550000 635200 550200 635400
rect 550400 635200 550600 635400
rect 550800 635200 551000 635400
rect 551200 635200 551400 635400
rect 551600 635200 551800 635400
rect 552000 635200 552200 635400
rect 552400 635200 552600 635400
rect 552800 635200 553000 635400
rect 550000 634800 550200 635000
rect 550400 634800 550600 635000
rect 550800 634800 551000 635000
rect 551200 634800 551400 635000
rect 551600 634800 551800 635000
rect 552000 634800 552200 635000
rect 552400 634800 552600 635000
rect 552800 634800 553000 635000
rect 550000 634400 550200 634600
rect 550400 634400 550600 634600
rect 550800 634400 551000 634600
rect 551200 634400 551400 634600
rect 551600 634400 551800 634600
rect 552000 634400 552200 634600
rect 552400 634400 552600 634600
rect 552800 634400 553000 634600
rect 550000 634000 550200 634200
rect 550400 634000 550600 634200
rect 550800 634000 551000 634200
rect 551200 634000 551400 634200
rect 551600 634000 551800 634200
rect 552000 634000 552200 634200
rect 552400 634000 552600 634200
rect 552800 634000 553000 634200
rect 550000 633600 550200 633800
rect 550400 633600 550600 633800
rect 550800 633600 551000 633800
rect 551200 633600 551400 633800
rect 551600 633600 551800 633800
rect 552000 633600 552200 633800
rect 552400 633600 552600 633800
rect 552800 633600 553000 633800
rect 550000 633200 550200 633400
rect 550400 633200 550600 633400
rect 550800 633200 551000 633400
rect 551200 633200 551400 633400
rect 551600 633200 551800 633400
rect 552000 633200 552200 633400
rect 552400 633200 552600 633400
rect 552800 633200 553000 633400
rect 550000 632800 550200 633000
rect 550400 632800 550600 633000
rect 550800 632800 551000 633000
rect 551200 632800 551400 633000
rect 551600 632800 551800 633000
rect 552000 632800 552200 633000
rect 552400 632800 552600 633000
rect 552800 632800 553000 633000
rect 550000 632400 550200 632600
rect 550400 632400 550600 632600
rect 550800 632400 551000 632600
rect 551200 632400 551400 632600
rect 551600 632400 551800 632600
rect 552000 632400 552200 632600
rect 552400 632400 552600 632600
rect 552800 632400 553000 632600
rect 550000 632000 550200 632200
rect 550400 632000 550600 632200
rect 550800 632000 551000 632200
rect 551200 632000 551400 632200
rect 551600 632000 551800 632200
rect 552000 632000 552200 632200
rect 552400 632000 552600 632200
rect 552800 632000 553000 632200
rect 550000 631600 550200 631800
rect 550400 631600 550600 631800
rect 550800 631600 551000 631800
rect 551200 631600 551400 631800
rect 551600 631600 551800 631800
rect 552000 631600 552200 631800
rect 552400 631600 552600 631800
rect 552800 631600 553000 631800
rect 550000 631200 550200 631400
rect 550400 631200 550600 631400
rect 550800 631200 551000 631400
rect 551200 631200 551400 631400
rect 551600 631200 551800 631400
rect 552000 631200 552200 631400
rect 552400 631200 552600 631400
rect 552800 631200 553000 631400
rect 550000 630800 550200 631000
rect 550400 630800 550600 631000
rect 550800 630800 551000 631000
rect 551200 630800 551400 631000
rect 551600 630800 551800 631000
rect 552000 630800 552200 631000
rect 552400 630800 552600 631000
rect 552800 630800 553000 631000
rect 550000 630500 550200 630700
rect 550400 630500 550600 630700
rect 550800 630500 551000 630700
rect 551200 630500 551400 630700
rect 551600 630500 551800 630700
rect 552000 630500 552200 630700
rect 552400 630500 552600 630700
rect 552800 630500 553000 630700
rect 550000 630200 550200 630400
rect 550400 630200 550600 630400
rect 550800 630200 551000 630400
rect 551200 630200 551400 630400
rect 551600 630200 551800 630400
rect 552000 630200 552200 630400
rect 552400 630200 552600 630400
rect 552800 630200 553000 630400
rect 550000 629800 550200 630000
rect 550400 629800 550600 630000
rect 550800 629800 551000 630000
rect 551200 629800 551400 630000
rect 551600 629800 551800 630000
rect 552000 629800 552200 630000
rect 552400 629800 552600 630000
rect 552800 629800 553000 630000
rect 32800 563900 33000 564100
rect 33200 563900 33400 564100
rect 33600 563900 33800 564100
rect 34000 563900 34200 564100
rect 34400 563900 34600 564100
rect 34800 563900 35000 564100
rect 35200 563900 35400 564100
rect 35600 563900 35800 564100
rect 36000 563900 36200 564100
rect 36400 563900 36600 564100
rect 36800 563900 37000 564100
rect 37200 563900 37400 564100
rect 37600 563900 37800 564100
rect 38000 563900 38200 564100
rect 38400 563900 38600 564100
rect 38800 563900 39000 564100
rect 39200 563900 39400 564100
rect 39600 563900 39800 564100
rect 40000 563900 40200 564100
rect 40400 563900 40600 564100
rect 32800 563500 33000 563700
rect 33200 563500 33400 563700
rect 33600 563500 33800 563700
rect 34000 563500 34200 563700
rect 34400 563500 34600 563700
rect 34800 563500 35000 563700
rect 35200 563500 35400 563700
rect 35600 563500 35800 563700
rect 36000 563500 36200 563700
rect 36400 563500 36600 563700
rect 36800 563500 37000 563700
rect 37200 563500 37400 563700
rect 37600 563500 37800 563700
rect 38000 563500 38200 563700
rect 38400 563500 38600 563700
rect 38800 563500 39000 563700
rect 39200 563500 39400 563700
rect 39600 563500 39800 563700
rect 40000 563500 40200 563700
rect 40400 563500 40600 563700
rect 32800 563100 33000 563300
rect 33200 563100 33400 563300
rect 33600 563100 33800 563300
rect 34000 563100 34200 563300
rect 34400 563100 34600 563300
rect 34800 563100 35000 563300
rect 35200 563100 35400 563300
rect 35600 563100 35800 563300
rect 36000 563100 36200 563300
rect 36400 563100 36600 563300
rect 36800 563100 37000 563300
rect 37200 563100 37400 563300
rect 37600 563100 37800 563300
rect 38000 563100 38200 563300
rect 38400 563100 38600 563300
rect 38800 563100 39000 563300
rect 39200 563100 39400 563300
rect 39600 563100 39800 563300
rect 40000 563100 40200 563300
rect 40400 563100 40600 563300
rect 32800 562700 33000 562900
rect 33200 562700 33400 562900
rect 33600 562700 33800 562900
rect 34000 562700 34200 562900
rect 34400 562700 34600 562900
rect 34800 562700 35000 562900
rect 35200 562700 35400 562900
rect 35600 562700 35800 562900
rect 36000 562700 36200 562900
rect 36400 562700 36600 562900
rect 36800 562700 37000 562900
rect 37200 562700 37400 562900
rect 37600 562700 37800 562900
rect 38000 562700 38200 562900
rect 38400 562700 38600 562900
rect 38800 562700 39000 562900
rect 39200 562700 39400 562900
rect 39600 562700 39800 562900
rect 40000 562700 40200 562900
rect 40400 562700 40600 562900
rect 32800 562300 33000 562500
rect 33200 562300 33400 562500
rect 33600 562300 33800 562500
rect 34000 562300 34200 562500
rect 34400 562300 34600 562500
rect 34800 562300 35000 562500
rect 35200 562300 35400 562500
rect 35600 562300 35800 562500
rect 36000 562300 36200 562500
rect 36400 562300 36600 562500
rect 36800 562300 37000 562500
rect 37200 562300 37400 562500
rect 37600 562300 37800 562500
rect 38000 562300 38200 562500
rect 38400 562300 38600 562500
rect 38800 562300 39000 562500
rect 39200 562300 39400 562500
rect 39600 562300 39800 562500
rect 40000 562300 40200 562500
rect 40400 562300 40600 562500
rect 32800 561900 33000 562100
rect 33200 561900 33400 562100
rect 33600 561900 33800 562100
rect 34000 561900 34200 562100
rect 34400 561900 34600 562100
rect 34800 561900 35000 562100
rect 35200 561900 35400 562100
rect 35600 561900 35800 562100
rect 36000 561900 36200 562100
rect 36400 561900 36600 562100
rect 36800 561900 37000 562100
rect 37200 561900 37400 562100
rect 37600 561900 37800 562100
rect 38000 561900 38200 562100
rect 38400 561900 38600 562100
rect 38800 561900 39000 562100
rect 39200 561900 39400 562100
rect 39600 561900 39800 562100
rect 40000 561900 40200 562100
rect 40400 561900 40600 562100
rect 32800 561500 33000 561700
rect 33200 561500 33400 561700
rect 33600 561500 33800 561700
rect 34000 561500 34200 561700
rect 34400 561500 34600 561700
rect 34800 561500 35000 561700
rect 35200 561500 35400 561700
rect 35600 561500 35800 561700
rect 36000 561500 36200 561700
rect 36400 561500 36600 561700
rect 36800 561500 37000 561700
rect 37200 561500 37400 561700
rect 37600 561500 37800 561700
rect 38000 561500 38200 561700
rect 38400 561500 38600 561700
rect 38800 561500 39000 561700
rect 39200 561500 39400 561700
rect 39600 561500 39800 561700
rect 40000 561500 40200 561700
rect 40400 561500 40600 561700
rect 32800 561100 33000 561300
rect 33200 561100 33400 561300
rect 33600 561100 33800 561300
rect 34000 561100 34200 561300
rect 34400 561100 34600 561300
rect 34800 561100 35000 561300
rect 35200 561100 35400 561300
rect 35600 561100 35800 561300
rect 36000 561100 36200 561300
rect 36400 561100 36600 561300
rect 36800 561100 37000 561300
rect 37200 561100 37400 561300
rect 37600 561100 37800 561300
rect 38000 561100 38200 561300
rect 38400 561100 38600 561300
rect 38800 561100 39000 561300
rect 39200 561100 39400 561300
rect 39600 561100 39800 561300
rect 40000 561100 40200 561300
rect 40400 561100 40600 561300
rect 32800 560700 33000 560900
rect 33200 560700 33400 560900
rect 33600 560700 33800 560900
rect 34000 560700 34200 560900
rect 34400 560700 34600 560900
rect 34800 560700 35000 560900
rect 35200 560700 35400 560900
rect 35600 560700 35800 560900
rect 36000 560700 36200 560900
rect 36400 560700 36600 560900
rect 36800 560700 37000 560900
rect 37200 560700 37400 560900
rect 37600 560700 37800 560900
rect 38000 560700 38200 560900
rect 38400 560700 38600 560900
rect 38800 560700 39000 560900
rect 39200 560700 39400 560900
rect 39600 560700 39800 560900
rect 40000 560700 40200 560900
rect 40400 560700 40600 560900
rect 32800 560300 33000 560500
rect 33200 560300 33400 560500
rect 33600 560300 33800 560500
rect 34000 560300 34200 560500
rect 34400 560300 34600 560500
rect 34800 560300 35000 560500
rect 35200 560300 35400 560500
rect 35600 560300 35800 560500
rect 36000 560300 36200 560500
rect 36400 560300 36600 560500
rect 36800 560300 37000 560500
rect 37200 560300 37400 560500
rect 37600 560300 37800 560500
rect 38000 560300 38200 560500
rect 38400 560300 38600 560500
rect 38800 560300 39000 560500
rect 39200 560300 39400 560500
rect 39600 560300 39800 560500
rect 40000 560300 40200 560500
rect 40400 560300 40600 560500
rect 32800 559900 33000 560100
rect 33200 559900 33400 560100
rect 33600 559900 33800 560100
rect 34000 559900 34200 560100
rect 34400 559900 34600 560100
rect 34800 559900 35000 560100
rect 35200 559900 35400 560100
rect 35600 559900 35800 560100
rect 36000 559900 36200 560100
rect 36400 559900 36600 560100
rect 36800 559900 37000 560100
rect 37200 559900 37400 560100
rect 37600 559900 37800 560100
rect 38000 559900 38200 560100
rect 38400 559900 38600 560100
rect 38800 559900 39000 560100
rect 39200 559900 39400 560100
rect 39600 559900 39800 560100
rect 40000 559900 40200 560100
rect 40400 559900 40600 560100
rect 32800 559500 33000 559700
rect 33200 559500 33400 559700
rect 33600 559500 33800 559700
rect 34000 559500 34200 559700
rect 34400 559500 34600 559700
rect 34800 559500 35000 559700
rect 35200 559500 35400 559700
rect 35600 559500 35800 559700
rect 36000 559500 36200 559700
rect 36400 559500 36600 559700
rect 36800 559500 37000 559700
rect 37200 559500 37400 559700
rect 37600 559500 37800 559700
rect 38000 559500 38200 559700
rect 38400 559500 38600 559700
rect 38800 559500 39000 559700
rect 39200 559500 39400 559700
rect 39600 559500 39800 559700
rect 40000 559500 40200 559700
rect 40400 559500 40600 559700
rect 32800 559100 33000 559300
rect 33200 559100 33400 559300
rect 33600 559100 33800 559300
rect 34000 559100 34200 559300
rect 34400 559100 34600 559300
rect 34800 559100 35000 559300
rect 35200 559100 35400 559300
rect 35600 559100 35800 559300
rect 36000 559100 36200 559300
rect 36400 559100 36600 559300
rect 36800 559100 37000 559300
rect 37200 559100 37400 559300
rect 37600 559100 37800 559300
rect 38000 559100 38200 559300
rect 38400 559100 38600 559300
rect 38800 559100 39000 559300
rect 39200 559100 39400 559300
rect 39600 559100 39800 559300
rect 40000 559100 40200 559300
rect 40400 559100 40600 559300
rect 32800 558700 33000 558900
rect 33200 558700 33400 558900
rect 33600 558700 33800 558900
rect 34000 558700 34200 558900
rect 34400 558700 34600 558900
rect 34800 558700 35000 558900
rect 35200 558700 35400 558900
rect 35600 558700 35800 558900
rect 36000 558700 36200 558900
rect 36400 558700 36600 558900
rect 36800 558700 37000 558900
rect 37200 558700 37400 558900
rect 37600 558700 37800 558900
rect 38000 558700 38200 558900
rect 38400 558700 38600 558900
rect 38800 558700 39000 558900
rect 39200 558700 39400 558900
rect 39600 558700 39800 558900
rect 40000 558700 40200 558900
rect 40400 558700 40600 558900
rect 32800 558300 33000 558500
rect 33200 558300 33400 558500
rect 33600 558300 33800 558500
rect 34000 558300 34200 558500
rect 34400 558300 34600 558500
rect 34800 558300 35000 558500
rect 35200 558300 35400 558500
rect 35600 558300 35800 558500
rect 36000 558300 36200 558500
rect 36400 558300 36600 558500
rect 36800 558300 37000 558500
rect 37200 558300 37400 558500
rect 37600 558300 37800 558500
rect 38000 558300 38200 558500
rect 38400 558300 38600 558500
rect 38800 558300 39000 558500
rect 39200 558300 39400 558500
rect 39600 558300 39800 558500
rect 40000 558300 40200 558500
rect 40400 558300 40600 558500
rect 32800 557900 33000 558100
rect 33200 557900 33400 558100
rect 33600 557900 33800 558100
rect 34000 557900 34200 558100
rect 34400 557900 34600 558100
rect 34800 557900 35000 558100
rect 35200 557900 35400 558100
rect 35600 557900 35800 558100
rect 36000 557900 36200 558100
rect 36400 557900 36600 558100
rect 36800 557900 37000 558100
rect 37200 557900 37400 558100
rect 37600 557900 37800 558100
rect 38000 557900 38200 558100
rect 38400 557900 38600 558100
rect 38800 557900 39000 558100
rect 39200 557900 39400 558100
rect 39600 557900 39800 558100
rect 40000 557900 40200 558100
rect 40400 557900 40600 558100
rect 32800 557500 33000 557700
rect 33200 557500 33400 557700
rect 33600 557500 33800 557700
rect 34000 557500 34200 557700
rect 34400 557500 34600 557700
rect 34800 557500 35000 557700
rect 35200 557500 35400 557700
rect 35600 557500 35800 557700
rect 36000 557500 36200 557700
rect 36400 557500 36600 557700
rect 36800 557500 37000 557700
rect 37200 557500 37400 557700
rect 37600 557500 37800 557700
rect 38000 557500 38200 557700
rect 38400 557500 38600 557700
rect 38800 557500 39000 557700
rect 39200 557500 39400 557700
rect 39600 557500 39800 557700
rect 40000 557500 40200 557700
rect 40400 557500 40600 557700
rect 32800 557100 33000 557300
rect 33200 557100 33400 557300
rect 33600 557100 33800 557300
rect 34000 557100 34200 557300
rect 34400 557100 34600 557300
rect 34800 557100 35000 557300
rect 35200 557100 35400 557300
rect 35600 557100 35800 557300
rect 36000 557100 36200 557300
rect 36400 557100 36600 557300
rect 36800 557100 37000 557300
rect 37200 557100 37400 557300
rect 37600 557100 37800 557300
rect 38000 557100 38200 557300
rect 38400 557100 38600 557300
rect 38800 557100 39000 557300
rect 39200 557100 39400 557300
rect 39600 557100 39800 557300
rect 40000 557100 40200 557300
rect 40400 557100 40600 557300
rect 32800 556700 33000 556900
rect 33200 556700 33400 556900
rect 33600 556700 33800 556900
rect 34000 556700 34200 556900
rect 34400 556700 34600 556900
rect 34800 556700 35000 556900
rect 35200 556700 35400 556900
rect 35600 556700 35800 556900
rect 36000 556700 36200 556900
rect 36400 556700 36600 556900
rect 36800 556700 37000 556900
rect 37200 556700 37400 556900
rect 37600 556700 37800 556900
rect 38000 556700 38200 556900
rect 38400 556700 38600 556900
rect 38800 556700 39000 556900
rect 39200 556700 39400 556900
rect 39600 556700 39800 556900
rect 40000 556700 40200 556900
rect 40400 556700 40600 556900
rect 32800 556300 33000 556500
rect 33200 556300 33400 556500
rect 33600 556300 33800 556500
rect 34000 556300 34200 556500
rect 34400 556300 34600 556500
rect 34800 556300 35000 556500
rect 35200 556300 35400 556500
rect 35600 556300 35800 556500
rect 36000 556300 36200 556500
rect 36400 556300 36600 556500
rect 36800 556300 37000 556500
rect 37200 556300 37400 556500
rect 37600 556300 37800 556500
rect 38000 556300 38200 556500
rect 38400 556300 38600 556500
rect 38800 556300 39000 556500
rect 39200 556300 39400 556500
rect 39600 556300 39800 556500
rect 40000 556300 40200 556500
rect 40400 556300 40600 556500
rect 32800 555900 33000 556100
rect 33200 555900 33400 556100
rect 33600 555900 33800 556100
rect 34000 555900 34200 556100
rect 34400 555900 34600 556100
rect 34800 555900 35000 556100
rect 35200 555900 35400 556100
rect 35600 555900 35800 556100
rect 36000 555900 36200 556100
rect 36400 555900 36600 556100
rect 36800 555900 37000 556100
rect 37200 555900 37400 556100
rect 37600 555900 37800 556100
rect 38000 555900 38200 556100
rect 38400 555900 38600 556100
rect 38800 555900 39000 556100
rect 39200 555900 39400 556100
rect 39600 555900 39800 556100
rect 40000 555900 40200 556100
rect 40400 555900 40600 556100
rect 32800 555500 33000 555700
rect 33200 555500 33400 555700
rect 33600 555500 33800 555700
rect 34000 555500 34200 555700
rect 34400 555500 34600 555700
rect 34800 555500 35000 555700
rect 35200 555500 35400 555700
rect 35600 555500 35800 555700
rect 36000 555500 36200 555700
rect 36400 555500 36600 555700
rect 36800 555500 37000 555700
rect 37200 555500 37400 555700
rect 37600 555500 37800 555700
rect 38000 555500 38200 555700
rect 38400 555500 38600 555700
rect 38800 555500 39000 555700
rect 39200 555500 39400 555700
rect 39600 555500 39800 555700
rect 40000 555500 40200 555700
rect 40400 555500 40600 555700
rect 32800 555100 33000 555300
rect 33200 555100 33400 555300
rect 33600 555100 33800 555300
rect 34000 555100 34200 555300
rect 34400 555100 34600 555300
rect 34800 555100 35000 555300
rect 35200 555100 35400 555300
rect 35600 555100 35800 555300
rect 36000 555100 36200 555300
rect 36400 555100 36600 555300
rect 36800 555100 37000 555300
rect 37200 555100 37400 555300
rect 37600 555100 37800 555300
rect 38000 555100 38200 555300
rect 38400 555100 38600 555300
rect 38800 555100 39000 555300
rect 39200 555100 39400 555300
rect 39600 555100 39800 555300
rect 40000 555100 40200 555300
rect 40400 555100 40600 555300
rect 32800 554700 33000 554900
rect 33200 554700 33400 554900
rect 33600 554700 33800 554900
rect 34000 554700 34200 554900
rect 34400 554700 34600 554900
rect 34800 554700 35000 554900
rect 35200 554700 35400 554900
rect 35600 554700 35800 554900
rect 36000 554700 36200 554900
rect 36400 554700 36600 554900
rect 36800 554700 37000 554900
rect 37200 554700 37400 554900
rect 37600 554700 37800 554900
rect 38000 554700 38200 554900
rect 38400 554700 38600 554900
rect 38800 554700 39000 554900
rect 39200 554700 39400 554900
rect 39600 554700 39800 554900
rect 40000 554700 40200 554900
rect 40400 554700 40600 554900
rect 32800 554300 33000 554500
rect 33200 554300 33400 554500
rect 33600 554300 33800 554500
rect 34000 554300 34200 554500
rect 34400 554300 34600 554500
rect 34800 554300 35000 554500
rect 35200 554300 35400 554500
rect 35600 554300 35800 554500
rect 36000 554300 36200 554500
rect 36400 554300 36600 554500
rect 36800 554300 37000 554500
rect 37200 554300 37400 554500
rect 37600 554300 37800 554500
rect 38000 554300 38200 554500
rect 38400 554300 38600 554500
rect 38800 554300 39000 554500
rect 39200 554300 39400 554500
rect 39600 554300 39800 554500
rect 40000 554300 40200 554500
rect 40400 554300 40600 554500
rect 32800 553900 33000 554100
rect 33200 553900 33400 554100
rect 33600 553900 33800 554100
rect 34000 553900 34200 554100
rect 34400 553900 34600 554100
rect 34800 553900 35000 554100
rect 35200 553900 35400 554100
rect 35600 553900 35800 554100
rect 36000 553900 36200 554100
rect 36400 553900 36600 554100
rect 36800 553900 37000 554100
rect 37200 553900 37400 554100
rect 37600 553900 37800 554100
rect 38000 553900 38200 554100
rect 38400 553900 38600 554100
rect 38800 553900 39000 554100
rect 39200 553900 39400 554100
rect 39600 553900 39800 554100
rect 40000 553900 40200 554100
rect 40400 553900 40600 554100
rect 32800 553500 33000 553700
rect 33200 553500 33400 553700
rect 33600 553500 33800 553700
rect 34000 553500 34200 553700
rect 34400 553500 34600 553700
rect 34800 553500 35000 553700
rect 35200 553500 35400 553700
rect 35600 553500 35800 553700
rect 36000 553500 36200 553700
rect 36400 553500 36600 553700
rect 36800 553500 37000 553700
rect 37200 553500 37400 553700
rect 37600 553500 37800 553700
rect 38000 553500 38200 553700
rect 38400 553500 38600 553700
rect 38800 553500 39000 553700
rect 39200 553500 39400 553700
rect 39600 553500 39800 553700
rect 40000 553500 40200 553700
rect 40400 553500 40600 553700
rect 32800 553100 33000 553300
rect 33200 553100 33400 553300
rect 33600 553100 33800 553300
rect 34000 553100 34200 553300
rect 34400 553100 34600 553300
rect 34800 553100 35000 553300
rect 35200 553100 35400 553300
rect 35600 553100 35800 553300
rect 36000 553100 36200 553300
rect 36400 553100 36600 553300
rect 36800 553100 37000 553300
rect 37200 553100 37400 553300
rect 37600 553100 37800 553300
rect 38000 553100 38200 553300
rect 38400 553100 38600 553300
rect 38800 553100 39000 553300
rect 39200 553100 39400 553300
rect 39600 553100 39800 553300
rect 40000 553100 40200 553300
rect 40400 553100 40600 553300
rect 32800 552700 33000 552900
rect 33200 552700 33400 552900
rect 33600 552700 33800 552900
rect 34000 552700 34200 552900
rect 34400 552700 34600 552900
rect 34800 552700 35000 552900
rect 35200 552700 35400 552900
rect 35600 552700 35800 552900
rect 36000 552700 36200 552900
rect 36400 552700 36600 552900
rect 36800 552700 37000 552900
rect 37200 552700 37400 552900
rect 37600 552700 37800 552900
rect 38000 552700 38200 552900
rect 38400 552700 38600 552900
rect 38800 552700 39000 552900
rect 39200 552700 39400 552900
rect 39600 552700 39800 552900
rect 40000 552700 40200 552900
rect 40400 552700 40600 552900
rect 32800 552300 33000 552500
rect 33200 552300 33400 552500
rect 33600 552300 33800 552500
rect 34000 552300 34200 552500
rect 34400 552300 34600 552500
rect 34800 552300 35000 552500
rect 35200 552300 35400 552500
rect 35600 552300 35800 552500
rect 36000 552300 36200 552500
rect 36400 552300 36600 552500
rect 36800 552300 37000 552500
rect 37200 552300 37400 552500
rect 37600 552300 37800 552500
rect 38000 552300 38200 552500
rect 38400 552300 38600 552500
rect 38800 552300 39000 552500
rect 39200 552300 39400 552500
rect 39600 552300 39800 552500
rect 40000 552300 40200 552500
rect 40400 552300 40600 552500
rect 32800 551900 33000 552100
rect 33200 551900 33400 552100
rect 33600 551900 33800 552100
rect 34000 551900 34200 552100
rect 34400 551900 34600 552100
rect 34800 551900 35000 552100
rect 35200 551900 35400 552100
rect 35600 551900 35800 552100
rect 36000 551900 36200 552100
rect 36400 551900 36600 552100
rect 36800 551900 37000 552100
rect 37200 551900 37400 552100
rect 37600 551900 37800 552100
rect 38000 551900 38200 552100
rect 38400 551900 38600 552100
rect 38800 551900 39000 552100
rect 39200 551900 39400 552100
rect 39600 551900 39800 552100
rect 40000 551900 40200 552100
rect 40400 551900 40600 552100
rect 32800 551500 33000 551700
rect 33200 551500 33400 551700
rect 33600 551500 33800 551700
rect 34000 551500 34200 551700
rect 34400 551500 34600 551700
rect 34800 551500 35000 551700
rect 35200 551500 35400 551700
rect 35600 551500 35800 551700
rect 36000 551500 36200 551700
rect 36400 551500 36600 551700
rect 36800 551500 37000 551700
rect 37200 551500 37400 551700
rect 37600 551500 37800 551700
rect 38000 551500 38200 551700
rect 38400 551500 38600 551700
rect 38800 551500 39000 551700
rect 39200 551500 39400 551700
rect 39600 551500 39800 551700
rect 40000 551500 40200 551700
rect 40400 551500 40600 551700
rect 32800 551100 33000 551300
rect 33200 551100 33400 551300
rect 33600 551100 33800 551300
rect 34000 551100 34200 551300
rect 34400 551100 34600 551300
rect 34800 551100 35000 551300
rect 35200 551100 35400 551300
rect 35600 551100 35800 551300
rect 36000 551100 36200 551300
rect 36400 551100 36600 551300
rect 36800 551100 37000 551300
rect 37200 551100 37400 551300
rect 37600 551100 37800 551300
rect 38000 551100 38200 551300
rect 38400 551100 38600 551300
rect 38800 551100 39000 551300
rect 39200 551100 39400 551300
rect 39600 551100 39800 551300
rect 40000 551100 40200 551300
rect 40400 551100 40600 551300
rect 32800 550700 33000 550900
rect 33200 550700 33400 550900
rect 33600 550700 33800 550900
rect 34000 550700 34200 550900
rect 34400 550700 34600 550900
rect 34800 550700 35000 550900
rect 35200 550700 35400 550900
rect 35600 550700 35800 550900
rect 36000 550700 36200 550900
rect 36400 550700 36600 550900
rect 36800 550700 37000 550900
rect 37200 550700 37400 550900
rect 37600 550700 37800 550900
rect 38000 550700 38200 550900
rect 38400 550700 38600 550900
rect 38800 550700 39000 550900
rect 39200 550700 39400 550900
rect 39600 550700 39800 550900
rect 40000 550700 40200 550900
rect 40400 550700 40600 550900
rect 32800 550300 33000 550500
rect 33200 550300 33400 550500
rect 33600 550300 33800 550500
rect 34000 550300 34200 550500
rect 34400 550300 34600 550500
rect 34800 550300 35000 550500
rect 35200 550300 35400 550500
rect 35600 550300 35800 550500
rect 36000 550300 36200 550500
rect 36400 550300 36600 550500
rect 36800 550300 37000 550500
rect 37200 550300 37400 550500
rect 37600 550300 37800 550500
rect 38000 550300 38200 550500
rect 38400 550300 38600 550500
rect 38800 550300 39000 550500
rect 39200 550300 39400 550500
rect 39600 550300 39800 550500
rect 40000 550300 40200 550500
rect 40400 550300 40600 550500
rect 32800 549900 33000 550100
rect 33200 549900 33400 550100
rect 33600 549900 33800 550100
rect 34000 549900 34200 550100
rect 34400 549900 34600 550100
rect 34800 549900 35000 550100
rect 35200 549900 35400 550100
rect 35600 549900 35800 550100
rect 36000 549900 36200 550100
rect 36400 549900 36600 550100
rect 36800 549900 37000 550100
rect 37200 549900 37400 550100
rect 37600 549900 37800 550100
rect 38000 549900 38200 550100
rect 38400 549900 38600 550100
rect 38800 549900 39000 550100
rect 39200 549900 39400 550100
rect 39600 549900 39800 550100
rect 40000 549900 40200 550100
rect 40400 549900 40600 550100
rect 32800 549500 33000 549700
rect 33200 549500 33400 549700
rect 33600 549500 33800 549700
rect 34000 549500 34200 549700
rect 34400 549500 34600 549700
rect 34800 549500 35000 549700
rect 35200 549500 35400 549700
rect 35600 549500 35800 549700
rect 36000 549500 36200 549700
rect 36400 549500 36600 549700
rect 36800 549500 37000 549700
rect 37200 549500 37400 549700
rect 37600 549500 37800 549700
rect 38000 549500 38200 549700
rect 38400 549500 38600 549700
rect 38800 549500 39000 549700
rect 39200 549500 39400 549700
rect 39600 549500 39800 549700
rect 40000 549500 40200 549700
rect 40400 549500 40600 549700
<< mimcap >>
rect 37350 700890 40550 700930
rect 37350 697770 37390 700890
rect 40510 697770 40550 700890
rect 37350 697730 40550 697770
rect 41150 700890 44350 700930
rect 41150 697770 41190 700890
rect 44310 697770 44350 700890
rect 41150 697730 44350 697770
rect 44950 700890 48150 700930
rect 44950 697770 44990 700890
rect 48110 697770 48150 700890
rect 44950 697730 48150 697770
rect 48750 700890 51950 700930
rect 48750 697770 48790 700890
rect 51910 697770 51950 700890
rect 48750 697730 51950 697770
rect 537269 694702 540469 694742
rect 537269 691582 537309 694702
rect 540429 691582 540469 694702
rect 537269 691542 540469 691582
rect 541069 694702 544269 694742
rect 541069 691582 541109 694702
rect 544229 691582 544269 694702
rect 541069 691542 544269 691582
rect 544869 694702 548069 694742
rect 544869 691582 544909 694702
rect 548029 691582 548069 694702
rect 544869 691542 548069 691582
rect 548669 694702 551869 694742
rect 548669 691582 548709 694702
rect 551829 691582 551869 694702
rect 548669 691542 551869 691582
<< mimcapcontact >>
rect 37390 697770 40510 700890
rect 41190 697770 44310 700890
rect 44990 697770 48110 700890
rect 48790 697770 51910 700890
rect 537309 691582 540429 694702
rect 541109 691582 544229 694702
rect 544909 691582 548029 694702
rect 548709 691582 551829 694702
<< metal4 >>
rect 16200 702200 21200 702300
rect 16200 702000 16400 702200
rect 16600 702000 16800 702200
rect 17000 702000 17200 702200
rect 17400 702000 17600 702200
rect 17800 702000 18000 702200
rect 18200 702000 18400 702200
rect 18600 702000 18800 702200
rect 19000 702000 19200 702200
rect 19400 702000 19600 702200
rect 19800 702000 20000 702200
rect 20200 702000 20400 702200
rect 20600 702000 20800 702200
rect 21000 702000 21200 702200
rect 16200 701800 21200 702000
rect 16200 701600 16400 701800
rect 16600 701600 16800 701800
rect 17000 701600 17200 701800
rect 17400 701600 17600 701800
rect 17800 701600 18000 701800
rect 18200 701600 18400 701800
rect 18600 701600 18800 701800
rect 19000 701600 19200 701800
rect 19400 701600 19600 701800
rect 19800 701600 20000 701800
rect 20200 701600 20400 701800
rect 20600 701600 20800 701800
rect 21000 701600 21200 701800
rect 16200 701400 21200 701600
rect 16200 701200 16400 701400
rect 16600 701200 16800 701400
rect 17000 701200 17200 701400
rect 17400 701200 17600 701400
rect 17800 701200 18000 701400
rect 18200 701200 18400 701400
rect 18600 701200 18800 701400
rect 19000 701200 19200 701400
rect 19400 701200 19600 701400
rect 19800 701200 20000 701400
rect 20200 701200 20400 701400
rect 20600 701200 20800 701400
rect 21000 701200 21200 701400
rect 68200 702200 73200 702300
rect 68200 702000 68400 702200
rect 68600 702000 68800 702200
rect 69000 702000 69200 702200
rect 69400 702000 69600 702200
rect 69800 702000 70000 702200
rect 70200 702000 70400 702200
rect 70600 702000 70800 702200
rect 71000 702000 71200 702200
rect 71400 702000 71600 702200
rect 71800 702000 72000 702200
rect 72200 702000 72400 702200
rect 72600 702000 72800 702200
rect 73000 702000 73200 702200
rect 68200 701800 73200 702000
rect 68200 701600 68400 701800
rect 68600 701600 68800 701800
rect 69000 701600 69200 701800
rect 69400 701600 69600 701800
rect 69800 701600 70000 701800
rect 70200 701600 70400 701800
rect 70600 701600 70800 701800
rect 71000 701600 71200 701800
rect 71400 701600 71600 701800
rect 71800 701600 72000 701800
rect 72200 701600 72400 701800
rect 72600 701600 72800 701800
rect 73000 701600 73200 701800
rect 68200 701400 73200 701600
rect 16200 701000 21200 701200
rect 16200 700800 16400 701000
rect 16600 700800 16800 701000
rect 17000 700800 17200 701000
rect 17400 700800 17600 701000
rect 17800 700800 18000 701000
rect 18200 700800 18400 701000
rect 18600 700800 18800 701000
rect 19000 700800 19200 701000
rect 19400 700800 19600 701000
rect 19800 700800 20000 701000
rect 20200 700800 20400 701000
rect 20600 700800 20800 701000
rect 21000 700800 21200 701000
rect 16200 700600 21200 700800
rect 16200 700400 16400 700600
rect 16600 700400 16800 700600
rect 17000 700400 17200 700600
rect 17400 700400 17600 700600
rect 17800 700400 18000 700600
rect 18200 700400 18400 700600
rect 18600 700400 18800 700600
rect 19000 700400 19200 700600
rect 19400 700400 19600 700600
rect 19800 700400 20000 700600
rect 20200 700400 20400 700600
rect 20600 700400 20800 700600
rect 21000 700400 21200 700600
rect 16200 700200 21200 700400
rect 16200 700000 16400 700200
rect 16600 700000 16800 700200
rect 17000 700000 17200 700200
rect 17400 700000 17600 700200
rect 17800 700000 18000 700200
rect 18200 700000 18400 700200
rect 18600 700000 18800 700200
rect 19000 700000 19200 700200
rect 19400 700000 19600 700200
rect 19800 700000 20000 700200
rect 20200 700000 20400 700200
rect 20600 700000 20800 700200
rect 21000 700000 21200 700200
rect 16200 688700 21200 700000
rect 36800 701109 52520 701260
rect 36800 701045 37278 701109
rect 40622 701045 41078 701109
rect 44422 701045 44878 701109
rect 48222 701045 48678 701109
rect 52022 701045 52520 701109
rect 36800 701020 52520 701045
rect 36800 694920 37020 701020
rect 37389 700890 40511 700891
rect 37389 697770 37390 700890
rect 40510 699550 40511 700890
rect 41189 700890 44311 700891
rect 41189 699550 41190 700890
rect 40510 699190 41190 699550
rect 40510 697770 40511 699190
rect 37389 697769 40511 697770
rect 36800 694850 36930 694920
rect 37000 694850 37020 694920
rect 36800 694810 37020 694850
rect 36800 694740 36820 694810
rect 36890 694740 37020 694810
rect 36800 694720 37020 694740
rect 40690 693960 41010 699190
rect 41189 697770 41190 699190
rect 44310 699550 44311 700890
rect 44989 700890 48111 700891
rect 44989 699550 44990 700890
rect 44310 699190 44990 699550
rect 44310 697770 44311 699190
rect 41189 697769 44311 697770
rect 44989 697770 44990 699190
rect 48110 699550 48111 700890
rect 48789 700890 51911 700891
rect 48789 699550 48790 700890
rect 48110 699190 48790 699550
rect 48110 697770 48111 699190
rect 44989 697769 48111 697770
rect 44009 695640 44281 695641
rect 44009 695370 44010 695640
rect 44280 695370 44281 695640
rect 44009 695369 44281 695370
rect 45059 695640 45331 695641
rect 45059 695370 45060 695640
rect 45330 695370 45331 695640
rect 45059 695369 45331 695370
rect 41839 695140 42091 695141
rect 41839 694890 41840 695140
rect 42090 694890 42091 695140
rect 41839 694889 42091 694890
rect 43739 695130 43991 695131
rect 43739 694880 43740 695130
rect 43990 694880 43991 695130
rect 43739 694879 43991 694880
rect 45319 695130 45571 695131
rect 45319 694880 45320 695130
rect 45570 694880 45571 695130
rect 45319 694879 45571 694880
rect 47219 695130 47471 695131
rect 47219 694880 47220 695130
rect 47470 694880 47471 695130
rect 47219 694879 47471 694880
rect 40690 693860 40710 693960
rect 40800 693860 40900 693960
rect 40990 693860 41010 693960
rect 40690 693840 41010 693860
rect 44009 694000 44281 694001
rect 44009 693730 44010 694000
rect 44280 693730 44281 694000
rect 44009 693729 44281 693730
rect 45059 694000 45331 694001
rect 45059 693730 45060 694000
rect 45330 693730 45331 694000
rect 48300 693960 48620 699190
rect 48789 697770 48790 699190
rect 51910 697770 51911 700890
rect 48789 697769 51911 697770
rect 52300 694920 52520 701020
rect 52300 694850 52320 694920
rect 52390 694850 52520 694920
rect 52300 694810 52520 694850
rect 52300 694740 52430 694810
rect 52500 694740 52520 694810
rect 52300 694720 52520 694740
rect 68200 701200 68400 701400
rect 68600 701200 68800 701400
rect 69000 701200 69200 701400
rect 69400 701200 69600 701400
rect 69800 701200 70000 701400
rect 70200 701200 70400 701400
rect 70600 701200 70800 701400
rect 71000 701200 71200 701400
rect 71400 701200 71600 701400
rect 71800 701200 72000 701400
rect 72200 701200 72400 701400
rect 72600 701200 72800 701400
rect 73000 701200 73200 701400
rect 68200 701000 73200 701200
rect 68200 700800 68400 701000
rect 68600 700800 68800 701000
rect 69000 700800 69200 701000
rect 69400 700800 69600 701000
rect 69800 700800 70000 701000
rect 70200 700800 70400 701000
rect 70600 700800 70800 701000
rect 71000 700800 71200 701000
rect 71400 700800 71600 701000
rect 71800 700800 72000 701000
rect 72200 700800 72400 701000
rect 72600 700800 72800 701000
rect 73000 700800 73200 701000
rect 68200 700600 73200 700800
rect 68200 700400 68400 700600
rect 68600 700400 68800 700600
rect 69000 700400 69200 700600
rect 69400 700400 69600 700600
rect 69800 700400 70000 700600
rect 70200 700400 70400 700600
rect 70600 700400 70800 700600
rect 71000 700400 71200 700600
rect 71400 700400 71600 700600
rect 71800 700400 72000 700600
rect 72200 700400 72400 700600
rect 72600 700400 72800 700600
rect 73000 700400 73200 700600
rect 68200 700200 73200 700400
rect 68200 700000 68400 700200
rect 68600 700000 68800 700200
rect 69000 700000 69200 700200
rect 69400 700000 69600 700200
rect 69800 700000 70000 700200
rect 70200 700000 70400 700200
rect 70600 700000 70800 700200
rect 71000 700000 71200 700200
rect 71400 700000 71600 700200
rect 71800 700000 72000 700200
rect 72200 700000 72400 700200
rect 72600 700000 72800 700200
rect 73000 700000 73200 700200
rect 48300 693860 48320 693960
rect 48410 693860 48510 693960
rect 48600 693860 48620 693960
rect 48300 693840 48620 693860
rect 45059 693729 45331 693730
rect 16200 688500 16400 688700
rect 16600 688500 16800 688700
rect 17000 688500 17200 688700
rect 17400 688500 17600 688700
rect 17800 688500 18000 688700
rect 18200 688500 18400 688700
rect 18600 688500 18800 688700
rect 19000 688500 19200 688700
rect 19400 688500 19600 688700
rect 19800 688500 20000 688700
rect 20200 688500 20400 688700
rect 20600 688500 20800 688700
rect 21000 688500 21200 688700
rect 16200 688300 21200 688500
rect 16200 688100 16400 688300
rect 16600 688100 16800 688300
rect 17000 688100 17200 688300
rect 17400 688100 17600 688300
rect 17800 688100 18000 688300
rect 18200 688100 18400 688300
rect 18600 688100 18800 688300
rect 19000 688100 19200 688300
rect 19400 688100 19600 688300
rect 19800 688100 20000 688300
rect 20200 688100 20400 688300
rect 20600 688100 20800 688300
rect 21000 688100 21200 688300
rect 16200 688000 21200 688100
rect 38670 693460 39330 693490
rect 38670 693360 38700 693460
rect 38880 693360 39120 693460
rect 39300 693360 39330 693460
rect 36600 687300 38400 687400
rect 36600 687100 36800 687300
rect 37000 687100 37200 687300
rect 37400 687100 37600 687300
rect 37800 687100 38000 687300
rect 38200 687100 38400 687300
rect 36600 685300 38400 687100
rect 36600 685100 36800 685300
rect 37000 685100 37200 685300
rect 37400 685100 37600 685300
rect 37800 685100 38000 685300
rect 38200 685100 38400 685300
rect 36600 684900 38400 685100
rect 36600 684700 36800 684900
rect 37000 684700 37200 684900
rect 37400 684700 37600 684900
rect 37800 684700 38000 684900
rect 38200 684700 38400 684900
rect 36600 684500 38400 684700
rect 36600 684300 36800 684500
rect 37000 684300 37200 684500
rect 37400 684300 37600 684500
rect 37800 684300 38000 684500
rect 38200 684300 38400 684500
rect 36600 684100 38400 684300
rect 36600 683900 36800 684100
rect 37000 683900 37200 684100
rect 37400 683900 37600 684100
rect 37800 683900 38000 684100
rect 38200 683900 38400 684100
rect 36600 683700 38400 683900
rect 36600 683500 36800 683700
rect 37000 683500 37200 683700
rect 37400 683500 37600 683700
rect 37800 683500 38000 683700
rect 38200 683500 38400 683700
rect 36600 683300 38400 683500
rect 36600 683100 36800 683300
rect 37000 683100 37200 683300
rect 37400 683100 37600 683300
rect 37800 683100 38000 683300
rect 38200 683100 38400 683300
rect 36600 682900 38400 683100
rect 36600 682700 36800 682900
rect 37000 682700 37200 682900
rect 37400 682700 37600 682900
rect 37800 682700 38000 682900
rect 38200 682700 38400 682900
rect 36600 682500 38400 682700
rect 36600 682300 36800 682500
rect 37000 682300 37200 682500
rect 37400 682300 37600 682500
rect 37800 682300 38000 682500
rect 38200 682300 38400 682500
rect 36600 682100 38400 682300
rect 36600 681900 36800 682100
rect 37000 681900 37200 682100
rect 37400 681900 37600 682100
rect 37800 681900 38000 682100
rect 38200 681900 38400 682100
rect 36600 681700 38400 681900
rect 36600 681500 36800 681700
rect 37000 681500 37200 681700
rect 37400 681500 37600 681700
rect 37800 681500 38000 681700
rect 38200 681500 38400 681700
rect 36600 681300 38400 681500
rect 36600 681100 36800 681300
rect 37000 681100 37200 681300
rect 37400 681100 37600 681300
rect 37800 681100 38000 681300
rect 38200 681100 38400 681300
rect 36600 680900 38400 681100
rect 36600 680700 36800 680900
rect 37000 680700 37200 680900
rect 37400 680700 37600 680900
rect 37800 680700 38000 680900
rect 38200 680700 38400 680900
rect 36600 680500 38400 680700
rect 36600 680300 36800 680500
rect 37000 680300 37200 680500
rect 37400 680300 37600 680500
rect 37800 680300 38000 680500
rect 38200 680300 38400 680500
rect 36600 680200 38400 680300
rect 38670 686020 39330 693360
rect 43339 693480 43601 693481
rect 43339 693220 43340 693480
rect 43600 693220 43601 693480
rect 43339 693219 43601 693220
rect 44609 693480 44871 693481
rect 44609 693220 44610 693480
rect 44870 693220 44871 693480
rect 44609 693219 44871 693220
rect 45869 693480 46131 693481
rect 45869 693220 45870 693480
rect 46130 693220 46131 693480
rect 45869 693219 46131 693220
rect 49920 693460 50580 693490
rect 49920 693360 49950 693460
rect 50130 693360 50370 693460
rect 50550 693360 50580 693460
rect 43779 692390 44041 692391
rect 43779 692130 43780 692390
rect 44040 692130 44041 692390
rect 43779 692129 44041 692130
rect 45279 692390 45541 692391
rect 45279 692130 45280 692390
rect 45540 692130 45541 692390
rect 45279 692129 45541 692130
rect 43339 691930 43601 691931
rect 43339 691670 43340 691930
rect 43600 691670 43601 691930
rect 43339 691669 43601 691670
rect 44609 691930 44871 691931
rect 44609 691670 44610 691930
rect 44870 691670 44871 691930
rect 44609 691669 44871 691670
rect 45869 691930 46131 691931
rect 45869 691670 45870 691930
rect 46130 691670 46131 691930
rect 45869 691669 46131 691670
rect 44519 689290 44781 689291
rect 44519 689030 44520 689290
rect 44780 689030 44781 689290
rect 44519 689029 44781 689030
rect 44519 687770 44781 687771
rect 44519 687510 44520 687770
rect 44780 687510 44781 687770
rect 44519 687509 44781 687510
rect 43499 686670 43751 686671
rect 43499 686420 43500 686670
rect 43750 686420 43751 686670
rect 43499 686419 43751 686420
rect 45559 686670 45811 686671
rect 45559 686420 45560 686670
rect 45810 686420 45811 686670
rect 45559 686419 45811 686420
rect 38670 685780 38700 686020
rect 38940 685780 39060 686020
rect 39300 685780 39330 686020
rect 44529 686250 44781 686251
rect 44529 686000 44530 686250
rect 44780 686000 44781 686250
rect 44529 685999 44781 686000
rect 49920 686020 50580 693360
rect 38670 685680 39330 685780
rect 38670 685440 38700 685680
rect 38940 685440 39060 685680
rect 39300 685440 39330 685680
rect 38670 675000 39330 685440
rect 49920 685780 49950 686020
rect 50190 685780 50310 686020
rect 50550 685780 50580 686020
rect 49920 685680 50580 685780
rect 49920 685440 49950 685680
rect 50190 685440 50310 685680
rect 50550 685440 50580 685680
rect 43239 685150 43491 685151
rect 43239 684900 43240 685150
rect 43490 684900 43491 685150
rect 43239 684899 43491 684900
rect 45819 685150 46071 685151
rect 45819 684900 45820 685150
rect 46070 684900 46071 685150
rect 45819 684899 46071 684900
rect 44529 684720 44781 684721
rect 44529 684470 44530 684720
rect 44780 684470 44781 684720
rect 44529 684469 44781 684470
rect 43570 683440 43750 683680
rect 45550 683440 45730 683680
rect 43570 682140 43790 683440
rect 43570 682060 43630 682140
rect 43710 682060 43790 682140
rect 43570 681920 43790 682060
rect 43570 681840 43630 681920
rect 43710 681840 43790 681920
rect 43570 681780 43790 681840
rect 43570 681700 43630 681780
rect 43710 681700 43790 681780
rect 43570 681680 43790 681700
rect 45510 682140 45730 683440
rect 45510 682060 45590 682140
rect 45670 682060 45730 682140
rect 45510 681920 45730 682060
rect 45510 681840 45590 681920
rect 45670 681840 45730 681920
rect 45510 681780 45730 681840
rect 45510 681700 45590 681780
rect 45670 681700 45730 681780
rect 45510 681680 45730 681700
rect 44130 680530 45090 680700
rect 44130 680520 44890 680530
rect 44130 680400 44270 680520
rect 44390 680410 44890 680520
rect 45010 680410 45090 680530
rect 44390 680400 45090 680410
rect 44130 679630 45090 680400
rect 44130 679540 44590 679630
rect 44680 679540 45090 679630
rect 44130 679250 45090 679540
rect 44130 679160 44580 679250
rect 44670 679160 45090 679250
rect 44130 677810 45090 679160
rect 44130 677720 44580 677810
rect 44670 677720 45090 677810
rect 32600 674000 40800 675000
rect 32600 673700 32800 674000
rect 33100 673700 33300 674000
rect 33600 673700 33800 674000
rect 34100 673700 34300 674000
rect 34600 673700 34800 674000
rect 35100 673700 35300 674000
rect 35600 673700 35800 674000
rect 36100 673700 36300 674000
rect 36600 673700 36800 674000
rect 37100 673700 37300 674000
rect 37600 673700 37800 674000
rect 38100 673700 38300 674000
rect 38600 673700 38800 674000
rect 39100 673700 39300 674000
rect 39600 673700 39800 674000
rect 40100 673700 40300 674000
rect 40600 673700 40800 674000
rect 32600 673200 40800 673700
rect 44130 674020 45090 677720
rect 44130 673780 44210 674020
rect 44450 673780 44770 674020
rect 45010 673780 45090 674020
rect 41199 673540 41441 673541
rect 41199 673300 41200 673540
rect 41440 673300 41441 673540
rect 41199 673299 41441 673300
rect 44130 673540 45090 673780
rect 49920 674000 50580 685440
rect 49920 673700 50100 674000
rect 50400 673700 50580 674000
rect 49920 673600 50580 673700
rect 44130 673300 44210 673540
rect 44450 673300 44770 673540
rect 45010 673300 45090 673540
rect 32600 672900 32800 673200
rect 33100 672900 33300 673200
rect 33600 672900 33800 673200
rect 34100 672900 34300 673200
rect 34600 672900 34800 673200
rect 35100 672900 35300 673200
rect 35600 672900 35800 673200
rect 36100 672900 36300 673200
rect 36600 672900 36800 673200
rect 37100 672900 37300 673200
rect 37600 672900 37800 673200
rect 38100 672900 38300 673200
rect 38600 672900 38800 673200
rect 39100 672900 39300 673200
rect 39600 672900 39800 673200
rect 40100 672900 40300 673200
rect 40600 672900 40800 673200
rect 32600 670700 40800 672900
rect 32600 670400 32800 670700
rect 33100 670400 33300 670700
rect 33600 670400 33800 670700
rect 34100 670400 34300 670700
rect 34600 670400 34800 670700
rect 35100 670400 35300 670700
rect 35600 670400 35800 670700
rect 36100 670400 36300 670700
rect 36600 670400 36800 670700
rect 37100 670400 37300 670700
rect 37600 670400 37800 670700
rect 38100 670400 38300 670700
rect 38600 670400 38800 670700
rect 39100 670400 39300 670700
rect 39600 670400 39800 670700
rect 40100 670400 40300 670700
rect 40600 670400 40800 670700
rect 32600 670000 40800 670400
rect 44130 673060 45090 673300
rect 47899 673540 48141 673541
rect 47899 673300 47900 673540
rect 48140 673300 48141 673540
rect 47899 673299 48141 673300
rect 49920 673300 50100 673600
rect 50400 673300 50580 673600
rect 44130 672820 44210 673060
rect 44450 672820 44770 673060
rect 45010 672820 45090 673060
rect 44130 670820 45090 672820
rect 49920 673200 50580 673300
rect 49920 672900 50100 673200
rect 50400 672900 50580 673200
rect 49920 672700 50580 672900
rect 57800 691900 62200 692200
rect 57800 691700 58000 691900
rect 58200 691700 58400 691900
rect 58600 691700 58800 691900
rect 59000 691700 59200 691900
rect 59400 691700 59600 691900
rect 59800 691700 60000 691900
rect 60200 691700 60400 691900
rect 60600 691700 60800 691900
rect 61000 691700 61200 691900
rect 61400 691700 61600 691900
rect 61800 691700 62200 691900
rect 57800 682200 62200 691700
rect 68200 690200 73200 700000
rect 534599 694992 554539 695052
rect 534599 694862 534639 694992
rect 534739 694862 534899 694992
rect 534999 694921 554129 694992
rect 534999 694862 537197 694921
rect 534599 694857 537197 694862
rect 540541 694857 540997 694921
rect 544341 694857 544797 694921
rect 548141 694857 548597 694921
rect 551941 694862 554129 694921
rect 554239 694862 554389 694992
rect 554499 694862 554539 694992
rect 551941 694857 554539 694862
rect 534599 694812 554539 694857
rect 537308 694702 540430 694703
rect 537308 691582 537309 694702
rect 540429 693552 540430 694702
rect 541108 694702 544230 694703
rect 541108 693552 541109 694702
rect 540429 693192 541109 693552
rect 540429 691582 540430 693192
rect 537308 691581 540430 691582
rect 540649 691372 540819 693192
rect 541108 691582 541109 693192
rect 544229 693552 544230 694702
rect 544908 694702 548030 694703
rect 544908 693552 544909 694702
rect 544229 693192 544909 693552
rect 544229 691582 544230 693192
rect 541108 691581 544230 691582
rect 544908 691582 544909 693192
rect 548029 693552 548030 694702
rect 548708 694702 551830 694703
rect 548708 693552 548709 694702
rect 548029 693192 548709 693552
rect 548029 691582 548030 693192
rect 544908 691581 548030 691582
rect 538849 691182 540819 691372
rect 548289 691392 548449 693192
rect 548708 691582 548709 693192
rect 551829 691582 551830 694702
rect 548708 691581 551830 691582
rect 548289 691262 549069 691392
rect 538849 690500 539139 691182
rect 541069 690682 541339 690812
rect 541069 690602 541089 690682
rect 541169 690602 541239 690682
rect 541319 690602 541339 690682
rect 68200 690000 68400 690200
rect 68600 690000 68800 690200
rect 69000 690000 69200 690200
rect 69400 690000 69600 690200
rect 69800 690000 70000 690200
rect 70200 690000 70400 690200
rect 70600 690000 70800 690200
rect 71000 690000 71200 690200
rect 71400 690000 71600 690200
rect 71800 690000 72000 690200
rect 72200 690000 72400 690200
rect 72600 690000 72800 690200
rect 73000 690000 73200 690200
rect 68200 689800 73200 690000
rect 68200 689600 68400 689800
rect 68600 689600 68800 689800
rect 69000 689600 69200 689800
rect 69400 689600 69600 689800
rect 69800 689600 70000 689800
rect 70200 689600 70400 689800
rect 70600 689600 70800 689800
rect 71000 689600 71200 689800
rect 71400 689600 71600 689800
rect 71800 689600 72000 689800
rect 72200 689600 72400 689800
rect 72600 689600 72800 689800
rect 73000 689600 73200 689800
rect 68200 689400 73200 689600
rect 532200 690400 539200 690500
rect 532200 690200 532300 690400
rect 532500 690200 532700 690400
rect 532900 690200 533100 690400
rect 533300 690200 533500 690400
rect 533700 690200 533900 690400
rect 534100 690200 539200 690400
rect 532200 690100 539200 690200
rect 532200 689900 532300 690100
rect 532500 689900 532700 690100
rect 532900 689900 533100 690100
rect 533300 689900 533500 690100
rect 533700 689900 533900 690100
rect 534100 689900 539200 690100
rect 532200 689700 539200 689900
rect 532200 689500 532300 689700
rect 532500 689500 532700 689700
rect 532900 689500 533100 689700
rect 533300 689500 533500 689700
rect 533700 689500 533900 689700
rect 534100 689500 539200 689700
rect 532200 689300 539200 689500
rect 532200 689100 532300 689300
rect 532500 689100 532700 689300
rect 532900 689100 533100 689300
rect 533300 689100 533500 689300
rect 533700 689100 533900 689300
rect 534100 689100 539200 689300
rect 532200 688900 539200 689100
rect 532200 688700 532300 688900
rect 532500 688700 532700 688900
rect 532900 688700 533100 688900
rect 533300 688700 533500 688900
rect 533700 688700 533900 688900
rect 534100 688700 539200 688900
rect 532200 688600 539200 688700
rect 541069 690142 541339 690602
rect 541069 690062 541089 690142
rect 541169 690062 541239 690142
rect 541319 690062 541339 690142
rect 541069 689602 541339 690062
rect 541069 689522 541089 689602
rect 541169 689522 541239 689602
rect 541319 689522 541339 689602
rect 538849 687652 539139 688600
rect 538849 687542 538869 687652
rect 538959 687542 539029 687652
rect 539119 687542 539139 687652
rect 538849 687322 539139 687542
rect 57800 682000 58000 682200
rect 58200 682000 58400 682200
rect 58600 682000 58800 682200
rect 59000 682000 59200 682200
rect 59400 682000 59600 682200
rect 59800 682000 60000 682200
rect 60200 682000 60400 682200
rect 60600 682000 60800 682200
rect 61000 682000 61200 682200
rect 61400 682000 61600 682200
rect 61800 682000 62200 682200
rect 44130 670580 44210 670820
rect 44450 670580 44770 670820
rect 45010 670580 45090 670820
rect 41199 670340 41441 670341
rect 41199 670100 41200 670340
rect 41440 670100 41441 670340
rect 41199 670099 41441 670100
rect 44130 670340 45090 670580
rect 44130 670100 44210 670340
rect 44450 670100 44770 670340
rect 45010 670100 45090 670340
rect 32600 669700 32800 670000
rect 33100 669700 33300 670000
rect 33600 669700 33800 670000
rect 34100 669700 34300 670000
rect 34600 669700 34800 670000
rect 35100 669700 35300 670000
rect 35600 669700 35800 670000
rect 36100 669700 36300 670000
rect 36600 669700 36800 670000
rect 37100 669700 37300 670000
rect 37600 669700 37800 670000
rect 38100 669700 38300 670000
rect 38600 669700 38800 670000
rect 39100 669700 39300 670000
rect 39600 669700 39800 670000
rect 40100 669700 40300 670000
rect 40600 669700 40800 670000
rect 32600 667400 40800 669700
rect 32600 667100 32800 667400
rect 33100 667100 33300 667400
rect 33600 667100 33800 667400
rect 34100 667100 34300 667400
rect 34600 667100 34800 667400
rect 35100 667100 35300 667400
rect 35600 667100 35800 667400
rect 36100 667100 36300 667400
rect 36600 667100 36800 667400
rect 37100 667100 37300 667400
rect 37600 667100 37800 667400
rect 38100 667100 38300 667400
rect 38600 667100 38800 667400
rect 39100 667100 39300 667400
rect 39600 667100 39800 667400
rect 40100 667100 40300 667400
rect 40600 667100 40800 667400
rect 32600 666700 40800 667100
rect 44130 669860 45090 670100
rect 47899 670340 48141 670341
rect 47899 670100 47900 670340
rect 48140 670100 48141 670340
rect 47899 670099 48141 670100
rect 44130 669620 44210 669860
rect 44450 669620 44770 669860
rect 45010 669620 45090 669860
rect 44130 667500 45090 669620
rect 44130 667260 44210 667500
rect 44450 667260 44770 667500
rect 45010 667260 45090 667500
rect 41199 667020 41441 667021
rect 41199 666780 41200 667020
rect 41440 666780 41441 667020
rect 41199 666779 41441 666780
rect 44130 667020 45090 667260
rect 44130 666780 44210 667020
rect 44450 666780 44770 667020
rect 45010 666780 45090 667020
rect 32600 666400 32800 666700
rect 33100 666400 33300 666700
rect 33600 666400 33800 666700
rect 34100 666400 34300 666700
rect 34600 666400 34800 666700
rect 35100 666400 35300 666700
rect 35600 666400 35800 666700
rect 36100 666400 36300 666700
rect 36600 666400 36800 666700
rect 37100 666400 37300 666700
rect 37600 666400 37800 666700
rect 38100 666400 38300 666700
rect 38600 666400 38800 666700
rect 39100 666400 39300 666700
rect 39600 666400 39800 666700
rect 40100 666400 40300 666700
rect 40600 666400 40800 666700
rect 32600 663300 40800 666400
rect 44130 666540 45090 666780
rect 47899 667020 48141 667021
rect 47899 666780 47900 667020
rect 48140 666780 48141 667020
rect 47899 666779 48141 666780
rect 44130 666300 44210 666540
rect 44450 666300 44770 666540
rect 45010 666300 45090 666540
rect 44130 666220 45090 666300
rect 32600 663000 32800 663300
rect 33100 663000 33300 663300
rect 33600 663000 33800 663300
rect 34100 663000 34300 663300
rect 34600 663000 34800 663300
rect 35100 663000 35300 663300
rect 35600 663000 35800 663300
rect 36100 663000 36300 663300
rect 36600 663000 36800 663300
rect 37100 663000 37300 663300
rect 37600 663000 37800 663300
rect 38100 663000 38300 663300
rect 38600 663000 38800 663300
rect 39100 663000 39300 663300
rect 39600 663000 39800 663300
rect 40100 663000 40300 663300
rect 40600 663000 40800 663300
rect 2499 648600 2801 648601
rect 2499 648300 2500 648600
rect 2800 648300 2801 648600
rect 2499 648299 2801 648300
rect 2999 648600 3301 648601
rect 2999 648300 3000 648600
rect 3300 648300 3301 648600
rect 2999 648299 3301 648300
rect 3499 648600 3801 648601
rect 3499 648300 3500 648600
rect 3800 648300 3801 648600
rect 3499 648299 3801 648300
rect 2499 648100 2801 648101
rect 2499 647800 2500 648100
rect 2800 647800 2801 648100
rect 2499 647799 2801 647800
rect 2999 648100 3301 648101
rect 2999 647800 3000 648100
rect 3300 647800 3301 648100
rect 2999 647799 3301 647800
rect 3499 648100 3801 648101
rect 3499 647800 3500 648100
rect 3800 647800 3801 648100
rect 3499 647799 3801 647800
rect 2499 647600 2801 647601
rect 2499 647300 2500 647600
rect 2800 647300 2801 647600
rect 2499 647299 2801 647300
rect 2999 647600 3301 647601
rect 2999 647300 3000 647600
rect 3300 647300 3301 647600
rect 2999 647299 3301 647300
rect 3499 647600 3801 647601
rect 3499 647300 3500 647600
rect 3800 647300 3801 647600
rect 3499 647299 3801 647300
rect 2499 647100 2801 647101
rect 2499 646800 2500 647100
rect 2800 646800 2801 647100
rect 2499 646799 2801 646800
rect 2999 647100 3301 647101
rect 2999 646800 3000 647100
rect 3300 646800 3301 647100
rect 2999 646799 3301 646800
rect 3499 647100 3801 647101
rect 3499 646800 3500 647100
rect 3800 646800 3801 647100
rect 3499 646799 3801 646800
rect 2499 646600 2801 646601
rect 2499 646300 2500 646600
rect 2800 646300 2801 646600
rect 2499 646299 2801 646300
rect 2999 646600 3301 646601
rect 2999 646300 3000 646600
rect 3300 646300 3301 646600
rect 2999 646299 3301 646300
rect 3499 646600 3801 646601
rect 3499 646300 3500 646600
rect 3800 646300 3801 646600
rect 3499 646299 3801 646300
rect 2499 646100 2801 646101
rect 2499 645800 2500 646100
rect 2800 645800 2801 646100
rect 2499 645799 2801 645800
rect 2999 646100 3301 646101
rect 2999 645800 3000 646100
rect 3300 645800 3301 646100
rect 2999 645799 3301 645800
rect 3499 646100 3801 646101
rect 3499 645800 3500 646100
rect 3800 645800 3801 646100
rect 3499 645799 3801 645800
rect 2499 645600 2801 645601
rect 2499 645300 2500 645600
rect 2800 645300 2801 645600
rect 2499 645299 2801 645300
rect 2999 645600 3301 645601
rect 2999 645300 3000 645600
rect 3300 645300 3301 645600
rect 2999 645299 3301 645300
rect 3499 645600 3801 645601
rect 3499 645300 3500 645600
rect 3800 645300 3801 645600
rect 3499 645299 3801 645300
rect 2499 645100 2801 645101
rect 2499 644800 2500 645100
rect 2800 644800 2801 645100
rect 2499 644799 2801 644800
rect 2999 645100 3301 645101
rect 2999 644800 3000 645100
rect 3300 644800 3301 645100
rect 2999 644799 3301 644800
rect 3499 645100 3801 645101
rect 3499 644800 3500 645100
rect 3800 644800 3801 645100
rect 3499 644799 3801 644800
rect 2499 644600 2801 644601
rect 2499 644300 2500 644600
rect 2800 644300 2801 644600
rect 2499 644299 2801 644300
rect 2999 644600 3301 644601
rect 2999 644300 3000 644600
rect 3300 644300 3301 644600
rect 2999 644299 3301 644300
rect 3499 644600 3801 644601
rect 3499 644300 3500 644600
rect 3800 644300 3801 644600
rect 3499 644299 3801 644300
rect 2499 644100 2801 644101
rect 2499 643800 2500 644100
rect 2800 643800 2801 644100
rect 2499 643799 2801 643800
rect 2999 644100 3301 644101
rect 2999 643800 3000 644100
rect 3300 643800 3301 644100
rect 2999 643799 3301 643800
rect 3499 644100 3801 644101
rect 3499 643800 3500 644100
rect 3800 643800 3801 644100
rect 3499 643799 3801 643800
rect 2499 643600 2801 643601
rect 2499 643300 2500 643600
rect 2800 643300 2801 643600
rect 2499 643299 2801 643300
rect 2999 643600 3301 643601
rect 2999 643300 3000 643600
rect 3300 643300 3301 643600
rect 2999 643299 3301 643300
rect 3499 643600 3801 643601
rect 3499 643300 3500 643600
rect 3800 643300 3801 643600
rect 3499 643299 3801 643300
rect 2499 643100 2801 643101
rect 2499 642800 2500 643100
rect 2800 642800 2801 643100
rect 2499 642799 2801 642800
rect 2999 643100 3301 643101
rect 2999 642800 3000 643100
rect 3300 642800 3301 643100
rect 2999 642799 3301 642800
rect 3499 643100 3801 643101
rect 3499 642800 3500 643100
rect 3800 642800 3801 643100
rect 3499 642799 3801 642800
rect 2499 642600 2801 642601
rect 2499 642300 2500 642600
rect 2800 642300 2801 642600
rect 2499 642299 2801 642300
rect 2999 642600 3301 642601
rect 2999 642300 3000 642600
rect 3300 642300 3301 642600
rect 2999 642299 3301 642300
rect 3499 642600 3801 642601
rect 3499 642300 3500 642600
rect 3800 642300 3801 642600
rect 3499 642299 3801 642300
rect 2499 642100 2801 642101
rect 2499 641800 2500 642100
rect 2800 641800 2801 642100
rect 2499 641799 2801 641800
rect 2999 642100 3301 642101
rect 2999 641800 3000 642100
rect 3300 641800 3301 642100
rect 2999 641799 3301 641800
rect 3499 642100 3801 642101
rect 3499 641800 3500 642100
rect 3800 641800 3801 642100
rect 3499 641799 3801 641800
rect 2499 641600 2801 641601
rect 2499 641300 2500 641600
rect 2800 641300 2801 641600
rect 2499 641299 2801 641300
rect 2999 641600 3301 641601
rect 2999 641300 3000 641600
rect 3300 641300 3301 641600
rect 2999 641299 3301 641300
rect 3499 641600 3801 641601
rect 3499 641300 3500 641600
rect 3800 641300 3801 641600
rect 3499 641299 3801 641300
rect 2499 641100 2801 641101
rect 2499 640800 2500 641100
rect 2800 640800 2801 641100
rect 2499 640799 2801 640800
rect 2999 641100 3301 641101
rect 2999 640800 3000 641100
rect 3300 640800 3301 641100
rect 2999 640799 3301 640800
rect 3499 641100 3801 641101
rect 3499 640800 3500 641100
rect 3800 640800 3801 641100
rect 3499 640799 3801 640800
rect 2499 640600 2801 640601
rect 2499 640300 2500 640600
rect 2800 640300 2801 640600
rect 2499 640299 2801 640300
rect 2999 640600 3301 640601
rect 2999 640300 3000 640600
rect 3300 640300 3301 640600
rect 2999 640299 3301 640300
rect 3499 640600 3801 640601
rect 3499 640300 3500 640600
rect 3800 640300 3801 640600
rect 3499 640299 3801 640300
rect 2499 640100 2801 640101
rect 2499 639800 2500 640100
rect 2800 639800 2801 640100
rect 2499 639799 2801 639800
rect 2999 640100 3301 640101
rect 2999 639800 3000 640100
rect 3300 639800 3301 640100
rect 2999 639799 3301 639800
rect 3499 640100 3801 640101
rect 3499 639800 3500 640100
rect 3800 639800 3801 640100
rect 3499 639799 3801 639800
rect 2499 639600 2801 639601
rect 2499 639300 2500 639600
rect 2800 639300 2801 639600
rect 2499 639299 2801 639300
rect 2999 639600 3301 639601
rect 2999 639300 3000 639600
rect 3300 639300 3301 639600
rect 2999 639299 3301 639300
rect 3499 639600 3801 639601
rect 3499 639300 3500 639600
rect 3800 639300 3801 639600
rect 3499 639299 3801 639300
rect 2499 639100 2801 639101
rect 2499 638800 2500 639100
rect 2800 638800 2801 639100
rect 2499 638799 2801 638800
rect 2999 639100 3301 639101
rect 2999 638800 3000 639100
rect 3300 638800 3301 639100
rect 2999 638799 3301 638800
rect 3499 639100 3801 639101
rect 3499 638800 3500 639100
rect 3800 638800 3801 639100
rect 3499 638799 3801 638800
rect 2499 638600 2801 638601
rect 2499 638300 2500 638600
rect 2800 638300 2801 638600
rect 2499 638299 2801 638300
rect 2999 638600 3301 638601
rect 2999 638300 3000 638600
rect 3300 638300 3301 638600
rect 2999 638299 3301 638300
rect 3499 638600 3801 638601
rect 3499 638300 3500 638600
rect 3800 638300 3801 638600
rect 3499 638299 3801 638300
rect 2499 638100 2801 638101
rect 2499 637800 2500 638100
rect 2800 637800 2801 638100
rect 2499 637799 2801 637800
rect 2999 638100 3301 638101
rect 2999 637800 3000 638100
rect 3300 637800 3301 638100
rect 2999 637799 3301 637800
rect 3499 638100 3801 638101
rect 3499 637800 3500 638100
rect 3800 637800 3801 638100
rect 3499 637799 3801 637800
rect 2499 637600 2801 637601
rect 2499 637300 2500 637600
rect 2800 637300 2801 637600
rect 2499 637299 2801 637300
rect 2999 637600 3301 637601
rect 2999 637300 3000 637600
rect 3300 637300 3301 637600
rect 2999 637299 3301 637300
rect 3499 637600 3801 637601
rect 3499 637300 3500 637600
rect 3800 637300 3801 637600
rect 3499 637299 3801 637300
rect 2499 637100 2801 637101
rect 2499 636800 2500 637100
rect 2800 636800 2801 637100
rect 2499 636799 2801 636800
rect 2999 637100 3301 637101
rect 2999 636800 3000 637100
rect 3300 636800 3301 637100
rect 2999 636799 3301 636800
rect 3499 637100 3801 637101
rect 3499 636800 3500 637100
rect 3800 636800 3801 637100
rect 3499 636799 3801 636800
rect 2499 636600 2801 636601
rect 2499 636300 2500 636600
rect 2800 636300 2801 636600
rect 2499 636299 2801 636300
rect 2999 636600 3301 636601
rect 2999 636300 3000 636600
rect 3300 636300 3301 636600
rect 2999 636299 3301 636300
rect 3499 636600 3801 636601
rect 3499 636300 3500 636600
rect 3800 636300 3801 636600
rect 3499 636299 3801 636300
rect 2499 636100 2801 636101
rect 2499 635800 2500 636100
rect 2800 635800 2801 636100
rect 2499 635799 2801 635800
rect 2999 636100 3301 636101
rect 2999 635800 3000 636100
rect 3300 635800 3301 636100
rect 2999 635799 3301 635800
rect 3499 636100 3801 636101
rect 3499 635800 3500 636100
rect 3800 635800 3801 636100
rect 3499 635799 3801 635800
rect 2499 635600 2801 635601
rect 2499 635300 2500 635600
rect 2800 635300 2801 635600
rect 2499 635299 2801 635300
rect 2999 635600 3301 635601
rect 2999 635300 3000 635600
rect 3300 635300 3301 635600
rect 2999 635299 3301 635300
rect 3499 635600 3801 635601
rect 3499 635300 3500 635600
rect 3800 635300 3801 635600
rect 3499 635299 3801 635300
rect 2499 635100 2801 635101
rect 2499 634800 2500 635100
rect 2800 634800 2801 635100
rect 2499 634799 2801 634800
rect 2999 635100 3301 635101
rect 2999 634800 3000 635100
rect 3300 634800 3301 635100
rect 2999 634799 3301 634800
rect 3499 635100 3801 635101
rect 3499 634800 3500 635100
rect 3800 634800 3801 635100
rect 3499 634799 3801 634800
rect 2499 634600 2801 634601
rect 2499 634300 2500 634600
rect 2800 634300 2801 634600
rect 2499 634299 2801 634300
rect 2999 634600 3301 634601
rect 2999 634300 3000 634600
rect 3300 634300 3301 634600
rect 2999 634299 3301 634300
rect 3499 634600 3801 634601
rect 3499 634300 3500 634600
rect 3800 634300 3801 634600
rect 3499 634299 3801 634300
rect 32600 564100 40800 663000
rect 57800 648600 62200 682000
rect 515500 684800 521000 685250
rect 515500 684600 515700 684800
rect 515900 684600 516100 684800
rect 516300 684600 516500 684800
rect 516700 684600 516900 684800
rect 517100 684600 517300 684800
rect 517500 684600 517700 684800
rect 517900 684600 518100 684800
rect 518300 684600 518500 684800
rect 518700 684600 518900 684800
rect 519100 684600 519300 684800
rect 519500 684600 519700 684800
rect 519900 684600 520100 684800
rect 520300 684600 520500 684800
rect 520700 684600 521000 684800
rect 515500 684400 521000 684600
rect 515500 684200 515700 684400
rect 515900 684200 516100 684400
rect 516300 684200 516500 684400
rect 516700 684200 516900 684400
rect 517100 684200 517300 684400
rect 517500 684200 517700 684400
rect 517900 684200 518100 684400
rect 518300 684200 518500 684400
rect 518700 684200 518900 684400
rect 519100 684200 519300 684400
rect 519500 684200 519700 684400
rect 519900 684200 520100 684400
rect 520300 684200 520500 684400
rect 520700 684200 521000 684400
rect 541069 684372 541339 689522
rect 543559 690682 543829 690862
rect 543559 690602 543579 690682
rect 543659 690602 543729 690682
rect 543809 690602 543829 690682
rect 543559 690142 543829 690602
rect 543559 690062 543579 690142
rect 543659 690062 543729 690142
rect 543809 690062 543829 690142
rect 543559 689602 543829 690062
rect 543559 689522 543579 689602
rect 543659 689522 543729 689602
rect 543809 689522 543829 689602
rect 542359 689002 542589 689022
rect 542359 688922 542379 689002
rect 542459 688922 542489 689002
rect 542569 688922 542589 689002
rect 542359 688392 542589 688922
rect 542359 688312 542379 688392
rect 542459 688312 542489 688392
rect 542569 688312 542589 688392
rect 542359 687880 542589 688312
rect 542350 687830 542600 687880
rect 542350 687750 542380 687830
rect 542460 687750 542500 687830
rect 542580 687750 542600 687830
rect 542350 687690 542600 687750
rect 542359 685132 542589 687690
rect 542359 685052 542379 685132
rect 542459 685052 542489 685132
rect 542569 685052 542589 685132
rect 542359 685032 542589 685052
rect 541069 684292 541089 684372
rect 541169 684292 541239 684372
rect 541319 684292 541339 684372
rect 543559 684392 543829 689522
rect 546039 690682 546309 690872
rect 546039 690602 546059 690682
rect 546139 690602 546209 690682
rect 546289 690602 546309 690682
rect 546039 690142 546309 690602
rect 546039 690062 546059 690142
rect 546139 690062 546209 690142
rect 546289 690062 546309 690142
rect 546039 689602 546309 690062
rect 546039 689522 546069 689602
rect 546149 689522 546209 689602
rect 546289 689522 546309 689602
rect 544769 689002 544999 689022
rect 544769 688922 544789 689002
rect 544869 688922 544899 689002
rect 544979 688922 544999 689002
rect 544769 688412 544999 688922
rect 544769 688332 544789 688412
rect 544869 688332 544899 688412
rect 544979 688332 544999 688412
rect 544769 687832 544999 688332
rect 544769 687752 544789 687832
rect 544869 687752 544899 687832
rect 544979 687752 544999 687832
rect 544769 685132 544999 687752
rect 544769 685052 544789 685132
rect 544869 685052 544899 685132
rect 544979 685052 544999 685132
rect 544769 685032 544999 685052
rect 543559 684312 543579 684392
rect 543659 684312 543729 684392
rect 543809 684312 543829 684392
rect 543559 684292 543829 684312
rect 546039 684392 546309 689522
rect 547229 688992 547459 689032
rect 547229 688912 547249 688992
rect 547329 688912 547359 688992
rect 547439 688912 547459 688992
rect 547229 688412 547459 688912
rect 547229 688332 547249 688412
rect 547329 688332 547359 688412
rect 547439 688332 547459 688412
rect 547229 687832 547459 688332
rect 547229 687752 547249 687832
rect 547329 687752 547359 687832
rect 547439 687752 547459 687832
rect 547229 685142 547459 687752
rect 548779 687602 549069 691262
rect 548779 687522 548799 687602
rect 548879 687522 548969 687602
rect 549049 687522 549069 687602
rect 548779 687112 549069 687522
rect 549700 687300 553100 687400
rect 549700 687200 551200 687300
rect 547229 685062 547249 685142
rect 547329 685062 547359 685142
rect 547439 685062 547459 685142
rect 547229 685042 547459 685062
rect 549700 687000 549900 687200
rect 550100 687000 550200 687200
rect 550400 687000 550500 687200
rect 550700 687000 550800 687200
rect 551000 687100 551200 687200
rect 551400 687100 553100 687300
rect 551000 687000 553100 687100
rect 549700 686800 551200 687000
rect 551400 686800 553100 687000
rect 549700 686700 553100 686800
rect 549700 686500 551200 686700
rect 551400 686500 553100 686700
rect 549700 686400 553100 686500
rect 549700 686200 551200 686400
rect 551400 686200 553100 686400
rect 549700 686100 553100 686200
rect 549700 685900 549800 686100
rect 550000 685900 550100 686100
rect 550300 685900 550400 686100
rect 550600 685900 550800 686100
rect 551000 685900 553100 686100
rect 546039 684312 546059 684392
rect 546139 684312 546199 684392
rect 546279 684312 546309 684392
rect 546039 684292 546309 684312
rect 541069 684262 541339 684292
rect 515500 684000 521000 684200
rect 515500 683800 515700 684000
rect 515900 683800 516100 684000
rect 516300 683800 516500 684000
rect 516700 683800 516900 684000
rect 517100 683800 517300 684000
rect 517500 683800 517700 684000
rect 517900 683800 518100 684000
rect 518300 683800 518500 684000
rect 518700 683800 518900 684000
rect 519100 683800 519300 684000
rect 519500 683800 519700 684000
rect 519900 683800 520100 684000
rect 520300 683800 520500 684000
rect 520700 683800 521000 684000
rect 515500 683600 521000 683800
rect 515500 683400 515700 683600
rect 515900 683400 516100 683600
rect 516300 683400 516500 683600
rect 516700 683400 516900 683600
rect 517100 683400 517300 683600
rect 517500 683400 517700 683600
rect 517900 683400 518100 683600
rect 518300 683400 518500 683600
rect 518700 683400 518900 683600
rect 519100 683400 519300 683600
rect 519500 683400 519700 683600
rect 519900 683400 520100 683600
rect 520300 683400 520500 683600
rect 520700 683400 521000 683600
rect 515500 683200 521000 683400
rect 515500 683000 515700 683200
rect 515900 683000 516100 683200
rect 516300 683000 516500 683200
rect 516700 683000 516900 683200
rect 517100 683000 517300 683200
rect 517500 683000 517700 683200
rect 517900 683000 518100 683200
rect 518300 683000 518500 683200
rect 518700 683000 518900 683200
rect 519100 683000 519300 683200
rect 519500 683000 519700 683200
rect 519900 683000 520100 683200
rect 520300 683000 520500 683200
rect 520700 683000 521000 683200
rect 515500 682800 521000 683000
rect 515500 682600 515700 682800
rect 515900 682600 516100 682800
rect 516300 682600 516500 682800
rect 516700 682600 516900 682800
rect 517100 682600 517300 682800
rect 517500 682600 517700 682800
rect 517900 682600 518100 682800
rect 518300 682600 518500 682800
rect 518700 682600 518900 682800
rect 519100 682600 519300 682800
rect 519500 682600 519700 682800
rect 519900 682600 520100 682800
rect 520300 682600 520500 682800
rect 520700 682600 521000 682800
rect 515500 679200 521000 682600
rect 546388 682442 546510 682443
rect 546388 682342 546389 682442
rect 546509 682342 546510 682442
rect 546388 682341 546510 682342
rect 515500 679000 515900 679200
rect 516100 679000 516300 679200
rect 516500 679000 516700 679200
rect 516900 679000 517100 679200
rect 517300 679000 517500 679200
rect 517700 679000 517900 679200
rect 518100 679000 518300 679200
rect 518500 679000 518700 679200
rect 518900 679000 519100 679200
rect 519300 679000 519500 679200
rect 519700 679000 519900 679200
rect 520100 679000 520300 679200
rect 520500 679000 520700 679200
rect 520900 679000 521000 679200
rect 515500 678800 521000 679000
rect 515500 678600 515900 678800
rect 516100 678600 516300 678800
rect 516500 678600 516700 678800
rect 516900 678600 517100 678800
rect 517300 678600 517500 678800
rect 517700 678600 517900 678800
rect 518100 678600 518300 678800
rect 518500 678600 518700 678800
rect 518900 678600 519100 678800
rect 519300 678600 519500 678800
rect 519700 678600 519900 678800
rect 520100 678600 520300 678800
rect 520500 678600 520700 678800
rect 520900 678600 521000 678800
rect 515500 678400 521000 678600
rect 515500 678200 515900 678400
rect 516100 678200 516300 678400
rect 516500 678200 516700 678400
rect 516900 678200 517100 678400
rect 517300 678200 517500 678400
rect 517700 678200 517900 678400
rect 518100 678200 518300 678400
rect 518500 678200 518700 678400
rect 518900 678200 519100 678400
rect 519300 678200 519500 678400
rect 519700 678200 519900 678400
rect 520100 678200 520300 678400
rect 520500 678200 520700 678400
rect 520900 678200 521000 678400
rect 515500 678000 521000 678200
rect 515500 677800 515900 678000
rect 516100 677800 516300 678000
rect 516500 677800 516700 678000
rect 516900 677800 517100 678000
rect 517300 677800 517500 678000
rect 517700 677800 517900 678000
rect 518100 677800 518300 678000
rect 518500 677800 518700 678000
rect 518900 677800 519100 678000
rect 519300 677800 519500 678000
rect 519700 677800 519900 678000
rect 520100 677800 520300 678000
rect 520500 677800 520700 678000
rect 520900 677800 521000 678000
rect 515500 677600 521000 677800
rect 515500 677400 515900 677600
rect 516100 677400 516300 677600
rect 516500 677400 516700 677600
rect 516900 677400 517100 677600
rect 517300 677400 517500 677600
rect 517700 677400 517900 677600
rect 518100 677400 518300 677600
rect 518500 677400 518700 677600
rect 518900 677400 519100 677600
rect 519300 677400 519500 677600
rect 519700 677400 519900 677600
rect 520100 677400 520300 677600
rect 520500 677400 520700 677600
rect 520900 677400 521000 677600
rect 515500 677200 521000 677400
rect 515500 677000 515900 677200
rect 516100 677000 516300 677200
rect 516500 677000 516700 677200
rect 516900 677000 517100 677200
rect 517300 677000 517500 677200
rect 517700 677000 517900 677200
rect 518100 677000 518300 677200
rect 518500 677000 518700 677200
rect 518900 677000 519100 677200
rect 519300 677000 519500 677200
rect 519700 677000 519900 677200
rect 520100 677000 520300 677200
rect 520500 677000 520700 677200
rect 520900 677000 521000 677200
rect 515500 676800 521000 677000
rect 515500 676600 515900 676800
rect 516100 676600 516300 676800
rect 516500 676600 516700 676800
rect 516900 676600 517100 676800
rect 517300 676600 517500 676800
rect 517700 676600 517900 676800
rect 518100 676600 518300 676800
rect 518500 676600 518700 676800
rect 518900 676600 519100 676800
rect 519300 676600 519500 676800
rect 519700 676600 519900 676800
rect 520100 676600 520300 676800
rect 520500 676600 520700 676800
rect 520900 676600 521000 676800
rect 515500 676460 521000 676600
rect 549700 681400 553100 685900
rect 549700 681200 549800 681400
rect 550000 681200 550200 681400
rect 550400 681200 550600 681400
rect 550800 681200 551000 681400
rect 551200 681200 551400 681400
rect 551600 681200 551800 681400
rect 552000 681200 552200 681400
rect 552400 681200 552600 681400
rect 552800 681200 553100 681400
rect 549700 681000 553100 681200
rect 549700 680800 549800 681000
rect 550000 680800 550200 681000
rect 550400 680800 550600 681000
rect 550800 680800 551000 681000
rect 551200 680800 551400 681000
rect 551600 680800 551800 681000
rect 552000 680800 552200 681000
rect 552400 680800 552600 681000
rect 552800 680800 553100 681000
rect 57800 648300 58000 648600
rect 58300 648300 58500 648600
rect 58800 648300 59000 648600
rect 59300 648300 59500 648600
rect 59800 648300 60000 648600
rect 60300 648300 60500 648600
rect 60800 648300 61000 648600
rect 61300 648300 61500 648600
rect 61800 648300 62200 648600
rect 57800 648100 62200 648300
rect 57800 647800 58000 648100
rect 58300 647800 58500 648100
rect 58800 647800 59000 648100
rect 59300 647800 59500 648100
rect 59800 647800 60000 648100
rect 60300 647800 60500 648100
rect 60800 647800 61000 648100
rect 61300 647800 61500 648100
rect 61800 647800 62200 648100
rect 57800 647600 62200 647800
rect 57800 647300 58000 647600
rect 58300 647300 58500 647600
rect 58800 647300 59000 647600
rect 59300 647300 59500 647600
rect 59800 647300 60000 647600
rect 60300 647300 60500 647600
rect 60800 647300 61000 647600
rect 61300 647300 61500 647600
rect 61800 647300 62200 647600
rect 57800 647100 62200 647300
rect 57800 646800 58000 647100
rect 58300 646800 58500 647100
rect 58800 646800 59000 647100
rect 59300 646800 59500 647100
rect 59800 646800 60000 647100
rect 60300 646800 60500 647100
rect 60800 646800 61000 647100
rect 61300 646800 61500 647100
rect 61800 646800 62200 647100
rect 57800 646600 62200 646800
rect 57800 646300 58000 646600
rect 58300 646300 58500 646600
rect 58800 646300 59000 646600
rect 59300 646300 59500 646600
rect 59800 646300 60000 646600
rect 60300 646300 60500 646600
rect 60800 646300 61000 646600
rect 61300 646300 61500 646600
rect 61800 646300 62200 646600
rect 57800 646100 62200 646300
rect 57800 645800 58000 646100
rect 58300 645800 58500 646100
rect 58800 645800 59000 646100
rect 59300 645800 59500 646100
rect 59800 645800 60000 646100
rect 60300 645800 60500 646100
rect 60800 645800 61000 646100
rect 61300 645800 61500 646100
rect 61800 645800 62200 646100
rect 57800 645600 62200 645800
rect 57800 645300 58000 645600
rect 58300 645300 58500 645600
rect 58800 645300 59000 645600
rect 59300 645300 59500 645600
rect 59800 645300 60000 645600
rect 60300 645300 60500 645600
rect 60800 645300 61000 645600
rect 61300 645300 61500 645600
rect 61800 645300 62200 645600
rect 57800 645100 62200 645300
rect 57800 644800 58000 645100
rect 58300 644800 58500 645100
rect 58800 644800 59000 645100
rect 59300 644800 59500 645100
rect 59800 644800 60000 645100
rect 60300 644800 60500 645100
rect 60800 644800 61000 645100
rect 61300 644800 61500 645100
rect 61800 644800 62200 645100
rect 57800 644600 62200 644800
rect 57800 644300 58000 644600
rect 58300 644300 58500 644600
rect 58800 644300 59000 644600
rect 59300 644300 59500 644600
rect 59800 644300 60000 644600
rect 60300 644300 60500 644600
rect 60800 644300 61000 644600
rect 61300 644300 61500 644600
rect 61800 644300 62200 644600
rect 57800 644100 62200 644300
rect 57800 643800 58000 644100
rect 58300 643800 58500 644100
rect 58800 643800 59000 644100
rect 59300 643800 59500 644100
rect 59800 643800 60000 644100
rect 60300 643800 60500 644100
rect 60800 643800 61000 644100
rect 61300 643800 61500 644100
rect 61800 643800 62200 644100
rect 57800 643600 62200 643800
rect 57800 643300 58000 643600
rect 58300 643300 58500 643600
rect 58800 643300 59000 643600
rect 59300 643300 59500 643600
rect 59800 643300 60000 643600
rect 60300 643300 60500 643600
rect 60800 643300 61000 643600
rect 61300 643300 61500 643600
rect 61800 643300 62200 643600
rect 57800 643100 62200 643300
rect 57800 642800 58000 643100
rect 58300 642800 58500 643100
rect 58800 642800 59000 643100
rect 59300 642800 59500 643100
rect 59800 642800 60000 643100
rect 60300 642800 60500 643100
rect 60800 642800 61000 643100
rect 61300 642800 61500 643100
rect 61800 642800 62200 643100
rect 57800 642600 62200 642800
rect 57800 642300 58000 642600
rect 58300 642300 58500 642600
rect 58800 642300 59000 642600
rect 59300 642300 59500 642600
rect 59800 642300 60000 642600
rect 60300 642300 60500 642600
rect 60800 642300 61000 642600
rect 61300 642300 61500 642600
rect 61800 642300 62200 642600
rect 57800 642100 62200 642300
rect 57800 641800 58000 642100
rect 58300 641800 58500 642100
rect 58800 641800 59000 642100
rect 59300 641800 59500 642100
rect 59800 641800 60000 642100
rect 60300 641800 60500 642100
rect 60800 641800 61000 642100
rect 61300 641800 61500 642100
rect 61800 641800 62200 642100
rect 57800 641600 62200 641800
rect 57800 641300 58000 641600
rect 58300 641300 58500 641600
rect 58800 641300 59000 641600
rect 59300 641300 59500 641600
rect 59800 641300 60000 641600
rect 60300 641300 60500 641600
rect 60800 641300 61000 641600
rect 61300 641300 61500 641600
rect 61800 641300 62200 641600
rect 57800 641100 62200 641300
rect 57800 640800 58000 641100
rect 58300 640800 58500 641100
rect 58800 640800 59000 641100
rect 59300 640800 59500 641100
rect 59800 640800 60000 641100
rect 60300 640800 60500 641100
rect 60800 640800 61000 641100
rect 61300 640800 61500 641100
rect 61800 640800 62200 641100
rect 57800 640600 62200 640800
rect 57800 640300 58000 640600
rect 58300 640300 58500 640600
rect 58800 640300 59000 640600
rect 59300 640300 59500 640600
rect 59800 640300 60000 640600
rect 60300 640300 60500 640600
rect 60800 640300 61000 640600
rect 61300 640300 61500 640600
rect 61800 640300 62200 640600
rect 57800 640100 62200 640300
rect 57800 639800 58000 640100
rect 58300 639800 58500 640100
rect 58800 639800 59000 640100
rect 59300 639800 59500 640100
rect 59800 639800 60000 640100
rect 60300 639800 60500 640100
rect 60800 639800 61000 640100
rect 61300 639800 61500 640100
rect 61800 639800 62200 640100
rect 57800 639600 62200 639800
rect 57800 639300 58000 639600
rect 58300 639300 58500 639600
rect 58800 639300 59000 639600
rect 59300 639300 59500 639600
rect 59800 639300 60000 639600
rect 60300 639300 60500 639600
rect 60800 639300 61000 639600
rect 61300 639300 61500 639600
rect 61800 639300 62200 639600
rect 57800 639100 62200 639300
rect 57800 638800 58000 639100
rect 58300 638800 58500 639100
rect 58800 638800 59000 639100
rect 59300 638800 59500 639100
rect 59800 638800 60000 639100
rect 60300 638800 60500 639100
rect 60800 638800 61000 639100
rect 61300 638800 61500 639100
rect 61800 638800 62200 639100
rect 57800 638600 62200 638800
rect 57800 638300 58000 638600
rect 58300 638300 58500 638600
rect 58800 638300 59000 638600
rect 59300 638300 59500 638600
rect 59800 638300 60000 638600
rect 60300 638300 60500 638600
rect 60800 638300 61000 638600
rect 61300 638300 61500 638600
rect 61800 638300 62200 638600
rect 57800 638100 62200 638300
rect 57800 637800 58000 638100
rect 58300 637800 58500 638100
rect 58800 637800 59000 638100
rect 59300 637800 59500 638100
rect 59800 637800 60000 638100
rect 60300 637800 60500 638100
rect 60800 637800 61000 638100
rect 61300 637800 61500 638100
rect 61800 637800 62200 638100
rect 57800 637600 62200 637800
rect 57800 637300 58000 637600
rect 58300 637300 58500 637600
rect 58800 637300 59000 637600
rect 59300 637300 59500 637600
rect 59800 637300 60000 637600
rect 60300 637300 60500 637600
rect 60800 637300 61000 637600
rect 61300 637300 61500 637600
rect 61800 637300 62200 637600
rect 57800 637100 62200 637300
rect 57800 636800 58000 637100
rect 58300 636800 58500 637100
rect 58800 636800 59000 637100
rect 59300 636800 59500 637100
rect 59800 636800 60000 637100
rect 60300 636800 60500 637100
rect 60800 636800 61000 637100
rect 61300 636800 61500 637100
rect 61800 636800 62200 637100
rect 57800 636600 62200 636800
rect 57800 636300 58000 636600
rect 58300 636300 58500 636600
rect 58800 636300 59000 636600
rect 59300 636300 59500 636600
rect 59800 636300 60000 636600
rect 60300 636300 60500 636600
rect 60800 636300 61000 636600
rect 61300 636300 61500 636600
rect 61800 636300 62200 636600
rect 57800 636100 62200 636300
rect 57800 635800 58000 636100
rect 58300 635800 58500 636100
rect 58800 635800 59000 636100
rect 59300 635800 59500 636100
rect 59800 635800 60000 636100
rect 60300 635800 60500 636100
rect 60800 635800 61000 636100
rect 61300 635800 61500 636100
rect 61800 635800 62200 636100
rect 57800 635600 62200 635800
rect 57800 635300 58000 635600
rect 58300 635300 58500 635600
rect 58800 635300 59000 635600
rect 59300 635300 59500 635600
rect 59800 635300 60000 635600
rect 60300 635300 60500 635600
rect 60800 635300 61000 635600
rect 61300 635300 61500 635600
rect 61800 635300 62200 635600
rect 57800 635100 62200 635300
rect 57800 634800 58000 635100
rect 58300 634800 58500 635100
rect 58800 634800 59000 635100
rect 59300 634800 59500 635100
rect 59800 634800 60000 635100
rect 60300 634800 60500 635100
rect 60800 634800 61000 635100
rect 61300 634800 61500 635100
rect 61800 634800 62200 635100
rect 57800 634600 62200 634800
rect 57800 634300 58000 634600
rect 58300 634300 58500 634600
rect 58800 634300 59000 634600
rect 59300 634300 59500 634600
rect 59800 634300 60000 634600
rect 60300 634300 60500 634600
rect 60800 634300 61000 634600
rect 61300 634300 61500 634600
rect 61800 634300 62200 634600
rect 57800 633800 62200 634300
rect 549700 644600 553100 680800
rect 549700 644400 550000 644600
rect 550200 644400 550400 644600
rect 550600 644400 550800 644600
rect 551000 644400 551200 644600
rect 551400 644400 551600 644600
rect 551800 644400 552000 644600
rect 552200 644400 552400 644600
rect 552600 644400 552800 644600
rect 553000 644400 553100 644600
rect 549700 644200 553100 644400
rect 549700 644000 550000 644200
rect 550200 644000 550400 644200
rect 550600 644000 550800 644200
rect 551000 644000 551200 644200
rect 551400 644000 551600 644200
rect 551800 644000 552000 644200
rect 552200 644000 552400 644200
rect 552600 644000 552800 644200
rect 553000 644000 553100 644200
rect 549700 643800 553100 644000
rect 549700 643600 550000 643800
rect 550200 643600 550400 643800
rect 550600 643600 550800 643800
rect 551000 643600 551200 643800
rect 551400 643600 551600 643800
rect 551800 643600 552000 643800
rect 552200 643600 552400 643800
rect 552600 643600 552800 643800
rect 553000 643600 553100 643800
rect 549700 643400 553100 643600
rect 549700 643200 550000 643400
rect 550200 643200 550400 643400
rect 550600 643200 550800 643400
rect 551000 643200 551200 643400
rect 551400 643200 551600 643400
rect 551800 643200 552000 643400
rect 552200 643200 552400 643400
rect 552600 643200 552800 643400
rect 553000 643200 553100 643400
rect 549700 643000 553100 643200
rect 549700 642800 550000 643000
rect 550200 642800 550400 643000
rect 550600 642800 550800 643000
rect 551000 642800 551200 643000
rect 551400 642800 551600 643000
rect 551800 642800 552000 643000
rect 552200 642800 552400 643000
rect 552600 642800 552800 643000
rect 553000 642800 553100 643000
rect 549700 642600 553100 642800
rect 549700 642400 550000 642600
rect 550200 642400 550400 642600
rect 550600 642400 550800 642600
rect 551000 642400 551200 642600
rect 551400 642400 551600 642600
rect 551800 642400 552000 642600
rect 552200 642400 552400 642600
rect 552600 642400 552800 642600
rect 553000 642400 553100 642600
rect 549700 642200 553100 642400
rect 549700 642000 550000 642200
rect 550200 642000 550400 642200
rect 550600 642000 550800 642200
rect 551000 642000 551200 642200
rect 551400 642000 551600 642200
rect 551800 642000 552000 642200
rect 552200 642000 552400 642200
rect 552600 642000 552800 642200
rect 553000 642000 553100 642200
rect 549700 641800 553100 642000
rect 549700 641600 550000 641800
rect 550200 641600 550400 641800
rect 550600 641600 550800 641800
rect 551000 641600 551200 641800
rect 551400 641600 551600 641800
rect 551800 641600 552000 641800
rect 552200 641600 552400 641800
rect 552600 641600 552800 641800
rect 553000 641600 553100 641800
rect 549700 641400 553100 641600
rect 549700 641200 550000 641400
rect 550200 641200 550400 641400
rect 550600 641200 550800 641400
rect 551000 641200 551200 641400
rect 551400 641200 551600 641400
rect 551800 641200 552000 641400
rect 552200 641200 552400 641400
rect 552600 641200 552800 641400
rect 553000 641200 553100 641400
rect 549700 641000 553100 641200
rect 549700 640800 550000 641000
rect 550200 640800 550400 641000
rect 550600 640800 550800 641000
rect 551000 640800 551200 641000
rect 551400 640800 551600 641000
rect 551800 640800 552000 641000
rect 552200 640800 552400 641000
rect 552600 640800 552800 641000
rect 553000 640800 553100 641000
rect 549700 640600 553100 640800
rect 549700 640400 550000 640600
rect 550200 640400 550400 640600
rect 550600 640400 550800 640600
rect 551000 640400 551200 640600
rect 551400 640400 551600 640600
rect 551800 640400 552000 640600
rect 552200 640400 552400 640600
rect 552600 640400 552800 640600
rect 553000 640400 553100 640600
rect 549700 640200 553100 640400
rect 549700 640000 550000 640200
rect 550200 640000 550400 640200
rect 550600 640000 550800 640200
rect 551000 640000 551200 640200
rect 551400 640000 551600 640200
rect 551800 640000 552000 640200
rect 552200 640000 552400 640200
rect 552600 640000 552800 640200
rect 553000 640000 553100 640200
rect 549700 639800 553100 640000
rect 549700 639600 550000 639800
rect 550200 639600 550400 639800
rect 550600 639600 550800 639800
rect 551000 639600 551200 639800
rect 551400 639600 551600 639800
rect 551800 639600 552000 639800
rect 552200 639600 552400 639800
rect 552600 639600 552800 639800
rect 553000 639600 553100 639800
rect 549700 639400 553100 639600
rect 549700 639200 550000 639400
rect 550200 639200 550400 639400
rect 550600 639200 550800 639400
rect 551000 639200 551200 639400
rect 551400 639200 551600 639400
rect 551800 639200 552000 639400
rect 552200 639200 552400 639400
rect 552600 639200 552800 639400
rect 553000 639200 553100 639400
rect 549700 639000 553100 639200
rect 549700 638800 550000 639000
rect 550200 638800 550400 639000
rect 550600 638800 550800 639000
rect 551000 638800 551200 639000
rect 551400 638800 551600 639000
rect 551800 638800 552000 639000
rect 552200 638800 552400 639000
rect 552600 638800 552800 639000
rect 553000 638800 553100 639000
rect 549700 638600 553100 638800
rect 549700 638400 550000 638600
rect 550200 638400 550400 638600
rect 550600 638400 550800 638600
rect 551000 638400 551200 638600
rect 551400 638400 551600 638600
rect 551800 638400 552000 638600
rect 552200 638400 552400 638600
rect 552600 638400 552800 638600
rect 553000 638400 553100 638600
rect 549700 638200 553100 638400
rect 549700 638000 550000 638200
rect 550200 638000 550400 638200
rect 550600 638000 550800 638200
rect 551000 638000 551200 638200
rect 551400 638000 551600 638200
rect 551800 638000 552000 638200
rect 552200 638000 552400 638200
rect 552600 638000 552800 638200
rect 553000 638000 553100 638200
rect 549700 637800 553100 638000
rect 549700 637600 550000 637800
rect 550200 637600 550400 637800
rect 550600 637600 550800 637800
rect 551000 637600 551200 637800
rect 551400 637600 551600 637800
rect 551800 637600 552000 637800
rect 552200 637600 552400 637800
rect 552600 637600 552800 637800
rect 553000 637600 553100 637800
rect 549700 637400 553100 637600
rect 549700 637200 550000 637400
rect 550200 637200 550400 637400
rect 550600 637200 550800 637400
rect 551000 637200 551200 637400
rect 551400 637200 551600 637400
rect 551800 637200 552000 637400
rect 552200 637200 552400 637400
rect 552600 637200 552800 637400
rect 553000 637200 553100 637400
rect 549700 637000 553100 637200
rect 549700 636800 550000 637000
rect 550200 636800 550400 637000
rect 550600 636800 550800 637000
rect 551000 636800 551200 637000
rect 551400 636800 551600 637000
rect 551800 636800 552000 637000
rect 552200 636800 552400 637000
rect 552600 636800 552800 637000
rect 553000 636800 553100 637000
rect 549700 636600 553100 636800
rect 549700 636400 550000 636600
rect 550200 636400 550400 636600
rect 550600 636400 550800 636600
rect 551000 636400 551200 636600
rect 551400 636400 551600 636600
rect 551800 636400 552000 636600
rect 552200 636400 552400 636600
rect 552600 636400 552800 636600
rect 553000 636400 553100 636600
rect 549700 636200 553100 636400
rect 549700 636000 550000 636200
rect 550200 636000 550400 636200
rect 550600 636000 550800 636200
rect 551000 636000 551200 636200
rect 551400 636000 551600 636200
rect 551800 636000 552000 636200
rect 552200 636000 552400 636200
rect 552600 636000 552800 636200
rect 553000 636000 553100 636200
rect 549700 635800 553100 636000
rect 549700 635600 550000 635800
rect 550200 635600 550400 635800
rect 550600 635600 550800 635800
rect 551000 635600 551200 635800
rect 551400 635600 551600 635800
rect 551800 635600 552000 635800
rect 552200 635600 552400 635800
rect 552600 635600 552800 635800
rect 553000 635600 553100 635800
rect 549700 635400 553100 635600
rect 549700 635200 550000 635400
rect 550200 635200 550400 635400
rect 550600 635200 550800 635400
rect 551000 635200 551200 635400
rect 551400 635200 551600 635400
rect 551800 635200 552000 635400
rect 552200 635200 552400 635400
rect 552600 635200 552800 635400
rect 553000 635200 553100 635400
rect 549700 635000 553100 635200
rect 549700 634800 550000 635000
rect 550200 634800 550400 635000
rect 550600 634800 550800 635000
rect 551000 634800 551200 635000
rect 551400 634800 551600 635000
rect 551800 634800 552000 635000
rect 552200 634800 552400 635000
rect 552600 634800 552800 635000
rect 553000 634800 553100 635000
rect 549700 634600 553100 634800
rect 549700 634400 550000 634600
rect 550200 634400 550400 634600
rect 550600 634400 550800 634600
rect 551000 634400 551200 634600
rect 551400 634400 551600 634600
rect 551800 634400 552000 634600
rect 552200 634400 552400 634600
rect 552600 634400 552800 634600
rect 553000 634400 553100 634600
rect 549700 634200 553100 634400
rect 549700 634000 550000 634200
rect 550200 634000 550400 634200
rect 550600 634000 550800 634200
rect 551000 634000 551200 634200
rect 551400 634000 551600 634200
rect 551800 634000 552000 634200
rect 552200 634000 552400 634200
rect 552600 634000 552800 634200
rect 553000 634000 553100 634200
rect 549700 633800 553100 634000
rect 549700 633600 550000 633800
rect 550200 633600 550400 633800
rect 550600 633600 550800 633800
rect 551000 633600 551200 633800
rect 551400 633600 551600 633800
rect 551800 633600 552000 633800
rect 552200 633600 552400 633800
rect 552600 633600 552800 633800
rect 553000 633600 553100 633800
rect 549700 633400 553100 633600
rect 549700 633200 550000 633400
rect 550200 633200 550400 633400
rect 550600 633200 550800 633400
rect 551000 633200 551200 633400
rect 551400 633200 551600 633400
rect 551800 633200 552000 633400
rect 552200 633200 552400 633400
rect 552600 633200 552800 633400
rect 553000 633200 553100 633400
rect 549700 633000 553100 633200
rect 549700 632800 550000 633000
rect 550200 632800 550400 633000
rect 550600 632800 550800 633000
rect 551000 632800 551200 633000
rect 551400 632800 551600 633000
rect 551800 632800 552000 633000
rect 552200 632800 552400 633000
rect 552600 632800 552800 633000
rect 553000 632800 553100 633000
rect 549700 632600 553100 632800
rect 549700 632400 550000 632600
rect 550200 632400 550400 632600
rect 550600 632400 550800 632600
rect 551000 632400 551200 632600
rect 551400 632400 551600 632600
rect 551800 632400 552000 632600
rect 552200 632400 552400 632600
rect 552600 632400 552800 632600
rect 553000 632400 553100 632600
rect 549700 632200 553100 632400
rect 549700 632000 550000 632200
rect 550200 632000 550400 632200
rect 550600 632000 550800 632200
rect 551000 632000 551200 632200
rect 551400 632000 551600 632200
rect 551800 632000 552000 632200
rect 552200 632000 552400 632200
rect 552600 632000 552800 632200
rect 553000 632000 553100 632200
rect 549700 631800 553100 632000
rect 549700 631600 550000 631800
rect 550200 631600 550400 631800
rect 550600 631600 550800 631800
rect 551000 631600 551200 631800
rect 551400 631600 551600 631800
rect 551800 631600 552000 631800
rect 552200 631600 552400 631800
rect 552600 631600 552800 631800
rect 553000 631600 553100 631800
rect 549700 631400 553100 631600
rect 549700 631200 550000 631400
rect 550200 631200 550400 631400
rect 550600 631200 550800 631400
rect 551000 631200 551200 631400
rect 551400 631200 551600 631400
rect 551800 631200 552000 631400
rect 552200 631200 552400 631400
rect 552600 631200 552800 631400
rect 553000 631200 553100 631400
rect 549700 631000 553100 631200
rect 549700 630800 550000 631000
rect 550200 630800 550400 631000
rect 550600 630800 550800 631000
rect 551000 630800 551200 631000
rect 551400 630800 551600 631000
rect 551800 630800 552000 631000
rect 552200 630800 552400 631000
rect 552600 630800 552800 631000
rect 553000 630800 553100 631000
rect 549700 630700 553100 630800
rect 549700 630500 550000 630700
rect 550200 630500 550400 630700
rect 550600 630500 550800 630700
rect 551000 630500 551200 630700
rect 551400 630500 551600 630700
rect 551800 630500 552000 630700
rect 552200 630500 552400 630700
rect 552600 630500 552800 630700
rect 553000 630500 553100 630700
rect 549700 630400 553100 630500
rect 549700 630200 550000 630400
rect 550200 630200 550400 630400
rect 550600 630200 550800 630400
rect 551000 630200 551200 630400
rect 551400 630200 551600 630400
rect 551800 630200 552000 630400
rect 552200 630200 552400 630400
rect 552600 630200 552800 630400
rect 553000 630200 553100 630400
rect 549700 630000 553100 630200
rect 549700 629800 550000 630000
rect 550200 629800 550400 630000
rect 550600 629800 550800 630000
rect 551000 629800 551200 630000
rect 551400 629800 551600 630000
rect 551800 629800 552000 630000
rect 552200 629800 552400 630000
rect 552600 629800 552800 630000
rect 553000 629800 553100 630000
rect 549700 629700 553100 629800
rect 32600 563900 32800 564100
rect 33000 563900 33200 564100
rect 33400 563900 33600 564100
rect 33800 563900 34000 564100
rect 34200 563900 34400 564100
rect 34600 563900 34800 564100
rect 35000 563900 35200 564100
rect 35400 563900 35600 564100
rect 35800 563900 36000 564100
rect 36200 563900 36400 564100
rect 36600 563900 36800 564100
rect 37000 563900 37200 564100
rect 37400 563900 37600 564100
rect 37800 563900 38000 564100
rect 38200 563900 38400 564100
rect 38600 563900 38800 564100
rect 39000 563900 39200 564100
rect 39400 563900 39600 564100
rect 39800 563900 40000 564100
rect 40200 563900 40400 564100
rect 40600 563900 40800 564100
rect 32600 563700 40800 563900
rect 32600 563500 32800 563700
rect 33000 563500 33200 563700
rect 33400 563500 33600 563700
rect 33800 563500 34000 563700
rect 34200 563500 34400 563700
rect 34600 563500 34800 563700
rect 35000 563500 35200 563700
rect 35400 563500 35600 563700
rect 35800 563500 36000 563700
rect 36200 563500 36400 563700
rect 36600 563500 36800 563700
rect 37000 563500 37200 563700
rect 37400 563500 37600 563700
rect 37800 563500 38000 563700
rect 38200 563500 38400 563700
rect 38600 563500 38800 563700
rect 39000 563500 39200 563700
rect 39400 563500 39600 563700
rect 39800 563500 40000 563700
rect 40200 563500 40400 563700
rect 40600 563500 40800 563700
rect 32600 563300 40800 563500
rect 32600 563100 32800 563300
rect 33000 563100 33200 563300
rect 33400 563100 33600 563300
rect 33800 563100 34000 563300
rect 34200 563100 34400 563300
rect 34600 563100 34800 563300
rect 35000 563100 35200 563300
rect 35400 563100 35600 563300
rect 35800 563100 36000 563300
rect 36200 563100 36400 563300
rect 36600 563100 36800 563300
rect 37000 563100 37200 563300
rect 37400 563100 37600 563300
rect 37800 563100 38000 563300
rect 38200 563100 38400 563300
rect 38600 563100 38800 563300
rect 39000 563100 39200 563300
rect 39400 563100 39600 563300
rect 39800 563100 40000 563300
rect 40200 563100 40400 563300
rect 40600 563100 40800 563300
rect 32600 562900 40800 563100
rect 32600 562700 32800 562900
rect 33000 562700 33200 562900
rect 33400 562700 33600 562900
rect 33800 562700 34000 562900
rect 34200 562700 34400 562900
rect 34600 562700 34800 562900
rect 35000 562700 35200 562900
rect 35400 562700 35600 562900
rect 35800 562700 36000 562900
rect 36200 562700 36400 562900
rect 36600 562700 36800 562900
rect 37000 562700 37200 562900
rect 37400 562700 37600 562900
rect 37800 562700 38000 562900
rect 38200 562700 38400 562900
rect 38600 562700 38800 562900
rect 39000 562700 39200 562900
rect 39400 562700 39600 562900
rect 39800 562700 40000 562900
rect 40200 562700 40400 562900
rect 40600 562700 40800 562900
rect 32600 562500 40800 562700
rect 32600 562300 32800 562500
rect 33000 562300 33200 562500
rect 33400 562300 33600 562500
rect 33800 562300 34000 562500
rect 34200 562300 34400 562500
rect 34600 562300 34800 562500
rect 35000 562300 35200 562500
rect 35400 562300 35600 562500
rect 35800 562300 36000 562500
rect 36200 562300 36400 562500
rect 36600 562300 36800 562500
rect 37000 562300 37200 562500
rect 37400 562300 37600 562500
rect 37800 562300 38000 562500
rect 38200 562300 38400 562500
rect 38600 562300 38800 562500
rect 39000 562300 39200 562500
rect 39400 562300 39600 562500
rect 39800 562300 40000 562500
rect 40200 562300 40400 562500
rect 40600 562300 40800 562500
rect 32600 562100 40800 562300
rect 32600 561900 32800 562100
rect 33000 561900 33200 562100
rect 33400 561900 33600 562100
rect 33800 561900 34000 562100
rect 34200 561900 34400 562100
rect 34600 561900 34800 562100
rect 35000 561900 35200 562100
rect 35400 561900 35600 562100
rect 35800 561900 36000 562100
rect 36200 561900 36400 562100
rect 36600 561900 36800 562100
rect 37000 561900 37200 562100
rect 37400 561900 37600 562100
rect 37800 561900 38000 562100
rect 38200 561900 38400 562100
rect 38600 561900 38800 562100
rect 39000 561900 39200 562100
rect 39400 561900 39600 562100
rect 39800 561900 40000 562100
rect 40200 561900 40400 562100
rect 40600 561900 40800 562100
rect 32600 561700 40800 561900
rect 32600 561500 32800 561700
rect 33000 561500 33200 561700
rect 33400 561500 33600 561700
rect 33800 561500 34000 561700
rect 34200 561500 34400 561700
rect 34600 561500 34800 561700
rect 35000 561500 35200 561700
rect 35400 561500 35600 561700
rect 35800 561500 36000 561700
rect 36200 561500 36400 561700
rect 36600 561500 36800 561700
rect 37000 561500 37200 561700
rect 37400 561500 37600 561700
rect 37800 561500 38000 561700
rect 38200 561500 38400 561700
rect 38600 561500 38800 561700
rect 39000 561500 39200 561700
rect 39400 561500 39600 561700
rect 39800 561500 40000 561700
rect 40200 561500 40400 561700
rect 40600 561500 40800 561700
rect 32600 561300 40800 561500
rect 32600 561100 32800 561300
rect 33000 561100 33200 561300
rect 33400 561100 33600 561300
rect 33800 561100 34000 561300
rect 34200 561100 34400 561300
rect 34600 561100 34800 561300
rect 35000 561100 35200 561300
rect 35400 561100 35600 561300
rect 35800 561100 36000 561300
rect 36200 561100 36400 561300
rect 36600 561100 36800 561300
rect 37000 561100 37200 561300
rect 37400 561100 37600 561300
rect 37800 561100 38000 561300
rect 38200 561100 38400 561300
rect 38600 561100 38800 561300
rect 39000 561100 39200 561300
rect 39400 561100 39600 561300
rect 39800 561100 40000 561300
rect 40200 561100 40400 561300
rect 40600 561100 40800 561300
rect 32600 560900 40800 561100
rect 32600 560700 32800 560900
rect 33000 560700 33200 560900
rect 33400 560700 33600 560900
rect 33800 560700 34000 560900
rect 34200 560700 34400 560900
rect 34600 560700 34800 560900
rect 35000 560700 35200 560900
rect 35400 560700 35600 560900
rect 35800 560700 36000 560900
rect 36200 560700 36400 560900
rect 36600 560700 36800 560900
rect 37000 560700 37200 560900
rect 37400 560700 37600 560900
rect 37800 560700 38000 560900
rect 38200 560700 38400 560900
rect 38600 560700 38800 560900
rect 39000 560700 39200 560900
rect 39400 560700 39600 560900
rect 39800 560700 40000 560900
rect 40200 560700 40400 560900
rect 40600 560700 40800 560900
rect 32600 560500 40800 560700
rect 32600 560300 32800 560500
rect 33000 560300 33200 560500
rect 33400 560300 33600 560500
rect 33800 560300 34000 560500
rect 34200 560300 34400 560500
rect 34600 560300 34800 560500
rect 35000 560300 35200 560500
rect 35400 560300 35600 560500
rect 35800 560300 36000 560500
rect 36200 560300 36400 560500
rect 36600 560300 36800 560500
rect 37000 560300 37200 560500
rect 37400 560300 37600 560500
rect 37800 560300 38000 560500
rect 38200 560300 38400 560500
rect 38600 560300 38800 560500
rect 39000 560300 39200 560500
rect 39400 560300 39600 560500
rect 39800 560300 40000 560500
rect 40200 560300 40400 560500
rect 40600 560300 40800 560500
rect 32600 560100 40800 560300
rect 32600 559900 32800 560100
rect 33000 559900 33200 560100
rect 33400 559900 33600 560100
rect 33800 559900 34000 560100
rect 34200 559900 34400 560100
rect 34600 559900 34800 560100
rect 35000 559900 35200 560100
rect 35400 559900 35600 560100
rect 35800 559900 36000 560100
rect 36200 559900 36400 560100
rect 36600 559900 36800 560100
rect 37000 559900 37200 560100
rect 37400 559900 37600 560100
rect 37800 559900 38000 560100
rect 38200 559900 38400 560100
rect 38600 559900 38800 560100
rect 39000 559900 39200 560100
rect 39400 559900 39600 560100
rect 39800 559900 40000 560100
rect 40200 559900 40400 560100
rect 40600 559900 40800 560100
rect 32600 559700 40800 559900
rect 32600 559500 32800 559700
rect 33000 559500 33200 559700
rect 33400 559500 33600 559700
rect 33800 559500 34000 559700
rect 34200 559500 34400 559700
rect 34600 559500 34800 559700
rect 35000 559500 35200 559700
rect 35400 559500 35600 559700
rect 35800 559500 36000 559700
rect 36200 559500 36400 559700
rect 36600 559500 36800 559700
rect 37000 559500 37200 559700
rect 37400 559500 37600 559700
rect 37800 559500 38000 559700
rect 38200 559500 38400 559700
rect 38600 559500 38800 559700
rect 39000 559500 39200 559700
rect 39400 559500 39600 559700
rect 39800 559500 40000 559700
rect 40200 559500 40400 559700
rect 40600 559500 40800 559700
rect 32600 559300 40800 559500
rect 32600 559100 32800 559300
rect 33000 559100 33200 559300
rect 33400 559100 33600 559300
rect 33800 559100 34000 559300
rect 34200 559100 34400 559300
rect 34600 559100 34800 559300
rect 35000 559100 35200 559300
rect 35400 559100 35600 559300
rect 35800 559100 36000 559300
rect 36200 559100 36400 559300
rect 36600 559100 36800 559300
rect 37000 559100 37200 559300
rect 37400 559100 37600 559300
rect 37800 559100 38000 559300
rect 38200 559100 38400 559300
rect 38600 559100 38800 559300
rect 39000 559100 39200 559300
rect 39400 559100 39600 559300
rect 39800 559100 40000 559300
rect 40200 559100 40400 559300
rect 40600 559100 40800 559300
rect 32600 558900 40800 559100
rect 32600 558700 32800 558900
rect 33000 558700 33200 558900
rect 33400 558700 33600 558900
rect 33800 558700 34000 558900
rect 34200 558700 34400 558900
rect 34600 558700 34800 558900
rect 35000 558700 35200 558900
rect 35400 558700 35600 558900
rect 35800 558700 36000 558900
rect 36200 558700 36400 558900
rect 36600 558700 36800 558900
rect 37000 558700 37200 558900
rect 37400 558700 37600 558900
rect 37800 558700 38000 558900
rect 38200 558700 38400 558900
rect 38600 558700 38800 558900
rect 39000 558700 39200 558900
rect 39400 558700 39600 558900
rect 39800 558700 40000 558900
rect 40200 558700 40400 558900
rect 40600 558700 40800 558900
rect 32600 558500 40800 558700
rect 32600 558300 32800 558500
rect 33000 558300 33200 558500
rect 33400 558300 33600 558500
rect 33800 558300 34000 558500
rect 34200 558300 34400 558500
rect 34600 558300 34800 558500
rect 35000 558300 35200 558500
rect 35400 558300 35600 558500
rect 35800 558300 36000 558500
rect 36200 558300 36400 558500
rect 36600 558300 36800 558500
rect 37000 558300 37200 558500
rect 37400 558300 37600 558500
rect 37800 558300 38000 558500
rect 38200 558300 38400 558500
rect 38600 558300 38800 558500
rect 39000 558300 39200 558500
rect 39400 558300 39600 558500
rect 39800 558300 40000 558500
rect 40200 558300 40400 558500
rect 40600 558300 40800 558500
rect 32600 558100 40800 558300
rect 32600 557900 32800 558100
rect 33000 557900 33200 558100
rect 33400 557900 33600 558100
rect 33800 557900 34000 558100
rect 34200 557900 34400 558100
rect 34600 557900 34800 558100
rect 35000 557900 35200 558100
rect 35400 557900 35600 558100
rect 35800 557900 36000 558100
rect 36200 557900 36400 558100
rect 36600 557900 36800 558100
rect 37000 557900 37200 558100
rect 37400 557900 37600 558100
rect 37800 557900 38000 558100
rect 38200 557900 38400 558100
rect 38600 557900 38800 558100
rect 39000 557900 39200 558100
rect 39400 557900 39600 558100
rect 39800 557900 40000 558100
rect 40200 557900 40400 558100
rect 40600 557900 40800 558100
rect 32600 557700 40800 557900
rect 32600 557500 32800 557700
rect 33000 557500 33200 557700
rect 33400 557500 33600 557700
rect 33800 557500 34000 557700
rect 34200 557500 34400 557700
rect 34600 557500 34800 557700
rect 35000 557500 35200 557700
rect 35400 557500 35600 557700
rect 35800 557500 36000 557700
rect 36200 557500 36400 557700
rect 36600 557500 36800 557700
rect 37000 557500 37200 557700
rect 37400 557500 37600 557700
rect 37800 557500 38000 557700
rect 38200 557500 38400 557700
rect 38600 557500 38800 557700
rect 39000 557500 39200 557700
rect 39400 557500 39600 557700
rect 39800 557500 40000 557700
rect 40200 557500 40400 557700
rect 40600 557500 40800 557700
rect 32600 557300 40800 557500
rect 32600 557100 32800 557300
rect 33000 557100 33200 557300
rect 33400 557100 33600 557300
rect 33800 557100 34000 557300
rect 34200 557100 34400 557300
rect 34600 557100 34800 557300
rect 35000 557100 35200 557300
rect 35400 557100 35600 557300
rect 35800 557100 36000 557300
rect 36200 557100 36400 557300
rect 36600 557100 36800 557300
rect 37000 557100 37200 557300
rect 37400 557100 37600 557300
rect 37800 557100 38000 557300
rect 38200 557100 38400 557300
rect 38600 557100 38800 557300
rect 39000 557100 39200 557300
rect 39400 557100 39600 557300
rect 39800 557100 40000 557300
rect 40200 557100 40400 557300
rect 40600 557100 40800 557300
rect 32600 556900 40800 557100
rect 32600 556700 32800 556900
rect 33000 556700 33200 556900
rect 33400 556700 33600 556900
rect 33800 556700 34000 556900
rect 34200 556700 34400 556900
rect 34600 556700 34800 556900
rect 35000 556700 35200 556900
rect 35400 556700 35600 556900
rect 35800 556700 36000 556900
rect 36200 556700 36400 556900
rect 36600 556700 36800 556900
rect 37000 556700 37200 556900
rect 37400 556700 37600 556900
rect 37800 556700 38000 556900
rect 38200 556700 38400 556900
rect 38600 556700 38800 556900
rect 39000 556700 39200 556900
rect 39400 556700 39600 556900
rect 39800 556700 40000 556900
rect 40200 556700 40400 556900
rect 40600 556700 40800 556900
rect 32600 556500 40800 556700
rect 32600 556300 32800 556500
rect 33000 556300 33200 556500
rect 33400 556300 33600 556500
rect 33800 556300 34000 556500
rect 34200 556300 34400 556500
rect 34600 556300 34800 556500
rect 35000 556300 35200 556500
rect 35400 556300 35600 556500
rect 35800 556300 36000 556500
rect 36200 556300 36400 556500
rect 36600 556300 36800 556500
rect 37000 556300 37200 556500
rect 37400 556300 37600 556500
rect 37800 556300 38000 556500
rect 38200 556300 38400 556500
rect 38600 556300 38800 556500
rect 39000 556300 39200 556500
rect 39400 556300 39600 556500
rect 39800 556300 40000 556500
rect 40200 556300 40400 556500
rect 40600 556300 40800 556500
rect 32600 556100 40800 556300
rect 32600 555900 32800 556100
rect 33000 555900 33200 556100
rect 33400 555900 33600 556100
rect 33800 555900 34000 556100
rect 34200 555900 34400 556100
rect 34600 555900 34800 556100
rect 35000 555900 35200 556100
rect 35400 555900 35600 556100
rect 35800 555900 36000 556100
rect 36200 555900 36400 556100
rect 36600 555900 36800 556100
rect 37000 555900 37200 556100
rect 37400 555900 37600 556100
rect 37800 555900 38000 556100
rect 38200 555900 38400 556100
rect 38600 555900 38800 556100
rect 39000 555900 39200 556100
rect 39400 555900 39600 556100
rect 39800 555900 40000 556100
rect 40200 555900 40400 556100
rect 40600 555900 40800 556100
rect 32600 555700 40800 555900
rect 32600 555500 32800 555700
rect 33000 555500 33200 555700
rect 33400 555500 33600 555700
rect 33800 555500 34000 555700
rect 34200 555500 34400 555700
rect 34600 555500 34800 555700
rect 35000 555500 35200 555700
rect 35400 555500 35600 555700
rect 35800 555500 36000 555700
rect 36200 555500 36400 555700
rect 36600 555500 36800 555700
rect 37000 555500 37200 555700
rect 37400 555500 37600 555700
rect 37800 555500 38000 555700
rect 38200 555500 38400 555700
rect 38600 555500 38800 555700
rect 39000 555500 39200 555700
rect 39400 555500 39600 555700
rect 39800 555500 40000 555700
rect 40200 555500 40400 555700
rect 40600 555500 40800 555700
rect 32600 555300 40800 555500
rect 32600 555100 32800 555300
rect 33000 555100 33200 555300
rect 33400 555100 33600 555300
rect 33800 555100 34000 555300
rect 34200 555100 34400 555300
rect 34600 555100 34800 555300
rect 35000 555100 35200 555300
rect 35400 555100 35600 555300
rect 35800 555100 36000 555300
rect 36200 555100 36400 555300
rect 36600 555100 36800 555300
rect 37000 555100 37200 555300
rect 37400 555100 37600 555300
rect 37800 555100 38000 555300
rect 38200 555100 38400 555300
rect 38600 555100 38800 555300
rect 39000 555100 39200 555300
rect 39400 555100 39600 555300
rect 39800 555100 40000 555300
rect 40200 555100 40400 555300
rect 40600 555100 40800 555300
rect 32600 554900 40800 555100
rect 32600 554700 32800 554900
rect 33000 554700 33200 554900
rect 33400 554700 33600 554900
rect 33800 554700 34000 554900
rect 34200 554700 34400 554900
rect 34600 554700 34800 554900
rect 35000 554700 35200 554900
rect 35400 554700 35600 554900
rect 35800 554700 36000 554900
rect 36200 554700 36400 554900
rect 36600 554700 36800 554900
rect 37000 554700 37200 554900
rect 37400 554700 37600 554900
rect 37800 554700 38000 554900
rect 38200 554700 38400 554900
rect 38600 554700 38800 554900
rect 39000 554700 39200 554900
rect 39400 554700 39600 554900
rect 39800 554700 40000 554900
rect 40200 554700 40400 554900
rect 40600 554700 40800 554900
rect 32600 554500 40800 554700
rect 32600 554300 32800 554500
rect 33000 554300 33200 554500
rect 33400 554300 33600 554500
rect 33800 554300 34000 554500
rect 34200 554300 34400 554500
rect 34600 554300 34800 554500
rect 35000 554300 35200 554500
rect 35400 554300 35600 554500
rect 35800 554300 36000 554500
rect 36200 554300 36400 554500
rect 36600 554300 36800 554500
rect 37000 554300 37200 554500
rect 37400 554300 37600 554500
rect 37800 554300 38000 554500
rect 38200 554300 38400 554500
rect 38600 554300 38800 554500
rect 39000 554300 39200 554500
rect 39400 554300 39600 554500
rect 39800 554300 40000 554500
rect 40200 554300 40400 554500
rect 40600 554300 40800 554500
rect 32600 554100 40800 554300
rect 32600 553900 32800 554100
rect 33000 553900 33200 554100
rect 33400 553900 33600 554100
rect 33800 553900 34000 554100
rect 34200 553900 34400 554100
rect 34600 553900 34800 554100
rect 35000 553900 35200 554100
rect 35400 553900 35600 554100
rect 35800 553900 36000 554100
rect 36200 553900 36400 554100
rect 36600 553900 36800 554100
rect 37000 553900 37200 554100
rect 37400 553900 37600 554100
rect 37800 553900 38000 554100
rect 38200 553900 38400 554100
rect 38600 553900 38800 554100
rect 39000 553900 39200 554100
rect 39400 553900 39600 554100
rect 39800 553900 40000 554100
rect 40200 553900 40400 554100
rect 40600 553900 40800 554100
rect 32600 553700 40800 553900
rect 32600 553500 32800 553700
rect 33000 553500 33200 553700
rect 33400 553500 33600 553700
rect 33800 553500 34000 553700
rect 34200 553500 34400 553700
rect 34600 553500 34800 553700
rect 35000 553500 35200 553700
rect 35400 553500 35600 553700
rect 35800 553500 36000 553700
rect 36200 553500 36400 553700
rect 36600 553500 36800 553700
rect 37000 553500 37200 553700
rect 37400 553500 37600 553700
rect 37800 553500 38000 553700
rect 38200 553500 38400 553700
rect 38600 553500 38800 553700
rect 39000 553500 39200 553700
rect 39400 553500 39600 553700
rect 39800 553500 40000 553700
rect 40200 553500 40400 553700
rect 40600 553500 40800 553700
rect 32600 553300 40800 553500
rect 32600 553100 32800 553300
rect 33000 553100 33200 553300
rect 33400 553100 33600 553300
rect 33800 553100 34000 553300
rect 34200 553100 34400 553300
rect 34600 553100 34800 553300
rect 35000 553100 35200 553300
rect 35400 553100 35600 553300
rect 35800 553100 36000 553300
rect 36200 553100 36400 553300
rect 36600 553100 36800 553300
rect 37000 553100 37200 553300
rect 37400 553100 37600 553300
rect 37800 553100 38000 553300
rect 38200 553100 38400 553300
rect 38600 553100 38800 553300
rect 39000 553100 39200 553300
rect 39400 553100 39600 553300
rect 39800 553100 40000 553300
rect 40200 553100 40400 553300
rect 40600 553100 40800 553300
rect 32600 552900 40800 553100
rect 32600 552700 32800 552900
rect 33000 552700 33200 552900
rect 33400 552700 33600 552900
rect 33800 552700 34000 552900
rect 34200 552700 34400 552900
rect 34600 552700 34800 552900
rect 35000 552700 35200 552900
rect 35400 552700 35600 552900
rect 35800 552700 36000 552900
rect 36200 552700 36400 552900
rect 36600 552700 36800 552900
rect 37000 552700 37200 552900
rect 37400 552700 37600 552900
rect 37800 552700 38000 552900
rect 38200 552700 38400 552900
rect 38600 552700 38800 552900
rect 39000 552700 39200 552900
rect 39400 552700 39600 552900
rect 39800 552700 40000 552900
rect 40200 552700 40400 552900
rect 40600 552700 40800 552900
rect 32600 552500 40800 552700
rect 32600 552300 32800 552500
rect 33000 552300 33200 552500
rect 33400 552300 33600 552500
rect 33800 552300 34000 552500
rect 34200 552300 34400 552500
rect 34600 552300 34800 552500
rect 35000 552300 35200 552500
rect 35400 552300 35600 552500
rect 35800 552300 36000 552500
rect 36200 552300 36400 552500
rect 36600 552300 36800 552500
rect 37000 552300 37200 552500
rect 37400 552300 37600 552500
rect 37800 552300 38000 552500
rect 38200 552300 38400 552500
rect 38600 552300 38800 552500
rect 39000 552300 39200 552500
rect 39400 552300 39600 552500
rect 39800 552300 40000 552500
rect 40200 552300 40400 552500
rect 40600 552300 40800 552500
rect 32600 552100 40800 552300
rect 32600 551900 32800 552100
rect 33000 551900 33200 552100
rect 33400 551900 33600 552100
rect 33800 551900 34000 552100
rect 34200 551900 34400 552100
rect 34600 551900 34800 552100
rect 35000 551900 35200 552100
rect 35400 551900 35600 552100
rect 35800 551900 36000 552100
rect 36200 551900 36400 552100
rect 36600 551900 36800 552100
rect 37000 551900 37200 552100
rect 37400 551900 37600 552100
rect 37800 551900 38000 552100
rect 38200 551900 38400 552100
rect 38600 551900 38800 552100
rect 39000 551900 39200 552100
rect 39400 551900 39600 552100
rect 39800 551900 40000 552100
rect 40200 551900 40400 552100
rect 40600 551900 40800 552100
rect 32600 551700 40800 551900
rect 32600 551500 32800 551700
rect 33000 551500 33200 551700
rect 33400 551500 33600 551700
rect 33800 551500 34000 551700
rect 34200 551500 34400 551700
rect 34600 551500 34800 551700
rect 35000 551500 35200 551700
rect 35400 551500 35600 551700
rect 35800 551500 36000 551700
rect 36200 551500 36400 551700
rect 36600 551500 36800 551700
rect 37000 551500 37200 551700
rect 37400 551500 37600 551700
rect 37800 551500 38000 551700
rect 38200 551500 38400 551700
rect 38600 551500 38800 551700
rect 39000 551500 39200 551700
rect 39400 551500 39600 551700
rect 39800 551500 40000 551700
rect 40200 551500 40400 551700
rect 40600 551500 40800 551700
rect 32600 551300 40800 551500
rect 32600 551100 32800 551300
rect 33000 551100 33200 551300
rect 33400 551100 33600 551300
rect 33800 551100 34000 551300
rect 34200 551100 34400 551300
rect 34600 551100 34800 551300
rect 35000 551100 35200 551300
rect 35400 551100 35600 551300
rect 35800 551100 36000 551300
rect 36200 551100 36400 551300
rect 36600 551100 36800 551300
rect 37000 551100 37200 551300
rect 37400 551100 37600 551300
rect 37800 551100 38000 551300
rect 38200 551100 38400 551300
rect 38600 551100 38800 551300
rect 39000 551100 39200 551300
rect 39400 551100 39600 551300
rect 39800 551100 40000 551300
rect 40200 551100 40400 551300
rect 40600 551100 40800 551300
rect 32600 550900 40800 551100
rect 32600 550700 32800 550900
rect 33000 550700 33200 550900
rect 33400 550700 33600 550900
rect 33800 550700 34000 550900
rect 34200 550700 34400 550900
rect 34600 550700 34800 550900
rect 35000 550700 35200 550900
rect 35400 550700 35600 550900
rect 35800 550700 36000 550900
rect 36200 550700 36400 550900
rect 36600 550700 36800 550900
rect 37000 550700 37200 550900
rect 37400 550700 37600 550900
rect 37800 550700 38000 550900
rect 38200 550700 38400 550900
rect 38600 550700 38800 550900
rect 39000 550700 39200 550900
rect 39400 550700 39600 550900
rect 39800 550700 40000 550900
rect 40200 550700 40400 550900
rect 40600 550700 40800 550900
rect 32600 550500 40800 550700
rect 32600 550300 32800 550500
rect 33000 550300 33200 550500
rect 33400 550300 33600 550500
rect 33800 550300 34000 550500
rect 34200 550300 34400 550500
rect 34600 550300 34800 550500
rect 35000 550300 35200 550500
rect 35400 550300 35600 550500
rect 35800 550300 36000 550500
rect 36200 550300 36400 550500
rect 36600 550300 36800 550500
rect 37000 550300 37200 550500
rect 37400 550300 37600 550500
rect 37800 550300 38000 550500
rect 38200 550300 38400 550500
rect 38600 550300 38800 550500
rect 39000 550300 39200 550500
rect 39400 550300 39600 550500
rect 39800 550300 40000 550500
rect 40200 550300 40400 550500
rect 40600 550300 40800 550500
rect 32600 550100 40800 550300
rect 32600 549900 32800 550100
rect 33000 549900 33200 550100
rect 33400 549900 33600 550100
rect 33800 549900 34000 550100
rect 34200 549900 34400 550100
rect 34600 549900 34800 550100
rect 35000 549900 35200 550100
rect 35400 549900 35600 550100
rect 35800 549900 36000 550100
rect 36200 549900 36400 550100
rect 36600 549900 36800 550100
rect 37000 549900 37200 550100
rect 37400 549900 37600 550100
rect 37800 549900 38000 550100
rect 38200 549900 38400 550100
rect 38600 549900 38800 550100
rect 39000 549900 39200 550100
rect 39400 549900 39600 550100
rect 39800 549900 40000 550100
rect 40200 549900 40400 550100
rect 40600 549900 40800 550100
rect 32600 549700 40800 549900
rect 32600 549500 32800 549700
rect 33000 549500 33200 549700
rect 33400 549500 33600 549700
rect 33800 549500 34000 549700
rect 34200 549500 34400 549700
rect 34600 549500 34800 549700
rect 35000 549500 35200 549700
rect 35400 549500 35600 549700
rect 35800 549500 36000 549700
rect 36200 549500 36400 549700
rect 36600 549500 36800 549700
rect 37000 549500 37200 549700
rect 37400 549500 37600 549700
rect 37800 549500 38000 549700
rect 38200 549500 38400 549700
rect 38600 549500 38800 549700
rect 39000 549500 39200 549700
rect 39400 549500 39600 549700
rect 39800 549500 40000 549700
rect 40200 549500 40400 549700
rect 40600 549500 40800 549700
rect 32600 549400 40800 549500
<< via4 >>
rect 44010 695370 44280 695640
rect 45060 695370 45330 695640
rect 41840 694890 42090 695140
rect 43740 694880 43990 695130
rect 45320 694880 45570 695130
rect 47220 694880 47470 695130
rect 44010 693730 44280 694000
rect 45060 693730 45330 694000
rect 43340 693220 43600 693480
rect 44610 693220 44870 693480
rect 45870 693220 46130 693480
rect 43780 692130 44040 692390
rect 45280 692130 45540 692390
rect 43340 691670 43600 691930
rect 44610 691670 44870 691930
rect 45870 691670 46130 691930
rect 44520 689030 44780 689290
rect 44520 687510 44780 687770
rect 43500 686420 43750 686670
rect 45560 686420 45810 686670
rect 38700 685780 38940 686020
rect 39060 685780 39300 686020
rect 44530 686000 44780 686250
rect 38700 685440 38940 685680
rect 39060 685440 39300 685680
rect 49950 685780 50190 686020
rect 50310 685780 50550 686020
rect 49950 685440 50190 685680
rect 50310 685440 50550 685680
rect 43240 684900 43490 685150
rect 45820 684900 46070 685150
rect 44530 684470 44780 684720
rect 43750 683620 43990 683680
rect 43750 683500 43810 683620
rect 43810 683500 43930 683620
rect 43930 683500 43990 683620
rect 43750 683440 43990 683500
rect 44270 683600 44510 683680
rect 44270 683520 44350 683600
rect 44350 683520 44430 683600
rect 44430 683520 44510 683600
rect 44270 683440 44510 683520
rect 44790 683600 45030 683680
rect 44790 683520 44870 683600
rect 44870 683520 44950 683600
rect 44950 683520 45030 683600
rect 44790 683440 45030 683520
rect 45310 683600 45550 683680
rect 45310 683520 45390 683600
rect 45390 683520 45470 683600
rect 45470 683520 45550 683600
rect 45310 683440 45550 683520
rect 32800 673700 33100 674000
rect 33300 673700 33600 674000
rect 33800 673700 34100 674000
rect 34300 673700 34600 674000
rect 34800 673700 35100 674000
rect 35300 673700 35600 674000
rect 35800 673700 36100 674000
rect 36300 673700 36600 674000
rect 36800 673700 37100 674000
rect 37300 673700 37600 674000
rect 37800 673700 38100 674000
rect 38300 673700 38600 674000
rect 38800 673700 39100 674000
rect 39300 673700 39600 674000
rect 39800 673700 40100 674000
rect 40300 673700 40600 674000
rect 44210 673780 44450 674020
rect 44770 673780 45010 674020
rect 41200 673300 41440 673540
rect 50100 673700 50400 674000
rect 44210 673300 44450 673540
rect 44770 673300 45010 673540
rect 32800 672900 33100 673200
rect 33300 672900 33600 673200
rect 33800 672900 34100 673200
rect 34300 672900 34600 673200
rect 34800 672900 35100 673200
rect 35300 672900 35600 673200
rect 35800 672900 36100 673200
rect 36300 672900 36600 673200
rect 36800 672900 37100 673200
rect 37300 672900 37600 673200
rect 37800 672900 38100 673200
rect 38300 672900 38600 673200
rect 38800 672900 39100 673200
rect 39300 672900 39600 673200
rect 39800 672900 40100 673200
rect 40300 672900 40600 673200
rect 32800 670400 33100 670700
rect 33300 670400 33600 670700
rect 33800 670400 34100 670700
rect 34300 670400 34600 670700
rect 34800 670400 35100 670700
rect 35300 670400 35600 670700
rect 35800 670400 36100 670700
rect 36300 670400 36600 670700
rect 36800 670400 37100 670700
rect 37300 670400 37600 670700
rect 37800 670400 38100 670700
rect 38300 670400 38600 670700
rect 38800 670400 39100 670700
rect 39300 670400 39600 670700
rect 39800 670400 40100 670700
rect 40300 670400 40600 670700
rect 47900 673300 48140 673540
rect 50100 673300 50400 673600
rect 44210 672820 44450 673060
rect 44770 672820 45010 673060
rect 50100 672900 50400 673200
rect 44210 670580 44450 670820
rect 44770 670580 45010 670820
rect 41200 670100 41440 670340
rect 44210 670100 44450 670340
rect 44770 670100 45010 670340
rect 32800 669700 33100 670000
rect 33300 669700 33600 670000
rect 33800 669700 34100 670000
rect 34300 669700 34600 670000
rect 34800 669700 35100 670000
rect 35300 669700 35600 670000
rect 35800 669700 36100 670000
rect 36300 669700 36600 670000
rect 36800 669700 37100 670000
rect 37300 669700 37600 670000
rect 37800 669700 38100 670000
rect 38300 669700 38600 670000
rect 38800 669700 39100 670000
rect 39300 669700 39600 670000
rect 39800 669700 40100 670000
rect 40300 669700 40600 670000
rect 32800 667100 33100 667400
rect 33300 667100 33600 667400
rect 33800 667100 34100 667400
rect 34300 667100 34600 667400
rect 34800 667100 35100 667400
rect 35300 667100 35600 667400
rect 35800 667100 36100 667400
rect 36300 667100 36600 667400
rect 36800 667100 37100 667400
rect 37300 667100 37600 667400
rect 37800 667100 38100 667400
rect 38300 667100 38600 667400
rect 38800 667100 39100 667400
rect 39300 667100 39600 667400
rect 39800 667100 40100 667400
rect 40300 667100 40600 667400
rect 47900 670100 48140 670340
rect 44210 669620 44450 669860
rect 44770 669620 45010 669860
rect 44210 667260 44450 667500
rect 44770 667260 45010 667500
rect 41200 666780 41440 667020
rect 44210 666780 44450 667020
rect 44770 666780 45010 667020
rect 32800 666400 33100 666700
rect 33300 666400 33600 666700
rect 33800 666400 34100 666700
rect 34300 666400 34600 666700
rect 34800 666400 35100 666700
rect 35300 666400 35600 666700
rect 35800 666400 36100 666700
rect 36300 666400 36600 666700
rect 36800 666400 37100 666700
rect 37300 666400 37600 666700
rect 37800 666400 38100 666700
rect 38300 666400 38600 666700
rect 38800 666400 39100 666700
rect 39300 666400 39600 666700
rect 39800 666400 40100 666700
rect 40300 666400 40600 666700
rect 47900 666780 48140 667020
rect 44210 666300 44450 666540
rect 44770 666300 45010 666540
rect 2500 648300 2800 648600
rect 3000 648300 3300 648600
rect 3500 648300 3800 648600
rect 2500 647800 2800 648100
rect 3000 647800 3300 648100
rect 3500 647800 3800 648100
rect 2500 647300 2800 647600
rect 3000 647300 3300 647600
rect 3500 647300 3800 647600
rect 2500 646800 2800 647100
rect 3000 646800 3300 647100
rect 3500 646800 3800 647100
rect 2500 646300 2800 646600
rect 3000 646300 3300 646600
rect 3500 646300 3800 646600
rect 2500 645800 2800 646100
rect 3000 645800 3300 646100
rect 3500 645800 3800 646100
rect 2500 645300 2800 645600
rect 3000 645300 3300 645600
rect 3500 645300 3800 645600
rect 2500 644800 2800 645100
rect 3000 644800 3300 645100
rect 3500 644800 3800 645100
rect 2500 644300 2800 644600
rect 3000 644300 3300 644600
rect 3500 644300 3800 644600
rect 2500 643800 2800 644100
rect 3000 643800 3300 644100
rect 3500 643800 3800 644100
rect 2500 643300 2800 643600
rect 3000 643300 3300 643600
rect 3500 643300 3800 643600
rect 2500 642800 2800 643100
rect 3000 642800 3300 643100
rect 3500 642800 3800 643100
rect 2500 642300 2800 642600
rect 3000 642300 3300 642600
rect 3500 642300 3800 642600
rect 2500 641800 2800 642100
rect 3000 641800 3300 642100
rect 3500 641800 3800 642100
rect 2500 641300 2800 641600
rect 3000 641300 3300 641600
rect 3500 641300 3800 641600
rect 2500 640800 2800 641100
rect 3000 640800 3300 641100
rect 3500 640800 3800 641100
rect 2500 640300 2800 640600
rect 3000 640300 3300 640600
rect 3500 640300 3800 640600
rect 2500 639800 2800 640100
rect 3000 639800 3300 640100
rect 3500 639800 3800 640100
rect 2500 639300 2800 639600
rect 3000 639300 3300 639600
rect 3500 639300 3800 639600
rect 2500 638800 2800 639100
rect 3000 638800 3300 639100
rect 3500 638800 3800 639100
rect 2500 638300 2800 638600
rect 3000 638300 3300 638600
rect 3500 638300 3800 638600
rect 2500 637800 2800 638100
rect 3000 637800 3300 638100
rect 3500 637800 3800 638100
rect 2500 637300 2800 637600
rect 3000 637300 3300 637600
rect 3500 637300 3800 637600
rect 2500 636800 2800 637100
rect 3000 636800 3300 637100
rect 3500 636800 3800 637100
rect 2500 636300 2800 636600
rect 3000 636300 3300 636600
rect 3500 636300 3800 636600
rect 2500 635800 2800 636100
rect 3000 635800 3300 636100
rect 3500 635800 3800 636100
rect 2500 635300 2800 635600
rect 3000 635300 3300 635600
rect 3500 635300 3800 635600
rect 2500 634800 2800 635100
rect 3000 634800 3300 635100
rect 3500 634800 3800 635100
rect 2500 634300 2800 634600
rect 3000 634300 3300 634600
rect 3500 634300 3800 634600
rect 58000 648300 58300 648600
rect 58500 648300 58800 648600
rect 59000 648300 59300 648600
rect 59500 648300 59800 648600
rect 60000 648300 60300 648600
rect 60500 648300 60800 648600
rect 61000 648300 61300 648600
rect 61500 648300 61800 648600
rect 58000 647800 58300 648100
rect 58500 647800 58800 648100
rect 59000 647800 59300 648100
rect 59500 647800 59800 648100
rect 60000 647800 60300 648100
rect 60500 647800 60800 648100
rect 61000 647800 61300 648100
rect 61500 647800 61800 648100
rect 58000 647300 58300 647600
rect 58500 647300 58800 647600
rect 59000 647300 59300 647600
rect 59500 647300 59800 647600
rect 60000 647300 60300 647600
rect 60500 647300 60800 647600
rect 61000 647300 61300 647600
rect 61500 647300 61800 647600
rect 58000 646800 58300 647100
rect 58500 646800 58800 647100
rect 59000 646800 59300 647100
rect 59500 646800 59800 647100
rect 60000 646800 60300 647100
rect 60500 646800 60800 647100
rect 61000 646800 61300 647100
rect 61500 646800 61800 647100
rect 58000 646300 58300 646600
rect 58500 646300 58800 646600
rect 59000 646300 59300 646600
rect 59500 646300 59800 646600
rect 60000 646300 60300 646600
rect 60500 646300 60800 646600
rect 61000 646300 61300 646600
rect 61500 646300 61800 646600
rect 58000 645800 58300 646100
rect 58500 645800 58800 646100
rect 59000 645800 59300 646100
rect 59500 645800 59800 646100
rect 60000 645800 60300 646100
rect 60500 645800 60800 646100
rect 61000 645800 61300 646100
rect 61500 645800 61800 646100
rect 58000 645300 58300 645600
rect 58500 645300 58800 645600
rect 59000 645300 59300 645600
rect 59500 645300 59800 645600
rect 60000 645300 60300 645600
rect 60500 645300 60800 645600
rect 61000 645300 61300 645600
rect 61500 645300 61800 645600
rect 58000 644800 58300 645100
rect 58500 644800 58800 645100
rect 59000 644800 59300 645100
rect 59500 644800 59800 645100
rect 60000 644800 60300 645100
rect 60500 644800 60800 645100
rect 61000 644800 61300 645100
rect 61500 644800 61800 645100
rect 58000 644300 58300 644600
rect 58500 644300 58800 644600
rect 59000 644300 59300 644600
rect 59500 644300 59800 644600
rect 60000 644300 60300 644600
rect 60500 644300 60800 644600
rect 61000 644300 61300 644600
rect 61500 644300 61800 644600
rect 58000 643800 58300 644100
rect 58500 643800 58800 644100
rect 59000 643800 59300 644100
rect 59500 643800 59800 644100
rect 60000 643800 60300 644100
rect 60500 643800 60800 644100
rect 61000 643800 61300 644100
rect 61500 643800 61800 644100
rect 58000 643300 58300 643600
rect 58500 643300 58800 643600
rect 59000 643300 59300 643600
rect 59500 643300 59800 643600
rect 60000 643300 60300 643600
rect 60500 643300 60800 643600
rect 61000 643300 61300 643600
rect 61500 643300 61800 643600
rect 58000 642800 58300 643100
rect 58500 642800 58800 643100
rect 59000 642800 59300 643100
rect 59500 642800 59800 643100
rect 60000 642800 60300 643100
rect 60500 642800 60800 643100
rect 61000 642800 61300 643100
rect 61500 642800 61800 643100
rect 58000 642300 58300 642600
rect 58500 642300 58800 642600
rect 59000 642300 59300 642600
rect 59500 642300 59800 642600
rect 60000 642300 60300 642600
rect 60500 642300 60800 642600
rect 61000 642300 61300 642600
rect 61500 642300 61800 642600
rect 58000 641800 58300 642100
rect 58500 641800 58800 642100
rect 59000 641800 59300 642100
rect 59500 641800 59800 642100
rect 60000 641800 60300 642100
rect 60500 641800 60800 642100
rect 61000 641800 61300 642100
rect 61500 641800 61800 642100
rect 58000 641300 58300 641600
rect 58500 641300 58800 641600
rect 59000 641300 59300 641600
rect 59500 641300 59800 641600
rect 60000 641300 60300 641600
rect 60500 641300 60800 641600
rect 61000 641300 61300 641600
rect 61500 641300 61800 641600
rect 58000 640800 58300 641100
rect 58500 640800 58800 641100
rect 59000 640800 59300 641100
rect 59500 640800 59800 641100
rect 60000 640800 60300 641100
rect 60500 640800 60800 641100
rect 61000 640800 61300 641100
rect 61500 640800 61800 641100
rect 58000 640300 58300 640600
rect 58500 640300 58800 640600
rect 59000 640300 59300 640600
rect 59500 640300 59800 640600
rect 60000 640300 60300 640600
rect 60500 640300 60800 640600
rect 61000 640300 61300 640600
rect 61500 640300 61800 640600
rect 58000 639800 58300 640100
rect 58500 639800 58800 640100
rect 59000 639800 59300 640100
rect 59500 639800 59800 640100
rect 60000 639800 60300 640100
rect 60500 639800 60800 640100
rect 61000 639800 61300 640100
rect 61500 639800 61800 640100
rect 58000 639300 58300 639600
rect 58500 639300 58800 639600
rect 59000 639300 59300 639600
rect 59500 639300 59800 639600
rect 60000 639300 60300 639600
rect 60500 639300 60800 639600
rect 61000 639300 61300 639600
rect 61500 639300 61800 639600
rect 58000 638800 58300 639100
rect 58500 638800 58800 639100
rect 59000 638800 59300 639100
rect 59500 638800 59800 639100
rect 60000 638800 60300 639100
rect 60500 638800 60800 639100
rect 61000 638800 61300 639100
rect 61500 638800 61800 639100
rect 58000 638300 58300 638600
rect 58500 638300 58800 638600
rect 59000 638300 59300 638600
rect 59500 638300 59800 638600
rect 60000 638300 60300 638600
rect 60500 638300 60800 638600
rect 61000 638300 61300 638600
rect 61500 638300 61800 638600
rect 58000 637800 58300 638100
rect 58500 637800 58800 638100
rect 59000 637800 59300 638100
rect 59500 637800 59800 638100
rect 60000 637800 60300 638100
rect 60500 637800 60800 638100
rect 61000 637800 61300 638100
rect 61500 637800 61800 638100
rect 58000 637300 58300 637600
rect 58500 637300 58800 637600
rect 59000 637300 59300 637600
rect 59500 637300 59800 637600
rect 60000 637300 60300 637600
rect 60500 637300 60800 637600
rect 61000 637300 61300 637600
rect 61500 637300 61800 637600
rect 58000 636800 58300 637100
rect 58500 636800 58800 637100
rect 59000 636800 59300 637100
rect 59500 636800 59800 637100
rect 60000 636800 60300 637100
rect 60500 636800 60800 637100
rect 61000 636800 61300 637100
rect 61500 636800 61800 637100
rect 58000 636300 58300 636600
rect 58500 636300 58800 636600
rect 59000 636300 59300 636600
rect 59500 636300 59800 636600
rect 60000 636300 60300 636600
rect 60500 636300 60800 636600
rect 61000 636300 61300 636600
rect 61500 636300 61800 636600
rect 58000 635800 58300 636100
rect 58500 635800 58800 636100
rect 59000 635800 59300 636100
rect 59500 635800 59800 636100
rect 60000 635800 60300 636100
rect 60500 635800 60800 636100
rect 61000 635800 61300 636100
rect 61500 635800 61800 636100
rect 58000 635300 58300 635600
rect 58500 635300 58800 635600
rect 59000 635300 59300 635600
rect 59500 635300 59800 635600
rect 60000 635300 60300 635600
rect 60500 635300 60800 635600
rect 61000 635300 61300 635600
rect 61500 635300 61800 635600
rect 58000 634800 58300 635100
rect 58500 634800 58800 635100
rect 59000 634800 59300 635100
rect 59500 634800 59800 635100
rect 60000 634800 60300 635100
rect 60500 634800 60800 635100
rect 61000 634800 61300 635100
rect 61500 634800 61800 635100
rect 58000 634300 58300 634600
rect 58500 634300 58800 634600
rect 59000 634300 59300 634600
rect 59500 634300 59800 634600
rect 60000 634300 60300 634600
rect 60500 634300 60800 634600
rect 61000 634300 61300 634600
rect 61500 634300 61800 634600
<< metal5 >>
rect 43980 695640 45360 695690
rect 43980 695370 44010 695640
rect 44280 695370 45060 695640
rect 45330 695370 45360 695640
rect 43980 695170 45360 695370
rect 41810 695140 47510 695170
rect 41810 694890 41840 695140
rect 42090 695130 47510 695140
rect 42090 694890 43740 695130
rect 41810 694880 43740 694890
rect 43990 694880 45320 695130
rect 45570 694880 47220 695130
rect 47470 694880 47510 695130
rect 41810 694840 47510 694880
rect 43980 694000 45360 694840
rect 43980 693730 44010 694000
rect 44280 693730 45060 694000
rect 45330 693730 45360 694000
rect 43980 693510 45360 693730
rect 43190 693480 46170 693510
rect 43190 693220 43340 693480
rect 43600 693220 44610 693480
rect 44870 693220 45870 693480
rect 46130 693220 46170 693480
rect 43190 693190 46170 693220
rect 43980 692420 45360 693190
rect 43750 692390 45570 692420
rect 43750 692130 43780 692390
rect 44040 692130 45280 692390
rect 45540 692130 45570 692390
rect 43750 691960 45570 692130
rect 43300 691930 46170 691960
rect 43300 691670 43340 691930
rect 43600 691670 44610 691930
rect 44870 691670 45870 691930
rect 46130 691670 46170 691930
rect 43300 691640 46170 691670
rect 44430 689290 44870 689330
rect 44430 689030 44520 689290
rect 44780 689030 44870 689290
rect 44430 687770 44870 689030
rect 44430 687510 44520 687770
rect 44780 687510 44870 687770
rect 44430 686710 44870 687510
rect 41820 686670 47460 686710
rect 41820 686420 43500 686670
rect 43750 686420 45560 686670
rect 45810 686420 47460 686670
rect 41820 686250 47460 686420
rect 41820 686050 44530 686250
rect 38670 686020 44530 686050
rect 38670 685780 38700 686020
rect 38940 685780 39060 686020
rect 39300 686000 44530 686020
rect 44780 686050 47460 686250
rect 44780 686020 50580 686050
rect 44780 686000 49950 686020
rect 39300 685780 49950 686000
rect 50190 685780 50310 686020
rect 50550 685780 50580 686020
rect 38670 685680 50580 685780
rect 38670 685440 38700 685680
rect 38940 685440 39060 685680
rect 39300 685440 49950 685680
rect 50190 685440 50310 685680
rect 50550 685440 50580 685680
rect 38670 685410 50580 685440
rect 41820 685150 47460 685410
rect 41820 684900 43240 685150
rect 43490 684900 45820 685150
rect 46070 684900 47460 685150
rect 41820 684860 47460 684900
rect 44440 684720 44880 684860
rect 44440 684470 44530 684720
rect 44780 684470 44880 684720
rect 44440 684400 44880 684470
rect 43490 683680 45850 684020
rect 43490 683440 43750 683680
rect 43990 683440 44270 683680
rect 44510 683440 44790 683680
rect 45030 683440 45310 683680
rect 45550 683440 45850 683680
rect 43490 683380 45850 683440
rect 32600 674020 51300 674200
rect 32600 674000 44210 674020
rect 32600 673700 32800 674000
rect 33100 673700 33300 674000
rect 33600 673700 33800 674000
rect 34100 673700 34300 674000
rect 34600 673700 34800 674000
rect 35100 673700 35300 674000
rect 35600 673700 35800 674000
rect 36100 673700 36300 674000
rect 36600 673700 36800 674000
rect 37100 673700 37300 674000
rect 37600 673700 37800 674000
rect 38100 673700 38300 674000
rect 38600 673700 38800 674000
rect 39100 673700 39300 674000
rect 39600 673700 39800 674000
rect 40100 673700 40300 674000
rect 40600 673780 44210 674000
rect 44450 673780 44770 674020
rect 45010 674000 51300 674020
rect 45010 673780 50100 674000
rect 40600 673700 50100 673780
rect 50400 673700 51300 674000
rect 32600 673600 51300 673700
rect 32600 673540 50100 673600
rect 32600 673300 41200 673540
rect 41440 673300 44210 673540
rect 44450 673300 44770 673540
rect 45010 673300 47900 673540
rect 48140 673300 50100 673540
rect 50400 673300 51300 673600
rect 32600 673200 51300 673300
rect 32600 672900 32800 673200
rect 33100 672900 33300 673200
rect 33600 672900 33800 673200
rect 34100 672900 34300 673200
rect 34600 672900 34800 673200
rect 35100 672900 35300 673200
rect 35600 672900 35800 673200
rect 36100 672900 36300 673200
rect 36600 672900 36800 673200
rect 37100 672900 37300 673200
rect 37600 672900 37800 673200
rect 38100 672900 38300 673200
rect 38600 672900 38800 673200
rect 39100 672900 39300 673200
rect 39600 672900 39800 673200
rect 40100 672900 40300 673200
rect 40600 673060 50100 673200
rect 40600 672900 44210 673060
rect 32600 672820 44210 672900
rect 44450 672820 44770 673060
rect 45010 672900 50100 673060
rect 50400 672900 51300 673200
rect 45010 672820 51300 672900
rect 32600 672700 51300 672820
rect 32600 670820 48300 670900
rect 32600 670700 44210 670820
rect 32600 670400 32800 670700
rect 33100 670400 33300 670700
rect 33600 670400 33800 670700
rect 34100 670400 34300 670700
rect 34600 670400 34800 670700
rect 35100 670400 35300 670700
rect 35600 670400 35800 670700
rect 36100 670400 36300 670700
rect 36600 670400 36800 670700
rect 37100 670400 37300 670700
rect 37600 670400 37800 670700
rect 38100 670400 38300 670700
rect 38600 670400 38800 670700
rect 39100 670400 39300 670700
rect 39600 670400 39800 670700
rect 40100 670400 40300 670700
rect 40600 670580 44210 670700
rect 44450 670580 44770 670820
rect 45010 670580 48300 670820
rect 40600 670400 48300 670580
rect 32600 670340 48300 670400
rect 32600 670100 41200 670340
rect 41440 670100 44210 670340
rect 44450 670100 44770 670340
rect 45010 670100 47900 670340
rect 48140 670100 48300 670340
rect 32600 670000 48300 670100
rect 32600 669700 32800 670000
rect 33100 669700 33300 670000
rect 33600 669700 33800 670000
rect 34100 669700 34300 670000
rect 34600 669700 34800 670000
rect 35100 669700 35300 670000
rect 35600 669700 35800 670000
rect 36100 669700 36300 670000
rect 36600 669700 36800 670000
rect 37100 669700 37300 670000
rect 37600 669700 37800 670000
rect 38100 669700 38300 670000
rect 38600 669700 38800 670000
rect 39100 669700 39300 670000
rect 39600 669700 39800 670000
rect 40100 669700 40300 670000
rect 40600 669860 48300 670000
rect 40600 669700 44210 669860
rect 32600 669620 44210 669700
rect 44450 669620 44770 669860
rect 45010 669620 48300 669860
rect 32600 669500 48300 669620
rect 32600 667500 48300 667600
rect 32600 667400 44210 667500
rect 32600 667100 32800 667400
rect 33100 667100 33300 667400
rect 33600 667100 33800 667400
rect 34100 667100 34300 667400
rect 34600 667100 34800 667400
rect 35100 667100 35300 667400
rect 35600 667100 35800 667400
rect 36100 667100 36300 667400
rect 36600 667100 36800 667400
rect 37100 667100 37300 667400
rect 37600 667100 37800 667400
rect 38100 667100 38300 667400
rect 38600 667100 38800 667400
rect 39100 667100 39300 667400
rect 39600 667100 39800 667400
rect 40100 667100 40300 667400
rect 40600 667260 44210 667400
rect 44450 667260 44770 667500
rect 45010 667260 48300 667500
rect 40600 667100 48300 667260
rect 32600 667020 48300 667100
rect 32600 666780 41200 667020
rect 41440 666780 44210 667020
rect 44450 666780 44770 667020
rect 45010 666780 47900 667020
rect 48140 666780 48300 667020
rect 32600 666700 48300 666780
rect 32600 666400 32800 666700
rect 33100 666400 33300 666700
rect 33600 666400 33800 666700
rect 34100 666400 34300 666700
rect 34600 666400 34800 666700
rect 35100 666400 35300 666700
rect 35600 666400 35800 666700
rect 36100 666400 36300 666700
rect 36600 666400 36800 666700
rect 37100 666400 37300 666700
rect 37600 666400 37800 666700
rect 38100 666400 38300 666700
rect 38600 666400 38800 666700
rect 39100 666400 39300 666700
rect 39600 666400 39800 666700
rect 40100 666400 40300 666700
rect 40600 666540 48300 666700
rect 40600 666400 44210 666540
rect 32600 666300 44210 666400
rect 44450 666300 44770 666540
rect 45010 666300 48300 666540
rect 32600 666200 48300 666300
rect 2300 648600 62200 648800
rect 2300 648300 2500 648600
rect 2800 648300 3000 648600
rect 3300 648300 3500 648600
rect 3800 648300 58000 648600
rect 58300 648300 58500 648600
rect 58800 648300 59000 648600
rect 59300 648300 59500 648600
rect 59800 648300 60000 648600
rect 60300 648300 60500 648600
rect 60800 648300 61000 648600
rect 61300 648300 61500 648600
rect 61800 648300 62200 648600
rect 2300 648100 62200 648300
rect 2300 647800 2500 648100
rect 2800 647800 3000 648100
rect 3300 647800 3500 648100
rect 3800 647800 58000 648100
rect 58300 647800 58500 648100
rect 58800 647800 59000 648100
rect 59300 647800 59500 648100
rect 59800 647800 60000 648100
rect 60300 647800 60500 648100
rect 60800 647800 61000 648100
rect 61300 647800 61500 648100
rect 61800 647800 62200 648100
rect 2300 647600 62200 647800
rect 2300 647300 2500 647600
rect 2800 647300 3000 647600
rect 3300 647300 3500 647600
rect 3800 647300 58000 647600
rect 58300 647300 58500 647600
rect 58800 647300 59000 647600
rect 59300 647300 59500 647600
rect 59800 647300 60000 647600
rect 60300 647300 60500 647600
rect 60800 647300 61000 647600
rect 61300 647300 61500 647600
rect 61800 647300 62200 647600
rect 2300 647100 62200 647300
rect 2300 646800 2500 647100
rect 2800 646800 3000 647100
rect 3300 646800 3500 647100
rect 3800 646800 58000 647100
rect 58300 646800 58500 647100
rect 58800 646800 59000 647100
rect 59300 646800 59500 647100
rect 59800 646800 60000 647100
rect 60300 646800 60500 647100
rect 60800 646800 61000 647100
rect 61300 646800 61500 647100
rect 61800 646800 62200 647100
rect 2300 646600 62200 646800
rect 2300 646300 2500 646600
rect 2800 646300 3000 646600
rect 3300 646300 3500 646600
rect 3800 646300 58000 646600
rect 58300 646300 58500 646600
rect 58800 646300 59000 646600
rect 59300 646300 59500 646600
rect 59800 646300 60000 646600
rect 60300 646300 60500 646600
rect 60800 646300 61000 646600
rect 61300 646300 61500 646600
rect 61800 646300 62200 646600
rect 2300 646100 62200 646300
rect 2300 645800 2500 646100
rect 2800 645800 3000 646100
rect 3300 645800 3500 646100
rect 3800 645800 58000 646100
rect 58300 645800 58500 646100
rect 58800 645800 59000 646100
rect 59300 645800 59500 646100
rect 59800 645800 60000 646100
rect 60300 645800 60500 646100
rect 60800 645800 61000 646100
rect 61300 645800 61500 646100
rect 61800 645800 62200 646100
rect 2300 645600 62200 645800
rect 2300 645300 2500 645600
rect 2800 645300 3000 645600
rect 3300 645300 3500 645600
rect 3800 645300 58000 645600
rect 58300 645300 58500 645600
rect 58800 645300 59000 645600
rect 59300 645300 59500 645600
rect 59800 645300 60000 645600
rect 60300 645300 60500 645600
rect 60800 645300 61000 645600
rect 61300 645300 61500 645600
rect 61800 645300 62200 645600
rect 2300 645100 62200 645300
rect 2300 644800 2500 645100
rect 2800 644800 3000 645100
rect 3300 644800 3500 645100
rect 3800 644800 58000 645100
rect 58300 644800 58500 645100
rect 58800 644800 59000 645100
rect 59300 644800 59500 645100
rect 59800 644800 60000 645100
rect 60300 644800 60500 645100
rect 60800 644800 61000 645100
rect 61300 644800 61500 645100
rect 61800 644800 62200 645100
rect 2300 644600 62200 644800
rect 2300 644300 2500 644600
rect 2800 644300 3000 644600
rect 3300 644300 3500 644600
rect 3800 644300 58000 644600
rect 58300 644300 58500 644600
rect 58800 644300 59000 644600
rect 59300 644300 59500 644600
rect 59800 644300 60000 644600
rect 60300 644300 60500 644600
rect 60800 644300 61000 644600
rect 61300 644300 61500 644600
rect 61800 644300 62200 644600
rect 2300 644100 62200 644300
rect 2300 643800 2500 644100
rect 2800 643800 3000 644100
rect 3300 643800 3500 644100
rect 3800 643800 58000 644100
rect 58300 643800 58500 644100
rect 58800 643800 59000 644100
rect 59300 643800 59500 644100
rect 59800 643800 60000 644100
rect 60300 643800 60500 644100
rect 60800 643800 61000 644100
rect 61300 643800 61500 644100
rect 61800 643800 62200 644100
rect 2300 643600 62200 643800
rect 2300 643300 2500 643600
rect 2800 643300 3000 643600
rect 3300 643300 3500 643600
rect 3800 643300 58000 643600
rect 58300 643300 58500 643600
rect 58800 643300 59000 643600
rect 59300 643300 59500 643600
rect 59800 643300 60000 643600
rect 60300 643300 60500 643600
rect 60800 643300 61000 643600
rect 61300 643300 61500 643600
rect 61800 643300 62200 643600
rect 2300 643100 62200 643300
rect 2300 642800 2500 643100
rect 2800 642800 3000 643100
rect 3300 642800 3500 643100
rect 3800 642800 58000 643100
rect 58300 642800 58500 643100
rect 58800 642800 59000 643100
rect 59300 642800 59500 643100
rect 59800 642800 60000 643100
rect 60300 642800 60500 643100
rect 60800 642800 61000 643100
rect 61300 642800 61500 643100
rect 61800 642800 62200 643100
rect 2300 642600 62200 642800
rect 2300 642300 2500 642600
rect 2800 642300 3000 642600
rect 3300 642300 3500 642600
rect 3800 642300 58000 642600
rect 58300 642300 58500 642600
rect 58800 642300 59000 642600
rect 59300 642300 59500 642600
rect 59800 642300 60000 642600
rect 60300 642300 60500 642600
rect 60800 642300 61000 642600
rect 61300 642300 61500 642600
rect 61800 642300 62200 642600
rect 2300 642100 62200 642300
rect 2300 641800 2500 642100
rect 2800 641800 3000 642100
rect 3300 641800 3500 642100
rect 3800 641800 58000 642100
rect 58300 641800 58500 642100
rect 58800 641800 59000 642100
rect 59300 641800 59500 642100
rect 59800 641800 60000 642100
rect 60300 641800 60500 642100
rect 60800 641800 61000 642100
rect 61300 641800 61500 642100
rect 61800 641800 62200 642100
rect 2300 641600 62200 641800
rect 2300 641300 2500 641600
rect 2800 641300 3000 641600
rect 3300 641300 3500 641600
rect 3800 641300 58000 641600
rect 58300 641300 58500 641600
rect 58800 641300 59000 641600
rect 59300 641300 59500 641600
rect 59800 641300 60000 641600
rect 60300 641300 60500 641600
rect 60800 641300 61000 641600
rect 61300 641300 61500 641600
rect 61800 641300 62200 641600
rect 2300 641100 62200 641300
rect 2300 640800 2500 641100
rect 2800 640800 3000 641100
rect 3300 640800 3500 641100
rect 3800 640800 58000 641100
rect 58300 640800 58500 641100
rect 58800 640800 59000 641100
rect 59300 640800 59500 641100
rect 59800 640800 60000 641100
rect 60300 640800 60500 641100
rect 60800 640800 61000 641100
rect 61300 640800 61500 641100
rect 61800 640800 62200 641100
rect 2300 640600 62200 640800
rect 2300 640300 2500 640600
rect 2800 640300 3000 640600
rect 3300 640300 3500 640600
rect 3800 640300 58000 640600
rect 58300 640300 58500 640600
rect 58800 640300 59000 640600
rect 59300 640300 59500 640600
rect 59800 640300 60000 640600
rect 60300 640300 60500 640600
rect 60800 640300 61000 640600
rect 61300 640300 61500 640600
rect 61800 640300 62200 640600
rect 2300 640100 62200 640300
rect 2300 639800 2500 640100
rect 2800 639800 3000 640100
rect 3300 639800 3500 640100
rect 3800 639800 58000 640100
rect 58300 639800 58500 640100
rect 58800 639800 59000 640100
rect 59300 639800 59500 640100
rect 59800 639800 60000 640100
rect 60300 639800 60500 640100
rect 60800 639800 61000 640100
rect 61300 639800 61500 640100
rect 61800 639800 62200 640100
rect 2300 639600 62200 639800
rect 2300 639300 2500 639600
rect 2800 639300 3000 639600
rect 3300 639300 3500 639600
rect 3800 639300 58000 639600
rect 58300 639300 58500 639600
rect 58800 639300 59000 639600
rect 59300 639300 59500 639600
rect 59800 639300 60000 639600
rect 60300 639300 60500 639600
rect 60800 639300 61000 639600
rect 61300 639300 61500 639600
rect 61800 639300 62200 639600
rect 2300 639100 62200 639300
rect 2300 638800 2500 639100
rect 2800 638800 3000 639100
rect 3300 638800 3500 639100
rect 3800 638800 58000 639100
rect 58300 638800 58500 639100
rect 58800 638800 59000 639100
rect 59300 638800 59500 639100
rect 59800 638800 60000 639100
rect 60300 638800 60500 639100
rect 60800 638800 61000 639100
rect 61300 638800 61500 639100
rect 61800 638800 62200 639100
rect 2300 638600 62200 638800
rect 2300 638300 2500 638600
rect 2800 638300 3000 638600
rect 3300 638300 3500 638600
rect 3800 638300 58000 638600
rect 58300 638300 58500 638600
rect 58800 638300 59000 638600
rect 59300 638300 59500 638600
rect 59800 638300 60000 638600
rect 60300 638300 60500 638600
rect 60800 638300 61000 638600
rect 61300 638300 61500 638600
rect 61800 638300 62200 638600
rect 2300 638100 62200 638300
rect 2300 637800 2500 638100
rect 2800 637800 3000 638100
rect 3300 637800 3500 638100
rect 3800 637800 58000 638100
rect 58300 637800 58500 638100
rect 58800 637800 59000 638100
rect 59300 637800 59500 638100
rect 59800 637800 60000 638100
rect 60300 637800 60500 638100
rect 60800 637800 61000 638100
rect 61300 637800 61500 638100
rect 61800 637800 62200 638100
rect 2300 637600 62200 637800
rect 2300 637300 2500 637600
rect 2800 637300 3000 637600
rect 3300 637300 3500 637600
rect 3800 637300 58000 637600
rect 58300 637300 58500 637600
rect 58800 637300 59000 637600
rect 59300 637300 59500 637600
rect 59800 637300 60000 637600
rect 60300 637300 60500 637600
rect 60800 637300 61000 637600
rect 61300 637300 61500 637600
rect 61800 637300 62200 637600
rect 2300 637100 62200 637300
rect 2300 636800 2500 637100
rect 2800 636800 3000 637100
rect 3300 636800 3500 637100
rect 3800 636800 58000 637100
rect 58300 636800 58500 637100
rect 58800 636800 59000 637100
rect 59300 636800 59500 637100
rect 59800 636800 60000 637100
rect 60300 636800 60500 637100
rect 60800 636800 61000 637100
rect 61300 636800 61500 637100
rect 61800 636800 62200 637100
rect 2300 636600 62200 636800
rect 2300 636300 2500 636600
rect 2800 636300 3000 636600
rect 3300 636300 3500 636600
rect 3800 636300 58000 636600
rect 58300 636300 58500 636600
rect 58800 636300 59000 636600
rect 59300 636300 59500 636600
rect 59800 636300 60000 636600
rect 60300 636300 60500 636600
rect 60800 636300 61000 636600
rect 61300 636300 61500 636600
rect 61800 636300 62200 636600
rect 2300 636100 62200 636300
rect 2300 635800 2500 636100
rect 2800 635800 3000 636100
rect 3300 635800 3500 636100
rect 3800 635800 58000 636100
rect 58300 635800 58500 636100
rect 58800 635800 59000 636100
rect 59300 635800 59500 636100
rect 59800 635800 60000 636100
rect 60300 635800 60500 636100
rect 60800 635800 61000 636100
rect 61300 635800 61500 636100
rect 61800 635800 62200 636100
rect 2300 635600 62200 635800
rect 2300 635300 2500 635600
rect 2800 635300 3000 635600
rect 3300 635300 3500 635600
rect 3800 635300 58000 635600
rect 58300 635300 58500 635600
rect 58800 635300 59000 635600
rect 59300 635300 59500 635600
rect 59800 635300 60000 635600
rect 60300 635300 60500 635600
rect 60800 635300 61000 635600
rect 61300 635300 61500 635600
rect 61800 635300 62200 635600
rect 2300 635100 62200 635300
rect 2300 634800 2500 635100
rect 2800 634800 3000 635100
rect 3300 634800 3500 635100
rect 3800 634800 58000 635100
rect 58300 634800 58500 635100
rect 58800 634800 59000 635100
rect 59300 634800 59500 635100
rect 59800 634800 60000 635100
rect 60300 634800 60500 635100
rect 60800 634800 61000 635100
rect 61300 634800 61500 635100
rect 61800 634800 62200 635100
rect 2300 634600 62200 634800
rect 2300 634300 2500 634600
rect 2800 634300 3000 634600
rect 3300 634300 3500 634600
rect 3800 634300 58000 634600
rect 58300 634300 58500 634600
rect 58800 634300 59000 634600
rect 59300 634300 59500 634600
rect 59800 634300 60000 634600
rect 60300 634300 60500 634600
rect 60800 634300 61000 634600
rect 61300 634300 61500 634600
rect 61800 634300 62200 634600
rect 2300 633800 62200 634300
<< res5p73 >>
rect 38123 694981 40127 696131
rect 49193 694981 51197 696131
rect 38123 693521 40127 694671
rect 49193 693521 51197 694671
rect 535152 686823 537156 687973
rect 552212 686823 554216 687973
rect 535152 685353 537156 686503
rect 552212 685353 554216 686503
rect 41720 663310 42870 677114
rect 43270 663310 44420 677114
rect 44810 663310 45960 677114
rect 46360 663310 47510 677114
rect 541759 663768 542909 677572
rect 543279 663768 544429 677572
rect 544789 663774 545939 677578
rect 546299 663774 547449 677578
<< labels >>
flabel metal3 s 582300 677984 584800 682984 0 FreeSans 1120 0 0 0 io_analog[0]
port 36 nsew signal bidirectional
flabel metal3 s 0 680242 1700 685242 0 FreeSans 1120 0 0 0 io_analog[10]
port 37 nsew signal bidirectional
flabel metal3 s 566594 702300 571594 704800 0 FreeSans 1920 180 0 0 io_analog[1]
port 38 nsew signal bidirectional
flabel metal3 s 465394 702300 470394 704800 0 FreeSans 1920 180 0 0 io_analog[2]
port 39 nsew signal bidirectional
flabel metal3 s 68194 702300 73194 704800 0 FreeSans 1920 180 0 0 io_analog[8]
port 45 nsew signal bidirectional
flabel metal3 s 16194 702300 21194 704800 0 FreeSans 1920 180 0 0 io_analog[9]
port 46 nsew signal bidirectional
flabel metal3 s 582340 639784 584800 644584 0 FreeSans 1120 0 0 0 vccd1
port 552 nsew signal bidirectional
flabel metal3 s 582340 629784 584800 634584 0 FreeSans 1120 0 0 0 vccd1
port 553 nsew signal bidirectional
flabel metal3 s 0 643842 1660 648642 0 FreeSans 1120 0 0 0 vccd2
port 554 nsew signal bidirectional
flabel metal3 s 0 633842 1660 638642 0 FreeSans 1120 0 0 0 vccd2
port 555 nsew signal bidirectional
flabel metal3 s 0 559442 1660 564242 0 FreeSans 1120 0 0 0 vssa2
port 566 nsew signal bidirectional
flabel metal3 s 0 549442 1660 554242 0 FreeSans 1120 0 0 0 vssa2
port 567 nsew signal bidirectional
rlabel metal5 43372 670040 43372 670040 1 constant_gm_fingers_0/VSS
rlabel metal3 44392 683084 44392 683084 1 constant_gm_fingers_0/Vout
rlabel metal5 44100 683900 44100 683900 1 constant_gm_fingers_0/VDD
<< end >>
