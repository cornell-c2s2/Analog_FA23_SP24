magic
tech sky130A
timestamp 1712710044
<< metal1 >>
rect -10 -5 50 60
<< labels >>
rlabel metal1 5 10 35 50 1 test
port 1 n
<< end >>
