** sch_path: /foss/designs/Analog_FA23_SP24/flashADC/xschem/flashADC_Testing_sym_v0p4p3.sch
.lib /foss/pdks/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.include /foss/pdks/sky130A/libs.ref/sky130_fd_sc_hd/spice/sky130_fd_sc_hd.spice

.subckt flashADC_Testing_sym_v0p4p3 VFS OUT3 OUT2 OUT1 OUT0 VDD VIN CLK GND VL
*.PININFO OUT3:O OUT2:O OUT1:O OUT0:O VDD:I GND:I VIN:I CLK:I VFS:I VL:I
XR1 VL net2 VL sky130_fd_pr__res_xhigh_po_5p73 L=2.865 mult=8 m=8
XR2 net2 net1 VL sky130_fd_pr__res_xhigh_po_5p73 L=2.865 mult=8 m=8
XR3 net1 net3 VL sky130_fd_pr__res_xhigh_po_5p73 L=2.865 mult=8 m=8
XR4 net3 net4 VL sky130_fd_pr__res_xhigh_po_5p73 L=2.865 mult=8 m=8
XR5 net4 net5 VL sky130_fd_pr__res_xhigh_po_5p73 L=2.865 mult=8 m=8
XR6 net5 net6 VL sky130_fd_pr__res_xhigh_po_5p73 L=2.865 mult=8 m=8
XR7 net6 net7 VL sky130_fd_pr__res_xhigh_po_5p73 L=2.865 mult=8 m=8
XR8 net7 net8 VL sky130_fd_pr__res_xhigh_po_5p73 L=2.865 mult=8 m=8
XR9 net8 net9 VL sky130_fd_pr__res_xhigh_po_5p73 L=2.865 mult=8 m=8
XR10 net9 net10 VL sky130_fd_pr__res_xhigh_po_5p73 L=2.865 mult=8 m=8
XR11 net10 net11 VL sky130_fd_pr__res_xhigh_po_5p73 L=2.865 mult=8 m=8
XR12 net11 net12 VL sky130_fd_pr__res_xhigh_po_5p73 L=2.865 mult=8 m=8
XR13 net12 net13 VL sky130_fd_pr__res_xhigh_po_5p73 L=2.865 mult=8 m=8
XR14 net13 net14 VL sky130_fd_pr__res_xhigh_po_5p73 L=2.865 mult=8 m=8
XR15 net14 net15 VL sky130_fd_pr__res_xhigh_po_5p73 L=2.865 mult=8 m=8
XR16 net15 net16 VL sky130_fd_pr__res_xhigh_po_5p73 L=2.865 mult=8 m=8
XR18 net16 VFS VL sky130_fd_pr__res_xhigh_po_5p73 L=2.865 mult=8 m=8
* noconn #net65
* noconn #net66
* noconn #net67
* noconn #net68
* noconn #net69
* noconn #net70
* noconn #net71
* noconn #net72
* noconn #net73
* noconn #net74
* noconn #net75
* noconn #net76
* noconn #net77
* noconn #net78
* noconn #net79
* noconn #net80
x64 net47 GND GND VDD VDD net81 sky130_fd_sc_hd__buf_1
x34 net48 GND GND VDD VDD net82 sky130_fd_sc_hd__buf_1
x35 net45 GND GND VDD VDD net83 sky130_fd_sc_hd__buf_1
x36 net46 GND GND VDD VDD net84 sky130_fd_sc_hd__buf_1
x37 net43 GND GND VDD VDD net85 sky130_fd_sc_hd__buf_1
x38 net44 GND GND VDD VDD net86 sky130_fd_sc_hd__buf_1
x39 net41 GND GND VDD VDD net87 sky130_fd_sc_hd__buf_1
x40 net42 GND GND VDD VDD net88 sky130_fd_sc_hd__buf_1
x41 net39 GND GND VDD VDD net89 sky130_fd_sc_hd__buf_1
x42 net40 GND GND VDD VDD net90 sky130_fd_sc_hd__buf_1
x43 net37 GND GND VDD VDD net91 sky130_fd_sc_hd__buf_1
x44 net38 GND GND VDD VDD net92 sky130_fd_sc_hd__buf_1
x45 net35 GND GND VDD VDD net93 sky130_fd_sc_hd__buf_1
x46 net36 GND GND VDD VDD net94 sky130_fd_sc_hd__buf_1
x47 net33 GND GND VDD VDD net95 sky130_fd_sc_hd__buf_1
x48 net34 GND GND VDD VDD net96 sky130_fd_sc_hd__buf_1
x49 net31 GND GND VDD VDD net97 sky130_fd_sc_hd__buf_1
x50 net32 GND GND VDD VDD net98 sky130_fd_sc_hd__buf_1
x51 net29 GND GND VDD VDD net99 sky130_fd_sc_hd__buf_1
x52 net30 GND GND VDD VDD net100 sky130_fd_sc_hd__buf_1
x53 net27 GND GND VDD VDD net101 sky130_fd_sc_hd__buf_1
x54 net28 GND GND VDD VDD net102 sky130_fd_sc_hd__buf_1
x55 net25 GND GND VDD VDD net103 sky130_fd_sc_hd__buf_1
x56 net26 GND GND VDD VDD net104 sky130_fd_sc_hd__buf_1
x57 net23 GND GND VDD VDD net105 sky130_fd_sc_hd__buf_1
x58 net24 GND GND VDD VDD net106 sky130_fd_sc_hd__buf_1
x59 net21 GND GND VDD VDD net107 sky130_fd_sc_hd__buf_1
x60 net22 GND GND VDD VDD net108 sky130_fd_sc_hd__buf_1
x61 net19 GND GND VDD VDD net109 sky130_fd_sc_hd__buf_1
x62 net20 GND GND VDD VDD net110 sky130_fd_sc_hd__buf_1
x63 net17 GND GND VDD VDD net111 sky130_fd_sc_hd__buf_1
x65 net18 GND GND VDD VDD net112 sky130_fd_sc_hd__buf_1
x19 VDD net81 net82 net59 net80 GND RSfetsym
x20 VDD net83 net84 net60 net79 GND RSfetsym
x21 VDD net85 net86 net61 net78 GND RSfetsym
x22 VDD net87 net88 net62 net77 GND RSfetsym
x23 VDD net89 net90 net63 net76 GND RSfetsym
x24 VDD net91 net92 net64 net75 GND RSfetsym
x25 VDD net93 net94 net49 net74 GND RSfetsym
x26 VDD net95 net96 net50 net73 GND RSfetsym
x27 VDD net97 net98 net51 net72 GND RSfetsym
x28 VDD net99 net100 net52 net71 GND RSfetsym
x29 VDD net101 net102 net53 net70 GND RSfetsym
x30 VDD net103 net104 net54 net69 GND RSfetsym
x31 VDD net105 net106 net55 net68 GND RSfetsym
x32 VDD net107 net108 net56 net67 GND RSfetsym
x33 VDD net109 net110 net57 net66 GND RSfetsym
x66 VDD net111 net112 net58 net65 GND RSfetsym
x1 OUT3 VDD net59 net60 net61 net62 net63 net64 OUT2 net49 net50 VDD net51 net52 net53 net54 OUT1 net55 net56 GND net57 net58 OUT0
+ 16to4_PriorityEncoder_v0p0p1
x2 VDD net47 net48 net16 VIN IB CLK GND class_AB_v4_sym
x3 VDD net45 net46 net15 VIN IB CLK GND class_AB_v4_sym
x4 VDD net43 net44 net14 VIN IB CLK GND class_AB_v4_sym
x5 VDD net41 net42 net13 VIN IB CLK GND class_AB_v4_sym
x6 VDD net39 net40 net12 VIN IB CLK GND class_AB_v4_sym
x7 VDD net37 net38 net11 VIN IB CLK GND class_AB_v4_sym
x8 VDD net35 net36 net10 VIN IB CLK GND class_AB_v4_sym
x9 VDD net33 net34 net9 VIN IB CLK GND class_AB_v4_sym
x10 VDD net31 net32 net8 VIN IB CLK GND class_AB_v4_sym
x11 VDD net29 net30 net7 VIN IB CLK GND class_AB_v4_sym
x12 VDD net27 net28 net6 VIN IB CLK GND class_AB_v4_sym
x13 VDD net25 net26 net5 VIN IB CLK GND class_AB_v4_sym
x14 VDD net23 net24 net4 VIN IB CLK GND class_AB_v4_sym
x15 VDD net21 net22 net3 VIN IB CLK GND class_AB_v4_sym
x16 VDD net19 net20 net1 VIN IB CLK GND class_AB_v4_sym
x17 VDD net17 net18 net2 VIN IB CLK GND class_AB_v4_sym
x18 VDD IB GND PTAT_v0p0p0
.ends


.GLOBAL GND
.GLOBAL VDD
.GLOBAL VIN
.GLOBAL CLK
.GLOBAL IB
.end
