magic
tech sky130A
magscale 1 2
timestamp 1716868724
<< error_p >>
rect -317 572 -259 578
rect -125 572 -67 578
rect 67 572 125 578
rect 259 572 317 578
rect -317 538 -305 572
rect -125 538 -113 572
rect 67 538 79 572
rect 259 538 271 572
rect -317 532 -259 538
rect -125 532 -67 538
rect 67 532 125 538
rect 259 532 317 538
rect -413 -538 -355 -532
rect -221 -538 -163 -532
rect -29 -538 29 -532
rect 163 -538 221 -532
rect 355 -538 413 -532
rect -413 -572 -401 -538
rect -221 -572 -209 -538
rect -29 -572 -17 -538
rect 163 -572 175 -538
rect 355 -572 367 -538
rect -413 -578 -355 -572
rect -221 -578 -163 -572
rect -29 -578 29 -572
rect 163 -578 221 -572
rect 355 -578 413 -572
<< pwell >>
rect -599 -710 599 710
<< nmos >>
rect -399 -500 -369 500
rect -303 -500 -273 500
rect -207 -500 -177 500
rect -111 -500 -81 500
rect -15 -500 15 500
rect 81 -500 111 500
rect 177 -500 207 500
rect 273 -500 303 500
rect 369 -500 399 500
<< ndiff >>
rect -461 488 -399 500
rect -461 -488 -449 488
rect -415 -488 -399 488
rect -461 -500 -399 -488
rect -369 488 -303 500
rect -369 -488 -353 488
rect -319 -488 -303 488
rect -369 -500 -303 -488
rect -273 488 -207 500
rect -273 -488 -257 488
rect -223 -488 -207 488
rect -273 -500 -207 -488
rect -177 488 -111 500
rect -177 -488 -161 488
rect -127 -488 -111 488
rect -177 -500 -111 -488
rect -81 488 -15 500
rect -81 -488 -65 488
rect -31 -488 -15 488
rect -81 -500 -15 -488
rect 15 488 81 500
rect 15 -488 31 488
rect 65 -488 81 488
rect 15 -500 81 -488
rect 111 488 177 500
rect 111 -488 127 488
rect 161 -488 177 488
rect 111 -500 177 -488
rect 207 488 273 500
rect 207 -488 223 488
rect 257 -488 273 488
rect 207 -500 273 -488
rect 303 488 369 500
rect 303 -488 319 488
rect 353 -488 369 488
rect 303 -500 369 -488
rect 399 488 461 500
rect 399 -488 415 488
rect 449 -488 461 488
rect 399 -500 461 -488
<< ndiffc >>
rect -449 -488 -415 488
rect -353 -488 -319 488
rect -257 -488 -223 488
rect -161 -488 -127 488
rect -65 -488 -31 488
rect 31 -488 65 488
rect 127 -488 161 488
rect 223 -488 257 488
rect 319 -488 353 488
rect 415 -488 449 488
<< psubdiff >>
rect -563 640 -467 674
rect 467 640 563 674
rect -563 578 -529 640
rect 529 578 563 640
rect -563 -640 -529 -578
rect 529 -640 563 -578
rect -563 -674 -467 -640
rect 467 -674 563 -640
<< psubdiffcont >>
rect -467 640 467 674
rect -563 -578 -529 578
rect 529 -578 563 578
rect -467 -674 467 -640
<< poly >>
rect -321 572 -255 588
rect -321 538 -305 572
rect -271 538 -255 572
rect -399 500 -369 526
rect -321 522 -255 538
rect -129 572 -63 588
rect -129 538 -113 572
rect -79 538 -63 572
rect -303 500 -273 522
rect -207 500 -177 526
rect -129 522 -63 538
rect 63 572 129 588
rect 63 538 79 572
rect 113 538 129 572
rect -111 500 -81 522
rect -15 500 15 526
rect 63 522 129 538
rect 255 572 321 588
rect 255 538 271 572
rect 305 538 321 572
rect 81 500 111 522
rect 177 500 207 526
rect 255 522 321 538
rect 273 500 303 522
rect 369 500 399 526
rect -399 -522 -369 -500
rect -417 -538 -351 -522
rect -303 -526 -273 -500
rect -207 -522 -177 -500
rect -417 -572 -401 -538
rect -367 -572 -351 -538
rect -417 -588 -351 -572
rect -225 -538 -159 -522
rect -111 -526 -81 -500
rect -15 -522 15 -500
rect -225 -572 -209 -538
rect -175 -572 -159 -538
rect -225 -588 -159 -572
rect -33 -538 33 -522
rect 81 -526 111 -500
rect 177 -522 207 -500
rect -33 -572 -17 -538
rect 17 -572 33 -538
rect -33 -588 33 -572
rect 159 -538 225 -522
rect 273 -526 303 -500
rect 369 -522 399 -500
rect 159 -572 175 -538
rect 209 -572 225 -538
rect 159 -588 225 -572
rect 351 -538 417 -522
rect 351 -572 367 -538
rect 401 -572 417 -538
rect 351 -588 417 -572
<< polycont >>
rect -305 538 -271 572
rect -113 538 -79 572
rect 79 538 113 572
rect 271 538 305 572
rect -401 -572 -367 -538
rect -209 -572 -175 -538
rect -17 -572 17 -538
rect 175 -572 209 -538
rect 367 -572 401 -538
<< locali >>
rect -563 640 -467 674
rect 467 640 563 674
rect -563 578 -529 640
rect 529 578 563 640
rect -321 538 -305 572
rect -271 538 -255 572
rect -129 538 -113 572
rect -79 538 -63 572
rect 63 538 79 572
rect 113 538 129 572
rect 255 538 271 572
rect 305 538 321 572
rect -449 488 -415 504
rect -449 -504 -415 -488
rect -353 488 -319 504
rect -353 -504 -319 -488
rect -257 488 -223 504
rect -257 -504 -223 -488
rect -161 488 -127 504
rect -161 -504 -127 -488
rect -65 488 -31 504
rect -65 -504 -31 -488
rect 31 488 65 504
rect 31 -504 65 -488
rect 127 488 161 504
rect 127 -504 161 -488
rect 223 488 257 504
rect 223 -504 257 -488
rect 319 488 353 504
rect 319 -504 353 -488
rect 415 488 449 504
rect 415 -504 449 -488
rect -417 -572 -401 -538
rect -367 -572 -351 -538
rect -225 -572 -209 -538
rect -175 -572 -159 -538
rect -33 -572 -17 -538
rect 17 -572 33 -538
rect 159 -572 175 -538
rect 209 -572 225 -538
rect 351 -572 367 -538
rect 401 -572 417 -538
rect -563 -640 -529 -578
rect 529 -640 563 -578
rect -563 -674 -467 -640
rect 467 -674 563 -640
<< viali >>
rect -305 538 -271 572
rect -113 538 -79 572
rect 79 538 113 572
rect 271 538 305 572
rect -449 -488 -415 488
rect -353 -488 -319 488
rect -257 -488 -223 488
rect -161 -488 -127 488
rect -65 -488 -31 488
rect 31 -488 65 488
rect 127 -488 161 488
rect 223 -488 257 488
rect 319 -488 353 488
rect 415 -488 449 488
rect -401 -572 -367 -538
rect -209 -572 -175 -538
rect -17 -572 17 -538
rect 175 -572 209 -538
rect 367 -572 401 -538
<< metal1 >>
rect -317 572 -259 578
rect -317 538 -305 572
rect -271 538 -259 572
rect -317 532 -259 538
rect -125 572 -67 578
rect -125 538 -113 572
rect -79 538 -67 572
rect -125 532 -67 538
rect 67 572 125 578
rect 67 538 79 572
rect 113 538 125 572
rect 67 532 125 538
rect 259 572 317 578
rect 259 538 271 572
rect 305 538 317 572
rect 259 532 317 538
rect -455 488 -409 500
rect -455 -488 -449 488
rect -415 -488 -409 488
rect -455 -500 -409 -488
rect -359 488 -313 500
rect -359 -488 -353 488
rect -319 -488 -313 488
rect -359 -500 -313 -488
rect -263 488 -217 500
rect -263 -488 -257 488
rect -223 -488 -217 488
rect -263 -500 -217 -488
rect -167 488 -121 500
rect -167 -488 -161 488
rect -127 -488 -121 488
rect -167 -500 -121 -488
rect -71 488 -25 500
rect -71 -488 -65 488
rect -31 -488 -25 488
rect -71 -500 -25 -488
rect 25 488 71 500
rect 25 -488 31 488
rect 65 -488 71 488
rect 25 -500 71 -488
rect 121 488 167 500
rect 121 -488 127 488
rect 161 -488 167 488
rect 121 -500 167 -488
rect 217 488 263 500
rect 217 -488 223 488
rect 257 -488 263 488
rect 217 -500 263 -488
rect 313 488 359 500
rect 313 -488 319 488
rect 353 -488 359 488
rect 313 -500 359 -488
rect 409 488 455 500
rect 409 -488 415 488
rect 449 -488 455 488
rect 409 -500 455 -488
rect -413 -538 -355 -532
rect -413 -572 -401 -538
rect -367 -572 -355 -538
rect -413 -578 -355 -572
rect -221 -538 -163 -532
rect -221 -572 -209 -538
rect -175 -572 -163 -538
rect -221 -578 -163 -572
rect -29 -538 29 -532
rect -29 -572 -17 -538
rect 17 -572 29 -538
rect -29 -578 29 -572
rect 163 -538 221 -532
rect 163 -572 175 -538
rect 209 -572 221 -538
rect 163 -578 221 -572
rect 355 -538 413 -532
rect 355 -572 367 -538
rect 401 -572 413 -538
rect 355 -578 413 -572
<< properties >>
string FIXED_BBOX -546 -657 546 657
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 5.0 l 0.15 m 1 nf 9 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
