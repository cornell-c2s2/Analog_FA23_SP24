magic
tech sky130A
magscale 1 2
timestamp 1717181165
<< metal1 >>
rect 5200 2400 6000 3200
rect 4600 2300 6600 2400
rect 4600 1900 4700 2300
rect 6500 1900 6600 2300
rect 4600 1800 6600 1900
rect 10247 1000 10600 1077
rect 10247 300 10400 1000
rect 10500 300 10600 1000
rect 10247 183 10600 300
rect 10900 800 11700 900
rect 10900 200 11000 800
rect 11600 200 11700 800
rect 10900 100 11700 200
rect 0 -100 4600 100
rect 6600 -100 10400 100
rect 0 -300 10400 -100
rect 0 -500 4600 -300
rect 6600 -500 10400 -300
rect 0 -800 177 -500
rect 0 -1600 180 -800
rect 0 -1800 4600 -1600
rect 6600 -1800 10400 -1600
rect 0 -1900 10400 -1800
rect 3800 -2200 7400 -1900
rect 4600 -2700 6600 -2200
<< via1 >>
rect 4700 1900 6500 2300
rect 10400 300 10500 1000
rect 11000 200 11600 800
<< metal2 >>
rect 4600 2300 6600 2400
rect 4600 1900 4700 2300
rect 6500 1900 6600 2300
rect 4600 1800 6600 1900
rect 10300 1000 12000 1100
rect 10300 300 10400 1000
rect 10500 800 12000 1000
rect 10500 300 11000 800
rect 10300 200 11000 300
rect 11600 200 12000 800
rect 10500 -500 12000 200
rect 10500 -1500 10600 -500
rect 11900 -1500 12000 -500
rect 10500 -1600 12000 -1500
<< via2 >>
rect 4700 1900 6500 2300
rect 10600 -1500 11900 -500
<< metal3 >>
rect 4600 2300 6600 2400
rect 4600 1900 4700 2300
rect 6500 1900 6600 2300
rect 4600 200 6600 1900
rect 4600 -500 12000 -400
rect 4600 -1500 10600 -500
rect 11900 -1500 12000 -500
rect 4600 -1600 12000 -1500
use diode_connected_nmos  diode_connected_nmos_0
timestamp 1717119771
transform 0 1 60 -1 0 -446
box -60 -60 1254 10360
use diode_connected_nmos  diode_connected_nmos_1
timestamp 1717119771
transform 0 1 60 -1 0 1254
box -60 -60 1254 10360
<< labels >>
flabel metal1 5200 -2700 6000 -1900 0 FreeSans 800 0 0 0 VSS
port 1 n
flabel metal1 5200 2400 6000 3200 0 FreeSans 800 0 0 0 VDD
port 3 n
flabel metal1 10900 100 11700 900 0 FreeSans 800 0 0 0 VIO
port 2 n
<< end >>
