* NGSPICE file created from frontAnalog_v0p0p1_flat.ext - technology: sky130A

.subckt frontAnalog_v0p0p1_flatten VDD GND VN VIN CLK Q IB
X0 RSfetsym_0.S a_5187_3971# GND.t29 GND.t21 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1 class_AB_v3_sym_0.VOP.t1 CLK.t0 class_AB_v3_sym_0.VON.t2 VDD.t19 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X2 class_AB_v3_sym_0.VOP.t3 class_AB_v3_sym_0.VON.t4 a_3332_2594# GND.t11 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X3 RSfetsym_0.R a_5187_2451# VDD.t3 VDD.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X4 RSfetsym_0.R a_5187_2451# GND.t22 GND.t21 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X5 GND.t10 RSfetsym_0.QN.t5 a_7641_3047# GND.t9 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X6 w_3064_2980# VIN.t0 a_1694_2534# GND.t42 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X7 VIN.t1 w_3064_3602# error sky130_fd_pr__cap_var_lvt w=2 l=0.18
X8 w_3064_3602# CLK.t1 class_AB_v3_sym_0.VOP.t0 VDD.t12 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X9 VDD.t11 RSfetsym_0.R RSfetsym_0.x1.Y VDD.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X10 VDD.t33 RSfetsym_0.S RSfetsym_0.QN.t4 VDD.t28 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.25
X11 RSfetsym_0.x1.Y RSfetsym_0.R VDD.t10 VDD.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12 class_AB_v3_sym_0.VON.t3 CLK.t2 w_3064_2980# VDD.t18 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X13 RSfetsym_0.QN.t1 Q.t5 VDD.t22 VDD.t0 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.3
X14 a_1694_2534# IB.t0 GND.t1 GND.t0 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X15 RSfetsym_0.QN.t0 RSfetsym_0.x1.Y GND.t20 GND.t19 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.25
X16 Q.t1 RSfetsym_0.QN.t6 VDD.t1 VDD.t0 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.3
X17 VDD.t9 RSfetsym_0.R RSfetsym_0.x1.Y VDD.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X18 a_1694_2534# VN.t0 w_3064_3602# GND.t4 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X19 GND.t31 Q.t6 a_7642_3560# GND.t30 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X20 VDD.t32 RSfetsym_0.S RSfetsym_0.x2.Y VDD.t26 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X21 RSfetsym_0.x2.Y RSfetsym_0.S VDD.t31 VDD.t26 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X22 VDD.t15 class_AB_v3_sym_0.VOP.t4 a_5187_3971# VDD.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X23 GND.t3 class_AB_v3_sym_0.VOP.t5 a_5187_3971# GND.t2 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X24 VDD.t30 RSfetsym_0.S RSfetsym_0.x2.Y VDD.t26 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X25 RSfetsym_0.QN.t3 RSfetsym_0.S VDD.t29 VDD.t28 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.25
X26 class_AB_v3_sym_0.VON.t0 class_AB_v3_sym_0.VOP.t6 a_3332_2594# GND.t8 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X27 GND.t40 RSfetsym_0.S RSfetsym_0.x2.Y GND.t39 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X28 GND.t28 RSfetsym_0.R RSfetsym_0.x1.Y GND.t23 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X29 GND.t5 class_AB_v3_sym_0.VON.t5 a_5187_2451# GND.t2 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X30 RSfetsym_0.x2.Y RSfetsym_0.S GND.t38 GND.t37 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X31 VDD.t25 class_AB_v3_sym_0.VON.t6 a_5187_2451# VDD.t24 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X32 RSfetsym_0.x1.Y RSfetsym_0.R GND.t27 GND.t23 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X33 VDD.t16 CLK.t3 w_3064_3602# GND.t6 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X34 VDD.t8 RSfetsym_0.R Q.t4 VDD.t4 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.25
X35 a_1694_2534# IB.t1 GND.t16 GND.t15 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X36 GND.t36 RSfetsym_0.S RSfetsym_0.x2.Y GND.t35 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X37 RSfetsym_0.x1.Y RSfetsym_0.R VDD.t7 VDD.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X38 GND.t26 RSfetsym_0.R RSfetsym_0.x1.Y GND.t23 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X39 a_7641_3047# RSfetsym_0.R Q.t2 GND.t25 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X40 VDD.t17 CLK.t4 w_3064_2980# GND.t14 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X41 RSfetsym_0.x2.Y RSfetsym_0.S VDD.t27 VDD.t26 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X42 class_AB_v3_sym_0.VON.t1 class_AB_v3_sym_0.VOP.t7 VDD.t13 VDD.t12 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X43 Q.t3 RSfetsym_0.R VDD.t5 VDD.t4 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.25
X44 VDD.t23 class_AB_v3_sym_0.VON.t7 class_AB_v3_sym_0.VOP.t2 VDD.t18 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X45 a_7642_3560# RSfetsym_0.S RSfetsym_0.QN.t2 GND.t34 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.315 ps=2.72 w=1 l=0.15
X46 VN.t1 w_3064_2980# error sky130_fd_pr__cap_var_lvt w=2 l=0.18
X47 Q.t0 RSfetsym_0.x2.Y GND.t18 GND.t17 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.25
X48 RSfetsym_0.x2.Y RSfetsym_0.S GND.t33 GND.t32 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X49 a_3332_2594# CLK.t5 GND.t13 GND.t12 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X50 RSfetsym_0.S a_5187_3971# VDD.t21 VDD.t20 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X51 RSfetsym_0.x1.Y RSfetsym_0.R GND.t24 GND.t23 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
R0 GND.n289 GND.n288 18594.9
R1 GND.t32 GND.n229 3790.39
R2 GND.t21 GND.n19 2572.31
R3 GND.n290 GND.n289 1839.93
R4 GND.n127 GND.n126 1773
R5 GND.n285 GND.n284 1559.14
R6 GND.n129 GND.n127 1384.79
R7 GND.n206 GND.n204 1384.79
R8 GND.n295 GND.n283 1153.03
R9 GND.n230 GND 1147.86
R10 GND.n62 GND.n57 1077.71
R11 GND.n62 GND.n58 1077.71
R12 GND.n41 GND.n36 1077.71
R13 GND.n40 GND.n37 1077.71
R14 GND.n63 GND.n56 1077.71
R15 GND GND.t23 1058.96
R16 GND.n63 GND.n55 1054.53
R17 GND.n151 GND.n149 915.471
R18 GND.n137 GND.n136 915.471
R19 GND.n198 GND.n197 915.471
R20 GND.n212 GND.n209 841.244
R21 GND.n317 GND.n310 778.15
R22 GND.n317 GND.n311 778.15
R23 GND.n278 GND.n274 778.15
R24 GND.n278 GND.n277 778.15
R25 GND.n151 GND.n150 521.471
R26 GND.n119 GND 484.329
R27 GND.n301 GND.n282 480.913
R28 GND.n212 GND.n210 473.865
R29 GND.n74 GND.n73 356.401
R30 GND.t39 GND.t37 352
R31 GND.t37 GND.t35 352
R32 GND.t35 GND.t32 352
R33 GND.t0 GND.n70 252.906
R34 GND.n73 GND.t0 226.601
R35 GND.n51 GND.t15 226.601
R36 GND.n47 GND.n46 225.946
R37 GND.n81 GND.n79 224.4
R38 GND.n54 GND.n53 209.695
R39 GND.n83 GND.n78 204.424
R40 GND.n293 GND.n287 203.294
R41 GND.n293 GND.n292 203.294
R42 GND.n94 GND.t28 193.933
R43 GND.n232 GND.t40 193.933
R44 GND.n103 GND.t24 192.982
R45 GND.n246 GND.t33 192.982
R46 GND.n263 GND.n262 185.514
R47 GND GND.t2 185.418
R48 GND.t19 GND.n119 185.314
R49 GND.t17 GND.n174 185.137
R50 GND.n89 GND.n83 183.47
R51 GND GND.t39 171.81
R52 GND.n308 GND.n281 153.601
R53 GND.n309 GND.n308 153.601
R54 GND.n35 GND.n34 137.827
R55 GND.n90 GND.n69 136.23
R56 GND.n157 GND.n156 135.422
R57 GND.n54 GND.n50 135.38
R58 GND.n20 GND.t21 123.612
R59 GND.n111 GND.n110 121.112
R60 GND.n243 GND.n242 121.112
R61 GND.t2 GND.n354 120.669
R62 GND.n181 GND.n180 115.201
R63 GND.n183 GND.n182 115.201
R64 GND.t8 GND.t12 111.784
R65 GND.n15 GND.n14 109.394
R66 GND.n5 GND.n4 107.24
R67 GND.t8 GND.n316 107.028
R68 GND.n81 GND.n80 92.4005
R69 GND.n148 GND.n147 90.3534
R70 GND.n208 GND.n207 90.3534
R71 GND.n169 GND.n168 86.1558
R72 GND.n227 GND.n226 86.1558
R73 GND.n34 GND.n33 78.6829
R74 GND.n280 GND.n273 78.6829
R75 GND.n50 GND.n49 78.6829
R76 GND.n320 GND.n319 78.6829
R77 GND.n294 GND.n293 74.9181
R78 GND.n319 GND.n309 70.7205
R79 GND.n61 GND.n59 70.024
R80 GND.n61 GND.n60 70.024
R81 GND.n42 GND.n35 70.024
R82 GND.n39 GND.n38 70.024
R83 GND.n64 GND.n54 70.024
R84 GND.n281 GND.n280 67.5205
R85 GND.t6 GND.n10 59.6186
R86 GND.n152 GND.n148 59.4829
R87 GND.n65 GND.n42 57.977
R88 GND.n65 GND.n64 57.224
R89 GND.n213 GND.n208 54.66
R90 GND.t14 GND.n23 51.7278
R91 GND.n319 GND.n318 50.5605
R92 GND.n280 GND.n279 50.5605
R93 GND.n27 GND.n26 46.2978
R94 GND.n323 GND.n322 45.1897
R95 GND.n90 GND.n89 44.6176
R96 GND.n344 GND.n13 42.8187
R97 GND.n66 GND.n30 39.6805
R98 GND.n153 GND.n152 33.8829
R99 GND.n14 GND.t22 33.462
R100 GND.n14 GND.t5 33.462
R101 GND.n4 GND.t29 33.462
R102 GND.n4 GND.t3 33.462
R103 GND.n214 GND.n213 30.7897
R104 GND.n330 GND.n325 28.9511
R105 GND.n202 GND.n201 28.8193
R106 GND.n143 GND.n142 26.7111
R107 GND.n110 GND.t27 24.9236
R108 GND.n110 GND.t26 24.9236
R109 GND.n242 GND.t38 24.9236
R110 GND.n242 GND.t36 24.9236
R111 GND.n47 GND.n45 23.7843
R112 GND.n66 GND.n65 23.4245
R113 GND.n215 GND.n214 22.9087
R114 GND.n184 GND.n183 22.4086
R115 GND.n154 GND.n153 22.0429
R116 GND.n95 GND.n94 21.8358
R117 GND.n300 GND.n299 20.6255
R118 GND.n13 GND.n12 19.2005
R119 GND.n118 GND.t31 17.475
R120 GND.n334 GND.t13 17.4601
R121 GND.n118 GND.t10 17.4528
R122 GND.n233 GND.n232 16.1887
R123 GND.n265 GND.n264 14.7755
R124 GND.n269 GND.n267 14.7755
R125 GND.n106 GND.n105 9.3005
R126 GND.n96 GND.n95 9.3005
R127 GND.n98 GND.n97 9.3005
R128 GND.n108 GND.n107 9.3005
R129 GND.n249 GND.n248 9.3005
R130 GND.n234 GND.n233 9.3005
R131 GND.n170 GND.n169 9.3005
R132 GND.n164 GND.n163 9.3005
R133 GND.n155 GND.n154 9.3005
R134 GND.n162 GND.n161 9.3005
R135 GND.n144 GND.n143 9.3005
R136 GND.n135 GND.n134 9.3005
R137 GND.n133 GND.n132 9.3005
R138 GND.n124 GND.n123 9.3005
R139 GND.n179 GND.n178 9.3005
R140 GND.n226 GND.n225 9.3005
R141 GND.n216 GND.n215 9.3005
R142 GND.n194 GND.n193 9.3005
R143 GND.n203 GND.n202 9.3005
R144 GND.n185 GND.n184 9.3005
R145 GND.n192 GND.n191 9.3005
R146 GND.n302 GND.n301 9.3005
R147 GND.n301 GND.n300 9.3005
R148 GND.n171 GND.t20 8.70904
R149 GND.n177 GND.t18 8.70236
R150 GND.t30 GND.t9 8.20945
R151 GND.n15 GND 8.05791
R152 GND.n26 GND.n25 7.90638
R153 GND.n308 GND.n307 6.5285
R154 GND.n349 GND 5.64756
R155 GND.n126 GND.n125 5.62907
R156 GND.n333 GND.n330 5.1205
R157 GND.n19 GND.n18 4.83274
R158 GND.n94 GND 4.66821
R159 GND.n104 GND.n103 4.6505
R160 GND.n232 GND.n231 4.6505
R161 GND.n247 GND.n246 4.6505
R162 GND.n100 GND.n99 4.5005
R163 GND.n109 GND.n102 4.5005
R164 GND.n238 GND.n237 4.5005
R165 GND.n251 GND.n245 4.5005
R166 GND.n91 GND.t1 4.41708
R167 GND.n92 GND.t16 4.35136
R168 GND.n112 GND.n111 3.03311
R169 GND.n253 GND.n243 3.03311
R170 GND.n6 GND.n5 3.03311
R171 GND.n350 GND.n349 3.03311
R172 GND.n17 GND 3.0005
R173 GND.n87 GND.n84 2.2005
R174 GND.n315 GND.n314 1.93119
R175 GND.n316 GND.n315 1.93119
R176 GND.n340 GND.n259 1.71871
R177 GND.n304 GND.n303 1.64041
R178 GND.n303 GND.n302 1.63319
R179 GND.n245 GND.n244 1.12991
R180 GND.n305 GND.n67 1.10116
R181 GND.n309 GND.n266 0.9605
R182 GND.n281 GND.n270 0.9605
R183 GND.n69 GND.n68 0.795337
R184 GND GND.n340 0.652549
R185 GND.n225 GND.n224 0.533636
R186 GND.n342 GND.n341 0.523375
R187 GND.n325 GND.n324 0.436742
R188 GND.n324 GND.n323 0.436742
R189 GND.n171 GND.n170 0.425574
R190 GND.n216 GND.n203 0.38056
R191 GND.n192 GND.n190 0.377583
R192 GND.n237 GND.n236 0.376971
R193 GND.n188 GND.n185 0.3755
R194 GND.n133 GND.n131 0.373417
R195 GND.n131 GND.n124 0.373417
R196 GND.n182 GND.n181 0.366214
R197 GND.n223 GND.n222 0.355857
R198 GND.n17 GND 0.354667
R199 GND.n165 GND.n122 0.345738
R200 GND.n27 GND.n22 0.321569
R201 GND.n345 GND.n344 0.321569
R202 GND.n343 GND.n342 0.314812
R203 GND.n155 GND.n144 0.313
R204 GND.n17 GND.n15 0.295052
R205 GND.n179 GND.n177 0.290381
R206 GND.n194 GND.n192 0.24425
R207 GND.n173 GND.n172 0.243155
R208 GND.n135 GND.n133 0.238893
R209 GND.n258 GND.n115 0.224247
R210 GND.n164 GND.n162 0.200996
R211 GND.n353 GND.n0 0.197423
R212 GND.n224 GND.n223 0.181736
R213 GND.n224 GND.n173 0.17675
R214 GND.n196 GND.n194 0.171333
R215 GND.n203 GND.n200 0.16925
R216 GND.n162 GND.n160 0.164786
R217 GND.n160 GND.n155 0.164786
R218 GND.n218 GND.n216 0.159429
R219 GND.n144 GND.n141 0.148714
R220 GND.n139 GND.n135 0.148714
R221 GND.n93 GND.n92 0.142154
R222 GND.n295 GND.n294 0.131784
R223 GND.n298 GND.n295 0.13084
R224 GND.n297 GND.n296 0.126877
R225 GND.n298 GND.n297 0.125988
R226 GND.n231 GND.n230 0.122064
R227 GND.n172 GND.n165 0.112135
R228 GND.n213 GND.n212 0.10956
R229 GND.n212 GND.n211 0.10956
R230 GND.n152 GND.n151 0.10956
R231 GND.n151 GND.t30 0.10956
R232 GND.n276 GND.n275 0.10956
R233 GND.t11 GND.n276 0.10956
R234 GND.n313 GND.n312 0.10956
R235 GND.t8 GND.n313 0.10956
R236 GND.n318 GND.n317 0.10956
R237 GND.n317 GND.t8 0.10956
R238 GND.n44 GND.n43 0.10956
R239 GND.n45 GND.n44 0.10956
R240 GND.n261 GND.n260 0.10956
R241 GND.n262 GND.n261 0.10956
R242 GND.n278 GND.t11 0.10956
R243 GND.n279 GND.n278 0.10956
R244 GND.n330 GND.n329 0.104537
R245 GND.n329 GND.n328 0.104537
R246 GND.n172 GND.n171 0.102333
R247 GND.n228 GND.n227 0.0944005
R248 GND.n229 GND.n228 0.0944005
R249 GND.n168 GND.n167 0.0944005
R250 GND.n167 GND.n166 0.0944005
R251 GND.n106 GND.n104 0.0921667
R252 GND.n249 GND.n247 0.0891364
R253 GND.n343 GND.n27 0.08745
R254 GND.n344 GND.n343 0.0868625
R255 GND.n259 GND.n258 0.0845572
R256 GND.n96 GND 0.0775833
R257 GND.n234 GND 0.0675455
R258 GND.n12 GND.n11 0.0636886
R259 GND.n11 GND.t6 0.0636886
R260 GND.n25 GND.n24 0.0636886
R261 GND.n24 GND.t14 0.0636886
R262 GND.n42 GND.n41 0.0636886
R263 GND.n41 GND.t42 0.0636886
R264 GND.n62 GND.n61 0.0636886
R265 GND.t4 GND.n62 0.0636886
R266 GND.t42 GND.n40 0.0636886
R267 GND.n40 GND.n39 0.0636886
R268 GND.n64 GND.n63 0.0636886
R269 GND.n63 GND.t4 0.0636886
R270 GND.n78 GND.n77 0.0636886
R271 GND.n77 GND.n76 0.0636886
R272 GND.n259 GND 0.060284
R273 GND.n21 GND.n20 0.0588369
R274 GND.n113 GND.n109 0.0582982
R275 GND.n240 GND.n239 0.05675
R276 GND.n253 GND.n252 0.0532741
R277 GND.n247 GND 0.0527727
R278 GND.n273 GND.n272 0.0525185
R279 GND.n272 GND.n271 0.0525185
R280 GND.n33 GND.n32 0.0525185
R281 GND.n32 GND.n31 0.0525185
R282 GND.n321 GND.n320 0.0525185
R283 GND.n322 GND.n321 0.0525185
R284 GND.n49 GND.n48 0.0525185
R285 GND.n48 GND.n47 0.0525185
R286 GND.n327 GND.n326 0.0525185
R287 GND.n328 GND.n327 0.0525185
R288 GND.n83 GND.n82 0.0523204
R289 GND.n82 GND.n81 0.0523204
R290 GND.n241 GND.n238 0.0516364
R291 GND.n173 GND.n118 0.0494583
R292 GND.n254 GND.n241 0.0493636
R293 GND.n114 GND.n101 0.0486039
R294 GND.n104 GND 0.0484167
R295 GND.n252 GND.n251 0.0483725
R296 GND.n93 GND.n91 0.0483051
R297 GND.n207 GND.n206 0.0425017
R298 GND.n206 GND.n205 0.0425017
R299 GND.n147 GND.n146 0.0425017
R300 GND.n146 GND.n145 0.0425017
R301 GND.n8 GND.n7 0.0415714
R302 GND.n345 GND.n9 0.0406786
R303 GND.n92 GND 0.0386944
R304 GND.n165 GND.n164 0.0345278
R305 GND.n118 GND.n115 0.0337917
R306 GND.n101 GND.n100 0.0335935
R307 GND.n335 GND.n334 0.0307537
R308 GND.n3 GND.n2 0.0208901
R309 GND.n6 GND.n3 0.0208901
R310 GND.n351 GND.n350 0.0208901
R311 GND.n21 GND.n17 0.0200011
R312 GND.n231 GND 0.0198182
R313 GND.n352 GND.n351 0.0195603
R314 GND.n235 GND.n234 0.0186818
R315 GND.n307 GND.n306 0.0176904
R316 GND.n341 GND 0.0172857
R317 GND.n100 GND.n98 0.0171667
R318 GND.n250 GND.n249 0.0164091
R319 GND.n339 GND.n337 0.0152059
R320 GND.n292 GND.n291 0.015169
R321 GND.n291 GND.n290 0.015169
R322 GND.n266 GND.n265 0.015169
R323 GND.n265 GND.n263 0.015169
R324 GND.n287 GND.n286 0.015169
R325 GND.n286 GND.n285 0.015169
R326 GND.n86 GND.n85 0.015169
R327 GND.n87 GND.n86 0.015169
R328 GND.n72 GND.n71 0.015169
R329 GND.n73 GND.n72 0.015169
R330 GND.n270 GND.n269 0.015169
R331 GND.n269 GND.n268 0.015169
R332 GND.n53 GND.n52 0.015169
R333 GND.n52 GND.n51 0.015169
R334 GND.n89 GND.n88 0.0144432
R335 GND.n88 GND.n87 0.0144432
R336 GND.n109 GND.n108 0.0140417
R337 GND.n348 GND.n347 0.0138596
R338 GND.n17 GND.n16 0.0120741
R339 GND.n223 GND.n179 0.0112143
R340 GND.n16 GND 0.0111481
R341 GND.n341 GND.n93 0.0097322
R342 GND.n350 GND.n348 0.00783909
R343 GND.n2 GND.n1 0.00739975
R344 GND.n141 GND.n139 0.00585714
R345 GND.n306 GND.n305 0.00507317
R346 GND.n108 GND.n106 0.00466667
R347 GND.n190 GND.n188 0.00466667
R348 GND.n255 GND.n117 0.00425
R349 GND.n333 GND.n332 0.00420666
R350 GND.n332 GND.n331 0.00420666
R351 GND.n139 GND.n138 0.00396756
R352 GND.n200 GND.n199 0.00396756
R353 GND.n258 GND.n257 0.00395031
R354 GND.n138 GND.n137 0.0039133
R355 GND.n137 GND.t34 0.0039133
R356 GND.n199 GND.n198 0.0039133
R357 GND.n198 GND.t25 0.0039133
R358 GND.n254 GND.n253 0.00390909
R359 GND.n251 GND.n250 0.00390909
R360 GND.n222 GND.n221 0.0034846
R361 GND.n221 GND.n220 0.00343883
R362 GND.n220 GND.n219 0.00343883
R363 GND.n159 GND.n158 0.00343883
R364 GND.n158 GND.n157 0.00343883
R365 GND.n113 GND.n112 0.00308428
R366 GND.n117 GND.n116 0.003
R367 GND.n200 GND.n196 0.00258333
R368 GND.n257 GND.n256 0.00245833
R369 GND.n222 GND.n218 0.00228571
R370 GND.n347 GND 0.00217027
R371 GND.n188 GND.n187 0.00183506
R372 GND.n187 GND.n186 0.00181454
R373 GND.n130 GND.n129 0.00181454
R374 GND.n129 GND.n128 0.00181454
R375 GND.n300 GND.n298 0.001708
R376 GND.n238 GND.n235 0.00163636
R377 GND.n98 GND.n96 0.00154167
R378 GND.n305 GND.n304 0.00150729
R379 GND.n335 GND.n333 0.00150234
R380 GND.n336 GND.n335 0.00150164
R381 GND.n345 GND.n8 0.00139286
R382 GND.n352 GND.n346 0.00138653
R383 GND.n176 GND.n175 0.00131092
R384 GND.n175 GND.t17 0.00131092
R385 GND.n121 GND.n120 0.00131092
R386 GND.n120 GND.t19 0.00131092
R387 GND.n22 GND.n21 0.00103916
R388 GND.n342 GND.n67 0.00101312
R389 GND.n67 GND.n66 0.00100714
R390 GND.n114 GND.n113 0.00100095
R391 GND.n339 GND.n338 0.00100064
R392 GND.n346 GND.n6 0.000943262
R393 GND.n90 GND.n75 0.000826763
R394 GND.n75 GND.n74 0.000826763
R395 GND.n30 GND.n29 0.000756235
R396 GND.n29 GND.n28 0.000756235
R397 GND.n241 GND.n240 0.000544755
R398 GND.n196 GND.n195 0.000530553
R399 GND.n218 GND.n217 0.00052846
R400 GND.n141 GND.n140 0.00052846
R401 GND.n160 GND.n159 0.0005264
R402 GND.n131 GND.n130 0.000512627
R403 GND.n190 GND.n189 0.000512369
R404 GND.n122 GND.n121 0.000507826
R405 GND.n177 GND.n176 0.000507826
R406 GND.n354 GND.n353 0.000505544
R407 GND.n115 GND.n114 0.000504863
R408 GND.n337 GND.n336 0.000504005
R409 GND.n340 GND.n339 0.000501449
R410 GND.n256 GND.n255 0.000501292
R411 GND.n255 GND.n254 0.000501292
R412 GND.n353 GND.n352 0.000500915
R413 GND.n91 GND.n90 0.000500526
R414 GND.n346 GND.n345 0.000500286
R415 CLK.t3 CLK.t2 344.122
R416 CLK.n2 CLK.t5 232.299
R417 CLK.n5 CLK.t4 182.915
R418 CLK.n5 CLK.t3 182.91
R419 CLK.t4 CLK.n4 182.769
R420 CLK.n0 CLK.t1 161.262
R421 CLK.n6 CLK.t0 159.958
R422 CLK.n6 CLK.n5 0.56781
R423 CLK.n7 CLK.n6 0.428385
R424 CLK.n7 CLK 0.12425
R425 CLK.n7 CLK 0.0636313
R426 CLK CLK.n7 0.0484798
R427 CLK.n1 CLK.n0 0.0178077
R428 CLK.n4 CLK.n1 0.00531334
R429 CLK.n4 CLK.n3 0.00224847
R430 CLK.n3 CLK.n2 0.00100535
R431 class_AB_v3_sym_0.VON.n2 class_AB_v3_sym_0.VON.t6 260.322
R432 class_AB_v3_sym_0.VON.n4 class_AB_v3_sym_0.VON.t4 233.888
R433 class_AB_v3_sym_0.VON.n2 class_AB_v3_sym_0.VON.t5 175.169
R434 class_AB_v3_sym_0.VON.n3 class_AB_v3_sym_0.VON.t7 159.725
R435 class_AB_v3_sym_0.VON.n1 class_AB_v3_sym_0.VON.t0 17.4109
R436 class_AB_v3_sym_0.VON.n0 class_AB_v3_sym_0.VON.n2 9.75129
R437 class_AB_v3_sym_0.VON.n1 class_AB_v3_sym_0.VON.t1 9.6027
R438 class_AB_v3_sym_0.VON.n0 class_AB_v3_sym_0.VON 2.33338
R439 class_AB_v3_sym_0.VON.n5 class_AB_v3_sym_0.VON.t2 8.40929
R440 class_AB_v3_sym_0.VON.n3 class_AB_v3_sym_0.VON.t3 8.06629
R441 class_AB_v3_sym_0.VON.n4 class_AB_v3_sym_0.VON.n3 1.73501
R442 class_AB_v3_sym_0.VON.n1 class_AB_v3_sym_0.VON.n4 0.99025
R443 class_AB_v3_sym_0.VON.n5 class_AB_v3_sym_0.VON.n1 0.853186
R444 class_AB_v3_sym_0.VON class_AB_v3_sym_0.VON.n0 0.349517
R445 class_AB_v3_sym_0.VON class_AB_v3_sym_0.VON.n5 0.24425
R446 class_AB_v3_sym_0.VOP.n1 class_AB_v3_sym_0.VOP.t4 260.322
R447 class_AB_v3_sym_0.VOP.n4 class_AB_v3_sym_0.VOP.t6 233.929
R448 class_AB_v3_sym_0.VOP.n1 class_AB_v3_sym_0.VOP.t5 175.169
R449 class_AB_v3_sym_0.VOP.n3 class_AB_v3_sym_0.VOP.t7 160.416
R450 class_AB_v3_sym_0.VOP.n2 class_AB_v3_sym_0.VOP.t3 17.4109
R451 class_AB_v3_sym_0.VOP.n2 class_AB_v3_sym_0.VOP.t2 10.2053
R452 class_AB_v3_sym_0.VOP.n0 class_AB_v3_sym_0.VOP 2.78715
R453 class_AB_v3_sym_0.VOP.n0 class_AB_v3_sym_0.VOP.n1 9.09103
R454 class_AB_v3_sym_0.VOP.n6 class_AB_v3_sym_0.VOP.t1 7.94569
R455 class_AB_v3_sym_0.VOP.n3 class_AB_v3_sym_0.VOP.t0 7.55846
R456 class_AB_v3_sym_0.VOP.n5 class_AB_v3_sym_0.VOP.n4 1.4614
R457 class_AB_v3_sym_0.VOP.n4 class_AB_v3_sym_0.VOP.n3 1.19626
R458 class_AB_v3_sym_0.VOP.n6 class_AB_v3_sym_0.VOP.n5 0.836961
R459 class_AB_v3_sym_0.VOP class_AB_v3_sym_0.VOP.n0 0.390342
R460 class_AB_v3_sym_0.VOP.n5 class_AB_v3_sym_0.VOP.n2 0.154668
R461 class_AB_v3_sym_0.VOP class_AB_v3_sym_0.VOP.n6 0.08175
R462 VDD.n138 VDD.n127 2565.88
R463 VDD.n143 VDD.n127 2565.88
R464 VDD.n160 VDD.n159 2565.88
R465 VDD.n192 VDD.n174 2565.88
R466 VDD.n192 VDD.n175 2565.88
R467 VDD.n90 VDD.n59 2082.55
R468 VDD.n40 VDD.n20 2080.64
R469 VDD.n88 VDD.n58 2015.29
R470 VDD.n44 VDD.n24 2015.29
R471 VDD.n147 VDD.n129 1997.65
R472 VDD.n147 VDD.n130 1997.65
R473 VDD.n183 VDD.n173 1997.65
R474 VDD.n178 VDD.n173 1997.65
R475 VDD.n160 VDD.n154 1814.12
R476 VDD.n163 VDD.n162 1598.82
R477 VDD.n44 VDD.n43 1514.12
R478 VDD.n135 VDD.n123 1440
R479 VDD.n148 VDD.n125 1440
R480 VDD.n194 VDD.n169 1422.35
R481 VDD.n179 VDD.n170 1422.35
R482 VDD.n59 VDD.n22 1231.76
R483 VDD.n111 VDD.n20 1228.24
R484 VDD.n111 VDD.n21 1224.71
R485 VDD.n22 VDD.n21 1224.71
R486 VDD.n64 VDD.n21 1153.33
R487 VDD.n181 VDD.n179 1143.53
R488 VDD.n141 VDD.n125 1125.88
R489 VDD.n102 VDD.n64 1072.94
R490 VDD.n64 VDD.n16 1069.41
R491 VDD.n135 VDD.n134 1051.76
R492 VDD.n185 VDD.n169 1051.76
R493 VDD.n105 VDD.n104 861.178
R494 VDD.n165 VDD.n154 751.765
R495 VDD.n60 VDD.n58 723.529
R496 VDD.n26 VDD.n24 720
R497 VDD.n41 VDD.t28 632.183
R498 VDD.n23 VDD.n20 593.144
R499 VDD.n26 VDD.n23 593.144
R500 VDD.n224 VDD.t7 584.644
R501 VDD.n210 VDD.t27 584.644
R502 VDD.n109 VDD.n59 576.668
R503 VDD.n109 VDD.n60 576.668
R504 VDD.n138 VDD.n129 568.236
R505 VDD.n141 VDD.n130 568.236
R506 VDD.n143 VDD.n130 568.236
R507 VDD.n134 VDD.n129 568.236
R508 VDD.n185 VDD.n183 568.236
R509 VDD.n178 VDD.n175 568.236
R510 VDD.n181 VDD.n178 568.236
R511 VDD.n183 VDD.n174 568.236
R512 VDD.n90 VDD.n89 481.226
R513 VDD.n136 VDD.n126 473.839
R514 VDD.t18 VDD.n128 473.839
R515 VDD.n193 VDD.n171 468.033
R516 VDD.t12 VDD.n172 468.033
R517 VDD.n55 VDD.n26 370.589
R518 VDD.n105 VDD.n60 370.589
R519 VDD.t0 VDD.t28 333.365
R520 VDD.t0 VDD.t4 333.365
R521 VDD.t0 VDD.n24 298.82
R522 VDD.t0 VDD.n58 298.82
R523 VDD.n140 VDD.n139 273.695
R524 VDD.n144 VDD.n140 273.695
R525 VDD.n158 VDD.n153 273.695
R526 VDD.n158 VDD.n157 273.695
R527 VDD.n191 VDD.n176 273.695
R528 VDD.n191 VDD.n190 273.695
R529 VDD.n146 VDD.n131 213.083
R530 VDD.n146 VDD.n145 213.083
R531 VDD.n188 VDD.n187 213.083
R532 VDD.n189 VDD.n188 213.083
R533 VDD.n180 VDD.n172 189.304
R534 VDD.n179 VDD.n177 185
R535 VDD.n179 VDD.n172 185
R536 VDD.n169 VDD.n167 185
R537 VDD.n171 VDD.n169 185
R538 VDD.n43 VDD.n28 185
R539 VDD.n142 VDD.n128 183.496
R540 VDD.n222 VDD.n221 180.994
R541 VDD.n219 VDD.n217 180.994
R542 VDD.t26 VDD.n232 174.632
R543 VDD.n157 VDD.n155 170.542
R544 VDD.n35 VDD.n19 167.234
R545 VDD.n92 VDD.n61 166.812
R546 VDD.n202 VDD.n201 165.767
R547 VDD.n2 VDD.n1 165.767
R548 VDD.n45 VDD.n28 161.506
R549 VDD.n87 VDD.n74 159.143
R550 VDD.n137 VDD.n136 159.108
R551 VDD.n184 VDD.n171 159.108
R552 VDD.n46 VDD.n45 158.776
R553 VDD.n25 VDD.n16 155.294
R554 VDD.n213 VDD.t11 151.123
R555 VDD.n215 VDD.t32 151.123
R556 VDD.n231 VDD.t6 146.691
R557 VDD.n87 VDD.n86 143.435
R558 VDD.t19 VDD.n156 136.591
R559 VDD.n43 VDD.n42 135.117
R560 VDD.n61 VDD.n18 131.388
R561 VDD.n112 VDD.n19 131.012
R562 VDD.n113 VDD.n18 130.636
R563 VDD.n113 VDD.n112 130.636
R564 VDD.n161 VDD.n159 129.691
R565 VDD.t14 VDD 126.02
R566 VDD.n182 VDD.n177 121.977
R567 VDD.n110 VDD.t0 121.114
R568 VDD.t0 VDD.n57 121.114
R569 VDD.n132 VDD.n124 120.094
R570 VDD.n114 VDD.n113 116.267
R571 VDD.n133 VDD.n122 112.189
R572 VDD.n186 VDD.n167 112.189
R573 VDD.n115 VDD.n114 102.721
R574 VDD.n101 VDD.n17 102.721
R575 VDD.t24 VDD 99.5973
R576 VDD.n79 VDD.n76 92.5005
R577 VDD.n194 VDD.n170 91.7652
R578 VDD.n166 VDD.n155 91.343
R579 VDD.n8 VDD.t14 89.1694
R580 VDD.n8 VDD.t20 81.2688
R581 VDD.n106 VDD.n63 80.5087
R582 VDD.n54 VDD.n15 80.2452
R583 VDD.n149 VDD.n124 76.5328
R584 VDD.n148 VDD.n123 74.1181
R585 VDD.n150 VDD.n122 71.6136
R586 VDD.n197 VDD.t24 70.4844
R587 VDD.n242 VDD.n153 66.2808
R588 VDD.n177 VDD.n168 65.0929
R589 VDD.n197 VDD.t2 64.3553
R590 VDD.n52 VDD.n19 63.2691
R591 VDD.n53 VDD.n52 63.2691
R592 VDD.n108 VDD.n61 61.5116
R593 VDD.n108 VDD.n107 61.5116
R594 VDD.n139 VDD.n131 60.6123
R595 VDD.n145 VDD.n132 60.6123
R596 VDD.n145 VDD.n144 60.6123
R597 VDD.n133 VDD.n131 60.6123
R598 VDD.n187 VDD.n176 60.6123
R599 VDD.n190 VDD.n189 60.6123
R600 VDD.n189 VDD.n182 60.6123
R601 VDD.n187 VDD.n186 60.6123
R602 VDD.n195 VDD.n167 58.0325
R603 VDD.n78 VDD.n77 55.4672
R604 VDD.n79 VDD.n75 55.4672
R605 VDD.n232 VDD 54.4858
R606 VDD.n242 VDD.n241 50.1034
R607 VDD.t6 VDD.n230 49.1183
R608 VDD.n46 VDD.n27 47.0405
R609 VDD.n51 VDD.n50 45.7605
R610 VDD.n35 VDD.n31 45.7605
R611 VDD.n30 VDD.n28 45.4405
R612 VDD.n54 VDD.n53 39.5299
R613 VDD.n107 VDD.n106 39.5299
R614 VDD.n240 VDD.n166 38.9491
R615 VDD.n92 VDD.n91 37.3765
R616 VDD.n74 VDD.n71 37.3765
R617 VDD.n201 VDD.t3 36.1587
R618 VDD.n201 VDD.t25 36.1587
R619 VDD.n1 VDD.t21 36.1587
R620 VDD.n1 VDD.t15 36.1587
R621 VDD VDD.n231 34.927
R622 VDD.n193 VDD.t12 30.1961
R623 VDD.n222 VDD.n211 28.2358
R624 VDD.n223 VDD.n222 28.2358
R625 VDD.n219 VDD.n216 28.2358
R626 VDD.n219 VDD.n218 28.2358
R627 VDD.n221 VDD.t10 26.5955
R628 VDD.n221 VDD.t9 26.5955
R629 VDD.n217 VDD.t31 26.5955
R630 VDD.n217 VDD.t30 26.5955
R631 VDD.t18 VDD.n126 24.3893
R632 VDD.n213 VDD.n211 22.2123
R633 VDD.n224 VDD.n223 22.2123
R634 VDD.n216 VDD.n215 22.2123
R635 VDD.n218 VDD.n210 22.2123
R636 VDD.n202 VDD.n200 22.2123
R637 VDD.n233 VDD.t26 20.9587
R638 VDD.n53 VDD.n51 20.5934
R639 VDD.n107 VDD.n62 17.109
R640 VDD.n32 VDD.t33 14.2962
R641 VDD.n12 VDD.t29 14.2955
R642 VDD.n95 VDD.t8 14.2865
R643 VDD.n83 VDD.t5 14.2864
R644 VDD.n117 VDD.t22 14.2849
R645 VDD.n99 VDD.t1 14.2849
R646 VDD.n115 VDD.n15 14.0805
R647 VDD.n101 VDD.n63 13.7605
R648 VDD.n195 VDD.n194 9.3005
R649 VDD.n194 VDD.n193 9.3005
R650 VDD.n93 VDD.n92 9.3005
R651 VDD.n74 VDD.n73 9.3005
R652 VDD.n77 VDD.n68 9.3005
R653 VDD.n51 VDD.n13 9.3005
R654 VDD.n36 VDD.n35 9.3005
R655 VDD.n80 VDD.n79 8.88939
R656 VDD.n241 VDD.n240 7.49764
R657 VDD.n196 VDD.t13 7.15136
R658 VDD.n151 VDD.t23 7.14897
R659 VDD.n200 VDD 6.4005
R660 VDD.n250 VDD 6.4005
R661 VDD.n225 VDD.n210 4.6505
R662 VDD.n225 VDD.n224 4.6505
R663 VDD.n220 VDD.n219 4.6505
R664 VDD.n222 VDD.n220 4.6505
R665 VDD.n218 VDD.n209 4.6505
R666 VDD.n216 VDD.n212 4.6505
R667 VDD.n215 VDD.n214 4.6505
R668 VDD.n223 VDD.n209 4.6505
R669 VDD.n212 VDD.n211 4.6505
R670 VDD.n214 VDD.n213 4.6505
R671 VDD.n200 VDD.n199 4.6505
R672 VDD.n251 VDD.n250 4.6505
R673 VDD.n3 VDD.n2 4.6505
R674 VDD.n97 VDD.n67 4.5005
R675 VDD.n97 VDD.n62 4.5005
R676 VDD.n97 VDD.n96 4.5005
R677 VDD.n206 VDD.n205 4.5005
R678 VDD.n229 VDD.n208 4.5005
R679 VDD.n229 VDD.n228 4.5005
R680 VDD.n226 VDD.n208 4.5005
R681 VDD.n244 VDD.t16 4.35136
R682 VDD.n238 VDD.t17 4.35136
R683 VDD.n203 VDD.n202 3.96837
R684 VDD.n40 VDD.n29 3.52991
R685 VDD.n47 VDD.n46 3.03311
R686 VDD.n252 VDD 3.0005
R687 VDD.n150 VDD.n149 2.98717
R688 VDD.n195 VDD.n168 2.72837
R689 VDD.n207 VDD.n206 2.2278
R690 VDD.n118 VDD.n117 1.51475
R691 VDD.n237 VDD.n196 1.49778
R692 VDD.n86 VDD.n75 1.42272
R693 VDD.n239 VDD.n238 1.25748
R694 VDD.n77 VDD.n62 1.06717
R695 VDD.n245 VDD.n151 1.00783
R696 VDD.n50 VDD.n27 0.9605
R697 VDD.n39 VDD.n31 0.6405
R698 VDD.n34 VDD.n33 0.590778
R699 VDD.n234 VDD.n233 0.589191
R700 VDD.n94 VDD.n69 0.514389
R701 VDD.n32 VDD.n11 0.471224
R702 VDD.n119 VDD.n12 0.467504
R703 VDD.n198 VDD 0.411214
R704 VDD.n99 VDD.n98 0.410606
R705 VDD.n84 VDD.n83 0.399706
R706 VDD.n95 VDD.n94 0.398914
R707 VDD.n83 VDD.n69 0.398403
R708 VDD.n33 VDD.n32 0.368458
R709 VDD.n34 VDD.n12 0.361663
R710 VDD.n96 VDD.n95 0.357683
R711 VDD.n80 VDD.n78 0.356056
R712 VDD.n5 VDD 0.355332
R713 VDD.n238 VDD.n237 0.349136
R714 VDD.n38 VDD.n33 0.340142
R715 VDD.n114 VDD.n17 0.3205
R716 VDD.n39 VDD.n30 0.3205
R717 VDD.n237 VDD.n236 0.314572
R718 VDD.n245 VDD.n244 0.311403
R719 VDD.n37 VDD.n36 0.296036
R720 VDD.n93 VDD.n70 0.261214
R721 VDD.n73 VDD.n72 0.261214
R722 VDD.n91 VDD.n71 0.2565
R723 VDD.n82 VDD.n81 0.251889
R724 VDD.n100 VDD.n65 0.248103
R725 VDD.n116 VDD.n14 0.247868
R726 VDD.n84 VDD.n67 0.232755
R727 VDD.n76 VDD.n68 0.217167
R728 VDD.n236 VDD.n235 0.215221
R729 VDD.n48 VDD.n47 0.204667
R730 VDD.n49 VDD.n13 0.199111
R731 VDD.n204 VDD.n203 0.192557
R732 VDD.n199 VDD.n198 0.192167
R733 VDD.n233 VDD.n205 0.180841
R734 VDD.n106 VDD.n105 0.164944
R735 VDD.n105 VDD.n57 0.164944
R736 VDD.n56 VDD.n55 0.159358
R737 VDD.n55 VDD.n54 0.15889
R738 VDD.n247 VDD.n121 0.141376
R739 VDD.n120 VDD.n119 0.117306
R740 VDD.n135 VDD.n122 0.104784
R741 VDD.n136 VDD.n135 0.104784
R742 VDD.n246 VDD.n245 0.0972991
R743 VDD.n199 VDD 0.0963333
R744 VDD VDD.n247 0.0948131
R745 VDD.n243 VDD.n152 0.0945934
R746 VDD.n5 VDD 0.0902606
R747 VDD.n226 VDD.n207 0.0864543
R748 VDD.n229 VDD.n207 0.0864543
R749 VDD.n120 VDD.n11 0.0855148
R750 VDD.n251 VDD.n249 0.0832206
R751 VDD.n73 VDD.n69 0.07913
R752 VDD.n94 VDD.n93 0.0773443
R753 VDD.n36 VDD.n34 0.0755586
R754 VDD.n247 VDD.n246 0.0710611
R755 VDD.n236 VDD.n204 0.0705353
R756 VDD.n125 VDD.n124 0.0694784
R757 VDD.n128 VDD.n125 0.0694784
R758 VDD.n234 VDD 0.064463
R759 VDD.n220 VDD.n212 0.0643889
R760 VDD.n220 VDD.n209 0.0643889
R761 VDD.n225 VDD.n209 0.0643889
R762 VDD.n118 VDD.n13 0.0588333
R763 VDD VDD.n212 0.0525833
R764 VDD.n228 VDD 0.0470278
R765 VDD.n235 VDD.n121 0.04574
R766 VDD.n252 VDD.n251 0.0409412
R767 VDD.n226 VDD.n205 0.0395625
R768 VDD.n5 VDD.n4 0.0372647
R769 VDD.n47 VDD.n11 0.0364409
R770 VDD.n7 VDD.n5 0.0361152
R771 VDD.n98 VDD.n97 0.0357224
R772 VDD.n30 VDD.n29 0.034445
R773 VDD VDD.n225 0.0324444
R774 VDD.n117 VDD.n116 0.0294474
R775 VDD.n100 VDD.n99 0.0287895
R776 VDD.n96 VDD.n66 0.0282778
R777 VDD.t0 VDD.n109 0.0282694
R778 VDD.n109 VDD.n108 0.0282694
R779 VDD.t0 VDD.n23 0.0282694
R780 VDD.n52 VDD.n23 0.0282694
R781 VDD.n139 VDD.n138 0.0265784
R782 VDD.n138 VDD.n137 0.0265784
R783 VDD.n141 VDD.n132 0.0265784
R784 VDD.n142 VDD.n141 0.0265784
R785 VDD.n144 VDD.n143 0.0265784
R786 VDD.n143 VDD.n142 0.0265784
R787 VDD.n137 VDD.n134 0.0265784
R788 VDD.n134 VDD.n133 0.0265784
R789 VDD.n160 VDD.n153 0.0265784
R790 VDD.t19 VDD.n160 0.0265784
R791 VDD.n162 VDD.n157 0.0265784
R792 VDD.n176 VDD.n174 0.0265784
R793 VDD.n184 VDD.n174 0.0265784
R794 VDD.n190 VDD.n175 0.0265784
R795 VDD.n180 VDD.n175 0.0265784
R796 VDD.n182 VDD.n181 0.0265784
R797 VDD.n181 VDD.n180 0.0265784
R798 VDD.n186 VDD.n185 0.0265784
R799 VDD.n185 VDD.n184 0.0265784
R800 VDD.n249 VDD.n248 0.0261194
R801 VDD.n42 VDD.n29 0.0257918
R802 VDD.n162 VDD.n161 0.02576
R803 VDD.n164 VDD.n163 0.0228205
R804 VDD.n163 VDD.n155 0.0223212
R805 VDD.n228 VDD.n227 0.0182941
R806 VDD.n208 VDD.n206 0.0178611
R807 VDD.n104 VDD.n103 0.0168386
R808 VDD.n56 VDD.n25 0.0168372
R809 VDD.n25 VDD.n15 0.0163404
R810 VDD.n104 VDD.n63 0.0163404
R811 VDD.n9 VDD.n8 0.0149834
R812 VDD.n239 VDD.n152 0.0145797
R813 VDD.n67 VDD.n66 0.0143889
R814 VDD.n248 VDD 0.0131689
R815 VDD.n214 VDD 0.0123056
R816 VDD.n246 VDD 0.0118881
R817 VDD.n244 VDD.n243 0.0111456
R818 VDD.n42 VDD.n41 0.0101514
R819 VDD.n165 VDD.n164 0.0101
R820 VDD.n149 VDD.n148 0.0096003
R821 VDD.n148 VDD.t18 0.0096003
R822 VDD.n166 VDD.n165 0.0096003
R823 VDD.t12 VDD.n170 0.00959985
R824 VDD.n170 VDD.n168 0.00959985
R825 VDD.n88 VDD.n87 0.0084202
R826 VDD.n45 VDD.n44 0.0084202
R827 VDD.n44 VDD.t28 0.0084202
R828 VDD.n22 VDD.n18 0.0084202
R829 VDD.n110 VDD.n22 0.0084202
R830 VDD.n112 VDD.n111 0.0084202
R831 VDD.n111 VDD.n110 0.0084202
R832 VDD.n89 VDD.n88 0.00702894
R833 VDD.n3 VDD.n0 0.00693382
R834 VDD.n85 VDD.n82 0.00605556
R835 VDD.n140 VDD.n127 0.00505015
R836 VDD.t18 VDD.n127 0.00505015
R837 VDD.n147 VDD.n146 0.00505015
R838 VDD.t18 VDD.n147 0.00505015
R839 VDD.n159 VDD.n158 0.00505015
R840 VDD.n192 VDD.n191 0.00505015
R841 VDD.t12 VDD.n192 0.00505015
R842 VDD.t12 VDD.n173 0.00505015
R843 VDD.n188 VDD.n173 0.00505015
R844 VDD.n97 VDD.n68 0.00466667
R845 VDD.n49 VDD.n48 0.00466667
R846 VDD.n38 VDD.n37 0.00466667
R847 VDD.n204 VDD.n197 0.00364862
R848 VDD.n89 VDD.t4 0.00289124
R849 VDD.n10 VDD.n7 0.00240766
R850 VDD.n249 VDD.n3 0.00233824
R851 VDD VDD.n252 0.00233824
R852 VDD.n161 VDD.t19 0.00231811
R853 VDD.n72 VDD.n70 0.00228571
R854 VDD.n40 VDD.n39 0.00221302
R855 VDD.n41 VDD.n40 0.00221302
R856 VDD.n39 VDD.n38 0.00221271
R857 VDD.n78 VDD.n76 0.00220611
R858 VDD.n48 VDD.n27 0.0022058
R859 VDD.n91 VDD.n70 0.0022058
R860 VDD.n91 VDD.n90 0.00212475
R861 VDD.n27 VDD.n24 0.00212475
R862 VDD.n78 VDD.n58 0.00212475
R863 VDD.n235 VDD.n234 0.00207613
R864 VDD.n103 VDD.n102 0.00194704
R865 VDD.n81 VDD.n76 0.00188889
R866 VDD.n232 VDD.n206 0.00175592
R867 VDD.n231 VDD.n206 0.00175592
R868 VDD.n249 VDD.n10 0.00162613
R869 VDD.n203 VDD.n198 0.00161113
R870 VDD.n230 VDD.n229 0.00151809
R871 VDD.n230 VDD.n206 0.00149567
R872 VDD.n196 VDD.n195 0.00148913
R873 VDD.n115 VDD.n16 0.00145131
R874 VDD.n57 VDD.n16 0.00145131
R875 VDD.n116 VDD.n115 0.00145112
R876 VDD.n102 VDD.n101 0.00144714
R877 VDD.n101 VDD.n100 0.00144695
R878 VDD.n65 VDD.n14 0.00139286
R879 VDD.n240 VDD.n154 0.00133663
R880 VDD.n156 VDD.n154 0.00133663
R881 VDD.n150 VDD.n123 0.00114565
R882 VDD.n126 VDD.n123 0.00114565
R883 VDD.n85 VDD.n84 0.00113805
R884 VDD.n227 VDD.n226 0.00108642
R885 VDD.n98 VDD.n66 0.00105202
R886 VDD.n57 VDD.n56 0.00100293
R887 VDD.n7 VDD.n6 0.00100132
R888 VDD.n227 VDD.n206 0.00100033
R889 VDD.n164 VDD.n156 0.00100021
R890 VDD.n103 VDD.n57 0.0010001
R891 VDD.n82 VDD.n75 0.000594432
R892 VDD.n119 VDD.n118 0.000558569
R893 VDD.n86 VDD.n85 0.000555817
R894 VDD.n114 VDD.n14 0.000534058
R895 VDD.n240 VDD.n239 0.000523376
R896 VDD.n50 VDD.n49 0.000516232
R897 VDD.n37 VDD.n31 0.000516232
R898 VDD.n81 VDD.n80 0.000515622
R899 VDD.n243 VDD.n242 0.000514451
R900 VDD.n72 VDD.n71 0.000505865
R901 VDD.n10 VDD.n9 0.000504381
R902 VDD.n65 VDD.n17 0.000503792
R903 VDD.n241 VDD.n152 0.000501164
R904 VDD.n151 VDD.n150 0.000500414
R905 VDD.n121 VDD.n120 0.000500121
R906 RSfetsym_0.QN.n1 RSfetsym_0.QN.t5 117.511
R907 RSfetsym_0.QN.n1 RSfetsym_0.QN.t6 110.698
R908 RSfetsym_0.QN.n2 RSfetsym_0.QN.t2 19.1963
R909 RSfetsym_0.QN.n3 RSfetsym_0.QN.t1 14.5206
R910 RSfetsym_0.QN.n0 RSfetsym_0.QN.t4 14.283
R911 RSfetsym_0.QN.n0 RSfetsym_0.QN.t3 14.283
R912 RSfetsym_0.QN RSfetsym_0.QN.t0 9.14075
R913 RSfetsym_0.QN.n2 RSfetsym_0.QN.n1 0.826818
R914 RSfetsym_0.QN RSfetsym_0.QN.n0 0.74645
R915 RSfetsym_0.QN.n0 RSfetsym_0.QN.n3 0.249509
R916 RSfetsym_0.QN.n3 RSfetsym_0.QN.n2 0.0968646
R917 VIN.n0 VIN.t1 167.326
R918 VIN.n0 VIN.t0 92.4649
R919 VIN.n1 VIN 4.6255
R920 VIN VIN.n1 1.6255
R921 VIN.n1 VIN.n0 1.49913
R922 Q.n0 Q.t6 117.314
R923 Q.n0 Q.t5 110.852
R924 Q.n1 Q.t2 17.6181
R925 Q.n3 Q.t1 14.2865
R926 Q.n5 Q.t4 14.283
R927 Q.n5 Q.t3 14.283
R928 Q.n7 Q.t0 8.77592
R929 Q.n7 Q.n6 1.20426
R930 Q Q.n7 0.405405
R931 Q.n4 Q.n3 0.300251
R932 Q.n2 Q.n0 0.159555
R933 Q.n6 Q.n5 0.106617
R934 Q.n4 Q.n2 0.0796167
R935 Q.n6 Q.n4 0.0480595
R936 Q.n2 Q.n1 0.000504658
R937 IB.n0 IB.t1 91.7714
R938 IB.n0 IB.t0 91.3136
R939 IB IB.n0 45.9747
R940 VN.n0 VN.t1 167.365
R941 VN.n0 VN.t0 92.4496
R942 VN.n1 VN.n0 2.07493
R943 VN.n1 VN 0.12425
R944 VN VN.n1 0.121824
C0 a_3332_2594# a_1694_2534# 0.015f
C1 IB w_3064_2980# 0.0217f
C2 w_3064_2980# class_AB_v3_sym_0.VOP 0.0988f
C3 VIN VN 0.108f
C4 RSfetsym_0.x2.Y VDD 0.926f
C5 RSfetsym_0.QN RSfetsym_0.S 2.28f
C6 IB class_AB_v3_sym_0.VOP 0.0352f
C7 w_3064_3602# VDD 0.679f
C8 CLK w_3064_3602# 0.57f
C9 a_1694_2534# VN 0.278f
C10 RSfetsym_0.R RSfetsym_0.S 0.143f
C11 a_1694_2534# VIN 0.265f
C12 RSfetsym_0.QN RSfetsym_0.x1.Y 0.17f
C13 w_3064_3602# class_AB_v3_sym_0.VON 0.0792f
C14 RSfetsym_0.R RSfetsym_0.x1.Y 0.883f
C15 a_3332_2594# w_3064_3602# 0.149f
C16 VDD RSfetsym_0.S 3.48f
C17 w_3064_2980# VDD 0.676f
C18 a_7641_3047# RSfetsym_0.QN 0.418f
C19 CLK w_3064_2980# 0.535f
C20 VDD RSfetsym_0.x1.Y 0.733f
C21 RSfetsym_0.R RSfetsym_0.QN 0.378f
C22 w_3064_3602# VN 0.795f
C23 a_5187_3971# RSfetsym_0.S 0.119f
C24 a_7641_3047# RSfetsym_0.R 0.28f
C25 VIN w_3064_3602# 0.864f
C26 IB VDD 0.151f
C27 w_3064_2980# class_AB_v3_sym_0.VON 0.659f
C28 CLK IB 0.0545f
C29 class_AB_v3_sym_0.VOP VDD 2.94f
C30 CLK class_AB_v3_sym_0.VOP 2.61f
C31 a_3332_2594# w_3064_2980# 0.12f
C32 IB class_AB_v3_sym_0.VON 0.0784f
C33 a_1694_2534# w_3064_3602# 0.359f
C34 class_AB_v3_sym_0.VOP class_AB_v3_sym_0.VON 3.16f
C35 a_5187_3971# class_AB_v3_sym_0.VOP 0.214f
C36 RSfetsym_0.QN VDD 2.54f
C37 a_3332_2594# IB 0.0848f
C38 a_7641_3047# VDD 0.0171f
C39 a_3332_2594# class_AB_v3_sym_0.VOP 0.461f
C40 RSfetsym_0.R a_5187_2451# 0.121f
C41 RSfetsym_0.R VDD 3.14f
C42 w_3064_2980# VN 0.75f
C43 w_3064_2980# VIN 0.73f
C44 RSfetsym_0.R class_AB_v3_sym_0.VON 0.0301f
C45 IB VN 0.0484f
C46 a_7642_3560# RSfetsym_0.S 0.436f
C47 IB VIN 0.0464f
C48 class_AB_v3_sym_0.VOP VN 0.22f
C49 VIN class_AB_v3_sym_0.VOP 0.626f
C50 a_1694_2534# w_3064_2980# 0.394f
C51 VDD a_5187_2451# 0.215f
C52 CLK VDD 2.47f
C53 IB a_1694_2534# 0.462f
C54 class_AB_v3_sym_0.VON a_5187_2451# 0.212f
C55 class_AB_v3_sym_0.VON VDD 3.18f
C56 a_5187_3971# VDD 0.215f
C57 CLK class_AB_v3_sym_0.VON 1.79f
C58 a_3332_2594# VDD 0.117f
C59 CLK a_3332_2594# 0.235f
C60 RSfetsym_0.x2.Y RSfetsym_0.S 0.526f
C61 RSfetsym_0.QN a_7642_3560# 0.255f
C62 a_3332_2594# class_AB_v3_sym_0.VON 1.24f
C63 RSfetsym_0.x2.Y RSfetsym_0.x1.Y 0.0254f
C64 w_3064_2980# w_3064_3602# 0.327f
C65 VN VDD 0.355f
C66 VIN VDD 0.453f
C67 CLK VN 0.588f
C68 CLK VIN 0.35f
C69 IB w_3064_3602# 0.0216f
C70 RSfetsym_0.R m3_6460_2180# 0.139f
C71 class_AB_v3_sym_0.VOP w_3064_3602# 0.658f
C72 class_AB_v3_sym_0.VON VN 0.577f
C73 VIN class_AB_v3_sym_0.VON 0.133f
C74 a_7642_3560# VDD 0.0207f
C75 a_1694_2534# VDD 0.0261f
C76 RSfetsym_0.QN RSfetsym_0.x2.Y 0.018f
C77 CLK a_1694_2534# 0.0136f
C78 a_3332_2594# VN 0.203f
C79 a_3332_2594# VIN 0.174f
C80 RSfetsym_0.S RSfetsym_0.x1.Y 0.182f
C81 RSfetsym_0.R RSfetsym_0.x2.Y 0.0923f
C82 VDD m3_6460_2180# 1.28f
C83 class_AB_v3_sym_0.VOP RSfetsym_0.S 0.0236f
C84 VN GND 2.25f
C85 VIN GND 2.03f
C86 CLK GND 4.33f
C87 IB GND 3.13f
C88 VDD GND 39.7f
C89 m3_6460_2180# GND 0.228f $ **FLOATING
C90 a_7641_3047# GND 0.561f
C91 a_5187_2451# GND 0.319f
C92 RSfetsym_0.x2.Y GND 1.53f
C93 RSfetsym_0.R GND 5.4f
C94 a_7642_3560# GND 0.555f
C95 RSfetsym_0.x1.Y GND 1.93f
C96 RSfetsym_0.QN GND 6.35f
C97 RSfetsym_0.S GND 5.09f
C98 a_5187_3971# GND 0.318f
C99 a_3332_2594# GND 1.18f
C100 a_1694_2534# GND 2.61f
C101 class_AB_v3_sym_0.VOP GND 2.65f
C102 class_AB_v3_sym_0.VON GND 2.47f
C103 w_3064_2980# GND 2.69f
C104 w_3064_3602# GND 2.69f
C105 Q.t6 GND 0.0237f
C106 Q.t5 GND 0.0725f
C107 Q.n0 GND 1.14f
C108 Q.t2 GND 0.0144f
C109 Q.n1 GND 0.341f
C110 Q.n2 GND 0.15f
C111 Q.t1 GND 0.0243f
C112 Q.n3 GND 0.226f
C113 Q.n4 GND 0.242f
C114 Q.t4 GND 0.0243f
C115 Q.t3 GND 0.0243f
C116 Q.n5 GND 0.333f
C117 Q.n6 GND 0.316f
C118 Q.t0 GND 0.0267f
C119 Q.n7 GND 0.864f
C120 RSfetsym_0.QN.n0 GND 0.993f
C121 RSfetsym_0.QN.t5 GND 0.0317f
C122 RSfetsym_0.QN.t6 GND 0.0933f
C123 RSfetsym_0.QN.n1 GND 1.47f
C124 RSfetsym_0.QN.n2 GND 0.587f
C125 RSfetsym_0.QN.t1 GND 0.0363f
C126 RSfetsym_0.QN.n3 GND 0.622f
C127 RSfetsym_0.QN.t4 GND 0.0317f
C128 RSfetsym_0.QN.t3 GND 0.0317f
C129 RSfetsym_0.QN.t0 GND 0.0558f
C130 VDD.n2 GND 0.0136f
C131 VDD.n4 GND 0.0105f
C132 VDD.n5 GND 0.101f
C133 VDD.n7 GND 0.0247f
C134 VDD.t20 GND 0.073f
C135 VDD.t14 GND 0.0275f
C136 VDD.n8 GND 0.0181f
C137 VDD.n9 GND 0.0509f
C138 VDD.n11 GND 0.0601f
C139 VDD.n12 GND 0.117f
C140 VDD.n14 GND 0.0223f
C141 VDD.n18 GND 0.0117f
C142 VDD.n19 GND 0.0164f
C143 VDD.n20 GND 0.0189f
C144 VDD.n21 GND 0.0184f
C145 VDD.n22 GND 0.0117f
C146 VDD.t28 GND 0.151f
C147 VDD.n24 GND 0.0889f
C148 VDD.n28 GND 0.0105f
C149 VDD.n32 GND 0.111f
C150 VDD.n33 GND 0.0385f
C151 VDD.n34 GND 0.0325f
C152 VDD.n35 GND 0.0108f
C153 VDD.n40 GND 0.0103f
C154 VDD.n41 GND 0.128f
C155 VDD.n43 GND 0.01f
C156 VDD.n44 GND 0.017f
C157 VDD.n45 GND 0.0144f
C158 VDD.n46 GND 0.0106f
C159 VDD.n57 GND 0.186f
C160 VDD.t4 GND 0.151f
C161 VDD.n58 GND 0.0889f
C162 VDD.n59 GND 0.0191f
C163 VDD.n61 GND 0.0165f
C164 VDD.n64 GND 0.0169f
C165 VDD.n65 GND 0.0223f
C166 VDD.n67 GND 0.125f
C167 VDD.n69 GND 0.0342f
C168 VDD.n74 GND 0.0113f
C169 VDD.n83 GND 0.123f
C170 VDD.n84 GND 0.148f
C171 VDD.n87 GND 0.0136f
C172 VDD.n88 GND 0.0195f
C173 VDD.n90 GND 0.148f
C174 VDD.n92 GND 0.0116f
C175 VDD.n94 GND 0.034f
C176 VDD.n95 GND 0.119f
C177 VDD.n96 GND 0.0167f
C178 VDD.n98 GND 0.0193f
C179 VDD.n99 GND 0.0734f
C180 VDD.n100 GND 0.0342f
C181 VDD.t0 GND 0.43f
C182 VDD.n110 GND 0.186f
C183 VDD.n111 GND 0.0116f
C184 VDD.n112 GND 0.0116f
C185 VDD.n113 GND 0.018f
C186 VDD.n114 GND 0.0121f
C187 VDD.n116 GND 0.0343f
C188 VDD.n117 GND 0.0728f
C189 VDD.n118 GND 0.0202f
C190 VDD.n119 GND 0.063f
C191 VDD.n120 GND 0.329f
C192 VDD.n121 GND 1.16f
C193 VDD.t23 GND 0.0116f
C194 VDD.n122 GND 0.0177f
C195 VDD.n124 GND 0.0167f
C196 VDD.n125 GND 0.0125f
C197 VDD.n126 GND 0.173f
C198 VDD.n127 GND 0.0246f
C199 VDD.n128 GND 0.228f
C200 VDD.n129 GND 0.0154f
C201 VDD.n130 GND 0.0154f
C202 VDD.n131 GND 0.0154f
C203 VDD.n135 GND 0.0121f
C204 VDD.n136 GND 0.22f
C205 VDD.n137 GND 0.0979f
C206 VDD.n138 GND 0.0153f
C207 VDD.n139 GND 0.0153f
C208 VDD.n140 GND 0.0246f
C209 VDD.n142 GND 0.106f
C210 VDD.n143 GND 0.0153f
C211 VDD.n144 GND 0.0153f
C212 VDD.n145 GND 0.0154f
C213 VDD.n146 GND 0.019f
C214 VDD.n147 GND 0.019f
C215 VDD.t18 GND 0.173f
C216 VDD.n149 GND 0.0217f
C217 VDD.n150 GND 0.0215f
C218 VDD.n151 GND 0.747f
C219 VDD.t16 GND 0.0114f
C220 VDD.n152 GND 0.0565f
C221 VDD.n153 GND 0.0157f
C222 VDD.n154 GND 0.0124f
C223 VDD.n155 GND 0.0121f
C224 VDD.n156 GND 0.173f
C225 VDD.n157 GND 0.0205f
C226 VDD.n158 GND 0.0246f
C227 VDD.n159 GND 0.198f
C228 VDD.n160 GND 0.0216f
C229 VDD.t19 GND 0.217f
C230 VDD.n162 GND 0.0205f
C231 VDD.n163 GND 0.0124f
C232 VDD.n166 GND 0.0144f
C233 VDD.t17 GND 0.0114f
C234 VDD.t13 GND 0.0118f
C235 VDD.n167 GND 0.0198f
C236 VDD.n168 GND 0.0307f
C237 VDD.n169 GND 0.012f
C238 VDD.n171 GND 0.218f
C239 VDD.n172 GND 0.228f
C240 VDD.n173 GND 0.019f
C241 VDD.n174 GND 0.0153f
C242 VDD.n175 GND 0.0153f
C243 VDD.n176 GND 0.0153f
C244 VDD.n177 GND 0.0177f
C245 VDD.n178 GND 0.0154f
C246 VDD.n179 GND 0.0125f
C247 VDD.n180 GND 0.108f
C248 VDD.n183 GND 0.0154f
C249 VDD.n184 GND 0.0979f
C250 VDD.n187 GND 0.0154f
C251 VDD.n188 GND 0.019f
C252 VDD.n189 GND 0.0154f
C253 VDD.n190 GND 0.0153f
C254 VDD.n191 GND 0.0246f
C255 VDD.n192 GND 0.0246f
C256 VDD.t12 GND 0.173f
C257 VDD.n193 GND 0.173f
C258 VDD.n195 GND 0.222f
C259 VDD.n196 GND 0.71f
C260 VDD.t2 GND 0.0971f
C261 VDD.t24 GND 0.0339f
C262 VDD.n197 GND 0.177f
C263 VDD.n198 GND 0.0113f
C264 VDD.n202 GND 0.0136f
C265 VDD.n203 GND 0.0116f
C266 VDD.n204 GND 0.147f
C267 VDD.n206 GND 0.0231f
C268 VDD.n208 GND 0.0137f
C269 VDD.n209 GND 0.0163f
C270 VDD.n212 GND 0.0148f
C271 VDD.t32 GND 0.0108f
C272 VDD.t11 GND 0.0108f
C273 VDD.n213 GND 0.0132f
C274 VDD.n214 GND 0.0111f
C275 VDD.n215 GND 0.0132f
C276 VDD.n220 GND 0.0163f
C277 VDD.n225 GND 0.0122f
C278 VDD.n230 GND 0.113f
C279 VDD.t6 GND 0.0474f
C280 VDD.n231 GND 0.0492f
C281 VDD.n232 GND 0.0606f
C282 VDD.t26 GND 0.0469f
C283 VDD.n233 GND 0.432f
C284 VDD.n234 GND 2.27f
C285 VDD.n235 GND 1.36f
C286 VDD.n236 GND 1.53f
C287 VDD.n237 GND 0.422f
C288 VDD.n238 GND 0.285f
C289 VDD.n239 GND 0.115f
C290 VDD.n241 GND 0.0109f
C291 VDD.n242 GND 0.015f
C292 VDD.n243 GND 0.0547f
C293 VDD.n244 GND 0.169f
C294 VDD.n245 GND 0.419f
C295 VDD.n246 GND 0.0969f
C296 VDD.n247 GND 1.07f
C297 VDD.n248 GND 0.0338f
C298 VDD.n249 GND 0.0269f
C299 class_AB_v3_sym_0.VOP.n0 GND 0.132f
C300 class_AB_v3_sym_0.VOP.t4 GND 0.0265f
C301 class_AB_v3_sym_0.VOP.t5 GND 0.0165f
C302 class_AB_v3_sym_0.VOP.n1 GND 0.0537f
C303 class_AB_v3_sym_0.VOP.t1 GND 0.141f
C304 class_AB_v3_sym_0.VOP.t2 GND 0.438f
C305 class_AB_v3_sym_0.VOP.t3 GND 0.0184f
C306 class_AB_v3_sym_0.VOP.n2 GND 1.51f
C307 class_AB_v3_sym_0.VOP.t6 GND 0.0301f
C308 class_AB_v3_sym_0.VOP.t0 GND 0.133f
C309 class_AB_v3_sym_0.VOP.t7 GND 0.208f
C310 class_AB_v3_sym_0.VOP.n3 GND 1.3f
C311 class_AB_v3_sym_0.VOP.n4 GND 0.849f
C312 class_AB_v3_sym_0.VOP.n5 GND 1.9f
C313 class_AB_v3_sym_0.VOP.n6 GND 1.63f
C314 class_AB_v3_sym_0.VON.n0 GND 0.111f
C315 class_AB_v3_sym_0.VON.n1 GND 2.06f
C316 class_AB_v3_sym_0.VON.t5 GND 0.013f
C317 class_AB_v3_sym_0.VON.t6 GND 0.0209f
C318 class_AB_v3_sym_0.VON.n2 GND 0.0431f
C319 class_AB_v3_sym_0.VON.t2 GND 0.14f
C320 class_AB_v3_sym_0.VON.t4 GND 0.0237f
C321 class_AB_v3_sym_0.VON.t3 GND 0.16f
C322 class_AB_v3_sym_0.VON.t7 GND 0.162f
C323 class_AB_v3_sym_0.VON.n3 GND 0.927f
C324 class_AB_v3_sym_0.VON.n4 GND 0.884f
C325 class_AB_v3_sym_0.VON.t0 GND 0.0145f
C326 class_AB_v3_sym_0.VON.t1 GND 0.31f
C327 class_AB_v3_sym_0.VON.n5 GND 1.16f
C328 CLK.t0 GND 0.108f
C329 CLK.t2 GND 0.624f
C330 CLK.t3 GND 0.631f
C331 CLK.t1 GND 0.114f
C332 CLK.n0 GND 0.889f
C333 CLK.n1 GND 0.0125f
C334 CLK.t5 GND 0.0163f
C335 CLK.n2 GND 0.549f
C336 CLK.n3 GND 0.0134f
C337 CLK.n4 GND 0.13f
C338 CLK.t4 GND 0.181f
C339 CLK.n5 GND 0.757f
C340 CLK.n6 GND 0.691f
C341 CLK.n7 GND 0.261f
.ends

