magic
tech sky130A
magscale 1 2
timestamp 1713499047
<< nwell >>
rect 12570 -540 13530 350
rect 8560 -1270 16750 -540
rect 8610 -2410 8980 -1850
rect 10660 -5770 19310 -5210
rect 10664 -9908 19314 -9348
rect 10660 -13560 19310 -13000
<< pwell >>
rect 8600 -1810 16750 -1310
rect 10870 -2160 11510 -1810
rect 15670 -1850 16710 -1810
rect 15390 -2090 16710 -1850
rect 15390 -2760 16350 -2090
rect 16560 -2140 16710 -2090
rect 10660 -6280 19310 -5810
rect 10664 -10418 19314 -9948
rect 10660 -14070 19310 -13600
<< psubdiff >>
rect 10360 -1640 10530 -1610
rect 9460 -1670 9630 -1640
rect 9460 -1780 9490 -1670
rect 9600 -1780 9630 -1670
rect 10360 -1750 10390 -1640
rect 10500 -1750 10530 -1640
rect 10360 -1780 10530 -1750
rect 11620 -1650 11790 -1620
rect 11620 -1760 11650 -1650
rect 11760 -1760 11790 -1650
rect 9460 -1810 9630 -1780
rect 11620 -1790 11790 -1760
rect 13030 -1640 13200 -1610
rect 13030 -1750 13060 -1640
rect 13170 -1750 13200 -1640
rect 13030 -1780 13200 -1750
rect 14190 -1650 14360 -1620
rect 14190 -1760 14220 -1650
rect 14330 -1760 14360 -1650
rect 14190 -1790 14360 -1760
rect 15260 -1640 15430 -1610
rect 15260 -1750 15290 -1640
rect 15400 -1750 15430 -1640
rect 15260 -1780 15430 -1750
rect 16370 -1630 16540 -1600
rect 16370 -1740 16400 -1630
rect 16510 -1740 16540 -1630
rect 16370 -1770 16540 -1740
rect 11350 -6110 11520 -6080
rect 11350 -6220 11380 -6110
rect 11490 -6220 11520 -6110
rect 11350 -6250 11520 -6220
rect 12990 -6120 13160 -6090
rect 12990 -6230 13020 -6120
rect 13130 -6230 13160 -6120
rect 12990 -6260 13160 -6230
rect 14400 -6110 14570 -6080
rect 14400 -6220 14430 -6110
rect 14540 -6220 14570 -6110
rect 14400 -6250 14570 -6220
rect 15780 -6110 15950 -6080
rect 15780 -6220 15810 -6110
rect 15920 -6220 15950 -6110
rect 15780 -6250 15950 -6220
rect 17320 -6120 17490 -6090
rect 17320 -6230 17350 -6120
rect 17460 -6230 17490 -6120
rect 17320 -6260 17490 -6230
rect 18600 -6120 18770 -6090
rect 18600 -6230 18630 -6120
rect 18740 -6230 18770 -6120
rect 18600 -6260 18770 -6230
rect 11354 -10248 11524 -10218
rect 11354 -10358 11384 -10248
rect 11494 -10358 11524 -10248
rect 11354 -10388 11524 -10358
rect 12994 -10258 13164 -10228
rect 12994 -10368 13024 -10258
rect 13134 -10368 13164 -10258
rect 12994 -10398 13164 -10368
rect 14404 -10248 14574 -10218
rect 14404 -10358 14434 -10248
rect 14544 -10358 14574 -10248
rect 14404 -10388 14574 -10358
rect 15784 -10248 15954 -10218
rect 15784 -10358 15814 -10248
rect 15924 -10358 15954 -10248
rect 15784 -10388 15954 -10358
rect 17324 -10258 17494 -10228
rect 17324 -10368 17354 -10258
rect 17464 -10368 17494 -10258
rect 17324 -10398 17494 -10368
rect 18604 -10258 18774 -10228
rect 18604 -10368 18634 -10258
rect 18744 -10368 18774 -10258
rect 18604 -10398 18774 -10368
rect 11350 -13900 11520 -13870
rect 11350 -14010 11380 -13900
rect 11490 -14010 11520 -13900
rect 11350 -14040 11520 -14010
rect 12990 -13910 13160 -13880
rect 12990 -14020 13020 -13910
rect 13130 -14020 13160 -13910
rect 12990 -14050 13160 -14020
rect 14400 -13900 14570 -13870
rect 14400 -14010 14430 -13900
rect 14540 -14010 14570 -13900
rect 14400 -14040 14570 -14010
rect 15780 -13900 15950 -13870
rect 15780 -14010 15810 -13900
rect 15920 -14010 15950 -13900
rect 15780 -14040 15950 -14010
rect 17320 -13910 17490 -13880
rect 17320 -14020 17350 -13910
rect 17460 -14020 17490 -13910
rect 17320 -14050 17490 -14020
rect 18600 -13910 18770 -13880
rect 18600 -14020 18630 -13910
rect 18740 -14020 18770 -13910
rect 18600 -14050 18770 -14020
<< nsubdiff >>
rect 8760 -690 8940 -660
rect 8760 -800 8790 -690
rect 8900 -800 8940 -690
rect 8760 -830 8940 -800
rect 9370 -690 9550 -660
rect 9370 -800 9410 -690
rect 9520 -800 9550 -690
rect 9370 -830 9550 -800
rect 9980 -700 10160 -670
rect 9980 -810 10010 -700
rect 10120 -810 10160 -700
rect 9980 -840 10160 -810
rect 10630 -710 10810 -680
rect 10630 -820 10660 -710
rect 10770 -820 10810 -710
rect 10630 -850 10810 -820
rect 11340 -700 11520 -670
rect 11340 -810 11380 -700
rect 11490 -810 11520 -700
rect 11340 -840 11520 -810
rect 12060 -700 12240 -670
rect 12060 -810 12090 -700
rect 12200 -810 12240 -700
rect 12060 -840 12240 -810
rect 13710 -720 13890 -690
rect 13710 -830 13750 -720
rect 13860 -830 13890 -720
rect 13710 -860 13890 -830
rect 15150 -730 15330 -700
rect 15150 -840 15190 -730
rect 15300 -840 15330 -730
rect 15150 -870 15330 -840
rect 8720 -2230 8890 -2200
rect 8720 -2340 8750 -2230
rect 8860 -2340 8890 -2230
rect 8720 -2370 8890 -2340
rect 11320 -5280 11490 -5250
rect 11320 -5390 11350 -5280
rect 11460 -5390 11490 -5280
rect 11320 -5420 11490 -5390
rect 13020 -5280 13190 -5250
rect 13020 -5390 13050 -5280
rect 13160 -5390 13190 -5280
rect 13020 -5420 13190 -5390
rect 14400 -5280 14570 -5250
rect 14400 -5390 14430 -5280
rect 14540 -5390 14570 -5280
rect 14400 -5420 14570 -5390
rect 15690 -5280 15860 -5250
rect 15690 -5390 15720 -5280
rect 15830 -5390 15860 -5280
rect 15690 -5420 15860 -5390
rect 17210 -5280 17380 -5250
rect 17210 -5390 17240 -5280
rect 17350 -5390 17380 -5280
rect 17210 -5420 17380 -5390
rect 18620 -5280 18790 -5250
rect 18620 -5390 18650 -5280
rect 18760 -5390 18790 -5280
rect 18620 -5420 18790 -5390
rect 11324 -9418 11494 -9388
rect 11324 -9528 11354 -9418
rect 11464 -9528 11494 -9418
rect 11324 -9558 11494 -9528
rect 13024 -9418 13194 -9388
rect 13024 -9528 13054 -9418
rect 13164 -9528 13194 -9418
rect 13024 -9558 13194 -9528
rect 14404 -9418 14574 -9388
rect 14404 -9528 14434 -9418
rect 14544 -9528 14574 -9418
rect 14404 -9558 14574 -9528
rect 15694 -9418 15864 -9388
rect 15694 -9528 15724 -9418
rect 15834 -9528 15864 -9418
rect 15694 -9558 15864 -9528
rect 17214 -9418 17384 -9388
rect 17214 -9528 17244 -9418
rect 17354 -9528 17384 -9418
rect 17214 -9558 17384 -9528
rect 18624 -9418 18794 -9388
rect 18624 -9528 18654 -9418
rect 18764 -9528 18794 -9418
rect 18624 -9558 18794 -9528
rect 11320 -13070 11490 -13040
rect 11320 -13180 11350 -13070
rect 11460 -13180 11490 -13070
rect 11320 -13210 11490 -13180
rect 13020 -13070 13190 -13040
rect 13020 -13180 13050 -13070
rect 13160 -13180 13190 -13070
rect 13020 -13210 13190 -13180
rect 14400 -13070 14570 -13040
rect 14400 -13180 14430 -13070
rect 14540 -13180 14570 -13070
rect 14400 -13210 14570 -13180
rect 15690 -13070 15860 -13040
rect 15690 -13180 15720 -13070
rect 15830 -13180 15860 -13070
rect 15690 -13210 15860 -13180
rect 17210 -13070 17380 -13040
rect 17210 -13180 17240 -13070
rect 17350 -13180 17380 -13070
rect 17210 -13210 17380 -13180
rect 18620 -13070 18790 -13040
rect 18620 -13180 18650 -13070
rect 18760 -13180 18790 -13070
rect 18620 -13210 18790 -13180
<< psubdiffcont >>
rect 9490 -1780 9600 -1670
rect 10390 -1750 10500 -1640
rect 11650 -1760 11760 -1650
rect 13060 -1750 13170 -1640
rect 14220 -1760 14330 -1650
rect 15290 -1750 15400 -1640
rect 16400 -1740 16510 -1630
rect 11380 -6220 11490 -6110
rect 13020 -6230 13130 -6120
rect 14430 -6220 14540 -6110
rect 15810 -6220 15920 -6110
rect 17350 -6230 17460 -6120
rect 18630 -6230 18740 -6120
rect 11384 -10358 11494 -10248
rect 13024 -10368 13134 -10258
rect 14434 -10358 14544 -10248
rect 15814 -10358 15924 -10248
rect 17354 -10368 17464 -10258
rect 18634 -10368 18744 -10258
rect 11380 -14010 11490 -13900
rect 13020 -14020 13130 -13910
rect 14430 -14010 14540 -13900
rect 15810 -14010 15920 -13900
rect 17350 -14020 17460 -13910
rect 18630 -14020 18740 -13910
<< nsubdiffcont >>
rect 8790 -800 8900 -690
rect 9410 -800 9520 -690
rect 10010 -810 10120 -700
rect 10660 -820 10770 -710
rect 11380 -810 11490 -700
rect 12090 -810 12200 -700
rect 13750 -830 13860 -720
rect 15190 -840 15300 -730
rect 8750 -2340 8860 -2230
rect 11350 -5390 11460 -5280
rect 13050 -5390 13160 -5280
rect 14430 -5390 14540 -5280
rect 15720 -5390 15830 -5280
rect 17240 -5390 17350 -5280
rect 18650 -5390 18760 -5280
rect 11354 -9528 11464 -9418
rect 13054 -9528 13164 -9418
rect 14434 -9528 14544 -9418
rect 15724 -9528 15834 -9418
rect 17244 -9528 17354 -9418
rect 18654 -9528 18764 -9418
rect 11350 -13180 11460 -13070
rect 13050 -13180 13160 -13070
rect 14430 -13180 14540 -13070
rect 15720 -13180 15830 -13070
rect 17240 -13180 17350 -13070
rect 18650 -13180 18760 -13070
<< locali >>
rect 10650 -1110 10690 -1100
rect 10640 -1150 10650 -1140
rect 10690 -1150 10700 -1140
rect 10640 -1190 10700 -1150
rect 8330 -1220 8620 -1200
rect 8330 -1380 8350 -1220
rect 8510 -1260 8620 -1220
rect 8780 -1260 8820 -1250
rect 9270 -1260 9320 -1250
rect 8510 -1270 8680 -1260
rect 8510 -1300 8730 -1270
rect 8510 -1380 8620 -1300
rect 8780 -1310 8980 -1260
rect 9270 -1310 9430 -1260
rect 8330 -1400 8620 -1380
rect 8330 -1670 8600 -1650
rect 8330 -1830 8350 -1670
rect 8510 -1820 8600 -1670
rect 8510 -1830 8780 -1820
rect 8330 -1860 8780 -1830
rect 11090 -5760 11190 -5740
rect 11090 -5800 11290 -5760
rect 11090 -5820 11190 -5800
rect 11340 -5810 11510 -5760
rect 11830 -5810 11970 -5760
rect 11090 -9900 11190 -9870
rect 11090 -9940 11290 -9900
rect 11340 -9910 11530 -9900
rect 11340 -9940 11570 -9910
rect 11090 -9980 11190 -9940
rect 11340 -9950 11530 -9940
rect 11830 -9950 11990 -9900
rect 11090 -13550 11190 -13500
rect 11090 -13590 11290 -13550
rect 11090 -13630 11190 -13590
rect 11340 -13600 11530 -13550
rect 11830 -13600 11980 -13550
<< viali >>
rect 8760 -690 8940 -660
rect 8760 -800 8790 -690
rect 8790 -800 8900 -690
rect 8900 -800 8940 -690
rect 8760 -830 8940 -800
rect 9370 -690 9550 -660
rect 9370 -800 9410 -690
rect 9410 -800 9520 -690
rect 9520 -800 9550 -690
rect 9370 -830 9550 -800
rect 9980 -700 10160 -670
rect 9980 -810 10010 -700
rect 10010 -810 10120 -700
rect 10120 -810 10160 -700
rect 9980 -840 10160 -810
rect 10630 -710 10810 -680
rect 10630 -820 10660 -710
rect 10660 -820 10770 -710
rect 10770 -820 10810 -710
rect 10630 -850 10810 -820
rect 11340 -700 11520 -670
rect 11340 -810 11380 -700
rect 11380 -810 11490 -700
rect 11490 -810 11520 -700
rect 11340 -840 11520 -810
rect 12060 -700 12240 -670
rect 12060 -810 12090 -700
rect 12090 -810 12200 -700
rect 12200 -810 12240 -700
rect 12060 -840 12240 -810
rect 13710 -720 13890 -690
rect 13710 -830 13750 -720
rect 13750 -830 13860 -720
rect 13860 -830 13890 -720
rect 13710 -860 13890 -830
rect 15150 -730 15330 -700
rect 15150 -840 15190 -730
rect 15190 -840 15300 -730
rect 15300 -840 15330 -730
rect 15150 -870 15330 -840
rect 10650 -1150 10690 -1110
rect 8350 -1380 8510 -1220
rect 10650 -1230 10690 -1190
rect 10650 -1310 10690 -1270
rect 11238 -1304 11643 -1264
rect 10650 -1400 10690 -1360
rect 12120 -1400 12160 -1130
rect 12740 -1307 13110 -1267
rect 13600 -1410 13640 -1140
rect 14199 -1304 14569 -1264
rect 15070 -1380 15110 -1110
rect 15339 -1305 15619 -1265
rect 16540 -1400 16580 -1130
rect 10360 -1640 10530 -1610
rect 8350 -1830 8510 -1670
rect 9460 -1670 9630 -1640
rect 9460 -1780 9490 -1670
rect 9490 -1780 9600 -1670
rect 9600 -1780 9630 -1670
rect 10360 -1750 10390 -1640
rect 10390 -1750 10500 -1640
rect 10500 -1750 10530 -1640
rect 10360 -1780 10530 -1750
rect 11620 -1650 11790 -1620
rect 11620 -1760 11650 -1650
rect 11650 -1760 11760 -1650
rect 11760 -1760 11790 -1650
rect 9460 -1810 9630 -1780
rect 11620 -1790 11790 -1760
rect 13030 -1640 13200 -1610
rect 13030 -1750 13060 -1640
rect 13060 -1750 13170 -1640
rect 13170 -1750 13200 -1640
rect 13030 -1780 13200 -1750
rect 14190 -1650 14360 -1620
rect 14190 -1760 14220 -1650
rect 14220 -1760 14330 -1650
rect 14330 -1760 14360 -1650
rect 14190 -1790 14360 -1760
rect 15260 -1640 15430 -1610
rect 15260 -1750 15290 -1640
rect 15290 -1750 15400 -1640
rect 15400 -1750 15430 -1640
rect 15260 -1780 15430 -1750
rect 16370 -1630 16540 -1600
rect 16370 -1740 16400 -1630
rect 16400 -1740 16510 -1630
rect 16510 -1740 16540 -1630
rect 16370 -1770 16540 -1740
rect 8810 -2030 8860 -1920
rect 8720 -2230 8890 -2200
rect 8720 -2340 8750 -2230
rect 8750 -2340 8860 -2230
rect 8860 -2340 8890 -2230
rect 8720 -2370 8890 -2340
rect 11320 -5280 11490 -5250
rect 11320 -5390 11350 -5280
rect 11350 -5390 11460 -5280
rect 11460 -5390 11490 -5280
rect 11320 -5420 11490 -5390
rect 13020 -5280 13190 -5250
rect 13020 -5390 13050 -5280
rect 13050 -5390 13160 -5280
rect 13160 -5390 13190 -5280
rect 13020 -5420 13190 -5390
rect 14400 -5280 14570 -5250
rect 14400 -5390 14430 -5280
rect 14430 -5390 14540 -5280
rect 14540 -5390 14570 -5280
rect 14400 -5420 14570 -5390
rect 15690 -5280 15860 -5250
rect 15690 -5390 15720 -5280
rect 15720 -5390 15830 -5280
rect 15830 -5390 15860 -5280
rect 15690 -5420 15860 -5390
rect 17210 -5280 17380 -5250
rect 17210 -5390 17240 -5280
rect 17240 -5390 17350 -5280
rect 17350 -5390 17380 -5280
rect 17210 -5420 17380 -5390
rect 18620 -5280 18790 -5250
rect 18620 -5390 18650 -5280
rect 18650 -5390 18760 -5280
rect 18760 -5390 18790 -5280
rect 18620 -5420 18790 -5390
rect 10750 -5860 10800 -5770
rect 10920 -5860 10960 -5780
rect 13200 -5860 13250 -5690
rect 13480 -5801 14341 -5767
rect 14680 -5860 14730 -5670
rect 14914 -5800 15775 -5766
rect 16150 -5860 16200 -5680
rect 16393 -5800 17254 -5766
rect 17620 -5870 17670 -5680
rect 17850 -5769 18617 -5767
rect 17848 -5803 18618 -5769
rect 19090 -5870 19140 -5680
rect 11350 -6110 11520 -6080
rect 11350 -6220 11380 -6110
rect 11380 -6220 11490 -6110
rect 11490 -6220 11520 -6110
rect 11350 -6250 11520 -6220
rect 12990 -6120 13160 -6090
rect 12990 -6230 13020 -6120
rect 13020 -6230 13130 -6120
rect 13130 -6230 13160 -6120
rect 12990 -6260 13160 -6230
rect 14400 -6110 14570 -6080
rect 14400 -6220 14430 -6110
rect 14430 -6220 14540 -6110
rect 14540 -6220 14570 -6110
rect 14400 -6250 14570 -6220
rect 15780 -6110 15950 -6080
rect 15780 -6220 15810 -6110
rect 15810 -6220 15920 -6110
rect 15920 -6220 15950 -6110
rect 15780 -6250 15950 -6220
rect 17320 -6120 17490 -6090
rect 17320 -6230 17350 -6120
rect 17350 -6230 17460 -6120
rect 17460 -6230 17490 -6120
rect 17320 -6260 17490 -6230
rect 18600 -6120 18770 -6090
rect 18600 -6230 18630 -6120
rect 18630 -6230 18740 -6120
rect 18740 -6230 18770 -6120
rect 18600 -6260 18770 -6230
rect 11324 -9418 11494 -9388
rect 11324 -9528 11354 -9418
rect 11354 -9528 11464 -9418
rect 11464 -9528 11494 -9418
rect 11324 -9558 11494 -9528
rect 13024 -9418 13194 -9388
rect 13024 -9528 13054 -9418
rect 13054 -9528 13164 -9418
rect 13164 -9528 13194 -9418
rect 13024 -9558 13194 -9528
rect 14404 -9418 14574 -9388
rect 14404 -9528 14434 -9418
rect 14434 -9528 14544 -9418
rect 14544 -9528 14574 -9418
rect 14404 -9558 14574 -9528
rect 15694 -9418 15864 -9388
rect 15694 -9528 15724 -9418
rect 15724 -9528 15834 -9418
rect 15834 -9528 15864 -9418
rect 15694 -9558 15864 -9528
rect 17214 -9418 17384 -9388
rect 17214 -9528 17244 -9418
rect 17244 -9528 17354 -9418
rect 17354 -9528 17384 -9418
rect 17214 -9558 17384 -9528
rect 18624 -9418 18794 -9388
rect 18624 -9528 18654 -9418
rect 18654 -9528 18764 -9418
rect 18764 -9528 18794 -9418
rect 18624 -9558 18794 -9528
rect 10740 -10000 10800 -9910
rect 10920 -10000 10960 -9910
rect 13204 -9998 13254 -9828
rect 13484 -9939 14345 -9905
rect 14684 -9998 14734 -9808
rect 14918 -9938 15779 -9904
rect 16154 -9998 16204 -9818
rect 16397 -9938 17258 -9904
rect 17624 -10008 17674 -9818
rect 17854 -9907 18621 -9905
rect 17852 -9941 18622 -9907
rect 19094 -10008 19144 -9818
rect 11354 -10248 11524 -10218
rect 11354 -10358 11384 -10248
rect 11384 -10358 11494 -10248
rect 11494 -10358 11524 -10248
rect 11354 -10388 11524 -10358
rect 12994 -10258 13164 -10228
rect 12994 -10368 13024 -10258
rect 13024 -10368 13134 -10258
rect 13134 -10368 13164 -10258
rect 12994 -10398 13164 -10368
rect 14404 -10248 14574 -10218
rect 14404 -10358 14434 -10248
rect 14434 -10358 14544 -10248
rect 14544 -10358 14574 -10248
rect 14404 -10388 14574 -10358
rect 15784 -10248 15954 -10218
rect 15784 -10358 15814 -10248
rect 15814 -10358 15924 -10248
rect 15924 -10358 15954 -10248
rect 15784 -10388 15954 -10358
rect 17324 -10258 17494 -10228
rect 17324 -10368 17354 -10258
rect 17354 -10368 17464 -10258
rect 17464 -10368 17494 -10258
rect 17324 -10398 17494 -10368
rect 18604 -10258 18774 -10228
rect 18604 -10368 18634 -10258
rect 18634 -10368 18744 -10258
rect 18744 -10368 18774 -10258
rect 18604 -10398 18774 -10368
rect 11320 -13070 11490 -13040
rect 11320 -13180 11350 -13070
rect 11350 -13180 11460 -13070
rect 11460 -13180 11490 -13070
rect 11320 -13210 11490 -13180
rect 13020 -13070 13190 -13040
rect 13020 -13180 13050 -13070
rect 13050 -13180 13160 -13070
rect 13160 -13180 13190 -13070
rect 13020 -13210 13190 -13180
rect 14400 -13070 14570 -13040
rect 14400 -13180 14430 -13070
rect 14430 -13180 14540 -13070
rect 14540 -13180 14570 -13070
rect 14400 -13210 14570 -13180
rect 15690 -13070 15860 -13040
rect 15690 -13180 15720 -13070
rect 15720 -13180 15830 -13070
rect 15830 -13180 15860 -13070
rect 15690 -13210 15860 -13180
rect 17210 -13070 17380 -13040
rect 17210 -13180 17240 -13070
rect 17240 -13180 17350 -13070
rect 17350 -13180 17380 -13070
rect 17210 -13210 17380 -13180
rect 18620 -13070 18790 -13040
rect 18620 -13180 18650 -13070
rect 18650 -13180 18760 -13070
rect 18760 -13180 18790 -13070
rect 18620 -13210 18790 -13180
rect 10740 -13650 10800 -13560
rect 10910 -13650 10960 -13560
rect 13200 -13650 13250 -13480
rect 13480 -13591 14341 -13557
rect 14680 -13650 14730 -13460
rect 14914 -13590 15775 -13556
rect 16150 -13650 16200 -13470
rect 16393 -13590 17254 -13556
rect 17620 -13660 17670 -13470
rect 17850 -13559 18617 -13557
rect 17848 -13593 18618 -13559
rect 19090 -13660 19140 -13470
rect 11350 -13900 11520 -13870
rect 11350 -14010 11380 -13900
rect 11380 -14010 11490 -13900
rect 11490 -14010 11520 -13900
rect 11350 -14040 11520 -14010
rect 12990 -13910 13160 -13880
rect 12990 -14020 13020 -13910
rect 13020 -14020 13130 -13910
rect 13130 -14020 13160 -13910
rect 12990 -14050 13160 -14020
rect 14400 -13900 14570 -13870
rect 14400 -14010 14430 -13900
rect 14430 -14010 14540 -13900
rect 14540 -14010 14570 -13900
rect 14400 -14040 14570 -14010
rect 15780 -13900 15950 -13870
rect 15780 -14010 15810 -13900
rect 15810 -14010 15920 -13900
rect 15920 -14010 15950 -13900
rect 15780 -14040 15950 -14010
rect 17320 -13910 17490 -13880
rect 17320 -14020 17350 -13910
rect 17350 -14020 17460 -13910
rect 17460 -14020 17490 -13910
rect 17320 -14050 17490 -14020
rect 18600 -13910 18770 -13880
rect 18600 -14020 18630 -13910
rect 18630 -14020 18740 -13910
rect 18740 -14020 18770 -13910
rect 18600 -14050 18770 -14020
<< metal1 >>
rect 12570 80 13530 350
rect 12570 -350 12830 80
rect 13270 -350 13530 80
rect 12570 -560 13530 -350
rect 15750 -260 16710 -10
rect 15750 -560 16020 -260
rect 480 -610 920 -600
rect 480 -790 690 -610
rect 910 -790 920 -610
rect 480 -800 920 -790
rect 8600 -660 16020 -560
rect 8600 -830 8760 -660
rect 8940 -830 9370 -660
rect 9550 -670 16020 -660
rect 9550 -830 9980 -670
rect 8600 -840 9980 -830
rect 10160 -680 11340 -670
rect 10160 -840 10630 -680
rect 8600 -850 10630 -840
rect 10810 -840 11340 -680
rect 11520 -840 12060 -670
rect 12240 -690 16020 -670
rect 16460 -690 16710 -260
rect 12240 -840 13710 -690
rect 10810 -850 13710 -840
rect 8600 -860 13710 -850
rect 13890 -700 16710 -690
rect 13890 -860 15150 -700
rect 8600 -870 15150 -860
rect 15330 -870 16710 -700
rect 480 -940 920 -930
rect 480 -1120 690 -940
rect 910 -1120 920 -940
rect 8600 -1030 16710 -870
rect 480 -1130 920 -1120
rect 10630 -1110 10780 -1100
rect 15040 -1110 15140 -1100
rect 10630 -1400 10650 -1110
rect 10690 -1140 10780 -1110
rect 10760 -1390 10780 -1140
rect 12090 -1120 12190 -1110
rect 11220 -1250 11660 -1240
rect 11220 -1264 11240 -1250
rect 11640 -1264 11660 -1250
rect 11220 -1304 11238 -1264
rect 11643 -1304 11660 -1264
rect 11220 -1320 11240 -1304
rect 11640 -1320 11660 -1304
rect 11220 -1330 11660 -1320
rect 10690 -1400 10780 -1390
rect 480 -1430 920 -1420
rect 10630 -1430 10780 -1400
rect 12090 -1410 12100 -1120
rect 12180 -1410 12190 -1120
rect 13570 -1130 13670 -1110
rect 12720 -1250 13130 -1240
rect 12720 -1320 12740 -1250
rect 13110 -1320 13130 -1250
rect 12720 -1330 13130 -1320
rect 12090 -1420 12190 -1410
rect 13570 -1420 13580 -1130
rect 13660 -1420 13670 -1130
rect 14180 -1250 14590 -1240
rect 14180 -1320 14190 -1250
rect 14580 -1320 14590 -1250
rect 14180 -1330 14590 -1320
rect 15040 -1380 15050 -1110
rect 15130 -1380 15140 -1110
rect 16510 -1120 16610 -1110
rect 15310 -1250 15640 -1240
rect 15310 -1320 15320 -1250
rect 15630 -1320 15640 -1250
rect 15310 -1330 15640 -1320
rect 15040 -1390 15140 -1380
rect 16510 -1410 16520 -1120
rect 16600 -1410 16610 -1120
rect 13570 -1430 13670 -1420
rect 480 -1610 690 -1430
rect 910 -1610 920 -1430
rect 19620 -1450 20030 -1420
rect 480 -1620 920 -1610
rect 8600 -1600 16710 -1470
rect 8600 -1610 16370 -1600
rect 8600 -1640 10360 -1610
rect 8600 -1650 9460 -1640
rect 480 -1710 920 -1700
rect 480 -1890 690 -1710
rect 910 -1890 920 -1710
rect 9350 -1810 9460 -1650
rect 9630 -1780 10360 -1640
rect 10530 -1620 13030 -1610
rect 10530 -1700 11620 -1620
rect 10530 -1780 11020 -1700
rect 9630 -1810 11020 -1780
rect 9350 -1850 11020 -1810
rect 480 -1900 920 -1890
rect 8380 -1920 8870 -1900
rect 8380 -1990 8810 -1920
rect 7640 -2000 8810 -1990
rect 480 -2170 920 -2160
rect 480 -2350 690 -2170
rect 910 -2350 920 -2170
rect 7640 -2240 7650 -2000
rect 7780 -2030 8810 -2000
rect 8860 -2030 8870 -1920
rect 7780 -2050 8870 -2030
rect 10870 -2050 11020 -1850
rect 11380 -1790 11620 -1700
rect 11790 -1780 13030 -1620
rect 13200 -1620 15260 -1610
rect 13200 -1780 14190 -1620
rect 11790 -1790 14190 -1780
rect 14360 -1780 15260 -1620
rect 15430 -1770 16370 -1610
rect 16540 -1770 16710 -1600
rect 15430 -1780 16710 -1770
rect 14360 -1790 16710 -1780
rect 11380 -1850 16710 -1790
rect 11380 -2050 11510 -1850
rect 7780 -2240 8560 -2050
rect 7640 -2250 8560 -2240
rect 8600 -2120 9470 -2090
rect 8600 -2200 9010 -2120
rect 480 -2360 920 -2350
rect 8600 -2370 8720 -2200
rect 8890 -2370 9010 -2200
rect 8600 -2380 9010 -2370
rect 9440 -2380 9470 -2120
rect 10870 -2160 11510 -2050
rect 15390 -2110 16710 -1850
rect 19620 -1830 19650 -1450
rect 20000 -1530 20030 -1450
rect 20000 -1730 20230 -1530
rect 20000 -1830 20030 -1730
rect 19620 -1860 20030 -1830
rect 8600 -2410 9470 -2380
rect 15390 -2460 15700 -2110
rect 16060 -2140 16710 -2110
rect 16060 -2460 16350 -2140
rect 480 -2530 920 -2520
rect 480 -2710 690 -2530
rect 910 -2710 920 -2530
rect 480 -2720 920 -2710
rect 15390 -2760 16350 -2460
rect 480 -2930 920 -2920
rect 480 -3110 690 -2930
rect 910 -3110 920 -2930
rect 480 -3120 920 -3110
rect 480 -3380 920 -3370
rect 480 -3560 690 -3380
rect 910 -3560 920 -3380
rect 480 -3570 920 -3560
rect 480 -3750 920 -3740
rect 480 -3930 690 -3750
rect 910 -3930 920 -3750
rect 480 -3940 920 -3930
rect 10660 -4610 19310 -4580
rect 10660 -5180 10690 -4610
rect 19280 -5180 19310 -4610
rect 10660 -5250 19310 -5180
rect 10660 -5420 11320 -5250
rect 11490 -5420 13020 -5250
rect 13190 -5420 14400 -5250
rect 14570 -5420 15690 -5250
rect 15860 -5420 17210 -5250
rect 17380 -5420 18620 -5250
rect 18790 -5420 19310 -5250
rect 10660 -5530 19310 -5420
rect 14660 -5660 14750 -5650
rect 13180 -5680 13270 -5670
rect 10330 -5760 10820 -5750
rect 10330 -5870 10340 -5760
rect 10420 -5770 10820 -5760
rect 10420 -5860 10750 -5770
rect 10800 -5860 10820 -5770
rect 10420 -5870 10820 -5860
rect 10330 -5880 10820 -5870
rect 10900 -5760 10980 -5750
rect 10900 -5870 10910 -5760
rect 10970 -5870 10980 -5760
rect 10900 -5880 10980 -5870
rect 13180 -5870 13190 -5680
rect 13260 -5870 13270 -5680
rect 13450 -5740 14360 -5730
rect 13450 -5820 13460 -5740
rect 14350 -5820 14360 -5740
rect 13450 -5830 14360 -5820
rect 13180 -5880 13270 -5870
rect 14660 -5870 14670 -5660
rect 14740 -5870 14750 -5660
rect 16130 -5670 16220 -5660
rect 14900 -5740 15800 -5730
rect 14900 -5820 14910 -5740
rect 15790 -5820 15800 -5740
rect 14900 -5830 15800 -5820
rect 14660 -5880 14750 -5870
rect 16130 -5870 16140 -5670
rect 16210 -5870 16220 -5670
rect 17600 -5670 17690 -5660
rect 16370 -5750 17270 -5740
rect 16370 -5820 16380 -5750
rect 17260 -5820 17270 -5750
rect 16370 -5830 17270 -5820
rect 16130 -5880 16220 -5870
rect 17600 -5880 17610 -5670
rect 17680 -5880 17690 -5670
rect 19070 -5670 19160 -5660
rect 17840 -5749 18640 -5740
rect 17840 -5767 17852 -5749
rect 17840 -5769 17850 -5767
rect 17840 -5803 17848 -5769
rect 17840 -5821 17852 -5803
rect 18632 -5821 18640 -5749
rect 17840 -5830 18640 -5821
rect 17600 -5890 17690 -5880
rect 19070 -5880 19080 -5670
rect 19150 -5880 19160 -5670
rect 19070 -5890 19160 -5880
rect 19620 -5950 20030 -5920
rect 10660 -6080 19310 -5970
rect 10660 -6250 11350 -6080
rect 11520 -6090 14400 -6080
rect 11520 -6250 12990 -6090
rect 10660 -6260 12990 -6250
rect 13160 -6250 14400 -6090
rect 14570 -6250 15780 -6080
rect 15950 -6090 19310 -6080
rect 15950 -6250 17320 -6090
rect 13160 -6260 17320 -6250
rect 17490 -6260 18600 -6090
rect 18770 -6260 19310 -6090
rect 10660 -6310 19310 -6260
rect 10660 -6880 10690 -6310
rect 19280 -6880 19310 -6310
rect 19620 -6330 19650 -5950
rect 20000 -6060 20030 -5950
rect 20000 -6260 20230 -6060
rect 20000 -6330 20030 -6260
rect 19620 -6360 20030 -6330
rect 10660 -6910 19310 -6880
rect 10664 -8748 19314 -8718
rect 680 -8770 920 -8760
rect 680 -8950 690 -8770
rect 910 -8950 920 -8770
rect 680 -8960 920 -8950
rect 470 -9100 920 -9090
rect 470 -9280 690 -9100
rect 910 -9280 920 -9100
rect 470 -9290 920 -9280
rect 10664 -9318 10694 -8748
rect 19284 -9318 19314 -8748
rect 10664 -9388 19314 -9318
rect 10664 -9558 11324 -9388
rect 11494 -9558 13024 -9388
rect 13194 -9558 14404 -9388
rect 14574 -9558 15694 -9388
rect 15864 -9558 17214 -9388
rect 17384 -9558 18624 -9388
rect 18794 -9558 19314 -9388
rect 470 -9590 920 -9580
rect 470 -9770 690 -9590
rect 910 -9770 920 -9590
rect 10664 -9668 19314 -9558
rect 470 -9780 920 -9770
rect 14664 -9798 14754 -9788
rect 13184 -9818 13274 -9808
rect 470 -9870 920 -9860
rect 470 -10050 690 -9870
rect 910 -10050 920 -9870
rect 9810 -9890 10820 -9880
rect 9810 -10010 9820 -9890
rect 9940 -9910 10820 -9890
rect 9940 -10000 10740 -9910
rect 10800 -10000 10820 -9910
rect 9940 -10010 10820 -10000
rect 9810 -10020 10820 -10010
rect 10900 -9890 10980 -9880
rect 10900 -10010 10910 -9890
rect 10970 -10010 10980 -9890
rect 10900 -10020 10980 -10010
rect 13184 -10008 13194 -9818
rect 13264 -10008 13274 -9818
rect 13454 -9878 14364 -9868
rect 13454 -9958 13464 -9878
rect 14354 -9958 14364 -9878
rect 13454 -9968 14364 -9958
rect 13184 -10018 13274 -10008
rect 14664 -10008 14674 -9798
rect 14744 -10008 14754 -9798
rect 16134 -9808 16224 -9798
rect 14904 -9878 15804 -9868
rect 14904 -9958 14914 -9878
rect 15794 -9958 15804 -9878
rect 14904 -9968 15804 -9958
rect 14664 -10018 14754 -10008
rect 16134 -10008 16144 -9808
rect 16214 -10008 16224 -9808
rect 17604 -9808 17694 -9798
rect 16374 -9888 17274 -9878
rect 16374 -9958 16384 -9888
rect 17264 -9958 17274 -9888
rect 16374 -9968 17274 -9958
rect 16134 -10018 16224 -10008
rect 17604 -10018 17614 -9808
rect 17684 -10018 17694 -9808
rect 19074 -9808 19164 -9798
rect 17844 -9887 18644 -9878
rect 17844 -9905 17856 -9887
rect 17844 -9907 17854 -9905
rect 17844 -9941 17852 -9907
rect 17844 -9959 17856 -9941
rect 18636 -9959 18644 -9887
rect 17844 -9968 18644 -9959
rect 17604 -10028 17694 -10018
rect 19074 -10018 19084 -9808
rect 19154 -10018 19164 -9808
rect 19074 -10028 19164 -10018
rect 470 -10060 920 -10050
rect 10664 -10218 19314 -10108
rect 470 -10330 920 -10320
rect 470 -10510 690 -10330
rect 910 -10510 920 -10330
rect 470 -10520 920 -10510
rect 10664 -10388 11354 -10218
rect 11524 -10228 14404 -10218
rect 11524 -10388 12994 -10228
rect 10664 -10398 12994 -10388
rect 13164 -10388 14404 -10228
rect 14574 -10388 15784 -10218
rect 15954 -10228 19314 -10218
rect 15954 -10388 17324 -10228
rect 13164 -10398 17324 -10388
rect 17494 -10398 18604 -10228
rect 18774 -10398 19314 -10228
rect 10664 -10448 19314 -10398
rect 470 -10690 920 -10680
rect 470 -10870 690 -10690
rect 910 -10870 920 -10690
rect 470 -10880 920 -10870
rect 10664 -11018 10694 -10448
rect 19284 -11018 19314 -10448
rect 19620 -10110 20030 -10080
rect 19620 -10490 19650 -10110
rect 20000 -10210 20030 -10110
rect 20000 -10410 20230 -10210
rect 20000 -10490 20030 -10410
rect 19620 -10520 20030 -10490
rect 10664 -11048 19314 -11018
rect 470 -11090 920 -11080
rect 470 -11270 690 -11090
rect 910 -11270 920 -11090
rect 470 -11280 920 -11270
rect 470 -11540 920 -11530
rect 470 -11720 690 -11540
rect 910 -11720 920 -11540
rect 470 -11730 920 -11720
rect 480 -11910 920 -11900
rect 480 -12090 690 -11910
rect 910 -12090 920 -11910
rect 480 -12100 920 -12090
rect 10660 -12400 19310 -12370
rect 10660 -12970 10690 -12400
rect 19280 -12970 19310 -12400
rect 10660 -13040 19310 -12970
rect 10660 -13210 11320 -13040
rect 11490 -13210 13020 -13040
rect 13190 -13210 14400 -13040
rect 14570 -13210 15690 -13040
rect 15860 -13210 17210 -13040
rect 17380 -13210 18620 -13040
rect 18790 -13210 19310 -13040
rect 10660 -13320 19310 -13210
rect 14660 -13450 14750 -13440
rect 13180 -13470 13270 -13460
rect 10150 -13550 10820 -13540
rect 10150 -13660 10160 -13550
rect 10310 -13560 10820 -13550
rect 10310 -13650 10740 -13560
rect 10800 -13650 10820 -13560
rect 10310 -13660 10820 -13650
rect 10150 -13670 10820 -13660
rect 10890 -13550 10980 -13540
rect 10890 -13660 10900 -13550
rect 10970 -13660 10980 -13550
rect 10890 -13670 10980 -13660
rect 13180 -13660 13190 -13470
rect 13260 -13660 13270 -13470
rect 13450 -13530 14360 -13520
rect 13450 -13610 13460 -13530
rect 14350 -13610 14360 -13530
rect 13450 -13620 14360 -13610
rect 13180 -13670 13270 -13660
rect 14660 -13660 14670 -13450
rect 14740 -13660 14750 -13450
rect 16130 -13460 16220 -13450
rect 14900 -13530 15800 -13520
rect 14900 -13610 14910 -13530
rect 15790 -13610 15800 -13530
rect 14900 -13620 15800 -13610
rect 14660 -13670 14750 -13660
rect 16130 -13660 16140 -13460
rect 16210 -13660 16220 -13460
rect 17600 -13460 17690 -13450
rect 16370 -13540 17270 -13530
rect 16370 -13610 16380 -13540
rect 17260 -13610 17270 -13540
rect 16370 -13620 17270 -13610
rect 16130 -13670 16220 -13660
rect 17600 -13670 17610 -13460
rect 17680 -13670 17690 -13460
rect 19070 -13460 19160 -13450
rect 17840 -13539 18640 -13530
rect 17840 -13557 17852 -13539
rect 17840 -13559 17850 -13557
rect 17840 -13593 17848 -13559
rect 17840 -13611 17852 -13593
rect 18632 -13611 18640 -13539
rect 17840 -13620 18640 -13611
rect 17600 -13680 17690 -13670
rect 19070 -13670 19080 -13460
rect 19150 -13670 19160 -13460
rect 19070 -13680 19160 -13670
rect 19620 -13740 20030 -13710
rect 10660 -13870 19310 -13760
rect 10660 -14040 11350 -13870
rect 11520 -13880 14400 -13870
rect 11520 -14040 12990 -13880
rect 10660 -14050 12990 -14040
rect 13160 -14040 14400 -13880
rect 14570 -14040 15780 -13870
rect 15950 -13880 19310 -13870
rect 15950 -14040 17320 -13880
rect 13160 -14050 17320 -14040
rect 17490 -14050 18600 -13880
rect 18770 -14050 19310 -13880
rect 10660 -14100 19310 -14050
rect 10660 -14670 10690 -14100
rect 19280 -14670 19310 -14100
rect 19620 -14120 19650 -13740
rect 20000 -13820 20030 -13740
rect 20000 -14020 20230 -13820
rect 20000 -14120 20030 -14020
rect 19620 -14150 20030 -14120
rect 10660 -14700 19310 -14670
<< via1 >>
rect 12830 -350 13270 80
rect 690 -790 910 -610
rect 16020 -690 16460 -260
rect 690 -1120 910 -940
rect 10650 -1150 10690 -1140
rect 10690 -1150 10760 -1140
rect 10650 -1190 10760 -1150
rect 10650 -1230 10690 -1190
rect 10690 -1230 10760 -1190
rect 10650 -1270 10760 -1230
rect 10650 -1310 10690 -1270
rect 10690 -1310 10760 -1270
rect 10650 -1360 10760 -1310
rect 10650 -1390 10690 -1360
rect 10690 -1390 10760 -1360
rect 11240 -1264 11640 -1250
rect 11240 -1304 11640 -1264
rect 11240 -1320 11640 -1304
rect 12100 -1130 12180 -1120
rect 12100 -1400 12120 -1130
rect 12120 -1400 12160 -1130
rect 12160 -1400 12180 -1130
rect 12100 -1410 12180 -1400
rect 12740 -1267 13110 -1250
rect 12740 -1307 13110 -1267
rect 12740 -1320 13110 -1307
rect 13580 -1140 13660 -1130
rect 13580 -1410 13600 -1140
rect 13600 -1410 13640 -1140
rect 13640 -1410 13660 -1140
rect 13580 -1420 13660 -1410
rect 14190 -1264 14580 -1250
rect 14190 -1304 14199 -1264
rect 14199 -1304 14569 -1264
rect 14569 -1304 14580 -1264
rect 14190 -1320 14580 -1304
rect 15050 -1380 15070 -1110
rect 15070 -1380 15110 -1110
rect 15110 -1380 15130 -1110
rect 15320 -1265 15630 -1250
rect 15320 -1305 15339 -1265
rect 15339 -1305 15619 -1265
rect 15619 -1305 15630 -1265
rect 15320 -1320 15630 -1305
rect 16520 -1130 16600 -1120
rect 16520 -1400 16540 -1130
rect 16540 -1400 16580 -1130
rect 16580 -1400 16600 -1130
rect 16520 -1410 16600 -1400
rect 690 -1610 910 -1430
rect 690 -1890 910 -1710
rect 690 -2350 910 -2170
rect 7650 -2240 7780 -2000
rect 11020 -2050 11380 -1700
rect 9010 -2380 9440 -2120
rect 19650 -1830 20000 -1450
rect 15700 -2460 16060 -2110
rect 690 -2710 910 -2530
rect 690 -3110 910 -2930
rect 690 -3560 910 -3380
rect 690 -3930 910 -3750
rect 10690 -5180 19280 -4610
rect 10340 -5870 10420 -5760
rect 10910 -5780 10970 -5760
rect 10910 -5860 10920 -5780
rect 10920 -5860 10960 -5780
rect 10960 -5860 10970 -5780
rect 10910 -5870 10970 -5860
rect 13190 -5690 13260 -5680
rect 13190 -5860 13200 -5690
rect 13200 -5860 13250 -5690
rect 13250 -5860 13260 -5690
rect 13190 -5870 13260 -5860
rect 13460 -5767 14350 -5740
rect 13460 -5801 13480 -5767
rect 13480 -5801 14341 -5767
rect 14341 -5801 14350 -5767
rect 13460 -5820 14350 -5801
rect 14670 -5670 14740 -5660
rect 14670 -5860 14680 -5670
rect 14680 -5860 14730 -5670
rect 14730 -5860 14740 -5670
rect 14670 -5870 14740 -5860
rect 14910 -5766 15790 -5740
rect 14910 -5800 14914 -5766
rect 14914 -5800 15775 -5766
rect 15775 -5800 15790 -5766
rect 14910 -5820 15790 -5800
rect 16140 -5680 16210 -5670
rect 16140 -5860 16150 -5680
rect 16150 -5860 16200 -5680
rect 16200 -5860 16210 -5680
rect 16140 -5870 16210 -5860
rect 16380 -5766 17260 -5750
rect 16380 -5800 16393 -5766
rect 16393 -5800 17254 -5766
rect 17254 -5800 17260 -5766
rect 16380 -5820 17260 -5800
rect 17610 -5680 17680 -5670
rect 17610 -5870 17620 -5680
rect 17620 -5870 17670 -5680
rect 17670 -5870 17680 -5680
rect 17610 -5880 17680 -5870
rect 17852 -5767 18632 -5749
rect 17852 -5769 18617 -5767
rect 18617 -5769 18632 -5767
rect 17852 -5803 18618 -5769
rect 18618 -5803 18632 -5769
rect 17852 -5821 18632 -5803
rect 19080 -5680 19150 -5670
rect 19080 -5870 19090 -5680
rect 19090 -5870 19140 -5680
rect 19140 -5870 19150 -5680
rect 19080 -5880 19150 -5870
rect 10690 -6880 19280 -6310
rect 19650 -6330 20000 -5950
rect 690 -8950 910 -8770
rect 690 -9280 910 -9100
rect 10694 -9318 19284 -8748
rect 690 -9770 910 -9590
rect 690 -10050 910 -9870
rect 9820 -10010 9940 -9890
rect 10910 -9910 10970 -9890
rect 10910 -10000 10920 -9910
rect 10920 -10000 10960 -9910
rect 10960 -10000 10970 -9910
rect 10910 -10010 10970 -10000
rect 13194 -9828 13264 -9818
rect 13194 -9998 13204 -9828
rect 13204 -9998 13254 -9828
rect 13254 -9998 13264 -9828
rect 13194 -10008 13264 -9998
rect 13464 -9905 14354 -9878
rect 13464 -9939 13484 -9905
rect 13484 -9939 14345 -9905
rect 14345 -9939 14354 -9905
rect 13464 -9958 14354 -9939
rect 14674 -9808 14744 -9798
rect 14674 -9998 14684 -9808
rect 14684 -9998 14734 -9808
rect 14734 -9998 14744 -9808
rect 14674 -10008 14744 -9998
rect 14914 -9904 15794 -9878
rect 14914 -9938 14918 -9904
rect 14918 -9938 15779 -9904
rect 15779 -9938 15794 -9904
rect 14914 -9958 15794 -9938
rect 16144 -9818 16214 -9808
rect 16144 -9998 16154 -9818
rect 16154 -9998 16204 -9818
rect 16204 -9998 16214 -9818
rect 16144 -10008 16214 -9998
rect 16384 -9904 17264 -9888
rect 16384 -9938 16397 -9904
rect 16397 -9938 17258 -9904
rect 17258 -9938 17264 -9904
rect 16384 -9958 17264 -9938
rect 17614 -9818 17684 -9808
rect 17614 -10008 17624 -9818
rect 17624 -10008 17674 -9818
rect 17674 -10008 17684 -9818
rect 17614 -10018 17684 -10008
rect 17856 -9905 18636 -9887
rect 17856 -9907 18621 -9905
rect 18621 -9907 18636 -9905
rect 17856 -9941 18622 -9907
rect 18622 -9941 18636 -9907
rect 17856 -9959 18636 -9941
rect 19084 -9818 19154 -9808
rect 19084 -10008 19094 -9818
rect 19094 -10008 19144 -9818
rect 19144 -10008 19154 -9818
rect 19084 -10018 19154 -10008
rect 690 -10510 910 -10330
rect 690 -10870 910 -10690
rect 10694 -11018 19284 -10448
rect 19650 -10490 20000 -10110
rect 690 -11270 910 -11090
rect 690 -11720 910 -11540
rect 690 -12090 910 -11910
rect 10690 -12970 19280 -12400
rect 10160 -13660 10310 -13550
rect 10900 -13560 10970 -13550
rect 10900 -13650 10910 -13560
rect 10910 -13650 10960 -13560
rect 10960 -13650 10970 -13560
rect 10900 -13660 10970 -13650
rect 13190 -13480 13260 -13470
rect 13190 -13650 13200 -13480
rect 13200 -13650 13250 -13480
rect 13250 -13650 13260 -13480
rect 13190 -13660 13260 -13650
rect 13460 -13557 14350 -13530
rect 13460 -13591 13480 -13557
rect 13480 -13591 14341 -13557
rect 14341 -13591 14350 -13557
rect 13460 -13610 14350 -13591
rect 14670 -13460 14740 -13450
rect 14670 -13650 14680 -13460
rect 14680 -13650 14730 -13460
rect 14730 -13650 14740 -13460
rect 14670 -13660 14740 -13650
rect 14910 -13556 15790 -13530
rect 14910 -13590 14914 -13556
rect 14914 -13590 15775 -13556
rect 15775 -13590 15790 -13556
rect 14910 -13610 15790 -13590
rect 16140 -13470 16210 -13460
rect 16140 -13650 16150 -13470
rect 16150 -13650 16200 -13470
rect 16200 -13650 16210 -13470
rect 16140 -13660 16210 -13650
rect 16380 -13556 17260 -13540
rect 16380 -13590 16393 -13556
rect 16393 -13590 17254 -13556
rect 17254 -13590 17260 -13556
rect 16380 -13610 17260 -13590
rect 17610 -13470 17680 -13460
rect 17610 -13660 17620 -13470
rect 17620 -13660 17670 -13470
rect 17670 -13660 17680 -13470
rect 17610 -13670 17680 -13660
rect 17852 -13557 18632 -13539
rect 17852 -13559 18617 -13557
rect 18617 -13559 18632 -13557
rect 17852 -13593 18618 -13559
rect 18618 -13593 18632 -13559
rect 17852 -13611 18632 -13593
rect 19080 -13470 19150 -13460
rect 19080 -13660 19090 -13470
rect 19090 -13660 19140 -13470
rect 19140 -13660 19150 -13470
rect 19080 -13670 19150 -13660
rect 10690 -14670 19280 -14100
rect 19650 -14120 20000 -13740
<< metal2 >>
rect 12570 80 13530 350
rect 12570 -350 12830 80
rect 13270 -350 13530 80
rect 12570 -560 13530 -350
rect 15750 -260 16710 -10
rect 680 -610 920 -600
rect 680 -790 690 -610
rect 910 -790 920 -610
rect 15750 -690 16020 -260
rect 16460 -690 16710 -260
rect 680 -800 920 -790
rect 10630 -880 10780 -860
rect 680 -940 920 -930
rect 680 -1120 690 -940
rect 910 -1120 920 -940
rect 10630 -970 10650 -880
rect 10760 -970 10780 -880
rect 680 -1130 920 -1120
rect 10630 -1140 10780 -970
rect 680 -1430 920 -1420
rect 680 -1610 690 -1430
rect 910 -1610 920 -1430
rect 680 -1620 920 -1610
rect 680 -1710 920 -1700
rect 680 -1890 690 -1710
rect 910 -1890 920 -1710
rect 680 -1900 920 -1890
rect 680 -2170 920 -2160
rect 680 -2350 690 -2170
rect 910 -2350 920 -2170
rect 680 -2360 920 -2350
rect 680 -2530 920 -2520
rect 680 -2710 690 -2530
rect 910 -2710 920 -2530
rect 680 -2720 920 -2710
rect 680 -2930 920 -2920
rect 680 -3110 690 -2930
rect 910 -3110 920 -2930
rect 680 -3120 920 -3110
rect 680 -3380 920 -3370
rect 680 -3560 690 -3380
rect 910 -3560 920 -3380
rect 680 -3570 920 -3560
rect 680 -3750 920 -3740
rect 680 -3930 690 -3750
rect 910 -3930 920 -3750
rect 680 -3940 920 -3930
rect 1080 -3770 1220 -1150
rect 10630 -1390 10650 -1140
rect 10760 -1390 10780 -1140
rect 11220 -880 11630 -860
rect 11220 -950 11240 -880
rect 11610 -950 11630 -880
rect 11220 -1240 11630 -950
rect 12720 -870 13130 -860
rect 12720 -940 12740 -870
rect 13110 -940 13130 -870
rect 12090 -1120 12190 -1110
rect 11220 -1250 11660 -1240
rect 11220 -1320 11240 -1250
rect 11640 -1320 11660 -1250
rect 11220 -1330 11660 -1320
rect 10630 -1430 10780 -1390
rect 12090 -1410 12100 -1120
rect 12180 -1410 12190 -1120
rect 12720 -1250 13130 -940
rect 14180 -870 14590 -860
rect 14180 -940 14200 -870
rect 14570 -940 14590 -870
rect 12720 -1320 12740 -1250
rect 13110 -1320 13130 -1250
rect 12720 -1330 13130 -1320
rect 13570 -1130 13670 -1110
rect 12090 -1570 12190 -1410
rect 10870 -1700 11510 -1570
rect 12090 -1680 12100 -1570
rect 12180 -1680 12190 -1570
rect 12090 -1690 12190 -1680
rect 13570 -1420 13580 -1130
rect 13660 -1420 13670 -1130
rect 14180 -1250 14590 -940
rect 15310 -870 15640 -860
rect 15310 -940 15330 -870
rect 15620 -940 15640 -870
rect 15750 -920 16710 -690
rect 14180 -1320 14190 -1250
rect 14580 -1320 14590 -1250
rect 14180 -1330 14590 -1320
rect 15040 -1110 15140 -1100
rect 13570 -1570 13670 -1420
rect 13570 -1680 13580 -1570
rect 13660 -1680 13670 -1570
rect 13570 -1690 13670 -1680
rect 15040 -1380 15050 -1110
rect 15130 -1380 15140 -1110
rect 15310 -1250 15640 -940
rect 15310 -1320 15320 -1250
rect 15630 -1320 15640 -1250
rect 15310 -1330 15640 -1320
rect 16510 -1120 16610 -1110
rect 15040 -1570 15140 -1380
rect 15040 -1680 15050 -1570
rect 15130 -1680 15140 -1570
rect 15040 -1690 15140 -1680
rect 16510 -1410 16520 -1120
rect 16600 -1410 16610 -1120
rect 16510 -1570 16610 -1410
rect 16510 -1680 16520 -1570
rect 16600 -1680 16610 -1570
rect 16510 -1690 16610 -1680
rect 19620 -1450 20030 -1420
rect 7600 -2000 7790 -1990
rect 7600 -2240 7650 -2000
rect 7780 -2240 7790 -2000
rect 10870 -2050 11020 -1700
rect 11380 -2050 11510 -1700
rect 19620 -1830 19650 -1450
rect 20000 -1830 20030 -1450
rect 1080 -3910 1090 -3770
rect 1210 -3910 1220 -3770
rect 1080 -3940 1220 -3910
rect 7600 -8060 7790 -2240
rect 8980 -2120 9470 -2090
rect 8980 -2380 9010 -2120
rect 9440 -2380 9470 -2120
rect 10870 -2160 11510 -2050
rect 15390 -2110 16350 -1850
rect 19620 -1860 20030 -1830
rect 8980 -2410 9470 -2380
rect 15390 -2460 15700 -2110
rect 16060 -2460 16350 -2110
rect 10300 -2780 10850 -2750
rect 15390 -2760 16350 -2460
rect 10300 -3160 10330 -2780
rect 10820 -3160 10850 -2780
rect 10300 -3190 10850 -3160
rect 9960 -4780 10390 -4750
rect 9960 -5160 9990 -4780
rect 10360 -5160 10390 -4780
rect 9960 -5190 10390 -5160
rect 9350 -7300 9830 -7270
rect 9350 -7680 9380 -7300
rect 9800 -7680 9830 -7300
rect 9350 -7710 9830 -7680
rect 7600 -8180 7610 -8060
rect 7780 -8180 7790 -8060
rect 7600 -8190 7790 -8180
rect 680 -8770 920 -8760
rect 680 -8950 690 -8770
rect 910 -8950 920 -8770
rect 680 -8960 920 -8950
rect 680 -9100 920 -9090
rect 680 -9280 690 -9100
rect 910 -9280 920 -9100
rect 680 -9290 920 -9280
rect 680 -9590 920 -9580
rect 680 -9770 690 -9590
rect 910 -9770 920 -9590
rect 680 -9780 920 -9770
rect 680 -9870 920 -9860
rect 680 -10050 690 -9870
rect 910 -10050 920 -9870
rect 680 -10060 920 -10050
rect 680 -10330 920 -10320
rect 680 -10510 690 -10330
rect 910 -10510 920 -10330
rect 680 -10520 920 -10510
rect 680 -10690 920 -10680
rect 680 -10870 690 -10690
rect 910 -10870 920 -10690
rect 680 -10880 920 -10870
rect 680 -11090 920 -11080
rect 680 -11270 690 -11090
rect 910 -11270 920 -11090
rect 680 -11280 920 -11270
rect 680 -11540 920 -11530
rect 680 -11720 690 -11540
rect 910 -11720 920 -11540
rect 680 -11730 920 -11720
rect 680 -11910 920 -11900
rect 680 -12090 690 -11910
rect 910 -12090 920 -11910
rect 680 -12100 920 -12090
rect 1080 -11930 1220 -9310
rect 1080 -12070 1090 -11930
rect 1210 -12070 1220 -11930
rect 1080 -12100 1220 -12070
rect 9500 -13550 9640 -7710
rect 9810 -9890 9950 -9880
rect 9810 -10010 9820 -9890
rect 9940 -10010 9950 -9890
rect 9810 -13010 9950 -10010
rect 10080 -9890 10220 -5190
rect 10080 -10010 10090 -9890
rect 10210 -10010 10220 -9890
rect 10080 -10020 10220 -10010
rect 10330 -5760 10430 -5750
rect 10330 -5870 10340 -5760
rect 10420 -5870 10430 -5760
rect 10330 -10790 10430 -5870
rect 10500 -5760 10600 -3190
rect 10680 -4610 19310 -4580
rect 10680 -5180 10690 -4610
rect 19280 -5180 19310 -4610
rect 10680 -5210 19310 -5180
rect 13180 -5320 13270 -5310
rect 13180 -5410 13190 -5320
rect 13260 -5410 13270 -5320
rect 13180 -5680 13270 -5410
rect 10500 -5870 10510 -5760
rect 10590 -5870 10600 -5760
rect 10500 -5880 10600 -5870
rect 10900 -5760 10980 -5750
rect 10900 -5870 10910 -5760
rect 10970 -5870 10980 -5760
rect 10900 -5880 10980 -5870
rect 13180 -5870 13190 -5680
rect 13260 -5870 13270 -5680
rect 13450 -5320 14360 -5310
rect 13450 -5410 13460 -5320
rect 14350 -5410 14360 -5320
rect 13450 -5740 14360 -5410
rect 14900 -5320 15800 -5310
rect 14900 -5410 14910 -5320
rect 15790 -5410 15800 -5320
rect 13450 -5820 13460 -5740
rect 14350 -5820 14360 -5740
rect 13450 -5830 14360 -5820
rect 14660 -5660 14750 -5650
rect 13180 -5880 13270 -5870
rect 14660 -5870 14670 -5660
rect 14740 -5870 14750 -5660
rect 14900 -5740 15800 -5410
rect 16370 -5320 17270 -5310
rect 16370 -5410 16380 -5320
rect 17260 -5410 17270 -5320
rect 14900 -5820 14910 -5740
rect 15790 -5820 15800 -5740
rect 14900 -5830 15800 -5820
rect 16130 -5670 16220 -5660
rect 14660 -6100 14750 -5870
rect 14660 -6180 14670 -6100
rect 14740 -6180 14750 -6100
rect 14660 -6190 14750 -6180
rect 16130 -5870 16140 -5670
rect 16210 -5870 16220 -5670
rect 16370 -5750 17270 -5410
rect 17840 -5320 18640 -5310
rect 17840 -5410 17850 -5320
rect 18630 -5410 18640 -5320
rect 16370 -5820 16380 -5750
rect 17260 -5820 17270 -5750
rect 16370 -5830 17270 -5820
rect 17610 -5670 17690 -5660
rect 16130 -6100 16220 -5870
rect 16130 -6180 16140 -6100
rect 16210 -6180 16220 -6100
rect 16130 -6190 16220 -6180
rect 17680 -5880 17690 -5670
rect 17840 -5749 18640 -5410
rect 17840 -5821 17852 -5749
rect 18632 -5821 18640 -5749
rect 17840 -5831 18640 -5821
rect 19070 -5670 19160 -5660
rect 17610 -6100 17690 -5880
rect 17610 -6180 17620 -6100
rect 17680 -6180 17690 -6100
rect 17610 -6190 17690 -6180
rect 19070 -5880 19080 -5670
rect 19150 -5880 19160 -5670
rect 19070 -6100 19160 -5880
rect 19070 -6180 19080 -6100
rect 19150 -6180 19160 -6100
rect 19070 -6190 19160 -6180
rect 19620 -5950 20030 -5920
rect 10660 -6310 19310 -6280
rect 10660 -6880 10690 -6310
rect 19280 -6880 19310 -6310
rect 19620 -6330 19650 -5950
rect 20000 -6330 20030 -5950
rect 19620 -6360 20030 -6330
rect 10660 -6910 19310 -6880
rect 10664 -8748 19314 -8718
rect 10664 -9318 10694 -8748
rect 19284 -9318 19314 -8748
rect 10664 -9348 19314 -9318
rect 13184 -9458 13274 -9448
rect 13184 -9548 13194 -9458
rect 13264 -9548 13274 -9458
rect 13184 -9818 13274 -9548
rect 10900 -9890 10980 -9880
rect 10900 -10010 10910 -9890
rect 10970 -10010 10980 -9890
rect 10900 -10020 10980 -10010
rect 13184 -10008 13194 -9818
rect 13264 -10008 13274 -9818
rect 13454 -9458 14364 -9448
rect 13454 -9548 13464 -9458
rect 14354 -9548 14364 -9458
rect 13454 -9878 14364 -9548
rect 14904 -9458 15804 -9448
rect 14904 -9548 14914 -9458
rect 15794 -9548 15804 -9458
rect 13454 -9958 13464 -9878
rect 14354 -9958 14364 -9878
rect 13454 -9968 14364 -9958
rect 14664 -9798 14754 -9788
rect 13184 -10018 13274 -10008
rect 14664 -10008 14674 -9798
rect 14744 -10008 14754 -9798
rect 14904 -9878 15804 -9548
rect 16374 -9458 17274 -9448
rect 16374 -9548 16384 -9458
rect 17264 -9548 17274 -9458
rect 14904 -9958 14914 -9878
rect 15794 -9958 15804 -9878
rect 14904 -9968 15804 -9958
rect 16134 -9808 16224 -9798
rect 14664 -10238 14754 -10008
rect 14664 -10318 14674 -10238
rect 14744 -10318 14754 -10238
rect 14664 -10328 14754 -10318
rect 16134 -10008 16144 -9808
rect 16214 -10008 16224 -9808
rect 16374 -9888 17274 -9548
rect 17844 -9458 18644 -9448
rect 17844 -9548 17854 -9458
rect 18634 -9548 18644 -9458
rect 16374 -9958 16384 -9888
rect 17264 -9958 17274 -9888
rect 16374 -9968 17274 -9958
rect 17614 -9808 17694 -9798
rect 16134 -10238 16224 -10008
rect 16134 -10318 16144 -10238
rect 16214 -10318 16224 -10238
rect 16134 -10328 16224 -10318
rect 17684 -10018 17694 -9808
rect 17844 -9887 18644 -9548
rect 17844 -9959 17856 -9887
rect 18636 -9959 18644 -9887
rect 17844 -9969 18644 -9959
rect 19074 -9808 19164 -9798
rect 17614 -10238 17694 -10018
rect 17614 -10318 17624 -10238
rect 17684 -10318 17694 -10238
rect 17614 -10328 17694 -10318
rect 19074 -10018 19084 -9808
rect 19154 -10018 19164 -9808
rect 19074 -10238 19164 -10018
rect 19074 -10318 19084 -10238
rect 19154 -10318 19164 -10238
rect 19074 -10328 19164 -10318
rect 19620 -10110 20030 -10080
rect 10664 -10448 19314 -10418
rect 10290 -10820 10510 -10790
rect 10290 -11200 10320 -10820
rect 10480 -11200 10510 -10820
rect 10664 -11018 10694 -10448
rect 19284 -11018 19314 -10448
rect 19620 -10490 19650 -10110
rect 20000 -10490 20030 -10110
rect 19620 -10520 20030 -10490
rect 10664 -11048 19314 -11018
rect 10290 -11230 10510 -11200
rect 10660 -12400 19310 -12370
rect 10660 -12970 10690 -12400
rect 19280 -12970 19310 -12400
rect 10660 -13000 19310 -12970
rect 9810 -13220 9820 -13010
rect 9940 -13220 9950 -13010
rect 9810 -13230 9950 -13220
rect 13180 -13110 13270 -13100
rect 13180 -13200 13190 -13110
rect 13260 -13200 13270 -13110
rect 13180 -13470 13270 -13200
rect 9500 -13660 9510 -13550
rect 9630 -13660 9640 -13550
rect 9500 -13670 9640 -13660
rect 10150 -13550 10320 -13540
rect 10150 -13660 10160 -13550
rect 10310 -13660 10320 -13550
rect 10150 -15310 10320 -13660
rect 10890 -13550 10980 -13540
rect 10890 -13660 10900 -13550
rect 10970 -13660 10980 -13550
rect 10890 -13670 10980 -13660
rect 13180 -13660 13190 -13470
rect 13260 -13660 13270 -13470
rect 13450 -13110 14360 -13100
rect 13450 -13200 13460 -13110
rect 14350 -13200 14360 -13110
rect 13450 -13530 14360 -13200
rect 14900 -13110 15800 -13100
rect 14900 -13200 14910 -13110
rect 15790 -13200 15800 -13110
rect 13450 -13610 13460 -13530
rect 14350 -13610 14360 -13530
rect 13450 -13620 14360 -13610
rect 14660 -13450 14750 -13440
rect 13180 -13670 13270 -13660
rect 14660 -13660 14670 -13450
rect 14740 -13660 14750 -13450
rect 14900 -13530 15800 -13200
rect 16370 -13110 17270 -13100
rect 16370 -13200 16380 -13110
rect 17260 -13200 17270 -13110
rect 14900 -13610 14910 -13530
rect 15790 -13610 15800 -13530
rect 14900 -13620 15800 -13610
rect 16130 -13460 16220 -13450
rect 14660 -13890 14750 -13660
rect 14660 -13970 14670 -13890
rect 14740 -13970 14750 -13890
rect 14660 -13980 14750 -13970
rect 16130 -13660 16140 -13460
rect 16210 -13660 16220 -13460
rect 16370 -13540 17270 -13200
rect 17840 -13110 18640 -13100
rect 17840 -13200 17850 -13110
rect 18630 -13200 18640 -13110
rect 16370 -13610 16380 -13540
rect 17260 -13610 17270 -13540
rect 16370 -13620 17270 -13610
rect 17610 -13460 17690 -13450
rect 16130 -13890 16220 -13660
rect 16130 -13970 16140 -13890
rect 16210 -13970 16220 -13890
rect 16130 -13980 16220 -13970
rect 17680 -13670 17690 -13460
rect 17840 -13539 18640 -13200
rect 17840 -13611 17852 -13539
rect 18632 -13611 18640 -13539
rect 17840 -13621 18640 -13611
rect 19070 -13460 19160 -13450
rect 17610 -13890 17690 -13670
rect 17610 -13970 17620 -13890
rect 17680 -13970 17690 -13890
rect 17610 -13980 17690 -13970
rect 19070 -13670 19080 -13460
rect 19150 -13670 19160 -13460
rect 19070 -13890 19160 -13670
rect 19070 -13970 19080 -13890
rect 19150 -13970 19160 -13890
rect 19070 -13980 19160 -13970
rect 19620 -13740 20030 -13710
rect 10660 -14100 19310 -14070
rect 10660 -14670 10690 -14100
rect 19280 -14670 19310 -14100
rect 19620 -14120 19650 -13740
rect 20000 -14120 20030 -13740
rect 19620 -14150 20030 -14120
rect 10660 -14700 19310 -14670
rect 9980 -15340 10650 -15310
rect 9980 -15720 10010 -15340
rect 10620 -15720 10650 -15340
rect 9980 -15750 10650 -15720
<< via2 >>
rect 12830 -350 13270 80
rect 690 -790 910 -610
rect 16020 -690 16460 -260
rect 3090 -890 3210 -790
rect 690 -1120 910 -940
rect 10650 -970 10760 -880
rect 2840 -1090 2960 -970
rect 690 -1610 910 -1430
rect 690 -1890 910 -1710
rect 690 -2350 910 -2170
rect 690 -2710 910 -2530
rect 690 -3110 910 -2930
rect 690 -3560 910 -3380
rect 690 -3930 910 -3750
rect 11240 -950 11610 -880
rect 12740 -940 13110 -870
rect 14200 -940 14570 -870
rect 2590 -1590 2710 -1450
rect 12100 -1680 12180 -1570
rect 15330 -940 15620 -870
rect 13580 -1680 13660 -1570
rect 15050 -1680 15130 -1570
rect 16520 -1680 16600 -1570
rect 2340 -1870 2460 -1730
rect 11020 -2050 11380 -1700
rect 19650 -1830 20000 -1450
rect 1840 -2690 1960 -2550
rect 1590 -3090 1710 -2960
rect 1340 -3540 1460 -3400
rect 1090 -3910 1210 -3770
rect 9010 -2380 9440 -2120
rect 15700 -2460 16060 -2110
rect 10330 -3160 10820 -2780
rect 9990 -5160 10360 -4780
rect 9380 -7680 9800 -7300
rect 7610 -8180 7780 -8060
rect 690 -8950 910 -8770
rect 3090 -9050 3210 -8950
rect 690 -9280 910 -9100
rect 2840 -9250 2960 -9130
rect 690 -9770 910 -9590
rect 690 -10050 910 -9870
rect 690 -10510 910 -10330
rect 690 -10870 910 -10690
rect 690 -11270 910 -11090
rect 690 -11720 910 -11540
rect 690 -12090 910 -11910
rect 2590 -9750 2710 -9610
rect 1840 -10850 1960 -10710
rect 1590 -11250 1710 -11110
rect 1340 -11700 1460 -11560
rect 1090 -12070 1210 -11930
rect 10090 -10010 10210 -9890
rect 10690 -5180 19280 -4610
rect 13190 -5410 13260 -5320
rect 10510 -5870 10590 -5760
rect 10910 -5870 10970 -5760
rect 13460 -5410 14350 -5320
rect 14910 -5410 15790 -5320
rect 16380 -5410 17260 -5320
rect 14670 -6180 14740 -6100
rect 17850 -5410 18630 -5320
rect 16140 -6180 16210 -6100
rect 17620 -6180 17680 -6100
rect 19080 -6180 19150 -6100
rect 10690 -6880 19280 -6310
rect 19650 -6330 20000 -5950
rect 10694 -9318 19284 -8748
rect 13194 -9548 13264 -9458
rect 10910 -10010 10970 -9890
rect 13464 -9548 14354 -9458
rect 14914 -9548 15794 -9458
rect 16384 -9548 17264 -9458
rect 14674 -10318 14744 -10238
rect 17854 -9548 18634 -9458
rect 16144 -10318 16214 -10238
rect 17624 -10318 17684 -10238
rect 19084 -10318 19154 -10238
rect 10320 -11200 10480 -10820
rect 10694 -11018 19284 -10448
rect 19650 -10490 20000 -10110
rect 10690 -12970 19280 -12400
rect 9820 -13220 9940 -13010
rect 13190 -13200 13260 -13110
rect 9510 -13660 9630 -13550
rect 10900 -13660 10970 -13550
rect 13460 -13200 14350 -13110
rect 14910 -13200 15790 -13110
rect 16380 -13200 17260 -13110
rect 14670 -13970 14740 -13890
rect 17850 -13200 18630 -13110
rect 16140 -13970 16210 -13890
rect 17620 -13970 17680 -13890
rect 19080 -13970 19150 -13890
rect 10690 -14670 19280 -14100
rect 19650 -14120 20000 -13740
rect 10010 -15720 10620 -15340
<< metal3 >>
rect 12570 80 13530 350
rect 12570 -350 12830 80
rect 13270 -350 13530 80
rect 12570 -560 13530 -350
rect 15750 -260 16710 -10
rect 680 -610 920 -600
rect 680 -790 690 -610
rect 910 -620 920 -610
rect 910 -780 1240 -620
rect 15750 -690 16020 -260
rect 16460 -690 16710 -260
rect 910 -790 920 -780
rect 680 -800 920 -790
rect 1080 -790 3220 -780
rect 1080 -890 3090 -790
rect 3210 -890 3220 -790
rect 1080 -900 3220 -890
rect 10630 -870 15640 -860
rect 10630 -880 12740 -870
rect 680 -940 920 -930
rect 680 -1120 690 -940
rect 910 -960 920 -940
rect 910 -970 2970 -960
rect 910 -1090 2840 -970
rect 2960 -1090 2970 -970
rect 10630 -970 10650 -880
rect 10760 -950 11240 -880
rect 11610 -940 12740 -880
rect 13110 -940 14200 -870
rect 14570 -940 15330 -870
rect 15620 -940 15640 -870
rect 15750 -920 16710 -690
rect 11610 -950 15640 -940
rect 10760 -960 15640 -950
rect 10760 -970 10780 -960
rect 10630 -990 10780 -970
rect 910 -1100 2970 -1090
rect 910 -1120 920 -1100
rect 680 -1130 920 -1120
rect 680 -1430 920 -1420
rect 680 -1610 690 -1430
rect 910 -1440 920 -1430
rect 910 -1450 2720 -1440
rect 910 -1590 2590 -1450
rect 2710 -1590 2720 -1450
rect 17450 -1450 20030 -1420
rect 17450 -1560 19650 -1450
rect 12090 -1570 19650 -1560
rect 910 -1600 2720 -1590
rect 910 -1610 920 -1600
rect 680 -1620 920 -1610
rect 10870 -1700 11510 -1570
rect 12090 -1680 12100 -1570
rect 12180 -1680 13580 -1570
rect 13660 -1680 15050 -1570
rect 15130 -1680 16520 -1570
rect 16600 -1680 19650 -1570
rect 12090 -1690 19650 -1680
rect 680 -1710 920 -1700
rect 680 -1890 690 -1710
rect 910 -1720 920 -1710
rect 910 -1730 2470 -1720
rect 910 -1870 2340 -1730
rect 2460 -1870 2470 -1730
rect 910 -1880 2470 -1870
rect 910 -1890 920 -1880
rect 680 -1900 920 -1890
rect 10870 -2050 11020 -1700
rect 11380 -2050 11510 -1700
rect 17450 -1830 19650 -1690
rect 20000 -1830 20030 -1450
rect 8980 -2120 9470 -2090
rect 680 -2170 920 -2160
rect 680 -2350 690 -2170
rect 910 -2180 920 -2170
rect 910 -2340 2220 -2180
rect 910 -2350 920 -2340
rect 680 -2360 920 -2350
rect 8980 -2380 9010 -2120
rect 9440 -2380 9470 -2120
rect 10870 -2160 11510 -2050
rect 15390 -2110 16350 -1850
rect 17450 -1860 20030 -1830
rect 8980 -2410 9470 -2380
rect 15390 -2460 15700 -2110
rect 16060 -2460 16350 -2110
rect 680 -2530 920 -2520
rect 680 -2710 690 -2530
rect 910 -2540 920 -2530
rect 910 -2550 1970 -2540
rect 910 -2690 1840 -2550
rect 1960 -2690 1970 -2550
rect 910 -2700 1970 -2690
rect 910 -2710 920 -2700
rect 680 -2720 920 -2710
rect 7920 -2780 10850 -2750
rect 15390 -2760 16350 -2460
rect 680 -2930 920 -2920
rect 680 -3110 690 -2930
rect 910 -2950 920 -2930
rect 910 -2960 1720 -2950
rect 910 -3090 1590 -2960
rect 1710 -3090 1720 -2960
rect 910 -3100 1720 -3090
rect 910 -3110 920 -3100
rect 680 -3120 920 -3110
rect 7920 -3160 10330 -2780
rect 10820 -3160 10850 -2780
rect 7920 -3190 10850 -3160
rect 680 -3380 920 -3370
rect 680 -3560 690 -3380
rect 910 -3390 920 -3380
rect 910 -3400 1470 -3390
rect 910 -3540 1340 -3400
rect 1460 -3540 1470 -3400
rect 910 -3550 1470 -3540
rect 910 -3560 920 -3550
rect 680 -3570 920 -3560
rect 680 -3750 920 -3740
rect 680 -3930 690 -3750
rect 910 -3760 920 -3750
rect 910 -3770 1220 -3760
rect 910 -3910 1090 -3770
rect 1210 -3910 1220 -3770
rect 910 -3920 1220 -3910
rect 910 -3930 920 -3920
rect 680 -3940 920 -3930
rect 10660 -4610 19310 -4580
rect 8230 -4780 10390 -4750
rect 8230 -5160 9990 -4780
rect 10360 -5160 10390 -4780
rect 8230 -5190 10390 -5160
rect 10660 -5180 10690 -4610
rect 19280 -5180 19310 -4610
rect 10660 -5210 19310 -5180
rect 13180 -5320 18640 -5310
rect 13180 -5410 13190 -5320
rect 13260 -5410 13460 -5320
rect 14350 -5410 14910 -5320
rect 15790 -5410 16380 -5320
rect 17260 -5410 17850 -5320
rect 18630 -5410 18640 -5320
rect 13180 -5420 18640 -5410
rect 10500 -5760 10980 -5750
rect 10500 -5870 10510 -5760
rect 10590 -5870 10910 -5760
rect 10970 -5870 10980 -5760
rect 10500 -5880 10980 -5870
rect 19620 -5950 20030 -5920
rect 19620 -6090 19650 -5950
rect 14660 -6100 19650 -6090
rect 14660 -6180 14670 -6100
rect 14740 -6180 16140 -6100
rect 16210 -6180 17620 -6100
rect 17680 -6180 19080 -6100
rect 19150 -6180 19650 -6100
rect 14660 -6190 19650 -6180
rect 10660 -6310 19310 -6280
rect 10660 -6880 10690 -6310
rect 19280 -6880 19310 -6310
rect 19620 -6330 19650 -6190
rect 20000 -6330 20030 -5950
rect 19620 -6360 20030 -6330
rect 10660 -6910 19310 -6880
rect 7850 -7300 9830 -7270
rect 7850 -7680 9380 -7300
rect 9800 -7680 9830 -7300
rect 7850 -7710 9830 -7680
rect 6630 -8060 7790 -8050
rect 6630 -8180 7610 -8060
rect 7780 -8180 7790 -8060
rect 6630 -8190 7790 -8180
rect 10664 -8748 19314 -8718
rect 680 -8770 920 -8760
rect 680 -8950 690 -8770
rect 910 -8780 920 -8770
rect 910 -8940 1240 -8780
rect 910 -8950 920 -8940
rect 680 -8960 920 -8950
rect 1080 -8950 3220 -8940
rect 1080 -9050 3090 -8950
rect 3210 -9050 3220 -8950
rect 1080 -9060 3220 -9050
rect 680 -9100 920 -9090
rect 680 -9280 690 -9100
rect 910 -9120 920 -9100
rect 910 -9130 2970 -9120
rect 910 -9250 2840 -9130
rect 2960 -9250 2970 -9130
rect 910 -9260 2970 -9250
rect 910 -9280 920 -9260
rect 680 -9290 920 -9280
rect 10664 -9318 10694 -8748
rect 19284 -9318 19314 -8748
rect 10664 -9348 19314 -9318
rect 13184 -9458 18644 -9448
rect 13184 -9548 13194 -9458
rect 13264 -9548 13464 -9458
rect 14354 -9548 14914 -9458
rect 15794 -9548 16384 -9458
rect 17264 -9548 17854 -9458
rect 18634 -9548 18644 -9458
rect 13184 -9558 18644 -9548
rect 680 -9590 920 -9580
rect 680 -9770 690 -9590
rect 910 -9600 920 -9590
rect 910 -9610 2720 -9600
rect 910 -9750 2590 -9610
rect 2710 -9750 2720 -9610
rect 910 -9760 2720 -9750
rect 910 -9770 920 -9760
rect 680 -9780 920 -9770
rect 680 -9870 920 -9860
rect 680 -10050 690 -9870
rect 910 -9880 920 -9870
rect 910 -10040 2470 -9880
rect 10080 -9890 10980 -9880
rect 10080 -10010 10090 -9890
rect 10210 -10010 10910 -9890
rect 10970 -10010 10980 -9890
rect 10080 -10020 10980 -10010
rect 910 -10050 920 -10040
rect 680 -10060 920 -10050
rect 2250 -10100 2470 -10040
rect 19620 -10110 20030 -10080
rect 19620 -10228 19650 -10110
rect 14664 -10238 19650 -10228
rect 14664 -10318 14674 -10238
rect 14744 -10318 16144 -10238
rect 16214 -10318 17624 -10238
rect 17684 -10318 19084 -10238
rect 19154 -10318 19650 -10238
rect 680 -10330 920 -10320
rect 14664 -10328 19650 -10318
rect 680 -10510 690 -10330
rect 910 -10340 920 -10330
rect 910 -10500 2220 -10340
rect 10664 -10448 19314 -10418
rect 910 -10510 920 -10500
rect 680 -10520 920 -10510
rect 680 -10690 920 -10680
rect 680 -10870 690 -10690
rect 910 -10700 920 -10690
rect 910 -10710 1970 -10700
rect 910 -10850 1840 -10710
rect 1960 -10850 1970 -10710
rect 910 -10860 1970 -10850
rect 8330 -10820 10510 -10790
rect 910 -10870 920 -10860
rect 680 -10880 920 -10870
rect 680 -11090 920 -11080
rect 680 -11270 690 -11090
rect 910 -11100 920 -11090
rect 910 -11110 1720 -11100
rect 910 -11250 1590 -11110
rect 1710 -11250 1720 -11110
rect 8330 -11200 10320 -10820
rect 10480 -11200 10510 -10820
rect 10664 -11018 10694 -10448
rect 19284 -11018 19314 -10448
rect 19620 -10490 19650 -10328
rect 20000 -10490 20030 -10110
rect 19620 -10520 20030 -10490
rect 10664 -11048 19314 -11018
rect 8330 -11230 10510 -11200
rect 910 -11260 1720 -11250
rect 910 -11270 920 -11260
rect 680 -11280 920 -11270
rect 680 -11540 920 -11530
rect 680 -11720 690 -11540
rect 910 -11550 920 -11540
rect 910 -11560 1470 -11550
rect 910 -11700 1340 -11560
rect 1460 -11700 1470 -11560
rect 910 -11710 1470 -11700
rect 910 -11720 920 -11710
rect 680 -11730 920 -11720
rect 680 -11910 920 -11900
rect 680 -12090 690 -11910
rect 910 -11920 920 -11910
rect 910 -11930 1220 -11920
rect 910 -12070 1090 -11930
rect 1210 -12070 1220 -11930
rect 910 -12080 1220 -12070
rect 910 -12090 920 -12080
rect 680 -12100 920 -12090
rect 10660 -12400 19310 -12370
rect 8250 -13010 9950 -12790
rect 10660 -12970 10690 -12400
rect 19280 -12970 19310 -12400
rect 10660 -13000 19310 -12970
rect 8250 -13220 9820 -13010
rect 9940 -13220 9950 -13010
rect 13180 -13110 18640 -13100
rect 13180 -13200 13190 -13110
rect 13260 -13200 13460 -13110
rect 14350 -13200 14910 -13110
rect 15790 -13200 16380 -13110
rect 17260 -13200 17850 -13110
rect 18630 -13200 18640 -13110
rect 13180 -13210 18640 -13200
rect 8250 -13230 9950 -13220
rect 9500 -13550 10980 -13540
rect 9500 -13660 9510 -13550
rect 9630 -13660 10900 -13550
rect 10970 -13660 10980 -13550
rect 9500 -13670 10980 -13660
rect 19620 -13740 20030 -13710
rect 19620 -13880 19650 -13740
rect 14660 -13890 19650 -13880
rect 14660 -13970 14670 -13890
rect 14740 -13970 16140 -13890
rect 16210 -13970 17620 -13890
rect 17680 -13970 19080 -13890
rect 19150 -13970 19650 -13890
rect 14660 -13980 19650 -13970
rect 10660 -14100 19310 -14070
rect 10660 -14670 10690 -14100
rect 19280 -14670 19310 -14100
rect 19620 -14120 19650 -13980
rect 20000 -14120 20030 -13740
rect 19620 -14150 20030 -14120
rect 10660 -14700 19310 -14670
rect 7850 -15340 10650 -15310
rect 7850 -15720 10010 -15340
rect 10620 -15720 10650 -15340
rect 7850 -15750 10650 -15720
<< via3 >>
rect 12830 -350 13270 80
rect 16020 -690 16460 -260
rect 11020 -2050 11380 -1700
rect 9010 -2380 9440 -2120
rect 15700 -2460 16060 -2110
rect 10690 -5180 19280 -4610
rect 10690 -6880 19280 -6310
rect 10694 -9318 19284 -8748
rect 10694 -11018 19284 -10448
rect 10690 -12970 19280 -12400
rect 10690 -14670 19280 -14100
<< metal4 >>
rect 4140 -500 8470 350
rect 4140 -15670 4950 -500
rect 7780 -1470 8470 -500
rect 12570 80 13530 350
rect 12570 -350 12830 80
rect 13270 -350 13530 80
rect 12570 -560 13530 -350
rect 15750 -260 16710 -10
rect 15750 -690 16020 -260
rect 16460 -690 16710 -260
rect 15750 -920 16710 -690
rect 7780 -1700 16350 -1470
rect 7780 -1850 11020 -1700
rect 7780 -6280 8470 -1850
rect 10870 -2050 11020 -1850
rect 11380 -1850 16350 -1700
rect 11380 -2050 11510 -1850
rect 8980 -2120 9470 -2090
rect 8980 -2380 9010 -2120
rect 9440 -2380 9470 -2120
rect 10870 -2160 11510 -2050
rect 15390 -2110 16350 -1850
rect 8980 -2410 9470 -2380
rect 15390 -2460 15700 -2110
rect 16060 -2460 16350 -2110
rect 15390 -2760 16350 -2460
rect 10660 -4610 19310 -4580
rect 10660 -5180 10690 -4610
rect 19280 -5180 19310 -4610
rect 10660 -5210 19310 -5180
rect 7780 -6310 19310 -6280
rect 7780 -6880 10690 -6310
rect 19280 -6880 19310 -6310
rect 7780 -6910 19310 -6880
rect 7780 -10410 8470 -6910
rect 10664 -8748 19314 -8718
rect 10664 -9318 10694 -8748
rect 19284 -9318 19314 -8748
rect 10664 -9348 19314 -9318
rect 7780 -10448 19320 -10410
rect 7780 -11018 10694 -10448
rect 19284 -11018 19320 -10448
rect 7780 -11050 19320 -11018
rect 7780 -14070 8470 -11050
rect 10660 -12400 19310 -12370
rect 10660 -12970 10690 -12400
rect 19280 -12970 19310 -12400
rect 10660 -13000 19310 -12970
rect 7780 -14100 19310 -14070
rect 7780 -14670 10690 -14100
rect 19280 -14670 19310 -14100
rect 7780 -14700 19310 -14670
<< via4 >>
rect 12830 -350 13270 80
rect 16020 -690 16460 -260
rect 9010 -2380 9440 -2120
rect 10690 -5180 19280 -4610
rect 10694 -9318 19284 -8748
rect 10690 -12970 19280 -12400
<< metal5 >>
rect 7160 80 13530 350
rect 7160 -350 12830 80
rect 13270 10 13530 80
rect 13270 -260 17310 10
rect 13270 -350 16020 -260
rect 7160 -690 16020 -350
rect 16460 -690 17310 -260
rect 7160 -1130 17310 -690
rect 7160 -1760 8400 -1130
rect 7160 -2120 9470 -1760
rect 7160 -2380 9010 -2120
rect 9440 -2380 9470 -2120
rect 7160 -2410 9470 -2380
rect 7160 -4580 8400 -2410
rect 7160 -4610 19310 -4580
rect 7160 -5180 10690 -4610
rect 19280 -5180 19310 -4610
rect 7160 -5210 19310 -5180
rect 7160 -8710 8400 -5210
rect 7160 -8748 19320 -8710
rect 7160 -9318 10694 -8748
rect 19284 -9318 19320 -8748
rect 7160 -9350 19320 -9318
rect 7160 -12370 8400 -9350
rect 7160 -12400 19310 -12370
rect 7160 -12970 10690 -12400
rect 19280 -12970 19310 -12400
rect 7160 -13000 19310 -12970
rect 7160 -15300 8400 -13000
use sky130_fd_sc_hd__or2_1  x1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 10708 0 1 -10162
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  x2
timestamp 1701704242
transform 1 0 10708 0 1 -13812
box -38 -48 498 592
use 8to3_Priority_Encoder_v0p2p0  x3
timestamp 1713495814
transform 1 0 4960 0 1 -8740
box -3910 -7130 3570 700
use sky130_fd_sc_hd__inv_16  x4 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 12288 0 1 -1522
box -38 -48 1510 592
use 8to3_Priority_Encoder_v0p2p0  x5
timestamp 1713495814
transform 1 0 4960 0 1 -700
box -3910 -7130 3570 700
use sky130_fd_sc_hd__inv_16  x6
timestamp 1701704242
transform 1 0 10816 0 1 -1522
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_1  x7 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 8658 0 -1 -1598
box -38 -48 314 592
use sky130_fd_sc_hd__inv_16  x8
timestamp 1701704242
transform 1 0 13760 0 1 -1522
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_16  x9
timestamp 1701704242
transform 1 0 15232 0 1 -1522
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_16  x10
timestamp 1701704242
transform 1 0 13376 0 1 -6022
box -38 -48 1510 592
use sky130_fd_sc_hd__or2_1  x11
timestamp 1701704242
transform 1 0 10708 0 1 -6022
box -38 -48 498 592
use sky130_fd_sc_hd__inv_16  x12
timestamp 1701704242
transform 1 0 14848 0 1 -6022
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_16  x13
timestamp 1701704242
transform 1 0 16320 0 1 -6022
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_16  x14
timestamp 1701704242
transform 1 0 17792 0 1 -6022
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_16  x15
timestamp 1701704242
transform 1 0 13376 0 1 -10162
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_16  x16
timestamp 1701704242
transform 1 0 14848 0 1 -10162
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_16  x17
timestamp 1701704242
transform 1 0 16320 0 1 -10162
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_16  x18
timestamp 1701704242
transform 1 0 17792 0 1 -10162
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_16  x19
timestamp 1701704242
transform 1 0 13376 0 1 -13812
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_1  x20
timestamp 1701704242
transform 1 0 11168 0 1 -13812
box -38 -48 314 592
use sky130_fd_sc_hd__inv_4  x21 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 11444 0 1 -13812
box -38 -48 498 592
use sky130_fd_sc_hd__inv_16  x22
timestamp 1701704242
transform 1 0 11904 0 1 -13812
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_16  x23
timestamp 1701704242
transform 1 0 14848 0 1 -13812
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_16  x24
timestamp 1701704242
transform 1 0 16320 0 1 -13812
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_16  x25
timestamp 1701704242
transform 1 0 17792 0 1 -13812
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_1  x27
timestamp 1701704242
transform 1 0 11168 0 1 -10162
box -38 -48 314 592
use sky130_fd_sc_hd__inv_4  x28
timestamp 1701704242
transform 1 0 11444 0 1 -10162
box -38 -48 498 592
use sky130_fd_sc_hd__inv_16  x29
timestamp 1701704242
transform 1 0 11904 0 1 -10162
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_1  x34
timestamp 1701704242
transform 1 0 11168 0 1 -6022
box -38 -48 314 592
use sky130_fd_sc_hd__inv_4  x35
timestamp 1701704242
transform 1 0 11444 0 1 -6022
box -38 -48 498 592
use sky130_fd_sc_hd__inv_16  x36
timestamp 1701704242
transform 1 0 11904 0 1 -6022
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_1  x41
timestamp 1701704242
transform 1 0 8608 0 1 -1522
box -38 -48 314 592
use sky130_fd_sc_hd__inv_4  x42
timestamp 1701704242
transform 1 0 8884 0 1 -1522
box -38 -48 498 592
use sky130_fd_sc_hd__inv_16  x43
timestamp 1701704242
transform 1 0 9344 0 1 -1522
box -38 -48 1510 592
<< labels >>
flabel metal1 480 -1130 680 -930 0 FreeSans 256 0 0 0 I15
port 2 nsew
flabel metal1 480 -800 680 -600 0 FreeSans 256 0 0 0 EI
port 1 nsew
flabel metal1 480 -1620 680 -1420 0 FreeSans 256 0 0 0 I14
port 3 nsew
flabel metal1 480 -1900 680 -1700 0 FreeSans 256 0 0 0 I13
port 4 nsew
flabel metal1 480 -2360 680 -2160 0 FreeSans 256 0 0 0 I12
port 5 nsew
flabel metal1 480 -2720 680 -2520 0 FreeSans 256 0 0 0 I11
port 6 nsew
flabel metal1 480 -3120 680 -2920 0 FreeSans 256 0 0 0 I10
port 7 nsew
flabel metal1 480 -3570 680 -3370 0 FreeSans 256 0 0 0 I9
port 9 nsew
flabel metal1 480 -3940 680 -3740 0 FreeSans 256 0 0 0 I8
port 10 nsew
flabel metal1 480 -12100 680 -11900 0 FreeSans 256 0 0 0 I0
port 19 nsew
flabel metal1 470 -11730 670 -11530 0 FreeSans 256 0 0 0 I1
port 18 nsew
flabel metal1 470 -11280 670 -11080 0 FreeSans 256 0 0 0 I2
port 17 nsew
flabel metal1 470 -10880 670 -10680 0 FreeSans 256 0 0 0 I3
port 16 nsew
flabel metal1 470 -10520 670 -10320 0 FreeSans 256 0 0 0 I4
port 14 nsew
flabel metal1 470 -10060 670 -9860 0 FreeSans 256 0 0 0 I5
port 13 nsew
flabel metal1 470 -9780 670 -9580 0 FreeSans 256 0 0 0 I6
port 12 nsew
flabel metal1 470 -9290 670 -9090 0 FreeSans 256 0 0 0 I7
port 11 nsew
flabel metal1 20030 -6260 20230 -6060 0 FreeSans 256 0 0 0 A2
port 8 nsew
flabel metal1 20030 -1730 20230 -1530 0 FreeSans 256 0 0 0 A3
port 0 nsew
flabel metal1 20030 -10410 20230 -10210 0 FreeSans 256 0 0 0 A1
port 15 nsew
flabel metal1 20030 -14020 20230 -13820 0 FreeSans 256 0 0 0 A0
port 20 nsew
flabel metal5 7160 -15300 8400 350 0 FreeSans 512 0 0 0 VDD
port 21 n
flabel metal4 4140 -15670 4950 350 1 FreeSans 512 0 0 0 GND
port 22 n
<< end >>
