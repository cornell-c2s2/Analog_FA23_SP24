magic
tech sky130A
magscale 1 2
timestamp 1713140669
<< nwell >>
rect -3327 -719 3327 719
<< pmos >>
rect -3131 -500 -3031 500
rect -2973 -500 -2873 500
rect -2815 -500 -2715 500
rect -2657 -500 -2557 500
rect -2499 -500 -2399 500
rect -2341 -500 -2241 500
rect -2183 -500 -2083 500
rect -2025 -500 -1925 500
rect -1867 -500 -1767 500
rect -1709 -500 -1609 500
rect -1551 -500 -1451 500
rect -1393 -500 -1293 500
rect -1235 -500 -1135 500
rect -1077 -500 -977 500
rect -919 -500 -819 500
rect -761 -500 -661 500
rect -603 -500 -503 500
rect -445 -500 -345 500
rect -287 -500 -187 500
rect -129 -500 -29 500
rect 29 -500 129 500
rect 187 -500 287 500
rect 345 -500 445 500
rect 503 -500 603 500
rect 661 -500 761 500
rect 819 -500 919 500
rect 977 -500 1077 500
rect 1135 -500 1235 500
rect 1293 -500 1393 500
rect 1451 -500 1551 500
rect 1609 -500 1709 500
rect 1767 -500 1867 500
rect 1925 -500 2025 500
rect 2083 -500 2183 500
rect 2241 -500 2341 500
rect 2399 -500 2499 500
rect 2557 -500 2657 500
rect 2715 -500 2815 500
rect 2873 -500 2973 500
rect 3031 -500 3131 500
<< pdiff >>
rect -3189 488 -3131 500
rect -3189 -488 -3177 488
rect -3143 -488 -3131 488
rect -3189 -500 -3131 -488
rect -3031 488 -2973 500
rect -3031 -488 -3019 488
rect -2985 -488 -2973 488
rect -3031 -500 -2973 -488
rect -2873 488 -2815 500
rect -2873 -488 -2861 488
rect -2827 -488 -2815 488
rect -2873 -500 -2815 -488
rect -2715 488 -2657 500
rect -2715 -488 -2703 488
rect -2669 -488 -2657 488
rect -2715 -500 -2657 -488
rect -2557 488 -2499 500
rect -2557 -488 -2545 488
rect -2511 -488 -2499 488
rect -2557 -500 -2499 -488
rect -2399 488 -2341 500
rect -2399 -488 -2387 488
rect -2353 -488 -2341 488
rect -2399 -500 -2341 -488
rect -2241 488 -2183 500
rect -2241 -488 -2229 488
rect -2195 -488 -2183 488
rect -2241 -500 -2183 -488
rect -2083 488 -2025 500
rect -2083 -488 -2071 488
rect -2037 -488 -2025 488
rect -2083 -500 -2025 -488
rect -1925 488 -1867 500
rect -1925 -488 -1913 488
rect -1879 -488 -1867 488
rect -1925 -500 -1867 -488
rect -1767 488 -1709 500
rect -1767 -488 -1755 488
rect -1721 -488 -1709 488
rect -1767 -500 -1709 -488
rect -1609 488 -1551 500
rect -1609 -488 -1597 488
rect -1563 -488 -1551 488
rect -1609 -500 -1551 -488
rect -1451 488 -1393 500
rect -1451 -488 -1439 488
rect -1405 -488 -1393 488
rect -1451 -500 -1393 -488
rect -1293 488 -1235 500
rect -1293 -488 -1281 488
rect -1247 -488 -1235 488
rect -1293 -500 -1235 -488
rect -1135 488 -1077 500
rect -1135 -488 -1123 488
rect -1089 -488 -1077 488
rect -1135 -500 -1077 -488
rect -977 488 -919 500
rect -977 -488 -965 488
rect -931 -488 -919 488
rect -977 -500 -919 -488
rect -819 488 -761 500
rect -819 -488 -807 488
rect -773 -488 -761 488
rect -819 -500 -761 -488
rect -661 488 -603 500
rect -661 -488 -649 488
rect -615 -488 -603 488
rect -661 -500 -603 -488
rect -503 488 -445 500
rect -503 -488 -491 488
rect -457 -488 -445 488
rect -503 -500 -445 -488
rect -345 488 -287 500
rect -345 -488 -333 488
rect -299 -488 -287 488
rect -345 -500 -287 -488
rect -187 488 -129 500
rect -187 -488 -175 488
rect -141 -488 -129 488
rect -187 -500 -129 -488
rect -29 488 29 500
rect -29 -488 -17 488
rect 17 -488 29 488
rect -29 -500 29 -488
rect 129 488 187 500
rect 129 -488 141 488
rect 175 -488 187 488
rect 129 -500 187 -488
rect 287 488 345 500
rect 287 -488 299 488
rect 333 -488 345 488
rect 287 -500 345 -488
rect 445 488 503 500
rect 445 -488 457 488
rect 491 -488 503 488
rect 445 -500 503 -488
rect 603 488 661 500
rect 603 -488 615 488
rect 649 -488 661 488
rect 603 -500 661 -488
rect 761 488 819 500
rect 761 -488 773 488
rect 807 -488 819 488
rect 761 -500 819 -488
rect 919 488 977 500
rect 919 -488 931 488
rect 965 -488 977 488
rect 919 -500 977 -488
rect 1077 488 1135 500
rect 1077 -488 1089 488
rect 1123 -488 1135 488
rect 1077 -500 1135 -488
rect 1235 488 1293 500
rect 1235 -488 1247 488
rect 1281 -488 1293 488
rect 1235 -500 1293 -488
rect 1393 488 1451 500
rect 1393 -488 1405 488
rect 1439 -488 1451 488
rect 1393 -500 1451 -488
rect 1551 488 1609 500
rect 1551 -488 1563 488
rect 1597 -488 1609 488
rect 1551 -500 1609 -488
rect 1709 488 1767 500
rect 1709 -488 1721 488
rect 1755 -488 1767 488
rect 1709 -500 1767 -488
rect 1867 488 1925 500
rect 1867 -488 1879 488
rect 1913 -488 1925 488
rect 1867 -500 1925 -488
rect 2025 488 2083 500
rect 2025 -488 2037 488
rect 2071 -488 2083 488
rect 2025 -500 2083 -488
rect 2183 488 2241 500
rect 2183 -488 2195 488
rect 2229 -488 2241 488
rect 2183 -500 2241 -488
rect 2341 488 2399 500
rect 2341 -488 2353 488
rect 2387 -488 2399 488
rect 2341 -500 2399 -488
rect 2499 488 2557 500
rect 2499 -488 2511 488
rect 2545 -488 2557 488
rect 2499 -500 2557 -488
rect 2657 488 2715 500
rect 2657 -488 2669 488
rect 2703 -488 2715 488
rect 2657 -500 2715 -488
rect 2815 488 2873 500
rect 2815 -488 2827 488
rect 2861 -488 2873 488
rect 2815 -500 2873 -488
rect 2973 488 3031 500
rect 2973 -488 2985 488
rect 3019 -488 3031 488
rect 2973 -500 3031 -488
rect 3131 488 3189 500
rect 3131 -488 3143 488
rect 3177 -488 3189 488
rect 3131 -500 3189 -488
<< pdiffc >>
rect -3177 -488 -3143 488
rect -3019 -488 -2985 488
rect -2861 -488 -2827 488
rect -2703 -488 -2669 488
rect -2545 -488 -2511 488
rect -2387 -488 -2353 488
rect -2229 -488 -2195 488
rect -2071 -488 -2037 488
rect -1913 -488 -1879 488
rect -1755 -488 -1721 488
rect -1597 -488 -1563 488
rect -1439 -488 -1405 488
rect -1281 -488 -1247 488
rect -1123 -488 -1089 488
rect -965 -488 -931 488
rect -807 -488 -773 488
rect -649 -488 -615 488
rect -491 -488 -457 488
rect -333 -488 -299 488
rect -175 -488 -141 488
rect -17 -488 17 488
rect 141 -488 175 488
rect 299 -488 333 488
rect 457 -488 491 488
rect 615 -488 649 488
rect 773 -488 807 488
rect 931 -488 965 488
rect 1089 -488 1123 488
rect 1247 -488 1281 488
rect 1405 -488 1439 488
rect 1563 -488 1597 488
rect 1721 -488 1755 488
rect 1879 -488 1913 488
rect 2037 -488 2071 488
rect 2195 -488 2229 488
rect 2353 -488 2387 488
rect 2511 -488 2545 488
rect 2669 -488 2703 488
rect 2827 -488 2861 488
rect 2985 -488 3019 488
rect 3143 -488 3177 488
<< nsubdiff >>
rect -3291 649 -3195 683
rect 3195 649 3291 683
rect -3291 587 -3257 649
rect 3257 587 3291 649
rect -3291 -649 -3257 -587
rect 3257 -649 3291 -587
rect -3291 -683 -3195 -649
rect 3195 -683 3291 -649
<< nsubdiffcont >>
rect -3195 649 3195 683
rect -3291 -587 -3257 587
rect 3257 -587 3291 587
rect -3195 -683 3195 -649
<< poly >>
rect -3131 581 -3031 597
rect -3131 547 -3115 581
rect -3047 547 -3031 581
rect -3131 500 -3031 547
rect -2973 581 -2873 597
rect -2973 547 -2957 581
rect -2889 547 -2873 581
rect -2973 500 -2873 547
rect -2815 581 -2715 597
rect -2815 547 -2799 581
rect -2731 547 -2715 581
rect -2815 500 -2715 547
rect -2657 581 -2557 597
rect -2657 547 -2641 581
rect -2573 547 -2557 581
rect -2657 500 -2557 547
rect -2499 581 -2399 597
rect -2499 547 -2483 581
rect -2415 547 -2399 581
rect -2499 500 -2399 547
rect -2341 581 -2241 597
rect -2341 547 -2325 581
rect -2257 547 -2241 581
rect -2341 500 -2241 547
rect -2183 581 -2083 597
rect -2183 547 -2167 581
rect -2099 547 -2083 581
rect -2183 500 -2083 547
rect -2025 581 -1925 597
rect -2025 547 -2009 581
rect -1941 547 -1925 581
rect -2025 500 -1925 547
rect -1867 581 -1767 597
rect -1867 547 -1851 581
rect -1783 547 -1767 581
rect -1867 500 -1767 547
rect -1709 581 -1609 597
rect -1709 547 -1693 581
rect -1625 547 -1609 581
rect -1709 500 -1609 547
rect -1551 581 -1451 597
rect -1551 547 -1535 581
rect -1467 547 -1451 581
rect -1551 500 -1451 547
rect -1393 581 -1293 597
rect -1393 547 -1377 581
rect -1309 547 -1293 581
rect -1393 500 -1293 547
rect -1235 581 -1135 597
rect -1235 547 -1219 581
rect -1151 547 -1135 581
rect -1235 500 -1135 547
rect -1077 581 -977 597
rect -1077 547 -1061 581
rect -993 547 -977 581
rect -1077 500 -977 547
rect -919 581 -819 597
rect -919 547 -903 581
rect -835 547 -819 581
rect -919 500 -819 547
rect -761 581 -661 597
rect -761 547 -745 581
rect -677 547 -661 581
rect -761 500 -661 547
rect -603 581 -503 597
rect -603 547 -587 581
rect -519 547 -503 581
rect -603 500 -503 547
rect -445 581 -345 597
rect -445 547 -429 581
rect -361 547 -345 581
rect -445 500 -345 547
rect -287 581 -187 597
rect -287 547 -271 581
rect -203 547 -187 581
rect -287 500 -187 547
rect -129 581 -29 597
rect -129 547 -113 581
rect -45 547 -29 581
rect -129 500 -29 547
rect 29 581 129 597
rect 29 547 45 581
rect 113 547 129 581
rect 29 500 129 547
rect 187 581 287 597
rect 187 547 203 581
rect 271 547 287 581
rect 187 500 287 547
rect 345 581 445 597
rect 345 547 361 581
rect 429 547 445 581
rect 345 500 445 547
rect 503 581 603 597
rect 503 547 519 581
rect 587 547 603 581
rect 503 500 603 547
rect 661 581 761 597
rect 661 547 677 581
rect 745 547 761 581
rect 661 500 761 547
rect 819 581 919 597
rect 819 547 835 581
rect 903 547 919 581
rect 819 500 919 547
rect 977 581 1077 597
rect 977 547 993 581
rect 1061 547 1077 581
rect 977 500 1077 547
rect 1135 581 1235 597
rect 1135 547 1151 581
rect 1219 547 1235 581
rect 1135 500 1235 547
rect 1293 581 1393 597
rect 1293 547 1309 581
rect 1377 547 1393 581
rect 1293 500 1393 547
rect 1451 581 1551 597
rect 1451 547 1467 581
rect 1535 547 1551 581
rect 1451 500 1551 547
rect 1609 581 1709 597
rect 1609 547 1625 581
rect 1693 547 1709 581
rect 1609 500 1709 547
rect 1767 581 1867 597
rect 1767 547 1783 581
rect 1851 547 1867 581
rect 1767 500 1867 547
rect 1925 581 2025 597
rect 1925 547 1941 581
rect 2009 547 2025 581
rect 1925 500 2025 547
rect 2083 581 2183 597
rect 2083 547 2099 581
rect 2167 547 2183 581
rect 2083 500 2183 547
rect 2241 581 2341 597
rect 2241 547 2257 581
rect 2325 547 2341 581
rect 2241 500 2341 547
rect 2399 581 2499 597
rect 2399 547 2415 581
rect 2483 547 2499 581
rect 2399 500 2499 547
rect 2557 581 2657 597
rect 2557 547 2573 581
rect 2641 547 2657 581
rect 2557 500 2657 547
rect 2715 581 2815 597
rect 2715 547 2731 581
rect 2799 547 2815 581
rect 2715 500 2815 547
rect 2873 581 2973 597
rect 2873 547 2889 581
rect 2957 547 2973 581
rect 2873 500 2973 547
rect 3031 581 3131 597
rect 3031 547 3047 581
rect 3115 547 3131 581
rect 3031 500 3131 547
rect -3131 -547 -3031 -500
rect -3131 -581 -3115 -547
rect -3047 -581 -3031 -547
rect -3131 -597 -3031 -581
rect -2973 -547 -2873 -500
rect -2973 -581 -2957 -547
rect -2889 -581 -2873 -547
rect -2973 -597 -2873 -581
rect -2815 -547 -2715 -500
rect -2815 -581 -2799 -547
rect -2731 -581 -2715 -547
rect -2815 -597 -2715 -581
rect -2657 -547 -2557 -500
rect -2657 -581 -2641 -547
rect -2573 -581 -2557 -547
rect -2657 -597 -2557 -581
rect -2499 -547 -2399 -500
rect -2499 -581 -2483 -547
rect -2415 -581 -2399 -547
rect -2499 -597 -2399 -581
rect -2341 -547 -2241 -500
rect -2341 -581 -2325 -547
rect -2257 -581 -2241 -547
rect -2341 -597 -2241 -581
rect -2183 -547 -2083 -500
rect -2183 -581 -2167 -547
rect -2099 -581 -2083 -547
rect -2183 -597 -2083 -581
rect -2025 -547 -1925 -500
rect -2025 -581 -2009 -547
rect -1941 -581 -1925 -547
rect -2025 -597 -1925 -581
rect -1867 -547 -1767 -500
rect -1867 -581 -1851 -547
rect -1783 -581 -1767 -547
rect -1867 -597 -1767 -581
rect -1709 -547 -1609 -500
rect -1709 -581 -1693 -547
rect -1625 -581 -1609 -547
rect -1709 -597 -1609 -581
rect -1551 -547 -1451 -500
rect -1551 -581 -1535 -547
rect -1467 -581 -1451 -547
rect -1551 -597 -1451 -581
rect -1393 -547 -1293 -500
rect -1393 -581 -1377 -547
rect -1309 -581 -1293 -547
rect -1393 -597 -1293 -581
rect -1235 -547 -1135 -500
rect -1235 -581 -1219 -547
rect -1151 -581 -1135 -547
rect -1235 -597 -1135 -581
rect -1077 -547 -977 -500
rect -1077 -581 -1061 -547
rect -993 -581 -977 -547
rect -1077 -597 -977 -581
rect -919 -547 -819 -500
rect -919 -581 -903 -547
rect -835 -581 -819 -547
rect -919 -597 -819 -581
rect -761 -547 -661 -500
rect -761 -581 -745 -547
rect -677 -581 -661 -547
rect -761 -597 -661 -581
rect -603 -547 -503 -500
rect -603 -581 -587 -547
rect -519 -581 -503 -547
rect -603 -597 -503 -581
rect -445 -547 -345 -500
rect -445 -581 -429 -547
rect -361 -581 -345 -547
rect -445 -597 -345 -581
rect -287 -547 -187 -500
rect -287 -581 -271 -547
rect -203 -581 -187 -547
rect -287 -597 -187 -581
rect -129 -547 -29 -500
rect -129 -581 -113 -547
rect -45 -581 -29 -547
rect -129 -597 -29 -581
rect 29 -547 129 -500
rect 29 -581 45 -547
rect 113 -581 129 -547
rect 29 -597 129 -581
rect 187 -547 287 -500
rect 187 -581 203 -547
rect 271 -581 287 -547
rect 187 -597 287 -581
rect 345 -547 445 -500
rect 345 -581 361 -547
rect 429 -581 445 -547
rect 345 -597 445 -581
rect 503 -547 603 -500
rect 503 -581 519 -547
rect 587 -581 603 -547
rect 503 -597 603 -581
rect 661 -547 761 -500
rect 661 -581 677 -547
rect 745 -581 761 -547
rect 661 -597 761 -581
rect 819 -547 919 -500
rect 819 -581 835 -547
rect 903 -581 919 -547
rect 819 -597 919 -581
rect 977 -547 1077 -500
rect 977 -581 993 -547
rect 1061 -581 1077 -547
rect 977 -597 1077 -581
rect 1135 -547 1235 -500
rect 1135 -581 1151 -547
rect 1219 -581 1235 -547
rect 1135 -597 1235 -581
rect 1293 -547 1393 -500
rect 1293 -581 1309 -547
rect 1377 -581 1393 -547
rect 1293 -597 1393 -581
rect 1451 -547 1551 -500
rect 1451 -581 1467 -547
rect 1535 -581 1551 -547
rect 1451 -597 1551 -581
rect 1609 -547 1709 -500
rect 1609 -581 1625 -547
rect 1693 -581 1709 -547
rect 1609 -597 1709 -581
rect 1767 -547 1867 -500
rect 1767 -581 1783 -547
rect 1851 -581 1867 -547
rect 1767 -597 1867 -581
rect 1925 -547 2025 -500
rect 1925 -581 1941 -547
rect 2009 -581 2025 -547
rect 1925 -597 2025 -581
rect 2083 -547 2183 -500
rect 2083 -581 2099 -547
rect 2167 -581 2183 -547
rect 2083 -597 2183 -581
rect 2241 -547 2341 -500
rect 2241 -581 2257 -547
rect 2325 -581 2341 -547
rect 2241 -597 2341 -581
rect 2399 -547 2499 -500
rect 2399 -581 2415 -547
rect 2483 -581 2499 -547
rect 2399 -597 2499 -581
rect 2557 -547 2657 -500
rect 2557 -581 2573 -547
rect 2641 -581 2657 -547
rect 2557 -597 2657 -581
rect 2715 -547 2815 -500
rect 2715 -581 2731 -547
rect 2799 -581 2815 -547
rect 2715 -597 2815 -581
rect 2873 -547 2973 -500
rect 2873 -581 2889 -547
rect 2957 -581 2973 -547
rect 2873 -597 2973 -581
rect 3031 -547 3131 -500
rect 3031 -581 3047 -547
rect 3115 -581 3131 -547
rect 3031 -597 3131 -581
<< polycont >>
rect -3115 547 -3047 581
rect -2957 547 -2889 581
rect -2799 547 -2731 581
rect -2641 547 -2573 581
rect -2483 547 -2415 581
rect -2325 547 -2257 581
rect -2167 547 -2099 581
rect -2009 547 -1941 581
rect -1851 547 -1783 581
rect -1693 547 -1625 581
rect -1535 547 -1467 581
rect -1377 547 -1309 581
rect -1219 547 -1151 581
rect -1061 547 -993 581
rect -903 547 -835 581
rect -745 547 -677 581
rect -587 547 -519 581
rect -429 547 -361 581
rect -271 547 -203 581
rect -113 547 -45 581
rect 45 547 113 581
rect 203 547 271 581
rect 361 547 429 581
rect 519 547 587 581
rect 677 547 745 581
rect 835 547 903 581
rect 993 547 1061 581
rect 1151 547 1219 581
rect 1309 547 1377 581
rect 1467 547 1535 581
rect 1625 547 1693 581
rect 1783 547 1851 581
rect 1941 547 2009 581
rect 2099 547 2167 581
rect 2257 547 2325 581
rect 2415 547 2483 581
rect 2573 547 2641 581
rect 2731 547 2799 581
rect 2889 547 2957 581
rect 3047 547 3115 581
rect -3115 -581 -3047 -547
rect -2957 -581 -2889 -547
rect -2799 -581 -2731 -547
rect -2641 -581 -2573 -547
rect -2483 -581 -2415 -547
rect -2325 -581 -2257 -547
rect -2167 -581 -2099 -547
rect -2009 -581 -1941 -547
rect -1851 -581 -1783 -547
rect -1693 -581 -1625 -547
rect -1535 -581 -1467 -547
rect -1377 -581 -1309 -547
rect -1219 -581 -1151 -547
rect -1061 -581 -993 -547
rect -903 -581 -835 -547
rect -745 -581 -677 -547
rect -587 -581 -519 -547
rect -429 -581 -361 -547
rect -271 -581 -203 -547
rect -113 -581 -45 -547
rect 45 -581 113 -547
rect 203 -581 271 -547
rect 361 -581 429 -547
rect 519 -581 587 -547
rect 677 -581 745 -547
rect 835 -581 903 -547
rect 993 -581 1061 -547
rect 1151 -581 1219 -547
rect 1309 -581 1377 -547
rect 1467 -581 1535 -547
rect 1625 -581 1693 -547
rect 1783 -581 1851 -547
rect 1941 -581 2009 -547
rect 2099 -581 2167 -547
rect 2257 -581 2325 -547
rect 2415 -581 2483 -547
rect 2573 -581 2641 -547
rect 2731 -581 2799 -547
rect 2889 -581 2957 -547
rect 3047 -581 3115 -547
<< locali >>
rect -3291 649 -3195 683
rect 3195 649 3291 683
rect -3291 587 -3257 649
rect 3257 587 3291 649
rect -3131 547 -3115 581
rect -3047 547 -3031 581
rect -2973 547 -2957 581
rect -2889 547 -2873 581
rect -2815 547 -2799 581
rect -2731 547 -2715 581
rect -2657 547 -2641 581
rect -2573 547 -2557 581
rect -2499 547 -2483 581
rect -2415 547 -2399 581
rect -2341 547 -2325 581
rect -2257 547 -2241 581
rect -2183 547 -2167 581
rect -2099 547 -2083 581
rect -2025 547 -2009 581
rect -1941 547 -1925 581
rect -1867 547 -1851 581
rect -1783 547 -1767 581
rect -1709 547 -1693 581
rect -1625 547 -1609 581
rect -1551 547 -1535 581
rect -1467 547 -1451 581
rect -1393 547 -1377 581
rect -1309 547 -1293 581
rect -1235 547 -1219 581
rect -1151 547 -1135 581
rect -1077 547 -1061 581
rect -993 547 -977 581
rect -919 547 -903 581
rect -835 547 -819 581
rect -761 547 -745 581
rect -677 547 -661 581
rect -603 547 -587 581
rect -519 547 -503 581
rect -445 547 -429 581
rect -361 547 -345 581
rect -287 547 -271 581
rect -203 547 -187 581
rect -129 547 -113 581
rect -45 547 -29 581
rect 29 547 45 581
rect 113 547 129 581
rect 187 547 203 581
rect 271 547 287 581
rect 345 547 361 581
rect 429 547 445 581
rect 503 547 519 581
rect 587 547 603 581
rect 661 547 677 581
rect 745 547 761 581
rect 819 547 835 581
rect 903 547 919 581
rect 977 547 993 581
rect 1061 547 1077 581
rect 1135 547 1151 581
rect 1219 547 1235 581
rect 1293 547 1309 581
rect 1377 547 1393 581
rect 1451 547 1467 581
rect 1535 547 1551 581
rect 1609 547 1625 581
rect 1693 547 1709 581
rect 1767 547 1783 581
rect 1851 547 1867 581
rect 1925 547 1941 581
rect 2009 547 2025 581
rect 2083 547 2099 581
rect 2167 547 2183 581
rect 2241 547 2257 581
rect 2325 547 2341 581
rect 2399 547 2415 581
rect 2483 547 2499 581
rect 2557 547 2573 581
rect 2641 547 2657 581
rect 2715 547 2731 581
rect 2799 547 2815 581
rect 2873 547 2889 581
rect 2957 547 2973 581
rect 3031 547 3047 581
rect 3115 547 3131 581
rect -3177 488 -3143 504
rect -3177 -504 -3143 -488
rect -3019 488 -2985 504
rect -3019 -504 -2985 -488
rect -2861 488 -2827 504
rect -2861 -504 -2827 -488
rect -2703 488 -2669 504
rect -2703 -504 -2669 -488
rect -2545 488 -2511 504
rect -2545 -504 -2511 -488
rect -2387 488 -2353 504
rect -2387 -504 -2353 -488
rect -2229 488 -2195 504
rect -2229 -504 -2195 -488
rect -2071 488 -2037 504
rect -2071 -504 -2037 -488
rect -1913 488 -1879 504
rect -1913 -504 -1879 -488
rect -1755 488 -1721 504
rect -1755 -504 -1721 -488
rect -1597 488 -1563 504
rect -1597 -504 -1563 -488
rect -1439 488 -1405 504
rect -1439 -504 -1405 -488
rect -1281 488 -1247 504
rect -1281 -504 -1247 -488
rect -1123 488 -1089 504
rect -1123 -504 -1089 -488
rect -965 488 -931 504
rect -965 -504 -931 -488
rect -807 488 -773 504
rect -807 -504 -773 -488
rect -649 488 -615 504
rect -649 -504 -615 -488
rect -491 488 -457 504
rect -491 -504 -457 -488
rect -333 488 -299 504
rect -333 -504 -299 -488
rect -175 488 -141 504
rect -175 -504 -141 -488
rect -17 488 17 504
rect -17 -504 17 -488
rect 141 488 175 504
rect 141 -504 175 -488
rect 299 488 333 504
rect 299 -504 333 -488
rect 457 488 491 504
rect 457 -504 491 -488
rect 615 488 649 504
rect 615 -504 649 -488
rect 773 488 807 504
rect 773 -504 807 -488
rect 931 488 965 504
rect 931 -504 965 -488
rect 1089 488 1123 504
rect 1089 -504 1123 -488
rect 1247 488 1281 504
rect 1247 -504 1281 -488
rect 1405 488 1439 504
rect 1405 -504 1439 -488
rect 1563 488 1597 504
rect 1563 -504 1597 -488
rect 1721 488 1755 504
rect 1721 -504 1755 -488
rect 1879 488 1913 504
rect 1879 -504 1913 -488
rect 2037 488 2071 504
rect 2037 -504 2071 -488
rect 2195 488 2229 504
rect 2195 -504 2229 -488
rect 2353 488 2387 504
rect 2353 -504 2387 -488
rect 2511 488 2545 504
rect 2511 -504 2545 -488
rect 2669 488 2703 504
rect 2669 -504 2703 -488
rect 2827 488 2861 504
rect 2827 -504 2861 -488
rect 2985 488 3019 504
rect 2985 -504 3019 -488
rect 3143 488 3177 504
rect 3143 -504 3177 -488
rect -3131 -581 -3115 -547
rect -3047 -581 -3031 -547
rect -2973 -581 -2957 -547
rect -2889 -581 -2873 -547
rect -2815 -581 -2799 -547
rect -2731 -581 -2715 -547
rect -2657 -581 -2641 -547
rect -2573 -581 -2557 -547
rect -2499 -581 -2483 -547
rect -2415 -581 -2399 -547
rect -2341 -581 -2325 -547
rect -2257 -581 -2241 -547
rect -2183 -581 -2167 -547
rect -2099 -581 -2083 -547
rect -2025 -581 -2009 -547
rect -1941 -581 -1925 -547
rect -1867 -581 -1851 -547
rect -1783 -581 -1767 -547
rect -1709 -581 -1693 -547
rect -1625 -581 -1609 -547
rect -1551 -581 -1535 -547
rect -1467 -581 -1451 -547
rect -1393 -581 -1377 -547
rect -1309 -581 -1293 -547
rect -1235 -581 -1219 -547
rect -1151 -581 -1135 -547
rect -1077 -581 -1061 -547
rect -993 -581 -977 -547
rect -919 -581 -903 -547
rect -835 -581 -819 -547
rect -761 -581 -745 -547
rect -677 -581 -661 -547
rect -603 -581 -587 -547
rect -519 -581 -503 -547
rect -445 -581 -429 -547
rect -361 -581 -345 -547
rect -287 -581 -271 -547
rect -203 -581 -187 -547
rect -129 -581 -113 -547
rect -45 -581 -29 -547
rect 29 -581 45 -547
rect 113 -581 129 -547
rect 187 -581 203 -547
rect 271 -581 287 -547
rect 345 -581 361 -547
rect 429 -581 445 -547
rect 503 -581 519 -547
rect 587 -581 603 -547
rect 661 -581 677 -547
rect 745 -581 761 -547
rect 819 -581 835 -547
rect 903 -581 919 -547
rect 977 -581 993 -547
rect 1061 -581 1077 -547
rect 1135 -581 1151 -547
rect 1219 -581 1235 -547
rect 1293 -581 1309 -547
rect 1377 -581 1393 -547
rect 1451 -581 1467 -547
rect 1535 -581 1551 -547
rect 1609 -581 1625 -547
rect 1693 -581 1709 -547
rect 1767 -581 1783 -547
rect 1851 -581 1867 -547
rect 1925 -581 1941 -547
rect 2009 -581 2025 -547
rect 2083 -581 2099 -547
rect 2167 -581 2183 -547
rect 2241 -581 2257 -547
rect 2325 -581 2341 -547
rect 2399 -581 2415 -547
rect 2483 -581 2499 -547
rect 2557 -581 2573 -547
rect 2641 -581 2657 -547
rect 2715 -581 2731 -547
rect 2799 -581 2815 -547
rect 2873 -581 2889 -547
rect 2957 -581 2973 -547
rect 3031 -581 3047 -547
rect 3115 -581 3131 -547
rect -3291 -649 -3257 -587
rect 3257 -649 3291 -587
rect -3291 -683 -3195 -649
rect 3195 -683 3291 -649
<< viali >>
rect -3115 547 -3047 581
rect -2957 547 -2889 581
rect -2799 547 -2731 581
rect -2641 547 -2573 581
rect -2483 547 -2415 581
rect -2325 547 -2257 581
rect -2167 547 -2099 581
rect -2009 547 -1941 581
rect -1851 547 -1783 581
rect -1693 547 -1625 581
rect -1535 547 -1467 581
rect -1377 547 -1309 581
rect -1219 547 -1151 581
rect -1061 547 -993 581
rect -903 547 -835 581
rect -745 547 -677 581
rect -587 547 -519 581
rect -429 547 -361 581
rect -271 547 -203 581
rect -113 547 -45 581
rect 45 547 113 581
rect 203 547 271 581
rect 361 547 429 581
rect 519 547 587 581
rect 677 547 745 581
rect 835 547 903 581
rect 993 547 1061 581
rect 1151 547 1219 581
rect 1309 547 1377 581
rect 1467 547 1535 581
rect 1625 547 1693 581
rect 1783 547 1851 581
rect 1941 547 2009 581
rect 2099 547 2167 581
rect 2257 547 2325 581
rect 2415 547 2483 581
rect 2573 547 2641 581
rect 2731 547 2799 581
rect 2889 547 2957 581
rect 3047 547 3115 581
rect -3177 -488 -3143 488
rect -3019 -488 -2985 488
rect -2861 -488 -2827 488
rect -2703 -488 -2669 488
rect -2545 -488 -2511 488
rect -2387 -488 -2353 488
rect -2229 -488 -2195 488
rect -2071 -488 -2037 488
rect -1913 -488 -1879 488
rect -1755 -488 -1721 488
rect -1597 -488 -1563 488
rect -1439 -488 -1405 488
rect -1281 -488 -1247 488
rect -1123 -488 -1089 488
rect -965 -488 -931 488
rect -807 -488 -773 488
rect -649 -488 -615 488
rect -491 -488 -457 488
rect -333 -488 -299 488
rect -175 -488 -141 488
rect -17 -488 17 488
rect 141 -488 175 488
rect 299 -488 333 488
rect 457 -488 491 488
rect 615 -488 649 488
rect 773 -488 807 488
rect 931 -488 965 488
rect 1089 -488 1123 488
rect 1247 -488 1281 488
rect 1405 -488 1439 488
rect 1563 -488 1597 488
rect 1721 -488 1755 488
rect 1879 -488 1913 488
rect 2037 -488 2071 488
rect 2195 -488 2229 488
rect 2353 -488 2387 488
rect 2511 -488 2545 488
rect 2669 -488 2703 488
rect 2827 -488 2861 488
rect 2985 -488 3019 488
rect 3143 -488 3177 488
rect -3115 -581 -3047 -547
rect -2957 -581 -2889 -547
rect -2799 -581 -2731 -547
rect -2641 -581 -2573 -547
rect -2483 -581 -2415 -547
rect -2325 -581 -2257 -547
rect -2167 -581 -2099 -547
rect -2009 -581 -1941 -547
rect -1851 -581 -1783 -547
rect -1693 -581 -1625 -547
rect -1535 -581 -1467 -547
rect -1377 -581 -1309 -547
rect -1219 -581 -1151 -547
rect -1061 -581 -993 -547
rect -903 -581 -835 -547
rect -745 -581 -677 -547
rect -587 -581 -519 -547
rect -429 -581 -361 -547
rect -271 -581 -203 -547
rect -113 -581 -45 -547
rect 45 -581 113 -547
rect 203 -581 271 -547
rect 361 -581 429 -547
rect 519 -581 587 -547
rect 677 -581 745 -547
rect 835 -581 903 -547
rect 993 -581 1061 -547
rect 1151 -581 1219 -547
rect 1309 -581 1377 -547
rect 1467 -581 1535 -547
rect 1625 -581 1693 -547
rect 1783 -581 1851 -547
rect 1941 -581 2009 -547
rect 2099 -581 2167 -547
rect 2257 -581 2325 -547
rect 2415 -581 2483 -547
rect 2573 -581 2641 -547
rect 2731 -581 2799 -547
rect 2889 -581 2957 -547
rect 3047 -581 3115 -547
<< metal1 >>
rect -3127 581 -3035 587
rect -3127 547 -3115 581
rect -3047 547 -3035 581
rect -3127 541 -3035 547
rect -2969 581 -2877 587
rect -2969 547 -2957 581
rect -2889 547 -2877 581
rect -2969 541 -2877 547
rect -2811 581 -2719 587
rect -2811 547 -2799 581
rect -2731 547 -2719 581
rect -2811 541 -2719 547
rect -2653 581 -2561 587
rect -2653 547 -2641 581
rect -2573 547 -2561 581
rect -2653 541 -2561 547
rect -2495 581 -2403 587
rect -2495 547 -2483 581
rect -2415 547 -2403 581
rect -2495 541 -2403 547
rect -2337 581 -2245 587
rect -2337 547 -2325 581
rect -2257 547 -2245 581
rect -2337 541 -2245 547
rect -2179 581 -2087 587
rect -2179 547 -2167 581
rect -2099 547 -2087 581
rect -2179 541 -2087 547
rect -2021 581 -1929 587
rect -2021 547 -2009 581
rect -1941 547 -1929 581
rect -2021 541 -1929 547
rect -1863 581 -1771 587
rect -1863 547 -1851 581
rect -1783 547 -1771 581
rect -1863 541 -1771 547
rect -1705 581 -1613 587
rect -1705 547 -1693 581
rect -1625 547 -1613 581
rect -1705 541 -1613 547
rect -1547 581 -1455 587
rect -1547 547 -1535 581
rect -1467 547 -1455 581
rect -1547 541 -1455 547
rect -1389 581 -1297 587
rect -1389 547 -1377 581
rect -1309 547 -1297 581
rect -1389 541 -1297 547
rect -1231 581 -1139 587
rect -1231 547 -1219 581
rect -1151 547 -1139 581
rect -1231 541 -1139 547
rect -1073 581 -981 587
rect -1073 547 -1061 581
rect -993 547 -981 581
rect -1073 541 -981 547
rect -915 581 -823 587
rect -915 547 -903 581
rect -835 547 -823 581
rect -915 541 -823 547
rect -757 581 -665 587
rect -757 547 -745 581
rect -677 547 -665 581
rect -757 541 -665 547
rect -599 581 -507 587
rect -599 547 -587 581
rect -519 547 -507 581
rect -599 541 -507 547
rect -441 581 -349 587
rect -441 547 -429 581
rect -361 547 -349 581
rect -441 541 -349 547
rect -283 581 -191 587
rect -283 547 -271 581
rect -203 547 -191 581
rect -283 541 -191 547
rect -125 581 -33 587
rect -125 547 -113 581
rect -45 547 -33 581
rect -125 541 -33 547
rect 33 581 125 587
rect 33 547 45 581
rect 113 547 125 581
rect 33 541 125 547
rect 191 581 283 587
rect 191 547 203 581
rect 271 547 283 581
rect 191 541 283 547
rect 349 581 441 587
rect 349 547 361 581
rect 429 547 441 581
rect 349 541 441 547
rect 507 581 599 587
rect 507 547 519 581
rect 587 547 599 581
rect 507 541 599 547
rect 665 581 757 587
rect 665 547 677 581
rect 745 547 757 581
rect 665 541 757 547
rect 823 581 915 587
rect 823 547 835 581
rect 903 547 915 581
rect 823 541 915 547
rect 981 581 1073 587
rect 981 547 993 581
rect 1061 547 1073 581
rect 981 541 1073 547
rect 1139 581 1231 587
rect 1139 547 1151 581
rect 1219 547 1231 581
rect 1139 541 1231 547
rect 1297 581 1389 587
rect 1297 547 1309 581
rect 1377 547 1389 581
rect 1297 541 1389 547
rect 1455 581 1547 587
rect 1455 547 1467 581
rect 1535 547 1547 581
rect 1455 541 1547 547
rect 1613 581 1705 587
rect 1613 547 1625 581
rect 1693 547 1705 581
rect 1613 541 1705 547
rect 1771 581 1863 587
rect 1771 547 1783 581
rect 1851 547 1863 581
rect 1771 541 1863 547
rect 1929 581 2021 587
rect 1929 547 1941 581
rect 2009 547 2021 581
rect 1929 541 2021 547
rect 2087 581 2179 587
rect 2087 547 2099 581
rect 2167 547 2179 581
rect 2087 541 2179 547
rect 2245 581 2337 587
rect 2245 547 2257 581
rect 2325 547 2337 581
rect 2245 541 2337 547
rect 2403 581 2495 587
rect 2403 547 2415 581
rect 2483 547 2495 581
rect 2403 541 2495 547
rect 2561 581 2653 587
rect 2561 547 2573 581
rect 2641 547 2653 581
rect 2561 541 2653 547
rect 2719 581 2811 587
rect 2719 547 2731 581
rect 2799 547 2811 581
rect 2719 541 2811 547
rect 2877 581 2969 587
rect 2877 547 2889 581
rect 2957 547 2969 581
rect 2877 541 2969 547
rect 3035 581 3127 587
rect 3035 547 3047 581
rect 3115 547 3127 581
rect 3035 541 3127 547
rect -3183 488 -3137 500
rect -3183 -488 -3177 488
rect -3143 -488 -3137 488
rect -3183 -500 -3137 -488
rect -3025 488 -2979 500
rect -3025 -488 -3019 488
rect -2985 -488 -2979 488
rect -3025 -500 -2979 -488
rect -2867 488 -2821 500
rect -2867 -488 -2861 488
rect -2827 -488 -2821 488
rect -2867 -500 -2821 -488
rect -2709 488 -2663 500
rect -2709 -488 -2703 488
rect -2669 -488 -2663 488
rect -2709 -500 -2663 -488
rect -2551 488 -2505 500
rect -2551 -488 -2545 488
rect -2511 -488 -2505 488
rect -2551 -500 -2505 -488
rect -2393 488 -2347 500
rect -2393 -488 -2387 488
rect -2353 -488 -2347 488
rect -2393 -500 -2347 -488
rect -2235 488 -2189 500
rect -2235 -488 -2229 488
rect -2195 -488 -2189 488
rect -2235 -500 -2189 -488
rect -2077 488 -2031 500
rect -2077 -488 -2071 488
rect -2037 -488 -2031 488
rect -2077 -500 -2031 -488
rect -1919 488 -1873 500
rect -1919 -488 -1913 488
rect -1879 -488 -1873 488
rect -1919 -500 -1873 -488
rect -1761 488 -1715 500
rect -1761 -488 -1755 488
rect -1721 -488 -1715 488
rect -1761 -500 -1715 -488
rect -1603 488 -1557 500
rect -1603 -488 -1597 488
rect -1563 -488 -1557 488
rect -1603 -500 -1557 -488
rect -1445 488 -1399 500
rect -1445 -488 -1439 488
rect -1405 -488 -1399 488
rect -1445 -500 -1399 -488
rect -1287 488 -1241 500
rect -1287 -488 -1281 488
rect -1247 -488 -1241 488
rect -1287 -500 -1241 -488
rect -1129 488 -1083 500
rect -1129 -488 -1123 488
rect -1089 -488 -1083 488
rect -1129 -500 -1083 -488
rect -971 488 -925 500
rect -971 -488 -965 488
rect -931 -488 -925 488
rect -971 -500 -925 -488
rect -813 488 -767 500
rect -813 -488 -807 488
rect -773 -488 -767 488
rect -813 -500 -767 -488
rect -655 488 -609 500
rect -655 -488 -649 488
rect -615 -488 -609 488
rect -655 -500 -609 -488
rect -497 488 -451 500
rect -497 -488 -491 488
rect -457 -488 -451 488
rect -497 -500 -451 -488
rect -339 488 -293 500
rect -339 -488 -333 488
rect -299 -488 -293 488
rect -339 -500 -293 -488
rect -181 488 -135 500
rect -181 -488 -175 488
rect -141 -488 -135 488
rect -181 -500 -135 -488
rect -23 488 23 500
rect -23 -488 -17 488
rect 17 -488 23 488
rect -23 -500 23 -488
rect 135 488 181 500
rect 135 -488 141 488
rect 175 -488 181 488
rect 135 -500 181 -488
rect 293 488 339 500
rect 293 -488 299 488
rect 333 -488 339 488
rect 293 -500 339 -488
rect 451 488 497 500
rect 451 -488 457 488
rect 491 -488 497 488
rect 451 -500 497 -488
rect 609 488 655 500
rect 609 -488 615 488
rect 649 -488 655 488
rect 609 -500 655 -488
rect 767 488 813 500
rect 767 -488 773 488
rect 807 -488 813 488
rect 767 -500 813 -488
rect 925 488 971 500
rect 925 -488 931 488
rect 965 -488 971 488
rect 925 -500 971 -488
rect 1083 488 1129 500
rect 1083 -488 1089 488
rect 1123 -488 1129 488
rect 1083 -500 1129 -488
rect 1241 488 1287 500
rect 1241 -488 1247 488
rect 1281 -488 1287 488
rect 1241 -500 1287 -488
rect 1399 488 1445 500
rect 1399 -488 1405 488
rect 1439 -488 1445 488
rect 1399 -500 1445 -488
rect 1557 488 1603 500
rect 1557 -488 1563 488
rect 1597 -488 1603 488
rect 1557 -500 1603 -488
rect 1715 488 1761 500
rect 1715 -488 1721 488
rect 1755 -488 1761 488
rect 1715 -500 1761 -488
rect 1873 488 1919 500
rect 1873 -488 1879 488
rect 1913 -488 1919 488
rect 1873 -500 1919 -488
rect 2031 488 2077 500
rect 2031 -488 2037 488
rect 2071 -488 2077 488
rect 2031 -500 2077 -488
rect 2189 488 2235 500
rect 2189 -488 2195 488
rect 2229 -488 2235 488
rect 2189 -500 2235 -488
rect 2347 488 2393 500
rect 2347 -488 2353 488
rect 2387 -488 2393 488
rect 2347 -500 2393 -488
rect 2505 488 2551 500
rect 2505 -488 2511 488
rect 2545 -488 2551 488
rect 2505 -500 2551 -488
rect 2663 488 2709 500
rect 2663 -488 2669 488
rect 2703 -488 2709 488
rect 2663 -500 2709 -488
rect 2821 488 2867 500
rect 2821 -488 2827 488
rect 2861 -488 2867 488
rect 2821 -500 2867 -488
rect 2979 488 3025 500
rect 2979 -488 2985 488
rect 3019 -488 3025 488
rect 2979 -500 3025 -488
rect 3137 488 3183 500
rect 3137 -488 3143 488
rect 3177 -488 3183 488
rect 3137 -500 3183 -488
rect -3127 -547 -3035 -541
rect -3127 -581 -3115 -547
rect -3047 -581 -3035 -547
rect -3127 -587 -3035 -581
rect -2969 -547 -2877 -541
rect -2969 -581 -2957 -547
rect -2889 -581 -2877 -547
rect -2969 -587 -2877 -581
rect -2811 -547 -2719 -541
rect -2811 -581 -2799 -547
rect -2731 -581 -2719 -547
rect -2811 -587 -2719 -581
rect -2653 -547 -2561 -541
rect -2653 -581 -2641 -547
rect -2573 -581 -2561 -547
rect -2653 -587 -2561 -581
rect -2495 -547 -2403 -541
rect -2495 -581 -2483 -547
rect -2415 -581 -2403 -547
rect -2495 -587 -2403 -581
rect -2337 -547 -2245 -541
rect -2337 -581 -2325 -547
rect -2257 -581 -2245 -547
rect -2337 -587 -2245 -581
rect -2179 -547 -2087 -541
rect -2179 -581 -2167 -547
rect -2099 -581 -2087 -547
rect -2179 -587 -2087 -581
rect -2021 -547 -1929 -541
rect -2021 -581 -2009 -547
rect -1941 -581 -1929 -547
rect -2021 -587 -1929 -581
rect -1863 -547 -1771 -541
rect -1863 -581 -1851 -547
rect -1783 -581 -1771 -547
rect -1863 -587 -1771 -581
rect -1705 -547 -1613 -541
rect -1705 -581 -1693 -547
rect -1625 -581 -1613 -547
rect -1705 -587 -1613 -581
rect -1547 -547 -1455 -541
rect -1547 -581 -1535 -547
rect -1467 -581 -1455 -547
rect -1547 -587 -1455 -581
rect -1389 -547 -1297 -541
rect -1389 -581 -1377 -547
rect -1309 -581 -1297 -547
rect -1389 -587 -1297 -581
rect -1231 -547 -1139 -541
rect -1231 -581 -1219 -547
rect -1151 -581 -1139 -547
rect -1231 -587 -1139 -581
rect -1073 -547 -981 -541
rect -1073 -581 -1061 -547
rect -993 -581 -981 -547
rect -1073 -587 -981 -581
rect -915 -547 -823 -541
rect -915 -581 -903 -547
rect -835 -581 -823 -547
rect -915 -587 -823 -581
rect -757 -547 -665 -541
rect -757 -581 -745 -547
rect -677 -581 -665 -547
rect -757 -587 -665 -581
rect -599 -547 -507 -541
rect -599 -581 -587 -547
rect -519 -581 -507 -547
rect -599 -587 -507 -581
rect -441 -547 -349 -541
rect -441 -581 -429 -547
rect -361 -581 -349 -547
rect -441 -587 -349 -581
rect -283 -547 -191 -541
rect -283 -581 -271 -547
rect -203 -581 -191 -547
rect -283 -587 -191 -581
rect -125 -547 -33 -541
rect -125 -581 -113 -547
rect -45 -581 -33 -547
rect -125 -587 -33 -581
rect 33 -547 125 -541
rect 33 -581 45 -547
rect 113 -581 125 -547
rect 33 -587 125 -581
rect 191 -547 283 -541
rect 191 -581 203 -547
rect 271 -581 283 -547
rect 191 -587 283 -581
rect 349 -547 441 -541
rect 349 -581 361 -547
rect 429 -581 441 -547
rect 349 -587 441 -581
rect 507 -547 599 -541
rect 507 -581 519 -547
rect 587 -581 599 -547
rect 507 -587 599 -581
rect 665 -547 757 -541
rect 665 -581 677 -547
rect 745 -581 757 -547
rect 665 -587 757 -581
rect 823 -547 915 -541
rect 823 -581 835 -547
rect 903 -581 915 -547
rect 823 -587 915 -581
rect 981 -547 1073 -541
rect 981 -581 993 -547
rect 1061 -581 1073 -547
rect 981 -587 1073 -581
rect 1139 -547 1231 -541
rect 1139 -581 1151 -547
rect 1219 -581 1231 -547
rect 1139 -587 1231 -581
rect 1297 -547 1389 -541
rect 1297 -581 1309 -547
rect 1377 -581 1389 -547
rect 1297 -587 1389 -581
rect 1455 -547 1547 -541
rect 1455 -581 1467 -547
rect 1535 -581 1547 -547
rect 1455 -587 1547 -581
rect 1613 -547 1705 -541
rect 1613 -581 1625 -547
rect 1693 -581 1705 -547
rect 1613 -587 1705 -581
rect 1771 -547 1863 -541
rect 1771 -581 1783 -547
rect 1851 -581 1863 -547
rect 1771 -587 1863 -581
rect 1929 -547 2021 -541
rect 1929 -581 1941 -547
rect 2009 -581 2021 -547
rect 1929 -587 2021 -581
rect 2087 -547 2179 -541
rect 2087 -581 2099 -547
rect 2167 -581 2179 -547
rect 2087 -587 2179 -581
rect 2245 -547 2337 -541
rect 2245 -581 2257 -547
rect 2325 -581 2337 -547
rect 2245 -587 2337 -581
rect 2403 -547 2495 -541
rect 2403 -581 2415 -547
rect 2483 -581 2495 -547
rect 2403 -587 2495 -581
rect 2561 -547 2653 -541
rect 2561 -581 2573 -547
rect 2641 -581 2653 -547
rect 2561 -587 2653 -581
rect 2719 -547 2811 -541
rect 2719 -581 2731 -547
rect 2799 -581 2811 -547
rect 2719 -587 2811 -581
rect 2877 -547 2969 -541
rect 2877 -581 2889 -547
rect 2957 -581 2969 -547
rect 2877 -587 2969 -581
rect 3035 -547 3127 -541
rect 3035 -581 3047 -547
rect 3115 -581 3127 -547
rect 3035 -587 3127 -581
<< properties >>
string FIXED_BBOX -3274 -666 3274 666
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 5.0 l 0.5 m 1 nf 40 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
