magic
tech sky130A
magscale 1 2
timestamp 1713199282
<< pwell >>
rect 41058 662788 48258 677598
<< metal1 >>
rect 47100 690276 47400 690400
rect 47100 690224 47224 690276
rect 47276 690224 47400 690276
rect 47100 690010 47400 690224
rect 43870 689830 43950 690010
rect 45350 689990 47400 690010
rect 45350 689938 47224 689990
rect 47276 689938 47400 689990
rect 45350 689926 47400 689938
rect 45350 689874 47224 689926
rect 47276 689874 47400 689926
rect 45350 689862 47400 689874
rect 45350 689830 47224 689862
rect 47100 689810 47224 689830
rect 47276 689810 47400 689862
rect 47100 689576 47400 689810
rect 47100 689524 47224 689576
rect 47276 689524 47400 689576
rect 47100 689400 47400 689524
rect 41900 688676 42200 688800
rect 41900 688624 42024 688676
rect 42076 688624 42200 688676
rect 41900 688490 42200 688624
rect 41900 688438 42024 688490
rect 42076 688438 43870 688490
rect 41900 688426 43870 688438
rect 41900 688374 42024 688426
rect 42076 688374 43870 688426
rect 41900 688362 43870 688374
rect 41900 688310 42024 688362
rect 42076 688310 43870 688362
rect 41900 688176 42200 688310
rect 41900 688124 42024 688176
rect 42076 688124 42200 688176
rect 41900 688000 42200 688124
rect 40920 662800 48300 663400
<< via1 >>
rect 47224 690224 47276 690276
rect 47224 689938 47276 689990
rect 47224 689874 47276 689926
rect 47224 689810 47276 689862
rect 47224 689524 47276 689576
rect 42024 688624 42076 688676
rect 42024 688438 42076 688490
rect 42024 688374 42076 688426
rect 42024 688310 42076 688362
rect 42024 688124 42076 688176
<< metal2 >>
rect 47200 690278 47300 690310
rect 47200 690222 47222 690278
rect 47278 690222 47300 690278
rect 47200 690190 47300 690222
rect 47200 689990 47300 690010
rect 47200 689968 47224 689990
rect 47276 689968 47300 689990
rect 47200 689912 47222 689968
rect 47278 689912 47300 689968
rect 47200 689888 47224 689912
rect 47276 689888 47300 689912
rect 47200 689832 47222 689888
rect 47278 689832 47300 689888
rect 47200 689810 47224 689832
rect 47276 689810 47300 689832
rect 47200 689790 47300 689810
rect 47200 689578 47300 689610
rect 47200 689522 47222 689578
rect 47278 689522 47300 689578
rect 47200 689490 47300 689522
rect 42000 688678 42100 688710
rect 42000 688622 42022 688678
rect 42078 688622 42100 688678
rect 42000 688590 42100 688622
rect 42000 688490 42100 688510
rect 42000 688468 42024 688490
rect 42076 688468 42100 688490
rect 42000 688412 42022 688468
rect 42078 688412 42100 688468
rect 42000 688388 42024 688412
rect 42076 688388 42100 688412
rect 42000 688332 42022 688388
rect 42078 688332 42100 688388
rect 42000 688310 42024 688332
rect 42076 688310 42100 688332
rect 42000 688290 42100 688310
rect 42000 688178 42100 688210
rect 42000 688122 42022 688178
rect 42078 688122 42100 688178
rect 42000 688090 42100 688122
rect 42240 683108 42640 684610
rect 42240 683052 42272 683108
rect 42328 683052 42412 683108
rect 42468 683052 42552 683108
rect 42608 683052 42640 683108
rect 42240 683020 42640 683052
rect 46640 683108 47040 684610
rect 46640 683052 46672 683108
rect 46728 683052 46812 683108
rect 46868 683052 46952 683108
rect 47008 683052 47040 683108
rect 46640 683020 47040 683052
<< via2 >>
rect 47222 690276 47278 690278
rect 47222 690224 47224 690276
rect 47224 690224 47276 690276
rect 47276 690224 47278 690276
rect 47222 690222 47278 690224
rect 47222 689938 47224 689968
rect 47224 689938 47276 689968
rect 47276 689938 47278 689968
rect 47222 689926 47278 689938
rect 47222 689912 47224 689926
rect 47224 689912 47276 689926
rect 47276 689912 47278 689926
rect 47222 689874 47224 689888
rect 47224 689874 47276 689888
rect 47276 689874 47278 689888
rect 47222 689862 47278 689874
rect 47222 689832 47224 689862
rect 47224 689832 47276 689862
rect 47276 689832 47278 689862
rect 47222 689576 47278 689578
rect 47222 689524 47224 689576
rect 47224 689524 47276 689576
rect 47276 689524 47278 689576
rect 47222 689522 47278 689524
rect 42022 688676 42078 688678
rect 42022 688624 42024 688676
rect 42024 688624 42076 688676
rect 42076 688624 42078 688676
rect 42022 688622 42078 688624
rect 42022 688438 42024 688468
rect 42024 688438 42076 688468
rect 42076 688438 42078 688468
rect 42022 688426 42078 688438
rect 42022 688412 42024 688426
rect 42024 688412 42076 688426
rect 42076 688412 42078 688426
rect 42022 688374 42024 688388
rect 42024 688374 42076 688388
rect 42076 688374 42078 688388
rect 42022 688362 42078 688374
rect 42022 688332 42024 688362
rect 42024 688332 42076 688362
rect 42076 688332 42078 688362
rect 42022 688176 42078 688178
rect 42022 688124 42024 688176
rect 42024 688124 42076 688176
rect 42076 688124 42078 688176
rect 42022 688122 42078 688124
rect 42272 683052 42328 683108
rect 42412 683052 42468 683108
rect 42552 683052 42608 683108
rect 46672 683052 46728 683108
rect 46812 683052 46868 683108
rect 46952 683052 47008 683108
<< metal3 >>
rect 46320 691800 56400 692040
rect 46320 691560 52800 691800
rect 46400 691400 52800 691560
rect 46600 691200 52800 691400
rect 53400 691200 54000 691800
rect 54600 691200 55200 691800
rect 55800 691200 56400 691800
rect 46600 691000 56400 691200
rect 47100 690278 57684 690400
rect 47100 690222 47222 690278
rect 47278 690222 57684 690278
rect 47100 689968 57684 690222
rect 47100 689912 47222 689968
rect 47278 689912 57684 689968
rect 47100 689888 57684 689912
rect 47100 689832 47222 689888
rect 47278 689832 57684 689888
rect 47100 689578 57684 689832
rect 47100 689522 47222 689578
rect 47278 689522 57684 689578
rect 47100 689400 57684 689522
rect 29796 688678 42200 688800
rect 29796 688622 42022 688678
rect 42078 688622 42200 688678
rect 29796 688468 42200 688622
rect 29796 688412 42022 688468
rect 42078 688412 42200 688468
rect 29796 688388 42200 688412
rect 29796 688332 42022 688388
rect 42078 688332 42200 688388
rect 29796 688178 42200 688332
rect 29796 688122 42022 688178
rect 42078 688122 42200 688178
rect 29796 687800 42200 688122
rect 29800 687000 47800 687400
rect 29800 686400 42900 687000
rect 42240 683108 43910 683140
rect 42240 683052 42272 683108
rect 42328 683052 42412 683108
rect 42468 683052 42552 683108
rect 42608 683052 43910 683108
rect 42240 683020 43910 683052
rect 45360 683108 47040 683140
rect 45360 683052 46672 683108
rect 46728 683052 46812 683108
rect 46868 683052 46952 683108
rect 47008 683052 47040 683108
rect 45360 683020 47040 683052
rect 45400 682400 56400 682600
rect 45400 681800 52800 682400
rect 53400 681800 54000 682400
rect 54600 681800 55200 682400
rect 55800 681800 56400 682400
rect 45400 681600 56400 681800
<< via3 >>
rect 52800 691200 53400 691800
rect 54000 691200 54600 691800
rect 55200 691200 55800 691800
rect 52800 681800 53400 682400
rect 54000 681800 54600 682400
rect 55200 681800 55800 682400
<< metal4 >>
rect 52400 691800 56400 692000
rect 52400 691200 52800 691800
rect 53400 691200 54000 691800
rect 54600 691200 55200 691800
rect 55800 691200 56400 691800
rect 38670 682003 39330 686050
rect 35200 673800 40000 682003
rect 35200 673000 35600 673800
rect 36400 673000 37200 673800
rect 38000 673000 38800 673800
rect 39600 673000 40000 673800
rect 35200 670600 40000 673000
rect 49920 673968 50580 686100
rect 52400 682400 56400 691200
rect 52400 681800 52800 682400
rect 53400 681800 54000 682400
rect 54600 681800 55200 682400
rect 55800 681800 56400 682400
rect 52400 680000 56400 681800
rect 49920 673732 50132 673968
rect 50368 673732 50580 673968
rect 49920 673568 50580 673732
rect 49920 673332 50132 673568
rect 50368 673332 50580 673568
rect 49920 673168 50580 673332
rect 49920 672932 50132 673168
rect 50368 672932 50580 673168
rect 49920 672700 50580 672932
rect 35200 669800 35600 670600
rect 36400 669800 37200 670600
rect 38000 669800 38800 670600
rect 39600 669800 40000 670600
rect 35200 667200 40000 669800
rect 35200 666400 35600 667200
rect 36400 666400 37200 667200
rect 38000 666400 38800 667200
rect 39600 666400 40000 667200
rect 35200 662800 40000 666400
<< via4 >>
rect 35600 673000 36400 673800
rect 37200 673000 38000 673800
rect 38800 673000 39600 673800
rect 50132 673732 50368 673968
rect 50132 673332 50368 673568
rect 50132 672932 50368 673168
rect 35600 669800 36400 670600
rect 37200 669800 38000 670600
rect 38800 669800 39600 670600
rect 35600 666400 36400 667200
rect 37200 666400 38000 667200
rect 38800 666400 39600 667200
<< metal5 >>
rect 35200 673968 51300 674200
rect 35200 673800 50132 673968
rect 35200 673000 35600 673800
rect 36400 673000 37200 673800
rect 38000 673000 38800 673800
rect 39600 673732 50132 673800
rect 50368 673732 51300 673968
rect 39600 673568 51300 673732
rect 39600 673332 50132 673568
rect 50368 673332 51300 673568
rect 39600 673168 51300 673332
rect 39600 673000 50132 673168
rect 35200 672932 50132 673000
rect 50368 672932 51300 673168
rect 35200 672700 51300 672932
rect 35200 670600 48300 670900
rect 35200 669800 35600 670600
rect 36400 669800 37200 670600
rect 38000 669800 38800 670600
rect 39600 669800 48300 670600
rect 35200 669500 48300 669800
rect 35200 667200 48300 667600
rect 35200 666400 35600 667200
rect 36400 666400 37200 667200
rect 38000 666400 38800 667200
rect 39600 666400 48300 667200
rect 35200 666200 48300 666400
use constant_gm_fingers  constant_gm_fingers_0
timestamp 1713140669
transform 1 0 43810 0 1 682900
box -2700 -20020 4420 1140
use OTA_fingers_031123_NON_FLAT  OTA_fingers_031123_NON_FLAT_0
timestamp 1713196850
transform 1 0 42740 0 1 684710
box -5940 -310 9780 16550
<< labels >>
rlabel metal3 56683 689400 57683 690400 1 VP
port 3 n
rlabel metal3 29800 687800 30800 688800 1 VN
port 2 n
rlabel metal4 35200 662800 40000 665000 1 VSS
port 4 n
rlabel metal3 29800 686400 30800 687400 1 OUT
port 0 n
rlabel metal4 52400 680000 56400 682800 1 VDD
port 1 n
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
