** sch_path: /foss/designs/Analog_FA23_SP24/PriorityEncoder/Priority_Encoder_Testing_v0p0p1.sch
.lib /foss/pdks/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.include /foss/pdks/sky130A/libs.ref/sky130_fd_sc_hd/spice/sky130_fd_sc_hd.spice

.subckt Priority_Encoder_Testing_v0p0p1

V0 IN0 GND pulse 0 1.8 '0.495/ 80E3 ' '0.01/80E3 ' '0.01/80E3 ' '0.49/80E3 ' '1/80E3 '
V1 IN1 GND pulse 0 1.8 '0.495/ 40E3 ' '0.01/40E3 ' '0.01/40E3 ' '0.49/40E3 ' '1/40E3 '
V2 IN2 GND pulse 0 1.8 '0.495/ 20E3 ' '0.01/20E3 ' '0.01/20E3 ' '0.49/20E3 ' '1/20E3 '
V3 IN3 GND pulse 0 1.8 '0.495/ 10E3 ' '0.01/10E3 ' '0.01/10E3 ' '0.49/10E3 ' '1/10E3 '
V4 IN4 GND pulse 0 1.8 '0.495/ 5E3 ' '0.01/5E3 ' '0.01/5E3 ' '0.49/5E3 ' '1/5E3 '
V5 IN5 GND pulse 0 1.8 '0.495/ 2.5E3 ' '0.01/2.5E3 ' '0.01/2.5E3 ' '0.49/2.5E3 ' '1/2.5E3 '
V6 IN6 GND pulse 0 1.8 '0.495/ 1.25E3 ' '0.01/1.25E3 ' '0.01/1.25E3 ' '0.49/1.25E3 ' '1/1.25E3 '
V7 IN7 GND pulse 0 1.8 '0.495/ 0.625E3 ' '0.01/0.625E3 ' '0.01/0.625E3 ' '0.49/0.625E3 ' '1/0.625E3 '
VDD VDD GND 1.8
x1 OUT0 IN0 IN1 IN2 IN3 OUT1 IN4 IN5 IN6 IN7 OUT2 Priority_Encoder_v0p0p1
**** begin user architecture code


.control
save all
tran 1u 2m
write Priority_Encoder_Testing_v0p0p1.raw

.endc


**** end user architecture code
.ends

* expanding   symbol:  /foss/designs/Analog_FA23_SP24/PriorityEncoder/Priority_Encoder_v0p0p1.sym # of pins=11
** sym_path: /foss/designs/Analog_FA23_SP24/PriorityEncoder/Priority_Encoder_v0p0p1.sym
** sch_path: /foss/designs/Analog_FA23_SP24/PriorityEncoder/Priority_Encoder_v0p0p1.sch
.subckt Priority_Encoder_v0p0p1 Q0 D0 D1 D2 D3 Q1 D4 D5 D6 D7 Q2
*.PININFO D2:I D3:I D4:I D5:I D6:I D7:I D1:I D0:I Q0:O Q1:O Q2:O
x0 D1 D3 D5 D7 GND GND VDD VDD Q0 sky130_fd_sc_hd__or4_4
x1 D2 D3 D6 D7 GND GND VDD VDD Q1 sky130_fd_sc_hd__or4_4
x2 D4 D5 D6 D7 GND GND VDD VDD Q2 sky130_fd_sc_hd__or4_4
VDD VDD GND 1.8
* noconn D0
.ends

.GLOBAL GND
.GLOBAL VDD
.end
