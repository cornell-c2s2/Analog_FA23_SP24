* NGSPICE file created from resistorDivider_v0p0p1.ext - technology: sky130A

.subckt sky130_fd_pr__res_xhigh_po_5p73_2GP8TG a_48_11780# a_3774_n8124# a_n4920_11780#
+ a_2532_2096# a_2532_n10168# a_n1194_n6616# a_1290_5648# a_n3678_3604# a_48_12316#
+ a_48_15868# a_n4920_15868# a_n3678_16404# a_n4920_12316# a_n2436_n14792# a_n2436_9736#
+ a_n4920_52# a_1290_n18344# a_n3678_n12212# a_2532_17912# a_3774_10272# a_48_n6616#
+ a_n2436_n16300# a_n4920_n6616# a_1290_n10704# a_n2436_n8124# a_3774_n16836# a_n1194_13824#
+ a_3774_n4572# a_n3678_7692# a_1290_6184# a_n3678_4140# a_n3678_8228# a_3774_52#
+ a_n2436_10272# a_n3678_52# a_1290_3604# a_48_13824# a_n4920_13824# a_1290_n6080#
+ a_n3678_17912# a_1290_n14792# a_n1194_n14256# a_1290_n1992# a_48_1560# a_n2436_n4572#
+ a_1290_n16300# a_3774_11780# a_n3678_n12748# a_n3678_n484# a_n2436_n16836# a_n1194_14360#
+ a_1290_n2528# a_48_5648# a_3774_15868# a_3774_12316# a_3774_2096# a_n1194_n8660#
+ a_1290_7692# a_1290_4140# a_48_14360# a_n4920_14360# a_2532_1560# a_3774_n6616#
+ a_n3678_9736# a_1290_8228# a_2532_n4036# a_n2436_11780# a_48_n8660# a_48_n14256#
+ a_2532_5648# a_n1194_n12212# a_n4920_n8660# a_n4920_n14256# a_48_6184# a_n2436_15868#
+ a_n2436_12316# a_n3678_n18344# a_1290_n8124# a_1290_n484# a_1290_n16836# a_n3678_n10704#
+ a_48_3604# a_n2436_n6616# a_3774_13824# a_n1194_16404# a_n3678_n4036# a_2532_6184#
+ a_3774_n10168# a_1290_10272# a_2532_n14256# a_48_52# a_1290_9736# a_48_16404# a_n4920_16404#
+ a_n3678_n14792# a_n1194_2096# a_2532_3604# a_48_n12212# a_n4920_n12212# a_48_7692#
+ a_1290_n4572# a_n1194_n12748# a_n2436_13824# a_48_4140# a_n3678_n16300# a_3774_14360#
+ a_48_8228# a_2532_52# a_n1194_17912# a_n2436_52# a_3774_1560# a_n4920_2096# a_3774_n8660#
+ a_2532_n6080# a_n2436_n10168# a_2532_n1992# a_2532_7692# a_3774_5648# a_1290_11780#
+ a_2532_4140# a_48_n484# a_2532_n12212# a_n2436_14360# a_2532_n2528# a_48_17912#
+ a_2532_8228# a_n4920_17912# a_1290_12316# a_n1194_n18344# a_1290_15868# a_48_n12748#
+ a_n4920_n12748# a_n1194_n10704# a_n2436_n8660# a_n3678_n16836# a_48_9736# a_1290_n6616#
+ a_n3678_n6080# a_2532_n484# a_n3678_n1992# a_3774_16404# a_3774_6184# a_1290_n10168#
+ a_n3678_n2528# a_3774_3604# a_2532_n8124# a_n1194_n14792# a_2532_n12748# a_2532_9736#
+ a_48_n18344# a_1290_13824# a_n4920_n18344# a_n1194_n16300# a_n1194_1560# a_n2436_16404#
+ a_48_n10704# a_n1194_n4036# a_n4920_n10704# a_n2436_2096# a_n1194_5648# a_2532_10272#
+ a_3774_17912# a_3774_7692# a_3774_4140# a_48_n4036# a_n4920_1560# a_n4920_n4036#
+ a_n3678_n8124# a_2532_n4572# a_3774_8228# a_3774_n14256# a_1290_14360# a_2532_n18344#
+ a_n4920_5648# a_48_n14792# a_n4920_n14792# a_2532_n10704# a_48_n16300# a_n1194_6184#
+ a_n5050_n18474# a_1290_n8660# a_n4920_n16300# a_n1194_n16836# a_n2436_17912# a_n3678_10272#
+ a_3774_n484# a_n1194_3604# a_2532_11780# a_n3678_n4572# a_n4920_6184# a_n3678_n10168#
+ a_2532_15868# a_2532_12316# a_2532_n14792# a_n2436_n14256# a_n1194_52# a_1290_52#
+ a_3774_9736# a_3774_n12212# a_2532_n16300# a_n4920_3604# a_n1194_n6080# a_2532_n6616#
+ a_n3678_2096# a_n1194_n1992# a_1290_16404# a_n1194_7692# a_n1194_4140# a_48_n16836#
+ a_3774_n4036# a_n4920_n16836# a_n3678_11780# a_n1194_n2528# a_n2436_1560# a_n1194_8228#
+ a_48_n6080# a_n3678_15868# a_n3678_12316# a_n4920_n6080# a_48_n1992# a_n2436_5648#
+ a_n4920_n1992# a_n4920_7692# a_n4920_4140# a_1290_n14256# a_2532_13824# a_48_n2528#
+ a_n2436_n12212# a_n4920_n2528# a_n3678_n6616# a_n1194_n484# a_n2436_n4036# a_n4920_8228#
+ a_3774_n12748# a_2532_n16836# a_1290_2096# a_1290_17912# a_n1194_n8124# a_n2436_6184#
+ a_n4920_n484# a_n1194_9736# a_2532_14360# a_n3678_13824# a_n1194_n10168# a_n2436_3604#
+ a_48_n8124# a_n4920_n8124# a_1290_n12212# a_n1194_10272# a_2532_n8660# a_n2436_n12748#
+ a_3774_n18344# a_n4920_9736# a_3774_n10704# a_3774_n6080# a_3774_n1992# a_n1194_n4572#
+ a_n3678_1560# a_48_10272# a_n4920_10272# a_n3678_14360# a_3774_n2528# a_n2436_7692#
+ a_n3678_5648# a_n2436_4140# a_48_n4572# a_48_n10168# a_n2436_8228# a_n4920_n4572#
+ a_n4920_n10168# a_n3678_n8660# a_48_2096# a_n2436_n6080# a_3774_n14792# a_n3678_n14256#
+ a_n2436_n1992# a_n2436_n18344# a_2532_16404# a_1290_n4036# a_n1194_11780# a_1290_n12748#
+ a_n2436_n10704# a_3774_n16300# a_n2436_n2528# a_n1194_12316# a_n1194_15868# a_n2436_n484#
+ a_n3678_6184# a_1290_1560#
X0 a_n4920_9736# a_n4920_8228# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X1 a_n1194_7692# a_n1194_6184# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X2 a_2532_7692# a_2532_6184# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X3 a_n3678_3604# a_n3678_2096# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X4 a_1290_17912# a_1290_16404# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X5 a_n4920_n6616# a_n4920_n8124# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X6 a_3774_9736# a_3774_8228# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X7 a_3774_n12748# a_3774_n14256# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X8 a_n3678_n2528# a_n3678_n4036# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X9 a_n2436_n8660# a_n2436_n10168# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X10 a_n4920_n16836# a_n4920_n18344# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X11 a_48_n10704# a_48_n12212# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X12 a_n1194_n10704# a_n1194_n12212# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X13 a_n2436_15868# a_n2436_14360# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X14 a_n2436_1560# a_n2436_52# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X15 a_3774_n14792# a_3774_n16300# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X16 a_n1194_11780# a_n1194_10272# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X17 a_n3678_n4572# a_n3678_n6080# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X18 a_3774_n6616# a_3774_n8124# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X19 a_n3678_17912# a_n3678_16404# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X20 a_n1194_n484# a_n1194_n1992# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X21 a_1290_n8660# a_1290_n10168# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X22 a_n3678_7692# a_n3678_6184# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X23 a_2532_5648# a_2532_4140# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X24 a_n1194_5648# a_n1194_4140# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X25 a_n1194_13824# a_n1194_12316# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X26 a_48_1560# a_48_52# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X27 a_1290_15868# a_1290_14360# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X28 a_48_n12748# a_48_n14256# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X29 a_n1194_n12748# a_n1194_n14256# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X30 a_3774_n16836# a_3774_n18344# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X31 a_48_11780# a_48_10272# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X32 a_n2436_n6616# a_n2436_n8124# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X33 a_48_n14792# a_48_n16300# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X34 a_n1194_n2528# a_n1194_n4036# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X35 a_48_n484# a_48_n1992# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X36 a_n1194_n14792# a_n1194_n16300# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X37 a_n2436_3604# a_n2436_2096# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X38 a_n2436_n10704# a_n2436_n12212# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X39 a_48_13824# a_48_12316# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X40 a_n3678_n8660# a_n3678_n10168# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X41 a_n3678_15868# a_n3678_14360# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X42 a_n1194_n4572# a_n1194_n6080# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X43 a_2532_11780# a_2532_10272# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X44 a_1290_n6616# a_1290_n8124# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X45 a_n1194_9736# a_n1194_8228# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X46 a_2532_9736# a_2532_8228# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X47 a_n4920_1560# a_n4920_52# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X48 a_1290_3604# a_1290_2096# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X49 a_n3678_5648# a_n3678_4140# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X50 a_n1194_1560# a_n1194_52# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X51 a_n1194_17912# a_n1194_16404# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X52 a_2532_1560# a_2532_52# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X53 a_2532_n484# a_2532_n1992# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X54 a_48_n16836# a_48_n18344# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X55 a_48_n2528# a_48_n4036# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X56 a_2532_13824# a_2532_12316# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X57 a_n1194_n16836# a_n1194_n18344# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X58 a_48_3604# a_48_2096# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X59 a_n2436_n12748# a_n2436_n14256# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X60 a_1290_n10704# a_1290_n12212# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X61 a_48_n4572# a_48_n6080# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X62 a_n2436_7692# a_n2436_6184# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X63 a_n4920_3604# a_n4920_2096# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X64 a_n2436_n14792# a_n2436_n16300# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X65 a_48_17912# a_48_16404# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X66 a_n4920_11780# a_n4920_10272# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X67 a_n3678_n6616# a_n3678_n8124# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X68 a_2532_n2528# a_2532_n4036# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X69 a_n1194_n8660# a_n1194_n10168# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X70 a_n4920_n484# a_n4920_n1992# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X71 a_n3678_9736# a_n3678_8228# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X72 a_1290_7692# a_1290_6184# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X73 a_3774_3604# a_3774_2096# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X74 a_n4920_13824# a_n4920_12316# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X75 a_n1194_15868# a_n1194_14360# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X76 a_2532_n4572# a_2532_n6080# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X77 a_1290_n12748# a_1290_n14256# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X78 a_3774_11780# a_3774_10272# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X79 a_2532_17912# a_2532_16404# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X80 a_48_7692# a_48_6184# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X81 a_n2436_n16836# a_n2436_n18344# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X82 a_3774_n484# a_3774_n1992# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X83 a_n3678_1560# a_n3678_52# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X84 a_n3678_n10704# a_n3678_n12212# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X85 a_1290_n14792# a_1290_n16300# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X86 a_1290_1560# a_1290_52# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X87 a_3774_13824# a_3774_12316# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X88 a_2532_n10704# a_2532_n12212# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X89 a_48_n8660# a_48_n10168# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X90 a_n4920_n2528# a_n4920_n4036# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X91 a_n4920_7692# a_n4920_6184# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X92 a_n2436_5648# a_n2436_4140# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X93 a_48_15868# a_48_14360# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X94 a_n4920_n4572# a_n4920_n6080# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X95 a_n2436_11780# a_n2436_10272# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X96 a_n1194_n6616# a_n1194_n8124# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X97 a_3774_7692# a_3774_6184# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X98 a_1290_5648# a_1290_4140# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X99 a_n4920_17912# a_n4920_16404# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X100 a_3774_n2528# a_3774_n4036# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X101 a_n3678_n12748# a_n3678_n14256# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X102 a_2532_n8660# a_2532_n10168# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X103 a_n2436_n484# a_n2436_n1992# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X104 a_1290_n16836# a_1290_n18344# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X105 a_n2436_13824# a_n2436_12316# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X106 a_2532_n12748# a_2532_n14256# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X107 a_2532_15868# a_2532_14360# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X108 a_48_5648# a_48_4140# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X109 a_1290_11780# a_1290_10272# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X110 a_3774_n4572# a_3774_n6080# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X111 a_n3678_n14792# a_n3678_n16300# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X112 a_3774_17912# a_3774_16404# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X113 a_n4920_n10704# a_n4920_n12212# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X114 a_1290_n484# a_1290_n1992# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X115 a_2532_n14792# a_2532_n16300# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X116 a_48_n6616# a_48_n8124# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X117 a_2532_3604# a_2532_2096# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X118 a_n2436_9736# a_n2436_8228# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X119 a_n1194_3604# a_n1194_2096# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X120 a_n4920_5648# a_n4920_4140# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X121 a_1290_13824# a_1290_12316# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X122 a_n2436_n2528# a_n2436_n4036# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X123 a_3774_1560# a_3774_52# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X124 a_n4920_n8660# a_n4920_n10168# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X125 a_1290_9736# a_1290_8228# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X126 a_3774_5648# a_3774_4140# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X127 a_n4920_15868# a_n4920_14360# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X128 a_n3678_n16836# a_n3678_n18344# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X129 a_n2436_n4572# a_n2436_n6080# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X130 a_2532_n6616# a_2532_n8124# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X131 a_n3678_11780# a_n3678_10272# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X132 a_n4920_n12748# a_n4920_n14256# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X133 a_1290_n2528# a_1290_n4036# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X134 a_n2436_17912# a_n2436_16404# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X135 a_2532_n16836# a_2532_n18344# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X136 a_48_9736# a_48_8228# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X137 a_3774_n10704# a_3774_n12212# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X138 a_n3678_n484# a_n3678_n1992# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X139 a_3774_n8660# a_3774_n10168# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X140 a_n3678_13824# a_n3678_12316# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X141 a_n4920_n14792# a_n4920_n16300# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X142 a_3774_15868# a_3774_14360# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
X143 a_1290_n4572# a_1290_n6080# a_n5050_n18474# sky130_fd_pr__res_xhigh_po_5p73 l=5.38
.ends

.subckt resistorDivider_v0p0p1
XXR1 m1_n4400_25950# m1_n4400_5500# m1_n4400_25950# m1_n4390_15730# m1_n4390_3420#
+ m1_n4400_7540# m1_n4400_19820# m1_n4390_17770# m1_n4400_25950# m1_n4410_30040# m1_n4410_30040#
+ m1_n4410_30040# m1_n4400_25950# m1_n4380_n670# m1_n4400_23900# m1_n4410_13680# m1_n4410_n4170#
+ m1_n4380_1370# m1_n4400_32090# m1_n4400_23900# m1_n4400_7540# m1_n4400_n2690# m1_n4400_7540#
+ m1_n4390_3420# m1_n4400_5500# m1_n4400_n2690# m1_n4400_27990# m1_n4400_9590# m1_n4400_21860#
+ m1_n4400_19820# m1_n4390_17770# m1_n4400_21860# m1_n4410_13680# m1_n4400_23900#
+ m1_n4410_13680# m1_n4390_17770# m1_n4400_27990# m1_n4400_27990# m1_n4400_7540# m1_n4400_32090#
+ m1_n4380_n670# m1_n4380_n670# m1_n4400_11630# m1_n4390_15730# m1_n4400_9590# m1_n4400_n2690#
+ m1_n4400_25950# m1_n4380_1370# m1_n4410_13680# m1_n4400_n2690# m1_n4400_27990# m1_n4400_11630#
+ m1_n4400_19820# m1_n4410_30040# m1_n4400_25950# m1_n4390_15730# m1_n4400_5500# m1_n4400_21860#
+ m1_n4390_17770# m1_n4400_27990# m1_n4400_27990# m1_n4390_15730# m1_n4400_7540# m1_n4400_23900#
+ m1_n4400_21860# m1_n4400_9590# m1_n4400_25950# m1_n4400_5500# m1_n4380_n670# m1_n4400_19820#
+ m1_n4380_1370# m1_n4400_5500# m1_n4380_n670# m1_n4400_19820# m1_n4410_30040# m1_n4400_25950#
+ m1_n4410_n4170# m1_n4400_5500# m1_n4410_13680# m1_n4400_n2690# m1_n4390_3420# m1_n4390_17770#
+ m1_n4400_7540# m1_n4400_27990# m1_n4410_30040# m1_n4400_9590# m1_n4400_19820# m1_n4390_3420#
+ m1_n4400_23900# m1_n4380_n670# m1_n4410_13680# m1_n4400_23900# m1_n4410_30040# m1_n4410_30040#
+ m1_n4380_n670# m1_n4390_15730# m1_n4390_17770# m1_n4380_1370# m1_n4380_1370# m1_n4400_21860#
+ m1_n4400_9590# m1_n4380_1370# m1_n4400_27990# m1_n4390_17770# m1_n4400_n2690# m1_n4400_27990#
+ m1_n4400_21860# m1_n4410_13680# m1_n4400_32090# m1_n4410_13680# m1_n4390_15730#
+ m1_n4390_15730# m1_n4400_5500# m1_n4400_7540# m1_n4390_3420# m1_n4400_11630# m1_n4400_21860#
+ m1_n4400_19820# m1_n4400_25950# m1_n4390_17770# m1_n4410_13680# m1_n4380_1370# m1_n4400_27990#
+ m1_n4400_11630# m1_n4400_32090# m1_n4400_21860# m1_n4400_32090# m1_n4400_25950#
+ m1_n4410_n4170# m1_n4410_30040# m1_n4380_1370# m1_n4380_1370# m1_n4390_3420# m1_n4400_5500#
+ m1_n4400_n2690# m1_n4400_23900# m1_n4400_7540# m1_n4400_7540# m1_n4410_13680# m1_n4400_11630#
+ m1_n4410_30040# m1_n4400_19820# m1_n4390_3420# m1_n4400_11630# m1_n4390_17770# m1_n4400_5500#
+ m1_n4380_n670# m1_n4380_1370# m1_n4400_23900# m1_n4410_n4170# m1_n4400_27990# m1_n4410_n4170#
+ m1_n4400_n2690# m1_n4390_15730# m1_n4410_30040# m1_n4390_3420# m1_n4400_9590# m1_n4390_3420#
+ m1_n4390_15730# m1_n4400_19820# m1_n4400_23900# m1_n4400_32090# m1_n4400_21860#
+ m1_n4390_17770# m1_n4400_9590# m1_n4390_15730# m1_n4400_9590# m1_n4400_5500# m1_n4400_9590#
+ m1_n4400_21860# m1_n4380_n670# m1_n4400_27990# m1_n4410_n4170# m1_n4400_19820# m1_n4380_n670#
+ m1_n4380_n670# m1_n4390_3420# m1_n4400_n2690# m1_n4400_19820# VSUBS m1_n4400_5500#
+ m1_n4400_n2690# m1_n4400_n2690# m1_n4400_32090# m1_n4400_23900# m1_n4410_13680#
+ m1_n4390_17770# m1_n4400_25950# m1_n4400_9590# m1_n4400_19820# m1_n4390_3420# m1_n4410_30040#
+ m1_n4400_25950# m1_n4380_n670# m1_n4380_n670# m1_n4410_13680# m1_n4410_13680# m1_n4400_23900#
+ m1_n4380_1370# m1_n4400_n2690# m1_n4390_17770# m1_n4400_7540# m1_n4400_7540# m1_n4390_15730#
+ m1_n4400_11630# m1_n4410_30040# m1_n4400_21860# m1_n4390_17770# m1_n4400_n2690#
+ m1_n4400_9590# m1_n4400_n2690# m1_n4400_25950# m1_n4400_11630# m1_n4390_15730# m1_n4400_21860#
+ m1_n4400_7540# m1_n4410_30040# m1_n4400_25950# m1_n4400_7540# m1_n4400_11630# m1_n4400_19820#
+ m1_n4400_11630# m1_n4400_21860# m1_n4390_17770# m1_n4380_n670# m1_n4400_27990# m1_n4400_11630#
+ m1_n4380_1370# m1_n4400_11630# m1_n4400_7540# m1_n4410_13680# m1_n4400_9590# m1_n4400_21860#
+ m1_n4380_1370# m1_n4400_n2690# m1_n4390_15730# m1_n4400_32090# m1_n4400_5500# m1_n4400_19820#
+ m1_n4410_13680# m1_n4400_23900# m1_n4400_27990# m1_n4400_27990# m1_n4390_3420# m1_n4390_17770#
+ m1_n4400_5500# m1_n4400_5500# m1_n4380_1370# m1_n4400_23900# m1_n4400_5500# m1_n4380_1370#
+ m1_n4410_n4170# m1_n4400_23900# m1_n4390_3420# m1_n4400_7540# m1_n4400_11630# m1_n4400_9590#
+ m1_n4390_15730# m1_n4400_23900# m1_n4400_23900# m1_n4400_27990# m1_n4400_11630#
+ m1_n4400_21860# m1_n4400_19820# m1_n4390_17770# m1_n4400_9590# m1_n4390_3420# m1_n4400_21860#
+ m1_n4400_9590# m1_n4390_3420# m1_n4400_5500# m1_n4390_15730# m1_n4400_7540# m1_n4380_n670#
+ m1_n4380_n670# m1_n4400_11630# m1_n4410_n4170# m1_n4410_30040# m1_n4400_9590# m1_n4400_25950#
+ m1_n4380_1370# m1_n4390_3420# m1_n4400_n2690# m1_n4400_11630# m1_n4400_25950# m1_n4410_30040#
+ m1_n4410_13680# m1_n4400_19820# m1_n4390_15730# sky130_fd_pr__res_xhigh_po_5p73_2GP8TG
.ends

