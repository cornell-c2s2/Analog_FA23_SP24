magic
tech sky130A
magscale 1 2
timestamp 1708718590
<< checkpaint >>
rect 5726 -978 8838 2962
<< error_s >>
rect 2034 1915 2069 1932
rect 2035 1914 2069 1915
rect 2035 1878 2105 1914
rect 3197 1878 3250 1879
rect 229 1847 287 1853
rect 421 1847 479 1853
rect 613 1847 671 1853
rect 805 1847 863 1853
rect 997 1847 1055 1853
rect 1189 1847 1247 1853
rect 1381 1847 1439 1853
rect 1573 1847 1631 1853
rect 1765 1847 1823 1853
rect 229 1813 241 1847
rect 421 1813 433 1847
rect 613 1813 625 1847
rect 805 1813 817 1847
rect 997 1813 1009 1847
rect 1189 1813 1201 1847
rect 1381 1813 1393 1847
rect 1573 1813 1585 1847
rect 1765 1813 1777 1847
rect 2052 1844 2123 1878
rect 3179 1844 3250 1878
rect 229 1807 287 1813
rect 421 1807 479 1813
rect 613 1807 671 1813
rect 805 1807 863 1813
rect 997 1807 1055 1813
rect 1189 1807 1247 1813
rect 1381 1807 1439 1813
rect 1573 1807 1631 1813
rect 1765 1807 1823 1813
rect 133 719 191 725
rect 325 719 383 725
rect 517 719 575 725
rect 709 719 767 725
rect 901 719 959 725
rect 1093 719 1151 725
rect 1285 719 1343 725
rect 1477 719 1535 725
rect 1669 719 1727 725
rect 1861 719 1919 725
rect 133 685 145 719
rect 325 685 337 719
rect 517 685 529 719
rect 709 685 721 719
rect 901 685 913 719
rect 1093 685 1105 719
rect 1285 685 1297 719
rect 1477 685 1489 719
rect 1669 685 1681 719
rect 1861 685 1873 719
rect 133 679 191 685
rect 325 679 383 685
rect 517 679 575 685
rect 709 679 767 685
rect 901 679 959 685
rect 1093 679 1151 685
rect 1285 679 1343 685
rect 1477 679 1535 685
rect 1669 679 1727 685
rect 1861 679 1919 685
rect 2052 583 2122 1844
rect 3180 1843 3250 1844
rect 3197 1809 3268 1843
rect 5284 1809 5319 1826
rect 2334 1776 2392 1782
rect 2526 1776 2584 1782
rect 2718 1776 2776 1782
rect 2910 1776 2968 1782
rect 2334 1742 2346 1776
rect 2526 1742 2538 1776
rect 2718 1742 2730 1776
rect 2910 1742 2922 1776
rect 2334 1736 2392 1742
rect 2526 1736 2584 1742
rect 2718 1736 2776 1742
rect 2910 1736 2968 1742
rect 2238 666 2296 672
rect 2430 666 2488 672
rect 2622 666 2680 672
rect 2814 666 2872 672
rect 3006 666 3064 672
rect 2238 632 2250 666
rect 2430 632 2442 666
rect 2622 632 2634 666
rect 2814 632 2826 666
rect 3006 632 3018 666
rect 2238 626 2296 632
rect 2430 626 2488 632
rect 2622 626 2680 632
rect 2814 626 2872 632
rect 3006 626 3064 632
rect 2052 547 2105 583
rect 3197 530 3267 1809
rect 5285 1808 5319 1809
rect 5285 1772 5355 1808
rect 6447 1772 6500 1773
rect 3479 1741 3537 1747
rect 3671 1741 3729 1747
rect 3863 1741 3921 1747
rect 4055 1741 4113 1747
rect 4247 1741 4305 1747
rect 4439 1741 4497 1747
rect 4631 1741 4689 1747
rect 4823 1741 4881 1747
rect 5015 1741 5073 1747
rect 3479 1707 3491 1741
rect 3671 1707 3683 1741
rect 3863 1707 3875 1741
rect 4055 1707 4067 1741
rect 4247 1707 4259 1741
rect 4439 1707 4451 1741
rect 4631 1707 4643 1741
rect 4823 1707 4835 1741
rect 5015 1707 5027 1741
rect 5302 1738 5373 1772
rect 6429 1738 6500 1772
rect 3479 1701 3537 1707
rect 3671 1701 3729 1707
rect 3863 1701 3921 1707
rect 4055 1701 4113 1707
rect 4247 1701 4305 1707
rect 4439 1701 4497 1707
rect 4631 1701 4689 1707
rect 4823 1701 4881 1707
rect 5015 1701 5073 1707
rect 3383 613 3441 619
rect 3575 613 3633 619
rect 3767 613 3825 619
rect 3959 613 4017 619
rect 4151 613 4209 619
rect 4343 613 4401 619
rect 4535 613 4593 619
rect 4727 613 4785 619
rect 4919 613 4977 619
rect 5111 613 5169 619
rect 3383 579 3395 613
rect 3575 579 3587 613
rect 3767 579 3779 613
rect 3959 579 3971 613
rect 4151 579 4163 613
rect 4343 579 4355 613
rect 4535 579 4547 613
rect 4727 579 4739 613
rect 4919 579 4931 613
rect 5111 579 5123 613
rect 3383 573 3441 579
rect 3575 573 3633 579
rect 3767 573 3825 579
rect 3959 573 4017 579
rect 4151 573 4209 579
rect 4343 573 4401 579
rect 4535 573 4593 579
rect 4727 573 4785 579
rect 4919 573 4977 579
rect 5111 573 5169 579
rect 3197 494 3250 530
rect 5302 477 5372 1738
rect 6430 1737 6500 1738
rect 6447 1703 6518 1737
rect 5584 1670 5642 1676
rect 5776 1670 5834 1676
rect 5968 1670 6026 1676
rect 6160 1670 6218 1676
rect 5584 1636 5596 1670
rect 5776 1636 5788 1670
rect 5968 1636 5980 1670
rect 6160 1636 6172 1670
rect 5584 1630 5642 1636
rect 5776 1630 5834 1636
rect 5968 1630 6026 1636
rect 6160 1630 6218 1636
rect 5488 560 5546 566
rect 5680 560 5738 566
rect 5872 560 5930 566
rect 6064 560 6122 566
rect 6256 560 6314 566
rect 5488 526 5500 560
rect 5680 526 5692 560
rect 5872 526 5884 560
rect 6064 526 6076 560
rect 6256 526 6268 560
rect 5488 520 5546 526
rect 5680 520 5738 526
rect 5872 520 5930 526
rect 6064 520 6122 526
rect 6256 520 6314 526
rect 5302 441 5355 477
rect 6447 424 6517 1703
rect 6447 388 6500 424
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
rect 0 -1600 200 -1400
rect 0 -2000 200 -1800
use sky130_fd_pr__pfet_01v8_BDZ9JN  XM1
timestamp 0
transform 1 0 1026 0 1 1266
box -1079 -719 1079 719
use sky130_fd_pr__nfet_01v8_KBNS5F  XM2
timestamp 0
transform 1 0 2651 0 1 1204
box -599 -710 599 710
use sky130_fd_pr__pfet_01v8_BDZ9JN  XM3
timestamp 0
transform 1 0 4276 0 1 1160
box -1079 -719 1079 719
use sky130_fd_pr__nfet_01v8_KBNS5F  XM4
timestamp 0
transform 1 0 5901 0 1 1098
box -599 -710 599 710
use sky130_fd_pr__nfet_01v8_MMMA4V  XM5
timestamp 0
transform 1 0 7282 0 1 992
box -296 -710 296 710
use sky130_fd_pr__pfet_01v8_3HZ9VM  XM8
timestamp 0
transform 1 0 6743 0 1 1054
box -296 -719 296 719
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 VREF_P
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 VDD
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 OUT
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 VIN
port 3 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 256 0 0 0 VSS
port 4 nsew
flabel metal1 0 -2000 200 -1800 0 FreeSans 256 0 0 0 VREF_N
port 5 nsew
<< end >>
