magic
tech sky130A
magscale 1 2
timestamp 1717026683
<< metal1 >>
rect 37800 2800 41600 3000
rect 37800 1400 38000 2800
rect 41400 1400 41600 2800
rect 37800 -400 41600 1400
rect 37800 -3600 37900 -400
rect 41500 -3600 41600 -400
rect 42800 2400 46600 2600
rect 42800 1000 43000 2400
rect 46400 1000 46600 2400
rect 42800 0 46600 1000
rect 42800 -1400 43000 0
rect 46400 -1400 46600 0
rect 50700 820 53300 2600
rect 50700 -20 50900 820
rect 53100 -20 53300 820
rect 50700 -100 53300 -20
rect 56720 1020 59220 2600
rect 56720 -40 56880 1020
rect 59080 -40 59220 1020
rect 56720 -100 59220 -40
rect 55300 -600 55800 -500
rect 55300 -1000 55400 -600
rect 55700 -1000 55800 -600
rect 55300 -1300 55800 -1000
rect 42800 -1600 46600 -1400
rect 53300 -1400 53800 -1300
rect 53300 -1600 53400 -1400
rect 53700 -1600 53800 -1400
rect 53300 -1700 53800 -1600
rect 53500 -1860 53800 -1700
rect 37800 -3700 41600 -3600
rect 59600 -4900 60500 -4700
rect 59600 -5200 59700 -4900
rect 60400 -5200 60500 -4900
rect 55500 -5300 56000 -5200
rect 59600 -5300 60500 -5200
rect 55500 -5600 55600 -5300
rect 55900 -5600 56000 -5300
rect 55500 -5700 56000 -5600
rect 55300 -6200 55800 -6100
rect 20800 -6600 22200 -6400
rect 55300 -6500 55400 -6200
rect 55700 -6500 55800 -6200
rect 55300 -6600 55800 -6500
rect 20800 -7400 21000 -6600
rect 22000 -7400 22200 -6600
rect 53500 -6860 53800 -6840
rect 53500 -7120 53520 -6860
rect 53780 -7120 53800 -6860
rect 53500 -7140 53800 -7120
rect 20800 -7600 22200 -7400
rect 59600 -10300 60500 -10100
rect 27000 -10600 34600 -10400
rect 27000 -13000 27200 -10600
rect 34400 -13000 34600 -10600
rect 55400 -10700 56100 -10600
rect 55400 -11100 55500 -10700
rect 56000 -11100 56100 -10700
rect 59600 -10700 59700 -10300
rect 60400 -10700 60500 -10300
rect 59600 -10800 60500 -10700
rect 55400 -11200 56100 -11100
rect 55320 -11660 55800 -11600
rect 55320 -11980 55380 -11660
rect 55740 -11980 55800 -11660
rect 55320 -12040 55800 -11980
rect 53460 -12340 53800 -12320
rect 53460 -12540 53480 -12340
rect 53780 -12540 53800 -12340
rect 53460 -12560 53800 -12540
rect 27000 -13200 34600 -13000
rect 59700 -15600 60400 -15400
rect 59700 -15900 59800 -15600
rect 60300 -15900 60400 -15600
rect 59700 -16000 60400 -15900
rect 55400 -16100 56100 -16000
rect 55400 -16500 55500 -16100
rect 56000 -16500 56100 -16100
rect 55400 -16600 56100 -16500
rect 55300 -17100 55800 -17000
rect 55300 -17400 55400 -17100
rect 55700 -17400 55800 -17100
rect 55300 -17500 55800 -17400
rect 53480 -17740 53800 -17720
rect 53480 -17940 53500 -17740
rect 53780 -17940 53800 -17740
rect 53480 -17960 53800 -17940
rect 59700 -21000 60400 -20800
rect 59700 -21300 59800 -21000
rect 60300 -21300 60400 -21000
rect 59700 -21400 60400 -21300
rect 55400 -21500 56200 -21400
rect 55400 -21900 55500 -21500
rect 56100 -21900 56200 -21500
rect 55400 -22000 56200 -21900
rect 55360 -22480 55800 -22400
rect 55360 -22760 55440 -22480
rect 55720 -22760 55800 -22480
rect 55360 -22840 55800 -22760
rect 53460 -23140 53800 -23120
rect 53460 -23340 53480 -23140
rect 53780 -23340 53800 -23140
rect 53460 -23360 53800 -23340
rect 14400 -26400 20000 -25800
rect 14400 -27200 15000 -26400
rect 10800 -30600 15000 -27200
rect 14400 -31200 15000 -30600
rect 19400 -31200 20000 -26400
rect 26000 -26400 35800 -25800
rect 26000 -30400 26600 -26400
rect 35200 -30400 35800 -26400
rect 59600 -26400 60500 -26200
rect 59600 -26800 59700 -26400
rect 60400 -26800 60500 -26400
rect 55400 -26900 56200 -26800
rect 59600 -26900 60500 -26800
rect 55400 -27300 55500 -26900
rect 56100 -27300 56200 -26900
rect 55400 -27400 56200 -27300
rect 55380 -27880 55800 -27800
rect 55380 -28160 55460 -27880
rect 55720 -28160 55800 -27880
rect 55380 -28240 55800 -28160
rect 53460 -28540 53800 -28520
rect 53460 -28740 53480 -28540
rect 53780 -28740 53800 -28540
rect 53460 -28760 53800 -28740
rect 26000 -31000 35800 -30400
rect 14400 -31800 20000 -31200
rect 59700 -31800 60400 -31600
rect 36000 -32200 37000 -32000
rect 59700 -32100 59800 -31800
rect 60300 -32100 60400 -31800
rect 59700 -32200 60400 -32100
rect 36000 -33000 36200 -32200
rect 36800 -33000 37000 -32200
rect 55400 -32300 56200 -32200
rect 55400 -32700 55500 -32300
rect 56100 -32700 56200 -32300
rect 55400 -32800 56200 -32700
rect 14000 -38000 25000 -33000
rect 36000 -33200 37000 -33000
rect 55380 -33280 55800 -33200
rect 55380 -33560 55460 -33280
rect 55720 -33560 55800 -33280
rect 35900 -33700 38200 -33600
rect 55380 -33640 55800 -33560
rect 35900 -34700 36000 -33700
rect 38100 -34700 38200 -33700
rect 53460 -33940 53800 -33920
rect 53460 -34140 53480 -33940
rect 53780 -34140 53800 -33940
rect 53460 -34160 53800 -34140
rect 71900 -34100 74100 -34000
rect 35900 -34800 38200 -34700
rect 35900 -35300 39100 -35200
rect 35900 -36300 36000 -35300
rect 39000 -36300 39100 -35300
rect 71900 -35500 72000 -34100
rect 74000 -35500 74100 -34100
rect 71900 -35600 74100 -35500
rect 35900 -36400 39100 -36300
rect 35900 -36900 40100 -36800
rect 35900 -37900 36000 -36900
rect 40000 -37900 40100 -36900
rect 59800 -37200 60300 -37000
rect 59800 -37400 59900 -37200
rect 60200 -37400 60300 -37200
rect 59800 -37500 60300 -37400
rect 35900 -38000 40100 -37900
rect 55300 -37700 56200 -37600
rect 14000 -49000 15000 -38000
rect 24000 -49000 25000 -38000
rect 55300 -38100 55400 -37700
rect 56100 -38100 56200 -37700
rect 55300 -38200 56200 -38100
rect 35900 -38500 41100 -38400
rect 35900 -39500 36000 -38500
rect 41000 -39500 41100 -38500
rect 55380 -38680 55800 -38600
rect 55380 -38960 55460 -38680
rect 55720 -38960 55800 -38680
rect 55380 -39040 55800 -38960
rect 35900 -39600 41100 -39500
rect 53460 -39340 53800 -39320
rect 53460 -39540 53480 -39340
rect 53780 -39540 53800 -39340
rect 53460 -39560 53800 -39540
rect 35900 -40100 42200 -40000
rect 35900 -41100 36000 -40100
rect 42100 -41100 42200 -40100
rect 92000 -40800 95800 -38600
rect 35900 -41200 42200 -41100
rect 35900 -41700 43200 -41600
rect 35900 -42700 36000 -41700
rect 43100 -42700 43200 -41700
rect 35900 -42800 43200 -42700
rect 59600 -42800 60600 -42400
rect 43100 -43200 44400 -43000
rect 35900 -43300 44400 -43200
rect 35900 -44300 36000 -43300
rect 44300 -44300 44400 -43300
rect 55400 -43100 56200 -43000
rect 55400 -43500 55500 -43100
rect 56100 -43500 56200 -43100
rect 55400 -43600 56200 -43500
rect 59600 -43400 59800 -42800
rect 60400 -43400 60600 -42800
rect 59600 -43600 60600 -43400
rect 35900 -44400 44400 -44300
rect 55420 -44080 55800 -44000
rect 55420 -44360 55500 -44080
rect 55720 -44360 55800 -44080
rect 55420 -44440 55800 -44360
rect 53460 -44740 53800 -44720
rect 35900 -44900 44400 -44800
rect 35900 -45900 36000 -44900
rect 44300 -45900 44400 -44900
rect 53460 -44940 53480 -44740
rect 53780 -44940 53800 -44740
rect 53460 -44960 53800 -44940
rect 92000 -45400 95800 -43200
rect 35900 -46000 44400 -45900
rect 35900 -46500 43500 -46400
rect 35900 -47500 36000 -46500
rect 43400 -47500 43500 -46500
rect 35900 -47600 43500 -47500
rect 14000 -55000 25000 -49000
rect 35900 -48100 42600 -48000
rect 35900 -49100 36000 -48100
rect 42500 -49100 42600 -48100
rect 55400 -48500 56200 -48400
rect 59600 -48500 60500 -47900
rect 55400 -48900 55500 -48500
rect 56100 -48900 56200 -48500
rect 55400 -49000 56200 -48900
rect 35900 -49200 42600 -49100
rect 92000 -49400 95800 -47200
rect 55380 -49480 55800 -49400
rect 35900 -49700 41700 -49600
rect 35900 -50700 36000 -49700
rect 41600 -50700 41700 -49700
rect 55380 -49760 55460 -49480
rect 55720 -49760 55800 -49480
rect 55380 -49840 55800 -49760
rect 53440 -50140 53800 -50120
rect 53440 -50340 53460 -50140
rect 53780 -50340 53800 -50140
rect 53440 -50360 53800 -50340
rect 35900 -50800 41700 -50700
rect 35900 -51300 40800 -51200
rect 35900 -52300 36000 -51300
rect 40700 -52300 40800 -51300
rect 35900 -52400 40800 -52300
rect 35900 -52900 39900 -52800
rect 35900 -53900 36000 -52900
rect 39800 -53900 39900 -52900
rect 92000 -53200 95800 -51000
rect 35900 -54000 39900 -53900
rect 55300 -53900 56200 -53800
rect 59600 -53900 60500 -53300
rect 55300 -54300 55400 -53900
rect 56100 -54300 56200 -53900
rect 55300 -54400 56200 -54300
rect 35900 -54500 38900 -54400
rect 35900 -55500 36000 -54500
rect 38800 -55500 38900 -54500
rect 55380 -54880 55800 -54800
rect 55380 -55160 55460 -54880
rect 55720 -55160 55800 -54880
rect 55380 -55240 55800 -55160
rect 35900 -55600 38900 -55500
rect 53460 -55540 53800 -55520
rect 53460 -55740 53480 -55540
rect 53780 -55740 53800 -55540
rect 53460 -55760 53800 -55740
rect 35900 -56100 37800 -56000
rect 35900 -57100 36000 -56100
rect 37700 -57100 37800 -56100
rect 35900 -57200 37800 -57100
rect 24400 -58800 36000 -58200
rect 14600 -60000 20200 -59400
rect 14600 -60800 15200 -60000
rect 10600 -64200 15200 -60800
rect 14600 -64800 15200 -64200
rect 19600 -64800 20200 -60000
rect 14600 -65400 20200 -64800
rect 24400 -64800 25000 -58800
rect 35400 -64800 36000 -58800
rect 55400 -59300 56200 -59200
rect 59600 -59300 60500 -58700
rect 55400 -59700 55500 -59300
rect 56100 -59700 56200 -59300
rect 55400 -59800 56200 -59700
rect 55380 -60280 55800 -60200
rect 55380 -60560 55460 -60280
rect 55720 -60560 55800 -60280
rect 55380 -60640 55800 -60560
rect 53460 -60940 53800 -60920
rect 53460 -61140 53480 -60940
rect 53780 -61140 53800 -60940
rect 53460 -61160 53800 -61140
rect 24400 -65400 36000 -64800
rect 55400 -64700 56200 -64600
rect 59600 -64700 60500 -64100
rect 55400 -65100 55500 -64700
rect 56100 -65100 56200 -64700
rect 55400 -65200 56200 -65100
rect 55360 -65680 55800 -65600
rect 55360 -65960 55440 -65680
rect 55720 -65960 55800 -65680
rect 55360 -66040 55800 -65960
rect 53460 -66340 53800 -66320
rect 53460 -66540 53480 -66340
rect 53780 -66540 53800 -66340
rect 53460 -66560 53800 -66540
rect 55400 -70100 56200 -70000
rect 59600 -70100 60500 -69500
rect 55400 -70500 55500 -70100
rect 56100 -70500 56200 -70100
rect 55400 -70600 56200 -70500
rect 55380 -71080 55800 -71000
rect 55380 -71360 55460 -71080
rect 55720 -71360 55800 -71080
rect 55380 -71440 55800 -71360
rect 53460 -71740 53800 -71720
rect 53460 -71940 53480 -71740
rect 53780 -71940 53800 -71740
rect 53460 -71960 53800 -71940
rect 55400 -75500 56200 -75400
rect 59600 -75500 60500 -74900
rect 55400 -75900 55500 -75500
rect 56100 -75900 56200 -75500
rect 55400 -76000 56200 -75900
rect 55320 -76480 55800 -76400
rect 55320 -76760 55400 -76480
rect 55720 -76760 55800 -76480
rect 55320 -76840 55800 -76760
rect 53460 -77140 53800 -77120
rect 53460 -77340 53480 -77140
rect 53780 -77340 53800 -77140
rect 53460 -77360 53800 -77340
rect 56580 -77892 57066 -77610
rect 56362 -79722 57006 -79558
rect 55400 -80900 56300 -80800
rect 59600 -80900 60500 -80300
rect 55400 -81300 55500 -80900
rect 56200 -81300 56300 -80900
rect 55400 -81400 56300 -81300
rect 55360 -81880 55800 -81800
rect 55360 -82160 55440 -81880
rect 55720 -82160 55800 -81880
rect 55360 -82240 55800 -82160
rect 53460 -82540 53800 -82520
rect 53460 -82740 53480 -82540
rect 53780 -82740 53800 -82540
rect 53460 -82760 53800 -82740
rect 56592 -83034 57024 -83024
rect 56584 -83258 57024 -83034
rect 56584 -83268 57016 -83258
rect 56374 -85082 57010 -84958
rect 55400 -86300 56200 -86200
rect 59600 -86300 60500 -85700
rect 55400 -86600 55500 -86300
rect 56100 -86600 56200 -86300
rect 55400 -86700 56200 -86600
<< via1 >>
rect 38000 1400 41400 2800
rect 37900 -3600 41500 -400
rect 43000 1000 46400 2400
rect 43000 -1400 46400 0
rect 50900 -20 53100 820
rect 56880 -40 59080 1020
rect 55400 -1000 55700 -600
rect 53400 -1600 53700 -1400
rect 59700 -5200 60400 -4900
rect 55600 -5600 55900 -5300
rect 55400 -6500 55700 -6200
rect 21000 -7400 22000 -6600
rect 53520 -7120 53780 -6860
rect 27200 -13000 34400 -10600
rect 55500 -11100 56000 -10700
rect 59700 -10700 60400 -10300
rect 55380 -11980 55740 -11660
rect 53480 -12540 53780 -12340
rect 59800 -15900 60300 -15600
rect 55500 -16500 56000 -16100
rect 55400 -17400 55700 -17100
rect 53500 -17940 53780 -17740
rect 59800 -21300 60300 -21000
rect 55500 -21900 56100 -21500
rect 55440 -22760 55720 -22480
rect 53480 -23340 53780 -23140
rect 15000 -31200 19400 -26400
rect 26600 -30400 35200 -26400
rect 59700 -26800 60400 -26400
rect 55500 -27300 56100 -26900
rect 55460 -28160 55720 -27880
rect 53480 -28740 53780 -28540
rect 59800 -32100 60300 -31800
rect 36200 -33000 36800 -32200
rect 55500 -32700 56100 -32300
rect 55460 -33560 55720 -33280
rect 36000 -34700 38100 -33700
rect 53480 -34140 53780 -33940
rect 36000 -36300 39000 -35300
rect 72000 -35500 74000 -34100
rect 36000 -37900 40000 -36900
rect 59900 -37400 60200 -37200
rect 15000 -49000 24000 -38000
rect 55400 -38100 56100 -37700
rect 36000 -39500 41000 -38500
rect 55460 -38960 55720 -38680
rect 53480 -39540 53780 -39340
rect 36000 -41100 42100 -40100
rect 36000 -42700 43100 -41700
rect 36000 -44300 44300 -43300
rect 55500 -43500 56100 -43100
rect 59800 -43400 60400 -42800
rect 55500 -44360 55720 -44080
rect 36000 -45900 44300 -44900
rect 53480 -44940 53780 -44740
rect 36000 -47500 43400 -46500
rect 36000 -49100 42500 -48100
rect 55500 -48900 56100 -48500
rect 36000 -50700 41600 -49700
rect 55460 -49760 55720 -49480
rect 53460 -50340 53780 -50140
rect 36000 -52300 40700 -51300
rect 36000 -53900 39800 -52900
rect 55400 -54300 56100 -53900
rect 36000 -55500 38800 -54500
rect 55460 -55160 55720 -54880
rect 53480 -55740 53780 -55540
rect 36000 -57100 37700 -56100
rect 15200 -64800 19600 -60000
rect 25000 -64800 35400 -58800
rect 55500 -59700 56100 -59300
rect 55460 -60560 55720 -60280
rect 53480 -61140 53780 -60940
rect 55500 -65100 56100 -64700
rect 55440 -65960 55720 -65680
rect 53480 -66540 53780 -66340
rect 55500 -70500 56100 -70100
rect 55460 -71360 55720 -71080
rect 53480 -71940 53780 -71740
rect 55500 -75900 56100 -75500
rect 55400 -76760 55720 -76480
rect 53480 -77340 53780 -77140
rect 55500 -81300 56200 -80900
rect 55440 -82160 55720 -81880
rect 53480 -82740 53780 -82540
rect 55500 -86600 56100 -86300
<< metal2 >>
rect 37800 2800 41600 3000
rect 37800 1400 38000 2800
rect 41400 1400 41600 2800
rect 37800 1200 41600 1400
rect 42800 2400 46600 2600
rect 42800 1000 43000 2400
rect 46400 1000 46600 2400
rect 42800 800 46600 1000
rect 56880 1020 59080 1030
rect 50800 820 53200 900
rect 42800 0 46600 200
rect 37800 -400 41600 -300
rect 37800 -3600 37900 -400
rect 41500 -3600 41600 -400
rect 42800 -1400 43000 0
rect 46400 -1400 46600 0
rect 50800 -20 50900 820
rect 53100 -20 53200 820
rect 50800 -100 53200 -20
rect 56880 -50 59080 -40
rect 51400 -800 52600 -100
rect 51400 -1000 51500 -800
rect 52500 -1000 52600 -800
rect 42800 -1600 46600 -1400
rect 47000 -1300 48100 -1100
rect 37800 -3700 41600 -3600
rect 47000 -1700 47700 -1300
rect 48000 -1700 48100 -1300
rect 36200 -5000 37200 -4800
rect 36200 -5800 36400 -5000
rect 37000 -5800 37200 -5000
rect 47000 -5300 48100 -1700
rect 20800 -6600 22200 -6400
rect 20800 -7400 21000 -6600
rect 22000 -7400 22200 -6600
rect 20800 -7600 22200 -7400
rect 24600 -8700 25800 -8600
rect 24600 -9400 24700 -8700
rect 25700 -9400 25800 -8700
rect 24600 -11800 25800 -9400
rect 27000 -10600 34600 -10400
rect 27000 -13000 27200 -10600
rect 34400 -13000 34600 -10600
rect 27000 -13200 34600 -13000
rect 14400 -26400 20000 -25800
rect 14400 -31200 15000 -26400
rect 19400 -31200 20000 -26400
rect 26000 -26400 35600 -25800
rect 26000 -30400 26600 -26400
rect 35200 -30400 35600 -26400
rect 26000 -31000 35600 -30400
rect 14400 -31800 20000 -31200
rect 36200 -32000 37200 -5800
rect 46400 -6780 48100 -5300
rect 46400 -7200 47640 -6780
rect 48080 -7200 48100 -6780
rect 46400 -8700 48100 -7200
rect 46400 -9400 46700 -8700
rect 47800 -9400 48100 -8700
rect 36000 -32200 37200 -32000
rect 36000 -33000 36200 -32200
rect 36800 -33000 37200 -32200
rect 36000 -33200 37200 -33000
rect 37500 -10700 38200 -10600
rect 37500 -11100 37600 -10700
rect 38100 -11100 38200 -10700
rect 37500 -33600 38200 -11100
rect 46400 -12220 48100 -9400
rect 46400 -12640 47700 -12220
rect 48080 -12640 48100 -12220
rect 35900 -33700 38200 -33600
rect 35900 -34700 36000 -33700
rect 38100 -34700 38200 -33700
rect 35900 -34800 38200 -34700
rect 38400 -16000 39100 -15900
rect 38400 -16600 38500 -16000
rect 39000 -16600 39100 -16000
rect 38400 -35200 39100 -16600
rect 46400 -17620 48100 -12640
rect 46400 -18100 47640 -17620
rect 48080 -18100 48100 -17620
rect 35900 -35300 39100 -35200
rect 35900 -36300 36000 -35300
rect 39000 -36300 39100 -35300
rect 35900 -36400 39100 -36300
rect 39400 -21400 40100 -21300
rect 39400 -22000 39500 -21400
rect 40000 -22000 40100 -21400
rect 39400 -36800 40100 -22000
rect 46400 -23020 48100 -18100
rect 46400 -23440 47680 -23020
rect 48080 -23440 48100 -23020
rect 35900 -36900 40100 -36800
rect 14000 -38000 25000 -37000
rect 35900 -37900 36000 -36900
rect 40000 -37900 40100 -36900
rect 35900 -38000 40100 -37900
rect 40300 -26800 41100 -26700
rect 40300 -27400 40400 -26800
rect 41000 -27400 41100 -26800
rect 14000 -49000 15000 -38000
rect 24000 -49000 25000 -38000
rect 40300 -38400 41100 -27400
rect 46400 -28460 48100 -23440
rect 46400 -28840 47800 -28460
rect 48080 -28840 48100 -28460
rect 35900 -38500 41100 -38400
rect 35900 -39500 36000 -38500
rect 41000 -39500 41100 -38500
rect 35900 -39600 41100 -39500
rect 41400 -32200 42200 -32100
rect 41400 -32800 41500 -32200
rect 42100 -32800 42200 -32200
rect 41400 -40000 42200 -32800
rect 46400 -33860 48100 -28840
rect 46400 -34200 47760 -33860
rect 48080 -34200 48100 -33860
rect 35900 -40100 42200 -40000
rect 35900 -41100 36000 -40100
rect 42100 -41100 42200 -40100
rect 35900 -41200 42200 -41100
rect 42400 -37600 43200 -37500
rect 42400 -38200 42500 -37600
rect 43100 -38200 43200 -37600
rect 42400 -41600 43200 -38200
rect 35900 -41700 43200 -41600
rect 35900 -42700 36000 -41700
rect 43100 -42700 43200 -41700
rect 35900 -42800 43200 -42700
rect 46400 -39220 48100 -34200
rect 46400 -39640 47760 -39220
rect 48080 -39640 48100 -39220
rect 43100 -43100 44400 -43000
rect 43100 -43200 43200 -43100
rect 35900 -43300 43200 -43200
rect 35900 -44300 36000 -43300
rect 44300 -44300 44400 -43100
rect 35900 -44400 44400 -44300
rect 46400 -44640 48100 -39640
rect 35900 -44900 44400 -44800
rect 35900 -45900 36000 -44900
rect 44300 -45900 44400 -44900
rect 35900 -46000 44400 -45900
rect 35900 -46500 43500 -46400
rect 35900 -47500 36000 -46500
rect 43400 -47500 43500 -46500
rect 35900 -47600 43500 -47500
rect 14000 -50000 25000 -49000
rect 35900 -48100 42600 -48000
rect 35900 -49100 36000 -48100
rect 42500 -49100 42600 -48100
rect 35900 -49200 42600 -49100
rect 35900 -49700 41700 -49600
rect 35900 -50700 36000 -49700
rect 41600 -50700 41700 -49700
rect 35900 -50800 41700 -50700
rect 35900 -51300 40800 -51200
rect 35900 -52300 36000 -51300
rect 40700 -52300 40800 -51300
rect 35900 -52400 40800 -52300
rect 35900 -52900 39900 -52800
rect 35900 -53900 36000 -52900
rect 39800 -53900 39900 -52900
rect 35900 -54000 39900 -53900
rect 35900 -54500 38900 -54400
rect 35900 -55500 36000 -54500
rect 38800 -55500 38900 -54500
rect 35900 -55600 38900 -55500
rect 35900 -56100 37800 -56000
rect 35900 -57100 36000 -56100
rect 37700 -57100 37800 -56100
rect 35900 -57200 37800 -57100
rect 24400 -58800 36000 -58200
rect 14600 -60000 20200 -59400
rect 14600 -64800 15200 -60000
rect 19600 -64800 20200 -60000
rect 14600 -65400 20200 -64800
rect 24400 -64800 25000 -58800
rect 35400 -64800 36000 -58800
rect 24400 -65400 36000 -64800
rect 37100 -86200 37800 -57200
rect 38200 -80800 38900 -55600
rect 39200 -75400 39900 -54000
rect 40100 -70000 40800 -52400
rect 41000 -64600 41700 -50800
rect 41900 -59200 42600 -49200
rect 42800 -53800 43500 -47600
rect 43700 -48400 44400 -46000
rect 43700 -49000 43800 -48400
rect 44300 -49000 44400 -48400
rect 43700 -49100 44400 -49000
rect 46400 -45060 47820 -44640
rect 48080 -45060 48100 -44640
rect 42800 -54400 42900 -53800
rect 43400 -54400 43500 -53800
rect 42800 -54500 43500 -54400
rect 46400 -49980 48100 -45060
rect 46400 -50480 47740 -49980
rect 48080 -50480 48100 -49980
rect 41900 -59800 42000 -59200
rect 42500 -59800 42600 -59200
rect 41900 -59900 42600 -59800
rect 46400 -55460 48100 -50480
rect 46400 -55820 47820 -55460
rect 48080 -55820 48100 -55460
rect 41000 -65200 41100 -64600
rect 41600 -65200 41700 -64600
rect 41000 -65300 41700 -65200
rect 46400 -60760 48100 -55820
rect 46400 -61300 47680 -60760
rect 48080 -61300 48100 -60760
rect 40100 -70600 40200 -70000
rect 40700 -70600 40800 -70000
rect 40100 -70700 40800 -70600
rect 46400 -66220 48100 -61300
rect 46400 -66660 47860 -66220
rect 48080 -66660 48100 -66220
rect 39200 -76000 39300 -75400
rect 39800 -76000 39900 -75400
rect 39200 -76100 39900 -76000
rect 46400 -71600 48100 -66660
rect 46400 -72060 47720 -71600
rect 48080 -72060 48100 -71600
rect 38200 -81400 38300 -80800
rect 38800 -81400 38900 -80800
rect 38200 -81500 38900 -81400
rect 46400 -76940 48100 -72060
rect 46400 -77500 47780 -76940
rect 48080 -77500 48100 -76940
rect 46400 -82380 48100 -77500
rect 46400 -82860 47800 -82380
rect 48080 -82860 48100 -82380
rect 46400 -82960 48100 -82860
rect 51400 -6300 52600 -1000
rect 55300 -600 55800 -500
rect 55300 -1000 55400 -600
rect 55700 -1000 55800 -600
rect 55300 -1100 55800 -1000
rect 53300 -1400 53800 -1300
rect 53300 -1600 53400 -1400
rect 53700 -1600 53800 -1400
rect 53300 -1700 53800 -1600
rect 57800 -3020 58240 -3010
rect 56900 -3140 57800 -3020
rect 57800 -3150 58240 -3140
rect 59600 -4900 60500 -4800
rect 59600 -5200 59700 -4900
rect 60400 -5200 60500 -4900
rect 55500 -5300 56000 -5200
rect 59600 -5300 60500 -5200
rect 68000 -4900 68700 -4800
rect 68000 -5200 68100 -4900
rect 68600 -5200 68700 -4900
rect 55500 -5600 55600 -5300
rect 55900 -5600 56000 -5300
rect 55500 -5700 56000 -5600
rect 51400 -6500 51500 -6300
rect 52500 -6500 52600 -6300
rect 51400 -11700 52600 -6500
rect 55300 -6200 55800 -6100
rect 55300 -6500 55400 -6200
rect 55700 -6500 55800 -6200
rect 55300 -6600 55800 -6500
rect 53500 -6860 53800 -6840
rect 53500 -7120 53520 -6860
rect 53780 -7120 53800 -6860
rect 53500 -7140 53800 -7120
rect 57800 -8420 58240 -8410
rect 56900 -8540 57800 -8420
rect 57800 -8550 58240 -8540
rect 59600 -10300 60500 -10200
rect 55400 -10700 56100 -10600
rect 55400 -11100 55500 -10700
rect 56000 -11100 56100 -10700
rect 59600 -10700 59700 -10300
rect 60400 -10700 60500 -10300
rect 59600 -10800 60500 -10700
rect 66800 -10300 67500 -10200
rect 66800 -10700 66900 -10300
rect 67400 -10700 67500 -10300
rect 55400 -11200 56100 -11100
rect 51400 -11900 51500 -11700
rect 52500 -11900 52600 -11700
rect 51400 -17100 52600 -11900
rect 55320 -11660 55800 -11600
rect 55320 -11980 55380 -11660
rect 55740 -11980 55800 -11660
rect 55320 -12040 55800 -11980
rect 53460 -12340 53800 -12320
rect 53460 -12540 53480 -12340
rect 53780 -12540 53800 -12340
rect 53460 -12560 53800 -12540
rect 57800 -13820 58240 -13810
rect 56900 -13940 57800 -13820
rect 57800 -13950 58240 -13940
rect 59700 -15600 60400 -15500
rect 59700 -15900 59800 -15600
rect 60300 -15900 60400 -15600
rect 59700 -16000 60400 -15900
rect 65800 -15600 66500 -15500
rect 65800 -15900 65900 -15600
rect 66400 -15900 66500 -15600
rect 55400 -16100 56100 -16000
rect 55400 -16500 55500 -16100
rect 56000 -16500 56100 -16100
rect 55400 -16600 56100 -16500
rect 51400 -17300 51500 -17100
rect 52500 -17300 52600 -17100
rect 51400 -22500 52600 -17300
rect 55360 -17100 55740 -17060
rect 55360 -17400 55400 -17100
rect 55700 -17400 55740 -17100
rect 55360 -17420 55740 -17400
rect 53480 -17740 53800 -17720
rect 53480 -17940 53500 -17740
rect 53780 -17940 53800 -17740
rect 53480 -17960 53800 -17940
rect 57800 -19220 58240 -19210
rect 56900 -19340 57800 -19220
rect 57800 -19350 58240 -19340
rect 59700 -21000 60400 -20900
rect 59700 -21300 59800 -21000
rect 60300 -21300 60400 -21000
rect 59700 -21400 60400 -21300
rect 64800 -21000 65500 -20900
rect 64800 -21300 64900 -21000
rect 65400 -21300 65500 -21000
rect 55400 -21500 56200 -21400
rect 55400 -21900 55500 -21500
rect 56100 -21900 56200 -21500
rect 55400 -22000 56200 -21900
rect 51400 -22700 51500 -22500
rect 52500 -22700 52600 -22500
rect 51400 -27900 52600 -22700
rect 55420 -22480 55740 -22460
rect 55420 -22760 55440 -22480
rect 55720 -22760 55740 -22480
rect 55420 -22780 55740 -22760
rect 53460 -23140 53800 -23120
rect 53460 -23340 53480 -23140
rect 53780 -23340 53800 -23140
rect 53460 -23360 53800 -23340
rect 57800 -24620 58240 -24610
rect 56900 -24740 57800 -24620
rect 57800 -24750 58240 -24740
rect 59600 -26400 60500 -26300
rect 59600 -26800 59700 -26400
rect 60400 -26800 60500 -26400
rect 55400 -26900 56200 -26800
rect 59600 -26900 60500 -26800
rect 63600 -26400 64200 -26300
rect 63600 -26800 63700 -26400
rect 64100 -26800 64200 -26400
rect 55400 -27300 55500 -26900
rect 56100 -27300 56200 -26900
rect 55400 -27400 56200 -27300
rect 51400 -28100 51500 -27900
rect 52500 -28100 52600 -27900
rect 51400 -33300 52600 -28100
rect 55440 -27880 55740 -27860
rect 55440 -28160 55460 -27880
rect 55720 -28160 55740 -27880
rect 55440 -28180 55740 -28160
rect 53460 -28540 53800 -28520
rect 53460 -28740 53480 -28540
rect 53780 -28740 53800 -28540
rect 53460 -28760 53800 -28740
rect 57800 -30020 58240 -30010
rect 56920 -30140 57800 -30020
rect 57800 -30150 58240 -30140
rect 59700 -31800 60400 -31700
rect 59700 -32100 59800 -31800
rect 60300 -32100 60400 -31800
rect 59700 -32200 60400 -32100
rect 62800 -31800 63400 -31700
rect 62800 -32100 62900 -31800
rect 63300 -32100 63400 -31800
rect 55400 -32300 56200 -32200
rect 55400 -32700 55500 -32300
rect 56100 -32700 56200 -32300
rect 55400 -32800 56200 -32700
rect 51400 -33500 51500 -33300
rect 52500 -33500 52600 -33300
rect 51400 -38700 52600 -33500
rect 55440 -33280 55740 -33260
rect 55440 -33560 55460 -33280
rect 55720 -33560 55740 -33280
rect 55440 -33580 55740 -33560
rect 53460 -33940 53800 -33920
rect 53460 -34140 53480 -33940
rect 53780 -34140 53800 -33940
rect 53460 -34160 53800 -34140
rect 57800 -35420 58240 -35410
rect 56900 -35540 57800 -35420
rect 57800 -35550 58240 -35540
rect 61900 -37100 62600 -37000
rect 59800 -37200 60300 -37100
rect 59800 -37400 59900 -37200
rect 60200 -37400 60300 -37200
rect 59800 -37500 60300 -37400
rect 55300 -37700 56200 -37600
rect 55300 -38100 55400 -37700
rect 56100 -38100 56200 -37700
rect 55300 -38200 56200 -38100
rect 61900 -37700 62000 -37100
rect 62500 -37700 62600 -37100
rect 51400 -38900 51500 -38700
rect 52500 -38900 52600 -38700
rect 51400 -44100 52600 -38900
rect 55440 -38680 55740 -38660
rect 55440 -38960 55460 -38680
rect 55720 -38960 55740 -38680
rect 55440 -38980 55740 -38960
rect 53460 -39340 53800 -39320
rect 53460 -39540 53480 -39340
rect 53780 -39540 53800 -39340
rect 53460 -39560 53800 -39540
rect 57800 -40820 58240 -40810
rect 56900 -40940 57800 -40820
rect 57800 -40950 58240 -40940
rect 61900 -41500 62600 -37700
rect 62800 -41000 63400 -32100
rect 63600 -40660 64200 -26800
rect 64800 -40200 65500 -21300
rect 65800 -39800 66500 -15900
rect 66800 -39400 67500 -10700
rect 68000 -39000 68700 -5200
rect 71900 -34100 74100 -34000
rect 71900 -35500 72000 -34100
rect 74000 -35500 74100 -34100
rect 71900 -35600 74100 -35500
rect 72800 -38900 73100 -35600
rect 68000 -39200 68100 -39000
rect 68600 -39200 68700 -39000
rect 68000 -39300 68700 -39200
rect 66800 -39600 66900 -39400
rect 67400 -39600 67500 -39400
rect 66800 -39800 67500 -39600
rect 65800 -40000 65900 -39800
rect 66400 -40000 66500 -39800
rect 65800 -40100 66500 -40000
rect 64800 -40400 64900 -40200
rect 65400 -40400 65500 -40200
rect 64800 -40500 65500 -40400
rect 63600 -40800 63640 -40660
rect 64160 -40800 64200 -40660
rect 63600 -40840 64200 -40800
rect 62800 -41300 62900 -41000
rect 63300 -41300 63400 -41000
rect 62800 -41400 63400 -41300
rect 61900 -41700 62000 -41500
rect 62500 -41700 62600 -41500
rect 61900 -41800 62600 -41700
rect 59600 -42800 60600 -42600
rect 55400 -43100 56200 -43000
rect 55400 -43500 55500 -43100
rect 56100 -43500 56200 -43100
rect 55400 -43600 56200 -43500
rect 59600 -43400 59800 -42800
rect 60400 -43400 60600 -42800
rect 59600 -43600 60600 -43400
rect 51400 -44300 51500 -44100
rect 52500 -44300 52600 -44100
rect 51400 -49500 52600 -44300
rect 55480 -44080 55740 -44060
rect 55480 -44360 55500 -44080
rect 55720 -44360 55740 -44080
rect 55480 -44380 55740 -44360
rect 53460 -44740 53800 -44720
rect 53460 -44940 53480 -44740
rect 53780 -44940 53800 -44740
rect 53460 -44960 53800 -44940
rect 57800 -46220 58240 -46210
rect 56920 -46340 57800 -46220
rect 57800 -46350 58240 -46340
rect 62400 -47200 63000 -47100
rect 62400 -47500 62500 -47200
rect 62900 -47500 63000 -47200
rect 59600 -48000 60500 -47900
rect 59600 -48400 59700 -48000
rect 60400 -48400 60500 -48000
rect 55400 -48500 56200 -48400
rect 59600 -48500 60500 -48400
rect 62400 -48000 63000 -47500
rect 62400 -48400 62500 -48000
rect 62900 -48400 63000 -48000
rect 62400 -48500 63000 -48400
rect 64100 -47700 64600 -47600
rect 64100 -47900 64200 -47700
rect 64500 -47900 64600 -47700
rect 55400 -48900 55500 -48500
rect 56100 -48900 56200 -48500
rect 55400 -49000 56200 -48900
rect 51400 -49700 51500 -49500
rect 52500 -49700 52600 -49500
rect 51400 -54900 52600 -49700
rect 55440 -49480 55740 -49460
rect 55440 -49760 55460 -49480
rect 55720 -49760 55740 -49480
rect 55440 -49780 55740 -49760
rect 53440 -50140 53800 -50120
rect 53440 -50340 53460 -50140
rect 53780 -50340 53800 -50140
rect 53440 -50360 53800 -50340
rect 57800 -51620 58240 -51610
rect 56900 -51740 57800 -51620
rect 57800 -51750 58240 -51740
rect 59600 -53400 60500 -53300
rect 59600 -53800 59700 -53400
rect 60400 -53800 60500 -53400
rect 55300 -53900 56200 -53800
rect 59600 -53900 60500 -53800
rect 64100 -53400 64600 -47900
rect 64100 -53800 64200 -53400
rect 64500 -53800 64600 -53400
rect 64100 -53900 64600 -53800
rect 65000 -48100 65500 -48000
rect 65000 -48300 65100 -48100
rect 65400 -48300 65500 -48100
rect 55300 -54300 55400 -53900
rect 56100 -54300 56200 -53900
rect 55300 -54400 56200 -54300
rect 51400 -55100 51500 -54900
rect 52500 -55100 52600 -54900
rect 51400 -60300 52600 -55100
rect 55440 -54880 55740 -54860
rect 55440 -55160 55460 -54880
rect 55720 -55160 55740 -54880
rect 55440 -55180 55740 -55160
rect 53460 -55540 53800 -55520
rect 53460 -55740 53480 -55540
rect 53780 -55740 53800 -55540
rect 53460 -55760 53800 -55740
rect 57800 -57020 58240 -57010
rect 56900 -57140 57800 -57020
rect 57800 -57150 58240 -57140
rect 59600 -58800 60500 -58700
rect 59600 -59200 59700 -58800
rect 60400 -59200 60500 -58800
rect 55400 -59300 56200 -59200
rect 59600 -59300 60500 -59200
rect 65000 -58800 65500 -48300
rect 65000 -59200 65100 -58800
rect 65400 -59200 65500 -58800
rect 65000 -59300 65500 -59200
rect 66000 -48500 66500 -48400
rect 66000 -48700 66100 -48500
rect 66400 -48700 66500 -48500
rect 55400 -59700 55500 -59300
rect 56100 -59700 56200 -59300
rect 55400 -59800 56200 -59700
rect 51400 -60500 51500 -60300
rect 52500 -60500 52600 -60300
rect 51400 -65700 52600 -60500
rect 55440 -60280 55740 -60260
rect 55440 -60560 55460 -60280
rect 55720 -60560 55740 -60280
rect 55440 -60580 55740 -60560
rect 53460 -60940 53800 -60920
rect 53460 -61140 53480 -60940
rect 53780 -61140 53800 -60940
rect 53460 -61160 53800 -61140
rect 57800 -62420 58240 -62410
rect 56920 -62540 57800 -62420
rect 57800 -62550 58240 -62540
rect 59600 -64200 60500 -64100
rect 59600 -64600 59700 -64200
rect 60400 -64600 60500 -64200
rect 55400 -64700 56200 -64600
rect 59600 -64700 60500 -64600
rect 66000 -64200 66500 -48700
rect 66000 -64600 66100 -64200
rect 66400 -64600 66500 -64200
rect 66000 -64700 66500 -64600
rect 67000 -48900 67500 -48800
rect 67000 -49100 67100 -48900
rect 67400 -49100 67500 -48900
rect 55400 -65100 55500 -64700
rect 56100 -65100 56200 -64700
rect 55400 -65200 56200 -65100
rect 51400 -65900 51500 -65700
rect 52500 -65900 52600 -65700
rect 51400 -71100 52600 -65900
rect 55420 -65680 55740 -65660
rect 55420 -65960 55440 -65680
rect 55720 -65960 55740 -65680
rect 55420 -65980 55740 -65960
rect 53460 -66340 53800 -66320
rect 53460 -66540 53480 -66340
rect 53780 -66540 53800 -66340
rect 53460 -66560 53800 -66540
rect 57800 -67820 58240 -67810
rect 56900 -67940 57800 -67820
rect 57800 -67950 58240 -67940
rect 59600 -69600 60500 -69500
rect 59600 -70000 59700 -69600
rect 60400 -70000 60500 -69600
rect 55400 -70100 56200 -70000
rect 59600 -70100 60500 -70000
rect 67000 -69600 67500 -49100
rect 67000 -70000 67100 -69600
rect 67400 -70000 67500 -69600
rect 67000 -70100 67500 -70000
rect 67900 -49300 68400 -49200
rect 67900 -49500 68000 -49300
rect 68300 -49500 68400 -49300
rect 55400 -70500 55500 -70100
rect 56100 -70500 56200 -70100
rect 55400 -70600 56200 -70500
rect 51400 -71300 51500 -71100
rect 52500 -71300 52600 -71100
rect 51400 -76500 52600 -71300
rect 55440 -71080 55740 -71060
rect 55440 -71360 55460 -71080
rect 55720 -71360 55740 -71080
rect 55440 -71380 55740 -71360
rect 53460 -71740 53800 -71720
rect 53460 -71940 53480 -71740
rect 53780 -71940 53800 -71740
rect 53460 -71960 53800 -71940
rect 57800 -73220 58240 -73210
rect 56900 -73340 57800 -73220
rect 57800 -73350 58240 -73340
rect 59600 -75000 60500 -74900
rect 59600 -75400 59700 -75000
rect 60400 -75400 60500 -75000
rect 55400 -75500 56200 -75400
rect 59600 -75500 60500 -75400
rect 67900 -75000 68400 -49500
rect 67900 -75400 68000 -75000
rect 68300 -75400 68400 -75000
rect 67900 -75500 68400 -75400
rect 68900 -49700 69400 -49600
rect 68900 -49900 69000 -49700
rect 69300 -49900 69400 -49700
rect 55400 -75900 55500 -75500
rect 56100 -75900 56200 -75500
rect 55400 -76000 56200 -75900
rect 51400 -76700 51500 -76500
rect 52500 -76700 52600 -76500
rect 51400 -81900 52600 -76700
rect 55380 -76480 55740 -76460
rect 55380 -76760 55400 -76480
rect 55720 -76760 55740 -76480
rect 55380 -76780 55740 -76760
rect 53460 -77140 53800 -77120
rect 53460 -77340 53480 -77140
rect 53780 -77340 53800 -77140
rect 53460 -77360 53800 -77340
rect 57800 -78620 58240 -78610
rect 56900 -78740 57800 -78620
rect 57800 -78750 58240 -78740
rect 59600 -80400 60500 -80300
rect 59600 -80800 59700 -80400
rect 60400 -80800 60500 -80400
rect 55400 -80900 56300 -80800
rect 59600 -80900 60500 -80800
rect 68900 -80400 69400 -49900
rect 68900 -80800 69000 -80400
rect 69300 -80800 69400 -80400
rect 68900 -80900 69400 -80800
rect 69900 -50100 70400 -50000
rect 69900 -50300 70000 -50100
rect 70300 -50300 70400 -50100
rect 55400 -81300 55500 -80900
rect 56200 -81300 56300 -80900
rect 55400 -81400 56300 -81300
rect 51400 -82100 51500 -81900
rect 52500 -82100 52600 -81900
rect 37100 -86700 37200 -86200
rect 37700 -86700 37800 -86200
rect 51400 -86700 52600 -82100
rect 55420 -81880 55740 -81860
rect 55420 -82160 55440 -81880
rect 55720 -82160 55740 -81880
rect 55420 -82180 55740 -82160
rect 53460 -82540 53800 -82520
rect 53460 -82740 53480 -82540
rect 53780 -82740 53800 -82540
rect 53460 -82760 53800 -82740
rect 57800 -84020 58240 -84010
rect 56900 -84140 57800 -84020
rect 57800 -84150 58240 -84140
rect 59600 -85800 60500 -85700
rect 59600 -86200 59700 -85800
rect 60400 -86200 60500 -85800
rect 55400 -86300 56200 -86200
rect 59600 -86300 60500 -86200
rect 69900 -85800 70400 -50300
rect 69900 -86200 70000 -85800
rect 70300 -86200 70400 -85800
rect 69900 -86300 70400 -86200
rect 55400 -86600 55500 -86300
rect 56100 -86600 56200 -86300
rect 55400 -86700 56200 -86600
rect 37100 -86800 37800 -86700
<< via2 >>
rect 38000 1400 41400 2800
rect 43000 1000 46400 2400
rect 37900 -3600 41500 -400
rect 43000 -1400 46400 0
rect 56880 -40 59080 1020
rect 51500 -1000 52500 -800
rect 47700 -1700 48000 -1300
rect 36400 -5800 37000 -5000
rect 21000 -7400 22000 -6600
rect 24700 -9400 25700 -8700
rect 27200 -13000 34400 -10600
rect 15000 -31200 19400 -26400
rect 26600 -30400 35200 -26400
rect 47640 -7200 48080 -6780
rect 46700 -9400 47800 -8700
rect 37600 -11100 38100 -10700
rect 47700 -12640 48080 -12220
rect 38500 -16600 39000 -16000
rect 47640 -18100 48080 -17620
rect 39500 -22000 40000 -21400
rect 47680 -23440 48080 -23020
rect 40400 -27400 41000 -26800
rect 15000 -49000 24000 -38000
rect 47800 -28840 48080 -28460
rect 41500 -32800 42100 -32200
rect 47760 -34200 48080 -33860
rect 42500 -38200 43100 -37600
rect 47760 -39640 48080 -39220
rect 43200 -43300 44300 -43100
rect 43200 -43800 44300 -43300
rect 15200 -64800 19600 -60000
rect 25000 -64800 35400 -58800
rect 43800 -49000 44300 -48400
rect 47820 -45060 48080 -44640
rect 42900 -54400 43400 -53800
rect 47740 -50480 48080 -49980
rect 42000 -59800 42500 -59200
rect 47820 -55820 48080 -55460
rect 41100 -65200 41600 -64600
rect 47680 -61300 48080 -60760
rect 40200 -70600 40700 -70000
rect 47860 -66660 48080 -66220
rect 39300 -76000 39800 -75400
rect 47720 -72060 48080 -71600
rect 38300 -81400 38800 -80800
rect 47780 -77500 48080 -76940
rect 47800 -82860 48080 -82380
rect 55400 -1000 55700 -600
rect 53400 -1600 53700 -1400
rect 57800 -3140 58240 -3020
rect 59700 -5200 60400 -4900
rect 68100 -5200 68600 -4900
rect 55600 -5600 55900 -5300
rect 51500 -6500 52500 -6300
rect 55400 -6500 55700 -6200
rect 53520 -7120 53780 -6860
rect 57800 -8540 58240 -8420
rect 55500 -11100 56000 -10700
rect 59700 -10700 60400 -10300
rect 66900 -10700 67400 -10300
rect 51500 -11900 52500 -11700
rect 55380 -11980 55740 -11660
rect 53480 -12540 53780 -12340
rect 57800 -13940 58240 -13820
rect 59800 -15900 60300 -15600
rect 65900 -15900 66400 -15600
rect 55500 -16500 56000 -16100
rect 51500 -17300 52500 -17100
rect 55400 -17400 55700 -17100
rect 53500 -17940 53780 -17740
rect 57800 -19340 58240 -19220
rect 59800 -21300 60300 -21000
rect 64900 -21300 65400 -21000
rect 55500 -21900 56100 -21500
rect 51500 -22700 52500 -22500
rect 55440 -22760 55720 -22480
rect 53480 -23340 53780 -23140
rect 57800 -24740 58240 -24620
rect 59700 -26800 60400 -26400
rect 63700 -26800 64100 -26400
rect 55500 -27300 56100 -26900
rect 51500 -28100 52500 -27900
rect 55460 -28160 55720 -27880
rect 53480 -28740 53780 -28540
rect 57800 -30140 58240 -30020
rect 59800 -32100 60300 -31800
rect 62900 -32100 63300 -31800
rect 55500 -32700 56100 -32300
rect 51500 -33500 52500 -33300
rect 55460 -33560 55720 -33280
rect 53480 -34140 53780 -33940
rect 57800 -35540 58240 -35420
rect 59900 -37400 60200 -37200
rect 55400 -38100 56100 -37700
rect 62000 -37700 62500 -37100
rect 51500 -38900 52500 -38700
rect 55460 -38960 55720 -38680
rect 53480 -39540 53780 -39340
rect 57800 -40940 58240 -40820
rect 72000 -35500 74000 -34100
rect 68100 -39200 68600 -39000
rect 66900 -39600 67400 -39400
rect 65900 -40000 66400 -39800
rect 64900 -40400 65400 -40200
rect 63640 -40800 64160 -40660
rect 62900 -41300 63300 -41000
rect 62000 -41700 62500 -41500
rect 55500 -43500 56100 -43100
rect 59800 -43400 60400 -42800
rect 51500 -44300 52500 -44100
rect 55500 -44360 55720 -44080
rect 53480 -44940 53780 -44740
rect 57800 -46340 58240 -46220
rect 62500 -47500 62900 -47200
rect 59700 -48400 60400 -48000
rect 62500 -48400 62900 -48000
rect 64200 -47900 64500 -47700
rect 55500 -48900 56100 -48500
rect 51500 -49700 52500 -49500
rect 55460 -49760 55720 -49480
rect 53460 -50340 53780 -50140
rect 57800 -51740 58240 -51620
rect 59700 -53800 60400 -53400
rect 64200 -53800 64500 -53400
rect 65100 -48300 65400 -48100
rect 55400 -54300 56100 -53900
rect 51500 -55100 52500 -54900
rect 55460 -55160 55720 -54880
rect 53480 -55740 53780 -55540
rect 57800 -57140 58240 -57020
rect 59700 -59200 60400 -58800
rect 65100 -59200 65400 -58800
rect 66100 -48700 66400 -48500
rect 55500 -59700 56100 -59300
rect 51500 -60500 52500 -60300
rect 55460 -60560 55720 -60280
rect 53480 -61140 53780 -60940
rect 57800 -62540 58240 -62420
rect 59700 -64600 60400 -64200
rect 66100 -64600 66400 -64200
rect 67100 -49100 67400 -48900
rect 55500 -65100 56100 -64700
rect 51500 -65900 52500 -65700
rect 55440 -65960 55720 -65680
rect 53480 -66540 53780 -66340
rect 57800 -67940 58240 -67820
rect 59700 -70000 60400 -69600
rect 67100 -70000 67400 -69600
rect 68000 -49500 68300 -49300
rect 55500 -70500 56100 -70100
rect 51500 -71300 52500 -71100
rect 55460 -71360 55720 -71080
rect 53480 -71940 53780 -71740
rect 57800 -73340 58240 -73220
rect 59700 -75400 60400 -75000
rect 68000 -75400 68300 -75000
rect 69000 -49900 69300 -49700
rect 55500 -75900 56100 -75500
rect 51500 -76700 52500 -76500
rect 55400 -76760 55720 -76480
rect 53480 -77340 53780 -77140
rect 57800 -78740 58240 -78620
rect 59700 -80800 60400 -80400
rect 69000 -80800 69300 -80400
rect 70000 -50300 70300 -50100
rect 55500 -81300 56200 -80900
rect 51500 -82100 52500 -81900
rect 37200 -86700 37700 -86200
rect 55440 -82160 55720 -81880
rect 53480 -82740 53780 -82540
rect 57800 -84140 58240 -84020
rect 59700 -86200 60400 -85800
rect 70000 -86200 70300 -85800
rect 55500 -86600 56100 -86300
<< metal3 >>
rect 10100 -2000 10500 -1500
rect 11000 -2000 11600 -1500
rect 12100 -2000 12700 -1500
rect 13200 -2000 13800 -1500
rect 14300 -2000 27500 -1500
rect 10100 -2500 27500 -2000
rect 10100 -3000 10500 -2500
rect 11000 -3000 11600 -2500
rect 12100 -3000 12700 -2500
rect 13200 -3000 13800 -2500
rect 14300 -3000 27500 -2500
rect 10100 -3500 27500 -3000
rect 10100 -4000 10500 -3500
rect 11000 -4000 11600 -3500
rect 12100 -4000 12700 -3500
rect 13200 -4000 13800 -3500
rect 14300 -4000 27500 -3500
rect 10100 -4500 27500 -4000
rect 10100 -5000 10500 -4500
rect 11000 -5000 11600 -4500
rect 12100 -5000 12700 -4500
rect 13200 -5000 13800 -4500
rect 14300 -5000 27500 -4500
rect 24300 -6000 27500 -5000
rect 35000 -6000 35600 5000
rect 37800 2800 41600 3000
rect 37800 1400 38000 2800
rect 41400 1400 41600 2800
rect 37800 1200 41600 1400
rect 42800 2400 46600 2600
rect 42800 1000 43000 2400
rect 46400 1000 46600 2400
rect 42800 800 46600 1000
rect 56870 1020 59090 1025
rect 42800 0 46600 200
rect 37800 -400 41600 -300
rect 37800 -3600 37900 -400
rect 41500 -3600 41600 -400
rect 42800 -1400 43000 0
rect 46400 -1400 46600 0
rect 56870 -40 56880 1020
rect 59080 -40 59090 1020
rect 56870 -45 59090 -40
rect 55300 -600 55800 -500
rect 55300 -700 55400 -600
rect 51400 -800 55400 -700
rect 51400 -1000 51500 -800
rect 52500 -1000 55400 -800
rect 55700 -1000 55800 -600
rect 51400 -1100 55800 -1000
rect 42800 -1600 46600 -1400
rect 47600 -1300 48100 -1200
rect 47600 -1700 47700 -1300
rect 48000 -1400 53800 -1300
rect 48000 -1600 53400 -1400
rect 53700 -1600 53800 -1400
rect 48000 -1700 53800 -1600
rect 47600 -1800 48100 -1700
rect 37800 -3700 41600 -3600
rect 57760 -3020 58280 -45
rect 57760 -3140 57800 -3020
rect 58240 -3140 58280 -3020
rect 36200 -5000 37200 -4800
rect 36200 -5800 36400 -5000
rect 37000 -5200 37200 -5000
rect 37000 -5300 56000 -5200
rect 37000 -5600 55600 -5300
rect 55900 -5600 56000 -5300
rect 37000 -5700 56000 -5600
rect 37000 -5800 37200 -5700
rect 36200 -6000 37200 -5800
rect 20800 -6600 22500 -6200
rect 20800 -7400 21000 -6600
rect 22000 -7400 22500 -6600
rect 20800 -7500 22500 -7400
rect 24300 -8600 35600 -6000
rect 55300 -6200 55800 -6100
rect 51400 -6300 55400 -6200
rect 51400 -6500 51500 -6300
rect 52500 -6500 55400 -6300
rect 55700 -6500 55800 -6200
rect 51400 -6600 55800 -6500
rect 47620 -6780 48100 -6760
rect 47620 -7200 47640 -6780
rect 48080 -6840 48100 -6780
rect 48080 -6860 53800 -6840
rect 48080 -7120 53520 -6860
rect 53780 -7120 53800 -6860
rect 48080 -7140 53800 -7120
rect 48080 -7200 48100 -7140
rect 47620 -7220 48100 -7200
rect 57760 -8420 58280 -3140
rect 59600 -4900 68700 -4800
rect 59600 -5200 59700 -4900
rect 60400 -5200 68100 -4900
rect 68600 -5200 68700 -4900
rect 59600 -5300 68700 -5200
rect 57760 -8540 57800 -8420
rect 58240 -8540 58280 -8420
rect 24300 -8700 47900 -8600
rect 24300 -9400 24700 -8700
rect 25700 -9400 46700 -8700
rect 47800 -9400 47900 -8700
rect 24300 -9500 47900 -9400
rect 31328 -9838 32878 -9500
rect 27000 -10600 34600 -10400
rect 27000 -13000 27200 -10600
rect 34400 -13000 34600 -10600
rect 37500 -10700 56100 -10600
rect 37500 -11100 37600 -10700
rect 38100 -11100 55500 -10700
rect 56000 -11100 56100 -10700
rect 37500 -11200 56100 -11100
rect 51400 -11660 55800 -11600
rect 51400 -11700 55380 -11660
rect 51400 -11900 51500 -11700
rect 52500 -11900 55380 -11700
rect 51400 -11980 55380 -11900
rect 55740 -11980 55800 -11660
rect 51400 -12000 55800 -11980
rect 55320 -12040 55800 -12000
rect 47680 -12220 48100 -12200
rect 47680 -12640 47700 -12220
rect 48080 -12320 48100 -12220
rect 48080 -12340 53800 -12320
rect 48080 -12540 53480 -12340
rect 53780 -12540 53800 -12340
rect 48080 -12560 53800 -12540
rect 48080 -12640 48100 -12560
rect 47680 -12660 48100 -12640
rect 27000 -13200 34600 -13000
rect 57760 -13820 58280 -8540
rect 59600 -10300 67500 -10200
rect 59600 -10700 59700 -10300
rect 60400 -10700 66900 -10300
rect 67400 -10700 67500 -10300
rect 59600 -10800 67500 -10700
rect 57760 -13940 57800 -13820
rect 58240 -13940 58280 -13820
rect 38400 -16000 39100 -15900
rect 38400 -16600 38500 -16000
rect 39000 -16100 56100 -16000
rect 39000 -16500 55500 -16100
rect 56000 -16500 56100 -16100
rect 39000 -16600 56100 -16500
rect 38400 -16700 39100 -16600
rect 51400 -17100 55800 -17000
rect 51400 -17300 51500 -17100
rect 52500 -17300 55400 -17100
rect 51400 -17400 55400 -17300
rect 55700 -17400 55800 -17100
rect 55300 -17500 55800 -17400
rect 47620 -17620 48100 -17600
rect 47620 -18100 47640 -17620
rect 48080 -17720 48100 -17620
rect 48080 -17740 53800 -17720
rect 48080 -17940 53500 -17740
rect 53780 -17940 53800 -17740
rect 48080 -17960 53800 -17940
rect 48080 -18100 48100 -17960
rect 47620 -18120 48100 -18100
rect 57760 -19220 58280 -13940
rect 59700 -15600 66500 -15500
rect 59700 -15900 59800 -15600
rect 60300 -15900 65900 -15600
rect 66400 -15900 66500 -15600
rect 59700 -16000 66500 -15900
rect 57760 -19340 57800 -19220
rect 58240 -19340 58280 -19220
rect 39400 -21400 40100 -21300
rect 39400 -22000 39500 -21400
rect 40000 -21500 56200 -21400
rect 40000 -21900 55500 -21500
rect 56100 -21900 56200 -21500
rect 40000 -22000 56200 -21900
rect 39400 -22100 40100 -22000
rect 51400 -22480 55800 -22400
rect 51400 -22500 55440 -22480
rect 51400 -22700 51500 -22500
rect 52500 -22700 55440 -22500
rect 51400 -22760 55440 -22700
rect 55720 -22760 55800 -22480
rect 51400 -22800 55800 -22760
rect 55360 -22840 55800 -22800
rect 47660 -23020 48100 -23000
rect 47660 -23440 47680 -23020
rect 48080 -23120 48100 -23020
rect 48080 -23140 53800 -23120
rect 48080 -23340 53480 -23140
rect 53780 -23340 53800 -23140
rect 48080 -23360 53800 -23340
rect 48080 -23440 48100 -23360
rect 47660 -23460 48100 -23440
rect 57760 -24620 58280 -19340
rect 59700 -21000 65500 -20900
rect 59700 -21300 59800 -21000
rect 60300 -21300 64900 -21000
rect 65400 -21300 65500 -21000
rect 59700 -21400 65500 -21300
rect 57760 -24740 57800 -24620
rect 58240 -24740 58280 -24620
rect 14400 -26400 36000 -25800
rect 14400 -31200 15000 -26400
rect 19400 -30400 26600 -26400
rect 35200 -30400 36000 -26400
rect 40300 -26800 41100 -26700
rect 40300 -27400 40400 -26800
rect 41000 -26900 56200 -26800
rect 41000 -27300 55500 -26900
rect 56100 -27300 56200 -26900
rect 41000 -27400 56200 -27300
rect 40300 -27500 41100 -27400
rect 51400 -27880 55800 -27800
rect 51400 -27900 55460 -27880
rect 51400 -28100 51500 -27900
rect 52500 -28100 55460 -27900
rect 51400 -28160 55460 -28100
rect 55720 -28160 55800 -27880
rect 51400 -28200 55800 -28160
rect 55380 -28240 55800 -28200
rect 47780 -28460 48100 -28440
rect 47780 -28840 47800 -28460
rect 48080 -28520 48100 -28460
rect 48080 -28540 53800 -28520
rect 48080 -28740 53480 -28540
rect 53780 -28740 53800 -28540
rect 48080 -28760 53800 -28740
rect 48080 -28840 48100 -28760
rect 47780 -28860 48100 -28840
rect 19400 -31200 36000 -30400
rect 14400 -31800 36000 -31200
rect 57760 -30020 58280 -24740
rect 59600 -26400 64200 -26300
rect 59600 -26800 59700 -26400
rect 60400 -26800 63700 -26400
rect 64100 -26800 64200 -26400
rect 59600 -26900 64200 -26800
rect 57760 -30140 57800 -30020
rect 58240 -30140 58280 -30020
rect 41400 -32200 42200 -32100
rect 41400 -32800 41500 -32200
rect 42100 -32300 56200 -32200
rect 42100 -32700 55500 -32300
rect 56100 -32700 56200 -32300
rect 42100 -32800 56200 -32700
rect 41400 -32900 42200 -32800
rect 51400 -33280 55800 -33200
rect 51400 -33300 55460 -33280
rect 51400 -33500 51500 -33300
rect 52500 -33500 55460 -33300
rect 51400 -33560 55460 -33500
rect 55720 -33560 55800 -33280
rect 51400 -33600 55800 -33560
rect 55380 -33640 55800 -33600
rect 47740 -33860 48100 -33840
rect 47740 -34200 47760 -33860
rect 48080 -33920 48100 -33860
rect 48080 -33940 53800 -33920
rect 48080 -34140 53480 -33940
rect 53780 -34140 53800 -33940
rect 48080 -34160 53800 -34140
rect 48080 -34200 48100 -34160
rect 47740 -34220 48100 -34200
rect 57760 -35420 58280 -30140
rect 59700 -31800 63400 -31700
rect 59700 -32100 59800 -31800
rect 60300 -32100 62900 -31800
rect 63300 -32100 63400 -31800
rect 59700 -32200 63400 -32100
rect 57760 -35540 57800 -35420
rect 58240 -35540 58280 -35420
rect 14000 -38000 25000 -37000
rect 14000 -49000 15000 -38000
rect 24000 -49000 25000 -38000
rect 42400 -37600 43200 -37500
rect 42400 -38200 42500 -37600
rect 43100 -37700 56200 -37600
rect 43100 -38100 55400 -37700
rect 56100 -38100 56200 -37700
rect 43100 -38200 56200 -38100
rect 42400 -38300 43200 -38200
rect 51400 -38680 55800 -38600
rect 51400 -38700 55460 -38680
rect 51400 -38900 51500 -38700
rect 52500 -38900 55460 -38700
rect 51400 -38960 55460 -38900
rect 55720 -38960 55800 -38680
rect 51400 -39000 55800 -38960
rect 55380 -39040 55800 -39000
rect 47740 -39220 48100 -39200
rect 47740 -39640 47760 -39220
rect 48080 -39320 48100 -39220
rect 48080 -39340 53800 -39320
rect 48080 -39540 53480 -39340
rect 53780 -39540 53800 -39340
rect 48080 -39560 53800 -39540
rect 48080 -39640 48100 -39560
rect 47740 -39660 48100 -39640
rect 57760 -40820 58280 -35540
rect 71900 -34100 74100 -34000
rect 71900 -35500 72000 -34100
rect 74000 -35500 74100 -34100
rect 71900 -35600 74100 -35500
rect 61900 -37100 62600 -37000
rect 59800 -37200 60300 -37100
rect 61900 -37200 62000 -37100
rect 59800 -37400 59900 -37200
rect 60200 -37400 62000 -37200
rect 59800 -37500 62000 -37400
rect 61900 -37700 62000 -37500
rect 62500 -37700 62600 -37100
rect 61900 -37800 62600 -37700
rect 68000 -39000 68700 -38900
rect 72600 -38920 73080 -38740
rect 68000 -39200 68100 -39000
rect 68600 -39060 68700 -39000
rect 68600 -39200 73080 -39060
rect 68000 -39240 73080 -39200
rect 68000 -39300 68700 -39240
rect 66800 -39400 67500 -39300
rect 66800 -39600 66900 -39400
rect 67400 -39560 67500 -39400
rect 67400 -39600 73200 -39560
rect 65800 -39800 66500 -39700
rect 66800 -39740 73200 -39600
rect 65800 -39839 65900 -39800
rect 65799 -40000 65900 -39839
rect 66400 -39839 66500 -39800
rect 66400 -39840 72399 -39839
rect 66400 -40000 73200 -39840
rect 65799 -40019 73200 -40000
rect 65800 -40100 66500 -40019
rect 66600 -40020 73200 -40019
rect 64800 -40200 65500 -40100
rect 64800 -40400 64900 -40200
rect 65400 -40300 65500 -40200
rect 65400 -40400 73200 -40300
rect 64800 -40480 73200 -40400
rect 64800 -40500 65500 -40480
rect 57760 -40940 57800 -40820
rect 58240 -40940 58280 -40820
rect 63600 -40660 64200 -40620
rect 63600 -40800 63640 -40660
rect 64160 -40800 73200 -40660
rect 63600 -40840 73200 -40800
rect 43100 -43100 56200 -43000
rect 43100 -43800 43200 -43100
rect 44300 -43500 55500 -43100
rect 56100 -43500 56200 -43100
rect 44300 -43600 56200 -43500
rect 44300 -43800 44400 -43600
rect 43100 -43900 44400 -43800
rect 51400 -44080 55800 -44000
rect 51400 -44100 55500 -44080
rect 51400 -44300 51500 -44100
rect 52500 -44300 55500 -44100
rect 51400 -44360 55500 -44300
rect 55720 -44360 55800 -44080
rect 51400 -44400 55800 -44360
rect 55420 -44440 55800 -44400
rect 47800 -44640 48100 -44620
rect 47800 -45060 47820 -44640
rect 48080 -44720 48100 -44640
rect 48080 -44740 53800 -44720
rect 48080 -44940 53480 -44740
rect 53780 -44940 53800 -44740
rect 48080 -44960 53800 -44940
rect 48080 -45060 48100 -44960
rect 47800 -45080 48100 -45060
rect 57760 -46220 58280 -40940
rect 62800 -41000 63400 -40900
rect 62800 -41300 62900 -41000
rect 63300 -41300 73200 -41000
rect 62800 -41400 63400 -41300
rect 61900 -41500 62600 -41400
rect 61900 -41700 62000 -41500
rect 62500 -41700 73100 -41500
rect 61900 -41800 62600 -41700
rect 72600 -42600 73200 -41900
rect 59600 -42800 73200 -42600
rect 59600 -43400 59800 -42800
rect 60400 -43400 73200 -42800
rect 59600 -43600 73200 -43400
rect 57760 -46340 57800 -46220
rect 58240 -46340 58280 -46220
rect 14000 -50000 25000 -49000
rect 43700 -48400 44400 -48300
rect 43700 -49000 43800 -48400
rect 44300 -48500 56200 -48400
rect 44300 -48900 55500 -48500
rect 56100 -48900 56200 -48500
rect 44300 -49000 56200 -48900
rect 43700 -49100 44400 -49000
rect 51400 -49480 55800 -49400
rect 51400 -49500 55460 -49480
rect 51400 -49700 51500 -49500
rect 52500 -49700 55460 -49500
rect 51400 -49760 55460 -49700
rect 55720 -49760 55800 -49480
rect 51400 -49800 55800 -49760
rect 55380 -49840 55800 -49800
rect 47720 -49980 48100 -49960
rect 47720 -50480 47740 -49980
rect 48080 -50120 48100 -49980
rect 48080 -50140 53800 -50120
rect 48080 -50340 53460 -50140
rect 53780 -50340 53800 -50140
rect 48080 -50360 53800 -50340
rect 48080 -50480 48100 -50360
rect 47720 -50500 48100 -50480
rect 57760 -51620 58280 -46340
rect 62400 -47200 63000 -47100
rect 63203 -47200 73103 -47199
rect 62400 -47500 62500 -47200
rect 62900 -47499 73103 -47200
rect 62900 -47500 63600 -47499
rect 62400 -47600 63000 -47500
rect 64100 -47700 73100 -47600
rect 64100 -47900 64200 -47700
rect 64500 -47900 73100 -47700
rect 59600 -48000 63000 -47900
rect 64100 -48000 64600 -47900
rect 59600 -48400 59700 -48000
rect 60400 -48400 62500 -48000
rect 62900 -48400 63000 -48000
rect 65000 -48100 73100 -48000
rect 65000 -48300 65100 -48100
rect 65400 -48300 73100 -48100
rect 65000 -48400 65500 -48300
rect 59600 -48500 63000 -48400
rect 66000 -48500 73100 -48400
rect 66000 -48700 66100 -48500
rect 66400 -48700 73100 -48500
rect 66000 -48800 66500 -48700
rect 67000 -48900 73100 -48800
rect 67000 -49100 67100 -48900
rect 67400 -49100 73100 -48900
rect 67000 -49200 67500 -49100
rect 67900 -49300 73100 -49200
rect 67900 -49500 68000 -49300
rect 68300 -49500 73100 -49300
rect 67900 -49600 68400 -49500
rect 68900 -49700 73100 -49600
rect 68900 -49900 69000 -49700
rect 69300 -49900 73100 -49700
rect 68900 -50000 69400 -49900
rect 69900 -50100 73100 -50000
rect 69900 -50300 70000 -50100
rect 70300 -50300 73100 -50100
rect 69900 -50400 70400 -50300
rect 57760 -51740 57800 -51620
rect 58240 -51740 58280 -51620
rect 42800 -53800 43500 -53700
rect 42800 -54400 42900 -53800
rect 43400 -53900 56200 -53800
rect 43400 -54300 55400 -53900
rect 56100 -54300 56200 -53900
rect 43400 -54400 56200 -54300
rect 42800 -54500 43500 -54400
rect 51400 -54880 55800 -54800
rect 51400 -54900 55460 -54880
rect 51400 -55100 51500 -54900
rect 52500 -55100 55460 -54900
rect 51400 -55160 55460 -55100
rect 55720 -55160 55800 -54880
rect 51400 -55200 55800 -55160
rect 55380 -55240 55800 -55200
rect 47800 -55460 48100 -55440
rect 47800 -55820 47820 -55460
rect 48080 -55520 48100 -55460
rect 48080 -55540 53800 -55520
rect 48080 -55740 53480 -55540
rect 53780 -55740 53800 -55540
rect 48080 -55760 53800 -55740
rect 48080 -55820 48100 -55760
rect 47800 -55840 48100 -55820
rect 57760 -57020 58280 -51740
rect 59600 -53400 64600 -53300
rect 59600 -53800 59700 -53400
rect 60400 -53800 64200 -53400
rect 64500 -53800 64600 -53400
rect 59600 -53900 64600 -53800
rect 57760 -57140 57800 -57020
rect 58240 -57140 58280 -57020
rect 24400 -58800 36000 -58200
rect 24400 -59400 25000 -58800
rect 14600 -60000 25000 -59400
rect 14600 -64800 15200 -60000
rect 19600 -64800 25000 -60000
rect 35400 -64800 36000 -58800
rect 41900 -59200 42600 -59100
rect 41900 -59800 42000 -59200
rect 42500 -59300 56200 -59200
rect 42500 -59700 55500 -59300
rect 56100 -59700 56200 -59300
rect 42500 -59800 56200 -59700
rect 41900 -59900 42600 -59800
rect 51400 -60280 55800 -60200
rect 51400 -60300 55460 -60280
rect 51400 -60500 51500 -60300
rect 52500 -60500 55460 -60300
rect 51400 -60560 55460 -60500
rect 55720 -60560 55800 -60280
rect 51400 -60600 55800 -60560
rect 55380 -60640 55800 -60600
rect 47660 -60760 48100 -60740
rect 47660 -61300 47680 -60760
rect 48080 -60920 48100 -60760
rect 48080 -60940 53800 -60920
rect 48080 -61140 53480 -60940
rect 53780 -61140 53800 -60940
rect 48080 -61160 53800 -61140
rect 48080 -61300 48100 -61160
rect 47660 -61320 48100 -61300
rect 57760 -62420 58280 -57140
rect 59600 -58800 65500 -58700
rect 59600 -59200 59700 -58800
rect 60400 -59200 65100 -58800
rect 65400 -59200 65500 -58800
rect 59600 -59300 65500 -59200
rect 57760 -62540 57800 -62420
rect 58240 -62540 58280 -62420
rect 14600 -65400 36000 -64800
rect 41000 -64600 41700 -64500
rect 41000 -65200 41100 -64600
rect 41600 -64700 56200 -64600
rect 41600 -65100 55500 -64700
rect 56100 -65100 56200 -64700
rect 41600 -65200 56200 -65100
rect 41000 -65300 41700 -65200
rect 51400 -65680 55800 -65600
rect 51400 -65700 55440 -65680
rect 51400 -65900 51500 -65700
rect 52500 -65900 55440 -65700
rect 51400 -65960 55440 -65900
rect 55720 -65960 55800 -65680
rect 51400 -66000 55800 -65960
rect 55360 -66040 55800 -66000
rect 47840 -66220 48100 -66200
rect 47840 -66660 47860 -66220
rect 48080 -66320 48100 -66220
rect 48080 -66340 53800 -66320
rect 48080 -66540 53480 -66340
rect 53780 -66540 53800 -66340
rect 48080 -66560 53800 -66540
rect 48080 -66660 48100 -66560
rect 47840 -66680 48100 -66660
rect 57760 -67820 58280 -62540
rect 59600 -64200 66500 -64100
rect 59600 -64600 59700 -64200
rect 60400 -64600 66100 -64200
rect 66400 -64600 66500 -64200
rect 59600 -64700 66500 -64600
rect 57760 -67940 57800 -67820
rect 58240 -67940 58280 -67820
rect 40100 -70000 40800 -69900
rect 40100 -70600 40200 -70000
rect 40700 -70100 56200 -70000
rect 40700 -70500 55500 -70100
rect 56100 -70500 56200 -70100
rect 40700 -70600 56200 -70500
rect 40100 -70700 40800 -70600
rect 51400 -71080 55800 -71000
rect 51400 -71100 55460 -71080
rect 51400 -71300 51500 -71100
rect 52500 -71300 55460 -71100
rect 51400 -71360 55460 -71300
rect 55720 -71360 55800 -71080
rect 51400 -71400 55800 -71360
rect 55380 -71440 55800 -71400
rect 47700 -71600 48100 -71580
rect 47700 -72060 47720 -71600
rect 48080 -71720 48100 -71600
rect 48080 -71740 53800 -71720
rect 48080 -71940 53480 -71740
rect 53780 -71940 53800 -71740
rect 48080 -71960 53800 -71940
rect 48080 -72060 48100 -71960
rect 47700 -72080 48100 -72060
rect 57760 -73220 58280 -67940
rect 59600 -69600 67500 -69500
rect 59600 -70000 59700 -69600
rect 60400 -70000 67100 -69600
rect 67400 -70000 67500 -69600
rect 59600 -70100 67500 -70000
rect 57760 -73340 57800 -73220
rect 58240 -73340 58280 -73220
rect 39200 -75400 39900 -75300
rect 39200 -76000 39300 -75400
rect 39800 -75500 56200 -75400
rect 39800 -75900 55500 -75500
rect 56100 -75900 56200 -75500
rect 39800 -76000 56200 -75900
rect 39200 -76100 39900 -76000
rect 51400 -76480 55800 -76400
rect 51400 -76500 55400 -76480
rect 51400 -76700 51500 -76500
rect 52500 -76700 55400 -76500
rect 51400 -76760 55400 -76700
rect 55720 -76760 55800 -76480
rect 51400 -76800 55800 -76760
rect 55320 -76840 55800 -76800
rect 47760 -76940 48100 -76920
rect 47760 -77500 47780 -76940
rect 48080 -77120 48100 -76940
rect 48080 -77140 53800 -77120
rect 48080 -77340 53480 -77140
rect 53780 -77340 53800 -77140
rect 48080 -77360 53800 -77340
rect 48080 -77500 48100 -77360
rect 47760 -77520 48100 -77500
rect 57760 -78620 58280 -73340
rect 59600 -75000 68400 -74900
rect 59600 -75400 59700 -75000
rect 60400 -75400 68000 -75000
rect 68300 -75400 68400 -75000
rect 59600 -75500 68400 -75400
rect 57760 -78740 57800 -78620
rect 58240 -78740 58280 -78620
rect 38200 -80800 38900 -80700
rect 38200 -81400 38300 -80800
rect 38800 -80900 56300 -80800
rect 38800 -81300 55500 -80900
rect 56200 -81300 56300 -80900
rect 38800 -81400 56300 -81300
rect 38200 -81500 38900 -81400
rect 51400 -81880 55800 -81800
rect 51400 -81900 55440 -81880
rect 51400 -82100 51500 -81900
rect 52500 -82100 55440 -81900
rect 51400 -82160 55440 -82100
rect 55720 -82160 55800 -81880
rect 51400 -82200 55800 -82160
rect 55360 -82240 55800 -82200
rect 47780 -82380 48100 -82360
rect 47780 -82860 47800 -82380
rect 48080 -82520 48100 -82380
rect 48080 -82540 53800 -82520
rect 48080 -82740 53480 -82540
rect 53780 -82740 53800 -82540
rect 48080 -82760 53800 -82740
rect 48080 -82860 48100 -82760
rect 47780 -82880 48100 -82860
rect 57760 -84020 58280 -78740
rect 59600 -80400 69400 -80300
rect 59600 -80800 59700 -80400
rect 60400 -80800 69000 -80400
rect 69300 -80800 69400 -80400
rect 59600 -80900 69400 -80800
rect 57760 -84140 57800 -84020
rect 58240 -84140 58280 -84020
rect 57790 -84145 58250 -84140
rect 59600 -85800 70400 -85700
rect 37100 -86200 37800 -86100
rect 59600 -86200 59700 -85800
rect 60400 -86200 70000 -85800
rect 70300 -86200 70400 -85800
rect 37100 -86700 37200 -86200
rect 37700 -86300 56200 -86200
rect 59600 -86300 70400 -86200
rect 37700 -86600 55500 -86300
rect 56100 -86600 56200 -86300
rect 37700 -86700 56200 -86600
rect 37100 -86800 37800 -86700
<< via3 >>
rect 10500 -2000 11000 -1500
rect 11600 -2000 12100 -1500
rect 12700 -2000 13200 -1500
rect 13800 -2000 14300 -1500
rect 10500 -3000 11000 -2500
rect 11600 -3000 12100 -2500
rect 12700 -3000 13200 -2500
rect 13800 -3000 14300 -2500
rect 10500 -4000 11000 -3500
rect 11600 -4000 12100 -3500
rect 12700 -4000 13200 -3500
rect 13800 -4000 14300 -3500
rect 10500 -5000 11000 -4500
rect 11600 -5000 12100 -4500
rect 12700 -5000 13200 -4500
rect 13800 -5000 14300 -4500
rect 38000 1400 41400 2800
rect 43000 1000 46400 2400
rect 37900 -3600 41500 -400
rect 43000 -1400 46400 0
rect 21000 -7400 22000 -6600
rect 27200 -13000 34400 -10600
rect 15000 -49000 24000 -38000
rect 72000 -35500 74000 -34100
<< metal4 >>
rect 35000 3000 69400 5000
rect 35000 2800 41600 3000
rect 35000 1400 38000 2800
rect 41400 1400 41600 2800
rect 35000 1200 41600 1400
rect 42800 2400 46600 2600
rect 10499 -1500 11001 -1499
rect 10499 -2000 10500 -1500
rect 11000 -2000 11001 -1500
rect 10499 -2001 11001 -2000
rect 11599 -1500 12101 -1499
rect 11599 -2000 11600 -1500
rect 12100 -2000 12101 -1500
rect 11599 -2001 12101 -2000
rect 12699 -1500 13201 -1499
rect 12699 -2000 12700 -1500
rect 13200 -2000 13201 -1500
rect 12699 -2001 13201 -2000
rect 13799 -1500 14301 -1499
rect 13799 -2000 13800 -1500
rect 14300 -2000 14301 -1500
rect 13799 -2001 14301 -2000
rect 10499 -2500 11001 -2499
rect 10499 -3000 10500 -2500
rect 11000 -3000 11001 -2500
rect 10499 -3001 11001 -3000
rect 11599 -2500 12101 -2499
rect 11599 -3000 11600 -2500
rect 12100 -3000 12101 -2500
rect 11599 -3001 12101 -3000
rect 12699 -2500 13201 -2499
rect 12699 -3000 12700 -2500
rect 13200 -3000 13201 -2500
rect 12699 -3001 13201 -3000
rect 13799 -2500 14301 -2499
rect 13799 -3000 13800 -2500
rect 14300 -3000 14301 -2500
rect 13799 -3001 14301 -3000
rect 10499 -3500 11001 -3499
rect 10499 -4000 10500 -3500
rect 11000 -4000 11001 -3500
rect 10499 -4001 11001 -4000
rect 11599 -3500 12101 -3499
rect 11599 -4000 11600 -3500
rect 12100 -4000 12101 -3500
rect 11599 -4001 12101 -4000
rect 12699 -3500 13201 -3499
rect 12699 -4000 12700 -3500
rect 13200 -4000 13201 -3500
rect 12699 -4001 13201 -4000
rect 13799 -3500 14301 -3499
rect 13799 -4000 13800 -3500
rect 14300 -4000 14301 -3500
rect 13799 -4001 14301 -4000
rect 10499 -4500 11001 -4499
rect 10499 -5000 10500 -4500
rect 11000 -5000 11001 -4500
rect 10499 -5001 11001 -5000
rect 11599 -4500 12101 -4499
rect 11599 -5000 11600 -4500
rect 12100 -5000 12101 -4500
rect 11599 -5001 12101 -5000
rect 12699 -4500 13201 -4499
rect 12699 -5000 12700 -4500
rect 13200 -5000 13201 -4500
rect 12699 -5001 13201 -5000
rect 13799 -4500 14301 -4499
rect 13799 -5000 13800 -4500
rect 14300 -5000 14301 -4500
rect 13799 -5001 14301 -5000
rect 35000 -6000 35600 1200
rect 42800 1000 43000 2400
rect 46400 1000 46600 2400
rect 42800 800 46600 1000
rect 42800 0 46600 200
rect 37800 -400 41600 -300
rect 37800 -3600 37900 -400
rect 41500 -2000 41600 -400
rect 42800 -1400 43000 0
rect 46400 -1400 46600 0
rect 42800 -1600 46600 -1400
rect 41500 -3600 56200 -2000
rect 20800 -6600 22200 -6400
rect 20800 -7400 21000 -6600
rect 22000 -7400 22200 -6600
rect 20800 -7600 22200 -7400
rect 37800 -10400 56200 -3600
rect 27000 -10600 56200 -10400
rect 27000 -13000 27200 -10600
rect 34400 -13000 56200 -10600
rect 27000 -13200 56200 -13000
rect 37800 -37000 56200 -13200
rect -33300 -38000 56200 -37000
rect -33300 -49000 15000 -38000
rect 24000 -49000 56200 -38000
rect -33300 -50000 56200 -49000
rect 37800 -86700 56200 -50000
rect 61820 -36800 69400 3000
rect 71900 -34100 74100 -34000
rect 71900 -35500 72000 -34100
rect 74000 -35500 74100 -34100
rect 71900 -35600 74100 -35500
rect 61820 -38000 80600 -36800
rect 61820 -54400 69400 -38000
rect 81400 -54400 91400 -52200
rect 61820 -56000 91400 -54400
rect 61820 -85940 69300 -56000
rect 53200 -86800 56200 -86700
<< via4 >>
rect 10500 -2000 11000 -1500
rect 11600 -2000 12100 -1500
rect 12700 -2000 13200 -1500
rect 13800 -2000 14300 -1500
rect 10500 -3000 11000 -2500
rect 11600 -3000 12100 -2500
rect 12700 -3000 13200 -2500
rect 13800 -3000 14300 -2500
rect 10500 -4000 11000 -3500
rect 11600 -4000 12100 -3500
rect 12700 -4000 13200 -3500
rect 13800 -4000 14300 -3500
rect 10500 -5000 11000 -4500
rect 11600 -5000 12100 -4500
rect 12700 -5000 13200 -4500
rect 13800 -5000 14300 -4500
rect 43000 1000 46400 2400
rect 43000 -1400 46400 0
rect 21000 -7400 22000 -6600
rect 72000 -35500 74000 -34100
<< metal5 >>
rect 42800 2400 65600 2600
rect 42800 1000 43000 2400
rect 46400 1000 65600 2400
rect 42800 800 65600 1000
rect 42800 0 46600 200
rect -30200 -1500 14400 -1100
rect -30200 -1800 10500 -1500
rect -30200 -2700 -29800 -1800
rect -23100 -2700 -22700 -1800
rect -16000 -2700 -15600 -1800
rect -8900 -2700 -8500 -1800
rect -1800 -2700 -1400 -1800
rect 5300 -1900 10500 -1800
rect 5300 -2700 5700 -1900
rect 10100 -2000 10500 -1900
rect 11000 -2000 11600 -1500
rect 12100 -2000 12700 -1500
rect 13200 -2000 13800 -1500
rect 14300 -2000 14400 -1500
rect 10100 -2500 14400 -2000
rect 10100 -3000 10500 -2500
rect 11000 -3000 11600 -2500
rect 12100 -3000 12700 -2500
rect 13200 -3000 13800 -2500
rect 14300 -3000 14400 -2500
rect 10100 -3500 14400 -3000
rect 10100 -4000 10500 -3500
rect 11000 -4000 11600 -3500
rect 12100 -4000 12700 -3500
rect 13200 -4000 13800 -3500
rect 14300 -4000 14400 -3500
rect 10100 -4500 14400 -4000
rect 10100 -5000 10500 -4500
rect 11000 -5000 11600 -4500
rect 12100 -5000 12700 -4500
rect 13200 -5000 13800 -4500
rect 14300 -5000 14400 -4500
rect 42800 -1400 43000 0
rect 46400 -1400 46600 0
rect 42800 -1500 46600 -1400
rect 42800 -4600 58900 -1500
rect 10476 -5024 11024 -5000
rect 11576 -5024 12124 -5000
rect 12676 -5024 13224 -5000
rect 13776 -5024 14324 -5000
rect 42800 -6400 53300 -4600
rect 20800 -6600 53300 -6400
rect 20800 -7400 21000 -6600
rect 22000 -6900 53300 -6600
rect 22000 -7400 58800 -6900
rect 20800 -7600 58800 -7400
rect 42700 -10000 58800 -7600
rect 42800 -12300 53300 -10000
rect 42800 -15400 58900 -12300
rect 42800 -17700 53300 -15400
rect 42800 -20800 58900 -17700
rect 42800 -23100 53300 -20800
rect 42800 -26200 58900 -23100
rect 42800 -28500 53300 -26200
rect 42800 -31600 58900 -28500
rect 42800 -33900 53300 -31600
rect 42800 -37000 58900 -33900
rect 63200 -34000 65600 800
rect 63200 -34100 89600 -34000
rect 63200 -35500 72000 -34100
rect 74000 -35500 89600 -34100
rect 63200 -35600 89600 -35500
rect 42800 -39300 53300 -37000
rect 42800 -42400 58900 -39300
rect 63200 -41000 65600 -35600
rect 79200 -38800 89600 -35600
rect 63200 -41792 69418 -41000
rect 72648 -41792 91400 -41000
rect 42800 -44700 53300 -42400
rect 63200 -42800 91400 -41792
rect 42800 -47800 58900 -44700
rect 63200 -45600 65600 -42800
rect 63200 -47400 91400 -45600
rect 42800 -50100 53300 -47800
rect 63200 -49600 65600 -47400
rect 42800 -53200 58900 -50100
rect 63200 -50492 69234 -49600
rect 73098 -50492 91400 -49600
rect 63200 -51400 91400 -50492
rect 42800 -55500 53300 -53200
rect 42800 -58600 58900 -55500
rect 42800 -60900 53300 -58600
rect 42800 -64000 58900 -60900
rect 42800 -66300 53300 -64000
rect 42800 -69400 58900 -66300
rect 42800 -71700 53300 -69400
rect 42800 -74800 58900 -71700
rect 42800 -77100 53300 -74800
rect 42800 -77520 58900 -77100
rect 42800 -78230 56224 -77520
rect 57194 -78230 58900 -77520
rect -30200 -79800 -29800 -78900
rect -23100 -79800 -22700 -78900
rect -16000 -79800 -15600 -78900
rect -8900 -79800 -8500 -78900
rect -1800 -79800 -1400 -78900
rect 5300 -79800 5700 -78900
rect -30200 -80200 5700 -79800
rect 42800 -79106 58900 -78230
rect 42800 -79798 56126 -79106
rect 57196 -79798 58900 -79106
rect 42800 -80200 58900 -79798
rect 42800 -82500 53300 -80200
rect 42800 -83000 58900 -82500
rect 42800 -83540 56342 -83000
rect 57110 -83540 58900 -83000
rect 42800 -84586 58900 -83540
rect 42800 -85078 56350 -84586
rect 57054 -85078 58900 -84586
rect 42800 -85600 58900 -85078
use 16to4_PriorityEncoder_v0p0p1  16to4_PriorityEncoder_v0p0p1_0 /foss/designs/Analog_FA23_SP24/PriorityEncoder/magic
timestamp 1717026683
transform 1 0 72130 0 1 -38130
box 470 -15870 20230 350
use frontAnalog_v0p0p1  frontAnalog_v0p0p1_0
timestamp 1717026683
transform 1 0 51936 0 1 -11930
box 1064 1130 10170 5492
use frontAnalog_v0p0p1  frontAnalog_v0p0p1_1
timestamp 1717026683
transform 1 0 51936 0 1 -44330
box 1064 1130 10170 5492
use frontAnalog_v0p0p1  frontAnalog_v0p0p1_2
timestamp 1717026683
transform 1 0 51936 0 1 -6530
box 1064 1130 10170 5492
use frontAnalog_v0p0p1  frontAnalog_v0p0p1_3
timestamp 1717026683
transform 1 0 51936 0 1 -17330
box 1064 1130 10170 5492
use frontAnalog_v0p0p1  frontAnalog_v0p0p1_4
timestamp 1717026683
transform 1 0 51936 0 1 -22730
box 1064 1130 10170 5492
use frontAnalog_v0p0p1  frontAnalog_v0p0p1_5
timestamp 1717026683
transform 1 0 51936 0 1 -28130
box 1064 1130 10170 5492
use frontAnalog_v0p0p1  frontAnalog_v0p0p1_6
timestamp 1717026683
transform 1 0 51936 0 1 -33530
box 1064 1130 10170 5492
use frontAnalog_v0p0p1  frontAnalog_v0p0p1_7
timestamp 1717026683
transform 1 0 51936 0 1 -38930
box 1064 1130 10170 5492
use frontAnalog_v0p0p1  frontAnalog_v0p0p1_8
timestamp 1717026683
transform 1 0 51936 0 1 -49730
box 1064 1130 10170 5492
use frontAnalog_v0p0p1  frontAnalog_v0p0p1_9
timestamp 1717026683
transform 1 0 51936 0 1 -55130
box 1064 1130 10170 5492
use frontAnalog_v0p0p1  frontAnalog_v0p0p1_10
timestamp 1717026683
transform 1 0 51936 0 1 -60530
box 1064 1130 10170 5492
use frontAnalog_v0p0p1  frontAnalog_v0p0p1_11
timestamp 1717026683
transform 1 0 51936 0 1 -65930
box 1064 1130 10170 5492
use frontAnalog_v0p0p1  frontAnalog_v0p0p1_12
timestamp 1717026683
transform 1 0 51936 0 1 -76730
box 1064 1130 10170 5492
use frontAnalog_v0p0p1  frontAnalog_v0p0p1_13
timestamp 1717026683
transform 1 0 51936 0 1 -71330
box 1064 1130 10170 5492
use frontAnalog_v0p0p1  frontAnalog_v0p0p1_14
timestamp 1717026683
transform 1 0 51936 0 1 -82130
box 1064 1130 10170 5492
use frontAnalog_v0p0p1  frontAnalog_v0p0p1_15
timestamp 1717026683
transform 1 0 51936 0 1 -87530
box 1064 1130 10170 5492
use PTAT_v0p0p0_mag  PTAT_v0p0p0_mag_0 /foss/designs/Analog_FA23_SP24/PTAT/magic
timestamp 1716869746
transform 1 0 18930 0 1 -12102
box -2530 -4098 15822 4693
use resistorDivider_v0p0p1  resistorDivider_v0p0p1_0
timestamp 1716869746
transform 1 0 40840 0 1 -44680
box -16460 -14720 -4458 14560
use sky130_fd_pr__cap_mim_m3_2_U5PCTN  sky130_fd_pr__cap_mim_m3_2_U5PCTN_0
timestamp 1716869746
transform 1 0 -12006 0 1 -40800
box -21094 -38400 21116 38400
<< labels >>
flabel metal1 12400 -29200 12600 -29000 0 FreeSans 256 0 0 0 VFS
port 0 nsew
flabel metal1 12400 -62800 12600 -62600 0 FreeSans 256 0 0 0 VL
port 9 nsew
flabel metal1 39700 600 39900 800 0 FreeSans 256 0 0 0 GND
port 8 nsew
flabel metal1 44600 400 44800 600 0 FreeSans 256 0 0 0 VDD
port 5 nsew
flabel metal1 52000 1100 52200 1300 0 FreeSans 256 0 0 0 VIN
port 6 nsew
flabel metal1 94000 -39800 94200 -39600 0 FreeSans 256 0 0 0 OUT3
port 1 nsew
flabel metal1 93800 -44400 94000 -44200 0 FreeSans 256 0 0 0 OUT2
port 2 nsew
flabel metal1 93800 -48400 94000 -48200 0 FreeSans 256 0 0 0 OUT1
port 3 nsew
flabel metal1 93800 -52200 94000 -52000 0 FreeSans 256 0 0 0 OUT0
port 4 nsew
flabel metal1 57920 1100 58120 1300 0 FreeSans 256 0 0 0 CLK
port 7 nsew
rlabel metal3 37700 -86700 55500 -86200 1 VV1
port 10 n
rlabel metal3 38800 -81400 55500 -80800 1 VV2
port 11 n
rlabel metal3 39800 -76000 55500 -75400 1 VV3
port 12 n
rlabel metal3 40700 -70600 55500 -70000 1 VV4
port 13 n
rlabel metal3 41600 -65200 55500 -64600 1 VV5
port 14 n
rlabel metal3 42500 -59800 55500 -59200 1 VV6
port 15 n
rlabel metal3 43400 -54400 55400 -53800 1 VV7
port 16 n
rlabel metal3 44300 -49000 55500 -48400 1 VV8
port 17 n
rlabel metal3 44300 -43600 55500 -43000 1 VV9
port 18 n
rlabel metal3 43100 -38200 55400 -37600 1 VV10
port 19 n
rlabel metal3 42100 -32800 55500 -32200 1 VV11
port 20 n
rlabel metal3 41000 -27400 55500 -26800 1 VV12
port 21 n
rlabel metal3 40000 -22000 55500 -21400 1 VV13
port 22 n
rlabel metal3 39000 -16600 55500 -16000 1 VV14
port 23 n
rlabel metal3 38100 -11200 55500 -10600 1 VV15
port 24 n
rlabel metal3 37000 -5700 55600 -5200 1 VV16
port 25 n
rlabel metal1 56374 -85082 57010 -84958 1 R0
port 26 n
flabel metal1 56592 -83258 57024 -83024 0 FreeSans 192 0 0 0 S0
port 27 n
rlabel metal1 56362 -79722 57006 -79558 1 R1
port 28 n
rlabel metal1 56580 -77892 57066 -77610 1 S1
port 29 n
rlabel metal3 68600 -39240 73080 -39060 1 I15
port 30 n
rlabel metal3 67400 -39740 73200 -39560 1 I14
port 31 n
rlabel metal3 66600 -40020 72399 -39839 1 I13
port 32 n
rlabel metal3 65400 -40480 73200 -40300 1 I12
port 33 n
rlabel metal3 64160 -40840 73200 -40660 1 I11
port 34 n
rlabel metal3 63300 -41300 73200 -41000 1 I10
port 35 n
rlabel metal3 62500 -41700 73100 -41500 1 I9
port 36 n
rlabel metal3 60400 -43600 73200 -42600 1 I8
port 37 n
rlabel metal3 63203 -47499 73103 -47199 1 I7
port 38 n
rlabel metal3 64500 -47900 73100 -47600 1 I6
port 39 n
rlabel metal3 65400 -48300 73100 -48000 1 I5
port 40 n
rlabel metal3 66400 -48700 73100 -48400 1 I4
port 41 n
rlabel metal3 67400 -49100 73100 -48800 1 I3
port 42 n
rlabel metal3 68300 -49500 73100 -49200 1 I2
port 43 n
rlabel metal3 69300 -49900 73100 -49600 1 I1
port 44 n
rlabel metal3 70300 -50300 73100 -50000 1 I0
port 45 n
rlabel metal3 31328 -9838 32878 -8600 1 IB
port 46 n
<< end >>
