magic
tech sky130A
magscale 1 2
timestamp 1709401415
<< error_p >>
rect -77 2081 -19 2087
rect 115 2081 173 2087
rect -77 2047 -65 2081
rect 115 2047 127 2081
rect -77 2041 -19 2047
rect 115 2041 173 2047
rect -173 -2047 -115 -2041
rect 19 -2047 77 -2041
rect -173 -2081 -161 -2047
rect 19 -2081 31 -2047
rect -173 -2087 -115 -2081
rect 19 -2087 77 -2081
<< nwell >>
rect -359 -2219 359 2219
<< pmos >>
rect -159 -2000 -129 2000
rect -63 -2000 -33 2000
rect 33 -2000 63 2000
rect 129 -2000 159 2000
<< pdiff >>
rect -221 1988 -159 2000
rect -221 -1988 -209 1988
rect -175 -1988 -159 1988
rect -221 -2000 -159 -1988
rect -129 1988 -63 2000
rect -129 -1988 -113 1988
rect -79 -1988 -63 1988
rect -129 -2000 -63 -1988
rect -33 1988 33 2000
rect -33 -1988 -17 1988
rect 17 -1988 33 1988
rect -33 -2000 33 -1988
rect 63 1988 129 2000
rect 63 -1988 79 1988
rect 113 -1988 129 1988
rect 63 -2000 129 -1988
rect 159 1988 221 2000
rect 159 -1988 175 1988
rect 209 -1988 221 1988
rect 159 -2000 221 -1988
<< pdiffc >>
rect -209 -1988 -175 1988
rect -113 -1988 -79 1988
rect -17 -1988 17 1988
rect 79 -1988 113 1988
rect 175 -1988 209 1988
<< nsubdiff >>
rect -323 2149 -227 2183
rect 227 2149 323 2183
rect -323 2087 -289 2149
rect 289 2087 323 2149
rect -323 -2149 -289 -2087
rect 289 -2149 323 -2087
rect -323 -2183 -227 -2149
rect 227 -2183 323 -2149
<< nsubdiffcont >>
rect -227 2149 227 2183
rect -323 -2087 -289 2087
rect 289 -2087 323 2087
rect -227 -2183 227 -2149
<< poly >>
rect -81 2081 -15 2097
rect -81 2047 -65 2081
rect -31 2047 -15 2081
rect -81 2031 -15 2047
rect 111 2081 177 2097
rect 111 2047 127 2081
rect 161 2047 177 2081
rect 111 2031 177 2047
rect -159 2000 -129 2026
rect -63 2000 -33 2031
rect 33 2000 63 2026
rect 129 2000 159 2031
rect -159 -2031 -129 -2000
rect -63 -2026 -33 -2000
rect 33 -2031 63 -2000
rect 129 -2026 159 -2000
rect -177 -2047 -111 -2031
rect -177 -2081 -161 -2047
rect -127 -2081 -111 -2047
rect -177 -2097 -111 -2081
rect 15 -2047 81 -2031
rect 15 -2081 31 -2047
rect 65 -2081 81 -2047
rect 15 -2097 81 -2081
<< polycont >>
rect -65 2047 -31 2081
rect 127 2047 161 2081
rect -161 -2081 -127 -2047
rect 31 -2081 65 -2047
<< locali >>
rect -323 2149 -227 2183
rect 227 2149 323 2183
rect -323 2087 -289 2149
rect 289 2087 323 2149
rect -81 2047 -65 2081
rect -31 2047 -15 2081
rect 111 2047 127 2081
rect 161 2047 177 2081
rect -209 1988 -175 2004
rect -209 -2004 -175 -1988
rect -113 1988 -79 2004
rect -113 -2004 -79 -1988
rect -17 1988 17 2004
rect -17 -2004 17 -1988
rect 79 1988 113 2004
rect 79 -2004 113 -1988
rect 175 1988 209 2004
rect 175 -2004 209 -1988
rect -177 -2081 -161 -2047
rect -127 -2081 -111 -2047
rect 15 -2081 31 -2047
rect 65 -2081 81 -2047
rect -323 -2149 -289 -2087
rect 289 -2149 323 -2087
rect -323 -2183 -227 -2149
rect 227 -2183 323 -2149
<< viali >>
rect -65 2047 -31 2081
rect 127 2047 161 2081
rect -209 -1988 -175 1988
rect -113 -1988 -79 1988
rect -17 -1988 17 1988
rect 79 -1988 113 1988
rect 175 -1988 209 1988
rect -161 -2081 -127 -2047
rect 31 -2081 65 -2047
<< metal1 >>
rect -77 2081 -19 2087
rect -77 2047 -65 2081
rect -31 2047 -19 2081
rect -77 2041 -19 2047
rect 115 2081 173 2087
rect 115 2047 127 2081
rect 161 2047 173 2081
rect 115 2041 173 2047
rect -215 1988 -169 2000
rect -215 -1988 -209 1988
rect -175 -1988 -169 1988
rect -215 -2000 -169 -1988
rect -119 1988 -73 2000
rect -119 -1988 -113 1988
rect -79 -1988 -73 1988
rect -119 -2000 -73 -1988
rect -23 1988 23 2000
rect -23 -1988 -17 1988
rect 17 -1988 23 1988
rect -23 -2000 23 -1988
rect 73 1988 119 2000
rect 73 -1988 79 1988
rect 113 -1988 119 1988
rect 73 -2000 119 -1988
rect 169 1988 215 2000
rect 169 -1988 175 1988
rect 209 -1988 215 1988
rect 169 -2000 215 -1988
rect -173 -2047 -115 -2041
rect -173 -2081 -161 -2047
rect -127 -2081 -115 -2047
rect -173 -2087 -115 -2081
rect 19 -2047 77 -2041
rect 19 -2081 31 -2047
rect 65 -2081 77 -2047
rect 19 -2087 77 -2081
<< properties >>
string FIXED_BBOX -306 -2166 306 2166
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 20 l 0.15 m 1 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
