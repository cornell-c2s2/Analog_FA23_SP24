magic
tech sky130A
magscale 1 2
timestamp 1709331665
<< metal1 >>
rect 8186 21652 8254 21700
rect 8186 21156 8256 21200
<< metal3 >>
rect 16562 22792 16872 22830
rect 16562 22648 16605 22792
rect 16829 22648 16872 22792
rect 16562 22610 16872 22648
rect 12832 17812 12986 17848
rect 12832 17748 12877 17812
rect 12941 17748 12986 17812
rect 12832 17712 12986 17748
rect 14600 16290 15536 19122
rect 14464 16238 15536 16290
rect 12894 15700 15536 16238
rect 14464 15642 15536 15700
rect 14464 15612 14854 15642
<< via3 >>
rect 16605 22648 16829 22792
rect 12877 17748 12941 17812
<< metal4 >>
rect 4330 25118 4480 25216
rect 16486 22792 16892 22854
rect 16486 22648 16605 22792
rect 16829 22648 16892 22792
rect 16486 17880 16892 22648
rect 12826 17812 16892 17880
rect 12826 17748 12877 17812
rect 12941 17748 16892 17812
rect 12826 17696 16892 17748
rect 16486 17486 16892 17696
use OTA_MULT_GM  OTA_MULT_GM_0
timestamp 1709331665
transform 1 0 10034 0 1 14648
box -10034 -14658 10202 17116
<< labels >>
rlabel metal4 s 16578 19274 16830 19502 4 VDD
port 1 nsew
rlabel metal4 s 4330 25118 4480 25216 4 Vout
port 2 nsew
rlabel metal3 s 14942 15832 15170 16212 4 VSS
port 3 nsew
rlabel metal1 s 8186 21652 8254 21700 4 Vp
port 4 nsew
rlabel metal1 s 8186 21156 8256 21200 4 Vn
port 5 nsew
<< end >>
