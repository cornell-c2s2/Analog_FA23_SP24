magic
tech sky130A
magscale 1 2
timestamp 1713142632
<< pwell >>
rect -1360 -14759 1360 14759
<< psubdiff >>
rect -1324 14689 -1228 14723
rect 1228 14689 1324 14723
rect -1324 14627 -1290 14689
rect 1290 14627 1324 14689
rect -1324 -14689 -1290 -14627
rect 1290 -14689 1324 -14627
rect -1324 -14723 -1228 -14689
rect 1228 -14723 1324 -14689
<< psubdiffcont >>
rect -1228 14689 1228 14723
rect -1324 -14627 -1290 14627
rect 1290 -14627 1324 14627
rect -1228 -14723 1228 -14689
<< xpolycontact >>
rect -1194 -14593 -48 -14161
rect 48 -14593 1194 -14161
<< xpolyres >>
rect -1194 13447 1194 14593
rect -1194 -14161 -48 13447
rect 48 -14161 1194 13447
<< locali >>
rect -1324 14689 -1228 14723
rect 1228 14689 1324 14723
rect -1324 14627 -1290 14689
rect 1290 14627 1324 14689
rect -1324 -14689 -1290 -14627
rect 1290 -14689 1324 -14627
rect -1324 -14723 -1228 -14689
rect 1228 -14723 1324 -14689
<< properties >>
string FIXED_BBOX -1307 -14706 1307 14706
string gencell sky130_fd_pr__res_xhigh_po_5p73
string library sky130
string parameters w 5.73 l 143.25 m 1 nx 2 wmin 5.730 lmin 0.50 rho 2000 val 102.065k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 5.730 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 1 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
