magic
tech sky130A
timestamp 1716868724
<< end >>
