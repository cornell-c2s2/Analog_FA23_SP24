magic
tech sky130A
magscale 1 2
timestamp 1714790421
<< pwell >>
rect -5086 -869 5086 869
<< psubdiff >>
rect -5050 799 -4954 833
rect 4954 799 5050 833
rect -5050 737 -5016 799
rect 5016 737 5050 799
rect -5050 -799 -5016 -737
rect 5016 -799 5050 -737
rect -5050 -833 -4954 -799
rect 4954 -833 5050 -799
<< psubdiffcont >>
rect -4954 799 4954 833
rect -5050 -737 -5016 737
rect 5016 -737 5050 737
rect -4954 -833 4954 -799
<< xpolycontact >>
rect -4920 271 -3774 703
rect -4920 -703 -3774 -271
rect -3678 271 -2532 703
rect -3678 -703 -2532 -271
rect -2436 271 -1290 703
rect -2436 -703 -1290 -271
rect -1194 271 -48 703
rect -1194 -703 -48 -271
rect 48 271 1194 703
rect 48 -703 1194 -271
rect 1290 271 2436 703
rect 1290 -703 2436 -271
rect 2532 271 3678 703
rect 2532 -703 3678 -271
rect 3774 271 4920 703
rect 3774 -703 4920 -271
<< xpolyres >>
rect -4920 -271 -3774 271
rect -3678 -271 -2532 271
rect -2436 -271 -1290 271
rect -1194 -271 -48 271
rect 48 -271 1194 271
rect 1290 -271 2436 271
rect 2532 -271 3678 271
rect 3774 -271 4920 271
<< locali >>
rect -5050 799 -4954 833
rect 4954 799 5050 833
rect -5050 737 -5016 799
rect 5016 737 5050 799
rect -5050 -799 -5016 -737
rect 5016 -799 5050 -737
rect -5050 -833 -4954 -799
rect 4954 -833 5050 -799
<< viali >>
rect -4904 288 -3790 685
rect -3662 288 -2548 685
rect -2420 288 -1306 685
rect -1178 288 -64 685
rect 64 288 1178 685
rect 1306 288 2420 685
rect 2548 288 3662 685
rect 3790 288 4904 685
rect -4904 -685 -3790 -288
rect -3662 -685 -2548 -288
rect -2420 -685 -1306 -288
rect -1178 -685 -64 -288
rect 64 -685 1178 -288
rect 1306 -685 2420 -288
rect 2548 -685 3662 -288
rect 3790 -685 4904 -288
<< metal1 >>
rect -4916 685 -3778 691
rect -4916 288 -4904 685
rect -3790 288 -3778 685
rect -4916 282 -3778 288
rect -3674 685 -2536 691
rect -3674 288 -3662 685
rect -2548 288 -2536 685
rect -3674 282 -2536 288
rect -2432 685 -1294 691
rect -2432 288 -2420 685
rect -1306 288 -1294 685
rect -2432 282 -1294 288
rect -1190 685 -52 691
rect -1190 288 -1178 685
rect -64 288 -52 685
rect -1190 282 -52 288
rect 52 685 1190 691
rect 52 288 64 685
rect 1178 288 1190 685
rect 52 282 1190 288
rect 1294 685 2432 691
rect 1294 288 1306 685
rect 2420 288 2432 685
rect 1294 282 2432 288
rect 2536 685 3674 691
rect 2536 288 2548 685
rect 3662 288 3674 685
rect 2536 282 3674 288
rect 3778 685 4916 691
rect 3778 288 3790 685
rect 4904 288 4916 685
rect 3778 282 4916 288
rect -4916 -288 -3778 -282
rect -4916 -685 -4904 -288
rect -3790 -685 -3778 -288
rect -4916 -691 -3778 -685
rect -3674 -288 -2536 -282
rect -3674 -685 -3662 -288
rect -2548 -685 -2536 -288
rect -3674 -691 -2536 -685
rect -2432 -288 -1294 -282
rect -2432 -685 -2420 -288
rect -1306 -685 -1294 -288
rect -2432 -691 -1294 -685
rect -1190 -288 -52 -282
rect -1190 -685 -1178 -288
rect -64 -685 -52 -288
rect -1190 -691 -52 -685
rect 52 -288 1190 -282
rect 52 -685 64 -288
rect 1178 -685 1190 -288
rect 52 -691 1190 -685
rect 1294 -288 2432 -282
rect 1294 -685 1306 -288
rect 2420 -685 2432 -288
rect 1294 -691 2432 -685
rect 2536 -288 3674 -282
rect 2536 -685 2548 -288
rect 3662 -685 3674 -288
rect 2536 -691 3674 -685
rect 3778 -288 4916 -282
rect 3778 -685 3790 -288
rect 4904 -685 4916 -288
rect 3778 -691 4916 -685
<< properties >>
string FIXED_BBOX -5033 -816 5033 816
string gencell sky130_fd_pr__res_xhigh_po_5p73
string library sky130
string parameters w 5.730 l 2.865 m 1 nx 8 wmin 5.730 lmin 0.50 rho 2000 val 1.065k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 5.730 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
