magic
tech sky130A
magscale 1 2
timestamp 1715635929
<< nwell >>
rect 1270 -630 1560 -620
rect 1258 -651 1560 -630
rect 1260 -1233 1560 -652
rect 1258 -1260 1560 -1233
rect 1880 -630 2170 -620
rect 1880 -1260 2182 -630
<< pwell >>
rect 1090 -620 2340 -480
rect 1090 -630 1270 -620
rect 1090 -1260 1258 -630
rect 1560 -1260 1880 -620
rect 2170 -630 2340 -620
rect 2182 -1260 2340 -630
rect 1090 -1320 2340 -1260
rect 1090 -1390 1260 -1320
rect 1740 -1330 1750 -1320
rect 2170 -1390 2340 -1320
rect 1090 -1426 1296 -1390
rect 2142 -1426 2340 -1390
<< psubdiff >>
rect 1150 -560 2290 -520
rect 1150 -1356 1190 -560
rect 1700 -660 1740 -560
rect 1150 -1360 1296 -1356
rect 1700 -1360 1740 -1100
rect 2250 -1356 2290 -560
rect 1150 -1380 1330 -1360
rect 1150 -1390 1296 -1380
rect 2142 -1390 2290 -1356
<< psubdiffcont >>
rect 1700 -1100 1740 -660
<< locali >>
rect 2820 -180 3050 -170
rect 530 -300 610 -220
rect 2820 -240 2890 -180
rect 3040 -240 3050 -180
rect 2820 -250 3050 -240
rect 540 -550 590 -300
rect 1670 -450 1770 -430
rect 1670 -520 1680 -450
rect 1760 -520 1770 -450
rect 1150 -560 2290 -520
rect 2840 -540 2900 -250
rect 1150 -1356 1190 -560
rect 1670 -660 1770 -560
rect 1670 -1100 1700 -660
rect 1740 -1100 1770 -660
rect 1670 -1150 1770 -1100
rect 1670 -1230 1680 -1150
rect 1760 -1230 1770 -1150
rect 1150 -1360 1296 -1356
rect 1150 -1380 1330 -1360
rect 1150 -1390 1296 -1380
rect 1670 -1430 1770 -1230
rect 2250 -1356 2290 -560
rect 2142 -1390 2290 -1356
<< viali >>
rect 1150 20 1780 90
rect 360 -300 530 -220
rect 2890 -240 3040 -180
rect 1680 -520 1760 -450
rect 1680 -1230 1760 -1150
rect 140 -2110 230 -1410
rect 3380 -940 3440 -790
rect 3220 -2110 3340 -1420
rect 800 -2930 2150 -2860
<< metal1 >>
rect 1610 760 1820 800
rect 900 490 1100 740
rect 1610 640 1650 760
rect 1780 640 1820 760
rect 1610 600 1820 640
rect 360 130 610 490
rect 900 400 1470 490
rect 890 330 900 400
rect 1030 350 1470 400
rect 1030 330 2110 350
rect 1320 300 2110 330
rect 1210 220 1220 290
rect 1280 220 1290 290
rect 2150 220 2160 290
rect 2220 220 2230 290
rect 1320 180 2110 210
rect 2390 180 2590 740
rect 1320 150 2400 180
rect 360 -70 390 130
rect 600 40 610 130
rect 1930 120 2400 150
rect 2520 120 2590 180
rect 2830 130 3090 170
rect 1138 90 1792 96
rect 1138 40 1150 90
rect 600 20 1150 40
rect 1780 40 1792 90
rect 2830 40 2840 130
rect 1780 20 2840 40
rect 600 -70 2840 20
rect 360 -90 2840 -70
rect 3040 -90 3090 130
rect 360 -140 3090 -90
rect 780 -200 2660 -140
rect 348 -220 542 -214
rect 348 -300 360 -220
rect 530 -300 542 -220
rect 780 -260 1560 -200
rect 1870 -260 2660 -200
rect 2878 -180 3052 -174
rect 2878 -240 2890 -180
rect 3040 -240 3052 -180
rect 2878 -246 3052 -240
rect 348 -306 542 -300
rect 640 -380 650 -290
rect 730 -380 740 -290
rect 1600 -380 1670 -290
rect 1760 -380 1840 -290
rect 2700 -380 2710 -290
rect 2790 -380 2800 -290
rect 760 -450 1560 -410
rect 1880 -440 2670 -410
rect 3830 -430 4030 -350
rect 1668 -450 1772 -444
rect 1870 -450 2670 -440
rect 760 -480 1590 -450
rect -330 -540 -130 -480
rect -330 -630 1440 -540
rect -330 -680 1170 -630
rect 1160 -720 1170 -680
rect 1270 -720 1440 -630
rect 440 -830 450 -740
rect 520 -750 1060 -740
rect 1530 -750 1590 -480
rect 1668 -520 1680 -450
rect 1760 -520 1772 -450
rect 1668 -526 1772 -520
rect 1840 -480 2670 -450
rect 520 -820 880 -750
rect 520 -830 590 -820
rect 870 -830 880 -820
rect 1050 -830 1060 -750
rect 1510 -760 1590 -750
rect 870 -850 1060 -830
rect 880 -860 1060 -850
rect 1480 -810 1590 -760
rect 1840 -750 1910 -480
rect 2900 -550 4030 -430
rect 2900 -580 3010 -550
rect 2180 -630 3010 -580
rect 2160 -640 2170 -630
rect 2000 -720 2170 -640
rect 2270 -690 3010 -630
rect 2270 -720 2280 -690
rect 3200 -730 3210 -650
rect 3300 -730 3310 -650
rect 1840 -760 1930 -750
rect 2380 -760 2880 -750
rect 1840 -810 1960 -760
rect 550 -970 560 -870
rect 630 -880 640 -870
rect 880 -880 1020 -860
rect 630 -940 840 -880
rect 630 -970 650 -940
rect 600 -1270 650 -970
rect 880 -1030 890 -940
rect 1060 -1030 1070 -940
rect 1480 -1060 1560 -810
rect 1870 -1060 1960 -810
rect 2380 -850 2390 -760
rect 2560 -850 2880 -760
rect 2970 -850 2990 -750
rect 2380 -870 2570 -850
rect 3150 -880 3220 -780
rect 3374 -790 3446 -778
rect 2600 -890 2840 -889
rect 2600 -949 2790 -890
rect 2370 -1040 2380 -950
rect 2550 -1040 2560 -950
rect 2780 -1020 2790 -949
rect 2850 -1020 2860 -890
rect 3050 -930 3220 -880
rect 1480 -1120 1570 -1060
rect 1640 -1120 1650 -1060
rect 1800 -1130 1960 -1060
rect 1668 -1150 1772 -1144
rect 1160 -1260 1170 -1170
rect 1270 -1250 1440 -1170
rect 1668 -1230 1680 -1150
rect 1760 -1230 1772 -1150
rect 1668 -1236 1772 -1230
rect 1270 -1260 1280 -1250
rect 350 -1340 650 -1270
rect 700 -1340 710 -1270
rect 800 -1340 810 -1270
rect 1800 -1300 1880 -1130
rect 2000 -1240 2170 -1170
rect 2160 -1260 2170 -1240
rect 2270 -1260 2280 -1170
rect 2790 -1279 2840 -1020
rect 3040 -1040 3050 -930
rect 3160 -970 3220 -930
rect 3280 -940 3360 -790
rect 3500 -940 3510 -790
rect 3280 -960 3510 -940
rect 3160 -980 3210 -970
rect 3160 -1040 3170 -980
rect -70 -1380 230 -1370
rect 600 -1380 650 -1340
rect 1340 -1360 1880 -1300
rect 2020 -1340 2030 -1280
rect 2100 -1340 2110 -1280
rect 2040 -1350 2110 -1340
rect 2620 -1350 2630 -1280
rect 2730 -1350 2740 -1280
rect 2790 -1349 3090 -1279
rect -70 -1400 330 -1380
rect 600 -1390 670 -1380
rect -70 -2110 -30 -1400
rect 210 -1410 330 -1400
rect 470 -1410 560 -1400
rect 230 -2110 330 -1410
rect -70 -2170 330 -2110
rect 430 -1510 470 -1410
rect 540 -1420 560 -1410
rect 550 -1510 560 -1420
rect 430 -1520 550 -1510
rect 430 -2170 520 -1520
rect 100 -2180 330 -2170
rect 600 -2180 680 -1390
rect 790 -1750 860 -1390
rect 1340 -1530 1400 -1360
rect 1460 -1420 1580 -1410
rect 1460 -1490 1470 -1420
rect 1560 -1490 1580 -1420
rect 1860 -1420 1980 -1410
rect 1860 -1490 1880 -1420
rect 1960 -1490 1980 -1420
rect 1860 -1500 1980 -1490
rect 2040 -1530 2100 -1350
rect 2790 -1380 2840 -1349
rect 2750 -1390 2840 -1380
rect 1340 -1540 1410 -1530
rect 2030 -1540 2100 -1530
rect 1340 -1550 1440 -1540
rect 1360 -1750 1440 -1550
rect 790 -1940 1440 -1750
rect 790 -2170 860 -1940
rect 600 -2210 670 -2180
rect 600 -2220 640 -2210
rect 350 -2290 640 -2220
rect 710 -2240 850 -2230
rect 710 -2310 730 -2240
rect 830 -2310 850 -2240
rect 710 -2320 850 -2310
rect 1360 -2320 1440 -1940
rect 1590 -2320 1850 -1540
rect 2000 -1550 2100 -1540
rect 2000 -1750 2080 -1550
rect 2580 -1750 2650 -1400
rect 2000 -1940 2650 -1750
rect 2000 -2320 2080 -1940
rect 2580 -2180 2650 -1940
rect 2740 -1402 2840 -1390
rect 2740 -2178 2746 -1402
rect 2760 -2178 2840 -1402
rect 2890 -1410 3010 -1400
rect 2890 -1520 2900 -1410
rect 2990 -1520 3010 -1410
rect 3110 -1410 3620 -1380
rect 3110 -1420 3320 -1410
rect 2890 -1530 3014 -1520
rect 2740 -2190 2840 -2178
rect 2920 -2180 3014 -1530
rect 3110 -2110 3220 -1420
rect 3110 -2120 3320 -2110
rect 3580 -2120 3620 -1410
rect 3110 -2160 3620 -2120
rect 3110 -2170 3340 -2160
rect 2770 -2219 2840 -2190
rect 2800 -2229 2840 -2219
rect 2600 -2250 2740 -2240
rect 2600 -2310 2640 -2250
rect 2720 -2310 2740 -2250
rect 2800 -2299 3090 -2229
rect 2600 -2320 2740 -2310
rect 1660 -2340 1770 -2320
rect 1150 -2400 1160 -2340
rect 1270 -2360 1280 -2340
rect 1270 -2400 1580 -2360
rect 1150 -2420 1580 -2400
rect 150 -2620 720 -2460
rect 1670 -2500 1760 -2340
rect 2160 -2360 2170 -2340
rect 1860 -2410 2170 -2360
rect 2280 -2410 2290 -2340
rect 1860 -2430 2290 -2410
rect 820 -2580 2620 -2500
rect 820 -2620 1600 -2580
rect 1840 -2620 2620 -2580
rect 150 -2740 490 -2620
rect 600 -2630 720 -2620
rect 600 -2740 770 -2630
rect 150 -2750 770 -2740
rect 1650 -2750 1790 -2630
rect 2670 -2750 2760 -2630
rect 2880 -2750 2890 -2630
rect 590 -2860 2620 -2780
rect 590 -2930 800 -2860
rect 2150 -2930 2620 -2860
rect 590 -3010 2620 -2930
rect 590 -3210 790 -3010
rect 2540 -3210 2620 -3010
rect 590 -3258 2620 -3210
rect 652 -3260 2620 -3258
<< via1 >>
rect 1650 640 1780 760
rect 900 330 1030 400
rect 1220 220 1280 290
rect 2160 220 2220 290
rect 390 -70 600 130
rect 2400 120 2520 180
rect 2840 -90 3040 130
rect 370 -300 520 -220
rect 2890 -240 3040 -180
rect 650 -380 730 -290
rect 1670 -380 1760 -290
rect 2710 -380 2790 -290
rect 1170 -720 1270 -630
rect 450 -830 520 -740
rect 1680 -520 1760 -450
rect 880 -830 1050 -750
rect 2170 -720 2270 -630
rect 3210 -730 3300 -650
rect 560 -970 630 -870
rect 890 -1030 1060 -940
rect 2390 -850 2560 -760
rect 2880 -850 2970 -750
rect 2380 -1040 2550 -950
rect 2790 -1020 2850 -890
rect 1570 -1120 1640 -1060
rect 1170 -1260 1270 -1170
rect 1680 -1230 1760 -1150
rect 710 -1340 800 -1270
rect 2170 -1260 2270 -1170
rect 3050 -1040 3160 -930
rect 3360 -940 3380 -790
rect 3380 -940 3440 -790
rect 3440 -940 3500 -790
rect 2030 -1340 2100 -1280
rect 2630 -1350 2730 -1280
rect -30 -1410 210 -1400
rect -30 -2110 140 -1410
rect 140 -2110 210 -1410
rect 470 -1420 540 -1410
rect 470 -1510 550 -1420
rect 1470 -1490 1560 -1420
rect 1880 -1490 1960 -1420
rect 730 -2310 830 -2240
rect 2900 -1520 2990 -1410
rect 3320 -1420 3580 -1410
rect 3320 -2110 3340 -1420
rect 3340 -2110 3580 -1420
rect 3320 -2120 3580 -2110
rect 2640 -2310 2720 -2250
rect 1160 -2400 1270 -2340
rect 2170 -2410 2280 -2340
rect 490 -2740 600 -2620
rect 2760 -2750 2880 -2630
rect 790 -3210 2540 -3010
<< metal2 >>
rect 1650 760 1780 780
rect 890 400 1040 410
rect 890 330 900 400
rect 1030 330 1040 400
rect 390 130 600 140
rect -40 -70 390 130
rect -40 -90 600 -70
rect -40 -1400 220 -90
rect 370 -220 520 -210
rect 370 -310 520 -300
rect 650 -290 680 -280
rect 730 -380 780 -290
rect 650 -410 780 -380
rect -40 -2110 -30 -1400
rect 210 -2110 220 -1400
rect 440 -740 520 -730
rect 440 -830 450 -740
rect 440 -1410 520 -830
rect 550 -860 640 -850
rect 550 -990 640 -980
rect 680 -1260 780 -410
rect 890 -550 1040 330
rect 1220 290 1280 300
rect 1220 210 1280 220
rect 1650 290 1780 640
rect 1650 220 1670 290
rect 1760 220 1780 290
rect 1650 -290 1780 220
rect 2160 290 2220 300
rect 2160 210 2220 220
rect 1650 -380 1670 -290
rect 1760 -380 1780 -290
rect 2400 180 2540 190
rect 2520 120 2540 180
rect 1670 -390 1760 -380
rect 890 -660 900 -550
rect 1030 -660 1040 -550
rect 1680 -450 1760 -440
rect 1170 -630 1270 -620
rect 890 -740 1040 -660
rect 1160 -720 1170 -660
rect 880 -750 1050 -740
rect 880 -840 1050 -830
rect 890 -940 1060 -930
rect 890 -1040 1060 -1030
rect 1160 -1170 1270 -720
rect 1160 -1260 1170 -1170
rect 680 -1270 800 -1260
rect 680 -1340 710 -1270
rect 680 -1350 800 -1340
rect 540 -1420 550 -1410
rect 470 -1520 550 -1510
rect -40 -2120 220 -2110
rect 680 -2230 780 -1350
rect 1160 -1410 1270 -1260
rect 1560 -1060 1640 -1050
rect 1560 -1120 1570 -1060
rect 1560 -1280 1640 -1120
rect 1680 -1140 1760 -520
rect 1680 -1250 1760 -1240
rect 2170 -630 2280 -620
rect 2270 -720 2280 -630
rect 2170 -1170 2280 -720
rect 2400 -750 2540 120
rect 2840 130 3040 140
rect 3040 -90 3750 130
rect 2840 -100 3040 -90
rect 2890 -180 3040 -170
rect 2890 -250 3040 -240
rect 2650 -290 3300 -280
rect 2650 -380 2710 -290
rect 2790 -380 3300 -290
rect 2650 -410 3300 -380
rect 2390 -760 2560 -750
rect 2390 -860 2560 -850
rect 2380 -950 2550 -940
rect 2380 -1050 2550 -1040
rect 2270 -1260 2280 -1170
rect 2030 -1280 2100 -1270
rect 1560 -1340 2030 -1280
rect 2030 -1350 2100 -1340
rect 2170 -1410 2280 -1260
rect 2650 -1270 2750 -410
rect 2810 -550 2910 -540
rect 2790 -640 2820 -550
rect 2790 -660 2910 -640
rect 3210 -650 3300 -410
rect 3570 -580 3750 -90
rect 2790 -880 2840 -660
rect 3210 -740 3300 -730
rect 2880 -750 2990 -740
rect 2970 -850 2990 -750
rect 2880 -860 2990 -850
rect 2790 -890 2850 -880
rect 2790 -1030 2850 -1020
rect 2630 -1280 2750 -1270
rect 2730 -1350 2750 -1280
rect 2630 -1360 2750 -1350
rect 1160 -1420 1560 -1410
rect 1160 -1490 1470 -1420
rect 680 -2240 830 -2230
rect 680 -2310 730 -2240
rect 680 -2320 830 -2310
rect 1160 -2340 1270 -1490
rect 1470 -1500 1560 -1490
rect 1880 -1420 2280 -1410
rect 1960 -1490 2280 -1420
rect 1880 -1500 1960 -1490
rect 1160 -2410 1270 -2400
rect 2170 -2340 2280 -1490
rect 2640 -2250 2750 -1360
rect 2900 -1410 2990 -860
rect 3360 -790 3500 -780
rect 3050 -930 3160 -920
rect 3360 -950 3500 -940
rect 3050 -1050 3160 -1040
rect 3580 -1400 3740 -580
rect 2900 -1530 2990 -1520
rect 3320 -1410 3740 -1400
rect 3580 -2120 3740 -1410
rect 3320 -2130 3740 -2120
rect 2720 -2310 2750 -2250
rect 2640 -2320 2750 -2310
rect 2170 -2420 2280 -2410
rect 490 -2620 600 -2610
rect 490 -2750 600 -2740
rect 2760 -2630 2880 -2620
rect 2760 -2760 2880 -2750
rect 790 -3010 2540 -3000
rect 790 -3220 2540 -3210
<< via2 >>
rect 370 -300 520 -220
rect 650 -380 730 -290
rect 550 -870 640 -860
rect 550 -970 560 -870
rect 560 -970 630 -870
rect 630 -970 640 -870
rect 550 -980 640 -970
rect 1220 220 1280 290
rect 1670 220 1760 290
rect 2160 220 2220 290
rect 1670 -380 1760 -290
rect 900 -660 1030 -550
rect 890 -1030 1060 -940
rect 1680 -1150 1760 -1140
rect 1680 -1230 1760 -1150
rect 1680 -1240 1760 -1230
rect 2890 -240 3040 -180
rect 2710 -380 2790 -290
rect 2390 -850 2560 -760
rect 2380 -1040 2550 -950
rect 2820 -640 2910 -550
rect 3050 -1040 3150 -940
rect 3360 -940 3500 -790
rect 490 -2740 600 -2620
rect 2760 -2750 2880 -2630
rect 790 -3210 2540 -3010
<< metal3 >>
rect 1210 290 1290 295
rect 1660 290 1770 295
rect 2150 290 2230 295
rect 1210 220 1220 290
rect 1280 220 1670 290
rect 1760 220 2160 290
rect 2220 220 2230 290
rect 1210 215 2230 220
rect 1220 210 2210 215
rect 570 -60 580 -40
rect 370 -200 580 -60
rect 740 -200 750 -40
rect 2690 -200 2700 -40
rect 2860 -60 2870 -40
rect 2860 -175 3040 -60
rect 2860 -180 3050 -175
rect 2860 -200 2890 -180
rect 370 -215 530 -200
rect 360 -220 530 -215
rect 360 -300 370 -220
rect 520 -300 530 -220
rect 2880 -240 2890 -200
rect 3040 -240 3050 -180
rect 2880 -245 3050 -240
rect 360 -305 530 -300
rect 640 -280 810 -270
rect 640 -290 1190 -280
rect 640 -380 650 -290
rect 730 -380 1190 -290
rect 640 -385 1190 -380
rect 690 -390 1190 -385
rect 1300 -290 2160 -280
rect 1300 -380 1670 -290
rect 1760 -380 2160 -290
rect 1300 -390 2160 -380
rect 2270 -285 2750 -280
rect 2270 -290 2800 -285
rect 2270 -380 2710 -290
rect 2790 -380 2800 -290
rect 2270 -385 2800 -380
rect 2270 -390 2750 -385
rect 890 -550 2920 -540
rect 890 -660 900 -550
rect 1030 -640 2820 -550
rect 2910 -640 2920 -550
rect 1030 -660 2920 -640
rect 890 -670 2920 -660
rect 2380 -760 2570 -750
rect 2380 -770 2390 -760
rect 540 -850 2390 -770
rect 2560 -850 2570 -760
rect 540 -855 2570 -850
rect 3350 -790 3510 -785
rect 540 -860 2550 -855
rect 540 -980 550 -860
rect 640 -980 650 -860
rect 540 -985 650 -980
rect 880 -940 1070 -935
rect 3040 -940 3160 -935
rect 880 -1030 890 -940
rect 1060 -950 1070 -940
rect 2470 -945 3050 -940
rect 2370 -950 3050 -945
rect 1060 -1030 2380 -950
rect 880 -1040 2380 -1030
rect 2550 -1040 3050 -950
rect 3150 -1040 3160 -940
rect 3350 -940 3360 -790
rect 3500 -940 3510 -790
rect 3350 -945 3510 -940
rect 2370 -1045 2560 -1040
rect 3040 -1045 3160 -1040
rect 1670 -1140 1770 -1135
rect 1670 -1240 1680 -1140
rect 1760 -1240 1770 -1140
rect 1670 -1245 1770 -1240
rect 480 -2620 610 -2615
rect 480 -2740 490 -2620
rect 600 -2630 610 -2620
rect 2750 -2630 2890 -2625
rect 600 -2740 2760 -2630
rect 480 -2745 2760 -2740
rect 490 -2750 2760 -2745
rect 2880 -2750 2890 -2630
rect 2750 -2755 2890 -2750
rect 780 -3010 2550 -3005
rect 780 -3210 790 -3010
rect 2540 -3210 2550 -3010
rect 780 -3215 2550 -3210
<< via3 >>
rect 580 -200 740 -40
rect 2700 -200 2860 -40
rect 3360 -940 3500 -790
rect 1680 -1240 1760 -1140
rect 790 -3210 2540 -3010
<< metal4 >>
rect 579 -40 741 -39
rect 2699 -40 2861 -39
rect 579 -200 580 -40
rect 740 -200 2700 -40
rect 2860 -200 2861 -40
rect 579 -201 741 -200
rect 1640 -1140 1800 -200
rect 2699 -201 2861 -200
rect 1640 -1240 1680 -1140
rect 1760 -1240 1800 -1140
rect 1640 -2970 1800 -1240
rect 3310 -790 3570 -750
rect 3310 -940 3360 -790
rect 3500 -940 3570 -790
rect 3310 -2970 3570 -940
rect 710 -3010 3570 -2970
rect 710 -3210 790 -3010
rect 2540 -3210 3570 -3010
rect 710 -3250 3570 -3210
use sky130_fd_pr__cap_var_lvt_CYVAFU  XC1
timestamp 1715635929
transform 1 0 1409 0 1 -942
box -151 -318 151 318
use sky130_fd_pr__cap_var_lvt_CYVAFU  XC2
timestamp 1715635929
transform 1 0 2031 0 1 -942
box -151 -318 151 318
use sky130_fd_pr__nfet_01v8_lvt_64Z3AY  XM1
timestamp 1715635929
transform 1 0 3251 0 1 -841
box -211 -279 211 279
use sky130_fd_pr__pfet_01v8_lvt_4QFHB3  XM2
timestamp 1715635929
transform 0 1 1719 -1 0 251
box -231 -619 231 619
use sky130_fd_pr__nfet_01v8_lvt_AWHWK2  XM3
timestamp 1715635929
transform 0 1 2274 -1 0 -334
box -256 -610 256 610
use sky130_fd_pr__nfet_01v8_lvt_AWHWK2  XM4
timestamp 1715635929
transform 0 1 1160 -1 0 -334
box -256 -610 256 610
use sky130_fd_pr__pfet_01v8_lvt_4QFHB3  XM6
timestamp 1715635929
transform 1 0 3057 0 1 -1791
box -231 -619 231 619
use sky130_fd_pr__pfet_01v8_lvt_4QFHB3  XM7
timestamp 1715635929
transform 1 0 385 0 1 -1781
box -231 -619 231 619
use sky130_fd_pr__pfet_01v8_lvt_4QFHB3  XM9
timestamp 1715635929
transform -1 0 2701 0 -1 -1791
box -231 -619 231 619
use sky130_fd_pr__nfet_01v8_lvt_64Z3AY  XM10
timestamp 1715635929
transform 0 -1 941 1 0 -909
box -211 -279 211 279
use sky130_fd_pr__nfet_01v8_lvt_64Z3AY  XM11
timestamp 1715635929
transform 0 1 2499 -1 0 -919
box -211 -279 211 279
use sky130_fd_pr__nfet_01v8_lvt_WJMR3R  XM13
timestamp 1715635929
transform 0 1 1719 -1 0 -2690
box -256 -1119 256 1119
use sky130_fd_pr__pfet_01v8_lvt_4QFHB3  XM14
timestamp 1715635929
transform -1 0 741 0 -1 -1781
box -231 -619 231 619
use sky130_fd_pr__nfet_01v8_lvt_AWHWK2  XM15
timestamp 1715635929
transform 1 0 1922 0 1 -1930
box -256 -610 256 610
use sky130_fd_pr__nfet_01v8_lvt_AWHWK2  XM17
timestamp 1715635929
transform 1 0 1516 0 1 -1930
box -256 -610 256 610
<< labels >>
flabel metal1 370 250 570 450 0 FreeSans 256 0 0 0 VDD
port 0 nsew
flabel metal4 1620 -3190 1820 -2990 0 FreeSans 256 0 0 0 VSS
port 7 nsew
flabel metal1 -330 -680 -130 -480 0 FreeSans 256 0 0 0 VIP
port 4 nsew
flabel metal1 900 540 1100 740 0 FreeSans 256 0 0 0 VOP
port 1 nsew
flabel metal1 2390 540 2590 740 0 FreeSans 256 0 0 0 VON
port 2 nsew
flabel metal1 1620 600 1820 800 0 FreeSans 256 0 0 0 CLK
port 6 nsew
flabel metal1 3830 -550 4030 -350 0 FreeSans 256 0 0 0 VIN
port 3 nsew
flabel metal1 150 -2670 350 -2470 0 FreeSans 256 0 0 0 IB
port 5 nsew
<< end >>
