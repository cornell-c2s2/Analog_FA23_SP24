magic
tech sky130A
magscale 1 2
timestamp 1716869746
<< nwell >>
rect -296 -2119 296 2119
<< pmoslvt >>
rect -100 -1900 100 1900
<< pdiff >>
rect -158 1888 -100 1900
rect -158 -1888 -146 1888
rect -112 -1888 -100 1888
rect -158 -1900 -100 -1888
rect 100 1888 158 1900
rect 100 -1888 112 1888
rect 146 -1888 158 1888
rect 100 -1900 158 -1888
<< pdiffc >>
rect -146 -1888 -112 1888
rect 112 -1888 146 1888
<< nsubdiff >>
rect -260 2049 -164 2083
rect 164 2049 260 2083
rect -260 1987 -226 2049
rect 226 1987 260 2049
rect -260 -2049 -226 -1987
rect 226 -2049 260 -1987
rect -260 -2083 -164 -2049
rect 164 -2083 260 -2049
<< nsubdiffcont >>
rect -164 2049 164 2083
rect -260 -1987 -226 1987
rect 226 -1987 260 1987
rect -164 -2083 164 -2049
<< poly >>
rect -100 1981 100 1997
rect -100 1947 -84 1981
rect 84 1947 100 1981
rect -100 1900 100 1947
rect -100 -1947 100 -1900
rect -100 -1981 -84 -1947
rect 84 -1981 100 -1947
rect -100 -1997 100 -1981
<< polycont >>
rect -84 1947 84 1981
rect -84 -1981 84 -1947
<< locali >>
rect -260 2049 -164 2083
rect 164 2049 260 2083
rect -260 1987 -226 2049
rect 226 1987 260 2049
rect -100 1947 -84 1981
rect 84 1947 100 1981
rect -146 1888 -112 1904
rect -146 -1904 -112 -1888
rect 112 1888 146 1904
rect 112 -1904 146 -1888
rect -100 -1981 -84 -1947
rect 84 -1981 100 -1947
rect -260 -2049 -226 -1987
rect 226 -2049 260 -1987
rect -260 -2083 -164 -2049
rect 164 -2083 260 -2049
<< viali >>
rect -84 1947 84 1981
rect -146 -1888 -112 1888
rect 112 -1888 146 1888
rect -84 -1981 84 -1947
<< metal1 >>
rect -96 1981 96 1987
rect -96 1947 -84 1981
rect 84 1947 96 1981
rect -96 1941 96 1947
rect -152 1888 -106 1900
rect -152 -1888 -146 1888
rect -112 -1888 -106 1888
rect -152 -1900 -106 -1888
rect 106 1888 152 1900
rect 106 -1888 112 1888
rect 146 -1888 152 1888
rect 106 -1900 152 -1888
rect -96 -1947 96 -1941
rect -96 -1981 -84 -1947
rect 84 -1981 96 -1947
rect -96 -1987 96 -1981
<< properties >>
string FIXED_BBOX -243 -2066 243 2066
string gencell sky130_fd_pr__pfet_01v8_lvt
string library sky130
string parameters w 19.0 l 1.0 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.35 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
