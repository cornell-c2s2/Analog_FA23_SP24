magic
tech sky130A
magscale 1 2
timestamp 1709401415
<< error_p >>
rect 19 1072 77 1078
rect 19 1038 31 1072
rect 19 1032 77 1038
rect -77 -1038 -19 -1032
rect -77 -1072 -65 -1038
rect -77 -1078 -19 -1072
<< pwell >>
rect -263 -1210 263 1210
<< nmos >>
rect -63 -1000 -33 1000
rect 33 -1000 63 1000
<< ndiff >>
rect -125 988 -63 1000
rect -125 -988 -113 988
rect -79 -988 -63 988
rect -125 -1000 -63 -988
rect -33 988 33 1000
rect -33 -988 -17 988
rect 17 -988 33 988
rect -33 -1000 33 -988
rect 63 988 125 1000
rect 63 -988 79 988
rect 113 -988 125 988
rect 63 -1000 125 -988
<< ndiffc >>
rect -113 -988 -79 988
rect -17 -988 17 988
rect 79 -988 113 988
<< psubdiff >>
rect -227 1140 -131 1174
rect 131 1140 227 1174
rect -227 1078 -193 1140
rect 193 1078 227 1140
rect -227 -1140 -193 -1078
rect 193 -1140 227 -1078
rect -227 -1174 -131 -1140
rect 131 -1174 227 -1140
<< psubdiffcont >>
rect -131 1140 131 1174
rect -227 -1078 -193 1078
rect 193 -1078 227 1078
rect -131 -1174 131 -1140
<< poly >>
rect 15 1072 81 1088
rect 15 1038 31 1072
rect 65 1038 81 1072
rect -63 1000 -33 1026
rect 15 1022 81 1038
rect 33 1000 63 1022
rect -63 -1022 -33 -1000
rect -81 -1038 -15 -1022
rect 33 -1026 63 -1000
rect -81 -1072 -65 -1038
rect -31 -1072 -15 -1038
rect -81 -1088 -15 -1072
<< polycont >>
rect 31 1038 65 1072
rect -65 -1072 -31 -1038
<< locali >>
rect -227 1140 -131 1174
rect 131 1140 227 1174
rect -227 1078 -193 1140
rect 193 1078 227 1140
rect 15 1038 31 1072
rect 65 1038 81 1072
rect -113 988 -79 1004
rect -113 -1004 -79 -988
rect -17 988 17 1004
rect -17 -1004 17 -988
rect 79 988 113 1004
rect 79 -1004 113 -988
rect -81 -1072 -65 -1038
rect -31 -1072 -15 -1038
rect -227 -1140 -193 -1078
rect 193 -1140 227 -1078
rect -227 -1174 -131 -1140
rect 131 -1174 227 -1140
<< viali >>
rect 31 1038 65 1072
rect -113 -988 -79 988
rect -17 -988 17 988
rect 79 -988 113 988
rect -65 -1072 -31 -1038
<< metal1 >>
rect 19 1072 77 1078
rect 19 1038 31 1072
rect 65 1038 77 1072
rect 19 1032 77 1038
rect -119 988 -73 1000
rect -119 -988 -113 988
rect -79 -988 -73 988
rect -119 -1000 -73 -988
rect -23 988 23 1000
rect -23 -988 -17 988
rect 17 -988 23 988
rect -23 -1000 23 -988
rect 73 988 119 1000
rect 73 -988 79 988
rect 113 -988 119 988
rect 73 -1000 119 -988
rect -77 -1038 -19 -1032
rect -77 -1072 -65 -1038
rect -31 -1072 -19 -1038
rect -77 -1078 -19 -1072
<< properties >>
string FIXED_BBOX -210 -1157 210 1157
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 10 l 0.150 m 1 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
