magic
tech sky130A
magscale 1 2
timestamp 1709390584
<< nwell >>
rect -296 -719 296 719
<< pmos >>
rect -100 -500 100 500
<< pdiff >>
rect -158 488 -100 500
rect -158 -488 -146 488
rect -112 -488 -100 488
rect -158 -500 -100 -488
rect 100 488 158 500
rect 100 -488 112 488
rect 146 -488 158 488
rect 100 -500 158 -488
<< pdiffc >>
rect -146 -488 -112 488
rect 112 -488 146 488
<< nsubdiff >>
rect -260 649 -164 683
rect 164 649 260 683
rect -260 587 -226 649
rect 226 587 260 649
rect -260 -649 -226 -587
rect 226 -649 260 -587
rect -260 -683 -164 -649
rect 164 -683 260 -649
<< nsubdiffcont >>
rect -164 649 164 683
rect -260 -587 -226 587
rect 226 -587 260 587
rect -164 -683 164 -649
<< poly >>
rect -100 581 100 597
rect -100 547 -84 581
rect 84 547 100 581
rect -100 500 100 547
rect -100 -547 100 -500
rect -100 -581 -84 -547
rect 84 -581 100 -547
rect -100 -597 100 -581
<< polycont >>
rect -84 547 84 581
rect -84 -581 84 -547
<< locali >>
rect -260 649 -164 683
rect 164 649 260 683
rect -260 587 -226 649
rect 226 587 260 649
rect -100 547 -84 581
rect 84 547 100 581
rect -146 488 -112 504
rect -146 -504 -112 -488
rect 112 488 146 504
rect 112 -504 146 -488
rect -100 -581 -84 -547
rect 84 -581 100 -547
rect -260 -649 -226 -587
rect 226 -649 260 -587
rect -260 -683 -164 -649
rect 164 -683 260 -649
<< viali >>
rect -84 547 84 581
rect -146 -488 -112 488
rect 112 -488 146 488
rect -84 -581 84 -547
<< metal1 >>
rect -96 581 96 587
rect -96 547 -84 581
rect 84 547 96 581
rect -96 541 96 547
rect -152 488 -106 500
rect -152 -488 -146 488
rect -112 -488 -106 488
rect -152 -500 -106 -488
rect 106 488 152 500
rect 106 -488 112 488
rect 146 -488 152 488
rect 106 -500 152 -488
rect -96 -547 96 -541
rect -96 -581 -84 -547
rect 84 -581 96 -547
rect -96 -587 96 -581
<< properties >>
string FIXED_BBOX -243 -666 243 666
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 5.0 l 1.0 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
