magic
tech sky130A
magscale 1 2
timestamp 1710000196
<< nwell >>
rect -3327 -719 3327 719
<< pmos >>
rect -3131 -500 -3031 500
rect -2973 -500 -2873 500
rect -2815 -500 -2715 500
rect -2657 -500 -2557 500
rect -2499 -500 -2399 500
rect -2341 -500 -2241 500
rect -2183 -500 -2083 500
rect -2025 -500 -1925 500
rect -1867 -500 -1767 500
rect -1709 -500 -1609 500
rect -1551 -500 -1451 500
rect -1393 -500 -1293 500
rect -1235 -500 -1135 500
rect -1077 -500 -977 500
rect -919 -500 -819 500
rect -761 -500 -661 500
rect -603 -500 -503 500
rect -445 -500 -345 500
rect -287 -500 -187 500
rect -129 -500 -29 500
rect 29 -500 129 500
rect 187 -500 287 500
rect 345 -500 445 500
rect 503 -500 603 500
rect 661 -500 761 500
rect 819 -500 919 500
rect 977 -500 1077 500
rect 1135 -500 1235 500
rect 1293 -500 1393 500
rect 1451 -500 1551 500
rect 1609 -500 1709 500
rect 1767 -500 1867 500
rect 1925 -500 2025 500
rect 2083 -500 2183 500
rect 2241 -500 2341 500
rect 2399 -500 2499 500
rect 2557 -500 2657 500
rect 2715 -500 2815 500
rect 2873 -500 2973 500
rect 3031 -500 3131 500
<< pdiff >>
rect -3189 459 -3131 500
rect -3189 425 -3177 459
rect -3143 425 -3131 459
rect -3189 391 -3131 425
rect -3189 357 -3177 391
rect -3143 357 -3131 391
rect -3189 323 -3131 357
rect -3189 289 -3177 323
rect -3143 289 -3131 323
rect -3189 255 -3131 289
rect -3189 221 -3177 255
rect -3143 221 -3131 255
rect -3189 187 -3131 221
rect -3189 153 -3177 187
rect -3143 153 -3131 187
rect -3189 119 -3131 153
rect -3189 85 -3177 119
rect -3143 85 -3131 119
rect -3189 51 -3131 85
rect -3189 17 -3177 51
rect -3143 17 -3131 51
rect -3189 -17 -3131 17
rect -3189 -51 -3177 -17
rect -3143 -51 -3131 -17
rect -3189 -85 -3131 -51
rect -3189 -119 -3177 -85
rect -3143 -119 -3131 -85
rect -3189 -153 -3131 -119
rect -3189 -187 -3177 -153
rect -3143 -187 -3131 -153
rect -3189 -221 -3131 -187
rect -3189 -255 -3177 -221
rect -3143 -255 -3131 -221
rect -3189 -289 -3131 -255
rect -3189 -323 -3177 -289
rect -3143 -323 -3131 -289
rect -3189 -357 -3131 -323
rect -3189 -391 -3177 -357
rect -3143 -391 -3131 -357
rect -3189 -425 -3131 -391
rect -3189 -459 -3177 -425
rect -3143 -459 -3131 -425
rect -3189 -500 -3131 -459
rect -3031 459 -2973 500
rect -3031 425 -3019 459
rect -2985 425 -2973 459
rect -3031 391 -2973 425
rect -3031 357 -3019 391
rect -2985 357 -2973 391
rect -3031 323 -2973 357
rect -3031 289 -3019 323
rect -2985 289 -2973 323
rect -3031 255 -2973 289
rect -3031 221 -3019 255
rect -2985 221 -2973 255
rect -3031 187 -2973 221
rect -3031 153 -3019 187
rect -2985 153 -2973 187
rect -3031 119 -2973 153
rect -3031 85 -3019 119
rect -2985 85 -2973 119
rect -3031 51 -2973 85
rect -3031 17 -3019 51
rect -2985 17 -2973 51
rect -3031 -17 -2973 17
rect -3031 -51 -3019 -17
rect -2985 -51 -2973 -17
rect -3031 -85 -2973 -51
rect -3031 -119 -3019 -85
rect -2985 -119 -2973 -85
rect -3031 -153 -2973 -119
rect -3031 -187 -3019 -153
rect -2985 -187 -2973 -153
rect -3031 -221 -2973 -187
rect -3031 -255 -3019 -221
rect -2985 -255 -2973 -221
rect -3031 -289 -2973 -255
rect -3031 -323 -3019 -289
rect -2985 -323 -2973 -289
rect -3031 -357 -2973 -323
rect -3031 -391 -3019 -357
rect -2985 -391 -2973 -357
rect -3031 -425 -2973 -391
rect -3031 -459 -3019 -425
rect -2985 -459 -2973 -425
rect -3031 -500 -2973 -459
rect -2873 459 -2815 500
rect -2873 425 -2861 459
rect -2827 425 -2815 459
rect -2873 391 -2815 425
rect -2873 357 -2861 391
rect -2827 357 -2815 391
rect -2873 323 -2815 357
rect -2873 289 -2861 323
rect -2827 289 -2815 323
rect -2873 255 -2815 289
rect -2873 221 -2861 255
rect -2827 221 -2815 255
rect -2873 187 -2815 221
rect -2873 153 -2861 187
rect -2827 153 -2815 187
rect -2873 119 -2815 153
rect -2873 85 -2861 119
rect -2827 85 -2815 119
rect -2873 51 -2815 85
rect -2873 17 -2861 51
rect -2827 17 -2815 51
rect -2873 -17 -2815 17
rect -2873 -51 -2861 -17
rect -2827 -51 -2815 -17
rect -2873 -85 -2815 -51
rect -2873 -119 -2861 -85
rect -2827 -119 -2815 -85
rect -2873 -153 -2815 -119
rect -2873 -187 -2861 -153
rect -2827 -187 -2815 -153
rect -2873 -221 -2815 -187
rect -2873 -255 -2861 -221
rect -2827 -255 -2815 -221
rect -2873 -289 -2815 -255
rect -2873 -323 -2861 -289
rect -2827 -323 -2815 -289
rect -2873 -357 -2815 -323
rect -2873 -391 -2861 -357
rect -2827 -391 -2815 -357
rect -2873 -425 -2815 -391
rect -2873 -459 -2861 -425
rect -2827 -459 -2815 -425
rect -2873 -500 -2815 -459
rect -2715 459 -2657 500
rect -2715 425 -2703 459
rect -2669 425 -2657 459
rect -2715 391 -2657 425
rect -2715 357 -2703 391
rect -2669 357 -2657 391
rect -2715 323 -2657 357
rect -2715 289 -2703 323
rect -2669 289 -2657 323
rect -2715 255 -2657 289
rect -2715 221 -2703 255
rect -2669 221 -2657 255
rect -2715 187 -2657 221
rect -2715 153 -2703 187
rect -2669 153 -2657 187
rect -2715 119 -2657 153
rect -2715 85 -2703 119
rect -2669 85 -2657 119
rect -2715 51 -2657 85
rect -2715 17 -2703 51
rect -2669 17 -2657 51
rect -2715 -17 -2657 17
rect -2715 -51 -2703 -17
rect -2669 -51 -2657 -17
rect -2715 -85 -2657 -51
rect -2715 -119 -2703 -85
rect -2669 -119 -2657 -85
rect -2715 -153 -2657 -119
rect -2715 -187 -2703 -153
rect -2669 -187 -2657 -153
rect -2715 -221 -2657 -187
rect -2715 -255 -2703 -221
rect -2669 -255 -2657 -221
rect -2715 -289 -2657 -255
rect -2715 -323 -2703 -289
rect -2669 -323 -2657 -289
rect -2715 -357 -2657 -323
rect -2715 -391 -2703 -357
rect -2669 -391 -2657 -357
rect -2715 -425 -2657 -391
rect -2715 -459 -2703 -425
rect -2669 -459 -2657 -425
rect -2715 -500 -2657 -459
rect -2557 459 -2499 500
rect -2557 425 -2545 459
rect -2511 425 -2499 459
rect -2557 391 -2499 425
rect -2557 357 -2545 391
rect -2511 357 -2499 391
rect -2557 323 -2499 357
rect -2557 289 -2545 323
rect -2511 289 -2499 323
rect -2557 255 -2499 289
rect -2557 221 -2545 255
rect -2511 221 -2499 255
rect -2557 187 -2499 221
rect -2557 153 -2545 187
rect -2511 153 -2499 187
rect -2557 119 -2499 153
rect -2557 85 -2545 119
rect -2511 85 -2499 119
rect -2557 51 -2499 85
rect -2557 17 -2545 51
rect -2511 17 -2499 51
rect -2557 -17 -2499 17
rect -2557 -51 -2545 -17
rect -2511 -51 -2499 -17
rect -2557 -85 -2499 -51
rect -2557 -119 -2545 -85
rect -2511 -119 -2499 -85
rect -2557 -153 -2499 -119
rect -2557 -187 -2545 -153
rect -2511 -187 -2499 -153
rect -2557 -221 -2499 -187
rect -2557 -255 -2545 -221
rect -2511 -255 -2499 -221
rect -2557 -289 -2499 -255
rect -2557 -323 -2545 -289
rect -2511 -323 -2499 -289
rect -2557 -357 -2499 -323
rect -2557 -391 -2545 -357
rect -2511 -391 -2499 -357
rect -2557 -425 -2499 -391
rect -2557 -459 -2545 -425
rect -2511 -459 -2499 -425
rect -2557 -500 -2499 -459
rect -2399 459 -2341 500
rect -2399 425 -2387 459
rect -2353 425 -2341 459
rect -2399 391 -2341 425
rect -2399 357 -2387 391
rect -2353 357 -2341 391
rect -2399 323 -2341 357
rect -2399 289 -2387 323
rect -2353 289 -2341 323
rect -2399 255 -2341 289
rect -2399 221 -2387 255
rect -2353 221 -2341 255
rect -2399 187 -2341 221
rect -2399 153 -2387 187
rect -2353 153 -2341 187
rect -2399 119 -2341 153
rect -2399 85 -2387 119
rect -2353 85 -2341 119
rect -2399 51 -2341 85
rect -2399 17 -2387 51
rect -2353 17 -2341 51
rect -2399 -17 -2341 17
rect -2399 -51 -2387 -17
rect -2353 -51 -2341 -17
rect -2399 -85 -2341 -51
rect -2399 -119 -2387 -85
rect -2353 -119 -2341 -85
rect -2399 -153 -2341 -119
rect -2399 -187 -2387 -153
rect -2353 -187 -2341 -153
rect -2399 -221 -2341 -187
rect -2399 -255 -2387 -221
rect -2353 -255 -2341 -221
rect -2399 -289 -2341 -255
rect -2399 -323 -2387 -289
rect -2353 -323 -2341 -289
rect -2399 -357 -2341 -323
rect -2399 -391 -2387 -357
rect -2353 -391 -2341 -357
rect -2399 -425 -2341 -391
rect -2399 -459 -2387 -425
rect -2353 -459 -2341 -425
rect -2399 -500 -2341 -459
rect -2241 459 -2183 500
rect -2241 425 -2229 459
rect -2195 425 -2183 459
rect -2241 391 -2183 425
rect -2241 357 -2229 391
rect -2195 357 -2183 391
rect -2241 323 -2183 357
rect -2241 289 -2229 323
rect -2195 289 -2183 323
rect -2241 255 -2183 289
rect -2241 221 -2229 255
rect -2195 221 -2183 255
rect -2241 187 -2183 221
rect -2241 153 -2229 187
rect -2195 153 -2183 187
rect -2241 119 -2183 153
rect -2241 85 -2229 119
rect -2195 85 -2183 119
rect -2241 51 -2183 85
rect -2241 17 -2229 51
rect -2195 17 -2183 51
rect -2241 -17 -2183 17
rect -2241 -51 -2229 -17
rect -2195 -51 -2183 -17
rect -2241 -85 -2183 -51
rect -2241 -119 -2229 -85
rect -2195 -119 -2183 -85
rect -2241 -153 -2183 -119
rect -2241 -187 -2229 -153
rect -2195 -187 -2183 -153
rect -2241 -221 -2183 -187
rect -2241 -255 -2229 -221
rect -2195 -255 -2183 -221
rect -2241 -289 -2183 -255
rect -2241 -323 -2229 -289
rect -2195 -323 -2183 -289
rect -2241 -357 -2183 -323
rect -2241 -391 -2229 -357
rect -2195 -391 -2183 -357
rect -2241 -425 -2183 -391
rect -2241 -459 -2229 -425
rect -2195 -459 -2183 -425
rect -2241 -500 -2183 -459
rect -2083 459 -2025 500
rect -2083 425 -2071 459
rect -2037 425 -2025 459
rect -2083 391 -2025 425
rect -2083 357 -2071 391
rect -2037 357 -2025 391
rect -2083 323 -2025 357
rect -2083 289 -2071 323
rect -2037 289 -2025 323
rect -2083 255 -2025 289
rect -2083 221 -2071 255
rect -2037 221 -2025 255
rect -2083 187 -2025 221
rect -2083 153 -2071 187
rect -2037 153 -2025 187
rect -2083 119 -2025 153
rect -2083 85 -2071 119
rect -2037 85 -2025 119
rect -2083 51 -2025 85
rect -2083 17 -2071 51
rect -2037 17 -2025 51
rect -2083 -17 -2025 17
rect -2083 -51 -2071 -17
rect -2037 -51 -2025 -17
rect -2083 -85 -2025 -51
rect -2083 -119 -2071 -85
rect -2037 -119 -2025 -85
rect -2083 -153 -2025 -119
rect -2083 -187 -2071 -153
rect -2037 -187 -2025 -153
rect -2083 -221 -2025 -187
rect -2083 -255 -2071 -221
rect -2037 -255 -2025 -221
rect -2083 -289 -2025 -255
rect -2083 -323 -2071 -289
rect -2037 -323 -2025 -289
rect -2083 -357 -2025 -323
rect -2083 -391 -2071 -357
rect -2037 -391 -2025 -357
rect -2083 -425 -2025 -391
rect -2083 -459 -2071 -425
rect -2037 -459 -2025 -425
rect -2083 -500 -2025 -459
rect -1925 459 -1867 500
rect -1925 425 -1913 459
rect -1879 425 -1867 459
rect -1925 391 -1867 425
rect -1925 357 -1913 391
rect -1879 357 -1867 391
rect -1925 323 -1867 357
rect -1925 289 -1913 323
rect -1879 289 -1867 323
rect -1925 255 -1867 289
rect -1925 221 -1913 255
rect -1879 221 -1867 255
rect -1925 187 -1867 221
rect -1925 153 -1913 187
rect -1879 153 -1867 187
rect -1925 119 -1867 153
rect -1925 85 -1913 119
rect -1879 85 -1867 119
rect -1925 51 -1867 85
rect -1925 17 -1913 51
rect -1879 17 -1867 51
rect -1925 -17 -1867 17
rect -1925 -51 -1913 -17
rect -1879 -51 -1867 -17
rect -1925 -85 -1867 -51
rect -1925 -119 -1913 -85
rect -1879 -119 -1867 -85
rect -1925 -153 -1867 -119
rect -1925 -187 -1913 -153
rect -1879 -187 -1867 -153
rect -1925 -221 -1867 -187
rect -1925 -255 -1913 -221
rect -1879 -255 -1867 -221
rect -1925 -289 -1867 -255
rect -1925 -323 -1913 -289
rect -1879 -323 -1867 -289
rect -1925 -357 -1867 -323
rect -1925 -391 -1913 -357
rect -1879 -391 -1867 -357
rect -1925 -425 -1867 -391
rect -1925 -459 -1913 -425
rect -1879 -459 -1867 -425
rect -1925 -500 -1867 -459
rect -1767 459 -1709 500
rect -1767 425 -1755 459
rect -1721 425 -1709 459
rect -1767 391 -1709 425
rect -1767 357 -1755 391
rect -1721 357 -1709 391
rect -1767 323 -1709 357
rect -1767 289 -1755 323
rect -1721 289 -1709 323
rect -1767 255 -1709 289
rect -1767 221 -1755 255
rect -1721 221 -1709 255
rect -1767 187 -1709 221
rect -1767 153 -1755 187
rect -1721 153 -1709 187
rect -1767 119 -1709 153
rect -1767 85 -1755 119
rect -1721 85 -1709 119
rect -1767 51 -1709 85
rect -1767 17 -1755 51
rect -1721 17 -1709 51
rect -1767 -17 -1709 17
rect -1767 -51 -1755 -17
rect -1721 -51 -1709 -17
rect -1767 -85 -1709 -51
rect -1767 -119 -1755 -85
rect -1721 -119 -1709 -85
rect -1767 -153 -1709 -119
rect -1767 -187 -1755 -153
rect -1721 -187 -1709 -153
rect -1767 -221 -1709 -187
rect -1767 -255 -1755 -221
rect -1721 -255 -1709 -221
rect -1767 -289 -1709 -255
rect -1767 -323 -1755 -289
rect -1721 -323 -1709 -289
rect -1767 -357 -1709 -323
rect -1767 -391 -1755 -357
rect -1721 -391 -1709 -357
rect -1767 -425 -1709 -391
rect -1767 -459 -1755 -425
rect -1721 -459 -1709 -425
rect -1767 -500 -1709 -459
rect -1609 459 -1551 500
rect -1609 425 -1597 459
rect -1563 425 -1551 459
rect -1609 391 -1551 425
rect -1609 357 -1597 391
rect -1563 357 -1551 391
rect -1609 323 -1551 357
rect -1609 289 -1597 323
rect -1563 289 -1551 323
rect -1609 255 -1551 289
rect -1609 221 -1597 255
rect -1563 221 -1551 255
rect -1609 187 -1551 221
rect -1609 153 -1597 187
rect -1563 153 -1551 187
rect -1609 119 -1551 153
rect -1609 85 -1597 119
rect -1563 85 -1551 119
rect -1609 51 -1551 85
rect -1609 17 -1597 51
rect -1563 17 -1551 51
rect -1609 -17 -1551 17
rect -1609 -51 -1597 -17
rect -1563 -51 -1551 -17
rect -1609 -85 -1551 -51
rect -1609 -119 -1597 -85
rect -1563 -119 -1551 -85
rect -1609 -153 -1551 -119
rect -1609 -187 -1597 -153
rect -1563 -187 -1551 -153
rect -1609 -221 -1551 -187
rect -1609 -255 -1597 -221
rect -1563 -255 -1551 -221
rect -1609 -289 -1551 -255
rect -1609 -323 -1597 -289
rect -1563 -323 -1551 -289
rect -1609 -357 -1551 -323
rect -1609 -391 -1597 -357
rect -1563 -391 -1551 -357
rect -1609 -425 -1551 -391
rect -1609 -459 -1597 -425
rect -1563 -459 -1551 -425
rect -1609 -500 -1551 -459
rect -1451 459 -1393 500
rect -1451 425 -1439 459
rect -1405 425 -1393 459
rect -1451 391 -1393 425
rect -1451 357 -1439 391
rect -1405 357 -1393 391
rect -1451 323 -1393 357
rect -1451 289 -1439 323
rect -1405 289 -1393 323
rect -1451 255 -1393 289
rect -1451 221 -1439 255
rect -1405 221 -1393 255
rect -1451 187 -1393 221
rect -1451 153 -1439 187
rect -1405 153 -1393 187
rect -1451 119 -1393 153
rect -1451 85 -1439 119
rect -1405 85 -1393 119
rect -1451 51 -1393 85
rect -1451 17 -1439 51
rect -1405 17 -1393 51
rect -1451 -17 -1393 17
rect -1451 -51 -1439 -17
rect -1405 -51 -1393 -17
rect -1451 -85 -1393 -51
rect -1451 -119 -1439 -85
rect -1405 -119 -1393 -85
rect -1451 -153 -1393 -119
rect -1451 -187 -1439 -153
rect -1405 -187 -1393 -153
rect -1451 -221 -1393 -187
rect -1451 -255 -1439 -221
rect -1405 -255 -1393 -221
rect -1451 -289 -1393 -255
rect -1451 -323 -1439 -289
rect -1405 -323 -1393 -289
rect -1451 -357 -1393 -323
rect -1451 -391 -1439 -357
rect -1405 -391 -1393 -357
rect -1451 -425 -1393 -391
rect -1451 -459 -1439 -425
rect -1405 -459 -1393 -425
rect -1451 -500 -1393 -459
rect -1293 459 -1235 500
rect -1293 425 -1281 459
rect -1247 425 -1235 459
rect -1293 391 -1235 425
rect -1293 357 -1281 391
rect -1247 357 -1235 391
rect -1293 323 -1235 357
rect -1293 289 -1281 323
rect -1247 289 -1235 323
rect -1293 255 -1235 289
rect -1293 221 -1281 255
rect -1247 221 -1235 255
rect -1293 187 -1235 221
rect -1293 153 -1281 187
rect -1247 153 -1235 187
rect -1293 119 -1235 153
rect -1293 85 -1281 119
rect -1247 85 -1235 119
rect -1293 51 -1235 85
rect -1293 17 -1281 51
rect -1247 17 -1235 51
rect -1293 -17 -1235 17
rect -1293 -51 -1281 -17
rect -1247 -51 -1235 -17
rect -1293 -85 -1235 -51
rect -1293 -119 -1281 -85
rect -1247 -119 -1235 -85
rect -1293 -153 -1235 -119
rect -1293 -187 -1281 -153
rect -1247 -187 -1235 -153
rect -1293 -221 -1235 -187
rect -1293 -255 -1281 -221
rect -1247 -255 -1235 -221
rect -1293 -289 -1235 -255
rect -1293 -323 -1281 -289
rect -1247 -323 -1235 -289
rect -1293 -357 -1235 -323
rect -1293 -391 -1281 -357
rect -1247 -391 -1235 -357
rect -1293 -425 -1235 -391
rect -1293 -459 -1281 -425
rect -1247 -459 -1235 -425
rect -1293 -500 -1235 -459
rect -1135 459 -1077 500
rect -1135 425 -1123 459
rect -1089 425 -1077 459
rect -1135 391 -1077 425
rect -1135 357 -1123 391
rect -1089 357 -1077 391
rect -1135 323 -1077 357
rect -1135 289 -1123 323
rect -1089 289 -1077 323
rect -1135 255 -1077 289
rect -1135 221 -1123 255
rect -1089 221 -1077 255
rect -1135 187 -1077 221
rect -1135 153 -1123 187
rect -1089 153 -1077 187
rect -1135 119 -1077 153
rect -1135 85 -1123 119
rect -1089 85 -1077 119
rect -1135 51 -1077 85
rect -1135 17 -1123 51
rect -1089 17 -1077 51
rect -1135 -17 -1077 17
rect -1135 -51 -1123 -17
rect -1089 -51 -1077 -17
rect -1135 -85 -1077 -51
rect -1135 -119 -1123 -85
rect -1089 -119 -1077 -85
rect -1135 -153 -1077 -119
rect -1135 -187 -1123 -153
rect -1089 -187 -1077 -153
rect -1135 -221 -1077 -187
rect -1135 -255 -1123 -221
rect -1089 -255 -1077 -221
rect -1135 -289 -1077 -255
rect -1135 -323 -1123 -289
rect -1089 -323 -1077 -289
rect -1135 -357 -1077 -323
rect -1135 -391 -1123 -357
rect -1089 -391 -1077 -357
rect -1135 -425 -1077 -391
rect -1135 -459 -1123 -425
rect -1089 -459 -1077 -425
rect -1135 -500 -1077 -459
rect -977 459 -919 500
rect -977 425 -965 459
rect -931 425 -919 459
rect -977 391 -919 425
rect -977 357 -965 391
rect -931 357 -919 391
rect -977 323 -919 357
rect -977 289 -965 323
rect -931 289 -919 323
rect -977 255 -919 289
rect -977 221 -965 255
rect -931 221 -919 255
rect -977 187 -919 221
rect -977 153 -965 187
rect -931 153 -919 187
rect -977 119 -919 153
rect -977 85 -965 119
rect -931 85 -919 119
rect -977 51 -919 85
rect -977 17 -965 51
rect -931 17 -919 51
rect -977 -17 -919 17
rect -977 -51 -965 -17
rect -931 -51 -919 -17
rect -977 -85 -919 -51
rect -977 -119 -965 -85
rect -931 -119 -919 -85
rect -977 -153 -919 -119
rect -977 -187 -965 -153
rect -931 -187 -919 -153
rect -977 -221 -919 -187
rect -977 -255 -965 -221
rect -931 -255 -919 -221
rect -977 -289 -919 -255
rect -977 -323 -965 -289
rect -931 -323 -919 -289
rect -977 -357 -919 -323
rect -977 -391 -965 -357
rect -931 -391 -919 -357
rect -977 -425 -919 -391
rect -977 -459 -965 -425
rect -931 -459 -919 -425
rect -977 -500 -919 -459
rect -819 459 -761 500
rect -819 425 -807 459
rect -773 425 -761 459
rect -819 391 -761 425
rect -819 357 -807 391
rect -773 357 -761 391
rect -819 323 -761 357
rect -819 289 -807 323
rect -773 289 -761 323
rect -819 255 -761 289
rect -819 221 -807 255
rect -773 221 -761 255
rect -819 187 -761 221
rect -819 153 -807 187
rect -773 153 -761 187
rect -819 119 -761 153
rect -819 85 -807 119
rect -773 85 -761 119
rect -819 51 -761 85
rect -819 17 -807 51
rect -773 17 -761 51
rect -819 -17 -761 17
rect -819 -51 -807 -17
rect -773 -51 -761 -17
rect -819 -85 -761 -51
rect -819 -119 -807 -85
rect -773 -119 -761 -85
rect -819 -153 -761 -119
rect -819 -187 -807 -153
rect -773 -187 -761 -153
rect -819 -221 -761 -187
rect -819 -255 -807 -221
rect -773 -255 -761 -221
rect -819 -289 -761 -255
rect -819 -323 -807 -289
rect -773 -323 -761 -289
rect -819 -357 -761 -323
rect -819 -391 -807 -357
rect -773 -391 -761 -357
rect -819 -425 -761 -391
rect -819 -459 -807 -425
rect -773 -459 -761 -425
rect -819 -500 -761 -459
rect -661 459 -603 500
rect -661 425 -649 459
rect -615 425 -603 459
rect -661 391 -603 425
rect -661 357 -649 391
rect -615 357 -603 391
rect -661 323 -603 357
rect -661 289 -649 323
rect -615 289 -603 323
rect -661 255 -603 289
rect -661 221 -649 255
rect -615 221 -603 255
rect -661 187 -603 221
rect -661 153 -649 187
rect -615 153 -603 187
rect -661 119 -603 153
rect -661 85 -649 119
rect -615 85 -603 119
rect -661 51 -603 85
rect -661 17 -649 51
rect -615 17 -603 51
rect -661 -17 -603 17
rect -661 -51 -649 -17
rect -615 -51 -603 -17
rect -661 -85 -603 -51
rect -661 -119 -649 -85
rect -615 -119 -603 -85
rect -661 -153 -603 -119
rect -661 -187 -649 -153
rect -615 -187 -603 -153
rect -661 -221 -603 -187
rect -661 -255 -649 -221
rect -615 -255 -603 -221
rect -661 -289 -603 -255
rect -661 -323 -649 -289
rect -615 -323 -603 -289
rect -661 -357 -603 -323
rect -661 -391 -649 -357
rect -615 -391 -603 -357
rect -661 -425 -603 -391
rect -661 -459 -649 -425
rect -615 -459 -603 -425
rect -661 -500 -603 -459
rect -503 459 -445 500
rect -503 425 -491 459
rect -457 425 -445 459
rect -503 391 -445 425
rect -503 357 -491 391
rect -457 357 -445 391
rect -503 323 -445 357
rect -503 289 -491 323
rect -457 289 -445 323
rect -503 255 -445 289
rect -503 221 -491 255
rect -457 221 -445 255
rect -503 187 -445 221
rect -503 153 -491 187
rect -457 153 -445 187
rect -503 119 -445 153
rect -503 85 -491 119
rect -457 85 -445 119
rect -503 51 -445 85
rect -503 17 -491 51
rect -457 17 -445 51
rect -503 -17 -445 17
rect -503 -51 -491 -17
rect -457 -51 -445 -17
rect -503 -85 -445 -51
rect -503 -119 -491 -85
rect -457 -119 -445 -85
rect -503 -153 -445 -119
rect -503 -187 -491 -153
rect -457 -187 -445 -153
rect -503 -221 -445 -187
rect -503 -255 -491 -221
rect -457 -255 -445 -221
rect -503 -289 -445 -255
rect -503 -323 -491 -289
rect -457 -323 -445 -289
rect -503 -357 -445 -323
rect -503 -391 -491 -357
rect -457 -391 -445 -357
rect -503 -425 -445 -391
rect -503 -459 -491 -425
rect -457 -459 -445 -425
rect -503 -500 -445 -459
rect -345 459 -287 500
rect -345 425 -333 459
rect -299 425 -287 459
rect -345 391 -287 425
rect -345 357 -333 391
rect -299 357 -287 391
rect -345 323 -287 357
rect -345 289 -333 323
rect -299 289 -287 323
rect -345 255 -287 289
rect -345 221 -333 255
rect -299 221 -287 255
rect -345 187 -287 221
rect -345 153 -333 187
rect -299 153 -287 187
rect -345 119 -287 153
rect -345 85 -333 119
rect -299 85 -287 119
rect -345 51 -287 85
rect -345 17 -333 51
rect -299 17 -287 51
rect -345 -17 -287 17
rect -345 -51 -333 -17
rect -299 -51 -287 -17
rect -345 -85 -287 -51
rect -345 -119 -333 -85
rect -299 -119 -287 -85
rect -345 -153 -287 -119
rect -345 -187 -333 -153
rect -299 -187 -287 -153
rect -345 -221 -287 -187
rect -345 -255 -333 -221
rect -299 -255 -287 -221
rect -345 -289 -287 -255
rect -345 -323 -333 -289
rect -299 -323 -287 -289
rect -345 -357 -287 -323
rect -345 -391 -333 -357
rect -299 -391 -287 -357
rect -345 -425 -287 -391
rect -345 -459 -333 -425
rect -299 -459 -287 -425
rect -345 -500 -287 -459
rect -187 459 -129 500
rect -187 425 -175 459
rect -141 425 -129 459
rect -187 391 -129 425
rect -187 357 -175 391
rect -141 357 -129 391
rect -187 323 -129 357
rect -187 289 -175 323
rect -141 289 -129 323
rect -187 255 -129 289
rect -187 221 -175 255
rect -141 221 -129 255
rect -187 187 -129 221
rect -187 153 -175 187
rect -141 153 -129 187
rect -187 119 -129 153
rect -187 85 -175 119
rect -141 85 -129 119
rect -187 51 -129 85
rect -187 17 -175 51
rect -141 17 -129 51
rect -187 -17 -129 17
rect -187 -51 -175 -17
rect -141 -51 -129 -17
rect -187 -85 -129 -51
rect -187 -119 -175 -85
rect -141 -119 -129 -85
rect -187 -153 -129 -119
rect -187 -187 -175 -153
rect -141 -187 -129 -153
rect -187 -221 -129 -187
rect -187 -255 -175 -221
rect -141 -255 -129 -221
rect -187 -289 -129 -255
rect -187 -323 -175 -289
rect -141 -323 -129 -289
rect -187 -357 -129 -323
rect -187 -391 -175 -357
rect -141 -391 -129 -357
rect -187 -425 -129 -391
rect -187 -459 -175 -425
rect -141 -459 -129 -425
rect -187 -500 -129 -459
rect -29 459 29 500
rect -29 425 -17 459
rect 17 425 29 459
rect -29 391 29 425
rect -29 357 -17 391
rect 17 357 29 391
rect -29 323 29 357
rect -29 289 -17 323
rect 17 289 29 323
rect -29 255 29 289
rect -29 221 -17 255
rect 17 221 29 255
rect -29 187 29 221
rect -29 153 -17 187
rect 17 153 29 187
rect -29 119 29 153
rect -29 85 -17 119
rect 17 85 29 119
rect -29 51 29 85
rect -29 17 -17 51
rect 17 17 29 51
rect -29 -17 29 17
rect -29 -51 -17 -17
rect 17 -51 29 -17
rect -29 -85 29 -51
rect -29 -119 -17 -85
rect 17 -119 29 -85
rect -29 -153 29 -119
rect -29 -187 -17 -153
rect 17 -187 29 -153
rect -29 -221 29 -187
rect -29 -255 -17 -221
rect 17 -255 29 -221
rect -29 -289 29 -255
rect -29 -323 -17 -289
rect 17 -323 29 -289
rect -29 -357 29 -323
rect -29 -391 -17 -357
rect 17 -391 29 -357
rect -29 -425 29 -391
rect -29 -459 -17 -425
rect 17 -459 29 -425
rect -29 -500 29 -459
rect 129 459 187 500
rect 129 425 141 459
rect 175 425 187 459
rect 129 391 187 425
rect 129 357 141 391
rect 175 357 187 391
rect 129 323 187 357
rect 129 289 141 323
rect 175 289 187 323
rect 129 255 187 289
rect 129 221 141 255
rect 175 221 187 255
rect 129 187 187 221
rect 129 153 141 187
rect 175 153 187 187
rect 129 119 187 153
rect 129 85 141 119
rect 175 85 187 119
rect 129 51 187 85
rect 129 17 141 51
rect 175 17 187 51
rect 129 -17 187 17
rect 129 -51 141 -17
rect 175 -51 187 -17
rect 129 -85 187 -51
rect 129 -119 141 -85
rect 175 -119 187 -85
rect 129 -153 187 -119
rect 129 -187 141 -153
rect 175 -187 187 -153
rect 129 -221 187 -187
rect 129 -255 141 -221
rect 175 -255 187 -221
rect 129 -289 187 -255
rect 129 -323 141 -289
rect 175 -323 187 -289
rect 129 -357 187 -323
rect 129 -391 141 -357
rect 175 -391 187 -357
rect 129 -425 187 -391
rect 129 -459 141 -425
rect 175 -459 187 -425
rect 129 -500 187 -459
rect 287 459 345 500
rect 287 425 299 459
rect 333 425 345 459
rect 287 391 345 425
rect 287 357 299 391
rect 333 357 345 391
rect 287 323 345 357
rect 287 289 299 323
rect 333 289 345 323
rect 287 255 345 289
rect 287 221 299 255
rect 333 221 345 255
rect 287 187 345 221
rect 287 153 299 187
rect 333 153 345 187
rect 287 119 345 153
rect 287 85 299 119
rect 333 85 345 119
rect 287 51 345 85
rect 287 17 299 51
rect 333 17 345 51
rect 287 -17 345 17
rect 287 -51 299 -17
rect 333 -51 345 -17
rect 287 -85 345 -51
rect 287 -119 299 -85
rect 333 -119 345 -85
rect 287 -153 345 -119
rect 287 -187 299 -153
rect 333 -187 345 -153
rect 287 -221 345 -187
rect 287 -255 299 -221
rect 333 -255 345 -221
rect 287 -289 345 -255
rect 287 -323 299 -289
rect 333 -323 345 -289
rect 287 -357 345 -323
rect 287 -391 299 -357
rect 333 -391 345 -357
rect 287 -425 345 -391
rect 287 -459 299 -425
rect 333 -459 345 -425
rect 287 -500 345 -459
rect 445 459 503 500
rect 445 425 457 459
rect 491 425 503 459
rect 445 391 503 425
rect 445 357 457 391
rect 491 357 503 391
rect 445 323 503 357
rect 445 289 457 323
rect 491 289 503 323
rect 445 255 503 289
rect 445 221 457 255
rect 491 221 503 255
rect 445 187 503 221
rect 445 153 457 187
rect 491 153 503 187
rect 445 119 503 153
rect 445 85 457 119
rect 491 85 503 119
rect 445 51 503 85
rect 445 17 457 51
rect 491 17 503 51
rect 445 -17 503 17
rect 445 -51 457 -17
rect 491 -51 503 -17
rect 445 -85 503 -51
rect 445 -119 457 -85
rect 491 -119 503 -85
rect 445 -153 503 -119
rect 445 -187 457 -153
rect 491 -187 503 -153
rect 445 -221 503 -187
rect 445 -255 457 -221
rect 491 -255 503 -221
rect 445 -289 503 -255
rect 445 -323 457 -289
rect 491 -323 503 -289
rect 445 -357 503 -323
rect 445 -391 457 -357
rect 491 -391 503 -357
rect 445 -425 503 -391
rect 445 -459 457 -425
rect 491 -459 503 -425
rect 445 -500 503 -459
rect 603 459 661 500
rect 603 425 615 459
rect 649 425 661 459
rect 603 391 661 425
rect 603 357 615 391
rect 649 357 661 391
rect 603 323 661 357
rect 603 289 615 323
rect 649 289 661 323
rect 603 255 661 289
rect 603 221 615 255
rect 649 221 661 255
rect 603 187 661 221
rect 603 153 615 187
rect 649 153 661 187
rect 603 119 661 153
rect 603 85 615 119
rect 649 85 661 119
rect 603 51 661 85
rect 603 17 615 51
rect 649 17 661 51
rect 603 -17 661 17
rect 603 -51 615 -17
rect 649 -51 661 -17
rect 603 -85 661 -51
rect 603 -119 615 -85
rect 649 -119 661 -85
rect 603 -153 661 -119
rect 603 -187 615 -153
rect 649 -187 661 -153
rect 603 -221 661 -187
rect 603 -255 615 -221
rect 649 -255 661 -221
rect 603 -289 661 -255
rect 603 -323 615 -289
rect 649 -323 661 -289
rect 603 -357 661 -323
rect 603 -391 615 -357
rect 649 -391 661 -357
rect 603 -425 661 -391
rect 603 -459 615 -425
rect 649 -459 661 -425
rect 603 -500 661 -459
rect 761 459 819 500
rect 761 425 773 459
rect 807 425 819 459
rect 761 391 819 425
rect 761 357 773 391
rect 807 357 819 391
rect 761 323 819 357
rect 761 289 773 323
rect 807 289 819 323
rect 761 255 819 289
rect 761 221 773 255
rect 807 221 819 255
rect 761 187 819 221
rect 761 153 773 187
rect 807 153 819 187
rect 761 119 819 153
rect 761 85 773 119
rect 807 85 819 119
rect 761 51 819 85
rect 761 17 773 51
rect 807 17 819 51
rect 761 -17 819 17
rect 761 -51 773 -17
rect 807 -51 819 -17
rect 761 -85 819 -51
rect 761 -119 773 -85
rect 807 -119 819 -85
rect 761 -153 819 -119
rect 761 -187 773 -153
rect 807 -187 819 -153
rect 761 -221 819 -187
rect 761 -255 773 -221
rect 807 -255 819 -221
rect 761 -289 819 -255
rect 761 -323 773 -289
rect 807 -323 819 -289
rect 761 -357 819 -323
rect 761 -391 773 -357
rect 807 -391 819 -357
rect 761 -425 819 -391
rect 761 -459 773 -425
rect 807 -459 819 -425
rect 761 -500 819 -459
rect 919 459 977 500
rect 919 425 931 459
rect 965 425 977 459
rect 919 391 977 425
rect 919 357 931 391
rect 965 357 977 391
rect 919 323 977 357
rect 919 289 931 323
rect 965 289 977 323
rect 919 255 977 289
rect 919 221 931 255
rect 965 221 977 255
rect 919 187 977 221
rect 919 153 931 187
rect 965 153 977 187
rect 919 119 977 153
rect 919 85 931 119
rect 965 85 977 119
rect 919 51 977 85
rect 919 17 931 51
rect 965 17 977 51
rect 919 -17 977 17
rect 919 -51 931 -17
rect 965 -51 977 -17
rect 919 -85 977 -51
rect 919 -119 931 -85
rect 965 -119 977 -85
rect 919 -153 977 -119
rect 919 -187 931 -153
rect 965 -187 977 -153
rect 919 -221 977 -187
rect 919 -255 931 -221
rect 965 -255 977 -221
rect 919 -289 977 -255
rect 919 -323 931 -289
rect 965 -323 977 -289
rect 919 -357 977 -323
rect 919 -391 931 -357
rect 965 -391 977 -357
rect 919 -425 977 -391
rect 919 -459 931 -425
rect 965 -459 977 -425
rect 919 -500 977 -459
rect 1077 459 1135 500
rect 1077 425 1089 459
rect 1123 425 1135 459
rect 1077 391 1135 425
rect 1077 357 1089 391
rect 1123 357 1135 391
rect 1077 323 1135 357
rect 1077 289 1089 323
rect 1123 289 1135 323
rect 1077 255 1135 289
rect 1077 221 1089 255
rect 1123 221 1135 255
rect 1077 187 1135 221
rect 1077 153 1089 187
rect 1123 153 1135 187
rect 1077 119 1135 153
rect 1077 85 1089 119
rect 1123 85 1135 119
rect 1077 51 1135 85
rect 1077 17 1089 51
rect 1123 17 1135 51
rect 1077 -17 1135 17
rect 1077 -51 1089 -17
rect 1123 -51 1135 -17
rect 1077 -85 1135 -51
rect 1077 -119 1089 -85
rect 1123 -119 1135 -85
rect 1077 -153 1135 -119
rect 1077 -187 1089 -153
rect 1123 -187 1135 -153
rect 1077 -221 1135 -187
rect 1077 -255 1089 -221
rect 1123 -255 1135 -221
rect 1077 -289 1135 -255
rect 1077 -323 1089 -289
rect 1123 -323 1135 -289
rect 1077 -357 1135 -323
rect 1077 -391 1089 -357
rect 1123 -391 1135 -357
rect 1077 -425 1135 -391
rect 1077 -459 1089 -425
rect 1123 -459 1135 -425
rect 1077 -500 1135 -459
rect 1235 459 1293 500
rect 1235 425 1247 459
rect 1281 425 1293 459
rect 1235 391 1293 425
rect 1235 357 1247 391
rect 1281 357 1293 391
rect 1235 323 1293 357
rect 1235 289 1247 323
rect 1281 289 1293 323
rect 1235 255 1293 289
rect 1235 221 1247 255
rect 1281 221 1293 255
rect 1235 187 1293 221
rect 1235 153 1247 187
rect 1281 153 1293 187
rect 1235 119 1293 153
rect 1235 85 1247 119
rect 1281 85 1293 119
rect 1235 51 1293 85
rect 1235 17 1247 51
rect 1281 17 1293 51
rect 1235 -17 1293 17
rect 1235 -51 1247 -17
rect 1281 -51 1293 -17
rect 1235 -85 1293 -51
rect 1235 -119 1247 -85
rect 1281 -119 1293 -85
rect 1235 -153 1293 -119
rect 1235 -187 1247 -153
rect 1281 -187 1293 -153
rect 1235 -221 1293 -187
rect 1235 -255 1247 -221
rect 1281 -255 1293 -221
rect 1235 -289 1293 -255
rect 1235 -323 1247 -289
rect 1281 -323 1293 -289
rect 1235 -357 1293 -323
rect 1235 -391 1247 -357
rect 1281 -391 1293 -357
rect 1235 -425 1293 -391
rect 1235 -459 1247 -425
rect 1281 -459 1293 -425
rect 1235 -500 1293 -459
rect 1393 459 1451 500
rect 1393 425 1405 459
rect 1439 425 1451 459
rect 1393 391 1451 425
rect 1393 357 1405 391
rect 1439 357 1451 391
rect 1393 323 1451 357
rect 1393 289 1405 323
rect 1439 289 1451 323
rect 1393 255 1451 289
rect 1393 221 1405 255
rect 1439 221 1451 255
rect 1393 187 1451 221
rect 1393 153 1405 187
rect 1439 153 1451 187
rect 1393 119 1451 153
rect 1393 85 1405 119
rect 1439 85 1451 119
rect 1393 51 1451 85
rect 1393 17 1405 51
rect 1439 17 1451 51
rect 1393 -17 1451 17
rect 1393 -51 1405 -17
rect 1439 -51 1451 -17
rect 1393 -85 1451 -51
rect 1393 -119 1405 -85
rect 1439 -119 1451 -85
rect 1393 -153 1451 -119
rect 1393 -187 1405 -153
rect 1439 -187 1451 -153
rect 1393 -221 1451 -187
rect 1393 -255 1405 -221
rect 1439 -255 1451 -221
rect 1393 -289 1451 -255
rect 1393 -323 1405 -289
rect 1439 -323 1451 -289
rect 1393 -357 1451 -323
rect 1393 -391 1405 -357
rect 1439 -391 1451 -357
rect 1393 -425 1451 -391
rect 1393 -459 1405 -425
rect 1439 -459 1451 -425
rect 1393 -500 1451 -459
rect 1551 459 1609 500
rect 1551 425 1563 459
rect 1597 425 1609 459
rect 1551 391 1609 425
rect 1551 357 1563 391
rect 1597 357 1609 391
rect 1551 323 1609 357
rect 1551 289 1563 323
rect 1597 289 1609 323
rect 1551 255 1609 289
rect 1551 221 1563 255
rect 1597 221 1609 255
rect 1551 187 1609 221
rect 1551 153 1563 187
rect 1597 153 1609 187
rect 1551 119 1609 153
rect 1551 85 1563 119
rect 1597 85 1609 119
rect 1551 51 1609 85
rect 1551 17 1563 51
rect 1597 17 1609 51
rect 1551 -17 1609 17
rect 1551 -51 1563 -17
rect 1597 -51 1609 -17
rect 1551 -85 1609 -51
rect 1551 -119 1563 -85
rect 1597 -119 1609 -85
rect 1551 -153 1609 -119
rect 1551 -187 1563 -153
rect 1597 -187 1609 -153
rect 1551 -221 1609 -187
rect 1551 -255 1563 -221
rect 1597 -255 1609 -221
rect 1551 -289 1609 -255
rect 1551 -323 1563 -289
rect 1597 -323 1609 -289
rect 1551 -357 1609 -323
rect 1551 -391 1563 -357
rect 1597 -391 1609 -357
rect 1551 -425 1609 -391
rect 1551 -459 1563 -425
rect 1597 -459 1609 -425
rect 1551 -500 1609 -459
rect 1709 459 1767 500
rect 1709 425 1721 459
rect 1755 425 1767 459
rect 1709 391 1767 425
rect 1709 357 1721 391
rect 1755 357 1767 391
rect 1709 323 1767 357
rect 1709 289 1721 323
rect 1755 289 1767 323
rect 1709 255 1767 289
rect 1709 221 1721 255
rect 1755 221 1767 255
rect 1709 187 1767 221
rect 1709 153 1721 187
rect 1755 153 1767 187
rect 1709 119 1767 153
rect 1709 85 1721 119
rect 1755 85 1767 119
rect 1709 51 1767 85
rect 1709 17 1721 51
rect 1755 17 1767 51
rect 1709 -17 1767 17
rect 1709 -51 1721 -17
rect 1755 -51 1767 -17
rect 1709 -85 1767 -51
rect 1709 -119 1721 -85
rect 1755 -119 1767 -85
rect 1709 -153 1767 -119
rect 1709 -187 1721 -153
rect 1755 -187 1767 -153
rect 1709 -221 1767 -187
rect 1709 -255 1721 -221
rect 1755 -255 1767 -221
rect 1709 -289 1767 -255
rect 1709 -323 1721 -289
rect 1755 -323 1767 -289
rect 1709 -357 1767 -323
rect 1709 -391 1721 -357
rect 1755 -391 1767 -357
rect 1709 -425 1767 -391
rect 1709 -459 1721 -425
rect 1755 -459 1767 -425
rect 1709 -500 1767 -459
rect 1867 459 1925 500
rect 1867 425 1879 459
rect 1913 425 1925 459
rect 1867 391 1925 425
rect 1867 357 1879 391
rect 1913 357 1925 391
rect 1867 323 1925 357
rect 1867 289 1879 323
rect 1913 289 1925 323
rect 1867 255 1925 289
rect 1867 221 1879 255
rect 1913 221 1925 255
rect 1867 187 1925 221
rect 1867 153 1879 187
rect 1913 153 1925 187
rect 1867 119 1925 153
rect 1867 85 1879 119
rect 1913 85 1925 119
rect 1867 51 1925 85
rect 1867 17 1879 51
rect 1913 17 1925 51
rect 1867 -17 1925 17
rect 1867 -51 1879 -17
rect 1913 -51 1925 -17
rect 1867 -85 1925 -51
rect 1867 -119 1879 -85
rect 1913 -119 1925 -85
rect 1867 -153 1925 -119
rect 1867 -187 1879 -153
rect 1913 -187 1925 -153
rect 1867 -221 1925 -187
rect 1867 -255 1879 -221
rect 1913 -255 1925 -221
rect 1867 -289 1925 -255
rect 1867 -323 1879 -289
rect 1913 -323 1925 -289
rect 1867 -357 1925 -323
rect 1867 -391 1879 -357
rect 1913 -391 1925 -357
rect 1867 -425 1925 -391
rect 1867 -459 1879 -425
rect 1913 -459 1925 -425
rect 1867 -500 1925 -459
rect 2025 459 2083 500
rect 2025 425 2037 459
rect 2071 425 2083 459
rect 2025 391 2083 425
rect 2025 357 2037 391
rect 2071 357 2083 391
rect 2025 323 2083 357
rect 2025 289 2037 323
rect 2071 289 2083 323
rect 2025 255 2083 289
rect 2025 221 2037 255
rect 2071 221 2083 255
rect 2025 187 2083 221
rect 2025 153 2037 187
rect 2071 153 2083 187
rect 2025 119 2083 153
rect 2025 85 2037 119
rect 2071 85 2083 119
rect 2025 51 2083 85
rect 2025 17 2037 51
rect 2071 17 2083 51
rect 2025 -17 2083 17
rect 2025 -51 2037 -17
rect 2071 -51 2083 -17
rect 2025 -85 2083 -51
rect 2025 -119 2037 -85
rect 2071 -119 2083 -85
rect 2025 -153 2083 -119
rect 2025 -187 2037 -153
rect 2071 -187 2083 -153
rect 2025 -221 2083 -187
rect 2025 -255 2037 -221
rect 2071 -255 2083 -221
rect 2025 -289 2083 -255
rect 2025 -323 2037 -289
rect 2071 -323 2083 -289
rect 2025 -357 2083 -323
rect 2025 -391 2037 -357
rect 2071 -391 2083 -357
rect 2025 -425 2083 -391
rect 2025 -459 2037 -425
rect 2071 -459 2083 -425
rect 2025 -500 2083 -459
rect 2183 459 2241 500
rect 2183 425 2195 459
rect 2229 425 2241 459
rect 2183 391 2241 425
rect 2183 357 2195 391
rect 2229 357 2241 391
rect 2183 323 2241 357
rect 2183 289 2195 323
rect 2229 289 2241 323
rect 2183 255 2241 289
rect 2183 221 2195 255
rect 2229 221 2241 255
rect 2183 187 2241 221
rect 2183 153 2195 187
rect 2229 153 2241 187
rect 2183 119 2241 153
rect 2183 85 2195 119
rect 2229 85 2241 119
rect 2183 51 2241 85
rect 2183 17 2195 51
rect 2229 17 2241 51
rect 2183 -17 2241 17
rect 2183 -51 2195 -17
rect 2229 -51 2241 -17
rect 2183 -85 2241 -51
rect 2183 -119 2195 -85
rect 2229 -119 2241 -85
rect 2183 -153 2241 -119
rect 2183 -187 2195 -153
rect 2229 -187 2241 -153
rect 2183 -221 2241 -187
rect 2183 -255 2195 -221
rect 2229 -255 2241 -221
rect 2183 -289 2241 -255
rect 2183 -323 2195 -289
rect 2229 -323 2241 -289
rect 2183 -357 2241 -323
rect 2183 -391 2195 -357
rect 2229 -391 2241 -357
rect 2183 -425 2241 -391
rect 2183 -459 2195 -425
rect 2229 -459 2241 -425
rect 2183 -500 2241 -459
rect 2341 459 2399 500
rect 2341 425 2353 459
rect 2387 425 2399 459
rect 2341 391 2399 425
rect 2341 357 2353 391
rect 2387 357 2399 391
rect 2341 323 2399 357
rect 2341 289 2353 323
rect 2387 289 2399 323
rect 2341 255 2399 289
rect 2341 221 2353 255
rect 2387 221 2399 255
rect 2341 187 2399 221
rect 2341 153 2353 187
rect 2387 153 2399 187
rect 2341 119 2399 153
rect 2341 85 2353 119
rect 2387 85 2399 119
rect 2341 51 2399 85
rect 2341 17 2353 51
rect 2387 17 2399 51
rect 2341 -17 2399 17
rect 2341 -51 2353 -17
rect 2387 -51 2399 -17
rect 2341 -85 2399 -51
rect 2341 -119 2353 -85
rect 2387 -119 2399 -85
rect 2341 -153 2399 -119
rect 2341 -187 2353 -153
rect 2387 -187 2399 -153
rect 2341 -221 2399 -187
rect 2341 -255 2353 -221
rect 2387 -255 2399 -221
rect 2341 -289 2399 -255
rect 2341 -323 2353 -289
rect 2387 -323 2399 -289
rect 2341 -357 2399 -323
rect 2341 -391 2353 -357
rect 2387 -391 2399 -357
rect 2341 -425 2399 -391
rect 2341 -459 2353 -425
rect 2387 -459 2399 -425
rect 2341 -500 2399 -459
rect 2499 459 2557 500
rect 2499 425 2511 459
rect 2545 425 2557 459
rect 2499 391 2557 425
rect 2499 357 2511 391
rect 2545 357 2557 391
rect 2499 323 2557 357
rect 2499 289 2511 323
rect 2545 289 2557 323
rect 2499 255 2557 289
rect 2499 221 2511 255
rect 2545 221 2557 255
rect 2499 187 2557 221
rect 2499 153 2511 187
rect 2545 153 2557 187
rect 2499 119 2557 153
rect 2499 85 2511 119
rect 2545 85 2557 119
rect 2499 51 2557 85
rect 2499 17 2511 51
rect 2545 17 2557 51
rect 2499 -17 2557 17
rect 2499 -51 2511 -17
rect 2545 -51 2557 -17
rect 2499 -85 2557 -51
rect 2499 -119 2511 -85
rect 2545 -119 2557 -85
rect 2499 -153 2557 -119
rect 2499 -187 2511 -153
rect 2545 -187 2557 -153
rect 2499 -221 2557 -187
rect 2499 -255 2511 -221
rect 2545 -255 2557 -221
rect 2499 -289 2557 -255
rect 2499 -323 2511 -289
rect 2545 -323 2557 -289
rect 2499 -357 2557 -323
rect 2499 -391 2511 -357
rect 2545 -391 2557 -357
rect 2499 -425 2557 -391
rect 2499 -459 2511 -425
rect 2545 -459 2557 -425
rect 2499 -500 2557 -459
rect 2657 459 2715 500
rect 2657 425 2669 459
rect 2703 425 2715 459
rect 2657 391 2715 425
rect 2657 357 2669 391
rect 2703 357 2715 391
rect 2657 323 2715 357
rect 2657 289 2669 323
rect 2703 289 2715 323
rect 2657 255 2715 289
rect 2657 221 2669 255
rect 2703 221 2715 255
rect 2657 187 2715 221
rect 2657 153 2669 187
rect 2703 153 2715 187
rect 2657 119 2715 153
rect 2657 85 2669 119
rect 2703 85 2715 119
rect 2657 51 2715 85
rect 2657 17 2669 51
rect 2703 17 2715 51
rect 2657 -17 2715 17
rect 2657 -51 2669 -17
rect 2703 -51 2715 -17
rect 2657 -85 2715 -51
rect 2657 -119 2669 -85
rect 2703 -119 2715 -85
rect 2657 -153 2715 -119
rect 2657 -187 2669 -153
rect 2703 -187 2715 -153
rect 2657 -221 2715 -187
rect 2657 -255 2669 -221
rect 2703 -255 2715 -221
rect 2657 -289 2715 -255
rect 2657 -323 2669 -289
rect 2703 -323 2715 -289
rect 2657 -357 2715 -323
rect 2657 -391 2669 -357
rect 2703 -391 2715 -357
rect 2657 -425 2715 -391
rect 2657 -459 2669 -425
rect 2703 -459 2715 -425
rect 2657 -500 2715 -459
rect 2815 459 2873 500
rect 2815 425 2827 459
rect 2861 425 2873 459
rect 2815 391 2873 425
rect 2815 357 2827 391
rect 2861 357 2873 391
rect 2815 323 2873 357
rect 2815 289 2827 323
rect 2861 289 2873 323
rect 2815 255 2873 289
rect 2815 221 2827 255
rect 2861 221 2873 255
rect 2815 187 2873 221
rect 2815 153 2827 187
rect 2861 153 2873 187
rect 2815 119 2873 153
rect 2815 85 2827 119
rect 2861 85 2873 119
rect 2815 51 2873 85
rect 2815 17 2827 51
rect 2861 17 2873 51
rect 2815 -17 2873 17
rect 2815 -51 2827 -17
rect 2861 -51 2873 -17
rect 2815 -85 2873 -51
rect 2815 -119 2827 -85
rect 2861 -119 2873 -85
rect 2815 -153 2873 -119
rect 2815 -187 2827 -153
rect 2861 -187 2873 -153
rect 2815 -221 2873 -187
rect 2815 -255 2827 -221
rect 2861 -255 2873 -221
rect 2815 -289 2873 -255
rect 2815 -323 2827 -289
rect 2861 -323 2873 -289
rect 2815 -357 2873 -323
rect 2815 -391 2827 -357
rect 2861 -391 2873 -357
rect 2815 -425 2873 -391
rect 2815 -459 2827 -425
rect 2861 -459 2873 -425
rect 2815 -500 2873 -459
rect 2973 459 3031 500
rect 2973 425 2985 459
rect 3019 425 3031 459
rect 2973 391 3031 425
rect 2973 357 2985 391
rect 3019 357 3031 391
rect 2973 323 3031 357
rect 2973 289 2985 323
rect 3019 289 3031 323
rect 2973 255 3031 289
rect 2973 221 2985 255
rect 3019 221 3031 255
rect 2973 187 3031 221
rect 2973 153 2985 187
rect 3019 153 3031 187
rect 2973 119 3031 153
rect 2973 85 2985 119
rect 3019 85 3031 119
rect 2973 51 3031 85
rect 2973 17 2985 51
rect 3019 17 3031 51
rect 2973 -17 3031 17
rect 2973 -51 2985 -17
rect 3019 -51 3031 -17
rect 2973 -85 3031 -51
rect 2973 -119 2985 -85
rect 3019 -119 3031 -85
rect 2973 -153 3031 -119
rect 2973 -187 2985 -153
rect 3019 -187 3031 -153
rect 2973 -221 3031 -187
rect 2973 -255 2985 -221
rect 3019 -255 3031 -221
rect 2973 -289 3031 -255
rect 2973 -323 2985 -289
rect 3019 -323 3031 -289
rect 2973 -357 3031 -323
rect 2973 -391 2985 -357
rect 3019 -391 3031 -357
rect 2973 -425 3031 -391
rect 2973 -459 2985 -425
rect 3019 -459 3031 -425
rect 2973 -500 3031 -459
rect 3131 459 3189 500
rect 3131 425 3143 459
rect 3177 425 3189 459
rect 3131 391 3189 425
rect 3131 357 3143 391
rect 3177 357 3189 391
rect 3131 323 3189 357
rect 3131 289 3143 323
rect 3177 289 3189 323
rect 3131 255 3189 289
rect 3131 221 3143 255
rect 3177 221 3189 255
rect 3131 187 3189 221
rect 3131 153 3143 187
rect 3177 153 3189 187
rect 3131 119 3189 153
rect 3131 85 3143 119
rect 3177 85 3189 119
rect 3131 51 3189 85
rect 3131 17 3143 51
rect 3177 17 3189 51
rect 3131 -17 3189 17
rect 3131 -51 3143 -17
rect 3177 -51 3189 -17
rect 3131 -85 3189 -51
rect 3131 -119 3143 -85
rect 3177 -119 3189 -85
rect 3131 -153 3189 -119
rect 3131 -187 3143 -153
rect 3177 -187 3189 -153
rect 3131 -221 3189 -187
rect 3131 -255 3143 -221
rect 3177 -255 3189 -221
rect 3131 -289 3189 -255
rect 3131 -323 3143 -289
rect 3177 -323 3189 -289
rect 3131 -357 3189 -323
rect 3131 -391 3143 -357
rect 3177 -391 3189 -357
rect 3131 -425 3189 -391
rect 3131 -459 3143 -425
rect 3177 -459 3189 -425
rect 3131 -500 3189 -459
<< pdiffc >>
rect -3177 425 -3143 459
rect -3177 357 -3143 391
rect -3177 289 -3143 323
rect -3177 221 -3143 255
rect -3177 153 -3143 187
rect -3177 85 -3143 119
rect -3177 17 -3143 51
rect -3177 -51 -3143 -17
rect -3177 -119 -3143 -85
rect -3177 -187 -3143 -153
rect -3177 -255 -3143 -221
rect -3177 -323 -3143 -289
rect -3177 -391 -3143 -357
rect -3177 -459 -3143 -425
rect -3019 425 -2985 459
rect -3019 357 -2985 391
rect -3019 289 -2985 323
rect -3019 221 -2985 255
rect -3019 153 -2985 187
rect -3019 85 -2985 119
rect -3019 17 -2985 51
rect -3019 -51 -2985 -17
rect -3019 -119 -2985 -85
rect -3019 -187 -2985 -153
rect -3019 -255 -2985 -221
rect -3019 -323 -2985 -289
rect -3019 -391 -2985 -357
rect -3019 -459 -2985 -425
rect -2861 425 -2827 459
rect -2861 357 -2827 391
rect -2861 289 -2827 323
rect -2861 221 -2827 255
rect -2861 153 -2827 187
rect -2861 85 -2827 119
rect -2861 17 -2827 51
rect -2861 -51 -2827 -17
rect -2861 -119 -2827 -85
rect -2861 -187 -2827 -153
rect -2861 -255 -2827 -221
rect -2861 -323 -2827 -289
rect -2861 -391 -2827 -357
rect -2861 -459 -2827 -425
rect -2703 425 -2669 459
rect -2703 357 -2669 391
rect -2703 289 -2669 323
rect -2703 221 -2669 255
rect -2703 153 -2669 187
rect -2703 85 -2669 119
rect -2703 17 -2669 51
rect -2703 -51 -2669 -17
rect -2703 -119 -2669 -85
rect -2703 -187 -2669 -153
rect -2703 -255 -2669 -221
rect -2703 -323 -2669 -289
rect -2703 -391 -2669 -357
rect -2703 -459 -2669 -425
rect -2545 425 -2511 459
rect -2545 357 -2511 391
rect -2545 289 -2511 323
rect -2545 221 -2511 255
rect -2545 153 -2511 187
rect -2545 85 -2511 119
rect -2545 17 -2511 51
rect -2545 -51 -2511 -17
rect -2545 -119 -2511 -85
rect -2545 -187 -2511 -153
rect -2545 -255 -2511 -221
rect -2545 -323 -2511 -289
rect -2545 -391 -2511 -357
rect -2545 -459 -2511 -425
rect -2387 425 -2353 459
rect -2387 357 -2353 391
rect -2387 289 -2353 323
rect -2387 221 -2353 255
rect -2387 153 -2353 187
rect -2387 85 -2353 119
rect -2387 17 -2353 51
rect -2387 -51 -2353 -17
rect -2387 -119 -2353 -85
rect -2387 -187 -2353 -153
rect -2387 -255 -2353 -221
rect -2387 -323 -2353 -289
rect -2387 -391 -2353 -357
rect -2387 -459 -2353 -425
rect -2229 425 -2195 459
rect -2229 357 -2195 391
rect -2229 289 -2195 323
rect -2229 221 -2195 255
rect -2229 153 -2195 187
rect -2229 85 -2195 119
rect -2229 17 -2195 51
rect -2229 -51 -2195 -17
rect -2229 -119 -2195 -85
rect -2229 -187 -2195 -153
rect -2229 -255 -2195 -221
rect -2229 -323 -2195 -289
rect -2229 -391 -2195 -357
rect -2229 -459 -2195 -425
rect -2071 425 -2037 459
rect -2071 357 -2037 391
rect -2071 289 -2037 323
rect -2071 221 -2037 255
rect -2071 153 -2037 187
rect -2071 85 -2037 119
rect -2071 17 -2037 51
rect -2071 -51 -2037 -17
rect -2071 -119 -2037 -85
rect -2071 -187 -2037 -153
rect -2071 -255 -2037 -221
rect -2071 -323 -2037 -289
rect -2071 -391 -2037 -357
rect -2071 -459 -2037 -425
rect -1913 425 -1879 459
rect -1913 357 -1879 391
rect -1913 289 -1879 323
rect -1913 221 -1879 255
rect -1913 153 -1879 187
rect -1913 85 -1879 119
rect -1913 17 -1879 51
rect -1913 -51 -1879 -17
rect -1913 -119 -1879 -85
rect -1913 -187 -1879 -153
rect -1913 -255 -1879 -221
rect -1913 -323 -1879 -289
rect -1913 -391 -1879 -357
rect -1913 -459 -1879 -425
rect -1755 425 -1721 459
rect -1755 357 -1721 391
rect -1755 289 -1721 323
rect -1755 221 -1721 255
rect -1755 153 -1721 187
rect -1755 85 -1721 119
rect -1755 17 -1721 51
rect -1755 -51 -1721 -17
rect -1755 -119 -1721 -85
rect -1755 -187 -1721 -153
rect -1755 -255 -1721 -221
rect -1755 -323 -1721 -289
rect -1755 -391 -1721 -357
rect -1755 -459 -1721 -425
rect -1597 425 -1563 459
rect -1597 357 -1563 391
rect -1597 289 -1563 323
rect -1597 221 -1563 255
rect -1597 153 -1563 187
rect -1597 85 -1563 119
rect -1597 17 -1563 51
rect -1597 -51 -1563 -17
rect -1597 -119 -1563 -85
rect -1597 -187 -1563 -153
rect -1597 -255 -1563 -221
rect -1597 -323 -1563 -289
rect -1597 -391 -1563 -357
rect -1597 -459 -1563 -425
rect -1439 425 -1405 459
rect -1439 357 -1405 391
rect -1439 289 -1405 323
rect -1439 221 -1405 255
rect -1439 153 -1405 187
rect -1439 85 -1405 119
rect -1439 17 -1405 51
rect -1439 -51 -1405 -17
rect -1439 -119 -1405 -85
rect -1439 -187 -1405 -153
rect -1439 -255 -1405 -221
rect -1439 -323 -1405 -289
rect -1439 -391 -1405 -357
rect -1439 -459 -1405 -425
rect -1281 425 -1247 459
rect -1281 357 -1247 391
rect -1281 289 -1247 323
rect -1281 221 -1247 255
rect -1281 153 -1247 187
rect -1281 85 -1247 119
rect -1281 17 -1247 51
rect -1281 -51 -1247 -17
rect -1281 -119 -1247 -85
rect -1281 -187 -1247 -153
rect -1281 -255 -1247 -221
rect -1281 -323 -1247 -289
rect -1281 -391 -1247 -357
rect -1281 -459 -1247 -425
rect -1123 425 -1089 459
rect -1123 357 -1089 391
rect -1123 289 -1089 323
rect -1123 221 -1089 255
rect -1123 153 -1089 187
rect -1123 85 -1089 119
rect -1123 17 -1089 51
rect -1123 -51 -1089 -17
rect -1123 -119 -1089 -85
rect -1123 -187 -1089 -153
rect -1123 -255 -1089 -221
rect -1123 -323 -1089 -289
rect -1123 -391 -1089 -357
rect -1123 -459 -1089 -425
rect -965 425 -931 459
rect -965 357 -931 391
rect -965 289 -931 323
rect -965 221 -931 255
rect -965 153 -931 187
rect -965 85 -931 119
rect -965 17 -931 51
rect -965 -51 -931 -17
rect -965 -119 -931 -85
rect -965 -187 -931 -153
rect -965 -255 -931 -221
rect -965 -323 -931 -289
rect -965 -391 -931 -357
rect -965 -459 -931 -425
rect -807 425 -773 459
rect -807 357 -773 391
rect -807 289 -773 323
rect -807 221 -773 255
rect -807 153 -773 187
rect -807 85 -773 119
rect -807 17 -773 51
rect -807 -51 -773 -17
rect -807 -119 -773 -85
rect -807 -187 -773 -153
rect -807 -255 -773 -221
rect -807 -323 -773 -289
rect -807 -391 -773 -357
rect -807 -459 -773 -425
rect -649 425 -615 459
rect -649 357 -615 391
rect -649 289 -615 323
rect -649 221 -615 255
rect -649 153 -615 187
rect -649 85 -615 119
rect -649 17 -615 51
rect -649 -51 -615 -17
rect -649 -119 -615 -85
rect -649 -187 -615 -153
rect -649 -255 -615 -221
rect -649 -323 -615 -289
rect -649 -391 -615 -357
rect -649 -459 -615 -425
rect -491 425 -457 459
rect -491 357 -457 391
rect -491 289 -457 323
rect -491 221 -457 255
rect -491 153 -457 187
rect -491 85 -457 119
rect -491 17 -457 51
rect -491 -51 -457 -17
rect -491 -119 -457 -85
rect -491 -187 -457 -153
rect -491 -255 -457 -221
rect -491 -323 -457 -289
rect -491 -391 -457 -357
rect -491 -459 -457 -425
rect -333 425 -299 459
rect -333 357 -299 391
rect -333 289 -299 323
rect -333 221 -299 255
rect -333 153 -299 187
rect -333 85 -299 119
rect -333 17 -299 51
rect -333 -51 -299 -17
rect -333 -119 -299 -85
rect -333 -187 -299 -153
rect -333 -255 -299 -221
rect -333 -323 -299 -289
rect -333 -391 -299 -357
rect -333 -459 -299 -425
rect -175 425 -141 459
rect -175 357 -141 391
rect -175 289 -141 323
rect -175 221 -141 255
rect -175 153 -141 187
rect -175 85 -141 119
rect -175 17 -141 51
rect -175 -51 -141 -17
rect -175 -119 -141 -85
rect -175 -187 -141 -153
rect -175 -255 -141 -221
rect -175 -323 -141 -289
rect -175 -391 -141 -357
rect -175 -459 -141 -425
rect -17 425 17 459
rect -17 357 17 391
rect -17 289 17 323
rect -17 221 17 255
rect -17 153 17 187
rect -17 85 17 119
rect -17 17 17 51
rect -17 -51 17 -17
rect -17 -119 17 -85
rect -17 -187 17 -153
rect -17 -255 17 -221
rect -17 -323 17 -289
rect -17 -391 17 -357
rect -17 -459 17 -425
rect 141 425 175 459
rect 141 357 175 391
rect 141 289 175 323
rect 141 221 175 255
rect 141 153 175 187
rect 141 85 175 119
rect 141 17 175 51
rect 141 -51 175 -17
rect 141 -119 175 -85
rect 141 -187 175 -153
rect 141 -255 175 -221
rect 141 -323 175 -289
rect 141 -391 175 -357
rect 141 -459 175 -425
rect 299 425 333 459
rect 299 357 333 391
rect 299 289 333 323
rect 299 221 333 255
rect 299 153 333 187
rect 299 85 333 119
rect 299 17 333 51
rect 299 -51 333 -17
rect 299 -119 333 -85
rect 299 -187 333 -153
rect 299 -255 333 -221
rect 299 -323 333 -289
rect 299 -391 333 -357
rect 299 -459 333 -425
rect 457 425 491 459
rect 457 357 491 391
rect 457 289 491 323
rect 457 221 491 255
rect 457 153 491 187
rect 457 85 491 119
rect 457 17 491 51
rect 457 -51 491 -17
rect 457 -119 491 -85
rect 457 -187 491 -153
rect 457 -255 491 -221
rect 457 -323 491 -289
rect 457 -391 491 -357
rect 457 -459 491 -425
rect 615 425 649 459
rect 615 357 649 391
rect 615 289 649 323
rect 615 221 649 255
rect 615 153 649 187
rect 615 85 649 119
rect 615 17 649 51
rect 615 -51 649 -17
rect 615 -119 649 -85
rect 615 -187 649 -153
rect 615 -255 649 -221
rect 615 -323 649 -289
rect 615 -391 649 -357
rect 615 -459 649 -425
rect 773 425 807 459
rect 773 357 807 391
rect 773 289 807 323
rect 773 221 807 255
rect 773 153 807 187
rect 773 85 807 119
rect 773 17 807 51
rect 773 -51 807 -17
rect 773 -119 807 -85
rect 773 -187 807 -153
rect 773 -255 807 -221
rect 773 -323 807 -289
rect 773 -391 807 -357
rect 773 -459 807 -425
rect 931 425 965 459
rect 931 357 965 391
rect 931 289 965 323
rect 931 221 965 255
rect 931 153 965 187
rect 931 85 965 119
rect 931 17 965 51
rect 931 -51 965 -17
rect 931 -119 965 -85
rect 931 -187 965 -153
rect 931 -255 965 -221
rect 931 -323 965 -289
rect 931 -391 965 -357
rect 931 -459 965 -425
rect 1089 425 1123 459
rect 1089 357 1123 391
rect 1089 289 1123 323
rect 1089 221 1123 255
rect 1089 153 1123 187
rect 1089 85 1123 119
rect 1089 17 1123 51
rect 1089 -51 1123 -17
rect 1089 -119 1123 -85
rect 1089 -187 1123 -153
rect 1089 -255 1123 -221
rect 1089 -323 1123 -289
rect 1089 -391 1123 -357
rect 1089 -459 1123 -425
rect 1247 425 1281 459
rect 1247 357 1281 391
rect 1247 289 1281 323
rect 1247 221 1281 255
rect 1247 153 1281 187
rect 1247 85 1281 119
rect 1247 17 1281 51
rect 1247 -51 1281 -17
rect 1247 -119 1281 -85
rect 1247 -187 1281 -153
rect 1247 -255 1281 -221
rect 1247 -323 1281 -289
rect 1247 -391 1281 -357
rect 1247 -459 1281 -425
rect 1405 425 1439 459
rect 1405 357 1439 391
rect 1405 289 1439 323
rect 1405 221 1439 255
rect 1405 153 1439 187
rect 1405 85 1439 119
rect 1405 17 1439 51
rect 1405 -51 1439 -17
rect 1405 -119 1439 -85
rect 1405 -187 1439 -153
rect 1405 -255 1439 -221
rect 1405 -323 1439 -289
rect 1405 -391 1439 -357
rect 1405 -459 1439 -425
rect 1563 425 1597 459
rect 1563 357 1597 391
rect 1563 289 1597 323
rect 1563 221 1597 255
rect 1563 153 1597 187
rect 1563 85 1597 119
rect 1563 17 1597 51
rect 1563 -51 1597 -17
rect 1563 -119 1597 -85
rect 1563 -187 1597 -153
rect 1563 -255 1597 -221
rect 1563 -323 1597 -289
rect 1563 -391 1597 -357
rect 1563 -459 1597 -425
rect 1721 425 1755 459
rect 1721 357 1755 391
rect 1721 289 1755 323
rect 1721 221 1755 255
rect 1721 153 1755 187
rect 1721 85 1755 119
rect 1721 17 1755 51
rect 1721 -51 1755 -17
rect 1721 -119 1755 -85
rect 1721 -187 1755 -153
rect 1721 -255 1755 -221
rect 1721 -323 1755 -289
rect 1721 -391 1755 -357
rect 1721 -459 1755 -425
rect 1879 425 1913 459
rect 1879 357 1913 391
rect 1879 289 1913 323
rect 1879 221 1913 255
rect 1879 153 1913 187
rect 1879 85 1913 119
rect 1879 17 1913 51
rect 1879 -51 1913 -17
rect 1879 -119 1913 -85
rect 1879 -187 1913 -153
rect 1879 -255 1913 -221
rect 1879 -323 1913 -289
rect 1879 -391 1913 -357
rect 1879 -459 1913 -425
rect 2037 425 2071 459
rect 2037 357 2071 391
rect 2037 289 2071 323
rect 2037 221 2071 255
rect 2037 153 2071 187
rect 2037 85 2071 119
rect 2037 17 2071 51
rect 2037 -51 2071 -17
rect 2037 -119 2071 -85
rect 2037 -187 2071 -153
rect 2037 -255 2071 -221
rect 2037 -323 2071 -289
rect 2037 -391 2071 -357
rect 2037 -459 2071 -425
rect 2195 425 2229 459
rect 2195 357 2229 391
rect 2195 289 2229 323
rect 2195 221 2229 255
rect 2195 153 2229 187
rect 2195 85 2229 119
rect 2195 17 2229 51
rect 2195 -51 2229 -17
rect 2195 -119 2229 -85
rect 2195 -187 2229 -153
rect 2195 -255 2229 -221
rect 2195 -323 2229 -289
rect 2195 -391 2229 -357
rect 2195 -459 2229 -425
rect 2353 425 2387 459
rect 2353 357 2387 391
rect 2353 289 2387 323
rect 2353 221 2387 255
rect 2353 153 2387 187
rect 2353 85 2387 119
rect 2353 17 2387 51
rect 2353 -51 2387 -17
rect 2353 -119 2387 -85
rect 2353 -187 2387 -153
rect 2353 -255 2387 -221
rect 2353 -323 2387 -289
rect 2353 -391 2387 -357
rect 2353 -459 2387 -425
rect 2511 425 2545 459
rect 2511 357 2545 391
rect 2511 289 2545 323
rect 2511 221 2545 255
rect 2511 153 2545 187
rect 2511 85 2545 119
rect 2511 17 2545 51
rect 2511 -51 2545 -17
rect 2511 -119 2545 -85
rect 2511 -187 2545 -153
rect 2511 -255 2545 -221
rect 2511 -323 2545 -289
rect 2511 -391 2545 -357
rect 2511 -459 2545 -425
rect 2669 425 2703 459
rect 2669 357 2703 391
rect 2669 289 2703 323
rect 2669 221 2703 255
rect 2669 153 2703 187
rect 2669 85 2703 119
rect 2669 17 2703 51
rect 2669 -51 2703 -17
rect 2669 -119 2703 -85
rect 2669 -187 2703 -153
rect 2669 -255 2703 -221
rect 2669 -323 2703 -289
rect 2669 -391 2703 -357
rect 2669 -459 2703 -425
rect 2827 425 2861 459
rect 2827 357 2861 391
rect 2827 289 2861 323
rect 2827 221 2861 255
rect 2827 153 2861 187
rect 2827 85 2861 119
rect 2827 17 2861 51
rect 2827 -51 2861 -17
rect 2827 -119 2861 -85
rect 2827 -187 2861 -153
rect 2827 -255 2861 -221
rect 2827 -323 2861 -289
rect 2827 -391 2861 -357
rect 2827 -459 2861 -425
rect 2985 425 3019 459
rect 2985 357 3019 391
rect 2985 289 3019 323
rect 2985 221 3019 255
rect 2985 153 3019 187
rect 2985 85 3019 119
rect 2985 17 3019 51
rect 2985 -51 3019 -17
rect 2985 -119 3019 -85
rect 2985 -187 3019 -153
rect 2985 -255 3019 -221
rect 2985 -323 3019 -289
rect 2985 -391 3019 -357
rect 2985 -459 3019 -425
rect 3143 425 3177 459
rect 3143 357 3177 391
rect 3143 289 3177 323
rect 3143 221 3177 255
rect 3143 153 3177 187
rect 3143 85 3177 119
rect 3143 17 3177 51
rect 3143 -51 3177 -17
rect 3143 -119 3177 -85
rect 3143 -187 3177 -153
rect 3143 -255 3177 -221
rect 3143 -323 3177 -289
rect 3143 -391 3177 -357
rect 3143 -459 3177 -425
<< nsubdiff >>
rect -3291 649 -3179 683
rect -3145 649 -3111 683
rect -3077 649 -3043 683
rect -3009 649 -2975 683
rect -2941 649 -2907 683
rect -2873 649 -2839 683
rect -2805 649 -2771 683
rect -2737 649 -2703 683
rect -2669 649 -2635 683
rect -2601 649 -2567 683
rect -2533 649 -2499 683
rect -2465 649 -2431 683
rect -2397 649 -2363 683
rect -2329 649 -2295 683
rect -2261 649 -2227 683
rect -2193 649 -2159 683
rect -2125 649 -2091 683
rect -2057 649 -2023 683
rect -1989 649 -1955 683
rect -1921 649 -1887 683
rect -1853 649 -1819 683
rect -1785 649 -1751 683
rect -1717 649 -1683 683
rect -1649 649 -1615 683
rect -1581 649 -1547 683
rect -1513 649 -1479 683
rect -1445 649 -1411 683
rect -1377 649 -1343 683
rect -1309 649 -1275 683
rect -1241 649 -1207 683
rect -1173 649 -1139 683
rect -1105 649 -1071 683
rect -1037 649 -1003 683
rect -969 649 -935 683
rect -901 649 -867 683
rect -833 649 -799 683
rect -765 649 -731 683
rect -697 649 -663 683
rect -629 649 -595 683
rect -561 649 -527 683
rect -493 649 -459 683
rect -425 649 -391 683
rect -357 649 -323 683
rect -289 649 -255 683
rect -221 649 -187 683
rect -153 649 -119 683
rect -85 649 -51 683
rect -17 649 17 683
rect 51 649 85 683
rect 119 649 153 683
rect 187 649 221 683
rect 255 649 289 683
rect 323 649 357 683
rect 391 649 425 683
rect 459 649 493 683
rect 527 649 561 683
rect 595 649 629 683
rect 663 649 697 683
rect 731 649 765 683
rect 799 649 833 683
rect 867 649 901 683
rect 935 649 969 683
rect 1003 649 1037 683
rect 1071 649 1105 683
rect 1139 649 1173 683
rect 1207 649 1241 683
rect 1275 649 1309 683
rect 1343 649 1377 683
rect 1411 649 1445 683
rect 1479 649 1513 683
rect 1547 649 1581 683
rect 1615 649 1649 683
rect 1683 649 1717 683
rect 1751 649 1785 683
rect 1819 649 1853 683
rect 1887 649 1921 683
rect 1955 649 1989 683
rect 2023 649 2057 683
rect 2091 649 2125 683
rect 2159 649 2193 683
rect 2227 649 2261 683
rect 2295 649 2329 683
rect 2363 649 2397 683
rect 2431 649 2465 683
rect 2499 649 2533 683
rect 2567 649 2601 683
rect 2635 649 2669 683
rect 2703 649 2737 683
rect 2771 649 2805 683
rect 2839 649 2873 683
rect 2907 649 2941 683
rect 2975 649 3009 683
rect 3043 649 3077 683
rect 3111 649 3145 683
rect 3179 649 3291 683
rect -3291 561 -3257 649
rect -3291 493 -3257 527
rect 3257 561 3291 649
rect -3291 425 -3257 459
rect -3291 357 -3257 391
rect -3291 289 -3257 323
rect -3291 221 -3257 255
rect -3291 153 -3257 187
rect -3291 85 -3257 119
rect -3291 17 -3257 51
rect -3291 -51 -3257 -17
rect -3291 -119 -3257 -85
rect -3291 -187 -3257 -153
rect -3291 -255 -3257 -221
rect -3291 -323 -3257 -289
rect -3291 -391 -3257 -357
rect -3291 -459 -3257 -425
rect -3291 -527 -3257 -493
rect 3257 493 3291 527
rect 3257 425 3291 459
rect 3257 357 3291 391
rect 3257 289 3291 323
rect 3257 221 3291 255
rect 3257 153 3291 187
rect 3257 85 3291 119
rect 3257 17 3291 51
rect 3257 -51 3291 -17
rect 3257 -119 3291 -85
rect 3257 -187 3291 -153
rect 3257 -255 3291 -221
rect 3257 -323 3291 -289
rect 3257 -391 3291 -357
rect 3257 -459 3291 -425
rect -3291 -649 -3257 -561
rect 3257 -527 3291 -493
rect 3257 -649 3291 -561
rect -3291 -683 -3179 -649
rect -3145 -683 -3111 -649
rect -3077 -683 -3043 -649
rect -3009 -683 -2975 -649
rect -2941 -683 -2907 -649
rect -2873 -683 -2839 -649
rect -2805 -683 -2771 -649
rect -2737 -683 -2703 -649
rect -2669 -683 -2635 -649
rect -2601 -683 -2567 -649
rect -2533 -683 -2499 -649
rect -2465 -683 -2431 -649
rect -2397 -683 -2363 -649
rect -2329 -683 -2295 -649
rect -2261 -683 -2227 -649
rect -2193 -683 -2159 -649
rect -2125 -683 -2091 -649
rect -2057 -683 -2023 -649
rect -1989 -683 -1955 -649
rect -1921 -683 -1887 -649
rect -1853 -683 -1819 -649
rect -1785 -683 -1751 -649
rect -1717 -683 -1683 -649
rect -1649 -683 -1615 -649
rect -1581 -683 -1547 -649
rect -1513 -683 -1479 -649
rect -1445 -683 -1411 -649
rect -1377 -683 -1343 -649
rect -1309 -683 -1275 -649
rect -1241 -683 -1207 -649
rect -1173 -683 -1139 -649
rect -1105 -683 -1071 -649
rect -1037 -683 -1003 -649
rect -969 -683 -935 -649
rect -901 -683 -867 -649
rect -833 -683 -799 -649
rect -765 -683 -731 -649
rect -697 -683 -663 -649
rect -629 -683 -595 -649
rect -561 -683 -527 -649
rect -493 -683 -459 -649
rect -425 -683 -391 -649
rect -357 -683 -323 -649
rect -289 -683 -255 -649
rect -221 -683 -187 -649
rect -153 -683 -119 -649
rect -85 -683 -51 -649
rect -17 -683 17 -649
rect 51 -683 85 -649
rect 119 -683 153 -649
rect 187 -683 221 -649
rect 255 -683 289 -649
rect 323 -683 357 -649
rect 391 -683 425 -649
rect 459 -683 493 -649
rect 527 -683 561 -649
rect 595 -683 629 -649
rect 663 -683 697 -649
rect 731 -683 765 -649
rect 799 -683 833 -649
rect 867 -683 901 -649
rect 935 -683 969 -649
rect 1003 -683 1037 -649
rect 1071 -683 1105 -649
rect 1139 -683 1173 -649
rect 1207 -683 1241 -649
rect 1275 -683 1309 -649
rect 1343 -683 1377 -649
rect 1411 -683 1445 -649
rect 1479 -683 1513 -649
rect 1547 -683 1581 -649
rect 1615 -683 1649 -649
rect 1683 -683 1717 -649
rect 1751 -683 1785 -649
rect 1819 -683 1853 -649
rect 1887 -683 1921 -649
rect 1955 -683 1989 -649
rect 2023 -683 2057 -649
rect 2091 -683 2125 -649
rect 2159 -683 2193 -649
rect 2227 -683 2261 -649
rect 2295 -683 2329 -649
rect 2363 -683 2397 -649
rect 2431 -683 2465 -649
rect 2499 -683 2533 -649
rect 2567 -683 2601 -649
rect 2635 -683 2669 -649
rect 2703 -683 2737 -649
rect 2771 -683 2805 -649
rect 2839 -683 2873 -649
rect 2907 -683 2941 -649
rect 2975 -683 3009 -649
rect 3043 -683 3077 -649
rect 3111 -683 3145 -649
rect 3179 -683 3291 -649
<< nsubdiffcont >>
rect -3179 649 -3145 683
rect -3111 649 -3077 683
rect -3043 649 -3009 683
rect -2975 649 -2941 683
rect -2907 649 -2873 683
rect -2839 649 -2805 683
rect -2771 649 -2737 683
rect -2703 649 -2669 683
rect -2635 649 -2601 683
rect -2567 649 -2533 683
rect -2499 649 -2465 683
rect -2431 649 -2397 683
rect -2363 649 -2329 683
rect -2295 649 -2261 683
rect -2227 649 -2193 683
rect -2159 649 -2125 683
rect -2091 649 -2057 683
rect -2023 649 -1989 683
rect -1955 649 -1921 683
rect -1887 649 -1853 683
rect -1819 649 -1785 683
rect -1751 649 -1717 683
rect -1683 649 -1649 683
rect -1615 649 -1581 683
rect -1547 649 -1513 683
rect -1479 649 -1445 683
rect -1411 649 -1377 683
rect -1343 649 -1309 683
rect -1275 649 -1241 683
rect -1207 649 -1173 683
rect -1139 649 -1105 683
rect -1071 649 -1037 683
rect -1003 649 -969 683
rect -935 649 -901 683
rect -867 649 -833 683
rect -799 649 -765 683
rect -731 649 -697 683
rect -663 649 -629 683
rect -595 649 -561 683
rect -527 649 -493 683
rect -459 649 -425 683
rect -391 649 -357 683
rect -323 649 -289 683
rect -255 649 -221 683
rect -187 649 -153 683
rect -119 649 -85 683
rect -51 649 -17 683
rect 17 649 51 683
rect 85 649 119 683
rect 153 649 187 683
rect 221 649 255 683
rect 289 649 323 683
rect 357 649 391 683
rect 425 649 459 683
rect 493 649 527 683
rect 561 649 595 683
rect 629 649 663 683
rect 697 649 731 683
rect 765 649 799 683
rect 833 649 867 683
rect 901 649 935 683
rect 969 649 1003 683
rect 1037 649 1071 683
rect 1105 649 1139 683
rect 1173 649 1207 683
rect 1241 649 1275 683
rect 1309 649 1343 683
rect 1377 649 1411 683
rect 1445 649 1479 683
rect 1513 649 1547 683
rect 1581 649 1615 683
rect 1649 649 1683 683
rect 1717 649 1751 683
rect 1785 649 1819 683
rect 1853 649 1887 683
rect 1921 649 1955 683
rect 1989 649 2023 683
rect 2057 649 2091 683
rect 2125 649 2159 683
rect 2193 649 2227 683
rect 2261 649 2295 683
rect 2329 649 2363 683
rect 2397 649 2431 683
rect 2465 649 2499 683
rect 2533 649 2567 683
rect 2601 649 2635 683
rect 2669 649 2703 683
rect 2737 649 2771 683
rect 2805 649 2839 683
rect 2873 649 2907 683
rect 2941 649 2975 683
rect 3009 649 3043 683
rect 3077 649 3111 683
rect 3145 649 3179 683
rect -3291 527 -3257 561
rect 3257 527 3291 561
rect -3291 459 -3257 493
rect -3291 391 -3257 425
rect -3291 323 -3257 357
rect -3291 255 -3257 289
rect -3291 187 -3257 221
rect -3291 119 -3257 153
rect -3291 51 -3257 85
rect -3291 -17 -3257 17
rect -3291 -85 -3257 -51
rect -3291 -153 -3257 -119
rect -3291 -221 -3257 -187
rect -3291 -289 -3257 -255
rect -3291 -357 -3257 -323
rect -3291 -425 -3257 -391
rect -3291 -493 -3257 -459
rect 3257 459 3291 493
rect 3257 391 3291 425
rect 3257 323 3291 357
rect 3257 255 3291 289
rect 3257 187 3291 221
rect 3257 119 3291 153
rect 3257 51 3291 85
rect 3257 -17 3291 17
rect 3257 -85 3291 -51
rect 3257 -153 3291 -119
rect 3257 -221 3291 -187
rect 3257 -289 3291 -255
rect 3257 -357 3291 -323
rect 3257 -425 3291 -391
rect 3257 -493 3291 -459
rect -3291 -561 -3257 -527
rect 3257 -561 3291 -527
rect -3179 -683 -3145 -649
rect -3111 -683 -3077 -649
rect -3043 -683 -3009 -649
rect -2975 -683 -2941 -649
rect -2907 -683 -2873 -649
rect -2839 -683 -2805 -649
rect -2771 -683 -2737 -649
rect -2703 -683 -2669 -649
rect -2635 -683 -2601 -649
rect -2567 -683 -2533 -649
rect -2499 -683 -2465 -649
rect -2431 -683 -2397 -649
rect -2363 -683 -2329 -649
rect -2295 -683 -2261 -649
rect -2227 -683 -2193 -649
rect -2159 -683 -2125 -649
rect -2091 -683 -2057 -649
rect -2023 -683 -1989 -649
rect -1955 -683 -1921 -649
rect -1887 -683 -1853 -649
rect -1819 -683 -1785 -649
rect -1751 -683 -1717 -649
rect -1683 -683 -1649 -649
rect -1615 -683 -1581 -649
rect -1547 -683 -1513 -649
rect -1479 -683 -1445 -649
rect -1411 -683 -1377 -649
rect -1343 -683 -1309 -649
rect -1275 -683 -1241 -649
rect -1207 -683 -1173 -649
rect -1139 -683 -1105 -649
rect -1071 -683 -1037 -649
rect -1003 -683 -969 -649
rect -935 -683 -901 -649
rect -867 -683 -833 -649
rect -799 -683 -765 -649
rect -731 -683 -697 -649
rect -663 -683 -629 -649
rect -595 -683 -561 -649
rect -527 -683 -493 -649
rect -459 -683 -425 -649
rect -391 -683 -357 -649
rect -323 -683 -289 -649
rect -255 -683 -221 -649
rect -187 -683 -153 -649
rect -119 -683 -85 -649
rect -51 -683 -17 -649
rect 17 -683 51 -649
rect 85 -683 119 -649
rect 153 -683 187 -649
rect 221 -683 255 -649
rect 289 -683 323 -649
rect 357 -683 391 -649
rect 425 -683 459 -649
rect 493 -683 527 -649
rect 561 -683 595 -649
rect 629 -683 663 -649
rect 697 -683 731 -649
rect 765 -683 799 -649
rect 833 -683 867 -649
rect 901 -683 935 -649
rect 969 -683 1003 -649
rect 1037 -683 1071 -649
rect 1105 -683 1139 -649
rect 1173 -683 1207 -649
rect 1241 -683 1275 -649
rect 1309 -683 1343 -649
rect 1377 -683 1411 -649
rect 1445 -683 1479 -649
rect 1513 -683 1547 -649
rect 1581 -683 1615 -649
rect 1649 -683 1683 -649
rect 1717 -683 1751 -649
rect 1785 -683 1819 -649
rect 1853 -683 1887 -649
rect 1921 -683 1955 -649
rect 1989 -683 2023 -649
rect 2057 -683 2091 -649
rect 2125 -683 2159 -649
rect 2193 -683 2227 -649
rect 2261 -683 2295 -649
rect 2329 -683 2363 -649
rect 2397 -683 2431 -649
rect 2465 -683 2499 -649
rect 2533 -683 2567 -649
rect 2601 -683 2635 -649
rect 2669 -683 2703 -649
rect 2737 -683 2771 -649
rect 2805 -683 2839 -649
rect 2873 -683 2907 -649
rect 2941 -683 2975 -649
rect 3009 -683 3043 -649
rect 3077 -683 3111 -649
rect 3145 -683 3179 -649
<< poly >>
rect -3131 581 -3031 597
rect -3131 547 -3098 581
rect -3064 547 -3031 581
rect -3131 500 -3031 547
rect -2973 581 -2873 597
rect -2973 547 -2940 581
rect -2906 547 -2873 581
rect -2973 500 -2873 547
rect -2815 581 -2715 597
rect -2815 547 -2782 581
rect -2748 547 -2715 581
rect -2815 500 -2715 547
rect -2657 581 -2557 597
rect -2657 547 -2624 581
rect -2590 547 -2557 581
rect -2657 500 -2557 547
rect -2499 581 -2399 597
rect -2499 547 -2466 581
rect -2432 547 -2399 581
rect -2499 500 -2399 547
rect -2341 581 -2241 597
rect -2341 547 -2308 581
rect -2274 547 -2241 581
rect -2341 500 -2241 547
rect -2183 581 -2083 597
rect -2183 547 -2150 581
rect -2116 547 -2083 581
rect -2183 500 -2083 547
rect -2025 581 -1925 597
rect -2025 547 -1992 581
rect -1958 547 -1925 581
rect -2025 500 -1925 547
rect -1867 581 -1767 597
rect -1867 547 -1834 581
rect -1800 547 -1767 581
rect -1867 500 -1767 547
rect -1709 581 -1609 597
rect -1709 547 -1676 581
rect -1642 547 -1609 581
rect -1709 500 -1609 547
rect -1551 581 -1451 597
rect -1551 547 -1518 581
rect -1484 547 -1451 581
rect -1551 500 -1451 547
rect -1393 581 -1293 597
rect -1393 547 -1360 581
rect -1326 547 -1293 581
rect -1393 500 -1293 547
rect -1235 581 -1135 597
rect -1235 547 -1202 581
rect -1168 547 -1135 581
rect -1235 500 -1135 547
rect -1077 581 -977 597
rect -1077 547 -1044 581
rect -1010 547 -977 581
rect -1077 500 -977 547
rect -919 581 -819 597
rect -919 547 -886 581
rect -852 547 -819 581
rect -919 500 -819 547
rect -761 581 -661 597
rect -761 547 -728 581
rect -694 547 -661 581
rect -761 500 -661 547
rect -603 581 -503 597
rect -603 547 -570 581
rect -536 547 -503 581
rect -603 500 -503 547
rect -445 581 -345 597
rect -445 547 -412 581
rect -378 547 -345 581
rect -445 500 -345 547
rect -287 581 -187 597
rect -287 547 -254 581
rect -220 547 -187 581
rect -287 500 -187 547
rect -129 581 -29 597
rect -129 547 -96 581
rect -62 547 -29 581
rect -129 500 -29 547
rect 29 581 129 597
rect 29 547 62 581
rect 96 547 129 581
rect 29 500 129 547
rect 187 581 287 597
rect 187 547 220 581
rect 254 547 287 581
rect 187 500 287 547
rect 345 581 445 597
rect 345 547 378 581
rect 412 547 445 581
rect 345 500 445 547
rect 503 581 603 597
rect 503 547 536 581
rect 570 547 603 581
rect 503 500 603 547
rect 661 581 761 597
rect 661 547 694 581
rect 728 547 761 581
rect 661 500 761 547
rect 819 581 919 597
rect 819 547 852 581
rect 886 547 919 581
rect 819 500 919 547
rect 977 581 1077 597
rect 977 547 1010 581
rect 1044 547 1077 581
rect 977 500 1077 547
rect 1135 581 1235 597
rect 1135 547 1168 581
rect 1202 547 1235 581
rect 1135 500 1235 547
rect 1293 581 1393 597
rect 1293 547 1326 581
rect 1360 547 1393 581
rect 1293 500 1393 547
rect 1451 581 1551 597
rect 1451 547 1484 581
rect 1518 547 1551 581
rect 1451 500 1551 547
rect 1609 581 1709 597
rect 1609 547 1642 581
rect 1676 547 1709 581
rect 1609 500 1709 547
rect 1767 581 1867 597
rect 1767 547 1800 581
rect 1834 547 1867 581
rect 1767 500 1867 547
rect 1925 581 2025 597
rect 1925 547 1958 581
rect 1992 547 2025 581
rect 1925 500 2025 547
rect 2083 581 2183 597
rect 2083 547 2116 581
rect 2150 547 2183 581
rect 2083 500 2183 547
rect 2241 581 2341 597
rect 2241 547 2274 581
rect 2308 547 2341 581
rect 2241 500 2341 547
rect 2399 581 2499 597
rect 2399 547 2432 581
rect 2466 547 2499 581
rect 2399 500 2499 547
rect 2557 581 2657 597
rect 2557 547 2590 581
rect 2624 547 2657 581
rect 2557 500 2657 547
rect 2715 581 2815 597
rect 2715 547 2748 581
rect 2782 547 2815 581
rect 2715 500 2815 547
rect 2873 581 2973 597
rect 2873 547 2906 581
rect 2940 547 2973 581
rect 2873 500 2973 547
rect 3031 581 3131 597
rect 3031 547 3064 581
rect 3098 547 3131 581
rect 3031 500 3131 547
rect -3131 -547 -3031 -500
rect -3131 -581 -3098 -547
rect -3064 -581 -3031 -547
rect -3131 -597 -3031 -581
rect -2973 -547 -2873 -500
rect -2973 -581 -2940 -547
rect -2906 -581 -2873 -547
rect -2973 -597 -2873 -581
rect -2815 -547 -2715 -500
rect -2815 -581 -2782 -547
rect -2748 -581 -2715 -547
rect -2815 -597 -2715 -581
rect -2657 -547 -2557 -500
rect -2657 -581 -2624 -547
rect -2590 -581 -2557 -547
rect -2657 -597 -2557 -581
rect -2499 -547 -2399 -500
rect -2499 -581 -2466 -547
rect -2432 -581 -2399 -547
rect -2499 -597 -2399 -581
rect -2341 -547 -2241 -500
rect -2341 -581 -2308 -547
rect -2274 -581 -2241 -547
rect -2341 -597 -2241 -581
rect -2183 -547 -2083 -500
rect -2183 -581 -2150 -547
rect -2116 -581 -2083 -547
rect -2183 -597 -2083 -581
rect -2025 -547 -1925 -500
rect -2025 -581 -1992 -547
rect -1958 -581 -1925 -547
rect -2025 -597 -1925 -581
rect -1867 -547 -1767 -500
rect -1867 -581 -1834 -547
rect -1800 -581 -1767 -547
rect -1867 -597 -1767 -581
rect -1709 -547 -1609 -500
rect -1709 -581 -1676 -547
rect -1642 -581 -1609 -547
rect -1709 -597 -1609 -581
rect -1551 -547 -1451 -500
rect -1551 -581 -1518 -547
rect -1484 -581 -1451 -547
rect -1551 -597 -1451 -581
rect -1393 -547 -1293 -500
rect -1393 -581 -1360 -547
rect -1326 -581 -1293 -547
rect -1393 -597 -1293 -581
rect -1235 -547 -1135 -500
rect -1235 -581 -1202 -547
rect -1168 -581 -1135 -547
rect -1235 -597 -1135 -581
rect -1077 -547 -977 -500
rect -1077 -581 -1044 -547
rect -1010 -581 -977 -547
rect -1077 -597 -977 -581
rect -919 -547 -819 -500
rect -919 -581 -886 -547
rect -852 -581 -819 -547
rect -919 -597 -819 -581
rect -761 -547 -661 -500
rect -761 -581 -728 -547
rect -694 -581 -661 -547
rect -761 -597 -661 -581
rect -603 -547 -503 -500
rect -603 -581 -570 -547
rect -536 -581 -503 -547
rect -603 -597 -503 -581
rect -445 -547 -345 -500
rect -445 -581 -412 -547
rect -378 -581 -345 -547
rect -445 -597 -345 -581
rect -287 -547 -187 -500
rect -287 -581 -254 -547
rect -220 -581 -187 -547
rect -287 -597 -187 -581
rect -129 -547 -29 -500
rect -129 -581 -96 -547
rect -62 -581 -29 -547
rect -129 -597 -29 -581
rect 29 -547 129 -500
rect 29 -581 62 -547
rect 96 -581 129 -547
rect 29 -597 129 -581
rect 187 -547 287 -500
rect 187 -581 220 -547
rect 254 -581 287 -547
rect 187 -597 287 -581
rect 345 -547 445 -500
rect 345 -581 378 -547
rect 412 -581 445 -547
rect 345 -597 445 -581
rect 503 -547 603 -500
rect 503 -581 536 -547
rect 570 -581 603 -547
rect 503 -597 603 -581
rect 661 -547 761 -500
rect 661 -581 694 -547
rect 728 -581 761 -547
rect 661 -597 761 -581
rect 819 -547 919 -500
rect 819 -581 852 -547
rect 886 -581 919 -547
rect 819 -597 919 -581
rect 977 -547 1077 -500
rect 977 -581 1010 -547
rect 1044 -581 1077 -547
rect 977 -597 1077 -581
rect 1135 -547 1235 -500
rect 1135 -581 1168 -547
rect 1202 -581 1235 -547
rect 1135 -597 1235 -581
rect 1293 -547 1393 -500
rect 1293 -581 1326 -547
rect 1360 -581 1393 -547
rect 1293 -597 1393 -581
rect 1451 -547 1551 -500
rect 1451 -581 1484 -547
rect 1518 -581 1551 -547
rect 1451 -597 1551 -581
rect 1609 -547 1709 -500
rect 1609 -581 1642 -547
rect 1676 -581 1709 -547
rect 1609 -597 1709 -581
rect 1767 -547 1867 -500
rect 1767 -581 1800 -547
rect 1834 -581 1867 -547
rect 1767 -597 1867 -581
rect 1925 -547 2025 -500
rect 1925 -581 1958 -547
rect 1992 -581 2025 -547
rect 1925 -597 2025 -581
rect 2083 -547 2183 -500
rect 2083 -581 2116 -547
rect 2150 -581 2183 -547
rect 2083 -597 2183 -581
rect 2241 -547 2341 -500
rect 2241 -581 2274 -547
rect 2308 -581 2341 -547
rect 2241 -597 2341 -581
rect 2399 -547 2499 -500
rect 2399 -581 2432 -547
rect 2466 -581 2499 -547
rect 2399 -597 2499 -581
rect 2557 -547 2657 -500
rect 2557 -581 2590 -547
rect 2624 -581 2657 -547
rect 2557 -597 2657 -581
rect 2715 -547 2815 -500
rect 2715 -581 2748 -547
rect 2782 -581 2815 -547
rect 2715 -597 2815 -581
rect 2873 -547 2973 -500
rect 2873 -581 2906 -547
rect 2940 -581 2973 -547
rect 2873 -597 2973 -581
rect 3031 -547 3131 -500
rect 3031 -581 3064 -547
rect 3098 -581 3131 -547
rect 3031 -597 3131 -581
<< polycont >>
rect -3098 547 -3064 581
rect -2940 547 -2906 581
rect -2782 547 -2748 581
rect -2624 547 -2590 581
rect -2466 547 -2432 581
rect -2308 547 -2274 581
rect -2150 547 -2116 581
rect -1992 547 -1958 581
rect -1834 547 -1800 581
rect -1676 547 -1642 581
rect -1518 547 -1484 581
rect -1360 547 -1326 581
rect -1202 547 -1168 581
rect -1044 547 -1010 581
rect -886 547 -852 581
rect -728 547 -694 581
rect -570 547 -536 581
rect -412 547 -378 581
rect -254 547 -220 581
rect -96 547 -62 581
rect 62 547 96 581
rect 220 547 254 581
rect 378 547 412 581
rect 536 547 570 581
rect 694 547 728 581
rect 852 547 886 581
rect 1010 547 1044 581
rect 1168 547 1202 581
rect 1326 547 1360 581
rect 1484 547 1518 581
rect 1642 547 1676 581
rect 1800 547 1834 581
rect 1958 547 1992 581
rect 2116 547 2150 581
rect 2274 547 2308 581
rect 2432 547 2466 581
rect 2590 547 2624 581
rect 2748 547 2782 581
rect 2906 547 2940 581
rect 3064 547 3098 581
rect -3098 -581 -3064 -547
rect -2940 -581 -2906 -547
rect -2782 -581 -2748 -547
rect -2624 -581 -2590 -547
rect -2466 -581 -2432 -547
rect -2308 -581 -2274 -547
rect -2150 -581 -2116 -547
rect -1992 -581 -1958 -547
rect -1834 -581 -1800 -547
rect -1676 -581 -1642 -547
rect -1518 -581 -1484 -547
rect -1360 -581 -1326 -547
rect -1202 -581 -1168 -547
rect -1044 -581 -1010 -547
rect -886 -581 -852 -547
rect -728 -581 -694 -547
rect -570 -581 -536 -547
rect -412 -581 -378 -547
rect -254 -581 -220 -547
rect -96 -581 -62 -547
rect 62 -581 96 -547
rect 220 -581 254 -547
rect 378 -581 412 -547
rect 536 -581 570 -547
rect 694 -581 728 -547
rect 852 -581 886 -547
rect 1010 -581 1044 -547
rect 1168 -581 1202 -547
rect 1326 -581 1360 -547
rect 1484 -581 1518 -547
rect 1642 -581 1676 -547
rect 1800 -581 1834 -547
rect 1958 -581 1992 -547
rect 2116 -581 2150 -547
rect 2274 -581 2308 -547
rect 2432 -581 2466 -547
rect 2590 -581 2624 -547
rect 2748 -581 2782 -547
rect 2906 -581 2940 -547
rect 3064 -581 3098 -547
<< locali >>
rect -3291 649 -3179 683
rect -3145 649 -3111 683
rect -3077 649 -3043 683
rect -3009 649 -2975 683
rect -2941 649 -2907 683
rect -2873 649 -2839 683
rect -2805 649 -2771 683
rect -2737 649 -2703 683
rect -2669 649 -2635 683
rect -2601 649 -2567 683
rect -2533 649 -2499 683
rect -2465 649 -2431 683
rect -2397 649 -2363 683
rect -2329 649 -2295 683
rect -2261 649 -2227 683
rect -2193 649 -2159 683
rect -2125 649 -2091 683
rect -2057 649 -2023 683
rect -1989 649 -1955 683
rect -1921 649 -1887 683
rect -1853 649 -1819 683
rect -1785 649 -1751 683
rect -1717 649 -1683 683
rect -1649 649 -1615 683
rect -1567 649 -1547 683
rect -1495 649 -1479 683
rect -1423 649 -1411 683
rect -1351 649 -1343 683
rect -1279 649 -1275 683
rect -1173 649 -1169 683
rect -1105 649 -1097 683
rect -1037 649 -1025 683
rect -969 649 -953 683
rect -901 649 -881 683
rect -833 649 -809 683
rect -765 649 -737 683
rect -697 649 -665 683
rect -629 649 -595 683
rect -559 649 -527 683
rect -487 649 -459 683
rect -415 649 -391 683
rect -343 649 -323 683
rect -271 649 -255 683
rect -199 649 -187 683
rect -127 649 -119 683
rect -55 649 -51 683
rect 51 649 55 683
rect 119 649 127 683
rect 187 649 199 683
rect 255 649 271 683
rect 323 649 343 683
rect 391 649 415 683
rect 459 649 487 683
rect 527 649 559 683
rect 595 649 629 683
rect 665 649 697 683
rect 737 649 765 683
rect 809 649 833 683
rect 881 649 901 683
rect 953 649 969 683
rect 1025 649 1037 683
rect 1097 649 1105 683
rect 1169 649 1173 683
rect 1275 649 1279 683
rect 1343 649 1351 683
rect 1411 649 1423 683
rect 1479 649 1495 683
rect 1547 649 1567 683
rect 1615 649 1649 683
rect 1683 649 1717 683
rect 1751 649 1785 683
rect 1819 649 1853 683
rect 1887 649 1921 683
rect 1955 649 1989 683
rect 2023 649 2057 683
rect 2091 649 2125 683
rect 2159 649 2193 683
rect 2227 649 2261 683
rect 2295 649 2329 683
rect 2363 649 2397 683
rect 2431 649 2465 683
rect 2499 649 2533 683
rect 2567 649 2601 683
rect 2635 649 2669 683
rect 2703 649 2737 683
rect 2771 649 2805 683
rect 2839 649 2873 683
rect 2907 649 2941 683
rect 2975 649 3009 683
rect 3043 649 3077 683
rect 3111 649 3145 683
rect 3179 649 3291 683
rect -3291 561 -3257 649
rect -3131 547 -3098 581
rect -3064 547 -3031 581
rect -2973 547 -2940 581
rect -2906 547 -2873 581
rect -2815 547 -2782 581
rect -2748 547 -2715 581
rect -2657 547 -2624 581
rect -2590 547 -2557 581
rect -2499 547 -2466 581
rect -2432 547 -2399 581
rect -2341 547 -2308 581
rect -2274 547 -2241 581
rect -2183 547 -2150 581
rect -2116 547 -2083 581
rect -2025 547 -1992 581
rect -1958 547 -1925 581
rect -1867 547 -1834 581
rect -1800 547 -1767 581
rect -1709 547 -1676 581
rect -1642 547 -1609 581
rect -1551 547 -1518 581
rect -1484 547 -1451 581
rect -1393 547 -1360 581
rect -1326 547 -1293 581
rect -1235 547 -1202 581
rect -1168 547 -1135 581
rect -1077 547 -1044 581
rect -1010 547 -977 581
rect -919 547 -886 581
rect -852 547 -819 581
rect -761 547 -728 581
rect -694 547 -661 581
rect -603 547 -570 581
rect -536 547 -503 581
rect -445 547 -412 581
rect -378 547 -345 581
rect -287 547 -254 581
rect -220 547 -187 581
rect -129 547 -96 581
rect -62 547 -29 581
rect 29 547 62 581
rect 96 547 129 581
rect 187 547 220 581
rect 254 547 287 581
rect 345 547 378 581
rect 412 547 445 581
rect 503 547 536 581
rect 570 547 603 581
rect 661 547 694 581
rect 728 547 761 581
rect 819 547 852 581
rect 886 547 919 581
rect 977 547 1010 581
rect 1044 547 1077 581
rect 1135 547 1168 581
rect 1202 547 1235 581
rect 1293 547 1326 581
rect 1360 547 1393 581
rect 1451 547 1484 581
rect 1518 547 1551 581
rect 1609 547 1642 581
rect 1676 547 1709 581
rect 1767 547 1800 581
rect 1834 547 1867 581
rect 1925 547 1958 581
rect 1992 547 2025 581
rect 2083 547 2116 581
rect 2150 547 2183 581
rect 2241 547 2274 581
rect 2308 547 2341 581
rect 2399 547 2432 581
rect 2466 547 2499 581
rect 2557 547 2590 581
rect 2624 547 2657 581
rect 2715 547 2748 581
rect 2782 547 2815 581
rect 2873 547 2906 581
rect 2940 547 2973 581
rect 3031 547 3064 581
rect 3098 547 3131 581
rect 3257 561 3291 649
rect -3291 493 -3257 527
rect -3291 425 -3257 459
rect -3291 357 -3257 391
rect -3291 289 -3257 323
rect -3291 221 -3257 255
rect -3291 153 -3257 187
rect -3291 85 -3257 119
rect -3291 17 -3257 51
rect -3291 -51 -3257 -17
rect -3291 -119 -3257 -85
rect -3291 -187 -3257 -153
rect -3291 -255 -3257 -221
rect -3291 -323 -3257 -289
rect -3291 -391 -3257 -357
rect -3291 -459 -3257 -425
rect -3291 -527 -3257 -493
rect -3177 485 -3143 504
rect -3177 413 -3143 425
rect -3177 341 -3143 357
rect -3177 269 -3143 289
rect -3177 197 -3143 221
rect -3177 125 -3143 153
rect -3177 53 -3143 85
rect -3177 -17 -3143 17
rect -3177 -85 -3143 -53
rect -3177 -153 -3143 -125
rect -3177 -221 -3143 -197
rect -3177 -289 -3143 -269
rect -3177 -357 -3143 -341
rect -3177 -425 -3143 -413
rect -3177 -504 -3143 -485
rect -3019 485 -2985 504
rect -3019 413 -2985 425
rect -3019 341 -2985 357
rect -3019 269 -2985 289
rect -3019 197 -2985 221
rect -3019 125 -2985 153
rect -3019 53 -2985 85
rect -3019 -17 -2985 17
rect -3019 -85 -2985 -53
rect -3019 -153 -2985 -125
rect -3019 -221 -2985 -197
rect -3019 -289 -2985 -269
rect -3019 -357 -2985 -341
rect -3019 -425 -2985 -413
rect -3019 -504 -2985 -485
rect -2861 485 -2827 504
rect -2861 413 -2827 425
rect -2861 341 -2827 357
rect -2861 269 -2827 289
rect -2861 197 -2827 221
rect -2861 125 -2827 153
rect -2861 53 -2827 85
rect -2861 -17 -2827 17
rect -2861 -85 -2827 -53
rect -2861 -153 -2827 -125
rect -2861 -221 -2827 -197
rect -2861 -289 -2827 -269
rect -2861 -357 -2827 -341
rect -2861 -425 -2827 -413
rect -2861 -504 -2827 -485
rect -2703 485 -2669 504
rect -2703 413 -2669 425
rect -2703 341 -2669 357
rect -2703 269 -2669 289
rect -2703 197 -2669 221
rect -2703 125 -2669 153
rect -2703 53 -2669 85
rect -2703 -17 -2669 17
rect -2703 -85 -2669 -53
rect -2703 -153 -2669 -125
rect -2703 -221 -2669 -197
rect -2703 -289 -2669 -269
rect -2703 -357 -2669 -341
rect -2703 -425 -2669 -413
rect -2703 -504 -2669 -485
rect -2545 485 -2511 504
rect -2545 413 -2511 425
rect -2545 341 -2511 357
rect -2545 269 -2511 289
rect -2545 197 -2511 221
rect -2545 125 -2511 153
rect -2545 53 -2511 85
rect -2545 -17 -2511 17
rect -2545 -85 -2511 -53
rect -2545 -153 -2511 -125
rect -2545 -221 -2511 -197
rect -2545 -289 -2511 -269
rect -2545 -357 -2511 -341
rect -2545 -425 -2511 -413
rect -2545 -504 -2511 -485
rect -2387 485 -2353 504
rect -2387 413 -2353 425
rect -2387 341 -2353 357
rect -2387 269 -2353 289
rect -2387 197 -2353 221
rect -2387 125 -2353 153
rect -2387 53 -2353 85
rect -2387 -17 -2353 17
rect -2387 -85 -2353 -53
rect -2387 -153 -2353 -125
rect -2387 -221 -2353 -197
rect -2387 -289 -2353 -269
rect -2387 -357 -2353 -341
rect -2387 -425 -2353 -413
rect -2387 -504 -2353 -485
rect -2229 485 -2195 504
rect -2229 413 -2195 425
rect -2229 341 -2195 357
rect -2229 269 -2195 289
rect -2229 197 -2195 221
rect -2229 125 -2195 153
rect -2229 53 -2195 85
rect -2229 -17 -2195 17
rect -2229 -85 -2195 -53
rect -2229 -153 -2195 -125
rect -2229 -221 -2195 -197
rect -2229 -289 -2195 -269
rect -2229 -357 -2195 -341
rect -2229 -425 -2195 -413
rect -2229 -504 -2195 -485
rect -2071 485 -2037 504
rect -2071 413 -2037 425
rect -2071 341 -2037 357
rect -2071 269 -2037 289
rect -2071 197 -2037 221
rect -2071 125 -2037 153
rect -2071 53 -2037 85
rect -2071 -17 -2037 17
rect -2071 -85 -2037 -53
rect -2071 -153 -2037 -125
rect -2071 -221 -2037 -197
rect -2071 -289 -2037 -269
rect -2071 -357 -2037 -341
rect -2071 -425 -2037 -413
rect -2071 -504 -2037 -485
rect -1913 485 -1879 504
rect -1913 413 -1879 425
rect -1913 341 -1879 357
rect -1913 269 -1879 289
rect -1913 197 -1879 221
rect -1913 125 -1879 153
rect -1913 53 -1879 85
rect -1913 -17 -1879 17
rect -1913 -85 -1879 -53
rect -1913 -153 -1879 -125
rect -1913 -221 -1879 -197
rect -1913 -289 -1879 -269
rect -1913 -357 -1879 -341
rect -1913 -425 -1879 -413
rect -1913 -504 -1879 -485
rect -1755 485 -1721 504
rect -1755 413 -1721 425
rect -1755 341 -1721 357
rect -1755 269 -1721 289
rect -1755 197 -1721 221
rect -1755 125 -1721 153
rect -1755 53 -1721 85
rect -1755 -17 -1721 17
rect -1755 -85 -1721 -53
rect -1755 -153 -1721 -125
rect -1755 -221 -1721 -197
rect -1755 -289 -1721 -269
rect -1755 -357 -1721 -341
rect -1755 -425 -1721 -413
rect -1755 -504 -1721 -485
rect -1597 485 -1563 504
rect -1597 413 -1563 425
rect -1597 341 -1563 357
rect -1597 269 -1563 289
rect -1597 197 -1563 221
rect -1597 125 -1563 153
rect -1597 53 -1563 85
rect -1597 -17 -1563 17
rect -1597 -85 -1563 -53
rect -1597 -153 -1563 -125
rect -1597 -221 -1563 -197
rect -1597 -289 -1563 -269
rect -1597 -357 -1563 -341
rect -1597 -425 -1563 -413
rect -1597 -504 -1563 -485
rect -1439 485 -1405 504
rect -1439 413 -1405 425
rect -1439 341 -1405 357
rect -1439 269 -1405 289
rect -1439 197 -1405 221
rect -1439 125 -1405 153
rect -1439 53 -1405 85
rect -1439 -17 -1405 17
rect -1439 -85 -1405 -53
rect -1439 -153 -1405 -125
rect -1439 -221 -1405 -197
rect -1439 -289 -1405 -269
rect -1439 -357 -1405 -341
rect -1439 -425 -1405 -413
rect -1439 -504 -1405 -485
rect -1281 485 -1247 504
rect -1281 413 -1247 425
rect -1281 341 -1247 357
rect -1281 269 -1247 289
rect -1281 197 -1247 221
rect -1281 125 -1247 153
rect -1281 53 -1247 85
rect -1281 -17 -1247 17
rect -1281 -85 -1247 -53
rect -1281 -153 -1247 -125
rect -1281 -221 -1247 -197
rect -1281 -289 -1247 -269
rect -1281 -357 -1247 -341
rect -1281 -425 -1247 -413
rect -1281 -504 -1247 -485
rect -1123 485 -1089 504
rect -1123 413 -1089 425
rect -1123 341 -1089 357
rect -1123 269 -1089 289
rect -1123 197 -1089 221
rect -1123 125 -1089 153
rect -1123 53 -1089 85
rect -1123 -17 -1089 17
rect -1123 -85 -1089 -53
rect -1123 -153 -1089 -125
rect -1123 -221 -1089 -197
rect -1123 -289 -1089 -269
rect -1123 -357 -1089 -341
rect -1123 -425 -1089 -413
rect -1123 -504 -1089 -485
rect -965 485 -931 504
rect -965 413 -931 425
rect -965 341 -931 357
rect -965 269 -931 289
rect -965 197 -931 221
rect -965 125 -931 153
rect -965 53 -931 85
rect -965 -17 -931 17
rect -965 -85 -931 -53
rect -965 -153 -931 -125
rect -965 -221 -931 -197
rect -965 -289 -931 -269
rect -965 -357 -931 -341
rect -965 -425 -931 -413
rect -965 -504 -931 -485
rect -807 485 -773 504
rect -807 413 -773 425
rect -807 341 -773 357
rect -807 269 -773 289
rect -807 197 -773 221
rect -807 125 -773 153
rect -807 53 -773 85
rect -807 -17 -773 17
rect -807 -85 -773 -53
rect -807 -153 -773 -125
rect -807 -221 -773 -197
rect -807 -289 -773 -269
rect -807 -357 -773 -341
rect -807 -425 -773 -413
rect -807 -504 -773 -485
rect -649 485 -615 504
rect -649 413 -615 425
rect -649 341 -615 357
rect -649 269 -615 289
rect -649 197 -615 221
rect -649 125 -615 153
rect -649 53 -615 85
rect -649 -17 -615 17
rect -649 -85 -615 -53
rect -649 -153 -615 -125
rect -649 -221 -615 -197
rect -649 -289 -615 -269
rect -649 -357 -615 -341
rect -649 -425 -615 -413
rect -649 -504 -615 -485
rect -491 485 -457 504
rect -491 413 -457 425
rect -491 341 -457 357
rect -491 269 -457 289
rect -491 197 -457 221
rect -491 125 -457 153
rect -491 53 -457 85
rect -491 -17 -457 17
rect -491 -85 -457 -53
rect -491 -153 -457 -125
rect -491 -221 -457 -197
rect -491 -289 -457 -269
rect -491 -357 -457 -341
rect -491 -425 -457 -413
rect -491 -504 -457 -485
rect -333 485 -299 504
rect -333 413 -299 425
rect -333 341 -299 357
rect -333 269 -299 289
rect -333 197 -299 221
rect -333 125 -299 153
rect -333 53 -299 85
rect -333 -17 -299 17
rect -333 -85 -299 -53
rect -333 -153 -299 -125
rect -333 -221 -299 -197
rect -333 -289 -299 -269
rect -333 -357 -299 -341
rect -333 -425 -299 -413
rect -333 -504 -299 -485
rect -175 485 -141 504
rect -175 413 -141 425
rect -175 341 -141 357
rect -175 269 -141 289
rect -175 197 -141 221
rect -175 125 -141 153
rect -175 53 -141 85
rect -175 -17 -141 17
rect -175 -85 -141 -53
rect -175 -153 -141 -125
rect -175 -221 -141 -197
rect -175 -289 -141 -269
rect -175 -357 -141 -341
rect -175 -425 -141 -413
rect -175 -504 -141 -485
rect -17 485 17 504
rect -17 413 17 425
rect -17 341 17 357
rect -17 269 17 289
rect -17 197 17 221
rect -17 125 17 153
rect -17 53 17 85
rect -17 -17 17 17
rect -17 -85 17 -53
rect -17 -153 17 -125
rect -17 -221 17 -197
rect -17 -289 17 -269
rect -17 -357 17 -341
rect -17 -425 17 -413
rect -17 -504 17 -485
rect 141 485 175 504
rect 141 413 175 425
rect 141 341 175 357
rect 141 269 175 289
rect 141 197 175 221
rect 141 125 175 153
rect 141 53 175 85
rect 141 -17 175 17
rect 141 -85 175 -53
rect 141 -153 175 -125
rect 141 -221 175 -197
rect 141 -289 175 -269
rect 141 -357 175 -341
rect 141 -425 175 -413
rect 141 -504 175 -485
rect 299 485 333 504
rect 299 413 333 425
rect 299 341 333 357
rect 299 269 333 289
rect 299 197 333 221
rect 299 125 333 153
rect 299 53 333 85
rect 299 -17 333 17
rect 299 -85 333 -53
rect 299 -153 333 -125
rect 299 -221 333 -197
rect 299 -289 333 -269
rect 299 -357 333 -341
rect 299 -425 333 -413
rect 299 -504 333 -485
rect 457 485 491 504
rect 457 413 491 425
rect 457 341 491 357
rect 457 269 491 289
rect 457 197 491 221
rect 457 125 491 153
rect 457 53 491 85
rect 457 -17 491 17
rect 457 -85 491 -53
rect 457 -153 491 -125
rect 457 -221 491 -197
rect 457 -289 491 -269
rect 457 -357 491 -341
rect 457 -425 491 -413
rect 457 -504 491 -485
rect 615 485 649 504
rect 615 413 649 425
rect 615 341 649 357
rect 615 269 649 289
rect 615 197 649 221
rect 615 125 649 153
rect 615 53 649 85
rect 615 -17 649 17
rect 615 -85 649 -53
rect 615 -153 649 -125
rect 615 -221 649 -197
rect 615 -289 649 -269
rect 615 -357 649 -341
rect 615 -425 649 -413
rect 615 -504 649 -485
rect 773 485 807 504
rect 773 413 807 425
rect 773 341 807 357
rect 773 269 807 289
rect 773 197 807 221
rect 773 125 807 153
rect 773 53 807 85
rect 773 -17 807 17
rect 773 -85 807 -53
rect 773 -153 807 -125
rect 773 -221 807 -197
rect 773 -289 807 -269
rect 773 -357 807 -341
rect 773 -425 807 -413
rect 773 -504 807 -485
rect 931 485 965 504
rect 931 413 965 425
rect 931 341 965 357
rect 931 269 965 289
rect 931 197 965 221
rect 931 125 965 153
rect 931 53 965 85
rect 931 -17 965 17
rect 931 -85 965 -53
rect 931 -153 965 -125
rect 931 -221 965 -197
rect 931 -289 965 -269
rect 931 -357 965 -341
rect 931 -425 965 -413
rect 931 -504 965 -485
rect 1089 485 1123 504
rect 1089 413 1123 425
rect 1089 341 1123 357
rect 1089 269 1123 289
rect 1089 197 1123 221
rect 1089 125 1123 153
rect 1089 53 1123 85
rect 1089 -17 1123 17
rect 1089 -85 1123 -53
rect 1089 -153 1123 -125
rect 1089 -221 1123 -197
rect 1089 -289 1123 -269
rect 1089 -357 1123 -341
rect 1089 -425 1123 -413
rect 1089 -504 1123 -485
rect 1247 485 1281 504
rect 1247 413 1281 425
rect 1247 341 1281 357
rect 1247 269 1281 289
rect 1247 197 1281 221
rect 1247 125 1281 153
rect 1247 53 1281 85
rect 1247 -17 1281 17
rect 1247 -85 1281 -53
rect 1247 -153 1281 -125
rect 1247 -221 1281 -197
rect 1247 -289 1281 -269
rect 1247 -357 1281 -341
rect 1247 -425 1281 -413
rect 1247 -504 1281 -485
rect 1405 485 1439 504
rect 1405 413 1439 425
rect 1405 341 1439 357
rect 1405 269 1439 289
rect 1405 197 1439 221
rect 1405 125 1439 153
rect 1405 53 1439 85
rect 1405 -17 1439 17
rect 1405 -85 1439 -53
rect 1405 -153 1439 -125
rect 1405 -221 1439 -197
rect 1405 -289 1439 -269
rect 1405 -357 1439 -341
rect 1405 -425 1439 -413
rect 1405 -504 1439 -485
rect 1563 485 1597 504
rect 1563 413 1597 425
rect 1563 341 1597 357
rect 1563 269 1597 289
rect 1563 197 1597 221
rect 1563 125 1597 153
rect 1563 53 1597 85
rect 1563 -17 1597 17
rect 1563 -85 1597 -53
rect 1563 -153 1597 -125
rect 1563 -221 1597 -197
rect 1563 -289 1597 -269
rect 1563 -357 1597 -341
rect 1563 -425 1597 -413
rect 1563 -504 1597 -485
rect 1721 485 1755 504
rect 1721 413 1755 425
rect 1721 341 1755 357
rect 1721 269 1755 289
rect 1721 197 1755 221
rect 1721 125 1755 153
rect 1721 53 1755 85
rect 1721 -17 1755 17
rect 1721 -85 1755 -53
rect 1721 -153 1755 -125
rect 1721 -221 1755 -197
rect 1721 -289 1755 -269
rect 1721 -357 1755 -341
rect 1721 -425 1755 -413
rect 1721 -504 1755 -485
rect 1879 485 1913 504
rect 1879 413 1913 425
rect 1879 341 1913 357
rect 1879 269 1913 289
rect 1879 197 1913 221
rect 1879 125 1913 153
rect 1879 53 1913 85
rect 1879 -17 1913 17
rect 1879 -85 1913 -53
rect 1879 -153 1913 -125
rect 1879 -221 1913 -197
rect 1879 -289 1913 -269
rect 1879 -357 1913 -341
rect 1879 -425 1913 -413
rect 1879 -504 1913 -485
rect 2037 485 2071 504
rect 2037 413 2071 425
rect 2037 341 2071 357
rect 2037 269 2071 289
rect 2037 197 2071 221
rect 2037 125 2071 153
rect 2037 53 2071 85
rect 2037 -17 2071 17
rect 2037 -85 2071 -53
rect 2037 -153 2071 -125
rect 2037 -221 2071 -197
rect 2037 -289 2071 -269
rect 2037 -357 2071 -341
rect 2037 -425 2071 -413
rect 2037 -504 2071 -485
rect 2195 485 2229 504
rect 2195 413 2229 425
rect 2195 341 2229 357
rect 2195 269 2229 289
rect 2195 197 2229 221
rect 2195 125 2229 153
rect 2195 53 2229 85
rect 2195 -17 2229 17
rect 2195 -85 2229 -53
rect 2195 -153 2229 -125
rect 2195 -221 2229 -197
rect 2195 -289 2229 -269
rect 2195 -357 2229 -341
rect 2195 -425 2229 -413
rect 2195 -504 2229 -485
rect 2353 485 2387 504
rect 2353 413 2387 425
rect 2353 341 2387 357
rect 2353 269 2387 289
rect 2353 197 2387 221
rect 2353 125 2387 153
rect 2353 53 2387 85
rect 2353 -17 2387 17
rect 2353 -85 2387 -53
rect 2353 -153 2387 -125
rect 2353 -221 2387 -197
rect 2353 -289 2387 -269
rect 2353 -357 2387 -341
rect 2353 -425 2387 -413
rect 2353 -504 2387 -485
rect 2511 485 2545 504
rect 2511 413 2545 425
rect 2511 341 2545 357
rect 2511 269 2545 289
rect 2511 197 2545 221
rect 2511 125 2545 153
rect 2511 53 2545 85
rect 2511 -17 2545 17
rect 2511 -85 2545 -53
rect 2511 -153 2545 -125
rect 2511 -221 2545 -197
rect 2511 -289 2545 -269
rect 2511 -357 2545 -341
rect 2511 -425 2545 -413
rect 2511 -504 2545 -485
rect 2669 485 2703 504
rect 2669 413 2703 425
rect 2669 341 2703 357
rect 2669 269 2703 289
rect 2669 197 2703 221
rect 2669 125 2703 153
rect 2669 53 2703 85
rect 2669 -17 2703 17
rect 2669 -85 2703 -53
rect 2669 -153 2703 -125
rect 2669 -221 2703 -197
rect 2669 -289 2703 -269
rect 2669 -357 2703 -341
rect 2669 -425 2703 -413
rect 2669 -504 2703 -485
rect 2827 485 2861 504
rect 2827 413 2861 425
rect 2827 341 2861 357
rect 2827 269 2861 289
rect 2827 197 2861 221
rect 2827 125 2861 153
rect 2827 53 2861 85
rect 2827 -17 2861 17
rect 2827 -85 2861 -53
rect 2827 -153 2861 -125
rect 2827 -221 2861 -197
rect 2827 -289 2861 -269
rect 2827 -357 2861 -341
rect 2827 -425 2861 -413
rect 2827 -504 2861 -485
rect 2985 485 3019 504
rect 2985 413 3019 425
rect 2985 341 3019 357
rect 2985 269 3019 289
rect 2985 197 3019 221
rect 2985 125 3019 153
rect 2985 53 3019 85
rect 2985 -17 3019 17
rect 2985 -85 3019 -53
rect 2985 -153 3019 -125
rect 2985 -221 3019 -197
rect 2985 -289 3019 -269
rect 2985 -357 3019 -341
rect 2985 -425 3019 -413
rect 2985 -504 3019 -485
rect 3143 485 3177 504
rect 3143 413 3177 425
rect 3143 341 3177 357
rect 3143 269 3177 289
rect 3143 197 3177 221
rect 3143 125 3177 153
rect 3143 53 3177 85
rect 3143 -17 3177 17
rect 3143 -85 3177 -53
rect 3143 -153 3177 -125
rect 3143 -221 3177 -197
rect 3143 -289 3177 -269
rect 3143 -357 3177 -341
rect 3143 -425 3177 -413
rect 3143 -504 3177 -485
rect 3257 493 3291 527
rect 3257 425 3291 459
rect 3257 357 3291 391
rect 3257 289 3291 323
rect 3257 221 3291 255
rect 3257 153 3291 187
rect 3257 85 3291 119
rect 3257 17 3291 51
rect 3257 -51 3291 -17
rect 3257 -119 3291 -85
rect 3257 -187 3291 -153
rect 3257 -255 3291 -221
rect 3257 -323 3291 -289
rect 3257 -391 3291 -357
rect 3257 -459 3291 -425
rect 3257 -527 3291 -493
rect -3291 -649 -3257 -561
rect -3131 -581 -3098 -547
rect -3064 -581 -3031 -547
rect -2973 -581 -2940 -547
rect -2906 -581 -2873 -547
rect -2815 -581 -2782 -547
rect -2748 -581 -2715 -547
rect -2657 -581 -2624 -547
rect -2590 -581 -2557 -547
rect -2499 -581 -2466 -547
rect -2432 -581 -2399 -547
rect -2341 -581 -2308 -547
rect -2274 -581 -2241 -547
rect -2183 -581 -2150 -547
rect -2116 -581 -2083 -547
rect -2025 -581 -1992 -547
rect -1958 -581 -1925 -547
rect -1867 -581 -1834 -547
rect -1800 -581 -1767 -547
rect -1709 -581 -1676 -547
rect -1642 -581 -1609 -547
rect -1551 -581 -1518 -547
rect -1484 -581 -1451 -547
rect -1393 -581 -1360 -547
rect -1326 -581 -1293 -547
rect -1235 -581 -1202 -547
rect -1168 -581 -1135 -547
rect -1077 -581 -1044 -547
rect -1010 -581 -977 -547
rect -919 -581 -886 -547
rect -852 -581 -819 -547
rect -761 -581 -728 -547
rect -694 -581 -661 -547
rect -603 -581 -570 -547
rect -536 -581 -503 -547
rect -445 -581 -412 -547
rect -378 -581 -345 -547
rect -287 -581 -254 -547
rect -220 -581 -187 -547
rect -129 -581 -96 -547
rect -62 -581 -29 -547
rect 29 -581 62 -547
rect 96 -581 129 -547
rect 187 -581 220 -547
rect 254 -581 287 -547
rect 345 -581 378 -547
rect 412 -581 445 -547
rect 503 -581 536 -547
rect 570 -581 603 -547
rect 661 -581 694 -547
rect 728 -581 761 -547
rect 819 -581 852 -547
rect 886 -581 919 -547
rect 977 -581 1010 -547
rect 1044 -581 1077 -547
rect 1135 -581 1168 -547
rect 1202 -581 1235 -547
rect 1293 -581 1326 -547
rect 1360 -581 1393 -547
rect 1451 -581 1484 -547
rect 1518 -581 1551 -547
rect 1609 -581 1642 -547
rect 1676 -581 1709 -547
rect 1767 -581 1800 -547
rect 1834 -581 1867 -547
rect 1925 -581 1958 -547
rect 1992 -581 2025 -547
rect 2083 -581 2116 -547
rect 2150 -581 2183 -547
rect 2241 -581 2274 -547
rect 2308 -581 2341 -547
rect 2399 -581 2432 -547
rect 2466 -581 2499 -547
rect 2557 -581 2590 -547
rect 2624 -581 2657 -547
rect 2715 -581 2748 -547
rect 2782 -581 2815 -547
rect 2873 -581 2906 -547
rect 2940 -581 2973 -547
rect 3031 -581 3064 -547
rect 3098 -581 3131 -547
rect 3257 -649 3291 -561
rect -3291 -683 -3179 -649
rect -3145 -683 -3111 -649
rect -3077 -683 -3043 -649
rect -3009 -683 -2975 -649
rect -2941 -683 -2907 -649
rect -2873 -683 -2839 -649
rect -2805 -683 -2771 -649
rect -2737 -683 -2703 -649
rect -2669 -683 -2635 -649
rect -2601 -683 -2567 -649
rect -2533 -683 -2499 -649
rect -2465 -683 -2431 -649
rect -2397 -683 -2363 -649
rect -2329 -683 -2295 -649
rect -2261 -683 -2227 -649
rect -2193 -683 -2159 -649
rect -2125 -683 -2091 -649
rect -2057 -683 -2023 -649
rect -1989 -683 -1955 -649
rect -1921 -683 -1887 -649
rect -1853 -683 -1819 -649
rect -1785 -683 -1751 -649
rect -1717 -683 -1683 -649
rect -1649 -683 -1615 -649
rect -1567 -683 -1547 -649
rect -1495 -683 -1479 -649
rect -1423 -683 -1411 -649
rect -1351 -683 -1343 -649
rect -1279 -683 -1275 -649
rect -1173 -683 -1169 -649
rect -1105 -683 -1097 -649
rect -1037 -683 -1025 -649
rect -969 -683 -953 -649
rect -901 -683 -881 -649
rect -833 -683 -809 -649
rect -765 -683 -737 -649
rect -697 -683 -665 -649
rect -629 -683 -595 -649
rect -559 -683 -527 -649
rect -487 -683 -459 -649
rect -415 -683 -391 -649
rect -343 -683 -323 -649
rect -271 -683 -255 -649
rect -199 -683 -187 -649
rect -127 -683 -119 -649
rect -55 -683 -51 -649
rect 51 -683 55 -649
rect 119 -683 127 -649
rect 187 -683 199 -649
rect 255 -683 271 -649
rect 323 -683 343 -649
rect 391 -683 415 -649
rect 459 -683 487 -649
rect 527 -683 559 -649
rect 595 -683 629 -649
rect 665 -683 697 -649
rect 737 -683 765 -649
rect 809 -683 833 -649
rect 881 -683 901 -649
rect 953 -683 969 -649
rect 1025 -683 1037 -649
rect 1097 -683 1105 -649
rect 1169 -683 1173 -649
rect 1275 -683 1279 -649
rect 1343 -683 1351 -649
rect 1411 -683 1423 -649
rect 1479 -683 1495 -649
rect 1547 -683 1567 -649
rect 1615 -683 1649 -649
rect 1683 -683 1717 -649
rect 1751 -683 1785 -649
rect 1819 -683 1853 -649
rect 1887 -683 1921 -649
rect 1955 -683 1989 -649
rect 2023 -683 2057 -649
rect 2091 -683 2125 -649
rect 2159 -683 2193 -649
rect 2227 -683 2261 -649
rect 2295 -683 2329 -649
rect 2363 -683 2397 -649
rect 2431 -683 2465 -649
rect 2499 -683 2533 -649
rect 2567 -683 2601 -649
rect 2635 -683 2669 -649
rect 2703 -683 2737 -649
rect 2771 -683 2805 -649
rect 2839 -683 2873 -649
rect 2907 -683 2941 -649
rect 2975 -683 3009 -649
rect 3043 -683 3077 -649
rect 3111 -683 3145 -649
rect 3179 -683 3291 -649
<< viali >>
rect -1601 649 -1581 683
rect -1581 649 -1567 683
rect -1529 649 -1513 683
rect -1513 649 -1495 683
rect -1457 649 -1445 683
rect -1445 649 -1423 683
rect -1385 649 -1377 683
rect -1377 649 -1351 683
rect -1313 649 -1309 683
rect -1309 649 -1279 683
rect -1241 649 -1207 683
rect -1169 649 -1139 683
rect -1139 649 -1135 683
rect -1097 649 -1071 683
rect -1071 649 -1063 683
rect -1025 649 -1003 683
rect -1003 649 -991 683
rect -953 649 -935 683
rect -935 649 -919 683
rect -881 649 -867 683
rect -867 649 -847 683
rect -809 649 -799 683
rect -799 649 -775 683
rect -737 649 -731 683
rect -731 649 -703 683
rect -665 649 -663 683
rect -663 649 -631 683
rect -593 649 -561 683
rect -561 649 -559 683
rect -521 649 -493 683
rect -493 649 -487 683
rect -449 649 -425 683
rect -425 649 -415 683
rect -377 649 -357 683
rect -357 649 -343 683
rect -305 649 -289 683
rect -289 649 -271 683
rect -233 649 -221 683
rect -221 649 -199 683
rect -161 649 -153 683
rect -153 649 -127 683
rect -89 649 -85 683
rect -85 649 -55 683
rect -17 649 17 683
rect 55 649 85 683
rect 85 649 89 683
rect 127 649 153 683
rect 153 649 161 683
rect 199 649 221 683
rect 221 649 233 683
rect 271 649 289 683
rect 289 649 305 683
rect 343 649 357 683
rect 357 649 377 683
rect 415 649 425 683
rect 425 649 449 683
rect 487 649 493 683
rect 493 649 521 683
rect 559 649 561 683
rect 561 649 593 683
rect 631 649 663 683
rect 663 649 665 683
rect 703 649 731 683
rect 731 649 737 683
rect 775 649 799 683
rect 799 649 809 683
rect 847 649 867 683
rect 867 649 881 683
rect 919 649 935 683
rect 935 649 953 683
rect 991 649 1003 683
rect 1003 649 1025 683
rect 1063 649 1071 683
rect 1071 649 1097 683
rect 1135 649 1139 683
rect 1139 649 1169 683
rect 1207 649 1241 683
rect 1279 649 1309 683
rect 1309 649 1313 683
rect 1351 649 1377 683
rect 1377 649 1385 683
rect 1423 649 1445 683
rect 1445 649 1457 683
rect 1495 649 1513 683
rect 1513 649 1529 683
rect 1567 649 1581 683
rect 1581 649 1601 683
rect -3098 547 -3064 581
rect -2940 547 -2906 581
rect -2782 547 -2748 581
rect -2624 547 -2590 581
rect -2466 547 -2432 581
rect -2308 547 -2274 581
rect -2150 547 -2116 581
rect -1992 547 -1958 581
rect -1834 547 -1800 581
rect -1676 547 -1642 581
rect -1518 547 -1484 581
rect -1360 547 -1326 581
rect -1202 547 -1168 581
rect -1044 547 -1010 581
rect -886 547 -852 581
rect -728 547 -694 581
rect -570 547 -536 581
rect -412 547 -378 581
rect -254 547 -220 581
rect -96 547 -62 581
rect 62 547 96 581
rect 220 547 254 581
rect 378 547 412 581
rect 536 547 570 581
rect 694 547 728 581
rect 852 547 886 581
rect 1010 547 1044 581
rect 1168 547 1202 581
rect 1326 547 1360 581
rect 1484 547 1518 581
rect 1642 547 1676 581
rect 1800 547 1834 581
rect 1958 547 1992 581
rect 2116 547 2150 581
rect 2274 547 2308 581
rect 2432 547 2466 581
rect 2590 547 2624 581
rect 2748 547 2782 581
rect 2906 547 2940 581
rect 3064 547 3098 581
rect -3177 459 -3143 485
rect -3177 451 -3143 459
rect -3177 391 -3143 413
rect -3177 379 -3143 391
rect -3177 323 -3143 341
rect -3177 307 -3143 323
rect -3177 255 -3143 269
rect -3177 235 -3143 255
rect -3177 187 -3143 197
rect -3177 163 -3143 187
rect -3177 119 -3143 125
rect -3177 91 -3143 119
rect -3177 51 -3143 53
rect -3177 19 -3143 51
rect -3177 -51 -3143 -19
rect -3177 -53 -3143 -51
rect -3177 -119 -3143 -91
rect -3177 -125 -3143 -119
rect -3177 -187 -3143 -163
rect -3177 -197 -3143 -187
rect -3177 -255 -3143 -235
rect -3177 -269 -3143 -255
rect -3177 -323 -3143 -307
rect -3177 -341 -3143 -323
rect -3177 -391 -3143 -379
rect -3177 -413 -3143 -391
rect -3177 -459 -3143 -451
rect -3177 -485 -3143 -459
rect -3019 459 -2985 485
rect -3019 451 -2985 459
rect -3019 391 -2985 413
rect -3019 379 -2985 391
rect -3019 323 -2985 341
rect -3019 307 -2985 323
rect -3019 255 -2985 269
rect -3019 235 -2985 255
rect -3019 187 -2985 197
rect -3019 163 -2985 187
rect -3019 119 -2985 125
rect -3019 91 -2985 119
rect -3019 51 -2985 53
rect -3019 19 -2985 51
rect -3019 -51 -2985 -19
rect -3019 -53 -2985 -51
rect -3019 -119 -2985 -91
rect -3019 -125 -2985 -119
rect -3019 -187 -2985 -163
rect -3019 -197 -2985 -187
rect -3019 -255 -2985 -235
rect -3019 -269 -2985 -255
rect -3019 -323 -2985 -307
rect -3019 -341 -2985 -323
rect -3019 -391 -2985 -379
rect -3019 -413 -2985 -391
rect -3019 -459 -2985 -451
rect -3019 -485 -2985 -459
rect -2861 459 -2827 485
rect -2861 451 -2827 459
rect -2861 391 -2827 413
rect -2861 379 -2827 391
rect -2861 323 -2827 341
rect -2861 307 -2827 323
rect -2861 255 -2827 269
rect -2861 235 -2827 255
rect -2861 187 -2827 197
rect -2861 163 -2827 187
rect -2861 119 -2827 125
rect -2861 91 -2827 119
rect -2861 51 -2827 53
rect -2861 19 -2827 51
rect -2861 -51 -2827 -19
rect -2861 -53 -2827 -51
rect -2861 -119 -2827 -91
rect -2861 -125 -2827 -119
rect -2861 -187 -2827 -163
rect -2861 -197 -2827 -187
rect -2861 -255 -2827 -235
rect -2861 -269 -2827 -255
rect -2861 -323 -2827 -307
rect -2861 -341 -2827 -323
rect -2861 -391 -2827 -379
rect -2861 -413 -2827 -391
rect -2861 -459 -2827 -451
rect -2861 -485 -2827 -459
rect -2703 459 -2669 485
rect -2703 451 -2669 459
rect -2703 391 -2669 413
rect -2703 379 -2669 391
rect -2703 323 -2669 341
rect -2703 307 -2669 323
rect -2703 255 -2669 269
rect -2703 235 -2669 255
rect -2703 187 -2669 197
rect -2703 163 -2669 187
rect -2703 119 -2669 125
rect -2703 91 -2669 119
rect -2703 51 -2669 53
rect -2703 19 -2669 51
rect -2703 -51 -2669 -19
rect -2703 -53 -2669 -51
rect -2703 -119 -2669 -91
rect -2703 -125 -2669 -119
rect -2703 -187 -2669 -163
rect -2703 -197 -2669 -187
rect -2703 -255 -2669 -235
rect -2703 -269 -2669 -255
rect -2703 -323 -2669 -307
rect -2703 -341 -2669 -323
rect -2703 -391 -2669 -379
rect -2703 -413 -2669 -391
rect -2703 -459 -2669 -451
rect -2703 -485 -2669 -459
rect -2545 459 -2511 485
rect -2545 451 -2511 459
rect -2545 391 -2511 413
rect -2545 379 -2511 391
rect -2545 323 -2511 341
rect -2545 307 -2511 323
rect -2545 255 -2511 269
rect -2545 235 -2511 255
rect -2545 187 -2511 197
rect -2545 163 -2511 187
rect -2545 119 -2511 125
rect -2545 91 -2511 119
rect -2545 51 -2511 53
rect -2545 19 -2511 51
rect -2545 -51 -2511 -19
rect -2545 -53 -2511 -51
rect -2545 -119 -2511 -91
rect -2545 -125 -2511 -119
rect -2545 -187 -2511 -163
rect -2545 -197 -2511 -187
rect -2545 -255 -2511 -235
rect -2545 -269 -2511 -255
rect -2545 -323 -2511 -307
rect -2545 -341 -2511 -323
rect -2545 -391 -2511 -379
rect -2545 -413 -2511 -391
rect -2545 -459 -2511 -451
rect -2545 -485 -2511 -459
rect -2387 459 -2353 485
rect -2387 451 -2353 459
rect -2387 391 -2353 413
rect -2387 379 -2353 391
rect -2387 323 -2353 341
rect -2387 307 -2353 323
rect -2387 255 -2353 269
rect -2387 235 -2353 255
rect -2387 187 -2353 197
rect -2387 163 -2353 187
rect -2387 119 -2353 125
rect -2387 91 -2353 119
rect -2387 51 -2353 53
rect -2387 19 -2353 51
rect -2387 -51 -2353 -19
rect -2387 -53 -2353 -51
rect -2387 -119 -2353 -91
rect -2387 -125 -2353 -119
rect -2387 -187 -2353 -163
rect -2387 -197 -2353 -187
rect -2387 -255 -2353 -235
rect -2387 -269 -2353 -255
rect -2387 -323 -2353 -307
rect -2387 -341 -2353 -323
rect -2387 -391 -2353 -379
rect -2387 -413 -2353 -391
rect -2387 -459 -2353 -451
rect -2387 -485 -2353 -459
rect -2229 459 -2195 485
rect -2229 451 -2195 459
rect -2229 391 -2195 413
rect -2229 379 -2195 391
rect -2229 323 -2195 341
rect -2229 307 -2195 323
rect -2229 255 -2195 269
rect -2229 235 -2195 255
rect -2229 187 -2195 197
rect -2229 163 -2195 187
rect -2229 119 -2195 125
rect -2229 91 -2195 119
rect -2229 51 -2195 53
rect -2229 19 -2195 51
rect -2229 -51 -2195 -19
rect -2229 -53 -2195 -51
rect -2229 -119 -2195 -91
rect -2229 -125 -2195 -119
rect -2229 -187 -2195 -163
rect -2229 -197 -2195 -187
rect -2229 -255 -2195 -235
rect -2229 -269 -2195 -255
rect -2229 -323 -2195 -307
rect -2229 -341 -2195 -323
rect -2229 -391 -2195 -379
rect -2229 -413 -2195 -391
rect -2229 -459 -2195 -451
rect -2229 -485 -2195 -459
rect -2071 459 -2037 485
rect -2071 451 -2037 459
rect -2071 391 -2037 413
rect -2071 379 -2037 391
rect -2071 323 -2037 341
rect -2071 307 -2037 323
rect -2071 255 -2037 269
rect -2071 235 -2037 255
rect -2071 187 -2037 197
rect -2071 163 -2037 187
rect -2071 119 -2037 125
rect -2071 91 -2037 119
rect -2071 51 -2037 53
rect -2071 19 -2037 51
rect -2071 -51 -2037 -19
rect -2071 -53 -2037 -51
rect -2071 -119 -2037 -91
rect -2071 -125 -2037 -119
rect -2071 -187 -2037 -163
rect -2071 -197 -2037 -187
rect -2071 -255 -2037 -235
rect -2071 -269 -2037 -255
rect -2071 -323 -2037 -307
rect -2071 -341 -2037 -323
rect -2071 -391 -2037 -379
rect -2071 -413 -2037 -391
rect -2071 -459 -2037 -451
rect -2071 -485 -2037 -459
rect -1913 459 -1879 485
rect -1913 451 -1879 459
rect -1913 391 -1879 413
rect -1913 379 -1879 391
rect -1913 323 -1879 341
rect -1913 307 -1879 323
rect -1913 255 -1879 269
rect -1913 235 -1879 255
rect -1913 187 -1879 197
rect -1913 163 -1879 187
rect -1913 119 -1879 125
rect -1913 91 -1879 119
rect -1913 51 -1879 53
rect -1913 19 -1879 51
rect -1913 -51 -1879 -19
rect -1913 -53 -1879 -51
rect -1913 -119 -1879 -91
rect -1913 -125 -1879 -119
rect -1913 -187 -1879 -163
rect -1913 -197 -1879 -187
rect -1913 -255 -1879 -235
rect -1913 -269 -1879 -255
rect -1913 -323 -1879 -307
rect -1913 -341 -1879 -323
rect -1913 -391 -1879 -379
rect -1913 -413 -1879 -391
rect -1913 -459 -1879 -451
rect -1913 -485 -1879 -459
rect -1755 459 -1721 485
rect -1755 451 -1721 459
rect -1755 391 -1721 413
rect -1755 379 -1721 391
rect -1755 323 -1721 341
rect -1755 307 -1721 323
rect -1755 255 -1721 269
rect -1755 235 -1721 255
rect -1755 187 -1721 197
rect -1755 163 -1721 187
rect -1755 119 -1721 125
rect -1755 91 -1721 119
rect -1755 51 -1721 53
rect -1755 19 -1721 51
rect -1755 -51 -1721 -19
rect -1755 -53 -1721 -51
rect -1755 -119 -1721 -91
rect -1755 -125 -1721 -119
rect -1755 -187 -1721 -163
rect -1755 -197 -1721 -187
rect -1755 -255 -1721 -235
rect -1755 -269 -1721 -255
rect -1755 -323 -1721 -307
rect -1755 -341 -1721 -323
rect -1755 -391 -1721 -379
rect -1755 -413 -1721 -391
rect -1755 -459 -1721 -451
rect -1755 -485 -1721 -459
rect -1597 459 -1563 485
rect -1597 451 -1563 459
rect -1597 391 -1563 413
rect -1597 379 -1563 391
rect -1597 323 -1563 341
rect -1597 307 -1563 323
rect -1597 255 -1563 269
rect -1597 235 -1563 255
rect -1597 187 -1563 197
rect -1597 163 -1563 187
rect -1597 119 -1563 125
rect -1597 91 -1563 119
rect -1597 51 -1563 53
rect -1597 19 -1563 51
rect -1597 -51 -1563 -19
rect -1597 -53 -1563 -51
rect -1597 -119 -1563 -91
rect -1597 -125 -1563 -119
rect -1597 -187 -1563 -163
rect -1597 -197 -1563 -187
rect -1597 -255 -1563 -235
rect -1597 -269 -1563 -255
rect -1597 -323 -1563 -307
rect -1597 -341 -1563 -323
rect -1597 -391 -1563 -379
rect -1597 -413 -1563 -391
rect -1597 -459 -1563 -451
rect -1597 -485 -1563 -459
rect -1439 459 -1405 485
rect -1439 451 -1405 459
rect -1439 391 -1405 413
rect -1439 379 -1405 391
rect -1439 323 -1405 341
rect -1439 307 -1405 323
rect -1439 255 -1405 269
rect -1439 235 -1405 255
rect -1439 187 -1405 197
rect -1439 163 -1405 187
rect -1439 119 -1405 125
rect -1439 91 -1405 119
rect -1439 51 -1405 53
rect -1439 19 -1405 51
rect -1439 -51 -1405 -19
rect -1439 -53 -1405 -51
rect -1439 -119 -1405 -91
rect -1439 -125 -1405 -119
rect -1439 -187 -1405 -163
rect -1439 -197 -1405 -187
rect -1439 -255 -1405 -235
rect -1439 -269 -1405 -255
rect -1439 -323 -1405 -307
rect -1439 -341 -1405 -323
rect -1439 -391 -1405 -379
rect -1439 -413 -1405 -391
rect -1439 -459 -1405 -451
rect -1439 -485 -1405 -459
rect -1281 459 -1247 485
rect -1281 451 -1247 459
rect -1281 391 -1247 413
rect -1281 379 -1247 391
rect -1281 323 -1247 341
rect -1281 307 -1247 323
rect -1281 255 -1247 269
rect -1281 235 -1247 255
rect -1281 187 -1247 197
rect -1281 163 -1247 187
rect -1281 119 -1247 125
rect -1281 91 -1247 119
rect -1281 51 -1247 53
rect -1281 19 -1247 51
rect -1281 -51 -1247 -19
rect -1281 -53 -1247 -51
rect -1281 -119 -1247 -91
rect -1281 -125 -1247 -119
rect -1281 -187 -1247 -163
rect -1281 -197 -1247 -187
rect -1281 -255 -1247 -235
rect -1281 -269 -1247 -255
rect -1281 -323 -1247 -307
rect -1281 -341 -1247 -323
rect -1281 -391 -1247 -379
rect -1281 -413 -1247 -391
rect -1281 -459 -1247 -451
rect -1281 -485 -1247 -459
rect -1123 459 -1089 485
rect -1123 451 -1089 459
rect -1123 391 -1089 413
rect -1123 379 -1089 391
rect -1123 323 -1089 341
rect -1123 307 -1089 323
rect -1123 255 -1089 269
rect -1123 235 -1089 255
rect -1123 187 -1089 197
rect -1123 163 -1089 187
rect -1123 119 -1089 125
rect -1123 91 -1089 119
rect -1123 51 -1089 53
rect -1123 19 -1089 51
rect -1123 -51 -1089 -19
rect -1123 -53 -1089 -51
rect -1123 -119 -1089 -91
rect -1123 -125 -1089 -119
rect -1123 -187 -1089 -163
rect -1123 -197 -1089 -187
rect -1123 -255 -1089 -235
rect -1123 -269 -1089 -255
rect -1123 -323 -1089 -307
rect -1123 -341 -1089 -323
rect -1123 -391 -1089 -379
rect -1123 -413 -1089 -391
rect -1123 -459 -1089 -451
rect -1123 -485 -1089 -459
rect -965 459 -931 485
rect -965 451 -931 459
rect -965 391 -931 413
rect -965 379 -931 391
rect -965 323 -931 341
rect -965 307 -931 323
rect -965 255 -931 269
rect -965 235 -931 255
rect -965 187 -931 197
rect -965 163 -931 187
rect -965 119 -931 125
rect -965 91 -931 119
rect -965 51 -931 53
rect -965 19 -931 51
rect -965 -51 -931 -19
rect -965 -53 -931 -51
rect -965 -119 -931 -91
rect -965 -125 -931 -119
rect -965 -187 -931 -163
rect -965 -197 -931 -187
rect -965 -255 -931 -235
rect -965 -269 -931 -255
rect -965 -323 -931 -307
rect -965 -341 -931 -323
rect -965 -391 -931 -379
rect -965 -413 -931 -391
rect -965 -459 -931 -451
rect -965 -485 -931 -459
rect -807 459 -773 485
rect -807 451 -773 459
rect -807 391 -773 413
rect -807 379 -773 391
rect -807 323 -773 341
rect -807 307 -773 323
rect -807 255 -773 269
rect -807 235 -773 255
rect -807 187 -773 197
rect -807 163 -773 187
rect -807 119 -773 125
rect -807 91 -773 119
rect -807 51 -773 53
rect -807 19 -773 51
rect -807 -51 -773 -19
rect -807 -53 -773 -51
rect -807 -119 -773 -91
rect -807 -125 -773 -119
rect -807 -187 -773 -163
rect -807 -197 -773 -187
rect -807 -255 -773 -235
rect -807 -269 -773 -255
rect -807 -323 -773 -307
rect -807 -341 -773 -323
rect -807 -391 -773 -379
rect -807 -413 -773 -391
rect -807 -459 -773 -451
rect -807 -485 -773 -459
rect -649 459 -615 485
rect -649 451 -615 459
rect -649 391 -615 413
rect -649 379 -615 391
rect -649 323 -615 341
rect -649 307 -615 323
rect -649 255 -615 269
rect -649 235 -615 255
rect -649 187 -615 197
rect -649 163 -615 187
rect -649 119 -615 125
rect -649 91 -615 119
rect -649 51 -615 53
rect -649 19 -615 51
rect -649 -51 -615 -19
rect -649 -53 -615 -51
rect -649 -119 -615 -91
rect -649 -125 -615 -119
rect -649 -187 -615 -163
rect -649 -197 -615 -187
rect -649 -255 -615 -235
rect -649 -269 -615 -255
rect -649 -323 -615 -307
rect -649 -341 -615 -323
rect -649 -391 -615 -379
rect -649 -413 -615 -391
rect -649 -459 -615 -451
rect -649 -485 -615 -459
rect -491 459 -457 485
rect -491 451 -457 459
rect -491 391 -457 413
rect -491 379 -457 391
rect -491 323 -457 341
rect -491 307 -457 323
rect -491 255 -457 269
rect -491 235 -457 255
rect -491 187 -457 197
rect -491 163 -457 187
rect -491 119 -457 125
rect -491 91 -457 119
rect -491 51 -457 53
rect -491 19 -457 51
rect -491 -51 -457 -19
rect -491 -53 -457 -51
rect -491 -119 -457 -91
rect -491 -125 -457 -119
rect -491 -187 -457 -163
rect -491 -197 -457 -187
rect -491 -255 -457 -235
rect -491 -269 -457 -255
rect -491 -323 -457 -307
rect -491 -341 -457 -323
rect -491 -391 -457 -379
rect -491 -413 -457 -391
rect -491 -459 -457 -451
rect -491 -485 -457 -459
rect -333 459 -299 485
rect -333 451 -299 459
rect -333 391 -299 413
rect -333 379 -299 391
rect -333 323 -299 341
rect -333 307 -299 323
rect -333 255 -299 269
rect -333 235 -299 255
rect -333 187 -299 197
rect -333 163 -299 187
rect -333 119 -299 125
rect -333 91 -299 119
rect -333 51 -299 53
rect -333 19 -299 51
rect -333 -51 -299 -19
rect -333 -53 -299 -51
rect -333 -119 -299 -91
rect -333 -125 -299 -119
rect -333 -187 -299 -163
rect -333 -197 -299 -187
rect -333 -255 -299 -235
rect -333 -269 -299 -255
rect -333 -323 -299 -307
rect -333 -341 -299 -323
rect -333 -391 -299 -379
rect -333 -413 -299 -391
rect -333 -459 -299 -451
rect -333 -485 -299 -459
rect -175 459 -141 485
rect -175 451 -141 459
rect -175 391 -141 413
rect -175 379 -141 391
rect -175 323 -141 341
rect -175 307 -141 323
rect -175 255 -141 269
rect -175 235 -141 255
rect -175 187 -141 197
rect -175 163 -141 187
rect -175 119 -141 125
rect -175 91 -141 119
rect -175 51 -141 53
rect -175 19 -141 51
rect -175 -51 -141 -19
rect -175 -53 -141 -51
rect -175 -119 -141 -91
rect -175 -125 -141 -119
rect -175 -187 -141 -163
rect -175 -197 -141 -187
rect -175 -255 -141 -235
rect -175 -269 -141 -255
rect -175 -323 -141 -307
rect -175 -341 -141 -323
rect -175 -391 -141 -379
rect -175 -413 -141 -391
rect -175 -459 -141 -451
rect -175 -485 -141 -459
rect -17 459 17 485
rect -17 451 17 459
rect -17 391 17 413
rect -17 379 17 391
rect -17 323 17 341
rect -17 307 17 323
rect -17 255 17 269
rect -17 235 17 255
rect -17 187 17 197
rect -17 163 17 187
rect -17 119 17 125
rect -17 91 17 119
rect -17 51 17 53
rect -17 19 17 51
rect -17 -51 17 -19
rect -17 -53 17 -51
rect -17 -119 17 -91
rect -17 -125 17 -119
rect -17 -187 17 -163
rect -17 -197 17 -187
rect -17 -255 17 -235
rect -17 -269 17 -255
rect -17 -323 17 -307
rect -17 -341 17 -323
rect -17 -391 17 -379
rect -17 -413 17 -391
rect -17 -459 17 -451
rect -17 -485 17 -459
rect 141 459 175 485
rect 141 451 175 459
rect 141 391 175 413
rect 141 379 175 391
rect 141 323 175 341
rect 141 307 175 323
rect 141 255 175 269
rect 141 235 175 255
rect 141 187 175 197
rect 141 163 175 187
rect 141 119 175 125
rect 141 91 175 119
rect 141 51 175 53
rect 141 19 175 51
rect 141 -51 175 -19
rect 141 -53 175 -51
rect 141 -119 175 -91
rect 141 -125 175 -119
rect 141 -187 175 -163
rect 141 -197 175 -187
rect 141 -255 175 -235
rect 141 -269 175 -255
rect 141 -323 175 -307
rect 141 -341 175 -323
rect 141 -391 175 -379
rect 141 -413 175 -391
rect 141 -459 175 -451
rect 141 -485 175 -459
rect 299 459 333 485
rect 299 451 333 459
rect 299 391 333 413
rect 299 379 333 391
rect 299 323 333 341
rect 299 307 333 323
rect 299 255 333 269
rect 299 235 333 255
rect 299 187 333 197
rect 299 163 333 187
rect 299 119 333 125
rect 299 91 333 119
rect 299 51 333 53
rect 299 19 333 51
rect 299 -51 333 -19
rect 299 -53 333 -51
rect 299 -119 333 -91
rect 299 -125 333 -119
rect 299 -187 333 -163
rect 299 -197 333 -187
rect 299 -255 333 -235
rect 299 -269 333 -255
rect 299 -323 333 -307
rect 299 -341 333 -323
rect 299 -391 333 -379
rect 299 -413 333 -391
rect 299 -459 333 -451
rect 299 -485 333 -459
rect 457 459 491 485
rect 457 451 491 459
rect 457 391 491 413
rect 457 379 491 391
rect 457 323 491 341
rect 457 307 491 323
rect 457 255 491 269
rect 457 235 491 255
rect 457 187 491 197
rect 457 163 491 187
rect 457 119 491 125
rect 457 91 491 119
rect 457 51 491 53
rect 457 19 491 51
rect 457 -51 491 -19
rect 457 -53 491 -51
rect 457 -119 491 -91
rect 457 -125 491 -119
rect 457 -187 491 -163
rect 457 -197 491 -187
rect 457 -255 491 -235
rect 457 -269 491 -255
rect 457 -323 491 -307
rect 457 -341 491 -323
rect 457 -391 491 -379
rect 457 -413 491 -391
rect 457 -459 491 -451
rect 457 -485 491 -459
rect 615 459 649 485
rect 615 451 649 459
rect 615 391 649 413
rect 615 379 649 391
rect 615 323 649 341
rect 615 307 649 323
rect 615 255 649 269
rect 615 235 649 255
rect 615 187 649 197
rect 615 163 649 187
rect 615 119 649 125
rect 615 91 649 119
rect 615 51 649 53
rect 615 19 649 51
rect 615 -51 649 -19
rect 615 -53 649 -51
rect 615 -119 649 -91
rect 615 -125 649 -119
rect 615 -187 649 -163
rect 615 -197 649 -187
rect 615 -255 649 -235
rect 615 -269 649 -255
rect 615 -323 649 -307
rect 615 -341 649 -323
rect 615 -391 649 -379
rect 615 -413 649 -391
rect 615 -459 649 -451
rect 615 -485 649 -459
rect 773 459 807 485
rect 773 451 807 459
rect 773 391 807 413
rect 773 379 807 391
rect 773 323 807 341
rect 773 307 807 323
rect 773 255 807 269
rect 773 235 807 255
rect 773 187 807 197
rect 773 163 807 187
rect 773 119 807 125
rect 773 91 807 119
rect 773 51 807 53
rect 773 19 807 51
rect 773 -51 807 -19
rect 773 -53 807 -51
rect 773 -119 807 -91
rect 773 -125 807 -119
rect 773 -187 807 -163
rect 773 -197 807 -187
rect 773 -255 807 -235
rect 773 -269 807 -255
rect 773 -323 807 -307
rect 773 -341 807 -323
rect 773 -391 807 -379
rect 773 -413 807 -391
rect 773 -459 807 -451
rect 773 -485 807 -459
rect 931 459 965 485
rect 931 451 965 459
rect 931 391 965 413
rect 931 379 965 391
rect 931 323 965 341
rect 931 307 965 323
rect 931 255 965 269
rect 931 235 965 255
rect 931 187 965 197
rect 931 163 965 187
rect 931 119 965 125
rect 931 91 965 119
rect 931 51 965 53
rect 931 19 965 51
rect 931 -51 965 -19
rect 931 -53 965 -51
rect 931 -119 965 -91
rect 931 -125 965 -119
rect 931 -187 965 -163
rect 931 -197 965 -187
rect 931 -255 965 -235
rect 931 -269 965 -255
rect 931 -323 965 -307
rect 931 -341 965 -323
rect 931 -391 965 -379
rect 931 -413 965 -391
rect 931 -459 965 -451
rect 931 -485 965 -459
rect 1089 459 1123 485
rect 1089 451 1123 459
rect 1089 391 1123 413
rect 1089 379 1123 391
rect 1089 323 1123 341
rect 1089 307 1123 323
rect 1089 255 1123 269
rect 1089 235 1123 255
rect 1089 187 1123 197
rect 1089 163 1123 187
rect 1089 119 1123 125
rect 1089 91 1123 119
rect 1089 51 1123 53
rect 1089 19 1123 51
rect 1089 -51 1123 -19
rect 1089 -53 1123 -51
rect 1089 -119 1123 -91
rect 1089 -125 1123 -119
rect 1089 -187 1123 -163
rect 1089 -197 1123 -187
rect 1089 -255 1123 -235
rect 1089 -269 1123 -255
rect 1089 -323 1123 -307
rect 1089 -341 1123 -323
rect 1089 -391 1123 -379
rect 1089 -413 1123 -391
rect 1089 -459 1123 -451
rect 1089 -485 1123 -459
rect 1247 459 1281 485
rect 1247 451 1281 459
rect 1247 391 1281 413
rect 1247 379 1281 391
rect 1247 323 1281 341
rect 1247 307 1281 323
rect 1247 255 1281 269
rect 1247 235 1281 255
rect 1247 187 1281 197
rect 1247 163 1281 187
rect 1247 119 1281 125
rect 1247 91 1281 119
rect 1247 51 1281 53
rect 1247 19 1281 51
rect 1247 -51 1281 -19
rect 1247 -53 1281 -51
rect 1247 -119 1281 -91
rect 1247 -125 1281 -119
rect 1247 -187 1281 -163
rect 1247 -197 1281 -187
rect 1247 -255 1281 -235
rect 1247 -269 1281 -255
rect 1247 -323 1281 -307
rect 1247 -341 1281 -323
rect 1247 -391 1281 -379
rect 1247 -413 1281 -391
rect 1247 -459 1281 -451
rect 1247 -485 1281 -459
rect 1405 459 1439 485
rect 1405 451 1439 459
rect 1405 391 1439 413
rect 1405 379 1439 391
rect 1405 323 1439 341
rect 1405 307 1439 323
rect 1405 255 1439 269
rect 1405 235 1439 255
rect 1405 187 1439 197
rect 1405 163 1439 187
rect 1405 119 1439 125
rect 1405 91 1439 119
rect 1405 51 1439 53
rect 1405 19 1439 51
rect 1405 -51 1439 -19
rect 1405 -53 1439 -51
rect 1405 -119 1439 -91
rect 1405 -125 1439 -119
rect 1405 -187 1439 -163
rect 1405 -197 1439 -187
rect 1405 -255 1439 -235
rect 1405 -269 1439 -255
rect 1405 -323 1439 -307
rect 1405 -341 1439 -323
rect 1405 -391 1439 -379
rect 1405 -413 1439 -391
rect 1405 -459 1439 -451
rect 1405 -485 1439 -459
rect 1563 459 1597 485
rect 1563 451 1597 459
rect 1563 391 1597 413
rect 1563 379 1597 391
rect 1563 323 1597 341
rect 1563 307 1597 323
rect 1563 255 1597 269
rect 1563 235 1597 255
rect 1563 187 1597 197
rect 1563 163 1597 187
rect 1563 119 1597 125
rect 1563 91 1597 119
rect 1563 51 1597 53
rect 1563 19 1597 51
rect 1563 -51 1597 -19
rect 1563 -53 1597 -51
rect 1563 -119 1597 -91
rect 1563 -125 1597 -119
rect 1563 -187 1597 -163
rect 1563 -197 1597 -187
rect 1563 -255 1597 -235
rect 1563 -269 1597 -255
rect 1563 -323 1597 -307
rect 1563 -341 1597 -323
rect 1563 -391 1597 -379
rect 1563 -413 1597 -391
rect 1563 -459 1597 -451
rect 1563 -485 1597 -459
rect 1721 459 1755 485
rect 1721 451 1755 459
rect 1721 391 1755 413
rect 1721 379 1755 391
rect 1721 323 1755 341
rect 1721 307 1755 323
rect 1721 255 1755 269
rect 1721 235 1755 255
rect 1721 187 1755 197
rect 1721 163 1755 187
rect 1721 119 1755 125
rect 1721 91 1755 119
rect 1721 51 1755 53
rect 1721 19 1755 51
rect 1721 -51 1755 -19
rect 1721 -53 1755 -51
rect 1721 -119 1755 -91
rect 1721 -125 1755 -119
rect 1721 -187 1755 -163
rect 1721 -197 1755 -187
rect 1721 -255 1755 -235
rect 1721 -269 1755 -255
rect 1721 -323 1755 -307
rect 1721 -341 1755 -323
rect 1721 -391 1755 -379
rect 1721 -413 1755 -391
rect 1721 -459 1755 -451
rect 1721 -485 1755 -459
rect 1879 459 1913 485
rect 1879 451 1913 459
rect 1879 391 1913 413
rect 1879 379 1913 391
rect 1879 323 1913 341
rect 1879 307 1913 323
rect 1879 255 1913 269
rect 1879 235 1913 255
rect 1879 187 1913 197
rect 1879 163 1913 187
rect 1879 119 1913 125
rect 1879 91 1913 119
rect 1879 51 1913 53
rect 1879 19 1913 51
rect 1879 -51 1913 -19
rect 1879 -53 1913 -51
rect 1879 -119 1913 -91
rect 1879 -125 1913 -119
rect 1879 -187 1913 -163
rect 1879 -197 1913 -187
rect 1879 -255 1913 -235
rect 1879 -269 1913 -255
rect 1879 -323 1913 -307
rect 1879 -341 1913 -323
rect 1879 -391 1913 -379
rect 1879 -413 1913 -391
rect 1879 -459 1913 -451
rect 1879 -485 1913 -459
rect 2037 459 2071 485
rect 2037 451 2071 459
rect 2037 391 2071 413
rect 2037 379 2071 391
rect 2037 323 2071 341
rect 2037 307 2071 323
rect 2037 255 2071 269
rect 2037 235 2071 255
rect 2037 187 2071 197
rect 2037 163 2071 187
rect 2037 119 2071 125
rect 2037 91 2071 119
rect 2037 51 2071 53
rect 2037 19 2071 51
rect 2037 -51 2071 -19
rect 2037 -53 2071 -51
rect 2037 -119 2071 -91
rect 2037 -125 2071 -119
rect 2037 -187 2071 -163
rect 2037 -197 2071 -187
rect 2037 -255 2071 -235
rect 2037 -269 2071 -255
rect 2037 -323 2071 -307
rect 2037 -341 2071 -323
rect 2037 -391 2071 -379
rect 2037 -413 2071 -391
rect 2037 -459 2071 -451
rect 2037 -485 2071 -459
rect 2195 459 2229 485
rect 2195 451 2229 459
rect 2195 391 2229 413
rect 2195 379 2229 391
rect 2195 323 2229 341
rect 2195 307 2229 323
rect 2195 255 2229 269
rect 2195 235 2229 255
rect 2195 187 2229 197
rect 2195 163 2229 187
rect 2195 119 2229 125
rect 2195 91 2229 119
rect 2195 51 2229 53
rect 2195 19 2229 51
rect 2195 -51 2229 -19
rect 2195 -53 2229 -51
rect 2195 -119 2229 -91
rect 2195 -125 2229 -119
rect 2195 -187 2229 -163
rect 2195 -197 2229 -187
rect 2195 -255 2229 -235
rect 2195 -269 2229 -255
rect 2195 -323 2229 -307
rect 2195 -341 2229 -323
rect 2195 -391 2229 -379
rect 2195 -413 2229 -391
rect 2195 -459 2229 -451
rect 2195 -485 2229 -459
rect 2353 459 2387 485
rect 2353 451 2387 459
rect 2353 391 2387 413
rect 2353 379 2387 391
rect 2353 323 2387 341
rect 2353 307 2387 323
rect 2353 255 2387 269
rect 2353 235 2387 255
rect 2353 187 2387 197
rect 2353 163 2387 187
rect 2353 119 2387 125
rect 2353 91 2387 119
rect 2353 51 2387 53
rect 2353 19 2387 51
rect 2353 -51 2387 -19
rect 2353 -53 2387 -51
rect 2353 -119 2387 -91
rect 2353 -125 2387 -119
rect 2353 -187 2387 -163
rect 2353 -197 2387 -187
rect 2353 -255 2387 -235
rect 2353 -269 2387 -255
rect 2353 -323 2387 -307
rect 2353 -341 2387 -323
rect 2353 -391 2387 -379
rect 2353 -413 2387 -391
rect 2353 -459 2387 -451
rect 2353 -485 2387 -459
rect 2511 459 2545 485
rect 2511 451 2545 459
rect 2511 391 2545 413
rect 2511 379 2545 391
rect 2511 323 2545 341
rect 2511 307 2545 323
rect 2511 255 2545 269
rect 2511 235 2545 255
rect 2511 187 2545 197
rect 2511 163 2545 187
rect 2511 119 2545 125
rect 2511 91 2545 119
rect 2511 51 2545 53
rect 2511 19 2545 51
rect 2511 -51 2545 -19
rect 2511 -53 2545 -51
rect 2511 -119 2545 -91
rect 2511 -125 2545 -119
rect 2511 -187 2545 -163
rect 2511 -197 2545 -187
rect 2511 -255 2545 -235
rect 2511 -269 2545 -255
rect 2511 -323 2545 -307
rect 2511 -341 2545 -323
rect 2511 -391 2545 -379
rect 2511 -413 2545 -391
rect 2511 -459 2545 -451
rect 2511 -485 2545 -459
rect 2669 459 2703 485
rect 2669 451 2703 459
rect 2669 391 2703 413
rect 2669 379 2703 391
rect 2669 323 2703 341
rect 2669 307 2703 323
rect 2669 255 2703 269
rect 2669 235 2703 255
rect 2669 187 2703 197
rect 2669 163 2703 187
rect 2669 119 2703 125
rect 2669 91 2703 119
rect 2669 51 2703 53
rect 2669 19 2703 51
rect 2669 -51 2703 -19
rect 2669 -53 2703 -51
rect 2669 -119 2703 -91
rect 2669 -125 2703 -119
rect 2669 -187 2703 -163
rect 2669 -197 2703 -187
rect 2669 -255 2703 -235
rect 2669 -269 2703 -255
rect 2669 -323 2703 -307
rect 2669 -341 2703 -323
rect 2669 -391 2703 -379
rect 2669 -413 2703 -391
rect 2669 -459 2703 -451
rect 2669 -485 2703 -459
rect 2827 459 2861 485
rect 2827 451 2861 459
rect 2827 391 2861 413
rect 2827 379 2861 391
rect 2827 323 2861 341
rect 2827 307 2861 323
rect 2827 255 2861 269
rect 2827 235 2861 255
rect 2827 187 2861 197
rect 2827 163 2861 187
rect 2827 119 2861 125
rect 2827 91 2861 119
rect 2827 51 2861 53
rect 2827 19 2861 51
rect 2827 -51 2861 -19
rect 2827 -53 2861 -51
rect 2827 -119 2861 -91
rect 2827 -125 2861 -119
rect 2827 -187 2861 -163
rect 2827 -197 2861 -187
rect 2827 -255 2861 -235
rect 2827 -269 2861 -255
rect 2827 -323 2861 -307
rect 2827 -341 2861 -323
rect 2827 -391 2861 -379
rect 2827 -413 2861 -391
rect 2827 -459 2861 -451
rect 2827 -485 2861 -459
rect 2985 459 3019 485
rect 2985 451 3019 459
rect 2985 391 3019 413
rect 2985 379 3019 391
rect 2985 323 3019 341
rect 2985 307 3019 323
rect 2985 255 3019 269
rect 2985 235 3019 255
rect 2985 187 3019 197
rect 2985 163 3019 187
rect 2985 119 3019 125
rect 2985 91 3019 119
rect 2985 51 3019 53
rect 2985 19 3019 51
rect 2985 -51 3019 -19
rect 2985 -53 3019 -51
rect 2985 -119 3019 -91
rect 2985 -125 3019 -119
rect 2985 -187 3019 -163
rect 2985 -197 3019 -187
rect 2985 -255 3019 -235
rect 2985 -269 3019 -255
rect 2985 -323 3019 -307
rect 2985 -341 3019 -323
rect 2985 -391 3019 -379
rect 2985 -413 3019 -391
rect 2985 -459 3019 -451
rect 2985 -485 3019 -459
rect 3143 459 3177 485
rect 3143 451 3177 459
rect 3143 391 3177 413
rect 3143 379 3177 391
rect 3143 323 3177 341
rect 3143 307 3177 323
rect 3143 255 3177 269
rect 3143 235 3177 255
rect 3143 187 3177 197
rect 3143 163 3177 187
rect 3143 119 3177 125
rect 3143 91 3177 119
rect 3143 51 3177 53
rect 3143 19 3177 51
rect 3143 -51 3177 -19
rect 3143 -53 3177 -51
rect 3143 -119 3177 -91
rect 3143 -125 3177 -119
rect 3143 -187 3177 -163
rect 3143 -197 3177 -187
rect 3143 -255 3177 -235
rect 3143 -269 3177 -255
rect 3143 -323 3177 -307
rect 3143 -341 3177 -323
rect 3143 -391 3177 -379
rect 3143 -413 3177 -391
rect 3143 -459 3177 -451
rect 3143 -485 3177 -459
rect -3098 -581 -3064 -547
rect -2940 -581 -2906 -547
rect -2782 -581 -2748 -547
rect -2624 -581 -2590 -547
rect -2466 -581 -2432 -547
rect -2308 -581 -2274 -547
rect -2150 -581 -2116 -547
rect -1992 -581 -1958 -547
rect -1834 -581 -1800 -547
rect -1676 -581 -1642 -547
rect -1518 -581 -1484 -547
rect -1360 -581 -1326 -547
rect -1202 -581 -1168 -547
rect -1044 -581 -1010 -547
rect -886 -581 -852 -547
rect -728 -581 -694 -547
rect -570 -581 -536 -547
rect -412 -581 -378 -547
rect -254 -581 -220 -547
rect -96 -581 -62 -547
rect 62 -581 96 -547
rect 220 -581 254 -547
rect 378 -581 412 -547
rect 536 -581 570 -547
rect 694 -581 728 -547
rect 852 -581 886 -547
rect 1010 -581 1044 -547
rect 1168 -581 1202 -547
rect 1326 -581 1360 -547
rect 1484 -581 1518 -547
rect 1642 -581 1676 -547
rect 1800 -581 1834 -547
rect 1958 -581 1992 -547
rect 2116 -581 2150 -547
rect 2274 -581 2308 -547
rect 2432 -581 2466 -547
rect 2590 -581 2624 -547
rect 2748 -581 2782 -547
rect 2906 -581 2940 -547
rect 3064 -581 3098 -547
rect -1601 -683 -1581 -649
rect -1581 -683 -1567 -649
rect -1529 -683 -1513 -649
rect -1513 -683 -1495 -649
rect -1457 -683 -1445 -649
rect -1445 -683 -1423 -649
rect -1385 -683 -1377 -649
rect -1377 -683 -1351 -649
rect -1313 -683 -1309 -649
rect -1309 -683 -1279 -649
rect -1241 -683 -1207 -649
rect -1169 -683 -1139 -649
rect -1139 -683 -1135 -649
rect -1097 -683 -1071 -649
rect -1071 -683 -1063 -649
rect -1025 -683 -1003 -649
rect -1003 -683 -991 -649
rect -953 -683 -935 -649
rect -935 -683 -919 -649
rect -881 -683 -867 -649
rect -867 -683 -847 -649
rect -809 -683 -799 -649
rect -799 -683 -775 -649
rect -737 -683 -731 -649
rect -731 -683 -703 -649
rect -665 -683 -663 -649
rect -663 -683 -631 -649
rect -593 -683 -561 -649
rect -561 -683 -559 -649
rect -521 -683 -493 -649
rect -493 -683 -487 -649
rect -449 -683 -425 -649
rect -425 -683 -415 -649
rect -377 -683 -357 -649
rect -357 -683 -343 -649
rect -305 -683 -289 -649
rect -289 -683 -271 -649
rect -233 -683 -221 -649
rect -221 -683 -199 -649
rect -161 -683 -153 -649
rect -153 -683 -127 -649
rect -89 -683 -85 -649
rect -85 -683 -55 -649
rect -17 -683 17 -649
rect 55 -683 85 -649
rect 85 -683 89 -649
rect 127 -683 153 -649
rect 153 -683 161 -649
rect 199 -683 221 -649
rect 221 -683 233 -649
rect 271 -683 289 -649
rect 289 -683 305 -649
rect 343 -683 357 -649
rect 357 -683 377 -649
rect 415 -683 425 -649
rect 425 -683 449 -649
rect 487 -683 493 -649
rect 493 -683 521 -649
rect 559 -683 561 -649
rect 561 -683 593 -649
rect 631 -683 663 -649
rect 663 -683 665 -649
rect 703 -683 731 -649
rect 731 -683 737 -649
rect 775 -683 799 -649
rect 799 -683 809 -649
rect 847 -683 867 -649
rect 867 -683 881 -649
rect 919 -683 935 -649
rect 935 -683 953 -649
rect 991 -683 1003 -649
rect 1003 -683 1025 -649
rect 1063 -683 1071 -649
rect 1071 -683 1097 -649
rect 1135 -683 1139 -649
rect 1139 -683 1169 -649
rect 1207 -683 1241 -649
rect 1279 -683 1309 -649
rect 1309 -683 1313 -649
rect 1351 -683 1377 -649
rect 1377 -683 1385 -649
rect 1423 -683 1445 -649
rect 1445 -683 1457 -649
rect 1495 -683 1513 -649
rect 1513 -683 1529 -649
rect 1567 -683 1581 -649
rect 1581 -683 1601 -649
<< metal1 >>
rect -1640 683 1640 689
rect -1640 649 -1601 683
rect -1567 649 -1529 683
rect -1495 649 -1457 683
rect -1423 649 -1385 683
rect -1351 649 -1313 683
rect -1279 649 -1241 683
rect -1207 649 -1169 683
rect -1135 649 -1097 683
rect -1063 649 -1025 683
rect -991 649 -953 683
rect -919 649 -881 683
rect -847 649 -809 683
rect -775 649 -737 683
rect -703 649 -665 683
rect -631 649 -593 683
rect -559 649 -521 683
rect -487 649 -449 683
rect -415 649 -377 683
rect -343 649 -305 683
rect -271 649 -233 683
rect -199 649 -161 683
rect -127 649 -89 683
rect -55 649 -17 683
rect 17 649 55 683
rect 89 649 127 683
rect 161 649 199 683
rect 233 649 271 683
rect 305 649 343 683
rect 377 649 415 683
rect 449 649 487 683
rect 521 649 559 683
rect 593 649 631 683
rect 665 649 703 683
rect 737 649 775 683
rect 809 649 847 683
rect 881 649 919 683
rect 953 649 991 683
rect 1025 649 1063 683
rect 1097 649 1135 683
rect 1169 649 1207 683
rect 1241 649 1279 683
rect 1313 649 1351 683
rect 1385 649 1423 683
rect 1457 649 1495 683
rect 1529 649 1567 683
rect 1601 649 1640 683
rect -1640 643 1640 649
rect -3127 581 -3035 587
rect -3127 547 -3098 581
rect -3064 547 -3035 581
rect -3127 541 -3035 547
rect -2969 581 -2877 587
rect -2969 547 -2940 581
rect -2906 547 -2877 581
rect -2969 541 -2877 547
rect -2811 581 -2719 587
rect -2811 547 -2782 581
rect -2748 547 -2719 581
rect -2811 541 -2719 547
rect -2653 581 -2561 587
rect -2653 547 -2624 581
rect -2590 547 -2561 581
rect -2653 541 -2561 547
rect -2495 581 -2403 587
rect -2495 547 -2466 581
rect -2432 547 -2403 581
rect -2495 541 -2403 547
rect -2337 581 -2245 587
rect -2337 547 -2308 581
rect -2274 547 -2245 581
rect -2337 541 -2245 547
rect -2179 581 -2087 587
rect -2179 547 -2150 581
rect -2116 547 -2087 581
rect -2179 541 -2087 547
rect -2021 581 -1929 587
rect -2021 547 -1992 581
rect -1958 547 -1929 581
rect -2021 541 -1929 547
rect -1863 581 -1771 587
rect -1863 547 -1834 581
rect -1800 547 -1771 581
rect -1863 541 -1771 547
rect -1705 581 -1613 587
rect -1705 547 -1676 581
rect -1642 547 -1613 581
rect -1705 541 -1613 547
rect -1547 581 -1455 587
rect -1547 547 -1518 581
rect -1484 547 -1455 581
rect -1547 541 -1455 547
rect -1389 581 -1297 587
rect -1389 547 -1360 581
rect -1326 547 -1297 581
rect -1389 541 -1297 547
rect -1231 581 -1139 587
rect -1231 547 -1202 581
rect -1168 547 -1139 581
rect -1231 541 -1139 547
rect -1073 581 -981 587
rect -1073 547 -1044 581
rect -1010 547 -981 581
rect -1073 541 -981 547
rect -915 581 -823 587
rect -915 547 -886 581
rect -852 547 -823 581
rect -915 541 -823 547
rect -757 581 -665 587
rect -757 547 -728 581
rect -694 547 -665 581
rect -757 541 -665 547
rect -599 581 -507 587
rect -599 547 -570 581
rect -536 547 -507 581
rect -599 541 -507 547
rect -441 581 -349 587
rect -441 547 -412 581
rect -378 547 -349 581
rect -441 541 -349 547
rect -283 581 -191 587
rect -283 547 -254 581
rect -220 547 -191 581
rect -283 541 -191 547
rect -125 581 -33 587
rect -125 547 -96 581
rect -62 547 -33 581
rect -125 541 -33 547
rect 33 581 125 587
rect 33 547 62 581
rect 96 547 125 581
rect 33 541 125 547
rect 191 581 283 587
rect 191 547 220 581
rect 254 547 283 581
rect 191 541 283 547
rect 349 581 441 587
rect 349 547 378 581
rect 412 547 441 581
rect 349 541 441 547
rect 507 581 599 587
rect 507 547 536 581
rect 570 547 599 581
rect 507 541 599 547
rect 665 581 757 587
rect 665 547 694 581
rect 728 547 757 581
rect 665 541 757 547
rect 823 581 915 587
rect 823 547 852 581
rect 886 547 915 581
rect 823 541 915 547
rect 981 581 1073 587
rect 981 547 1010 581
rect 1044 547 1073 581
rect 981 541 1073 547
rect 1139 581 1231 587
rect 1139 547 1168 581
rect 1202 547 1231 581
rect 1139 541 1231 547
rect 1297 581 1389 587
rect 1297 547 1326 581
rect 1360 547 1389 581
rect 1297 541 1389 547
rect 1455 581 1547 587
rect 1455 547 1484 581
rect 1518 547 1547 581
rect 1455 541 1547 547
rect 1613 581 1705 587
rect 1613 547 1642 581
rect 1676 547 1705 581
rect 1613 541 1705 547
rect 1771 581 1863 587
rect 1771 547 1800 581
rect 1834 547 1863 581
rect 1771 541 1863 547
rect 1929 581 2021 587
rect 1929 547 1958 581
rect 1992 547 2021 581
rect 1929 541 2021 547
rect 2087 581 2179 587
rect 2087 547 2116 581
rect 2150 547 2179 581
rect 2087 541 2179 547
rect 2245 581 2337 587
rect 2245 547 2274 581
rect 2308 547 2337 581
rect 2245 541 2337 547
rect 2403 581 2495 587
rect 2403 547 2432 581
rect 2466 547 2495 581
rect 2403 541 2495 547
rect 2561 581 2653 587
rect 2561 547 2590 581
rect 2624 547 2653 581
rect 2561 541 2653 547
rect 2719 581 2811 587
rect 2719 547 2748 581
rect 2782 547 2811 581
rect 2719 541 2811 547
rect 2877 581 2969 587
rect 2877 547 2906 581
rect 2940 547 2969 581
rect 2877 541 2969 547
rect 3035 581 3127 587
rect 3035 547 3064 581
rect 3098 547 3127 581
rect 3035 541 3127 547
rect -3183 485 -3137 500
rect -3183 451 -3177 485
rect -3143 451 -3137 485
rect -3183 413 -3137 451
rect -3183 379 -3177 413
rect -3143 379 -3137 413
rect -3183 341 -3137 379
rect -3183 307 -3177 341
rect -3143 307 -3137 341
rect -3183 269 -3137 307
rect -3183 235 -3177 269
rect -3143 235 -3137 269
rect -3183 197 -3137 235
rect -3183 163 -3177 197
rect -3143 163 -3137 197
rect -3183 125 -3137 163
rect -3183 91 -3177 125
rect -3143 91 -3137 125
rect -3183 53 -3137 91
rect -3183 19 -3177 53
rect -3143 19 -3137 53
rect -3183 -19 -3137 19
rect -3183 -53 -3177 -19
rect -3143 -53 -3137 -19
rect -3183 -91 -3137 -53
rect -3183 -125 -3177 -91
rect -3143 -125 -3137 -91
rect -3183 -163 -3137 -125
rect -3183 -197 -3177 -163
rect -3143 -197 -3137 -163
rect -3183 -235 -3137 -197
rect -3183 -269 -3177 -235
rect -3143 -269 -3137 -235
rect -3183 -307 -3137 -269
rect -3183 -341 -3177 -307
rect -3143 -341 -3137 -307
rect -3183 -379 -3137 -341
rect -3183 -413 -3177 -379
rect -3143 -413 -3137 -379
rect -3183 -451 -3137 -413
rect -3183 -485 -3177 -451
rect -3143 -485 -3137 -451
rect -3183 -500 -3137 -485
rect -3025 485 -2979 500
rect -3025 451 -3019 485
rect -2985 451 -2979 485
rect -3025 413 -2979 451
rect -3025 379 -3019 413
rect -2985 379 -2979 413
rect -3025 341 -2979 379
rect -3025 307 -3019 341
rect -2985 307 -2979 341
rect -3025 269 -2979 307
rect -3025 235 -3019 269
rect -2985 235 -2979 269
rect -3025 197 -2979 235
rect -3025 163 -3019 197
rect -2985 163 -2979 197
rect -3025 125 -2979 163
rect -3025 91 -3019 125
rect -2985 91 -2979 125
rect -3025 53 -2979 91
rect -3025 19 -3019 53
rect -2985 19 -2979 53
rect -3025 -19 -2979 19
rect -3025 -53 -3019 -19
rect -2985 -53 -2979 -19
rect -3025 -91 -2979 -53
rect -3025 -125 -3019 -91
rect -2985 -125 -2979 -91
rect -3025 -163 -2979 -125
rect -3025 -197 -3019 -163
rect -2985 -197 -2979 -163
rect -3025 -235 -2979 -197
rect -3025 -269 -3019 -235
rect -2985 -269 -2979 -235
rect -3025 -307 -2979 -269
rect -3025 -341 -3019 -307
rect -2985 -341 -2979 -307
rect -3025 -379 -2979 -341
rect -3025 -413 -3019 -379
rect -2985 -413 -2979 -379
rect -3025 -451 -2979 -413
rect -3025 -485 -3019 -451
rect -2985 -485 -2979 -451
rect -3025 -500 -2979 -485
rect -2867 485 -2821 500
rect -2867 451 -2861 485
rect -2827 451 -2821 485
rect -2867 413 -2821 451
rect -2867 379 -2861 413
rect -2827 379 -2821 413
rect -2867 341 -2821 379
rect -2867 307 -2861 341
rect -2827 307 -2821 341
rect -2867 269 -2821 307
rect -2867 235 -2861 269
rect -2827 235 -2821 269
rect -2867 197 -2821 235
rect -2867 163 -2861 197
rect -2827 163 -2821 197
rect -2867 125 -2821 163
rect -2867 91 -2861 125
rect -2827 91 -2821 125
rect -2867 53 -2821 91
rect -2867 19 -2861 53
rect -2827 19 -2821 53
rect -2867 -19 -2821 19
rect -2867 -53 -2861 -19
rect -2827 -53 -2821 -19
rect -2867 -91 -2821 -53
rect -2867 -125 -2861 -91
rect -2827 -125 -2821 -91
rect -2867 -163 -2821 -125
rect -2867 -197 -2861 -163
rect -2827 -197 -2821 -163
rect -2867 -235 -2821 -197
rect -2867 -269 -2861 -235
rect -2827 -269 -2821 -235
rect -2867 -307 -2821 -269
rect -2867 -341 -2861 -307
rect -2827 -341 -2821 -307
rect -2867 -379 -2821 -341
rect -2867 -413 -2861 -379
rect -2827 -413 -2821 -379
rect -2867 -451 -2821 -413
rect -2867 -485 -2861 -451
rect -2827 -485 -2821 -451
rect -2867 -500 -2821 -485
rect -2709 485 -2663 500
rect -2709 451 -2703 485
rect -2669 451 -2663 485
rect -2709 413 -2663 451
rect -2709 379 -2703 413
rect -2669 379 -2663 413
rect -2709 341 -2663 379
rect -2709 307 -2703 341
rect -2669 307 -2663 341
rect -2709 269 -2663 307
rect -2709 235 -2703 269
rect -2669 235 -2663 269
rect -2709 197 -2663 235
rect -2709 163 -2703 197
rect -2669 163 -2663 197
rect -2709 125 -2663 163
rect -2709 91 -2703 125
rect -2669 91 -2663 125
rect -2709 53 -2663 91
rect -2709 19 -2703 53
rect -2669 19 -2663 53
rect -2709 -19 -2663 19
rect -2709 -53 -2703 -19
rect -2669 -53 -2663 -19
rect -2709 -91 -2663 -53
rect -2709 -125 -2703 -91
rect -2669 -125 -2663 -91
rect -2709 -163 -2663 -125
rect -2709 -197 -2703 -163
rect -2669 -197 -2663 -163
rect -2709 -235 -2663 -197
rect -2709 -269 -2703 -235
rect -2669 -269 -2663 -235
rect -2709 -307 -2663 -269
rect -2709 -341 -2703 -307
rect -2669 -341 -2663 -307
rect -2709 -379 -2663 -341
rect -2709 -413 -2703 -379
rect -2669 -413 -2663 -379
rect -2709 -451 -2663 -413
rect -2709 -485 -2703 -451
rect -2669 -485 -2663 -451
rect -2709 -500 -2663 -485
rect -2551 485 -2505 500
rect -2551 451 -2545 485
rect -2511 451 -2505 485
rect -2551 413 -2505 451
rect -2551 379 -2545 413
rect -2511 379 -2505 413
rect -2551 341 -2505 379
rect -2551 307 -2545 341
rect -2511 307 -2505 341
rect -2551 269 -2505 307
rect -2551 235 -2545 269
rect -2511 235 -2505 269
rect -2551 197 -2505 235
rect -2551 163 -2545 197
rect -2511 163 -2505 197
rect -2551 125 -2505 163
rect -2551 91 -2545 125
rect -2511 91 -2505 125
rect -2551 53 -2505 91
rect -2551 19 -2545 53
rect -2511 19 -2505 53
rect -2551 -19 -2505 19
rect -2551 -53 -2545 -19
rect -2511 -53 -2505 -19
rect -2551 -91 -2505 -53
rect -2551 -125 -2545 -91
rect -2511 -125 -2505 -91
rect -2551 -163 -2505 -125
rect -2551 -197 -2545 -163
rect -2511 -197 -2505 -163
rect -2551 -235 -2505 -197
rect -2551 -269 -2545 -235
rect -2511 -269 -2505 -235
rect -2551 -307 -2505 -269
rect -2551 -341 -2545 -307
rect -2511 -341 -2505 -307
rect -2551 -379 -2505 -341
rect -2551 -413 -2545 -379
rect -2511 -413 -2505 -379
rect -2551 -451 -2505 -413
rect -2551 -485 -2545 -451
rect -2511 -485 -2505 -451
rect -2551 -500 -2505 -485
rect -2393 485 -2347 500
rect -2393 451 -2387 485
rect -2353 451 -2347 485
rect -2393 413 -2347 451
rect -2393 379 -2387 413
rect -2353 379 -2347 413
rect -2393 341 -2347 379
rect -2393 307 -2387 341
rect -2353 307 -2347 341
rect -2393 269 -2347 307
rect -2393 235 -2387 269
rect -2353 235 -2347 269
rect -2393 197 -2347 235
rect -2393 163 -2387 197
rect -2353 163 -2347 197
rect -2393 125 -2347 163
rect -2393 91 -2387 125
rect -2353 91 -2347 125
rect -2393 53 -2347 91
rect -2393 19 -2387 53
rect -2353 19 -2347 53
rect -2393 -19 -2347 19
rect -2393 -53 -2387 -19
rect -2353 -53 -2347 -19
rect -2393 -91 -2347 -53
rect -2393 -125 -2387 -91
rect -2353 -125 -2347 -91
rect -2393 -163 -2347 -125
rect -2393 -197 -2387 -163
rect -2353 -197 -2347 -163
rect -2393 -235 -2347 -197
rect -2393 -269 -2387 -235
rect -2353 -269 -2347 -235
rect -2393 -307 -2347 -269
rect -2393 -341 -2387 -307
rect -2353 -341 -2347 -307
rect -2393 -379 -2347 -341
rect -2393 -413 -2387 -379
rect -2353 -413 -2347 -379
rect -2393 -451 -2347 -413
rect -2393 -485 -2387 -451
rect -2353 -485 -2347 -451
rect -2393 -500 -2347 -485
rect -2235 485 -2189 500
rect -2235 451 -2229 485
rect -2195 451 -2189 485
rect -2235 413 -2189 451
rect -2235 379 -2229 413
rect -2195 379 -2189 413
rect -2235 341 -2189 379
rect -2235 307 -2229 341
rect -2195 307 -2189 341
rect -2235 269 -2189 307
rect -2235 235 -2229 269
rect -2195 235 -2189 269
rect -2235 197 -2189 235
rect -2235 163 -2229 197
rect -2195 163 -2189 197
rect -2235 125 -2189 163
rect -2235 91 -2229 125
rect -2195 91 -2189 125
rect -2235 53 -2189 91
rect -2235 19 -2229 53
rect -2195 19 -2189 53
rect -2235 -19 -2189 19
rect -2235 -53 -2229 -19
rect -2195 -53 -2189 -19
rect -2235 -91 -2189 -53
rect -2235 -125 -2229 -91
rect -2195 -125 -2189 -91
rect -2235 -163 -2189 -125
rect -2235 -197 -2229 -163
rect -2195 -197 -2189 -163
rect -2235 -235 -2189 -197
rect -2235 -269 -2229 -235
rect -2195 -269 -2189 -235
rect -2235 -307 -2189 -269
rect -2235 -341 -2229 -307
rect -2195 -341 -2189 -307
rect -2235 -379 -2189 -341
rect -2235 -413 -2229 -379
rect -2195 -413 -2189 -379
rect -2235 -451 -2189 -413
rect -2235 -485 -2229 -451
rect -2195 -485 -2189 -451
rect -2235 -500 -2189 -485
rect -2077 485 -2031 500
rect -2077 451 -2071 485
rect -2037 451 -2031 485
rect -2077 413 -2031 451
rect -2077 379 -2071 413
rect -2037 379 -2031 413
rect -2077 341 -2031 379
rect -2077 307 -2071 341
rect -2037 307 -2031 341
rect -2077 269 -2031 307
rect -2077 235 -2071 269
rect -2037 235 -2031 269
rect -2077 197 -2031 235
rect -2077 163 -2071 197
rect -2037 163 -2031 197
rect -2077 125 -2031 163
rect -2077 91 -2071 125
rect -2037 91 -2031 125
rect -2077 53 -2031 91
rect -2077 19 -2071 53
rect -2037 19 -2031 53
rect -2077 -19 -2031 19
rect -2077 -53 -2071 -19
rect -2037 -53 -2031 -19
rect -2077 -91 -2031 -53
rect -2077 -125 -2071 -91
rect -2037 -125 -2031 -91
rect -2077 -163 -2031 -125
rect -2077 -197 -2071 -163
rect -2037 -197 -2031 -163
rect -2077 -235 -2031 -197
rect -2077 -269 -2071 -235
rect -2037 -269 -2031 -235
rect -2077 -307 -2031 -269
rect -2077 -341 -2071 -307
rect -2037 -341 -2031 -307
rect -2077 -379 -2031 -341
rect -2077 -413 -2071 -379
rect -2037 -413 -2031 -379
rect -2077 -451 -2031 -413
rect -2077 -485 -2071 -451
rect -2037 -485 -2031 -451
rect -2077 -500 -2031 -485
rect -1919 485 -1873 500
rect -1919 451 -1913 485
rect -1879 451 -1873 485
rect -1919 413 -1873 451
rect -1919 379 -1913 413
rect -1879 379 -1873 413
rect -1919 341 -1873 379
rect -1919 307 -1913 341
rect -1879 307 -1873 341
rect -1919 269 -1873 307
rect -1919 235 -1913 269
rect -1879 235 -1873 269
rect -1919 197 -1873 235
rect -1919 163 -1913 197
rect -1879 163 -1873 197
rect -1919 125 -1873 163
rect -1919 91 -1913 125
rect -1879 91 -1873 125
rect -1919 53 -1873 91
rect -1919 19 -1913 53
rect -1879 19 -1873 53
rect -1919 -19 -1873 19
rect -1919 -53 -1913 -19
rect -1879 -53 -1873 -19
rect -1919 -91 -1873 -53
rect -1919 -125 -1913 -91
rect -1879 -125 -1873 -91
rect -1919 -163 -1873 -125
rect -1919 -197 -1913 -163
rect -1879 -197 -1873 -163
rect -1919 -235 -1873 -197
rect -1919 -269 -1913 -235
rect -1879 -269 -1873 -235
rect -1919 -307 -1873 -269
rect -1919 -341 -1913 -307
rect -1879 -341 -1873 -307
rect -1919 -379 -1873 -341
rect -1919 -413 -1913 -379
rect -1879 -413 -1873 -379
rect -1919 -451 -1873 -413
rect -1919 -485 -1913 -451
rect -1879 -485 -1873 -451
rect -1919 -500 -1873 -485
rect -1761 485 -1715 500
rect -1761 451 -1755 485
rect -1721 451 -1715 485
rect -1761 413 -1715 451
rect -1761 379 -1755 413
rect -1721 379 -1715 413
rect -1761 341 -1715 379
rect -1761 307 -1755 341
rect -1721 307 -1715 341
rect -1761 269 -1715 307
rect -1761 235 -1755 269
rect -1721 235 -1715 269
rect -1761 197 -1715 235
rect -1761 163 -1755 197
rect -1721 163 -1715 197
rect -1761 125 -1715 163
rect -1761 91 -1755 125
rect -1721 91 -1715 125
rect -1761 53 -1715 91
rect -1761 19 -1755 53
rect -1721 19 -1715 53
rect -1761 -19 -1715 19
rect -1761 -53 -1755 -19
rect -1721 -53 -1715 -19
rect -1761 -91 -1715 -53
rect -1761 -125 -1755 -91
rect -1721 -125 -1715 -91
rect -1761 -163 -1715 -125
rect -1761 -197 -1755 -163
rect -1721 -197 -1715 -163
rect -1761 -235 -1715 -197
rect -1761 -269 -1755 -235
rect -1721 -269 -1715 -235
rect -1761 -307 -1715 -269
rect -1761 -341 -1755 -307
rect -1721 -341 -1715 -307
rect -1761 -379 -1715 -341
rect -1761 -413 -1755 -379
rect -1721 -413 -1715 -379
rect -1761 -451 -1715 -413
rect -1761 -485 -1755 -451
rect -1721 -485 -1715 -451
rect -1761 -500 -1715 -485
rect -1603 485 -1557 500
rect -1603 451 -1597 485
rect -1563 451 -1557 485
rect -1603 413 -1557 451
rect -1603 379 -1597 413
rect -1563 379 -1557 413
rect -1603 341 -1557 379
rect -1603 307 -1597 341
rect -1563 307 -1557 341
rect -1603 269 -1557 307
rect -1603 235 -1597 269
rect -1563 235 -1557 269
rect -1603 197 -1557 235
rect -1603 163 -1597 197
rect -1563 163 -1557 197
rect -1603 125 -1557 163
rect -1603 91 -1597 125
rect -1563 91 -1557 125
rect -1603 53 -1557 91
rect -1603 19 -1597 53
rect -1563 19 -1557 53
rect -1603 -19 -1557 19
rect -1603 -53 -1597 -19
rect -1563 -53 -1557 -19
rect -1603 -91 -1557 -53
rect -1603 -125 -1597 -91
rect -1563 -125 -1557 -91
rect -1603 -163 -1557 -125
rect -1603 -197 -1597 -163
rect -1563 -197 -1557 -163
rect -1603 -235 -1557 -197
rect -1603 -269 -1597 -235
rect -1563 -269 -1557 -235
rect -1603 -307 -1557 -269
rect -1603 -341 -1597 -307
rect -1563 -341 -1557 -307
rect -1603 -379 -1557 -341
rect -1603 -413 -1597 -379
rect -1563 -413 -1557 -379
rect -1603 -451 -1557 -413
rect -1603 -485 -1597 -451
rect -1563 -485 -1557 -451
rect -1603 -500 -1557 -485
rect -1445 485 -1399 500
rect -1445 451 -1439 485
rect -1405 451 -1399 485
rect -1445 413 -1399 451
rect -1445 379 -1439 413
rect -1405 379 -1399 413
rect -1445 341 -1399 379
rect -1445 307 -1439 341
rect -1405 307 -1399 341
rect -1445 269 -1399 307
rect -1445 235 -1439 269
rect -1405 235 -1399 269
rect -1445 197 -1399 235
rect -1445 163 -1439 197
rect -1405 163 -1399 197
rect -1445 125 -1399 163
rect -1445 91 -1439 125
rect -1405 91 -1399 125
rect -1445 53 -1399 91
rect -1445 19 -1439 53
rect -1405 19 -1399 53
rect -1445 -19 -1399 19
rect -1445 -53 -1439 -19
rect -1405 -53 -1399 -19
rect -1445 -91 -1399 -53
rect -1445 -125 -1439 -91
rect -1405 -125 -1399 -91
rect -1445 -163 -1399 -125
rect -1445 -197 -1439 -163
rect -1405 -197 -1399 -163
rect -1445 -235 -1399 -197
rect -1445 -269 -1439 -235
rect -1405 -269 -1399 -235
rect -1445 -307 -1399 -269
rect -1445 -341 -1439 -307
rect -1405 -341 -1399 -307
rect -1445 -379 -1399 -341
rect -1445 -413 -1439 -379
rect -1405 -413 -1399 -379
rect -1445 -451 -1399 -413
rect -1445 -485 -1439 -451
rect -1405 -485 -1399 -451
rect -1445 -500 -1399 -485
rect -1287 485 -1241 500
rect -1287 451 -1281 485
rect -1247 451 -1241 485
rect -1287 413 -1241 451
rect -1287 379 -1281 413
rect -1247 379 -1241 413
rect -1287 341 -1241 379
rect -1287 307 -1281 341
rect -1247 307 -1241 341
rect -1287 269 -1241 307
rect -1287 235 -1281 269
rect -1247 235 -1241 269
rect -1287 197 -1241 235
rect -1287 163 -1281 197
rect -1247 163 -1241 197
rect -1287 125 -1241 163
rect -1287 91 -1281 125
rect -1247 91 -1241 125
rect -1287 53 -1241 91
rect -1287 19 -1281 53
rect -1247 19 -1241 53
rect -1287 -19 -1241 19
rect -1287 -53 -1281 -19
rect -1247 -53 -1241 -19
rect -1287 -91 -1241 -53
rect -1287 -125 -1281 -91
rect -1247 -125 -1241 -91
rect -1287 -163 -1241 -125
rect -1287 -197 -1281 -163
rect -1247 -197 -1241 -163
rect -1287 -235 -1241 -197
rect -1287 -269 -1281 -235
rect -1247 -269 -1241 -235
rect -1287 -307 -1241 -269
rect -1287 -341 -1281 -307
rect -1247 -341 -1241 -307
rect -1287 -379 -1241 -341
rect -1287 -413 -1281 -379
rect -1247 -413 -1241 -379
rect -1287 -451 -1241 -413
rect -1287 -485 -1281 -451
rect -1247 -485 -1241 -451
rect -1287 -500 -1241 -485
rect -1129 485 -1083 500
rect -1129 451 -1123 485
rect -1089 451 -1083 485
rect -1129 413 -1083 451
rect -1129 379 -1123 413
rect -1089 379 -1083 413
rect -1129 341 -1083 379
rect -1129 307 -1123 341
rect -1089 307 -1083 341
rect -1129 269 -1083 307
rect -1129 235 -1123 269
rect -1089 235 -1083 269
rect -1129 197 -1083 235
rect -1129 163 -1123 197
rect -1089 163 -1083 197
rect -1129 125 -1083 163
rect -1129 91 -1123 125
rect -1089 91 -1083 125
rect -1129 53 -1083 91
rect -1129 19 -1123 53
rect -1089 19 -1083 53
rect -1129 -19 -1083 19
rect -1129 -53 -1123 -19
rect -1089 -53 -1083 -19
rect -1129 -91 -1083 -53
rect -1129 -125 -1123 -91
rect -1089 -125 -1083 -91
rect -1129 -163 -1083 -125
rect -1129 -197 -1123 -163
rect -1089 -197 -1083 -163
rect -1129 -235 -1083 -197
rect -1129 -269 -1123 -235
rect -1089 -269 -1083 -235
rect -1129 -307 -1083 -269
rect -1129 -341 -1123 -307
rect -1089 -341 -1083 -307
rect -1129 -379 -1083 -341
rect -1129 -413 -1123 -379
rect -1089 -413 -1083 -379
rect -1129 -451 -1083 -413
rect -1129 -485 -1123 -451
rect -1089 -485 -1083 -451
rect -1129 -500 -1083 -485
rect -971 485 -925 500
rect -971 451 -965 485
rect -931 451 -925 485
rect -971 413 -925 451
rect -971 379 -965 413
rect -931 379 -925 413
rect -971 341 -925 379
rect -971 307 -965 341
rect -931 307 -925 341
rect -971 269 -925 307
rect -971 235 -965 269
rect -931 235 -925 269
rect -971 197 -925 235
rect -971 163 -965 197
rect -931 163 -925 197
rect -971 125 -925 163
rect -971 91 -965 125
rect -931 91 -925 125
rect -971 53 -925 91
rect -971 19 -965 53
rect -931 19 -925 53
rect -971 -19 -925 19
rect -971 -53 -965 -19
rect -931 -53 -925 -19
rect -971 -91 -925 -53
rect -971 -125 -965 -91
rect -931 -125 -925 -91
rect -971 -163 -925 -125
rect -971 -197 -965 -163
rect -931 -197 -925 -163
rect -971 -235 -925 -197
rect -971 -269 -965 -235
rect -931 -269 -925 -235
rect -971 -307 -925 -269
rect -971 -341 -965 -307
rect -931 -341 -925 -307
rect -971 -379 -925 -341
rect -971 -413 -965 -379
rect -931 -413 -925 -379
rect -971 -451 -925 -413
rect -971 -485 -965 -451
rect -931 -485 -925 -451
rect -971 -500 -925 -485
rect -813 485 -767 500
rect -813 451 -807 485
rect -773 451 -767 485
rect -813 413 -767 451
rect -813 379 -807 413
rect -773 379 -767 413
rect -813 341 -767 379
rect -813 307 -807 341
rect -773 307 -767 341
rect -813 269 -767 307
rect -813 235 -807 269
rect -773 235 -767 269
rect -813 197 -767 235
rect -813 163 -807 197
rect -773 163 -767 197
rect -813 125 -767 163
rect -813 91 -807 125
rect -773 91 -767 125
rect -813 53 -767 91
rect -813 19 -807 53
rect -773 19 -767 53
rect -813 -19 -767 19
rect -813 -53 -807 -19
rect -773 -53 -767 -19
rect -813 -91 -767 -53
rect -813 -125 -807 -91
rect -773 -125 -767 -91
rect -813 -163 -767 -125
rect -813 -197 -807 -163
rect -773 -197 -767 -163
rect -813 -235 -767 -197
rect -813 -269 -807 -235
rect -773 -269 -767 -235
rect -813 -307 -767 -269
rect -813 -341 -807 -307
rect -773 -341 -767 -307
rect -813 -379 -767 -341
rect -813 -413 -807 -379
rect -773 -413 -767 -379
rect -813 -451 -767 -413
rect -813 -485 -807 -451
rect -773 -485 -767 -451
rect -813 -500 -767 -485
rect -655 485 -609 500
rect -655 451 -649 485
rect -615 451 -609 485
rect -655 413 -609 451
rect -655 379 -649 413
rect -615 379 -609 413
rect -655 341 -609 379
rect -655 307 -649 341
rect -615 307 -609 341
rect -655 269 -609 307
rect -655 235 -649 269
rect -615 235 -609 269
rect -655 197 -609 235
rect -655 163 -649 197
rect -615 163 -609 197
rect -655 125 -609 163
rect -655 91 -649 125
rect -615 91 -609 125
rect -655 53 -609 91
rect -655 19 -649 53
rect -615 19 -609 53
rect -655 -19 -609 19
rect -655 -53 -649 -19
rect -615 -53 -609 -19
rect -655 -91 -609 -53
rect -655 -125 -649 -91
rect -615 -125 -609 -91
rect -655 -163 -609 -125
rect -655 -197 -649 -163
rect -615 -197 -609 -163
rect -655 -235 -609 -197
rect -655 -269 -649 -235
rect -615 -269 -609 -235
rect -655 -307 -609 -269
rect -655 -341 -649 -307
rect -615 -341 -609 -307
rect -655 -379 -609 -341
rect -655 -413 -649 -379
rect -615 -413 -609 -379
rect -655 -451 -609 -413
rect -655 -485 -649 -451
rect -615 -485 -609 -451
rect -655 -500 -609 -485
rect -497 485 -451 500
rect -497 451 -491 485
rect -457 451 -451 485
rect -497 413 -451 451
rect -497 379 -491 413
rect -457 379 -451 413
rect -497 341 -451 379
rect -497 307 -491 341
rect -457 307 -451 341
rect -497 269 -451 307
rect -497 235 -491 269
rect -457 235 -451 269
rect -497 197 -451 235
rect -497 163 -491 197
rect -457 163 -451 197
rect -497 125 -451 163
rect -497 91 -491 125
rect -457 91 -451 125
rect -497 53 -451 91
rect -497 19 -491 53
rect -457 19 -451 53
rect -497 -19 -451 19
rect -497 -53 -491 -19
rect -457 -53 -451 -19
rect -497 -91 -451 -53
rect -497 -125 -491 -91
rect -457 -125 -451 -91
rect -497 -163 -451 -125
rect -497 -197 -491 -163
rect -457 -197 -451 -163
rect -497 -235 -451 -197
rect -497 -269 -491 -235
rect -457 -269 -451 -235
rect -497 -307 -451 -269
rect -497 -341 -491 -307
rect -457 -341 -451 -307
rect -497 -379 -451 -341
rect -497 -413 -491 -379
rect -457 -413 -451 -379
rect -497 -451 -451 -413
rect -497 -485 -491 -451
rect -457 -485 -451 -451
rect -497 -500 -451 -485
rect -339 485 -293 500
rect -339 451 -333 485
rect -299 451 -293 485
rect -339 413 -293 451
rect -339 379 -333 413
rect -299 379 -293 413
rect -339 341 -293 379
rect -339 307 -333 341
rect -299 307 -293 341
rect -339 269 -293 307
rect -339 235 -333 269
rect -299 235 -293 269
rect -339 197 -293 235
rect -339 163 -333 197
rect -299 163 -293 197
rect -339 125 -293 163
rect -339 91 -333 125
rect -299 91 -293 125
rect -339 53 -293 91
rect -339 19 -333 53
rect -299 19 -293 53
rect -339 -19 -293 19
rect -339 -53 -333 -19
rect -299 -53 -293 -19
rect -339 -91 -293 -53
rect -339 -125 -333 -91
rect -299 -125 -293 -91
rect -339 -163 -293 -125
rect -339 -197 -333 -163
rect -299 -197 -293 -163
rect -339 -235 -293 -197
rect -339 -269 -333 -235
rect -299 -269 -293 -235
rect -339 -307 -293 -269
rect -339 -341 -333 -307
rect -299 -341 -293 -307
rect -339 -379 -293 -341
rect -339 -413 -333 -379
rect -299 -413 -293 -379
rect -339 -451 -293 -413
rect -339 -485 -333 -451
rect -299 -485 -293 -451
rect -339 -500 -293 -485
rect -181 485 -135 500
rect -181 451 -175 485
rect -141 451 -135 485
rect -181 413 -135 451
rect -181 379 -175 413
rect -141 379 -135 413
rect -181 341 -135 379
rect -181 307 -175 341
rect -141 307 -135 341
rect -181 269 -135 307
rect -181 235 -175 269
rect -141 235 -135 269
rect -181 197 -135 235
rect -181 163 -175 197
rect -141 163 -135 197
rect -181 125 -135 163
rect -181 91 -175 125
rect -141 91 -135 125
rect -181 53 -135 91
rect -181 19 -175 53
rect -141 19 -135 53
rect -181 -19 -135 19
rect -181 -53 -175 -19
rect -141 -53 -135 -19
rect -181 -91 -135 -53
rect -181 -125 -175 -91
rect -141 -125 -135 -91
rect -181 -163 -135 -125
rect -181 -197 -175 -163
rect -141 -197 -135 -163
rect -181 -235 -135 -197
rect -181 -269 -175 -235
rect -141 -269 -135 -235
rect -181 -307 -135 -269
rect -181 -341 -175 -307
rect -141 -341 -135 -307
rect -181 -379 -135 -341
rect -181 -413 -175 -379
rect -141 -413 -135 -379
rect -181 -451 -135 -413
rect -181 -485 -175 -451
rect -141 -485 -135 -451
rect -181 -500 -135 -485
rect -23 485 23 500
rect -23 451 -17 485
rect 17 451 23 485
rect -23 413 23 451
rect -23 379 -17 413
rect 17 379 23 413
rect -23 341 23 379
rect -23 307 -17 341
rect 17 307 23 341
rect -23 269 23 307
rect -23 235 -17 269
rect 17 235 23 269
rect -23 197 23 235
rect -23 163 -17 197
rect 17 163 23 197
rect -23 125 23 163
rect -23 91 -17 125
rect 17 91 23 125
rect -23 53 23 91
rect -23 19 -17 53
rect 17 19 23 53
rect -23 -19 23 19
rect -23 -53 -17 -19
rect 17 -53 23 -19
rect -23 -91 23 -53
rect -23 -125 -17 -91
rect 17 -125 23 -91
rect -23 -163 23 -125
rect -23 -197 -17 -163
rect 17 -197 23 -163
rect -23 -235 23 -197
rect -23 -269 -17 -235
rect 17 -269 23 -235
rect -23 -307 23 -269
rect -23 -341 -17 -307
rect 17 -341 23 -307
rect -23 -379 23 -341
rect -23 -413 -17 -379
rect 17 -413 23 -379
rect -23 -451 23 -413
rect -23 -485 -17 -451
rect 17 -485 23 -451
rect -23 -500 23 -485
rect 135 485 181 500
rect 135 451 141 485
rect 175 451 181 485
rect 135 413 181 451
rect 135 379 141 413
rect 175 379 181 413
rect 135 341 181 379
rect 135 307 141 341
rect 175 307 181 341
rect 135 269 181 307
rect 135 235 141 269
rect 175 235 181 269
rect 135 197 181 235
rect 135 163 141 197
rect 175 163 181 197
rect 135 125 181 163
rect 135 91 141 125
rect 175 91 181 125
rect 135 53 181 91
rect 135 19 141 53
rect 175 19 181 53
rect 135 -19 181 19
rect 135 -53 141 -19
rect 175 -53 181 -19
rect 135 -91 181 -53
rect 135 -125 141 -91
rect 175 -125 181 -91
rect 135 -163 181 -125
rect 135 -197 141 -163
rect 175 -197 181 -163
rect 135 -235 181 -197
rect 135 -269 141 -235
rect 175 -269 181 -235
rect 135 -307 181 -269
rect 135 -341 141 -307
rect 175 -341 181 -307
rect 135 -379 181 -341
rect 135 -413 141 -379
rect 175 -413 181 -379
rect 135 -451 181 -413
rect 135 -485 141 -451
rect 175 -485 181 -451
rect 135 -500 181 -485
rect 293 485 339 500
rect 293 451 299 485
rect 333 451 339 485
rect 293 413 339 451
rect 293 379 299 413
rect 333 379 339 413
rect 293 341 339 379
rect 293 307 299 341
rect 333 307 339 341
rect 293 269 339 307
rect 293 235 299 269
rect 333 235 339 269
rect 293 197 339 235
rect 293 163 299 197
rect 333 163 339 197
rect 293 125 339 163
rect 293 91 299 125
rect 333 91 339 125
rect 293 53 339 91
rect 293 19 299 53
rect 333 19 339 53
rect 293 -19 339 19
rect 293 -53 299 -19
rect 333 -53 339 -19
rect 293 -91 339 -53
rect 293 -125 299 -91
rect 333 -125 339 -91
rect 293 -163 339 -125
rect 293 -197 299 -163
rect 333 -197 339 -163
rect 293 -235 339 -197
rect 293 -269 299 -235
rect 333 -269 339 -235
rect 293 -307 339 -269
rect 293 -341 299 -307
rect 333 -341 339 -307
rect 293 -379 339 -341
rect 293 -413 299 -379
rect 333 -413 339 -379
rect 293 -451 339 -413
rect 293 -485 299 -451
rect 333 -485 339 -451
rect 293 -500 339 -485
rect 451 485 497 500
rect 451 451 457 485
rect 491 451 497 485
rect 451 413 497 451
rect 451 379 457 413
rect 491 379 497 413
rect 451 341 497 379
rect 451 307 457 341
rect 491 307 497 341
rect 451 269 497 307
rect 451 235 457 269
rect 491 235 497 269
rect 451 197 497 235
rect 451 163 457 197
rect 491 163 497 197
rect 451 125 497 163
rect 451 91 457 125
rect 491 91 497 125
rect 451 53 497 91
rect 451 19 457 53
rect 491 19 497 53
rect 451 -19 497 19
rect 451 -53 457 -19
rect 491 -53 497 -19
rect 451 -91 497 -53
rect 451 -125 457 -91
rect 491 -125 497 -91
rect 451 -163 497 -125
rect 451 -197 457 -163
rect 491 -197 497 -163
rect 451 -235 497 -197
rect 451 -269 457 -235
rect 491 -269 497 -235
rect 451 -307 497 -269
rect 451 -341 457 -307
rect 491 -341 497 -307
rect 451 -379 497 -341
rect 451 -413 457 -379
rect 491 -413 497 -379
rect 451 -451 497 -413
rect 451 -485 457 -451
rect 491 -485 497 -451
rect 451 -500 497 -485
rect 609 485 655 500
rect 609 451 615 485
rect 649 451 655 485
rect 609 413 655 451
rect 609 379 615 413
rect 649 379 655 413
rect 609 341 655 379
rect 609 307 615 341
rect 649 307 655 341
rect 609 269 655 307
rect 609 235 615 269
rect 649 235 655 269
rect 609 197 655 235
rect 609 163 615 197
rect 649 163 655 197
rect 609 125 655 163
rect 609 91 615 125
rect 649 91 655 125
rect 609 53 655 91
rect 609 19 615 53
rect 649 19 655 53
rect 609 -19 655 19
rect 609 -53 615 -19
rect 649 -53 655 -19
rect 609 -91 655 -53
rect 609 -125 615 -91
rect 649 -125 655 -91
rect 609 -163 655 -125
rect 609 -197 615 -163
rect 649 -197 655 -163
rect 609 -235 655 -197
rect 609 -269 615 -235
rect 649 -269 655 -235
rect 609 -307 655 -269
rect 609 -341 615 -307
rect 649 -341 655 -307
rect 609 -379 655 -341
rect 609 -413 615 -379
rect 649 -413 655 -379
rect 609 -451 655 -413
rect 609 -485 615 -451
rect 649 -485 655 -451
rect 609 -500 655 -485
rect 767 485 813 500
rect 767 451 773 485
rect 807 451 813 485
rect 767 413 813 451
rect 767 379 773 413
rect 807 379 813 413
rect 767 341 813 379
rect 767 307 773 341
rect 807 307 813 341
rect 767 269 813 307
rect 767 235 773 269
rect 807 235 813 269
rect 767 197 813 235
rect 767 163 773 197
rect 807 163 813 197
rect 767 125 813 163
rect 767 91 773 125
rect 807 91 813 125
rect 767 53 813 91
rect 767 19 773 53
rect 807 19 813 53
rect 767 -19 813 19
rect 767 -53 773 -19
rect 807 -53 813 -19
rect 767 -91 813 -53
rect 767 -125 773 -91
rect 807 -125 813 -91
rect 767 -163 813 -125
rect 767 -197 773 -163
rect 807 -197 813 -163
rect 767 -235 813 -197
rect 767 -269 773 -235
rect 807 -269 813 -235
rect 767 -307 813 -269
rect 767 -341 773 -307
rect 807 -341 813 -307
rect 767 -379 813 -341
rect 767 -413 773 -379
rect 807 -413 813 -379
rect 767 -451 813 -413
rect 767 -485 773 -451
rect 807 -485 813 -451
rect 767 -500 813 -485
rect 925 485 971 500
rect 925 451 931 485
rect 965 451 971 485
rect 925 413 971 451
rect 925 379 931 413
rect 965 379 971 413
rect 925 341 971 379
rect 925 307 931 341
rect 965 307 971 341
rect 925 269 971 307
rect 925 235 931 269
rect 965 235 971 269
rect 925 197 971 235
rect 925 163 931 197
rect 965 163 971 197
rect 925 125 971 163
rect 925 91 931 125
rect 965 91 971 125
rect 925 53 971 91
rect 925 19 931 53
rect 965 19 971 53
rect 925 -19 971 19
rect 925 -53 931 -19
rect 965 -53 971 -19
rect 925 -91 971 -53
rect 925 -125 931 -91
rect 965 -125 971 -91
rect 925 -163 971 -125
rect 925 -197 931 -163
rect 965 -197 971 -163
rect 925 -235 971 -197
rect 925 -269 931 -235
rect 965 -269 971 -235
rect 925 -307 971 -269
rect 925 -341 931 -307
rect 965 -341 971 -307
rect 925 -379 971 -341
rect 925 -413 931 -379
rect 965 -413 971 -379
rect 925 -451 971 -413
rect 925 -485 931 -451
rect 965 -485 971 -451
rect 925 -500 971 -485
rect 1083 485 1129 500
rect 1083 451 1089 485
rect 1123 451 1129 485
rect 1083 413 1129 451
rect 1083 379 1089 413
rect 1123 379 1129 413
rect 1083 341 1129 379
rect 1083 307 1089 341
rect 1123 307 1129 341
rect 1083 269 1129 307
rect 1083 235 1089 269
rect 1123 235 1129 269
rect 1083 197 1129 235
rect 1083 163 1089 197
rect 1123 163 1129 197
rect 1083 125 1129 163
rect 1083 91 1089 125
rect 1123 91 1129 125
rect 1083 53 1129 91
rect 1083 19 1089 53
rect 1123 19 1129 53
rect 1083 -19 1129 19
rect 1083 -53 1089 -19
rect 1123 -53 1129 -19
rect 1083 -91 1129 -53
rect 1083 -125 1089 -91
rect 1123 -125 1129 -91
rect 1083 -163 1129 -125
rect 1083 -197 1089 -163
rect 1123 -197 1129 -163
rect 1083 -235 1129 -197
rect 1083 -269 1089 -235
rect 1123 -269 1129 -235
rect 1083 -307 1129 -269
rect 1083 -341 1089 -307
rect 1123 -341 1129 -307
rect 1083 -379 1129 -341
rect 1083 -413 1089 -379
rect 1123 -413 1129 -379
rect 1083 -451 1129 -413
rect 1083 -485 1089 -451
rect 1123 -485 1129 -451
rect 1083 -500 1129 -485
rect 1241 485 1287 500
rect 1241 451 1247 485
rect 1281 451 1287 485
rect 1241 413 1287 451
rect 1241 379 1247 413
rect 1281 379 1287 413
rect 1241 341 1287 379
rect 1241 307 1247 341
rect 1281 307 1287 341
rect 1241 269 1287 307
rect 1241 235 1247 269
rect 1281 235 1287 269
rect 1241 197 1287 235
rect 1241 163 1247 197
rect 1281 163 1287 197
rect 1241 125 1287 163
rect 1241 91 1247 125
rect 1281 91 1287 125
rect 1241 53 1287 91
rect 1241 19 1247 53
rect 1281 19 1287 53
rect 1241 -19 1287 19
rect 1241 -53 1247 -19
rect 1281 -53 1287 -19
rect 1241 -91 1287 -53
rect 1241 -125 1247 -91
rect 1281 -125 1287 -91
rect 1241 -163 1287 -125
rect 1241 -197 1247 -163
rect 1281 -197 1287 -163
rect 1241 -235 1287 -197
rect 1241 -269 1247 -235
rect 1281 -269 1287 -235
rect 1241 -307 1287 -269
rect 1241 -341 1247 -307
rect 1281 -341 1287 -307
rect 1241 -379 1287 -341
rect 1241 -413 1247 -379
rect 1281 -413 1287 -379
rect 1241 -451 1287 -413
rect 1241 -485 1247 -451
rect 1281 -485 1287 -451
rect 1241 -500 1287 -485
rect 1399 485 1445 500
rect 1399 451 1405 485
rect 1439 451 1445 485
rect 1399 413 1445 451
rect 1399 379 1405 413
rect 1439 379 1445 413
rect 1399 341 1445 379
rect 1399 307 1405 341
rect 1439 307 1445 341
rect 1399 269 1445 307
rect 1399 235 1405 269
rect 1439 235 1445 269
rect 1399 197 1445 235
rect 1399 163 1405 197
rect 1439 163 1445 197
rect 1399 125 1445 163
rect 1399 91 1405 125
rect 1439 91 1445 125
rect 1399 53 1445 91
rect 1399 19 1405 53
rect 1439 19 1445 53
rect 1399 -19 1445 19
rect 1399 -53 1405 -19
rect 1439 -53 1445 -19
rect 1399 -91 1445 -53
rect 1399 -125 1405 -91
rect 1439 -125 1445 -91
rect 1399 -163 1445 -125
rect 1399 -197 1405 -163
rect 1439 -197 1445 -163
rect 1399 -235 1445 -197
rect 1399 -269 1405 -235
rect 1439 -269 1445 -235
rect 1399 -307 1445 -269
rect 1399 -341 1405 -307
rect 1439 -341 1445 -307
rect 1399 -379 1445 -341
rect 1399 -413 1405 -379
rect 1439 -413 1445 -379
rect 1399 -451 1445 -413
rect 1399 -485 1405 -451
rect 1439 -485 1445 -451
rect 1399 -500 1445 -485
rect 1557 485 1603 500
rect 1557 451 1563 485
rect 1597 451 1603 485
rect 1557 413 1603 451
rect 1557 379 1563 413
rect 1597 379 1603 413
rect 1557 341 1603 379
rect 1557 307 1563 341
rect 1597 307 1603 341
rect 1557 269 1603 307
rect 1557 235 1563 269
rect 1597 235 1603 269
rect 1557 197 1603 235
rect 1557 163 1563 197
rect 1597 163 1603 197
rect 1557 125 1603 163
rect 1557 91 1563 125
rect 1597 91 1603 125
rect 1557 53 1603 91
rect 1557 19 1563 53
rect 1597 19 1603 53
rect 1557 -19 1603 19
rect 1557 -53 1563 -19
rect 1597 -53 1603 -19
rect 1557 -91 1603 -53
rect 1557 -125 1563 -91
rect 1597 -125 1603 -91
rect 1557 -163 1603 -125
rect 1557 -197 1563 -163
rect 1597 -197 1603 -163
rect 1557 -235 1603 -197
rect 1557 -269 1563 -235
rect 1597 -269 1603 -235
rect 1557 -307 1603 -269
rect 1557 -341 1563 -307
rect 1597 -341 1603 -307
rect 1557 -379 1603 -341
rect 1557 -413 1563 -379
rect 1597 -413 1603 -379
rect 1557 -451 1603 -413
rect 1557 -485 1563 -451
rect 1597 -485 1603 -451
rect 1557 -500 1603 -485
rect 1715 485 1761 500
rect 1715 451 1721 485
rect 1755 451 1761 485
rect 1715 413 1761 451
rect 1715 379 1721 413
rect 1755 379 1761 413
rect 1715 341 1761 379
rect 1715 307 1721 341
rect 1755 307 1761 341
rect 1715 269 1761 307
rect 1715 235 1721 269
rect 1755 235 1761 269
rect 1715 197 1761 235
rect 1715 163 1721 197
rect 1755 163 1761 197
rect 1715 125 1761 163
rect 1715 91 1721 125
rect 1755 91 1761 125
rect 1715 53 1761 91
rect 1715 19 1721 53
rect 1755 19 1761 53
rect 1715 -19 1761 19
rect 1715 -53 1721 -19
rect 1755 -53 1761 -19
rect 1715 -91 1761 -53
rect 1715 -125 1721 -91
rect 1755 -125 1761 -91
rect 1715 -163 1761 -125
rect 1715 -197 1721 -163
rect 1755 -197 1761 -163
rect 1715 -235 1761 -197
rect 1715 -269 1721 -235
rect 1755 -269 1761 -235
rect 1715 -307 1761 -269
rect 1715 -341 1721 -307
rect 1755 -341 1761 -307
rect 1715 -379 1761 -341
rect 1715 -413 1721 -379
rect 1755 -413 1761 -379
rect 1715 -451 1761 -413
rect 1715 -485 1721 -451
rect 1755 -485 1761 -451
rect 1715 -500 1761 -485
rect 1873 485 1919 500
rect 1873 451 1879 485
rect 1913 451 1919 485
rect 1873 413 1919 451
rect 1873 379 1879 413
rect 1913 379 1919 413
rect 1873 341 1919 379
rect 1873 307 1879 341
rect 1913 307 1919 341
rect 1873 269 1919 307
rect 1873 235 1879 269
rect 1913 235 1919 269
rect 1873 197 1919 235
rect 1873 163 1879 197
rect 1913 163 1919 197
rect 1873 125 1919 163
rect 1873 91 1879 125
rect 1913 91 1919 125
rect 1873 53 1919 91
rect 1873 19 1879 53
rect 1913 19 1919 53
rect 1873 -19 1919 19
rect 1873 -53 1879 -19
rect 1913 -53 1919 -19
rect 1873 -91 1919 -53
rect 1873 -125 1879 -91
rect 1913 -125 1919 -91
rect 1873 -163 1919 -125
rect 1873 -197 1879 -163
rect 1913 -197 1919 -163
rect 1873 -235 1919 -197
rect 1873 -269 1879 -235
rect 1913 -269 1919 -235
rect 1873 -307 1919 -269
rect 1873 -341 1879 -307
rect 1913 -341 1919 -307
rect 1873 -379 1919 -341
rect 1873 -413 1879 -379
rect 1913 -413 1919 -379
rect 1873 -451 1919 -413
rect 1873 -485 1879 -451
rect 1913 -485 1919 -451
rect 1873 -500 1919 -485
rect 2031 485 2077 500
rect 2031 451 2037 485
rect 2071 451 2077 485
rect 2031 413 2077 451
rect 2031 379 2037 413
rect 2071 379 2077 413
rect 2031 341 2077 379
rect 2031 307 2037 341
rect 2071 307 2077 341
rect 2031 269 2077 307
rect 2031 235 2037 269
rect 2071 235 2077 269
rect 2031 197 2077 235
rect 2031 163 2037 197
rect 2071 163 2077 197
rect 2031 125 2077 163
rect 2031 91 2037 125
rect 2071 91 2077 125
rect 2031 53 2077 91
rect 2031 19 2037 53
rect 2071 19 2077 53
rect 2031 -19 2077 19
rect 2031 -53 2037 -19
rect 2071 -53 2077 -19
rect 2031 -91 2077 -53
rect 2031 -125 2037 -91
rect 2071 -125 2077 -91
rect 2031 -163 2077 -125
rect 2031 -197 2037 -163
rect 2071 -197 2077 -163
rect 2031 -235 2077 -197
rect 2031 -269 2037 -235
rect 2071 -269 2077 -235
rect 2031 -307 2077 -269
rect 2031 -341 2037 -307
rect 2071 -341 2077 -307
rect 2031 -379 2077 -341
rect 2031 -413 2037 -379
rect 2071 -413 2077 -379
rect 2031 -451 2077 -413
rect 2031 -485 2037 -451
rect 2071 -485 2077 -451
rect 2031 -500 2077 -485
rect 2189 485 2235 500
rect 2189 451 2195 485
rect 2229 451 2235 485
rect 2189 413 2235 451
rect 2189 379 2195 413
rect 2229 379 2235 413
rect 2189 341 2235 379
rect 2189 307 2195 341
rect 2229 307 2235 341
rect 2189 269 2235 307
rect 2189 235 2195 269
rect 2229 235 2235 269
rect 2189 197 2235 235
rect 2189 163 2195 197
rect 2229 163 2235 197
rect 2189 125 2235 163
rect 2189 91 2195 125
rect 2229 91 2235 125
rect 2189 53 2235 91
rect 2189 19 2195 53
rect 2229 19 2235 53
rect 2189 -19 2235 19
rect 2189 -53 2195 -19
rect 2229 -53 2235 -19
rect 2189 -91 2235 -53
rect 2189 -125 2195 -91
rect 2229 -125 2235 -91
rect 2189 -163 2235 -125
rect 2189 -197 2195 -163
rect 2229 -197 2235 -163
rect 2189 -235 2235 -197
rect 2189 -269 2195 -235
rect 2229 -269 2235 -235
rect 2189 -307 2235 -269
rect 2189 -341 2195 -307
rect 2229 -341 2235 -307
rect 2189 -379 2235 -341
rect 2189 -413 2195 -379
rect 2229 -413 2235 -379
rect 2189 -451 2235 -413
rect 2189 -485 2195 -451
rect 2229 -485 2235 -451
rect 2189 -500 2235 -485
rect 2347 485 2393 500
rect 2347 451 2353 485
rect 2387 451 2393 485
rect 2347 413 2393 451
rect 2347 379 2353 413
rect 2387 379 2393 413
rect 2347 341 2393 379
rect 2347 307 2353 341
rect 2387 307 2393 341
rect 2347 269 2393 307
rect 2347 235 2353 269
rect 2387 235 2393 269
rect 2347 197 2393 235
rect 2347 163 2353 197
rect 2387 163 2393 197
rect 2347 125 2393 163
rect 2347 91 2353 125
rect 2387 91 2393 125
rect 2347 53 2393 91
rect 2347 19 2353 53
rect 2387 19 2393 53
rect 2347 -19 2393 19
rect 2347 -53 2353 -19
rect 2387 -53 2393 -19
rect 2347 -91 2393 -53
rect 2347 -125 2353 -91
rect 2387 -125 2393 -91
rect 2347 -163 2393 -125
rect 2347 -197 2353 -163
rect 2387 -197 2393 -163
rect 2347 -235 2393 -197
rect 2347 -269 2353 -235
rect 2387 -269 2393 -235
rect 2347 -307 2393 -269
rect 2347 -341 2353 -307
rect 2387 -341 2393 -307
rect 2347 -379 2393 -341
rect 2347 -413 2353 -379
rect 2387 -413 2393 -379
rect 2347 -451 2393 -413
rect 2347 -485 2353 -451
rect 2387 -485 2393 -451
rect 2347 -500 2393 -485
rect 2505 485 2551 500
rect 2505 451 2511 485
rect 2545 451 2551 485
rect 2505 413 2551 451
rect 2505 379 2511 413
rect 2545 379 2551 413
rect 2505 341 2551 379
rect 2505 307 2511 341
rect 2545 307 2551 341
rect 2505 269 2551 307
rect 2505 235 2511 269
rect 2545 235 2551 269
rect 2505 197 2551 235
rect 2505 163 2511 197
rect 2545 163 2551 197
rect 2505 125 2551 163
rect 2505 91 2511 125
rect 2545 91 2551 125
rect 2505 53 2551 91
rect 2505 19 2511 53
rect 2545 19 2551 53
rect 2505 -19 2551 19
rect 2505 -53 2511 -19
rect 2545 -53 2551 -19
rect 2505 -91 2551 -53
rect 2505 -125 2511 -91
rect 2545 -125 2551 -91
rect 2505 -163 2551 -125
rect 2505 -197 2511 -163
rect 2545 -197 2551 -163
rect 2505 -235 2551 -197
rect 2505 -269 2511 -235
rect 2545 -269 2551 -235
rect 2505 -307 2551 -269
rect 2505 -341 2511 -307
rect 2545 -341 2551 -307
rect 2505 -379 2551 -341
rect 2505 -413 2511 -379
rect 2545 -413 2551 -379
rect 2505 -451 2551 -413
rect 2505 -485 2511 -451
rect 2545 -485 2551 -451
rect 2505 -500 2551 -485
rect 2663 485 2709 500
rect 2663 451 2669 485
rect 2703 451 2709 485
rect 2663 413 2709 451
rect 2663 379 2669 413
rect 2703 379 2709 413
rect 2663 341 2709 379
rect 2663 307 2669 341
rect 2703 307 2709 341
rect 2663 269 2709 307
rect 2663 235 2669 269
rect 2703 235 2709 269
rect 2663 197 2709 235
rect 2663 163 2669 197
rect 2703 163 2709 197
rect 2663 125 2709 163
rect 2663 91 2669 125
rect 2703 91 2709 125
rect 2663 53 2709 91
rect 2663 19 2669 53
rect 2703 19 2709 53
rect 2663 -19 2709 19
rect 2663 -53 2669 -19
rect 2703 -53 2709 -19
rect 2663 -91 2709 -53
rect 2663 -125 2669 -91
rect 2703 -125 2709 -91
rect 2663 -163 2709 -125
rect 2663 -197 2669 -163
rect 2703 -197 2709 -163
rect 2663 -235 2709 -197
rect 2663 -269 2669 -235
rect 2703 -269 2709 -235
rect 2663 -307 2709 -269
rect 2663 -341 2669 -307
rect 2703 -341 2709 -307
rect 2663 -379 2709 -341
rect 2663 -413 2669 -379
rect 2703 -413 2709 -379
rect 2663 -451 2709 -413
rect 2663 -485 2669 -451
rect 2703 -485 2709 -451
rect 2663 -500 2709 -485
rect 2821 485 2867 500
rect 2821 451 2827 485
rect 2861 451 2867 485
rect 2821 413 2867 451
rect 2821 379 2827 413
rect 2861 379 2867 413
rect 2821 341 2867 379
rect 2821 307 2827 341
rect 2861 307 2867 341
rect 2821 269 2867 307
rect 2821 235 2827 269
rect 2861 235 2867 269
rect 2821 197 2867 235
rect 2821 163 2827 197
rect 2861 163 2867 197
rect 2821 125 2867 163
rect 2821 91 2827 125
rect 2861 91 2867 125
rect 2821 53 2867 91
rect 2821 19 2827 53
rect 2861 19 2867 53
rect 2821 -19 2867 19
rect 2821 -53 2827 -19
rect 2861 -53 2867 -19
rect 2821 -91 2867 -53
rect 2821 -125 2827 -91
rect 2861 -125 2867 -91
rect 2821 -163 2867 -125
rect 2821 -197 2827 -163
rect 2861 -197 2867 -163
rect 2821 -235 2867 -197
rect 2821 -269 2827 -235
rect 2861 -269 2867 -235
rect 2821 -307 2867 -269
rect 2821 -341 2827 -307
rect 2861 -341 2867 -307
rect 2821 -379 2867 -341
rect 2821 -413 2827 -379
rect 2861 -413 2867 -379
rect 2821 -451 2867 -413
rect 2821 -485 2827 -451
rect 2861 -485 2867 -451
rect 2821 -500 2867 -485
rect 2979 485 3025 500
rect 2979 451 2985 485
rect 3019 451 3025 485
rect 2979 413 3025 451
rect 2979 379 2985 413
rect 3019 379 3025 413
rect 2979 341 3025 379
rect 2979 307 2985 341
rect 3019 307 3025 341
rect 2979 269 3025 307
rect 2979 235 2985 269
rect 3019 235 3025 269
rect 2979 197 3025 235
rect 2979 163 2985 197
rect 3019 163 3025 197
rect 2979 125 3025 163
rect 2979 91 2985 125
rect 3019 91 3025 125
rect 2979 53 3025 91
rect 2979 19 2985 53
rect 3019 19 3025 53
rect 2979 -19 3025 19
rect 2979 -53 2985 -19
rect 3019 -53 3025 -19
rect 2979 -91 3025 -53
rect 2979 -125 2985 -91
rect 3019 -125 3025 -91
rect 2979 -163 3025 -125
rect 2979 -197 2985 -163
rect 3019 -197 3025 -163
rect 2979 -235 3025 -197
rect 2979 -269 2985 -235
rect 3019 -269 3025 -235
rect 2979 -307 3025 -269
rect 2979 -341 2985 -307
rect 3019 -341 3025 -307
rect 2979 -379 3025 -341
rect 2979 -413 2985 -379
rect 3019 -413 3025 -379
rect 2979 -451 3025 -413
rect 2979 -485 2985 -451
rect 3019 -485 3025 -451
rect 2979 -500 3025 -485
rect 3137 485 3183 500
rect 3137 451 3143 485
rect 3177 451 3183 485
rect 3137 413 3183 451
rect 3137 379 3143 413
rect 3177 379 3183 413
rect 3137 341 3183 379
rect 3137 307 3143 341
rect 3177 307 3183 341
rect 3137 269 3183 307
rect 3137 235 3143 269
rect 3177 235 3183 269
rect 3137 197 3183 235
rect 3137 163 3143 197
rect 3177 163 3183 197
rect 3137 125 3183 163
rect 3137 91 3143 125
rect 3177 91 3183 125
rect 3137 53 3183 91
rect 3137 19 3143 53
rect 3177 19 3183 53
rect 3137 -19 3183 19
rect 3137 -53 3143 -19
rect 3177 -53 3183 -19
rect 3137 -91 3183 -53
rect 3137 -125 3143 -91
rect 3177 -125 3183 -91
rect 3137 -163 3183 -125
rect 3137 -197 3143 -163
rect 3177 -197 3183 -163
rect 3137 -235 3183 -197
rect 3137 -269 3143 -235
rect 3177 -269 3183 -235
rect 3137 -307 3183 -269
rect 3137 -341 3143 -307
rect 3177 -341 3183 -307
rect 3137 -379 3183 -341
rect 3137 -413 3143 -379
rect 3177 -413 3183 -379
rect 3137 -451 3183 -413
rect 3137 -485 3143 -451
rect 3177 -485 3183 -451
rect 3137 -500 3183 -485
rect -3127 -547 -3035 -541
rect -3127 -581 -3098 -547
rect -3064 -581 -3035 -547
rect -3127 -587 -3035 -581
rect -2969 -547 -2877 -541
rect -2969 -581 -2940 -547
rect -2906 -581 -2877 -547
rect -2969 -587 -2877 -581
rect -2811 -547 -2719 -541
rect -2811 -581 -2782 -547
rect -2748 -581 -2719 -547
rect -2811 -587 -2719 -581
rect -2653 -547 -2561 -541
rect -2653 -581 -2624 -547
rect -2590 -581 -2561 -547
rect -2653 -587 -2561 -581
rect -2495 -547 -2403 -541
rect -2495 -581 -2466 -547
rect -2432 -581 -2403 -547
rect -2495 -587 -2403 -581
rect -2337 -547 -2245 -541
rect -2337 -581 -2308 -547
rect -2274 -581 -2245 -547
rect -2337 -587 -2245 -581
rect -2179 -547 -2087 -541
rect -2179 -581 -2150 -547
rect -2116 -581 -2087 -547
rect -2179 -587 -2087 -581
rect -2021 -547 -1929 -541
rect -2021 -581 -1992 -547
rect -1958 -581 -1929 -547
rect -2021 -587 -1929 -581
rect -1863 -547 -1771 -541
rect -1863 -581 -1834 -547
rect -1800 -581 -1771 -547
rect -1863 -587 -1771 -581
rect -1705 -547 -1613 -541
rect -1705 -581 -1676 -547
rect -1642 -581 -1613 -547
rect -1705 -587 -1613 -581
rect -1547 -547 -1455 -541
rect -1547 -581 -1518 -547
rect -1484 -581 -1455 -547
rect -1547 -587 -1455 -581
rect -1389 -547 -1297 -541
rect -1389 -581 -1360 -547
rect -1326 -581 -1297 -547
rect -1389 -587 -1297 -581
rect -1231 -547 -1139 -541
rect -1231 -581 -1202 -547
rect -1168 -581 -1139 -547
rect -1231 -587 -1139 -581
rect -1073 -547 -981 -541
rect -1073 -581 -1044 -547
rect -1010 -581 -981 -547
rect -1073 -587 -981 -581
rect -915 -547 -823 -541
rect -915 -581 -886 -547
rect -852 -581 -823 -547
rect -915 -587 -823 -581
rect -757 -547 -665 -541
rect -757 -581 -728 -547
rect -694 -581 -665 -547
rect -757 -587 -665 -581
rect -599 -547 -507 -541
rect -599 -581 -570 -547
rect -536 -581 -507 -547
rect -599 -587 -507 -581
rect -441 -547 -349 -541
rect -441 -581 -412 -547
rect -378 -581 -349 -547
rect -441 -587 -349 -581
rect -283 -547 -191 -541
rect -283 -581 -254 -547
rect -220 -581 -191 -547
rect -283 -587 -191 -581
rect -125 -547 -33 -541
rect -125 -581 -96 -547
rect -62 -581 -33 -547
rect -125 -587 -33 -581
rect 33 -547 125 -541
rect 33 -581 62 -547
rect 96 -581 125 -547
rect 33 -587 125 -581
rect 191 -547 283 -541
rect 191 -581 220 -547
rect 254 -581 283 -547
rect 191 -587 283 -581
rect 349 -547 441 -541
rect 349 -581 378 -547
rect 412 -581 441 -547
rect 349 -587 441 -581
rect 507 -547 599 -541
rect 507 -581 536 -547
rect 570 -581 599 -547
rect 507 -587 599 -581
rect 665 -547 757 -541
rect 665 -581 694 -547
rect 728 -581 757 -547
rect 665 -587 757 -581
rect 823 -547 915 -541
rect 823 -581 852 -547
rect 886 -581 915 -547
rect 823 -587 915 -581
rect 981 -547 1073 -541
rect 981 -581 1010 -547
rect 1044 -581 1073 -547
rect 981 -587 1073 -581
rect 1139 -547 1231 -541
rect 1139 -581 1168 -547
rect 1202 -581 1231 -547
rect 1139 -587 1231 -581
rect 1297 -547 1389 -541
rect 1297 -581 1326 -547
rect 1360 -581 1389 -547
rect 1297 -587 1389 -581
rect 1455 -547 1547 -541
rect 1455 -581 1484 -547
rect 1518 -581 1547 -547
rect 1455 -587 1547 -581
rect 1613 -547 1705 -541
rect 1613 -581 1642 -547
rect 1676 -581 1705 -547
rect 1613 -587 1705 -581
rect 1771 -547 1863 -541
rect 1771 -581 1800 -547
rect 1834 -581 1863 -547
rect 1771 -587 1863 -581
rect 1929 -547 2021 -541
rect 1929 -581 1958 -547
rect 1992 -581 2021 -547
rect 1929 -587 2021 -581
rect 2087 -547 2179 -541
rect 2087 -581 2116 -547
rect 2150 -581 2179 -547
rect 2087 -587 2179 -581
rect 2245 -547 2337 -541
rect 2245 -581 2274 -547
rect 2308 -581 2337 -547
rect 2245 -587 2337 -581
rect 2403 -547 2495 -541
rect 2403 -581 2432 -547
rect 2466 -581 2495 -547
rect 2403 -587 2495 -581
rect 2561 -547 2653 -541
rect 2561 -581 2590 -547
rect 2624 -581 2653 -547
rect 2561 -587 2653 -581
rect 2719 -547 2811 -541
rect 2719 -581 2748 -547
rect 2782 -581 2811 -547
rect 2719 -587 2811 -581
rect 2877 -547 2969 -541
rect 2877 -581 2906 -547
rect 2940 -581 2969 -547
rect 2877 -587 2969 -581
rect 3035 -547 3127 -541
rect 3035 -581 3064 -547
rect 3098 -581 3127 -547
rect 3035 -587 3127 -581
rect -1640 -649 1640 -643
rect -1640 -683 -1601 -649
rect -1567 -683 -1529 -649
rect -1495 -683 -1457 -649
rect -1423 -683 -1385 -649
rect -1351 -683 -1313 -649
rect -1279 -683 -1241 -649
rect -1207 -683 -1169 -649
rect -1135 -683 -1097 -649
rect -1063 -683 -1025 -649
rect -991 -683 -953 -649
rect -919 -683 -881 -649
rect -847 -683 -809 -649
rect -775 -683 -737 -649
rect -703 -683 -665 -649
rect -631 -683 -593 -649
rect -559 -683 -521 -649
rect -487 -683 -449 -649
rect -415 -683 -377 -649
rect -343 -683 -305 -649
rect -271 -683 -233 -649
rect -199 -683 -161 -649
rect -127 -683 -89 -649
rect -55 -683 -17 -649
rect 17 -683 55 -649
rect 89 -683 127 -649
rect 161 -683 199 -649
rect 233 -683 271 -649
rect 305 -683 343 -649
rect 377 -683 415 -649
rect 449 -683 487 -649
rect 521 -683 559 -649
rect 593 -683 631 -649
rect 665 -683 703 -649
rect 737 -683 775 -649
rect 809 -683 847 -649
rect 881 -683 919 -649
rect 953 -683 991 -649
rect 1025 -683 1063 -649
rect 1097 -683 1135 -649
rect 1169 -683 1207 -649
rect 1241 -683 1279 -649
rect 1313 -683 1351 -649
rect 1385 -683 1423 -649
rect 1457 -683 1495 -649
rect 1529 -683 1567 -649
rect 1601 -683 1640 -649
rect -1640 -689 1640 -683
<< properties >>
string FIXED_BBOX -3274 -666 3274 666
<< end >>
