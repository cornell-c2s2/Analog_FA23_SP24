magic
tech sky130A
magscale 1 2
timestamp 1713140669
<< pwell >>
rect -1715 -710 1715 710
<< nmos >>
rect -1519 -500 -1319 500
rect -1261 -500 -1061 500
rect -1003 -500 -803 500
rect -745 -500 -545 500
rect -487 -500 -287 500
rect -229 -500 -29 500
rect 29 -500 229 500
rect 287 -500 487 500
rect 545 -500 745 500
rect 803 -500 1003 500
rect 1061 -500 1261 500
rect 1319 -500 1519 500
<< ndiff >>
rect -1577 488 -1519 500
rect -1577 -488 -1565 488
rect -1531 -488 -1519 488
rect -1577 -500 -1519 -488
rect -1319 488 -1261 500
rect -1319 -488 -1307 488
rect -1273 -488 -1261 488
rect -1319 -500 -1261 -488
rect -1061 488 -1003 500
rect -1061 -488 -1049 488
rect -1015 -488 -1003 488
rect -1061 -500 -1003 -488
rect -803 488 -745 500
rect -803 -488 -791 488
rect -757 -488 -745 488
rect -803 -500 -745 -488
rect -545 488 -487 500
rect -545 -488 -533 488
rect -499 -488 -487 488
rect -545 -500 -487 -488
rect -287 488 -229 500
rect -287 -488 -275 488
rect -241 -488 -229 488
rect -287 -500 -229 -488
rect -29 488 29 500
rect -29 -488 -17 488
rect 17 -488 29 488
rect -29 -500 29 -488
rect 229 488 287 500
rect 229 -488 241 488
rect 275 -488 287 488
rect 229 -500 287 -488
rect 487 488 545 500
rect 487 -488 499 488
rect 533 -488 545 488
rect 487 -500 545 -488
rect 745 488 803 500
rect 745 -488 757 488
rect 791 -488 803 488
rect 745 -500 803 -488
rect 1003 488 1061 500
rect 1003 -488 1015 488
rect 1049 -488 1061 488
rect 1003 -500 1061 -488
rect 1261 488 1319 500
rect 1261 -488 1273 488
rect 1307 -488 1319 488
rect 1261 -500 1319 -488
rect 1519 488 1577 500
rect 1519 -488 1531 488
rect 1565 -488 1577 488
rect 1519 -500 1577 -488
<< ndiffc >>
rect -1565 -488 -1531 488
rect -1307 -488 -1273 488
rect -1049 -488 -1015 488
rect -791 -488 -757 488
rect -533 -488 -499 488
rect -275 -488 -241 488
rect -17 -488 17 488
rect 241 -488 275 488
rect 499 -488 533 488
rect 757 -488 791 488
rect 1015 -488 1049 488
rect 1273 -488 1307 488
rect 1531 -488 1565 488
<< psubdiff >>
rect -1679 640 -1583 674
rect 1583 640 1679 674
rect -1679 578 -1645 640
rect 1645 578 1679 640
rect -1679 -640 -1645 -578
rect 1645 -640 1679 -578
rect -1679 -674 -1583 -640
rect 1583 -674 1679 -640
<< psubdiffcont >>
rect -1583 640 1583 674
rect -1679 -578 -1645 578
rect 1645 -578 1679 578
rect -1583 -674 1583 -640
<< poly >>
rect -1519 572 -1319 588
rect -1519 538 -1503 572
rect -1335 538 -1319 572
rect -1519 500 -1319 538
rect -1261 572 -1061 588
rect -1261 538 -1245 572
rect -1077 538 -1061 572
rect -1261 500 -1061 538
rect -1003 572 -803 588
rect -1003 538 -987 572
rect -819 538 -803 572
rect -1003 500 -803 538
rect -745 572 -545 588
rect -745 538 -729 572
rect -561 538 -545 572
rect -745 500 -545 538
rect -487 572 -287 588
rect -487 538 -471 572
rect -303 538 -287 572
rect -487 500 -287 538
rect -229 572 -29 588
rect -229 538 -213 572
rect -45 538 -29 572
rect -229 500 -29 538
rect 29 572 229 588
rect 29 538 45 572
rect 213 538 229 572
rect 29 500 229 538
rect 287 572 487 588
rect 287 538 303 572
rect 471 538 487 572
rect 287 500 487 538
rect 545 572 745 588
rect 545 538 561 572
rect 729 538 745 572
rect 545 500 745 538
rect 803 572 1003 588
rect 803 538 819 572
rect 987 538 1003 572
rect 803 500 1003 538
rect 1061 572 1261 588
rect 1061 538 1077 572
rect 1245 538 1261 572
rect 1061 500 1261 538
rect 1319 572 1519 588
rect 1319 538 1335 572
rect 1503 538 1519 572
rect 1319 500 1519 538
rect -1519 -538 -1319 -500
rect -1519 -572 -1503 -538
rect -1335 -572 -1319 -538
rect -1519 -588 -1319 -572
rect -1261 -538 -1061 -500
rect -1261 -572 -1245 -538
rect -1077 -572 -1061 -538
rect -1261 -588 -1061 -572
rect -1003 -538 -803 -500
rect -1003 -572 -987 -538
rect -819 -572 -803 -538
rect -1003 -588 -803 -572
rect -745 -538 -545 -500
rect -745 -572 -729 -538
rect -561 -572 -545 -538
rect -745 -588 -545 -572
rect -487 -538 -287 -500
rect -487 -572 -471 -538
rect -303 -572 -287 -538
rect -487 -588 -287 -572
rect -229 -538 -29 -500
rect -229 -572 -213 -538
rect -45 -572 -29 -538
rect -229 -588 -29 -572
rect 29 -538 229 -500
rect 29 -572 45 -538
rect 213 -572 229 -538
rect 29 -588 229 -572
rect 287 -538 487 -500
rect 287 -572 303 -538
rect 471 -572 487 -538
rect 287 -588 487 -572
rect 545 -538 745 -500
rect 545 -572 561 -538
rect 729 -572 745 -538
rect 545 -588 745 -572
rect 803 -538 1003 -500
rect 803 -572 819 -538
rect 987 -572 1003 -538
rect 803 -588 1003 -572
rect 1061 -538 1261 -500
rect 1061 -572 1077 -538
rect 1245 -572 1261 -538
rect 1061 -588 1261 -572
rect 1319 -538 1519 -500
rect 1319 -572 1335 -538
rect 1503 -572 1519 -538
rect 1319 -588 1519 -572
<< polycont >>
rect -1503 538 -1335 572
rect -1245 538 -1077 572
rect -987 538 -819 572
rect -729 538 -561 572
rect -471 538 -303 572
rect -213 538 -45 572
rect 45 538 213 572
rect 303 538 471 572
rect 561 538 729 572
rect 819 538 987 572
rect 1077 538 1245 572
rect 1335 538 1503 572
rect -1503 -572 -1335 -538
rect -1245 -572 -1077 -538
rect -987 -572 -819 -538
rect -729 -572 -561 -538
rect -471 -572 -303 -538
rect -213 -572 -45 -538
rect 45 -572 213 -538
rect 303 -572 471 -538
rect 561 -572 729 -538
rect 819 -572 987 -538
rect 1077 -572 1245 -538
rect 1335 -572 1503 -538
<< locali >>
rect -1679 640 -1583 674
rect 1583 640 1679 674
rect -1679 578 -1645 640
rect 1645 578 1679 640
rect -1519 538 -1503 572
rect -1335 538 -1319 572
rect -1261 538 -1245 572
rect -1077 538 -1061 572
rect -1003 538 -987 572
rect -819 538 -803 572
rect -745 538 -729 572
rect -561 538 -545 572
rect -487 538 -471 572
rect -303 538 -287 572
rect -229 538 -213 572
rect -45 538 -29 572
rect 29 538 45 572
rect 213 538 229 572
rect 287 538 303 572
rect 471 538 487 572
rect 545 538 561 572
rect 729 538 745 572
rect 803 538 819 572
rect 987 538 1003 572
rect 1061 538 1077 572
rect 1245 538 1261 572
rect 1319 538 1335 572
rect 1503 538 1519 572
rect -1565 488 -1531 504
rect -1565 -504 -1531 -488
rect -1307 488 -1273 504
rect -1307 -504 -1273 -488
rect -1049 488 -1015 504
rect -1049 -504 -1015 -488
rect -791 488 -757 504
rect -791 -504 -757 -488
rect -533 488 -499 504
rect -533 -504 -499 -488
rect -275 488 -241 504
rect -275 -504 -241 -488
rect -17 488 17 504
rect -17 -504 17 -488
rect 241 488 275 504
rect 241 -504 275 -488
rect 499 488 533 504
rect 499 -504 533 -488
rect 757 488 791 504
rect 757 -504 791 -488
rect 1015 488 1049 504
rect 1015 -504 1049 -488
rect 1273 488 1307 504
rect 1273 -504 1307 -488
rect 1531 488 1565 504
rect 1531 -504 1565 -488
rect -1519 -572 -1503 -538
rect -1335 -572 -1319 -538
rect -1261 -572 -1245 -538
rect -1077 -572 -1061 -538
rect -1003 -572 -987 -538
rect -819 -572 -803 -538
rect -745 -572 -729 -538
rect -561 -572 -545 -538
rect -487 -572 -471 -538
rect -303 -572 -287 -538
rect -229 -572 -213 -538
rect -45 -572 -29 -538
rect 29 -572 45 -538
rect 213 -572 229 -538
rect 287 -572 303 -538
rect 471 -572 487 -538
rect 545 -572 561 -538
rect 729 -572 745 -538
rect 803 -572 819 -538
rect 987 -572 1003 -538
rect 1061 -572 1077 -538
rect 1245 -572 1261 -538
rect 1319 -572 1335 -538
rect 1503 -572 1519 -538
rect -1679 -640 -1645 -578
rect 1645 -640 1679 -578
rect -1679 -674 -1583 -640
rect 1583 -674 1679 -640
<< viali >>
rect -1503 538 -1335 572
rect -1245 538 -1077 572
rect -987 538 -819 572
rect -729 538 -561 572
rect -471 538 -303 572
rect -213 538 -45 572
rect 45 538 213 572
rect 303 538 471 572
rect 561 538 729 572
rect 819 538 987 572
rect 1077 538 1245 572
rect 1335 538 1503 572
rect -1565 -488 -1531 488
rect -1307 -488 -1273 488
rect -1049 -488 -1015 488
rect -791 -488 -757 488
rect -533 -488 -499 488
rect -275 -488 -241 488
rect -17 -488 17 488
rect 241 -488 275 488
rect 499 -488 533 488
rect 757 -488 791 488
rect 1015 -488 1049 488
rect 1273 -488 1307 488
rect 1531 -488 1565 488
rect -1503 -572 -1335 -538
rect -1245 -572 -1077 -538
rect -987 -572 -819 -538
rect -729 -572 -561 -538
rect -471 -572 -303 -538
rect -213 -572 -45 -538
rect 45 -572 213 -538
rect 303 -572 471 -538
rect 561 -572 729 -538
rect 819 -572 987 -538
rect 1077 -572 1245 -538
rect 1335 -572 1503 -538
<< metal1 >>
rect -1515 572 -1323 578
rect -1515 538 -1503 572
rect -1335 538 -1323 572
rect -1515 532 -1323 538
rect -1257 572 -1065 578
rect -1257 538 -1245 572
rect -1077 538 -1065 572
rect -1257 532 -1065 538
rect -999 572 -807 578
rect -999 538 -987 572
rect -819 538 -807 572
rect -999 532 -807 538
rect -741 572 -549 578
rect -741 538 -729 572
rect -561 538 -549 572
rect -741 532 -549 538
rect -483 572 -291 578
rect -483 538 -471 572
rect -303 538 -291 572
rect -483 532 -291 538
rect -225 572 -33 578
rect -225 538 -213 572
rect -45 538 -33 572
rect -225 532 -33 538
rect 33 572 225 578
rect 33 538 45 572
rect 213 538 225 572
rect 33 532 225 538
rect 291 572 483 578
rect 291 538 303 572
rect 471 538 483 572
rect 291 532 483 538
rect 549 572 741 578
rect 549 538 561 572
rect 729 538 741 572
rect 549 532 741 538
rect 807 572 999 578
rect 807 538 819 572
rect 987 538 999 572
rect 807 532 999 538
rect 1065 572 1257 578
rect 1065 538 1077 572
rect 1245 538 1257 572
rect 1065 532 1257 538
rect 1323 572 1515 578
rect 1323 538 1335 572
rect 1503 538 1515 572
rect 1323 532 1515 538
rect -1571 488 -1525 500
rect -1571 -488 -1565 488
rect -1531 -488 -1525 488
rect -1571 -500 -1525 -488
rect -1313 488 -1267 500
rect -1313 -488 -1307 488
rect -1273 -488 -1267 488
rect -1313 -500 -1267 -488
rect -1055 488 -1009 500
rect -1055 -488 -1049 488
rect -1015 -488 -1009 488
rect -1055 -500 -1009 -488
rect -797 488 -751 500
rect -797 -488 -791 488
rect -757 -488 -751 488
rect -797 -500 -751 -488
rect -539 488 -493 500
rect -539 -488 -533 488
rect -499 -488 -493 488
rect -539 -500 -493 -488
rect -281 488 -235 500
rect -281 -488 -275 488
rect -241 -488 -235 488
rect -281 -500 -235 -488
rect -23 488 23 500
rect -23 -488 -17 488
rect 17 -488 23 488
rect -23 -500 23 -488
rect 235 488 281 500
rect 235 -488 241 488
rect 275 -488 281 488
rect 235 -500 281 -488
rect 493 488 539 500
rect 493 -488 499 488
rect 533 -488 539 488
rect 493 -500 539 -488
rect 751 488 797 500
rect 751 -488 757 488
rect 791 -488 797 488
rect 751 -500 797 -488
rect 1009 488 1055 500
rect 1009 -488 1015 488
rect 1049 -488 1055 488
rect 1009 -500 1055 -488
rect 1267 488 1313 500
rect 1267 -488 1273 488
rect 1307 -488 1313 488
rect 1267 -500 1313 -488
rect 1525 488 1571 500
rect 1525 -488 1531 488
rect 1565 -488 1571 488
rect 1525 -500 1571 -488
rect -1515 -538 -1323 -532
rect -1515 -572 -1503 -538
rect -1335 -572 -1323 -538
rect -1515 -578 -1323 -572
rect -1257 -538 -1065 -532
rect -1257 -572 -1245 -538
rect -1077 -572 -1065 -538
rect -1257 -578 -1065 -572
rect -999 -538 -807 -532
rect -999 -572 -987 -538
rect -819 -572 -807 -538
rect -999 -578 -807 -572
rect -741 -538 -549 -532
rect -741 -572 -729 -538
rect -561 -572 -549 -538
rect -741 -578 -549 -572
rect -483 -538 -291 -532
rect -483 -572 -471 -538
rect -303 -572 -291 -538
rect -483 -578 -291 -572
rect -225 -538 -33 -532
rect -225 -572 -213 -538
rect -45 -572 -33 -538
rect -225 -578 -33 -572
rect 33 -538 225 -532
rect 33 -572 45 -538
rect 213 -572 225 -538
rect 33 -578 225 -572
rect 291 -538 483 -532
rect 291 -572 303 -538
rect 471 -572 483 -538
rect 291 -578 483 -572
rect 549 -538 741 -532
rect 549 -572 561 -538
rect 729 -572 741 -538
rect 549 -578 741 -572
rect 807 -538 999 -532
rect 807 -572 819 -538
rect 987 -572 999 -538
rect 807 -578 999 -572
rect 1065 -538 1257 -532
rect 1065 -572 1077 -538
rect 1245 -572 1257 -538
rect 1065 -578 1257 -572
rect 1323 -538 1515 -532
rect 1323 -572 1335 -538
rect 1503 -572 1515 -538
rect 1323 -578 1515 -572
<< properties >>
string FIXED_BBOX -1662 -657 1662 657
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 5.0 l 1.0 m 1 nf 12 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
