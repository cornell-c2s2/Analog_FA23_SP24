magic
tech sky130A
magscale 1 2
timestamp 1712606724
<< pwell >>
rect 3560 -2640 3640 -2600
<< locali >>
rect 1550 -25 1600 25
rect 2125 -25 2150 25
<< viali >>
rect 2640 100 2680 140
rect 3040 100 3080 140
rect 3440 100 3480 140
rect 3840 100 3880 140
rect 4240 100 4280 140
rect 5040 100 5080 140
rect 5440 100 5480 140
rect 5840 100 5880 140
rect 6240 100 6280 140
rect 6640 100 6680 140
rect 1600 -25 1650 25
rect 2075 -25 2125 25
rect 1798 -2740 1952 -2684
rect 3520 -2720 3560 -2680
rect 3840 -2720 3880 -2680
rect 4160 -2720 4200 -2680
rect 4480 -2720 4520 -2680
rect 4800 -2720 4840 -2680
rect 5120 -2720 5160 -2680
rect 5440 -2720 5480 -2680
rect 5760 -2720 5800 -2680
<< metal1 >>
rect 2200 140 6775 150
rect 2200 100 2640 140
rect 2680 100 3040 140
rect 3080 100 3440 140
rect 3480 100 3840 140
rect 3880 100 4240 140
rect 4280 100 5040 140
rect 5080 100 5440 140
rect 5480 100 5840 140
rect 5880 100 6240 140
rect 6280 100 6640 140
rect 6680 100 6775 140
rect 2200 50 2400 100
rect 2628 94 2692 100
rect 3028 94 3092 100
rect 3428 94 3492 100
rect 3828 94 3892 100
rect 4228 94 4292 100
rect 5028 94 5092 100
rect 5428 94 5492 100
rect 5828 94 5892 100
rect 6228 94 6292 100
rect 6628 94 6692 100
rect 1550 25 2400 50
rect 1550 -25 1600 25
rect 1650 -25 2075 25
rect 2125 -25 2400 25
rect 1550 -50 2400 -25
rect 2500 -50 3450 50
rect 3550 -50 4550 50
rect 4800 -50 5750 50
rect 5850 -50 6800 50
rect 2290 -600 2300 -500
rect 2400 -600 4550 -500
rect 1650 -650 1850 -600
rect 1650 -750 1750 -650
rect 1850 -750 2100 -650
rect 4590 -750 4600 -650
rect 4700 -750 6700 -650
rect 1650 -800 1850 -750
rect 1700 -1250 1950 -1150
rect 2650 -1250 6700 -1150
rect 1850 -1300 1950 -1250
rect 1850 -1400 2300 -1300
rect 2400 -1400 2410 -1300
rect 4550 -1400 4750 -1250
rect 1800 -1500 1950 -1400
rect 3450 -1500 5850 -1400
rect 1700 -1950 1750 -1850
rect 1850 -1950 4500 -1850
rect 4590 -2100 4600 -2000
rect 4700 -2100 5700 -2000
rect 2200 -2600 2400 -2550
rect 1700 -2680 2400 -2600
rect 3430 -2640 3450 -2574
rect 3550 -2640 4500 -2574
rect 4720 -2640 5750 -2574
rect 5850 -2640 5856 -2574
rect 3508 -2680 3572 -2674
rect 3828 -2680 3892 -2674
rect 4148 -2680 4212 -2674
rect 4468 -2680 4532 -2674
rect 4788 -2680 4852 -2674
rect 5108 -2680 5172 -2674
rect 5428 -2680 5492 -2674
rect 5748 -2680 5812 -2674
rect 1700 -2684 3520 -2680
rect 1700 -2700 1798 -2684
rect 1786 -2740 1798 -2700
rect 1952 -2700 3520 -2684
rect 1952 -2740 1964 -2700
rect 1786 -2746 1964 -2740
rect 2200 -2720 3520 -2700
rect 3560 -2720 3840 -2680
rect 3880 -2720 4160 -2680
rect 4200 -2720 4480 -2680
rect 4520 -2720 4800 -2680
rect 4840 -2720 5120 -2680
rect 5160 -2720 5440 -2680
rect 5480 -2720 5760 -2680
rect 5800 -2720 5840 -2680
rect 2200 -2760 5840 -2720
<< via1 >>
rect 3450 -50 3550 50
rect 5750 -50 5850 50
rect 2300 -600 2400 -500
rect 1750 -750 1850 -650
rect 4600 -750 4700 -650
rect 2300 -1400 2400 -1300
rect 1750 -1950 1850 -1850
rect 4600 -2100 4700 -2000
rect 3450 -2640 3550 -2574
rect 5750 -2640 5850 -2574
<< metal2 >>
rect 3450 50 3550 60
rect 2300 -500 2400 -490
rect 1750 -650 1850 -640
rect 1750 -760 1850 -750
rect 2300 -1300 2400 -600
rect 3450 -1115 3550 -50
rect 5750 50 5850 60
rect 4600 -650 4700 -640
rect 4600 -760 4700 -750
rect 3390 -1215 3580 -1115
rect 1750 -1850 1850 -1840
rect 1750 -1960 1850 -1950
rect 2300 -2000 2400 -1400
rect 2300 -2110 2400 -2100
rect 3450 -2550 3550 -1215
rect 4600 -2000 4700 -1990
rect 4600 -2110 4700 -2100
rect 3444 -2574 3556 -2550
rect 3444 -2640 3450 -2574
rect 3550 -2640 3556 -2574
rect 3444 -2650 3556 -2640
rect 5750 -2574 5850 -50
rect 5750 -2656 5850 -2640
<< via2 >>
rect 1750 -750 1850 -650
rect 4600 -750 4700 -650
rect 1750 -1950 1850 -1850
rect 2300 -2100 2400 -2000
rect 4600 -2100 4700 -2000
<< metal3 >>
rect 1740 -650 1860 -645
rect 4590 -650 4710 -645
rect 1740 -750 1750 -650
rect 1850 -750 4600 -650
rect 4700 -750 4710 -650
rect 1740 -755 1860 -750
rect 4590 -755 4710 -750
rect 1750 -1845 1850 -755
rect 1740 -1850 1860 -1845
rect 1740 -1950 1750 -1850
rect 1850 -1950 1860 -1850
rect 1740 -1955 1860 -1950
rect 2290 -2000 2410 -1995
rect 4590 -2000 4710 -1995
rect 2290 -2100 2300 -2000
rect 2400 -2100 4600 -2000
rect 4700 -2100 4710 -2000
rect 2290 -2105 2410 -2100
rect 4590 -2105 4710 -2100
use sky130_fd_pr__nfet_01v8_6H2JYD  sky130_fd_pr__nfet_01v8_6H2JYD_0
timestamp 1710000826
transform 1 0 1813 0 1 -2040
box -263 -710 263 710
use sky130_fd_pr__pfet_01v8_UJHYGH  sky130_fd_pr__pfet_01v8_UJHYGH_0
timestamp 1709401415
transform 1 0 1859 0 1 -581
box -359 -719 359 719
use sky130_fd_pr__pfet_01v8_BDZ9JN  XM1
timestamp 1709390584
transform 1 0 3579 0 1 -581
box -1079 -719 1079 719
use sky130_fd_pr__nfet_01v8_KBNS5F  XM2
timestamp 1709392794
transform 1 0 4049 0 1 -2040
box -599 -710 599 710
use sky130_fd_pr__pfet_01v8_BDZ9JN  XM3
timestamp 1709390584
transform 1 0 5729 0 1 -581
box -1079 -719 1079 719
use sky130_fd_pr__nfet_01v8_KBNS5F  XM4
timestamp 1709392794
transform 1 0 5249 0 1 -2040
box -599 -710 599 710
<< labels >>
flabel metal1 2200 -2750 2400 -2550 0 FreeSans 256 0 0 0 VSS
port 4 nsew
flabel metal1 4550 -1350 4750 -1150 0 FreeSans 256 0 0 0 OUT
port 2 nsew
flabel metal1 1650 -800 1850 -600 0 FreeSans 256 0 0 0 VIN
port 3 nsew
flabel metal1 2200 -50 2400 150 0 FreeSans 256 0 0 0 VDD
port 1 nsew
flabel metal1 4450 -50 4550 50 0 FreeSans 256 0 0 0 VREF_P
port 6 nsew
rlabel metal1 4800 -50 4900 50 1 VREF_N
port 7 n
<< end >>
