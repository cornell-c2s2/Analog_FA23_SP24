magic
tech sky130A
magscale 1 2
timestamp 1717181351
<< metal1 >>
rect 402894 693024 402900 693624
rect 403500 693024 403506 693624
rect 446000 689400 446800 689406
rect 446000 688594 446800 688600
rect 539000 688600 539800 688606
rect 539000 687794 539800 687800
rect 386062 683484 406370 684600
rect 408370 683484 408376 684600
rect 402900 678100 403500 678106
rect 386200 677500 402900 678100
rect 402900 677494 403500 677500
rect 82390 676000 82400 676800
rect 83200 676000 83210 676800
rect 131590 676000 131600 676800
rect 132400 676000 132410 676800
rect 154390 676000 154400 676800
rect 155200 676000 155210 676800
rect 456100 675300 457100 675400
rect 456100 675100 456200 675300
rect 456400 675100 456500 675300
rect 456700 675100 456800 675300
rect 457000 675100 457100 675300
rect 456100 675000 457100 675100
rect 456100 674800 456200 675000
rect 456400 674800 456500 675000
rect 456700 674800 456800 675000
rect 457000 674800 457100 675000
rect 53190 670800 53200 671600
rect 54000 670800 54010 671600
rect 58190 670800 58200 671600
rect 59000 670800 59010 671600
rect 82390 670800 82400 671600
rect 83200 670800 83210 671600
rect 131590 670800 131600 671600
rect 132400 670800 132410 671600
rect 154390 670800 154400 671600
rect 155200 670800 155210 671600
rect 456100 665600 457100 674800
rect 560700 668400 561300 668406
rect 560700 667794 561300 667800
rect 456100 665400 456200 665600
rect 456400 665400 456500 665600
rect 456700 665400 456800 665600
rect 457000 665400 457100 665600
rect 456100 665300 457100 665400
rect 456100 665100 456200 665300
rect 456400 665100 456500 665300
rect 456700 665100 456800 665300
rect 457000 665100 457100 665300
rect 456100 665000 457100 665100
rect 391400 650000 395000 651000
rect 391400 649400 392000 650000
rect 392600 649400 393800 650000
rect 394400 649400 395000 650000
rect 391400 649200 395000 649400
rect 391400 648600 393000 649200
rect 393600 648600 395000 649200
rect 391400 648200 395000 648600
rect 391400 647600 392000 648200
rect 392600 647600 393800 648200
rect 394400 647600 395000 648200
rect 391400 647000 395000 647600
rect 44800 625200 46000 625206
rect 44800 623994 46000 624000
rect 44800 620600 46000 620606
rect 44800 619394 46000 619400
rect 44800 616600 46000 616606
rect 44800 615394 46000 615400
rect 44795 612810 46005 612816
rect 44795 611594 46005 611600
rect 10190 601400 10200 602200
rect 11000 601400 11010 602200
rect 15190 601400 15200 602200
rect 16000 601400 16010 602200
rect 19190 601400 19200 602200
rect 20000 601400 20010 602200
rect 24190 601400 24200 602200
rect 25000 601400 25010 602200
rect 28390 601400 28400 602200
rect 29200 601400 29210 602200
rect 33390 601400 33400 602200
rect 34200 601400 34210 602200
rect 37590 601400 37600 602200
rect 38400 601400 38410 602200
rect 42590 601400 42600 602200
rect 43400 601400 43410 602200
<< via1 >>
rect 402900 693024 403500 693624
rect 446000 688600 446800 689400
rect 451400 688562 452200 689362
rect 539000 687800 539800 688600
rect 406370 683484 408370 684600
rect 402900 677500 403500 678100
rect 82400 676000 83200 676800
rect 131600 676000 132400 676800
rect 154400 676000 155200 676800
rect 456200 675100 456400 675300
rect 456500 675100 456700 675300
rect 456800 675100 457000 675300
rect 456200 674800 456400 675000
rect 456500 674800 456700 675000
rect 456800 674800 457000 675000
rect 53200 670800 54000 671600
rect 58200 670800 59000 671600
rect 82400 670800 83200 671600
rect 131600 670800 132400 671600
rect 154400 670800 155200 671600
rect 560700 667800 561300 668400
rect 456200 665400 456400 665600
rect 456500 665400 456700 665600
rect 456800 665400 457000 665600
rect 456200 665100 456400 665300
rect 456500 665100 456700 665300
rect 456800 665100 457000 665300
rect 392000 649400 392600 650000
rect 393800 649400 394400 650000
rect 393000 648600 393600 649200
rect 392000 647600 392600 648200
rect 393800 647600 394400 648200
rect 392800 642200 394400 642400
rect 44800 624000 46000 625200
rect 44800 619400 46000 620600
rect 44800 615400 46000 616600
rect 44795 611600 46005 612810
rect 10200 601400 11000 602200
rect 15200 601400 16000 602200
rect 19200 601400 20000 602200
rect 24200 601400 25000 602200
rect 28400 601400 29200 602200
rect 33400 601400 34200 602200
rect 37600 601400 38400 602200
rect 42600 601400 43400 602200
<< metal2 >>
rect 17600 703600 18800 703609
rect 17600 688395 18800 702400
rect 69600 703600 70800 703609
rect 69600 697795 70800 702400
rect 122200 703600 123400 703609
rect 100200 697800 101400 697809
rect 69596 696605 69605 697795
rect 70795 696605 70804 697795
rect 69600 696600 70800 696605
rect 17600 687205 17605 688395
rect 18795 687205 18800 688395
rect 17600 687200 18800 687205
rect 87991 687200 88000 688400
rect 89200 687200 89209 688400
rect 17605 687196 18795 687200
rect 3200 681200 4400 681209
rect 3200 665795 4400 680000
rect 82400 676800 83200 676810
rect 82400 675990 83200 676000
rect 53200 671600 54000 671610
rect 53200 670790 54000 670800
rect 58200 671600 59000 671610
rect 58200 670790 59000 670800
rect 82400 671600 83200 671610
rect 82400 670790 83200 670800
rect 3196 664605 3205 665795
rect 4395 664605 4404 665795
rect 3200 664600 4400 664605
rect 88000 662600 89200 687200
rect 100200 676995 101400 696600
rect 122200 690595 123400 702400
rect 402900 693624 403500 693630
rect 122200 689405 122205 690595
rect 123395 689405 123400 690595
rect 122200 689400 123400 689405
rect 147800 690600 149000 690609
rect 122205 689396 123395 689400
rect 100200 675805 100205 676995
rect 101395 675805 101400 676995
rect 100200 675800 101400 675805
rect 125600 677000 126800 677009
rect 131600 676800 132400 676810
rect 131600 675990 132400 676000
rect 100205 675796 101395 675800
rect 125600 633600 126800 675800
rect 131600 671600 132400 671610
rect 131600 670790 132400 670800
rect 44805 625200 45995 625204
rect 8400 625195 9600 625200
rect 8396 624005 8405 625195
rect 9595 624005 9604 625195
rect 8400 608200 9600 624005
rect 44794 624000 44800 625200
rect 46000 624000 46006 625200
rect 44805 623996 45995 624000
rect 17600 620600 18800 621200
rect 44805 620600 45995 620604
rect 44794 619400 44800 620600
rect 46000 619400 46006 620600
rect 17600 608200 18800 619400
rect 44805 619396 45995 619400
rect 26805 616600 27995 616604
rect 44805 616600 45995 616604
rect 26800 616595 28000 616600
rect 26800 615405 26805 616595
rect 27995 615405 28000 616595
rect 26800 608200 28000 615405
rect 44794 615400 44800 616600
rect 46000 615400 46006 616600
rect 44805 615396 45995 615400
rect 36000 612810 37200 612814
rect 44800 612810 46000 612814
rect 35995 612805 37205 612810
rect 35995 611605 36000 612805
rect 37200 611605 37205 612805
rect 35995 608200 37205 611605
rect 44789 611600 44795 612810
rect 46005 611600 46011 612810
rect 44800 611596 46000 611600
rect 8400 606800 13400 608200
rect 17600 606800 22400 608200
rect 26800 606800 31600 608200
rect 35995 606800 40800 608200
rect 8400 512400 9600 606800
rect 10200 602200 11000 602210
rect 10200 601390 11000 601400
rect 15200 602200 16000 602210
rect 15200 601390 16000 601400
rect 8400 511191 9600 511200
rect 17600 468995 18800 606800
rect 19200 602200 20000 602210
rect 19200 601390 20000 601400
rect 24200 602200 25000 602210
rect 24200 601390 25000 601400
rect 17600 467805 17605 468995
rect 18795 467805 18800 468995
rect 17600 467800 18800 467805
rect 17605 467796 18795 467800
rect 26800 425800 28000 606800
rect 28400 602200 29200 602210
rect 28400 601390 29200 601400
rect 33400 602200 34200 602210
rect 33400 601390 34200 601400
rect 26800 424591 28000 424600
rect 35995 382405 37205 606800
rect 37600 602200 38400 602210
rect 37600 601390 38400 601400
rect 42600 602200 43400 602210
rect 42600 601390 43400 601400
rect 147800 601195 149000 689400
rect 154400 676800 155200 676810
rect 154400 675990 155200 676000
rect 392650 675550 393350 680900
rect 402900 678100 403500 693024
rect 407800 685490 408400 694800
rect 445994 688600 446000 689400
rect 446800 688600 446806 689400
rect 451400 689362 452200 689400
rect 406370 684600 408400 685490
rect 402894 677500 402900 678100
rect 403500 677500 403506 678100
rect 392650 674841 393350 674850
rect 154400 671600 155200 671610
rect 154400 670790 155200 670800
rect 391400 650000 395000 651000
rect 391400 649400 392000 650000
rect 392600 649400 393800 650000
rect 394400 649400 395000 650000
rect 391400 649200 395000 649400
rect 391400 648600 393000 649200
rect 393600 648600 395000 649200
rect 391400 648200 395000 648600
rect 391400 647600 392000 648200
rect 392600 647600 393800 648200
rect 394400 647600 395000 648200
rect 391400 647000 395000 647600
rect 392600 642400 394600 642600
rect 392600 642200 392800 642400
rect 394400 642200 394600 642400
rect 392600 641800 394600 642200
rect 398600 641200 400000 645800
rect 402900 643571 403500 677500
rect 406370 669195 408370 683484
rect 406366 667205 406375 669195
rect 408365 667205 408374 669195
rect 406370 667200 408370 667205
rect 446000 643800 446800 688600
rect 539005 688600 539795 688604
rect 451400 668600 452200 688562
rect 538994 687800 539000 688600
rect 539800 687800 539806 688600
rect 539005 687796 539795 687800
rect 456200 675300 456400 675310
rect 456200 675090 456400 675100
rect 456500 675300 456700 675310
rect 456500 675090 456700 675100
rect 456800 675300 457000 675310
rect 456800 675090 457000 675100
rect 456200 675000 456400 675010
rect 456200 674790 456400 674800
rect 456500 675000 456700 675010
rect 456500 674790 456700 674800
rect 456800 675000 457000 675010
rect 456800 674790 457000 674800
rect 544000 674300 544600 689800
rect 543991 673700 544000 674300
rect 544600 673700 544609 674300
rect 541105 670500 541695 670504
rect 544000 670500 544600 673700
rect 451400 667791 452200 667800
rect 541100 670495 541700 670500
rect 541100 669905 541105 670495
rect 541695 669905 541700 670495
rect 538600 666390 538800 666610
rect 539000 666390 539200 666610
rect 538600 665990 538800 666210
rect 539000 665990 539200 666210
rect 456200 665600 456400 665610
rect 456200 665390 456400 665400
rect 456500 665600 456700 665610
rect 456500 665390 456700 665400
rect 456800 665600 457000 665610
rect 538600 665590 538800 665810
rect 539000 665590 539200 665810
rect 456800 665390 457000 665400
rect 456200 665300 456400 665310
rect 456200 665090 456400 665100
rect 456500 665300 456700 665310
rect 456500 665090 456700 665100
rect 456800 665300 457000 665310
rect 456800 665090 457000 665100
rect 402896 642981 402905 643571
rect 403495 642981 403504 643571
rect 446000 642991 446800 643000
rect 402900 642976 403500 642981
rect 398600 640200 398800 641200
rect 399800 640200 400000 641200
rect 398600 640000 400000 640200
rect 541100 631900 541700 669905
rect 543991 669900 544000 670500
rect 544600 669900 544609 670500
rect 560694 667800 560700 668400
rect 561300 667800 561306 668400
rect 541091 631300 541100 631900
rect 541700 631300 541709 631900
rect 147800 600005 147805 601195
rect 148995 600005 149000 601195
rect 147800 600000 149000 600005
rect 147805 599996 148995 600000
rect 35995 381205 36000 382405
rect 37200 381205 37205 382405
rect 35995 381195 37205 381205
rect 524 -800 636 480
rect 1706 -800 1818 480
rect 2888 -800 3000 480
rect 4070 -800 4182 480
rect 5252 -800 5364 480
rect 6434 -800 6546 480
rect 7616 -800 7728 480
rect 8798 -800 8910 480
rect 9980 -800 10092 480
rect 11162 -800 11274 480
rect 12344 -800 12456 480
rect 13526 -800 13638 480
rect 14708 -800 14820 480
rect 15890 -800 16002 480
rect 17072 -800 17184 480
rect 18254 -800 18366 480
rect 19436 -800 19548 480
rect 20618 -800 20730 480
rect 21800 -800 21912 480
rect 22982 -800 23094 480
rect 24164 -800 24276 480
rect 25346 -800 25458 480
rect 26528 -800 26640 480
rect 27710 -800 27822 480
rect 28892 -800 29004 480
rect 30074 -800 30186 480
rect 31256 -800 31368 480
rect 32438 -800 32550 480
rect 33620 -800 33732 480
rect 34802 -800 34914 480
rect 35984 -800 36096 480
rect 37166 -800 37278 480
rect 38348 -800 38460 480
rect 39530 -800 39642 480
rect 40712 -800 40824 480
rect 41894 -800 42006 480
rect 43076 -800 43188 480
rect 44258 -800 44370 480
rect 45440 -800 45552 480
rect 46622 -800 46734 480
rect 47804 -800 47916 480
rect 48986 -800 49098 480
rect 50168 -800 50280 480
rect 51350 -800 51462 480
rect 52532 -800 52644 480
rect 53714 -800 53826 480
rect 54896 -800 55008 480
rect 56078 -800 56190 480
rect 57260 -800 57372 480
rect 58442 -800 58554 480
rect 59624 -800 59736 480
rect 60806 -800 60918 480
rect 61988 -800 62100 480
rect 63170 -800 63282 480
rect 64352 -800 64464 480
rect 65534 -800 65646 480
rect 66716 -800 66828 480
rect 67898 -800 68010 480
rect 69080 -800 69192 480
rect 70262 -800 70374 480
rect 71444 -800 71556 480
rect 72626 -800 72738 480
rect 73808 -800 73920 480
rect 74990 -800 75102 480
rect 76172 -800 76284 480
rect 77354 -800 77466 480
rect 78536 -800 78648 480
rect 79718 -800 79830 480
rect 80900 -800 81012 480
rect 82082 -800 82194 480
rect 83264 -800 83376 480
rect 84446 -800 84558 480
rect 85628 -800 85740 480
rect 86810 -800 86922 480
rect 87992 -800 88104 480
rect 89174 -800 89286 480
rect 90356 -800 90468 480
rect 91538 -800 91650 480
rect 92720 -800 92832 480
rect 93902 -800 94014 480
rect 95084 -800 95196 480
rect 96266 -800 96378 480
rect 97448 -800 97560 480
rect 98630 -800 98742 480
rect 99812 -800 99924 480
rect 100994 -800 101106 480
rect 102176 -800 102288 480
rect 103358 -800 103470 480
rect 104540 -800 104652 480
rect 105722 -800 105834 480
rect 106904 -800 107016 480
rect 108086 -800 108198 480
rect 109268 -800 109380 480
rect 110450 -800 110562 480
rect 111632 -800 111744 480
rect 112814 -800 112926 480
rect 113996 -800 114108 480
rect 115178 -800 115290 480
rect 116360 -800 116472 480
rect 117542 -800 117654 480
rect 118724 -800 118836 480
rect 119906 -800 120018 480
rect 121088 -800 121200 480
rect 122270 -800 122382 480
rect 123452 -800 123564 480
rect 124634 -800 124746 480
rect 125816 -800 125928 480
rect 126998 -800 127110 480
rect 128180 -800 128292 480
rect 129362 -800 129474 480
rect 130544 -800 130656 480
rect 131726 -800 131838 480
rect 132908 -800 133020 480
rect 134090 -800 134202 480
rect 135272 -800 135384 480
rect 136454 -800 136566 480
rect 137636 -800 137748 480
rect 138818 -800 138930 480
rect 140000 -800 140112 480
rect 141182 -800 141294 480
rect 142364 -800 142476 480
rect 143546 -800 143658 480
rect 144728 -800 144840 480
rect 145910 -800 146022 480
rect 147092 -800 147204 480
rect 148274 -800 148386 480
rect 149456 -800 149568 480
rect 150638 -800 150750 480
rect 151820 -800 151932 480
rect 153002 -800 153114 480
rect 154184 -800 154296 480
rect 155366 -800 155478 480
rect 156548 -800 156660 480
rect 157730 -800 157842 480
rect 158912 -800 159024 480
rect 160094 -800 160206 480
rect 161276 -800 161388 480
rect 162458 -800 162570 480
rect 163640 -800 163752 480
rect 164822 -800 164934 480
rect 166004 -800 166116 480
rect 167186 -800 167298 480
rect 168368 -800 168480 480
rect 169550 -800 169662 480
rect 170732 -800 170844 480
rect 171914 -800 172026 480
rect 173096 -800 173208 480
rect 174278 -800 174390 480
rect 175460 -800 175572 480
rect 176642 -800 176754 480
rect 177824 -800 177936 480
rect 179006 -800 179118 480
rect 180188 -800 180300 480
rect 181370 -800 181482 480
rect 182552 -800 182664 480
rect 183734 -800 183846 480
rect 184916 -800 185028 480
rect 186098 -800 186210 480
rect 187280 -800 187392 480
rect 188462 -800 188574 480
rect 189644 -800 189756 480
rect 190826 -800 190938 480
rect 192008 -800 192120 480
rect 193190 -800 193302 480
rect 194372 -800 194484 480
rect 195554 -800 195666 480
rect 196736 -800 196848 480
rect 197918 -800 198030 480
rect 199100 -800 199212 480
rect 200282 -800 200394 480
rect 201464 -800 201576 480
rect 202646 -800 202758 480
rect 203828 -800 203940 480
rect 205010 -800 205122 480
rect 206192 -800 206304 480
rect 207374 -800 207486 480
rect 208556 -800 208668 480
rect 209738 -800 209850 480
rect 210920 -800 211032 480
rect 212102 -800 212214 480
rect 213284 -800 213396 480
rect 214466 -800 214578 480
rect 215648 -800 215760 480
rect 216830 -800 216942 480
rect 218012 -800 218124 480
rect 219194 -800 219306 480
rect 220376 -800 220488 480
rect 221558 -800 221670 480
rect 222740 -800 222852 480
rect 223922 -800 224034 480
rect 225104 -800 225216 480
rect 226286 -800 226398 480
rect 227468 -800 227580 480
rect 228650 -800 228762 480
rect 229832 -800 229944 480
rect 231014 -800 231126 480
rect 232196 -800 232308 480
rect 233378 -800 233490 480
rect 234560 -800 234672 480
rect 235742 -800 235854 480
rect 236924 -800 237036 480
rect 238106 -800 238218 480
rect 239288 -800 239400 480
rect 240470 -800 240582 480
rect 241652 -800 241764 480
rect 242834 -800 242946 480
rect 244016 -800 244128 480
rect 245198 -800 245310 480
rect 246380 -800 246492 480
rect 247562 -800 247674 480
rect 248744 -800 248856 480
rect 249926 -800 250038 480
rect 251108 -800 251220 480
rect 252290 -800 252402 480
rect 253472 -800 253584 480
rect 254654 -800 254766 480
rect 255836 -800 255948 480
rect 257018 -800 257130 480
rect 258200 -800 258312 480
rect 259382 -800 259494 480
rect 260564 -800 260676 480
rect 261746 -800 261858 480
rect 262928 -800 263040 480
rect 264110 -800 264222 480
rect 265292 -800 265404 480
rect 266474 -800 266586 480
rect 267656 -800 267768 480
rect 268838 -800 268950 480
rect 270020 -800 270132 480
rect 271202 -800 271314 480
rect 272384 -800 272496 480
rect 273566 -800 273678 480
rect 274748 -800 274860 480
rect 275930 -800 276042 480
rect 277112 -800 277224 480
rect 278294 -800 278406 480
rect 279476 -800 279588 480
rect 280658 -800 280770 480
rect 281840 -800 281952 480
rect 283022 -800 283134 480
rect 284204 -800 284316 480
rect 285386 -800 285498 480
rect 286568 -800 286680 480
rect 287750 -800 287862 480
rect 288932 -800 289044 480
rect 290114 -800 290226 480
rect 291296 -800 291408 480
rect 292478 -800 292590 480
rect 293660 -800 293772 480
rect 294842 -800 294954 480
rect 296024 -800 296136 480
rect 297206 -800 297318 480
rect 298388 -800 298500 480
rect 299570 -800 299682 480
rect 300752 -800 300864 480
rect 301934 -800 302046 480
rect 303116 -800 303228 480
rect 304298 -800 304410 480
rect 305480 -800 305592 480
rect 306662 -800 306774 480
rect 307844 -800 307956 480
rect 309026 -800 309138 480
rect 310208 -800 310320 480
rect 311390 -800 311502 480
rect 312572 -800 312684 480
rect 313754 -800 313866 480
rect 314936 -800 315048 480
rect 316118 -800 316230 480
rect 317300 -800 317412 480
rect 318482 -800 318594 480
rect 319664 -800 319776 480
rect 320846 -800 320958 480
rect 322028 -800 322140 480
rect 323210 -800 323322 480
rect 324392 -800 324504 480
rect 325574 -800 325686 480
rect 326756 -800 326868 480
rect 327938 -800 328050 480
rect 329120 -800 329232 480
rect 330302 -800 330414 480
rect 331484 -800 331596 480
rect 332666 -800 332778 480
rect 333848 -800 333960 480
rect 335030 -800 335142 480
rect 336212 -800 336324 480
rect 337394 -800 337506 480
rect 338576 -800 338688 480
rect 339758 -800 339870 480
rect 340940 -800 341052 480
rect 342122 -800 342234 480
rect 343304 -800 343416 480
rect 344486 -800 344598 480
rect 345668 -800 345780 480
rect 346850 -800 346962 480
rect 348032 -800 348144 480
rect 349214 -800 349326 480
rect 350396 -800 350508 480
rect 351578 -800 351690 480
rect 352760 -800 352872 480
rect 353942 -800 354054 480
rect 355124 -800 355236 480
rect 356306 -800 356418 480
rect 357488 -800 357600 480
rect 358670 -800 358782 480
rect 359852 -800 359964 480
rect 361034 -800 361146 480
rect 362216 -800 362328 480
rect 363398 -800 363510 480
rect 364580 -800 364692 480
rect 365762 -800 365874 480
rect 366944 -800 367056 480
rect 368126 -800 368238 480
rect 369308 -800 369420 480
rect 370490 -800 370602 480
rect 371672 -800 371784 480
rect 372854 -800 372966 480
rect 374036 -800 374148 480
rect 375218 -800 375330 480
rect 376400 -800 376512 480
rect 377582 -800 377694 480
rect 378764 -800 378876 480
rect 379946 -800 380058 480
rect 381128 -800 381240 480
rect 382310 -800 382422 480
rect 383492 -800 383604 480
rect 384674 -800 384786 480
rect 385856 -800 385968 480
rect 387038 -800 387150 480
rect 388220 -800 388332 480
rect 389402 -800 389514 480
rect 390584 -800 390696 480
rect 391766 -800 391878 480
rect 392948 -800 393060 480
rect 394130 -800 394242 480
rect 395312 -800 395424 480
rect 396494 -800 396606 480
rect 397676 -800 397788 480
rect 398858 -800 398970 480
rect 400040 -800 400152 480
rect 401222 -800 401334 480
rect 402404 -800 402516 480
rect 403586 -800 403698 480
rect 404768 -800 404880 480
rect 405950 -800 406062 480
rect 407132 -800 407244 480
rect 408314 -800 408426 480
rect 409496 -800 409608 480
rect 410678 -800 410790 480
rect 411860 -800 411972 480
rect 413042 -800 413154 480
rect 414224 -800 414336 480
rect 415406 -800 415518 480
rect 416588 -800 416700 480
rect 417770 -800 417882 480
rect 418952 -800 419064 480
rect 420134 -800 420246 480
rect 421316 -800 421428 480
rect 422498 -800 422610 480
rect 423680 -800 423792 480
rect 424862 -800 424974 480
rect 426044 -800 426156 480
rect 427226 -800 427338 480
rect 428408 -800 428520 480
rect 429590 -800 429702 480
rect 430772 -800 430884 480
rect 431954 -800 432066 480
rect 433136 -800 433248 480
rect 434318 -800 434430 480
rect 435500 -800 435612 480
rect 436682 -800 436794 480
rect 437864 -800 437976 480
rect 439046 -800 439158 480
rect 440228 -800 440340 480
rect 441410 -800 441522 480
rect 442592 -800 442704 480
rect 443774 -800 443886 480
rect 444956 -800 445068 480
rect 446138 -800 446250 480
rect 447320 -800 447432 480
rect 448502 -800 448614 480
rect 449684 -800 449796 480
rect 450866 -800 450978 480
rect 452048 -800 452160 480
rect 453230 -800 453342 480
rect 454412 -800 454524 480
rect 455594 -800 455706 480
rect 456776 -800 456888 480
rect 457958 -800 458070 480
rect 459140 -800 459252 480
rect 460322 -800 460434 480
rect 461504 -800 461616 480
rect 462686 -800 462798 480
rect 463868 -800 463980 480
rect 465050 -800 465162 480
rect 466232 -800 466344 480
rect 467414 -800 467526 480
rect 468596 -800 468708 480
rect 469778 -800 469890 480
rect 470960 -800 471072 480
rect 472142 -800 472254 480
rect 473324 -800 473436 480
rect 474506 -800 474618 480
rect 475688 -800 475800 480
rect 476870 -800 476982 480
rect 478052 -800 478164 480
rect 479234 -800 479346 480
rect 480416 -800 480528 480
rect 481598 -800 481710 480
rect 482780 -800 482892 480
rect 483962 -800 484074 480
rect 485144 -800 485256 480
rect 486326 -800 486438 480
rect 487508 -800 487620 480
rect 488690 -800 488802 480
rect 489872 -800 489984 480
rect 491054 -800 491166 480
rect 492236 -800 492348 480
rect 493418 -800 493530 480
rect 494600 -800 494712 480
rect 495782 -800 495894 480
rect 496964 -800 497076 480
rect 498146 -800 498258 480
rect 499328 -800 499440 480
rect 500510 -800 500622 480
rect 501692 -800 501804 480
rect 502874 -800 502986 480
rect 504056 -800 504168 480
rect 505238 -800 505350 480
rect 506420 -800 506532 480
rect 507602 -800 507714 480
rect 508784 -800 508896 480
rect 509966 -800 510078 480
rect 511148 -800 511260 480
rect 512330 -800 512442 480
rect 513512 -800 513624 480
rect 514694 -800 514806 480
rect 515876 -800 515988 480
rect 517058 -800 517170 480
rect 518240 -800 518352 480
rect 519422 -800 519534 480
rect 520604 -800 520716 480
rect 521786 -800 521898 480
rect 522968 -800 523080 480
rect 524150 -800 524262 480
rect 525332 -800 525444 480
rect 526514 -800 526626 480
rect 527696 -800 527808 480
rect 528878 -800 528990 480
rect 530060 -800 530172 480
rect 531242 -800 531354 480
rect 532424 -800 532536 480
rect 533606 -800 533718 480
rect 534788 -800 534900 480
rect 535970 -800 536082 480
rect 537152 -800 537264 480
rect 538334 -800 538446 480
rect 539516 -800 539628 480
rect 540698 -800 540810 480
rect 541880 -800 541992 480
rect 543062 -800 543174 480
rect 544244 -800 544356 480
rect 545426 -800 545538 480
rect 546608 -800 546720 480
rect 547790 -800 547902 480
rect 548972 -800 549084 480
rect 550154 -800 550266 480
rect 551336 -800 551448 480
rect 552518 -800 552630 480
rect 553700 -800 553812 480
rect 554882 -800 554994 480
rect 556064 -800 556176 480
rect 557246 -800 557358 480
rect 558428 -800 558540 480
rect 559610 -800 559722 480
rect 560792 -800 560904 480
rect 561974 -800 562086 480
rect 563156 -800 563268 480
rect 564338 -800 564450 480
rect 565520 -800 565632 480
rect 566702 -800 566814 480
rect 567884 -800 567996 480
rect 569066 -800 569178 480
rect 570248 -800 570360 480
rect 571430 -800 571542 480
rect 572612 -800 572724 480
rect 573794 -800 573906 480
rect 574976 -800 575088 480
rect 576158 -800 576270 480
rect 577340 -800 577452 480
rect 578522 -800 578634 480
rect 579704 -800 579816 480
rect 580886 -800 580998 480
rect 582068 -800 582180 480
rect 583250 -800 583362 480
<< via2 >>
rect 17600 702400 18800 703600
rect 69600 702400 70800 703600
rect 122200 702400 123400 703600
rect 69605 696605 70795 697795
rect 100200 696600 101400 697800
rect 17605 687205 18795 688395
rect 88000 687200 89200 688400
rect 3200 680000 4400 681200
rect 82400 676000 83200 676800
rect 53200 670800 54000 671600
rect 58200 670800 59000 671600
rect 82400 670800 83200 671600
rect 3205 664605 4395 665795
rect 122205 689405 123395 690595
rect 147800 689400 149000 690600
rect 100205 675805 101395 676995
rect 125600 675800 126800 677000
rect 131600 676000 132400 676800
rect 131600 670800 132400 671600
rect 8405 624005 9595 625195
rect 44805 624005 45995 625195
rect 17600 619400 18800 620600
rect 44805 619405 45995 620595
rect 26805 615405 27995 616595
rect 44805 615405 45995 616595
rect 36000 611605 37200 612805
rect 44800 611605 46000 612805
rect 10200 601400 11000 602200
rect 15200 601400 16000 602200
rect 8400 511200 9600 512400
rect 19200 601400 20000 602200
rect 24200 601400 25000 602200
rect 17605 467805 18795 468995
rect 28400 601400 29200 602200
rect 33400 601400 34200 602200
rect 26800 424600 28000 425800
rect 37600 601400 38400 602200
rect 42600 601400 43400 602200
rect 154400 676000 155200 676800
rect 392650 674850 393350 675550
rect 154400 670800 155200 671600
rect 392000 649400 392600 650000
rect 393800 649400 394400 650000
rect 393000 648600 393600 649200
rect 392000 647600 392600 648200
rect 393800 647600 394400 648200
rect 392800 642200 394400 642400
rect 406375 667205 408365 669195
rect 539005 687805 539795 688595
rect 456200 675100 456400 675300
rect 456500 675100 456700 675300
rect 456800 675100 457000 675300
rect 456200 674800 456400 675000
rect 456500 674800 456700 675000
rect 456800 674800 457000 675000
rect 544000 673700 544600 674300
rect 451400 667800 452200 668600
rect 541105 669905 541695 670495
rect 456200 665400 456400 665600
rect 456500 665400 456700 665600
rect 456800 665400 457000 665600
rect 456200 665100 456400 665300
rect 456500 665100 456700 665300
rect 456800 665100 457000 665300
rect 402905 642981 403495 643571
rect 446000 643000 446800 643800
rect 398800 640200 399800 641200
rect 544000 669900 544600 670500
rect 560705 667805 561295 668395
rect 541100 631300 541700 631900
rect 147805 600005 148995 601195
rect 36000 381205 37200 382405
<< metal3 >>
rect 16194 703600 21194 704800
rect 16194 702400 17600 703600
rect 18800 702400 21194 703600
rect 16194 702300 21194 702400
rect 68194 703600 73194 704800
rect 68194 702400 69600 703600
rect 70800 702400 73194 703600
rect 68194 702300 73194 702400
rect 120194 703600 125194 704800
rect 120194 702400 122200 703600
rect 123400 702400 125194 703600
rect 120194 702300 125194 702400
rect 165594 702300 170594 704800
rect 170894 702300 173094 704800
rect 173394 702300 175594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 222594 702300 224794 704800
rect 225094 702300 227294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 324294 702300 326494 704800
rect 326794 702300 328994 704800
rect 329294 702300 334294 704800
rect 413394 702400 418394 704800
rect 465394 704000 470394 704800
rect 510594 704000 515394 704800
rect 520594 704000 525394 704800
rect 413394 702300 418400 702400
rect 100195 697800 101405 697805
rect 69600 697795 100200 697800
rect 69600 696605 69605 697795
rect 70795 696605 100200 697795
rect 69600 696600 100200 696605
rect 101400 696600 101405 697800
rect 100195 696595 101405 696600
rect 147795 690600 149005 690605
rect 122200 690595 147800 690600
rect 122200 689405 122205 690595
rect 123395 689405 147800 690595
rect 122200 689400 147800 689405
rect 149000 689400 149005 690600
rect 147795 689395 149005 689400
rect 87995 688400 89205 688405
rect 17600 688395 88000 688400
rect 17600 687205 17605 688395
rect 18795 687205 88000 688395
rect 17600 687200 88000 687205
rect 89200 687200 89205 688400
rect 413400 688200 418400 702300
rect 465000 700000 471000 704000
rect 510594 702800 525394 704000
rect 566594 703000 571594 704800
rect 510594 702340 525400 702800
rect 510600 701200 525400 702340
rect 566594 702300 571600 703000
rect 405200 687400 418400 688200
rect 87995 687195 89205 687200
rect -800 681200 1700 685242
rect 3195 681200 4405 681205
rect -800 680242 3200 681200
rect 0 680000 3200 680242
rect 4400 680000 4405 681200
rect 3195 679995 4405 680000
rect 125595 677000 126805 677005
rect 100200 676995 125600 677000
rect 82390 676800 83210 676805
rect 82390 676000 82400 676800
rect 83200 676000 83210 676800
rect 82390 675995 83210 676000
rect 100200 675805 100205 676995
rect 101395 675805 125600 676995
rect 100200 675800 125600 675805
rect 126800 675800 126805 677000
rect 131590 676800 132410 676805
rect 131590 676000 131600 676800
rect 132400 676000 132410 676800
rect 131590 675995 132410 676000
rect 154390 676800 155210 676805
rect 154390 676000 154400 676800
rect 155200 676000 155210 676800
rect 154390 675995 155210 676000
rect 125595 675795 126805 675800
rect 392645 675555 393355 675561
rect 392645 674850 392650 674855
rect 393350 674850 393355 674855
rect 392645 674845 393355 674850
rect 413400 673400 418400 687400
rect 456100 698900 471000 700000
rect 456100 683400 457100 698900
rect 448000 682600 457100 683400
rect 456100 675300 457100 682600
rect 520600 688600 525400 701200
rect 566600 695800 571600 702300
rect 545900 694500 571600 695800
rect 520600 688595 539800 688600
rect 520600 687805 539005 688595
rect 539795 687805 539800 688595
rect 520600 687800 539800 687805
rect 456100 675100 456200 675300
rect 456400 675100 456500 675300
rect 456700 675100 456800 675300
rect 457000 675100 457100 675300
rect 456100 675000 457100 675100
rect 456100 674800 456200 675000
rect 456400 674800 456500 675000
rect 456700 674800 456800 675000
rect 457000 674800 457100 675000
rect 463700 676300 465100 676400
rect 463700 676000 463800 676300
rect 464100 676000 464300 676300
rect 464600 676000 465100 676300
rect 463700 675800 465100 676000
rect 463700 675500 463800 675800
rect 464100 675500 464300 675800
rect 464600 675500 465100 675800
rect 463700 675300 465100 675500
rect 463700 675000 463800 675300
rect 464100 675000 464300 675300
rect 464600 675000 465100 675300
rect 463700 674900 465100 675000
rect 456100 674700 457100 674800
rect 520600 674200 525400 687800
rect 545900 683000 547900 694500
rect 541000 682400 547900 683000
rect 545900 678500 547900 682400
rect 545900 678200 546000 678500
rect 546300 678200 546500 678500
rect 546800 678200 547000 678500
rect 547300 678200 547500 678500
rect 547800 678200 547900 678500
rect 545900 678000 547900 678200
rect 545900 677700 546000 678000
rect 546300 677700 546500 678000
rect 546800 677700 547000 678000
rect 547300 677700 547500 678000
rect 547800 677700 547900 678000
rect 545900 677500 547900 677700
rect 545900 677200 546000 677500
rect 546300 677200 546500 677500
rect 546800 677200 547000 677500
rect 547300 677200 547500 677500
rect 547800 677200 547900 677500
rect 545900 677100 547900 677200
rect 575800 682984 582600 683000
rect 575800 678000 584800 682984
rect 520600 673600 520800 674200
rect 521400 673600 521800 674200
rect 522400 673600 522800 674200
rect 523400 673600 523800 674200
rect 524400 673600 525400 674200
rect 543995 674300 544605 674305
rect 543995 673700 544000 674300
rect 544600 673700 561100 674300
rect 543995 673695 544605 673700
rect 53190 671600 54010 671605
rect 53190 670800 53200 671600
rect 54000 670800 54010 671600
rect 53190 670795 54010 670800
rect 58190 671600 59010 671605
rect 58190 670800 58200 671600
rect 59000 670800 59010 671600
rect 58190 670795 59010 670800
rect 82390 671600 83210 671605
rect 82390 670800 82400 671600
rect 83200 670800 83210 671600
rect 82390 670795 83210 670800
rect 131590 671600 132410 671605
rect 131590 670800 131600 671600
rect 132400 670800 132410 671600
rect 131590 670795 132410 670800
rect 154390 671600 155210 671605
rect 154390 670800 154400 671600
rect 155200 670800 155210 671600
rect 154390 670795 155210 670800
rect 413400 670400 450400 673400
rect 520600 673200 525400 673600
rect 520600 672600 520800 673200
rect 521400 672600 521800 673200
rect 522400 672600 522800 673200
rect 523400 672600 523800 673200
rect 524400 672600 525400 673200
rect 560500 673100 561100 673700
rect 520600 672200 525400 672600
rect 520600 671600 520800 672200
rect 521400 671600 521800 672200
rect 522400 671600 522800 672200
rect 523400 671600 523800 672200
rect 524400 671600 525400 672200
rect 520600 671200 525400 671600
rect 520600 670600 520800 671200
rect 521400 670600 521800 671200
rect 522400 670600 522800 671200
rect 523400 670600 523800 671200
rect 524400 670600 525400 671200
rect 520600 670400 525400 670600
rect 543995 670500 544605 670505
rect 541100 670495 544000 670500
rect 541100 669905 541105 670495
rect 541695 669905 544000 670495
rect 541100 669900 544000 669905
rect 544600 669900 544605 670500
rect 543995 669895 544605 669900
rect 406370 669199 408370 669200
rect 406365 667201 406371 669199
rect 408369 667201 408375 669199
rect 451395 668600 451405 668605
rect 451395 667800 451400 668600
rect 451395 667795 451405 667800
rect 452205 667795 452211 668605
rect 535694 667800 535700 668400
rect 536300 668395 561300 668400
rect 536300 667805 560705 668395
rect 561295 667805 561300 668395
rect 536300 667800 561300 667805
rect 406370 667200 408370 667201
rect 565900 666800 567300 670700
rect 575800 666800 579000 678000
rect 582300 677984 584800 678000
rect 3200 665795 81600 665800
rect 3200 664605 3205 665795
rect 4395 664605 81600 665795
rect 3200 664600 81600 664605
rect 456100 665600 457100 665700
rect 456100 665400 456200 665600
rect 456400 665400 456500 665600
rect 456700 665400 456800 665600
rect 457000 665400 457100 665600
rect 456100 665300 457100 665400
rect 456100 665100 456200 665300
rect 456400 665100 456500 665300
rect 456700 665100 456800 665300
rect 457000 665100 457100 665300
rect 456100 654000 457100 665100
rect 543600 665400 579000 666800
rect 391400 650000 395000 651000
rect 543600 650300 544700 665400
rect 391400 649400 392000 650000
rect 392600 649400 393800 650000
rect 394400 649400 395000 650000
rect 391400 649200 395000 649400
rect -800 648600 1660 648642
rect 391400 648600 393000 649200
rect 393600 648600 395000 649200
rect -800 644000 4700 648600
rect 391400 648200 395000 648600
rect 391400 647600 392000 648200
rect 392600 647600 393800 648200
rect 394400 647600 395000 648200
rect 391400 647000 395000 647600
rect -800 643842 2400 644000
rect 1600 643700 2400 643842
rect 1700 643400 2400 643700
rect 3000 643400 3600 644000
rect 4200 643400 4700 644000
rect 577800 644584 583100 644600
rect 445995 643805 446805 643811
rect 402900 643575 403500 643576
rect 1700 642800 4700 643400
rect 402895 642977 402901 643575
rect 403499 642977 403505 643575
rect 445995 643000 446000 643005
rect 446800 643000 446805 643005
rect 445995 642995 446805 643000
rect 402900 642976 403500 642977
rect 1700 642200 2400 642800
rect 3000 642200 3600 642800
rect 4200 642200 4700 642800
rect 1700 641600 4700 642200
rect 392600 642400 394600 642600
rect 392600 642200 392800 642400
rect 394400 642200 394600 642400
rect 401200 642400 402200 642600
rect 401200 642200 401400 642400
rect 392600 642000 401400 642200
rect 402000 642000 402200 642400
rect 392600 641800 402200 642000
rect 1700 641000 2400 641600
rect 3000 641000 3600 641600
rect 4200 641000 4700 641600
rect 1700 640400 4700 641000
rect 1700 639800 2400 640400
rect 3000 639800 3600 640400
rect 4200 639800 4700 640400
rect 398600 641200 400000 641400
rect 398600 640200 398800 641200
rect 399800 640200 400000 641200
rect 398600 640000 400000 640200
rect 1700 638800 4700 639800
rect 1600 638642 4700 638800
rect -800 633900 4700 638642
rect 577800 639784 584800 644584
rect 577800 634584 584000 639784
rect -800 633842 1660 633900
rect 577800 633500 584800 634584
rect 577800 633200 577900 633500
rect 578200 633200 578400 633500
rect 578700 633200 584800 633500
rect 577800 633000 584800 633200
rect 577800 632700 577900 633000
rect 578200 632700 578400 633000
rect 578700 632700 584800 633000
rect 577800 632500 584800 632700
rect 577800 632200 577900 632500
rect 578200 632200 578400 632500
rect 578700 632200 584800 632500
rect 577800 632000 584800 632200
rect 541089 631295 541095 631905
rect 541695 631900 541705 631905
rect 541700 631300 541705 631900
rect 541695 631295 541705 631300
rect 577800 631700 577900 632000
rect 578200 631700 578400 632000
rect 578700 631700 584800 632000
rect 577800 631500 584800 631700
rect 577800 631200 577900 631500
rect 578200 631200 578400 631500
rect 578700 631200 584800 631500
rect 577800 631000 584800 631200
rect 577800 630700 577900 631000
rect 578200 630700 578400 631000
rect 578700 630700 584800 631000
rect 577800 630500 584800 630700
rect 577800 630200 577900 630500
rect 578200 630200 578400 630500
rect 578700 630200 584800 630500
rect 577800 629800 584800 630200
rect 582340 629784 584800 629800
rect 8400 625195 46000 625200
rect 8400 624005 8405 625195
rect 9595 624005 44805 625195
rect 45995 624005 46000 625195
rect 8400 624000 46000 624005
rect 17595 620600 18805 620605
rect 17595 619400 17600 620600
rect 18800 620595 46000 620600
rect 18800 619405 44805 620595
rect 45995 619405 46000 620595
rect 18800 619400 46000 619405
rect 17595 619395 18805 619400
rect 26800 616595 46000 616600
rect 26800 615405 26805 616595
rect 27995 615405 44805 616595
rect 45995 615405 46000 616595
rect 26800 615400 46000 615405
rect 35995 612805 46005 612810
rect 35995 611605 36000 612805
rect 37200 611605 44800 612805
rect 46000 611605 46005 612805
rect 35995 611600 46005 611605
rect 10190 602200 11010 602205
rect 10190 601400 10200 602200
rect 11000 601400 11010 602200
rect 10190 601395 11010 601400
rect 15190 602200 16010 602205
rect 15190 601400 15200 602200
rect 16000 601400 16010 602200
rect 15190 601395 16010 601400
rect 19190 602200 20010 602205
rect 19190 601400 19200 602200
rect 20000 601400 20010 602200
rect 19190 601395 20010 601400
rect 24190 602200 25010 602205
rect 24190 601400 24200 602200
rect 25000 601400 25010 602200
rect 24190 601395 25010 601400
rect 28390 602200 29210 602205
rect 28390 601400 28400 602200
rect 29200 601400 29210 602200
rect 28390 601395 29210 601400
rect 33390 602200 34210 602205
rect 33390 601400 33400 602200
rect 34200 601400 34210 602200
rect 33390 601395 34210 601400
rect 37590 602200 38410 602205
rect 37590 601400 37600 602200
rect 38400 601400 38410 602200
rect 37590 601395 38410 601400
rect 42590 602200 43410 602205
rect 42590 601400 42600 602200
rect 43400 601400 43410 602200
rect 42590 601395 43410 601400
rect 123600 601195 149000 601200
rect 123600 600005 147805 601195
rect 148995 600005 149000 601195
rect 123600 600000 149000 600005
rect 583520 589472 584800 589584
rect 583520 588290 584800 588402
rect 583520 587108 584800 587220
rect 583520 585926 584800 586038
rect 583520 584744 584800 584856
rect 583520 583562 584800 583674
rect -800 559442 1660 564242
rect -800 549442 1660 554242
rect 582340 550562 584800 555362
rect 582340 540562 584800 545362
rect 8395 512400 9605 512405
rect 0 511642 8400 512400
rect -800 511530 8400 511642
rect 0 511200 8400 511530
rect 9600 511200 9605 512400
rect 8395 511195 9605 511200
rect -800 510348 480 510460
rect -800 509166 480 509278
rect -800 507984 480 508096
rect -800 506802 480 506914
rect -800 505620 480 505732
rect 583520 500050 584800 500162
rect 583520 498868 584800 498980
rect 583520 497686 584800 497798
rect 583520 496504 584800 496616
rect 583520 495322 584800 495434
rect 583520 494140 584800 494252
rect 0 468995 18800 469000
rect 0 468420 17605 468995
rect -800 468308 17605 468420
rect 0 467805 17605 468308
rect 18795 467805 18800 468995
rect 0 467800 18800 467805
rect -800 467126 480 467238
rect -800 465944 480 466056
rect -800 464762 480 464874
rect -800 463580 480 463692
rect -800 462398 480 462510
rect 583520 455628 584800 455740
rect 583520 454446 584800 454558
rect 583520 453264 584800 453376
rect 583520 452082 584800 452194
rect 583520 450900 584800 451012
rect 583520 449718 584800 449830
rect 26795 425800 28005 425805
rect 0 425198 26800 425800
rect -800 425086 26800 425198
rect 0 424600 26800 425086
rect 28000 424600 28005 425800
rect 26795 424595 28005 424600
rect -800 423904 480 424016
rect -800 422722 480 422834
rect -800 421540 480 421652
rect -800 420358 480 420470
rect -800 419176 480 419288
rect 583520 411206 584800 411318
rect 583520 410024 584800 410136
rect 583520 408842 584800 408954
rect 583520 407660 584800 407772
rect 583520 406478 584800 406590
rect 583520 405296 584800 405408
rect 0 382405 37205 382410
rect 0 381976 36000 382405
rect -800 381864 36000 381976
rect 0 381205 36000 381864
rect 37200 381205 37205 382405
rect 0 381200 37205 381205
rect -800 380682 480 380794
rect -800 379500 480 379612
rect -800 378318 480 378430
rect -800 377136 480 377248
rect -800 375954 480 376066
rect 583520 364784 584800 364896
rect 583520 363602 584800 363714
rect 583520 362420 584800 362532
rect 583520 361238 584800 361350
rect 583520 360056 584800 360168
rect 583520 358874 584800 358986
rect -800 338642 480 338754
rect -800 337460 480 337572
rect -800 336278 480 336390
rect -800 335096 480 335208
rect -800 333914 480 334026
rect -800 332732 480 332844
rect 583520 319562 584800 319674
rect 583520 318380 584800 318492
rect 583520 317198 584800 317310
rect 583520 316016 584800 316128
rect 583520 314834 584800 314946
rect 583520 313652 584800 313764
rect -800 295420 480 295532
rect -800 294238 480 294350
rect -800 293056 480 293168
rect -800 291874 480 291986
rect -800 290692 480 290804
rect -800 289510 480 289622
rect 583520 275140 584800 275252
rect 583520 273958 584800 274070
rect 583520 272776 584800 272888
rect 583520 271594 584800 271706
rect 583520 270412 584800 270524
rect 583520 269230 584800 269342
rect -800 252398 480 252510
rect -800 251216 480 251328
rect -800 250034 480 250146
rect -800 248852 480 248964
rect -800 247670 480 247782
rect -800 246488 480 246600
rect 582340 235230 584800 240030
rect 582340 225230 584800 230030
rect -800 214888 1660 219688
rect -800 204888 1660 209688
rect 582340 191430 584800 196230
rect 582340 181430 584800 186230
rect -800 172888 1660 177688
rect -800 162888 1660 167688
rect 582340 146830 584800 151630
rect 582340 136830 584800 141630
rect -800 124776 480 124888
rect -800 123594 480 123706
rect -800 122412 480 122524
rect -800 121230 480 121342
rect -800 120048 480 120160
rect -800 118866 480 118978
rect 583520 95118 584800 95230
rect 583520 93936 584800 94048
rect 583520 92754 584800 92866
rect 583520 91572 584800 91684
rect -800 81554 480 81666
rect -800 80372 480 80484
rect -800 79190 480 79302
rect -800 78008 480 78120
rect -800 76826 480 76938
rect -800 75644 480 75756
rect 583520 50460 584800 50572
rect 583520 49278 584800 49390
rect 583520 48096 584800 48208
rect 583520 46914 584800 47026
rect -800 38332 480 38444
rect -800 37150 480 37262
rect -800 35968 480 36080
rect -800 34786 480 34898
rect -800 33604 480 33716
rect -800 32422 480 32534
rect 583520 24002 584800 24114
rect 583520 22820 584800 22932
rect 583520 21638 584800 21750
rect 583520 20456 584800 20568
rect 583520 19274 584800 19386
rect 583520 18092 584800 18204
rect -800 16910 480 17022
rect 583520 16910 584800 17022
rect -800 15728 480 15840
rect 583520 15728 584800 15840
rect -800 14546 480 14658
rect 583520 14546 584800 14658
rect -800 13364 480 13476
rect 583520 13364 584800 13476
rect -800 12182 480 12294
rect 583520 12182 584800 12294
rect -800 11000 480 11112
rect 583520 11000 584800 11112
rect -800 9818 480 9930
rect 583520 9818 584800 9930
rect -800 8636 480 8748
rect 583520 8636 584800 8748
rect -800 7454 480 7566
rect 583520 7454 584800 7566
rect -800 6272 480 6384
rect 583520 6272 584800 6384
rect -800 5090 480 5202
rect 583520 5090 584800 5202
rect -800 3908 480 4020
rect 583520 3908 584800 4020
rect -800 2726 480 2838
rect 583520 2726 584800 2838
rect -800 1544 480 1656
rect 583520 1544 584800 1656
<< via3 >>
rect 82400 676000 83200 676800
rect 131600 676000 132400 676800
rect 154400 676000 155200 676800
rect 392645 675550 393355 675555
rect 392645 674855 392650 675550
rect 392650 674855 393350 675550
rect 393350 674855 393355 675550
rect 463800 676000 464100 676300
rect 464300 676000 464600 676300
rect 463800 675500 464100 675800
rect 464300 675500 464600 675800
rect 463800 675000 464100 675300
rect 464300 675000 464600 675300
rect 546000 678200 546300 678500
rect 546500 678200 546800 678500
rect 547000 678200 547300 678500
rect 547500 678200 547800 678500
rect 546000 677700 546300 678000
rect 546500 677700 546800 678000
rect 547000 677700 547300 678000
rect 547500 677700 547800 678000
rect 546000 677200 546300 677500
rect 546500 677200 546800 677500
rect 547000 677200 547300 677500
rect 547500 677200 547800 677500
rect 520800 673600 521400 674200
rect 521800 673600 522400 674200
rect 522800 673600 523400 674200
rect 523800 673600 524400 674200
rect 53200 670800 54000 671600
rect 58200 670800 59000 671600
rect 82400 670800 83200 671600
rect 131600 670800 132400 671600
rect 154400 670800 155200 671600
rect 520800 672600 521400 673200
rect 521800 672600 522400 673200
rect 522800 672600 523400 673200
rect 523800 672600 524400 673200
rect 520800 671600 521400 672200
rect 521800 671600 522400 672200
rect 522800 671600 523400 672200
rect 523800 671600 524400 672200
rect 520800 670600 521400 671200
rect 521800 670600 522400 671200
rect 522800 670600 523400 671200
rect 523800 670600 524400 671200
rect 406371 669195 408369 669199
rect 406371 667205 406375 669195
rect 406375 667205 408365 669195
rect 408365 667205 408369 669195
rect 406371 667201 408369 667205
rect 451405 668600 452205 668605
rect 451405 667800 452200 668600
rect 452200 667800 452205 668600
rect 451405 667795 452205 667800
rect 535700 667800 536300 668400
rect 392000 649400 392600 650000
rect 393800 649400 394400 650000
rect 393000 648600 393600 649200
rect 392000 647600 392600 648200
rect 393800 647600 394400 648200
rect 2400 643400 3000 644000
rect 3600 643400 4200 644000
rect 445995 643800 446805 643805
rect 402901 643571 403499 643575
rect 402901 642981 402905 643571
rect 402905 642981 403495 643571
rect 403495 642981 403499 643571
rect 402901 642977 403499 642981
rect 445995 643005 446000 643800
rect 446000 643005 446800 643800
rect 446800 643005 446805 643800
rect 2400 642200 3000 642800
rect 3600 642200 4200 642800
rect 401400 642000 402000 642400
rect 2400 641000 3000 641600
rect 3600 641000 4200 641600
rect 2400 639800 3000 640400
rect 3600 639800 4200 640400
rect 398800 640200 399800 641200
rect 577900 633200 578200 633500
rect 578400 633200 578700 633500
rect 577900 632700 578200 633000
rect 578400 632700 578700 633000
rect 577900 632200 578200 632500
rect 578400 632200 578700 632500
rect 541095 631900 541695 631905
rect 541095 631300 541100 631900
rect 541100 631300 541695 631900
rect 541095 631295 541695 631300
rect 577900 631700 578200 632000
rect 578400 631700 578700 632000
rect 577900 631200 578200 631500
rect 578400 631200 578700 631500
rect 577900 630700 578200 631000
rect 578400 630700 578700 631000
rect 577900 630200 578200 630500
rect 578400 630200 578700 630500
rect 10200 601400 11000 602200
rect 15200 601400 16000 602200
rect 19200 601400 20000 602200
rect 24200 601400 25000 602200
rect 28400 601400 29200 602200
rect 33400 601400 34200 602200
rect 37600 601400 38400 602200
rect 42600 601400 43400 602200
<< metal4 >>
rect 165594 702300 170594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 329294 702300 334294 704800
rect 545999 678500 546301 678501
rect 545999 678200 546000 678500
rect 546300 678200 546301 678500
rect 545999 678199 546301 678200
rect 546499 678500 546801 678501
rect 546499 678200 546500 678500
rect 546800 678200 546801 678500
rect 546499 678199 546801 678200
rect 546999 678500 547301 678501
rect 546999 678200 547000 678500
rect 547300 678200 547301 678500
rect 546999 678199 547301 678200
rect 547499 678500 547801 678501
rect 547499 678200 547500 678500
rect 547800 678200 547801 678500
rect 547499 678199 547801 678200
rect 545999 678000 546301 678001
rect 545999 677700 546000 678000
rect 546300 677700 546301 678000
rect 545999 677699 546301 677700
rect 546499 678000 546801 678001
rect 546499 677700 546500 678000
rect 546800 677700 546801 678000
rect 546499 677699 546801 677700
rect 546999 678000 547301 678001
rect 546999 677700 547000 678000
rect 547300 677700 547301 678000
rect 546999 677699 547301 677700
rect 547499 678000 547801 678001
rect 547499 677700 547500 678000
rect 547800 677700 547801 678000
rect 547499 677699 547801 677700
rect 545999 677500 546301 677501
rect 545999 677200 546000 677500
rect 546300 677200 546301 677500
rect 545999 677199 546301 677200
rect 546499 677500 546801 677501
rect 546499 677200 546500 677500
rect 546800 677200 546801 677500
rect 546499 677199 546801 677200
rect 546999 677500 547301 677501
rect 546999 677200 547000 677500
rect 547300 677200 547301 677500
rect 546999 677199 547301 677200
rect 547499 677500 547801 677501
rect 547499 677200 547500 677500
rect 547800 677200 547801 677500
rect 547499 677199 547801 677200
rect 82399 676800 83201 676801
rect 82399 676000 82400 676800
rect 83200 676000 83201 676800
rect 82399 675999 83201 676000
rect 131599 676800 132401 676801
rect 131599 676000 131600 676800
rect 132400 676000 132401 676800
rect 131599 675999 132401 676000
rect 154399 676800 155201 676801
rect 154399 676000 154400 676800
rect 155200 676000 155201 676800
rect 154399 675999 155201 676000
rect 329300 676400 465100 676500
rect 329300 676100 329500 676400
rect 329800 676100 330000 676400
rect 330300 676100 330500 676400
rect 330800 676100 331000 676400
rect 331300 676100 331500 676400
rect 331800 676100 332000 676400
rect 332300 676100 332500 676400
rect 332800 676100 333000 676400
rect 333300 676100 333500 676400
rect 333800 676300 465100 676400
rect 333800 676100 463800 676300
rect 329300 676000 463800 676100
rect 464100 676000 464300 676300
rect 464600 676000 465100 676300
rect 329300 675900 465100 676000
rect 329300 675600 329500 675900
rect 329800 675600 330000 675900
rect 330300 675600 330500 675900
rect 330800 675600 331000 675900
rect 331300 675600 331500 675900
rect 331800 675600 332000 675900
rect 332300 675600 332500 675900
rect 332800 675600 333000 675900
rect 333300 675600 333500 675900
rect 333800 675800 465100 675900
rect 333800 675600 463800 675800
rect 329300 675555 463800 675600
rect 329300 675400 392645 675555
rect 329300 675100 329500 675400
rect 329800 675100 330000 675400
rect 330300 675100 330500 675400
rect 330800 675100 331000 675400
rect 331300 675100 331500 675400
rect 331800 675100 332000 675400
rect 332300 675100 332500 675400
rect 332800 675100 333000 675400
rect 333300 675100 333500 675400
rect 333800 675100 392645 675400
rect 329300 674900 392645 675100
rect 392644 674855 392645 674900
rect 393355 675500 463800 675555
rect 464100 675500 464300 675800
rect 464600 675500 465100 675800
rect 393355 675300 465100 675500
rect 393355 675000 463800 675300
rect 464100 675000 464300 675300
rect 464600 675000 465100 675300
rect 393355 674900 465100 675000
rect 393355 674855 393356 674900
rect 392644 674854 393356 674855
rect 520799 674200 521401 674201
rect 520799 673600 520800 674200
rect 521400 673600 521401 674200
rect 520799 673599 521401 673600
rect 521799 674200 522401 674201
rect 521799 673600 521800 674200
rect 522400 673600 522401 674200
rect 521799 673599 522401 673600
rect 522799 674200 523401 674201
rect 522799 673600 522800 674200
rect 523400 673600 523401 674200
rect 522799 673599 523401 673600
rect 523799 674200 524401 674201
rect 523799 673600 523800 674200
rect 524400 673600 524401 674200
rect 523799 673599 524401 673600
rect 520799 673200 521401 673201
rect 520799 672600 520800 673200
rect 521400 672600 521401 673200
rect 520799 672599 521401 672600
rect 521799 673200 522401 673201
rect 521799 672600 521800 673200
rect 522400 672600 522401 673200
rect 521799 672599 522401 672600
rect 522799 673200 523401 673201
rect 522799 672600 522800 673200
rect 523400 672600 523401 673200
rect 522799 672599 523401 672600
rect 523799 673200 524401 673201
rect 523799 672600 523800 673200
rect 524400 672600 524401 673200
rect 523799 672599 524401 672600
rect 520799 672200 521401 672201
rect 53199 671600 54001 671601
rect 53199 670800 53200 671600
rect 54000 670800 54001 671600
rect 53199 670799 54001 670800
rect 58199 671600 59001 671601
rect 82399 671600 83201 671601
rect 131599 671600 132401 671601
rect 154399 671600 155201 671601
rect 58199 670800 58200 671600
rect 59000 670800 82400 671600
rect 83200 670800 131600 671600
rect 132400 670800 154400 671600
rect 155200 670800 155201 671600
rect 520799 671600 520800 672200
rect 521400 671600 521401 672200
rect 520799 671599 521401 671600
rect 521799 672200 522401 672201
rect 521799 671600 521800 672200
rect 522400 671600 522401 672200
rect 521799 671599 522401 671600
rect 522799 672200 523401 672201
rect 522799 671600 522800 672200
rect 523400 671600 523401 672200
rect 522799 671599 523401 671600
rect 523799 672200 524401 672201
rect 523799 671600 523800 672200
rect 524400 671600 524401 672200
rect 523799 671599 524401 671600
rect 58199 670799 59001 670800
rect 82399 670799 83201 670800
rect 82400 669400 83200 670799
rect 99400 668200 102800 670800
rect 131599 670799 132401 670800
rect 154399 670799 155201 670800
rect 520799 671200 521401 671201
rect 520799 670600 520800 671200
rect 521400 670600 521401 671200
rect 520799 670599 521401 670600
rect 521799 671200 522401 671201
rect 521799 670600 521800 671200
rect 522400 670600 522401 671200
rect 521799 670599 522401 670600
rect 522799 671200 523401 671201
rect 522799 670600 522800 671200
rect 523400 670600 523401 671200
rect 522799 670599 523401 670600
rect 523799 671200 524401 671201
rect 523799 670600 523800 671200
rect 524400 670600 524401 671200
rect 523799 670599 524401 670600
rect 406370 669199 408370 669200
rect 406370 667201 406371 669199
rect 408369 667201 408370 669199
rect 451404 667795 451405 667806
rect 452205 667795 452206 667806
rect 535699 668400 536301 668401
rect 535699 667800 535700 668400
rect 536300 667800 536301 668400
rect 535699 667799 536301 667800
rect 451404 667794 452206 667795
rect 406370 667200 408370 667201
rect 391400 650000 395000 651000
rect 391400 649400 392000 650000
rect 392600 649400 393800 650000
rect 394400 649400 395000 650000
rect 391400 649200 395000 649400
rect 391400 648600 393000 649200
rect 393600 648600 395000 649200
rect 391400 648200 395000 648600
rect 391400 647600 392000 648200
rect 392600 647600 393800 648200
rect 394400 647600 395000 648200
rect 447000 650000 456000 651000
rect 447000 649000 448000 650000
rect 449000 649000 456000 650000
rect 447000 648000 456000 649000
rect 391400 647000 395000 647600
rect 2399 644000 3001 644001
rect 2399 643400 2400 644000
rect 3000 643400 3001 644000
rect 2399 643399 3001 643400
rect 3599 644000 4201 644001
rect 3599 643400 3600 644000
rect 4200 643400 4201 644000
rect 3599 643399 4201 643400
rect 401200 643600 402200 643800
rect 401200 643000 401400 643600
rect 402000 643000 402200 643600
rect 2399 642800 3001 642801
rect 2399 642200 2400 642800
rect 3000 642200 3001 642800
rect 2399 642199 3001 642200
rect 3599 642800 4201 642801
rect 3599 642200 3600 642800
rect 4200 642200 4201 642800
rect 3599 642199 4201 642200
rect 401200 642400 402200 643000
rect 445994 643005 445995 643006
rect 446805 643005 446806 643006
rect 445994 643004 446806 643005
rect 457600 643400 459800 643800
rect 402900 642977 402901 643000
rect 403499 642977 403500 643000
rect 402900 642976 403500 642977
rect 401200 642000 401400 642400
rect 402000 642000 402200 642400
rect 457600 642400 458000 643400
rect 459400 642400 459800 643400
rect 457600 642000 459800 642400
rect 401200 641800 402200 642000
rect 2399 641600 3001 641601
rect 2399 641000 2400 641600
rect 3000 641000 3001 641600
rect 2399 640999 3001 641000
rect 3599 641600 4201 641601
rect 3599 641000 3600 641600
rect 4200 641000 4201 641600
rect 3599 640999 4201 641000
rect 323600 641400 332600 641500
rect 411700 641400 424300 641500
rect 323600 641100 323700 641400
rect 324000 641100 324200 641400
rect 324500 641100 324700 641400
rect 325000 641100 330600 641400
rect 330900 641100 331100 641400
rect 331400 641100 332600 641400
rect 323600 640900 332600 641100
rect 323600 640600 323700 640900
rect 324000 640600 324200 640900
rect 324500 640600 324700 640900
rect 325000 640600 330600 640900
rect 330900 640600 331100 640900
rect 331400 640600 332600 640900
rect 2399 640400 3001 640401
rect 2399 639800 2400 640400
rect 3000 639800 3001 640400
rect 2399 639799 3001 639800
rect 3599 640400 4201 640401
rect 3599 639800 3600 640400
rect 4200 639800 4201 640400
rect 323600 640400 332600 640600
rect 323600 640100 323700 640400
rect 324000 640100 324200 640400
rect 324500 640100 324700 640400
rect 325000 640100 330600 640400
rect 330900 640100 331100 640400
rect 331400 640100 332600 640400
rect 323600 640000 332600 640100
rect 398600 641200 400000 641400
rect 398600 640200 398800 641200
rect 399800 640200 400000 641200
rect 398600 640000 400000 640200
rect 411700 641100 411800 641400
rect 412100 641100 412300 641400
rect 412600 641100 422900 641400
rect 423200 641100 423400 641400
rect 423700 641100 424300 641400
rect 411700 640900 424300 641100
rect 411700 640600 411800 640900
rect 412100 640600 412300 640900
rect 412600 640600 422900 640900
rect 423200 640600 423400 640900
rect 423700 640600 424300 640900
rect 411700 640400 424300 640600
rect 411700 640100 411800 640400
rect 412100 640100 412300 640400
rect 412600 640100 422900 640400
rect 423200 640100 423400 640400
rect 423700 640100 424300 640400
rect 411700 640000 424300 640100
rect 3599 639799 4201 639800
rect 577899 633500 578201 633501
rect 577899 633200 577900 633500
rect 578200 633200 578201 633500
rect 577899 633199 578201 633200
rect 578399 633500 578701 633501
rect 578399 633200 578400 633500
rect 578700 633200 578701 633500
rect 578399 633199 578701 633200
rect 577899 633000 578201 633001
rect 577899 632700 577900 633000
rect 578200 632700 578201 633000
rect 577899 632699 578201 632700
rect 578399 633000 578701 633001
rect 578399 632700 578400 633000
rect 578700 632700 578701 633000
rect 578399 632699 578701 632700
rect 577899 632500 578201 632501
rect 577899 632200 577900 632500
rect 578200 632200 578201 632500
rect 577899 632199 578201 632200
rect 578399 632500 578701 632501
rect 578399 632200 578400 632500
rect 578700 632200 578701 632500
rect 578399 632199 578701 632200
rect 577899 632000 578201 632001
rect 541094 631905 541096 631906
rect 541094 631295 541095 631905
rect 577899 631700 577900 632000
rect 578200 631700 578201 632000
rect 577899 631699 578201 631700
rect 578399 632000 578701 632001
rect 578399 631700 578400 632000
rect 578700 631700 578701 632000
rect 578399 631699 578701 631700
rect 541094 631294 541096 631295
rect 577899 631500 578201 631501
rect 577899 631200 577900 631500
rect 578200 631200 578201 631500
rect 577899 631199 578201 631200
rect 578399 631500 578701 631501
rect 578399 631200 578400 631500
rect 578700 631200 578701 631500
rect 578399 631199 578701 631200
rect 577899 631000 578201 631001
rect 577899 630700 577900 631000
rect 578200 630700 578201 631000
rect 577899 630699 578201 630700
rect 578399 631000 578701 631001
rect 578399 630700 578400 631000
rect 578700 630700 578701 631000
rect 578399 630699 578701 630700
rect 577899 630500 578201 630501
rect 577899 630200 577900 630500
rect 578200 630200 578201 630500
rect 577899 630199 578201 630200
rect 578399 630500 578701 630501
rect 578399 630200 578400 630500
rect 578700 630200 578701 630500
rect 578399 630199 578701 630200
rect 49200 603800 50000 610200
rect 15200 603000 50000 603800
rect 15200 602800 43400 603000
rect 15200 602201 16000 602800
rect 24200 602201 25000 602800
rect 33400 602201 34200 602800
rect 42600 602201 43400 602800
rect 10199 602200 11001 602201
rect 10199 601400 10200 602200
rect 11000 601400 11001 602200
rect 10199 601399 11001 601400
rect 15199 602200 16001 602201
rect 15199 601400 15200 602200
rect 16000 601400 16001 602200
rect 15199 601399 16001 601400
rect 19199 602200 20001 602201
rect 19199 601400 19200 602200
rect 20000 601400 20001 602200
rect 19199 601399 20001 601400
rect 24199 602200 25001 602201
rect 24199 601400 24200 602200
rect 25000 601400 25001 602200
rect 24199 601399 25001 601400
rect 28399 602200 29201 602201
rect 28399 601400 28400 602200
rect 29200 601400 29201 602200
rect 28399 601399 29201 601400
rect 33399 602200 34201 602201
rect 33399 601400 33400 602200
rect 34200 601400 34201 602200
rect 33399 601399 34201 601400
rect 37599 602200 38401 602201
rect 37599 601400 37600 602200
rect 38400 601400 38401 602200
rect 37599 601399 38401 601400
rect 42599 602200 43401 602201
rect 42599 601400 42600 602200
rect 43400 601400 43401 602200
rect 42599 601399 43401 601400
<< via4 >>
rect 546000 678200 546300 678500
rect 546500 678200 546800 678500
rect 547000 678200 547300 678500
rect 547500 678200 547800 678500
rect 546000 677700 546300 678000
rect 546500 677700 546800 678000
rect 547000 677700 547300 678000
rect 547500 677700 547800 678000
rect 546000 677200 546300 677500
rect 546500 677200 546800 677500
rect 547000 677200 547300 677500
rect 547500 677200 547800 677500
rect 82400 676000 83200 676800
rect 131600 676000 132400 676800
rect 154400 676000 155200 676800
rect 329500 676100 329800 676400
rect 330000 676100 330300 676400
rect 330500 676100 330800 676400
rect 331000 676100 331300 676400
rect 331500 676100 331800 676400
rect 332000 676100 332300 676400
rect 332500 676100 332800 676400
rect 333000 676100 333300 676400
rect 333500 676100 333800 676400
rect 329500 675600 329800 675900
rect 330000 675600 330300 675900
rect 330500 675600 330800 675900
rect 331000 675600 331300 675900
rect 331500 675600 331800 675900
rect 332000 675600 332300 675900
rect 332500 675600 332800 675900
rect 333000 675600 333300 675900
rect 333500 675600 333800 675900
rect 329500 675100 329800 675400
rect 330000 675100 330300 675400
rect 330500 675100 330800 675400
rect 331000 675100 331300 675400
rect 331500 675100 331800 675400
rect 332000 675100 332300 675400
rect 332500 675100 332800 675400
rect 333000 675100 333300 675400
rect 333500 675100 333800 675400
rect 520800 673600 521400 674200
rect 521800 673600 522400 674200
rect 522800 673600 523400 674200
rect 523800 673600 524400 674200
rect 520800 672600 521400 673200
rect 521800 672600 522400 673200
rect 522800 672600 523400 673200
rect 523800 672600 524400 673200
rect 53200 670800 54000 671600
rect 520800 671600 521400 672200
rect 521800 671600 522400 672200
rect 522800 671600 523400 672200
rect 523800 671600 524400 672200
rect 520800 670600 521400 671200
rect 521800 670600 522400 671200
rect 522800 670600 523400 671200
rect 523800 670600 524400 671200
rect 406394 667224 408346 669176
rect 451404 668605 452206 668606
rect 451404 667806 451405 668605
rect 451405 667806 452205 668605
rect 452205 667806 452206 668605
rect 392000 649400 392600 650000
rect 393800 649400 394400 650000
rect 393000 648600 393600 649200
rect 392000 647600 392600 648200
rect 393800 647600 394400 648200
rect 448000 649000 449000 650000
rect 2400 643400 3000 644000
rect 3600 643400 4200 644000
rect 445994 643805 446806 643806
rect 401400 643000 402000 643600
rect 2400 642200 3000 642800
rect 3600 642200 4200 642800
rect 402900 643575 403500 643600
rect 402900 643000 402901 643575
rect 402901 643000 403499 643575
rect 403499 643000 403500 643575
rect 445994 643006 445995 643805
rect 445995 643006 446805 643805
rect 446805 643006 446806 643805
rect 458000 642400 459400 643400
rect 2400 641000 3000 641600
rect 3600 641000 4200 641600
rect 323700 641100 324000 641400
rect 324200 641100 324500 641400
rect 324700 641100 325000 641400
rect 330600 641100 330900 641400
rect 331100 641100 331400 641400
rect 323700 640600 324000 640900
rect 324200 640600 324500 640900
rect 324700 640600 325000 640900
rect 330600 640600 330900 640900
rect 331100 640600 331400 640900
rect 2400 639800 3000 640400
rect 3600 639800 4200 640400
rect 323700 640100 324000 640400
rect 324200 640100 324500 640400
rect 324700 640100 325000 640400
rect 330600 640100 330900 640400
rect 331100 640100 331400 640400
rect 398800 640200 399800 641200
rect 411800 641100 412100 641400
rect 412300 641100 412600 641400
rect 422900 641100 423200 641400
rect 423400 641100 423700 641400
rect 411800 640600 412100 640900
rect 412300 640600 412600 640900
rect 422900 640600 423200 640900
rect 423400 640600 423700 640900
rect 411800 640100 412100 640400
rect 412300 640100 412600 640400
rect 422900 640100 423200 640400
rect 423400 640100 423700 640400
rect 577900 633200 578200 633500
rect 578400 633200 578700 633500
rect 577900 632700 578200 633000
rect 578400 632700 578700 633000
rect 577900 632200 578200 632500
rect 578400 632200 578700 632500
rect 541096 631905 541696 631906
rect 541096 631295 541695 631905
rect 541695 631295 541696 631905
rect 577900 631700 578200 632000
rect 578400 631700 578700 632000
rect 541096 631294 541696 631295
rect 577900 631200 578200 631500
rect 578400 631200 578700 631500
rect 577900 630700 578200 631000
rect 578400 630700 578700 631000
rect 577900 630200 578200 630500
rect 578400 630200 578700 630500
rect 10200 601400 11000 602200
rect 19200 601400 20000 602200
rect 28400 601400 29200 602200
rect 37600 601400 38400 602200
<< metal5 >>
rect 165594 702300 170594 704800
rect 175894 702300 180894 704800
rect 217294 704000 222294 704800
rect 227594 704000 232594 704800
rect 217294 703100 232594 704000
rect 318994 704000 324000 704800
rect 329300 704000 334294 704800
rect 217294 702300 232600 703100
rect 318994 702800 334294 704000
rect 318994 702300 334300 702800
rect 217300 702000 232600 702300
rect 82376 676800 83224 676824
rect 131576 676800 132424 676824
rect 154376 676800 155224 676824
rect 82376 676000 82400 676800
rect 83200 676000 131600 676800
rect 132400 676000 154400 676800
rect 155200 676000 155224 676800
rect 82376 675976 83224 676000
rect 53176 671600 54024 671624
rect 53176 670800 53200 671600
rect 54000 670800 54024 671600
rect 53176 670776 54024 670800
rect 53200 667400 54000 670776
rect 53200 666600 75800 667400
rect 91400 666600 92400 676000
rect 131576 675976 132424 676000
rect 154376 675976 155224 676000
rect 2200 644000 77200 644200
rect 2200 643400 2400 644000
rect 3000 643400 3600 644000
rect 4200 643400 77200 644000
rect 2200 642800 77200 643400
rect 2200 642200 2400 642800
rect 3000 642200 3600 642800
rect 4200 642200 77200 642800
rect 2200 641600 77200 642200
rect 2200 641000 2400 641600
rect 3000 641000 3600 641600
rect 4200 641000 77200 641600
rect 2200 640400 77200 641000
rect 2200 639800 2400 640400
rect 3000 639800 3600 640400
rect 4200 639800 77200 640400
rect 227600 641500 232600 702000
rect 319000 701900 334300 702300
rect 329300 676400 334300 701900
rect 502500 678500 547900 678600
rect 502500 678200 546000 678500
rect 546300 678200 546500 678500
rect 546800 678200 547000 678500
rect 547300 678200 547500 678500
rect 547800 678200 547900 678500
rect 502500 678000 547900 678200
rect 502500 677700 546000 678000
rect 546300 677700 546500 678000
rect 546800 677700 547000 678000
rect 547300 677700 547500 678000
rect 547800 677700 547900 678000
rect 502500 677500 547900 677700
rect 502500 677200 546000 677500
rect 546300 677200 546500 677500
rect 546800 677200 547000 677500
rect 547300 677200 547500 677500
rect 547800 677200 547900 677500
rect 502500 677100 547900 677200
rect 329300 676100 329500 676400
rect 329800 676100 330000 676400
rect 330300 676100 330500 676400
rect 330800 676100 331000 676400
rect 331300 676100 331500 676400
rect 331800 676100 332000 676400
rect 332300 676100 332500 676400
rect 332800 676100 333000 676400
rect 333300 676100 333500 676400
rect 333800 676100 334300 676400
rect 329300 675900 334300 676100
rect 329300 675600 329500 675900
rect 329800 675600 330000 675900
rect 330300 675600 330500 675900
rect 330800 675600 331000 675900
rect 331300 675600 331500 675900
rect 331800 675600 332000 675900
rect 332300 675600 332500 675900
rect 332800 675600 333000 675900
rect 333300 675600 333500 675900
rect 333800 675600 334300 675900
rect 329300 675400 334300 675600
rect 329300 675100 329500 675400
rect 329800 675100 330000 675400
rect 330300 675100 330500 675400
rect 330800 675100 331000 675400
rect 331300 675100 331500 675400
rect 331800 675100 332000 675400
rect 332300 675100 332500 675400
rect 332800 675100 333000 675400
rect 333300 675100 333500 675400
rect 333800 675100 334300 675400
rect 329300 674900 334300 675100
rect 520776 674200 521424 674224
rect 520776 673600 520800 674200
rect 521400 673600 521424 674200
rect 520776 673576 521424 673600
rect 521776 674200 522424 674224
rect 521776 673600 521800 674200
rect 522400 673600 522424 674200
rect 521776 673576 522424 673600
rect 522776 674200 523424 674224
rect 522776 673600 522800 674200
rect 523400 673600 523424 674200
rect 522776 673576 523424 673600
rect 523776 674200 524424 674224
rect 523776 673600 523800 674200
rect 524400 673600 524424 674200
rect 523776 673576 524424 673600
rect 520776 673200 521424 673224
rect 520776 672600 520800 673200
rect 521400 672600 521424 673200
rect 520776 672576 521424 672600
rect 521776 673200 522424 673224
rect 521776 672600 521800 673200
rect 522400 672600 522424 673200
rect 521776 672576 522424 672600
rect 522776 673200 523424 673224
rect 522776 672600 522800 673200
rect 523400 672600 523424 673200
rect 522776 672576 523424 672600
rect 523776 673200 524424 673224
rect 523776 672600 523800 673200
rect 524400 672600 524424 673200
rect 523776 672576 524424 672600
rect 520776 672200 521424 672224
rect 520776 671600 520800 672200
rect 521400 671600 521424 672200
rect 520776 671576 521424 671600
rect 521776 672200 522424 672224
rect 521776 671600 521800 672200
rect 522400 671600 522424 672200
rect 521776 671576 522424 671600
rect 522776 672200 523424 672224
rect 522776 671600 522800 672200
rect 523400 671600 523424 672200
rect 522776 671576 523424 671600
rect 523776 672200 524424 672224
rect 523776 671600 523800 672200
rect 524400 671600 524424 672200
rect 523776 671576 524424 671600
rect 520776 671200 521424 671224
rect 520776 670600 520800 671200
rect 521400 670600 521424 671200
rect 520776 670576 521424 670600
rect 521776 671200 522424 671224
rect 521776 670600 521800 671200
rect 522400 670600 522424 671200
rect 521776 670576 522424 670600
rect 522776 671200 523424 671224
rect 522776 670600 522800 671200
rect 523400 670600 523424 671200
rect 522776 670576 523424 670600
rect 523776 671200 524424 671224
rect 523776 670600 523800 671200
rect 524400 670600 524424 671200
rect 523776 670576 524424 670600
rect 406370 669176 455800 669200
rect 406370 667224 406394 669176
rect 408346 668606 455800 669176
rect 408346 667806 451404 668606
rect 452206 667806 455800 668606
rect 408346 667224 455800 667806
rect 406370 667200 455800 667224
rect 391400 650000 450000 651000
rect 391400 649400 392000 650000
rect 392600 649400 393800 650000
rect 394400 649400 448000 650000
rect 391400 649200 448000 649400
rect 391400 648600 393000 649200
rect 393600 649000 448000 649200
rect 449000 649000 450000 650000
rect 393600 648600 450000 649000
rect 391400 648200 450000 648600
rect 391400 647600 392000 648200
rect 392600 647600 393800 648200
rect 394400 648000 450000 648200
rect 394400 647600 395000 648000
rect 391400 647000 395000 647600
rect 445970 643806 446830 643830
rect 401200 643600 402200 643800
rect 402876 643600 403524 643624
rect 445970 643600 445994 643806
rect 401200 643000 401400 643600
rect 402000 643000 402900 643600
rect 403500 643006 445994 643600
rect 446806 643600 446830 643806
rect 446806 643400 459600 643600
rect 446806 643006 458000 643400
rect 403500 643000 458000 643006
rect 401200 642800 402200 643000
rect 402876 642976 403524 643000
rect 445970 642982 446830 643000
rect 457800 642400 458000 643000
rect 459400 642400 459600 643400
rect 457800 642200 459600 642400
rect 227600 641400 325500 641500
rect 227600 641100 323700 641400
rect 324000 641100 324200 641400
rect 324500 641100 324700 641400
rect 325000 641100 325500 641400
rect 227600 640900 325500 641100
rect 227600 640600 323700 640900
rect 324000 640600 324200 640900
rect 324500 640600 324700 640900
rect 325000 640600 325500 640900
rect 227600 640400 325500 640600
rect 227600 640100 323700 640400
rect 324000 640100 324200 640400
rect 324500 640100 324700 640400
rect 325000 640100 325500 640400
rect 227600 640000 325500 640100
rect 330400 641400 412800 641500
rect 330400 641100 330600 641400
rect 330900 641100 331100 641400
rect 331400 641200 411800 641400
rect 331400 641100 398800 641200
rect 330400 640900 398800 641100
rect 330400 640600 330600 640900
rect 330900 640600 331100 640900
rect 331400 640600 398800 640900
rect 330400 640400 398800 640600
rect 330400 640100 330600 640400
rect 330900 640100 331100 640400
rect 331400 640200 398800 640400
rect 399800 641100 411800 641200
rect 412100 641100 412300 641400
rect 412600 641100 412800 641400
rect 399800 640900 412800 641100
rect 399800 640600 411800 640900
rect 412100 640600 412300 640900
rect 412600 640600 412800 640900
rect 399800 640400 412800 640600
rect 399800 640200 411800 640400
rect 331400 640100 411800 640200
rect 412100 640100 412300 640400
rect 412600 640100 412800 640400
rect 330400 640000 412800 640100
rect 422800 641400 457300 641500
rect 422800 641100 422900 641400
rect 423200 641100 423400 641400
rect 423700 641100 457300 641400
rect 422800 640900 457300 641100
rect 422800 640600 422900 640900
rect 423200 640600 423400 640900
rect 423700 640600 457300 640900
rect 422800 640400 457300 640600
rect 422800 640100 422900 640400
rect 423200 640100 423400 640400
rect 423700 640100 457300 640400
rect 422800 640000 457300 640100
rect 2200 639600 77200 639800
rect 514200 633500 580000 634000
rect 514200 633200 577900 633500
rect 578200 633200 578400 633500
rect 578700 633200 580000 633500
rect 514200 633000 580000 633200
rect 514200 632700 577900 633000
rect 578200 632700 578400 633000
rect 578700 632700 580000 633000
rect 514200 632500 580000 632700
rect 514200 632200 577900 632500
rect 578200 632200 578400 632500
rect 578700 632200 580000 632500
rect 514200 632000 580000 632200
rect 514200 631906 577900 632000
rect 514200 631294 541096 631906
rect 541696 631700 577900 631906
rect 578200 631700 578400 632000
rect 578700 631700 580000 632000
rect 541696 631500 580000 631700
rect 541696 631294 577900 631500
rect 514200 631200 577900 631294
rect 578200 631200 578400 631500
rect 578700 631200 580000 631500
rect 514200 631000 580000 631200
rect 514200 630700 577900 631000
rect 578200 630700 578400 631000
rect 578700 630700 580000 631000
rect 514200 630500 580000 630700
rect 514200 630200 577900 630500
rect 578200 630200 578400 630500
rect 578700 630200 580000 630500
rect 514200 630100 580000 630200
rect 515000 630000 521000 630100
rect 10176 602200 11024 602224
rect 19176 602200 20024 602224
rect 28376 602200 29224 602224
rect 37576 602200 38424 602224
rect 49200 602200 50000 614600
rect 10176 601400 10200 602200
rect 11000 601400 19200 602200
rect 20000 601400 28400 602200
rect 29200 601400 37600 602200
rect 38400 601400 50000 602200
rect 10176 601376 11024 601400
rect 19176 601376 20024 601400
rect 28376 601376 29224 601400
rect 37576 601376 38424 601400
<< comment >>
rect -100 704000 584100 704100
rect -100 0 0 704000
rect 584000 0 584100 704000
rect -100 -100 584100 0
use chip_art  chip_art_0
timestamp 1717028336
transform 1 0 61200 0 1 40000
box -1200 0 201200 200000
use chip_art_inv  chip_art_inv_0
timestamp 1717029187
transform 1 0 321200 0 1 40000
box -1200 0 201200 200000
use DS_2024_2p2  DS_2024_2p2_0
timestamp 1717179484
transform -1 0 685396 0 -1 626372
box 135892 -55212 236396 -3628
use ESD  ESD_0
timestamp 1717181165
transform 1 0 388066 0 1 644880
box 0 -2700 12000 3200
use ESD  ESD_1
timestamp 1717181165
transform 0 -1 56400 -1 0 676800
box 0 -2700 12000 3200
use ESD  ESD_2
timestamp 1717181165
transform 1 0 381600 0 1 680700
box 0 -2700 12000 3200
use ESD  ESD_3
timestamp 1717181165
transform 0 1 405992 -1 0 699456
box 0 -2700 12000 3200
use ESD  ESD_4
timestamp 1717181165
transform 0 1 449036 -1 0 694562
box 0 -2700 12000 3200
use ESD  ESD_5
timestamp 1717181165
transform 1 0 555200 0 1 671100
box 0 -2700 12000 3200
use ESD  ESD_6
timestamp 1717181165
transform 0 1 542100 -1 0 694400
box 0 -2700 12000 3200
use ESD  ESD_7
timestamp 1717181165
transform 0 -1 13400 1 0 596200
box 0 -2700 12000 3200
use ESD  ESD_8
timestamp 1717181165
transform -1 0 160400 0 1 673500
box 0 -2700 12000 3200
use ESD  ESD_9
timestamp 1717181165
transform -1 0 137600 0 1 673500
box 0 -2700 12000 3200
use ESD  ESD_10
timestamp 1717181165
transform 0 -1 40800 1 0 596200
box 0 -2700 12000 3200
use ESD  ESD_11
timestamp 1717181165
transform 0 -1 31600 1 0 596200
box 0 -2700 12000 3200
use ESD  ESD_12
timestamp 1717181165
transform 0 -1 22400 1 0 596200
box 0 -2700 12000 3200
use ESD  ESD_13
timestamp 1717181165
transform 1 0 77200 0 1 673500
box 0 -2700 12000 3200
use flashADC  flashADC_0
timestamp 1717179484
transform -1 0 140600 0 1 664800
box -33300 -86800 95800 5000
<< labels >>
flabel metal3 s 583520 269230 584800 269342 0 FreeSans 1120 0 0 0 gpio_analog[0]
port 0 nsew signal bidirectional
flabel metal3 s -800 381864 480 381976 0 FreeSans 1120 0 0 0 gpio_analog[10]
port 1 nsew signal bidirectional
flabel metal3 s -800 338642 480 338754 0 FreeSans 1120 0 0 0 gpio_analog[11]
port 2 nsew signal bidirectional
flabel metal3 s -800 295420 480 295532 0 FreeSans 1120 0 0 0 gpio_analog[12]
port 3 nsew signal bidirectional
flabel metal3 s -800 252398 480 252510 0 FreeSans 1120 0 0 0 gpio_analog[13]
port 4 nsew signal bidirectional
flabel metal3 s -800 124776 480 124888 0 FreeSans 1120 0 0 0 gpio_analog[14]
port 5 nsew signal bidirectional
flabel metal3 s -800 81554 480 81666 0 FreeSans 1120 0 0 0 gpio_analog[15]
port 6 nsew signal bidirectional
flabel metal3 s -800 38332 480 38444 0 FreeSans 1120 0 0 0 gpio_analog[16]
port 7 nsew signal bidirectional
flabel metal3 s -800 16910 480 17022 0 FreeSans 1120 0 0 0 gpio_analog[17]
port 8 nsew signal bidirectional
flabel metal3 s 583520 313652 584800 313764 0 FreeSans 1120 0 0 0 gpio_analog[1]
port 9 nsew signal bidirectional
flabel metal3 s 583520 358874 584800 358986 0 FreeSans 1120 0 0 0 gpio_analog[2]
port 10 nsew signal bidirectional
flabel metal3 s 583520 405296 584800 405408 0 FreeSans 1120 0 0 0 gpio_analog[3]
port 11 nsew signal bidirectional
flabel metal3 s 583520 449718 584800 449830 0 FreeSans 1120 0 0 0 gpio_analog[4]
port 12 nsew signal bidirectional
flabel metal3 s 583520 494140 584800 494252 0 FreeSans 1120 0 0 0 gpio_analog[5]
port 13 nsew signal bidirectional
flabel metal3 s 583520 583562 584800 583674 0 FreeSans 1120 0 0 0 gpio_analog[6]
port 14 nsew signal bidirectional
flabel metal3 s -800 511530 480 511642 0 FreeSans 1120 0 0 0 gpio_analog[7]
port 15 nsew signal bidirectional
flabel metal3 s -800 468308 480 468420 0 FreeSans 1120 0 0 0 gpio_analog[8]
port 16 nsew signal bidirectional
flabel metal3 s -800 425086 480 425198 0 FreeSans 1120 0 0 0 gpio_analog[9]
port 17 nsew signal bidirectional
flabel metal3 s 583520 270412 584800 270524 0 FreeSans 1120 0 0 0 gpio_noesd[0]
port 18 nsew signal bidirectional
flabel metal3 s -800 380682 480 380794 0 FreeSans 1120 0 0 0 gpio_noesd[10]
port 19 nsew signal bidirectional
flabel metal3 s -800 337460 480 337572 0 FreeSans 1120 0 0 0 gpio_noesd[11]
port 20 nsew signal bidirectional
flabel metal3 s -800 294238 480 294350 0 FreeSans 1120 0 0 0 gpio_noesd[12]
port 21 nsew signal bidirectional
flabel metal3 s -800 251216 480 251328 0 FreeSans 1120 0 0 0 gpio_noesd[13]
port 22 nsew signal bidirectional
flabel metal3 s -800 123594 480 123706 0 FreeSans 1120 0 0 0 gpio_noesd[14]
port 23 nsew signal bidirectional
flabel metal3 s -800 80372 480 80484 0 FreeSans 1120 0 0 0 gpio_noesd[15]
port 24 nsew signal bidirectional
flabel metal3 s -800 37150 480 37262 0 FreeSans 1120 0 0 0 gpio_noesd[16]
port 25 nsew signal bidirectional
flabel metal3 s -800 15728 480 15840 0 FreeSans 1120 0 0 0 gpio_noesd[17]
port 26 nsew signal bidirectional
flabel metal3 s 583520 314834 584800 314946 0 FreeSans 1120 0 0 0 gpio_noesd[1]
port 27 nsew signal bidirectional
flabel metal3 s 583520 360056 584800 360168 0 FreeSans 1120 0 0 0 gpio_noesd[2]
port 28 nsew signal bidirectional
flabel metal3 s 583520 406478 584800 406590 0 FreeSans 1120 0 0 0 gpio_noesd[3]
port 29 nsew signal bidirectional
flabel metal3 s 583520 450900 584800 451012 0 FreeSans 1120 0 0 0 gpio_noesd[4]
port 30 nsew signal bidirectional
flabel metal3 s 583520 495322 584800 495434 0 FreeSans 1120 0 0 0 gpio_noesd[5]
port 31 nsew signal bidirectional
flabel metal3 s 583520 584744 584800 584856 0 FreeSans 1120 0 0 0 gpio_noesd[6]
port 32 nsew signal bidirectional
flabel metal3 s -800 510348 480 510460 0 FreeSans 1120 0 0 0 gpio_noesd[7]
port 33 nsew signal bidirectional
flabel metal3 s -800 467126 480 467238 0 FreeSans 1120 0 0 0 gpio_noesd[8]
port 34 nsew signal bidirectional
flabel metal3 s -800 423904 480 424016 0 FreeSans 1120 0 0 0 gpio_noesd[9]
port 35 nsew signal bidirectional
flabel metal3 s 582300 677984 584800 682984 0 FreeSans 1120 0 0 0 io_analog[0]
port 36 nsew signal bidirectional
flabel metal3 s 0 680242 1700 685242 0 FreeSans 1120 0 0 0 io_analog[10]
port 37 nsew signal bidirectional
flabel metal3 s 566594 702300 571594 704800 0 FreeSans 1920 180 0 0 io_analog[1]
port 38 nsew signal bidirectional
flabel metal3 s 465394 702300 470394 704800 0 FreeSans 1920 180 0 0 io_analog[2]
port 39 nsew signal bidirectional
flabel metal3 s 413394 702300 418394 704800 0 FreeSans 1920 180 0 0 io_analog[3]
port 40 nsew signal bidirectional
flabel metal3 s 329294 702300 334294 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 41 nsew signal bidirectional
flabel metal5 s 329294 702300 334294 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 41 nsew signal bidirectional
flabel metal3 s 227594 702300 232594 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 42 nsew signal bidirectional
flabel metal4 s 227594 702300 232594 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 42 nsew signal bidirectional
flabel metal5 s 227594 702300 232594 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 42 nsew signal bidirectional
flabel metal3 s 175894 702300 180894 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 43 nsew signal bidirectional
flabel metal4 s 175894 702300 180894 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 43 nsew signal bidirectional
flabel metal5 s 175894 702300 180894 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 43 nsew signal bidirectional
flabel metal3 s 120194 702300 125194 704800 0 FreeSans 1920 180 0 0 io_analog[7]
port 44 nsew signal bidirectional
flabel metal3 s 68194 702300 73194 704800 0 FreeSans 1920 180 0 0 io_analog[8]
port 45 nsew signal bidirectional
flabel metal3 s 16194 702300 21194 704800 0 FreeSans 1920 180 0 0 io_analog[9]
port 46 nsew signal bidirectional
flabel metal3 s 318994 702300 323994 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 47 nsew signal bidirectional
flabel metal5 s 318994 702300 323994 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 47 nsew signal bidirectional
flabel metal3 s 217294 702300 222294 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 48 nsew signal bidirectional
flabel metal4 s 217294 702300 222294 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 48 nsew signal bidirectional
flabel metal5 s 217294 702300 222294 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 48 nsew signal bidirectional
flabel metal3 s 165594 702300 170594 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 49 nsew signal bidirectional
flabel metal4 s 165594 702300 170594 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 49 nsew signal bidirectional
flabel metal5 s 165594 702300 170594 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 49 nsew signal bidirectional
flabel metal3 s 326794 702300 328994 704800 0 FreeSans 1920 180 0 0 io_clamp_high[0]
port 50 nsew signal bidirectional
flabel metal3 s 225094 702300 227294 704800 0 FreeSans 1920 180 0 0 io_clamp_high[1]
port 51 nsew signal bidirectional
flabel metal3 s 173394 702300 175594 704800 0 FreeSans 1920 180 0 0 io_clamp_high[2]
port 52 nsew signal bidirectional
flabel metal3 s 324294 702300 326494 704800 0 FreeSans 1920 180 0 0 io_clamp_low[0]
port 53 nsew signal bidirectional
flabel metal3 s 222594 702300 224794 704800 0 FreeSans 1920 180 0 0 io_clamp_low[1]
port 54 nsew signal bidirectional
flabel metal3 s 170894 702300 173094 704800 0 FreeSans 1920 180 0 0 io_clamp_low[2]
port 55 nsew signal bidirectional
flabel metal3 s 583520 2726 584800 2838 0 FreeSans 1120 0 0 0 io_in[0]
port 56 nsew signal input
flabel metal3 s 583520 408842 584800 408954 0 FreeSans 1120 0 0 0 io_in[10]
port 57 nsew signal input
flabel metal3 s 583520 453264 584800 453376 0 FreeSans 1120 0 0 0 io_in[11]
port 58 nsew signal input
flabel metal3 s 583520 497686 584800 497798 0 FreeSans 1120 0 0 0 io_in[12]
port 59 nsew signal input
flabel metal3 s 583520 587108 584800 587220 0 FreeSans 1120 0 0 0 io_in[13]
port 60 nsew signal input
flabel metal3 s -800 507984 480 508096 0 FreeSans 1120 0 0 0 io_in[14]
port 61 nsew signal input
flabel metal3 s -800 464762 480 464874 0 FreeSans 1120 0 0 0 io_in[15]
port 62 nsew signal input
flabel metal3 s -800 421540 480 421652 0 FreeSans 1120 0 0 0 io_in[16]
port 63 nsew signal input
flabel metal3 s -800 378318 480 378430 0 FreeSans 1120 0 0 0 io_in[17]
port 64 nsew signal input
flabel metal3 s -800 335096 480 335208 0 FreeSans 1120 0 0 0 io_in[18]
port 65 nsew signal input
flabel metal3 s -800 291874 480 291986 0 FreeSans 1120 0 0 0 io_in[19]
port 66 nsew signal input
flabel metal3 s 583520 7454 584800 7566 0 FreeSans 1120 0 0 0 io_in[1]
port 67 nsew signal input
flabel metal3 s -800 248852 480 248964 0 FreeSans 1120 0 0 0 io_in[20]
port 68 nsew signal input
flabel metal3 s -800 121230 480 121342 0 FreeSans 1120 0 0 0 io_in[21]
port 69 nsew signal input
flabel metal3 s -800 78008 480 78120 0 FreeSans 1120 0 0 0 io_in[22]
port 70 nsew signal input
flabel metal3 s -800 34786 480 34898 0 FreeSans 1120 0 0 0 io_in[23]
port 71 nsew signal input
flabel metal3 s -800 13364 480 13476 0 FreeSans 1120 0 0 0 io_in[24]
port 72 nsew signal input
flabel metal3 s -800 8636 480 8748 0 FreeSans 1120 0 0 0 io_in[25]
port 73 nsew signal input
flabel metal3 s -800 3908 480 4020 0 FreeSans 1120 0 0 0 io_in[26]
port 74 nsew signal input
flabel metal3 s 583520 12182 584800 12294 0 FreeSans 1120 0 0 0 io_in[2]
port 75 nsew signal input
flabel metal3 s 583520 16910 584800 17022 0 FreeSans 1120 0 0 0 io_in[3]
port 76 nsew signal input
flabel metal3 s 583520 21638 584800 21750 0 FreeSans 1120 0 0 0 io_in[4]
port 77 nsew signal input
flabel metal3 s 583520 48096 584800 48208 0 FreeSans 1120 0 0 0 io_in[5]
port 78 nsew signal input
flabel metal3 s 583520 92754 584800 92866 0 FreeSans 1120 0 0 0 io_in[6]
port 79 nsew signal input
flabel metal3 s 583520 272776 584800 272888 0 FreeSans 1120 0 0 0 io_in[7]
port 80 nsew signal input
flabel metal3 s 583520 317198 584800 317310 0 FreeSans 1120 0 0 0 io_in[8]
port 81 nsew signal input
flabel metal3 s 583520 362420 584800 362532 0 FreeSans 1120 0 0 0 io_in[9]
port 82 nsew signal input
flabel metal3 s 583520 1544 584800 1656 0 FreeSans 1120 0 0 0 io_in_3v3[0]
port 83 nsew signal input
flabel metal3 s 583520 407660 584800 407772 0 FreeSans 1120 0 0 0 io_in_3v3[10]
port 84 nsew signal input
flabel metal3 s 583520 452082 584800 452194 0 FreeSans 1120 0 0 0 io_in_3v3[11]
port 85 nsew signal input
flabel metal3 s 583520 496504 584800 496616 0 FreeSans 1120 0 0 0 io_in_3v3[12]
port 86 nsew signal input
flabel metal3 s 583520 585926 584800 586038 0 FreeSans 1120 0 0 0 io_in_3v3[13]
port 87 nsew signal input
flabel metal3 s -800 509166 480 509278 0 FreeSans 1120 0 0 0 io_in_3v3[14]
port 88 nsew signal input
flabel metal3 s -800 465944 480 466056 0 FreeSans 1120 0 0 0 io_in_3v3[15]
port 89 nsew signal input
flabel metal3 s -800 422722 480 422834 0 FreeSans 1120 0 0 0 io_in_3v3[16]
port 90 nsew signal input
flabel metal3 s -800 379500 480 379612 0 FreeSans 1120 0 0 0 io_in_3v3[17]
port 91 nsew signal input
flabel metal3 s -800 336278 480 336390 0 FreeSans 1120 0 0 0 io_in_3v3[18]
port 92 nsew signal input
flabel metal3 s -800 293056 480 293168 0 FreeSans 1120 0 0 0 io_in_3v3[19]
port 93 nsew signal input
flabel metal3 s 583520 6272 584800 6384 0 FreeSans 1120 0 0 0 io_in_3v3[1]
port 94 nsew signal input
flabel metal3 s -800 250034 480 250146 0 FreeSans 1120 0 0 0 io_in_3v3[20]
port 95 nsew signal input
flabel metal3 s -800 122412 480 122524 0 FreeSans 1120 0 0 0 io_in_3v3[21]
port 96 nsew signal input
flabel metal3 s -800 79190 480 79302 0 FreeSans 1120 0 0 0 io_in_3v3[22]
port 97 nsew signal input
flabel metal3 s -800 35968 480 36080 0 FreeSans 1120 0 0 0 io_in_3v3[23]
port 98 nsew signal input
flabel metal3 s -800 14546 480 14658 0 FreeSans 1120 0 0 0 io_in_3v3[24]
port 99 nsew signal input
flabel metal3 s -800 9818 480 9930 0 FreeSans 1120 0 0 0 io_in_3v3[25]
port 100 nsew signal input
flabel metal3 s -800 5090 480 5202 0 FreeSans 1120 0 0 0 io_in_3v3[26]
port 101 nsew signal input
flabel metal3 s 583520 11000 584800 11112 0 FreeSans 1120 0 0 0 io_in_3v3[2]
port 102 nsew signal input
flabel metal3 s 583520 15728 584800 15840 0 FreeSans 1120 0 0 0 io_in_3v3[3]
port 103 nsew signal input
flabel metal3 s 583520 20456 584800 20568 0 FreeSans 1120 0 0 0 io_in_3v3[4]
port 104 nsew signal input
flabel metal3 s 583520 46914 584800 47026 0 FreeSans 1120 0 0 0 io_in_3v3[5]
port 105 nsew signal input
flabel metal3 s 583520 91572 584800 91684 0 FreeSans 1120 0 0 0 io_in_3v3[6]
port 106 nsew signal input
flabel metal3 s 583520 271594 584800 271706 0 FreeSans 1120 0 0 0 io_in_3v3[7]
port 107 nsew signal input
flabel metal3 s 583520 316016 584800 316128 0 FreeSans 1120 0 0 0 io_in_3v3[8]
port 108 nsew signal input
flabel metal3 s 583520 361238 584800 361350 0 FreeSans 1120 0 0 0 io_in_3v3[9]
port 109 nsew signal input
flabel metal3 s 583520 5090 584800 5202 0 FreeSans 1120 0 0 0 io_oeb[0]
port 110 nsew signal tristate
flabel metal3 s 583520 411206 584800 411318 0 FreeSans 1120 0 0 0 io_oeb[10]
port 111 nsew signal tristate
flabel metal3 s 583520 455628 584800 455740 0 FreeSans 1120 0 0 0 io_oeb[11]
port 112 nsew signal tristate
flabel metal3 s 583520 500050 584800 500162 0 FreeSans 1120 0 0 0 io_oeb[12]
port 113 nsew signal tristate
flabel metal3 s 583520 589472 584800 589584 0 FreeSans 1120 0 0 0 io_oeb[13]
port 114 nsew signal tristate
flabel metal3 s -800 505620 480 505732 0 FreeSans 1120 0 0 0 io_oeb[14]
port 115 nsew signal tristate
flabel metal3 s -800 462398 480 462510 0 FreeSans 1120 0 0 0 io_oeb[15]
port 116 nsew signal tristate
flabel metal3 s -800 419176 480 419288 0 FreeSans 1120 0 0 0 io_oeb[16]
port 117 nsew signal tristate
flabel metal3 s -800 375954 480 376066 0 FreeSans 1120 0 0 0 io_oeb[17]
port 118 nsew signal tristate
flabel metal3 s -800 332732 480 332844 0 FreeSans 1120 0 0 0 io_oeb[18]
port 119 nsew signal tristate
flabel metal3 s -800 289510 480 289622 0 FreeSans 1120 0 0 0 io_oeb[19]
port 120 nsew signal tristate
flabel metal3 s 583520 9818 584800 9930 0 FreeSans 1120 0 0 0 io_oeb[1]
port 121 nsew signal tristate
flabel metal3 s -800 246488 480 246600 0 FreeSans 1120 0 0 0 io_oeb[20]
port 122 nsew signal tristate
flabel metal3 s -800 118866 480 118978 0 FreeSans 1120 0 0 0 io_oeb[21]
port 123 nsew signal tristate
flabel metal3 s -800 75644 480 75756 0 FreeSans 1120 0 0 0 io_oeb[22]
port 124 nsew signal tristate
flabel metal3 s -800 32422 480 32534 0 FreeSans 1120 0 0 0 io_oeb[23]
port 125 nsew signal tristate
flabel metal3 s -800 11000 480 11112 0 FreeSans 1120 0 0 0 io_oeb[24]
port 126 nsew signal tristate
flabel metal3 s -800 6272 480 6384 0 FreeSans 1120 0 0 0 io_oeb[25]
port 127 nsew signal tristate
flabel metal3 s -800 1544 480 1656 0 FreeSans 1120 0 0 0 io_oeb[26]
port 128 nsew signal tristate
flabel metal3 s 583520 14546 584800 14658 0 FreeSans 1120 0 0 0 io_oeb[2]
port 129 nsew signal tristate
flabel metal3 s 583520 19274 584800 19386 0 FreeSans 1120 0 0 0 io_oeb[3]
port 130 nsew signal tristate
flabel metal3 s 583520 24002 584800 24114 0 FreeSans 1120 0 0 0 io_oeb[4]
port 131 nsew signal tristate
flabel metal3 s 583520 50460 584800 50572 0 FreeSans 1120 0 0 0 io_oeb[5]
port 132 nsew signal tristate
flabel metal3 s 583520 95118 584800 95230 0 FreeSans 1120 0 0 0 io_oeb[6]
port 133 nsew signal tristate
flabel metal3 s 583520 275140 584800 275252 0 FreeSans 1120 0 0 0 io_oeb[7]
port 134 nsew signal tristate
flabel metal3 s 583520 319562 584800 319674 0 FreeSans 1120 0 0 0 io_oeb[8]
port 135 nsew signal tristate
flabel metal3 s 583520 364784 584800 364896 0 FreeSans 1120 0 0 0 io_oeb[9]
port 136 nsew signal tristate
flabel metal3 s 583520 3908 584800 4020 0 FreeSans 1120 0 0 0 io_out[0]
port 137 nsew signal tristate
flabel metal3 s 583520 410024 584800 410136 0 FreeSans 1120 0 0 0 io_out[10]
port 138 nsew signal tristate
flabel metal3 s 583520 454446 584800 454558 0 FreeSans 1120 0 0 0 io_out[11]
port 139 nsew signal tristate
flabel metal3 s 583520 498868 584800 498980 0 FreeSans 1120 0 0 0 io_out[12]
port 140 nsew signal tristate
flabel metal3 s 583520 588290 584800 588402 0 FreeSans 1120 0 0 0 io_out[13]
port 141 nsew signal tristate
flabel metal3 s -800 506802 480 506914 0 FreeSans 1120 0 0 0 io_out[14]
port 142 nsew signal tristate
flabel metal3 s -800 463580 480 463692 0 FreeSans 1120 0 0 0 io_out[15]
port 143 nsew signal tristate
flabel metal3 s -800 420358 480 420470 0 FreeSans 1120 0 0 0 io_out[16]
port 144 nsew signal tristate
flabel metal3 s -800 377136 480 377248 0 FreeSans 1120 0 0 0 io_out[17]
port 145 nsew signal tristate
flabel metal3 s -800 333914 480 334026 0 FreeSans 1120 0 0 0 io_out[18]
port 146 nsew signal tristate
flabel metal3 s -800 290692 480 290804 0 FreeSans 1120 0 0 0 io_out[19]
port 147 nsew signal tristate
flabel metal3 s 583520 8636 584800 8748 0 FreeSans 1120 0 0 0 io_out[1]
port 148 nsew signal tristate
flabel metal3 s -800 247670 480 247782 0 FreeSans 1120 0 0 0 io_out[20]
port 149 nsew signal tristate
flabel metal3 s -800 120048 480 120160 0 FreeSans 1120 0 0 0 io_out[21]
port 150 nsew signal tristate
flabel metal3 s -800 76826 480 76938 0 FreeSans 1120 0 0 0 io_out[22]
port 151 nsew signal tristate
flabel metal3 s -800 33604 480 33716 0 FreeSans 1120 0 0 0 io_out[23]
port 152 nsew signal tristate
flabel metal3 s -800 12182 480 12294 0 FreeSans 1120 0 0 0 io_out[24]
port 153 nsew signal tristate
flabel metal3 s -800 7454 480 7566 0 FreeSans 1120 0 0 0 io_out[25]
port 154 nsew signal tristate
flabel metal3 s -800 2726 480 2838 0 FreeSans 1120 0 0 0 io_out[26]
port 155 nsew signal tristate
flabel metal3 s 583520 13364 584800 13476 0 FreeSans 1120 0 0 0 io_out[2]
port 156 nsew signal tristate
flabel metal3 s 583520 18092 584800 18204 0 FreeSans 1120 0 0 0 io_out[3]
port 157 nsew signal tristate
flabel metal3 s 583520 22820 584800 22932 0 FreeSans 1120 0 0 0 io_out[4]
port 158 nsew signal tristate
flabel metal3 s 583520 49278 584800 49390 0 FreeSans 1120 0 0 0 io_out[5]
port 159 nsew signal tristate
flabel metal3 s 583520 93936 584800 94048 0 FreeSans 1120 0 0 0 io_out[6]
port 160 nsew signal tristate
flabel metal3 s 583520 273958 584800 274070 0 FreeSans 1120 0 0 0 io_out[7]
port 161 nsew signal tristate
flabel metal3 s 583520 318380 584800 318492 0 FreeSans 1120 0 0 0 io_out[8]
port 162 nsew signal tristate
flabel metal3 s 583520 363602 584800 363714 0 FreeSans 1120 0 0 0 io_out[9]
port 163 nsew signal tristate
flabel metal2 s 125816 -800 125928 480 0 FreeSans 1120 90 0 0 la_data_in[0]
port 164 nsew signal input
flabel metal2 s 480416 -800 480528 480 0 FreeSans 1120 90 0 0 la_data_in[100]
port 165 nsew signal input
flabel metal2 s 483962 -800 484074 480 0 FreeSans 1120 90 0 0 la_data_in[101]
port 166 nsew signal input
flabel metal2 s 487508 -800 487620 480 0 FreeSans 1120 90 0 0 la_data_in[102]
port 167 nsew signal input
flabel metal2 s 491054 -800 491166 480 0 FreeSans 1120 90 0 0 la_data_in[103]
port 168 nsew signal input
flabel metal2 s 494600 -800 494712 480 0 FreeSans 1120 90 0 0 la_data_in[104]
port 169 nsew signal input
flabel metal2 s 498146 -800 498258 480 0 FreeSans 1120 90 0 0 la_data_in[105]
port 170 nsew signal input
flabel metal2 s 501692 -800 501804 480 0 FreeSans 1120 90 0 0 la_data_in[106]
port 171 nsew signal input
flabel metal2 s 505238 -800 505350 480 0 FreeSans 1120 90 0 0 la_data_in[107]
port 172 nsew signal input
flabel metal2 s 508784 -800 508896 480 0 FreeSans 1120 90 0 0 la_data_in[108]
port 173 nsew signal input
flabel metal2 s 512330 -800 512442 480 0 FreeSans 1120 90 0 0 la_data_in[109]
port 174 nsew signal input
flabel metal2 s 161276 -800 161388 480 0 FreeSans 1120 90 0 0 la_data_in[10]
port 175 nsew signal input
flabel metal2 s 515876 -800 515988 480 0 FreeSans 1120 90 0 0 la_data_in[110]
port 176 nsew signal input
flabel metal2 s 519422 -800 519534 480 0 FreeSans 1120 90 0 0 la_data_in[111]
port 177 nsew signal input
flabel metal2 s 522968 -800 523080 480 0 FreeSans 1120 90 0 0 la_data_in[112]
port 178 nsew signal input
flabel metal2 s 526514 -800 526626 480 0 FreeSans 1120 90 0 0 la_data_in[113]
port 179 nsew signal input
flabel metal2 s 530060 -800 530172 480 0 FreeSans 1120 90 0 0 la_data_in[114]
port 180 nsew signal input
flabel metal2 s 533606 -800 533718 480 0 FreeSans 1120 90 0 0 la_data_in[115]
port 181 nsew signal input
flabel metal2 s 537152 -800 537264 480 0 FreeSans 1120 90 0 0 la_data_in[116]
port 182 nsew signal input
flabel metal2 s 540698 -800 540810 480 0 FreeSans 1120 90 0 0 la_data_in[117]
port 183 nsew signal input
flabel metal2 s 544244 -800 544356 480 0 FreeSans 1120 90 0 0 la_data_in[118]
port 184 nsew signal input
flabel metal2 s 547790 -800 547902 480 0 FreeSans 1120 90 0 0 la_data_in[119]
port 185 nsew signal input
flabel metal2 s 164822 -800 164934 480 0 FreeSans 1120 90 0 0 la_data_in[11]
port 186 nsew signal input
flabel metal2 s 551336 -800 551448 480 0 FreeSans 1120 90 0 0 la_data_in[120]
port 187 nsew signal input
flabel metal2 s 554882 -800 554994 480 0 FreeSans 1120 90 0 0 la_data_in[121]
port 188 nsew signal input
flabel metal2 s 558428 -800 558540 480 0 FreeSans 1120 90 0 0 la_data_in[122]
port 189 nsew signal input
flabel metal2 s 561974 -800 562086 480 0 FreeSans 1120 90 0 0 la_data_in[123]
port 190 nsew signal input
flabel metal2 s 565520 -800 565632 480 0 FreeSans 1120 90 0 0 la_data_in[124]
port 191 nsew signal input
flabel metal2 s 569066 -800 569178 480 0 FreeSans 1120 90 0 0 la_data_in[125]
port 192 nsew signal input
flabel metal2 s 572612 -800 572724 480 0 FreeSans 1120 90 0 0 la_data_in[126]
port 193 nsew signal input
flabel metal2 s 576158 -800 576270 480 0 FreeSans 1120 90 0 0 la_data_in[127]
port 194 nsew signal input
flabel metal2 s 168368 -800 168480 480 0 FreeSans 1120 90 0 0 la_data_in[12]
port 195 nsew signal input
flabel metal2 s 171914 -800 172026 480 0 FreeSans 1120 90 0 0 la_data_in[13]
port 196 nsew signal input
flabel metal2 s 175460 -800 175572 480 0 FreeSans 1120 90 0 0 la_data_in[14]
port 197 nsew signal input
flabel metal2 s 179006 -800 179118 480 0 FreeSans 1120 90 0 0 la_data_in[15]
port 198 nsew signal input
flabel metal2 s 182552 -800 182664 480 0 FreeSans 1120 90 0 0 la_data_in[16]
port 199 nsew signal input
flabel metal2 s 186098 -800 186210 480 0 FreeSans 1120 90 0 0 la_data_in[17]
port 200 nsew signal input
flabel metal2 s 189644 -800 189756 480 0 FreeSans 1120 90 0 0 la_data_in[18]
port 201 nsew signal input
flabel metal2 s 193190 -800 193302 480 0 FreeSans 1120 90 0 0 la_data_in[19]
port 202 nsew signal input
flabel metal2 s 129362 -800 129474 480 0 FreeSans 1120 90 0 0 la_data_in[1]
port 203 nsew signal input
flabel metal2 s 196736 -800 196848 480 0 FreeSans 1120 90 0 0 la_data_in[20]
port 204 nsew signal input
flabel metal2 s 200282 -800 200394 480 0 FreeSans 1120 90 0 0 la_data_in[21]
port 205 nsew signal input
flabel metal2 s 203828 -800 203940 480 0 FreeSans 1120 90 0 0 la_data_in[22]
port 206 nsew signal input
flabel metal2 s 207374 -800 207486 480 0 FreeSans 1120 90 0 0 la_data_in[23]
port 207 nsew signal input
flabel metal2 s 210920 -800 211032 480 0 FreeSans 1120 90 0 0 la_data_in[24]
port 208 nsew signal input
flabel metal2 s 214466 -800 214578 480 0 FreeSans 1120 90 0 0 la_data_in[25]
port 209 nsew signal input
flabel metal2 s 218012 -800 218124 480 0 FreeSans 1120 90 0 0 la_data_in[26]
port 210 nsew signal input
flabel metal2 s 221558 -800 221670 480 0 FreeSans 1120 90 0 0 la_data_in[27]
port 211 nsew signal input
flabel metal2 s 225104 -800 225216 480 0 FreeSans 1120 90 0 0 la_data_in[28]
port 212 nsew signal input
flabel metal2 s 228650 -800 228762 480 0 FreeSans 1120 90 0 0 la_data_in[29]
port 213 nsew signal input
flabel metal2 s 132908 -800 133020 480 0 FreeSans 1120 90 0 0 la_data_in[2]
port 214 nsew signal input
flabel metal2 s 232196 -800 232308 480 0 FreeSans 1120 90 0 0 la_data_in[30]
port 215 nsew signal input
flabel metal2 s 235742 -800 235854 480 0 FreeSans 1120 90 0 0 la_data_in[31]
port 216 nsew signal input
flabel metal2 s 239288 -800 239400 480 0 FreeSans 1120 90 0 0 la_data_in[32]
port 217 nsew signal input
flabel metal2 s 242834 -800 242946 480 0 FreeSans 1120 90 0 0 la_data_in[33]
port 218 nsew signal input
flabel metal2 s 246380 -800 246492 480 0 FreeSans 1120 90 0 0 la_data_in[34]
port 219 nsew signal input
flabel metal2 s 249926 -800 250038 480 0 FreeSans 1120 90 0 0 la_data_in[35]
port 220 nsew signal input
flabel metal2 s 253472 -800 253584 480 0 FreeSans 1120 90 0 0 la_data_in[36]
port 221 nsew signal input
flabel metal2 s 257018 -800 257130 480 0 FreeSans 1120 90 0 0 la_data_in[37]
port 222 nsew signal input
flabel metal2 s 260564 -800 260676 480 0 FreeSans 1120 90 0 0 la_data_in[38]
port 223 nsew signal input
flabel metal2 s 264110 -800 264222 480 0 FreeSans 1120 90 0 0 la_data_in[39]
port 224 nsew signal input
flabel metal2 s 136454 -800 136566 480 0 FreeSans 1120 90 0 0 la_data_in[3]
port 225 nsew signal input
flabel metal2 s 267656 -800 267768 480 0 FreeSans 1120 90 0 0 la_data_in[40]
port 226 nsew signal input
flabel metal2 s 271202 -800 271314 480 0 FreeSans 1120 90 0 0 la_data_in[41]
port 227 nsew signal input
flabel metal2 s 274748 -800 274860 480 0 FreeSans 1120 90 0 0 la_data_in[42]
port 228 nsew signal input
flabel metal2 s 278294 -800 278406 480 0 FreeSans 1120 90 0 0 la_data_in[43]
port 229 nsew signal input
flabel metal2 s 281840 -800 281952 480 0 FreeSans 1120 90 0 0 la_data_in[44]
port 230 nsew signal input
flabel metal2 s 285386 -800 285498 480 0 FreeSans 1120 90 0 0 la_data_in[45]
port 231 nsew signal input
flabel metal2 s 288932 -800 289044 480 0 FreeSans 1120 90 0 0 la_data_in[46]
port 232 nsew signal input
flabel metal2 s 292478 -800 292590 480 0 FreeSans 1120 90 0 0 la_data_in[47]
port 233 nsew signal input
flabel metal2 s 296024 -800 296136 480 0 FreeSans 1120 90 0 0 la_data_in[48]
port 234 nsew signal input
flabel metal2 s 299570 -800 299682 480 0 FreeSans 1120 90 0 0 la_data_in[49]
port 235 nsew signal input
flabel metal2 s 140000 -800 140112 480 0 FreeSans 1120 90 0 0 la_data_in[4]
port 236 nsew signal input
flabel metal2 s 303116 -800 303228 480 0 FreeSans 1120 90 0 0 la_data_in[50]
port 237 nsew signal input
flabel metal2 s 306662 -800 306774 480 0 FreeSans 1120 90 0 0 la_data_in[51]
port 238 nsew signal input
flabel metal2 s 310208 -800 310320 480 0 FreeSans 1120 90 0 0 la_data_in[52]
port 239 nsew signal input
flabel metal2 s 313754 -800 313866 480 0 FreeSans 1120 90 0 0 la_data_in[53]
port 240 nsew signal input
flabel metal2 s 317300 -800 317412 480 0 FreeSans 1120 90 0 0 la_data_in[54]
port 241 nsew signal input
flabel metal2 s 320846 -800 320958 480 0 FreeSans 1120 90 0 0 la_data_in[55]
port 242 nsew signal input
flabel metal2 s 324392 -800 324504 480 0 FreeSans 1120 90 0 0 la_data_in[56]
port 243 nsew signal input
flabel metal2 s 327938 -800 328050 480 0 FreeSans 1120 90 0 0 la_data_in[57]
port 244 nsew signal input
flabel metal2 s 331484 -800 331596 480 0 FreeSans 1120 90 0 0 la_data_in[58]
port 245 nsew signal input
flabel metal2 s 335030 -800 335142 480 0 FreeSans 1120 90 0 0 la_data_in[59]
port 246 nsew signal input
flabel metal2 s 143546 -800 143658 480 0 FreeSans 1120 90 0 0 la_data_in[5]
port 247 nsew signal input
flabel metal2 s 338576 -800 338688 480 0 FreeSans 1120 90 0 0 la_data_in[60]
port 248 nsew signal input
flabel metal2 s 342122 -800 342234 480 0 FreeSans 1120 90 0 0 la_data_in[61]
port 249 nsew signal input
flabel metal2 s 345668 -800 345780 480 0 FreeSans 1120 90 0 0 la_data_in[62]
port 250 nsew signal input
flabel metal2 s 349214 -800 349326 480 0 FreeSans 1120 90 0 0 la_data_in[63]
port 251 nsew signal input
flabel metal2 s 352760 -800 352872 480 0 FreeSans 1120 90 0 0 la_data_in[64]
port 252 nsew signal input
flabel metal2 s 356306 -800 356418 480 0 FreeSans 1120 90 0 0 la_data_in[65]
port 253 nsew signal input
flabel metal2 s 359852 -800 359964 480 0 FreeSans 1120 90 0 0 la_data_in[66]
port 254 nsew signal input
flabel metal2 s 363398 -800 363510 480 0 FreeSans 1120 90 0 0 la_data_in[67]
port 255 nsew signal input
flabel metal2 s 366944 -800 367056 480 0 FreeSans 1120 90 0 0 la_data_in[68]
port 256 nsew signal input
flabel metal2 s 370490 -800 370602 480 0 FreeSans 1120 90 0 0 la_data_in[69]
port 257 nsew signal input
flabel metal2 s 147092 -800 147204 480 0 FreeSans 1120 90 0 0 la_data_in[6]
port 258 nsew signal input
flabel metal2 s 374036 -800 374148 480 0 FreeSans 1120 90 0 0 la_data_in[70]
port 259 nsew signal input
flabel metal2 s 377582 -800 377694 480 0 FreeSans 1120 90 0 0 la_data_in[71]
port 260 nsew signal input
flabel metal2 s 381128 -800 381240 480 0 FreeSans 1120 90 0 0 la_data_in[72]
port 261 nsew signal input
flabel metal2 s 384674 -800 384786 480 0 FreeSans 1120 90 0 0 la_data_in[73]
port 262 nsew signal input
flabel metal2 s 388220 -800 388332 480 0 FreeSans 1120 90 0 0 la_data_in[74]
port 263 nsew signal input
flabel metal2 s 391766 -800 391878 480 0 FreeSans 1120 90 0 0 la_data_in[75]
port 264 nsew signal input
flabel metal2 s 395312 -800 395424 480 0 FreeSans 1120 90 0 0 la_data_in[76]
port 265 nsew signal input
flabel metal2 s 398858 -800 398970 480 0 FreeSans 1120 90 0 0 la_data_in[77]
port 266 nsew signal input
flabel metal2 s 402404 -800 402516 480 0 FreeSans 1120 90 0 0 la_data_in[78]
port 267 nsew signal input
flabel metal2 s 405950 -800 406062 480 0 FreeSans 1120 90 0 0 la_data_in[79]
port 268 nsew signal input
flabel metal2 s 150638 -800 150750 480 0 FreeSans 1120 90 0 0 la_data_in[7]
port 269 nsew signal input
flabel metal2 s 409496 -800 409608 480 0 FreeSans 1120 90 0 0 la_data_in[80]
port 270 nsew signal input
flabel metal2 s 413042 -800 413154 480 0 FreeSans 1120 90 0 0 la_data_in[81]
port 271 nsew signal input
flabel metal2 s 416588 -800 416700 480 0 FreeSans 1120 90 0 0 la_data_in[82]
port 272 nsew signal input
flabel metal2 s 420134 -800 420246 480 0 FreeSans 1120 90 0 0 la_data_in[83]
port 273 nsew signal input
flabel metal2 s 423680 -800 423792 480 0 FreeSans 1120 90 0 0 la_data_in[84]
port 274 nsew signal input
flabel metal2 s 427226 -800 427338 480 0 FreeSans 1120 90 0 0 la_data_in[85]
port 275 nsew signal input
flabel metal2 s 430772 -800 430884 480 0 FreeSans 1120 90 0 0 la_data_in[86]
port 276 nsew signal input
flabel metal2 s 434318 -800 434430 480 0 FreeSans 1120 90 0 0 la_data_in[87]
port 277 nsew signal input
flabel metal2 s 437864 -800 437976 480 0 FreeSans 1120 90 0 0 la_data_in[88]
port 278 nsew signal input
flabel metal2 s 441410 -800 441522 480 0 FreeSans 1120 90 0 0 la_data_in[89]
port 279 nsew signal input
flabel metal2 s 154184 -800 154296 480 0 FreeSans 1120 90 0 0 la_data_in[8]
port 280 nsew signal input
flabel metal2 s 444956 -800 445068 480 0 FreeSans 1120 90 0 0 la_data_in[90]
port 281 nsew signal input
flabel metal2 s 448502 -800 448614 480 0 FreeSans 1120 90 0 0 la_data_in[91]
port 282 nsew signal input
flabel metal2 s 452048 -800 452160 480 0 FreeSans 1120 90 0 0 la_data_in[92]
port 283 nsew signal input
flabel metal2 s 455594 -800 455706 480 0 FreeSans 1120 90 0 0 la_data_in[93]
port 284 nsew signal input
flabel metal2 s 459140 -800 459252 480 0 FreeSans 1120 90 0 0 la_data_in[94]
port 285 nsew signal input
flabel metal2 s 462686 -800 462798 480 0 FreeSans 1120 90 0 0 la_data_in[95]
port 286 nsew signal input
flabel metal2 s 466232 -800 466344 480 0 FreeSans 1120 90 0 0 la_data_in[96]
port 287 nsew signal input
flabel metal2 s 469778 -800 469890 480 0 FreeSans 1120 90 0 0 la_data_in[97]
port 288 nsew signal input
flabel metal2 s 473324 -800 473436 480 0 FreeSans 1120 90 0 0 la_data_in[98]
port 289 nsew signal input
flabel metal2 s 476870 -800 476982 480 0 FreeSans 1120 90 0 0 la_data_in[99]
port 290 nsew signal input
flabel metal2 s 157730 -800 157842 480 0 FreeSans 1120 90 0 0 la_data_in[9]
port 291 nsew signal input
flabel metal2 s 126998 -800 127110 480 0 FreeSans 1120 90 0 0 la_data_out[0]
port 292 nsew signal tristate
flabel metal2 s 481598 -800 481710 480 0 FreeSans 1120 90 0 0 la_data_out[100]
port 293 nsew signal tristate
flabel metal2 s 485144 -800 485256 480 0 FreeSans 1120 90 0 0 la_data_out[101]
port 294 nsew signal tristate
flabel metal2 s 488690 -800 488802 480 0 FreeSans 1120 90 0 0 la_data_out[102]
port 295 nsew signal tristate
flabel metal2 s 492236 -800 492348 480 0 FreeSans 1120 90 0 0 la_data_out[103]
port 296 nsew signal tristate
flabel metal2 s 495782 -800 495894 480 0 FreeSans 1120 90 0 0 la_data_out[104]
port 297 nsew signal tristate
flabel metal2 s 499328 -800 499440 480 0 FreeSans 1120 90 0 0 la_data_out[105]
port 298 nsew signal tristate
flabel metal2 s 502874 -800 502986 480 0 FreeSans 1120 90 0 0 la_data_out[106]
port 299 nsew signal tristate
flabel metal2 s 506420 -800 506532 480 0 FreeSans 1120 90 0 0 la_data_out[107]
port 300 nsew signal tristate
flabel metal2 s 509966 -800 510078 480 0 FreeSans 1120 90 0 0 la_data_out[108]
port 301 nsew signal tristate
flabel metal2 s 513512 -800 513624 480 0 FreeSans 1120 90 0 0 la_data_out[109]
port 302 nsew signal tristate
flabel metal2 s 162458 -800 162570 480 0 FreeSans 1120 90 0 0 la_data_out[10]
port 303 nsew signal tristate
flabel metal2 s 517058 -800 517170 480 0 FreeSans 1120 90 0 0 la_data_out[110]
port 304 nsew signal tristate
flabel metal2 s 520604 -800 520716 480 0 FreeSans 1120 90 0 0 la_data_out[111]
port 305 nsew signal tristate
flabel metal2 s 524150 -800 524262 480 0 FreeSans 1120 90 0 0 la_data_out[112]
port 306 nsew signal tristate
flabel metal2 s 527696 -800 527808 480 0 FreeSans 1120 90 0 0 la_data_out[113]
port 307 nsew signal tristate
flabel metal2 s 531242 -800 531354 480 0 FreeSans 1120 90 0 0 la_data_out[114]
port 308 nsew signal tristate
flabel metal2 s 534788 -800 534900 480 0 FreeSans 1120 90 0 0 la_data_out[115]
port 309 nsew signal tristate
flabel metal2 s 538334 -800 538446 480 0 FreeSans 1120 90 0 0 la_data_out[116]
port 310 nsew signal tristate
flabel metal2 s 541880 -800 541992 480 0 FreeSans 1120 90 0 0 la_data_out[117]
port 311 nsew signal tristate
flabel metal2 s 545426 -800 545538 480 0 FreeSans 1120 90 0 0 la_data_out[118]
port 312 nsew signal tristate
flabel metal2 s 548972 -800 549084 480 0 FreeSans 1120 90 0 0 la_data_out[119]
port 313 nsew signal tristate
flabel metal2 s 166004 -800 166116 480 0 FreeSans 1120 90 0 0 la_data_out[11]
port 314 nsew signal tristate
flabel metal2 s 552518 -800 552630 480 0 FreeSans 1120 90 0 0 la_data_out[120]
port 315 nsew signal tristate
flabel metal2 s 556064 -800 556176 480 0 FreeSans 1120 90 0 0 la_data_out[121]
port 316 nsew signal tristate
flabel metal2 s 559610 -800 559722 480 0 FreeSans 1120 90 0 0 la_data_out[122]
port 317 nsew signal tristate
flabel metal2 s 563156 -800 563268 480 0 FreeSans 1120 90 0 0 la_data_out[123]
port 318 nsew signal tristate
flabel metal2 s 566702 -800 566814 480 0 FreeSans 1120 90 0 0 la_data_out[124]
port 319 nsew signal tristate
flabel metal2 s 570248 -800 570360 480 0 FreeSans 1120 90 0 0 la_data_out[125]
port 320 nsew signal tristate
flabel metal2 s 573794 -800 573906 480 0 FreeSans 1120 90 0 0 la_data_out[126]
port 321 nsew signal tristate
flabel metal2 s 577340 -800 577452 480 0 FreeSans 1120 90 0 0 la_data_out[127]
port 322 nsew signal tristate
flabel metal2 s 169550 -800 169662 480 0 FreeSans 1120 90 0 0 la_data_out[12]
port 323 nsew signal tristate
flabel metal2 s 173096 -800 173208 480 0 FreeSans 1120 90 0 0 la_data_out[13]
port 324 nsew signal tristate
flabel metal2 s 176642 -800 176754 480 0 FreeSans 1120 90 0 0 la_data_out[14]
port 325 nsew signal tristate
flabel metal2 s 180188 -800 180300 480 0 FreeSans 1120 90 0 0 la_data_out[15]
port 326 nsew signal tristate
flabel metal2 s 183734 -800 183846 480 0 FreeSans 1120 90 0 0 la_data_out[16]
port 327 nsew signal tristate
flabel metal2 s 187280 -800 187392 480 0 FreeSans 1120 90 0 0 la_data_out[17]
port 328 nsew signal tristate
flabel metal2 s 190826 -800 190938 480 0 FreeSans 1120 90 0 0 la_data_out[18]
port 329 nsew signal tristate
flabel metal2 s 194372 -800 194484 480 0 FreeSans 1120 90 0 0 la_data_out[19]
port 330 nsew signal tristate
flabel metal2 s 130544 -800 130656 480 0 FreeSans 1120 90 0 0 la_data_out[1]
port 331 nsew signal tristate
flabel metal2 s 197918 -800 198030 480 0 FreeSans 1120 90 0 0 la_data_out[20]
port 332 nsew signal tristate
flabel metal2 s 201464 -800 201576 480 0 FreeSans 1120 90 0 0 la_data_out[21]
port 333 nsew signal tristate
flabel metal2 s 205010 -800 205122 480 0 FreeSans 1120 90 0 0 la_data_out[22]
port 334 nsew signal tristate
flabel metal2 s 208556 -800 208668 480 0 FreeSans 1120 90 0 0 la_data_out[23]
port 335 nsew signal tristate
flabel metal2 s 212102 -800 212214 480 0 FreeSans 1120 90 0 0 la_data_out[24]
port 336 nsew signal tristate
flabel metal2 s 215648 -800 215760 480 0 FreeSans 1120 90 0 0 la_data_out[25]
port 337 nsew signal tristate
flabel metal2 s 219194 -800 219306 480 0 FreeSans 1120 90 0 0 la_data_out[26]
port 338 nsew signal tristate
flabel metal2 s 222740 -800 222852 480 0 FreeSans 1120 90 0 0 la_data_out[27]
port 339 nsew signal tristate
flabel metal2 s 226286 -800 226398 480 0 FreeSans 1120 90 0 0 la_data_out[28]
port 340 nsew signal tristate
flabel metal2 s 229832 -800 229944 480 0 FreeSans 1120 90 0 0 la_data_out[29]
port 341 nsew signal tristate
flabel metal2 s 134090 -800 134202 480 0 FreeSans 1120 90 0 0 la_data_out[2]
port 342 nsew signal tristate
flabel metal2 s 233378 -800 233490 480 0 FreeSans 1120 90 0 0 la_data_out[30]
port 343 nsew signal tristate
flabel metal2 s 236924 -800 237036 480 0 FreeSans 1120 90 0 0 la_data_out[31]
port 344 nsew signal tristate
flabel metal2 s 240470 -800 240582 480 0 FreeSans 1120 90 0 0 la_data_out[32]
port 345 nsew signal tristate
flabel metal2 s 244016 -800 244128 480 0 FreeSans 1120 90 0 0 la_data_out[33]
port 346 nsew signal tristate
flabel metal2 s 247562 -800 247674 480 0 FreeSans 1120 90 0 0 la_data_out[34]
port 347 nsew signal tristate
flabel metal2 s 251108 -800 251220 480 0 FreeSans 1120 90 0 0 la_data_out[35]
port 348 nsew signal tristate
flabel metal2 s 254654 -800 254766 480 0 FreeSans 1120 90 0 0 la_data_out[36]
port 349 nsew signal tristate
flabel metal2 s 258200 -800 258312 480 0 FreeSans 1120 90 0 0 la_data_out[37]
port 350 nsew signal tristate
flabel metal2 s 261746 -800 261858 480 0 FreeSans 1120 90 0 0 la_data_out[38]
port 351 nsew signal tristate
flabel metal2 s 265292 -800 265404 480 0 FreeSans 1120 90 0 0 la_data_out[39]
port 352 nsew signal tristate
flabel metal2 s 137636 -800 137748 480 0 FreeSans 1120 90 0 0 la_data_out[3]
port 353 nsew signal tristate
flabel metal2 s 268838 -800 268950 480 0 FreeSans 1120 90 0 0 la_data_out[40]
port 354 nsew signal tristate
flabel metal2 s 272384 -800 272496 480 0 FreeSans 1120 90 0 0 la_data_out[41]
port 355 nsew signal tristate
flabel metal2 s 275930 -800 276042 480 0 FreeSans 1120 90 0 0 la_data_out[42]
port 356 nsew signal tristate
flabel metal2 s 279476 -800 279588 480 0 FreeSans 1120 90 0 0 la_data_out[43]
port 357 nsew signal tristate
flabel metal2 s 283022 -800 283134 480 0 FreeSans 1120 90 0 0 la_data_out[44]
port 358 nsew signal tristate
flabel metal2 s 286568 -800 286680 480 0 FreeSans 1120 90 0 0 la_data_out[45]
port 359 nsew signal tristate
flabel metal2 s 290114 -800 290226 480 0 FreeSans 1120 90 0 0 la_data_out[46]
port 360 nsew signal tristate
flabel metal2 s 293660 -800 293772 480 0 FreeSans 1120 90 0 0 la_data_out[47]
port 361 nsew signal tristate
flabel metal2 s 297206 -800 297318 480 0 FreeSans 1120 90 0 0 la_data_out[48]
port 362 nsew signal tristate
flabel metal2 s 300752 -800 300864 480 0 FreeSans 1120 90 0 0 la_data_out[49]
port 363 nsew signal tristate
flabel metal2 s 141182 -800 141294 480 0 FreeSans 1120 90 0 0 la_data_out[4]
port 364 nsew signal tristate
flabel metal2 s 304298 -800 304410 480 0 FreeSans 1120 90 0 0 la_data_out[50]
port 365 nsew signal tristate
flabel metal2 s 307844 -800 307956 480 0 FreeSans 1120 90 0 0 la_data_out[51]
port 366 nsew signal tristate
flabel metal2 s 311390 -800 311502 480 0 FreeSans 1120 90 0 0 la_data_out[52]
port 367 nsew signal tristate
flabel metal2 s 314936 -800 315048 480 0 FreeSans 1120 90 0 0 la_data_out[53]
port 368 nsew signal tristate
flabel metal2 s 318482 -800 318594 480 0 FreeSans 1120 90 0 0 la_data_out[54]
port 369 nsew signal tristate
flabel metal2 s 322028 -800 322140 480 0 FreeSans 1120 90 0 0 la_data_out[55]
port 370 nsew signal tristate
flabel metal2 s 325574 -800 325686 480 0 FreeSans 1120 90 0 0 la_data_out[56]
port 371 nsew signal tristate
flabel metal2 s 329120 -800 329232 480 0 FreeSans 1120 90 0 0 la_data_out[57]
port 372 nsew signal tristate
flabel metal2 s 332666 -800 332778 480 0 FreeSans 1120 90 0 0 la_data_out[58]
port 373 nsew signal tristate
flabel metal2 s 336212 -800 336324 480 0 FreeSans 1120 90 0 0 la_data_out[59]
port 374 nsew signal tristate
flabel metal2 s 144728 -800 144840 480 0 FreeSans 1120 90 0 0 la_data_out[5]
port 375 nsew signal tristate
flabel metal2 s 339758 -800 339870 480 0 FreeSans 1120 90 0 0 la_data_out[60]
port 376 nsew signal tristate
flabel metal2 s 343304 -800 343416 480 0 FreeSans 1120 90 0 0 la_data_out[61]
port 377 nsew signal tristate
flabel metal2 s 346850 -800 346962 480 0 FreeSans 1120 90 0 0 la_data_out[62]
port 378 nsew signal tristate
flabel metal2 s 350396 -800 350508 480 0 FreeSans 1120 90 0 0 la_data_out[63]
port 379 nsew signal tristate
flabel metal2 s 353942 -800 354054 480 0 FreeSans 1120 90 0 0 la_data_out[64]
port 380 nsew signal tristate
flabel metal2 s 357488 -800 357600 480 0 FreeSans 1120 90 0 0 la_data_out[65]
port 381 nsew signal tristate
flabel metal2 s 361034 -800 361146 480 0 FreeSans 1120 90 0 0 la_data_out[66]
port 382 nsew signal tristate
flabel metal2 s 364580 -800 364692 480 0 FreeSans 1120 90 0 0 la_data_out[67]
port 383 nsew signal tristate
flabel metal2 s 368126 -800 368238 480 0 FreeSans 1120 90 0 0 la_data_out[68]
port 384 nsew signal tristate
flabel metal2 s 371672 -800 371784 480 0 FreeSans 1120 90 0 0 la_data_out[69]
port 385 nsew signal tristate
flabel metal2 s 148274 -800 148386 480 0 FreeSans 1120 90 0 0 la_data_out[6]
port 386 nsew signal tristate
flabel metal2 s 375218 -800 375330 480 0 FreeSans 1120 90 0 0 la_data_out[70]
port 387 nsew signal tristate
flabel metal2 s 378764 -800 378876 480 0 FreeSans 1120 90 0 0 la_data_out[71]
port 388 nsew signal tristate
flabel metal2 s 382310 -800 382422 480 0 FreeSans 1120 90 0 0 la_data_out[72]
port 389 nsew signal tristate
flabel metal2 s 385856 -800 385968 480 0 FreeSans 1120 90 0 0 la_data_out[73]
port 390 nsew signal tristate
flabel metal2 s 389402 -800 389514 480 0 FreeSans 1120 90 0 0 la_data_out[74]
port 391 nsew signal tristate
flabel metal2 s 392948 -800 393060 480 0 FreeSans 1120 90 0 0 la_data_out[75]
port 392 nsew signal tristate
flabel metal2 s 396494 -800 396606 480 0 FreeSans 1120 90 0 0 la_data_out[76]
port 393 nsew signal tristate
flabel metal2 s 400040 -800 400152 480 0 FreeSans 1120 90 0 0 la_data_out[77]
port 394 nsew signal tristate
flabel metal2 s 403586 -800 403698 480 0 FreeSans 1120 90 0 0 la_data_out[78]
port 395 nsew signal tristate
flabel metal2 s 407132 -800 407244 480 0 FreeSans 1120 90 0 0 la_data_out[79]
port 396 nsew signal tristate
flabel metal2 s 151820 -800 151932 480 0 FreeSans 1120 90 0 0 la_data_out[7]
port 397 nsew signal tristate
flabel metal2 s 410678 -800 410790 480 0 FreeSans 1120 90 0 0 la_data_out[80]
port 398 nsew signal tristate
flabel metal2 s 414224 -800 414336 480 0 FreeSans 1120 90 0 0 la_data_out[81]
port 399 nsew signal tristate
flabel metal2 s 417770 -800 417882 480 0 FreeSans 1120 90 0 0 la_data_out[82]
port 400 nsew signal tristate
flabel metal2 s 421316 -800 421428 480 0 FreeSans 1120 90 0 0 la_data_out[83]
port 401 nsew signal tristate
flabel metal2 s 424862 -800 424974 480 0 FreeSans 1120 90 0 0 la_data_out[84]
port 402 nsew signal tristate
flabel metal2 s 428408 -800 428520 480 0 FreeSans 1120 90 0 0 la_data_out[85]
port 403 nsew signal tristate
flabel metal2 s 431954 -800 432066 480 0 FreeSans 1120 90 0 0 la_data_out[86]
port 404 nsew signal tristate
flabel metal2 s 435500 -800 435612 480 0 FreeSans 1120 90 0 0 la_data_out[87]
port 405 nsew signal tristate
flabel metal2 s 439046 -800 439158 480 0 FreeSans 1120 90 0 0 la_data_out[88]
port 406 nsew signal tristate
flabel metal2 s 442592 -800 442704 480 0 FreeSans 1120 90 0 0 la_data_out[89]
port 407 nsew signal tristate
flabel metal2 s 155366 -800 155478 480 0 FreeSans 1120 90 0 0 la_data_out[8]
port 408 nsew signal tristate
flabel metal2 s 446138 -800 446250 480 0 FreeSans 1120 90 0 0 la_data_out[90]
port 409 nsew signal tristate
flabel metal2 s 449684 -800 449796 480 0 FreeSans 1120 90 0 0 la_data_out[91]
port 410 nsew signal tristate
flabel metal2 s 453230 -800 453342 480 0 FreeSans 1120 90 0 0 la_data_out[92]
port 411 nsew signal tristate
flabel metal2 s 456776 -800 456888 480 0 FreeSans 1120 90 0 0 la_data_out[93]
port 412 nsew signal tristate
flabel metal2 s 460322 -800 460434 480 0 FreeSans 1120 90 0 0 la_data_out[94]
port 413 nsew signal tristate
flabel metal2 s 463868 -800 463980 480 0 FreeSans 1120 90 0 0 la_data_out[95]
port 414 nsew signal tristate
flabel metal2 s 467414 -800 467526 480 0 FreeSans 1120 90 0 0 la_data_out[96]
port 415 nsew signal tristate
flabel metal2 s 470960 -800 471072 480 0 FreeSans 1120 90 0 0 la_data_out[97]
port 416 nsew signal tristate
flabel metal2 s 474506 -800 474618 480 0 FreeSans 1120 90 0 0 la_data_out[98]
port 417 nsew signal tristate
flabel metal2 s 478052 -800 478164 480 0 FreeSans 1120 90 0 0 la_data_out[99]
port 418 nsew signal tristate
flabel metal2 s 158912 -800 159024 480 0 FreeSans 1120 90 0 0 la_data_out[9]
port 419 nsew signal tristate
flabel metal2 s 128180 -800 128292 480 0 FreeSans 1120 90 0 0 la_oenb[0]
port 420 nsew signal input
flabel metal2 s 482780 -800 482892 480 0 FreeSans 1120 90 0 0 la_oenb[100]
port 421 nsew signal input
flabel metal2 s 486326 -800 486438 480 0 FreeSans 1120 90 0 0 la_oenb[101]
port 422 nsew signal input
flabel metal2 s 489872 -800 489984 480 0 FreeSans 1120 90 0 0 la_oenb[102]
port 423 nsew signal input
flabel metal2 s 493418 -800 493530 480 0 FreeSans 1120 90 0 0 la_oenb[103]
port 424 nsew signal input
flabel metal2 s 496964 -800 497076 480 0 FreeSans 1120 90 0 0 la_oenb[104]
port 425 nsew signal input
flabel metal2 s 500510 -800 500622 480 0 FreeSans 1120 90 0 0 la_oenb[105]
port 426 nsew signal input
flabel metal2 s 504056 -800 504168 480 0 FreeSans 1120 90 0 0 la_oenb[106]
port 427 nsew signal input
flabel metal2 s 507602 -800 507714 480 0 FreeSans 1120 90 0 0 la_oenb[107]
port 428 nsew signal input
flabel metal2 s 511148 -800 511260 480 0 FreeSans 1120 90 0 0 la_oenb[108]
port 429 nsew signal input
flabel metal2 s 514694 -800 514806 480 0 FreeSans 1120 90 0 0 la_oenb[109]
port 430 nsew signal input
flabel metal2 s 163640 -800 163752 480 0 FreeSans 1120 90 0 0 la_oenb[10]
port 431 nsew signal input
flabel metal2 s 518240 -800 518352 480 0 FreeSans 1120 90 0 0 la_oenb[110]
port 432 nsew signal input
flabel metal2 s 521786 -800 521898 480 0 FreeSans 1120 90 0 0 la_oenb[111]
port 433 nsew signal input
flabel metal2 s 525332 -800 525444 480 0 FreeSans 1120 90 0 0 la_oenb[112]
port 434 nsew signal input
flabel metal2 s 528878 -800 528990 480 0 FreeSans 1120 90 0 0 la_oenb[113]
port 435 nsew signal input
flabel metal2 s 532424 -800 532536 480 0 FreeSans 1120 90 0 0 la_oenb[114]
port 436 nsew signal input
flabel metal2 s 535970 -800 536082 480 0 FreeSans 1120 90 0 0 la_oenb[115]
port 437 nsew signal input
flabel metal2 s 539516 -800 539628 480 0 FreeSans 1120 90 0 0 la_oenb[116]
port 438 nsew signal input
flabel metal2 s 543062 -800 543174 480 0 FreeSans 1120 90 0 0 la_oenb[117]
port 439 nsew signal input
flabel metal2 s 546608 -800 546720 480 0 FreeSans 1120 90 0 0 la_oenb[118]
port 440 nsew signal input
flabel metal2 s 550154 -800 550266 480 0 FreeSans 1120 90 0 0 la_oenb[119]
port 441 nsew signal input
flabel metal2 s 167186 -800 167298 480 0 FreeSans 1120 90 0 0 la_oenb[11]
port 442 nsew signal input
flabel metal2 s 553700 -800 553812 480 0 FreeSans 1120 90 0 0 la_oenb[120]
port 443 nsew signal input
flabel metal2 s 557246 -800 557358 480 0 FreeSans 1120 90 0 0 la_oenb[121]
port 444 nsew signal input
flabel metal2 s 560792 -800 560904 480 0 FreeSans 1120 90 0 0 la_oenb[122]
port 445 nsew signal input
flabel metal2 s 564338 -800 564450 480 0 FreeSans 1120 90 0 0 la_oenb[123]
port 446 nsew signal input
flabel metal2 s 567884 -800 567996 480 0 FreeSans 1120 90 0 0 la_oenb[124]
port 447 nsew signal input
flabel metal2 s 571430 -800 571542 480 0 FreeSans 1120 90 0 0 la_oenb[125]
port 448 nsew signal input
flabel metal2 s 574976 -800 575088 480 0 FreeSans 1120 90 0 0 la_oenb[126]
port 449 nsew signal input
flabel metal2 s 578522 -800 578634 480 0 FreeSans 1120 90 0 0 la_oenb[127]
port 450 nsew signal input
flabel metal2 s 170732 -800 170844 480 0 FreeSans 1120 90 0 0 la_oenb[12]
port 451 nsew signal input
flabel metal2 s 174278 -800 174390 480 0 FreeSans 1120 90 0 0 la_oenb[13]
port 452 nsew signal input
flabel metal2 s 177824 -800 177936 480 0 FreeSans 1120 90 0 0 la_oenb[14]
port 453 nsew signal input
flabel metal2 s 181370 -800 181482 480 0 FreeSans 1120 90 0 0 la_oenb[15]
port 454 nsew signal input
flabel metal2 s 184916 -800 185028 480 0 FreeSans 1120 90 0 0 la_oenb[16]
port 455 nsew signal input
flabel metal2 s 188462 -800 188574 480 0 FreeSans 1120 90 0 0 la_oenb[17]
port 456 nsew signal input
flabel metal2 s 192008 -800 192120 480 0 FreeSans 1120 90 0 0 la_oenb[18]
port 457 nsew signal input
flabel metal2 s 195554 -800 195666 480 0 FreeSans 1120 90 0 0 la_oenb[19]
port 458 nsew signal input
flabel metal2 s 131726 -800 131838 480 0 FreeSans 1120 90 0 0 la_oenb[1]
port 459 nsew signal input
flabel metal2 s 199100 -800 199212 480 0 FreeSans 1120 90 0 0 la_oenb[20]
port 460 nsew signal input
flabel metal2 s 202646 -800 202758 480 0 FreeSans 1120 90 0 0 la_oenb[21]
port 461 nsew signal input
flabel metal2 s 206192 -800 206304 480 0 FreeSans 1120 90 0 0 la_oenb[22]
port 462 nsew signal input
flabel metal2 s 209738 -800 209850 480 0 FreeSans 1120 90 0 0 la_oenb[23]
port 463 nsew signal input
flabel metal2 s 213284 -800 213396 480 0 FreeSans 1120 90 0 0 la_oenb[24]
port 464 nsew signal input
flabel metal2 s 216830 -800 216942 480 0 FreeSans 1120 90 0 0 la_oenb[25]
port 465 nsew signal input
flabel metal2 s 220376 -800 220488 480 0 FreeSans 1120 90 0 0 la_oenb[26]
port 466 nsew signal input
flabel metal2 s 223922 -800 224034 480 0 FreeSans 1120 90 0 0 la_oenb[27]
port 467 nsew signal input
flabel metal2 s 227468 -800 227580 480 0 FreeSans 1120 90 0 0 la_oenb[28]
port 468 nsew signal input
flabel metal2 s 231014 -800 231126 480 0 FreeSans 1120 90 0 0 la_oenb[29]
port 469 nsew signal input
flabel metal2 s 135272 -800 135384 480 0 FreeSans 1120 90 0 0 la_oenb[2]
port 470 nsew signal input
flabel metal2 s 234560 -800 234672 480 0 FreeSans 1120 90 0 0 la_oenb[30]
port 471 nsew signal input
flabel metal2 s 238106 -800 238218 480 0 FreeSans 1120 90 0 0 la_oenb[31]
port 472 nsew signal input
flabel metal2 s 241652 -800 241764 480 0 FreeSans 1120 90 0 0 la_oenb[32]
port 473 nsew signal input
flabel metal2 s 245198 -800 245310 480 0 FreeSans 1120 90 0 0 la_oenb[33]
port 474 nsew signal input
flabel metal2 s 248744 -800 248856 480 0 FreeSans 1120 90 0 0 la_oenb[34]
port 475 nsew signal input
flabel metal2 s 252290 -800 252402 480 0 FreeSans 1120 90 0 0 la_oenb[35]
port 476 nsew signal input
flabel metal2 s 255836 -800 255948 480 0 FreeSans 1120 90 0 0 la_oenb[36]
port 477 nsew signal input
flabel metal2 s 259382 -800 259494 480 0 FreeSans 1120 90 0 0 la_oenb[37]
port 478 nsew signal input
flabel metal2 s 262928 -800 263040 480 0 FreeSans 1120 90 0 0 la_oenb[38]
port 479 nsew signal input
flabel metal2 s 266474 -800 266586 480 0 FreeSans 1120 90 0 0 la_oenb[39]
port 480 nsew signal input
flabel metal2 s 138818 -800 138930 480 0 FreeSans 1120 90 0 0 la_oenb[3]
port 481 nsew signal input
flabel metal2 s 270020 -800 270132 480 0 FreeSans 1120 90 0 0 la_oenb[40]
port 482 nsew signal input
flabel metal2 s 273566 -800 273678 480 0 FreeSans 1120 90 0 0 la_oenb[41]
port 483 nsew signal input
flabel metal2 s 277112 -800 277224 480 0 FreeSans 1120 90 0 0 la_oenb[42]
port 484 nsew signal input
flabel metal2 s 280658 -800 280770 480 0 FreeSans 1120 90 0 0 la_oenb[43]
port 485 nsew signal input
flabel metal2 s 284204 -800 284316 480 0 FreeSans 1120 90 0 0 la_oenb[44]
port 486 nsew signal input
flabel metal2 s 287750 -800 287862 480 0 FreeSans 1120 90 0 0 la_oenb[45]
port 487 nsew signal input
flabel metal2 s 291296 -800 291408 480 0 FreeSans 1120 90 0 0 la_oenb[46]
port 488 nsew signal input
flabel metal2 s 294842 -800 294954 480 0 FreeSans 1120 90 0 0 la_oenb[47]
port 489 nsew signal input
flabel metal2 s 298388 -800 298500 480 0 FreeSans 1120 90 0 0 la_oenb[48]
port 490 nsew signal input
flabel metal2 s 301934 -800 302046 480 0 FreeSans 1120 90 0 0 la_oenb[49]
port 491 nsew signal input
flabel metal2 s 142364 -800 142476 480 0 FreeSans 1120 90 0 0 la_oenb[4]
port 492 nsew signal input
flabel metal2 s 305480 -800 305592 480 0 FreeSans 1120 90 0 0 la_oenb[50]
port 493 nsew signal input
flabel metal2 s 309026 -800 309138 480 0 FreeSans 1120 90 0 0 la_oenb[51]
port 494 nsew signal input
flabel metal2 s 312572 -800 312684 480 0 FreeSans 1120 90 0 0 la_oenb[52]
port 495 nsew signal input
flabel metal2 s 316118 -800 316230 480 0 FreeSans 1120 90 0 0 la_oenb[53]
port 496 nsew signal input
flabel metal2 s 319664 -800 319776 480 0 FreeSans 1120 90 0 0 la_oenb[54]
port 497 nsew signal input
flabel metal2 s 323210 -800 323322 480 0 FreeSans 1120 90 0 0 la_oenb[55]
port 498 nsew signal input
flabel metal2 s 326756 -800 326868 480 0 FreeSans 1120 90 0 0 la_oenb[56]
port 499 nsew signal input
flabel metal2 s 330302 -800 330414 480 0 FreeSans 1120 90 0 0 la_oenb[57]
port 500 nsew signal input
flabel metal2 s 333848 -800 333960 480 0 FreeSans 1120 90 0 0 la_oenb[58]
port 501 nsew signal input
flabel metal2 s 337394 -800 337506 480 0 FreeSans 1120 90 0 0 la_oenb[59]
port 502 nsew signal input
flabel metal2 s 145910 -800 146022 480 0 FreeSans 1120 90 0 0 la_oenb[5]
port 503 nsew signal input
flabel metal2 s 340940 -800 341052 480 0 FreeSans 1120 90 0 0 la_oenb[60]
port 504 nsew signal input
flabel metal2 s 344486 -800 344598 480 0 FreeSans 1120 90 0 0 la_oenb[61]
port 505 nsew signal input
flabel metal2 s 348032 -800 348144 480 0 FreeSans 1120 90 0 0 la_oenb[62]
port 506 nsew signal input
flabel metal2 s 351578 -800 351690 480 0 FreeSans 1120 90 0 0 la_oenb[63]
port 507 nsew signal input
flabel metal2 s 355124 -800 355236 480 0 FreeSans 1120 90 0 0 la_oenb[64]
port 508 nsew signal input
flabel metal2 s 358670 -800 358782 480 0 FreeSans 1120 90 0 0 la_oenb[65]
port 509 nsew signal input
flabel metal2 s 362216 -800 362328 480 0 FreeSans 1120 90 0 0 la_oenb[66]
port 510 nsew signal input
flabel metal2 s 365762 -800 365874 480 0 FreeSans 1120 90 0 0 la_oenb[67]
port 511 nsew signal input
flabel metal2 s 369308 -800 369420 480 0 FreeSans 1120 90 0 0 la_oenb[68]
port 512 nsew signal input
flabel metal2 s 372854 -800 372966 480 0 FreeSans 1120 90 0 0 la_oenb[69]
port 513 nsew signal input
flabel metal2 s 149456 -800 149568 480 0 FreeSans 1120 90 0 0 la_oenb[6]
port 514 nsew signal input
flabel metal2 s 376400 -800 376512 480 0 FreeSans 1120 90 0 0 la_oenb[70]
port 515 nsew signal input
flabel metal2 s 379946 -800 380058 480 0 FreeSans 1120 90 0 0 la_oenb[71]
port 516 nsew signal input
flabel metal2 s 383492 -800 383604 480 0 FreeSans 1120 90 0 0 la_oenb[72]
port 517 nsew signal input
flabel metal2 s 387038 -800 387150 480 0 FreeSans 1120 90 0 0 la_oenb[73]
port 518 nsew signal input
flabel metal2 s 390584 -800 390696 480 0 FreeSans 1120 90 0 0 la_oenb[74]
port 519 nsew signal input
flabel metal2 s 394130 -800 394242 480 0 FreeSans 1120 90 0 0 la_oenb[75]
port 520 nsew signal input
flabel metal2 s 397676 -800 397788 480 0 FreeSans 1120 90 0 0 la_oenb[76]
port 521 nsew signal input
flabel metal2 s 401222 -800 401334 480 0 FreeSans 1120 90 0 0 la_oenb[77]
port 522 nsew signal input
flabel metal2 s 404768 -800 404880 480 0 FreeSans 1120 90 0 0 la_oenb[78]
port 523 nsew signal input
flabel metal2 s 408314 -800 408426 480 0 FreeSans 1120 90 0 0 la_oenb[79]
port 524 nsew signal input
flabel metal2 s 153002 -800 153114 480 0 FreeSans 1120 90 0 0 la_oenb[7]
port 525 nsew signal input
flabel metal2 s 411860 -800 411972 480 0 FreeSans 1120 90 0 0 la_oenb[80]
port 526 nsew signal input
flabel metal2 s 415406 -800 415518 480 0 FreeSans 1120 90 0 0 la_oenb[81]
port 527 nsew signal input
flabel metal2 s 418952 -800 419064 480 0 FreeSans 1120 90 0 0 la_oenb[82]
port 528 nsew signal input
flabel metal2 s 422498 -800 422610 480 0 FreeSans 1120 90 0 0 la_oenb[83]
port 529 nsew signal input
flabel metal2 s 426044 -800 426156 480 0 FreeSans 1120 90 0 0 la_oenb[84]
port 530 nsew signal input
flabel metal2 s 429590 -800 429702 480 0 FreeSans 1120 90 0 0 la_oenb[85]
port 531 nsew signal input
flabel metal2 s 433136 -800 433248 480 0 FreeSans 1120 90 0 0 la_oenb[86]
port 532 nsew signal input
flabel metal2 s 436682 -800 436794 480 0 FreeSans 1120 90 0 0 la_oenb[87]
port 533 nsew signal input
flabel metal2 s 440228 -800 440340 480 0 FreeSans 1120 90 0 0 la_oenb[88]
port 534 nsew signal input
flabel metal2 s 443774 -800 443886 480 0 FreeSans 1120 90 0 0 la_oenb[89]
port 535 nsew signal input
flabel metal2 s 156548 -800 156660 480 0 FreeSans 1120 90 0 0 la_oenb[8]
port 536 nsew signal input
flabel metal2 s 447320 -800 447432 480 0 FreeSans 1120 90 0 0 la_oenb[90]
port 537 nsew signal input
flabel metal2 s 450866 -800 450978 480 0 FreeSans 1120 90 0 0 la_oenb[91]
port 538 nsew signal input
flabel metal2 s 454412 -800 454524 480 0 FreeSans 1120 90 0 0 la_oenb[92]
port 539 nsew signal input
flabel metal2 s 457958 -800 458070 480 0 FreeSans 1120 90 0 0 la_oenb[93]
port 540 nsew signal input
flabel metal2 s 461504 -800 461616 480 0 FreeSans 1120 90 0 0 la_oenb[94]
port 541 nsew signal input
flabel metal2 s 465050 -800 465162 480 0 FreeSans 1120 90 0 0 la_oenb[95]
port 542 nsew signal input
flabel metal2 s 468596 -800 468708 480 0 FreeSans 1120 90 0 0 la_oenb[96]
port 543 nsew signal input
flabel metal2 s 472142 -800 472254 480 0 FreeSans 1120 90 0 0 la_oenb[97]
port 544 nsew signal input
flabel metal2 s 475688 -800 475800 480 0 FreeSans 1120 90 0 0 la_oenb[98]
port 545 nsew signal input
flabel metal2 s 479234 -800 479346 480 0 FreeSans 1120 90 0 0 la_oenb[99]
port 546 nsew signal input
flabel metal2 s 160094 -800 160206 480 0 FreeSans 1120 90 0 0 la_oenb[9]
port 547 nsew signal input
flabel metal2 s 579704 -800 579816 480 0 FreeSans 1120 90 0 0 user_clock2
port 548 nsew signal input
flabel metal2 s 580886 -800 580998 480 0 FreeSans 1120 90 0 0 user_irq[0]
port 549 nsew signal tristate
flabel metal2 s 582068 -800 582180 480 0 FreeSans 1120 90 0 0 user_irq[1]
port 550 nsew signal tristate
flabel metal2 s 583250 -800 583362 480 0 FreeSans 1120 90 0 0 user_irq[2]
port 551 nsew signal tristate
flabel metal3 s 582340 639784 584800 644584 0 FreeSans 1120 0 0 0 vccd1
port 552 nsew signal bidirectional
flabel metal3 s 582340 629784 584800 634584 0 FreeSans 1120 0 0 0 vccd1
port 553 nsew signal bidirectional
flabel metal3 s 0 643842 1660 648642 0 FreeSans 1120 0 0 0 vccd2
port 554 nsew signal bidirectional
flabel metal3 s 0 633842 1660 638642 0 FreeSans 1120 0 0 0 vccd2
port 555 nsew signal bidirectional
flabel metal3 s 582340 540562 584800 545362 0 FreeSans 1120 0 0 0 vdda1
port 556 nsew signal bidirectional
flabel metal3 s 582340 550562 584800 555362 0 FreeSans 1120 0 0 0 vdda1
port 557 nsew signal bidirectional
flabel metal3 s 582340 235230 584800 240030 0 FreeSans 1120 0 0 0 vdda1
port 558 nsew signal bidirectional
flabel metal3 s 582340 225230 584800 230030 0 FreeSans 1120 0 0 0 vdda1
port 559 nsew signal bidirectional
flabel metal3 s 0 204888 1660 209688 0 FreeSans 1120 0 0 0 vdda2
port 560 nsew signal bidirectional
flabel metal3 s 0 214888 1660 219688 0 FreeSans 1120 0 0 0 vdda2
port 561 nsew signal bidirectional
flabel metal3 s 520594 702340 525394 704800 0 FreeSans 1920 180 0 0 vssa1
port 562 nsew signal bidirectional
flabel metal3 s 510594 702340 515394 704800 0 FreeSans 1920 180 0 0 vssa1
port 563 nsew signal bidirectional
flabel metal3 s 582340 146830 584800 151630 0 FreeSans 1120 0 0 0 vssa1
port 564 nsew signal bidirectional
flabel metal3 s 582340 136830 584800 141630 0 FreeSans 1120 0 0 0 vssa1
port 565 nsew signal bidirectional
flabel metal3 s 0 559442 1660 564242 0 FreeSans 1120 0 0 0 vssa2
port 566 nsew signal bidirectional
flabel metal3 s 0 549442 1660 554242 0 FreeSans 1120 0 0 0 vssa2
port 567 nsew signal bidirectional
flabel metal3 s 582340 191430 584800 196230 0 FreeSans 1120 0 0 0 vssd1
port 568 nsew signal bidirectional
flabel metal3 s 582340 181430 584800 186230 0 FreeSans 1120 0 0 0 vssd1
port 569 nsew signal bidirectional
flabel metal3 s 0 172888 1660 177688 0 FreeSans 1120 0 0 0 vssd2
port 570 nsew signal bidirectional
flabel metal3 s 0 162888 1660 167688 0 FreeSans 1120 0 0 0 vssd2
port 571 nsew signal bidirectional
flabel metal2 s 524 -800 636 480 0 FreeSans 1120 90 0 0 wb_clk_i
port 572 nsew signal input
flabel metal2 s 1706 -800 1818 480 0 FreeSans 1120 90 0 0 wb_rst_i
port 573 nsew signal input
flabel metal2 s 2888 -800 3000 480 0 FreeSans 1120 90 0 0 wbs_ack_o
port 574 nsew signal tristate
flabel metal2 s 7616 -800 7728 480 0 FreeSans 1120 90 0 0 wbs_adr_i[0]
port 575 nsew signal input
flabel metal2 s 47804 -800 47916 480 0 FreeSans 1120 90 0 0 wbs_adr_i[10]
port 576 nsew signal input
flabel metal2 s 51350 -800 51462 480 0 FreeSans 1120 90 0 0 wbs_adr_i[11]
port 577 nsew signal input
flabel metal2 s 54896 -800 55008 480 0 FreeSans 1120 90 0 0 wbs_adr_i[12]
port 578 nsew signal input
flabel metal2 s 58442 -800 58554 480 0 FreeSans 1120 90 0 0 wbs_adr_i[13]
port 579 nsew signal input
flabel metal2 s 61988 -800 62100 480 0 FreeSans 1120 90 0 0 wbs_adr_i[14]
port 580 nsew signal input
flabel metal2 s 65534 -800 65646 480 0 FreeSans 1120 90 0 0 wbs_adr_i[15]
port 581 nsew signal input
flabel metal2 s 69080 -800 69192 480 0 FreeSans 1120 90 0 0 wbs_adr_i[16]
port 582 nsew signal input
flabel metal2 s 72626 -800 72738 480 0 FreeSans 1120 90 0 0 wbs_adr_i[17]
port 583 nsew signal input
flabel metal2 s 76172 -800 76284 480 0 FreeSans 1120 90 0 0 wbs_adr_i[18]
port 584 nsew signal input
flabel metal2 s 79718 -800 79830 480 0 FreeSans 1120 90 0 0 wbs_adr_i[19]
port 585 nsew signal input
flabel metal2 s 12344 -800 12456 480 0 FreeSans 1120 90 0 0 wbs_adr_i[1]
port 586 nsew signal input
flabel metal2 s 83264 -800 83376 480 0 FreeSans 1120 90 0 0 wbs_adr_i[20]
port 587 nsew signal input
flabel metal2 s 86810 -800 86922 480 0 FreeSans 1120 90 0 0 wbs_adr_i[21]
port 588 nsew signal input
flabel metal2 s 90356 -800 90468 480 0 FreeSans 1120 90 0 0 wbs_adr_i[22]
port 589 nsew signal input
flabel metal2 s 93902 -800 94014 480 0 FreeSans 1120 90 0 0 wbs_adr_i[23]
port 590 nsew signal input
flabel metal2 s 97448 -800 97560 480 0 FreeSans 1120 90 0 0 wbs_adr_i[24]
port 591 nsew signal input
flabel metal2 s 100994 -800 101106 480 0 FreeSans 1120 90 0 0 wbs_adr_i[25]
port 592 nsew signal input
flabel metal2 s 104540 -800 104652 480 0 FreeSans 1120 90 0 0 wbs_adr_i[26]
port 593 nsew signal input
flabel metal2 s 108086 -800 108198 480 0 FreeSans 1120 90 0 0 wbs_adr_i[27]
port 594 nsew signal input
flabel metal2 s 111632 -800 111744 480 0 FreeSans 1120 90 0 0 wbs_adr_i[28]
port 595 nsew signal input
flabel metal2 s 115178 -800 115290 480 0 FreeSans 1120 90 0 0 wbs_adr_i[29]
port 596 nsew signal input
flabel metal2 s 17072 -800 17184 480 0 FreeSans 1120 90 0 0 wbs_adr_i[2]
port 597 nsew signal input
flabel metal2 s 118724 -800 118836 480 0 FreeSans 1120 90 0 0 wbs_adr_i[30]
port 598 nsew signal input
flabel metal2 s 122270 -800 122382 480 0 FreeSans 1120 90 0 0 wbs_adr_i[31]
port 599 nsew signal input
flabel metal2 s 21800 -800 21912 480 0 FreeSans 1120 90 0 0 wbs_adr_i[3]
port 600 nsew signal input
flabel metal2 s 26528 -800 26640 480 0 FreeSans 1120 90 0 0 wbs_adr_i[4]
port 601 nsew signal input
flabel metal2 s 30074 -800 30186 480 0 FreeSans 1120 90 0 0 wbs_adr_i[5]
port 602 nsew signal input
flabel metal2 s 33620 -800 33732 480 0 FreeSans 1120 90 0 0 wbs_adr_i[6]
port 603 nsew signal input
flabel metal2 s 37166 -800 37278 480 0 FreeSans 1120 90 0 0 wbs_adr_i[7]
port 604 nsew signal input
flabel metal2 s 40712 -800 40824 480 0 FreeSans 1120 90 0 0 wbs_adr_i[8]
port 605 nsew signal input
flabel metal2 s 44258 -800 44370 480 0 FreeSans 1120 90 0 0 wbs_adr_i[9]
port 606 nsew signal input
flabel metal2 s 4070 -800 4182 480 0 FreeSans 1120 90 0 0 wbs_cyc_i
port 607 nsew signal input
flabel metal2 s 8798 -800 8910 480 0 FreeSans 1120 90 0 0 wbs_dat_i[0]
port 608 nsew signal input
flabel metal2 s 48986 -800 49098 480 0 FreeSans 1120 90 0 0 wbs_dat_i[10]
port 609 nsew signal input
flabel metal2 s 52532 -800 52644 480 0 FreeSans 1120 90 0 0 wbs_dat_i[11]
port 610 nsew signal input
flabel metal2 s 56078 -800 56190 480 0 FreeSans 1120 90 0 0 wbs_dat_i[12]
port 611 nsew signal input
flabel metal2 s 59624 -800 59736 480 0 FreeSans 1120 90 0 0 wbs_dat_i[13]
port 612 nsew signal input
flabel metal2 s 63170 -800 63282 480 0 FreeSans 1120 90 0 0 wbs_dat_i[14]
port 613 nsew signal input
flabel metal2 s 66716 -800 66828 480 0 FreeSans 1120 90 0 0 wbs_dat_i[15]
port 614 nsew signal input
flabel metal2 s 70262 -800 70374 480 0 FreeSans 1120 90 0 0 wbs_dat_i[16]
port 615 nsew signal input
flabel metal2 s 73808 -800 73920 480 0 FreeSans 1120 90 0 0 wbs_dat_i[17]
port 616 nsew signal input
flabel metal2 s 77354 -800 77466 480 0 FreeSans 1120 90 0 0 wbs_dat_i[18]
port 617 nsew signal input
flabel metal2 s 80900 -800 81012 480 0 FreeSans 1120 90 0 0 wbs_dat_i[19]
port 618 nsew signal input
flabel metal2 s 13526 -800 13638 480 0 FreeSans 1120 90 0 0 wbs_dat_i[1]
port 619 nsew signal input
flabel metal2 s 84446 -800 84558 480 0 FreeSans 1120 90 0 0 wbs_dat_i[20]
port 620 nsew signal input
flabel metal2 s 87992 -800 88104 480 0 FreeSans 1120 90 0 0 wbs_dat_i[21]
port 621 nsew signal input
flabel metal2 s 91538 -800 91650 480 0 FreeSans 1120 90 0 0 wbs_dat_i[22]
port 622 nsew signal input
flabel metal2 s 95084 -800 95196 480 0 FreeSans 1120 90 0 0 wbs_dat_i[23]
port 623 nsew signal input
flabel metal2 s 98630 -800 98742 480 0 FreeSans 1120 90 0 0 wbs_dat_i[24]
port 624 nsew signal input
flabel metal2 s 102176 -800 102288 480 0 FreeSans 1120 90 0 0 wbs_dat_i[25]
port 625 nsew signal input
flabel metal2 s 105722 -800 105834 480 0 FreeSans 1120 90 0 0 wbs_dat_i[26]
port 626 nsew signal input
flabel metal2 s 109268 -800 109380 480 0 FreeSans 1120 90 0 0 wbs_dat_i[27]
port 627 nsew signal input
flabel metal2 s 112814 -800 112926 480 0 FreeSans 1120 90 0 0 wbs_dat_i[28]
port 628 nsew signal input
flabel metal2 s 116360 -800 116472 480 0 FreeSans 1120 90 0 0 wbs_dat_i[29]
port 629 nsew signal input
flabel metal2 s 18254 -800 18366 480 0 FreeSans 1120 90 0 0 wbs_dat_i[2]
port 630 nsew signal input
flabel metal2 s 119906 -800 120018 480 0 FreeSans 1120 90 0 0 wbs_dat_i[30]
port 631 nsew signal input
flabel metal2 s 123452 -800 123564 480 0 FreeSans 1120 90 0 0 wbs_dat_i[31]
port 632 nsew signal input
flabel metal2 s 22982 -800 23094 480 0 FreeSans 1120 90 0 0 wbs_dat_i[3]
port 633 nsew signal input
flabel metal2 s 27710 -800 27822 480 0 FreeSans 1120 90 0 0 wbs_dat_i[4]
port 634 nsew signal input
flabel metal2 s 31256 -800 31368 480 0 FreeSans 1120 90 0 0 wbs_dat_i[5]
port 635 nsew signal input
flabel metal2 s 34802 -800 34914 480 0 FreeSans 1120 90 0 0 wbs_dat_i[6]
port 636 nsew signal input
flabel metal2 s 38348 -800 38460 480 0 FreeSans 1120 90 0 0 wbs_dat_i[7]
port 637 nsew signal input
flabel metal2 s 41894 -800 42006 480 0 FreeSans 1120 90 0 0 wbs_dat_i[8]
port 638 nsew signal input
flabel metal2 s 45440 -800 45552 480 0 FreeSans 1120 90 0 0 wbs_dat_i[9]
port 639 nsew signal input
flabel metal2 s 9980 -800 10092 480 0 FreeSans 1120 90 0 0 wbs_dat_o[0]
port 640 nsew signal tristate
flabel metal2 s 50168 -800 50280 480 0 FreeSans 1120 90 0 0 wbs_dat_o[10]
port 641 nsew signal tristate
flabel metal2 s 53714 -800 53826 480 0 FreeSans 1120 90 0 0 wbs_dat_o[11]
port 642 nsew signal tristate
flabel metal2 s 57260 -800 57372 480 0 FreeSans 1120 90 0 0 wbs_dat_o[12]
port 643 nsew signal tristate
flabel metal2 s 60806 -800 60918 480 0 FreeSans 1120 90 0 0 wbs_dat_o[13]
port 644 nsew signal tristate
flabel metal2 s 64352 -800 64464 480 0 FreeSans 1120 90 0 0 wbs_dat_o[14]
port 645 nsew signal tristate
flabel metal2 s 67898 -800 68010 480 0 FreeSans 1120 90 0 0 wbs_dat_o[15]
port 646 nsew signal tristate
flabel metal2 s 71444 -800 71556 480 0 FreeSans 1120 90 0 0 wbs_dat_o[16]
port 647 nsew signal tristate
flabel metal2 s 74990 -800 75102 480 0 FreeSans 1120 90 0 0 wbs_dat_o[17]
port 648 nsew signal tristate
flabel metal2 s 78536 -800 78648 480 0 FreeSans 1120 90 0 0 wbs_dat_o[18]
port 649 nsew signal tristate
flabel metal2 s 82082 -800 82194 480 0 FreeSans 1120 90 0 0 wbs_dat_o[19]
port 650 nsew signal tristate
flabel metal2 s 14708 -800 14820 480 0 FreeSans 1120 90 0 0 wbs_dat_o[1]
port 651 nsew signal tristate
flabel metal2 s 85628 -800 85740 480 0 FreeSans 1120 90 0 0 wbs_dat_o[20]
port 652 nsew signal tristate
flabel metal2 s 89174 -800 89286 480 0 FreeSans 1120 90 0 0 wbs_dat_o[21]
port 653 nsew signal tristate
flabel metal2 s 92720 -800 92832 480 0 FreeSans 1120 90 0 0 wbs_dat_o[22]
port 654 nsew signal tristate
flabel metal2 s 96266 -800 96378 480 0 FreeSans 1120 90 0 0 wbs_dat_o[23]
port 655 nsew signal tristate
flabel metal2 s 99812 -800 99924 480 0 FreeSans 1120 90 0 0 wbs_dat_o[24]
port 656 nsew signal tristate
flabel metal2 s 103358 -800 103470 480 0 FreeSans 1120 90 0 0 wbs_dat_o[25]
port 657 nsew signal tristate
flabel metal2 s 106904 -800 107016 480 0 FreeSans 1120 90 0 0 wbs_dat_o[26]
port 658 nsew signal tristate
flabel metal2 s 110450 -800 110562 480 0 FreeSans 1120 90 0 0 wbs_dat_o[27]
port 659 nsew signal tristate
flabel metal2 s 113996 -800 114108 480 0 FreeSans 1120 90 0 0 wbs_dat_o[28]
port 660 nsew signal tristate
flabel metal2 s 117542 -800 117654 480 0 FreeSans 1120 90 0 0 wbs_dat_o[29]
port 661 nsew signal tristate
flabel metal2 s 19436 -800 19548 480 0 FreeSans 1120 90 0 0 wbs_dat_o[2]
port 662 nsew signal tristate
flabel metal2 s 121088 -800 121200 480 0 FreeSans 1120 90 0 0 wbs_dat_o[30]
port 663 nsew signal tristate
flabel metal2 s 124634 -800 124746 480 0 FreeSans 1120 90 0 0 wbs_dat_o[31]
port 664 nsew signal tristate
flabel metal2 s 24164 -800 24276 480 0 FreeSans 1120 90 0 0 wbs_dat_o[3]
port 665 nsew signal tristate
flabel metal2 s 28892 -800 29004 480 0 FreeSans 1120 90 0 0 wbs_dat_o[4]
port 666 nsew signal tristate
flabel metal2 s 32438 -800 32550 480 0 FreeSans 1120 90 0 0 wbs_dat_o[5]
port 667 nsew signal tristate
flabel metal2 s 35984 -800 36096 480 0 FreeSans 1120 90 0 0 wbs_dat_o[6]
port 668 nsew signal tristate
flabel metal2 s 39530 -800 39642 480 0 FreeSans 1120 90 0 0 wbs_dat_o[7]
port 669 nsew signal tristate
flabel metal2 s 43076 -800 43188 480 0 FreeSans 1120 90 0 0 wbs_dat_o[8]
port 670 nsew signal tristate
flabel metal2 s 46622 -800 46734 480 0 FreeSans 1120 90 0 0 wbs_dat_o[9]
port 671 nsew signal tristate
flabel metal2 s 11162 -800 11274 480 0 FreeSans 1120 90 0 0 wbs_sel_i[0]
port 672 nsew signal input
flabel metal2 s 15890 -800 16002 480 0 FreeSans 1120 90 0 0 wbs_sel_i[1]
port 673 nsew signal input
flabel metal2 s 20618 -800 20730 480 0 FreeSans 1120 90 0 0 wbs_sel_i[2]
port 674 nsew signal input
flabel metal2 s 25346 -800 25458 480 0 FreeSans 1120 90 0 0 wbs_sel_i[3]
port 675 nsew signal input
flabel metal2 s 5252 -800 5364 480 0 FreeSans 1120 90 0 0 wbs_stb_i
port 676 nsew signal input
flabel metal2 s 6434 -800 6546 480 0 FreeSans 1120 90 0 0 wbs_we_i
port 677 nsew signal input
flabel metal4 s 318994 702300 323994 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 47 nsew signal bidirectional
flabel metal4 s 329294 702300 334294 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 41 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
