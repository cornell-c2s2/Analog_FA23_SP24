magic
tech sky130A
magscale 1 2
timestamp 1709399651
<< error_p >>
rect 19 1081 77 1087
rect 19 1047 31 1081
rect 19 1041 77 1047
rect -77 -1047 -19 -1041
rect -77 -1081 -65 -1047
rect -77 -1087 -19 -1081
<< nwell >>
rect -263 -1219 263 1219
<< pmos >>
rect -63 -1000 -33 1000
rect 33 -1000 63 1000
<< pdiff >>
rect -125 988 -63 1000
rect -125 -988 -113 988
rect -79 -988 -63 988
rect -125 -1000 -63 -988
rect -33 988 33 1000
rect -33 -988 -17 988
rect 17 -988 33 988
rect -33 -1000 33 -988
rect 63 988 125 1000
rect 63 -988 79 988
rect 113 -988 125 988
rect 63 -1000 125 -988
<< pdiffc >>
rect -113 -988 -79 988
rect -17 -988 17 988
rect 79 -988 113 988
<< nsubdiff >>
rect -227 1149 -131 1183
rect 131 1149 227 1183
rect -227 1087 -193 1149
rect 193 1087 227 1149
rect -227 -1149 -193 -1087
rect 193 -1149 227 -1087
rect -227 -1183 -131 -1149
rect 131 -1183 227 -1149
<< nsubdiffcont >>
rect -131 1149 131 1183
rect -227 -1087 -193 1087
rect 193 -1087 227 1087
rect -131 -1183 131 -1149
<< poly >>
rect 15 1081 81 1097
rect 15 1047 31 1081
rect 65 1047 81 1081
rect 15 1031 81 1047
rect -63 1000 -33 1026
rect 33 1000 63 1031
rect -63 -1031 -33 -1000
rect 33 -1026 63 -1000
rect -81 -1047 -15 -1031
rect -81 -1081 -65 -1047
rect -31 -1081 -15 -1047
rect -81 -1097 -15 -1081
<< polycont >>
rect 31 1047 65 1081
rect -65 -1081 -31 -1047
<< locali >>
rect -227 1149 -131 1183
rect 131 1149 227 1183
rect -227 1087 -193 1149
rect 193 1087 227 1149
rect 15 1047 31 1081
rect 65 1047 81 1081
rect -113 988 -79 1004
rect -113 -1004 -79 -988
rect -17 988 17 1004
rect -17 -1004 17 -988
rect 79 988 113 1004
rect 79 -1004 113 -988
rect -81 -1081 -65 -1047
rect -31 -1081 -15 -1047
rect -227 -1149 -193 -1087
rect 193 -1149 227 -1087
rect -227 -1183 -131 -1149
rect 131 -1183 227 -1149
<< viali >>
rect 31 1047 65 1081
rect -113 -988 -79 988
rect -17 -988 17 988
rect 79 -988 113 988
rect -65 -1081 -31 -1047
<< metal1 >>
rect 19 1081 77 1087
rect 19 1047 31 1081
rect 65 1047 77 1081
rect 19 1041 77 1047
rect -119 988 -73 1000
rect -119 -988 -113 988
rect -79 -988 -73 988
rect -119 -1000 -73 -988
rect -23 988 23 1000
rect -23 -988 -17 988
rect 17 -988 23 988
rect -23 -1000 23 -988
rect 73 988 119 1000
rect 73 -988 79 988
rect 113 -988 119 988
rect 73 -1000 119 -988
rect -77 -1047 -19 -1041
rect -77 -1081 -65 -1047
rect -31 -1081 -19 -1047
rect -77 -1087 -19 -1081
<< properties >>
string FIXED_BBOX -210 -1166 210 1166
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 10 l 0.15 m 1 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
