* NGSPICE file created from class_AB_v3_sym_flatten.ext - technology: sky130A

.subckt class_AB_v3_sym_flatten VDD VOP VON VIN VIP IB CLK VSS
X0 a_810_n2630# IB.t2 VSS.t15 VSS.t14 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1 w_1880_n1260# CLK.t0 VON.t2 VDD.t8 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X2 VIP.t0 w_1258_n1260# error sky130_fd_pr__cap_var_lvt w=2 l=0.18
X3 VSS.t13 IB.t0 IB.t1 VSS.t12 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X4 VOP.t3 CLK.t1 w_1258_n1260# VDD.t7 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X5 a_810_n2630# IB.t3 VSS.t11 VSS.t10 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X6 a_810_n2630# VIP.t1 w_1880_n1260# VSS.t4 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X7 VOP.t2 CLK.t2 VON.t3 VDD.t6 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X8 VDD.t4 CLK.t3 w_1880_n1260# VSS.t7 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X9 VDD.t5 CLK.t4 w_1258_n1260# VSS.t8 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X10 VSS.t3 CLK.t5 a_872_n982# VSS.t2 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X11 VOP.t1 VON.t4 a_872_n982# VSS.t5 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X12 VIN.t0 w_1880_n1260# error sky130_fd_pr__cap_var_lvt w=2 l=0.18
X13 VON.t0 VOP.t4 a_872_n982# VSS.t0 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X14 w_1258_n1260# VIN.t1 a_810_n2630# VSS.t9 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X15 VDD.t3 VOP.t5 VON.t1 VDD.t2 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X16 VOP.t0 VON.t5 VDD.t1 VDD.t0 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
R0 IB.t2 IB.t3 365.654
R1 IB.n0 IB.t2 183.337
R2 IB.n0 IB.t0 91.8423
R3 IB.n1 IB.t1 4.35136
R4 IB.n1 IB.n0 0.508078
R5 IB IB.n1 0.0332381
R6 VSS.n79 VSS.n73 1176.21
R7 VSS.n151 VSS.n148 1176.21
R8 VSS.n78 VSS.n75 1176.21
R9 VSS.n147 VSS.n142 1176.21
R10 VSS.n147 VSS.n143 1176.21
R11 VSS.n128 VSS.n125 1088.07
R12 VSS.n79 VSS.n74 1054.53
R13 VSS.n8 VSS.n5 1054.53
R14 VSS.n23 VSS.n22 811.506
R15 VSS.n31 VSS.n27 778.15
R16 VSS.n31 VSS.n28 778.15
R17 VSS.n56 VSS.n43 778.15
R18 VSS.n56 VSS.n44 778.15
R19 VSS.n140 VSS.n138 556.236
R20 VSS.n11 VSS.n1 382.413
R21 VSS.n156 VSS.n155 298.243
R22 VSS.n132 VSS.n131 279.719
R23 VSS.n37 VSS.n25 279.154
R24 VSS.n62 VSS.n41 278.815
R25 VSS.t2 VSS.n89 247.315
R26 VSS.n118 VSS.n113 204.424
R27 VSS.n72 VSS.n71 203.294
R28 VSS.t7 VSS.n42 191.946
R29 VSS.n69 VSS.t10 189.624
R30 VSS.n155 VSS.t14 189.624
R31 VSS.n116 VSS.n115 187.782
R32 VSS.n124 VSS.n118 183.47
R33 VSS.t8 VSS.n33 167.513
R34 VSS.n64 VSS.n38 160
R35 VSS.n64 VSS.n63 160
R36 VSS.n93 VSS.n88 138.166
R37 VSS.n20 VSS.n15 138.166
R38 VSS.n53 VSS.n50 138.166
R39 VSS.n137 VSS.n133 136.758
R40 VSS.n158 VSS.n141 136.23
R41 VSS.n18 VSS.t5 115.398
R42 VSS.t14 VSS.n152 114.837
R43 VSS.n51 VSS.t0 114.43
R44 VSS.n94 VSS.n93 91.8593
R45 VSS.n21 VSS.n20 78.6829
R46 VSS.n54 VSS.n53 78.6829
R47 VSS.n47 VSS.n46 78.6829
R48 VSS.n116 VSS.n114 77.3227
R49 VSS.n80 VSS.n72 76.424
R50 VSS.n150 VSS.n149 76.424
R51 VSS.n77 VSS.n76 76.424
R52 VSS.n146 VSS.n144 76.424
R53 VSS.n146 VSS.n145 76.424
R54 VSS.n156 VSS.t4 75.4817
R55 VSS.n133 VSS.n132 70.6977
R56 VSS.n7 VSS.n6 68.5181
R57 VSS.n38 VSS.n21 61.1205
R58 VSS.n81 VSS.n80 57.224
R59 VSS.n137 VSS.n136 54.668
R60 VSS.n30 VSS.n29 50.5605
R61 VSS.n55 VSS.n47 50.5605
R62 VSS.n55 VSS.n54 50.5605
R63 VSS.n36 VSS.n26 49.2505
R64 VSS.n158 VSS.n124 44.6176
R65 VSS.n82 VSS.n68 39.6805
R66 VSS.n141 VSS.n137 36.1417
R67 VSS.n82 VSS.n81 23.4245
R68 VSS.n10 VSS.n2 20.6255
R69 VSS.n61 VSS.n60 19.7005
R70 VSS.n84 VSS.t3 17.4601
R71 VSS.n1 VSS.n0 14.7755
R72 VSS.n32 VSS.n31 13.3929
R73 VSS.t8 VSS.n32 11.8519
R74 VSS.n12 VSS.n11 9.3005
R75 VSS.n11 VSS.n10 9.3005
R76 VSS.n65 VSS.n64 6.52902
R77 VSS.n160 VSS.t11 4.49301
R78 VSS.n110 VSS.t13 4.45895
R79 VSS.n110 VSS.t15 4.35136
R80 VSS.n38 VSS.n37 3.2005
R81 VSS.n57 VSS.n56 2.10052
R82 VSS.n95 VSS.n94 1.93119
R83 VSS.n102 VSS.n95 1.9252
R84 VSS.n122 VSS.n119 1.8415
R85 VSS.n65 VSS.n12 1.7464
R86 VSS.t7 VSS.n57 1.68204
R87 VSS.n63 VSS.n62 1.2805
R88 VSS.n83 VSS.n65 1.1024
R89 VSS.n141 VSS.n140 0.795337
R90 VSS.n140 VSS.n139 0.795337
R91 VSS.n109 VSS.n108 0.669735
R92 VSS.n109 VSS.n83 0.52389
R93 VSS.n100 VSS.n99 0.436831
R94 VSS.n99 VSS.n98 0.436742
R95 VSS.n8 VSS.n7 0.131784
R96 VSS.n9 VSS.n8 0.13084
R97 VSS.n4 VSS.n3 0.126877
R98 VSS.n9 VSS.n4 0.125988
R99 VSS.n91 VSS.n90 0.10956
R100 VSS.t2 VSS.n91 0.10956
R101 VSS.n92 VSS.t2 0.10956
R102 VSS.n93 VSS.n92 0.10956
R103 VSS.n15 VSS.n14 0.10956
R104 VSS.n14 VSS.n13 0.10956
R105 VSS.n31 VSS.n30 0.10956
R106 VSS.n50 VSS.n49 0.10956
R107 VSS.n49 VSS.n48 0.10956
R108 VSS.n56 VSS.n55 0.10956
R109 VSS.n100 VSS.n97 0.104939
R110 VSS.n97 VSS.n96 0.104537
R111 VSS.n159 VSS.n110 0.0662242
R112 VSS.n80 VSS.n79 0.0636886
R113 VSS.n79 VSS.t9 0.0636886
R114 VSS.n25 VSS.n24 0.0636886
R115 VSS.n24 VSS.n23 0.0636886
R116 VSS.n41 VSS.n40 0.0636886
R117 VSS.n40 VSS.n39 0.0636886
R118 VSS.n151 VSS.n150 0.0636886
R119 VSS.t4 VSS.n151 0.0636886
R120 VSS.n132 VSS.n128 0.0636886
R121 VSS.n128 VSS.t12 0.0636886
R122 VSS.t12 VSS.n127 0.0636886
R123 VSS.n127 VSS.n126 0.0636886
R124 VSS.n113 VSS.n112 0.0636886
R125 VSS.n112 VSS.n111 0.0636886
R126 VSS.t9 VSS.n78 0.0636886
R127 VSS.n78 VSS.n77 0.0636886
R128 VSS.t4 VSS.n147 0.0636886
R129 VSS.n147 VSS.n146 0.0636886
R130 VSS.n88 VSS.n87 0.0525185
R131 VSS.n87 VSS.n86 0.0525185
R132 VSS.n17 VSS.n16 0.0525185
R133 VSS.n18 VSS.n17 0.0525185
R134 VSS.n19 VSS.n18 0.0525185
R135 VSS.n20 VSS.n19 0.0525185
R136 VSS.n46 VSS.n45 0.0525185
R137 VSS.n53 VSS.n52 0.0525185
R138 VSS.n52 VSS.n51 0.0525185
R139 VSS.n118 VSS.n117 0.0523204
R140 VSS.n117 VSS.n116 0.0523204
R141 VSS.n160 VSS.n159 0.0483051
R142 VSS.n85 VSS.n84 0.0296391
R143 VSS.n108 VSS.n107 0.0152059
R144 VSS.n71 VSS.n70 0.015169
R145 VSS.n70 VSS.n69 0.015169
R146 VSS.n59 VSS.n58 0.015169
R147 VSS.t7 VSS.n59 0.015169
R148 VSS.n35 VSS.n34 0.015169
R149 VSS.t8 VSS.n35 0.015169
R150 VSS.n36 VSS.t8 0.015169
R151 VSS.n37 VSS.n36 0.015169
R152 VSS.n61 VSS.t7 0.015169
R153 VSS.n62 VSS.n61 0.015169
R154 VSS.n154 VSS.n153 0.015169
R155 VSS.n155 VSS.n154 0.015169
R156 VSS.n131 VSS.n130 0.015169
R157 VSS.n130 VSS.n129 0.015169
R158 VSS.n136 VSS.n135 0.015169
R159 VSS.n135 VSS.n134 0.015169
R160 VSS.n121 VSS.n120 0.015169
R161 VSS.n122 VSS.n121 0.015169
R162 VSS.n124 VSS.n123 0.0144432
R163 VSS.n123 VSS.n122 0.0144432
R164 VSS.n161 VSS.n109 0.00973214
R165 VSS VSS.n161 0.00805357
R166 VSS.n103 VSS.n102 0.0046942
R167 VSS.n104 VSS.n103 0.00420666
R168 VSS.n106 VSS.n85 0.00174202
R169 VSS.n10 VSS.n9 0.001708
R170 VSS.n101 VSS.n100 0.00107905
R171 VSS.n83 VSS.n82 0.00101351
R172 VSS.n102 VSS.n101 0.00101243
R173 VSS.n105 VSS.n104 0.001004
R174 VSS.n106 VSS.n105 0.00100001
R175 VSS.n158 VSS.n157 0.000826763
R176 VSS.n157 VSS.n156 0.000826763
R177 VSS.n68 VSS.n67 0.000756235
R178 VSS.n67 VSS.n66 0.000756235
R179 VSS.n107 VSS.n106 0.000504005
R180 VSS.n159 VSS.n158 0.000500526
R181 VSS.n161 VSS.n160 0.000500059
R182 CLK.n2 CLK.t1 319.637
R183 CLK.n6 CLK.t0 319.635
R184 CLK.n5 CLK.t5 232.303
R185 CLK.t4 CLK.n10 183.964
R186 CLK.n11 CLK.t3 182.915
R187 CLK.n11 CLK.t4 182.91
R188 CLK.t3 CLK.n5 182.769
R189 CLK.n12 CLK.t2 159.959
R190 CLK.n5 CLK.n4 1.15949
R191 CLK.n12 CLK.n11 0.56781
R192 CLK CLK.n12 0.487909
R193 CLK.n3 CLK.n2 0.0382423
R194 CLK.n7 CLK.n6 0.0255
R195 CLK.n9 CLK.n8 0.0255
R196 CLK.n1 CLK.n0 0.0232273
R197 CLK.n10 CLK.n9 0.0160001
R198 CLK.n4 CLK.n1 0.0146364
R199 CLK.n10 CLK.n7 0.00101096
R200 CLK.n4 CLK.n3 0.00100868
R201 VON.n1 VON.t4 233.888
R202 VON.n0 VON.t5 159.725
R203 VON.n2 VON.t0 17.4109
R204 VON.n2 VON.t1 9.60468
R205 VON.n4 VON.t3 8.40929
R206 VON.n0 VON.t2 8.06629
R207 VON.n1 VON.n0 1.73501
R208 VON.n3 VON.n1 0.991249
R209 VON.n4 VON.n3 0.853186
R210 VON VON.n4 0.24425
R211 VON.n3 VON.n2 0.000500726
R212 VDD.n20 VDD.n11 628.236
R213 VDD.n19 VDD.n15 628.236
R214 VDD.n49 VDD.n40 628.236
R215 VDD.n48 VDD.n44 628.236
R216 VDD.n64 VDD.n61 170.542
R217 VDD.t0 VDD.n14 136.591
R218 VDD.t2 VDD.n43 136.591
R219 VDD.n7 VDD.n5 129.692
R220 VDD.n36 VDD.n34 129.691
R221 VDD.n22 VDD.n21 112.189
R222 VDD.n51 VDD.n50 112.189
R223 VDD.n68 VDD.n64 91.343
R224 VDD.n77 VDD.n76 69.036
R225 VDD.n10 VDD.n9 67.0123
R226 VDD.n21 VDD.n10 67.0123
R227 VDD.n17 VDD.n16 67.0123
R228 VDD.n18 VDD.n17 67.0123
R229 VDD.n50 VDD.n39 67.0123
R230 VDD.n39 VDD.n38 67.0123
R231 VDD.n47 VDD.n46 67.0123
R232 VDD.n46 VDD.n45 67.0123
R233 VDD.n71 VDD.n68 38.9491
R234 VDD.n57 VDD.n29 8.85536
R235 VDD.n58 VDD.t3 7.14934
R236 VDD.n28 VDD.t1 7.14897
R237 VDD.n79 VDD.t5 4.35136
R238 VDD.n59 VDD.t4 4.35136
R239 VDD.n57 VDD.n56 2.72837
R240 VDD.n59 VDD.n58 1.81738
R241 VDD.n72 VDD.n59 1.25748
R242 VDD.n80 VDD.n28 1.00708
R243 VDD.n53 VDD.n32 0.597135
R244 VDD.n80 VDD.n79 0.311403
R245 VDD VDD.n80 0.1105
R246 VDD.n23 VDD.n22 0.104784
R247 VDD.n24 VDD.n23 0.104784
R248 VDD.n52 VDD.n51 0.104784
R249 VDD.n53 VDD.n52 0.104784
R250 VDD.n78 VDD.n74 0.0945934
R251 VDD.n3 VDD.n2 0.0694784
R252 VDD.n24 VDD.n3 0.0694784
R253 VDD.n54 VDD.n31 0.0648339
R254 VDD.n31 VDD.n30 0.0643371
R255 VDD.n21 VDD.n20 0.0265784
R256 VDD.n20 VDD.t0 0.0265784
R257 VDD.n9 VDD.n8 0.0265784
R258 VDD.t8 VDD.n6 0.0265784
R259 VDD.t0 VDD.n19 0.0265784
R260 VDD.n19 VDD.n18 0.0265784
R261 VDD.n61 VDD.n60 0.0265784
R262 VDD.n76 VDD.n75 0.0265784
R263 VDD.n50 VDD.n49 0.0265784
R264 VDD.n49 VDD.t2 0.0265784
R265 VDD.n38 VDD.n37 0.0265784
R266 VDD.n37 VDD.t7 0.0265784
R267 VDD.t2 VDD.n48 0.0265784
R268 VDD.n48 VDD.n47 0.0265784
R269 VDD.n8 VDD.n7 0.0257725
R270 VDD.n36 VDD.n35 0.02576
R271 VDD.n64 VDD.n63 0.0223212
R272 VDD.n63 VDD.n62 0.0168633
R273 VDD.n74 VDD.n72 0.0145797
R274 VDD.n79 VDD.n78 0.0111456
R275 VDD.n78 VDD.n77 0.0105432
R276 VDD.n55 VDD.n54 0.0100998
R277 VDD.n25 VDD.n1 0.0100991
R278 VDD.n1 VDD.n0 0.0096003
R279 VDD.n68 VDD.n67 0.0096003
R280 VDD.n67 VDD.t6 0.0096003
R281 VDD.n56 VDD.n55 0.0096003
R282 VDD.n5 VDD.n4 0.00505015
R283 VDD.n13 VDD.n12 0.00505015
R284 VDD.n14 VDD.n13 0.00505015
R285 VDD.n66 VDD.n65 0.00505015
R286 VDD.t6 VDD.n66 0.00505015
R287 VDD.n42 VDD.n41 0.00505015
R288 VDD.n43 VDD.n42 0.00505015
R289 VDD.n34 VDD.n33 0.00505015
R290 VDD.n7 VDD.t8 0.00255322
R291 VDD.t7 VDD.n36 0.00231811
R292 VDD.n26 VDD.n25 0.00164557
R293 VDD.n70 VDD.n69 0.00159754
R294 VDD.n72 VDD.n71 0.00133663
R295 VDD.n71 VDD.n70 0.00133663
R296 VDD.n27 VDD.n26 0.00114565
R297 VDD.n58 VDD.n57 0.00100098
R298 VDD.n54 VDD.n53 0.00100041
R299 VDD.n25 VDD.n24 0.00100008
R300 VDD.n74 VDD.n73 0.000501102
R301 VDD.n28 VDD.n27 0.000500414
R302 VIP.n0 VIP.t0 167.326
R303 VIP.n0 VIP.t1 92.4649
R304 VIP VIP.n0 1.62592
R305 VOP.n1 VOP.t4 233.929
R306 VOP.n0 VOP.t5 160.416
R307 VOP.n2 VOP.t1 17.4109
R308 VOP.n2 VOP.t0 10.2055
R309 VOP.n4 VOP.t2 7.98684
R310 VOP.n0 VOP.t3 7.55846
R311 VOP.n3 VOP.n1 1.4614
R312 VOP.n1 VOP.n0 1.19626
R313 VOP.n4 VOP.n3 0.808836
R314 VOP.n3 VOP.n2 0.154668
R315 VOP VOP.n4 0.0203171
R316 VIN.n0 VIN.t0 167.365
R317 VIN.n0 VIN.t1 92.4511
R318 VIN VIN.n0 2.11118
C0 w_1880_n1260# a_810_n2630# 0.394f
C1 w_1258_n1260# a_872_n982# 0.149f
C2 w_1880_n1260# a_872_n982# 0.12f
C3 IB a_810_n2630# 0.256f
C4 VIP VDD 0.448f
C5 VDD VON 2.93f
C6 VOP VDD 2.71f
C7 VIP a_810_n2630# 0.265f
C8 VIP a_872_n982# 0.174f
C9 w_1258_n1260# w_1880_n1260# 0.327f
C10 a_872_n982# VON 1.24f
C11 a_872_n982# VOP 0.461f
C12 VDD CLK 2.42f
C13 a_810_n2630# CLK 0.0136f
C14 VIN VDD 0.336f
C15 w_1258_n1260# VIP 0.864f
C16 w_1258_n1260# VON 0.0792f
C17 a_872_n982# CLK 0.235f
C18 w_1880_n1260# VIP 0.73f
C19 w_1880_n1260# VON 0.659f
C20 w_1258_n1260# VOP 0.658f
C21 VIN a_810_n2630# 0.278f
C22 IB VON 0.0548f
C23 w_1880_n1260# VOP 0.0988f
C24 VIN a_872_n982# 0.203f
C25 w_1258_n1260# CLK 0.57f
C26 VIP VON 0.133f
C27 w_1880_n1260# CLK 0.535f
C28 VIP VOP 0.625f
C29 IB CLK 0.0319f
C30 VOP VON 3.16f
C31 w_1258_n1260# VIN 0.795f
C32 w_1880_n1260# VIN 0.75f
C33 VIP CLK 0.35f
C34 CLK VON 1.79f
C35 VOP CLK 2.6f
C36 VIN VIP 0.108f
C37 VIN VON 0.577f
C38 VIN VOP 0.22f
C39 VDD a_810_n2630# 0.0261f
C40 a_872_n982# VDD 0.109f
C41 a_872_n982# a_810_n2630# 0.015f
C42 VIN CLK 0.588f
C43 w_1258_n1260# VDD 0.679f
C44 w_1880_n1260# VDD 0.676f
C45 IB VDD 0.0948f
C46 w_1258_n1260# a_810_n2630# 0.359f
.ends

