magic
tech sky130A
timestamp 1711205355
<< checkpaint >>
rect -649 1202 787 1226
rect -649 1178 1082 1202
rect -649 1154 1377 1178
rect -649 1130 1626 1154
rect -649 1106 1875 1130
rect -649 1082 2124 1106
rect -649 1058 2373 1082
rect -649 1034 2622 1058
rect -649 1010 2871 1034
rect -649 986 3166 1010
rect -649 962 3461 986
rect -649 938 3802 962
rect -649 914 4143 938
rect -649 890 4484 914
rect -649 866 4825 890
rect -649 842 5074 866
rect -649 818 5323 842
rect -649 794 5618 818
rect -649 770 5775 794
rect -649 746 5932 770
rect -649 722 6089 746
rect -649 -354 6246 722
rect -630 -474 6246 -354
rect -630 -3230 730 -474
rect 845 -498 6246 -474
rect 1094 -522 6246 -498
rect 1343 -546 6246 -522
rect 1592 -570 6246 -546
rect 1887 -594 6246 -570
rect 2182 -618 6246 -594
rect 2523 -642 6246 -618
rect 2864 -666 6246 -642
rect 3205 -690 6246 -666
rect 3546 -714 6246 -690
rect 3795 -738 6246 -714
rect 4044 -762 6246 -738
rect 4339 -786 6246 -762
rect 4496 -810 6246 -786
rect 4653 -834 6246 -810
rect 4810 -858 6246 -834
<< metal1 >>
rect 0 0 100 100
rect 0 -200 100 -100
rect 0 -400 100 -300
rect 0 -600 100 -500
rect 0 -800 100 -700
rect 0 -1000 100 -900
rect 0 -1200 100 -1100
rect 0 -1400 100 -1300
rect 0 -1600 100 -1500
rect 0 -1800 100 -1700
rect 0 -2000 100 -1900
rect 0 -2200 100 -2100
rect 0 -2400 100 -2300
rect 0 -2600 100 -2500
use sky130_fd_sc_hd__or4_1  x1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 157 0 1 276
box -19 -24 295 296
use sky130_fd_sc_hd__or4_1  x2
timestamp 1701704242
transform 1 0 452 0 1 252
box -19 -24 295 296
use sky130_fd_sc_hd__inv_1  x3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 4988 0 1 -132
box -19 -24 157 296
use sky130_fd_sc_hd__or3_1  x4 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 747 0 1 228
box -19 -24 249 296
use sky130_fd_sc_hd__inv_1  x5
timestamp 1701704242
transform 1 0 5145 0 1 -156
box -19 -24 157 296
use sky130_fd_sc_hd__inv_1  x6
timestamp 1701704242
transform 1 0 5302 0 1 -180
box -19 -24 157 296
use sky130_fd_sc_hd__inv_1  x7
timestamp 1701704242
transform 1 0 5459 0 1 -204
box -19 -24 157 296
use sky130_fd_sc_hd__and2_1  x8 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 996 0 1 204
box -19 -24 249 296
use sky130_fd_sc_hd__inv_1  x9
timestamp 1701704242
transform 1 0 0 0 1 300
box -19 -24 157 296
use sky130_fd_sc_hd__and2_1  x10
timestamp 1701704242
transform 1 0 1245 0 1 180
box -19 -24 249 296
use sky130_fd_sc_hd__and2_1  x11
timestamp 1701704242
transform 1 0 1494 0 1 156
box -19 -24 249 296
use sky130_fd_sc_hd__and2_1  x12
timestamp 1701704242
transform 1 0 1743 0 1 132
box -19 -24 249 296
use sky130_fd_sc_hd__and2_1  x13
timestamp 1701704242
transform 1 0 1992 0 1 108
box -19 -24 249 296
use sky130_fd_sc_hd__or4_1  x14
timestamp 1701704242
transform 1 0 2241 0 1 84
box -19 -24 295 296
use sky130_fd_sc_hd__and4_1  x15 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 2831 0 1 36
box -19 -24 341 296
use sky130_fd_sc_hd__and4_1  x16
timestamp 1701704242
transform 1 0 3172 0 1 12
box -19 -24 341 296
use sky130_fd_sc_hd__or4_1  x17
timestamp 1701704242
transform 1 0 2536 0 1 60
box -19 -24 295 296
use sky130_fd_sc_hd__and4_1  x18
timestamp 1701704242
transform 1 0 3513 0 1 -12
box -19 -24 341 296
use sky130_fd_sc_hd__and4_1  x19
timestamp 1701704242
transform 1 0 3854 0 1 -36
box -19 -24 341 296
use sky130_fd_sc_hd__and3_1  x20 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 4195 0 1 -60
box -19 -24 249 296
use sky130_fd_sc_hd__and2_1  x21
timestamp 1701704242
transform 1 0 4444 0 1 -84
box -19 -24 249 296
use sky130_fd_sc_hd__or4_1  x22
timestamp 1701704242
transform 1 0 4693 0 1 -108
box -19 -24 295 296
<< labels >>
flabel metal1 0 0 100 100 0 FreeSans 128 0 0 0 I1
port 0 nsew
flabel metal1 0 -200 100 -100 0 FreeSans 128 0 0 0 I5
port 1 nsew
flabel metal1 0 -400 100 -300 0 FreeSans 128 0 0 0 I3
port 2 nsew
flabel metal1 0 -600 100 -500 0 FreeSans 128 0 0 0 I0
port 3 nsew
flabel metal1 0 -800 100 -700 0 FreeSans 128 0 0 0 I2
port 4 nsew
flabel metal1 0 -1000 100 -900 0 FreeSans 128 0 0 0 I6
port 5 nsew
flabel metal1 0 -1200 100 -1100 0 FreeSans 128 0 0 0 I7
port 6 nsew
flabel metal1 0 -1400 100 -1300 0 FreeSans 128 0 0 0 I4
port 7 nsew
flabel metal1 0 -1600 100 -1500 0 FreeSans 128 0 0 0 EO
port 8 nsew
flabel metal1 0 -1800 100 -1700 0 FreeSans 128 0 0 0 GS
port 9 nsew
flabel metal1 0 -2000 100 -1900 0 FreeSans 128 0 0 0 A2
port 10 nsew
flabel metal1 0 -2200 100 -2100 0 FreeSans 128 0 0 0 A1
port 11 nsew
flabel metal1 0 -2400 100 -2300 0 FreeSans 128 0 0 0 A0
port 12 nsew
flabel metal1 0 -2600 100 -2500 0 FreeSans 128 0 0 0 EI
port 13 nsew
<< end >>
