* NGSPICE file created from user_analog_project_wrapper.ext - technology: sky130A

.subckt user_analog_project_wrapper io_analog[0] io_analog[10] io_analog[1] io_analog[2]
+ io_analog[8] io_analog[9] vssa2 vccd2 vccd1
X0 vccd1.t114 a_540271_687858.t5 a_540271_687858.t6 vccd1.t66 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X1 vccd1.t113 a_540271_687858.t49 a_537154_685355.t27 vccd1.t79 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X2 io_analog[10].t49 a_40125_693523.t32 vccd2.t138 vccd2.t137 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X3 a_42818_684860.t20 io_analog[9].t0 a_43026_690892.t42 vssa2.t116 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X4 a_40125_693523.t19 a_43026_690892.t49 vccd2.t57 vccd2.t20 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X5 a_43026_690892.t41 a_43026_690892.t40 vccd2.t21 vccd2.t20 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X6 a_537154_685355.t30 a_534722_685355.t6 vssa2.t140 sky130_fd_pr__res_xhigh_po_5p73 l=1e+07u
X7 vccd1.t40 a_540916_680434.t22 a_540371_681998.t5 vccd1.t10 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X8 a_40125_693523.t20 a_43026_690892.t50 vccd2.t58 vccd2.t39 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X9 a_43026_690892.t39 a_43026_690892.t38 vccd2.t40 vccd2.t39 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X10 a_534722_685355.t4 a_537154_685355.t6 vssa2.t128 sky130_fd_pr__res_xhigh_po_5p73 l=1e+07u
X11 vccd1.t112 a_540271_687858.t50 a_537154_685355.t26 vccd1.t77 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X12 a_43026_690892.t37 a_43026_690892.t36 vccd2.t19 vccd2.t6 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X13 vccd1.t111 a_540271_687858.t25 a_540271_687858.t26 vccd1.t79 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X14 a_42818_684860.t6 constant_gm_fingers_0/Vout.t14 vssa2.t50 vssa2.t49 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X15 a_40125_693523.t2 a_43026_690892.t51 vccd2.t7 vccd2.t6 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X16 vssa2.t38 constant_gm_fingers_0/Vout.t15 a_42818_684860.t4 vssa2.t37 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X17 io_analog[2].t51 a_540371_681998.t16 vssa2.t29 vssa2.t28 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X18 vssa2.t40 constant_gm_fingers_0/Vout.t16 a_42818_684860.t5 vssa2.t39 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X19 vccd1.t9 a_540916_680434.t23 a_540371_681998.t4 vccd1.t8 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X20 a_42818_684860.t0 io_analog[8].t0 a_40125_693523.t4 vssa2.t11 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X21 vccd2.t136 a_40125_693523.t33 io_analog[10].t48 vccd2.t135 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X22 io_analog[10].t52 a_37693_693523.t6 sky130_fd_pr__cap_mim_m3_1 l=1.6e+07u w=1.6e+07u
X23 vssa2.t30 a_540371_681998.t17 a_540459_681940.t27 vssa2 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X24 io_analog[10].t47 a_40125_693523.t34 vccd2.t134 vccd2.t133 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X25 vccd1.t110 a_540271_687858.t51 a_537154_685355.t25 vccd1.t71 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X26 a_40125_693523.t3 a_43026_690892.t52 vccd2.t9 vccd2.t8 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X27 a_43026_690892.t35 a_43026_690892.t34 vccd2.t29 vccd2.t8 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X28 vccd1.t48 a_540916_680434.t18 a_540916_680434.t19 vccd1.t47 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X29 vssa2.t97 a_540371_681998.t18 a_540459_681940.t26 vssa2 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X30 vccd2.t145 a_43026_690892.t32 a_43026_690892.t33 vccd2.t41 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X31 vccd2.t42 a_43026_690892.t53 a_40125_693523.t8 vccd2.t41 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X32 vccd1.t109 a_540271_687858.t45 a_540271_687858.t46 vccd1.t71 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X33 a_537154_685355.t3 io_analog[1].t0 a_540459_681940.t5 vssa2.t43 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X34 a_540916_680434.t3 a_540371_681998.t19 a_541059_678436.t9 vssa2.t98 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X35 vssa2.t4 constant_gm_fingers_0/Vout.t10 constant_gm_fingers_0/Vout.t11 vssa2.t3 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=1e+06u
X36 io_analog[2].t50 a_540371_681998.t20 vssa2.t83 vssa2.t82 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X37 io_analog[10].t46 a_40125_693523.t35 vccd2.t132 vccd2.t131 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X38 vccd1.t50 a_537154_685355.t32 io_analog[2].t39 vccd1.t31 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X39 io_analog[10].t53 a_37693_693523.t5 sky130_fd_pr__cap_mim_m3_1 l=1.6e+07u w=1.6e+07u
X40 vssa2.t127 a_41722_677112.t9 vssa2 sky130_fd_pr__res_xhigh_po_5p73 l=6.9e+07u
X41 a_43833_677960.t5 constant_gm_fingers_0/Vout.t17 a_41722_677112.t5 vssa2.t137 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X42 vccd2.t33 a_43833_677960.t20 a_43833_677960.t21 vccd2.t32 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X43 vccd2.t130 a_40125_693523.t36 io_analog[10].t45 vccd2.t129 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X44 vccd1.t108 a_540271_687858.t52 a_537154_685355.t24 vccd1.t66 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X45 a_40125_693523.t9 a_43026_690892.t54 vccd2.t44 vccd2.t43 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X46 a_43026_690892.t31 a_43026_690892.t30 vccd2.t50 vccd2.t43 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X47 a_42818_684860.t25 constant_gm_fingers_0/Vout.t18 vssa2.t139 vssa2.t138 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X48 vccd2.t160 a_43026_690892.t28 a_43026_690892.t29 vccd2.t47 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X49 vccd2.t48 a_43026_690892.t55 a_40125_693523.t11 vccd2.t47 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X50 vccd1.t51 a_537154_685355.t33 io_analog[2].t38 vccd1.t31 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X51 vccd1.t107 a_540271_687858.t43 a_540271_687858.t44 vccd1.t66 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X52 vccd1.t106 a_540271_687858.t53 a_537154_685355.t23 vccd1.t93 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X53 vccd1.t105 a_540271_687858.t54 a_537154_685355.t22 vccd1.t79 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X54 vccd1.t52 a_537154_685355.t34 io_analog[2].t37 vccd1.t14 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X55 io_analog[10].t5 constant_gm_fingers_0/Vout.t19 vssa2.t76 vssa2.t75 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X56 io_analog[2].t52 a_534722_685355.t2 sky130_fd_pr__cap_mim_m3_1 l=1.6e+07u w=1.6e+07u
X57 io_analog[10].t44 a_40125_693523.t37 vccd2.t128 vccd2.t127 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X58 a_43026_690892.t48 io_analog[9].t1 a_42818_684860.t19 vssa2.t115 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X59 vssa2.t78 constant_gm_fingers_0/Vout.t20 io_analog[10].t6 vssa2.t77 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X60 vssa2.t151 a_541059_678436.t3 vssa2 sky130_fd_pr__res_xhigh_po_5p73 l=6.9e+07u
X61 vssa2.t7 a_41722_677112.t1 vssa2 sky130_fd_pr__res_xhigh_po_5p73 l=6.9e+07u
X62 a_540459_681940.t10 io_analog[0].t0 a_540271_687858.t4 vssa2.t100 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X63 vccd2.t49 a_43026_690892.t56 a_40125_693523.t12 vccd2.t10 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X64 vccd2.t11 a_43026_690892.t26 a_43026_690892.t27 vccd2.t10 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X65 io_analog[10].t43 a_40125_693523.t38 vccd2.t108 vccd2.t107 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X66 vccd1.t104 a_540271_687858.t37 a_540271_687858.t38 vccd1.t93 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X67 a_540916_680434.t7 a_540916_680434.t6 a_540371_681998.t7 vssa2.t85 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.5e+06u l=500000u
X68 vccd1.t53 a_537154_685355.t35 io_analog[2].t36 vccd1.t14 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X69 vccd2.t139 a_43833_677960.t22 constant_gm_fingers_0/Vout.t3 vccd2.t16 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X70 constant_gm_fingers_0/Vout.t1 a_43833_677960.t23 vccd2.t28 vccd2.t24 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X71 vccd1.t103 a_540271_687858.t35 a_540271_687858.t36 vccd1.t93 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X72 vccd2.t106 a_40125_693523.t39 io_analog[10].t42 vccd2.t105 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X73 a_537154_685355.t5 io_analog[1].t1 a_540459_681940.t9 vssa2.t99 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X74 a_43833_677960.t4 constant_gm_fingers_0/Vout.t21 a_41722_677112.t2 vssa2.t156 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X75 a_41722_677112.t6 constant_gm_fingers_0/Vout.t22 a_43833_677960.t3 vssa2.t157 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X76 io_analog[2].t49 a_540371_681998.t21 vssa2.t84 vssa2 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X77 a_40125_693523.t10 io_analog[8].t1 a_42818_684860.t11 vssa2.t73 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X78 io_analog[10].t54 a_37693_693523.t4 sky130_fd_pr__cap_mim_m3_1 l=1.6e+07u w=1.6e+07u
X79 a_43833_677960.t19 a_43833_677960.t18 vccd2.t15 vccd2.t14 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X80 a_540459_681940.t11 io_analog[0].t1 a_540271_687858.t47 vssa2.t133 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X81 a_40125_693523.t21 io_analog[8].t2 a_42818_684860.t21 vssa2.t123 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X82 io_analog[2].t53 a_534722_685355.t3 sky130_fd_pr__cap_mim_m3_1 l=1.6e+07u w=1.6e+07u
X83 io_analog[10].t41 a_40125_693523.t40 vccd2.t126 vccd2.t125 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X84 io_analog[10].t40 a_40125_693523.t41 vccd2.t124 vccd2.t123 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X85 vccd1.t102 a_540271_687858.t55 a_537154_685355.t21 vccd1.t71 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X86 vssa2.t142 a_540371_681998.t22 a_540459_681940.t25 vssa2 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X87 a_40125_693523.t28 a_43026_690892.t57 vccd2.t156 vccd2.t45 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X88 a_43026_690892.t25 a_43026_690892.t24 vccd2.t46 vccd2.t45 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X89 vssa2.t65 constant_gm_fingers_0/Vout.t23 a_42818_684860.t9 vssa2.t64 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X90 a_42818_684860.t10 constant_gm_fingers_0/Vout.t24 vssa2.t67 vssa2.t66 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X91 vccd2.t122 a_40125_693523.t42 io_analog[10].t39 vccd2.t121 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X92 a_43026_690892.t23 a_43026_690892.t22 vccd2.t143 vccd2.t142 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X93 vccd1.t115 a_540916_680434.t16 a_540916_680434.t17 vccd1.t33 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X94 a_40125_693523.t29 a_43026_690892.t58 vccd2.t157 vccd2.t142 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X95 vssa2.t143 a_540371_681998.t23 a_540459_681940.t24 vssa2.t46 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X96 vccd2.t110 a_40125_693523.t43 io_analog[10].t38 vccd2.t109 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X97 io_analog[10].t37 a_40125_693523.t44 vccd2.t120 vccd2.t119 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X98 vccd1.t101 a_540271_687858.t56 a_537154_685355.t20 vccd1.t66 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X99 vccd1.t29 a_537154_685355.t36 io_analog[2].t35 vccd1.t2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X100 constant_gm_fingers_0/Vout.t9 constant_gm_fingers_0/Vout.t8 vssa2.t94 vssa2.t93 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=1e+06u
X101 constant_gm_fingers_0/Vout.t3 a_43833_677960.t24 vccd2.t38 vccd2.t37 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X102 vccd2.t118 a_40125_693523.t45 io_analog[10].t36 vccd2.t117 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X103 a_42818_684860.t22 io_analog[8].t3 a_40125_693523.t22 vssa2.t124 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X104 io_analog[2].t48 a_540371_681998.t24 vssa2.t45 vssa2.t35 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X105 vccd2.t31 a_43026_690892.t20 a_43026_690892.t21 vccd2.t30 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X106 vccd2.t51 a_43026_690892.t59 a_40125_693523.t13 vccd2.t30 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X107 vccd2.t152 a_43026_690892.t18 a_43026_690892.t19 vccd2.t52 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X108 a_537154_685355.t28 a_534722_685355.t5 vssa2.t140 sky130_fd_pr__res_xhigh_po_5p73 l=1e+07u
X109 vssa2.t47 a_540371_681998.t25 a_540459_681940.t23 vssa2.t46 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X110 io_analog[10].t35 a_40125_693523.t46 vccd2.t116 vccd2.t115 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X111 vccd2.t53 a_43026_690892.t60 a_40125_693523.t14 vccd2.t52 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X112 a_534722_685355.t7 a_537154_685355.t31 vssa2.t128 sky130_fd_pr__res_xhigh_po_5p73 l=1e+07u
X113 vccd1.t30 a_537154_685355.t37 io_analog[2].t34 vccd1.t2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X114 vccd1.t22 a_540916_680434.t14 a_540916_680434.t15 vccd1.t21 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X115 vccd1.t100 a_540271_687858.t57 a_537154_685355.t19 vccd1.t93 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X116 io_analog[2].t54 a_534722_685355.t0 sky130_fd_pr__cap_mim_m3_1 l=1.6e+07u w=1.6e+07u
X117 vssa2.t54 constant_gm_fingers_0/Vout.t25 a_42818_684860.t7 vssa2.t53 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X118 vccd2.t114 a_40125_693523.t47 io_analog[10].t34 vccd2.t113 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X119 a_540916_680434.t0 a_540371_681998.t26 a_541059_678436.t8 vssa2.t79 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X120 a_540371_681998.t15 a_540371_681998.t14 vssa2.t52 vssa2.t51 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=1e+06u
X121 a_42818_684860.t18 io_analog[9].t2 a_43026_690892.t47 vssa2.t114 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X122 a_42818_684860.t17 io_analog[9].t3 a_43026_690892.t44 vssa2.t113 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X123 vccd1.t32 a_537154_685355.t38 io_analog[2].t33 vccd1.t31 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X124 io_analog[10].t33 a_40125_693523.t48 vccd2.t112 vccd2.t111 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X125 vccd1.t36 a_537154_685355.t39 io_analog[2].t32 vccd1.t35 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X126 vccd1.t99 a_540271_687858.t11 a_540271_687858.t12 vccd1.t93 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X127 a_537154_685355.t29 io_analog[1].t2 a_540459_681940.t13 vssa2.t141 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X128 io_analog[2].t47 a_540371_681998.t27 vssa2.t81 vssa2.t80 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X129 io_analog[10].t2 constant_gm_fingers_0/Vout.t26 vssa2.t56 vssa2.t55 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X130 a_540459_681940.t12 io_analog[0].t2 a_540271_687858.t48 vssa2.t134 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X131 io_analog[10].t9 constant_gm_fingers_0/Vout.t27 vssa2.t120 vssa2.t119 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X132 vccd1.t37 a_537154_685355.t40 io_analog[2].t31 vccd1.t31 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X133 vssa2.t6 constant_gm_fingers_0/Vout.t6 constant_gm_fingers_0/Vout.t7 vssa2.t5 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=1e+06u
X134 vccd1.t16 a_540916_680434.t24 a_540371_681998.t3 vccd1.t0 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X135 a_42818_684860.t23 io_analog[8].t4 a_40125_693523.t23 vssa2.t126 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X136 vccd1.t38 a_537154_685355.t41 io_analog[2].t30 vccd1.t35 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X137 io_analog[10].t32 a_40125_693523.t49 vccd2.t104 vccd2.t103 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X138 vccd1.t63 a_537154_685355.t42 io_analog[2].t29 vccd1.t27 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X139 a_43833_677960.t2 constant_gm_fingers_0/Vout.t28 a_41722_677112.t7 vssa2.t121 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X140 vccd2.t102 a_40125_693523.t50 io_analog[10].t31 vccd2.t101 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X141 vccd1.t98 a_540271_687858.t58 a_537154_685355.t18 vccd1.t68 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X142 vssa2.t0 a_41722_677112.t0 vssa2 sky130_fd_pr__res_xhigh_po_5p73 l=6.9e+07u
X143 io_analog[10].t30 a_40125_693523.t51 vccd2.t100 vccd2.t99 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X144 vccd2.t1 a_43026_690892.t16 a_43026_690892.t17 vccd2.t0 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X145 a_43026_690892.t43 io_analog[9].t4 a_42818_684860.t16 vssa2.t112 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X146 vccd2.t54 a_43026_690892.t61 a_40125_693523.t15 vccd2.t0 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X147 vccd1.t64 a_537154_685355.t43 io_analog[2].t28 vccd1.t27 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X148 a_37693_693523.t2 a_40125_693523.t17 vssa2.t44 sky130_fd_pr__res_xhigh_po_5p73 l=1e+07u
X149 vccd2.t98 a_40125_693523.t52 io_analog[10].t29 vccd2.t97 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X150 vccd1.t95 a_540271_687858.t31 a_540271_687858.t32 vccd1.t68 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X151 vssa2.t145 constant_gm_fingers_0/Vout.t29 a_42818_684860.t26 vssa2.t144 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X152 a_540459_681940.t8 io_analog[0].t3 a_540271_687858.t3 vssa2.t59 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X153 a_43833_677960.t9 a_43833_677960.t8 constant_gm_fingers_0/Vout.t12 vssa2.t86 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.5e+06u l=500000u
X154 vccd1.t97 a_540271_687858.t33 a_540271_687858.t34 vccd1.t68 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X155 vssa2.t68 a_540371_681998.t28 a_540459_681940.t22 vssa2 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X156 io_analog[2].t46 a_540371_681998.t29 vssa2.t70 vssa2.t69 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X157 vssa2.t41 a_541059_678436.t0 vssa2 sky130_fd_pr__res_xhigh_po_5p73 l=6.9e+07u
X158 io_analog[10].t28 a_40125_693523.t53 vccd2.t96 vccd2.t95 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X159 vssa2.t147 constant_gm_fingers_0/Vout.t30 io_analog[10].t51 vssa2.t146 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X160 vssa2.t125 a_41722_677112.t8 vssa2 sky130_fd_pr__res_xhigh_po_5p73 l=6.9e+07u
X161 vccd1.t11 a_540916_680434.t12 a_540916_680434.t13 vccd1.t10 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X162 vccd1.t96 a_540271_687858.t59 a_537154_685355.t17 vccd1.t74 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X163 vssa2.t154 a_540371_681998.t30 a_540459_681940.t21 vssa2.t46 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X164 io_analog[10].t27 a_40125_693523.t54 vccd2.t94 vccd2.t93 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X165 vccd2.t92 a_40125_693523.t55 io_analog[10].t26 vccd2.t91 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X166 a_540371_681998.t13 a_540371_681998.t12 vssa2.t153 vssa2.t152 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=1e+06u
X167 a_43026_690892.t15 a_43026_690892.t14 vccd2.t149 vccd2.t55 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X168 a_40125_693523.t16 a_43026_690892.t62 vccd2.t56 vccd2.t55 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X169 vccd1.t65 a_537154_685355.t44 io_analog[2].t27 vccd1.t18 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X170 vssa2.t155 a_540371_681998.t31 a_540459_681940.t20 vssa2 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X171 vccd2.t158 a_43833_677960.t25 constant_gm_fingers_0/Vout.t1 vccd2.t32 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X172 vccd1.t94 a_540271_687858.t60 a_537154_685355.t16 vccd1.t93 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X173 vccd1.t49 a_540916_680434.t10 a_540916_680434.t11 vccd1.t8 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X174 vccd2.t3 a_43026_690892.t63 a_40125_693523.t0 vccd2.t2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X175 vccd2.t148 a_43026_690892.t12 a_43026_690892.t13 vccd2.t2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X176 vccd1.t92 a_540271_687858.t29 a_540271_687858.t30 vccd1.t74 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X177 vccd2.t155 a_43833_677960.t16 a_43833_677960.t17 vccd2.t26 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X178 vccd1.t91 a_540271_687858.t27 a_540271_687858.t28 vccd1.t74 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X179 a_540916_680434.t2 a_540371_681998.t32 a_541059_678436.t7 vssa2.t95 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X180 constant_gm_fingers_0/Vout.t13 a_43833_677960.t6 a_43833_677960.t7 vssa2.t122 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.5e+06u l=500000u
X181 io_analog[10].t25 a_40125_693523.t56 vccd2.t90 vccd2.t89 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X182 a_41722_677112.t3 constant_gm_fingers_0/Vout.t31 a_43833_677960.t1 vssa2.t148 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X183 vccd1.t116 a_540916_680434.t25 a_540371_681998.t2 vccd1.t47 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X184 io_analog[2].t45 a_540371_681998.t33 vssa2.t96 vssa2.t28 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X185 a_43026_690892.t46 io_analog[9].t5 a_42818_684860.t15 vssa2.t111 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X186 vccd1.t17 a_537154_685355.t45 io_analog[2].t26 vccd1.t2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X187 a_42818_684860.t27 constant_gm_fingers_0/Vout.t32 vssa2.t150 vssa2.t149 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X188 vccd1.t19 a_537154_685355.t46 io_analog[2].t25 vccd1.t18 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X189 vccd2.t88 a_40125_693523.t57 io_analog[10].t24 vccd2.t87 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X190 vccd2.t86 a_40125_693523.t58 io_analog[10].t23 vccd2.t85 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X191 a_42818_684860.t8 io_analog[8].t5 a_40125_693523.t7 vssa2.t57 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X192 vccd1.t20 a_537154_685355.t47 io_analog[2].t24 vccd1.t4 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X193 a_37693_693523.t1 a_40125_693523.t6 vssa2.t44 sky130_fd_pr__res_xhigh_po_5p73 l=1e+07u
X194 a_42818_684860.t24 constant_gm_fingers_0/Vout.t33 vssa2.t130 vssa2.t129 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X195 vssa2.t92 a_540371_681998.t34 a_540459_681940.t19 vssa2.t91 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X196 io_analog[10].t22 a_40125_693523.t59 vccd2.t84 vccd2.t83 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X197 io_analog[10].t55 a_37693_693523.t3 sky130_fd_pr__cap_mim_m3_1 l=1.6e+07u w=1.6e+07u
X198 vccd1.t3 a_537154_685355.t48 io_analog[2].t23 vccd1.t2 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X199 vssa2.t132 constant_gm_fingers_0/Vout.t34 io_analog[10].t50 vssa2.t131 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X200 vccd1.t5 a_537154_685355.t49 io_analog[2].t22 vccd1.t4 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X201 vccd1.t7 a_537154_685355.t50 io_analog[2].t21 vccd1.t6 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X202 vccd2.t82 a_40125_693523.t60 io_analog[10].t21 vccd2.t81 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X203 vccd1.t90 a_540271_687858.t61 a_537154_685355.t15 vccd1.t68 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X204 vssa2.t17 constant_gm_fingers_0/Vout.t35 io_analog[10].t0 vssa2.t16 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X205 vccd1.t89 a_540271_687858.t62 a_537154_685355.t14 vccd1.t77 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X206 a_537154_685355.t4 io_analog[1].t3 a_540459_681940.t6 vssa2.t48 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X207 a_540916_680434.t1 a_540371_681998.t35 a_541059_678436.t6 vssa2 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X208 constant_gm_fingers_0/Vout.t5 constant_gm_fingers_0/Vout.t4 vssa2.t10 vssa2.t9 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=1e+06u
X209 io_analog[2].t44 a_540371_681998.t36 vssa2.t12 vssa2 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X210 vccd2.t80 a_40125_693523.t61 io_analog[10].t20 vccd2.t79 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X211 a_540459_681940.t1 io_analog[0].t4 a_540271_687858.t1 vssa2.t2 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X212 vccd1.t54 a_537154_685355.t51 io_analog[2].t20 vccd1.t35 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X213 constant_gm_fingers_0/Vout.t2 a_43833_677960.t26 vccd2.t36 vccd2.t14 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X214 vccd1.t55 a_537154_685355.t52 io_analog[2].t19 vccd1.t6 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X215 vccd1.t56 a_537154_685355.t53 io_analog[2].t18 vccd1.t23 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X216 vccd1.t44 a_537154_685355.t54 io_analog[2].t17 vccd1.t25 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X217 a_40125_693523.t5 a_37693_693523.t0 vssa2.t32 sky130_fd_pr__res_xhigh_po_5p73 l=1e+07u
X218 vccd1.t88 a_540271_687858.t21 a_540271_687858.t22 vccd1.t77 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X219 vccd1.t87 a_540271_687858.t19 a_540271_687858.t20 vccd1.t68 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X220 vccd1.t86 a_540271_687858.t17 a_540271_687858.t18 vccd1.t77 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X221 a_537154_685355.t0 io_analog[1].t4 a_540459_681940.t2 vssa2.t20 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X222 vccd2.t78 a_40125_693523.t62 io_analog[10].t19 vccd2.t77 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X223 a_42818_684860.t1 constant_gm_fingers_0/Vout.t36 vssa2.t19 vssa2.t18 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X224 vccd1.t85 a_540271_687858.t63 a_537154_685355.t13 vccd1.t74 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X225 vccd1.t45 a_537154_685355.t55 io_analog[2].t16 vccd1.t35 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X226 vccd1.t46 a_537154_685355.t56 io_analog[2].t15 vccd1.t27 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X227 vccd1.t24 a_537154_685355.t57 io_analog[2].t14 vccd1.t23 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X228 io_analog[10].t18 a_40125_693523.t63 vccd2.t76 vccd2.t75 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X229 vccd1.t26 a_537154_685355.t58 io_analog[2].t13 vccd1.t25 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X230 vssa2.t13 a_540371_681998.t37 a_540459_681940.t18 vssa2 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X231 io_analog[2].t55 a_534722_685355.t1 sky130_fd_pr__cap_mim_m3_1 l=1.6e+07u w=1.6e+07u
X232 vccd2.t18 a_43026_690892.t10 a_43026_690892.t11 vccd2.t4 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X233 a_43026_690892.t45 io_analog[9].t6 a_42818_684860.t14 vssa2.t110 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X234 vccd2.t5 a_43026_690892.t64 a_40125_693523.t1 vccd2.t4 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X235 io_analog[10].t1 constant_gm_fingers_0/Vout.t37 vssa2.t22 vssa2.t21 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X236 a_540916_680434.t5 a_540916_680434.t4 a_540371_681998.t6 vssa2.t8 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=2.5e+06u l=500000u
X237 a_40125_693523.t24 a_43026_690892.t65 vccd2.t140 vccd2.t12 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X238 a_43026_690892.t9 a_43026_690892.t8 vccd2.t13 vccd2.t12 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X239 vccd1.t84 a_540271_687858.t41 a_540271_687858.t42 vccd1.t74 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X240 vccd1.t28 a_537154_685355.t59 io_analog[2].t12 vccd1.t27 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X241 vssa2.t107 a_540371_681998.t38 a_540459_681940.t17 vssa2.t46 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X242 vccd1.t34 a_540916_680434.t26 a_540371_681998.t1 vccd1.t33 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X243 vccd2.t74 a_40125_693523.t64 io_analog[10].t17 vccd2.t73 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X244 a_540459_681940.t7 io_analog[0].t5 a_540271_687858.t2 vssa2.t58 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X245 io_analog[10].t16 a_40125_693523.t65 vccd2.t72 vccd2.t71 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X246 a_40125_693523.t30 a_37693_693523.t7 vssa2.t32 sky130_fd_pr__res_xhigh_po_5p73 l=1e+07u
X247 vccd2.t17 a_43833_677960.t14 a_43833_677960.t15 vccd2.t16 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X248 a_43833_677960.t13 a_43833_677960.t12 vccd2.t25 vccd2.t24 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X249 vssa2.t109 a_540371_681998.t39 a_540459_681940.t16 vssa2.t108 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X250 io_analog[2].t43 a_540371_681998.t40 vssa2.t34 vssa2.t33 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X251 vccd1.t83 a_540271_687858.t64 a_537154_685355.t12 vccd1.t79 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X252 a_540371_681998.t11 a_540371_681998.t10 vssa2.t72 vssa2.t71 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=1e+06u
X253 a_40125_693523.t25 a_43026_690892.t66 vccd2.t141 vccd2.t22 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X254 a_43026_690892.t7 a_43026_690892.t6 vccd2.t23 vccd2.t22 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X255 vccd1.t57 a_537154_685355.t60 io_analog[2].t11 vccd1.t18 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X256 a_42818_684860.t2 constant_gm_fingers_0/Vout.t38 vssa2.t24 vssa2.t23 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X257 vssa2.t88 constant_gm_fingers_0/Vout.t39 a_42818_684860.t12 vssa2.t87 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X258 vccd1.t69 a_540271_687858.t65 a_537154_685355.t11 vccd1.t68 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X259 vccd1.t82 a_540271_687858.t39 a_540271_687858.t40 vccd1.t79 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X260 vccd1.t81 a_540271_687858.t66 a_537154_685355.t10 vccd1.t77 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X261 vccd1.t80 a_540271_687858.t15 a_540271_687858.t16 vccd1.t79 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X262 vssa2.t74 a_541059_678436.t1 vssa2 sky130_fd_pr__res_xhigh_po_5p73 l=6.9e+07u
X263 vccd2.t70 a_40125_693523.t66 io_analog[10].t15 vccd2.t69 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X264 a_43026_690892.t5 a_43026_690892.t4 vccd2.t151 vccd2.t150 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X265 a_40125_693523.t18 io_analog[8].t6 a_42818_684860.t13 vssa2.t105 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X266 vccd1.t58 a_537154_685355.t61 io_analog[2].t10 vccd1.t18 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X267 vccd1.t59 a_537154_685355.t62 io_analog[2].t9 vccd1.t4 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X268 vccd1.t39 a_540916_680434.t27 a_540371_681998.t0 vccd1.t21 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X269 a_40125_693523.t26 a_43026_690892.t67 vccd2.t153 vccd2.t150 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X270 io_analog[10].t7 constant_gm_fingers_0/Vout.t40 vssa2.t90 vssa2.t89 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X271 a_537154_685355.t1 io_analog[1].t5 a_540459_681940.t3 vssa2.t31 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X272 vccd2.t68 a_40125_693523.t67 io_analog[10].t14 vccd2.t67 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X273 io_analog[2].t42 a_540371_681998.t41 vssa2.t36 vssa2.t35 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X274 vccd1.t78 a_540271_687858.t13 a_540271_687858.t14 vccd1.t77 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X275 vccd1.t76 a_540271_687858.t67 a_537154_685355.t9 vccd1.t71 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X276 vssa2.t106 a_541059_678436.t2 vssa2 sky130_fd_pr__res_xhigh_po_5p73 l=6.9e+07u
X277 a_540371_681998.t9 a_540371_681998.t8 vssa2.t15 vssa2.t14 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.25e+06u l=1e+06u
X278 vssa2.t135 a_540371_681998.t42 a_540459_681940.t15 vssa2.t46 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X279 vccd1.t75 a_540271_687858.t68 a_537154_685355.t8 vccd1.t74 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X280 vccd1.t12 a_537154_685355.t63 io_analog[2].t8 vccd1.t4 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X281 vccd1.t13 a_537154_685355.t64 io_analog[2].t7 vccd1.t6 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X282 vccd1.t15 a_537154_685355.t65 io_analog[2].t6 vccd1.t14 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X283 a_41722_677112.t4 constant_gm_fingers_0/Vout.t41 a_43833_677960.t0 vssa2.t25 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X284 a_43833_677960.t11 a_43833_677960.t10 vccd2.t144 vccd2.t37 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X285 vccd2.t66 a_40125_693523.t68 io_analog[10].t13 vccd2.t65 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X286 vccd1.t73 a_540271_687858.t9 a_540271_687858.t10 vccd1.t71 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X287 a_540916_680434.t21 a_540371_681998.t43 a_541059_678436.t5 vssa2.t136 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X288 vccd1.t72 a_540271_687858.t7 a_540271_687858.t8 vccd1.t71 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X289 io_analog[10].t12 a_40125_693523.t69 vccd2.t64 vccd2.t63 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X290 vccd1.t41 a_537154_685355.t66 io_analog[2].t5 vccd1.t6 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X291 vssa2.t27 constant_gm_fingers_0/Vout.t42 a_42818_684860.t3 vssa2.t26 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X292 a_540916_680434.t20 a_540371_681998.t44 a_541059_678436.t4 vssa2.t103 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X293 vccd1.t1 a_540916_680434.t8 a_540916_680434.t9 vccd1.t0 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X294 vccd2.t154 a_43026_690892.t68 a_40125_693523.t27 vccd2.t34 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X295 vccd2.t35 a_43026_690892.t2 a_43026_690892.t3 vccd2.t34 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X296 vccd1.t70 a_540271_687858.t69 a_537154_685355.t7 vccd1.t66 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X297 vccd1.t42 a_537154_685355.t67 io_analog[2].t4 vccd1.t25 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X298 vccd1.t43 a_537154_685355.t68 io_analog[2].t3 vccd1.t23 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X299 vccd1.t60 a_537154_685355.t69 io_analog[2].t2 vccd1.t14 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X300 a_537154_685355.t2 io_analog[1].t6 a_540459_681940.t4 vssa2.t42 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X301 io_analog[2].t41 a_540371_681998.t45 vssa2.t104 vssa2 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X302 io_analog[2].t40 a_540371_681998.t46 vssa2.t101 vssa2 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X303 vccd2.t159 a_43026_690892.t69 a_40125_693523.t31 vccd2.t146 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X304 vccd2.t147 a_43026_690892.t0 a_43026_690892.t1 vccd2.t146 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X305 a_540459_681940.t0 io_analog[0].t6 a_540271_687858.t0 vssa2.t1 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X306 vssa2.t61 constant_gm_fingers_0/Vout.t43 io_analog[10].t3 vssa2.t60 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X307 vssa2.t102 a_540371_681998.t47 a_540459_681940.t14 vssa2 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X308 vssa2.t63 constant_gm_fingers_0/Vout.t44 io_analog[10].t4 vssa2.t62 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X309 vccd2.t62 a_40125_693523.t70 io_analog[10].t11 vccd2.t61 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X310 io_analog[10].t10 a_40125_693523.t71 vccd2.t60 vccd2.t59 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X311 vccd1.t67 a_540271_687858.t23 a_540271_687858.t24 vccd1.t66 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X312 io_analog[10].t8 constant_gm_fingers_0/Vout.t45 vssa2.t118 vssa2.t117 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
X313 vccd1.t61 a_537154_685355.t70 io_analog[2].t1 vccd1.t25 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X314 vccd1.t62 a_537154_685355.t71 io_analog[2].t0 vccd1.t23 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=500000u
X315 vccd2.t27 a_43833_677960.t27 constant_gm_fingers_0/Vout.t0 vccd2.t26 sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=5e+06u l=1e+06u
R0 a_540271_687858.n7 a_540271_687858.t7 271.872
R1 a_540271_687858.n30 a_540271_687858.t17 271.872
R2 a_540271_687858.n131 a_540271_687858.t21 271.872
R3 a_540271_687858.n42 a_540271_687858.t9 271.872
R4 a_540271_687858.n59 a_540271_687858.t31 271.872
R5 a_540271_687858.n64 a_540271_687858.t39 271.872
R6 a_540271_687858.n26 a_540271_687858.t37 271.872
R7 a_540271_687858.n28 a_540271_687858.t29 271.872
R8 a_540271_687858.n123 a_540271_687858.t41 271.872
R9 a_540271_687858.n115 a_540271_687858.t11 271.872
R10 a_540271_687858.n66 a_540271_687858.t25 271.872
R11 a_540271_687858.n68 a_540271_687858.t19 271.872
R12 a_540271_687858.n77 a_540271_687858.t45 271.872
R13 a_540271_687858.n110 a_540271_687858.t35 271.872
R14 a_540271_687858.n111 a_540271_687858.t27 271.872
R15 a_540271_687858.n47 a_540271_687858.t15 271.872
R16 a_540271_687858.n45 a_540271_687858.t33 271.872
R17 a_540271_687858.n23 a_540271_687858.t13 271.872
R18 a_540271_687858.n98 a_540271_687858.t43 271.872
R19 a_540271_687858.n48 a_540271_687858.t5 271.872
R20 a_540271_687858.n65 a_540271_687858.t23 271.872
R21 a_540271_687858.n18 a_540271_687858.t50 136.729
R22 a_540271_687858.n19 a_540271_687858.t66 136.729
R23 a_540271_687858.n25 a_540271_687858.t62 136.729
R24 a_540271_687858.n119 a_540271_687858.t68 136.727
R25 a_540271_687858.n122 a_540271_687858.t59 136.724
R26 a_540271_687858.n120 a_540271_687858.t63 136.724
R27 a_540271_687858.n93 a_540271_687858.t56 135.244
R28 a_540271_687858.n90 a_540271_687858.t69 135.244
R29 a_540271_687858.n72 a_540271_687858.t55 135.243
R30 a_540271_687858.n118 a_540271_687858.t60 135.243
R31 a_540271_687858.n121 a_540271_687858.t53 135.243
R32 a_540271_687858.n92 a_540271_687858.t52 135.243
R33 a_540271_687858.n117 a_540271_687858.t57 135.243
R34 a_540271_687858.n74 a_540271_687858.t51 135.243
R35 a_540271_687858.n75 a_540271_687858.t67 135.243
R36 a_540271_687858.n94 a_540271_687858.t54 135.243
R37 a_540271_687858.n91 a_540271_687858.t64 135.243
R38 a_540271_687858.n85 a_540271_687858.t65 135.242
R39 a_540271_687858.n83 a_540271_687858.t58 135.242
R40 a_540271_687858.n87 a_540271_687858.t61 135.242
R41 a_540271_687858.n96 a_540271_687858.t49 135.242
R42 a_540271_687858.n113 a_540271_687858.n112 9.3
R43 a_540271_687858.n11 a_540271_687858.n37 9.3
R44 a_540271_687858.n13 a_540271_687858.n102 9.3
R45 a_540271_687858.n127 a_540271_687858.n126 9.3
R46 a_540271_687858.n109 a_540271_687858.n108 9.3
R47 a_540271_687858.n5 a_540271_687858.n52 9.3
R48 a_540271_687858.n54 a_540271_687858.n53 9.3
R49 a_540271_687858.n34 a_540271_687858.n43 9.3
R50 a_540271_687858.n26 a_540271_687858.t38 6.215
R51 a_540271_687858.n110 a_540271_687858.t36 6.215
R52 a_540271_687858.n80 a_540271_687858.t47 6.131
R53 a_540271_687858.n39 a_540271_687858.t34 5.713
R54 a_540271_687858.n29 a_540271_687858.t8 5.713
R55 a_540271_687858.n130 a_540271_687858.t22 5.713
R56 a_540271_687858.n41 a_540271_687858.t10 5.713
R57 a_540271_687858.n57 a_540271_687858.t32 5.713
R58 a_540271_687858.n63 a_540271_687858.t40 5.713
R59 a_540271_687858.n50 a_540271_687858.t24 5.713
R60 a_540271_687858.n106 a_540271_687858.t30 5.713
R61 a_540271_687858.n124 a_540271_687858.t42 5.713
R62 a_540271_687858.n114 a_540271_687858.t12 5.713
R63 a_540271_687858.n100 a_540271_687858.t44 5.713
R64 a_540271_687858.n89 a_540271_687858.t26 5.713
R65 a_540271_687858.n70 a_540271_687858.t20 5.713
R66 a_540271_687858.n76 a_540271_687858.t46 5.713
R67 a_540271_687858.n1 a_540271_687858.t6 5.713
R68 a_540271_687858.n46 a_540271_687858.t16 5.713
R69 a_540271_687858.n21 a_540271_687858.t14 5.713
R70 a_540271_687858.n128 a_540271_687858.t3 3.753
R71 a_540271_687858.n105 a_540271_687858.t48 3.48
R72 a_540271_687858.n103 a_540271_687858.t4 3.48
R73 a_540271_687858.n81 a_540271_687858.t1 3.48
R74 a_540271_687858.n80 a_540271_687858.t2 3.48
R75 a_540271_687858.t0 a_540271_687858.n129 3.48
R76 a_540271_687858.n129 a_540271_687858.n105 2.661
R77 a_540271_687858.n129 a_540271_687858.n128 1.972
R78 a_540271_687858.n104 a_540271_687858.n103 1.879
R79 a_540271_687858.n82 a_540271_687858.n80 1.831
R80 a_540271_687858.n122 a_540271_687858.n121 1.484
R81 a_540271_687858.n16 a_540271_687858.n74 1.483
R82 a_540271_687858.n95 a_540271_687858.n94 1.483
R83 a_540271_687858.n120 a_540271_687858.n117 1.483
R84 a_540271_687858.n73 a_540271_687858.n72 1.483
R85 a_540271_687858.n97 a_540271_687858.n91 1.483
R86 a_540271_687858.n86 a_540271_687858.n85 1.482
R87 a_540271_687858.n119 a_540271_687858.n118 1.482
R88 a_540271_687858.n17 a_540271_687858.n75 1.482
R89 a_540271_687858.n0 a_540271_687858.n83 1.482
R90 a_540271_687858.n2 a_540271_687858.n87 1.482
R91 a_540271_687858.n15 a_540271_687858.n92 1.481
R92 a_540271_687858.n114 a_540271_687858.n133 1.481
R93 a_540271_687858.n95 a_540271_687858.n93 1.476
R94 a_540271_687858.n97 a_540271_687858.n90 1.474
R95 a_540271_687858.n15 a_540271_687858.n96 1.393
R96 a_540271_687858.n128 a_540271_687858.n10 0.91
R97 a_540271_687858.n104 a_540271_687858.n14 0.907
R98 a_540271_687858.n9 a_540271_687858.n82 0.907
R99 a_540271_687858.n46 a_540271_687858.n45 0.592
R100 a_540271_687858.n41 a_540271_687858.n131 0.592
R101 a_540271_687858.n76 a_540271_687858.n24 0.545
R102 a_540271_687858.n47 a_540271_687858.n46 0.503
R103 a_540271_687858.n66 a_540271_687858.n89 0.503
R104 a_540271_687858.n64 a_540271_687858.n63 0.503
R105 a_540271_687858.n115 a_540271_687858.n114 0.502
R106 a_540271_687858.n89 a_540271_687858.n88 0.502
R107 a_540271_687858.n63 a_540271_687858.n62 0.502
R108 a_540271_687858.n32 a_540271_687858.n29 0.502
R109 a_540271_687858.n77 a_540271_687858.n76 0.502
R110 a_540271_687858.n42 a_540271_687858.n41 0.502
R111 a_540271_687858.n29 a_540271_687858.n7 0.502
R112 a_540271_687858.n15 a_540271_687858.n95 0.484
R113 a_540271_687858.n133 a_540271_687858.n132 0.483
R114 a_540271_687858.n2 a_540271_687858.n86 0.483
R115 a_540271_687858.n17 a_540271_687858.n16 0.483
R116 a_540271_687858.n16 a_540271_687858.n73 0.482
R117 a_540271_687858.n122 a_540271_687858.n120 0.482
R118 a_540271_687858.n120 a_540271_687858.n119 0.482
R119 a_540271_687858.n82 a_540271_687858.n81 0.464
R120 a_540271_687858.n0 a_540271_687858.n2 0.454
R121 a_540271_687858.n116 a_540271_687858.n122 0.449
R122 a_540271_687858.n67 a_540271_687858.n97 0.448
R123 a_540271_687858.n25 a_540271_687858.n24 0.448
R124 a_540271_687858.n68 a_540271_687858.n71 0.446
R125 a_540271_687858.n45 a_540271_687858.n40 0.446
R126 a_540271_687858.n59 a_540271_687858.n58 0.446
R127 a_540271_687858.n78 a_540271_687858.n17 0.445
R128 a_540271_687858.n23 a_540271_687858.n22 0.425
R129 a_540271_687858.n131 a_540271_687858.n130 0.501
R130 a_540271_687858.n105 a_540271_687858.n104 0.381
R131 a_540271_687858.n8 a_540271_687858.n7 0.202
R132 a_540271_687858.n8 a_540271_687858.n42 0.297
R133 a_540271_687858.n71 a_540271_687858.n9 0.195
R134 a_540271_687858.n3 a_540271_687858.n111 0.136
R135 a_540271_687858.n4 a_540271_687858.n28 0.136
R136 a_540271_687858.n10 a_540271_687858.n123 0.135
R137 a_540271_687858.n6 a_540271_687858.n65 0.12
R138 a_540271_687858.n12 a_540271_687858.n48 0.119
R139 a_540271_687858.n14 a_540271_687858.n98 0.119
R140 a_540271_687858.n127 a_540271_687858.n125 0.107
R141 a_540271_687858.n109 a_540271_687858.n107 0.107
R142 a_540271_687858.n3 a_540271_687858.n113 0.098
R143 a_540271_687858.n10 a_540271_687858.n127 0.098
R144 a_540271_687858.n4 a_540271_687858.n109 0.098
R145 a_540271_687858.n12 a_540271_687858.n6 0.094
R146 a_540271_687858.n14 a_540271_687858.n12 0.094
R147 a_540271_687858.n111 a_540271_687858.n110 0.09
R148 a_540271_687858.n32 a_540271_687858.n30 0.089
R149 a_540271_687858.n65 a_540271_687858.n64 0.088
R150 a_540271_687858.n48 a_540271_687858.n47 0.086
R151 a_540271_687858.n11 a_540271_687858.n1 0.157
R152 a_540271_687858.n13 a_540271_687858.n101 0.084
R153 a_540271_687858.n5 a_540271_687858.n51 0.084
R154 a_540271_687858.n56 a_540271_687858.n54 0.08
R155 a_540271_687858.n36 a_540271_687858.n34 0.08
R156 a_540271_687858.n101 a_540271_687858.n100 0.077
R157 a_540271_687858.n51 a_540271_687858.n50 0.077
R158 a_540271_687858.n22 a_540271_687858.n21 0.076
R159 a_540271_687858.n30 a_540271_687858.t18 6.214
R160 a_540271_687858.n28 a_540271_687858.n27 0.072
R161 a_540271_687858.n58 a_540271_687858.n57 0.056
R162 a_540271_687858.n40 a_540271_687858.n39 0.056
R163 a_540271_687858.n71 a_540271_687858.n70 0.056
R164 a_540271_687858.n67 a_540271_687858.n66 0.046
R165 a_540271_687858.n61 a_540271_687858.n59 0.046
R166 a_540271_687858.n79 a_540271_687858.n78 0.046
R167 a_540271_687858.n116 a_540271_687858.n115 0.046
R168 a_540271_687858.n28 a_540271_687858.n26 0.046
R169 a_540271_687858.n24 a_540271_687858.n23 0.046
R170 a_540271_687858.n62 a_540271_687858.n61 0.045
R171 a_540271_687858.n88 a_540271_687858.n69 0.045
R172 a_540271_687858.n69 a_540271_687858.n68 0.045
R173 a_540271_687858.n123 a_540271_687858.n116 0.044
R174 a_540271_687858.n78 a_540271_687858.n77 0.042
R175 a_540271_687858.n98 a_540271_687858.n67 0.041
R176 a_540271_687858.n61 a_540271_687858.n60 0.029
R177 a_540271_687858.n125 a_540271_687858.n124 0.028
R178 a_540271_687858.n107 a_540271_687858.n106 0.028
R179 a_540271_687858.n32 a_540271_687858.n31 0.028
R180 a_540271_687858.n36 a_540271_687858.n35 0.012
R181 a_540271_687858.n56 a_540271_687858.n55 0.01
R182 a_540271_687858.n36 a_540271_687858.n33 0.01
R183 a_540271_687858.n101 a_540271_687858.n99 0.01
R184 a_540271_687858.n51 a_540271_687858.n49 0.01
R185 a_540271_687858.n58 a_540271_687858.n56 0.004
R186 a_540271_687858.n22 a_540271_687858.n20 0.004
R187 a_540271_687858.n38 a_540271_687858.n44 0.004
R188 a_540271_687858.n38 a_540271_687858.n36 0.002
R189 a_540271_687858.n40 a_540271_687858.n38 0.001
R190 a_540271_687858.n25 a_540271_687858.n19 0.483
R191 a_540271_687858.n19 a_540271_687858.n18 0.483
R192 a_540271_687858.n97 a_540271_687858.n15 0.482
R193 a_540271_687858.n9 a_540271_687858.n79 0.114
R194 a_540271_687858.n10 a_540271_687858.n3 0.095
R195 a_540271_687858.n3 a_540271_687858.n4 0.095
R196 a_540271_687858.n2 a_540271_687858.n84 0.093
R197 a_540271_687858.n6 a_540271_687858.n5 0.085
R198 a_540271_687858.n14 a_540271_687858.n13 0.085
R199 a_540271_687858.n12 a_540271_687858.n11 0.085
R200 a_540271_687858.n34 a_540271_687858.n8 0.081
R201 a_540271_687858.n113 a_540271_687858.t28 5.848
R202 a_540271_687858.n69 a_540271_687858.n0 0.478
R203 vccd1.n248 vccd1.n208 397.746
R204 vccd1.n265 vccd1.n207 394.638
R205 vccd1.n290 vccd1.n266 325.116
R206 vccd1.n247 vccd1.n228 323.618
R207 vccd1.n145 vccd1.n143 246.592
R208 vccd1.n145 vccd1.n144 246.592
R209 vccd1.n298 vccd1.n296 246.592
R210 vccd1.n298 vccd1.n297 246.592
R211 vccd1.n117 vccd1.n115 211.952
R212 vccd1.n113 vccd1.n110 211.952
R213 vccd1.n242 vccd1.t25 205.018
R214 vccd1.n89 vccd1.n21 202.541
R215 vccd1.n53 vccd1.n51 201.034
R216 vccd1.n58 vccd1.n55 201.034
R217 vccd1.n35 vccd1.n34 196.141
R218 vccd1.n35 vccd1.n29 196.141
R219 vccd1.n244 vccd1.n243 185
R220 vccd1.n277 vccd1.n276 185
R221 vccd1.n1 vccd1.t21 173.631
R222 vccd1.n73 vccd1.t10 172.101
R223 vccd1.n90 vccd1.n13 127.427
R224 vccd1.n82 vccd1.n44 125.545
R225 vccd1.n206 vccd1.n205 116.309
R226 vccd1.n295 vccd1.t23 116.305
R227 vccd1.t25 vccd1.n239 116.305
R228 vccd1.n227 vccd1.n226 116.173
R229 vccd1.t77 vccd1.t14 110.367
R230 vccd1.t2 vccd1.n157 109.669
R231 vccd1.t35 vccd1.n202 109.145
R232 vccd1.t6 vccd1.t68 105.477
R233 vccd1.t74 vccd1.t27 105.477
R234 vccd1.n102 vccd1.n93 103.529
R235 vccd1.n118 vccd1.n113 97.129
R236 vccd1.n118 vccd1.n117 97.129
R237 vccd1.n224 vccd1.t18 96.397
R238 vccd1.n278 vccd1.t4 96.222
R239 vccd1.n251 vccd1.t6 93.253
R240 vccd1.n158 vccd1.t2 92.904
R241 vccd1.n65 vccd1.n63 92.611
R242 vccd1.n203 vccd1.t35 89.935
R243 vccd1.n245 vccd1.t31 89.761
R244 vccd1.n72 vccd1.n71 87.905
R245 vccd1.n59 vccd1.n53 86.211
R246 vccd1.n59 vccd1.n58 86.211
R247 vccd1.n100 vccd1.n99 82.144
R248 vccd1.t31 vccd1.n244 65.487
R249 vccd1.t4 vccd1.n277 59.375
R250 vccd1.n277 vccd1.t77 46.102
R251 vccd1.n244 vccd1.t74 44.88
R252 vccd1.n47 vccd1.t47 37.479
R253 vccd1.n161 vccd1.n160 36.407
R254 vccd1.n203 vccd1.n201 14.843
R255 vccd1.n278 vccd1.t71 14.145
R256 vccd1.n224 vccd1.t93 13.97
R257 vccd1.n22 vccd1.t0 13.003
R258 vccd1.t79 vccd1.n158 12.573
R259 vccd1.t27 vccd1.n242 10.827
R260 vccd1.n225 vccd1.n224 9.3
R261 vccd1.n247 vccd1.n246 9.3
R262 vccd1.n246 vccd1.n245 9.3
R263 vccd1.n290 vccd1.n279 9.3
R264 vccd1.n279 vccd1.n278 9.3
R265 vccd1.n204 vccd1.n203 9.3
R266 vccd1.n264 vccd1.n252 9.3
R267 vccd1.n252 vccd1.n251 9.3
R268 vccd1.n250 vccd1.n249 8.457
R269 vccd1.n283 vccd1.t86 8.382
R270 vccd1.n198 vccd1.t78 8.382
R271 vccd1.n288 vccd1.t88 8.382
R272 vccd1.n210 vccd1.t92 8.348
R273 vccd1.n213 vccd1.t91 8.347
R274 vccd1.n214 vccd1.t84 8.347
R275 vccd1.n168 vccd1.t112 8.095
R276 vccd1.n166 vccd1.t81 8.095
R277 vccd1.n171 vccd1.t89 8.095
R278 vccd1.n155 vccd1.t75 8.087
R279 vccd1.n176 vccd1.t85 8.087
R280 vccd1.n177 vccd1.t96 8.087
R281 vccd1.n136 vccd1.t61 7.864
R282 vccd1.n300 vccd1.t44 7.672
R283 vccd1.n135 vccd1.t42 7.669
R284 vccd1.n302 vccd1.t26 7.669
R285 vccd1.n105 vccd1.t8 6.884
R286 vccd1.n91 vccd1.n4 6.4
R287 vccd1.n91 vccd1.n6 6.4
R288 vccd1.n89 vccd1.n36 6.4
R289 vccd1.n89 vccd1.n35 6.4
R290 vccd1.n87 vccd1.n86 6.4
R291 vccd1.n87 vccd1.n84 6.4
R292 vccd1.n81 vccd1.n79 6.4
R293 vccd1.n81 vccd1.n78 6.4
R294 vccd1.n65 vccd1.n46 6.4
R295 vccd1.n65 vccd1.n59 6.4
R296 vccd1.n119 vccd1.n118 6.4
R297 vccd1.n119 vccd1.n104 6.4
R298 vccd1.t14 vccd1.n275 5.937
R299 vccd1.n136 vccd1.t28 5.794
R300 vccd1.n300 vccd1.t63 5.788
R301 vccd1.n302 vccd1.t64 5.787
R302 vccd1.n135 vccd1.t46 5.787
R303 vccd1.n124 vccd1.t12 5.775
R304 vccd1.n318 vccd1.t5 5.771
R305 vccd1.n316 vccd1.t20 5.771
R306 vccd1.n122 vccd1.t59 5.771
R307 vccd1.n155 vccd1.t94 5.769
R308 vccd1.n176 vccd1.t100 5.769
R309 vccd1.n177 vccd1.t106 5.769
R310 vccd1.n168 vccd1.t102 5.769
R311 vccd1.n166 vccd1.t110 5.769
R312 vccd1.n171 vccd1.t76 5.769
R313 vccd1.n153 vccd1.t105 5.766
R314 vccd1.n173 vccd1.t113 5.766
R315 vccd1.n175 vccd1.t83 5.766
R316 vccd1.n307 vccd1.t65 5.763
R317 vccd1.n128 vccd1.t41 5.761
R318 vccd1.n313 vccd1.t7 5.759
R319 vccd1.n311 vccd1.t55 5.759
R320 vccd1.n126 vccd1.t13 5.757
R321 vccd1.n305 vccd1.t19 5.756
R322 vccd1.n323 vccd1.t56 5.75
R323 vccd1.n134 vccd1.t58 5.749
R324 vccd1.n131 vccd1.t57 5.748
R325 vccd1.n149 vccd1.t62 5.746
R326 vccd1.n147 vccd1.t43 5.746
R327 vccd1.n321 vccd1.t24 5.746
R328 vccd1.n102 vccd1.t49 5.717
R329 vccd1.n119 vccd1.t9 5.717
R330 vccd1.n3 vccd1.t39 5.713
R331 vccd1.n64 vccd1.t48 5.713
R332 vccd1.n75 vccd1.t11 5.713
R333 vccd1.n87 vccd1.t115 5.713
R334 vccd1.n14 vccd1.t1 5.713
R335 vccd1.n0 vccd1.t22 5.713
R336 vccd1.n88 vccd1.t16 5.713
R337 vccd1.n87 vccd1.t34 5.713
R338 vccd1.n80 vccd1.t40 5.713
R339 vccd1.n45 vccd1.t116 5.713
R340 vccd1.n280 vccd1.t95 5.713
R341 vccd1.n254 vccd1.t82 5.713
R342 vccd1.n253 vccd1.t67 5.713
R343 vccd1.n257 vccd1.t80 5.713
R344 vccd1.n256 vccd1.t114 5.713
R345 vccd1.n211 vccd1.t103 5.713
R346 vccd1.n284 vccd1.t97 5.713
R347 vccd1.n282 vccd1.t72 5.713
R348 vccd1.n188 vccd1.t107 5.713
R349 vccd1.n215 vccd1.t99 5.713
R350 vccd1.n189 vccd1.t111 5.713
R351 vccd1.n195 vccd1.t87 5.713
R352 vccd1.n197 vccd1.t109 5.713
R353 vccd1.n317 vccd1.t38 5.713
R354 vccd1.n310 vccd1.t30 5.713
R355 vccd1.n304 vccd1.t51 5.713
R356 vccd1.n129 vccd1.t32 5.713
R357 vccd1.n125 vccd1.t17 5.713
R358 vccd1.n127 vccd1.t3 5.713
R359 vccd1.n306 vccd1.t50 5.713
R360 vccd1.n312 vccd1.t29 5.713
R361 vccd1.n315 vccd1.t36 5.713
R362 vccd1.n322 vccd1.t15 5.713
R363 vccd1.n133 vccd1.t37 5.713
R364 vccd1.n123 vccd1.t45 5.713
R365 vccd1.n148 vccd1.t53 5.713
R366 vccd1.n121 vccd1.t54 5.713
R367 vccd1.n146 vccd1.t52 5.713
R368 vccd1.n320 vccd1.t60 5.713
R369 vccd1.n167 vccd1.t69 5.713
R370 vccd1.n152 vccd1.t101 5.713
R371 vccd1.n165 vccd1.t90 5.713
R372 vccd1.n172 vccd1.t108 5.713
R373 vccd1.n170 vccd1.t98 5.713
R374 vccd1.n174 vccd1.t70 5.713
R375 vccd1.n209 vccd1.t104 5.713
R376 vccd1.n287 vccd1.t73 5.713
R377 vccd1.n227 vccd1.n225 5.528
R378 vccd1.n206 vccd1.n204 5.524
R379 vccd1.t79 vccd1.n162 4.894
R380 vccd1.n301 vccd1.n299 4.425
R381 vccd1.n324 vccd1.n298 4.425
R382 vccd1.n150 vccd1.n145 4.425
R383 vccd1.n138 vccd1.n137 4.425
R384 vccd1.n179 vccd1.n178 4.1
R385 vccd1.n185 vccd1.n184 4.085
R386 vccd1.n200 vccd1.n186 4.085
R387 vccd1.n219 vccd1.n218 3.744
R388 vccd1.n156 vccd1.n154 3.649
R389 vccd1.n290 vccd1.n206 3.606
R390 vccd1.n247 vccd1.n227 3.602
R391 vccd1.n34 vccd1.n32 3.388
R392 vccd1.n29 vccd1.n27 3.388
R393 vccd1.n21 vccd1.n16 3.388
R394 vccd1.n169 vccd1.n164 3.368
R395 vccd1.n255 vccd1.n253 2.674
R396 vccd1.n258 vccd1.n256 2.673
R397 vccd1.n190 vccd1.n188 2.668
R398 vccd1.n285 vccd1.n284 2.653
R399 vccd1.n196 vccd1.n195 2.653
R400 vccd1.n281 vccd1.n280 2.653
R401 vccd1.n153 vccd1.n152 2.386
R402 vccd1.n173 vccd1.n172 2.386
R403 vccd1.n175 vccd1.n174 2.386
R404 vccd1.n168 vccd1.n167 2.367
R405 vccd1.n166 vccd1.n165 2.367
R406 vccd1.n171 vccd1.n170 2.367
R407 vccd1.n163 vccd1.t79 2.365
R408 vccd1.n149 vccd1.n148 2.305
R409 vccd1.n134 vccd1.n133 2.297
R410 vccd1.n128 vccd1.n127 2.275
R411 vccd1.n124 vccd1.n123 2.235
R412 vccd1.n323 vccd1.n322 2.094
R413 vccd1.n147 vccd1.n146 2.091
R414 vccd1.n321 vccd1.n320 2.091
R415 vccd1.n130 vccd1.n129 2.084
R416 vccd1.n305 vccd1.n304 2.068
R417 vccd1.n313 vccd1.n312 2.065
R418 vccd1.n311 vccd1.n310 2.065
R419 vccd1.n126 vccd1.n125 2.062
R420 vccd1.n307 vccd1.n306 2.049
R421 vccd1.n316 vccd1.n315 2.03
R422 vccd1.n122 vccd1.n121 2.03
R423 vccd1.n318 vccd1.n317 2.03
R424 vccd1.n161 vccd1.n159 1.976
R425 vccd1.n293 vccd1.n169 1.034
R426 vccd1.t93 vccd1.n223 0.873
R427 vccd1.n292 vccd1.n185 0.846
R428 vccd1.n291 vccd1.n200 0.809
R429 vccd1.n37 vccd1.t33 0.764
R430 vccd1.n157 vccd1.t66 0.698
R431 vccd1.n291 vccd1.n290 0.65
R432 vccd1.n163 vccd1.n156 0.603
R433 vccd1.n169 vccd1.n163 0.596
R434 vccd1.n327 vccd1.n325 0.587
R435 vccd1.n264 vccd1.n250 0.534
R436 vccd1.n180 vccd1.n179 0.508
R437 vccd1.n183 vccd1.n182 0.504
R438 vccd1.n200 vccd1.n194 0.467
R439 vccd1.t79 vccd1.n161 0.447
R440 vccd1.n308 vccd1.n303 0.325
R441 vccd1.n319 vccd1.n314 0.317
R442 vccd1.n139 vccd1.n138 0.307
R443 vccd1.n142 vccd1.n141 0.299
R444 vccd1.n324 vccd1.n319 0.293
R445 vccd1.n151 vccd1.n142 0.29
R446 vccd1.n175 vccd1.n173 0.25
R447 vccd1.n177 vccd1.n176 0.25
R448 vccd1.n102 vccd1.n100 0.25
R449 vccd1.n309 vccd1.n308 0.243
R450 vccd1.n263 vccd1.n261 0.231
R451 vccd1.n140 vccd1.n139 0.229
R452 vccd1.n222 vccd1.n220 0.229
R453 vccd1.n289 vccd1.n286 0.227
R454 vccd1.n169 vccd1.n166 0.196
R455 vccd1.n139 vccd1.n134 0.176
R456 vccd1.n308 vccd1.n305 0.176
R457 vccd1.n141 vccd1.n128 0.176
R458 vccd1.n314 vccd1.n311 0.176
R459 vccd1.n142 vccd1.n124 0.176
R460 vccd1.n319 vccd1.n318 0.176
R461 vccd1.n150 vccd1.n149 0.176
R462 vccd1.n324 vccd1.n321 0.176
R463 vccd1.n138 vccd1.n136 0.169
R464 vccd1.n220 vccd1.n219 0.169
R465 vccd1.n303 vccd1.n302 0.166
R466 vccd1.n248 vccd1.n247 0.151
R467 vccd1.n264 vccd1.n248 0.151
R468 vccd1.n265 vccd1.n264 0.15
R469 vccd1.n290 vccd1.n265 0.149
R470 vccd1.n326 vccd1 0.141
R471 vccd1.n293 vccd1.n292 0.13
R472 vccd1.n283 vccd1.n282 0.13
R473 vccd1.n198 vccd1.n197 0.13
R474 vccd1.n288 vccd1.n287 0.13
R475 vccd1.n325 vccd1.n120 0.123
R476 vccd1.n258 vccd1.n257 0.116
R477 vccd1.n255 vccd1.n254 0.115
R478 vccd1.n190 vccd1.n189 0.111
R479 vccd1.n212 vccd1.n211 0.111
R480 vccd1.n216 vccd1.n215 0.111
R481 vccd1.n91 vccd1.n0 0.109
R482 vccd1.n81 vccd1.n80 0.109
R483 vccd1.n91 vccd1.n3 0.109
R484 vccd1.n81 vccd1.n75 0.108
R485 vccd1.n294 vccd1.n293 0.107
R486 vccd1.n328 vccd1.n327 0.094
R487 vccd1.n326 vccd1 0.08
R488 vccd1.n314 vccd1.n309 0.077
R489 vccd1.n141 vccd1.n140 0.072
R490 vccd1.n292 vccd1.n291 0.067
R491 vccd1.n210 vccd1.n209 0.066
R492 vccd1.n179 vccd1.n177 0.066
R493 vccd1.n200 vccd1.n199 0.066
R494 vccd1.n120 vccd1.n119 0.064
R495 vccd1.n325 vccd1.n324 0.064
R496 vccd1.n183 vccd1.n171 0.063
R497 vccd1.n324 vccd1.n323 0.06
R498 vccd1.n219 vccd1.n217 0.059
R499 vccd1.n181 vccd1.n175 0.059
R500 vccd1.n192 vccd1.n191 0.057
R501 vccd1.n314 vccd1.n313 0.056
R502 vccd1.n142 vccd1.n122 0.056
R503 vccd1.n319 vccd1.n316 0.056
R504 vccd1.n150 vccd1.n147 0.056
R505 vccd1.n156 vccd1.n155 0.056
R506 vccd1.n169 vccd1.n168 0.053
R507 vccd1.n120 vccd1.n103 0.052
R508 vccd1.n301 vccd1.n300 0.052
R509 vccd1.n139 vccd1.n132 0.051
R510 vccd1.n308 vccd1.n307 0.051
R511 vccd1.n141 vccd1.n126 0.051
R512 vccd1.n290 vccd1.n289 0.051
R513 vccd1.n328 vccd1 0.051
R514 vccd1.n163 vccd1.n153 0.049
R515 vccd1.n138 vccd1.n135 0.048
R516 vccd1.n327 vccd1 0.048
R517 vccd1 vccd1.n326 0.047
R518 vccd1.n264 vccd1.n263 0.046
R519 vccd1.n247 vccd1.n222 0.046
R520 vccd1 vccd1.n328 0.045
R521 vccd1.n89 vccd1.n87 0.043
R522 vccd1.n296 vccd1.n295 0.041
R523 vccd1.n275 vccd1.n267 0.041
R524 vccd1.n275 vccd1.n268 0.041
R525 vccd1.n275 vccd1.n269 0.041
R526 vccd1.n275 vccd1.n272 0.041
R527 vccd1.n239 vccd1.n237 0.041
R528 vccd1.n239 vccd1.n235 0.041
R529 vccd1.n239 vccd1.n236 0.041
R530 vccd1.n239 vccd1.n238 0.041
R531 vccd1.n242 vccd1.n234 0.041
R532 vccd1.n242 vccd1.n233 0.041
R533 vccd1.n242 vccd1.n232 0.041
R534 vccd1.n242 vccd1.n229 0.041
R535 vccd1.n103 vccd1.n91 0.035
R536 vccd1.n90 vccd1.n89 0.029
R537 vccd1.n91 vccd1.n90 0.029
R538 vccd1.n87 vccd1.n82 0.028
R539 vccd1.n82 vccd1.n81 0.028
R540 vccd1.n65 vccd1.n64 0.023
R541 vccd1.n65 vccd1.n45 0.023
R542 vccd1.n231 vccd1.n230 0.022
R543 vccd1.n242 vccd1.n231 0.022
R544 vccd1.n271 vccd1.n270 0.022
R545 vccd1.n275 vccd1.n271 0.022
R546 vccd1.n242 vccd1.n241 0.022
R547 vccd1.n275 vccd1.n274 0.022
R548 vccd1.n72 vccd1.n65 0.02
R549 vccd1.n81 vccd1.n72 0.02
R550 vccd1.n274 vccd1.n273 0.02
R551 vccd1.n241 vccd1.n240 0.02
R552 vccd1.n222 vccd1.n221 0.02
R553 vccd1.n53 vccd1.n52 0.02
R554 vccd1.n58 vccd1.n57 0.02
R555 vccd1.n57 vccd1.n56 0.02
R556 vccd1.n63 vccd1.n62 0.02
R557 vccd1.n93 vccd1.n92 0.017
R558 vccd1.n113 vccd1.n112 0.017
R559 vccd1.n112 vccd1.n111 0.017
R560 vccd1.n117 vccd1.n116 0.017
R561 vccd1.n103 vccd1.n102 0.016
R562 vccd1.n185 vccd1.n183 0.015
R563 vccd1.n51 vccd1.n50 0.015
R564 vccd1.n50 vccd1.n49 0.015
R565 vccd1.n115 vccd1.n114 0.015
R566 vccd1.n55 vccd1.n54 0.015
R567 vccd1.n110 vccd1.n109 0.015
R568 vccd1.n109 vccd1.n108 0.015
R569 vccd1.n181 vccd1.n180 0.014
R570 vccd1.n182 vccd1.n181 0.014
R571 vccd1.n324 vccd1.n294 0.014
R572 vccd1.n97 vccd1.n96 0.01
R573 vccd1.n98 vccd1.n97 0.01
R574 vccd1.n95 vccd1.n94 0.01
R575 vccd1.n98 vccd1.n95 0.01
R576 vccd1.n99 vccd1.n98 0.01
R577 vccd1.n67 vccd1.n66 0.009
R578 vccd1.n70 vccd1.n67 0.009
R579 vccd1.n69 vccd1.n68 0.009
R580 vccd1.n70 vccd1.n69 0.009
R581 vccd1.n71 vccd1.n70 0.009
R582 vccd1.n89 vccd1.n14 0.008
R583 vccd1.n89 vccd1.n88 0.008
R584 vccd1.n32 vccd1.n31 0.008
R585 vccd1.n31 vccd1.n30 0.008
R586 vccd1.n27 vccd1.n26 0.008
R587 vccd1.n16 vccd1.n15 0.008
R588 vccd1.n9 vccd1.n8 0.006
R589 vccd1.n12 vccd1.n9 0.006
R590 vccd1.n11 vccd1.n10 0.006
R591 vccd1.n12 vccd1.n11 0.006
R592 vccd1.n40 vccd1.n39 0.006
R593 vccd1.n43 vccd1.n40 0.006
R594 vccd1.n42 vccd1.n41 0.006
R595 vccd1.n43 vccd1.n42 0.006
R596 vccd1.n44 vccd1.n43 0.006
R597 vccd1.n13 vccd1.n12 0.006
R598 vccd1.n303 vccd1.n301 0.005
R599 vccd1.n132 vccd1.n131 0.004
R600 vccd1.n89 vccd1.n25 0.003
R601 vccd1.n89 vccd1.n24 0.003
R602 vccd1.n87 vccd1.n85 0.003
R603 vccd1.n87 vccd1.n83 0.003
R604 vccd1.n81 vccd1.n77 0.003
R605 vccd1.n81 vccd1.n76 0.003
R606 vccd1.n65 vccd1.n48 0.003
R607 vccd1.n48 vccd1.n47 0.003
R608 vccd1.n65 vccd1.n60 0.003
R609 vccd1.n65 vccd1.n61 0.003
R610 vccd1.n81 vccd1.n74 0.003
R611 vccd1.n74 vccd1.n73 0.003
R612 vccd1.n87 vccd1.n38 0.003
R613 vccd1.n38 vccd1.n37 0.003
R614 vccd1.n89 vccd1.n23 0.003
R615 vccd1.n23 vccd1.n22 0.003
R616 vccd1.n91 vccd1.n2 0.003
R617 vccd1.n2 vccd1.n1 0.003
R618 vccd1.n102 vccd1.n101 0.003
R619 vccd1.n119 vccd1.n106 0.003
R620 vccd1.n106 vccd1.n105 0.003
R621 vccd1.n119 vccd1.n107 0.003
R622 vccd1.n91 vccd1.n5 0.003
R623 vccd1.n91 vccd1.n7 0.003
R624 vccd1.n194 vccd1.n193 0.003
R625 vccd1.n193 vccd1.n192 0.002
R626 vccd1.n131 vccd1.n130 0.001
R627 vccd1.n151 vccd1.n150 0.001
R628 vccd1.n260 vccd1.n259 0.001
R629 vccd1.n34 vccd1.n33 0.001
R630 vccd1.n29 vccd1.n28 0.001
R631 vccd1.n21 vccd1.n20 0.001
R632 vccd1.n20 vccd1.n19 0.001
R633 vccd1.n294 vccd1.n151 0.001
R634 vccd1.n286 vccd1.n285 0.001
R635 vccd1.n199 vccd1.n196 0.001
R636 vccd1.n289 vccd1.n281 0.001
R637 vccd1.n286 vccd1.n283 0.001
R638 vccd1.n289 vccd1.n288 0.001
R639 vccd1.n199 vccd1.n198 0.001
R640 vccd1.n220 vccd1.n213 0.001
R641 vccd1.n217 vccd1.n214 0.001
R642 vccd1.n263 vccd1.n262 0.001
R643 vccd1.n191 vccd1.n187 0.001
R644 vccd1.n261 vccd1.n258 0.001
R645 vccd1.n263 vccd1.n255 0.001
R646 vccd1.n220 vccd1.n212 0.001
R647 vccd1.n217 vccd1.n216 0.001
R648 vccd1.n191 vccd1.n190 0.001
R649 vccd1.n222 vccd1.n210 0.001
R650 vccd1.n18 vccd1.n17 0.001
R651 vccd1.n19 vccd1.n18 0.001
R652 vccd1.n261 vccd1.n260 0.001
R653 a_537154_685355.n39 a_537154_685355.t67 271.866
R654 a_537154_685355.n18 a_537154_685355.t56 271.859
R655 a_537154_685355.n15 a_537154_685355.t58 135.085
R656 a_537154_685355.n248 a_537154_685355.t54 135.079
R657 a_537154_685355.n54 a_537154_685355.t70 135.078
R658 a_537154_685355.n197 a_537154_685355.t57 135.077
R659 a_537154_685355.n212 a_537154_685355.t53 135.077
R660 a_537154_685355.n179 a_537154_685355.t71 135.077
R661 a_537154_685355.n25 a_537154_685355.t38 135.077
R662 a_537154_685355.n139 a_537154_685355.t64 135.077
R663 a_537154_685355.n170 a_537154_685355.t62 135.077
R664 a_537154_685355.n172 a_537154_685355.t49 135.077
R665 a_537154_685355.n142 a_537154_685355.t52 135.077
R666 a_537154_685355.n6 a_537154_685355.t33 135.077
R667 a_537154_685355.n47 a_537154_685355.t40 135.077
R668 a_537154_685355.n137 a_537154_685355.t66 135.077
R669 a_537154_685355.n167 a_537154_685355.t63 135.077
R670 a_537154_685355.n175 a_537154_685355.t47 135.077
R671 a_537154_685355.n145 a_537154_685355.t50 135.077
R672 a_537154_685355.n243 a_537154_685355.t32 135.077
R673 a_537154_685355.n153 a_537154_685355.t51 135.076
R674 a_537154_685355.n155 a_537154_685355.t41 135.076
R675 a_537154_685355.n9 a_537154_685355.t43 135.076
R676 a_537154_685355.n49 a_537154_685355.t59 135.076
R677 a_537154_685355.n149 a_537154_685355.t55 135.076
R678 a_537154_685355.n161 a_537154_685355.t39 135.076
R679 a_537154_685355.n246 a_537154_685355.t42 135.076
R680 a_537154_685355.n19 a_537154_685355.t60 135.076
R681 a_537154_685355.n120 a_537154_685355.t45 135.076
R682 a_537154_685355.n191 a_537154_685355.t34 135.076
R683 a_537154_685355.n206 a_537154_685355.t69 135.076
R684 a_537154_685355.n126 a_537154_685355.t37 135.076
R685 a_537154_685355.n0 a_537154_685355.t46 135.076
R686 a_537154_685355.n42 a_537154_685355.t61 135.076
R687 a_537154_685355.n115 a_537154_685355.t48 135.076
R688 a_537154_685355.n183 a_537154_685355.t35 135.076
R689 a_537154_685355.n215 a_537154_685355.t65 135.076
R690 a_537154_685355.n132 a_537154_685355.t36 135.076
R691 a_537154_685355.n237 a_537154_685355.t44 135.076
R692 a_537154_685355.n187 a_537154_685355.t68 135.056
R693 a_537154_685355.n74 a_537154_685355.t14 5.767
R694 a_537154_685355.n78 a_537154_685355.t10 5.767
R695 a_537154_685355.n80 a_537154_685355.t26 5.765
R696 a_537154_685355.n61 a_537154_685355.t8 5.765
R697 a_537154_685355.n58 a_537154_685355.t17 5.757
R698 a_537154_685355.n59 a_537154_685355.t13 5.756
R699 a_537154_685355.n92 a_537154_685355.t9 5.713
R700 a_537154_685355.n95 a_537154_685355.t18 5.713
R701 a_537154_685355.n64 a_537154_685355.t12 5.713
R702 a_537154_685355.n65 a_537154_685355.t7 5.713
R703 a_537154_685355.n69 a_537154_685355.t23 5.713
R704 a_537154_685355.n110 a_537154_685355.t19 5.713
R705 a_537154_685355.n106 a_537154_685355.t24 5.713
R706 a_537154_685355.n105 a_537154_685355.t27 5.713
R707 a_537154_685355.n85 a_537154_685355.t11 5.713
R708 a_537154_685355.n88 a_537154_685355.t22 5.713
R709 a_537154_685355.n89 a_537154_685355.t20 5.713
R710 a_537154_685355.n62 a_537154_685355.t16 5.713
R711 a_537154_685355.n82 a_537154_685355.t21 5.713
R712 a_537154_685355.n102 a_537154_685355.t15 5.713
R713 a_537154_685355.n99 a_537154_685355.t25 5.713
R714 a_537154_685355.n221 a_537154_685355.t0 3.482
R715 a_537154_685355.n236 a_537154_685355.t2 3.48
R716 a_537154_685355.n234 a_537154_685355.t29 3.48
R717 a_537154_685355.n231 a_537154_685355.t1 3.48
R718 a_537154_685355.n229 a_537154_685355.t4 3.48
R719 a_537154_685355.n226 a_537154_685355.t3 3.48
R720 a_537154_685355.n225 a_537154_685355.t5 3.48
R721 a_537154_685355.n29 a_537154_685355.n28 3.439
R722 a_537154_685355.n39 a_537154_685355.n38 3.422
R723 a_537154_685355.n212 a_537154_685355.n211 2.948
R724 a_537154_685355.n55 a_537154_685355.n54 2.827
R725 a_537154_685355.n249 a_537154_685355.n248 2.765
R726 a_537154_685355.n57 a_537154_685355.n15 2.712
R727 a_537154_685355.n226 a_537154_685355.n225 2.695
R728 a_537154_685355.n231 a_537154_685355.n230 2.678
R729 a_537154_685355.n236 a_537154_685355.n235 2.629
R730 a_537154_685355.n107 a_537154_685355.n105 2.61
R731 a_537154_685355.n66 a_537154_685355.n64 2.609
R732 a_537154_685355.n93 a_537154_685355.n92 2.571
R733 a_537154_685355.n100 a_537154_685355.n99 2.566
R734 a_537154_685355.n208 a_537154_685355.t28 2.419
R735 a_537154_685355.n211 a_537154_685355.t30 2.412
R736 a_537154_685355.n55 a_537154_685355.t31 2.407
R737 a_537154_685355.n62 a_537154_685355.n61 2.37
R738 a_537154_685355.n90 a_537154_685355.n88 2.35
R739 a_537154_685355.n83 a_537154_685355.n82 2.318
R740 a_537154_685355.n228 a_537154_685355.n227 1.98
R741 a_537154_685355.n222 a_537154_685355.n221 1.966
R742 a_537154_685355.n75 a_537154_685355.n74 1.869
R743 a_537154_685355.n233 a_537154_685355.n232 1.856
R744 a_537154_685355.n215 a_537154_685355.n214 1.819
R745 a_537154_685355.n206 a_537154_685355.n205 1.818
R746 a_537154_685355.n247 a_537154_685355.n246 1.818
R747 a_537154_685355.n154 a_537154_685355.n153 1.817
R748 a_537154_685355.n116 a_537154_685355.n115 1.817
R749 a_537154_685355.n207 a_537154_685355.n206 1.817
R750 a_537154_685355.n49 a_537154_685355.n48 1.817
R751 a_537154_685355.n150 a_537154_685355.n149 1.817
R752 a_537154_685355.n162 a_537154_685355.n161 1.817
R753 a_537154_685355.n50 a_537154_685355.n49 1.817
R754 a_537154_685355.n10 a_537154_685355.n9 1.817
R755 a_537154_685355.n156 a_537154_685355.n155 1.817
R756 a_537154_685355.n97 a_537154_685355.n96 1.817
R757 a_537154_685355.n216 a_537154_685355.n215 1.816
R758 a_537154_685355.n184 a_537154_685355.n183 1.816
R759 a_537154_685355.n238 a_537154_685355.n237 1.816
R760 a_537154_685355.n43 a_537154_685355.n42 1.816
R761 a_537154_685355.n1 a_537154_685355.n0 1.816
R762 a_537154_685355.n192 a_537154_685355.n191 1.816
R763 a_537154_685355.n20 a_537154_685355.n19 1.816
R764 a_537154_685355.n246 a_537154_685355.n245 1.816
R765 a_537154_685355.n9 a_537154_685355.n8 1.816
R766 a_537154_685355.n48 a_537154_685355.n47 1.814
R767 a_537154_685355.n171 a_537154_685355.n170 1.814
R768 a_537154_685355.n168 a_537154_685355.n167 1.813
R769 a_537154_685355.n244 a_537154_685355.n243 1.813
R770 a_537154_685355.n176 a_537154_685355.n175 1.813
R771 a_537154_685355.n7 a_537154_685355.n6 1.813
R772 a_537154_685355.n26 a_537154_685355.n25 1.813
R773 a_537154_685355.n214 a_537154_685355.n212 1.812
R774 a_537154_685355.n180 a_537154_685355.n179 1.811
R775 a_537154_685355.n173 a_537154_685355.n172 1.811
R776 a_537154_685355.n138 a_537154_685355.n137 1.809
R777 a_537154_685355.n146 a_537154_685355.n145 1.809
R778 a_537154_685355.n143 a_537154_685355.n142 1.809
R779 a_537154_685355.n47 a_537154_685355.n46 1.808
R780 a_537154_685355.n140 a_537154_685355.n139 1.807
R781 a_537154_685355.n54 a_537154_685355.n53 1.806
R782 a_537154_685355.n248 a_537154_685355.n247 1.805
R783 a_537154_685355.n104 a_537154_685355.n103 1.8
R784 a_537154_685355.n188 a_537154_685355.n187 1.766
R785 a_537154_685355.n191 a_537154_685355.n190 1.727
R786 a_537154_685355.n183 a_537154_685355.n182 1.727
R787 a_537154_685355.n133 a_537154_685355.n132 1.727
R788 a_537154_685355.n127 a_537154_685355.n126 1.727
R789 a_537154_685355.n121 a_537154_685355.n120 1.727
R790 a_537154_685355.n81 a_537154_685355.n80 1.723
R791 a_537154_685355.n25 a_537154_685355.n24 1.722
R792 a_537154_685355.n243 a_537154_685355.n242 1.722
R793 a_537154_685355.n6 a_537154_685355.n5 1.722
R794 a_537154_685355.n198 a_537154_685355.n197 1.722
R795 a_537154_685355.n15 a_537154_685355.n14 1.705
R796 a_537154_685355.n87 a_537154_685355.n86 1.669
R797 a_537154_685355.n70 a_537154_685355.n68 1.641
R798 a_537154_685355.n111 a_537154_685355.n109 1.633
R799 a_537154_685355.n36 a_537154_685355.n35 1.505
R800 a_537154_685355.n18 a_537154_685355.n17 1.505
R801 a_537154_685355.n56 a_537154_685355.n39 1.011
R802 a_537154_685355.n244 a_537154_685355.n236 0.629
R803 a_537154_685355.n70 a_537154_685355.n69 0.592
R804 a_537154_685355.n111 a_537154_685355.n110 0.588
R805 a_537154_685355.n221 a_537154_685355.n220 0.58
R806 a_537154_685355.n233 a_537154_685355.n112 0.552
R807 a_537154_685355.n230 a_537154_685355.n146 0.546
R808 a_537154_685355.n232 a_537154_685355.n136 0.546
R809 a_537154_685355.n227 a_537154_685355.n166 0.545
R810 a_537154_685355.n224 a_537154_685355.n176 0.534
R811 a_537154_685355.n63 a_537154_685355.n62 0.517
R812 a_537154_685355.n105 a_537154_685355.n104 0.462
R813 a_537154_685355.n144 a_537154_685355.n143 0.449
R814 a_537154_685355.n131 a_537154_685355.n130 0.449
R815 a_537154_685355.n204 a_537154_685355.n203 0.449
R816 a_537154_685355.n125 a_537154_685355.n124 0.449
R817 a_537154_685355.n169 a_537154_685355.n168 0.449
R818 a_537154_685355.n140 a_537154_685355.n138 0.449
R819 a_537154_685355.n163 a_537154_685355.n160 0.448
R820 a_537154_685355.n207 a_537154_685355.n196 0.448
R821 a_537154_685355.n202 a_537154_685355.n201 0.448
R822 a_537154_685355.n173 a_537154_685355.n171 0.448
R823 a_537154_685355.n141 a_537154_685355.n140 0.448
R824 a_537154_685355.n157 a_537154_685355.n154 0.448
R825 a_537154_685355.n174 a_537154_685355.n173 0.448
R826 a_537154_685355.n217 a_537154_685355.n207 0.448
R827 a_537154_685355.n214 a_537154_685355.n213 0.421
R828 a_537154_685355.n119 a_537154_685355.n118 0.42
R829 a_537154_685355.n154 a_537154_685355.n152 0.42
R830 a_537154_685355.n193 a_537154_685355.n186 0.42
R831 a_537154_685355.n88 a_537154_685355.n87 0.407
R832 a_537154_685355.n234 a_537154_685355.n233 0.402
R833 a_537154_685355.n82 a_537154_685355.n81 0.386
R834 a_537154_685355.n229 a_537154_685355.n228 0.332
R835 a_537154_685355.n224 a_537154_685355.n223 0.33
R836 a_537154_685355.n61 a_537154_685355.n60 0.258
R837 a_537154_685355.n60 a_537154_685355.n58 0.246
R838 a_537154_685355.n80 a_537154_685355.n79 0.246
R839 a_537154_685355.n108 a_537154_685355.n91 0.216
R840 a_537154_685355.n209 a_537154_685355.n208 0.159
R841 a_537154_685355.n210 a_537154_685355.n209 0.141
R842 a_537154_685355.n57 a_537154_685355.n56 0.14
R843 a_537154_685355.n56 a_537154_685355.n55 0.127
R844 a_537154_685355.n111 a_537154_685355.n70 0.125
R845 a_537154_685355.n66 a_537154_685355.n65 0.123
R846 a_537154_685355.n107 a_537154_685355.n106 0.122
R847 a_537154_685355.n98 a_537154_685355.n97 0.121
R848 a_537154_685355.n76 a_537154_685355.n75 0.119
R849 a_537154_685355.n77 a_537154_685355.n76 0.118
R850 a_537154_685355.n90 a_537154_685355.n89 0.114
R851 a_537154_685355.n112 a_537154_685355.n111 0.114
R852 a_537154_685355.n96 a_537154_685355.n95 0.109
R853 a_537154_685355.n86 a_537154_685355.n85 0.104
R854 a_537154_685355.n103 a_537154_685355.n102 0.104
R855 a_537154_685355.n28 a_537154_685355.n27 0.095
R856 a_537154_685355.n135 a_537154_685355.n133 0.091
R857 a_537154_685355.n135 a_537154_685355.n134 0.091
R858 a_537154_685355.n182 a_537154_685355.n181 0.091
R859 a_537154_685355.n129 a_537154_685355.n127 0.091
R860 a_537154_685355.n129 a_537154_685355.n128 0.091
R861 a_537154_685355.n199 a_537154_685355.n198 0.091
R862 a_537154_685355.n189 a_537154_685355.n188 0.091
R863 a_537154_685355.n190 a_537154_685355.n189 0.091
R864 a_537154_685355.n123 a_537154_685355.n121 0.091
R865 a_537154_685355.n123 a_537154_685355.n122 0.091
R866 a_537154_685355.n165 a_537154_685355.n164 0.089
R867 a_537154_685355.n14 a_537154_685355.n13 0.089
R868 a_537154_685355.n159 a_537154_685355.n158 0.089
R869 a_537154_685355.n34 a_537154_685355.n33 0.089
R870 a_537154_685355.t6 a_537154_685355.n249 0.089
R871 a_537154_685355.n32 a_537154_685355.n31 0.088
R872 a_537154_685355.n242 a_537154_685355.n241 0.087
R873 a_537154_685355.n219 a_537154_685355.n218 0.087
R874 a_537154_685355.n5 a_537154_685355.n4 0.087
R875 a_537154_685355.n195 a_537154_685355.n194 0.087
R876 a_537154_685355.n24 a_537154_685355.n23 0.087
R877 a_537154_685355.n211 a_537154_685355.n210 0.085
R878 a_537154_685355.n249 a_537154_685355.n57 0.083
R879 a_537154_685355.n235 a_537154_685355.n234 0.075
R880 a_537154_685355.n232 a_537154_685355.n231 0.053
R881 a_537154_685355.n45 a_537154_685355.n44 0.028
R882 a_537154_685355.n118 a_537154_685355.n117 0.028
R883 a_537154_685355.n152 a_537154_685355.n151 0.028
R884 a_537154_685355.n186 a_537154_685355.n185 0.028
R885 a_537154_685355.n52 a_537154_685355.n51 0.028
R886 a_537154_685355.n38 a_537154_685355.n37 0.026
R887 a_537154_685355.n30 a_537154_685355.n29 0.023
R888 a_537154_685355.n230 a_537154_685355.n229 0.019
R889 a_537154_685355.n225 a_537154_685355.n224 0.015
R890 a_537154_685355.n30 a_537154_685355.n18 0.012
R891 a_537154_685355.n37 a_537154_685355.n36 0.012
R892 a_537154_685355.n227 a_537154_685355.n226 0.009
R893 a_537154_685355.n31 a_537154_685355.n30 0.007
R894 a_537154_685355.n37 a_537154_685355.n34 0.003
R895 a_537154_685355.n33 a_537154_685355.n32 0.003
R896 a_537154_685355.n146 a_537154_685355.n144 0.001
R897 a_537154_685355.n143 a_537154_685355.n141 0.001
R898 a_537154_685355.n245 a_537154_685355.n244 0.001
R899 a_537154_685355.n176 a_537154_685355.n174 0.001
R900 a_537154_685355.n8 a_537154_685355.n7 0.001
R901 a_537154_685355.n27 a_537154_685355.n26 0.001
R902 a_537154_685355.n32 a_537154_685355.n16 0.001
R903 a_537154_685355.n223 a_537154_685355.n222 0.001
R904 a_537154_685355.n60 a_537154_685355.n59 0.001
R905 a_537154_685355.n79 a_537154_685355.n78 0.001
R906 a_537154_685355.n94 a_537154_685355.n93 0.001
R907 a_537154_685355.n109 a_537154_685355.n108 0.001
R908 a_537154_685355.n68 a_537154_685355.n67 0.001
R909 a_537154_685355.n101 a_537154_685355.n100 0.001
R910 a_537154_685355.n67 a_537154_685355.n66 0.001
R911 a_537154_685355.n108 a_537154_685355.n107 0.001
R912 a_537154_685355.n96 a_537154_685355.n94 0.001
R913 a_537154_685355.n103 a_537154_685355.n101 0.001
R914 a_537154_685355.n84 a_537154_685355.n83 0.001
R915 a_537154_685355.n91 a_537154_685355.n71 0.001
R916 a_537154_685355.n91 a_537154_685355.n90 0.001
R917 a_537154_685355.n86 a_537154_685355.n84 0.001
R918 a_537154_685355.n104 a_537154_685355.n98 0.001
R919 a_537154_685355.n171 a_537154_685355.n169 0.001
R920 a_537154_685355.n87 a_537154_685355.n72 0.001
R921 a_537154_685355.n76 a_537154_685355.n73 0.001
R922 a_537154_685355.n81 a_537154_685355.n77 0.001
R923 a_537154_685355.n112 a_537154_685355.n63 0.001
R924 a_537154_685355.n240 a_537154_685355.n239 0.001
R925 a_537154_685355.n241 a_537154_685355.n240 0.001
R926 a_537154_685355.n239 a_537154_685355.n238 0.001
R927 a_537154_685355.n136 a_537154_685355.n135 0.001
R928 a_537154_685355.n136 a_537154_685355.n131 0.001
R929 a_537154_685355.n166 a_537154_685355.n163 0.001
R930 a_537154_685355.n166 a_537154_685355.n165 0.001
R931 a_537154_685355.n163 a_537154_685355.n162 0.001
R932 a_537154_685355.n220 a_537154_685355.n217 0.001
R933 a_537154_685355.n220 a_537154_685355.n219 0.001
R934 a_537154_685355.n217 a_537154_685355.n216 0.001
R935 a_537154_685355.n181 a_537154_685355.n180 0.001
R936 a_537154_685355.n201 a_537154_685355.n200 0.001
R937 a_537154_685355.n185 a_537154_685355.n184 0.001
R938 a_537154_685355.n185 a_537154_685355.n178 0.001
R939 a_537154_685355.n178 a_537154_685355.n177 0.001
R940 a_537154_685355.n151 a_537154_685355.n150 0.001
R941 a_537154_685355.n151 a_537154_685355.n148 0.001
R942 a_537154_685355.n148 a_537154_685355.n147 0.001
R943 a_537154_685355.n117 a_537154_685355.n116 0.001
R944 a_537154_685355.n117 a_537154_685355.n114 0.001
R945 a_537154_685355.n114 a_537154_685355.n113 0.001
R946 a_537154_685355.n45 a_537154_685355.n43 0.001
R947 a_537154_685355.n46 a_537154_685355.n45 0.001
R948 a_537154_685355.n46 a_537154_685355.n41 0.001
R949 a_537154_685355.n52 a_537154_685355.n50 0.001
R950 a_537154_685355.n53 a_537154_685355.n52 0.001
R951 a_537154_685355.n53 a_537154_685355.n40 0.001
R952 a_537154_685355.n12 a_537154_685355.n11 0.001
R953 a_537154_685355.n13 a_537154_685355.n12 0.001
R954 a_537154_685355.n11 a_537154_685355.n10 0.001
R955 a_537154_685355.n3 a_537154_685355.n2 0.001
R956 a_537154_685355.n4 a_537154_685355.n3 0.001
R957 a_537154_685355.n2 a_537154_685355.n1 0.001
R958 a_537154_685355.n130 a_537154_685355.n129 0.001
R959 a_537154_685355.n130 a_537154_685355.n125 0.001
R960 a_537154_685355.n160 a_537154_685355.n157 0.001
R961 a_537154_685355.n160 a_537154_685355.n159 0.001
R962 a_537154_685355.n157 a_537154_685355.n156 0.001
R963 a_537154_685355.n205 a_537154_685355.n199 0.001
R964 a_537154_685355.n205 a_537154_685355.n204 0.001
R965 a_537154_685355.n203 a_537154_685355.n202 0.001
R966 a_537154_685355.n196 a_537154_685355.n193 0.001
R967 a_537154_685355.n196 a_537154_685355.n195 0.001
R968 a_537154_685355.n193 a_537154_685355.n192 0.001
R969 a_537154_685355.n124 a_537154_685355.n123 0.001
R970 a_537154_685355.n124 a_537154_685355.n119 0.001
R971 a_537154_685355.n22 a_537154_685355.n21 0.001
R972 a_537154_685355.n23 a_537154_685355.n22 0.001
R973 a_537154_685355.n21 a_537154_685355.n20 0.001
R974 a_40125_693523.n74 a_40125_693523.t57 271.872
R975 a_40125_693523.n47 a_40125_693523.t71 271.872
R976 a_40125_693523.n64 a_40125_693523.t65 271.866
R977 a_40125_693523.n63 a_40125_693523.t67 271.866
R978 a_40125_693523.n62 a_40125_693523.t34 271.866
R979 a_40125_693523.n61 a_40125_693523.t52 271.866
R980 a_40125_693523.n60 a_40125_693523.t40 271.866
R981 a_40125_693523.n59 a_40125_693523.t50 271.866
R982 a_40125_693523.n58 a_40125_693523.t54 271.866
R983 a_40125_693523.n46 a_40125_693523.t33 271.866
R984 a_40125_693523.n45 a_40125_693523.t41 271.866
R985 a_40125_693523.n44 a_40125_693523.t45 271.866
R986 a_40125_693523.n43 a_40125_693523.t49 271.866
R987 a_40125_693523.n42 a_40125_693523.t60 271.866
R988 a_40125_693523.n41 a_40125_693523.t63 271.866
R989 a_40125_693523.n40 a_40125_693523.t68 271.866
R990 a_40125_693523.n39 a_40125_693523.t32 271.866
R991 a_40125_693523.n38 a_40125_693523.t55 271.866
R992 a_40125_693523.n37 a_40125_693523.t59 271.866
R993 a_40125_693523.n36 a_40125_693523.t47 271.866
R994 a_40125_693523.n35 a_40125_693523.t56 271.866
R995 a_40125_693523.n34 a_40125_693523.t61 271.866
R996 a_40125_693523.n33 a_40125_693523.t37 271.866
R997 a_40125_693523.n32 a_40125_693523.t42 271.866
R998 a_40125_693523.n65 a_40125_693523.t51 271.866
R999 a_40125_693523.n66 a_40125_693523.t39 271.866
R1000 a_40125_693523.n67 a_40125_693523.t44 271.866
R1001 a_40125_693523.n68 a_40125_693523.t66 271.866
R1002 a_40125_693523.n69 a_40125_693523.t69 271.866
R1003 a_40125_693523.n70 a_40125_693523.t36 271.866
R1004 a_40125_693523.n71 a_40125_693523.t38 271.866
R1005 a_40125_693523.n72 a_40125_693523.t70 271.866
R1006 a_40125_693523.n73 a_40125_693523.t53 271.866
R1007 a_40125_693523.n31 a_40125_693523.t62 271.866
R1008 a_40125_693523.n30 a_40125_693523.t35 271.866
R1009 a_40125_693523.n29 a_40125_693523.t43 271.866
R1010 a_40125_693523.n28 a_40125_693523.t48 271.866
R1011 a_40125_693523.n27 a_40125_693523.t58 271.866
R1012 a_40125_693523.n26 a_40125_693523.t46 271.866
R1013 a_40125_693523.n25 a_40125_693523.t64 271.866
R1014 a_40125_693523.n97 a_40125_693523.t3 6.245
R1015 a_40125_693523.n77 a_40125_693523.t31 5.713
R1016 a_40125_693523.n77 a_40125_693523.t2 5.713
R1017 a_40125_693523.n79 a_40125_693523.t0 5.713
R1018 a_40125_693523.n79 a_40125_693523.t24 5.713
R1019 a_40125_693523.n81 a_40125_693523.t27 5.713
R1020 a_40125_693523.n81 a_40125_693523.t9 5.713
R1021 a_40125_693523.n83 a_40125_693523.t8 5.713
R1022 a_40125_693523.n83 a_40125_693523.t26 5.713
R1023 a_40125_693523.n85 a_40125_693523.t15 5.713
R1024 a_40125_693523.n85 a_40125_693523.t20 5.713
R1025 a_40125_693523.n87 a_40125_693523.t12 5.713
R1026 a_40125_693523.n87 a_40125_693523.t29 5.713
R1027 a_40125_693523.n89 a_40125_693523.t14 5.713
R1028 a_40125_693523.n89 a_40125_693523.t19 5.713
R1029 a_40125_693523.n91 a_40125_693523.t1 5.713
R1030 a_40125_693523.n91 a_40125_693523.t25 5.713
R1031 a_40125_693523.n93 a_40125_693523.t13 5.713
R1032 a_40125_693523.n93 a_40125_693523.t16 5.713
R1033 a_40125_693523.n95 a_40125_693523.t11 5.713
R1034 a_40125_693523.n95 a_40125_693523.t28 5.713
R1035 a_40125_693523.n98 a_40125_693523.t22 3.797
R1036 a_40125_693523.n99 a_40125_693523.t4 3.48
R1037 a_40125_693523.n99 a_40125_693523.t21 3.48
R1038 a_40125_693523.n101 a_40125_693523.t23 3.48
R1039 a_40125_693523.n101 a_40125_693523.t18 3.48
R1040 a_40125_693523.n103 a_40125_693523.t7 3.48
R1041 a_40125_693523.n103 a_40125_693523.t10 3.48
R1042 a_40125_693523.n48 a_40125_693523.t17 2.639
R1043 a_40125_693523.n115 a_40125_693523.t30 2.591
R1044 a_40125_693523.n48 a_40125_693523.t6 2.576
R1045 a_40125_693523.n105 a_40125_693523.n104 2.006
R1046 a_40125_693523.n114 a_40125_693523.n113 1.109
R1047 a_40125_693523.n58 a_40125_693523.n57 1.094
R1048 a_40125_693523.n114 a_40125_693523.n31 1.062
R1049 a_40125_693523.n57 a_40125_693523.n56 1.047
R1050 a_40125_693523.n106 a_40125_693523.n105 1.008
R1051 a_40125_693523.n76 a_40125_693523.n75 1.008
R1052 a_40125_693523.n80 a_40125_693523.n79 0.532
R1053 a_40125_693523.n82 a_40125_693523.n81 0.532
R1054 a_40125_693523.n84 a_40125_693523.n83 0.532
R1055 a_40125_693523.n86 a_40125_693523.n85 0.532
R1056 a_40125_693523.n88 a_40125_693523.n87 0.532
R1057 a_40125_693523.n90 a_40125_693523.n89 0.532
R1058 a_40125_693523.n92 a_40125_693523.n91 0.532
R1059 a_40125_693523.n94 a_40125_693523.n93 0.532
R1060 a_40125_693523.n96 a_40125_693523.n95 0.532
R1061 a_40125_693523.n78 a_40125_693523.n77 0.532
R1062 a_40125_693523.n113 a_40125_693523.n112 0.395
R1063 a_40125_693523.n112 a_40125_693523.n111 0.395
R1064 a_40125_693523.n111 a_40125_693523.n110 0.395
R1065 a_40125_693523.n110 a_40125_693523.n109 0.395
R1066 a_40125_693523.n109 a_40125_693523.n108 0.395
R1067 a_40125_693523.n108 a_40125_693523.n107 0.395
R1068 a_40125_693523.n46 a_40125_693523.n45 0.395
R1069 a_40125_693523.n45 a_40125_693523.n44 0.395
R1070 a_40125_693523.n44 a_40125_693523.n43 0.395
R1071 a_40125_693523.n43 a_40125_693523.n42 0.395
R1072 a_40125_693523.n42 a_40125_693523.n41 0.395
R1073 a_40125_693523.n41 a_40125_693523.n40 0.395
R1074 a_40125_693523.n40 a_40125_693523.n39 0.395
R1075 a_40125_693523.n39 a_40125_693523.n38 0.395
R1076 a_40125_693523.n38 a_40125_693523.n37 0.395
R1077 a_40125_693523.n37 a_40125_693523.n36 0.395
R1078 a_40125_693523.n36 a_40125_693523.n35 0.395
R1079 a_40125_693523.n35 a_40125_693523.n34 0.395
R1080 a_40125_693523.n34 a_40125_693523.n33 0.395
R1081 a_40125_693523.n33 a_40125_693523.n32 0.395
R1082 a_40125_693523.n66 a_40125_693523.n65 0.395
R1083 a_40125_693523.n67 a_40125_693523.n66 0.395
R1084 a_40125_693523.n68 a_40125_693523.n67 0.395
R1085 a_40125_693523.n69 a_40125_693523.n68 0.395
R1086 a_40125_693523.n70 a_40125_693523.n69 0.395
R1087 a_40125_693523.n71 a_40125_693523.n70 0.395
R1088 a_40125_693523.n72 a_40125_693523.n71 0.395
R1089 a_40125_693523.n73 a_40125_693523.n72 0.395
R1090 a_40125_693523.n64 a_40125_693523.n63 0.395
R1091 a_40125_693523.n63 a_40125_693523.n62 0.395
R1092 a_40125_693523.n62 a_40125_693523.n61 0.395
R1093 a_40125_693523.n61 a_40125_693523.n60 0.395
R1094 a_40125_693523.n60 a_40125_693523.n59 0.395
R1095 a_40125_693523.n59 a_40125_693523.n58 0.395
R1096 a_40125_693523.n31 a_40125_693523.n30 0.395
R1097 a_40125_693523.n30 a_40125_693523.n29 0.395
R1098 a_40125_693523.n29 a_40125_693523.n28 0.395
R1099 a_40125_693523.n28 a_40125_693523.n27 0.395
R1100 a_40125_693523.n27 a_40125_693523.n26 0.395
R1101 a_40125_693523.n26 a_40125_693523.n25 0.395
R1102 a_40125_693523.n25 a_40125_693523.n24 0.395
R1103 a_40125_693523.n24 a_40125_693523.n23 0.395
R1104 a_40125_693523.n23 a_40125_693523.n22 0.395
R1105 a_40125_693523.n22 a_40125_693523.n21 0.395
R1106 a_40125_693523.n21 a_40125_693523.n20 0.395
R1107 a_40125_693523.n20 a_40125_693523.n19 0.395
R1108 a_40125_693523.n19 a_40125_693523.n18 0.395
R1109 a_40125_693523.n18 a_40125_693523.n17 0.395
R1110 a_40125_693523.n17 a_40125_693523.n16 0.395
R1111 a_40125_693523.n16 a_40125_693523.n15 0.395
R1112 a_40125_693523.n15 a_40125_693523.n14 0.395
R1113 a_40125_693523.n14 a_40125_693523.n13 0.395
R1114 a_40125_693523.n13 a_40125_693523.n12 0.395
R1115 a_40125_693523.n12 a_40125_693523.n11 0.395
R1116 a_40125_693523.n11 a_40125_693523.n10 0.395
R1117 a_40125_693523.n10 a_40125_693523.n9 0.395
R1118 a_40125_693523.n9 a_40125_693523.n8 0.395
R1119 a_40125_693523.n8 a_40125_693523.n7 0.395
R1120 a_40125_693523.n7 a_40125_693523.n6 0.395
R1121 a_40125_693523.n6 a_40125_693523.n5 0.395
R1122 a_40125_693523.n5 a_40125_693523.n4 0.395
R1123 a_40125_693523.n4 a_40125_693523.n3 0.395
R1124 a_40125_693523.n3 a_40125_693523.n2 0.395
R1125 a_40125_693523.n2 a_40125_693523.n1 0.395
R1126 a_40125_693523.n1 a_40125_693523.n0 0.395
R1127 a_40125_693523.n50 a_40125_693523.n49 0.395
R1128 a_40125_693523.n51 a_40125_693523.n50 0.395
R1129 a_40125_693523.n52 a_40125_693523.n51 0.395
R1130 a_40125_693523.n53 a_40125_693523.n52 0.395
R1131 a_40125_693523.n54 a_40125_693523.n53 0.395
R1132 a_40125_693523.n55 a_40125_693523.n54 0.395
R1133 a_40125_693523.n56 a_40125_693523.n55 0.395
R1134 a_40125_693523.n74 a_40125_693523.n73 0.37
R1135 a_40125_693523.n47 a_40125_693523.n46 0.351
R1136 a_40125_693523.n57 a_40125_693523.n48 0.349
R1137 a_40125_693523.n115 a_40125_693523.n114 0.349
R1138 a_40125_693523.t5 a_40125_693523.n115 0.344
R1139 a_40125_693523.n102 a_40125_693523.n101 0.317
R1140 a_40125_693523.n100 a_40125_693523.n99 0.317
R1141 a_40125_693523.n104 a_40125_693523.n103 0.317
R1142 a_40125_693523.n107 a_40125_693523.n106 0.166
R1143 a_40125_693523.n75 a_40125_693523.n64 0.13
R1144 a_40125_693523.n78 a_40125_693523.n76 0.083
R1145 a_40125_693523.n75 a_40125_693523.n74 0.071
R1146 a_40125_693523.n105 a_40125_693523.n97 0.057
R1147 a_40125_693523.n106 a_40125_693523.n47 0.054
R1148 a_40125_693523.n96 a_40125_693523.n94 0.05
R1149 a_40125_693523.n94 a_40125_693523.n92 0.05
R1150 a_40125_693523.n90 a_40125_693523.n88 0.05
R1151 a_40125_693523.n86 a_40125_693523.n84 0.05
R1152 a_40125_693523.n84 a_40125_693523.n82 0.05
R1153 a_40125_693523.n80 a_40125_693523.n78 0.05
R1154 a_40125_693523.n97 a_40125_693523.n96 0.048
R1155 a_40125_693523.n92 a_40125_693523.n90 0.048
R1156 a_40125_693523.n88 a_40125_693523.n86 0.048
R1157 a_40125_693523.n82 a_40125_693523.n80 0.048
R1158 a_40125_693523.n104 a_40125_693523.n102 0.039
R1159 a_40125_693523.n100 a_40125_693523.n98 0.039
R1160 a_40125_693523.n102 a_40125_693523.n100 0.038
R1161 vccd2.n177 vccd2.n174 185
R1162 vccd2.n49 vccd2.n34 185
R1163 vccd2.n33 vccd2.n32 127.623
R1164 vccd2.n160 vccd2.n159 126.117
R1165 vccd2.t26 vccd2.t14 83.367
R1166 vccd2.t14 vccd2.t16 83.367
R1167 vccd2.t32 vccd2.t37 83.367
R1168 vccd2.t24 vccd2.t32 83.367
R1169 vccd2.n14 vccd2.t26 78.52
R1170 vccd2.n224 vccd2.t24 78.52
R1171 vccd2.t37 vccd2.n210 41.683
R1172 vccd2.t77 vccd2.n163 38.604
R1173 vccd2.t93 vccd2.n38 38.604
R1174 vccd2.t131 vccd2.t77 31.6
R1175 vccd2.t109 vccd2.t131 31.6
R1176 vccd2.t111 vccd2.t109 31.6
R1177 vccd2.t85 vccd2.t111 31.6
R1178 vccd2.t73 vccd2.t115 31.6
R1179 vccd2.t59 vccd2.t73 31.6
R1180 vccd2.t135 vccd2.t59 31.6
R1181 vccd2.t95 vccd2.t87 31.6
R1182 vccd2.t87 vccd2.t71 31.6
R1183 vccd2.t71 vccd2.t67 31.6
R1184 vccd2.t133 vccd2.t97 31.6
R1185 vccd2.t97 vccd2.t125 31.6
R1186 vccd2.t125 vccd2.t101 31.6
R1187 vccd2.t101 vccd2.t93 31.6
R1188 vccd2.t67 vccd2.n41 24.2
R1189 vccd2.t115 vccd2.n168 24
R1190 vccd2.t61 vccd2.n46 23
R1191 vccd2.t123 vccd2.n173 22.6
R1192 vccd2.t8 vccd2.t123 16
R1193 vccd2.t47 vccd2.t117 16
R1194 vccd2.t30 vccd2.t81 16
R1195 vccd2.t55 vccd2.t75 16
R1196 vccd2.t4 vccd2.t65 16
R1197 vccd2.t137 vccd2.t22 16
R1198 vccd2.t91 vccd2.t52 16
R1199 vccd2.t10 vccd2.t113 16
R1200 vccd2.t79 vccd2.t0 16
R1201 vccd2.t127 vccd2.t39 16
R1202 vccd2.t41 vccd2.t121 16
R1203 vccd2.t150 vccd2.t99 16
R1204 vccd2.t119 vccd2.t43 16
R1205 vccd2.t69 vccd2.t2 16
R1206 vccd2.t63 vccd2.t12 16
R1207 vccd2.t107 vccd2.t6 16
R1208 vccd2.t117 vccd2.t8 15.6
R1209 vccd2.t81 vccd2.t45 15.6
R1210 vccd2.t75 vccd2.t30 15.6
R1211 vccd2.t65 vccd2.t55 15.6
R1212 vccd2.t22 vccd2.t91 15.6
R1213 vccd2.t52 vccd2.t83 15.6
R1214 vccd2.t113 vccd2.t20 15.6
R1215 vccd2.t89 vccd2.t10 15.6
R1216 vccd2.t142 vccd2.t79 15.6
R1217 vccd2.t0 vccd2.t127 15.6
R1218 vccd2.t99 vccd2.t41 15.6
R1219 vccd2.t105 vccd2.t150 15.6
R1220 vccd2.t34 vccd2.t119 15.6
R1221 vccd2.t43 vccd2.t69 15.6
R1222 vccd2.t2 vccd2.t63 15.6
R1223 vccd2.t146 vccd2.t107 15.6
R1224 vccd2.t6 vccd2.t61 15.6
R1225 vccd2.n97 vccd2.t89 15.2
R1226 vccd2.n90 vccd2.n87 14.117
R1227 vccd2.n49 vccd2.t146 13.4
R1228 vccd2.n177 vccd2.t47 12.6
R1229 vccd2.n55 vccd2.t34 11.8
R1230 vccd2.n180 vccd2.t103 11.6
R1231 vccd2.n52 vccd2.t129 11.2
R1232 vccd2.n182 vccd2.t4 10.2
R1233 vccd2.n173 vccd2.t135 9
R1234 vccd2.n46 vccd2.t95 8.6
R1235 vccd2.n168 vccd2.t85 7.6
R1236 vccd2.n41 vccd2.t133 7.4
R1237 vccd2.n197 vccd2.t25 6.413
R1238 vccd2.n23 vccd2.t155 6.413
R1239 vccd2.n77 vccd2.t7 6.3
R1240 vccd2.n58 vccd2.t19 6.273
R1241 vccd2.n101 vccd2.t94 6.215
R1242 vccd2.n121 vccd2.t78 6.214
R1243 vccd2.n228 vccd2.t28 5.713
R1244 vccd2.n193 vccd2.t38 5.713
R1245 vccd2.n193 vccd2.t158 5.713
R1246 vccd2.n191 vccd2.t36 5.713
R1247 vccd2.n191 vccd2.t139 5.713
R1248 vccd2.n20 vccd2.t27 5.713
R1249 vccd2.n195 vccd2.t144 5.713
R1250 vccd2.n195 vccd2.t33 5.713
R1251 vccd2.n21 vccd2.t15 5.713
R1252 vccd2.n21 vccd2.t17 5.713
R1253 vccd2.n29 vccd2.t149 5.713
R1254 vccd2.n29 vccd2.t18 5.713
R1255 vccd2.n27 vccd2.t23 5.713
R1256 vccd2.n27 vccd2.t152 5.713
R1257 vccd2.n154 vccd2.t21 5.713
R1258 vccd2.n154 vccd2.t11 5.713
R1259 vccd2.n151 vccd2.t143 5.713
R1260 vccd2.n151 vccd2.t1 5.713
R1261 vccd2.n149 vccd2.t40 5.713
R1262 vccd2.n149 vccd2.t145 5.713
R1263 vccd2.n147 vccd2.t151 5.713
R1264 vccd2.n147 vccd2.t35 5.713
R1265 vccd2.n59 vccd2.t50 5.713
R1266 vccd2.n59 vccd2.t148 5.713
R1267 vccd2.n57 vccd2.t13 5.713
R1268 vccd2.n57 vccd2.t147 5.713
R1269 vccd2.n25 vccd2.t29 5.713
R1270 vccd2.n25 vccd2.t160 5.713
R1271 vccd2.n26 vccd2.t46 5.713
R1272 vccd2.n26 vccd2.t31 5.713
R1273 vccd2.n68 vccd2.t56 5.713
R1274 vccd2.n68 vccd2.t5 5.713
R1275 vccd2.n70 vccd2.t141 5.713
R1276 vccd2.n70 vccd2.t53 5.713
R1277 vccd2.n72 vccd2.t57 5.713
R1278 vccd2.n72 vccd2.t49 5.713
R1279 vccd2.n65 vccd2.t157 5.713
R1280 vccd2.n65 vccd2.t54 5.713
R1281 vccd2.n63 vccd2.t58 5.713
R1282 vccd2.n63 vccd2.t42 5.713
R1283 vccd2.n78 vccd2.t153 5.713
R1284 vccd2.n78 vccd2.t154 5.713
R1285 vccd2.n80 vccd2.t44 5.713
R1286 vccd2.n80 vccd2.t3 5.713
R1287 vccd2.n76 vccd2.t140 5.713
R1288 vccd2.n76 vccd2.t159 5.713
R1289 vccd2.n85 vccd2.t9 5.713
R1290 vccd2.n85 vccd2.t48 5.713
R1291 vccd2.n83 vccd2.t156 5.713
R1292 vccd2.n83 vccd2.t51 5.713
R1293 vccd2.n123 vccd2.t116 5.713
R1294 vccd2.n123 vccd2.t74 5.713
R1295 vccd2.n125 vccd2.t60 5.713
R1296 vccd2.n125 vccd2.t136 5.713
R1297 vccd2.n127 vccd2.t124 5.713
R1298 vccd2.n127 vccd2.t118 5.713
R1299 vccd2.n129 vccd2.t104 5.713
R1300 vccd2.n129 vccd2.t82 5.713
R1301 vccd2.n131 vccd2.t76 5.713
R1302 vccd2.n131 vccd2.t66 5.713
R1303 vccd2.n137 vccd2.t138 5.713
R1304 vccd2.n137 vccd2.t92 5.713
R1305 vccd2.n135 vccd2.t84 5.713
R1306 vccd2.n135 vccd2.t114 5.713
R1307 vccd2.n133 vccd2.t90 5.713
R1308 vccd2.n133 vccd2.t80 5.713
R1309 vccd2.n103 vccd2.t128 5.713
R1310 vccd2.n103 vccd2.t122 5.713
R1311 vccd2.n105 vccd2.t100 5.713
R1312 vccd2.n105 vccd2.t106 5.713
R1313 vccd2.n115 vccd2.t120 5.713
R1314 vccd2.n115 vccd2.t70 5.713
R1315 vccd2.n113 vccd2.t64 5.713
R1316 vccd2.n113 vccd2.t130 5.713
R1317 vccd2.n111 vccd2.t108 5.713
R1318 vccd2.n111 vccd2.t62 5.713
R1319 vccd2.n109 vccd2.t96 5.713
R1320 vccd2.n109 vccd2.t88 5.713
R1321 vccd2.n107 vccd2.t72 5.713
R1322 vccd2.n107 vccd2.t68 5.713
R1323 vccd2.n98 vccd2.t134 5.713
R1324 vccd2.n98 vccd2.t98 5.713
R1325 vccd2.n100 vccd2.t126 5.713
R1326 vccd2.n100 vccd2.t102 5.713
R1327 vccd2.n120 vccd2.t132 5.713
R1328 vccd2.n120 vccd2.t110 5.713
R1329 vccd2.n118 vccd2.t112 5.713
R1330 vccd2.n118 vccd2.t86 5.713
R1331 vccd2.n182 vccd2.t137 5.4
R1332 vccd2.n55 vccd2.n54 4.65
R1333 vccd2.n182 vccd2.n181 4.65
R1334 vccd2.n183 vccd2.n161 4.593
R1335 vccd2.n55 vccd2.n53 4.591
R1336 vccd2.t45 vccd2.n180 4.4
R1337 vccd2.t12 vccd2.n52 4.4
R1338 vccd2.n55 vccd2.t105 4.2
R1339 vccd2.n56 vccd2.n33 3.798
R1340 vccd2.n184 vccd2.n160 3.797
R1341 vccd2.t103 vccd2.n177 3
R1342 vccd2.t129 vccd2.n49 2.6
R1343 vccd2.n89 vccd2.n88 1.505
R1344 vccd2.n188 vccd2.n187 1.282
R1345 vccd2.n189 vccd2.n188 1.274
R1346 vccd2.n196 vccd2.n195 0.7
R1347 vccd2.n22 vccd2.n21 0.7
R1348 vccd2.t142 vccd2.n97 0.6
R1349 vccd2.n194 vccd2.n193 0.593
R1350 vccd2.n192 vccd2.n191 0.593
R1351 vccd2.n86 vccd2.n85 0.565
R1352 vccd2.n73 vccd2.n72 0.542
R1353 vccd2.n64 vccd2.n63 0.541
R1354 vccd2.n71 vccd2.n70 0.541
R1355 vccd2.n77 vccd2.n76 0.541
R1356 vccd2.n81 vccd2.n80 0.54
R1357 vccd2.n84 vccd2.n83 0.539
R1358 vccd2.n66 vccd2.n65 0.537
R1359 vccd2.n79 vccd2.n78 0.537
R1360 vccd2.n69 vccd2.n68 0.537
R1361 vccd2.n155 vccd2.n154 0.515
R1362 vccd2.n150 vccd2.n149 0.514
R1363 vccd2.n58 vccd2.n57 0.514
R1364 vccd2.n187 vccd2.n25 0.514
R1365 vccd2.n60 vccd2.n59 0.513
R1366 vccd2.n31 vccd2.n26 0.513
R1367 vccd2.n28 vccd2.n27 0.511
R1368 vccd2.n152 vccd2.n151 0.511
R1369 vccd2.n148 vccd2.n147 0.511
R1370 vccd2.n30 vccd2.n29 0.511
R1371 vccd2.n188 vccd2.n24 0.464
R1372 vccd2.n114 vccd2.n113 0.461
R1373 vccd2.n104 vccd2.n103 0.461
R1374 vccd2.n136 vccd2.n135 0.461
R1375 vccd2.n130 vccd2.n129 0.461
R1376 vccd2.n126 vccd2.n125 0.461
R1377 vccd2.n121 vccd2.n120 0.461
R1378 vccd2.n101 vccd2.n100 0.459
R1379 vccd2.n128 vccd2.n127 0.457
R1380 vccd2.n132 vccd2.n131 0.457
R1381 vccd2.n138 vccd2.n137 0.457
R1382 vccd2.n134 vccd2.n133 0.457
R1383 vccd2.n106 vccd2.n105 0.457
R1384 vccd2.n116 vccd2.n115 0.457
R1385 vccd2.n112 vccd2.n111 0.457
R1386 vccd2.n110 vccd2.n109 0.457
R1387 vccd2.n108 vccd2.n107 0.457
R1388 vccd2.n99 vccd2.n98 0.457
R1389 vccd2.n124 vccd2.n123 0.457
R1390 vccd2.n119 vccd2.n118 0.457
R1391 vccd2.n190 vccd2.n20 0.336
R1392 vccd2.n229 vccd2.n228 0.335
R1393 vccd2.n190 vccd2.n189 0.323
R1394 vccd2.n230 vccd2.n198 0.321
R1395 vccd2.n23 vccd2.n22 0.203
R1396 vccd2.n197 vccd2.n196 0.199
R1397 vccd2.n117 vccd2.n102 0.168
R1398 vccd2.n139 vccd2.n122 0.166
R1399 vccd2.n144 vccd2.t142 0.084
R1400 vccd2.n198 vccd2.n197 0.082
R1401 vccd2.n186 vccd2.n185 0.069
R1402 vccd2.n145 vccd2.n86 0.058
R1403 vccd2.n185 vccd2.n61 0.054
R1404 vccd2.n31 vccd2.n30 0.05
R1405 vccd2.n30 vccd2.n28 0.05
R1406 vccd2.n150 vccd2.n148 0.05
R1407 vccd2.n73 vccd2.n71 0.05
R1408 vccd2.n81 vccd2.n79 0.05
R1409 vccd2.n71 vccd2.n69 0.048
R1410 vccd2.n66 vccd2.n64 0.048
R1411 vccd2.n152 vccd2.n150 0.048
R1412 vccd2.n145 vccd2.n82 0.047
R1413 vccd2.n128 vccd2.n126 0.045
R1414 vccd2.n132 vccd2.n130 0.045
R1415 vccd2.n136 vccd2.n134 0.045
R1416 vccd2.n106 vccd2.n104 0.045
R1417 vccd2.n114 vccd2.n112 0.045
R1418 vccd2.n112 vccd2.n110 0.045
R1419 vccd2.n126 vccd2.n124 0.044
R1420 vccd2.n130 vccd2.n128 0.044
R1421 vccd2.n138 vccd2.n136 0.044
R1422 vccd2.n116 vccd2.n114 0.044
R1423 vccd2.n110 vccd2.n108 0.044
R1424 vccd2.n185 vccd2.n184 0.031
R1425 vccd2.n185 vccd2.n56 0.029
R1426 vccd2.n82 vccd2.n77 0.027
R1427 vccd2.n185 vccd2.n145 0.027
R1428 vccd2.n61 vccd2.n60 0.026
R1429 vccd2.n82 vccd2.n81 0.026
R1430 vccd2.n67 vccd2.n66 0.025
R1431 vccd2.n153 vccd2.n152 0.025
R1432 vccd2.n187 vccd2.n186 0.025
R1433 vccd2.n86 vccd2.n84 0.025
R1434 vccd2.n186 vccd2.n31 0.025
R1435 vccd2.n192 vccd2.n190 0.024
R1436 vccd2.n102 vccd2.n101 0.023
R1437 vccd2.n61 vccd2.n58 0.023
R1438 vccd2.n144 vccd2.n143 0.023
R1439 vccd2.n102 vccd2.n99 0.023
R1440 vccd2.n189 vccd2.n23 0.022
R1441 vccd2.n122 vccd2.n121 0.022
R1442 vccd2.n122 vccd2.n119 0.022
R1443 vccd2.n139 vccd2.n132 0.022
R1444 vccd2.n139 vccd2.n138 0.022
R1445 vccd2.n117 vccd2.n106 0.022
R1446 vccd2.n117 vccd2.n116 0.022
R1447 vccd2.n194 vccd2.n192 0.021
R1448 vccd2.n157 vccd2.n156 0.02
R1449 vccd2.n219 vccd2.n218 0.02
R1450 vccd2.n224 vccd2.n219 0.02
R1451 vccd2.n11 vccd2.n10 0.02
R1452 vccd2.n14 vccd2.n11 0.02
R1453 vccd2.n17 vccd2.n16 0.019
R1454 vccd2.n4 vccd2.n3 0.019
R1455 vccd2.n75 vccd2.n74 0.019
R1456 vccd2.n3 vccd2.n2 0.019
R1457 vccd2.n16 vccd2.n15 0.019
R1458 vccd2.n223 vccd2.n222 0.019
R1459 vccd2.n224 vccd2.n223 0.019
R1460 vccd2.n212 vccd2.n211 0.019
R1461 vccd2.n224 vccd2.n212 0.019
R1462 vccd2.n13 vccd2.n12 0.018
R1463 vccd2.n14 vccd2.n13 0.018
R1464 vccd2.n221 vccd2.n220 0.018
R1465 vccd2.n224 vccd2.n221 0.018
R1466 vccd2.n158 vccd2.n146 0.017
R1467 vccd2.n145 vccd2.n62 0.017
R1468 vccd2.n48 vccd2.n47 0.013
R1469 vccd2.n49 vccd2.n48 0.013
R1470 vccd2.n176 vccd2.n175 0.013
R1471 vccd2.n177 vccd2.n176 0.013
R1472 vccd2 vccd2.n194 0.012
R1473 vccd2.n52 vccd2.n51 0.01
R1474 vccd2.n180 vccd2.n179 0.01
R1475 vccd2.n143 vccd2.n117 0.01
R1476 vccd2.n143 vccd2.n142 0.01
R1477 vccd2.n145 vccd2.n144 0.01
R1478 vccd2.n51 vccd2.n50 0.01
R1479 vccd2.n179 vccd2.n178 0.01
R1480 vccd2.n96 vccd2.n95 0.009
R1481 vccd2.n97 vccd2.n96 0.009
R1482 vccd2.n184 vccd2.n183 0.008
R1483 vccd2.n4 vccd2.n1 0.007
R1484 vccd2.n217 vccd2.n214 0.007
R1485 vccd2.n9 vccd2.n6 0.007
R1486 vccd2.n225 vccd2.n201 0.007
R1487 vccd2.n201 vccd2.n200 0.007
R1488 vccd2.n1 vccd2.n0 0.007
R1489 vccd2.n214 vccd2.n213 0.007
R1490 vccd2.n6 vccd2.n5 0.007
R1491 vccd2.n143 vccd2.n139 0.007
R1492 vccd2.n56 vccd2.n55 0.007
R1493 vccd2 vccd2.n231 0.006
R1494 vccd2.n156 vccd2.n155 0.006
R1495 vccd2.n74 vccd2.n73 0.005
R1496 vccd2.n165 vccd2.n164 0.005
R1497 vccd2.n36 vccd2.n35 0.005
R1498 vccd2.n24 vccd2 0.005
R1499 vccd2.n41 vccd2.n36 0.005
R1500 vccd2.n168 vccd2.n165 0.005
R1501 vccd2.n167 vccd2.n166 0.005
R1502 vccd2.n168 vccd2.n167 0.005
R1503 vccd2.n40 vccd2.n39 0.005
R1504 vccd2.n41 vccd2.n40 0.005
R1505 vccd2.n231 vccd2.n230 0.005
R1506 vccd2.n185 vccd2.n158 0.004
R1507 vccd2.n230 vccd2.n229 0.004
R1508 vccd2.n45 vccd2.n44 0.004
R1509 vccd2.n46 vccd2.n45 0.004
R1510 vccd2.n172 vccd2.n171 0.004
R1511 vccd2.n173 vccd2.n172 0.004
R1512 vccd2.n43 vccd2.n42 0.004
R1513 vccd2.n46 vccd2.n43 0.004
R1514 vccd2.n170 vccd2.n169 0.004
R1515 vccd2.n173 vccd2.n170 0.004
R1516 vccd2.n38 vccd2.n37 0.004
R1517 vccd2.n163 vccd2.n162 0.004
R1518 vccd2.n209 vccd2.n208 0.003
R1519 vccd2.n210 vccd2.n209 0.003
R1520 vccd2.n207 vccd2.n206 0.003
R1521 vccd2.n210 vccd2.n207 0.003
R1522 vccd2.n205 vccd2.n204 0.003
R1523 vccd2.n210 vccd2.n205 0.003
R1524 vccd2.n203 vccd2.n202 0.003
R1525 vccd2.n210 vccd2.n203 0.003
R1526 vccd2.n18 vccd2.n17 0.002
R1527 vccd2.n217 vccd2.n216 0.002
R1528 vccd2.n9 vccd2.n8 0.002
R1529 vccd2.n226 vccd2.n225 0.002
R1530 vccd2.n227 vccd2.n226 0.002
R1531 vccd2.n19 vccd2.n18 0.002
R1532 vccd2.n216 vccd2.n215 0.002
R1533 vccd2.n8 vccd2.n7 0.002
R1534 vccd2.n94 vccd2.n93 0.002
R1535 vccd2.t142 vccd2.n94 0.002
R1536 vccd2.n90 vccd2.n89 0.002
R1537 vccd2.t142 vccd2.n90 0.002
R1538 vccd2.n20 vccd2.n19 0.002
R1539 vccd2.n228 vccd2.n227 0.002
R1540 vccd2.n145 vccd2.n75 0.001
R1541 vccd2.n183 vccd2.n182 0.001
R1542 vccd2.n92 vccd2.n91 0.001
R1543 vccd2.t142 vccd2.n92 0.001
R1544 vccd2.n24 vccd2 0.001
R1545 vccd2.n142 vccd2.n141 0.001
R1546 vccd2.n142 vccd2.n140 0.001
R1547 vccd2.n229 vccd2.n199 0.001
R1548 vccd2.n75 vccd2.n67 0.001
R1549 vccd2.n225 vccd2.n224 0.001
R1550 vccd2.n224 vccd2.n217 0.001
R1551 vccd2.n14 vccd2.n9 0.001
R1552 vccd2.n14 vccd2.n4 0.001
R1553 vccd2.n17 vccd2.n14 0.001
R1554 vccd2.n157 vccd2.n153 0.001
R1555 vccd2.n158 vccd2.n157 0.001
R1556 io_analog[10].n5 io_analog[10].n4 6.526
R1557 io_analog[10].n56 io_analog[10].n55 6.355
R1558 io_analog[10].n2 io_analog[10].t19 5.713
R1559 io_analog[10].n2 io_analog[10].t46 5.713
R1560 io_analog[10].n49 io_analog[10].t29 5.713
R1561 io_analog[10].n49 io_analog[10].t41 5.713
R1562 io_analog[10].n47 io_analog[10].t14 5.713
R1563 io_analog[10].n47 io_analog[10].t47 5.713
R1564 io_analog[10].n45 io_analog[10].t24 5.713
R1565 io_analog[10].n45 io_analog[10].t16 5.713
R1566 io_analog[10].n43 io_analog[10].t11 5.713
R1567 io_analog[10].n43 io_analog[10].t28 5.713
R1568 io_analog[10].n41 io_analog[10].t45 5.713
R1569 io_analog[10].n41 io_analog[10].t43 5.713
R1570 io_analog[10].n39 io_analog[10].t15 5.713
R1571 io_analog[10].n39 io_analog[10].t12 5.713
R1572 io_analog[10].n37 io_analog[10].t42 5.713
R1573 io_analog[10].n37 io_analog[10].t37 5.713
R1574 io_analog[10].n35 io_analog[10].t39 5.713
R1575 io_analog[10].n35 io_analog[10].t30 5.713
R1576 io_analog[10].n33 io_analog[10].t20 5.713
R1577 io_analog[10].n33 io_analog[10].t44 5.713
R1578 io_analog[10].n31 io_analog[10].t34 5.713
R1579 io_analog[10].n31 io_analog[10].t25 5.713
R1580 io_analog[10].n29 io_analog[10].t26 5.713
R1581 io_analog[10].n29 io_analog[10].t22 5.713
R1582 io_analog[10].n27 io_analog[10].t13 5.713
R1583 io_analog[10].n27 io_analog[10].t49 5.713
R1584 io_analog[10].n25 io_analog[10].t21 5.713
R1585 io_analog[10].n25 io_analog[10].t18 5.713
R1586 io_analog[10].n23 io_analog[10].t36 5.713
R1587 io_analog[10].n23 io_analog[10].t32 5.713
R1588 io_analog[10].n21 io_analog[10].t48 5.713
R1589 io_analog[10].n21 io_analog[10].t40 5.713
R1590 io_analog[10].n19 io_analog[10].t17 5.713
R1591 io_analog[10].n19 io_analog[10].t10 5.713
R1592 io_analog[10].n17 io_analog[10].t23 5.713
R1593 io_analog[10].n17 io_analog[10].t35 5.713
R1594 io_analog[10].n0 io_analog[10].t38 5.713
R1595 io_analog[10].n0 io_analog[10].t33 5.713
R1596 io_analog[10].n51 io_analog[10].t31 5.713
R1597 io_analog[10].n51 io_analog[10].t27 5.713
R1598 io_analog[10].n16 io_analog[10].t51 4.096
R1599 io_analog[10].n5 io_analog[10].t7 4.096
R1600 io_analog[10].n14 io_analog[10].t6 3.48
R1601 io_analog[10].n14 io_analog[10].t2 3.48
R1602 io_analog[10].n12 io_analog[10].t3 3.48
R1603 io_analog[10].n12 io_analog[10].t8 3.48
R1604 io_analog[10].n10 io_analog[10].t0 3.48
R1605 io_analog[10].n10 io_analog[10].t1 3.48
R1606 io_analog[10].n8 io_analog[10].t50 3.48
R1607 io_analog[10].n8 io_analog[10].t9 3.48
R1608 io_analog[10].n6 io_analog[10].t4 3.48
R1609 io_analog[10].n6 io_analog[10].t5 3.48
R1610 io_analog[10].n55 io_analog[10].n54 1.013
R1611 io_analog[10] io_analog[10].n56 0.802
R1612 io_analog[10].n15 io_analog[10].n14 0.616
R1613 io_analog[10].n13 io_analog[10].n12 0.616
R1614 io_analog[10].n11 io_analog[10].n10 0.616
R1615 io_analog[10].n9 io_analog[10].n8 0.616
R1616 io_analog[10].n7 io_analog[10].n6 0.616
R1617 io_analog[10].n3 io_analog[10].n2 0.451
R1618 io_analog[10].n48 io_analog[10].n47 0.451
R1619 io_analog[10].n44 io_analog[10].n43 0.451
R1620 io_analog[10].n40 io_analog[10].n39 0.451
R1621 io_analog[10].n36 io_analog[10].n35 0.451
R1622 io_analog[10].n32 io_analog[10].n31 0.451
R1623 io_analog[10].n28 io_analog[10].n27 0.451
R1624 io_analog[10].n24 io_analog[10].n23 0.451
R1625 io_analog[10].n20 io_analog[10].n19 0.451
R1626 io_analog[10].n1 io_analog[10].n0 0.451
R1627 io_analog[10].n50 io_analog[10].n49 0.451
R1628 io_analog[10].n46 io_analog[10].n45 0.451
R1629 io_analog[10].n42 io_analog[10].n41 0.451
R1630 io_analog[10].n38 io_analog[10].n37 0.451
R1631 io_analog[10].n34 io_analog[10].n33 0.451
R1632 io_analog[10].n30 io_analog[10].n29 0.451
R1633 io_analog[10].n26 io_analog[10].n25 0.451
R1634 io_analog[10].n22 io_analog[10].n21 0.451
R1635 io_analog[10].n18 io_analog[10].n17 0.451
R1636 io_analog[10].n52 io_analog[10].n51 0.451
R1637 io_analog[10].n55 io_analog[10].n52 0.355
R1638 io_analog[10].n4 io_analog[10].n3 0.355
R1639 io_analog[10].n56 io_analog[10].n16 0.17
R1640 io_analog[10].t55 io_analog[10].t53 0.134
R1641 io_analog[10].t53 io_analog[10].n53 0.068
R1642 io_analog[10].n54 io_analog[10].t52 0.067
R1643 io_analog[10].n54 io_analog[10].t55 0.067
R1644 io_analog[10].n53 io_analog[10].t54 0.065
R1645 io_analog[10].n7 io_analog[10].n5 0.061
R1646 io_analog[10].n9 io_analog[10].n7 0.061
R1647 io_analog[10].n13 io_analog[10].n11 0.061
R1648 io_analog[10].n16 io_analog[10].n15 0.061
R1649 io_analog[10].n11 io_analog[10].n9 0.059
R1650 io_analog[10].n15 io_analog[10].n13 0.059
R1651 io_analog[10].n3 io_analog[10].n1 0.045
R1652 io_analog[10].n22 io_analog[10].n20 0.045
R1653 io_analog[10].n24 io_analog[10].n22 0.045
R1654 io_analog[10].n28 io_analog[10].n26 0.045
R1655 io_analog[10].n32 io_analog[10].n30 0.045
R1656 io_analog[10].n34 io_analog[10].n32 0.045
R1657 io_analog[10].n38 io_analog[10].n36 0.045
R1658 io_analog[10].n40 io_analog[10].n38 0.045
R1659 io_analog[10].n44 io_analog[10].n42 0.045
R1660 io_analog[10].n48 io_analog[10].n46 0.045
R1661 io_analog[10].n50 io_analog[10].n48 0.045
R1662 io_analog[10].n20 io_analog[10].n18 0.044
R1663 io_analog[10].n26 io_analog[10].n24 0.044
R1664 io_analog[10].n30 io_analog[10].n28 0.044
R1665 io_analog[10].n36 io_analog[10].n34 0.044
R1666 io_analog[10].n42 io_analog[10].n40 0.044
R1667 io_analog[10].n46 io_analog[10].n44 0.044
R1668 io_analog[10].n52 io_analog[10].n50 0.044
R1669 io_analog[9].n8 io_analog[9].t5 267.528
R1670 io_analog[9].n7 io_analog[9].t3 267.528
R1671 io_analog[9].n3 io_analog[9].t0 267.528
R1672 io_analog[9].n4 io_analog[9].t1 267.528
R1673 io_analog[9].n5 io_analog[9].t2 267.528
R1674 io_analog[9].n6 io_analog[9].t4 267.528
R1675 io_analog[9].n0 io_analog[9].t6 133.054
R1676 io_analog[9] io_analog[9].n13 2.539
R1677 io_analog[9].n1 io_analog[9].n0 1.817
R1678 io_analog[9].n13 io_analog[9].n12 1.293
R1679 io_analog[9].n13 io_analog[9].n6 1.293
R1680 io_analog[9].n8 io_analog[9].n7 0.395
R1681 io_analog[9].n9 io_analog[9].n8 0.395
R1682 io_analog[9].n10 io_analog[9].n9 0.395
R1683 io_analog[9].n11 io_analog[9].n10 0.395
R1684 io_analog[9].n12 io_analog[9].n11 0.395
R1685 io_analog[9].n2 io_analog[9].n1 0.395
R1686 io_analog[9].n3 io_analog[9].n2 0.395
R1687 io_analog[9].n4 io_analog[9].n3 0.395
R1688 io_analog[9].n5 io_analog[9].n4 0.395
R1689 io_analog[9].n6 io_analog[9].n5 0.395
R1690 a_43026_690892.n70 a_43026_690892.t34 272.261
R1691 a_43026_690892.n29 a_43026_690892.t36 272.261
R1692 a_43026_690892.n69 a_43026_690892.t24 271.866
R1693 a_43026_690892.n100 a_43026_690892.t20 271.866
R1694 a_43026_690892.n94 a_43026_690892.t26 271.866
R1695 a_43026_690892.n95 a_43026_690892.t40 271.866
R1696 a_43026_690892.n96 a_43026_690892.t18 271.866
R1697 a_43026_690892.n97 a_43026_690892.t6 271.866
R1698 a_43026_690892.n98 a_43026_690892.t10 271.866
R1699 a_43026_690892.n99 a_43026_690892.t14 271.866
R1700 a_43026_690892.n37 a_43026_690892.t16 271.866
R1701 a_43026_690892.n38 a_43026_690892.t38 271.866
R1702 a_43026_690892.n39 a_43026_690892.t32 271.866
R1703 a_43026_690892.n40 a_43026_690892.t4 271.866
R1704 a_43026_690892.n41 a_43026_690892.t2 271.866
R1705 a_43026_690892.n31 a_43026_690892.t12 271.866
R1706 a_43026_690892.n35 a_43026_690892.t30 271.866
R1707 a_43026_690892.n29 a_43026_690892.t0 271.866
R1708 a_43026_690892.n24 a_43026_690892.t69 271.866
R1709 a_43026_690892.n13 a_43026_690892.t65 271.866
R1710 a_43026_690892.n12 a_43026_690892.t63 271.866
R1711 a_43026_690892.n11 a_43026_690892.t54 271.866
R1712 a_43026_690892.n10 a_43026_690892.t68 271.866
R1713 a_43026_690892.n9 a_43026_690892.t67 271.866
R1714 a_43026_690892.n44 a_43026_690892.t53 271.866
R1715 a_43026_690892.n45 a_43026_690892.t50 271.866
R1716 a_43026_690892.n46 a_43026_690892.t61 271.866
R1717 a_43026_690892.n49 a_43026_690892.t58 271.866
R1718 a_43026_690892.n48 a_43026_690892.t56 271.866
R1719 a_43026_690892.n47 a_43026_690892.t49 271.866
R1720 a_43026_690892.n72 a_43026_690892.t60 271.866
R1721 a_43026_690892.n73 a_43026_690892.t66 271.866
R1722 a_43026_690892.n74 a_43026_690892.t64 271.866
R1723 a_43026_690892.n75 a_43026_690892.t62 271.866
R1724 a_43026_690892.n76 a_43026_690892.t59 271.866
R1725 a_43026_690892.n77 a_43026_690892.t57 271.866
R1726 a_43026_690892.n89 a_43026_690892.t55 271.866
R1727 a_43026_690892.n70 a_43026_690892.t28 271.866
R1728 a_43026_690892.n30 a_43026_690892.t8 271.866
R1729 a_43026_690892.n36 a_43026_690892.t22 271.866
R1730 a_43026_690892.n88 a_43026_690892.t52 135.324
R1731 a_43026_690892.n23 a_43026_690892.t51 135.322
R1732 a_43026_690892.n2 a_43026_690892.t35 6.295
R1733 a_43026_690892.n8 a_43026_690892.t1 5.713
R1734 a_43026_690892.n8 a_43026_690892.t37 5.713
R1735 a_43026_690892.n58 a_43026_690892.t33 5.713
R1736 a_43026_690892.n58 a_43026_690892.t5 5.713
R1737 a_43026_690892.n60 a_43026_690892.t17 5.713
R1738 a_43026_690892.n60 a_43026_690892.t39 5.713
R1739 a_43026_690892.n62 a_43026_690892.t27 5.713
R1740 a_43026_690892.n62 a_43026_690892.t23 5.713
R1741 a_43026_690892.n110 a_43026_690892.t11 5.713
R1742 a_43026_690892.n110 a_43026_690892.t7 5.713
R1743 a_43026_690892.n7 a_43026_690892.t21 5.713
R1744 a_43026_690892.n7 a_43026_690892.t15 5.713
R1745 a_43026_690892.n6 a_43026_690892.t3 5.713
R1746 a_43026_690892.n6 a_43026_690892.t31 5.713
R1747 a_43026_690892.n4 a_43026_690892.t13 5.713
R1748 a_43026_690892.n4 a_43026_690892.t9 5.713
R1749 a_43026_690892.n5 a_43026_690892.t29 5.713
R1750 a_43026_690892.n5 a_43026_690892.t25 5.713
R1751 a_43026_690892.n113 a_43026_690892.t19 5.713
R1752 a_43026_690892.t41 a_43026_690892.n113 5.713
R1753 a_43026_690892.n68 a_43026_690892.t45 3.802
R1754 a_43026_690892.n33 a_43026_690892.t47 3.48
R1755 a_43026_690892.n33 a_43026_690892.t43 3.48
R1756 a_43026_690892.n64 a_43026_690892.t42 3.48
R1757 a_43026_690892.n64 a_43026_690892.t48 3.48
R1758 a_43026_690892.n66 a_43026_690892.t44 3.48
R1759 a_43026_690892.n66 a_43026_690892.t46 3.48
R1760 a_43026_690892.n2 a_43026_690892.n68 2.808
R1761 a_43026_690892.n3 a_43026_690892.n34 2.807
R1762 a_43026_690892.n23 a_43026_690892.n22 1.617
R1763 a_43026_690892.n88 a_43026_690892.n87 1.615
R1764 a_43026_690892.n24 a_43026_690892.n23 1.222
R1765 a_43026_690892.n89 a_43026_690892.n88 1.22
R1766 a_43026_690892.n7 a_43026_690892.n108 1.177
R1767 a_43026_690892.n6 a_43026_690892.n57 1.177
R1768 a_43026_690892.n4 a_43026_690892.n28 1.177
R1769 a_43026_690892.n5 a_43026_690892.n93 1.125
R1770 a_43026_690892.n3 a_43026_690892.n8 0.582
R1771 a_43026_690892.n59 a_43026_690892.n58 0.532
R1772 a_43026_690892.n61 a_43026_690892.n60 0.532
R1773 a_43026_690892.n63 a_43026_690892.n62 0.532
R1774 a_43026_690892.n111 a_43026_690892.n110 0.532
R1775 a_43026_690892.n113 a_43026_690892.n112 0.53
R1776 a_43026_690892.n0 a_43026_690892.n7 0.421
R1777 a_43026_690892.n1 a_43026_690892.n6 0.421
R1778 a_43026_690892.n2 a_43026_690892.n5 0.421
R1779 a_43026_690892.n3 a_43026_690892.n4 0.421
R1780 a_43026_690892.n46 a_43026_690892.n45 0.395
R1781 a_43026_690892.n45 a_43026_690892.n44 0.395
R1782 a_43026_690892.n10 a_43026_690892.n9 0.395
R1783 a_43026_690892.n11 a_43026_690892.n10 0.395
R1784 a_43026_690892.n12 a_43026_690892.n11 0.395
R1785 a_43026_690892.n13 a_43026_690892.n12 0.395
R1786 a_43026_690892.n77 a_43026_690892.n76 0.395
R1787 a_43026_690892.n76 a_43026_690892.n75 0.395
R1788 a_43026_690892.n75 a_43026_690892.n74 0.395
R1789 a_43026_690892.n74 a_43026_690892.n73 0.395
R1790 a_43026_690892.n73 a_43026_690892.n72 0.395
R1791 a_43026_690892.n48 a_43026_690892.n47 0.395
R1792 a_43026_690892.n87 a_43026_690892.n86 0.395
R1793 a_43026_690892.n86 a_43026_690892.n85 0.395
R1794 a_43026_690892.n85 a_43026_690892.n84 0.395
R1795 a_43026_690892.n84 a_43026_690892.n83 0.395
R1796 a_43026_690892.n83 a_43026_690892.n82 0.395
R1797 a_43026_690892.n82 a_43026_690892.n81 0.395
R1798 a_43026_690892.n81 a_43026_690892.n80 0.395
R1799 a_43026_690892.n80 a_43026_690892.n79 0.395
R1800 a_43026_690892.n79 a_43026_690892.n78 0.395
R1801 a_43026_690892.n15 a_43026_690892.n14 0.395
R1802 a_43026_690892.n16 a_43026_690892.n15 0.395
R1803 a_43026_690892.n17 a_43026_690892.n16 0.395
R1804 a_43026_690892.n18 a_43026_690892.n17 0.395
R1805 a_43026_690892.n19 a_43026_690892.n18 0.395
R1806 a_43026_690892.n20 a_43026_690892.n19 0.395
R1807 a_43026_690892.n21 a_43026_690892.n20 0.395
R1808 a_43026_690892.n22 a_43026_690892.n21 0.395
R1809 a_43026_690892.n30 a_43026_690892.n29 0.395
R1810 a_43026_690892.n53 a_43026_690892.n52 0.395
R1811 a_43026_690892.n54 a_43026_690892.n53 0.395
R1812 a_43026_690892.n55 a_43026_690892.n54 0.395
R1813 a_43026_690892.n56 a_43026_690892.n55 0.395
R1814 a_43026_690892.n99 a_43026_690892.n98 0.395
R1815 a_43026_690892.n98 a_43026_690892.n97 0.395
R1816 a_43026_690892.n97 a_43026_690892.n96 0.395
R1817 a_43026_690892.n96 a_43026_690892.n95 0.395
R1818 a_43026_690892.n95 a_43026_690892.n94 0.395
R1819 a_43026_690892.n37 a_43026_690892.n36 0.395
R1820 a_43026_690892.n38 a_43026_690892.n37 0.395
R1821 a_43026_690892.n39 a_43026_690892.n38 0.395
R1822 a_43026_690892.n40 a_43026_690892.n39 0.395
R1823 a_43026_690892.n41 a_43026_690892.n40 0.395
R1824 a_43026_690892.n106 a_43026_690892.n105 0.395
R1825 a_43026_690892.n105 a_43026_690892.n104 0.395
R1826 a_43026_690892.n104 a_43026_690892.n103 0.395
R1827 a_43026_690892.n103 a_43026_690892.n102 0.395
R1828 a_43026_690892.n65 a_43026_690892.n64 0.322
R1829 a_43026_690892.n34 a_43026_690892.n33 0.322
R1830 a_43026_690892.n67 a_43026_690892.n66 0.322
R1831 a_43026_690892.n1 a_43026_690892.n42 0.27
R1832 a_43026_690892.n2 a_43026_690892.n71 0.268
R1833 a_43026_690892.n3 a_43026_690892.n32 0.267
R1834 a_43026_690892.n0 a_43026_690892.n101 0.271
R1835 a_43026_690892.n24 a_43026_690892.n13 0.255
R1836 a_43026_690892.n26 a_43026_690892.n25 0.255
R1837 a_43026_690892.n89 a_43026_690892.n77 0.25
R1838 a_43026_690892.n93 a_43026_690892.n92 0.2
R1839 a_43026_690892.n93 a_43026_690892.n91 0.195
R1840 a_43026_690892.n91 a_43026_690892.n90 0.192
R1841 a_43026_690892.n25 a_43026_690892.n24 0.189
R1842 a_43026_690892.n51 a_43026_690892.n49 0.189
R1843 a_43026_690892.n90 a_43026_690892.n89 0.178
R1844 a_43026_690892.n42 a_43026_690892.n35 0.13
R1845 a_43026_690892.n57 a_43026_690892.n43 0.13
R1846 a_43026_690892.n108 a_43026_690892.n107 0.13
R1847 a_43026_690892.n101 a_43026_690892.n100 0.13
R1848 a_43026_690892.n32 a_43026_690892.n31 0.125
R1849 a_43026_690892.n28 a_43026_690892.n27 0.125
R1850 a_43026_690892.n71 a_43026_690892.n69 0.125
R1851 a_43026_690892.n28 a_43026_690892.n26 0.12
R1852 a_43026_690892.n32 a_43026_690892.n30 0.12
R1853 a_43026_690892.n71 a_43026_690892.n70 0.12
R1854 a_43026_690892.n57 a_43026_690892.n56 0.115
R1855 a_43026_690892.n101 a_43026_690892.n99 0.115
R1856 a_43026_690892.n42 a_43026_690892.n41 0.115
R1857 a_43026_690892.n108 a_43026_690892.n106 0.115
R1858 a_43026_690892.n49 a_43026_690892.n48 0.06
R1859 a_43026_690892.n51 a_43026_690892.n50 0.06
R1860 a_43026_690892.n49 a_43026_690892.n46 0.055
R1861 a_43026_690892.n52 a_43026_690892.n51 0.055
R1862 a_43026_690892.n111 a_43026_690892.n0 0.05
R1863 a_43026_690892.n112 a_43026_690892.n63 0.05
R1864 a_43026_690892.n63 a_43026_690892.n61 0.05
R1865 a_43026_690892.n59 a_43026_690892.n1 0.05
R1866 a_43026_690892.n1 a_43026_690892.n3 0.049
R1867 a_43026_690892.n0 a_43026_690892.n2 0.049
R1868 a_43026_690892.n112 a_43026_690892.n111 0.048
R1869 a_43026_690892.n61 a_43026_690892.n59 0.048
R1870 a_43026_690892.n68 a_43026_690892.n67 0.039
R1871 a_43026_690892.n67 a_43026_690892.n65 0.039
R1872 a_43026_690892.n0 a_43026_690892.n109 0.006
R1873 a_42818_684860.n19 a_42818_684860.t3 4.1
R1874 a_42818_684860.n6 a_42818_684860.t1 4.096
R1875 a_42818_684860.n9 a_42818_684860.t8 3.802
R1876 a_42818_684860.n25 a_42818_684860.t16 3.797
R1877 a_42818_684860.n26 a_42818_684860.t19 3.48
R1878 a_42818_684860.n26 a_42818_684860.t18 3.48
R1879 a_42818_684860.n11 a_42818_684860.t14 3.48
R1880 a_42818_684860.n11 a_42818_684860.t17 3.48
R1881 a_42818_684860.n20 a_42818_684860.t13 3.48
R1882 a_42818_684860.n20 a_42818_684860.t0 3.48
R1883 a_42818_684860.n7 a_42818_684860.t11 3.48
R1884 a_42818_684860.n7 a_42818_684860.t23 3.48
R1885 a_42818_684860.n22 a_42818_684860.t21 3.48
R1886 a_42818_684860.n22 a_42818_684860.t22 3.48
R1887 a_42818_684860.n17 a_42818_684860.t4 3.48
R1888 a_42818_684860.n17 a_42818_684860.t25 3.48
R1889 a_42818_684860.n15 a_42818_684860.t9 3.48
R1890 a_42818_684860.n15 a_42818_684860.t2 3.48
R1891 a_42818_684860.n13 a_42818_684860.t7 3.48
R1892 a_42818_684860.n13 a_42818_684860.t27 3.48
R1893 a_42818_684860.n0 a_42818_684860.t5 3.48
R1894 a_42818_684860.n0 a_42818_684860.t10 3.48
R1895 a_42818_684860.n2 a_42818_684860.t12 3.48
R1896 a_42818_684860.n2 a_42818_684860.t6 3.48
R1897 a_42818_684860.n4 a_42818_684860.t26 3.48
R1898 a_42818_684860.n4 a_42818_684860.t24 3.48
R1899 a_42818_684860.n29 a_42818_684860.t15 3.48
R1900 a_42818_684860.t20 a_42818_684860.n29 3.48
R1901 a_42818_684860.n24 a_42818_684860.n19 2.175
R1902 a_42818_684860.n10 a_42818_684860.n6 2.175
R1903 a_42818_684860.n24 a_42818_684860.n23 0.75
R1904 a_42818_684860.n10 a_42818_684860.n9 0.73
R1905 a_42818_684860.n18 a_42818_684860.n17 0.616
R1906 a_42818_684860.n16 a_42818_684860.n15 0.616
R1907 a_42818_684860.n14 a_42818_684860.n13 0.616
R1908 a_42818_684860.n1 a_42818_684860.n0 0.616
R1909 a_42818_684860.n3 a_42818_684860.n2 0.616
R1910 a_42818_684860.n5 a_42818_684860.n4 0.616
R1911 a_42818_684860.n23 a_42818_684860.n22 0.323
R1912 a_42818_684860.n8 a_42818_684860.n7 0.322
R1913 a_42818_684860.n21 a_42818_684860.n20 0.322
R1914 a_42818_684860.n27 a_42818_684860.n26 0.321
R1915 a_42818_684860.n12 a_42818_684860.n11 0.317
R1916 a_42818_684860.n29 a_42818_684860.n28 0.316
R1917 a_42818_684860.n12 a_42818_684860.n10 0.172
R1918 a_42818_684860.n25 a_42818_684860.n24 0.152
R1919 a_42818_684860.n5 a_42818_684860.n3 0.09
R1920 a_42818_684860.n3 a_42818_684860.n1 0.09
R1921 a_42818_684860.n16 a_42818_684860.n14 0.09
R1922 a_42818_684860.n19 a_42818_684860.n18 0.09
R1923 a_42818_684860.n6 a_42818_684860.n5 0.088
R1924 a_42818_684860.n18 a_42818_684860.n16 0.088
R1925 a_42818_684860.n9 a_42818_684860.n8 0.039
R1926 a_42818_684860.n28 a_42818_684860.n12 0.039
R1927 a_42818_684860.n27 a_42818_684860.n25 0.039
R1928 a_42818_684860.n23 a_42818_684860.n21 0.038
R1929 a_42818_684860.n28 a_42818_684860.n27 0.038
R1930 vssa2.n4 vssa2.t31 3613.01
R1931 vssa2.n5 vssa2.t134 3613.01
R1932 vssa2.n119 vssa2.n118 3505.44
R1933 vssa2.t59 vssa2.t1 3317.89
R1934 vssa2.t42 vssa2.t141 3317.89
R1935 vssa2.n200 vssa2.n184 3302.65
R1936 vssa2 vssa2.t79 2616.22
R1937 vssa2 vssa2.t98 2579.05
R1938 vssa2.t99 vssa2.n69 1922.76
R1939 vssa2.t58 vssa2.n70 1922.76
R1940 vssa2.t2 vssa2.t58 3872.36
R1941 vssa2.t43 vssa2.t99 3872.36
R1942 vssa2 vssa2.t69 1797.69
R1943 vssa2 vssa2.t82 1797.69
R1944 vssa2 vssa2.t33 1797.69
R1945 vssa2 vssa2.t80 1797.69
R1946 vssa2.n200 vssa2.n199 1749.82
R1947 vssa2.t46 vssa2.n122 1708.05
R1948 vssa2 vssa2.n137 1708.05
R1949 vssa2.n122 vssa2.t91 1708.05
R1950 vssa2.n137 vssa2.t108 1708.05
R1951 vssa2.t20 vssa2.n47 1689.22
R1952 vssa2.t133 vssa2.n58 1689.22
R1953 vssa2.n47 vssa2.t42 1689.22
R1954 vssa2.n58 vssa2.t59 1689.22
R1955 vssa2.n196 vssa2.n194 1478.78
R1956 vssa2.n194 vssa2.n189 1478.78
R1957 vssa2 vssa2.n284 1367.57
R1958 vssa2.n240 vssa2.t8 1252.03
R1959 vssa2.n256 vssa2.t85 1234.15
R1960 vssa2.n288 vssa2.n285 1066.12
R1961 vssa2.n444 vssa2.t93 847.164
R1962 vssa2.t62 vssa2.t75 799.436
R1963 vssa2.t119 vssa2.t131 799.436
R1964 vssa2.t16 vssa2.t119 799.436
R1965 vssa2.t21 vssa2.t60 799.436
R1966 vssa2.t60 vssa2.t117 799.436
R1967 vssa2.t55 vssa2.t77 799.436
R1968 vssa2.t144 vssa2.t18 799.436
R1969 vssa2.t129 vssa2.t87 799.436
R1970 vssa2.t39 vssa2.t49 799.436
R1971 vssa2.t66 vssa2.t39 799.436
R1972 vssa2.t53 vssa2.t149 799.436
R1973 vssa2.t149 vssa2.t64 799.436
R1974 vssa2.t37 vssa2.t23 799.436
R1975 vssa2.t138 vssa2.t26 799.436
R1976 vssa2 vssa2.n89 763.858
R1977 vssa2 vssa2.t5 761.791
R1978 vssa2.n369 vssa2.t129 728.169
R1979 vssa2.n361 vssa2.t37 728.169
R1980 vssa2.n114 vssa2.n109 709.647
R1981 vssa2.n114 vssa2.n113 709.647
R1982 vssa2 vssa2.n19 692.328
R1983 vssa2 vssa2.n24 692.328
R1984 vssa2.n305 vssa2.n302 688.563
R1985 vssa2.n419 vssa2.t89 672.394
R1986 vssa2.n377 vssa2.t146 669.295
R1987 vssa2.n347 vssa2.n346 662.21
R1988 vssa2.n496 vssa2.t156 585.633
R1989 vssa2.n149 vssa2.n148 585
R1990 vssa2 vssa2.n149 585
R1991 vssa2.n134 vssa2.n133 585
R1992 vssa2 vssa2.n134 585
R1993 vssa2.n139 vssa2.n138 585
R1994 vssa2.n120 vssa2.n119 585
R1995 vssa2.n141 vssa2.n140 585
R1996 vssa2 vssa2.n141 585
R1997 vssa2.n124 vssa2.n123 585
R1998 vssa2.t46 vssa2.n124 585
R1999 vssa2 vssa2.n142 585
R2000 vssa2.n144 vssa2.n143 585
R2001 vssa2 vssa2.n144 585
R2002 vssa2.n126 vssa2.n125 585
R2003 vssa2.t46 vssa2.n126 585
R2004 vssa2.n147 vssa2.n146 585
R2005 vssa2 vssa2.n147 585
R2006 vssa2.n132 vssa2.n131 585
R2007 vssa2 vssa2.n132 585
R2008 vssa2.n51 vssa2.n50 585
R2009 vssa2.n36 vssa2.n35 585
R2010 vssa2.n35 vssa2.n34 585
R2011 vssa2.n29 vssa2.n28 585
R2012 vssa2.n28 vssa2.n27 585
R2013 vssa2.n72 vssa2.n71 585
R2014 vssa2.n4 vssa2.n72 585
R2015 vssa2.n74 vssa2.n73 585
R2016 vssa2.n5 vssa2.n74 585
R2017 vssa2.n54 vssa2.n53 585
R2018 vssa2.n53 vssa2.n52 585
R2019 vssa2.n43 vssa2.n42 585
R2020 vssa2.n42 vssa2.n41 585
R2021 vssa2.n65 vssa2.n64 585
R2022 vssa2.n60 vssa2.n59 585
R2023 vssa2.n49 vssa2.n48 585
R2024 vssa2 vssa2.n91 585
R2025 vssa2.n0 vssa2.n104 585
R2026 vssa2.n21 vssa2.n20 585
R2027 vssa2.t128 vssa2.n14 585
R2028 vssa2 vssa2.n183 585
R2029 vssa2.n199 vssa2.n197 585
R2030 vssa2.n187 vssa2.n186 585
R2031 vssa2.n288 vssa2.n287 585
R2032 vssa2 vssa2.n288 585
R2033 vssa2 vssa2.n174 585
R2034 vssa2.n272 vssa2.n271 585
R2035 vssa2.n244 vssa2.n243 585
R2036 vssa2.n243 vssa2.n242 585
R2037 vssa2.n207 vssa2.n206 585
R2038 vssa2.n206 vssa2.n205 585
R2039 vssa2.n277 vssa2.n276 585
R2040 vssa2.n276 vssa2.n275 585
R2041 vssa2.n260 vssa2.n259 585
R2042 vssa2.n259 vssa2.n258 585
R2043 vssa2.n263 vssa2.n262 585
R2044 vssa2.n262 vssa2.n261 585
R2045 vssa2.n250 vssa2.n249 585
R2046 vssa2.n249 vssa2.n248 585
R2047 vssa2.n247 vssa2.n246 585
R2048 vssa2.n246 vssa2.n245 585
R2049 vssa2.n10 vssa2.n9 575.622
R2050 vssa2.n0 vssa2.n103 541.74
R2051 vssa2.n489 vssa2.t148 532.957
R2052 vssa2 vssa2.n90 530.069
R2053 vssa2.n305 vssa2.n304 490.916
R2054 vssa2.t105 vssa2.t126 489.577
R2055 vssa2.t105 vssa2.t11 489.577
R2056 vssa2.t116 vssa2.t111 489.577
R2057 vssa2.t116 vssa2.t115 489.577
R2058 vssa2 vssa2.n201 483.108
R2059 vssa2 vssa2.n21 483.01
R2060 vssa2.n3 vssa2.n350 477.363
R2061 vssa2 vssa2.t51 453.378
R2062 vssa2.n371 vssa2.n368 438.211
R2063 vssa2.n363 vssa2.n360 438.211
R2064 vssa2.n394 vssa2.t123 436.901
R2065 vssa2.n383 vssa2.t114 436.901
R2066 vssa2.n402 vssa2.t73 433.802
R2067 vssa2.n413 vssa2.t113 433.802
R2068 vssa2.n269 vssa2.n268 416.794
R2069 vssa2.n421 vssa2.n418 414.117
R2070 vssa2.n379 vssa2.n374 413.741
R2071 vssa2.n498 vssa2.n493 403.576
R2072 vssa2.n430 vssa2.t137 399.718
R2073 vssa2.n423 vssa2.t16 399.718
R2074 vssa2.n423 vssa2.t21 399.718
R2075 vssa2.n423 vssa2.t66 399.718
R2076 vssa2.n423 vssa2.t53 399.718
R2077 vssa2.n491 vssa2.n486 397.176
R2078 vssa2.n439 vssa2.t3 380.895
R2079 vssa2.n454 vssa2.t86 377.826
R2080 vssa2.n454 vssa2.t122 377.826
R2081 vssa2 vssa2.t157 350.14
R2082 vssa2.t46 vssa2.n120 326.776
R2083 vssa2 vssa2.n139 326.776
R2084 vssa2.n358 vssa2.n357 324.544
R2085 vssa2.n364 vssa2.n363 324.48
R2086 vssa2.n358 vssa2.n355 323.788
R2087 vssa2.n372 vssa2.n371 323.722
R2088 vssa2.n404 vssa2.n399 320.376
R2089 vssa2.n415 vssa2.n412 320.376
R2090 vssa2.n396 vssa2.n391 319.999
R2091 vssa2.n385 vssa2.n382 319.999
R2092 vssa2.n199 vssa2.n198 305.227
R2093 vssa2.t20 vssa2.n49 300.422
R2094 vssa2.t133 vssa2.n51 300.422
R2095 vssa2.n186 vssa2.n185 300.071
R2096 vssa2 vssa2.n25 299.367
R2097 vssa2.n436 vssa2.t9 295.522
R2098 vssa2.n372 vssa2.n366 275.361
R2099 vssa2.n422 vssa2.n421 275.36
R2100 vssa2.n380 vssa2.n379 272.564
R2101 vssa2.n489 vssa2.t121 266.478
R2102 vssa2 vssa2.t103 260.135
R2103 vssa2.t32 vssa2.n1 232.13
R2104 vssa2.n261 vssa2.t136 215.54
R2105 vssa2.n496 vssa2.t25 213.802
R2106 vssa2.n189 vssa2.n187 213.458
R2107 vssa2.t128 vssa2.n16 208.955
R2108 vssa2 vssa2.t14 200.675
R2109 vssa2.n197 vssa2.n196 194.258
R2110 vssa2 vssa2.t71 185.81
R2111 vssa2.n100 vssa2.n92 173.823
R2112 vssa2.n457 vssa2.n456 164.894
R2113 vssa2.n16 vssa2.n15 156.716
R2114 vssa2 vssa2.t152 156.081
R2115 vssa2 vssa2.n491 146.536
R2116 vssa2.n66 vssa2.n65 144.941
R2117 vssa2.n61 vssa2.n60 144.941
R2118 vssa2.n499 vssa2.n498 143.717
R2119 vssa2.n37 vssa2.n36 141.176
R2120 vssa2.n30 vssa2.n29 141.176
R2121 vssa2.n377 vssa2.t55 130.14
R2122 vssa2.n218 vssa2.n215 127.623
R2123 vssa2.n419 vssa2.t62 127.042
R2124 vssa2.n272 vssa2.n270 120.846
R2125 vssa2.n446 vssa2.n441 117.816
R2126 vssa2 vssa2.n438 117.082
R2127 vssa2.n24 vssa2.n23 107.294
R2128 vssa2.n19 vssa2.t128 107.294
R2129 vssa2.n264 vssa2.n263 101.647
R2130 vssa2.n408 vssa2.n404 86.452
R2131 vssa2.n397 vssa2.n396 86.45
R2132 vssa2.n386 vssa2.n385 86.45
R2133 vssa2.n407 vssa2.n406 86.211
R2134 vssa2.n389 vssa2.n388 86.211
R2135 vssa2.n416 vssa2.n415 86.211
R2136 vssa2.n55 vssa2.n54 81.317
R2137 vssa2.n44 vssa2.n43 81.317
R2138 vssa2.n251 vssa2.n250 77.176
R2139 vssa2.n369 vssa2.t144 71.267
R2140 vssa2.n361 vssa2.t138 71.267
R2141 vssa2.n251 vssa2.n244 71.152
R2142 vssa2.n264 vssa2.n260 70.776
R2143 vssa2.n287 vssa2.n286 69.27
R2144 vssa2.n280 vssa2.n279 67.906
R2145 vssa2 vssa2.n128 66.891
R2146 vssa2.n219 vssa2.n213 66.258
R2147 vssa2 vssa2.n267 62.117
R2148 vssa2.n280 vssa2.n277 62.117
R2149 vssa2.n208 vssa2.n207 56.47
R2150 vssa2.n208 vssa2.n204 56.47
R2151 vssa2.n402 vssa2.t57 55.774
R2152 vssa2.n413 vssa2.t110 55.774
R2153 vssa2.n394 vssa2.t124 52.676
R2154 vssa2.n383 vssa2.t112 52.676
R2155 vssa2.n132 vssa2.n129 52.147
R2156 vssa2.n346 vssa2.n345 46.592
R2157 vssa2.t140 vssa2.n99 44.776
R2158 vssa2.n302 vssa2.n301 39.424
R2159 vssa2.n182 vssa2.n178 37.647
R2160 vssa2.n182 vssa2.n181 37.647
R2161 vssa2.n234 vssa2.n233 37.27
R2162 vssa2.n234 vssa2.n224 36.517
R2163 vssa2.n250 vssa2.n247 33.882
R2164 vssa2.n245 vssa2.t95 29.729
R2165 vssa2.n301 vssa2.n289 28.16
R2166 vssa2.n219 vssa2.n218 27.314
R2167 vssa2.t46 vssa2.n127 23.176
R2168 vssa2 vssa2.n145 23.176
R2169 vssa2.n339 vssa2.n338 22.199
R2170 vssa2.n345 vssa2.n336 20.992
R2171 vssa2 vssa2.t52 13.954
R2172 vssa2 vssa2.t72 13.95
R2173 vssa2 vssa2.t153 13.948
R2174 vssa2 vssa2.t15 13.948
R2175 vssa2.n484 vssa2.t10 13.926
R2176 vssa2.n474 vssa2.t4 13.924
R2177 vssa2 vssa2.t94 13.92
R2178 vssa2 vssa2.t6 13.92
R2179 vssa2.n89 vssa2.n88 13.575
R2180 vssa2 vssa2.n272 13.532
R2181 vssa2.n102 vssa2.n101 11.294
R2182 vssa2.n295 vssa2.n294 9.952
R2183 vssa2 vssa2.n102 9.833
R2184 vssa2 vssa2.n499 9.383
R2185 vssa2 vssa2.n154 9.3
R2186 vssa2 vssa2.n151 9.3
R2187 vssa2 vssa2.n157 9.3
R2188 vssa2 vssa2.n159 9.3
R2189 vssa2 vssa2.n161 9.3
R2190 vssa2 vssa2.n155 9.3
R2191 vssa2 vssa2.n163 9.3
R2192 vssa2 vssa2.n165 9.3
R2193 vssa2 vssa2.n171 9.3
R2194 vssa2 vssa2.n172 9.3
R2195 vssa2.n33 vssa2.n32 9.3
R2196 vssa2.n32 vssa2.n31 9.3
R2197 vssa2.n40 vssa2.n39 9.3
R2198 vssa2.n39 vssa2.n38 9.3
R2199 vssa2.n78 vssa2.n77 9.3
R2200 vssa2.n77 vssa2.n76 9.3
R2201 vssa2.n82 vssa2.n81 9.3
R2202 vssa2.n81 vssa2.n80 9.3
R2203 vssa2.n63 vssa2.n62 9.3
R2204 vssa2.n68 vssa2.n67 9.3
R2205 vssa2 vssa2.n105 9.3
R2206 vssa2 vssa2.n26 9.3
R2207 vssa2.n201 vssa2.n200 9.3
R2208 vssa2 vssa2.n283 9.3
R2209 vssa2.n283 vssa2.n282 9.3
R2210 vssa2.n211 vssa2.n210 9.3
R2211 vssa2 vssa2.n236 9.3
R2212 vssa2.n236 vssa2.n235 9.3
R2213 vssa2 vssa2.n177 9.3
R2214 vssa2.n177 vssa2.n176 9.3
R2215 vssa2.n281 vssa2.n274 9.3
R2216 vssa2 vssa2.n257 9.3
R2217 vssa2.n257 vssa2.n256 9.3
R2218 vssa2 vssa2.n254 9.3
R2219 vssa2.n254 vssa2.n253 9.3
R2220 vssa2 vssa2.n241 9.3
R2221 vssa2.n241 vssa2.n240 9.3
R2222 vssa2 vssa2.n239 9.3
R2223 vssa2.n239 vssa2.n238 9.3
R2224 vssa2.n105 vssa2.n0 9.3
R2225 vssa2.n231 vssa2.n226 8.943
R2226 vssa2 vssa2.n234 8.138
R2227 vssa2 vssa2.n237 8.138
R2228 vssa2 vssa2.n175 8.138
R2229 vssa2 vssa2.n182 8.138
R2230 vssa2.n128 vssa2.t46 7.432
R2231 vssa2 vssa2.n264 6.658
R2232 vssa2 vssa2.n255 6.658
R2233 vssa2 vssa2.n252 6.658
R2234 vssa2 vssa2.n251 6.658
R2235 vssa2 vssa2.n87 6.476
R2236 vssa2 vssa2.n114 6.476
R2237 vssa2.n296 vssa2.n295 6.247
R2238 vssa2.n274 vssa2.n273 5.984
R2239 vssa2 vssa2.t84 5.911
R2240 vssa2 vssa2.t104 5.911
R2241 vssa2.n232 vssa2.n225 5.794
R2242 vssa2.n230 vssa2.n227 5.794
R2243 vssa2.n210 vssa2.n209 5.78
R2244 vssa2.n168 vssa2.t109 5.763
R2245 vssa2 vssa2.n117 5.189
R2246 vssa2 vssa2.n135 5.189
R2247 vssa2 vssa2.n153 5.189
R2248 vssa2 vssa2.n156 5.189
R2249 vssa2 vssa2.n162 5.189
R2250 vssa2 vssa2.n160 5.189
R2251 vssa2 vssa2.n166 5.189
R2252 vssa2 vssa2.n164 5.189
R2253 vssa2 vssa2.n173 5.189
R2254 vssa2 vssa2.n167 5.189
R2255 vssa2 vssa2.n435 5.12
R2256 vssa2 vssa2.t92 4.374
R2257 vssa2 vssa2.n158 4.324
R2258 vssa2.n340 vssa2.n339 4.245
R2259 vssa2 vssa2.n446 4.16
R2260 vssa2 vssa2.n150 3.632
R2261 vssa2.n433 vssa2.n432 3.52
R2262 vssa2 vssa2.n211 3.507
R2263 vssa2 vssa2.t155 3.482
R2264 vssa2 vssa2.t47 3.482
R2265 vssa2.n325 vssa2.t118 3.48
R2266 vssa2.n325 vssa2.t78 3.48
R2267 vssa2.n323 vssa2.t22 3.48
R2268 vssa2.n323 vssa2.t61 3.48
R2269 vssa2.n318 vssa2.t120 3.48
R2270 vssa2.n318 vssa2.t17 3.48
R2271 vssa2.n320 vssa2.t76 3.48
R2272 vssa2.n320 vssa2.t132 3.48
R2273 vssa2.n317 vssa2.t90 3.48
R2274 vssa2.n317 vssa2.t63 3.48
R2275 vssa2.n322 vssa2.t56 3.48
R2276 vssa2.n322 vssa2.t147 3.48
R2277 vssa2.n316 vssa2.t19 3.48
R2278 vssa2.n316 vssa2.t145 3.48
R2279 vssa2.n331 vssa2.t139 3.48
R2280 vssa2.n331 vssa2.t27 3.48
R2281 vssa2.n329 vssa2.t24 3.48
R2282 vssa2.n329 vssa2.t38 3.48
R2283 vssa2.n327 vssa2.t150 3.48
R2284 vssa2.n327 vssa2.t65 3.48
R2285 vssa2.n310 vssa2.t67 3.48
R2286 vssa2.n310 vssa2.t54 3.48
R2287 vssa2.n312 vssa2.t50 3.48
R2288 vssa2.n312 vssa2.t40 3.48
R2289 vssa2.n314 vssa2.t130 3.48
R2290 vssa2.n314 vssa2.t88 3.48
R2291 vssa2 vssa2.t30 3.48
R2292 vssa2 vssa2.t135 3.48
R2293 vssa2 vssa2.t107 3.48
R2294 vssa2 vssa2.t143 3.48
R2295 vssa2 vssa2.t13 3.48
R2296 vssa2.n168 vssa2.t142 3.48
R2297 vssa2.n170 vssa2.t68 3.48
R2298 vssa2.n169 vssa2.t102 3.48
R2299 vssa2.n152 vssa2.t97 3.48
R2300 vssa2 vssa2.t154 3.48
R2301 vssa2 vssa2.t12 3.48
R2302 vssa2.n84 vssa2.t83 3.48
R2303 vssa2.n83 vssa2.t96 3.48
R2304 vssa2.n116 vssa2.t29 3.48
R2305 vssa2 vssa2.t34 3.48
R2306 vssa2.n115 vssa2.t45 3.48
R2307 vssa2.n85 vssa2.t36 3.48
R2308 vssa2.n86 vssa2.t81 3.48
R2309 vssa2 vssa2.t101 3.48
R2310 vssa2 vssa2.t70 3.48
R2311 vssa2 vssa2.n78 3.451
R2312 vssa2 vssa2.n40 3.45
R2313 vssa2 vssa2.t133 3.45
R2314 vssa2 vssa2.n63 3.45
R2315 vssa2 vssa2.n68 3.45
R2316 vssa2 vssa2.n82 3.45
R2317 vssa2 vssa2.n33 3.45
R2318 vssa2 vssa2.t20 3.45
R2319 vssa2 vssa2.t2 3.45
R2320 vssa2 vssa2.t43 3.45
R2321 vssa2 vssa2.n5 3.45
R2322 vssa2 vssa2.n4 3.45
R2323 vssa2.n131 vssa2.n130 3.388
R2324 vssa2 vssa2.n281 2.566
R2325 vssa2.n211 vssa2.n208 2.515
R2326 vssa2.n86 vssa2.n85 2.465
R2327 vssa2.n84 vssa2.n83 2.465
R2328 vssa2 vssa2.n86 2.445
R2329 vssa2 vssa2.n84 2.444
R2330 vssa2 vssa2.n115 2.428
R2331 vssa2 vssa2.n116 2.427
R2332 vssa2 vssa2.t41 2.413
R2333 vssa2 vssa2.t0 2.412
R2334 vssa2 vssa2.t125 2.412
R2335 vssa2 vssa2.t127 2.412
R2336 vssa2 vssa2.t7 2.412
R2337 vssa2 vssa2.t106 2.412
R2338 vssa2 vssa2.t74 2.412
R2339 vssa2 vssa2.t151 2.412
R2340 vssa2.n170 vssa2.n169 2.283
R2341 vssa2 vssa2.n170 2.261
R2342 vssa2 vssa2.n152 2.243
R2343 vssa2 vssa2.n168 2.24
R2344 vssa2 vssa2.n219 2.201
R2345 vssa2 vssa2.n433 1.6
R2346 vssa2.n33 vssa2.n30 1.163
R2347 vssa2.n78 vssa2.n75 1.163
R2348 vssa2.n63 vssa2.n61 1.163
R2349 vssa2.n281 vssa2.n280 1.066
R2350 vssa2.n40 vssa2.n37 1.047
R2351 vssa2.n82 vssa2.n79 1.047
R2352 vssa2.n68 vssa2.n66 1.047
R2353 vssa2.n386 vssa2.n380 0.908
R2354 vssa2 vssa2.n429 0.876
R2355 vssa2.n218 vssa2.n217 0.794
R2356 vssa2.n352 vssa2.n331 0.661
R2357 vssa2.n424 vssa2.n317 0.661
R2358 vssa2.n353 vssa2.n322 0.661
R2359 vssa2.n425 vssa2.n316 0.659
R2360 vssa2.n324 vssa2.n323 0.616
R2361 vssa2.n321 vssa2.n320 0.616
R2362 vssa2.n330 vssa2.n329 0.616
R2363 vssa2.n328 vssa2.n327 0.616
R2364 vssa2.n311 vssa2.n310 0.616
R2365 vssa2.n313 vssa2.n312 0.616
R2366 vssa2.n315 vssa2.n314 0.616
R2367 vssa2.n326 vssa2.n325 0.616
R2368 vssa2.n319 vssa2.n318 0.616
R2369 vssa2.n217 vssa2.n216 0.557
R2370 vssa2.n351 vssa2.n3 0.539
R2371 vssa2.n309 vssa2.n2 0.534
R2372 vssa2.n229 vssa2.n228 0.376
R2373 vssa2.n422 vssa2.n416 0.242
R2374 vssa2.n408 vssa2.n407 0.242
R2375 vssa2.n397 vssa2.n389 0.24
R2376 vssa2.n481 vssa2.n480 0.218
R2377 vssa2.n471 vssa2.n470 0.218
R2378 vssa2.n477 vssa2.n476 0.218
R2379 vssa2.n480 vssa2.n479 0.218
R2380 vssa2.n476 vssa2.n475 0.218
R2381 vssa2.n470 vssa2.n469 0.218
R2382 vssa2.n467 vssa2.n464 0.201
R2383 vssa2.n464 vssa2.n463 0.201
R2384 vssa2 vssa2.n484 0.189
R2385 vssa2 vssa2.n474 0.188
R2386 vssa2.n181 vssa2.n180 0.162
R2387 vssa2.n180 vssa2.n179 0.162
R2388 vssa2 vssa2.n458 0.155
R2389 vssa2.n462 vssa2.n461 0.155
R2390 vssa2 vssa2.n462 0.155
R2391 vssa2.n458 vssa2.n457 0.155
R2392 vssa2.n352 vssa2.n351 0.147
R2393 vssa2 vssa2.n449 0.146
R2394 vssa2.n449 vssa2.n448 0.146
R2395 vssa2.n460 vssa2.n459 0.146
R2396 vssa2 vssa2.n460 0.146
R2397 vssa2.n426 vssa2.n425 0.141
R2398 vssa2.n474 vssa2.n473 0.14
R2399 vssa2.n338 vssa2.n337 0.131
R2400 vssa2.n294 vssa2.n293 0.131
R2401 vssa2.n484 vssa2.n483 0.126
R2402 vssa2 vssa2.n447 0.121
R2403 vssa2.n394 vssa2.n393 0.118
R2404 vssa2.n402 vssa2.n401 0.118
R2405 vssa2.n396 vssa2.n395 0.118
R2406 vssa2.n395 vssa2.n394 0.118
R2407 vssa2.n404 vssa2.n403 0.118
R2408 vssa2.n403 vssa2.n402 0.118
R2409 vssa2.n388 vssa2.n387 0.118
R2410 vssa2.n406 vssa2.n405 0.118
R2411 vssa2.n385 vssa2.n384 0.118
R2412 vssa2.n384 vssa2.n383 0.118
R2413 vssa2.n415 vssa2.n414 0.118
R2414 vssa2.n414 vssa2.n413 0.118
R2415 vssa2.n401 vssa2.n400 0.111
R2416 vssa2.n393 vssa2.n392 0.111
R2417 vssa2.n204 vssa2.n203 0.101
R2418 vssa2.n203 vssa2.n202 0.101
R2419 vssa2.n267 vssa2.n266 0.091
R2420 vssa2.n266 vssa2.n265 0.091
R2421 vssa2.n326 vssa2.n324 0.09
R2422 vssa2.n315 vssa2.n313 0.09
R2423 vssa2.n330 vssa2.n328 0.09
R2424 vssa2.n321 vssa2.n319 0.088
R2425 vssa2.n313 vssa2.n311 0.088
R2426 vssa2.n467 vssa2.n466 0.072
R2427 vssa2.n466 vssa2.n465 0.072
R2428 vssa2.n438 vssa2.n437 0.07
R2429 vssa2.n437 vssa2.n436 0.07
R2430 vssa2.n213 vssa2.n212 0.07
R2431 vssa2.n279 vssa2.n278 0.07
R2432 vssa2.t105 vssa2.n397 0.067
R2433 vssa2.t116 vssa2.n386 0.067
R2434 vssa2.t105 vssa2.n408 0.066
R2435 vssa2.n441 vssa2.n440 0.065
R2436 vssa2.n440 vssa2.n439 0.065
R2437 vssa2.n423 vssa2.n372 0.064
R2438 vssa2.n423 vssa2.n422 0.064
R2439 vssa2.n423 vssa2.n364 0.063
R2440 vssa2.n196 vssa2.n195 0.046
R2441 vssa2.n189 vssa2.n188 0.046
R2442 vssa2.n270 vssa2.n269 0.046
R2443 vssa2.n215 vssa2.n214 0.046
R2444 vssa2.n424 vssa2.n321 0.045
R2445 vssa2.n425 vssa2.n315 0.045
R2446 vssa2 vssa2.n451 0.043
R2447 vssa2.n353 vssa2.n326 0.043
R2448 vssa2.n352 vssa2.n330 0.043
R2449 vssa2.n451 vssa2.n450 0.043
R2450 vssa2.n491 vssa2.n490 0.042
R2451 vssa2.n490 vssa2.n489 0.042
R2452 vssa2.n488 vssa2.n487 0.042
R2453 vssa2.n489 vssa2.n488 0.042
R2454 vssa2.n495 vssa2.n494 0.04
R2455 vssa2.n496 vssa2.n495 0.04
R2456 vssa2.n498 vssa2.n497 0.04
R2457 vssa2.n497 vssa2.n496 0.04
R2458 vssa2.n456 vssa2.n455 0.038
R2459 vssa2.n455 vssa2.n454 0.038
R2460 vssa2.n453 vssa2.n452 0.038
R2461 vssa2.n454 vssa2.n453 0.038
R2462 vssa2.n379 vssa2.n378 0.037
R2463 vssa2.n378 vssa2.n377 0.037
R2464 vssa2.n421 vssa2.n420 0.037
R2465 vssa2.n420 vssa2.n419 0.037
R2466 vssa2.n376 vssa2.n375 0.037
R2467 vssa2.n377 vssa2.n376 0.037
R2468 vssa2.n366 vssa2.n365 0.037
R2469 vssa2.n363 vssa2.n362 0.031
R2470 vssa2.n362 vssa2.n361 0.031
R2471 vssa2.n371 vssa2.n370 0.031
R2472 vssa2.n370 vssa2.n369 0.031
R2473 vssa2.n357 vssa2.n356 0.031
R2474 vssa2.n355 vssa2.n354 0.031
R2475 vssa2.n350 vssa2.n349 0.026
R2476 vssa2.n304 vssa2.n303 0.025
R2477 vssa2.n446 vssa2.n445 0.025
R2478 vssa2.n445 vssa2.n444 0.025
R2479 vssa2.n292 vssa2.n291 0.022
R2480 vssa2.n1 vssa2.n292 0.022
R2481 vssa2.n335 vssa2.n334 0.021
R2482 vssa2.n3 vssa2.n335 0.021
R2483 vssa2.n233 vssa2.n232 0.02
R2484 vssa2.n232 vssa2.n231 0.02
R2485 vssa2.n231 vssa2.n230 0.02
R2486 vssa2.n230 vssa2.n229 0.02
R2487 vssa2.n435 vssa2.n434 0.017
R2488 vssa2.n432 vssa2.n431 0.017
R2489 vssa2.n431 vssa2.n430 0.017
R2490 vssa2.n424 vssa2.n423 0.016
R2491 vssa2.n423 vssa2.n353 0.016
R2492 vssa2.n429 vssa2.n428 0.016
R2493 vssa2.n224 vssa2.n223 0.015
R2494 vssa2.n223 vssa2.n222 0.015
R2495 vssa2.n443 vssa2.n442 0.013
R2496 vssa2.n444 vssa2.n443 0.013
R2497 vssa2.n486 vssa2.n485 0.012
R2498 vssa2.n493 vssa2.n492 0.012
R2499 vssa2.n399 vssa2.n398 0.012
R2500 vssa2.n391 vssa2.n390 0.012
R2501 vssa2.n412 vssa2.n411 0.012
R2502 vssa2.n382 vssa2.n381 0.012
R2503 vssa2.n418 vssa2.n417 0.012
R2504 vssa2.n374 vssa2.n373 0.012
R2505 vssa2.n368 vssa2.n367 0.012
R2506 vssa2.n360 vssa2.n359 0.012
R2507 vssa2 vssa2.n8 0.012
R2508 vssa2.n348 vssa2.n347 0.011
R2509 vssa2.n3 vssa2.n348 0.011
R2510 vssa2.n333 vssa2.n332 0.011
R2511 vssa2.n308 vssa2.n307 0.011
R2512 vssa2.n306 vssa2.n305 0.011
R2513 vssa2.n2 vssa2.n306 0.011
R2514 vssa2.n13 vssa2.n12 0.011
R2515 vssa2.t128 vssa2.n13 0.011
R2516 vssa2.t128 vssa2.n11 0.011
R2517 vssa2.n11 vssa2.n10 0.011
R2518 vssa2.n3 vssa2.n333 0.011
R2519 vssa2.n2 vssa2.n308 0.011
R2520 vssa2.n1 vssa2.n290 0.011
R2521 vssa2 vssa2.n7 0.011
R2522 vssa2.n427 vssa2.n309 0.01
R2523 vssa2.n472 vssa2.n471 0.009
R2524 vssa2.t44 vssa2.n340 0.009
R2525 vssa2.t32 vssa2.n296 0.009
R2526 vssa2.n473 vssa2.n472 0.009
R2527 vssa2.n102 vssa2.n100 0.009
R2528 vssa2.n100 vssa2.t140 0.009
R2529 vssa2.n18 vssa2.n17 0.009
R2530 vssa2.t128 vssa2.n18 0.009
R2531 vssa2.n221 vssa2.n220 0.008
R2532 vssa2.n222 vssa2.n221 0.008
R2533 vssa2.n482 vssa2.n481 0.007
R2534 vssa2.n483 vssa2.n482 0.006
R2535 vssa2.n429 vssa2.n427 0.005
R2536 vssa2.n427 vssa2.n426 0.005
R2537 vssa2.n342 vssa2.n341 0.005
R2538 vssa2.t44 vssa2.n342 0.005
R2539 vssa2.n343 vssa2.t44 0.005
R2540 vssa2.n345 vssa2.n343 0.005
R2541 vssa2.n345 vssa2.n344 0.005
R2542 vssa2.n298 vssa2.n297 0.005
R2543 vssa2.t32 vssa2.n298 0.005
R2544 vssa2.n299 vssa2.t32 0.005
R2545 vssa2.n301 vssa2.n299 0.005
R2546 vssa2.n301 vssa2.n300 0.005
R2547 vssa2.n94 vssa2.n93 0.005
R2548 vssa2.t140 vssa2.n94 0.005
R2549 vssa2.n96 vssa2.n95 0.005
R2550 vssa2.t140 vssa2.n96 0.005
R2551 vssa2.t140 vssa2.n98 0.005
R2552 vssa2.n98 vssa2.n97 0.005
R2553 vssa2.n23 vssa2.n22 0.005
R2554 vssa2.n425 vssa2.n424 0.004
R2555 vssa2.n353 vssa2.n352 0.004
R2556 vssa2.n7 vssa2.n6 0.004
R2557 vssa2.n56 vssa2.n55 0.003
R2558 vssa2.t100 vssa2.n56 0.003
R2559 vssa2.n45 vssa2.n44 0.003
R2560 vssa2.t48 vssa2.n45 0.003
R2561 vssa2.n191 vssa2.n190 0.003
R2562 vssa2.n192 vssa2.n191 0.003
R2563 vssa2.n122 vssa2.n121 0.002
R2564 vssa2.n137 vssa2.n136 0.002
R2565 vssa2.n47 vssa2.n46 0.002
R2566 vssa2.n46 vssa2.t48 0.002
R2567 vssa2.n58 vssa2.n57 0.002
R2568 vssa2.n57 vssa2.t100 0.002
R2569 vssa2.n111 vssa2.n110 0.002
R2570 vssa2.t28 vssa2.n111 0.002
R2571 vssa2.n109 vssa2.n108 0.002
R2572 vssa2.n108 vssa2.t35 0.002
R2573 vssa2.n113 vssa2.n112 0.002
R2574 vssa2.n112 vssa2.t28 0.002
R2575 vssa2.t35 vssa2.n107 0.002
R2576 vssa2.n107 vssa2.n106 0.002
R2577 vssa2.n194 vssa2.n193 0.002
R2578 vssa2.n193 vssa2.n192 0.002
R2579 vssa2.n423 vssa2.n410 0.001
R2580 vssa2.n423 vssa2.n358 0.001
R2581 vssa2.n409 vssa2.t105 0.001
R2582 vssa2.t116 vssa2.n409 0.001
R2583 vssa2.n478 vssa2.n477 0.001
R2584 vssa2.n468 vssa2.n467 0.001
R2585 vssa2.n471 vssa2.n468 0.001
R2586 vssa2.n481 vssa2.n478 0.001
R2587 vssa2.n410 vssa2.t116 0.001
R2588 a_534722_685355.n0 a_534722_685355.t6 2.767
R2589 a_534722_685355.n5 a_534722_685355.t7 2.412
R2590 a_534722_685355.n0 a_534722_685355.t5 2.401
R2591 a_534722_685355.n1 a_534722_685355.n0 1.709
R2592 a_534722_685355.n5 a_534722_685355.n4 1.66
R2593 a_534722_685355.n2 a_534722_685355.n1 0.744
R2594 a_534722_685355.n3 a_534722_685355.n2 0.744
R2595 a_534722_685355.n4 a_534722_685355.n3 0.744
R2596 a_534722_685355.t4 a_534722_685355.n5 0.462
R2597 a_534722_685355.n4 a_534722_685355.t2 0.024
R2598 a_534722_685355.n3 a_534722_685355.t1 0.024
R2599 a_534722_685355.n2 a_534722_685355.t3 0.024
R2600 a_534722_685355.n1 a_534722_685355.t0 0.024
R2601 a_540916_680434.n9 a_540916_680434.t4 147.028
R2602 a_540916_680434.n6 a_540916_680434.t6 147.028
R2603 a_540916_680434.n37 a_540916_680434.t12 135.928
R2604 a_540916_680434.n33 a_540916_680434.t16 135.928
R2605 a_540916_680434.n30 a_540916_680434.t8 135.928
R2606 a_540916_680434.n27 a_540916_680434.t14 135.928
R2607 a_540916_680434.n20 a_540916_680434.t27 135.928
R2608 a_540916_680434.n3 a_540916_680434.t22 135.928
R2609 a_540916_680434.n15 a_540916_680434.t25 68.504
R2610 a_540916_680434.n21 a_540916_680434.t23 68.504
R2611 a_540916_680434.n38 a_540916_680434.t18 67.965
R2612 a_540916_680434.n23 a_540916_680434.t10 67.964
R2613 a_540916_680434.n2 a_540916_680434.t26 67.575
R2614 a_540916_680434.n1 a_540916_680434.t24 67.575
R2615 a_540916_680434.n19 a_540916_680434.n18 9.306
R2616 a_540916_680434.n8 a_540916_680434.t5 6.96
R2617 a_540916_680434.n5 a_540916_680434.t7 6.96
R2618 a_540916_680434.t19 a_540916_680434.n38 5.88
R2619 a_540916_680434.n23 a_540916_680434.t11 5.88
R2620 a_540916_680434.n25 a_540916_680434.t15 5.713
R2621 a_540916_680434.n29 a_540916_680434.t9 5.713
R2622 a_540916_680434.n32 a_540916_680434.t17 5.713
R2623 a_540916_680434.n36 a_540916_680434.t13 5.713
R2624 a_540916_680434.n10 a_540916_680434.t1 5.185
R2625 a_540916_680434.n17 a_540916_680434.t20 5.185
R2626 a_540916_680434.n10 a_540916_680434.t3 3.48
R2627 a_540916_680434.n12 a_540916_680434.t2 3.48
R2628 a_540916_680434.n11 a_540916_680434.t21 3.48
R2629 a_540916_680434.n17 a_540916_680434.t0 3.48
R2630 a_540916_680434.n2 a_540916_680434.n1 1.708
R2631 a_540916_680434.n12 a_540916_680434.n11 1.707
R2632 a_540916_680434.n13 a_540916_680434.n12 1.22
R2633 a_540916_680434.n16 a_540916_680434.n15 1.019
R2634 a_540916_680434.n22 a_540916_680434.n21 0.947
R2635 a_540916_680434.n3 a_540916_680434.n2 0.929
R2636 a_540916_680434.n22 a_540916_680434.n0 0.603
R2637 a_540916_680434.n14 a_540916_680434.n9 0.555
R2638 a_540916_680434.n16 a_540916_680434.n14 0.477
R2639 a_540916_680434.n25 a_540916_680434.n24 0.332
R2640 a_540916_680434.n29 a_540916_680434.n28 0.332
R2641 a_540916_680434.n30 a_540916_680434.n29 0.332
R2642 a_540916_680434.n32 a_540916_680434.n31 0.332
R2643 a_540916_680434.n33 a_540916_680434.n32 0.332
R2644 a_540916_680434.n37 a_540916_680434.n36 0.332
R2645 a_540916_680434.n22 a_540916_680434.n20 0.286
R2646 a_540916_680434.n16 a_540916_680434.n3 0.241
R2647 a_540916_680434.n24 a_540916_680434.n23 0.229
R2648 a_540916_680434.n38 a_540916_680434.n37 0.229
R2649 a_540916_680434.n35 a_540916_680434.n16 0.223
R2650 a_540916_680434.n5 a_540916_680434.n4 0.211
R2651 a_540916_680434.n6 a_540916_680434.n5 0.211
R2652 a_540916_680434.n8 a_540916_680434.n7 0.211
R2653 a_540916_680434.n9 a_540916_680434.n8 0.211
R2654 a_540916_680434.n26 a_540916_680434.n22 0.21
R2655 a_540916_680434.n13 a_540916_680434.n10 0.192
R2656 a_540916_680434.n14 a_540916_680434.n13 0.162
R2657 a_540916_680434.n0 a_540916_680434.n19 0.151
R2658 a_540916_680434.n0 a_540916_680434.n17 0.124
R2659 a_540916_680434.n27 a_540916_680434.n26 0.121
R2660 a_540916_680434.n35 a_540916_680434.n34 0.102
R2661 a_540916_680434.n36 a_540916_680434.n35 0.1
R2662 a_540916_680434.n7 a_540916_680434.n6 0.075
R2663 a_540916_680434.n26 a_540916_680434.n25 0.069
R2664 a_540916_680434.n28 a_540916_680434.n27 0.063
R2665 a_540916_680434.n31 a_540916_680434.n30 0.063
R2666 a_540916_680434.n34 a_540916_680434.n33 0.063
R2667 a_540371_681998.n4 a_540371_681998.t16 133.764
R2668 a_540371_681998.n45 a_540371_681998.t28 133.759
R2669 a_540371_681998.n43 a_540371_681998.t18 133.759
R2670 a_540371_681998.n60 a_540371_681998.t42 133.759
R2671 a_540371_681998.n55 a_540371_681998.t17 133.759
R2672 a_540371_681998.n57 a_540371_681998.t23 133.759
R2673 a_540371_681998.n46 a_540371_681998.t22 133.759
R2674 a_540371_681998.n28 a_540371_681998.t27 133.759
R2675 a_540371_681998.n30 a_540371_681998.t24 133.759
R2676 a_540371_681998.n39 a_540371_681998.t20 133.759
R2677 a_540371_681998.n10 a_540371_681998.t43 133.759
R2678 a_540371_681998.n11 a_540371_681998.t32 133.759
R2679 a_540371_681998.n12 a_540371_681998.t35 68.256
R2680 a_540371_681998.n21 a_540371_681998.t44 68.256
R2681 a_540371_681998.n26 a_540371_681998.t21 67.856
R2682 a_540371_681998.n53 a_540371_681998.t34 67.28
R2683 a_540371_681998.n51 a_540371_681998.t39 67.28
R2684 a_540371_681998.n36 a_540371_681998.t46 67.28
R2685 a_540371_681998.n58 a_540371_681998.t25 67.28
R2686 a_540371_681998.n41 a_540371_681998.t31 67.28
R2687 a_540371_681998.n50 a_540371_681998.t36 67.233
R2688 a_540371_681998.n32 a_540371_681998.t45 67.146
R2689 a_540371_681998.n33 a_540371_681998.t29 66.592
R2690 a_540371_681998.n47 a_540371_681998.t37 66.592
R2691 a_540371_681998.n44 a_540371_681998.t47 66.592
R2692 a_540371_681998.n56 a_540371_681998.t30 66.592
R2693 a_540371_681998.n61 a_540371_681998.t38 66.592
R2694 a_540371_681998.n29 a_540371_681998.t41 66.592
R2695 a_540371_681998.n26 a_540371_681998.t40 66.592
R2696 a_540371_681998.n40 a_540371_681998.t33 66.592
R2697 a_540371_681998.n12 a_540371_681998.t19 66.475
R2698 a_540371_681998.n21 a_540371_681998.t26 66.475
R2699 a_540371_681998.n5 a_540371_681998.t12 43.389
R2700 a_540371_681998.n1 a_540371_681998.t14 43.388
R2701 a_540371_681998.n0 a_540371_681998.t8 43.387
R2702 a_540371_681998.n0 a_540371_681998.t10 43.387
R2703 a_540371_681998.n7 a_540371_681998.t13 13.925
R2704 a_540371_681998.n20 a_540371_681998.t15 13.923
R2705 a_540371_681998.n17 a_540371_681998.t11 13.923
R2706 a_540371_681998.n6 a_540371_681998.t9 13.922
R2707 a_540371_681998.n2 a_540371_681998.n66 9.37
R2708 a_540371_681998.n9 a_540371_681998.n8 9.3
R2709 a_540371_681998.n65 a_540371_681998.t2 7.331
R2710 a_540371_681998.n18 a_540371_681998.t4 7.331
R2711 a_540371_681998.n15 a_540371_681998.t6 6.96
R2712 a_540371_681998.n24 a_540371_681998.t7 6.96
R2713 a_540371_681998.n64 a_540371_681998.t1 5.713
R2714 a_540371_681998.n19 a_540371_681998.t3 5.713
R2715 a_540371_681998.n18 a_540371_681998.t0 5.713
R2716 a_540371_681998.t5 a_540371_681998.n65 5.713
R2717 a_540371_681998.n19 a_540371_681998.n18 1.617
R2718 a_540371_681998.n65 a_540371_681998.n64 1.616
R2719 a_540371_681998.n22 a_540371_681998.n21 0.97
R2720 a_540371_681998.n13 a_540371_681998.n12 0.97
R2721 a_540371_681998.n35 a_540371_681998.n31 0.968
R2722 a_540371_681998.n38 a_540371_681998.n37 0.968
R2723 a_540371_681998.n23 a_540371_681998.n22 0.939
R2724 a_540371_681998.n14 a_540371_681998.n13 0.939
R2725 a_540371_681998.n5 a_540371_681998.n63 0.688
R2726 a_540371_681998.n34 a_540371_681998.n33 0.688
R2727 a_540371_681998.n47 a_540371_681998.n46 0.688
R2728 a_540371_681998.n45 a_540371_681998.n44 0.688
R2729 a_540371_681998.n56 a_540371_681998.n55 0.688
R2730 a_540371_681998.n62 a_540371_681998.n61 0.688
R2731 a_540371_681998.n61 a_540371_681998.n60 0.688
R2732 a_540371_681998.n57 a_540371_681998.n56 0.688
R2733 a_540371_681998.n44 a_540371_681998.n43 0.688
R2734 a_540371_681998.n48 a_540371_681998.n47 0.688
R2735 a_540371_681998.n29 a_540371_681998.n28 0.688
R2736 a_540371_681998.n27 a_540371_681998.n26 0.688
R2737 a_540371_681998.n30 a_540371_681998.n29 0.688
R2738 a_540371_681998.n40 a_540371_681998.n39 0.688
R2739 a_540371_681998.n4 a_540371_681998.n40 0.674
R2740 a_540371_681998.n33 a_540371_681998.n32 0.667
R2741 a_540371_681998.n37 a_540371_681998.n36 0.601
R2742 a_540371_681998.n31 a_540371_681998.n27 0.582
R2743 a_540371_681998.n35 a_540371_681998.n34 0.582
R2744 a_540371_681998.n31 a_540371_681998.n30 0.573
R2745 a_540371_681998.n49 a_540371_681998.n48 0.568
R2746 a_540371_681998.n60 a_540371_681998.n59 0.562
R2747 a_540371_681998.n43 a_540371_681998.n42 0.562
R2748 a_540371_681998.n39 a_540371_681998.n38 0.555
R2749 a_540371_681998.n54 a_540371_681998.n53 0.554
R2750 a_540371_681998.n52 a_540371_681998.n51 0.554
R2751 a_540371_681998.n14 a_540371_681998.n11 0.53
R2752 a_540371_681998.n55 a_540371_681998.n54 0.477
R2753 a_540371_681998.n59 a_540371_681998.n58 0.468
R2754 a_540371_681998.n42 a_540371_681998.n41 0.468
R2755 a_540371_681998.n4 a_540371_681998.n35 0.464
R2756 a_540371_681998.n63 a_540371_681998.n62 0.462
R2757 a_540371_681998.n49 a_540371_681998.n45 0.462
R2758 a_540371_681998.n1 a_540371_681998.n25 0.431
R2759 a_540371_681998.n0 a_540371_681998.n16 0.424
R2760 a_540371_681998.n63 a_540371_681998.n57 0.422
R2761 a_540371_681998.n49 a_540371_681998.n4 0.363
R2762 a_540371_681998.n52 a_540371_681998.n50 0.357
R2763 a_540371_681998.n54 a_540371_681998.n52 0.357
R2764 a_540371_681998.n63 a_540371_681998.n49 0.33
R2765 a_540371_681998.n3 a_540371_681998.n0 0.327
R2766 a_540371_681998.n1 a_540371_681998.n2 0.319
R2767 a_540371_681998.n16 a_540371_681998.n14 0.251
R2768 a_540371_681998.n25 a_540371_681998.n23 0.251
R2769 a_540371_681998.n11 a_540371_681998.n10 0.158
R2770 a_540371_681998.n2 a_540371_681998.n19 0.118
R2771 a_540371_681998.n0 a_540371_681998.n17 0.116
R2772 a_540371_681998.n64 a_540371_681998.n3 0.104
R2773 a_540371_681998.n1 a_540371_681998.n20 0.102
R2774 a_540371_681998.n7 a_540371_681998.n1 0.098
R2775 a_540371_681998.n0 a_540371_681998.n6 0.083
R2776 a_540371_681998.n3 a_540371_681998.n9 0.082
R2777 a_540371_681998.n25 a_540371_681998.n24 0.069
R2778 a_540371_681998.n16 a_540371_681998.n15 0.067
R2779 a_540371_681998.n5 a_540371_681998.n7 0.051
R2780 a_540371_681998.n6 a_540371_681998.n5 0.041
R2781 constant_gm_fingers_0/Vout.n37 constant_gm_fingers_0/Vout.t17 133.759
R2782 constant_gm_fingers_0/Vout.n52 constant_gm_fingers_0/Vout.t22 133.759
R2783 constant_gm_fingers_0/Vout.n74 constant_gm_fingers_0/Vout.t26 133.759
R2784 constant_gm_fingers_0/Vout.n73 constant_gm_fingers_0/Vout.t20 133.759
R2785 constant_gm_fingers_0/Vout.n72 constant_gm_fingers_0/Vout.t45 133.759
R2786 constant_gm_fingers_0/Vout.n71 constant_gm_fingers_0/Vout.t43 133.759
R2787 constant_gm_fingers_0/Vout.n70 constant_gm_fingers_0/Vout.t37 133.759
R2788 constant_gm_fingers_0/Vout.n13 constant_gm_fingers_0/Vout.t35 133.759
R2789 constant_gm_fingers_0/Vout.n14 constant_gm_fingers_0/Vout.t27 133.759
R2790 constant_gm_fingers_0/Vout.n15 constant_gm_fingers_0/Vout.t34 133.759
R2791 constant_gm_fingers_0/Vout.n16 constant_gm_fingers_0/Vout.t19 133.759
R2792 constant_gm_fingers_0/Vout.n17 constant_gm_fingers_0/Vout.t44 133.759
R2793 constant_gm_fingers_0/Vout.n18 constant_gm_fingers_0/Vout.t40 133.759
R2794 constant_gm_fingers_0/Vout.n75 constant_gm_fingers_0/Vout.t30 133.759
R2795 constant_gm_fingers_0/Vout.n63 constant_gm_fingers_0/Vout.t42 133.759
R2796 constant_gm_fingers_0/Vout.n62 constant_gm_fingers_0/Vout.t18 133.759
R2797 constant_gm_fingers_0/Vout.n61 constant_gm_fingers_0/Vout.t15 133.759
R2798 constant_gm_fingers_0/Vout.n60 constant_gm_fingers_0/Vout.t38 133.759
R2799 constant_gm_fingers_0/Vout.n59 constant_gm_fingers_0/Vout.t23 133.759
R2800 constant_gm_fingers_0/Vout.n58 constant_gm_fingers_0/Vout.t32 133.759
R2801 constant_gm_fingers_0/Vout.n57 constant_gm_fingers_0/Vout.t25 133.759
R2802 constant_gm_fingers_0/Vout.n26 constant_gm_fingers_0/Vout.t24 133.759
R2803 constant_gm_fingers_0/Vout.n27 constant_gm_fingers_0/Vout.t16 133.759
R2804 constant_gm_fingers_0/Vout.n28 constant_gm_fingers_0/Vout.t14 133.759
R2805 constant_gm_fingers_0/Vout.n29 constant_gm_fingers_0/Vout.t39 133.759
R2806 constant_gm_fingers_0/Vout.n30 constant_gm_fingers_0/Vout.t33 133.759
R2807 constant_gm_fingers_0/Vout.n31 constant_gm_fingers_0/Vout.t29 133.759
R2808 constant_gm_fingers_0/Vout.n32 constant_gm_fingers_0/Vout.t36 133.759
R2809 constant_gm_fingers_0/Vout.n2 constant_gm_fingers_0/Vout.t41 133.758
R2810 constant_gm_fingers_0/Vout.n3 constant_gm_fingers_0/Vout.t28 133.758
R2811 constant_gm_fingers_0/Vout.n36 constant_gm_fingers_0/Vout.t21 66.052
R2812 constant_gm_fingers_0/Vout.n51 constant_gm_fingers_0/Vout.t31 66.049
R2813 constant_gm_fingers_0/Vout.n56 constant_gm_fingers_0/Vout.t4 43.387
R2814 constant_gm_fingers_0/Vout.n47 constant_gm_fingers_0/Vout.t6 43.384
R2815 constant_gm_fingers_0/Vout.n41 constant_gm_fingers_0/Vout.t8 43.384
R2816 constant_gm_fingers_0/Vout.n43 constant_gm_fingers_0/Vout.t10 43.384
R2817 constant_gm_fingers_0/Vout.n4 constant_gm_fingers_0/Vout.t7 13.92
R2818 constant_gm_fingers_0/Vout.n4 constant_gm_fingers_0/Vout.t5 13.92
R2819 constant_gm_fingers_0/Vout.n5 constant_gm_fingers_0/Vout.t11 13.92
R2820 constant_gm_fingers_0/Vout.n5 constant_gm_fingers_0/Vout.t9 13.92
R2821 constant_gm_fingers_0/Vout.n45 constant_gm_fingers_0/Vout.t12 6.96
R2822 constant_gm_fingers_0/Vout.n45 constant_gm_fingers_0/Vout.t13 6.96
R2823 constant_gm_fingers_0/Vout.n6 constant_gm_fingers_0/Vout.t0 5.713
R2824 constant_gm_fingers_0/Vout.n6 constant_gm_fingers_0/Vout.t2 5.713
R2825 constant_gm_fingers_0/Vout.n44 constant_gm_fingers_0/Vout.n43 4.431
R2826 constant_gm_fingers_0/Vout.t1 constant_gm_fingers_0/Vout.n56 4.348
R2827 constant_gm_fingers_0/Vout.n51 constant_gm_fingers_0/Vout.n50 2.308
R2828 constant_gm_fingers_0/Vout.n36 constant_gm_fingers_0/Vout.n35 2.303
R2829 constant_gm_fingers_0/Vout.n3 constant_gm_fingers_0/Vout.n51 2.28
R2830 constant_gm_fingers_0/Vout.n2 constant_gm_fingers_0/Vout.n36 2.276
R2831 constant_gm_fingers_0/Vout.n0 constant_gm_fingers_0/Vout.n69 1.934
R2832 constant_gm_fingers_0/Vout.n1 constant_gm_fingers_0/Vout.n12 1.859
R2833 constant_gm_fingers_0/Vout.n0 constant_gm_fingers_0/Vout.n75 1.588
R2834 constant_gm_fingers_0/Vout.n1 constant_gm_fingers_0/Vout.n18 1.513
R2835 constant_gm_fingers_0/Vout.t1 constant_gm_fingers_0/Vout.n83 1.146
R2836 constant_gm_fingers_0/Vout.n44 constant_gm_fingers_0/Vout.n33 1.138
R2837 constant_gm_fingers_0/Vout.n46 constant_gm_fingers_0/Vout.n45 1.054
R2838 constant_gm_fingers_0/Vout.n0 constant_gm_fingers_0/Vout.n82 0.938
R2839 constant_gm_fingers_0/Vout.n83 constant_gm_fingers_0/Vout.n63 0.938
R2840 constant_gm_fingers_0/Vout.n1 constant_gm_fingers_0/Vout.n25 0.873
R2841 constant_gm_fingers_0/Vout.n33 constant_gm_fingers_0/Vout.n32 0.873
R2842 constant_gm_fingers_0/Vout.n35 constant_gm_fingers_0/Vout.n34 0.645
R2843 constant_gm_fingers_0/Vout.n50 constant_gm_fingers_0/Vout.n49 0.645
R2844 constant_gm_fingers_0/Vout.n18 constant_gm_fingers_0/Vout.n17 0.645
R2845 constant_gm_fingers_0/Vout.n17 constant_gm_fingers_0/Vout.n16 0.645
R2846 constant_gm_fingers_0/Vout.n16 constant_gm_fingers_0/Vout.n15 0.645
R2847 constant_gm_fingers_0/Vout.n15 constant_gm_fingers_0/Vout.n14 0.645
R2848 constant_gm_fingers_0/Vout.n14 constant_gm_fingers_0/Vout.n13 0.645
R2849 constant_gm_fingers_0/Vout.n71 constant_gm_fingers_0/Vout.n70 0.645
R2850 constant_gm_fingers_0/Vout.n72 constant_gm_fingers_0/Vout.n71 0.645
R2851 constant_gm_fingers_0/Vout.n73 constant_gm_fingers_0/Vout.n72 0.645
R2852 constant_gm_fingers_0/Vout.n74 constant_gm_fingers_0/Vout.n73 0.645
R2853 constant_gm_fingers_0/Vout.n75 constant_gm_fingers_0/Vout.n74 0.645
R2854 constant_gm_fingers_0/Vout.n25 constant_gm_fingers_0/Vout.n24 0.645
R2855 constant_gm_fingers_0/Vout.n24 constant_gm_fingers_0/Vout.n23 0.645
R2856 constant_gm_fingers_0/Vout.n23 constant_gm_fingers_0/Vout.n22 0.645
R2857 constant_gm_fingers_0/Vout.n22 constant_gm_fingers_0/Vout.n21 0.645
R2858 constant_gm_fingers_0/Vout.n21 constant_gm_fingers_0/Vout.n20 0.645
R2859 constant_gm_fingers_0/Vout.n20 constant_gm_fingers_0/Vout.n19 0.645
R2860 constant_gm_fingers_0/Vout.n77 constant_gm_fingers_0/Vout.n76 0.645
R2861 constant_gm_fingers_0/Vout.n78 constant_gm_fingers_0/Vout.n77 0.645
R2862 constant_gm_fingers_0/Vout.n79 constant_gm_fingers_0/Vout.n78 0.645
R2863 constant_gm_fingers_0/Vout.n80 constant_gm_fingers_0/Vout.n79 0.645
R2864 constant_gm_fingers_0/Vout.n81 constant_gm_fingers_0/Vout.n80 0.645
R2865 constant_gm_fingers_0/Vout.n82 constant_gm_fingers_0/Vout.n81 0.645
R2866 constant_gm_fingers_0/Vout.n32 constant_gm_fingers_0/Vout.n31 0.645
R2867 constant_gm_fingers_0/Vout.n31 constant_gm_fingers_0/Vout.n30 0.645
R2868 constant_gm_fingers_0/Vout.n30 constant_gm_fingers_0/Vout.n29 0.645
R2869 constant_gm_fingers_0/Vout.n29 constant_gm_fingers_0/Vout.n28 0.645
R2870 constant_gm_fingers_0/Vout.n28 constant_gm_fingers_0/Vout.n27 0.645
R2871 constant_gm_fingers_0/Vout.n27 constant_gm_fingers_0/Vout.n26 0.645
R2872 constant_gm_fingers_0/Vout.n58 constant_gm_fingers_0/Vout.n57 0.645
R2873 constant_gm_fingers_0/Vout.n59 constant_gm_fingers_0/Vout.n58 0.645
R2874 constant_gm_fingers_0/Vout.n60 constant_gm_fingers_0/Vout.n59 0.645
R2875 constant_gm_fingers_0/Vout.n61 constant_gm_fingers_0/Vout.n60 0.645
R2876 constant_gm_fingers_0/Vout.n62 constant_gm_fingers_0/Vout.n61 0.645
R2877 constant_gm_fingers_0/Vout.n63 constant_gm_fingers_0/Vout.n62 0.645
R2878 constant_gm_fingers_0/Vout.n12 constant_gm_fingers_0/Vout.n11 0.645
R2879 constant_gm_fingers_0/Vout.n11 constant_gm_fingers_0/Vout.n10 0.645
R2880 constant_gm_fingers_0/Vout.n10 constant_gm_fingers_0/Vout.n9 0.645
R2881 constant_gm_fingers_0/Vout.n9 constant_gm_fingers_0/Vout.n8 0.645
R2882 constant_gm_fingers_0/Vout.n8 constant_gm_fingers_0/Vout.n7 0.645
R2883 constant_gm_fingers_0/Vout.n65 constant_gm_fingers_0/Vout.n64 0.645
R2884 constant_gm_fingers_0/Vout.n66 constant_gm_fingers_0/Vout.n65 0.645
R2885 constant_gm_fingers_0/Vout.n67 constant_gm_fingers_0/Vout.n66 0.645
R2886 constant_gm_fingers_0/Vout.n68 constant_gm_fingers_0/Vout.n67 0.645
R2887 constant_gm_fingers_0/Vout.n69 constant_gm_fingers_0/Vout.n68 0.645
R2888 constant_gm_fingers_0/Vout.n3 constant_gm_fingers_0/Vout.n52 0.599
R2889 constant_gm_fingers_0/Vout.n2 constant_gm_fingers_0/Vout.n37 0.594
R2890 constant_gm_fingers_0/Vout.n44 constant_gm_fingers_0/Vout.n6 0.587
R2891 constant_gm_fingers_0/Vout.n38 constant_gm_fingers_0/Vout.n2 0.586
R2892 constant_gm_fingers_0/Vout.n53 constant_gm_fingers_0/Vout.n3 0.583
R2893 constant_gm_fingers_0/Vout.n33 constant_gm_fingers_0/Vout.n1 0.474
R2894 constant_gm_fingers_0/Vout.n83 constant_gm_fingers_0/Vout.n0 0.474
R2895 constant_gm_fingers_0/Vout.n55 constant_gm_fingers_0/Vout.n4 0.415
R2896 constant_gm_fingers_0/Vout.n42 constant_gm_fingers_0/Vout.n5 0.414
R2897 constant_gm_fingers_0/Vout.n5 constant_gm_fingers_0/Vout.n40 0.414
R2898 constant_gm_fingers_0/Vout.n4 constant_gm_fingers_0/Vout.n54 0.412
R2899 constant_gm_fingers_0/Vout.n42 constant_gm_fingers_0/Vout.n41 0.332
R2900 constant_gm_fingers_0/Vout.n40 constant_gm_fingers_0/Vout.n39 0.332
R2901 constant_gm_fingers_0/Vout.n56 constant_gm_fingers_0/Vout.n55 0.323
R2902 constant_gm_fingers_0/Vout.n55 constant_gm_fingers_0/Vout.n47 0.322
R2903 constant_gm_fingers_0/Vout.n54 constant_gm_fingers_0/Vout.n48 0.322
R2904 constant_gm_fingers_0/Vout.n43 constant_gm_fingers_0/Vout.n42 0.312
R2905 constant_gm_fingers_0/Vout.n54 constant_gm_fingers_0/Vout.n53 0.283
R2906 constant_gm_fingers_0/Vout.n40 constant_gm_fingers_0/Vout.n38 0.283
R2907 constant_gm_fingers_0/Vout.n47 constant_gm_fingers_0/Vout.n46 0.277
R2908 constant_gm_fingers_0/Vout.t1 constant_gm_fingers_0/Vout.t3 0.203
R2909 constant_gm_fingers_0/Vout.t3 constant_gm_fingers_0/Vout.n44 0.203
R2910 io_analog[2].n33 io_analog[2].n32 21.976
R2911 io_analog[2].n37 io_analog[2].n36 17.091
R2912 io_analog[2].n67 io_analog[2].t14 7.884
R2913 io_analog[2].n20 io_analog[2].t0 7.884
R2914 io_analog[2].n68 io_analog[2].t3 7.884
R2915 io_analog[2].n65 io_analog[2].t18 7.88
R2916 io_analog[2].n25 io_analog[2].t44 6.315
R2917 io_analog[2].n80 io_analog[2].t4 5.78
R2918 io_analog[2].n53 io_analog[2].t17 5.779
R2919 io_analog[2].n41 io_analog[2].t13 5.779
R2920 io_analog[2].n1 io_analog[2].t1 5.779
R2921 io_analog[2].n63 io_analog[2].t32 5.778
R2922 io_analog[2].n70 io_analog[2].t20 5.775
R2923 io_analog[2].n17 io_analog[2].t16 5.774
R2924 io_analog[2].n67 io_analog[2].t2 5.769
R2925 io_analog[2].n20 io_analog[2].t36 5.769
R2926 io_analog[2].n68 io_analog[2].t37 5.769
R2927 io_analog[2].n5 io_analog[2].t30 5.769
R2928 io_analog[2].n65 io_analog[2].t6 5.767
R2929 io_analog[2].n69 io_analog[2].t9 5.713
R2930 io_analog[2].n71 io_analog[2].t7 5.713
R2931 io_analog[2].n73 io_analog[2].t26 5.713
R2932 io_analog[2].n75 io_analog[2].t11 5.713
R2933 io_analog[2].n77 io_analog[2].t33 5.713
R2934 io_analog[2].n79 io_analog[2].t15 5.713
R2935 io_analog[2].n8 io_analog[2].t12 5.713
R2936 io_analog[2].n10 io_analog[2].t31 5.713
R2937 io_analog[2].n12 io_analog[2].t10 5.713
R2938 io_analog[2].n14 io_analog[2].t23 5.713
R2939 io_analog[2].n16 io_analog[2].t5 5.713
R2940 io_analog[2].n23 io_analog[2].t39 5.713
R2941 io_analog[2].n54 io_analog[2].t29 5.713
R2942 io_analog[2].n58 io_analog[2].t27 5.713
R2943 io_analog[2].n60 io_analog[2].t35 5.713
R2944 io_analog[2].n62 io_analog[2].t21 5.713
R2945 io_analog[2].n64 io_analog[2].t24 5.713
R2946 io_analog[2].n44 io_analog[2].t38 5.713
R2947 io_analog[2].n42 io_analog[2].t28 5.713
R2948 io_analog[2].n50 io_analog[2].t25 5.713
R2949 io_analog[2].n48 io_analog[2].t34 5.713
R2950 io_analog[2].n46 io_analog[2].t19 5.713
R2951 io_analog[2].n66 io_analog[2].t22 5.713
R2952 io_analog[2].n19 io_analog[2].t8 5.713
R2953 io_analog[2].n40 io_analog[2].t40 3.531
R2954 io_analog[2].n30 io_analog[2].t41 3.481
R2955 io_analog[2].n29 io_analog[2].t46 3.48
R2956 io_analog[2].n28 io_analog[2].t51 3.48
R2957 io_analog[2].n37 io_analog[2].t42 3.48
R2958 io_analog[2].n39 io_analog[2].t47 3.48
R2959 io_analog[2].n35 io_analog[2].t48 3.48
R2960 io_analog[2].n33 io_analog[2].t43 3.48
R2961 io_analog[2].n26 io_analog[2].t45 3.48
R2962 io_analog[2].n25 io_analog[2].t50 3.48
R2963 io_analog[2].n31 io_analog[2].t49 3.48
R2964 io_analog[2].n29 io_analog[2].n28 2.835
R2965 io_analog[2].n35 io_analog[2].n34 2.831
R2966 io_analog[2].n39 io_analog[2].n38 2.821
R2967 io_analog[2].n26 io_analog[2].n25 2.819
R2968 io_analog[2].n30 io_analog[2].n29 2.815
R2969 io_analog[2].n28 io_analog[2].n27 2.722
R2970 io_analog[2].n36 io_analog[2].n35 2.701
R2971 io_analog[2].n32 io_analog[2].n31 2.396
R2972 io_analog[2].n40 io_analog[2].n39 2.375
R2973 io_analog[2].n8 io_analog[2].n1 2.213
R2974 io_analog[2].n42 io_analog[2].n41 2.213
R2975 io_analog[2].n54 io_analog[2].n53 2.213
R2976 io_analog[2].n80 io_analog[2].n79 2.212
R2977 io_analog[2].n75 io_analog[2].n74 2.21
R2978 io_analog[2].n59 io_analog[2].n58 2.209
R2979 io_analog[2].n50 io_analog[2].n49 2.209
R2980 io_analog[2].n13 io_analog[2].n12 2.209
R2981 io_analog[2].n46 io_analog[2].n5 2.203
R2982 io_analog[2].n67 io_analog[2].n66 2.2
R2983 io_analog[2].n20 io_analog[2].n19 2.2
R2984 io_analog[2].n69 io_analog[2].n68 2.2
R2985 io_analog[2].n65 io_analog[2].n64 2.196
R2986 io_analog[2].n63 io_analog[2].n62 2.185
R2987 io_analog[2].n17 io_analog[2].n16 2.185
R2988 io_analog[2].n71 io_analog[2].n70 2.185
R2989 io_analog[2].n12 io_analog[2].n11 2.181
R2990 io_analog[2].n76 io_analog[2].n75 2.18
R2991 io_analog[2].n66 io_analog[2].n5 2.167
R2992 io_analog[2].n19 io_analog[2].n17 2.167
R2993 io_analog[2].n70 io_analog[2].n69 2.167
R2994 io_analog[2].n51 io_analog[2].n50 2.162
R2995 io_analog[2].n58 io_analog[2].n57 2.16
R2996 io_analog[2].n64 io_analog[2].n63 2.15
R2997 io_analog[2].n47 io_analog[2].n46 2.149
R2998 io_analog[2].n16 io_analog[2].n15 2.149
R2999 io_analog[2].n62 io_analog[2].n61 2.131
R3000 io_analog[2].n72 io_analog[2].n71 2.13
R3001 io_analog[2].n79 io_analog[2].n78 2.107
R3002 io_analog[2].n9 io_analog[2].n8 2.106
R3003 io_analog[2].n43 io_analog[2].n42 2.088
R3004 io_analog[2].n55 io_analog[2].n54 2.085
R3005 io_analog[2] io_analog[2].n83 1.8
R3006 io_analog[2].n20 io_analog[2].n18 1.418
R3007 io_analog[2].n31 io_analog[2].n30 1.027
R3008 io_analog[2].n83 io_analog[2].n0 1.022
R3009 io_analog[2].n27 io_analog[2].n24 0.957
R3010 io_analog[2].n57 io_analog[2].n40 0.917
R3011 io_analog[2].n63 io_analog[2].n21 0.851
R3012 io_analog[2].n24 io_analog[2].n22 0.665
R3013 io_analog[2].n83 io_analog[2].n82 0.314
R3014 io_analog[2].n67 io_analog[2].n65 0.237
R3015 io_analog[2].n53 io_analog[2].n2 0.233
R3016 io_analog[2].n70 io_analog[2].n17 0.232
R3017 io_analog[2].n70 io_analog[2].n5 0.232
R3018 io_analog[2].n68 io_analog[2].n20 0.232
R3019 io_analog[2].n68 io_analog[2].n67 0.232
R3020 io_analog[2].n45 io_analog[2].n22 0.232
R3021 io_analog[2].n82 io_analog[2].n81 0.232
R3022 io_analog[2].n81 io_analog[2].n2 0.232
R3023 io_analog[2].n45 io_analog[2].n4 0.231
R3024 io_analog[2].n6 io_analog[2].n4 0.231
R3025 io_analog[2].n63 io_analog[2].n5 0.23
R3026 io_analog[2].n44 io_analog[2].n43 0.22
R3027 io_analog[2].n55 io_analog[2].n23 0.214
R3028 io_analog[2].n52 io_analog[2].n3 0.21
R3029 io_analog[2].n7 io_analog[2].n3 0.209
R3030 io_analog[2].n10 io_analog[2].n9 0.202
R3031 io_analog[2].n78 io_analog[2].n77 0.201
R3032 io_analog[2].n73 io_analog[2].n72 0.177
R3033 io_analog[2].n61 io_analog[2].n60 0.176
R3034 io_analog[2].n56 io_analog[2].n52 0.166
R3035 io_analog[2].n15 io_analog[2].n14 0.158
R3036 io_analog[2].n48 io_analog[2].n47 0.158
R3037 io_analog[2].n51 io_analog[2].n44 0.144
R3038 io_analog[2].n57 io_analog[2].n23 0.139
R3039 io_analog[2].t53 io_analog[2].t55 0.134
R3040 io_analog[2].n77 io_analog[2].n76 0.126
R3041 io_analog[2].n11 io_analog[2].n10 0.125
R3042 io_analog[2].n60 io_analog[2].n59 0.098
R3043 io_analog[2].n49 io_analog[2].n48 0.098
R3044 io_analog[2].n14 io_analog[2].n13 0.098
R3045 io_analog[2].n74 io_analog[2].n73 0.097
R3046 io_analog[2].t55 io_analog[2].n0 0.071
R3047 io_analog[2].n18 io_analog[2].t54 0.067
R3048 io_analog[2].n18 io_analog[2].t53 0.067
R3049 io_analog[2].n0 io_analog[2].t52 0.062
R3050 io_analog[2].n57 io_analog[2].n56 0.057
R3051 io_analog[2].n56 io_analog[2].n55 0.057
R3052 io_analog[2].n34 io_analog[2].n21 0.051
R3053 io_analog[2].n27 io_analog[2].n26 0.049
R3054 io_analog[2].n38 io_analog[2].n24 0.049
R3055 io_analog[2].n36 io_analog[2].n24 0.021
R3056 io_analog[2].n9 io_analog[2].n7 0.002
R3057 io_analog[2].n13 io_analog[2].n6 0.002
R3058 io_analog[2].n32 io_analog[2].n21 0.001
R3059 io_analog[2].n82 io_analog[2].n1 0.001
R3060 io_analog[2].n41 io_analog[2].n2 0.001
R3061 io_analog[2].n52 io_analog[2].n43 0.001
R3062 io_analog[2].n78 io_analog[2].n3 0.001
R3063 io_analog[2].n72 io_analog[2].n4 0.001
R3064 io_analog[2].n61 io_analog[2].n22 0.001
R3065 io_analog[2].n52 io_analog[2].n51 0.001
R3066 io_analog[2].n47 io_analog[2].n45 0.001
R3067 io_analog[2].n15 io_analog[2].n6 0.001
R3068 io_analog[2].n76 io_analog[2].n3 0.001
R3069 io_analog[2].n11 io_analog[2].n7 0.001
R3070 io_analog[2].n59 io_analog[2].n22 0.001
R3071 io_analog[2].n49 io_analog[2].n45 0.001
R3072 io_analog[2].n74 io_analog[2].n4 0.001
R3073 io_analog[2].n81 io_analog[2].n80 0.001
R3074 io_analog[2].n38 io_analog[2].n37 0.001
R3075 io_analog[2].n34 io_analog[2].n33 0.001
R3076 io_analog[8].n7 io_analog[8].t2 267.528
R3077 io_analog[8].n8 io_analog[8].t0 267.528
R3078 io_analog[8].n6 io_analog[8].t5 267.528
R3079 io_analog[8].n5 io_analog[8].t1 267.528
R3080 io_analog[8].n4 io_analog[8].t4 267.528
R3081 io_analog[8].n3 io_analog[8].t6 267.528
R3082 io_analog[8].n0 io_analog[8].t3 133.051
R3083 io_analog[8] io_analog[8].n13 2.289
R3084 io_analog[8].n1 io_analog[8].n0 1.822
R3085 io_analog[8].n13 io_analog[8].n12 1.288
R3086 io_analog[8].n13 io_analog[8].n6 1.288
R3087 io_analog[8].n12 io_analog[8].n11 0.395
R3088 io_analog[8].n11 io_analog[8].n10 0.395
R3089 io_analog[8].n10 io_analog[8].n9 0.395
R3090 io_analog[8].n9 io_analog[8].n8 0.395
R3091 io_analog[8].n8 io_analog[8].n7 0.395
R3092 io_analog[8].n6 io_analog[8].n5 0.395
R3093 io_analog[8].n5 io_analog[8].n4 0.395
R3094 io_analog[8].n4 io_analog[8].n3 0.395
R3095 io_analog[8].n3 io_analog[8].n2 0.395
R3096 io_analog[8].n2 io_analog[8].n1 0.395
R3097 a_37693_693523.n0 a_37693_693523.t1 2.62
R3098 a_37693_693523.n0 a_37693_693523.t2 2.618
R3099 a_37693_693523.n5 a_37693_693523.t7 2.609
R3100 a_37693_693523.n5 a_37693_693523.n4 2.124
R3101 a_37693_693523.n1 a_37693_693523.n0 2.12
R3102 a_37693_693523.n4 a_37693_693523.n3 0.744
R3103 a_37693_693523.n3 a_37693_693523.n2 0.744
R3104 a_37693_693523.n2 a_37693_693523.n1 0.744
R3105 a_37693_693523.t0 a_37693_693523.n5 0.295
R3106 a_37693_693523.n1 a_37693_693523.t6 0.024
R3107 a_37693_693523.n2 a_37693_693523.t3 0.024
R3108 a_37693_693523.n3 a_37693_693523.t5 0.024
R3109 a_37693_693523.n4 a_37693_693523.t4 0.024
R3110 a_540459_681940.n32 a_540459_681940.t11 6.281
R3111 a_540459_681940.n22 a_540459_681940.t2 6.193
R3112 a_540459_681940.n15 a_540459_681940.t23 5.945
R3113 a_540459_681940.n36 a_540459_681940.t20 5.945
R3114 a_540459_681940.n6 a_540459_681940.n34 4.5
R3115 a_540459_681940.n5 a_540459_681940.n21 4.5
R3116 a_540459_681940.n2 a_540459_681940.t4 3.502
R3117 a_540459_681940.n14 a_540459_681940.t14 3.48
R3118 a_540459_681940.n13 a_540459_681940.t22 3.48
R3119 a_540459_681940.n12 a_540459_681940.t18 3.48
R3120 a_540459_681940.n11 a_540459_681940.t25 3.48
R3121 a_540459_681940.n24 a_540459_681940.t13 3.48
R3122 a_540459_681940.n25 a_540459_681940.t3 3.48
R3123 a_540459_681940.n26 a_540459_681940.t6 3.48
R3124 a_540459_681940.n20 a_540459_681940.t17 3.48
R3125 a_540459_681940.n19 a_540459_681940.t24 3.48
R3126 a_540459_681940.n18 a_540459_681940.t21 3.48
R3127 a_540459_681940.n17 a_540459_681940.t27 3.48
R3128 a_540459_681940.n16 a_540459_681940.t19 3.48
R3129 a_540459_681940.n15 a_540459_681940.t15 3.48
R3130 a_540459_681940.n5 a_540459_681940.t5 3.48
R3131 a_540459_681940.n22 a_540459_681940.t9 3.48
R3132 a_540459_681940.n6 a_540459_681940.t1 3.48
R3133 a_540459_681940.n32 a_540459_681940.t7 3.48
R3134 a_540459_681940.n30 a_540459_681940.t10 3.48
R3135 a_540459_681940.n29 a_540459_681940.t12 3.48
R3136 a_540459_681940.n28 a_540459_681940.t0 3.48
R3137 a_540459_681940.n4 a_540459_681940.t8 3.498
R3138 a_540459_681940.n10 a_540459_681940.t16 3.48
R3139 a_540459_681940.t26 a_540459_681940.n36 3.48
R3140 a_540459_681940.n29 a_540459_681940.n28 2.783
R3141 a_540459_681940.n30 a_540459_681940.n29 2.759
R3142 a_540459_681940.n26 a_540459_681940.n25 2.722
R3143 a_540459_681940.n25 a_540459_681940.n24 2.71
R3144 a_540459_681940.n18 a_540459_681940.n17 2.465
R3145 a_540459_681940.n19 a_540459_681940.n18 2.465
R3146 a_540459_681940.n12 a_540459_681940.n11 2.465
R3147 a_540459_681940.n13 a_540459_681940.n12 2.465
R3148 a_540459_681940.n11 a_540459_681940.n10 2.448
R3149 a_540459_681940.n17 a_540459_681940.n16 2.438
R3150 a_540459_681940.n8 a_540459_681940.n19 2.412
R3151 a_540459_681940.n0 a_540459_681940.n13 2.412
R3152 a_540459_681940.n36 a_540459_681940.n0 2.223
R3153 a_540459_681940.n8 a_540459_681940.n15 2.223
R3154 a_540459_681940.n31 a_540459_681940.n30 2.2
R3155 a_540459_681940.n27 a_540459_681940.n26 2.19
R3156 a_540459_681940.n23 a_540459_681940.n22 2.08
R3157 a_540459_681940.n33 a_540459_681940.n32 2.051
R3158 a_540459_681940.n4 a_540459_681940.n3 1.115
R3159 a_540459_681940.n0 a_540459_681940.n35 1.092
R3160 a_540459_681940.n4 a_540459_681940.n1 0.783
R3161 a_540459_681940.n9 a_540459_681940.n27 0.734
R3162 a_540459_681940.n7 a_540459_681940.n31 0.687
R3163 a_540459_681940.n9 a_540459_681940.n23 0.624
R3164 a_540459_681940.n7 a_540459_681940.n33 0.573
R3165 a_540459_681940.n0 a_540459_681940.n8 0.318
R3166 a_540459_681940.n4 a_540459_681940.n2 0.084
R3167 a_540459_681940.n7 a_540459_681940.n9 0.08
R3168 a_540459_681940.n0 a_540459_681940.n14 0.032
R3169 a_540459_681940.n8 a_540459_681940.n20 0.027
R3170 a_540459_681940.n10 a_540459_681940.n3 0.02
R3171 a_540459_681940.n7 a_540459_681940.n6 0.018
R3172 a_540459_681940.n9 a_540459_681940.n5 0.018
R3173 a_540459_681940.n35 a_540459_681940.n7 0.015
R3174 io_analog[1].n0 io_analog[1].t6 136.549
R3175 io_analog[1].n5 io_analog[1].t4 132.921
R3176 io_analog[1].n0 io_analog[1].t2 132.921
R3177 io_analog[1].n4 io_analog[1].t1 132.92
R3178 io_analog[1].n3 io_analog[1].t0 132.918
R3179 io_analog[1].n2 io_analog[1].t3 132.918
R3180 io_analog[1].n1 io_analog[1].t5 132.918
R3181 io_analog[1] io_analog[1].n5 11.861
R3182 io_analog[1].n2 io_analog[1].n1 3.578
R3183 io_analog[1].n3 io_analog[1].n2 3.578
R3184 io_analog[1].n4 io_analog[1].n3 3.575
R3185 io_analog[1].n1 io_analog[1].n0 3.574
R3186 io_analog[1].n5 io_analog[1].n4 3.569
R3187 a_541059_678436.n2 a_541059_678436.t4 4.732
R3188 a_541059_678436.n9 a_541059_678436.t6 4.731
R3189 a_541059_678436.n5 a_541059_678436.t5 3.504
R3190 a_541059_678436.n0 a_541059_678436.t9 3.48
R3191 a_541059_678436.n6 a_541059_678436.t7 3.48
R3192 a_541059_678436.n1 a_541059_678436.t8 3.48
R3193 a_541059_678436.n2 a_541059_678436.t3 2.458
R3194 a_541059_678436.n8 a_541059_678436.t1 2.401
R3195 a_541059_678436.n3 a_541059_678436.t2 2.401
R3196 a_541059_678436.n9 a_541059_678436.n8 0.26
R3197 a_541059_678436.n3 a_541059_678436.n2 0.257
R3198 a_541059_678436.n7 a_541059_678436.n5 0.222
R3199 a_541059_678436.t0 a_541059_678436.n9 0.056
R3200 a_541059_678436.n9 a_541059_678436.n0 0.055
R3201 a_541059_678436.n2 a_541059_678436.n1 0.053
R3202 a_541059_678436.n8 a_541059_678436.n7 0.031
R3203 a_541059_678436.n4 a_541059_678436.n3 0.012
R3204 a_541059_678436.n5 a_541059_678436.n4 0.005
R3205 a_541059_678436.n7 a_541059_678436.n6 0.002
R3206 a_41722_677112.n4 a_41722_677112.t7 3.48
R3207 a_41722_677112.n4 a_41722_677112.t3 3.48
R3208 a_41722_677112.n5 a_41722_677112.t5 3.48
R3209 a_41722_677112.n5 a_41722_677112.t6 3.48
R3210 a_41722_677112.n1 a_41722_677112.t2 3.48
R3211 a_41722_677112.n1 a_41722_677112.t4 3.48
R3212 a_41722_677112.n0 a_41722_677112.t1 2.841
R3213 a_41722_677112.n0 a_41722_677112.t9 2.401
R3214 a_41722_677112.n9 a_41722_677112.t8 2.401
R3215 a_41722_677112.n8 a_41722_677112.n7 0.937
R3216 a_41722_677112.n3 a_41722_677112.n2 0.937
R3217 a_41722_677112.n6 a_41722_677112.n5 0.532
R3218 a_41722_677112.n2 a_41722_677112.n1 0.532
R3219 a_41722_677112.n7 a_41722_677112.n4 0.532
R3220 a_41722_677112.t0 a_41722_677112.n9 0.446
R3221 a_41722_677112.n7 a_41722_677112.n6 0.305
R3222 a_41722_677112.n8 a_41722_677112.n3 0.292
R3223 a_41722_677112.n9 a_41722_677112.n8 0.078
R3224 a_41722_677112.n3 a_41722_677112.n0 0.066
R3225 a_43833_677960.n27 a_43833_677960.t6 147.028
R3226 a_43833_677960.n30 a_43833_677960.t8 147.028
R3227 a_43833_677960.n33 a_43833_677960.t16 135.931
R3228 a_43833_677960.n16 a_43833_677960.t23 135.931
R3229 a_43833_677960.n1 a_43833_677960.t27 135.931
R3230 a_43833_677960.n40 a_43833_677960.t10 135.931
R3231 a_43833_677960.n37 a_43833_677960.t14 135.928
R3232 a_43833_677960.n36 a_43833_677960.t18 135.928
R3233 a_43833_677960.n41 a_43833_677960.t20 135.928
R3234 a_43833_677960.n48 a_43833_677960.t12 135.928
R3235 a_43833_677960.n15 a_43833_677960.t25 135.928
R3236 a_43833_677960.n4 a_43833_677960.t24 135.928
R3237 a_43833_677960.n3 a_43833_677960.t22 135.928
R3238 a_43833_677960.n2 a_43833_677960.t26 135.928
R3239 a_43833_677960.n29 a_43833_677960.t9 6.96
R3240 a_43833_677960.n26 a_43833_677960.t7 6.96
R3241 a_43833_677960.n32 a_43833_677960.t15 5.713
R3242 a_43833_677960.n32 a_43833_677960.t11 5.713
R3243 a_43833_677960.n34 a_43833_677960.t17 5.713
R3244 a_43833_677960.n34 a_43833_677960.t19 5.713
R3245 a_43833_677960.t21 a_43833_677960.n50 5.713
R3246 a_43833_677960.n50 a_43833_677960.t13 5.713
R3247 a_43833_677960.n47 a_43833_677960.t1 3.985
R3248 a_43833_677960.n44 a_43833_677960.t4 3.985
R3249 a_43833_677960.n7 a_43833_677960.n6 3.522
R3250 a_43833_677960.n43 a_43833_677960.t0 3.48
R3251 a_43833_677960.n43 a_43833_677960.t5 3.48
R3252 a_43833_677960.n42 a_43833_677960.t3 3.48
R3253 a_43833_677960.n42 a_43833_677960.t2 3.48
R3254 a_43833_677960.n22 a_43833_677960.n21 3.474
R3255 a_43833_677960.n48 a_43833_677960.n47 2.547
R3256 a_43833_677960.n50 a_43833_677960.n24 1.435
R3257 a_43833_677960.n35 a_43833_677960.n34 1.429
R3258 a_43833_677960.n50 a_43833_677960.n49 1.429
R3259 a_43833_677960.n38 a_43833_677960.n32 1.413
R3260 a_43833_677960.n26 a_43833_677960.n25 0.954
R3261 a_43833_677960.n29 a_43833_677960.n28 0.954
R3262 a_43833_677960.n27 a_43833_677960.n26 0.921
R3263 a_43833_677960.n30 a_43833_677960.n29 0.921
R3264 a_43833_677960.n16 a_43833_677960.n15 0.646
R3265 a_43833_677960.n14 a_43833_677960.n13 0.645
R3266 a_43833_677960.n3 a_43833_677960.n2 0.645
R3267 a_43833_677960.n18 a_43833_677960.n17 0.645
R3268 a_43833_677960.n19 a_43833_677960.n18 0.645
R3269 a_43833_677960.n20 a_43833_677960.n19 0.645
R3270 a_43833_677960.n21 a_43833_677960.n20 0.645
R3271 a_43833_677960.n37 a_43833_677960.n36 0.645
R3272 a_43833_677960.n11 a_43833_677960.n10 0.645
R3273 a_43833_677960.n2 a_43833_677960.n1 0.645
R3274 a_43833_677960.n41 a_43833_677960.n40 0.635
R3275 a_43833_677960.n39 a_43833_677960.n31 0.61
R3276 a_43833_677960.n46 a_43833_677960.n42 0.505
R3277 a_43833_677960.n23 a_43833_677960.n0 0.46
R3278 a_43833_677960.n8 a_43833_677960.n7 0.455
R3279 a_43833_677960.n45 a_43833_677960.n43 0.45
R3280 a_43833_677960.n12 a_43833_677960.n5 0.375
R3281 a_43833_677960.n35 a_43833_677960.n33 0.328
R3282 a_43833_677960.n9 a_43833_677960.n8 0.328
R3283 a_43833_677960.n24 a_43833_677960.n23 0.323
R3284 a_43833_677960.n24 a_43833_677960.n14 0.322
R3285 a_43833_677960.n49 a_43833_677960.n41 0.322
R3286 a_43833_677960.n49 a_43833_677960.n48 0.322
R3287 a_43833_677960.n36 a_43833_677960.n35 0.317
R3288 a_43833_677960.n10 a_43833_677960.n9 0.317
R3289 a_43833_677960.n47 a_43833_677960.n46 0.305
R3290 a_43833_677960.n13 a_43833_677960.n12 0.29
R3291 a_43833_677960.n5 a_43833_677960.n4 0.29
R3292 a_43833_677960.n38 a_43833_677960.n37 0.289
R3293 a_43833_677960.n46 a_43833_677960.n45 0.287
R3294 a_43833_677960.n45 a_43833_677960.n44 0.287
R3295 a_43833_677960.n5 a_43833_677960.n3 0.27
R3296 a_43833_677960.n12 a_43833_677960.n11 0.27
R3297 a_43833_677960.n40 a_43833_677960.n39 0.233
R3298 a_43833_677960.n31 a_43833_677960.n27 0.147
R3299 a_43833_677960.n31 a_43833_677960.n30 0.147
R3300 a_43833_677960.n0 a_43833_677960.n16 0.084
R3301 a_43833_677960.n0 a_43833_677960.n22 0.053
R3302 a_43833_677960.n39 a_43833_677960.n38 0.031
R3303 io_analog[0].n0 io_analog[0].t3 136.549
R3304 io_analog[0].n5 io_analog[0].t1 132.921
R3305 io_analog[0].n0 io_analog[0].t6 132.921
R3306 io_analog[0].n4 io_analog[0].t5 132.92
R3307 io_analog[0].n3 io_analog[0].t4 132.918
R3308 io_analog[0].n2 io_analog[0].t0 132.918
R3309 io_analog[0].n1 io_analog[0].t2 132.918
R3310 io_analog[0] io_analog[0].n5 5.818
R3311 io_analog[0].n2 io_analog[0].n1 3.578
R3312 io_analog[0].n3 io_analog[0].n2 3.578
R3313 io_analog[0].n4 io_analog[0].n3 3.575
R3314 io_analog[0].n1 io_analog[0].n0 3.574
R3315 io_analog[0].n5 io_analog[0].n4 3.569
C0 io_analog[10] io_analog[9] 2.02fF
C1 vccd1 io_analog[2] 51.50fF
C2 vccd1 io_analog[0] 1.08fF
C3 io_analog[2] io_analog[1] 0.85fF
C4 io_analog[10] io_analog[8] 0.77fF
C5 io_analog[10] vccd2 31.93fF
C6 io_analog[1] io_analog[0] 0.94fF
C7 io_analog[8] io_analog[9] 0.24fF
C8 vccd1 io_analog[1] 1.51fF
C9 io_analog[2] io_analog[0] 0.60fF
C10 io_analog[8] vccd2 13.23fF
C11 io_analog[0] vssa2 175.84fF
C12 io_analog[1] vssa2 143.75fF
C13 io_analog[2] vssa2 272.06fF
C14 io_analog[9] vssa2 104.20fF
C15 io_analog[8] vssa2 114.04fF
C16 io_analog[10] vssa2 240.56fF
C17 vccd1 vssa2 497.18fF
C18 vccd2 vssa2 593.03fF
C19 io_analog[0].t1 vssa2 0.03fF
C20 io_analog[0].t5 vssa2 0.03fF
C21 io_analog[0].t4 vssa2 0.03fF
C22 io_analog[0].t0 vssa2 0.03fF
C23 io_analog[0].t2 vssa2 0.03fF
C24 io_analog[0].t6 vssa2 0.03fF
C25 io_analog[0].t3 vssa2 0.03fF
C26 io_analog[0].n0 vssa2 0.14fF $ **FLOATING
C27 io_analog[0].n1 vssa2 0.07fF $ **FLOATING
C28 io_analog[0].n2 vssa2 0.07fF $ **FLOATING
C29 io_analog[0].n3 vssa2 0.07fF $ **FLOATING
C30 io_analog[0].n4 vssa2 0.07fF $ **FLOATING
C31 io_analog[0].n5 vssa2 2.70fF $ **FLOATING
C32 a_43833_677960.n0 vssa2 0.18fF $ **FLOATING
C33 a_43833_677960.t27 vssa2 0.60fF
C34 a_43833_677960.n1 vssa2 0.40fF $ **FLOATING
C35 a_43833_677960.t26 vssa2 0.60fF
C36 a_43833_677960.n2 vssa2 0.44fF $ **FLOATING
C37 a_43833_677960.t22 vssa2 0.60fF
C38 a_43833_677960.n3 vssa2 0.42fF $ **FLOATING
C39 a_43833_677960.t24 vssa2 0.60fF
C40 a_43833_677960.n4 vssa2 0.42fF $ **FLOATING
C41 a_43833_677960.n5 vssa2 0.17fF $ **FLOATING
C42 a_43833_677960.n6 vssa2 0.70fF $ **FLOATING
C43 a_43833_677960.n7 vssa2 0.49fF $ **FLOATING
C44 a_43833_677960.n8 vssa2 0.52fF $ **FLOATING
C45 a_43833_677960.n9 vssa2 0.11fF $ **FLOATING
C46 a_43833_677960.n10 vssa2 0.42fF $ **FLOATING
C47 a_43833_677960.n11 vssa2 0.42fF $ **FLOATING
C48 a_43833_677960.n12 vssa2 0.25fF $ **FLOATING
C49 a_43833_677960.n13 vssa2 0.42fF $ **FLOATING
C50 a_43833_677960.n14 vssa2 0.42fF $ **FLOATING
C51 a_43833_677960.t25 vssa2 0.60fF
C52 a_43833_677960.n15 vssa2 0.44fF $ **FLOATING
C53 a_43833_677960.t23 vssa2 0.60fF
C54 a_43833_677960.n16 vssa2 0.40fF $ **FLOATING
C55 a_43833_677960.n17 vssa2 0.44fF $ **FLOATING
C56 a_43833_677960.n18 vssa2 0.44fF $ **FLOATING
C57 a_43833_677960.n19 vssa2 0.44fF $ **FLOATING
C58 a_43833_677960.n20 vssa2 0.44fF $ **FLOATING
C59 a_43833_677960.n21 vssa2 0.70fF $ **FLOATING
C60 a_43833_677960.n22 vssa2 0.32fF $ **FLOATING
C61 a_43833_677960.n23 vssa2 0.52fF $ **FLOATING
C62 a_43833_677960.n24 vssa2 0.11fF $ **FLOATING
C63 a_43833_677960.t10 vssa2 0.60fF
C64 a_43833_677960.t6 vssa2 0.16fF
C65 a_43833_677960.t7 vssa2 0.04fF
C66 a_43833_677960.n25 vssa2 0.19fF $ **FLOATING
C67 a_43833_677960.n26 vssa2 0.30fF $ **FLOATING
C68 a_43833_677960.n27 vssa2 0.18fF $ **FLOATING
C69 a_43833_677960.t9 vssa2 0.04fF
C70 a_43833_677960.n28 vssa2 0.19fF $ **FLOATING
C71 a_43833_677960.n29 vssa2 0.30fF $ **FLOATING
C72 a_43833_677960.t8 vssa2 0.16fF
C73 a_43833_677960.n30 vssa2 0.18fF $ **FLOATING
C74 a_43833_677960.n31 vssa2 0.17fF $ **FLOATING
C75 a_43833_677960.t15 vssa2 0.08fF
C76 a_43833_677960.t11 vssa2 0.08fF
C77 a_43833_677960.n32 vssa2 0.47fF $ **FLOATING
C78 a_43833_677960.t16 vssa2 0.60fF
C79 a_43833_677960.n33 vssa2 1.42fF $ **FLOATING
C80 a_43833_677960.t17 vssa2 0.08fF
C81 a_43833_677960.t19 vssa2 0.08fF
C82 a_43833_677960.n34 vssa2 0.47fF $ **FLOATING
C83 a_43833_677960.n35 vssa2 0.11fF $ **FLOATING
C84 a_43833_677960.t18 vssa2 0.60fF
C85 a_43833_677960.n36 vssa2 0.42fF $ **FLOATING
C86 a_43833_677960.t14 vssa2 0.60fF
C87 a_43833_677960.n37 vssa2 0.42fF $ **FLOATING
C88 a_43833_677960.n38 vssa2 0.10fF $ **FLOATING
C89 a_43833_677960.n39 vssa2 0.16fF $ **FLOATING
C90 a_43833_677960.n40 vssa2 0.42fF $ **FLOATING
C91 a_43833_677960.t20 vssa2 0.60fF
C92 a_43833_677960.n41 vssa2 0.43fF $ **FLOATING
C93 a_43833_677960.t12 vssa2 0.60fF
C94 a_43833_677960.t1 vssa2 0.14fF
C95 a_43833_677960.t2 vssa2 0.08fF
C96 a_43833_677960.t3 vssa2 0.08fF
C97 a_43833_677960.n42 vssa2 0.41fF $ **FLOATING
C98 a_43833_677960.t5 vssa2 0.08fF
C99 a_43833_677960.t0 vssa2 0.08fF
C100 a_43833_677960.n43 vssa2 0.41fF $ **FLOATING
C101 a_43833_677960.t4 vssa2 0.14fF
C102 a_43833_677960.n44 vssa2 1.80fF $ **FLOATING
C103 a_43833_677960.n45 vssa2 0.58fF $ **FLOATING
C104 a_43833_677960.n46 vssa2 0.43fF $ **FLOATING
C105 a_43833_677960.n47 vssa2 1.84fF $ **FLOATING
C106 a_43833_677960.n48 vssa2 1.39fF $ **FLOATING
C107 a_43833_677960.n49 vssa2 0.10fF $ **FLOATING
C108 a_43833_677960.t13 vssa2 0.08fF
C109 a_43833_677960.n50 vssa2 0.47fF $ **FLOATING
C110 a_43833_677960.t21 vssa2 0.08fF
C111 a_41722_677112.t8 vssa2 0.20fF
C112 a_41722_677112.t9 vssa2 0.20fF
C113 a_41722_677112.t1 vssa2 0.45fF
C114 a_41722_677112.n0 vssa2 3.38fF $ **FLOATING
C115 a_41722_677112.t4 vssa2 0.02fF
C116 a_41722_677112.t2 vssa2 0.02fF
C117 a_41722_677112.n1 vssa2 0.12fF $ **FLOATING
C118 a_41722_677112.n2 vssa2 0.19fF $ **FLOATING
C119 a_41722_677112.n3 vssa2 0.57fF $ **FLOATING
C120 a_41722_677112.t3 vssa2 0.02fF
C121 a_41722_677112.t7 vssa2 0.02fF
C122 a_41722_677112.n4 vssa2 0.12fF $ **FLOATING
C123 a_41722_677112.t6 vssa2 0.02fF
C124 a_41722_677112.t5 vssa2 0.02fF
C125 a_41722_677112.n5 vssa2 0.12fF $ **FLOATING
C126 a_41722_677112.n6 vssa2 0.13fF $ **FLOATING
C127 a_41722_677112.n7 vssa2 0.19fF $ **FLOATING
C128 a_41722_677112.n8 vssa2 0.59fF $ **FLOATING
C129 a_41722_677112.n9 vssa2 2.05fF $ **FLOATING
C130 a_41722_677112.t0 vssa2 2.50fF
C131 a_541059_678436.t9 vssa2 0.03fF
C132 a_541059_678436.n0 vssa2 0.35fF $ **FLOATING
C133 a_541059_678436.t6 vssa2 0.12fF
C134 a_541059_678436.t1 vssa2 0.25fF
C135 a_541059_678436.t2 vssa2 0.25fF
C136 a_541059_678436.t4 vssa2 0.12fF
C137 a_541059_678436.t8 vssa2 0.03fF
C138 a_541059_678436.n1 vssa2 0.35fF $ **FLOATING
C139 a_541059_678436.t3 vssa2 0.32fF
C140 a_541059_678436.n2 vssa2 4.27fF $ **FLOATING
C141 a_541059_678436.n3 vssa2 2.58fF $ **FLOATING
C142 a_541059_678436.n4 vssa2 1.11fF $ **FLOATING
C143 a_541059_678436.t5 vssa2 0.03fF
C144 a_541059_678436.n5 vssa2 0.37fF $ **FLOATING
C145 a_541059_678436.t7 vssa2 0.03fF
C146 a_541059_678436.n6 vssa2 0.40fF $ **FLOATING
C147 a_541059_678436.n7 vssa2 1.14fF $ **FLOATING
C148 a_541059_678436.n8 vssa2 2.65fF $ **FLOATING
C149 a_541059_678436.n9 vssa2 1.49fF $ **FLOATING
C150 a_541059_678436.t0 vssa2 3.10fF
C151 io_analog[1].t4 vssa2 0.03fF
C152 io_analog[1].t1 vssa2 0.03fF
C153 io_analog[1].t0 vssa2 0.03fF
C154 io_analog[1].t3 vssa2 0.03fF
C155 io_analog[1].t5 vssa2 0.03fF
C156 io_analog[1].t2 vssa2 0.03fF
C157 io_analog[1].t6 vssa2 0.04fF
C158 io_analog[1].n0 vssa2 0.15fF $ **FLOATING
C159 io_analog[1].n1 vssa2 0.07fF $ **FLOATING
C160 io_analog[1].n2 vssa2 0.07fF $ **FLOATING
C161 io_analog[1].n3 vssa2 0.07fF $ **FLOATING
C162 io_analog[1].n4 vssa2 0.07fF $ **FLOATING
C163 io_analog[1].n5 vssa2 1.69fF $ **FLOATING
C164 a_540459_681940.n0 vssa2 3.68fF $ **FLOATING
C165 a_540459_681940.n1 vssa2 0.40fF $ **FLOATING
C166 a_540459_681940.t8 vssa2 0.13fF
C167 a_540459_681940.t4 vssa2 0.14fF
C168 a_540459_681940.n2 vssa2 1.72fF $ **FLOATING
C169 a_540459_681940.n3 vssa2 3.32fF $ **FLOATING
C170 a_540459_681940.n4 vssa2 3.62fF $ **FLOATING
C171 a_540459_681940.n5 vssa2 0.56fF $ **FLOATING
C172 a_540459_681940.n6 vssa2 0.55fF $ **FLOATING
C173 a_540459_681940.n7 vssa2 0.75fF $ **FLOATING
C174 a_540459_681940.n8 vssa2 1.67fF $ **FLOATING
C175 a_540459_681940.n9 vssa2 0.65fF $ **FLOATING
C176 a_540459_681940.t20 vssa2 0.70fF
C177 a_540459_681940.t22 vssa2 0.13fF
C178 a_540459_681940.t18 vssa2 0.13fF
C179 a_540459_681940.t25 vssa2 0.13fF
C180 a_540459_681940.t16 vssa2 0.13fF
C181 a_540459_681940.n10 vssa2 0.91fF $ **FLOATING
C182 a_540459_681940.n11 vssa2 1.42fF $ **FLOATING
C183 a_540459_681940.n12 vssa2 1.41fF $ **FLOATING
C184 a_540459_681940.n13 vssa2 1.42fF $ **FLOATING
C185 a_540459_681940.t14 vssa2 0.13fF
C186 a_540459_681940.n14 vssa2 0.49fF $ **FLOATING
C187 a_540459_681940.t15 vssa2 0.13fF
C188 a_540459_681940.t23 vssa2 0.70fF
C189 a_540459_681940.n15 vssa2 2.18fF $ **FLOATING
C190 a_540459_681940.t24 vssa2 0.13fF
C191 a_540459_681940.t21 vssa2 0.13fF
C192 a_540459_681940.t27 vssa2 0.13fF
C193 a_540459_681940.t19 vssa2 0.13fF
C194 a_540459_681940.n16 vssa2 2.09fF $ **FLOATING
C195 a_540459_681940.n17 vssa2 1.42fF $ **FLOATING
C196 a_540459_681940.n18 vssa2 1.41fF $ **FLOATING
C197 a_540459_681940.n19 vssa2 1.42fF $ **FLOATING
C198 a_540459_681940.t17 vssa2 0.13fF
C199 a_540459_681940.n20 vssa2 0.49fF $ **FLOATING
C200 a_540459_681940.t5 vssa2 0.13fF
C201 a_540459_681940.n21 vssa2 0.05fF $ **FLOATING
C202 a_540459_681940.t9 vssa2 0.13fF
C203 a_540459_681940.t2 vssa2 0.71fF
C204 a_540459_681940.n22 vssa2 1.99fF $ **FLOATING
C205 a_540459_681940.n23 vssa2 0.35fF $ **FLOATING
C206 a_540459_681940.t6 vssa2 0.13fF
C207 a_540459_681940.t3 vssa2 0.13fF
C208 a_540459_681940.t13 vssa2 0.13fF
C209 a_540459_681940.n24 vssa2 1.34fF $ **FLOATING
C210 a_540459_681940.n25 vssa2 1.37fF $ **FLOATING
C211 a_540459_681940.n26 vssa2 1.25fF $ **FLOATING
C212 a_540459_681940.n27 vssa2 0.40fF $ **FLOATING
C213 a_540459_681940.t10 vssa2 0.13fF
C214 a_540459_681940.t12 vssa2 0.13fF
C215 a_540459_681940.t0 vssa2 0.13fF
C216 a_540459_681940.n28 vssa2 1.30fF $ **FLOATING
C217 a_540459_681940.n29 vssa2 1.29fF $ **FLOATING
C218 a_540459_681940.n30 vssa2 1.31fF $ **FLOATING
C219 a_540459_681940.n31 vssa2 0.39fF $ **FLOATING
C220 a_540459_681940.t7 vssa2 0.13fF
C221 a_540459_681940.t11 vssa2 0.69fF
C222 a_540459_681940.n32 vssa2 1.99fF $ **FLOATING
C223 a_540459_681940.n33 vssa2 0.33fF $ **FLOATING
C224 a_540459_681940.t1 vssa2 0.13fF
C225 a_540459_681940.n34 vssa2 0.05fF $ **FLOATING
C226 a_540459_681940.n35 vssa2 2.11fF $ **FLOATING
C227 a_540459_681940.n36 vssa2 2.18fF $ **FLOATING
C228 a_540459_681940.t26 vssa2 0.13fF
C229 a_37693_693523.t4 vssa2 19.79fF
C230 a_37693_693523.t5 vssa2 19.79fF
C231 a_37693_693523.t3 vssa2 19.79fF
C232 a_37693_693523.t6 vssa2 19.79fF
C233 a_37693_693523.t2 vssa2 0.51fF
C234 a_37693_693523.t1 vssa2 0.51fF
C235 a_37693_693523.n0 vssa2 8.33fF $ **FLOATING
C236 a_37693_693523.n1 vssa2 10.84fF $ **FLOATING
C237 a_37693_693523.n2 vssa2 9.18fF $ **FLOATING
C238 a_37693_693523.n3 vssa2 9.18fF $ **FLOATING
C239 a_37693_693523.n4 vssa2 10.85fF $ **FLOATING
C240 a_37693_693523.t7 vssa2 0.51fF
C241 a_37693_693523.n5 vssa2 6.62fF $ **FLOATING
C242 a_37693_693523.t0 vssa2 2.22fF
C243 io_analog[8].t5 vssa2 0.03fF
C244 io_analog[8].t1 vssa2 0.03fF
C245 io_analog[8].t4 vssa2 0.03fF
C246 io_analog[8].t6 vssa2 0.03fF
C247 io_analog[8].t3 vssa2 0.03fF
C248 io_analog[8].n0 vssa2 0.02fF $ **FLOATING
C249 io_analog[8].n1 vssa2 0.07fF $ **FLOATING
C250 io_analog[8].n2 vssa2 0.02fF $ **FLOATING
C251 io_analog[8].n3 vssa2 0.02fF $ **FLOATING
C252 io_analog[8].n4 vssa2 0.02fF $ **FLOATING
C253 io_analog[8].n5 vssa2 0.02fF $ **FLOATING
C254 io_analog[8].n6 vssa2 0.03fF $ **FLOATING
C255 io_analog[8].t0 vssa2 0.03fF
C256 io_analog[8].t2 vssa2 0.03fF
C257 io_analog[8].n7 vssa2 0.07fF $ **FLOATING
C258 io_analog[8].n8 vssa2 0.02fF $ **FLOATING
C259 io_analog[8].n9 vssa2 0.02fF $ **FLOATING
C260 io_analog[8].n10 vssa2 0.02fF $ **FLOATING
C261 io_analog[8].n11 vssa2 0.02fF $ **FLOATING
C262 io_analog[8].n12 vssa2 0.03fF $ **FLOATING
C263 io_analog[8].n13 vssa2 4.22fF $ **FLOATING
C264 io_analog[2].t52 vssa2 19.75fF
C265 io_analog[2].n0 vssa2 2.28fF $ **FLOATING
C266 io_analog[2].t1 vssa2 0.02fF
C267 io_analog[2].n1 vssa2 0.10fF $ **FLOATING
C268 io_analog[2].n2 vssa2 0.23fF $ **FLOATING
C269 io_analog[2].t15 vssa2 0.01fF
C270 io_analog[2].n3 vssa2 0.21fF $ **FLOATING
C271 io_analog[2].t11 vssa2 0.01fF
C272 io_analog[2].n4 vssa2 0.19fF $ **FLOATING
C273 io_analog[2].t7 vssa2 0.01fF
C274 io_analog[2].t30 vssa2 0.02fF
C275 io_analog[2].n5 vssa2 0.34fF $ **FLOATING
C276 io_analog[2].t16 vssa2 0.02fF
C277 io_analog[2].t5 vssa2 0.01fF
C278 io_analog[2].n6 vssa2 0.12fF $ **FLOATING
C279 io_analog[2].t10 vssa2 0.01fF
C280 io_analog[2].n7 vssa2 0.12fF $ **FLOATING
C281 io_analog[2].t12 vssa2 0.01fF
C282 io_analog[2].n8 vssa2 0.16fF $ **FLOATING
C283 io_analog[2].n9 vssa2 0.07fF $ **FLOATING
C284 io_analog[2].t31 vssa2 0.01fF
C285 io_analog[2].n10 vssa2 0.06fF $ **FLOATING
C286 io_analog[2].n11 vssa2 0.04fF $ **FLOATING
C287 io_analog[2].n12 vssa2 0.16fF $ **FLOATING
C288 io_analog[2].n13 vssa2 0.07fF $ **FLOATING
C289 io_analog[2].t23 vssa2 0.01fF
C290 io_analog[2].n14 vssa2 0.06fF $ **FLOATING
C291 io_analog[2].n15 vssa2 0.04fF $ **FLOATING
C292 io_analog[2].n16 vssa2 0.16fF $ **FLOATING
C293 io_analog[2].n17 vssa2 0.30fF $ **FLOATING
C294 io_analog[2].t9 vssa2 0.01fF
C295 io_analog[2].t3 vssa2 0.06fF
C296 io_analog[2].t37 vssa2 0.02fF
C297 io_analog[2].t54 vssa2 19.82fF
C298 io_analog[2].t55 vssa2 20.00fF
C299 io_analog[2].t53 vssa2 19.95fF
C300 io_analog[2].n18 vssa2 2.57fF $ **FLOATING
C301 io_analog[2].t0 vssa2 0.06fF
C302 io_analog[2].t36 vssa2 0.02fF
C303 io_analog[2].t8 vssa2 0.01fF
C304 io_analog[2].n19 vssa2 0.16fF $ **FLOATING
C305 io_analog[2].n20 vssa2 1.50fF $ **FLOATING
C306 io_analog[2].t24 vssa2 0.01fF
C307 io_analog[2].n21 vssa2 0.21fF $ **FLOATING
C308 io_analog[2].t21 vssa2 0.01fF
C309 io_analog[2].n22 vssa2 0.34fF $ **FLOATING
C310 io_analog[2].t27 vssa2 0.01fF
C311 io_analog[2].t39 vssa2 0.01fF
C312 io_analog[2].n23 vssa2 0.09fF $ **FLOATING
C313 io_analog[2].t47 vssa2 0.01fF
C314 io_analog[2].n24 vssa2 0.27fF $ **FLOATING
C315 io_analog[2].t42 vssa2 0.01fF
C316 io_analog[2].t48 vssa2 0.01fF
C317 io_analog[2].t43 vssa2 0.01fF
C318 io_analog[2].t49 vssa2 0.01fF
C319 io_analog[2].t46 vssa2 0.01fF
C320 io_analog[2].t51 vssa2 0.01fF
C321 io_analog[2].t45 vssa2 0.01fF
C322 io_analog[2].t50 vssa2 0.01fF
C323 io_analog[2].t44 vssa2 0.08fF
C324 io_analog[2].n25 vssa2 0.23fF $ **FLOATING
C325 io_analog[2].n26 vssa2 0.10fF $ **FLOATING
C326 io_analog[2].n27 vssa2 0.08fF $ **FLOATING
C327 io_analog[2].n28 vssa2 0.15fF $ **FLOATING
C328 io_analog[2].n29 vssa2 0.15fF $ **FLOATING
C329 io_analog[2].t41 vssa2 0.01fF
C330 io_analog[2].n30 vssa2 0.18fF $ **FLOATING
C331 io_analog[2].n31 vssa2 0.16fF $ **FLOATING
C332 io_analog[2].n32 vssa2 0.04fF $ **FLOATING
C333 io_analog[2].n33 vssa2 0.05fF $ **FLOATING
C334 io_analog[2].n34 vssa2 0.05fF $ **FLOATING
C335 io_analog[2].n35 vssa2 0.15fF $ **FLOATING
C336 io_analog[2].n36 vssa2 0.04fF $ **FLOATING
C337 io_analog[2].n37 vssa2 0.05fF $ **FLOATING
C338 io_analog[2].n38 vssa2 0.05fF $ **FLOATING
C339 io_analog[2].n39 vssa2 0.15fF $ **FLOATING
C340 io_analog[2].t40 vssa2 0.02fF
C341 io_analog[2].n40 vssa2 0.32fF $ **FLOATING
C342 io_analog[2].t28 vssa2 0.01fF
C343 io_analog[2].t13 vssa2 0.02fF
C344 io_analog[2].n41 vssa2 0.10fF $ **FLOATING
C345 io_analog[2].n42 vssa2 0.16fF $ **FLOATING
C346 io_analog[2].n43 vssa2 0.04fF $ **FLOATING
C347 io_analog[2].t38 vssa2 0.01fF
C348 io_analog[2].n44 vssa2 0.06fF $ **FLOATING
C349 io_analog[2].t25 vssa2 0.01fF
C350 io_analog[2].n45 vssa2 0.19fF $ **FLOATING
C351 io_analog[2].t19 vssa2 0.01fF
C352 io_analog[2].n46 vssa2 0.16fF $ **FLOATING
C353 io_analog[2].n47 vssa2 0.04fF $ **FLOATING
C354 io_analog[2].t34 vssa2 0.01fF
C355 io_analog[2].n48 vssa2 0.06fF $ **FLOATING
C356 io_analog[2].n49 vssa2 0.04fF $ **FLOATING
C357 io_analog[2].n50 vssa2 0.16fF $ **FLOATING
C358 io_analog[2].n51 vssa2 0.04fF $ **FLOATING
C359 io_analog[2].n52 vssa2 0.19fF $ **FLOATING
C360 io_analog[2].t29 vssa2 0.01fF
C361 io_analog[2].t17 vssa2 0.02fF
C362 io_analog[2].n53 vssa2 0.26fF $ **FLOATING
C363 io_analog[2].n54 vssa2 0.16fF $ **FLOATING
C364 io_analog[2].n55 vssa2 0.07fF $ **FLOATING
C365 io_analog[2].n56 vssa2 0.10fF $ **FLOATING
C366 io_analog[2].n57 vssa2 0.23fF $ **FLOATING
C367 io_analog[2].n58 vssa2 0.16fF $ **FLOATING
C368 io_analog[2].n59 vssa2 0.04fF $ **FLOATING
C369 io_analog[2].t35 vssa2 0.01fF
C370 io_analog[2].n60 vssa2 0.06fF $ **FLOATING
C371 io_analog[2].n61 vssa2 0.04fF $ **FLOATING
C372 io_analog[2].n62 vssa2 0.16fF $ **FLOATING
C373 io_analog[2].t32 vssa2 0.02fF
C374 io_analog[2].n63 vssa2 0.44fF $ **FLOATING
C375 io_analog[2].n64 vssa2 0.16fF $ **FLOATING
C376 io_analog[2].t18 vssa2 0.06fF
C377 io_analog[2].t6 vssa2 0.02fF
C378 io_analog[2].n65 vssa2 0.39fF $ **FLOATING
C379 io_analog[2].t14 vssa2 0.06fF
C380 io_analog[2].t2 vssa2 0.02fF
C381 io_analog[2].t22 vssa2 0.01fF
C382 io_analog[2].n66 vssa2 0.16fF $ **FLOATING
C383 io_analog[2].n67 vssa2 0.46fF $ **FLOATING
C384 io_analog[2].n68 vssa2 0.45fF $ **FLOATING
C385 io_analog[2].n69 vssa2 0.16fF $ **FLOATING
C386 io_analog[2].t20 vssa2 0.02fF
C387 io_analog[2].n70 vssa2 0.34fF $ **FLOATING
C388 io_analog[2].n71 vssa2 0.16fF $ **FLOATING
C389 io_analog[2].n72 vssa2 0.04fF $ **FLOATING
C390 io_analog[2].t26 vssa2 0.01fF
C391 io_analog[2].n73 vssa2 0.06fF $ **FLOATING
C392 io_analog[2].n74 vssa2 0.04fF $ **FLOATING
C393 io_analog[2].n75 vssa2 0.16fF $ **FLOATING
C394 io_analog[2].n76 vssa2 0.04fF $ **FLOATING
C395 io_analog[2].t33 vssa2 0.01fF
C396 io_analog[2].n77 vssa2 0.06fF $ **FLOATING
C397 io_analog[2].n78 vssa2 0.04fF $ **FLOATING
C398 io_analog[2].n79 vssa2 0.16fF $ **FLOATING
C399 io_analog[2].t4 vssa2 0.02fF
C400 io_analog[2].n80 vssa2 0.10fF $ **FLOATING
C401 io_analog[2].n81 vssa2 0.23fF $ **FLOATING
C402 io_analog[2].n82 vssa2 0.39fF $ **FLOATING
C403 io_analog[2].n83 vssa2 78.50fF $ **FLOATING
C404 constant_gm_fingers_0/Vout.n0 vssa2 4.61fF $ **FLOATING
C405 constant_gm_fingers_0/Vout.n1 vssa2 4.59fF $ **FLOATING
C406 constant_gm_fingers_0/Vout.n2 vssa2 0.89fF $ **FLOATING
C407 constant_gm_fingers_0/Vout.n3 vssa2 0.89fF $ **FLOATING
C408 constant_gm_fingers_0/Vout.n4 vssa2 0.11fF $ **FLOATING
C409 constant_gm_fingers_0/Vout.n5 vssa2 0.11fF $ **FLOATING
C410 constant_gm_fingers_0/Vout.t2 vssa2 0.07fF
C411 constant_gm_fingers_0/Vout.t0 vssa2 0.07fF
C412 constant_gm_fingers_0/Vout.n6 vssa2 0.37fF $ **FLOATING
C413 constant_gm_fingers_0/Vout.n7 vssa2 0.39fF $ **FLOATING
C414 constant_gm_fingers_0/Vout.n8 vssa2 0.39fF $ **FLOATING
C415 constant_gm_fingers_0/Vout.n9 vssa2 0.39fF $ **FLOATING
C416 constant_gm_fingers_0/Vout.n10 vssa2 0.39fF $ **FLOATING
C417 constant_gm_fingers_0/Vout.n11 vssa2 0.39fF $ **FLOATING
C418 constant_gm_fingers_0/Vout.n12 vssa2 0.73fF $ **FLOATING
C419 constant_gm_fingers_0/Vout.t40 vssa2 0.52fF
C420 constant_gm_fingers_0/Vout.t44 vssa2 0.52fF
C421 constant_gm_fingers_0/Vout.t19 vssa2 0.52fF
C422 constant_gm_fingers_0/Vout.t34 vssa2 0.52fF
C423 constant_gm_fingers_0/Vout.t27 vssa2 0.52fF
C424 constant_gm_fingers_0/Vout.t35 vssa2 0.52fF
C425 constant_gm_fingers_0/Vout.n13 vssa2 0.39fF $ **FLOATING
C426 constant_gm_fingers_0/Vout.n14 vssa2 0.39fF $ **FLOATING
C427 constant_gm_fingers_0/Vout.n15 vssa2 0.39fF $ **FLOATING
C428 constant_gm_fingers_0/Vout.n16 vssa2 0.39fF $ **FLOATING
C429 constant_gm_fingers_0/Vout.n17 vssa2 0.39fF $ **FLOATING
C430 constant_gm_fingers_0/Vout.n18 vssa2 0.43fF $ **FLOATING
C431 constant_gm_fingers_0/Vout.n19 vssa2 0.39fF $ **FLOATING
C432 constant_gm_fingers_0/Vout.n20 vssa2 0.39fF $ **FLOATING
C433 constant_gm_fingers_0/Vout.n21 vssa2 0.39fF $ **FLOATING
C434 constant_gm_fingers_0/Vout.n22 vssa2 0.39fF $ **FLOATING
C435 constant_gm_fingers_0/Vout.n23 vssa2 0.39fF $ **FLOATING
C436 constant_gm_fingers_0/Vout.n24 vssa2 0.39fF $ **FLOATING
C437 constant_gm_fingers_0/Vout.n25 vssa2 0.40fF $ **FLOATING
C438 constant_gm_fingers_0/Vout.t36 vssa2 0.52fF
C439 constant_gm_fingers_0/Vout.t29 vssa2 0.52fF
C440 constant_gm_fingers_0/Vout.t33 vssa2 0.52fF
C441 constant_gm_fingers_0/Vout.t39 vssa2 0.52fF
C442 constant_gm_fingers_0/Vout.t14 vssa2 0.52fF
C443 constant_gm_fingers_0/Vout.t16 vssa2 0.52fF
C444 constant_gm_fingers_0/Vout.t24 vssa2 0.52fF
C445 constant_gm_fingers_0/Vout.n26 vssa2 0.39fF $ **FLOATING
C446 constant_gm_fingers_0/Vout.n27 vssa2 0.39fF $ **FLOATING
C447 constant_gm_fingers_0/Vout.n28 vssa2 0.39fF $ **FLOATING
C448 constant_gm_fingers_0/Vout.n29 vssa2 0.39fF $ **FLOATING
C449 constant_gm_fingers_0/Vout.n30 vssa2 0.39fF $ **FLOATING
C450 constant_gm_fingers_0/Vout.n31 vssa2 0.39fF $ **FLOATING
C451 constant_gm_fingers_0/Vout.n32 vssa2 0.40fF $ **FLOATING
C452 constant_gm_fingers_0/Vout.n33 vssa2 4.12fF $ **FLOATING
C453 constant_gm_fingers_0/Vout.t10 vssa2 0.17fF
C454 constant_gm_fingers_0/Vout.n34 vssa2 0.39fF $ **FLOATING
C455 constant_gm_fingers_0/Vout.n35 vssa2 0.80fF $ **FLOATING
C456 constant_gm_fingers_0/Vout.t21 vssa2 0.52fF
C457 constant_gm_fingers_0/Vout.n36 vssa2 0.31fF $ **FLOATING
C458 constant_gm_fingers_0/Vout.t41 vssa2 0.52fF
C459 constant_gm_fingers_0/Vout.t17 vssa2 0.52fF
C460 constant_gm_fingers_0/Vout.n37 vssa2 0.39fF $ **FLOATING
C461 constant_gm_fingers_0/Vout.n38 vssa2 0.27fF $ **FLOATING
C462 constant_gm_fingers_0/Vout.n39 vssa2 0.19fF $ **FLOATING
C463 constant_gm_fingers_0/Vout.n40 vssa2 0.05fF $ **FLOATING
C464 constant_gm_fingers_0/Vout.t11 vssa2 0.02fF
C465 constant_gm_fingers_0/Vout.t9 vssa2 0.02fF
C466 constant_gm_fingers_0/Vout.t8 vssa2 0.17fF
C467 constant_gm_fingers_0/Vout.n41 vssa2 0.18fF $ **FLOATING
C468 constant_gm_fingers_0/Vout.n42 vssa2 0.05fF $ **FLOATING
C469 constant_gm_fingers_0/Vout.n43 vssa2 0.97fF $ **FLOATING
C470 constant_gm_fingers_0/Vout.n44 vssa2 2.73fF $ **FLOATING
C471 constant_gm_fingers_0/Vout.t3 vssa2 1.00fF
C472 constant_gm_fingers_0/Vout.t4 vssa2 0.17fF
C473 constant_gm_fingers_0/Vout.t13 vssa2 0.03fF
C474 constant_gm_fingers_0/Vout.t12 vssa2 0.03fF
C475 constant_gm_fingers_0/Vout.n45 vssa2 0.34fF $ **FLOATING
C476 constant_gm_fingers_0/Vout.n46 vssa2 0.22fF $ **FLOATING
C477 constant_gm_fingers_0/Vout.t6 vssa2 0.17fF
C478 constant_gm_fingers_0/Vout.n47 vssa2 0.18fF $ **FLOATING
C479 constant_gm_fingers_0/Vout.t7 vssa2 0.02fF
C480 constant_gm_fingers_0/Vout.t5 vssa2 0.02fF
C481 constant_gm_fingers_0/Vout.n48 vssa2 0.19fF $ **FLOATING
C482 constant_gm_fingers_0/Vout.t28 vssa2 0.52fF
C483 constant_gm_fingers_0/Vout.n49 vssa2 0.39fF $ **FLOATING
C484 constant_gm_fingers_0/Vout.n50 vssa2 0.80fF $ **FLOATING
C485 constant_gm_fingers_0/Vout.t31 vssa2 0.52fF
C486 constant_gm_fingers_0/Vout.n51 vssa2 0.31fF $ **FLOATING
C487 constant_gm_fingers_0/Vout.t22 vssa2 0.52fF
C488 constant_gm_fingers_0/Vout.n52 vssa2 0.39fF $ **FLOATING
C489 constant_gm_fingers_0/Vout.n53 vssa2 0.28fF $ **FLOATING
C490 constant_gm_fingers_0/Vout.n54 vssa2 0.05fF $ **FLOATING
C491 constant_gm_fingers_0/Vout.n55 vssa2 0.05fF $ **FLOATING
C492 constant_gm_fingers_0/Vout.n56 vssa2 0.97fF $ **FLOATING
C493 constant_gm_fingers_0/Vout.t25 vssa2 0.52fF
C494 constant_gm_fingers_0/Vout.n57 vssa2 0.39fF $ **FLOATING
C495 constant_gm_fingers_0/Vout.t32 vssa2 0.52fF
C496 constant_gm_fingers_0/Vout.n58 vssa2 0.39fF $ **FLOATING
C497 constant_gm_fingers_0/Vout.t23 vssa2 0.52fF
C498 constant_gm_fingers_0/Vout.n59 vssa2 0.39fF $ **FLOATING
C499 constant_gm_fingers_0/Vout.t38 vssa2 0.52fF
C500 constant_gm_fingers_0/Vout.n60 vssa2 0.39fF $ **FLOATING
C501 constant_gm_fingers_0/Vout.t15 vssa2 0.52fF
C502 constant_gm_fingers_0/Vout.n61 vssa2 0.39fF $ **FLOATING
C503 constant_gm_fingers_0/Vout.t18 vssa2 0.52fF
C504 constant_gm_fingers_0/Vout.n62 vssa2 0.39fF $ **FLOATING
C505 constant_gm_fingers_0/Vout.t42 vssa2 0.52fF
C506 constant_gm_fingers_0/Vout.n63 vssa2 0.40fF $ **FLOATING
C507 constant_gm_fingers_0/Vout.n64 vssa2 0.39fF $ **FLOATING
C508 constant_gm_fingers_0/Vout.n65 vssa2 0.39fF $ **FLOATING
C509 constant_gm_fingers_0/Vout.n66 vssa2 0.39fF $ **FLOATING
C510 constant_gm_fingers_0/Vout.n67 vssa2 0.39fF $ **FLOATING
C511 constant_gm_fingers_0/Vout.n68 vssa2 0.39fF $ **FLOATING
C512 constant_gm_fingers_0/Vout.n69 vssa2 0.72fF $ **FLOATING
C513 constant_gm_fingers_0/Vout.t37 vssa2 0.52fF
C514 constant_gm_fingers_0/Vout.n70 vssa2 0.39fF $ **FLOATING
C515 constant_gm_fingers_0/Vout.t43 vssa2 0.52fF
C516 constant_gm_fingers_0/Vout.n71 vssa2 0.39fF $ **FLOATING
C517 constant_gm_fingers_0/Vout.t45 vssa2 0.52fF
C518 constant_gm_fingers_0/Vout.n72 vssa2 0.39fF $ **FLOATING
C519 constant_gm_fingers_0/Vout.t20 vssa2 0.52fF
C520 constant_gm_fingers_0/Vout.n73 vssa2 0.39fF $ **FLOATING
C521 constant_gm_fingers_0/Vout.t26 vssa2 0.52fF
C522 constant_gm_fingers_0/Vout.n74 vssa2 0.39fF $ **FLOATING
C523 constant_gm_fingers_0/Vout.t30 vssa2 0.52fF
C524 constant_gm_fingers_0/Vout.n75 vssa2 0.43fF $ **FLOATING
C525 constant_gm_fingers_0/Vout.n76 vssa2 0.39fF $ **FLOATING
C526 constant_gm_fingers_0/Vout.n77 vssa2 0.39fF $ **FLOATING
C527 constant_gm_fingers_0/Vout.n78 vssa2 0.39fF $ **FLOATING
C528 constant_gm_fingers_0/Vout.n79 vssa2 0.39fF $ **FLOATING
C529 constant_gm_fingers_0/Vout.n80 vssa2 0.39fF $ **FLOATING
C530 constant_gm_fingers_0/Vout.n81 vssa2 0.39fF $ **FLOATING
C531 constant_gm_fingers_0/Vout.n82 vssa2 0.40fF $ **FLOATING
C532 constant_gm_fingers_0/Vout.n83 vssa2 4.13fF $ **FLOATING
C533 constant_gm_fingers_0/Vout.t1 vssa2 3.22fF
C534 a_540371_681998.n0 vssa2 1.85fF $ **FLOATING
C535 a_540371_681998.n1 vssa2 1.82fF $ **FLOATING
C536 a_540371_681998.n2 vssa2 0.94fF $ **FLOATING
C537 a_540371_681998.n3 vssa2 0.90fF $ **FLOATING
C538 a_540371_681998.n4 vssa2 2.10fF $ **FLOATING
C539 a_540371_681998.n5 vssa2 4.12fF $ **FLOATING
C540 a_540371_681998.n6 vssa2 0.28fF $ **FLOATING
C541 a_540371_681998.n7 vssa2 0.33fF $ **FLOATING
C542 a_540371_681998.n8 vssa2 0.02fF $ **FLOATING
C543 a_540371_681998.n9 vssa2 0.04fF $ **FLOATING
C544 a_540371_681998.t43 vssa2 0.74fF
C545 a_540371_681998.n10 vssa2 0.56fF $ **FLOATING
C546 a_540371_681998.t32 vssa2 0.74fF
C547 a_540371_681998.n11 vssa2 0.56fF $ **FLOATING
C548 a_540371_681998.t35 vssa2 0.78fF
C549 a_540371_681998.t19 vssa2 0.74fF
C550 a_540371_681998.n12 vssa2 2.40fF $ **FLOATING
C551 a_540371_681998.n13 vssa2 1.29fF $ **FLOATING
C552 a_540371_681998.n14 vssa2 0.83fF $ **FLOATING
C553 a_540371_681998.t6 vssa2 0.05fF
C554 a_540371_681998.n15 vssa2 0.47fF $ **FLOATING
C555 a_540371_681998.n16 vssa2 1.09fF $ **FLOATING
C556 a_540371_681998.t11 vssa2 0.02fF
C557 a_540371_681998.n17 vssa2 0.75fF $ **FLOATING
C558 a_540371_681998.t10 vssa2 0.24fF
C559 a_540371_681998.t12 vssa2 0.24fF
C560 a_540371_681998.t13 vssa2 0.02fF
C561 a_540371_681998.t0 vssa2 0.10fF
C562 a_540371_681998.t4 vssa2 0.38fF
C563 a_540371_681998.n18 vssa2 2.31fF $ **FLOATING
C564 a_540371_681998.t3 vssa2 0.10fF
C565 a_540371_681998.n19 vssa2 0.83fF $ **FLOATING
C566 a_540371_681998.t15 vssa2 0.02fF
C567 a_540371_681998.n20 vssa2 0.78fF $ **FLOATING
C568 a_540371_681998.t14 vssa2 0.24fF
C569 a_540371_681998.t44 vssa2 0.78fF
C570 a_540371_681998.t26 vssa2 0.74fF
C571 a_540371_681998.n21 vssa2 2.40fF $ **FLOATING
C572 a_540371_681998.n22 vssa2 1.29fF $ **FLOATING
C573 a_540371_681998.n23 vssa2 0.81fF $ **FLOATING
C574 a_540371_681998.t7 vssa2 0.05fF
C575 a_540371_681998.n24 vssa2 0.47fF $ **FLOATING
C576 a_540371_681998.n25 vssa2 1.11fF $ **FLOATING
C577 a_540371_681998.t21 vssa2 0.78fF
C578 a_540371_681998.t40 vssa2 0.74fF
C579 a_540371_681998.n26 vssa2 2.88fF $ **FLOATING
C580 a_540371_681998.n27 vssa2 1.49fF $ **FLOATING
C581 a_540371_681998.t24 vssa2 0.74fF
C582 a_540371_681998.t27 vssa2 0.74fF
C583 a_540371_681998.n28 vssa2 1.48fF $ **FLOATING
C584 a_540371_681998.t41 vssa2 0.74fF
C585 a_540371_681998.n29 vssa2 0.30fF $ **FLOATING
C586 a_540371_681998.n30 vssa2 1.48fF $ **FLOATING
C587 a_540371_681998.n31 vssa2 0.65fF $ **FLOATING
C588 a_540371_681998.t45 vssa2 0.75fF
C589 a_540371_681998.n32 vssa2 3.18fF $ **FLOATING
C590 a_540371_681998.t29 vssa2 0.74fF
C591 a_540371_681998.n33 vssa2 0.28fF $ **FLOATING
C592 a_540371_681998.n34 vssa2 1.49fF $ **FLOATING
C593 a_540371_681998.n35 vssa2 0.60fF $ **FLOATING
C594 a_540371_681998.t20 vssa2 0.74fF
C595 a_540371_681998.t46 vssa2 0.76fF
C596 a_540371_681998.n36 vssa2 2.55fF $ **FLOATING
C597 a_540371_681998.n37 vssa2 0.65fF $ **FLOATING
C598 a_540371_681998.n38 vssa2 0.60fF $ **FLOATING
C599 a_540371_681998.n39 vssa2 1.48fF $ **FLOATING
C600 a_540371_681998.t33 vssa2 0.74fF
C601 a_540371_681998.n40 vssa2 0.29fF $ **FLOATING
C602 a_540371_681998.t16 vssa2 0.74fF
C603 a_540371_681998.t31 vssa2 0.76fF
C604 a_540371_681998.n41 vssa2 2.49fF $ **FLOATING
C605 a_540371_681998.n42 vssa2 1.34fF $ **FLOATING
C606 a_540371_681998.t18 vssa2 0.74fF
C607 a_540371_681998.n43 vssa2 1.48fF $ **FLOATING
C608 a_540371_681998.t47 vssa2 0.74fF
C609 a_540371_681998.n44 vssa2 0.30fF $ **FLOATING
C610 a_540371_681998.t28 vssa2 0.74fF
C611 a_540371_681998.n45 vssa2 1.44fF $ **FLOATING
C612 a_540371_681998.t22 vssa2 0.74fF
C613 a_540371_681998.n46 vssa2 1.45fF $ **FLOATING
C614 a_540371_681998.t37 vssa2 0.74fF
C615 a_540371_681998.n47 vssa2 0.30fF $ **FLOATING
C616 a_540371_681998.n48 vssa2 1.48fF $ **FLOATING
C617 a_540371_681998.n49 vssa2 1.32fF $ **FLOATING
C618 a_540371_681998.t23 vssa2 0.74fF
C619 a_540371_681998.t17 vssa2 0.74fF
C620 a_540371_681998.t36 vssa2 0.75fF
C621 a_540371_681998.n50 vssa2 3.11fF $ **FLOATING
C622 a_540371_681998.t39 vssa2 0.76fF
C623 a_540371_681998.n51 vssa2 2.53fF $ **FLOATING
C624 a_540371_681998.n52 vssa2 1.34fF $ **FLOATING
C625 a_540371_681998.t34 vssa2 0.76fF
C626 a_540371_681998.n53 vssa2 2.52fF $ **FLOATING
C627 a_540371_681998.n54 vssa2 0.99fF $ **FLOATING
C628 a_540371_681998.n55 vssa2 1.45fF $ **FLOATING
C629 a_540371_681998.t30 vssa2 0.74fF
C630 a_540371_681998.n56 vssa2 0.30fF $ **FLOATING
C631 a_540371_681998.n57 vssa2 1.43fF $ **FLOATING
C632 a_540371_681998.t25 vssa2 0.76fF
C633 a_540371_681998.n58 vssa2 2.49fF $ **FLOATING
C634 a_540371_681998.n59 vssa2 0.99fF $ **FLOATING
C635 a_540371_681998.t42 vssa2 0.74fF
C636 a_540371_681998.n60 vssa2 1.48fF $ **FLOATING
C637 a_540371_681998.t38 vssa2 0.74fF
C638 a_540371_681998.n61 vssa2 0.30fF $ **FLOATING
C639 a_540371_681998.n62 vssa2 1.44fF $ **FLOATING
C640 a_540371_681998.n63 vssa2 4.08fF $ **FLOATING
C641 a_540371_681998.t9 vssa2 0.02fF
C642 a_540371_681998.t8 vssa2 0.24fF
C643 a_540371_681998.t1 vssa2 0.10fF
C644 a_540371_681998.n64 vssa2 0.83fF $ **FLOATING
C645 a_540371_681998.t2 vssa2 0.38fF
C646 a_540371_681998.n65 vssa2 2.32fF $ **FLOATING
C647 a_540371_681998.t5 vssa2 0.10fF
C648 a_540371_681998.n66 vssa2 0.02fF $ **FLOATING
C649 a_540916_680434.n0 vssa2 2.92fF $ **FLOATING
C650 a_540916_680434.t13 vssa2 0.08fF
C651 a_540916_680434.t24 vssa2 0.65fF
C652 a_540916_680434.n1 vssa2 0.81fF $ **FLOATING
C653 a_540916_680434.t26 vssa2 0.65fF
C654 a_540916_680434.n2 vssa2 0.81fF $ **FLOATING
C655 a_540916_680434.t22 vssa2 0.65fF
C656 a_540916_680434.n3 vssa2 1.04fF $ **FLOATING
C657 a_540916_680434.t5 vssa2 0.04fF
C658 a_540916_680434.t7 vssa2 0.04fF
C659 a_540916_680434.n4 vssa2 0.71fF $ **FLOATING
C660 a_540916_680434.n5 vssa2 0.54fF $ **FLOATING
C661 a_540916_680434.t6 vssa2 0.18fF
C662 a_540916_680434.n6 vssa2 0.34fF $ **FLOATING
C663 a_540916_680434.n7 vssa2 0.34fF $ **FLOATING
C664 a_540916_680434.n8 vssa2 0.54fF $ **FLOATING
C665 a_540916_680434.t4 vssa2 0.18fF
C666 a_540916_680434.n9 vssa2 0.70fF $ **FLOATING
C667 a_540916_680434.t3 vssa2 0.08fF
C668 a_540916_680434.t1 vssa2 0.43fF
C669 a_540916_680434.n10 vssa2 1.41fF $ **FLOATING
C670 a_540916_680434.t2 vssa2 0.08fF
C671 a_540916_680434.t21 vssa2 0.08fF
C672 a_540916_680434.n11 vssa2 1.00fF $ **FLOATING
C673 a_540916_680434.n12 vssa2 1.00fF $ **FLOATING
C674 a_540916_680434.n13 vssa2 0.94fF $ **FLOATING
C675 a_540916_680434.n14 vssa2 2.55fF $ **FLOATING
C676 a_540916_680434.t25 vssa2 0.66fF
C677 a_540916_680434.n15 vssa2 1.97fF $ **FLOATING
C678 a_540916_680434.n16 vssa2 2.12fF $ **FLOATING
C679 a_540916_680434.t17 vssa2 0.08fF
C680 a_540916_680434.t9 vssa2 0.08fF
C681 a_540916_680434.t0 vssa2 0.08fF
C682 a_540916_680434.t20 vssa2 0.43fF
C683 a_540916_680434.n17 vssa2 1.39fF $ **FLOATING
C684 a_540916_680434.n18 vssa2 0.03fF $ **FLOATING
C685 a_540916_680434.n19 vssa2 0.06fF $ **FLOATING
C686 a_540916_680434.t27 vssa2 0.65fF
C687 a_540916_680434.n20 vssa2 1.05fF $ **FLOATING
C688 a_540916_680434.t23 vssa2 0.66fF
C689 a_540916_680434.n21 vssa2 1.96fF $ **FLOATING
C690 a_540916_680434.n22 vssa2 2.93fF $ **FLOATING
C691 a_540916_680434.t15 vssa2 0.08fF
C692 a_540916_680434.t11 vssa2 0.14fF
C693 a_540916_680434.t10 vssa2 0.66fF
C694 a_540916_680434.n23 vssa2 2.10fF $ **FLOATING
C695 a_540916_680434.n24 vssa2 1.39fF $ **FLOATING
C696 a_540916_680434.n25 vssa2 0.87fF $ **FLOATING
C697 a_540916_680434.n26 vssa2 1.18fF $ **FLOATING
C698 a_540916_680434.t14 vssa2 0.65fF
C699 a_540916_680434.n27 vssa2 0.58fF $ **FLOATING
C700 a_540916_680434.n28 vssa2 0.80fF $ **FLOATING
C701 a_540916_680434.n29 vssa2 1.14fF $ **FLOATING
C702 a_540916_680434.t8 vssa2 0.65fF
C703 a_540916_680434.n30 vssa2 0.80fF $ **FLOATING
C704 a_540916_680434.n31 vssa2 0.80fF $ **FLOATING
C705 a_540916_680434.n32 vssa2 1.14fF $ **FLOATING
C706 a_540916_680434.t16 vssa2 0.65fF
C707 a_540916_680434.n33 vssa2 0.80fF $ **FLOATING
C708 a_540916_680434.n34 vssa2 0.56fF $ **FLOATING
C709 a_540916_680434.n35 vssa2 1.11fF $ **FLOATING
C710 a_540916_680434.n36 vssa2 0.90fF $ **FLOATING
C711 a_540916_680434.t12 vssa2 0.65fF
C712 a_540916_680434.n37 vssa2 1.39fF $ **FLOATING
C713 a_540916_680434.t18 vssa2 0.66fF
C714 a_540916_680434.n38 vssa2 2.07fF $ **FLOATING
C715 a_540916_680434.t19 vssa2 0.14fF
C716 a_534722_685355.t7 vssa2 0.28fF
C717 a_534722_685355.t2 vssa2 19.73fF
C718 a_534722_685355.t1 vssa2 19.73fF
C719 a_534722_685355.t3 vssa2 19.73fF
C720 a_534722_685355.t0 vssa2 19.73fF
C721 a_534722_685355.t5 vssa2 0.28fF
C722 a_534722_685355.t6 vssa2 0.73fF
C723 a_534722_685355.n0 vssa2 11.89fF $ **FLOATING
C724 a_534722_685355.n1 vssa2 12.23fF $ **FLOATING
C725 a_534722_685355.n2 vssa2 9.15fF $ **FLOATING
C726 a_534722_685355.n3 vssa2 9.15fF $ **FLOATING
C727 a_534722_685355.n4 vssa2 12.15fF $ **FLOATING
C728 a_534722_685355.n5 vssa2 9.95fF $ **FLOATING
C729 a_534722_685355.t4 vssa2 2.90fF
C730 a_42818_684860.t10 vssa2 0.07fF
C731 a_42818_684860.t5 vssa2 0.07fF
C732 a_42818_684860.n0 vssa2 0.38fF $ **FLOATING
C733 a_42818_684860.n1 vssa2 0.91fF $ **FLOATING
C734 a_42818_684860.t6 vssa2 0.07fF
C735 a_42818_684860.t12 vssa2 0.07fF
C736 a_42818_684860.n2 vssa2 0.38fF $ **FLOATING
C737 a_42818_684860.n3 vssa2 0.92fF $ **FLOATING
C738 a_42818_684860.t24 vssa2 0.07fF
C739 a_42818_684860.t26 vssa2 0.07fF
C740 a_42818_684860.n4 vssa2 0.38fF $ **FLOATING
C741 a_42818_684860.n5 vssa2 0.91fF $ **FLOATING
C742 a_42818_684860.t1 vssa2 0.14fF
C743 a_42818_684860.n6 vssa2 2.18fF $ **FLOATING
C744 a_42818_684860.t23 vssa2 0.07fF
C745 a_42818_684860.t11 vssa2 0.07fF
C746 a_42818_684860.n7 vssa2 0.36fF $ **FLOATING
C747 a_42818_684860.n8 vssa2 0.85fF $ **FLOATING
C748 a_42818_684860.t8 vssa2 0.11fF
C749 a_42818_684860.n9 vssa2 3.50fF $ **FLOATING
C750 a_42818_684860.n10 vssa2 3.33fF $ **FLOATING
C751 a_42818_684860.t17 vssa2 0.07fF
C752 a_42818_684860.t14 vssa2 0.07fF
C753 a_42818_684860.n11 vssa2 0.36fF $ **FLOATING
C754 a_42818_684860.n12 vssa2 1.83fF $ **FLOATING
C755 a_42818_684860.t27 vssa2 0.07fF
C756 a_42818_684860.t7 vssa2 0.07fF
C757 a_42818_684860.n13 vssa2 0.38fF $ **FLOATING
C758 a_42818_684860.n14 vssa2 0.91fF $ **FLOATING
C759 a_42818_684860.t2 vssa2 0.07fF
C760 a_42818_684860.t9 vssa2 0.07fF
C761 a_42818_684860.n15 vssa2 0.38fF $ **FLOATING
C762 a_42818_684860.n16 vssa2 0.91fF $ **FLOATING
C763 a_42818_684860.t25 vssa2 0.07fF
C764 a_42818_684860.t4 vssa2 0.07fF
C765 a_42818_684860.n17 vssa2 0.38fF $ **FLOATING
C766 a_42818_684860.n18 vssa2 0.91fF $ **FLOATING
C767 a_42818_684860.t3 vssa2 0.14fF
C768 a_42818_684860.n19 vssa2 2.18fF $ **FLOATING
C769 a_42818_684860.t0 vssa2 0.07fF
C770 a_42818_684860.t13 vssa2 0.07fF
C771 a_42818_684860.n20 vssa2 0.36fF $ **FLOATING
C772 a_42818_684860.n21 vssa2 0.84fF $ **FLOATING
C773 a_42818_684860.t22 vssa2 0.07fF
C774 a_42818_684860.t21 vssa2 0.07fF
C775 a_42818_684860.n22 vssa2 0.36fF $ **FLOATING
C776 a_42818_684860.n23 vssa2 3.32fF $ **FLOATING
C777 a_42818_684860.n24 vssa2 3.25fF $ **FLOATING
C778 a_42818_684860.t16 vssa2 0.11fF
C779 a_42818_684860.n25 vssa2 2.08fF $ **FLOATING
C780 a_42818_684860.t18 vssa2 0.07fF
C781 a_42818_684860.t19 vssa2 0.07fF
C782 a_42818_684860.n26 vssa2 0.36fF $ **FLOATING
C783 a_42818_684860.n27 vssa2 0.84fF $ **FLOATING
C784 a_42818_684860.n28 vssa2 0.84fF $ **FLOATING
C785 a_42818_684860.t15 vssa2 0.07fF
C786 a_42818_684860.n29 vssa2 0.36fF $ **FLOATING
C787 a_42818_684860.t20 vssa2 0.07fF
C788 a_43026_690892.n0 vssa2 0.71fF $ **FLOATING
C789 a_43026_690892.n1 vssa2 0.74fF $ **FLOATING
C790 a_43026_690892.n2 vssa2 2.79fF $ **FLOATING
C791 a_43026_690892.n3 vssa2 2.56fF $ **FLOATING
C792 a_43026_690892.n4 vssa2 0.35fF $ **FLOATING
C793 a_43026_690892.n5 vssa2 0.34fF $ **FLOATING
C794 a_43026_690892.n6 vssa2 0.35fF $ **FLOATING
C795 a_43026_690892.n7 vssa2 0.35fF $ **FLOATING
C796 a_43026_690892.t37 vssa2 0.07fF
C797 a_43026_690892.t1 vssa2 0.07fF
C798 a_43026_690892.n8 vssa2 0.46fF $ **FLOATING
C799 a_43026_690892.t9 vssa2 0.07fF
C800 a_43026_690892.t13 vssa2 0.07fF
C801 a_43026_690892.t67 vssa2 0.28fF
C802 a_43026_690892.n9 vssa2 0.21fF $ **FLOATING
C803 a_43026_690892.t68 vssa2 0.28fF
C804 a_43026_690892.n10 vssa2 0.21fF $ **FLOATING
C805 a_43026_690892.t54 vssa2 0.28fF
C806 a_43026_690892.n11 vssa2 0.21fF $ **FLOATING
C807 a_43026_690892.t63 vssa2 0.28fF
C808 a_43026_690892.n12 vssa2 0.21fF $ **FLOATING
C809 a_43026_690892.t65 vssa2 0.28fF
C810 a_43026_690892.n13 vssa2 0.21fF $ **FLOATING
C811 a_43026_690892.t69 vssa2 0.28fF
C812 a_43026_690892.n14 vssa2 0.21fF $ **FLOATING
C813 a_43026_690892.n15 vssa2 0.21fF $ **FLOATING
C814 a_43026_690892.n16 vssa2 0.21fF $ **FLOATING
C815 a_43026_690892.n17 vssa2 0.21fF $ **FLOATING
C816 a_43026_690892.n18 vssa2 0.21fF $ **FLOATING
C817 a_43026_690892.n19 vssa2 0.21fF $ **FLOATING
C818 a_43026_690892.n20 vssa2 0.21fF $ **FLOATING
C819 a_43026_690892.n21 vssa2 0.21fF $ **FLOATING
C820 a_43026_690892.n22 vssa2 0.56fF $ **FLOATING
C821 a_43026_690892.t51 vssa2 0.28fF
C822 a_43026_690892.n23 vssa2 0.11fF $ **FLOATING
C823 a_43026_690892.n24 vssa2 0.95fF $ **FLOATING
C824 a_43026_690892.n25 vssa2 0.67fF $ **FLOATING
C825 a_43026_690892.n26 vssa2 0.19fF $ **FLOATING
C826 a_43026_690892.n27 vssa2 0.20fF $ **FLOATING
C827 a_43026_690892.n28 vssa2 0.12fF $ **FLOATING
C828 a_43026_690892.t8 vssa2 0.28fF
C829 a_43026_690892.t0 vssa2 0.28fF
C830 a_43026_690892.t36 vssa2 0.28fF
C831 a_43026_690892.n29 vssa2 0.42fF $ **FLOATING
C832 a_43026_690892.n30 vssa2 0.20fF $ **FLOATING
C833 a_43026_690892.t12 vssa2 0.28fF
C834 a_43026_690892.n31 vssa2 0.20fF $ **FLOATING
C835 a_43026_690892.n32 vssa2 0.04fF $ **FLOATING
C836 a_43026_690892.t43 vssa2 0.07fF
C837 a_43026_690892.t47 vssa2 0.07fF
C838 a_43026_690892.n33 vssa2 0.37fF $ **FLOATING
C839 a_43026_690892.n34 vssa2 3.23fF $ **FLOATING
C840 a_43026_690892.t30 vssa2 0.28fF
C841 a_43026_690892.n35 vssa2 0.20fF $ **FLOATING
C842 a_43026_690892.t22 vssa2 0.28fF
C843 a_43026_690892.n36 vssa2 0.21fF $ **FLOATING
C844 a_43026_690892.t16 vssa2 0.28fF
C845 a_43026_690892.n37 vssa2 0.21fF $ **FLOATING
C846 a_43026_690892.t38 vssa2 0.28fF
C847 a_43026_690892.n38 vssa2 0.21fF $ **FLOATING
C848 a_43026_690892.t32 vssa2 0.28fF
C849 a_43026_690892.n39 vssa2 0.21fF $ **FLOATING
C850 a_43026_690892.t4 vssa2 0.28fF
C851 a_43026_690892.n40 vssa2 0.21fF $ **FLOATING
C852 a_43026_690892.t2 vssa2 0.28fF
C853 a_43026_690892.n41 vssa2 0.20fF $ **FLOATING
C854 a_43026_690892.n42 vssa2 0.04fF $ **FLOATING
C855 a_43026_690892.t31 vssa2 0.07fF
C856 a_43026_690892.t3 vssa2 0.07fF
C857 a_43026_690892.n43 vssa2 0.20fF $ **FLOATING
C858 a_43026_690892.t61 vssa2 0.28fF
C859 a_43026_690892.t50 vssa2 0.28fF
C860 a_43026_690892.t53 vssa2 0.28fF
C861 a_43026_690892.n44 vssa2 0.21fF $ **FLOATING
C862 a_43026_690892.n45 vssa2 0.21fF $ **FLOATING
C863 a_43026_690892.n46 vssa2 0.20fF $ **FLOATING
C864 a_43026_690892.t49 vssa2 0.28fF
C865 a_43026_690892.n47 vssa2 0.21fF $ **FLOATING
C866 a_43026_690892.t56 vssa2 0.28fF
C867 a_43026_690892.n48 vssa2 0.20fF $ **FLOATING
C868 a_43026_690892.t58 vssa2 0.28fF
C869 a_43026_690892.n49 vssa2 0.49fF $ **FLOATING
C870 a_43026_690892.n50 vssa2 0.20fF $ **FLOATING
C871 a_43026_690892.n51 vssa2 0.49fF $ **FLOATING
C872 a_43026_690892.n52 vssa2 0.20fF $ **FLOATING
C873 a_43026_690892.n53 vssa2 0.21fF $ **FLOATING
C874 a_43026_690892.n54 vssa2 0.21fF $ **FLOATING
C875 a_43026_690892.n55 vssa2 0.21fF $ **FLOATING
C876 a_43026_690892.n56 vssa2 0.20fF $ **FLOATING
C877 a_43026_690892.n57 vssa2 0.12fF $ **FLOATING
C878 a_43026_690892.t5 vssa2 0.07fF
C879 a_43026_690892.t33 vssa2 0.07fF
C880 a_43026_690892.n58 vssa2 0.39fF $ **FLOATING
C881 a_43026_690892.n59 vssa2 0.73fF $ **FLOATING
C882 a_43026_690892.t39 vssa2 0.07fF
C883 a_43026_690892.t17 vssa2 0.07fF
C884 a_43026_690892.n60 vssa2 0.39fF $ **FLOATING
C885 a_43026_690892.n61 vssa2 0.73fF $ **FLOATING
C886 a_43026_690892.t23 vssa2 0.07fF
C887 a_43026_690892.t27 vssa2 0.07fF
C888 a_43026_690892.n62 vssa2 0.39fF $ **FLOATING
C889 a_43026_690892.n63 vssa2 0.74fF $ **FLOATING
C890 a_43026_690892.t35 vssa2 0.12fF
C891 a_43026_690892.t48 vssa2 0.07fF
C892 a_43026_690892.t42 vssa2 0.07fF
C893 a_43026_690892.n64 vssa2 0.37fF $ **FLOATING
C894 a_43026_690892.n65 vssa2 0.87fF $ **FLOATING
C895 a_43026_690892.t46 vssa2 0.07fF
C896 a_43026_690892.t44 vssa2 0.07fF
C897 a_43026_690892.n66 vssa2 0.37fF $ **FLOATING
C898 a_43026_690892.n67 vssa2 0.88fF $ **FLOATING
C899 a_43026_690892.t45 vssa2 0.11fF
C900 a_43026_690892.n68 vssa2 3.67fF $ **FLOATING
C901 a_43026_690892.t24 vssa2 0.28fF
C902 a_43026_690892.n69 vssa2 0.20fF $ **FLOATING
C903 a_43026_690892.t34 vssa2 0.28fF
C904 a_43026_690892.t28 vssa2 0.28fF
C905 a_43026_690892.n70 vssa2 0.41fF $ **FLOATING
C906 a_43026_690892.n71 vssa2 0.04fF $ **FLOATING
C907 a_43026_690892.t25 vssa2 0.07fF
C908 a_43026_690892.t29 vssa2 0.07fF
C909 a_43026_690892.t57 vssa2 0.28fF
C910 a_43026_690892.t59 vssa2 0.28fF
C911 a_43026_690892.t62 vssa2 0.28fF
C912 a_43026_690892.t64 vssa2 0.28fF
C913 a_43026_690892.t66 vssa2 0.28fF
C914 a_43026_690892.t60 vssa2 0.28fF
C915 a_43026_690892.n72 vssa2 0.21fF $ **FLOATING
C916 a_43026_690892.n73 vssa2 0.21fF $ **FLOATING
C917 a_43026_690892.n74 vssa2 0.21fF $ **FLOATING
C918 a_43026_690892.n75 vssa2 0.21fF $ **FLOATING
C919 a_43026_690892.n76 vssa2 0.21fF $ **FLOATING
C920 a_43026_690892.n77 vssa2 0.21fF $ **FLOATING
C921 a_43026_690892.t52 vssa2 0.28fF
C922 a_43026_690892.n78 vssa2 0.21fF $ **FLOATING
C923 a_43026_690892.n79 vssa2 0.21fF $ **FLOATING
C924 a_43026_690892.n80 vssa2 0.21fF $ **FLOATING
C925 a_43026_690892.n81 vssa2 0.21fF $ **FLOATING
C926 a_43026_690892.n82 vssa2 0.21fF $ **FLOATING
C927 a_43026_690892.n83 vssa2 0.21fF $ **FLOATING
C928 a_43026_690892.n84 vssa2 0.21fF $ **FLOATING
C929 a_43026_690892.n85 vssa2 0.21fF $ **FLOATING
C930 a_43026_690892.n86 vssa2 0.21fF $ **FLOATING
C931 a_43026_690892.n87 vssa2 0.56fF $ **FLOATING
C932 a_43026_690892.n88 vssa2 0.11fF $ **FLOATING
C933 a_43026_690892.t55 vssa2 0.28fF
C934 a_43026_690892.n89 vssa2 0.94fF $ **FLOATING
C935 a_43026_690892.n90 vssa2 0.48fF $ **FLOATING
C936 a_43026_690892.n91 vssa2 0.19fF $ **FLOATING
C937 a_43026_690892.n92 vssa2 0.20fF $ **FLOATING
C938 a_43026_690892.n93 vssa2 0.12fF $ **FLOATING
C939 a_43026_690892.t14 vssa2 0.28fF
C940 a_43026_690892.t10 vssa2 0.28fF
C941 a_43026_690892.t6 vssa2 0.28fF
C942 a_43026_690892.t18 vssa2 0.28fF
C943 a_43026_690892.t40 vssa2 0.28fF
C944 a_43026_690892.t26 vssa2 0.28fF
C945 a_43026_690892.n94 vssa2 0.21fF $ **FLOATING
C946 a_43026_690892.n95 vssa2 0.21fF $ **FLOATING
C947 a_43026_690892.n96 vssa2 0.21fF $ **FLOATING
C948 a_43026_690892.n97 vssa2 0.21fF $ **FLOATING
C949 a_43026_690892.n98 vssa2 0.21fF $ **FLOATING
C950 a_43026_690892.n99 vssa2 0.20fF $ **FLOATING
C951 a_43026_690892.t20 vssa2 0.28fF
C952 a_43026_690892.n100 vssa2 0.20fF $ **FLOATING
C953 a_43026_690892.n101 vssa2 0.04fF $ **FLOATING
C954 a_43026_690892.t15 vssa2 0.07fF
C955 a_43026_690892.t21 vssa2 0.07fF
C956 a_43026_690892.n102 vssa2 0.21fF $ **FLOATING
C957 a_43026_690892.n103 vssa2 0.21fF $ **FLOATING
C958 a_43026_690892.n104 vssa2 0.21fF $ **FLOATING
C959 a_43026_690892.n105 vssa2 0.21fF $ **FLOATING
C960 a_43026_690892.n106 vssa2 0.20fF $ **FLOATING
C961 a_43026_690892.n107 vssa2 0.20fF $ **FLOATING
C962 a_43026_690892.n108 vssa2 0.12fF $ **FLOATING
C963 a_43026_690892.n109 vssa2 0.03fF $ **FLOATING
C964 a_43026_690892.t7 vssa2 0.07fF
C965 a_43026_690892.t11 vssa2 0.07fF
C966 a_43026_690892.n110 vssa2 0.39fF $ **FLOATING
C967 a_43026_690892.n111 vssa2 0.73fF $ **FLOATING
C968 a_43026_690892.n112 vssa2 0.73fF $ **FLOATING
C969 a_43026_690892.t19 vssa2 0.07fF
C970 a_43026_690892.n113 vssa2 0.39fF $ **FLOATING
C971 a_43026_690892.t41 vssa2 0.07fF
C972 io_analog[9].t6 vssa2 0.03fF
C973 io_analog[9].n0 vssa2 0.02fF $ **FLOATING
C974 io_analog[9].n1 vssa2 0.06fF $ **FLOATING
C975 io_analog[9].n2 vssa2 0.02fF $ **FLOATING
C976 io_analog[9].t0 vssa2 0.03fF
C977 io_analog[9].n3 vssa2 0.02fF $ **FLOATING
C978 io_analog[9].t1 vssa2 0.03fF
C979 io_analog[9].n4 vssa2 0.02fF $ **FLOATING
C980 io_analog[9].t2 vssa2 0.03fF
C981 io_analog[9].n5 vssa2 0.02fF $ **FLOATING
C982 io_analog[9].t4 vssa2 0.03fF
C983 io_analog[9].n6 vssa2 0.03fF $ **FLOATING
C984 io_analog[9].t3 vssa2 0.03fF
C985 io_analog[9].n7 vssa2 0.06fF $ **FLOATING
C986 io_analog[9].t5 vssa2 0.03fF
C987 io_analog[9].n8 vssa2 0.02fF $ **FLOATING
C988 io_analog[9].n9 vssa2 0.02fF $ **FLOATING
C989 io_analog[9].n10 vssa2 0.02fF $ **FLOATING
C990 io_analog[9].n11 vssa2 0.02fF $ **FLOATING
C991 io_analog[9].n12 vssa2 0.03fF $ **FLOATING
C992 io_analog[9].n13 vssa2 3.30fF $ **FLOATING
C993 io_analog[10].t33 vssa2 0.01fF
C994 io_analog[10].t38 vssa2 0.01fF
C995 io_analog[10].n0 vssa2 0.06fF $ **FLOATING
C996 io_analog[10].n1 vssa2 0.13fF $ **FLOATING
C997 io_analog[10].t46 vssa2 0.01fF
C998 io_analog[10].t19 vssa2 0.01fF
C999 io_analog[10].n2 vssa2 0.06fF $ **FLOATING
C1000 io_analog[10].n3 vssa2 0.18fF $ **FLOATING
C1001 io_analog[10].n4 vssa2 1.04fF $ **FLOATING
C1002 io_analog[10].t7 vssa2 0.02fF
C1003 io_analog[10].n5 vssa2 1.08fF $ **FLOATING
C1004 io_analog[10].t5 vssa2 0.01fF
C1005 io_analog[10].t4 vssa2 0.01fF
C1006 io_analog[10].n6 vssa2 0.06fF $ **FLOATING
C1007 io_analog[10].n7 vssa2 0.21fF $ **FLOATING
C1008 io_analog[10].t9 vssa2 0.01fF
C1009 io_analog[10].t50 vssa2 0.01fF
C1010 io_analog[10].n8 vssa2 0.06fF $ **FLOATING
C1011 io_analog[10].n9 vssa2 0.21fF $ **FLOATING
C1012 io_analog[10].t1 vssa2 0.01fF
C1013 io_analog[10].t0 vssa2 0.01fF
C1014 io_analog[10].n10 vssa2 0.06fF $ **FLOATING
C1015 io_analog[10].n11 vssa2 0.21fF $ **FLOATING
C1016 io_analog[10].t8 vssa2 0.01fF
C1017 io_analog[10].t3 vssa2 0.01fF
C1018 io_analog[10].n12 vssa2 0.06fF $ **FLOATING
C1019 io_analog[10].n13 vssa2 0.21fF $ **FLOATING
C1020 io_analog[10].t2 vssa2 0.01fF
C1021 io_analog[10].t6 vssa2 0.01fF
C1022 io_analog[10].n14 vssa2 0.06fF $ **FLOATING
C1023 io_analog[10].n15 vssa2 0.21fF $ **FLOATING
C1024 io_analog[10].t51 vssa2 0.02fF
C1025 io_analog[10].n16 vssa2 0.43fF $ **FLOATING
C1026 io_analog[10].t35 vssa2 0.01fF
C1027 io_analog[10].t23 vssa2 0.01fF
C1028 io_analog[10].n17 vssa2 0.06fF $ **FLOATING
C1029 io_analog[10].n18 vssa2 0.13fF $ **FLOATING
C1030 io_analog[10].t10 vssa2 0.01fF
C1031 io_analog[10].t17 vssa2 0.01fF
C1032 io_analog[10].n19 vssa2 0.06fF $ **FLOATING
C1033 io_analog[10].n20 vssa2 0.13fF $ **FLOATING
C1034 io_analog[10].t40 vssa2 0.01fF
C1035 io_analog[10].t48 vssa2 0.01fF
C1036 io_analog[10].n21 vssa2 0.06fF $ **FLOATING
C1037 io_analog[10].n22 vssa2 0.13fF $ **FLOATING
C1038 io_analog[10].t32 vssa2 0.01fF
C1039 io_analog[10].t36 vssa2 0.01fF
C1040 io_analog[10].n23 vssa2 0.06fF $ **FLOATING
C1041 io_analog[10].n24 vssa2 0.13fF $ **FLOATING
C1042 io_analog[10].t18 vssa2 0.01fF
C1043 io_analog[10].t21 vssa2 0.01fF
C1044 io_analog[10].n25 vssa2 0.06fF $ **FLOATING
C1045 io_analog[10].n26 vssa2 0.13fF $ **FLOATING
C1046 io_analog[10].t49 vssa2 0.01fF
C1047 io_analog[10].t13 vssa2 0.01fF
C1048 io_analog[10].n27 vssa2 0.06fF $ **FLOATING
C1049 io_analog[10].n28 vssa2 0.13fF $ **FLOATING
C1050 io_analog[10].t22 vssa2 0.01fF
C1051 io_analog[10].t26 vssa2 0.01fF
C1052 io_analog[10].n29 vssa2 0.06fF $ **FLOATING
C1053 io_analog[10].n30 vssa2 0.13fF $ **FLOATING
C1054 io_analog[10].t25 vssa2 0.01fF
C1055 io_analog[10].t34 vssa2 0.01fF
C1056 io_analog[10].n31 vssa2 0.06fF $ **FLOATING
C1057 io_analog[10].n32 vssa2 0.13fF $ **FLOATING
C1058 io_analog[10].t44 vssa2 0.01fF
C1059 io_analog[10].t20 vssa2 0.01fF
C1060 io_analog[10].n33 vssa2 0.06fF $ **FLOATING
C1061 io_analog[10].n34 vssa2 0.13fF $ **FLOATING
C1062 io_analog[10].t30 vssa2 0.01fF
C1063 io_analog[10].t39 vssa2 0.01fF
C1064 io_analog[10].n35 vssa2 0.06fF $ **FLOATING
C1065 io_analog[10].n36 vssa2 0.13fF $ **FLOATING
C1066 io_analog[10].t37 vssa2 0.01fF
C1067 io_analog[10].t42 vssa2 0.01fF
C1068 io_analog[10].n37 vssa2 0.06fF $ **FLOATING
C1069 io_analog[10].n38 vssa2 0.13fF $ **FLOATING
C1070 io_analog[10].t12 vssa2 0.01fF
C1071 io_analog[10].t15 vssa2 0.01fF
C1072 io_analog[10].n39 vssa2 0.06fF $ **FLOATING
C1073 io_analog[10].n40 vssa2 0.13fF $ **FLOATING
C1074 io_analog[10].t43 vssa2 0.01fF
C1075 io_analog[10].t45 vssa2 0.01fF
C1076 io_analog[10].n41 vssa2 0.06fF $ **FLOATING
C1077 io_analog[10].n42 vssa2 0.13fF $ **FLOATING
C1078 io_analog[10].t28 vssa2 0.01fF
C1079 io_analog[10].t11 vssa2 0.01fF
C1080 io_analog[10].n43 vssa2 0.06fF $ **FLOATING
C1081 io_analog[10].n44 vssa2 0.13fF $ **FLOATING
C1082 io_analog[10].t16 vssa2 0.01fF
C1083 io_analog[10].t24 vssa2 0.01fF
C1084 io_analog[10].n45 vssa2 0.06fF $ **FLOATING
C1085 io_analog[10].n46 vssa2 0.13fF $ **FLOATING
C1086 io_analog[10].t47 vssa2 0.01fF
C1087 io_analog[10].t14 vssa2 0.01fF
C1088 io_analog[10].n47 vssa2 0.06fF $ **FLOATING
C1089 io_analog[10].n48 vssa2 0.13fF $ **FLOATING
C1090 io_analog[10].t41 vssa2 0.01fF
C1091 io_analog[10].t29 vssa2 0.01fF
C1092 io_analog[10].n49 vssa2 0.06fF $ **FLOATING
C1093 io_analog[10].n50 vssa2 0.13fF $ **FLOATING
C1094 io_analog[10].t27 vssa2 0.01fF
C1095 io_analog[10].t31 vssa2 0.01fF
C1096 io_analog[10].n51 vssa2 0.06fF $ **FLOATING
C1097 io_analog[10].n52 vssa2 0.18fF $ **FLOATING
C1098 io_analog[10].t54 vssa2 15.79fF
C1099 io_analog[10].n53 vssa2 2.40fF $ **FLOATING
C1100 io_analog[10].t53 vssa2 15.92fF
C1101 io_analog[10].t55 vssa2 15.91fF
C1102 io_analog[10].t52 vssa2 15.81fF
C1103 io_analog[10].n54 vssa2 2.39fF $ **FLOATING
C1104 io_analog[10].n55 vssa2 1.02fF $ **FLOATING
C1105 io_analog[10].n56 vssa2 41.75fF $ **FLOATING
C1106 vccd2.t27 vssa2 0.01fF
C1107 vccd2.n0 vssa2 0.00fF $ **FLOATING
C1108 vccd2.n1 vssa2 0.00fF $ **FLOATING
C1109 vccd2.n2 vssa2 0.01fF $ **FLOATING
C1110 vccd2.n3 vssa2 0.02fF $ **FLOATING
C1111 vccd2.n5 vssa2 0.00fF $ **FLOATING
C1112 vccd2.n6 vssa2 0.00fF $ **FLOATING
C1113 vccd2.n7 vssa2 0.03fF $ **FLOATING
C1114 vccd2.n8 vssa2 0.00fF $ **FLOATING
C1115 vccd2.n10 vssa2 0.01fF $ **FLOATING
C1116 vccd2.n11 vssa2 0.01fF $ **FLOATING
C1117 vccd2.t16 vssa2 0.32fF
C1118 vccd2.t14 vssa2 0.43fF
C1119 vccd2.t26 vssa2 0.42fF
C1120 vccd2.n12 vssa2 0.01fF $ **FLOATING
C1121 vccd2.n13 vssa2 0.02fF $ **FLOATING
C1122 vccd2.n14 vssa2 0.30fF $ **FLOATING
C1123 vccd2.n15 vssa2 0.01fF $ **FLOATING
C1124 vccd2.n16 vssa2 0.02fF $ **FLOATING
C1125 vccd2.n18 vssa2 0.00fF $ **FLOATING
C1126 vccd2.n19 vssa2 0.03fF $ **FLOATING
C1127 vccd2.n20 vssa2 0.04fF $ **FLOATING
C1128 vccd2.t155 vssa2 0.01fF
C1129 vccd2.t17 vssa2 0.01fF
C1130 vccd2.t15 vssa2 0.01fF
C1131 vccd2.n21 vssa2 0.05fF $ **FLOATING
C1132 vccd2.n22 vssa2 0.06fF $ **FLOATING
C1133 vccd2.n23 vssa2 0.11fF $ **FLOATING
C1134 vccd2.n24 vssa2 549.95fF $ **FLOATING
C1135 vccd2.t160 vssa2 0.01fF
C1136 vccd2.t29 vssa2 0.01fF
C1137 vccd2.n25 vssa2 0.04fF $ **FLOATING
C1138 vccd2.t31 vssa2 0.01fF
C1139 vccd2.t46 vssa2 0.01fF
C1140 vccd2.n26 vssa2 0.04fF $ **FLOATING
C1141 vccd2.t152 vssa2 0.01fF
C1142 vccd2.t23 vssa2 0.01fF
C1143 vccd2.n27 vssa2 0.04fF $ **FLOATING
C1144 vccd2.n28 vssa2 0.08fF $ **FLOATING
C1145 vccd2.t18 vssa2 0.01fF
C1146 vccd2.t149 vssa2 0.01fF
C1147 vccd2.n29 vssa2 0.04fF $ **FLOATING
C1148 vccd2.n30 vssa2 0.08fF $ **FLOATING
C1149 vccd2.n31 vssa2 0.07fF $ **FLOATING
C1150 vccd2.n32 vssa2 0.01fF $ **FLOATING
C1151 vccd2.n33 vssa2 0.01fF $ **FLOATING
C1152 vccd2.n34 vssa2 0.02fF $ **FLOATING
C1153 vccd2.n35 vssa2 0.04fF $ **FLOATING
C1154 vccd2.n36 vssa2 0.04fF $ **FLOATING
C1155 vccd2.n37 vssa2 0.03fF $ **FLOATING
C1156 vccd2.n38 vssa2 0.43fF $ **FLOATING
C1157 vccd2.t93 vssa2 0.47fF
C1158 vccd2.t101 vssa2 0.43fF
C1159 vccd2.t125 vssa2 0.43fF
C1160 vccd2.t97 vssa2 0.43fF
C1161 vccd2.t133 vssa2 0.26fF
C1162 vccd2.n39 vssa2 0.03fF $ **FLOATING
C1163 vccd2.n40 vssa2 0.04fF $ **FLOATING
C1164 vccd2.n41 vssa2 0.21fF $ **FLOATING
C1165 vccd2.t67 vssa2 0.38fF
C1166 vccd2.t71 vssa2 0.43fF
C1167 vccd2.t87 vssa2 0.43fF
C1168 vccd2.t95 vssa2 0.27fF
C1169 vccd2.n42 vssa2 0.03fF $ **FLOATING
C1170 vccd2.n43 vssa2 0.03fF $ **FLOATING
C1171 vccd2.n44 vssa2 0.02fF $ **FLOATING
C1172 vccd2.n45 vssa2 0.02fF $ **FLOATING
C1173 vccd2.n46 vssa2 0.21fF $ **FLOATING
C1174 vccd2.t61 vssa2 0.26fF
C1175 vccd2.t6 vssa2 0.21fF
C1176 vccd2.t107 vssa2 0.21fF
C1177 vccd2.t146 vssa2 0.20fF
C1178 vccd2.n47 vssa2 0.01fF $ **FLOATING
C1179 vccd2.n48 vssa2 0.02fF $ **FLOATING
C1180 vccd2.n49 vssa2 0.11fF $ **FLOATING
C1181 vccd2.t129 vssa2 0.09fF
C1182 vccd2.n50 vssa2 0.02fF $ **FLOATING
C1183 vccd2.n51 vssa2 0.02fF $ **FLOATING
C1184 vccd2.n52 vssa2 0.10fF $ **FLOATING
C1185 vccd2.t12 vssa2 0.14fF
C1186 vccd2.t63 vssa2 0.21fF
C1187 vccd2.t2 vssa2 0.21fF
C1188 vccd2.t69 vssa2 0.21fF
C1189 vccd2.t43 vssa2 0.21fF
C1190 vccd2.t119 vssa2 0.21fF
C1191 vccd2.t34 vssa2 0.18fF
C1192 vccd2.t121 vssa2 0.21fF
C1193 vccd2.t41 vssa2 0.21fF
C1194 vccd2.t99 vssa2 0.21fF
C1195 vccd2.t150 vssa2 0.21fF
C1196 vccd2.t105 vssa2 0.13fF
C1197 vccd2.n53 vssa2 0.02fF $ **FLOATING
C1198 vccd2.n54 vssa2 0.01fF $ **FLOATING
C1199 vccd2.n55 vssa2 0.20fF $ **FLOATING
C1200 vccd2.n56 vssa2 0.23fF $ **FLOATING
C1201 vccd2.t19 vssa2 0.01fF
C1202 vccd2.t147 vssa2 0.01fF
C1203 vccd2.t13 vssa2 0.01fF
C1204 vccd2.n57 vssa2 0.04fF $ **FLOATING
C1205 vccd2.n58 vssa2 0.18fF $ **FLOATING
C1206 vccd2.t148 vssa2 0.01fF
C1207 vccd2.t50 vssa2 0.01fF
C1208 vccd2.n59 vssa2 0.04fF $ **FLOATING
C1209 vccd2.n60 vssa2 0.07fF $ **FLOATING
C1210 vccd2.n61 vssa2 0.15fF $ **FLOATING
C1211 vccd2.n62 vssa2 0.01fF $ **FLOATING
C1212 vccd2.t42 vssa2 0.01fF
C1213 vccd2.t58 vssa2 0.01fF
C1214 vccd2.n63 vssa2 0.04fF $ **FLOATING
C1215 vccd2.n64 vssa2 0.08fF $ **FLOATING
C1216 vccd2.t54 vssa2 0.01fF
C1217 vccd2.t157 vssa2 0.01fF
C1218 vccd2.n65 vssa2 0.04fF $ **FLOATING
C1219 vccd2.n66 vssa2 0.07fF $ **FLOATING
C1220 vccd2.n67 vssa2 0.03fF $ **FLOATING
C1221 vccd2.t5 vssa2 0.01fF
C1222 vccd2.t56 vssa2 0.01fF
C1223 vccd2.n68 vssa2 0.04fF $ **FLOATING
C1224 vccd2.n69 vssa2 0.08fF $ **FLOATING
C1225 vccd2.t53 vssa2 0.01fF
C1226 vccd2.t141 vssa2 0.01fF
C1227 vccd2.n70 vssa2 0.04fF $ **FLOATING
C1228 vccd2.n71 vssa2 0.08fF $ **FLOATING
C1229 vccd2.t49 vssa2 0.01fF
C1230 vccd2.t57 vssa2 0.01fF
C1231 vccd2.n72 vssa2 0.04fF $ **FLOATING
C1232 vccd2.n73 vssa2 0.06fF $ **FLOATING
C1233 vccd2.n74 vssa2 0.01fF $ **FLOATING
C1234 vccd2.n75 vssa2 0.00fF $ **FLOATING
C1235 vccd2.t7 vssa2 0.01fF
C1236 vccd2.t159 vssa2 0.01fF
C1237 vccd2.t140 vssa2 0.01fF
C1238 vccd2.n76 vssa2 0.04fF $ **FLOATING
C1239 vccd2.n77 vssa2 0.18fF $ **FLOATING
C1240 vccd2.t154 vssa2 0.01fF
C1241 vccd2.t153 vssa2 0.01fF
C1242 vccd2.n78 vssa2 0.04fF $ **FLOATING
C1243 vccd2.n79 vssa2 0.08fF $ **FLOATING
C1244 vccd2.t3 vssa2 0.01fF
C1245 vccd2.t44 vssa2 0.01fF
C1246 vccd2.n80 vssa2 0.04fF $ **FLOATING
C1247 vccd2.n81 vssa2 0.07fF $ **FLOATING
C1248 vccd2.n82 vssa2 0.16fF $ **FLOATING
C1249 vccd2.t51 vssa2 0.01fF
C1250 vccd2.t156 vssa2 0.01fF
C1251 vccd2.n83 vssa2 0.04fF $ **FLOATING
C1252 vccd2.n84 vssa2 0.07fF $ **FLOATING
C1253 vccd2.t48 vssa2 0.01fF
C1254 vccd2.t9 vssa2 0.01fF
C1255 vccd2.n85 vssa2 0.05fF $ **FLOATING
C1256 vccd2.n86 vssa2 0.23fF $ **FLOATING
C1257 vccd2.n87 vssa2 0.01fF $ **FLOATING
C1258 vccd2.n88 vssa2 0.00fF $ **FLOATING
C1259 vccd2.n89 vssa2 0.00fF $ **FLOATING
C1260 vccd2.n90 vssa2 0.01fF $ **FLOATING
C1261 vccd2.t39 vssa2 0.21fF
C1262 vccd2.t127 vssa2 0.21fF
C1263 vccd2.t0 vssa2 0.21fF
C1264 vccd2.t79 vssa2 0.21fF
C1265 vccd2.n91 vssa2 0.05fF $ **FLOATING
C1266 vccd2.n92 vssa2 0.05fF $ **FLOATING
C1267 vccd2.n93 vssa2 0.00fF $ **FLOATING
C1268 vccd2.n94 vssa2 0.01fF $ **FLOATING
C1269 vccd2.t20 vssa2 0.21fF
C1270 vccd2.t113 vssa2 0.21fF
C1271 vccd2.t10 vssa2 0.21fF
C1272 vccd2.t89 vssa2 0.21fF
C1273 vccd2.n95 vssa2 0.00fF $ **FLOATING
C1274 vccd2.n96 vssa2 0.01fF $ **FLOATING
C1275 vccd2.n97 vssa2 0.11fF $ **FLOATING
C1276 vccd2.t142 vssa2 0.53fF
C1277 vccd2.t98 vssa2 0.01fF
C1278 vccd2.t134 vssa2 0.01fF
C1279 vccd2.n98 vssa2 0.04fF $ **FLOATING
C1280 vccd2.n99 vssa2 0.08fF $ **FLOATING
C1281 vccd2.t94 vssa2 0.01fF
C1282 vccd2.t102 vssa2 0.01fF
C1283 vccd2.t126 vssa2 0.01fF
C1284 vccd2.n100 vssa2 0.04fF $ **FLOATING
C1285 vccd2.n101 vssa2 0.18fF $ **FLOATING
C1286 vccd2.n102 vssa2 0.27fF $ **FLOATING
C1287 vccd2.t122 vssa2 0.01fF
C1288 vccd2.t128 vssa2 0.01fF
C1289 vccd2.n103 vssa2 0.04fF $ **FLOATING
C1290 vccd2.n104 vssa2 0.09fF $ **FLOATING
C1291 vccd2.t106 vssa2 0.01fF
C1292 vccd2.t100 vssa2 0.01fF
C1293 vccd2.n105 vssa2 0.04fF $ **FLOATING
C1294 vccd2.n106 vssa2 0.07fF $ **FLOATING
C1295 vccd2.t68 vssa2 0.01fF
C1296 vccd2.t72 vssa2 0.01fF
C1297 vccd2.n107 vssa2 0.04fF $ **FLOATING
C1298 vccd2.n108 vssa2 0.09fF $ **FLOATING
C1299 vccd2.t88 vssa2 0.01fF
C1300 vccd2.t96 vssa2 0.01fF
C1301 vccd2.n109 vssa2 0.04fF $ **FLOATING
C1302 vccd2.n110 vssa2 0.09fF $ **FLOATING
C1303 vccd2.t62 vssa2 0.01fF
C1304 vccd2.t108 vssa2 0.01fF
C1305 vccd2.n111 vssa2 0.04fF $ **FLOATING
C1306 vccd2.n112 vssa2 0.09fF $ **FLOATING
C1307 vccd2.t130 vssa2 0.01fF
C1308 vccd2.t64 vssa2 0.01fF
C1309 vccd2.n113 vssa2 0.04fF $ **FLOATING
C1310 vccd2.n114 vssa2 0.09fF $ **FLOATING
C1311 vccd2.t70 vssa2 0.01fF
C1312 vccd2.t120 vssa2 0.01fF
C1313 vccd2.n115 vssa2 0.04fF $ **FLOATING
C1314 vccd2.n116 vssa2 0.07fF $ **FLOATING
C1315 vccd2.n117 vssa2 0.26fF $ **FLOATING
C1316 vccd2.t86 vssa2 0.01fF
C1317 vccd2.t112 vssa2 0.01fF
C1318 vccd2.n118 vssa2 0.04fF $ **FLOATING
C1319 vccd2.n119 vssa2 0.07fF $ **FLOATING
C1320 vccd2.t78 vssa2 0.01fF
C1321 vccd2.t110 vssa2 0.01fF
C1322 vccd2.t132 vssa2 0.01fF
C1323 vccd2.n120 vssa2 0.04fF $ **FLOATING
C1324 vccd2.n121 vssa2 0.18fF $ **FLOATING
C1325 vccd2.n122 vssa2 0.27fF $ **FLOATING
C1326 vccd2.t74 vssa2 0.01fF
C1327 vccd2.t116 vssa2 0.01fF
C1328 vccd2.n123 vssa2 0.04fF $ **FLOATING
C1329 vccd2.n124 vssa2 0.09fF $ **FLOATING
C1330 vccd2.t136 vssa2 0.01fF
C1331 vccd2.t60 vssa2 0.01fF
C1332 vccd2.n125 vssa2 0.04fF $ **FLOATING
C1333 vccd2.n126 vssa2 0.09fF $ **FLOATING
C1334 vccd2.t118 vssa2 0.01fF
C1335 vccd2.t124 vssa2 0.01fF
C1336 vccd2.n127 vssa2 0.04fF $ **FLOATING
C1337 vccd2.n128 vssa2 0.09fF $ **FLOATING
C1338 vccd2.t82 vssa2 0.01fF
C1339 vccd2.t104 vssa2 0.01fF
C1340 vccd2.n129 vssa2 0.04fF $ **FLOATING
C1341 vccd2.n130 vssa2 0.09fF $ **FLOATING
C1342 vccd2.t66 vssa2 0.01fF
C1343 vccd2.t76 vssa2 0.01fF
C1344 vccd2.n131 vssa2 0.04fF $ **FLOATING
C1345 vccd2.n132 vssa2 0.07fF $ **FLOATING
C1346 vccd2.t80 vssa2 0.01fF
C1347 vccd2.t90 vssa2 0.01fF
C1348 vccd2.n133 vssa2 0.04fF $ **FLOATING
C1349 vccd2.n134 vssa2 0.09fF $ **FLOATING
C1350 vccd2.t114 vssa2 0.01fF
C1351 vccd2.t84 vssa2 0.01fF
C1352 vccd2.n135 vssa2 0.04fF $ **FLOATING
C1353 vccd2.n136 vssa2 0.09fF $ **FLOATING
C1354 vccd2.t92 vssa2 0.01fF
C1355 vccd2.t138 vssa2 0.01fF
C1356 vccd2.n137 vssa2 0.04fF $ **FLOATING
C1357 vccd2.n138 vssa2 0.07fF $ **FLOATING
C1358 vccd2.n139 vssa2 0.25fF $ **FLOATING
C1359 vccd2.n140 vssa2 0.03fF $ **FLOATING
C1360 vccd2.n141 vssa2 0.03fF $ **FLOATING
C1361 vccd2.n142 vssa2 0.82fF $ **FLOATING
C1362 vccd2.n143 vssa2 0.66fF $ **FLOATING
C1363 vccd2.n144 vssa2 1.15fF $ **FLOATING
C1364 vccd2.n145 vssa2 0.85fF $ **FLOATING
C1365 vccd2.n146 vssa2 0.01fF $ **FLOATING
C1366 vccd2.t35 vssa2 0.01fF
C1367 vccd2.t151 vssa2 0.01fF
C1368 vccd2.n147 vssa2 0.04fF $ **FLOATING
C1369 vccd2.n148 vssa2 0.08fF $ **FLOATING
C1370 vccd2.t145 vssa2 0.01fF
C1371 vccd2.t40 vssa2 0.01fF
C1372 vccd2.n149 vssa2 0.04fF $ **FLOATING
C1373 vccd2.n150 vssa2 0.08fF $ **FLOATING
C1374 vccd2.t1 vssa2 0.01fF
C1375 vccd2.t143 vssa2 0.01fF
C1376 vccd2.n151 vssa2 0.04fF $ **FLOATING
C1377 vccd2.n152 vssa2 0.07fF $ **FLOATING
C1378 vccd2.n153 vssa2 0.01fF $ **FLOATING
C1379 vccd2.t11 vssa2 0.01fF
C1380 vccd2.t21 vssa2 0.01fF
C1381 vccd2.n154 vssa2 0.04fF $ **FLOATING
C1382 vccd2.n155 vssa2 0.06fF $ **FLOATING
C1383 vccd2.n156 vssa2 0.01fF $ **FLOATING
C1384 vccd2.n157 vssa2 0.01fF $ **FLOATING
C1385 vccd2.n158 vssa2 0.24fF $ **FLOATING
C1386 vccd2.n159 vssa2 0.01fF $ **FLOATING
C1387 vccd2.n160 vssa2 0.01fF $ **FLOATING
C1388 vccd2.n161 vssa2 0.02fF $ **FLOATING
C1389 vccd2.t83 vssa2 0.21fF
C1390 vccd2.t52 vssa2 0.21fF
C1391 vccd2.t91 vssa2 0.21fF
C1392 vccd2.t22 vssa2 0.21fF
C1393 vccd2.t137 vssa2 0.14fF
C1394 vccd2.n162 vssa2 0.03fF $ **FLOATING
C1395 vccd2.n163 vssa2 0.45fF $ **FLOATING
C1396 vccd2.t77 vssa2 0.47fF
C1397 vccd2.t131 vssa2 0.43fF
C1398 vccd2.t109 vssa2 0.43fF
C1399 vccd2.t111 vssa2 0.43fF
C1400 vccd2.t85 vssa2 0.26fF
C1401 vccd2.n164 vssa2 0.04fF $ **FLOATING
C1402 vccd2.n165 vssa2 0.04fF $ **FLOATING
C1403 vccd2.n166 vssa2 0.03fF $ **FLOATING
C1404 vccd2.n167 vssa2 0.04fF $ **FLOATING
C1405 vccd2.n168 vssa2 0.21fF $ **FLOATING
C1406 vccd2.t115 vssa2 0.37fF
C1407 vccd2.t73 vssa2 0.43fF
C1408 vccd2.t59 vssa2 0.43fF
C1409 vccd2.t135 vssa2 0.27fF
C1410 vccd2.n169 vssa2 0.03fF $ **FLOATING
C1411 vccd2.n170 vssa2 0.03fF $ **FLOATING
C1412 vccd2.n171 vssa2 0.02fF $ **FLOATING
C1413 vccd2.n172 vssa2 0.02fF $ **FLOATING
C1414 vccd2.n173 vssa2 0.21fF $ **FLOATING
C1415 vccd2.t123 vssa2 0.26fF
C1416 vccd2.t8 vssa2 0.21fF
C1417 vccd2.t117 vssa2 0.21fF
C1418 vccd2.t47 vssa2 0.19fF
C1419 vccd2.n174 vssa2 0.02fF $ **FLOATING
C1420 vccd2.n175 vssa2 0.01fF $ **FLOATING
C1421 vccd2.n176 vssa2 0.02fF $ **FLOATING
C1422 vccd2.n177 vssa2 0.10fF $ **FLOATING
C1423 vccd2.t103 vssa2 0.10fF
C1424 vccd2.n178 vssa2 0.02fF $ **FLOATING
C1425 vccd2.n179 vssa2 0.02fF $ **FLOATING
C1426 vccd2.n180 vssa2 0.11fF $ **FLOATING
C1427 vccd2.t45 vssa2 0.13fF
C1428 vccd2.t81 vssa2 0.21fF
C1429 vccd2.t30 vssa2 0.21fF
C1430 vccd2.t75 vssa2 0.21fF
C1431 vccd2.t55 vssa2 0.21fF
C1432 vccd2.t65 vssa2 0.21fF
C1433 vccd2.t4 vssa2 0.18fF
C1434 vccd2.n181 vssa2 0.01fF $ **FLOATING
C1435 vccd2.n182 vssa2 0.13fF $ **FLOATING
C1436 vccd2.n183 vssa2 0.06fF $ **FLOATING
C1437 vccd2.n184 vssa2 0.23fF $ **FLOATING
C1438 vccd2.n185 vssa2 0.73fF $ **FLOATING
C1439 vccd2.n186 vssa2 0.17fF $ **FLOATING
C1440 vccd2.n187 vssa2 2.91fF $ **FLOATING
C1441 vccd2.n188 vssa2 149.18fF $ **FLOATING
C1442 vccd2.n189 vssa2 1.83fF $ **FLOATING
C1443 vccd2.n190 vssa2 0.39fF $ **FLOATING
C1444 vccd2.t139 vssa2 0.01fF
C1445 vccd2.t36 vssa2 0.01fF
C1446 vccd2.n191 vssa2 0.04fF $ **FLOATING
C1447 vccd2.n192 vssa2 0.31fF $ **FLOATING
C1448 vccd2.t158 vssa2 0.01fF
C1449 vccd2.t38 vssa2 0.01fF
C1450 vccd2.n193 vssa2 0.04fF $ **FLOATING
C1451 vccd2.n194 vssa2 0.24fF $ **FLOATING
C1452 vccd2.t25 vssa2 0.01fF
C1453 vccd2.t33 vssa2 0.01fF
C1454 vccd2.t144 vssa2 0.01fF
C1455 vccd2.n195 vssa2 0.05fF $ **FLOATING
C1456 vccd2.n196 vssa2 0.06fF $ **FLOATING
C1457 vccd2.n197 vssa2 0.10fF $ **FLOATING
C1458 vccd2.n198 vssa2 0.15fF $ **FLOATING
C1459 vccd2.n199 vssa2 0.03fF $ **FLOATING
C1460 vccd2.t28 vssa2 0.01fF
C1461 vccd2.n200 vssa2 0.00fF $ **FLOATING
C1462 vccd2.n201 vssa2 0.00fF $ **FLOATING
C1463 vccd2.n202 vssa2 0.02fF $ **FLOATING
C1464 vccd2.n203 vssa2 0.02fF $ **FLOATING
C1465 vccd2.n204 vssa2 0.02fF $ **FLOATING
C1466 vccd2.n205 vssa2 0.02fF $ **FLOATING
C1467 vccd2.n206 vssa2 0.02fF $ **FLOATING
C1468 vccd2.n207 vssa2 0.02fF $ **FLOATING
C1469 vccd2.n208 vssa2 0.02fF $ **FLOATING
C1470 vccd2.n209 vssa2 0.02fF $ **FLOATING
C1471 vccd2.n210 vssa2 0.21fF $ **FLOATING
C1472 vccd2.t37 vssa2 0.32fF
C1473 vccd2.t32 vssa2 0.43fF
C1474 vccd2.t24 vssa2 0.42fF
C1475 vccd2.n211 vssa2 0.01fF $ **FLOATING
C1476 vccd2.n212 vssa2 0.02fF $ **FLOATING
C1477 vccd2.n213 vssa2 0.00fF $ **FLOATING
C1478 vccd2.n214 vssa2 0.00fF $ **FLOATING
C1479 vccd2.n215 vssa2 0.08fF $ **FLOATING
C1480 vccd2.n216 vssa2 0.00fF $ **FLOATING
C1481 vccd2.n218 vssa2 0.01fF $ **FLOATING
C1482 vccd2.n219 vssa2 0.01fF $ **FLOATING
C1483 vccd2.n220 vssa2 0.01fF $ **FLOATING
C1484 vccd2.n221 vssa2 0.02fF $ **FLOATING
C1485 vccd2.n222 vssa2 0.01fF $ **FLOATING
C1486 vccd2.n223 vssa2 0.02fF $ **FLOATING
C1487 vccd2.n224 vssa2 0.29fF $ **FLOATING
C1488 vccd2.n226 vssa2 0.00fF $ **FLOATING
C1489 vccd2.n227 vssa2 0.03fF $ **FLOATING
C1490 vccd2.n228 vssa2 0.04fF $ **FLOATING
C1491 vccd2.n229 vssa2 0.03fF $ **FLOATING
C1492 vccd2.n230 vssa2 0.24fF $ **FLOATING
C1493 vccd2.n231 vssa2 0.07fF $ **FLOATING
C1494 a_40125_693523.t62 vssa2 0.24fF
C1495 a_40125_693523.t35 vssa2 0.24fF
C1496 a_40125_693523.t43 vssa2 0.24fF
C1497 a_40125_693523.t48 vssa2 0.24fF
C1498 a_40125_693523.t58 vssa2 0.24fF
C1499 a_40125_693523.t46 vssa2 0.24fF
C1500 a_40125_693523.t64 vssa2 0.24fF
C1501 a_40125_693523.n0 vssa2 0.18fF $ **FLOATING
C1502 a_40125_693523.n1 vssa2 0.18fF $ **FLOATING
C1503 a_40125_693523.n2 vssa2 0.18fF $ **FLOATING
C1504 a_40125_693523.n3 vssa2 0.18fF $ **FLOATING
C1505 a_40125_693523.n4 vssa2 0.18fF $ **FLOATING
C1506 a_40125_693523.n5 vssa2 0.18fF $ **FLOATING
C1507 a_40125_693523.n6 vssa2 0.18fF $ **FLOATING
C1508 a_40125_693523.n7 vssa2 0.18fF $ **FLOATING
C1509 a_40125_693523.n8 vssa2 0.18fF $ **FLOATING
C1510 a_40125_693523.n9 vssa2 0.18fF $ **FLOATING
C1511 a_40125_693523.n10 vssa2 0.18fF $ **FLOATING
C1512 a_40125_693523.n11 vssa2 0.18fF $ **FLOATING
C1513 a_40125_693523.n12 vssa2 0.18fF $ **FLOATING
C1514 a_40125_693523.n13 vssa2 0.18fF $ **FLOATING
C1515 a_40125_693523.n14 vssa2 0.18fF $ **FLOATING
C1516 a_40125_693523.n15 vssa2 0.18fF $ **FLOATING
C1517 a_40125_693523.n16 vssa2 0.18fF $ **FLOATING
C1518 a_40125_693523.n17 vssa2 0.18fF $ **FLOATING
C1519 a_40125_693523.n18 vssa2 0.18fF $ **FLOATING
C1520 a_40125_693523.n19 vssa2 0.18fF $ **FLOATING
C1521 a_40125_693523.n20 vssa2 0.18fF $ **FLOATING
C1522 a_40125_693523.n21 vssa2 0.18fF $ **FLOATING
C1523 a_40125_693523.n22 vssa2 0.18fF $ **FLOATING
C1524 a_40125_693523.n23 vssa2 0.18fF $ **FLOATING
C1525 a_40125_693523.n24 vssa2 0.18fF $ **FLOATING
C1526 a_40125_693523.n25 vssa2 0.18fF $ **FLOATING
C1527 a_40125_693523.n26 vssa2 0.18fF $ **FLOATING
C1528 a_40125_693523.n27 vssa2 0.18fF $ **FLOATING
C1529 a_40125_693523.n28 vssa2 0.18fF $ **FLOATING
C1530 a_40125_693523.n29 vssa2 0.18fF $ **FLOATING
C1531 a_40125_693523.n30 vssa2 0.18fF $ **FLOATING
C1532 a_40125_693523.n31 vssa2 0.24fF $ **FLOATING
C1533 a_40125_693523.t33 vssa2 0.24fF
C1534 a_40125_693523.t41 vssa2 0.24fF
C1535 a_40125_693523.t45 vssa2 0.24fF
C1536 a_40125_693523.t49 vssa2 0.24fF
C1537 a_40125_693523.t60 vssa2 0.24fF
C1538 a_40125_693523.t63 vssa2 0.24fF
C1539 a_40125_693523.t68 vssa2 0.24fF
C1540 a_40125_693523.t32 vssa2 0.24fF
C1541 a_40125_693523.t55 vssa2 0.24fF
C1542 a_40125_693523.t59 vssa2 0.24fF
C1543 a_40125_693523.t47 vssa2 0.24fF
C1544 a_40125_693523.t56 vssa2 0.24fF
C1545 a_40125_693523.t61 vssa2 0.24fF
C1546 a_40125_693523.t37 vssa2 0.24fF
C1547 a_40125_693523.t42 vssa2 0.24fF
C1548 a_40125_693523.n32 vssa2 0.18fF $ **FLOATING
C1549 a_40125_693523.n33 vssa2 0.18fF $ **FLOATING
C1550 a_40125_693523.n34 vssa2 0.18fF $ **FLOATING
C1551 a_40125_693523.n35 vssa2 0.18fF $ **FLOATING
C1552 a_40125_693523.n36 vssa2 0.18fF $ **FLOATING
C1553 a_40125_693523.n37 vssa2 0.18fF $ **FLOATING
C1554 a_40125_693523.n38 vssa2 0.18fF $ **FLOATING
C1555 a_40125_693523.n39 vssa2 0.18fF $ **FLOATING
C1556 a_40125_693523.n40 vssa2 0.18fF $ **FLOATING
C1557 a_40125_693523.n41 vssa2 0.18fF $ **FLOATING
C1558 a_40125_693523.n42 vssa2 0.18fF $ **FLOATING
C1559 a_40125_693523.n43 vssa2 0.18fF $ **FLOATING
C1560 a_40125_693523.n44 vssa2 0.18fF $ **FLOATING
C1561 a_40125_693523.n45 vssa2 0.18fF $ **FLOATING
C1562 a_40125_693523.n46 vssa2 0.18fF $ **FLOATING
C1563 a_40125_693523.t71 vssa2 0.24fF
C1564 a_40125_693523.n47 vssa2 0.18fF $ **FLOATING
C1565 a_40125_693523.t65 vssa2 0.24fF
C1566 a_40125_693523.t67 vssa2 0.24fF
C1567 a_40125_693523.t34 vssa2 0.24fF
C1568 a_40125_693523.t52 vssa2 0.24fF
C1569 a_40125_693523.t40 vssa2 0.24fF
C1570 a_40125_693523.t50 vssa2 0.24fF
C1571 a_40125_693523.t54 vssa2 0.24fF
C1572 a_40125_693523.t17 vssa2 1.01fF
C1573 a_40125_693523.t6 vssa2 0.87fF
C1574 a_40125_693523.n48 vssa2 11.68fF $ **FLOATING
C1575 a_40125_693523.n49 vssa2 0.18fF $ **FLOATING
C1576 a_40125_693523.n50 vssa2 0.18fF $ **FLOATING
C1577 a_40125_693523.n51 vssa2 0.18fF $ **FLOATING
C1578 a_40125_693523.n52 vssa2 0.18fF $ **FLOATING
C1579 a_40125_693523.n53 vssa2 0.18fF $ **FLOATING
C1580 a_40125_693523.n54 vssa2 0.18fF $ **FLOATING
C1581 a_40125_693523.n55 vssa2 0.18fF $ **FLOATING
C1582 a_40125_693523.n56 vssa2 0.24fF $ **FLOATING
C1583 a_40125_693523.n57 vssa2 0.75fF $ **FLOATING
C1584 a_40125_693523.n58 vssa2 0.24fF $ **FLOATING
C1585 a_40125_693523.n59 vssa2 0.18fF $ **FLOATING
C1586 a_40125_693523.n60 vssa2 0.18fF $ **FLOATING
C1587 a_40125_693523.n61 vssa2 0.18fF $ **FLOATING
C1588 a_40125_693523.n62 vssa2 0.18fF $ **FLOATING
C1589 a_40125_693523.n63 vssa2 0.18fF $ **FLOATING
C1590 a_40125_693523.n64 vssa2 0.18fF $ **FLOATING
C1591 a_40125_693523.t51 vssa2 0.24fF
C1592 a_40125_693523.n65 vssa2 0.18fF $ **FLOATING
C1593 a_40125_693523.t39 vssa2 0.24fF
C1594 a_40125_693523.n66 vssa2 0.18fF $ **FLOATING
C1595 a_40125_693523.t44 vssa2 0.24fF
C1596 a_40125_693523.n67 vssa2 0.18fF $ **FLOATING
C1597 a_40125_693523.t66 vssa2 0.24fF
C1598 a_40125_693523.n68 vssa2 0.18fF $ **FLOATING
C1599 a_40125_693523.t69 vssa2 0.24fF
C1600 a_40125_693523.n69 vssa2 0.18fF $ **FLOATING
C1601 a_40125_693523.t36 vssa2 0.24fF
C1602 a_40125_693523.n70 vssa2 0.18fF $ **FLOATING
C1603 a_40125_693523.t38 vssa2 0.24fF
C1604 a_40125_693523.n71 vssa2 0.18fF $ **FLOATING
C1605 a_40125_693523.t70 vssa2 0.24fF
C1606 a_40125_693523.n72 vssa2 0.18fF $ **FLOATING
C1607 a_40125_693523.t53 vssa2 0.24fF
C1608 a_40125_693523.n73 vssa2 0.18fF $ **FLOATING
C1609 a_40125_693523.t57 vssa2 0.24fF
C1610 a_40125_693523.n74 vssa2 0.18fF $ **FLOATING
C1611 a_40125_693523.n75 vssa2 0.52fF $ **FLOATING
C1612 a_40125_693523.n76 vssa2 1.96fF $ **FLOATING
C1613 a_40125_693523.t2 vssa2 0.06fF
C1614 a_40125_693523.t31 vssa2 0.06fF
C1615 a_40125_693523.n77 vssa2 0.32fF $ **FLOATING
C1616 a_40125_693523.n78 vssa2 0.75fF $ **FLOATING
C1617 a_40125_693523.t24 vssa2 0.06fF
C1618 a_40125_693523.t0 vssa2 0.06fF
C1619 a_40125_693523.n79 vssa2 0.32fF $ **FLOATING
C1620 a_40125_693523.n80 vssa2 0.61fF $ **FLOATING
C1621 a_40125_693523.t9 vssa2 0.06fF
C1622 a_40125_693523.t27 vssa2 0.06fF
C1623 a_40125_693523.n81 vssa2 0.32fF $ **FLOATING
C1624 a_40125_693523.n82 vssa2 0.61fF $ **FLOATING
C1625 a_40125_693523.t26 vssa2 0.06fF
C1626 a_40125_693523.t8 vssa2 0.06fF
C1627 a_40125_693523.n83 vssa2 0.32fF $ **FLOATING
C1628 a_40125_693523.n84 vssa2 0.61fF $ **FLOATING
C1629 a_40125_693523.t20 vssa2 0.06fF
C1630 a_40125_693523.t15 vssa2 0.06fF
C1631 a_40125_693523.n85 vssa2 0.32fF $ **FLOATING
C1632 a_40125_693523.n86 vssa2 0.61fF $ **FLOATING
C1633 a_40125_693523.t29 vssa2 0.06fF
C1634 a_40125_693523.t12 vssa2 0.06fF
C1635 a_40125_693523.n87 vssa2 0.32fF $ **FLOATING
C1636 a_40125_693523.n88 vssa2 0.61fF $ **FLOATING
C1637 a_40125_693523.t19 vssa2 0.06fF
C1638 a_40125_693523.t14 vssa2 0.06fF
C1639 a_40125_693523.n89 vssa2 0.32fF $ **FLOATING
C1640 a_40125_693523.n90 vssa2 0.61fF $ **FLOATING
C1641 a_40125_693523.t25 vssa2 0.06fF
C1642 a_40125_693523.t1 vssa2 0.06fF
C1643 a_40125_693523.n91 vssa2 0.32fF $ **FLOATING
C1644 a_40125_693523.n92 vssa2 0.61fF $ **FLOATING
C1645 a_40125_693523.t16 vssa2 0.06fF
C1646 a_40125_693523.t13 vssa2 0.06fF
C1647 a_40125_693523.n93 vssa2 0.32fF $ **FLOATING
C1648 a_40125_693523.n94 vssa2 0.61fF $ **FLOATING
C1649 a_40125_693523.t28 vssa2 0.06fF
C1650 a_40125_693523.t11 vssa2 0.06fF
C1651 a_40125_693523.n95 vssa2 0.32fF $ **FLOATING
C1652 a_40125_693523.n96 vssa2 0.61fF $ **FLOATING
C1653 a_40125_693523.t3 vssa2 0.09fF
C1654 a_40125_693523.n97 vssa2 0.98fF $ **FLOATING
C1655 a_40125_693523.t22 vssa2 0.09fF
C1656 a_40125_693523.n98 vssa2 4.05fF $ **FLOATING
C1657 a_40125_693523.t21 vssa2 0.06fF
C1658 a_40125_693523.t4 vssa2 0.06fF
C1659 a_40125_693523.n99 vssa2 0.31fF $ **FLOATING
C1660 a_40125_693523.n100 vssa2 0.72fF $ **FLOATING
C1661 a_40125_693523.t18 vssa2 0.06fF
C1662 a_40125_693523.t23 vssa2 0.06fF
C1663 a_40125_693523.n101 vssa2 0.31fF $ **FLOATING
C1664 a_40125_693523.n102 vssa2 0.72fF $ **FLOATING
C1665 a_40125_693523.t10 vssa2 0.06fF
C1666 a_40125_693523.t7 vssa2 0.06fF
C1667 a_40125_693523.n103 vssa2 0.31fF $ **FLOATING
C1668 a_40125_693523.n104 vssa2 3.93fF $ **FLOATING
C1669 a_40125_693523.n105 vssa2 1.89fF $ **FLOATING
C1670 a_40125_693523.n106 vssa2 0.52fF $ **FLOATING
C1671 a_40125_693523.n107 vssa2 0.18fF $ **FLOATING
C1672 a_40125_693523.n108 vssa2 0.18fF $ **FLOATING
C1673 a_40125_693523.n109 vssa2 0.18fF $ **FLOATING
C1674 a_40125_693523.n110 vssa2 0.18fF $ **FLOATING
C1675 a_40125_693523.n111 vssa2 0.18fF $ **FLOATING
C1676 a_40125_693523.n112 vssa2 0.18fF $ **FLOATING
C1677 a_40125_693523.n113 vssa2 0.24fF $ **FLOATING
C1678 a_40125_693523.n114 vssa2 0.75fF $ **FLOATING
C1679 a_40125_693523.t30 vssa2 0.88fF
C1680 a_40125_693523.n115 vssa2 8.36fF $ **FLOATING
C1681 a_40125_693523.t5 vssa2 4.20fF
C1682 a_537154_685355.t43 vssa2 0.42fF
C1683 a_537154_685355.t33 vssa2 0.42fF
C1684 a_537154_685355.t46 vssa2 0.42fF
C1685 a_537154_685355.n0 vssa2 0.02fF $ **FLOATING
C1686 a_537154_685355.n1 vssa2 0.43fF $ **FLOATING
C1687 a_537154_685355.n2 vssa2 0.32fF $ **FLOATING
C1688 a_537154_685355.n3 vssa2 0.28fF $ **FLOATING
C1689 a_537154_685355.n4 vssa2 0.01fF $ **FLOATING
C1690 a_537154_685355.n5 vssa2 0.43fF $ **FLOATING
C1691 a_537154_685355.n6 vssa2 0.02fF $ **FLOATING
C1692 a_537154_685355.n7 vssa2 0.70fF $ **FLOATING
C1693 a_537154_685355.n8 vssa2 0.74fF $ **FLOATING
C1694 a_537154_685355.n9 vssa2 0.05fF $ **FLOATING
C1695 a_537154_685355.n10 vssa2 0.42fF $ **FLOATING
C1696 a_537154_685355.n11 vssa2 0.32fF $ **FLOATING
C1697 a_537154_685355.n12 vssa2 0.28fF $ **FLOATING
C1698 a_537154_685355.n13 vssa2 0.02fF $ **FLOATING
C1699 a_537154_685355.n14 vssa2 0.43fF $ **FLOATING
C1700 a_537154_685355.t58 vssa2 0.42fF
C1701 a_537154_685355.n15 vssa2 0.30fF $ **FLOATING
C1702 a_537154_685355.n16 vssa2 0.30fF $ **FLOATING
C1703 a_537154_685355.n17 vssa2 0.01fF $ **FLOATING
C1704 a_537154_685355.t56 vssa2 0.42fF
C1705 a_537154_685355.n18 vssa2 0.24fF $ **FLOATING
C1706 a_537154_685355.t38 vssa2 0.42fF
C1707 a_537154_685355.t60 vssa2 0.42fF
C1708 a_537154_685355.n19 vssa2 0.02fF $ **FLOATING
C1709 a_537154_685355.n20 vssa2 0.43fF $ **FLOATING
C1710 a_537154_685355.n21 vssa2 0.30fF $ **FLOATING
C1711 a_537154_685355.n22 vssa2 0.28fF $ **FLOATING
C1712 a_537154_685355.n23 vssa2 0.01fF $ **FLOATING
C1713 a_537154_685355.n24 vssa2 0.43fF $ **FLOATING
C1714 a_537154_685355.n25 vssa2 0.02fF $ **FLOATING
C1715 a_537154_685355.n26 vssa2 0.70fF $ **FLOATING
C1716 a_537154_685355.n27 vssa2 0.33fF $ **FLOATING
C1717 a_537154_685355.n28 vssa2 0.43fF $ **FLOATING
C1718 a_537154_685355.n29 vssa2 0.17fF $ **FLOATING
C1719 a_537154_685355.n30 vssa2 0.02fF $ **FLOATING
C1720 a_537154_685355.n31 vssa2 0.01fF $ **FLOATING
C1721 a_537154_685355.n32 vssa2 0.01fF $ **FLOATING
C1722 a_537154_685355.n33 vssa2 0.29fF $ **FLOATING
C1723 a_537154_685355.n34 vssa2 0.01fF $ **FLOATING
C1724 a_537154_685355.n35 vssa2 0.01fF $ **FLOATING
C1725 a_537154_685355.n36 vssa2 0.24fF $ **FLOATING
C1726 a_537154_685355.n37 vssa2 0.02fF $ **FLOATING
C1727 a_537154_685355.n38 vssa2 0.17fF $ **FLOATING
C1728 a_537154_685355.t67 vssa2 0.42fF
C1729 a_537154_685355.n39 vssa2 0.79fF $ **FLOATING
C1730 a_537154_685355.n40 vssa2 0.02fF $ **FLOATING
C1731 a_537154_685355.t59 vssa2 0.42fF
C1732 a_537154_685355.t40 vssa2 0.42fF
C1733 a_537154_685355.n41 vssa2 0.01fF $ **FLOATING
C1734 a_537154_685355.t61 vssa2 0.42fF
C1735 a_537154_685355.n42 vssa2 0.05fF $ **FLOATING
C1736 a_537154_685355.n43 vssa2 0.43fF $ **FLOATING
C1737 a_537154_685355.n44 vssa2 0.30fF $ **FLOATING
C1738 a_537154_685355.n45 vssa2 0.09fF $ **FLOATING
C1739 a_537154_685355.n46 vssa2 0.41fF $ **FLOATING
C1740 a_537154_685355.n47 vssa2 0.04fF $ **FLOATING
C1741 a_537154_685355.n48 vssa2 1.23fF $ **FLOATING
C1742 a_537154_685355.n49 vssa2 0.05fF $ **FLOATING
C1743 a_537154_685355.n50 vssa2 0.42fF $ **FLOATING
C1744 a_537154_685355.n51 vssa2 0.29fF $ **FLOATING
C1745 a_537154_685355.n52 vssa2 0.09fF $ **FLOATING
C1746 a_537154_685355.n53 vssa2 0.41fF $ **FLOATING
C1747 a_537154_685355.t70 vssa2 0.42fF
C1748 a_537154_685355.n54 vssa2 0.32fF $ **FLOATING
C1749 a_537154_685355.t31 vssa2 0.93fF
C1750 a_537154_685355.n55 vssa2 9.84fF $ **FLOATING
C1751 a_537154_685355.n56 vssa2 2.34fF $ **FLOATING
C1752 a_537154_685355.n57 vssa2 2.58fF $ **FLOATING
C1753 a_537154_685355.t42 vssa2 0.42fF
C1754 a_537154_685355.t16 vssa2 0.11fF
C1755 a_537154_685355.t17 vssa2 0.11fF
C1756 a_537154_685355.n58 vssa2 1.89fF $ **FLOATING
C1757 a_537154_685355.t13 vssa2 0.11fF
C1758 a_537154_685355.n59 vssa2 0.69fF $ **FLOATING
C1759 a_537154_685355.n60 vssa2 1.68fF $ **FLOATING
C1760 a_537154_685355.t8 vssa2 0.11fF
C1761 a_537154_685355.n61 vssa2 1.94fF $ **FLOATING
C1762 a_537154_685355.n62 vssa2 0.83fF $ **FLOATING
C1763 a_537154_685355.n63 vssa2 0.16fF $ **FLOATING
C1764 a_537154_685355.t12 vssa2 0.11fF
C1765 a_537154_685355.n64 vssa2 0.77fF $ **FLOATING
C1766 a_537154_685355.t7 vssa2 0.11fF
C1767 a_537154_685355.n65 vssa2 0.39fF $ **FLOATING
C1768 a_537154_685355.n66 vssa2 0.30fF $ **FLOATING
C1769 a_537154_685355.n67 vssa2 1.14fF $ **FLOATING
C1770 a_537154_685355.n68 vssa2 0.20fF $ **FLOATING
C1771 a_537154_685355.t23 vssa2 0.11fF
C1772 a_537154_685355.n69 vssa2 0.80fF $ **FLOATING
C1773 a_537154_685355.n70 vssa2 1.40fF $ **FLOATING
C1774 a_537154_685355.n71 vssa2 0.29fF $ **FLOATING
C1775 a_537154_685355.n72 vssa2 3.31fF $ **FLOATING
C1776 a_537154_685355.n73 vssa2 0.25fF $ **FLOATING
C1777 a_537154_685355.t14 vssa2 0.11fF
C1778 a_537154_685355.n74 vssa2 1.93fF $ **FLOATING
C1779 a_537154_685355.n75 vssa2 1.40fF $ **FLOATING
C1780 a_537154_685355.n76 vssa2 1.51fF $ **FLOATING
C1781 a_537154_685355.n77 vssa2 3.30fF $ **FLOATING
C1782 a_537154_685355.t10 vssa2 0.11fF
C1783 a_537154_685355.n78 vssa2 0.61fF $ **FLOATING
C1784 a_537154_685355.n79 vssa2 1.67fF $ **FLOATING
C1785 a_537154_685355.t26 vssa2 0.11fF
C1786 a_537154_685355.n80 vssa2 1.82fF $ **FLOATING
C1787 a_537154_685355.n81 vssa2 0.26fF $ **FLOATING
C1788 a_537154_685355.t21 vssa2 0.11fF
C1789 a_537154_685355.n82 vssa2 0.81fF $ **FLOATING
C1790 a_537154_685355.n83 vssa2 0.32fF $ **FLOATING
C1791 a_537154_685355.n84 vssa2 0.93fF $ **FLOATING
C1792 a_537154_685355.t11 vssa2 0.11fF
C1793 a_537154_685355.n85 vssa2 0.40fF $ **FLOATING
C1794 a_537154_685355.n86 vssa2 0.24fF $ **FLOATING
C1795 a_537154_685355.n87 vssa2 0.25fF $ **FLOATING
C1796 a_537154_685355.t22 vssa2 0.11fF
C1797 a_537154_685355.n88 vssa2 0.82fF $ **FLOATING
C1798 a_537154_685355.t20 vssa2 0.11fF
C1799 a_537154_685355.n89 vssa2 0.40fF $ **FLOATING
C1800 a_537154_685355.n90 vssa2 0.32fF $ **FLOATING
C1801 a_537154_685355.n91 vssa2 1.14fF $ **FLOATING
C1802 a_537154_685355.t9 vssa2 0.11fF
C1803 a_537154_685355.n92 vssa2 0.76fF $ **FLOATING
C1804 a_537154_685355.n93 vssa2 0.29fF $ **FLOATING
C1805 a_537154_685355.n94 vssa2 1.01fF $ **FLOATING
C1806 a_537154_685355.t18 vssa2 0.11fF
C1807 a_537154_685355.n95 vssa2 0.39fF $ **FLOATING
C1808 a_537154_685355.n96 vssa2 0.22fF $ **FLOATING
C1809 a_537154_685355.n97 vssa2 1.33fF $ **FLOATING
C1810 a_537154_685355.n98 vssa2 1.52fF $ **FLOATING
C1811 a_537154_685355.t25 vssa2 0.11fF
C1812 a_537154_685355.n99 vssa2 0.76fF $ **FLOATING
C1813 a_537154_685355.n100 vssa2 0.29fF $ **FLOATING
C1814 a_537154_685355.n101 vssa2 1.44fF $ **FLOATING
C1815 a_537154_685355.t15 vssa2 0.11fF
C1816 a_537154_685355.n102 vssa2 0.39fF $ **FLOATING
C1817 a_537154_685355.n103 vssa2 0.21fF $ **FLOATING
C1818 a_537154_685355.n104 vssa2 0.24fF $ **FLOATING
C1819 a_537154_685355.t27 vssa2 0.11fF
C1820 a_537154_685355.n105 vssa2 0.77fF $ **FLOATING
C1821 a_537154_685355.t24 vssa2 0.11fF
C1822 a_537154_685355.n106 vssa2 0.39fF $ **FLOATING
C1823 a_537154_685355.n107 vssa2 0.30fF $ **FLOATING
C1824 a_537154_685355.n108 vssa2 1.62fF $ **FLOATING
C1825 a_537154_685355.n109 vssa2 0.20fF $ **FLOATING
C1826 a_537154_685355.t19 vssa2 0.11fF
C1827 a_537154_685355.n110 vssa2 0.90fF $ **FLOATING
C1828 a_537154_685355.n111 vssa2 1.67fF $ **FLOATING
C1829 a_537154_685355.n112 vssa2 3.52fF $ **FLOATING
C1830 a_537154_685355.n113 vssa2 0.03fF $ **FLOATING
C1831 a_537154_685355.n114 vssa2 0.41fF $ **FLOATING
C1832 a_537154_685355.t48 vssa2 0.42fF
C1833 a_537154_685355.n115 vssa2 0.05fF $ **FLOATING
C1834 a_537154_685355.n116 vssa2 0.41fF $ **FLOATING
C1835 a_537154_685355.n117 vssa2 0.09fF $ **FLOATING
C1836 a_537154_685355.n118 vssa2 0.30fF $ **FLOATING
C1837 a_537154_685355.n119 vssa2 0.30fF $ **FLOATING
C1838 a_537154_685355.t45 vssa2 0.42fF
C1839 a_537154_685355.n120 vssa2 0.02fF $ **FLOATING
C1840 a_537154_685355.n121 vssa2 0.43fF $ **FLOATING
C1841 a_537154_685355.n122 vssa2 0.43fF $ **FLOATING
C1842 a_537154_685355.n123 vssa2 0.03fF $ **FLOATING
C1843 a_537154_685355.n124 vssa2 0.28fF $ **FLOATING
C1844 a_537154_685355.n125 vssa2 0.32fF $ **FLOATING
C1845 a_537154_685355.t37 vssa2 0.42fF
C1846 a_537154_685355.n126 vssa2 0.02fF $ **FLOATING
C1847 a_537154_685355.n127 vssa2 0.43fF $ **FLOATING
C1848 a_537154_685355.n128 vssa2 0.43fF $ **FLOATING
C1849 a_537154_685355.n129 vssa2 0.03fF $ **FLOATING
C1850 a_537154_685355.n130 vssa2 0.28fF $ **FLOATING
C1851 a_537154_685355.n131 vssa2 0.32fF $ **FLOATING
C1852 a_537154_685355.t36 vssa2 0.42fF
C1853 a_537154_685355.n132 vssa2 0.02fF $ **FLOATING
C1854 a_537154_685355.n133 vssa2 0.43fF $ **FLOATING
C1855 a_537154_685355.n134 vssa2 0.43fF $ **FLOATING
C1856 a_537154_685355.n135 vssa2 0.03fF $ **FLOATING
C1857 a_537154_685355.n136 vssa2 0.34fF $ **FLOATING
C1858 a_537154_685355.t1 vssa2 0.11fF
C1859 a_537154_685355.t66 vssa2 0.42fF
C1860 a_537154_685355.n137 vssa2 0.04fF $ **FLOATING
C1861 a_537154_685355.n138 vssa2 1.21fF $ **FLOATING
C1862 a_537154_685355.t64 vssa2 0.42fF
C1863 a_537154_685355.n139 vssa2 0.04fF $ **FLOATING
C1864 a_537154_685355.n140 vssa2 1.45fF $ **FLOATING
C1865 a_537154_685355.n141 vssa2 0.74fF $ **FLOATING
C1866 a_537154_685355.t52 vssa2 0.42fF
C1867 a_537154_685355.n142 vssa2 0.02fF $ **FLOATING
C1868 a_537154_685355.n143 vssa2 0.70fF $ **FLOATING
C1869 a_537154_685355.n144 vssa2 0.75fF $ **FLOATING
C1870 a_537154_685355.t50 vssa2 0.42fF
C1871 a_537154_685355.n145 vssa2 0.02fF $ **FLOATING
C1872 a_537154_685355.n146 vssa2 0.77fF $ **FLOATING
C1873 a_537154_685355.n147 vssa2 0.02fF $ **FLOATING
C1874 a_537154_685355.n148 vssa2 0.41fF $ **FLOATING
C1875 a_537154_685355.t55 vssa2 0.42fF
C1876 a_537154_685355.n149 vssa2 0.05fF $ **FLOATING
C1877 a_537154_685355.n150 vssa2 0.42fF $ **FLOATING
C1878 a_537154_685355.n151 vssa2 0.09fF $ **FLOATING
C1879 a_537154_685355.n152 vssa2 0.30fF $ **FLOATING
C1880 a_537154_685355.t51 vssa2 0.42fF
C1881 a_537154_685355.n153 vssa2 0.05fF $ **FLOATING
C1882 a_537154_685355.n154 vssa2 1.43fF $ **FLOATING
C1883 a_537154_685355.t41 vssa2 0.42fF
C1884 a_537154_685355.n155 vssa2 0.05fF $ **FLOATING
C1885 a_537154_685355.n156 vssa2 0.42fF $ **FLOATING
C1886 a_537154_685355.n157 vssa2 0.32fF $ **FLOATING
C1887 a_537154_685355.n158 vssa2 0.43fF $ **FLOATING
C1888 a_537154_685355.n159 vssa2 0.02fF $ **FLOATING
C1889 a_537154_685355.n160 vssa2 0.28fF $ **FLOATING
C1890 a_537154_685355.t39 vssa2 0.42fF
C1891 a_537154_685355.n161 vssa2 0.05fF $ **FLOATING
C1892 a_537154_685355.n162 vssa2 0.42fF $ **FLOATING
C1893 a_537154_685355.n163 vssa2 0.32fF $ **FLOATING
C1894 a_537154_685355.n164 vssa2 0.43fF $ **FLOATING
C1895 a_537154_685355.n165 vssa2 0.02fF $ **FLOATING
C1896 a_537154_685355.n166 vssa2 0.34fF $ **FLOATING
C1897 a_537154_685355.t3 vssa2 0.11fF
C1898 a_537154_685355.t63 vssa2 0.42fF
C1899 a_537154_685355.n167 vssa2 0.04fF $ **FLOATING
C1900 a_537154_685355.n168 vssa2 1.24fF $ **FLOATING
C1901 a_537154_685355.n169 vssa2 0.74fF $ **FLOATING
C1902 a_537154_685355.t62 vssa2 0.42fF
C1903 a_537154_685355.n170 vssa2 0.02fF $ **FLOATING
C1904 a_537154_685355.n171 vssa2 0.70fF $ **FLOATING
C1905 a_537154_685355.t49 vssa2 0.42fF
C1906 a_537154_685355.n172 vssa2 0.04fF $ **FLOATING
C1907 a_537154_685355.n173 vssa2 1.45fF $ **FLOATING
C1908 a_537154_685355.n174 vssa2 0.74fF $ **FLOATING
C1909 a_537154_685355.t47 vssa2 0.42fF
C1910 a_537154_685355.n175 vssa2 0.02fF $ **FLOATING
C1911 a_537154_685355.n176 vssa2 0.76fF $ **FLOATING
C1912 a_537154_685355.n177 vssa2 0.01fF $ **FLOATING
C1913 a_537154_685355.n178 vssa2 0.41fF $ **FLOATING
C1914 a_537154_685355.t35 vssa2 0.42fF
C1915 a_537154_685355.t71 vssa2 0.42fF
C1916 a_537154_685355.n179 vssa2 0.34fF $ **FLOATING
C1917 a_537154_685355.n180 vssa2 0.41fF $ **FLOATING
C1918 a_537154_685355.n181 vssa2 0.03fF $ **FLOATING
C1919 a_537154_685355.n182 vssa2 0.43fF $ **FLOATING
C1920 a_537154_685355.n183 vssa2 0.02fF $ **FLOATING
C1921 a_537154_685355.n184 vssa2 0.43fF $ **FLOATING
C1922 a_537154_685355.n185 vssa2 0.10fF $ **FLOATING
C1923 a_537154_685355.n186 vssa2 0.30fF $ **FLOATING
C1924 a_537154_685355.t34 vssa2 0.42fF
C1925 a_537154_685355.t68 vssa2 0.42fF
C1926 a_537154_685355.n187 vssa2 0.32fF $ **FLOATING
C1927 a_537154_685355.n188 vssa2 0.44fF $ **FLOATING
C1928 a_537154_685355.n189 vssa2 0.03fF $ **FLOATING
C1929 a_537154_685355.n190 vssa2 0.43fF $ **FLOATING
C1930 a_537154_685355.n191 vssa2 0.02fF $ **FLOATING
C1931 a_537154_685355.n192 vssa2 0.43fF $ **FLOATING
C1932 a_537154_685355.n193 vssa2 0.30fF $ **FLOATING
C1933 a_537154_685355.n194 vssa2 0.43fF $ **FLOATING
C1934 a_537154_685355.n195 vssa2 0.01fF $ **FLOATING
C1935 a_537154_685355.n196 vssa2 0.28fF $ **FLOATING
C1936 a_537154_685355.t69 vssa2 0.42fF
C1937 a_537154_685355.t57 vssa2 0.42fF
C1938 a_537154_685355.n197 vssa2 0.32fF $ **FLOATING
C1939 a_537154_685355.n198 vssa2 0.43fF $ **FLOATING
C1940 a_537154_685355.n199 vssa2 0.03fF $ **FLOATING
C1941 a_537154_685355.n200 vssa2 0.10fF $ **FLOATING
C1942 a_537154_685355.n201 vssa2 0.28fF $ **FLOATING
C1943 a_537154_685355.n202 vssa2 0.32fF $ **FLOATING
C1944 a_537154_685355.n203 vssa2 0.28fF $ **FLOATING
C1945 a_537154_685355.n204 vssa2 0.32fF $ **FLOATING
C1946 a_537154_685355.n205 vssa2 0.41fF $ **FLOATING
C1947 a_537154_685355.n206 vssa2 0.05fF $ **FLOATING
C1948 a_537154_685355.n207 vssa2 1.45fF $ **FLOATING
C1949 a_537154_685355.t53 vssa2 0.42fF
C1950 a_537154_685355.t30 vssa2 0.91fF
C1951 a_537154_685355.t28 vssa2 0.94fF
C1952 a_537154_685355.n208 vssa2 10.66fF $ **FLOATING
C1953 a_537154_685355.n209 vssa2 2.54fF $ **FLOATING
C1954 a_537154_685355.n210 vssa2 2.54fF $ **FLOATING
C1955 a_537154_685355.n211 vssa2 9.95fF $ **FLOATING
C1956 a_537154_685355.n212 vssa2 0.38fF $ **FLOATING
C1957 a_537154_685355.n213 vssa2 0.30fF $ **FLOATING
C1958 a_537154_685355.n214 vssa2 1.20fF $ **FLOATING
C1959 a_537154_685355.t65 vssa2 0.42fF
C1960 a_537154_685355.n215 vssa2 0.05fF $ **FLOATING
C1961 a_537154_685355.n216 vssa2 0.43fF $ **FLOATING
C1962 a_537154_685355.n217 vssa2 0.32fF $ **FLOATING
C1963 a_537154_685355.n218 vssa2 0.43fF $ **FLOATING
C1964 a_537154_685355.n219 vssa2 0.01fF $ **FLOATING
C1965 a_537154_685355.n220 vssa2 0.39fF $ **FLOATING
C1966 a_537154_685355.t0 vssa2 0.11fF
C1967 a_537154_685355.n221 vssa2 1.39fF $ **FLOATING
C1968 a_537154_685355.n222 vssa2 0.26fF $ **FLOATING
C1969 a_537154_685355.n223 vssa2 2.90fF $ **FLOATING
C1970 a_537154_685355.n224 vssa2 0.55fF $ **FLOATING
C1971 a_537154_685355.t5 vssa2 0.11fF
C1972 a_537154_685355.n225 vssa2 0.77fF $ **FLOATING
C1973 a_537154_685355.n226 vssa2 0.73fF $ **FLOATING
C1974 a_537154_685355.n227 vssa2 0.71fF $ **FLOATING
C1975 a_537154_685355.n228 vssa2 3.18fF $ **FLOATING
C1976 a_537154_685355.t4 vssa2 0.11fF
C1977 a_537154_685355.n229 vssa2 0.45fF $ **FLOATING
C1978 a_537154_685355.n230 vssa2 0.88fF $ **FLOATING
C1979 a_537154_685355.n231 vssa2 0.72fF $ **FLOATING
C1980 a_537154_685355.n232 vssa2 0.81fF $ **FLOATING
C1981 a_537154_685355.n233 vssa2 3.13fF $ **FLOATING
C1982 a_537154_685355.t29 vssa2 0.11fF
C1983 a_537154_685355.n234 vssa2 0.46fF $ **FLOATING
C1984 a_537154_685355.n235 vssa2 0.86fF $ **FLOATING
C1985 a_537154_685355.t2 vssa2 0.11fF
C1986 a_537154_685355.n236 vssa2 1.37fF $ **FLOATING
C1987 a_537154_685355.t32 vssa2 0.42fF
C1988 a_537154_685355.t44 vssa2 0.42fF
C1989 a_537154_685355.n237 vssa2 0.02fF $ **FLOATING
C1990 a_537154_685355.n238 vssa2 0.43fF $ **FLOATING
C1991 a_537154_685355.n239 vssa2 0.32fF $ **FLOATING
C1992 a_537154_685355.n240 vssa2 0.34fF $ **FLOATING
C1993 a_537154_685355.n241 vssa2 0.01fF $ **FLOATING
C1994 a_537154_685355.n242 vssa2 0.43fF $ **FLOATING
C1995 a_537154_685355.n243 vssa2 0.02fF $ **FLOATING
C1996 a_537154_685355.n244 vssa2 0.87fF $ **FLOATING
C1997 a_537154_685355.n245 vssa2 0.74fF $ **FLOATING
C1998 a_537154_685355.n246 vssa2 0.05fF $ **FLOATING
C1999 a_537154_685355.n247 vssa2 1.23fF $ **FLOATING
C2000 a_537154_685355.t54 vssa2 0.42fF
C2001 a_537154_685355.n248 vssa2 0.36fF $ **FLOATING
C2002 a_537154_685355.n249 vssa2 10.87fF $ **FLOATING
C2003 a_537154_685355.t6 vssa2 0.03fF
C2004 vccd1.t22 vssa2 0.01fF
C2005 vccd1.n0 vssa2 0.24fF $ **FLOATING
C2006 vccd1.t21 vssa2 0.42fF
C2007 vccd1.n1 vssa2 0.41fF $ **FLOATING
C2008 vccd1.n2 vssa2 0.02fF $ **FLOATING
C2009 vccd1.t39 vssa2 0.01fF
C2010 vccd1.n3 vssa2 0.24fF $ **FLOATING
C2011 vccd1.n4 vssa2 0.02fF $ **FLOATING
C2012 vccd1.n5 vssa2 0.02fF $ **FLOATING
C2013 vccd1.n6 vssa2 0.03fF $ **FLOATING
C2014 vccd1.n7 vssa2 0.02fF $ **FLOATING
C2015 vccd1.n8 vssa2 0.02fF $ **FLOATING
C2016 vccd1.n9 vssa2 0.02fF $ **FLOATING
C2017 vccd1.n10 vssa2 0.02fF $ **FLOATING
C2018 vccd1.n11 vssa2 0.02fF $ **FLOATING
C2019 vccd1.n12 vssa2 0.70fF $ **FLOATING
C2020 vccd1.n13 vssa2 0.04fF $ **FLOATING
C2021 vccd1.t1 vssa2 0.01fF
C2022 vccd1.n14 vssa2 0.22fF $ **FLOATING
C2023 vccd1.n15 vssa2 0.01fF $ **FLOATING
C2024 vccd1.n16 vssa2 0.01fF $ **FLOATING
C2025 vccd1.n17 vssa2 0.12fF $ **FLOATING
C2026 vccd1.n18 vssa2 0.12fF $ **FLOATING
C2027 vccd1.n19 vssa2 0.35fF $ **FLOATING
C2028 vccd1.n20 vssa2 0.01fF $ **FLOATING
C2029 vccd1.n21 vssa2 0.01fF $ **FLOATING
C2030 vccd1.t0 vssa2 0.42fF
C2031 vccd1.n22 vssa2 0.35fF $ **FLOATING
C2032 vccd1.n23 vssa2 0.02fF $ **FLOATING
C2033 vccd1.n24 vssa2 0.02fF $ **FLOATING
C2034 vccd1.n25 vssa2 0.02fF $ **FLOATING
C2035 vccd1.n26 vssa2 0.01fF $ **FLOATING
C2036 vccd1.n27 vssa2 0.01fF $ **FLOATING
C2037 vccd1.n28 vssa2 0.01fF $ **FLOATING
C2038 vccd1.n29 vssa2 0.01fF $ **FLOATING
C2039 vccd1.n30 vssa2 0.35fF $ **FLOATING
C2040 vccd1.n31 vssa2 0.01fF $ **FLOATING
C2041 vccd1.n32 vssa2 0.01fF $ **FLOATING
C2042 vccd1.n33 vssa2 0.01fF $ **FLOATING
C2043 vccd1.n34 vssa2 0.01fF $ **FLOATING
C2044 vccd1.n35 vssa2 0.02fF $ **FLOATING
C2045 vccd1.n36 vssa2 0.03fF $ **FLOATING
C2046 vccd1.t33 vssa2 0.35fF
C2047 vccd1.n37 vssa2 0.41fF $ **FLOATING
C2048 vccd1.n38 vssa2 0.02fF $ **FLOATING
C2049 vccd1.n39 vssa2 0.02fF $ **FLOATING
C2050 vccd1.n40 vssa2 0.02fF $ **FLOATING
C2051 vccd1.n41 vssa2 0.02fF $ **FLOATING
C2052 vccd1.n42 vssa2 0.02fF $ **FLOATING
C2053 vccd1.n43 vssa2 0.70fF $ **FLOATING
C2054 vccd1.n44 vssa2 0.04fF $ **FLOATING
C2055 vccd1.t116 vssa2 0.01fF
C2056 vccd1.n45 vssa2 0.19fF $ **FLOATING
C2057 vccd1.n46 vssa2 0.02fF $ **FLOATING
C2058 vccd1.t47 vssa2 0.30fF
C2059 vccd1.n47 vssa2 0.20fF $ **FLOATING
C2060 vccd1.n48 vssa2 0.01fF $ **FLOATING
C2061 vccd1.n49 vssa2 -0.17fF $ **FLOATING
C2062 vccd1.n50 vssa2 0.07fF $ **FLOATING
C2063 vccd1.n51 vssa2 0.07fF $ **FLOATING
C2064 vccd1.n52 vssa2 0.01fF $ **FLOATING
C2065 vccd1.n53 vssa2 0.01fF $ **FLOATING
C2066 vccd1.n54 vssa2 0.02fF $ **FLOATING
C2067 vccd1.n55 vssa2 0.02fF $ **FLOATING
C2068 vccd1.n56 vssa2 0.35fF $ **FLOATING
C2069 vccd1.n57 vssa2 0.01fF $ **FLOATING
C2070 vccd1.n58 vssa2 0.01fF $ **FLOATING
C2071 vccd1.n59 vssa2 0.01fF $ **FLOATING
C2072 vccd1.n60 vssa2 0.01fF $ **FLOATING
C2073 vccd1.n61 vssa2 0.01fF $ **FLOATING
C2074 vccd1.n62 vssa2 0.01fF $ **FLOATING
C2075 vccd1.n63 vssa2 0.01fF $ **FLOATING
C2076 vccd1.t48 vssa2 0.01fF
C2077 vccd1.n64 vssa2 0.19fF $ **FLOATING
C2078 vccd1.n65 vssa2 1.04fF $ **FLOATING
C2079 vccd1.n66 vssa2 0.01fF $ **FLOATING
C2080 vccd1.n67 vssa2 0.02fF $ **FLOATING
C2081 vccd1.n68 vssa2 0.01fF $ **FLOATING
C2082 vccd1.n69 vssa2 0.02fF $ **FLOATING
C2083 vccd1.n70 vssa2 0.57fF $ **FLOATING
C2084 vccd1.n71 vssa2 0.03fF $ **FLOATING
C2085 vccd1.n72 vssa2 0.00fF $ **FLOATING
C2086 vccd1.t10 vssa2 0.41fF
C2087 vccd1.n73 vssa2 0.43fF $ **FLOATING
C2088 vccd1.n74 vssa2 0.02fF $ **FLOATING
C2089 vccd1.t11 vssa2 0.01fF
C2090 vccd1.n75 vssa2 0.23fF $ **FLOATING
C2091 vccd1.n76 vssa2 0.02fF $ **FLOATING
C2092 vccd1.n77 vssa2 0.02fF $ **FLOATING
C2093 vccd1.n78 vssa2 0.02fF $ **FLOATING
C2094 vccd1.n79 vssa2 0.03fF $ **FLOATING
C2095 vccd1.t40 vssa2 0.01fF
C2096 vccd1.n80 vssa2 0.24fF $ **FLOATING
C2097 vccd1.n81 vssa2 1.78fF $ **FLOATING
C2098 vccd1.n82 vssa2 0.00fF $ **FLOATING
C2099 vccd1.t115 vssa2 0.01fF
C2100 vccd1.n83 vssa2 0.02fF $ **FLOATING
C2101 vccd1.n84 vssa2 0.03fF $ **FLOATING
C2102 vccd1.n85 vssa2 0.02fF $ **FLOATING
C2103 vccd1.n86 vssa2 0.02fF $ **FLOATING
C2104 vccd1.t34 vssa2 0.01fF
C2105 vccd1.n87 vssa2 2.30fF $ **FLOATING
C2106 vccd1.t16 vssa2 0.01fF
C2107 vccd1.n88 vssa2 0.22fF $ **FLOATING
C2108 vccd1.n89 vssa2 1.90fF $ **FLOATING
C2109 vccd1.n90 vssa2 0.00fF $ **FLOATING
C2110 vccd1.n91 vssa2 1.71fF $ **FLOATING
C2111 vccd1.t49 vssa2 0.01fF
C2112 vccd1.n92 vssa2 0.01fF $ **FLOATING
C2113 vccd1.n93 vssa2 0.01fF $ **FLOATING
C2114 vccd1.n94 vssa2 0.01fF $ **FLOATING
C2115 vccd1.n95 vssa2 0.02fF $ **FLOATING
C2116 vccd1.n96 vssa2 0.01fF $ **FLOATING
C2117 vccd1.n97 vssa2 0.02fF $ **FLOATING
C2118 vccd1.n98 vssa2 0.57fF $ **FLOATING
C2119 vccd1.n99 vssa2 0.03fF $ **FLOATING
C2120 vccd1.n100 vssa2 0.00fF $ **FLOATING
C2121 vccd1.n101 vssa2 0.01fF $ **FLOATING
C2122 vccd1.n102 vssa2 0.47fF $ **FLOATING
C2123 vccd1.n103 vssa2 0.54fF $ **FLOATING
C2124 vccd1.n104 vssa2 0.02fF $ **FLOATING
C2125 vccd1.t8 vssa2 0.19fF
C2126 vccd1.n105 vssa2 0.29fF $ **FLOATING
C2127 vccd1.n106 vssa2 0.01fF $ **FLOATING
C2128 vccd1.n107 vssa2 0.01fF $ **FLOATING
C2129 vccd1.n108 vssa2 -0.01fF $ **FLOATING
C2130 vccd1.n109 vssa2 0.02fF $ **FLOATING
C2131 vccd1.n110 vssa2 0.02fF $ **FLOATING
C2132 vccd1.n111 vssa2 0.38fF $ **FLOATING
C2133 vccd1.n112 vssa2 0.01fF $ **FLOATING
C2134 vccd1.n113 vssa2 0.01fF $ **FLOATING
C2135 vccd1.n114 vssa2 0.07fF $ **FLOATING
C2136 vccd1.n115 vssa2 0.07fF $ **FLOATING
C2137 vccd1.n116 vssa2 0.01fF $ **FLOATING
C2138 vccd1.n117 vssa2 0.01fF $ **FLOATING
C2139 vccd1.n118 vssa2 0.01fF $ **FLOATING
C2140 vccd1.t9 vssa2 0.01fF
C2141 vccd1.n119 vssa2 0.39fF $ **FLOATING
C2142 vccd1.n120 vssa2 0.81fF $ **FLOATING
C2143 vccd1.t59 vssa2 0.01fF
C2144 vccd1.t54 vssa2 0.01fF
C2145 vccd1.n121 vssa2 0.15fF $ **FLOATING
C2146 vccd1.n122 vssa2 0.26fF $ **FLOATING
C2147 vccd1.t12 vssa2 0.01fF
C2148 vccd1.t45 vssa2 0.01fF
C2149 vccd1.n123 vssa2 0.14fF $ **FLOATING
C2150 vccd1.n124 vssa2 0.23fF $ **FLOATING
C2151 vccd1.t13 vssa2 0.01fF
C2152 vccd1.t17 vssa2 0.01fF
C2153 vccd1.n125 vssa2 0.15fF $ **FLOATING
C2154 vccd1.n126 vssa2 0.26fF $ **FLOATING
C2155 vccd1.t41 vssa2 0.01fF
C2156 vccd1.t3 vssa2 0.01fF
C2157 vccd1.n127 vssa2 0.14fF $ **FLOATING
C2158 vccd1.n128 vssa2 0.24fF $ **FLOATING
C2159 vccd1.t57 vssa2 0.01fF
C2160 vccd1.t32 vssa2 0.01fF
C2161 vccd1.n129 vssa2 0.15fF $ **FLOATING
C2162 vccd1.n130 vssa2 0.12fF $ **FLOATING
C2163 vccd1.n131 vssa2 0.08fF $ **FLOATING
C2164 vccd1.n132 vssa2 0.06fF $ **FLOATING
C2165 vccd1.t37 vssa2 0.01fF
C2166 vccd1.n133 vssa2 0.14fF $ **FLOATING
C2167 vccd1.t58 vssa2 0.01fF
C2168 vccd1.n134 vssa2 0.23fF $ **FLOATING
C2169 vccd1.t46 vssa2 0.01fF
C2170 vccd1.t42 vssa2 0.05fF
C2171 vccd1.n135 vssa2 0.37fF $ **FLOATING
C2172 vccd1.t28 vssa2 0.01fF
C2173 vccd1.t61 vssa2 0.05fF
C2174 vccd1.n136 vssa2 0.34fF $ **FLOATING
C2175 vccd1.n137 vssa2 0.06fF $ **FLOATING
C2176 vccd1.n138 vssa2 1.42fF $ **FLOATING
C2177 vccd1.n139 vssa2 1.08fF $ **FLOATING
C2178 vccd1.n141 vssa2 1.03fF $ **FLOATING
C2179 vccd1.n142 vssa2 1.07fF $ **FLOATING
C2180 vccd1.n143 vssa2 0.22fF $ **FLOATING
C2181 vccd1.n144 vssa2 0.22fF $ **FLOATING
C2182 vccd1.n145 vssa2 0.03fF $ **FLOATING
C2183 vccd1.t43 vssa2 0.01fF
C2184 vccd1.t52 vssa2 0.01fF
C2185 vccd1.n146 vssa2 0.15fF $ **FLOATING
C2186 vccd1.n147 vssa2 0.25fF $ **FLOATING
C2187 vccd1.t62 vssa2 0.01fF
C2188 vccd1.t53 vssa2 0.01fF
C2189 vccd1.n148 vssa2 0.14fF $ **FLOATING
C2190 vccd1.n149 vssa2 0.22fF $ **FLOATING
C2191 vccd1.n150 vssa2 0.27fF $ **FLOATING
C2192 vccd1.t101 vssa2 0.01fF
C2193 vccd1.n152 vssa2 0.14fF $ **FLOATING
C2194 vccd1.t105 vssa2 0.01fF
C2195 vccd1.n153 vssa2 0.19fF $ **FLOATING
C2196 vccd1.n154 vssa2 0.07fF $ **FLOATING
C2197 vccd1.t94 vssa2 0.01fF
C2198 vccd1.t75 vssa2 0.05fF
C2199 vccd1.n155 vssa2 0.28fF $ **FLOATING
C2200 vccd1.n156 vssa2 0.77fF $ **FLOATING
C2201 vccd1.t66 vssa2 1.51fF
C2202 vccd1.n157 vssa2 1.57fF $ **FLOATING
C2203 vccd1.t2 vssa2 2.87fF
C2204 vccd1.n158 vssa2 1.50fF $ **FLOATING
C2205 vccd1.n159 vssa2 2.76fF $ **FLOATING
C2206 vccd1.n160 vssa2 0.00fF $ **FLOATING
C2207 vccd1.n161 vssa2 0.00fF $ **FLOATING
C2208 vccd1.n162 vssa2 0.00fF $ **FLOATING
C2209 vccd1.t79 vssa2 2.52fF
C2210 vccd1.n163 vssa2 0.68fF $ **FLOATING
C2211 vccd1.n164 vssa2 0.07fF $ **FLOATING
C2212 vccd1.t90 vssa2 0.01fF
C2213 vccd1.n165 vssa2 0.14fF $ **FLOATING
C2214 vccd1.t81 vssa2 0.05fF
C2215 vccd1.t110 vssa2 0.01fF
C2216 vccd1.n166 vssa2 0.39fF $ **FLOATING
C2217 vccd1.t112 vssa2 0.05fF
C2218 vccd1.t102 vssa2 0.01fF
C2219 vccd1.t69 vssa2 0.01fF
C2220 vccd1.n167 vssa2 0.14fF $ **FLOATING
C2221 vccd1.n168 vssa2 0.28fF $ **FLOATING
C2222 vccd1.n169 vssa2 0.75fF $ **FLOATING
C2223 vccd1.t89 vssa2 0.05fF
C2224 vccd1.t98 vssa2 0.01fF
C2225 vccd1.n170 vssa2 0.14fF $ **FLOATING
C2226 vccd1.t76 vssa2 0.01fF
C2227 vccd1.n171 vssa2 0.35fF $ **FLOATING
C2228 vccd1.t113 vssa2 0.01fF
C2229 vccd1.t108 vssa2 0.01fF
C2230 vccd1.n172 vssa2 0.14fF $ **FLOATING
C2231 vccd1.n173 vssa2 0.30fF $ **FLOATING
C2232 vccd1.t83 vssa2 0.01fF
C2233 vccd1.t70 vssa2 0.01fF
C2234 vccd1.n174 vssa2 0.14fF $ **FLOATING
C2235 vccd1.n175 vssa2 0.25fF $ **FLOATING
C2236 vccd1.t100 vssa2 0.01fF
C2237 vccd1.t85 vssa2 0.05fF
C2238 vccd1.n176 vssa2 0.39fF $ **FLOATING
C2239 vccd1.t106 vssa2 0.01fF
C2240 vccd1.t96 vssa2 0.05fF
C2241 vccd1.n177 vssa2 0.35fF $ **FLOATING
C2242 vccd1.n178 vssa2 0.07fF $ **FLOATING
C2243 vccd1.n179 vssa2 0.79fF $ **FLOATING
C2244 vccd1.n180 vssa2 0.36fF $ **FLOATING
C2245 vccd1.n181 vssa2 0.01fF $ **FLOATING
C2246 vccd1.n182 vssa2 0.36fF $ **FLOATING
C2247 vccd1.n183 vssa2 0.35fF $ **FLOATING
C2248 vccd1.n184 vssa2 0.07fF $ **FLOATING
C2249 vccd1.n185 vssa2 0.45fF $ **FLOATING
C2250 vccd1.n186 vssa2 0.07fF $ **FLOATING
C2251 vccd1.n187 vssa2 0.03fF $ **FLOATING
C2252 vccd1.t107 vssa2 0.01fF
C2253 vccd1.n188 vssa2 0.13fF $ **FLOATING
C2254 vccd1.t111 vssa2 0.01fF
C2255 vccd1.n189 vssa2 0.05fF $ **FLOATING
C2256 vccd1.n190 vssa2 0.03fF $ **FLOATING
C2257 vccd1.n191 vssa2 0.06fF $ **FLOATING
C2258 vccd1.n192 vssa2 0.38fF $ **FLOATING
C2259 vccd1.n194 vssa2 0.40fF $ **FLOATING
C2260 vccd1.t87 vssa2 0.01fF
C2261 vccd1.n195 vssa2 0.13fF $ **FLOATING
C2262 vccd1.n196 vssa2 0.03fF $ **FLOATING
C2263 vccd1.t109 vssa2 0.01fF
C2264 vccd1.n197 vssa2 0.05fF $ **FLOATING
C2265 vccd1.t78 vssa2 0.05fF
C2266 vccd1.n198 vssa2 0.12fF $ **FLOATING
C2267 vccd1.n199 vssa2 0.12fF $ **FLOATING
C2268 vccd1.n200 vssa2 0.89fF $ **FLOATING
C2269 vccd1.n201 vssa2 0.22fF $ **FLOATING
C2270 vccd1.n202 vssa2 1.57fF $ **FLOATING
C2271 vccd1.t35 vssa2 2.83fF
C2272 vccd1.n203 vssa2 1.49fF $ **FLOATING
C2273 vccd1.n204 vssa2 0.02fF $ **FLOATING
C2274 vccd1.n205 vssa2 0.00fF $ **FLOATING
C2275 vccd1.n207 vssa2 0.05fF $ **FLOATING
C2276 vccd1.n208 vssa2 0.05fF $ **FLOATING
C2277 vccd1.t92 vssa2 0.05fF
C2278 vccd1.t104 vssa2 0.01fF
C2279 vccd1.n209 vssa2 0.05fF $ **FLOATING
C2280 vccd1.n210 vssa2 0.12fF $ **FLOATING
C2281 vccd1.t103 vssa2 0.01fF
C2282 vccd1.n211 vssa2 0.05fF $ **FLOATING
C2283 vccd1.n212 vssa2 0.03fF $ **FLOATING
C2284 vccd1.t91 vssa2 0.05fF
C2285 vccd1.n213 vssa2 0.12fF $ **FLOATING
C2286 vccd1.t84 vssa2 0.05fF
C2287 vccd1.n214 vssa2 0.12fF $ **FLOATING
C2288 vccd1.t99 vssa2 0.01fF
C2289 vccd1.n215 vssa2 0.05fF $ **FLOATING
C2290 vccd1.n216 vssa2 0.03fF $ **FLOATING
C2291 vccd1.n217 vssa2 0.06fF $ **FLOATING
C2292 vccd1.n218 vssa2 0.06fF $ **FLOATING
C2293 vccd1.n219 vssa2 0.98fF $ **FLOATING
C2294 vccd1.n220 vssa2 0.15fF $ **FLOATING
C2295 vccd1.n221 vssa2 0.04fF $ **FLOATING
C2296 vccd1.n222 vssa2 0.11fF $ **FLOATING
C2297 vccd1.t18 vssa2 2.86fF
C2298 vccd1.n223 vssa2 0.22fF $ **FLOATING
C2299 vccd1.t93 vssa2 0.21fF
C2300 vccd1.n224 vssa2 1.57fF $ **FLOATING
C2301 vccd1.n225 vssa2 0.02fF $ **FLOATING
C2302 vccd1.n226 vssa2 0.00fF $ **FLOATING
C2303 vccd1.n228 vssa2 0.03fF $ **FLOATING
C2304 vccd1.n229 vssa2 0.18fF $ **FLOATING
C2305 vccd1.n230 vssa2 0.06fF $ **FLOATING
C2306 vccd1.n231 vssa2 0.14fF $ **FLOATING
C2307 vccd1.n232 vssa2 0.18fF $ **FLOATING
C2308 vccd1.n233 vssa2 0.18fF $ **FLOATING
C2309 vccd1.n234 vssa2 0.18fF $ **FLOATING
C2310 vccd1.n235 vssa2 0.24fF $ **FLOATING
C2311 vccd1.n236 vssa2 0.24fF $ **FLOATING
C2312 vccd1.n237 vssa2 0.24fF $ **FLOATING
C2313 vccd1.n238 vssa2 0.24fF $ **FLOATING
C2314 vccd1.n239 vssa2 2.38fF $ **FLOATING
C2315 vccd1.t25 vssa2 4.56fF
C2316 vccd1.n240 vssa2 0.09fF $ **FLOATING
C2317 vccd1.n241 vssa2 0.09fF $ **FLOATING
C2318 vccd1.n242 vssa2 3.32fF $ **FLOATING
C2319 vccd1.t27 vssa2 1.65fF
C2320 vccd1.t74 vssa2 2.13fF
C2321 vccd1.n243 vssa2 0.03fF $ **FLOATING
C2322 vccd1.n244 vssa2 1.57fF $ **FLOATING
C2323 vccd1.t31 vssa2 2.20fF
C2324 vccd1.n245 vssa2 1.48fF $ **FLOATING
C2325 vccd1.n246 vssa2 0.02fF $ **FLOATING
C2326 vccd1.n247 vssa2 1.22fF $ **FLOATING
C2327 vccd1.n248 vssa2 0.02fF $ **FLOATING
C2328 vccd1.n249 vssa2 0.02fF $ **FLOATING
C2329 vccd1.t68 vssa2 1.51fF
C2330 vccd1.t6 vssa2 2.82fF
C2331 vccd1.n251 vssa2 1.53fF $ **FLOATING
C2332 vccd1.n252 vssa2 0.02fF $ **FLOATING
C2333 vccd1.t67 vssa2 0.01fF
C2334 vccd1.n253 vssa2 0.13fF $ **FLOATING
C2335 vccd1.t82 vssa2 0.01fF
C2336 vccd1.n254 vssa2 0.05fF $ **FLOATING
C2337 vccd1.n255 vssa2 0.03fF $ **FLOATING
C2338 vccd1.t114 vssa2 0.01fF
C2339 vccd1.n256 vssa2 0.13fF $ **FLOATING
C2340 vccd1.t80 vssa2 0.01fF
C2341 vccd1.n257 vssa2 0.05fF $ **FLOATING
C2342 vccd1.n258 vssa2 0.03fF $ **FLOATING
C2343 vccd1.n259 vssa2 0.04fF $ **FLOATING
C2344 vccd1.n260 vssa2 0.05fF $ **FLOATING
C2345 vccd1.n261 vssa2 0.09fF $ **FLOATING
C2346 vccd1.n262 vssa2 0.03fF $ **FLOATING
C2347 vccd1.n263 vssa2 0.11fF $ **FLOATING
C2348 vccd1.n264 vssa2 0.91fF $ **FLOATING
C2349 vccd1.n265 vssa2 0.02fF $ **FLOATING
C2350 vccd1.n266 vssa2 0.03fF $ **FLOATING
C2351 vccd1.n267 vssa2 0.18fF $ **FLOATING
C2352 vccd1.n268 vssa2 0.18fF $ **FLOATING
C2353 vccd1.n269 vssa2 0.18fF $ **FLOATING
C2354 vccd1.n270 vssa2 0.06fF $ **FLOATING
C2355 vccd1.n271 vssa2 0.14fF $ **FLOATING
C2356 vccd1.n272 vssa2 0.18fF $ **FLOATING
C2357 vccd1.n273 vssa2 0.09fF $ **FLOATING
C2358 vccd1.n274 vssa2 0.09fF $ **FLOATING
C2359 vccd1.n275 vssa2 3.33fF $ **FLOATING
C2360 vccd1.t14 vssa2 1.65fF
C2361 vccd1.t77 vssa2 2.22fF
C2362 vccd1.n276 vssa2 0.03fF $ **FLOATING
C2363 vccd1.n277 vssa2 1.50fF $ **FLOATING
C2364 vccd1.t4 vssa2 2.21fF
C2365 vccd1.t71 vssa2 0.21fF
C2366 vccd1.n278 vssa2 1.57fF $ **FLOATING
C2367 vccd1.n279 vssa2 0.02fF $ **FLOATING
C2368 vccd1.t95 vssa2 0.01fF
C2369 vccd1.n280 vssa2 0.13fF $ **FLOATING
C2370 vccd1.n281 vssa2 0.03fF $ **FLOATING
C2371 vccd1.t72 vssa2 0.01fF
C2372 vccd1.n282 vssa2 0.05fF $ **FLOATING
C2373 vccd1.t86 vssa2 0.05fF
C2374 vccd1.n283 vssa2 0.12fF $ **FLOATING
C2375 vccd1.t97 vssa2 0.01fF
C2376 vccd1.n284 vssa2 0.13fF $ **FLOATING
C2377 vccd1.n285 vssa2 0.03fF $ **FLOATING
C2378 vccd1.n286 vssa2 0.15fF $ **FLOATING
C2379 vccd1.t73 vssa2 0.01fF
C2380 vccd1.n287 vssa2 0.05fF $ **FLOATING
C2381 vccd1.t88 vssa2 0.05fF
C2382 vccd1.n288 vssa2 0.12fF $ **FLOATING
C2383 vccd1.n289 vssa2 0.11fF $ **FLOATING
C2384 vccd1.n290 vssa2 1.37fF $ **FLOATING
C2385 vccd1.n291 vssa2 1.48fF $ **FLOATING
C2386 vccd1.n292 vssa2 0.72fF $ **FLOATING
C2387 vccd1.n293 vssa2 0.71fF $ **FLOATING
C2388 vccd1.n294 vssa2 3.63fF $ **FLOATING
C2389 vccd1.t23 vssa2 4.63fF
C2390 vccd1.n295 vssa2 2.47fF $ **FLOATING
C2391 vccd1.n296 vssa2 0.22fF $ **FLOATING
C2392 vccd1.n297 vssa2 0.22fF $ **FLOATING
C2393 vccd1.n298 vssa2 0.03fF $ **FLOATING
C2394 vccd1.n299 vssa2 0.06fF $ **FLOATING
C2395 vccd1.t63 vssa2 0.01fF
C2396 vccd1.t44 vssa2 0.05fF
C2397 vccd1.n300 vssa2 0.31fF $ **FLOATING
C2398 vccd1.n301 vssa2 0.72fF $ **FLOATING
C2399 vccd1.t26 vssa2 0.05fF
C2400 vccd1.t64 vssa2 0.01fF
C2401 vccd1.n302 vssa2 0.41fF $ **FLOATING
C2402 vccd1.n303 vssa2 0.52fF $ **FLOATING
C2403 vccd1.t51 vssa2 0.01fF
C2404 vccd1.n304 vssa2 0.15fF $ **FLOATING
C2405 vccd1.t19 vssa2 0.01fF
C2406 vccd1.n305 vssa2 0.29fF $ **FLOATING
C2407 vccd1.t65 vssa2 0.01fF
C2408 vccd1.t50 vssa2 0.01fF
C2409 vccd1.n306 vssa2 0.15fF $ **FLOATING
C2410 vccd1.n307 vssa2 0.20fF $ **FLOATING
C2411 vccd1.n308 vssa2 1.03fF $ **FLOATING
C2412 vccd1.t30 vssa2 0.01fF
C2413 vccd1.n310 vssa2 0.15fF $ **FLOATING
C2414 vccd1.t55 vssa2 0.01fF
C2415 vccd1.n311 vssa2 0.29fF $ **FLOATING
C2416 vccd1.t7 vssa2 0.01fF
C2417 vccd1.t29 vssa2 0.01fF
C2418 vccd1.n312 vssa2 0.15fF $ **FLOATING
C2419 vccd1.n313 vssa2 0.20fF $ **FLOATING
C2420 vccd1.n314 vssa2 0.98fF $ **FLOATING
C2421 vccd1.t36 vssa2 0.01fF
C2422 vccd1.n315 vssa2 0.15fF $ **FLOATING
C2423 vccd1.t20 vssa2 0.01fF
C2424 vccd1.n316 vssa2 0.26fF $ **FLOATING
C2425 vccd1.t38 vssa2 0.01fF
C2426 vccd1.n317 vssa2 0.15fF $ **FLOATING
C2427 vccd1.t5 vssa2 0.01fF
C2428 vccd1.n318 vssa2 0.29fF $ **FLOATING
C2429 vccd1.n319 vssa2 1.01fF $ **FLOATING
C2430 vccd1.t60 vssa2 0.01fF
C2431 vccd1.n320 vssa2 0.15fF $ **FLOATING
C2432 vccd1.t24 vssa2 0.01fF
C2433 vccd1.n321 vssa2 0.28fF $ **FLOATING
C2434 vccd1.t56 vssa2 0.01fF
C2435 vccd1.t15 vssa2 0.01fF
C2436 vccd1.n322 vssa2 0.15fF $ **FLOATING
C2437 vccd1.n323 vssa2 0.19fF $ **FLOATING
C2438 vccd1.n324 vssa2 10.32fF $ **FLOATING
C2439 vccd1.n325 vssa2 115.38fF $ **FLOATING
C2440 vccd1.n326 vssa2 15.53fF $ **FLOATING
C2441 vccd1.n327 vssa2 479.87fF $ **FLOATING
C2442 vccd1.n328 vssa2 15.67fF $ **FLOATING
C2443 a_540271_687858.n0 vssa2 1.35fF $ **FLOATING
C2444 a_540271_687858.n1 vssa2 1.19fF $ **FLOATING
C2445 a_540271_687858.n2 vssa2 0.95fF $ **FLOATING
C2446 a_540271_687858.n3 vssa2 1.56fF $ **FLOATING
C2447 a_540271_687858.n4 vssa2 1.38fF $ **FLOATING
C2448 a_540271_687858.n5 vssa2 0.09fF $ **FLOATING
C2449 a_540271_687858.n6 vssa2 1.43fF $ **FLOATING
C2450 a_540271_687858.n7 vssa2 1.16fF $ **FLOATING
C2451 a_540271_687858.n8 vssa2 2.94fF $ **FLOATING
C2452 a_540271_687858.n9 vssa2 5.71fF $ **FLOATING
C2453 a_540271_687858.n10 vssa2 5.64fF $ **FLOATING
C2454 a_540271_687858.n11 vssa2 0.79fF $ **FLOATING
C2455 a_540271_687858.n12 vssa2 1.52fF $ **FLOATING
C2456 a_540271_687858.n13 vssa2 0.09fF $ **FLOATING
C2457 a_540271_687858.n14 vssa2 5.57fF $ **FLOATING
C2458 a_540271_687858.n15 vssa2 1.38fF $ **FLOATING
C2459 a_540271_687858.n16 vssa2 1.38fF $ **FLOATING
C2460 a_540271_687858.n17 vssa2 1.36fF $ **FLOATING
C2461 a_540271_687858.n18 vssa2 1.56fF $ **FLOATING
C2462 a_540271_687858.n19 vssa2 1.81fF $ **FLOATING
C2463 a_540271_687858.t62 vssa2 0.37fF
C2464 a_540271_687858.t50 vssa2 0.37fF
C2465 a_540271_687858.t66 vssa2 0.37fF
C2466 a_540271_687858.n20 vssa2 1.09fF $ **FLOATING
C2467 a_540271_687858.n21 vssa2 0.38fF $ **FLOATING
C2468 a_540271_687858.n22 vssa2 0.68fF $ **FLOATING
C2469 a_540271_687858.t14 vssa2 0.09fF
C2470 a_540271_687858.t13 vssa2 0.36fF
C2471 a_540271_687858.n23 vssa2 0.50fF $ **FLOATING
C2472 a_540271_687858.n24 vssa2 1.01fF $ **FLOATING
C2473 a_540271_687858.n25 vssa2 1.78fF $ **FLOATING
C2474 a_540271_687858.n26 vssa2 2.71fF $ **FLOATING
C2475 a_540271_687858.n27 vssa2 0.26fF $ **FLOATING
C2476 a_540271_687858.n28 vssa2 0.47fF $ **FLOATING
C2477 a_540271_687858.t8 vssa2 0.09fF
C2478 a_540271_687858.t7 vssa2 0.36fF
C2479 a_540271_687858.n29 vssa2 1.01fF $ **FLOATING
C2480 a_540271_687858.n30 vssa2 2.93fF $ **FLOATING
C2481 a_540271_687858.n31 vssa2 0.26fF $ **FLOATING
C2482 a_540271_687858.n32 vssa2 0.82fF $ **FLOATING
C2483 a_540271_687858.t18 vssa2 0.28fF
C2484 a_540271_687858.t17 vssa2 0.36fF
C2485 a_540271_687858.n33 vssa2 0.02fF $ **FLOATING
C2486 a_540271_687858.n34 vssa2 0.08fF $ **FLOATING
C2487 a_540271_687858.n35 vssa2 0.50fF $ **FLOATING
C2488 a_540271_687858.n36 vssa2 0.11fF $ **FLOATING
C2489 a_540271_687858.t6 vssa2 0.09fF
C2490 a_540271_687858.n37 vssa2 0.02fF $ **FLOATING
C2491 a_540271_687858.t5 vssa2 0.36fF
C2492 a_540271_687858.t16 vssa2 0.09fF
C2493 a_540271_687858.n38 vssa2 0.06fF $ **FLOATING
C2494 a_540271_687858.n39 vssa2 0.38fF $ **FLOATING
C2495 a_540271_687858.n40 vssa2 0.28fF $ **FLOATING
C2496 a_540271_687858.t10 vssa2 0.09fF
C2497 a_540271_687858.n41 vssa2 1.11fF $ **FLOATING
C2498 a_540271_687858.t9 vssa2 0.36fF
C2499 a_540271_687858.n42 vssa2 1.51fF $ **FLOATING
C2500 a_540271_687858.n43 vssa2 0.02fF $ **FLOATING
C2501 a_540271_687858.n44 vssa2 0.56fF $ **FLOATING
C2502 a_540271_687858.t34 vssa2 0.09fF
C2503 a_540271_687858.t33 vssa2 0.36fF
C2504 a_540271_687858.n45 vssa2 1.44fF $ **FLOATING
C2505 a_540271_687858.n46 vssa2 1.12fF $ **FLOATING
C2506 a_540271_687858.t15 vssa2 0.36fF
C2507 a_540271_687858.n47 vssa2 0.77fF $ **FLOATING
C2508 a_540271_687858.n48 vssa2 0.62fF $ **FLOATING
C2509 a_540271_687858.n49 vssa2 0.02fF $ **FLOATING
C2510 a_540271_687858.n50 vssa2 0.41fF $ **FLOATING
C2511 a_540271_687858.n51 vssa2 1.34fF $ **FLOATING
C2512 a_540271_687858.t24 vssa2 0.09fF
C2513 a_540271_687858.n52 vssa2 0.02fF $ **FLOATING
C2514 a_540271_687858.t40 vssa2 0.09fF
C2515 a_540271_687858.n53 vssa2 0.02fF $ **FLOATING
C2516 a_540271_687858.n54 vssa2 0.08fF $ **FLOATING
C2517 a_540271_687858.n55 vssa2 0.02fF $ **FLOATING
C2518 a_540271_687858.n56 vssa2 0.76fF $ **FLOATING
C2519 a_540271_687858.n57 vssa2 0.38fF $ **FLOATING
C2520 a_540271_687858.n58 vssa2 0.62fF $ **FLOATING
C2521 a_540271_687858.t32 vssa2 0.09fF
C2522 a_540271_687858.t31 vssa2 0.36fF
C2523 a_540271_687858.n59 vssa2 0.51fF $ **FLOATING
C2524 a_540271_687858.n60 vssa2 0.26fF $ **FLOATING
C2525 a_540271_687858.n61 vssa2 0.15fF $ **FLOATING
C2526 a_540271_687858.n62 vssa2 0.50fF $ **FLOATING
C2527 a_540271_687858.n63 vssa2 1.01fF $ **FLOATING
C2528 a_540271_687858.t39 vssa2 0.36fF
C2529 a_540271_687858.n64 vssa2 0.69fF $ **FLOATING
C2530 a_540271_687858.n65 vssa2 0.52fF $ **FLOATING
C2531 a_540271_687858.t23 vssa2 0.36fF
C2532 a_540271_687858.t43 vssa2 0.36fF
C2533 a_540271_687858.n66 vssa2 0.50fF $ **FLOATING
C2534 a_540271_687858.n67 vssa2 0.57fF $ **FLOATING
C2535 a_540271_687858.t26 vssa2 0.09fF
C2536 a_540271_687858.n68 vssa2 0.50fF $ **FLOATING
C2537 a_540271_687858.n69 vssa2 0.57fF $ **FLOATING
C2538 a_540271_687858.n70 vssa2 0.38fF $ **FLOATING
C2539 a_540271_687858.n71 vssa2 1.10fF $ **FLOATING
C2540 a_540271_687858.t55 vssa2 0.36fF
C2541 a_540271_687858.n72 vssa2 0.05fF $ **FLOATING
C2542 a_540271_687858.n73 vssa2 1.17fF $ **FLOATING
C2543 a_540271_687858.t51 vssa2 0.36fF
C2544 a_540271_687858.n74 vssa2 0.03fF $ **FLOATING
C2545 a_540271_687858.t67 vssa2 0.36fF
C2546 a_540271_687858.n75 vssa2 0.03fF $ **FLOATING
C2547 a_540271_687858.t46 vssa2 0.09fF
C2548 a_540271_687858.n76 vssa2 1.04fF $ **FLOATING
C2549 a_540271_687858.t45 vssa2 0.36fF
C2550 a_540271_687858.n77 vssa2 0.50fF $ **FLOATING
C2551 a_540271_687858.n78 vssa2 0.59fF $ **FLOATING
C2552 a_540271_687858.n79 vssa2 0.32fF $ **FLOATING
C2553 a_540271_687858.t2 vssa2 0.09fF
C2554 a_540271_687858.t47 vssa2 0.51fF
C2555 a_540271_687858.n80 vssa2 1.45fF $ **FLOATING
C2556 a_540271_687858.t1 vssa2 0.09fF
C2557 a_540271_687858.n81 vssa2 0.73fF $ **FLOATING
C2558 a_540271_687858.n82 vssa2 5.27fF $ **FLOATING
C2559 a_540271_687858.t20 vssa2 0.09fF
C2560 a_540271_687858.t19 vssa2 0.36fF
C2561 a_540271_687858.t58 vssa2 0.36fF
C2562 a_540271_687858.n83 vssa2 0.03fF $ **FLOATING
C2563 a_540271_687858.n84 vssa2 0.41fF $ **FLOATING
C2564 a_540271_687858.t65 vssa2 0.36fF
C2565 a_540271_687858.n85 vssa2 0.03fF $ **FLOATING
C2566 a_540271_687858.n86 vssa2 1.14fF $ **FLOATING
C2567 a_540271_687858.t61 vssa2 0.36fF
C2568 a_540271_687858.n87 vssa2 0.03fF $ **FLOATING
C2569 a_540271_687858.n88 vssa2 0.50fF $ **FLOATING
C2570 a_540271_687858.n89 vssa2 1.01fF $ **FLOATING
C2571 a_540271_687858.t25 vssa2 0.36fF
C2572 a_540271_687858.t69 vssa2 0.36fF
C2573 a_540271_687858.n90 vssa2 0.05fF $ **FLOATING
C2574 a_540271_687858.t64 vssa2 0.36fF
C2575 a_540271_687858.n91 vssa2 0.05fF $ **FLOATING
C2576 a_540271_687858.t52 vssa2 0.36fF
C2577 a_540271_687858.n92 vssa2 0.05fF $ **FLOATING
C2578 a_540271_687858.t56 vssa2 0.36fF
C2579 a_540271_687858.n93 vssa2 0.05fF $ **FLOATING
C2580 a_540271_687858.t54 vssa2 0.36fF
C2581 a_540271_687858.n94 vssa2 0.05fF $ **FLOATING
C2582 a_540271_687858.n95 vssa2 1.14fF $ **FLOATING
C2583 a_540271_687858.t49 vssa2 0.36fF
C2584 a_540271_687858.n96 vssa2 0.00fF $ **FLOATING
C2585 a_540271_687858.n97 vssa2 1.34fF $ **FLOATING
C2586 a_540271_687858.n98 vssa2 0.31fF $ **FLOATING
C2587 a_540271_687858.n99 vssa2 0.02fF $ **FLOATING
C2588 a_540271_687858.t44 vssa2 0.09fF
C2589 a_540271_687858.n100 vssa2 0.42fF $ **FLOATING
C2590 a_540271_687858.n101 vssa2 1.04fF $ **FLOATING
C2591 a_540271_687858.n102 vssa2 0.02fF $ **FLOATING
C2592 a_540271_687858.t4 vssa2 0.09fF
C2593 a_540271_687858.n103 vssa2 0.92fF $ **FLOATING
C2594 a_540271_687858.n104 vssa2 5.28fF $ **FLOATING
C2595 a_540271_687858.t48 vssa2 0.09fF
C2596 a_540271_687858.n105 vssa2 0.72fF $ **FLOATING
C2597 a_540271_687858.t3 vssa2 0.15fF
C2598 a_540271_687858.t30 vssa2 0.09fF
C2599 a_540271_687858.n106 vssa2 0.38fF $ **FLOATING
C2600 a_540271_687858.n107 vssa2 1.55fF $ **FLOATING
C2601 a_540271_687858.n108 vssa2 0.03fF $ **FLOATING
C2602 a_540271_687858.n109 vssa2 0.23fF $ **FLOATING
C2603 a_540271_687858.t37 vssa2 0.36fF
C2604 a_540271_687858.t38 vssa2 0.29fF
C2605 a_540271_687858.t29 vssa2 0.36fF
C2606 a_540271_687858.n110 vssa2 3.14fF $ **FLOATING
C2607 a_540271_687858.n111 vssa2 0.61fF $ **FLOATING
C2608 a_540271_687858.t36 vssa2 0.30fF
C2609 a_540271_687858.t35 vssa2 0.36fF
C2610 a_540271_687858.t27 vssa2 0.36fF
C2611 a_540271_687858.t28 vssa2 0.13fF
C2612 a_540271_687858.n112 vssa2 0.03fF $ **FLOATING
C2613 a_540271_687858.n113 vssa2 2.39fF $ **FLOATING
C2614 a_540271_687858.t41 vssa2 0.36fF
C2615 a_540271_687858.t12 vssa2 0.09fF
C2616 a_540271_687858.n114 vssa2 2.45fF $ **FLOATING
C2617 a_540271_687858.t11 vssa2 0.36fF
C2618 a_540271_687858.n115 vssa2 0.51fF $ **FLOATING
C2619 a_540271_687858.n116 vssa2 0.56fF $ **FLOATING
C2620 a_540271_687858.t63 vssa2 0.37fF
C2621 a_540271_687858.t57 vssa2 0.36fF
C2622 a_540271_687858.n117 vssa2 0.05fF $ **FLOATING
C2623 a_540271_687858.t68 vssa2 0.37fF
C2624 a_540271_687858.t60 vssa2 0.36fF
C2625 a_540271_687858.n118 vssa2 0.05fF $ **FLOATING
C2626 a_540271_687858.n119 vssa2 1.57fF $ **FLOATING
C2627 a_540271_687858.n120 vssa2 1.78fF $ **FLOATING
C2628 a_540271_687858.t53 vssa2 0.36fF
C2629 a_540271_687858.n121 vssa2 0.05fF $ **FLOATING
C2630 a_540271_687858.t59 vssa2 0.37fF
C2631 a_540271_687858.n122 vssa2 1.76fF $ **FLOATING
C2632 a_540271_687858.n123 vssa2 0.32fF $ **FLOATING
C2633 a_540271_687858.t42 vssa2 0.09fF
C2634 a_540271_687858.n124 vssa2 0.38fF $ **FLOATING
C2635 a_540271_687858.n125 vssa2 1.41fF $ **FLOATING
C2636 a_540271_687858.n126 vssa2 0.03fF $ **FLOATING
C2637 a_540271_687858.n127 vssa2 0.22fF $ **FLOATING
C2638 a_540271_687858.n128 vssa2 6.04fF $ **FLOATING
C2639 a_540271_687858.n129 vssa2 0.91fF $ **FLOATING
C2640 a_540271_687858.t0 vssa2 0.09fF
C2641 a_540271_687858.n130 vssa2 2.27fF $ **FLOATING
C2642 a_540271_687858.t22 vssa2 0.09fF
C2643 a_540271_687858.n131 vssa2 1.60fF $ **FLOATING
C2644 a_540271_687858.t21 vssa2 0.36fF
C2645 a_540271_687858.n132 vssa2 1.19fF $ **FLOATING
C2646 a_540271_687858.n133 vssa2 2.82fF $ **FLOATING
.ends

