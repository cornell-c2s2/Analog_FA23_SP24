magic
tech sky130A
magscale 1 2
timestamp 1713929811
<< pwell >>
rect -256 -10281 256 10281
<< nmoslvt >>
rect -60 9271 60 10071
rect -60 8253 60 9053
rect -60 7235 60 8035
rect -60 6217 60 7017
rect -60 5199 60 5999
rect -60 4181 60 4981
rect -60 3163 60 3963
rect -60 2145 60 2945
rect -60 1127 60 1927
rect -60 109 60 909
rect -60 -909 60 -109
rect -60 -1927 60 -1127
rect -60 -2945 60 -2145
rect -60 -3963 60 -3163
rect -60 -4981 60 -4181
rect -60 -5999 60 -5199
rect -60 -7017 60 -6217
rect -60 -8035 60 -7235
rect -60 -9053 60 -8253
rect -60 -10071 60 -9271
<< ndiff >>
rect -118 10059 -60 10071
rect -118 9283 -106 10059
rect -72 9283 -60 10059
rect -118 9271 -60 9283
rect 60 10059 118 10071
rect 60 9283 72 10059
rect 106 9283 118 10059
rect 60 9271 118 9283
rect -118 9041 -60 9053
rect -118 8265 -106 9041
rect -72 8265 -60 9041
rect -118 8253 -60 8265
rect 60 9041 118 9053
rect 60 8265 72 9041
rect 106 8265 118 9041
rect 60 8253 118 8265
rect -118 8023 -60 8035
rect -118 7247 -106 8023
rect -72 7247 -60 8023
rect -118 7235 -60 7247
rect 60 8023 118 8035
rect 60 7247 72 8023
rect 106 7247 118 8023
rect 60 7235 118 7247
rect -118 7005 -60 7017
rect -118 6229 -106 7005
rect -72 6229 -60 7005
rect -118 6217 -60 6229
rect 60 7005 118 7017
rect 60 6229 72 7005
rect 106 6229 118 7005
rect 60 6217 118 6229
rect -118 5987 -60 5999
rect -118 5211 -106 5987
rect -72 5211 -60 5987
rect -118 5199 -60 5211
rect 60 5987 118 5999
rect 60 5211 72 5987
rect 106 5211 118 5987
rect 60 5199 118 5211
rect -118 4969 -60 4981
rect -118 4193 -106 4969
rect -72 4193 -60 4969
rect -118 4181 -60 4193
rect 60 4969 118 4981
rect 60 4193 72 4969
rect 106 4193 118 4969
rect 60 4181 118 4193
rect -118 3951 -60 3963
rect -118 3175 -106 3951
rect -72 3175 -60 3951
rect -118 3163 -60 3175
rect 60 3951 118 3963
rect 60 3175 72 3951
rect 106 3175 118 3951
rect 60 3163 118 3175
rect -118 2933 -60 2945
rect -118 2157 -106 2933
rect -72 2157 -60 2933
rect -118 2145 -60 2157
rect 60 2933 118 2945
rect 60 2157 72 2933
rect 106 2157 118 2933
rect 60 2145 118 2157
rect -118 1915 -60 1927
rect -118 1139 -106 1915
rect -72 1139 -60 1915
rect -118 1127 -60 1139
rect 60 1915 118 1927
rect 60 1139 72 1915
rect 106 1139 118 1915
rect 60 1127 118 1139
rect -118 897 -60 909
rect -118 121 -106 897
rect -72 121 -60 897
rect -118 109 -60 121
rect 60 897 118 909
rect 60 121 72 897
rect 106 121 118 897
rect 60 109 118 121
rect -118 -121 -60 -109
rect -118 -897 -106 -121
rect -72 -897 -60 -121
rect -118 -909 -60 -897
rect 60 -121 118 -109
rect 60 -897 72 -121
rect 106 -897 118 -121
rect 60 -909 118 -897
rect -118 -1139 -60 -1127
rect -118 -1915 -106 -1139
rect -72 -1915 -60 -1139
rect -118 -1927 -60 -1915
rect 60 -1139 118 -1127
rect 60 -1915 72 -1139
rect 106 -1915 118 -1139
rect 60 -1927 118 -1915
rect -118 -2157 -60 -2145
rect -118 -2933 -106 -2157
rect -72 -2933 -60 -2157
rect -118 -2945 -60 -2933
rect 60 -2157 118 -2145
rect 60 -2933 72 -2157
rect 106 -2933 118 -2157
rect 60 -2945 118 -2933
rect -118 -3175 -60 -3163
rect -118 -3951 -106 -3175
rect -72 -3951 -60 -3175
rect -118 -3963 -60 -3951
rect 60 -3175 118 -3163
rect 60 -3951 72 -3175
rect 106 -3951 118 -3175
rect 60 -3963 118 -3951
rect -118 -4193 -60 -4181
rect -118 -4969 -106 -4193
rect -72 -4969 -60 -4193
rect -118 -4981 -60 -4969
rect 60 -4193 118 -4181
rect 60 -4969 72 -4193
rect 106 -4969 118 -4193
rect 60 -4981 118 -4969
rect -118 -5211 -60 -5199
rect -118 -5987 -106 -5211
rect -72 -5987 -60 -5211
rect -118 -5999 -60 -5987
rect 60 -5211 118 -5199
rect 60 -5987 72 -5211
rect 106 -5987 118 -5211
rect 60 -5999 118 -5987
rect -118 -6229 -60 -6217
rect -118 -7005 -106 -6229
rect -72 -7005 -60 -6229
rect -118 -7017 -60 -7005
rect 60 -6229 118 -6217
rect 60 -7005 72 -6229
rect 106 -7005 118 -6229
rect 60 -7017 118 -7005
rect -118 -7247 -60 -7235
rect -118 -8023 -106 -7247
rect -72 -8023 -60 -7247
rect -118 -8035 -60 -8023
rect 60 -7247 118 -7235
rect 60 -8023 72 -7247
rect 106 -8023 118 -7247
rect 60 -8035 118 -8023
rect -118 -8265 -60 -8253
rect -118 -9041 -106 -8265
rect -72 -9041 -60 -8265
rect -118 -9053 -60 -9041
rect 60 -8265 118 -8253
rect 60 -9041 72 -8265
rect 106 -9041 118 -8265
rect 60 -9053 118 -9041
rect -118 -9283 -60 -9271
rect -118 -10059 -106 -9283
rect -72 -10059 -60 -9283
rect -118 -10071 -60 -10059
rect 60 -9283 118 -9271
rect 60 -10059 72 -9283
rect 106 -10059 118 -9283
rect 60 -10071 118 -10059
<< ndiffc >>
rect -106 9283 -72 10059
rect 72 9283 106 10059
rect -106 8265 -72 9041
rect 72 8265 106 9041
rect -106 7247 -72 8023
rect 72 7247 106 8023
rect -106 6229 -72 7005
rect 72 6229 106 7005
rect -106 5211 -72 5987
rect 72 5211 106 5987
rect -106 4193 -72 4969
rect 72 4193 106 4969
rect -106 3175 -72 3951
rect 72 3175 106 3951
rect -106 2157 -72 2933
rect 72 2157 106 2933
rect -106 1139 -72 1915
rect 72 1139 106 1915
rect -106 121 -72 897
rect 72 121 106 897
rect -106 -897 -72 -121
rect 72 -897 106 -121
rect -106 -1915 -72 -1139
rect 72 -1915 106 -1139
rect -106 -2933 -72 -2157
rect 72 -2933 106 -2157
rect -106 -3951 -72 -3175
rect 72 -3951 106 -3175
rect -106 -4969 -72 -4193
rect 72 -4969 106 -4193
rect -106 -5987 -72 -5211
rect 72 -5987 106 -5211
rect -106 -7005 -72 -6229
rect 72 -7005 106 -6229
rect -106 -8023 -72 -7247
rect 72 -8023 106 -7247
rect -106 -9041 -72 -8265
rect 72 -9041 106 -8265
rect -106 -10059 -72 -9283
rect 72 -10059 106 -9283
<< psubdiff >>
rect -220 10211 -124 10245
rect 124 10211 220 10245
rect -220 10149 -186 10211
rect 186 10149 220 10211
rect -220 -10211 -186 -10149
rect 186 -10211 220 -10149
rect -220 -10245 -124 -10211
rect 124 -10245 220 -10211
<< psubdiffcont >>
rect -124 10211 124 10245
rect -220 -10149 -186 10149
rect 186 -10149 220 10149
rect -124 -10245 124 -10211
<< poly >>
rect -60 10143 60 10159
rect -60 10109 -44 10143
rect 44 10109 60 10143
rect -60 10071 60 10109
rect -60 9233 60 9271
rect -60 9199 -44 9233
rect 44 9199 60 9233
rect -60 9183 60 9199
rect -60 9125 60 9141
rect -60 9091 -44 9125
rect 44 9091 60 9125
rect -60 9053 60 9091
rect -60 8215 60 8253
rect -60 8181 -44 8215
rect 44 8181 60 8215
rect -60 8165 60 8181
rect -60 8107 60 8123
rect -60 8073 -44 8107
rect 44 8073 60 8107
rect -60 8035 60 8073
rect -60 7197 60 7235
rect -60 7163 -44 7197
rect 44 7163 60 7197
rect -60 7147 60 7163
rect -60 7089 60 7105
rect -60 7055 -44 7089
rect 44 7055 60 7089
rect -60 7017 60 7055
rect -60 6179 60 6217
rect -60 6145 -44 6179
rect 44 6145 60 6179
rect -60 6129 60 6145
rect -60 6071 60 6087
rect -60 6037 -44 6071
rect 44 6037 60 6071
rect -60 5999 60 6037
rect -60 5161 60 5199
rect -60 5127 -44 5161
rect 44 5127 60 5161
rect -60 5111 60 5127
rect -60 5053 60 5069
rect -60 5019 -44 5053
rect 44 5019 60 5053
rect -60 4981 60 5019
rect -60 4143 60 4181
rect -60 4109 -44 4143
rect 44 4109 60 4143
rect -60 4093 60 4109
rect -60 4035 60 4051
rect -60 4001 -44 4035
rect 44 4001 60 4035
rect -60 3963 60 4001
rect -60 3125 60 3163
rect -60 3091 -44 3125
rect 44 3091 60 3125
rect -60 3075 60 3091
rect -60 3017 60 3033
rect -60 2983 -44 3017
rect 44 2983 60 3017
rect -60 2945 60 2983
rect -60 2107 60 2145
rect -60 2073 -44 2107
rect 44 2073 60 2107
rect -60 2057 60 2073
rect -60 1999 60 2015
rect -60 1965 -44 1999
rect 44 1965 60 1999
rect -60 1927 60 1965
rect -60 1089 60 1127
rect -60 1055 -44 1089
rect 44 1055 60 1089
rect -60 1039 60 1055
rect -60 981 60 997
rect -60 947 -44 981
rect 44 947 60 981
rect -60 909 60 947
rect -60 71 60 109
rect -60 37 -44 71
rect 44 37 60 71
rect -60 21 60 37
rect -60 -37 60 -21
rect -60 -71 -44 -37
rect 44 -71 60 -37
rect -60 -109 60 -71
rect -60 -947 60 -909
rect -60 -981 -44 -947
rect 44 -981 60 -947
rect -60 -997 60 -981
rect -60 -1055 60 -1039
rect -60 -1089 -44 -1055
rect 44 -1089 60 -1055
rect -60 -1127 60 -1089
rect -60 -1965 60 -1927
rect -60 -1999 -44 -1965
rect 44 -1999 60 -1965
rect -60 -2015 60 -1999
rect -60 -2073 60 -2057
rect -60 -2107 -44 -2073
rect 44 -2107 60 -2073
rect -60 -2145 60 -2107
rect -60 -2983 60 -2945
rect -60 -3017 -44 -2983
rect 44 -3017 60 -2983
rect -60 -3033 60 -3017
rect -60 -3091 60 -3075
rect -60 -3125 -44 -3091
rect 44 -3125 60 -3091
rect -60 -3163 60 -3125
rect -60 -4001 60 -3963
rect -60 -4035 -44 -4001
rect 44 -4035 60 -4001
rect -60 -4051 60 -4035
rect -60 -4109 60 -4093
rect -60 -4143 -44 -4109
rect 44 -4143 60 -4109
rect -60 -4181 60 -4143
rect -60 -5019 60 -4981
rect -60 -5053 -44 -5019
rect 44 -5053 60 -5019
rect -60 -5069 60 -5053
rect -60 -5127 60 -5111
rect -60 -5161 -44 -5127
rect 44 -5161 60 -5127
rect -60 -5199 60 -5161
rect -60 -6037 60 -5999
rect -60 -6071 -44 -6037
rect 44 -6071 60 -6037
rect -60 -6087 60 -6071
rect -60 -6145 60 -6129
rect -60 -6179 -44 -6145
rect 44 -6179 60 -6145
rect -60 -6217 60 -6179
rect -60 -7055 60 -7017
rect -60 -7089 -44 -7055
rect 44 -7089 60 -7055
rect -60 -7105 60 -7089
rect -60 -7163 60 -7147
rect -60 -7197 -44 -7163
rect 44 -7197 60 -7163
rect -60 -7235 60 -7197
rect -60 -8073 60 -8035
rect -60 -8107 -44 -8073
rect 44 -8107 60 -8073
rect -60 -8123 60 -8107
rect -60 -8181 60 -8165
rect -60 -8215 -44 -8181
rect 44 -8215 60 -8181
rect -60 -8253 60 -8215
rect -60 -9091 60 -9053
rect -60 -9125 -44 -9091
rect 44 -9125 60 -9091
rect -60 -9141 60 -9125
rect -60 -9199 60 -9183
rect -60 -9233 -44 -9199
rect 44 -9233 60 -9199
rect -60 -9271 60 -9233
rect -60 -10109 60 -10071
rect -60 -10143 -44 -10109
rect 44 -10143 60 -10109
rect -60 -10159 60 -10143
<< polycont >>
rect -44 10109 44 10143
rect -44 9199 44 9233
rect -44 9091 44 9125
rect -44 8181 44 8215
rect -44 8073 44 8107
rect -44 7163 44 7197
rect -44 7055 44 7089
rect -44 6145 44 6179
rect -44 6037 44 6071
rect -44 5127 44 5161
rect -44 5019 44 5053
rect -44 4109 44 4143
rect -44 4001 44 4035
rect -44 3091 44 3125
rect -44 2983 44 3017
rect -44 2073 44 2107
rect -44 1965 44 1999
rect -44 1055 44 1089
rect -44 947 44 981
rect -44 37 44 71
rect -44 -71 44 -37
rect -44 -981 44 -947
rect -44 -1089 44 -1055
rect -44 -1999 44 -1965
rect -44 -2107 44 -2073
rect -44 -3017 44 -2983
rect -44 -3125 44 -3091
rect -44 -4035 44 -4001
rect -44 -4143 44 -4109
rect -44 -5053 44 -5019
rect -44 -5161 44 -5127
rect -44 -6071 44 -6037
rect -44 -6179 44 -6145
rect -44 -7089 44 -7055
rect -44 -7197 44 -7163
rect -44 -8107 44 -8073
rect -44 -8215 44 -8181
rect -44 -9125 44 -9091
rect -44 -9233 44 -9199
rect -44 -10143 44 -10109
<< locali >>
rect -220 10211 -124 10245
rect 124 10211 220 10245
rect -220 10149 -186 10211
rect 186 10149 220 10211
rect -60 10109 -44 10143
rect 44 10109 60 10143
rect -106 10059 -72 10075
rect -106 9267 -72 9283
rect 72 10059 106 10075
rect 72 9267 106 9283
rect -60 9199 -44 9233
rect 44 9199 60 9233
rect -60 9091 -44 9125
rect 44 9091 60 9125
rect -106 9041 -72 9057
rect -106 8249 -72 8265
rect 72 9041 106 9057
rect 72 8249 106 8265
rect -60 8181 -44 8215
rect 44 8181 60 8215
rect -60 8073 -44 8107
rect 44 8073 60 8107
rect -106 8023 -72 8039
rect -106 7231 -72 7247
rect 72 8023 106 8039
rect 72 7231 106 7247
rect -60 7163 -44 7197
rect 44 7163 60 7197
rect -60 7055 -44 7089
rect 44 7055 60 7089
rect -106 7005 -72 7021
rect -106 6213 -72 6229
rect 72 7005 106 7021
rect 72 6213 106 6229
rect -60 6145 -44 6179
rect 44 6145 60 6179
rect -60 6037 -44 6071
rect 44 6037 60 6071
rect -106 5987 -72 6003
rect -106 5195 -72 5211
rect 72 5987 106 6003
rect 72 5195 106 5211
rect -60 5127 -44 5161
rect 44 5127 60 5161
rect -60 5019 -44 5053
rect 44 5019 60 5053
rect -106 4969 -72 4985
rect -106 4177 -72 4193
rect 72 4969 106 4985
rect 72 4177 106 4193
rect -60 4109 -44 4143
rect 44 4109 60 4143
rect -60 4001 -44 4035
rect 44 4001 60 4035
rect -106 3951 -72 3967
rect -106 3159 -72 3175
rect 72 3951 106 3967
rect 72 3159 106 3175
rect -60 3091 -44 3125
rect 44 3091 60 3125
rect -60 2983 -44 3017
rect 44 2983 60 3017
rect -106 2933 -72 2949
rect -106 2141 -72 2157
rect 72 2933 106 2949
rect 72 2141 106 2157
rect -60 2073 -44 2107
rect 44 2073 60 2107
rect -60 1965 -44 1999
rect 44 1965 60 1999
rect -106 1915 -72 1931
rect -106 1123 -72 1139
rect 72 1915 106 1931
rect 72 1123 106 1139
rect -60 1055 -44 1089
rect 44 1055 60 1089
rect -60 947 -44 981
rect 44 947 60 981
rect -106 897 -72 913
rect -106 105 -72 121
rect 72 897 106 913
rect 72 105 106 121
rect -60 37 -44 71
rect 44 37 60 71
rect -60 -71 -44 -37
rect 44 -71 60 -37
rect -106 -121 -72 -105
rect -106 -913 -72 -897
rect 72 -121 106 -105
rect 72 -913 106 -897
rect -60 -981 -44 -947
rect 44 -981 60 -947
rect -60 -1089 -44 -1055
rect 44 -1089 60 -1055
rect -106 -1139 -72 -1123
rect -106 -1931 -72 -1915
rect 72 -1139 106 -1123
rect 72 -1931 106 -1915
rect -60 -1999 -44 -1965
rect 44 -1999 60 -1965
rect -60 -2107 -44 -2073
rect 44 -2107 60 -2073
rect -106 -2157 -72 -2141
rect -106 -2949 -72 -2933
rect 72 -2157 106 -2141
rect 72 -2949 106 -2933
rect -60 -3017 -44 -2983
rect 44 -3017 60 -2983
rect -60 -3125 -44 -3091
rect 44 -3125 60 -3091
rect -106 -3175 -72 -3159
rect -106 -3967 -72 -3951
rect 72 -3175 106 -3159
rect 72 -3967 106 -3951
rect -60 -4035 -44 -4001
rect 44 -4035 60 -4001
rect -60 -4143 -44 -4109
rect 44 -4143 60 -4109
rect -106 -4193 -72 -4177
rect -106 -4985 -72 -4969
rect 72 -4193 106 -4177
rect 72 -4985 106 -4969
rect -60 -5053 -44 -5019
rect 44 -5053 60 -5019
rect -60 -5161 -44 -5127
rect 44 -5161 60 -5127
rect -106 -5211 -72 -5195
rect -106 -6003 -72 -5987
rect 72 -5211 106 -5195
rect 72 -6003 106 -5987
rect -60 -6071 -44 -6037
rect 44 -6071 60 -6037
rect -60 -6179 -44 -6145
rect 44 -6179 60 -6145
rect -106 -6229 -72 -6213
rect -106 -7021 -72 -7005
rect 72 -6229 106 -6213
rect 72 -7021 106 -7005
rect -60 -7089 -44 -7055
rect 44 -7089 60 -7055
rect -60 -7197 -44 -7163
rect 44 -7197 60 -7163
rect -106 -7247 -72 -7231
rect -106 -8039 -72 -8023
rect 72 -7247 106 -7231
rect 72 -8039 106 -8023
rect -60 -8107 -44 -8073
rect 44 -8107 60 -8073
rect -60 -8215 -44 -8181
rect 44 -8215 60 -8181
rect -106 -8265 -72 -8249
rect -106 -9057 -72 -9041
rect 72 -8265 106 -8249
rect 72 -9057 106 -9041
rect -60 -9125 -44 -9091
rect 44 -9125 60 -9091
rect -60 -9233 -44 -9199
rect 44 -9233 60 -9199
rect -106 -9283 -72 -9267
rect -106 -10075 -72 -10059
rect 72 -9283 106 -9267
rect 72 -10075 106 -10059
rect -60 -10143 -44 -10109
rect 44 -10143 60 -10109
rect -220 -10211 -186 -10149
rect 186 -10211 220 -10149
rect -220 -10245 -124 -10211
rect 124 -10245 220 -10211
<< viali >>
rect -44 10109 44 10143
rect -106 9283 -72 10059
rect 72 9283 106 10059
rect -44 9199 44 9233
rect -44 9091 44 9125
rect -106 8265 -72 9041
rect 72 8265 106 9041
rect -44 8181 44 8215
rect -44 8073 44 8107
rect -106 7247 -72 8023
rect 72 7247 106 8023
rect -44 7163 44 7197
rect -44 7055 44 7089
rect -106 6229 -72 7005
rect 72 6229 106 7005
rect -44 6145 44 6179
rect -44 6037 44 6071
rect -106 5211 -72 5987
rect 72 5211 106 5987
rect -44 5127 44 5161
rect -44 5019 44 5053
rect -106 4193 -72 4969
rect 72 4193 106 4969
rect -44 4109 44 4143
rect -44 4001 44 4035
rect -106 3175 -72 3951
rect 72 3175 106 3951
rect -44 3091 44 3125
rect -44 2983 44 3017
rect -106 2157 -72 2933
rect 72 2157 106 2933
rect -44 2073 44 2107
rect -44 1965 44 1999
rect -106 1139 -72 1915
rect 72 1139 106 1915
rect -44 1055 44 1089
rect -44 947 44 981
rect -106 121 -72 897
rect 72 121 106 897
rect -44 37 44 71
rect -44 -71 44 -37
rect -106 -897 -72 -121
rect 72 -897 106 -121
rect -44 -981 44 -947
rect -44 -1089 44 -1055
rect -106 -1915 -72 -1139
rect 72 -1915 106 -1139
rect -44 -1999 44 -1965
rect -44 -2107 44 -2073
rect -106 -2933 -72 -2157
rect 72 -2933 106 -2157
rect -44 -3017 44 -2983
rect -44 -3125 44 -3091
rect -106 -3951 -72 -3175
rect 72 -3951 106 -3175
rect -44 -4035 44 -4001
rect -44 -4143 44 -4109
rect -106 -4969 -72 -4193
rect 72 -4969 106 -4193
rect -44 -5053 44 -5019
rect -44 -5161 44 -5127
rect -106 -5987 -72 -5211
rect 72 -5987 106 -5211
rect -44 -6071 44 -6037
rect -44 -6179 44 -6145
rect -106 -7005 -72 -6229
rect 72 -7005 106 -6229
rect -44 -7089 44 -7055
rect -44 -7197 44 -7163
rect -106 -8023 -72 -7247
rect 72 -8023 106 -7247
rect -44 -8107 44 -8073
rect -44 -8215 44 -8181
rect -106 -9041 -72 -8265
rect 72 -9041 106 -8265
rect -44 -9125 44 -9091
rect -44 -9233 44 -9199
rect -106 -10059 -72 -9283
rect 72 -10059 106 -9283
rect -44 -10143 44 -10109
<< metal1 >>
rect -56 10143 56 10149
rect -56 10109 -44 10143
rect 44 10109 56 10143
rect -56 10103 56 10109
rect -112 10059 -66 10071
rect -112 9283 -106 10059
rect -72 9283 -66 10059
rect -112 9271 -66 9283
rect 66 10059 112 10071
rect 66 9283 72 10059
rect 106 9283 112 10059
rect 66 9271 112 9283
rect -56 9233 56 9239
rect -56 9199 -44 9233
rect 44 9199 56 9233
rect -56 9193 56 9199
rect -56 9125 56 9131
rect -56 9091 -44 9125
rect 44 9091 56 9125
rect -56 9085 56 9091
rect -112 9041 -66 9053
rect -112 8265 -106 9041
rect -72 8265 -66 9041
rect -112 8253 -66 8265
rect 66 9041 112 9053
rect 66 8265 72 9041
rect 106 8265 112 9041
rect 66 8253 112 8265
rect -56 8215 56 8221
rect -56 8181 -44 8215
rect 44 8181 56 8215
rect -56 8175 56 8181
rect -56 8107 56 8113
rect -56 8073 -44 8107
rect 44 8073 56 8107
rect -56 8067 56 8073
rect -112 8023 -66 8035
rect -112 7247 -106 8023
rect -72 7247 -66 8023
rect -112 7235 -66 7247
rect 66 8023 112 8035
rect 66 7247 72 8023
rect 106 7247 112 8023
rect 66 7235 112 7247
rect -56 7197 56 7203
rect -56 7163 -44 7197
rect 44 7163 56 7197
rect -56 7157 56 7163
rect -56 7089 56 7095
rect -56 7055 -44 7089
rect 44 7055 56 7089
rect -56 7049 56 7055
rect -112 7005 -66 7017
rect -112 6229 -106 7005
rect -72 6229 -66 7005
rect -112 6217 -66 6229
rect 66 7005 112 7017
rect 66 6229 72 7005
rect 106 6229 112 7005
rect 66 6217 112 6229
rect -56 6179 56 6185
rect -56 6145 -44 6179
rect 44 6145 56 6179
rect -56 6139 56 6145
rect -56 6071 56 6077
rect -56 6037 -44 6071
rect 44 6037 56 6071
rect -56 6031 56 6037
rect -112 5987 -66 5999
rect -112 5211 -106 5987
rect -72 5211 -66 5987
rect -112 5199 -66 5211
rect 66 5987 112 5999
rect 66 5211 72 5987
rect 106 5211 112 5987
rect 66 5199 112 5211
rect -56 5161 56 5167
rect -56 5127 -44 5161
rect 44 5127 56 5161
rect -56 5121 56 5127
rect -56 5053 56 5059
rect -56 5019 -44 5053
rect 44 5019 56 5053
rect -56 5013 56 5019
rect -112 4969 -66 4981
rect -112 4193 -106 4969
rect -72 4193 -66 4969
rect -112 4181 -66 4193
rect 66 4969 112 4981
rect 66 4193 72 4969
rect 106 4193 112 4969
rect 66 4181 112 4193
rect -56 4143 56 4149
rect -56 4109 -44 4143
rect 44 4109 56 4143
rect -56 4103 56 4109
rect -56 4035 56 4041
rect -56 4001 -44 4035
rect 44 4001 56 4035
rect -56 3995 56 4001
rect -112 3951 -66 3963
rect -112 3175 -106 3951
rect -72 3175 -66 3951
rect -112 3163 -66 3175
rect 66 3951 112 3963
rect 66 3175 72 3951
rect 106 3175 112 3951
rect 66 3163 112 3175
rect -56 3125 56 3131
rect -56 3091 -44 3125
rect 44 3091 56 3125
rect -56 3085 56 3091
rect -56 3017 56 3023
rect -56 2983 -44 3017
rect 44 2983 56 3017
rect -56 2977 56 2983
rect -112 2933 -66 2945
rect -112 2157 -106 2933
rect -72 2157 -66 2933
rect -112 2145 -66 2157
rect 66 2933 112 2945
rect 66 2157 72 2933
rect 106 2157 112 2933
rect 66 2145 112 2157
rect -56 2107 56 2113
rect -56 2073 -44 2107
rect 44 2073 56 2107
rect -56 2067 56 2073
rect -56 1999 56 2005
rect -56 1965 -44 1999
rect 44 1965 56 1999
rect -56 1959 56 1965
rect -112 1915 -66 1927
rect -112 1139 -106 1915
rect -72 1139 -66 1915
rect -112 1127 -66 1139
rect 66 1915 112 1927
rect 66 1139 72 1915
rect 106 1139 112 1915
rect 66 1127 112 1139
rect -56 1089 56 1095
rect -56 1055 -44 1089
rect 44 1055 56 1089
rect -56 1049 56 1055
rect -56 981 56 987
rect -56 947 -44 981
rect 44 947 56 981
rect -56 941 56 947
rect -112 897 -66 909
rect -112 121 -106 897
rect -72 121 -66 897
rect -112 109 -66 121
rect 66 897 112 909
rect 66 121 72 897
rect 106 121 112 897
rect 66 109 112 121
rect -56 71 56 77
rect -56 37 -44 71
rect 44 37 56 71
rect -56 31 56 37
rect -56 -37 56 -31
rect -56 -71 -44 -37
rect 44 -71 56 -37
rect -56 -77 56 -71
rect -112 -121 -66 -109
rect -112 -897 -106 -121
rect -72 -897 -66 -121
rect -112 -909 -66 -897
rect 66 -121 112 -109
rect 66 -897 72 -121
rect 106 -897 112 -121
rect 66 -909 112 -897
rect -56 -947 56 -941
rect -56 -981 -44 -947
rect 44 -981 56 -947
rect -56 -987 56 -981
rect -56 -1055 56 -1049
rect -56 -1089 -44 -1055
rect 44 -1089 56 -1055
rect -56 -1095 56 -1089
rect -112 -1139 -66 -1127
rect -112 -1915 -106 -1139
rect -72 -1915 -66 -1139
rect -112 -1927 -66 -1915
rect 66 -1139 112 -1127
rect 66 -1915 72 -1139
rect 106 -1915 112 -1139
rect 66 -1927 112 -1915
rect -56 -1965 56 -1959
rect -56 -1999 -44 -1965
rect 44 -1999 56 -1965
rect -56 -2005 56 -1999
rect -56 -2073 56 -2067
rect -56 -2107 -44 -2073
rect 44 -2107 56 -2073
rect -56 -2113 56 -2107
rect -112 -2157 -66 -2145
rect -112 -2933 -106 -2157
rect -72 -2933 -66 -2157
rect -112 -2945 -66 -2933
rect 66 -2157 112 -2145
rect 66 -2933 72 -2157
rect 106 -2933 112 -2157
rect 66 -2945 112 -2933
rect -56 -2983 56 -2977
rect -56 -3017 -44 -2983
rect 44 -3017 56 -2983
rect -56 -3023 56 -3017
rect -56 -3091 56 -3085
rect -56 -3125 -44 -3091
rect 44 -3125 56 -3091
rect -56 -3131 56 -3125
rect -112 -3175 -66 -3163
rect -112 -3951 -106 -3175
rect -72 -3951 -66 -3175
rect -112 -3963 -66 -3951
rect 66 -3175 112 -3163
rect 66 -3951 72 -3175
rect 106 -3951 112 -3175
rect 66 -3963 112 -3951
rect -56 -4001 56 -3995
rect -56 -4035 -44 -4001
rect 44 -4035 56 -4001
rect -56 -4041 56 -4035
rect -56 -4109 56 -4103
rect -56 -4143 -44 -4109
rect 44 -4143 56 -4109
rect -56 -4149 56 -4143
rect -112 -4193 -66 -4181
rect -112 -4969 -106 -4193
rect -72 -4969 -66 -4193
rect -112 -4981 -66 -4969
rect 66 -4193 112 -4181
rect 66 -4969 72 -4193
rect 106 -4969 112 -4193
rect 66 -4981 112 -4969
rect -56 -5019 56 -5013
rect -56 -5053 -44 -5019
rect 44 -5053 56 -5019
rect -56 -5059 56 -5053
rect -56 -5127 56 -5121
rect -56 -5161 -44 -5127
rect 44 -5161 56 -5127
rect -56 -5167 56 -5161
rect -112 -5211 -66 -5199
rect -112 -5987 -106 -5211
rect -72 -5987 -66 -5211
rect -112 -5999 -66 -5987
rect 66 -5211 112 -5199
rect 66 -5987 72 -5211
rect 106 -5987 112 -5211
rect 66 -5999 112 -5987
rect -56 -6037 56 -6031
rect -56 -6071 -44 -6037
rect 44 -6071 56 -6037
rect -56 -6077 56 -6071
rect -56 -6145 56 -6139
rect -56 -6179 -44 -6145
rect 44 -6179 56 -6145
rect -56 -6185 56 -6179
rect -112 -6229 -66 -6217
rect -112 -7005 -106 -6229
rect -72 -7005 -66 -6229
rect -112 -7017 -66 -7005
rect 66 -6229 112 -6217
rect 66 -7005 72 -6229
rect 106 -7005 112 -6229
rect 66 -7017 112 -7005
rect -56 -7055 56 -7049
rect -56 -7089 -44 -7055
rect 44 -7089 56 -7055
rect -56 -7095 56 -7089
rect -56 -7163 56 -7157
rect -56 -7197 -44 -7163
rect 44 -7197 56 -7163
rect -56 -7203 56 -7197
rect -112 -7247 -66 -7235
rect -112 -8023 -106 -7247
rect -72 -8023 -66 -7247
rect -112 -8035 -66 -8023
rect 66 -7247 112 -7235
rect 66 -8023 72 -7247
rect 106 -8023 112 -7247
rect 66 -8035 112 -8023
rect -56 -8073 56 -8067
rect -56 -8107 -44 -8073
rect 44 -8107 56 -8073
rect -56 -8113 56 -8107
rect -56 -8181 56 -8175
rect -56 -8215 -44 -8181
rect 44 -8215 56 -8181
rect -56 -8221 56 -8215
rect -112 -8265 -66 -8253
rect -112 -9041 -106 -8265
rect -72 -9041 -66 -8265
rect -112 -9053 -66 -9041
rect 66 -8265 112 -8253
rect 66 -9041 72 -8265
rect 106 -9041 112 -8265
rect 66 -9053 112 -9041
rect -56 -9091 56 -9085
rect -56 -9125 -44 -9091
rect 44 -9125 56 -9091
rect -56 -9131 56 -9125
rect -56 -9199 56 -9193
rect -56 -9233 -44 -9199
rect 44 -9233 56 -9199
rect -56 -9239 56 -9233
rect -112 -9283 -66 -9271
rect -112 -10059 -106 -9283
rect -72 -10059 -66 -9283
rect -112 -10071 -66 -10059
rect 66 -9283 112 -9271
rect 66 -10059 72 -9283
rect 106 -10059 112 -9283
rect 66 -10071 112 -10059
rect -56 -10109 56 -10103
rect -56 -10143 -44 -10109
rect 44 -10143 56 -10109
rect -56 -10149 56 -10143
<< properties >>
string FIXED_BBOX -203 -10228 203 10228
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 4.0 l 0.6 m 20 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
