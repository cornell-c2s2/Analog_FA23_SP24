magic
tech sky130A
magscale 1 2
timestamp 1714790421
<< error_p >>
rect -4920 34 -3774 36
rect -3678 34 -2532 36
rect -2436 34 -1290 36
rect -1194 34 -48 36
rect 48 34 1194 36
rect 1290 34 2436 36
rect 2532 34 3678 36
rect 3774 34 4920 36
<< pwell >>
rect -5086 -632 5086 632
<< psubdiff >>
rect -5050 562 -4954 596
rect 4954 562 5050 596
rect -5050 500 -5016 562
rect 5016 500 5050 562
rect -5050 -562 -5016 -500
rect 5016 -562 5050 -500
rect -5050 -596 -4954 -562
rect 4954 -596 5050 -562
<< psubdiffcont >>
rect -4954 562 4954 596
rect -5050 -500 -5016 500
rect 5016 -500 5050 500
rect -4954 -596 4954 -562
<< xpolycontact >>
rect -4920 34 -3774 466
rect -4920 -466 -3774 -34
rect -3678 34 -2532 466
rect -3678 -466 -2532 -34
rect -2436 34 -1290 466
rect -2436 -466 -1290 -34
rect -1194 34 -48 466
rect -1194 -466 -48 -34
rect 48 34 1194 466
rect 48 -466 1194 -34
rect 1290 34 2436 466
rect 1290 -466 2436 -34
rect 2532 34 3678 466
rect 2532 -466 3678 -34
rect 3774 34 4920 466
rect 3774 -466 4920 -34
<< xpolyres >>
rect -4920 -34 -3774 34
rect -3678 -34 -2532 34
rect -2436 -34 -1290 34
rect -1194 -34 -48 34
rect 48 -34 1194 34
rect 1290 -34 2436 34
rect 2532 -34 3678 34
rect 3774 -34 4920 34
<< locali >>
rect -5050 562 -4954 596
rect 4954 562 5050 596
rect -5050 500 -5016 562
rect 5016 500 5050 562
rect -5050 -562 -5016 -500
rect 5016 -562 5050 -500
rect -5050 -596 -4954 -562
rect 4954 -596 5050 -562
<< viali >>
rect -4904 51 -3790 448
rect -3662 51 -2548 448
rect -2420 51 -1306 448
rect -1178 51 -64 448
rect 64 51 1178 448
rect 1306 51 2420 448
rect 2548 51 3662 448
rect 3790 51 4904 448
rect -4904 -448 -3790 -51
rect -3662 -448 -2548 -51
rect -2420 -448 -1306 -51
rect -1178 -448 -64 -51
rect 64 -448 1178 -51
rect 1306 -448 2420 -51
rect 2548 -448 3662 -51
rect 3790 -448 4904 -51
<< metal1 >>
rect -4916 448 -3778 454
rect -4916 51 -4904 448
rect -3790 51 -3778 448
rect -4916 45 -3778 51
rect -3674 448 -2536 454
rect -3674 51 -3662 448
rect -2548 51 -2536 448
rect -3674 45 -2536 51
rect -2432 448 -1294 454
rect -2432 51 -2420 448
rect -1306 51 -1294 448
rect -2432 45 -1294 51
rect -1190 448 -52 454
rect -1190 51 -1178 448
rect -64 51 -52 448
rect -1190 45 -52 51
rect 52 448 1190 454
rect 52 51 64 448
rect 1178 51 1190 448
rect 52 45 1190 51
rect 1294 448 2432 454
rect 1294 51 1306 448
rect 2420 51 2432 448
rect 1294 45 2432 51
rect 2536 448 3674 454
rect 2536 51 2548 448
rect 3662 51 3674 448
rect 2536 45 3674 51
rect 3778 448 4916 454
rect 3778 51 3790 448
rect 4904 51 4916 448
rect 3778 45 4916 51
rect -4916 -51 -3778 -45
rect -4916 -448 -4904 -51
rect -3790 -448 -3778 -51
rect -4916 -454 -3778 -448
rect -3674 -51 -2536 -45
rect -3674 -448 -3662 -51
rect -2548 -448 -2536 -51
rect -3674 -454 -2536 -448
rect -2432 -51 -1294 -45
rect -2432 -448 -2420 -51
rect -1306 -448 -1294 -51
rect -2432 -454 -1294 -448
rect -1190 -51 -52 -45
rect -1190 -448 -1178 -51
rect -64 -448 -52 -51
rect -1190 -454 -52 -448
rect 52 -51 1190 -45
rect 52 -448 64 -51
rect 1178 -448 1190 -51
rect 52 -454 1190 -448
rect 1294 -51 2432 -45
rect 1294 -448 1306 -51
rect 2420 -448 2432 -51
rect 1294 -454 2432 -448
rect 2536 -51 3674 -45
rect 2536 -448 2548 -51
rect 3662 -448 3674 -51
rect 2536 -454 3674 -448
rect 3778 -51 4916 -45
rect 3778 -448 3790 -51
rect 4904 -448 4916 -51
rect 3778 -454 4916 -448
<< properties >>
string FIXED_BBOX -5033 -579 5033 579
string gencell sky130_fd_pr__res_xhigh_po_5p73
string library sky130
string parameters w 5.73 l 0.50 m 1 nx 8 wmin 5.730 lmin 0.50 rho 2000 val 240.209 dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 5.730 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
