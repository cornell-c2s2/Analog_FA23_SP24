* NGSPICE file created from RSfetsym-ext_flat.ext - technology: sky130A

.subckt RSfetsym-ext_flat VDD S R QN Q GND
X0 VDD.t23 S.t0 Q.t3 VDD.t22 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.25
X1 VDD.t3 Q.t5 QN.t1 VDD.t2 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.3
X2 x1.Y R.t0 GND.t9 GND.t8 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X3 x2.Y S.t1 GND.t19 GND.t18 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 x2.Y S.t2 VDD.t21 VDD.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 QN.t0 R.t1 VDD.t1 VDD.t0 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.25
X6 GND.t7 R.t2 x1.Y GND.t6 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X7 GND.t23 x2.Y QN.t4 GND.t22 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.25
X8 Q.t1 S.t3 VDD.t19 VDD.t18 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.25
X9 Q.t2 S.t4 a_1070_n1178# GND.t10 sky130_fd_pr__nfet_01v8 ad=0.315 pd=2.72 as=0.29 ps=2.58 w=1 l=0.15
X10 x1.Y R.t3 GND.t5 GND.t4 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11 GND.t3 R.t4 x1.Y GND.t2 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X12 VDD.t20 S.t5 x2.Y VDD.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13 GND.t17 S.t6 x2.Y GND.t16 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X14 x2.Y S.t7 GND.t15 GND.t14 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X15 GND.t13 S.t8 x2.Y GND.t12 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X16 x2.Y S.t9 VDD.t17 VDD.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X17 VDD.t16 S.t10 x2.Y VDD.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X18 a_1070_n1178# QN.t5 GND.t11 GND.t10 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X19 x1.Y R.t5 VDD.t7 VDD.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X20 a_1583_n1177# Q.t6 GND.t1 GND.t0 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X21 VDD.t5 R.t6 x1.Y VDD.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X22 x1.Y R.t7 VDD.t13 VDD.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X23 VDD.t11 R.t8 x1.Y VDD.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X24 QN.t2 R.t9 a_1583_n1177# GND.t0 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X25 VDD.t15 QN.t6 Q.t0 VDD.t14 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.3
X26 VDD.t9 R.t10 QN.t3 VDD.t8 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.25
X27 GND.t21 x1.Y Q.t4 GND.t20 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.25
R0 S.n19 S.t3 258.589
R1 S.n15 S.t0 258.58
R2 S.n40 S.t10 212.081
R3 S.n41 S.t2 212.081
R4 S.n33 S.t5 212.081
R5 S.n7 S.t9 212.081
R6 S.n40 S.t8 139.78
R7 S.n41 S.t1 139.78
R8 S.n33 S.t6 139.78
R9 S.n7 S.t7 139.78
R10 S.n20 S.t4 117.227
R11 S.n42 S.n40 30.6732
R12 S.n42 S.n41 30.6732
R13 S.n34 S.n33 30.6732
R14 S.n8 S.n7 29.9429
R15 S S.n26 12.8005
R16 S.n6 S.n5 11.6853
R17 S.n9 S.n8 9.3005
R18 S.n32 S.n31 9.3005
R19 S.n43 S.n42 8.75567
R20 S.n35 S.n34 8.28655
R21 S.n24 S.n10 4.6085
R22 S.n36 S.n1 4.3525
R23 S.n35 S 4.3525
R24 S.n28 S.n27 4.3525
R25 S.n26 S.n25 4.3525
R26 S.n4 S.n3 4.0965
R27 S S.n44 2.8165
R28 S.n22 S.n21 1.83593
R29 S S.n43 1.79306
R30 S.n17 S.n16 1.35797
R31 S.n10 S 1.2805
R32 S.n27 S 1.0245
R33 S.n28 S.n9 0.7685
R34 S.n8 S.n6 0.730803
R35 S.n36 S.n35 0.5125
R36 S.n25 S.n24 0.5125
R37 S.n21 S.n18 0.429669
R38 S S.n32 0.2565
R39 S.n9 S.n4 0.2565
R40 S.n18 S.n17 0.215426
R41 S.n20 S.n19 0.12975
R42 S.n18 S 0.0828355
R43 S.n31 S.n30 0.0766364
R44 S.n11 S.n2 0.0618636
R45 S.n39 S.n38 0.0516364
R46 S.n14 S.n13 0.034875
R47 S.n43 S.n39 0.0220871
R48 S.n31 S.n0 0.0209545
R49 S.n23 S.n22 0.0209545
R50 S.n38 S.n37 0.0198182
R51 S.n29 S.n2 0.0198182
R52 S.n12 S.n11 0.0198182
R53 S.n17 S.n14 0.0130265
R54 S.n16 S.n15 0.00883333
R55 S.n30 S.n29 0.00390909
R56 S.n21 S.n20 0.0028536
R57 S.n37 S.n0 0.00277273
R58 S.n23 S.n12 0.00277273
R59 S.n29 S.n28 0.00119109
R60 S.n37 S.n36 0.00119109
R61 S.n24 S.n23 0.00119109
R62 Q.n0 Q.t6 117.522
R63 Q.n0 Q.t5 110.698
R64 Q.n3 Q.t2 19.1973
R65 Q.n5 Q.t0 14.2842
R66 Q.n9 Q.t3 14.283
R67 Q.n9 Q.t1 14.283
R68 Q.n11 Q.t4 9.14126
R69 Q.n5 Q.n4 7.90638
R70 Q.n11 Q.n10 0.746571
R71 Q.n1 Q.n0 0.685831
R72 Q.n10 Q.n8 0.2402
R73 Q.n8 Q.n7 0.237833
R74 Q Q.n11 0.132261
R75 Q.n3 Q.n2 0.132187
R76 Q.n8 Q.n3 0.0968646
R77 Q.n7 Q.n6 0.0272537
R78 Q.n10 Q.n9 0.0107755
R79 Q.n2 Q.n1 0.00981526
R80 Q.n7 Q.n5 0.00225338
R81 VDD.n89 VDD.n86 1224.71
R82 VDD.n94 VDD.n92 1069.41
R83 VDD.n104 VDD.n102 593.144
R84 VDD.n5 VDD.t16 584.644
R85 VDD.n6 VDD.t11 584.644
R86 VDD.n54 VDD.n52 576.668
R87 VDD.n100 VDD.n98 370.589
R88 VDD.n49 VDD.n47 370.589
R89 VDD.t10 VDD.n147 286.462
R90 VDD.n118 VDD.n117 185
R91 VDD.n16 VDD.n15 174.595
R92 VDD.n14 VDD.n13 174.595
R93 VDD.n135 VDD.n134 158.457
R94 VDD.n7 VDD.t17 151.123
R95 VDD.n8 VDD.t13 151.123
R96 VDD.n63 VDD.n62 143.435
R97 VDD.n88 VDD.n87 131.012
R98 VDD.t6 VDD.t10 122.769
R99 VDD.t4 VDD.t6 122.769
R100 VDD.t12 VDD.t4 122.769
R101 VDD.n84 VDD.n83 116.267
R102 VDD.t18 VDD.n116 110.177
R103 VDD VDD.t12 109.615
R104 VDD.n106 VDD.n105 63.2691
R105 VDD.n56 VDD.n55 61.5116
R106 VDD.n55 VDD.n51 61.5116
R107 VDD.n128 VDD.t22 61.2177
R108 VDD.n128 VDD.t18 61.2177
R109 VDD.n41 VDD.t8 61.2177
R110 VDD.n41 VDD.t0 61.2177
R111 VDD.n126 VDD.n118 45.817
R112 VDD.n106 VDD.n101 39.5299
R113 VDD.n56 VDD.n50 39.5299
R114 VDD.n15 VDD.t21 26.5955
R115 VDD.n15 VDD.t20 26.5955
R116 VDD.n13 VDD.t7 26.5955
R117 VDD.n13 VDD.t5 26.5955
R118 VDD.n107 VDD.n106 20.9134
R119 VDD.n57 VDD.n56 17.109
R120 VDD.n111 VDD.t19 14.2962
R121 VDD.n25 VDD.t23 14.2955
R122 VDD.n59 VDD.t1 14.2865
R123 VDD.n60 VDD.t9 14.2864
R124 VDD.n97 VDD.t15 14.2849
R125 VDD.n72 VDD.t3 14.2849
R126 VDD.n95 VDD.n91 14.0805
R127 VDD.n79 VDD.n76 13.7605
R128 VDD.n121 VDD.n120 9.3005
R129 VDD.n37 VDD.n36 9.3005
R130 VDD.n32 VDD.n31 9.3005
R131 VDD.n108 VDD.n107 9.3005
R132 VDD.n27 VDD.n26 4.66685
R133 VDD.n9 VDD.n8 4.6505
R134 VDD.n12 VDD.n10 4.6505
R135 VDD.n17 VDD.n14 4.6505
R136 VDD.n20 VDD.n18 4.6505
R137 VDD.n21 VDD.n6 4.6505
R138 VDD.n9 VDD.n7 4.6505
R139 VDD.n12 VDD.n11 4.6505
R140 VDD.n17 VDD.n16 4.6505
R141 VDD.n20 VDD.n19 4.6505
R142 VDD.n21 VDD.n5 4.6505
R143 VDD.n58 VDD.n57 4.5005
R144 VDD.n137 VDD.n136 4.5005
R145 VDD.n109 VDD.n97 1.51475
R146 VDD.n57 VDD.n46 1.06717
R147 VDD.n130 VDD.n115 0.6405
R148 VDD.n146 VDD.n145 0.599115
R149 VDD.n110 VDD.n25 0.467504
R150 VDD.n112 VDD.n111 0.456265
R151 VDD.n67 VDD.n60 0.399688
R152 VDD.n72 VDD.n71 0.39626
R153 VDD.n69 VDD.n59 0.38579
R154 VDD.n125 VDD.n124 0.338059
R155 VDD.n136 VDD.n135 0.3205
R156 VDD.n123 VDD.n121 0.29425
R157 VDD.n34 VDD.n32 0.261214
R158 VDD.n38 VDD.n37 0.261214
R159 VDD.n82 VDD.n80 0.248103
R160 VDD.n96 VDD.n85 0.247868
R161 VDD.n68 VDD.n67 0.232774
R162 VDD.n45 VDD.n44 0.217167
R163 VDD.n137 VDD.n132 0.201889
R164 VDD.n50 VDD.n49 0.164944
R165 VDD.n49 VDD.n48 0.164944
R166 VDD.n101 VDD.n100 0.15889
R167 VDD.n100 VDD.n99 0.15889
R168 VDD.n140 VDD.n110 0.117306
R169 VDD.n140 VDD.n139 0.0856364
R170 VDD.n32 VDD.n30 0.07913
R171 VDD.n22 VDD.n21 0.0789722
R172 VDD.n121 VDD.n119 0.0773443
R173 VDD.n37 VDD.n35 0.0773443
R174 VDD.n21 VDD.n20 0.0643889
R175 VDD.n20 VDD.n17 0.0643889
R176 VDD.n17 VDD.n12 0.0643889
R177 VDD.n12 VDD.n9 0.0643889
R178 VDD.n142 VDD 0.0630006
R179 VDD.n109 VDD.n108 0.0602222
R180 VDD.n141 VDD.n140 0.0464453
R181 VDD.n29 VDD.n27 0.0352222
R182 VDD.n70 VDD.n58 0.0352222
R183 VDD.n139 VDD.n138 0.0349477
R184 VDD.n97 VDD.n96 0.0294474
R185 VDD.n80 VDD.n72 0.0287895
R186 VDD.n105 VDD.n104 0.0282694
R187 VDD.n104 VDD.n103 0.0282694
R188 VDD.n55 VDD.n54 0.0282694
R189 VDD.n54 VDD.n53 0.0282694
R190 VDD.n23 VDD.n22 0.0178611
R191 VDD.n76 VDD.n75 0.0163404
R192 VDD.n75 VDD.t2 0.0163404
R193 VDD.n91 VDD.n90 0.0163404
R194 VDD.n90 VDD.t14 0.0163404
R195 VDD.n139 VDD.n112 0.0153419
R196 VDD.n69 VDD.n68 0.0148892
R197 VDD.n71 VDD.n70 0.0143889
R198 VDD.n9 VDD 0.0123056
R199 VDD.n65 VDD.n64 0.0114541
R200 VDD.n134 VDD.n133 0.0084202
R201 VDD.n89 VDD.n88 0.0084202
R202 VDD.t14 VDD.n89 0.0084202
R203 VDD.n74 VDD.n73 0.0084202
R204 VDD.t2 VDD.n74 0.0084202
R205 VDD.n62 VDD.n61 0.0084202
R206 VDD.n125 VDD.n123 0.00675
R207 VDD.n66 VDD.n65 0.00605556
R208 VDD.n58 VDD.n45 0.00466667
R209 VDD.n131 VDD.n114 0.00466667
R210 VDD.n85 VDD.n84 0.00445072
R211 VDD.n132 VDD.n131 0.00327778
R212 VDD.n147 VDD.n146 0.00281774
R213 VDD.n38 VDD.n34 0.00228571
R214 VDD.n126 VDD.n125 0.00221302
R215 VDD.n39 VDD.n38 0.00220642
R216 VDD.n44 VDD.n43 0.00220642
R217 VDD.n131 VDD.n130 0.00220642
R218 VDD.n127 VDD.n126 0.00213073
R219 VDD.n128 VDD.n127 0.00213073
R220 VDD.n130 VDD.n129 0.00212475
R221 VDD.n40 VDD.n39 0.00212475
R222 VDD.n41 VDD.n40 0.00212475
R223 VDD.n43 VDD.n42 0.00212475
R224 VDD.n42 VDD.n41 0.00212475
R225 VDD.n129 VDD.n128 0.00212475
R226 VDD.n44 VDD.n29 0.00188889
R227 VDD.n138 VDD.n137 0.00188889
R228 VDD.n24 VDD.n23 0.00160338
R229 VDD.n23 VDD.n4 0.0014897
R230 VDD.n96 VDD.n95 0.00145131
R231 VDD.n95 VDD.n94 0.00145131
R232 VDD.n94 VDD.n93 0.00145131
R233 VDD.n80 VDD.n79 0.00144714
R234 VDD.n79 VDD.n78 0.00144714
R235 VDD.n78 VDD.n77 0.00144714
R236 VDD.n85 VDD.n82 0.00139286
R237 VDD.n1 VDD.n0 0.00133311
R238 VDD.n143 VDD.n141 0.00121484
R239 VDD.n67 VDD.n66 0.00113805
R240 VDD.n23 VDD.n3 0.001086
R241 VDD.n145 VDD.n144 0.00107785
R242 VDD.n70 VDD.n69 0.00105186
R243 VDD.n147 VDD.n24 0.0010245
R244 VDD.n23 VDD.n1 0.00100128
R245 VDD.n145 VDD.n143 0.00100103
R246 VDD.n3 VDD.n2 0.00100075
R247 VDD.n110 VDD.n109 0.000558569
R248 VDD.n66 VDD.n63 0.000555817
R249 VDD.n114 VDD.n113 0.000516232
R250 VDD.n123 VDD.n122 0.000516232
R251 VDD.n29 VDD.n28 0.000515622
R252 VDD.n34 VDD.n33 0.000505865
R253 VDD.n82 VDD.n81 0.000503792
R254 VDD.n143 VDD.n142 0.000500084
R255 QN.n2 QN.t5 117.314
R256 QN.n2 QN.t6 110.852
R257 QN.n1 QN.t2 17.6182
R258 QN.n4 QN.t1 14.2865
R259 QN.n0 QN.t3 14.283
R260 QN.n0 QN.t0 14.283
R261 QN.n7 QN.t4 8.77813
R262 QN.n7 QN.n6 1.20426
R263 QN QN.n7 0.364385
R264 QN.n5 QN.n4 0.299268
R265 QN.n3 QN.n2 0.159555
R266 QN.n6 QN.n0 0.107614
R267 QN.n5 QN.n3 0.0796167
R268 QN.n6 QN.n5 0.0480595
R269 QN.n3 QN.n1 0.000504658
R270 R.n13 R.t10 258.584
R271 R.n23 R.t1 258.58
R272 R.n46 R.t8 212.081
R273 R.n47 R.t5 212.081
R274 R.n39 R.t6 212.081
R275 R.n7 R.t7 212.081
R276 R.n46 R.t4 139.78
R277 R.n47 R.t0 139.78
R278 R.n39 R.t2 139.78
R279 R.n7 R.t3 139.78
R280 R.n19 R.t9 110.734
R281 R.n48 R.n46 30.6732
R282 R.n48 R.n47 30.6732
R283 R.n40 R.n39 30.6732
R284 R.n8 R.n7 29.9429
R285 R R.n32 12.8005
R286 R.n6 R.n5 11.6853
R287 R.n9 R.n8 9.3005
R288 R.n38 R.n37 9.3005
R289 R.n49 R.n48 8.75567
R290 R.n41 R.n40 8.28655
R291 R.n30 R.n10 4.6085
R292 R.n42 R.n1 4.3525
R293 R.n41 R 4.3525
R294 R.n34 R.n33 4.3525
R295 R.n32 R.n31 4.3525
R296 R.n4 R.n3 4.0965
R297 R R.n50 2.8165
R298 R R.n49 1.79306
R299 R.n28 R.n27 1.54944
R300 R.n10 R 1.2805
R301 R.n33 R 1.0245
R302 R.n34 R.n9 0.7685
R303 R.n8 R.n6 0.730803
R304 R.n42 R.n41 0.5125
R305 R.n31 R.n30 0.5125
R306 R.n27 R.n18 0.44229
R307 R R.n38 0.2565
R308 R.n9 R.n4 0.2565
R309 R.n18 R.n17 0.178789
R310 R.n27 R.n26 0.14376
R311 R.n37 R.n36 0.105187
R312 R.n18 R 0.0926682
R313 R.n11 R.n2 0.0844489
R314 R.n45 R.n44 0.0708125
R315 R.n26 R.n25 0.0475
R316 R.n49 R.n45 0.0297575
R317 R.n37 R.n0 0.028625
R318 R.n44 R.n43 0.0270625
R319 R.n35 R.n2 0.0270625
R320 R.n16 R.n15 0.0255
R321 R.n29 R.n28 0.0209545
R322 R.n12 R.n11 0.0198182
R323 R.n21 R.n20 0.0172791
R324 R.n22 R.n19 0.0133182
R325 R.n24 R.n23 0.00951733
R326 R.n14 R.n13 0.00583593
R327 R.n36 R.n35 0.0051875
R328 R.n17 R.n16 0.00390909
R329 R.n43 R.n0 0.003625
R330 R.n29 R.n12 0.00277273
R331 R.n25 R.n22 0.00263636
R332 R.n43 R.n42 0.00119109
R333 R.n35 R.n34 0.00119109
R334 R.n30 R.n29 0.00119109
R335 R.n22 R.n21 0.000747155
R336 R.n25 R.n24 0.000588765
R337 R.n17 R.n14 0.000588763
R338 GND.n25 GND.t12 1878.21
R339 GND.n1 GND.n0 1773
R340 GND.n49 GND.n48 1773
R341 GND.n52 GND.n49 1384.79
R342 GND.n2 GND.n1 1384.79
R343 GND.n27 GND.n23 841.244
R344 GND.n82 GND.n79 816.971
R345 GND.n37 GND.n35 816.971
R346 GND.t12 GND.t18 551.643
R347 GND.t18 GND.t16 551.643
R348 GND.t16 GND.t14 551.643
R349 GND.t14 GND 492.538
R350 GND.n27 GND.n22 473.865
R351 GND.n147 GND 440
R352 GND.n82 GND.n78 422.971
R353 GND.t0 GND.t2 411.332
R354 GND.t6 GND.t8 349.01
R355 GND.t4 GND.t6 349.01
R356 GND GND.t4 311.615
R357 GND GND.n147 278.377
R358 GND.n78 GND.n77 197
R359 GND.n114 GND.t3 196.756
R360 GND.n3 GND.t13 196.633
R361 GND.n115 GND.t5 193.933
R362 GND.n140 GND.t15 193.933
R363 GND.n26 GND.n25 154.464
R364 GND.n81 GND.n80 121.365
R365 GND.n58 GND.n57 115.201
R366 GND.n125 GND.n124 114.713
R367 GND.n6 GND.n5 114.713
R368 GND.n26 GND.n24 103.712
R369 GND.n145 GND.n144 96.7534
R370 GND.n51 GND.n50 90.3534
R371 GND.n145 GND.n143 90.3427
R372 GND.t10 GND.n142 55.4632
R373 GND.n29 GND.n28 30.7897
R374 GND.n85 GND.n84 28.4429
R375 GND.n84 GND.n83 27.4829
R376 GND.n147 GND.t10 25.5893
R377 GND.n124 GND.t9 24.9236
R378 GND.n124 GND.t7 24.9236
R379 GND.n5 GND.t19 24.9236
R380 GND.n5 GND.t17 24.9236
R381 GND.n30 GND.n29 22.9087
R382 GND.n33 GND.n32 22.0993
R383 GND.n59 GND.n58 22.0886
R384 GND.n75 GND.n74 20.3111
R385 GND.n113 GND.t11 17.474
R386 GND.n113 GND.t1 17.4535
R387 GND.n118 GND.n117 9.3005
R388 GND.n120 GND.n119 9.3005
R389 GND.n139 GND.n138 9.3005
R390 GND.n93 GND.n92 9.3005
R391 GND.n86 GND.n85 9.3005
R392 GND.n68 GND.n67 9.3005
R393 GND.n76 GND.n75 9.3005
R394 GND.n66 GND.n65 9.3005
R395 GND.n62 GND.n61 9.3005
R396 GND.n45 GND.n44 9.3005
R397 GND.n60 GND.n59 9.3005
R398 GND.n43 GND.n42 9.3005
R399 GND.n34 GND.n33 9.3005
R400 GND.n31 GND.n30 9.3005
R401 GND.n107 GND.n106 9.3005
R402 GND.n110 GND.n109 9.3005
R403 GND.n13 GND.n12 9.3005
R404 GND.n95 GND.n94 9.3005
R405 GND.n142 GND 9.21319
R406 GND.n14 GND.t21 8.70904
R407 GND.n105 GND.t23 8.70236
R408 GND.n116 GND.n115 4.6505
R409 GND.n141 GND.n140 4.6505
R410 GND.n122 GND.n121 4.5005
R411 GND.n126 GND.n125 3.03311
R412 GND.n137 GND.n136 3.03311
R413 GND.n7 GND.n6 3.03311
R414 GND.n111 GND.n110 0.533636
R415 GND.n14 GND.n13 0.425574
R416 GND.n34 GND.n31 0.378476
R417 GND.n60 GND.n55 0.377583
R418 GND.n47 GND.n45 0.3755
R419 GND.n64 GND.n62 0.373417
R420 GND.n66 GND.n64 0.373417
R421 GND.n57 GND.n56 0.366214
R422 GND.n100 GND.n99 0.345738
R423 GND.n62 GND.n60 0.31925
R424 GND.n86 GND.n76 0.313
R425 GND.n127 GND.n114 0.301442
R426 GND.n107 GND.n105 0.290381
R427 GND.n4 GND.n3 0.284578
R428 GND.n45 GND.n43 0.248417
R429 GND.n68 GND.n66 0.238893
R430 GND.n130 GND.n129 0.224247
R431 GND.n112 GND.n101 0.219655
R432 GND.n95 GND.n93 0.200996
R433 GND.n111 GND.n108 0.181736
R434 GND.n112 GND.n111 0.17675
R435 GND.n39 GND.n34 0.171333
R436 GND.n43 GND.n41 0.16925
R437 GND.n91 GND.n86 0.164786
R438 GND.n93 GND.n91 0.164786
R439 GND.n31 GND.n21 0.159429
R440 GND.n71 GND.n68 0.148714
R441 GND.n76 GND.n73 0.148714
R442 GND.n130 GND 0.142351
R443 GND.n101 GND.n100 0.135635
R444 GND.n83 GND.n82 0.10956
R445 GND.n82 GND.n81 0.10956
R446 GND.n28 GND.n27 0.10956
R447 GND.n27 GND.n26 0.10956
R448 GND.t22 GND.n16 0.0944005
R449 GND.n16 GND.n15 0.0944005
R450 GND.t20 GND.n88 0.0944005
R451 GND.n88 GND.n87 0.0944005
R452 GND.n118 GND.n116 0.09425
R453 GND.n141 GND.n139 0.0857273
R454 GND.n101 GND.n14 0.0788333
R455 GND.n7 GND.n4 0.0768735
R456 GND.n11 GND.n10 0.058
R457 GND.n133 GND.n11 0.05425
R458 GND.n137 GND.n135 0.0527727
R459 GND.n113 GND.n112 0.0494583
R460 GND.n135 GND.n134 0.0493636
R461 GND.n126 GND.n123 0.0432584
R462 GND.t0 GND.n52 0.0425017
R463 GND.n52 GND.n51 0.0425017
R464 GND.t10 GND.n146 0.0425017
R465 GND.n146 GND.n145 0.0425017
R466 GND.n123 GND.n122 0.0392297
R467 GND.n100 GND.n95 0.0345278
R468 GND.n129 GND.n113 0.0337917
R469 GND.n139 GND.n137 0.0198182
R470 GND GND.n141 0.0198182
R471 GND.n116 GND 0.0182083
R472 GND.n122 GND.n120 0.016125
R473 GND.n108 GND.n107 0.0112143
R474 GND.n73 GND.n71 0.00585714
R475 GND.n55 GND.n47 0.00466667
R476 GND.n133 GND.n9 0.00425
R477 GND.n71 GND.n70 0.00396627
R478 GND.n39 GND.n38 0.00396498
R479 GND.n131 GND.n130 0.00395031
R480 GND.n70 GND.n69 0.0039133
R481 GND.n38 GND.n37 0.0039133
R482 GND.n37 GND.n36 0.0039133
R483 GND.n134 GND.n7 0.00390909
R484 GND.n19 GND.n18 0.00348555
R485 GND.n90 GND.n89 0.00343883
R486 GND.n89 GND.t20 0.00343883
R487 GND.n18 GND.n17 0.00343883
R488 GND.n17 GND.t22 0.00343883
R489 GND.n127 GND.n126 0.00308338
R490 GND.n9 GND.n8 0.003
R491 GND.n120 GND.n118 0.00258333
R492 GND.n41 GND.n39 0.00258333
R493 GND.n132 GND.n131 0.00245833
R494 GND.n21 GND.n19 0.00228571
R495 GND.n55 GND.n54 0.00183544
R496 GND.n54 GND.n53 0.00181454
R497 GND.n53 GND.t0 0.00181454
R498 GND.n63 GND.n2 0.00181454
R499 GND.t10 GND.n2 0.00181454
R500 GND.n104 GND.n103 0.00131092
R501 GND.n103 GND.n102 0.00131092
R502 GND.n98 GND.n97 0.00131092
R503 GND.n97 GND.n96 0.00131092
R504 GND.n128 GND.n127 0.00100184
R505 GND.n41 GND.n40 0.000530554
R506 GND.n73 GND.n72 0.00052846
R507 GND.n21 GND.n20 0.00052846
R508 GND.n91 GND.n90 0.0005264
R509 GND.n64 GND.n63 0.000512627
R510 GND.n47 GND.n46 0.000512368
R511 GND.n99 GND.n98 0.000507826
R512 GND.n105 GND.n104 0.000507826
R513 GND.n129 GND.n128 0.000504863
R514 GND.n133 GND.n132 0.000501292
R515 GND.n134 GND.n133 0.000501292
C0 S VDD 2.9f
C1 x1.Y S 0.182f
C2 a_1583_n1177# QN 0.29f
C3 R QN 1.55f
C4 a_1070_n1178# QN 0.42f
C5 Q a_1583_n1177# 0.418f
C6 Q R 0.379f
C7 a_1583_n1177# VDD 0.0171f
C8 Q a_1070_n1178# 0.255f
C9 x2.Y QN 0.182f
C10 R VDD 2.62f
C11 a_1070_n1178# VDD 0.0207f
C12 x1.Y R 0.882f
C13 Q x2.Y 0.0178f
C14 x2.Y VDD 0.902f
C15 R S 0.136f
C16 x1.Y x2.Y 0.0254f
C17 S a_1070_n1178# 0.436f
C18 QN m3_2150_n210# 0.0416f
C19 x2.Y S 0.526f
C20 R a_1583_n1177# 0.28f
C21 m3_2150_n210# VDD 1.21f
C22 x2.Y R 0.0934f
C23 Q QN 2.02f
C24 QN VDD 2.6f
C25 x1.Y QN 0.0386f
C26 Q VDD 2.52f
C27 R m3_2150_n210# 0.114f
C28 Q x1.Y 0.17f
C29 S QN 0.444f
C30 x1.Y VDD 0.733f
C31 Q S 2.28f
C32 R GND 4.32f
C33 QN GND 4.31f
C34 Q GND 3.75f
C35 S GND 4.87f
C36 VDD GND 16.2f
C37 m3_2150_n210# GND 0.252f $ **FLOATING
C38 x2.Y GND 1.5f
C39 x1.Y GND 1.93f
C40 a_1583_n1177# GND 0.561f
C41 a_1070_n1178# GND 0.555f
C42 R.n7 GND 0.0157f
C43 R.t10 GND 0.035f
C44 R.n13 GND 0.033f
C45 R.n15 GND 0.0313f
C46 R.n17 GND 0.0489f
C47 R.n18 GND 0.296f
C48 R.t9 GND 0.0117f
C49 R.n19 GND 0.237f
C50 R.t1 GND 0.035f
C51 R.n23 GND 0.0312f
C52 R.n24 GND 0.0142f
C53 R.n25 GND 0.0142f
C54 R.n26 GND 0.0956f
C55 R.n27 GND 0.524f
C56 R.n28 GND 0.496f
C57 R.n39 GND 0.0124f
C58 R.n46 GND 0.0127f
C59 R.n47 GND 0.0136f
C60 R.n49 GND 0.0109f
C61 QN.t3 GND 0.0243f
C62 QN.t0 GND 0.0243f
C63 QN.n0 GND 0.331f
C64 QN.t2 GND 0.0144f
C65 QN.n1 GND 0.341f
C66 QN.t6 GND 0.0725f
C67 QN.t5 GND 0.0237f
C68 QN.n2 GND 1.14f
C69 QN.n3 GND 0.15f
C70 QN.t1 GND 0.0243f
C71 QN.n4 GND 0.227f
C72 QN.n5 GND 0.242f
C73 QN.n6 GND 0.318f
C74 QN.t4 GND 0.0267f
C75 QN.n7 GND 0.803f
C76 VDD.n1 GND 0.0161f
C77 VDD.t16 GND 0.0104f
C78 VDD.t11 GND 0.0104f
C79 VDD.t17 GND 0.0127f
C80 VDD.n7 GND 0.0155f
C81 VDD.t13 GND 0.0127f
C82 VDD.n8 GND 0.0155f
C83 VDD.n9 GND 0.0113f
C84 VDD.n12 GND 0.0191f
C85 VDD.n17 GND 0.0191f
C86 VDD.n20 GND 0.0191f
C87 VDD.n21 GND 0.0213f
C88 VDD.n22 GND 0.0143f
C89 VDD.n23 GND 0.0271f
C90 VDD.n25 GND 0.138f
C91 VDD.t8 GND 0.107f
C92 VDD.t0 GND 0.108f
C93 VDD.n30 GND 0.04f
C94 VDD.n31 GND 0.0132f
C95 VDD.n35 GND 0.0398f
C96 VDD.n36 GND 0.0136f
C97 VDD.n40 GND 0.0236f
C98 VDD.n41 GND 0.0523f
C99 VDD.n42 GND 0.0156f
C100 VDD.n47 GND 0.0104f
C101 VDD.n48 GND 0.0943f
C102 VDD.n51 GND 0.0193f
C103 VDD.n52 GND 0.0224f
C104 VDD.n53 GND 0.138f
C105 VDD.n59 GND 0.141f
C106 VDD.n60 GND 0.144f
C107 VDD.n61 GND 0.156f
C108 VDD.n62 GND 0.016f
C109 VDD.n67 GND 0.173f
C110 VDD.n68 GND 0.146f
C111 VDD.n69 GND 0.0196f
C112 VDD.n71 GND 0.0216f
C113 VDD.n72 GND 0.0853f
C114 VDD.n73 GND 0.0137f
C115 VDD.n74 GND 0.0137f
C116 VDD.t2 GND 0.0749f
C117 VDD.n77 GND 0.179f
C118 VDD.n80 GND 0.0401f
C119 VDD.n82 GND 0.0262f
C120 VDD.n83 GND 0.0211f
C121 VDD.n84 GND 0.0142f
C122 VDD.n85 GND 0.0262f
C123 VDD.n86 GND 0.0215f
C124 VDD.n87 GND 0.0192f
C125 VDD.n88 GND 0.0136f
C126 VDD.n89 GND 0.0136f
C127 VDD.t14 GND 0.0749f
C128 VDD.n92 GND 0.0198f
C129 VDD.n93 GND 0.179f
C130 VDD.n96 GND 0.0403f
C131 VDD.n97 GND 0.0854f
C132 VDD.n98 GND 0.0103f
C133 VDD.n99 GND 0.0946f
C134 VDD.n102 GND 0.0222f
C135 VDD.n103 GND 0.138f
C136 VDD.n109 GND 0.0237f
C137 VDD.n110 GND 0.0739f
C138 VDD.n111 GND 0.129f
C139 VDD.n112 GND 0.02f
C140 VDD.t22 GND 0.107f
C141 VDD.n116 GND 0.0745f
C142 VDD.t18 GND 0.0761f
C143 VDD.n117 GND 0.0118f
C144 VDD.n118 GND 0.0122f
C145 VDD.n119 GND 0.0381f
C146 VDD.n120 GND 0.0126f
C147 VDD.n124 GND 0.0451f
C148 VDD.n127 GND 0.0148f
C149 VDD.n128 GND 0.0523f
C150 VDD.n129 GND 0.0156f
C151 VDD.n133 GND 0.11f
C152 VDD.n134 GND 0.0169f
C153 VDD.n139 GND 0.0509f
C154 VDD.n140 GND 1.28f
C155 VDD.n141 GND 1.14f
C156 VDD.n142 GND 0.315f
C157 VDD.n143 GND 0.0556f
C158 VDD.n144 GND 0.0573f
C159 VDD.n145 GND 2.33f
C160 VDD.n146 GND 0.378f
C161 VDD.n147 GND 0.202f
C162 VDD.t10 GND 0.105f
C163 VDD.t6 GND 0.0628f
C164 VDD.t4 GND 0.0628f
C165 VDD.t12 GND 0.0597f
C166 Q.t4 GND 0.0559f
C167 Q.t5 GND 0.0933f
C168 Q.t6 GND 0.0317f
C169 Q.n0 GND 1.44f
C170 Q.n1 GND 0.0773f
C171 Q.n2 GND 0.1f
C172 Q.n3 GND 0.439f
C173 Q.n4 GND 0.0129f
C174 Q.t0 GND 0.0317f
C175 Q.n5 GND 0.107f
C176 Q.n6 GND 0.0336f
C177 Q.n7 GND 0.129f
C178 Q.n8 GND 0.345f
C179 Q.t3 GND 0.0317f
C180 Q.t1 GND 0.0317f
C181 Q.n9 GND 0.147f
C182 Q.n10 GND 0.846f
C183 Q.n11 GND 2.6f
C184 S.n2 GND 0.0165f
C185 S.t9 GND 0.0177f
C186 S.t7 GND 0.0104f
C187 S.n7 GND 0.0295f
C188 S.n11 GND 0.0165f
C189 S.n13 GND 0.0496f
C190 S.t0 GND 0.0658f
C191 S.n15 GND 0.0569f
C192 S.n16 GND 0.0106f
C193 S.n17 GND 0.103f
C194 S.n18 GND 0.648f
C195 S.t4 GND 0.0239f
C196 S.t3 GND 0.0658f
C197 S.n19 GND 0.277f
C198 S.n20 GND 0.676f
C199 S.n21 GND 0.966f
C200 S.n22 GND 0.949f
C201 S.n25 GND 0.0152f
C202 S.n30 GND 0.0162f
C203 S.n31 GND 0.0197f
C204 S.t5 GND 0.0177f
C205 S.t6 GND 0.0104f
C206 S.n33 GND 0.0233f
C207 S.n34 GND 0.0117f
C208 S.n38 GND 0.0144f
C209 S.n39 GND 0.0159f
C210 S.t10 GND 0.0177f
C211 S.t8 GND 0.0104f
C212 S.n40 GND 0.0239f
C213 S.t2 GND 0.0177f
C214 S.t1 GND 0.0104f
C215 S.n41 GND 0.0255f
C216 S.n42 GND 0.012f
C217 S.n43 GND 0.0293f
.ends

