* NGSPICE file created from flashADC_flat.ext - technology: sky130A

.subckt flashADC_flat VL VV11 VV12 VV15 S0 S1 I0 VV16 I3 VV6 VV8 VV10 I13 VV14 I5
+ VV3 I4 VV9 I11 VV4 VV1 I10 I1 I2 I6 OUT3 OUT2 VV7 VV2 I12 I9 R1 OUT1 VFS I14 VV5
+ VV13 I8 OUT0 R0 CLK I15 VIN GND VDD I7
X0 GND.t1270 frontAnalog_v0p0p1_7.x65.X frontAnalog_v0p0p1_7.RSfetsym_0.x2.Y GND.t1269 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 OUT3.t127 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD.t332 VDD.t331 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 VDD.t132 R0.t4 a_57123_n85079# VDD.t131 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X3 GND.t986 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t63 GND.t985 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 VDD.t790 frontAnalog_v0p0p1_10.x63.X I5.t3 VDD.t785 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.25
X5 VDD.t1054 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t127 VDD.t1053 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 VFS.t4 VV16.t9 GND.t122 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X7 a_78315_n41309# 16to4_PriorityEncoder_v0p0p1_0.x5.x11.X a_78243_n41309# VDD.t410 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X8 a_16719_n13117.t23 a_16599_n13205.t4 a_16541_n13117.t21 GND.t729 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X9 w_55000_n56928# CLK.t0 frontAnalog_v0p0p1_10.x65.A.t1 VDD.t562 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X10 VV4.t8 VV3.t7 GND.t106 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X11 frontAnalog_v0p0p1_3.x65.X a_57123_n13359# VDD.t1298 VDD.t1297 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X12 VDD.t1104 frontAnalog_v0p0p1_9.x63.X frontAnalog_v0p0p1_9.RSfetsym_0.x1.Y VDD.t1097 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13 OUT3.t63 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND.t343 GND.t342 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X14 S1.t2 R1.t4 a_55268_n79536# GND.t819 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X15 OUT2.t63 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND.t1114 GND.t1113 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X16 frontAnalog_v0p0p1_5.RSfetsym_0.QN.t1 frontAnalog_v0p0p1_5.RSfetsym_0.x1.Y GND.t1247 GND.t1196 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.25
X17 16to4_PriorityEncoder_v0p0p1_0.x29.A 16to4_PriorityEncoder_v0p0p1_0.x28.A VDD.t1080 VDD.t1079 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X18 VV11.t10 VV10.t9 GND.t24 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X19 frontAnalog_v0p0p1_6.x63.X a_57123_n31079# GND.t720 GND.t719 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X20 GND.t341 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t62 GND.t340 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X21 GND.t814 frontAnalog_v0p0p1_8.x63.X frontAnalog_v0p0p1_8.RSfetsym_0.x1.Y GND.t809 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X22 GND.t1112 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t62 GND.t1111 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X23 OUT3.t126 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD.t330 VDD.t329 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X24 VV2.t10 VV1.t12 GND.t52 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X25 a_53630_n84996# VV1.t16 w_55000_n83928# GND.t1239 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X26 16to4_PriorityEncoder_v0p0p1_0.x29.Y 16to4_PriorityEncoder_v0p0p1_0.x29.A GND.t565 GND.t564 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X27 GND.t1140 I0.t5 a_77605_n47345# GND.t154 sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X28 VDD.t926 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t127 VDD.t925 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X29 VDD.t328 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t125 VDD.t327 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X30 a_55268_n63336# CLK.t1 GND.t589 GND.t588 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X31 GND.t1388 16to4_PriorityEncoder_v0p0p1_0.x5.x17.A a_78349_n43045# GND.t175 sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X32 frontAnalog_v0p0p1_14.RSfetsym_0.x1.Y frontAnalog_v0p0p1_14.x63.X VDD.t354 VDD.t347 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X33 a_77605_n51335# I2.t5 VDD.t334 VDD.t333 sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.109 ps=1.36 w=0.42 l=0.15
X34 frontAnalog_v0p0p1_5.RSfetsym_0.x1.Y frontAnalog_v0p0p1_5.x63.X GND.t30 GND.t26 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X35 VDD.t789 frontAnalog_v0p0p1_10.x63.X frontAnalog_v0p0p1_10.RSfetsym_0.x1.Y VDD.t783 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X36 VDD.t1181 VDD.t1179 a_77605_n43295# VDD.t1180 sky130_fd_pr__pfet_01v8_hvt ad=0.312 pd=1.68 as=0.0588 ps=0.7 w=0.42 l=0.15
X37 VDD.t1464 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t127 VDD.t1463 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X38 GND.t339 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t61 GND.t338 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X39 GND.t683 frontAnalog_v0p0p1_8.RSfetsym_0.QN.t5 a_59577_n46683# GND.t682 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X40 GND.t1110 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t61 GND.t1109 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X41 GND.t745 I5.t5 a_59578_n56970# GND.t744 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X42 a_53630_n41796# VV9.t16 w_55000_n40728# GND.t162 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X43 VDD.t1052 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t126 VDD.t1051 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X44 VV16.t7 VV15.t9 GND.t51 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X45 OUT1.t63 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND.t1528 GND.t1527 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X46 GND.t199 frontAnalog_v0p0p1_12.x65.X frontAnalog_v0p0p1_12.RSfetsym_0.x2.Y GND.t198 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X47 OUT2.t125 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD.t1050 VDD.t1049 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X48 GND.t563 16to4_PriorityEncoder_v0p0p1_0.x29.A 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND.t562 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X49 frontAnalog_v0p0p1_7.RSfetsym_0.x1.Y frontAnalog_v0p0p1_7.x63.X VDD.t555 VDD.t548 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X50 OUT0.t62 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND.t984 GND.t983 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X51 a_77637_n50057# 16to4_PriorityEncoder_v0p0p1_0.x3.EI VDD.t1249 VDD.t459 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X52 frontAnalog_v0p0p1_2.x65.A.t2 frontAnalog_v0p0p1_2.x63.A.t4 a_55268_n3936# GND.t70 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X53 VDD.t199 frontAnalog_v0p0p1_15.x65.X frontAnalog_v0p0p1_15.RSfetsym_0.QN.t1 VDD.t195 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.25
X54 GND.t337 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t60 GND.t336 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X55 GND.t982 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t61 GND.t981 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X56 a_82906_n51645# 16to4_PriorityEncoder_v0p0p1_0.x3.A0 GND.t167 GND.t166 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X57 OUT3.t124 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD.t326 VDD.t325 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X58 VV6.t13 VV5.t11 GND.t24 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X59 frontAnalog_v0p0p1_6.RSfetsym_0.QN.t4 I10.t5 VDD.t126 VDD.t125 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.3
X60 a_77881_n44527# 16to4_PriorityEncoder_v0p0p1_0.x5.x18.C a_77775_n44527# GND.t528 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X61 GND.t775 I13.t5 a_59578_n13770# GND.t774 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X62 OUT3.t59 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND.t335 GND.t334 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X63 16to4_PriorityEncoder_v0p0p1_0.x36.Y 16to4_PriorityEncoder_v0p0p1_0.x36.A GND.t1565 GND.t1564 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X64 a_53630_n9396# frontAnalog_v0p0p1_10.IB.t3 GND.t385 GND.t384 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X65 VDD.t324 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t123 VDD.t323 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X66 VDD.t55 frontAnalog_v0p0p1_2.x63.A.t5 a_57123_n4079# VDD.t54 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X67 frontAnalog_v0p0p1_11.x63.X a_57123_n63479# VDD.t489 VDD.t488 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X68 a_77723_n41087# VDD.t1502 a_77637_n41087# GND.t695 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X69 VV14.t5 VV13.t3 GND.t24 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X70 GND.t12 frontAnalog_v0p0p1_6.x65.X frontAnalog_v0p0p1_6.RSfetsym_0.x2.Y GND.t11 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X71 GND.t1355 16to4_PriorityEncoder_v0p0p1_0.x21.A 16to4_PriorityEncoder_v0p0p1_0.x22.A GND.t1354 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X72 w_55000_n79150# VIN.t0 a_53630_n79596# GND.t854 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X73 GND.t502 frontAnalog_v0p0p1_15.x63.X frontAnalog_v0p0p1_15.RSfetsym_0.x1.Y GND.t497 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X74 VIN.t1 w_55000_n51528# error sky130_fd_pr__cap_var_lvt w=2 l=0.18
X75 GND.t1526 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t62 GND.t1525 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X76 16to4_PriorityEncoder_v0p0p1_0.x5.x19.X a_77605_n44779# VDD.t1321 VDD.t1320 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.312 ps=1.68 w=1 l=0.15
X77 OUT2.t124 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD.t1048 VDD.t1047 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X78 VV4.t6 VV3.t6 GND.t77 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X79 16to4_PriorityEncoder_v0p0p1_0.x43.Y 16to4_PriorityEncoder_v0p0p1_0.x43.A VDD.t644 VDD.t643 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X80 VDD.t1145 frontAnalog_v0p0p1_4.x65.A.t4 a_57123_n18759# VDD.t1144 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X81 VV10.t14 VV9.t13 GND.t52 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X82 OUT0.t126 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD.t924 VDD.t923 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X83 a_78065_n41309# 16to4_PriorityEncoder_v0p0p1_0.x5.x22.A GND.t427 GND.t426 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X84 OUT0.t60 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND.t980 GND.t979 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X85 GND.t978 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t59 GND.t977 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X86 VV3.t5 VV2.t4 GND.t422 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X87 VDD.t1248 16to4_PriorityEncoder_v0p0p1_0.x3.EI a_77605_n51335# VDD.t1247 sky130_fd_pr__pfet_01v8_hvt ad=0.312 pd=1.68 as=0.0588 ps=0.7 w=0.42 l=0.15
X88 VV13.t2 VV12.t2 GND.t52 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X89 VDD.t922 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t125 VDD.t921 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X90 OUT3.t58 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND.t333 GND.t332 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X91 frontAnalog_v0p0p1_9.x65.A.t2 CLK.t2 frontAnalog_v0p0p1_9.x63.A.t1 VDD.t142 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X92 OUT2.t60 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND.t1108 GND.t1107 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X93 frontAnalog_v0p0p1_12.RSfetsym_0.x2.Y frontAnalog_v0p0p1_12.x65.X VDD.t190 VDD.t185 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X94 VDD.t322 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t122 VDD.t321 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X95 frontAnalog_v0p0p1_4.x63.X a_57123_n20279# VDD.t500 VDD.t499 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X96 GND.t1524 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t61 GND.t1523 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X97 w_55000_n35950# VIN.t2 a_53630_n36396# GND.t127 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X98 GND.t182 frontAnalog_v0p0p1_1.x63.X frontAnalog_v0p0p1_1.RSfetsym_0.x1.Y GND.t177 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X99 frontAnalog_v0p0p1_10.RSfetsym_0.x2.Y frontAnalog_v0p0p1_10.x65.X GND.t103 GND.t102 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X100 GND.t331 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t57 GND.t330 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X101 VDD.t699 I5.t6 a_77637_n49127# VDD.t698 sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X102 GND.t1563 16to4_PriorityEncoder_v0p0p1_0.x36.A 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND.t1562 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X103 VDD.t1296 16to4_PriorityEncoder_v0p0p1_0.x21.A 16to4_PriorityEncoder_v0p0p1_0.x22.A VDD.t1295 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X104 frontAnalog_v0p0p1_2.RSfetsym_0.x1.Y frontAnalog_v0p0p1_2.x63.X GND.t58 GND.t53 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X105 VDD.t1499 16to4_PriorityEncoder_v0p0p1_0.x36.A 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD.t1498 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X106 a_16541_n13117.t1 GND.t1271 GND.t392 sky130_fd_pr__res_xhigh_po_5p73 l=85.8
X107 I1.t3 frontAnalog_v0p0p1_14.RSfetsym_0.x2.Y GND.t437 GND.t436 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.25
X108 GND.t691 frontAnalog_v0p0p1_9.x65.A.t4 a_57123_n51159# GND.t690 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X109 VV3.t11 VV2.t11 GND.t214 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X110 VDD.t732 I13.t6 a_77605_n45765# VDD.t731 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X111 a_77881_n52567# 16to4_PriorityEncoder_v0p0p1_0.x3.x18.C a_77775_n52567# GND.t153 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X112 16to4_PriorityEncoder_v0p0p1_0.x22.Y 16to4_PriorityEncoder_v0p0p1_0.x22.A GND.t469 GND.t468 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X113 frontAnalog_v0p0p1_9.x63.A.t2 frontAnalog_v0p0p1_9.x65.A.t5 a_55268_n52536# GND.t692 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X114 OUT2.t123 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD.t1046 VDD.t1045 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X115 OUT0.t124 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD.t920 VDD.t919 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X116 VDD.t918 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t123 VDD.t917 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X117 I6.t0 frontAnalog_v0p0p1_9.RSfetsym_0.QN.t5 VDD.t1143 VDD.t1141 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.3
X118 frontAnalog_v0p0p1_6.RSfetsym_0.x2.Y frontAnalog_v0p0p1_6.x65.X VDD.t13 VDD.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X119 GND.t653 16to4_PriorityEncoder_v0p0p1_0.x43.A 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND.t652 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X120 GND.t1522 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t60 GND.t1521 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X121 OUT2.t122 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD.t1044 VDD.t1043 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X122 frontAnalog_v0p0p1_3.RSfetsym_0.x2.Y frontAnalog_v0p0p1_3.x65.X GND.t574 GND.t573 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X123 a_77639_n42341# VDD.t1176 VDD.t1178 VDD.t1177 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X124 frontAnalog_v0p0p1_13.RSfetsym_0.x1.Y frontAnalog_v0p0p1_13.x63.X GND.t383 GND.t379 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X125 a_59577_n57483# frontAnalog_v0p0p1_10.x63.X I5.t1 GND.t847 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X126 a_59578_n67770# frontAnalog_v0p0p1_13.x65.X frontAnalog_v0p0p1_13.RSfetsym_0.QN.t1 GND.t1208 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.315 ps=2.72 w=1 l=0.15
X127 a_77687_n45765# I13.t7 a_77605_n45765# GND.t1175 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X128 16to4_PriorityEncoder_v0p0p1_0.x42.A 16to4_PriorityEncoder_v0p0p1_0.x5.GS VDD.t394 VDD.t393 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X129 16to4_PriorityEncoder_v0p0p1_0.x3.x19.X a_77605_n52819# VDD.t381 VDD.t380 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.312 ps=1.68 w=1 l=0.15
X130 VV2.t7 VV1.t5 GND.t202 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X131 VDD.t1042 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t121 VDD.t1041 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X132 OUT1.t59 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND.t1520 GND.t1519 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X133 frontAnalog_v0p0p1_7.x63.A.t3 frontAnalog_v0p0p1_7.x65.A.t4 VDD.t1301 VDD.t1186 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X134 I9.t4 frontAnalog_v0p0p1_7.RSfetsym_0.x2.Y GND.t674 GND.t183 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.25
X135 VV7.t16 w_55000_n52150# error sky130_fd_pr__cap_var_lvt w=2 l=0.18
X136 a_16719_n13117.t22 a_16599_n13205.t5 a_16541_n13117.t7 GND.t730 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X137 16to4_PriorityEncoder_v0p0p1_0.x5.x11.X a_77637_n41087# GND.t69 GND.t68 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.112 ps=1.04 w=0.65 l=0.15
X138 OUT0.t58 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND.t976 GND.t975 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X139 GND.t1210 16to4_PriorityEncoder_v0p0p1_0.x3.x14.A a_78065_n49349# GND.t1209 sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X140 a_78703_n45515# 16to4_PriorityEncoder_v0p0p1_0.x5.x19.X a_78607_n45515# VDD.t456 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X141 frontAnalog_v0p0p1_2.x65.X a_57123_n2559# GND.t396 GND.t395 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X142 16to4_PriorityEncoder_v0p0p1_0.x22.Y 16to4_PriorityEncoder_v0p0p1_0.x22.A VDD.t455 VDD.t454 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X143 a_16719_n13117.t3 a_16719_n13117.t2 a_16599_n13205.t0 GND.t1246 sky130_fd_pr__nfet_01v8_lvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X144 VDD.t1336 frontAnalog_v0p0p1_8.x65.X frontAnalog_v0p0p1_8.RSfetsym_0.x2.Y VDD.t1329 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X145 GND.t329 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t56 GND.t328 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X146 GND.t467 16to4_PriorityEncoder_v0p0p1_0.x22.A 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND.t466 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X147 VDD.t1040 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t120 VDD.t1039 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X148 VDD.t580 frontAnalog_v0p0p1_13.x63.A.t4 a_57123_n68879# VDD.t579 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X149 a_59577_n14283# frontAnalog_v0p0p1_3.x63.X I13.t1 GND.t487 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X150 a_59578_n24570# frontAnalog_v0p0p1_5.x65.X frontAnalog_v0p0p1_5.RSfetsym_0.QN.t4 GND.t1380 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.315 ps=2.72 w=1 l=0.15
X151 16to4_PriorityEncoder_v0p0p1_0.x29.Y 16to4_PriorityEncoder_v0p0p1_0.x29.A GND.t561 GND.t560 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X152 VV7.t1 VV6.t1 GND.t33 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X153 I6.t3 frontAnalog_v0p0p1_9.x63.X VDD.t1103 VDD.t1100 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.25
X154 a_53630_n63396# frontAnalog_v0p0p1_10.IB.t4 GND.t386 GND.t36 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X155 16to4_PriorityEncoder_v0p0p1_0.x5.x22.A a_77639_n42341# VDD.t341 VDD.t340 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.167 ps=1.39 w=1 l=0.15
X156 frontAnalog_v0p0p1_0.RSfetsym_0.x1.Y frontAnalog_v0p0p1_0.x63.X GND.t373 GND.t369 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X157 16to4_PriorityEncoder_v0p0p1_0.x43.Y 16to4_PriorityEncoder_v0p0p1_0.x43.A GND.t651 GND.t650 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X158 VDD.t564 frontAnalog_v0p0p1_10.x63.A.t4 frontAnalog_v0p0p1_10.x65.A.t2 VDD.t563 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X159 OUT2.t59 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND.t1106 GND.t1105 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X160 frontAnalog_v0p0p1_0.RSfetsym_0.x2.Y frontAnalog_v0p0p1_0.x65.X GND.t50 GND.t49 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X161 OUT1.t126 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD.t1462 VDD.t1461 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X162 w_55000_n8950# VIN.t3 a_53630_n9396# GND.t818 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X163 VDD.t701 I5.t7 a_77605_n53805# VDD.t700 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X164 frontAnalog_v0p0p1_12.x65.X a_57123_n72759# GND.t620 GND.t619 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X165 VDD.t1460 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t125 VDD.t1459 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X166 OUT0.t122 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD.t916 VDD.t915 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X167 frontAnalog_v0p0p1_4.RSfetsym_0.x2.Y frontAnalog_v0p0p1_4.x65.X GND.t496 GND.t495 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X168 GND.t327 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t55 GND.t326 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X169 VDD.t404 frontAnalog_v0p0p1_5.x63.A.t4 a_57123_n25679# VDD.t403 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X170 GND.t974 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t57 GND.t973 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X171 a_53630_n20196# frontAnalog_v0p0p1_10.IB.t5 GND.t387 GND.t36 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X172 a_77639_n50381# 16to4_PriorityEncoder_v0p0p1_0.x3.EI VDD.t1246 VDD.t1245 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X173 VDD.t1497 16to4_PriorityEncoder_v0p0p1_0.x36.A 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD.t1496 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X174 VDD.t453 16to4_PriorityEncoder_v0p0p1_0.x22.A 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD.t452 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X175 VDD.t104 frontAnalog_v0p0p1_3.x63.A.t4 frontAnalog_v0p0p1_3.x65.A.t3 VDD.t103 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X176 OUT3.t54 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND.t325 GND.t324 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X177 VDD.t134 S0.t4 a_57123_n83559# VDD.t133 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X178 GND.t820 R1.t5 a_57123_n79679# GND.t608 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X179 a_55268_n47136# CLK.t3 GND.t159 GND.t158 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X180 frontAnalog_v0p0p1_1.RSfetsym_0.x2.Y frontAnalog_v0p0p1_1.x65.X GND.t756 GND.t755 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X181 VDD.t189 frontAnalog_v0p0p1_12.x65.X frontAnalog_v0p0p1_12.RSfetsym_0.x2.Y VDD.t185 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X182 GND.t1341 16to4_PriorityEncoder_v0p0p1_0.x3.x15.X a_78349_n51085# GND.t14 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X183 frontAnalog_v0p0p1_4.x65.A.t2 frontAnalog_v0p0p1_4.x63.A.t4 a_55268_n20136# GND.t806 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X184 frontAnalog_v0p0p1_9.RSfetsym_0.QN.t1 I6.t5 VDD.t1142 VDD.t1141 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.3
X185 OUT3.t121 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD.t320 VDD.t319 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X186 VV10.t15 VV9.t14 GND.t202 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X187 a_78703_n53555# 16to4_PriorityEncoder_v0p0p1_0.x3.x19.X a_78607_n53555# VDD.t86 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X188 GND.t972 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t56 GND.t971 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X189 OUT1.t58 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND.t1518 GND.t1517 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X190 VV12.t1 VV11.t0 GND.t123 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X191 VV3.t4 VV2.t2 GND.t394 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X192 a_77775_n51335# 16to4_PriorityEncoder_v0p0p1_0.x3.x19.C a_77687_n51335# GND.t346 sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
X193 16to4_PriorityEncoder_v0p0p1_0.x43.A 16to4_PriorityEncoder_v0p0p1_0.x42.A VDD.t402 VDD.t401 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X194 a_53630_n25596# VV12.t16 w_55000_n24528# GND.t606 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X195 VV13.t6 VV12.t5 GND.t202 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X196 OUT3.t53 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND.t323 GND.t322 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X197 16to4_PriorityEncoder_v0p0p1_0.x28.A 16to4_PriorityEncoder_v0p0p1_0.x1.X GND.t681 GND.t680 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X198 VDD.t914 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t121 VDD.t913 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X199 VDD.t1038 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t119 VDD.t1037 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X200 frontAnalog_v0p0p1_9.RSfetsym_0.x2.Y frontAnalog_v0p0p1_9.x65.X VDD.t1275 VDD.t1270 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X201 VDD.t158 frontAnalog_v0p0p1_1.x65.A.t4 a_57123_n40359# VDD.t157 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X202 GND.t1279 frontAnalog_v0p0p1_7.x63.A.t4 a_57123_n36479# GND.t1278 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X203 frontAnalog_v0p0p1_10.RSfetsym_0.QN.t3 frontAnalog_v0p0p1_10.x65.X VDD.t85 VDD.t81 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.25
X204 frontAnalog_v0p0p1_9.RSfetsym_0.x1.Y frontAnalog_v0p0p1_9.x63.X GND.t1193 GND.t1188 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X205 VDD.t12 frontAnalog_v0p0p1_6.x65.X frontAnalog_v0p0p1_6.RSfetsym_0.x2.Y VDD.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X206 16to4_PriorityEncoder_v0p0p1_0.x36.Y 16to4_PriorityEncoder_v0p0p1_0.x36.A VDD.t1495 VDD.t1494 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X207 VDD.t458 I4.t5 a_77637_n48817# VDD.t457 sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X208 VDD.t1458 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t124 VDD.t1457 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X209 VDD.t1116 frontAnalog_v0p0p1_13.x65.X frontAnalog_v0p0p1_13.RSfetsym_0.QN.t3 VDD.t1112 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.25
X210 GND.t970 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t55 GND.t969 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X211 VDD.t912 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t120 VDD.t911 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X212 frontAnalog_v0p0p1_11.RSfetsym_0.x1.Y frontAnalog_v0p0p1_11.x63.X VDD.t497 VDD.t492 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X213 OUT0.t54 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND.t968 GND.t967 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X214 VFS.t3 VV16.t8 GND.t59 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X215 frontAnalog_v0p0p1_3.RSfetsym_0.QN.t2 frontAnalog_v0p0p1_3.x65.X VDD.t545 VDD.t541 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.25
X216 VDD.t400 16to4_PriorityEncoder_v0p0p1_0.x42.A 16to4_PriorityEncoder_v0p0p1_0.x43.A VDD.t399 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X217 VDD.t1456 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t123 VDD.t1455 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X218 VV4.t3 VV3.t3 GND.t51 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X219 VV15.t16 w_55000_n8950# error sky130_fd_pr__cap_var_lvt w=2 l=0.18
X220 16to4_PriorityEncoder_v0p0p1_0.x5.x17.A a_77637_n42017# GND.t352 GND.t351 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.112 ps=1.04 w=0.65 l=0.15
X221 VDD.t1313 frontAnalog_v0p0p1_5.x65.X frontAnalog_v0p0p1_5.RSfetsym_0.QN.t3 VDD.t1309 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.25
X222 VV15.t14 VV14.t15 GND.t106 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X223 GND.t372 frontAnalog_v0p0p1_0.x63.X frontAnalog_v0p0p1_0.RSfetsym_0.x1.Y GND.t369 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X224 VDD.t318 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t120 VDD.t317 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X225 16to4_PriorityEncoder_v0p0p1_0.x22.Y 16to4_PriorityEncoder_v0p0p1_0.x22.A GND.t465 GND.t464 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X226 VDD.t910 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t119 VDD.t909 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X227 a_16719_n13117.t21 a_16599_n13205.t6 a_16541_n13117.t6 GND.t731 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X228 frontAnalog_v0p0p1_7.x65.A.t3 CLK.t4 frontAnalog_v0p0p1_7.x63.A.t1 VDD.t143 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X229 VV7.t6 VV6.t7 GND.t78 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X230 VDD.t353 frontAnalog_v0p0p1_14.x63.X frontAnalog_v0p0p1_14.RSfetsym_0.x1.Y VDD.t347 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X231 frontAnalog_v0p0p1_6.x63.A.t3 CLK.t5 w_55000_n30550# VDD.t144 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X232 GND.t29 frontAnalog_v0p0p1_5.x63.X frontAnalog_v0p0p1_5.RSfetsym_0.x1.Y GND.t26 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X233 OUT2.t118 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD.t1036 VDD.t1035 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X234 OUT0.t118 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD.t908 VDD.t907 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X235 a_78607_n45515# 16to4_PriorityEncoder_v0p0p1_0.x5.x20.X a_78525_n45515# VDD.t728 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X236 VDD.t358 frontAnalog_v0p0p1_2.x65.A.t4 a_57123_n2559# VDD.t357 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X237 frontAnalog_v0p0p1_11.x65.X a_57123_n61959# VDD.t719 VDD.t718 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X238 GND.t494 frontAnalog_v0p0p1_4.x65.X frontAnalog_v0p0p1_4.RSfetsym_0.x2.Y GND.t493 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X239 frontAnalog_v0p0p1_10.x63.X a_57123_n58079# GND.t675 GND.t75 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X240 OUT1.t122 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD.t1454 VDD.t1453 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X241 frontAnalog_v0p0p1_9.x63.A.t0 CLK.t6 w_55000_n52150# VDD.t145 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X242 VDD.t146 CLK.t7 w_55000_n73128# GND.t160 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X243 GND.t1366 frontAnalog_v0p0p1_7.x65.A.t5 a_57123_n34959# GND.t1278 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X244 frontAnalog_v0p0p1_12.RSfetsym_0.QN.t3 frontAnalog_v0p0p1_12.RSfetsym_0.x1.Y GND.t503 GND.t187 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.25
X245 GND.t1104 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t58 GND.t1103 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X246 16to4_PriorityEncoder_v0p0p1_0.x5.x16.X a_77605_n43545# GND.t857 GND.t856 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.196 ps=1.33 w=0.65 l=0.15
X247 GND.t1516 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t57 GND.t1515 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X248 GND.t754 frontAnalog_v0p0p1_1.x65.X frontAnalog_v0p0p1_1.RSfetsym_0.x2.Y GND.t753 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X249 frontAnalog_v0p0p1_15.RSfetsym_0.x2.Y frontAnalog_v0p0p1_15.x65.X GND.t213 GND.t212 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X250 frontAnalog_v0p0p1_3.RSfetsym_0.x2.Y frontAnalog_v0p0p1_3.x65.X VDD.t544 VDD.t538 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X251 VDD.t554 frontAnalog_v0p0p1_7.x63.X frontAnalog_v0p0p1_7.RSfetsym_0.x1.Y VDD.t548 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X252 VDD.t496 frontAnalog_v0p0p1_11.x63.X I4.t3 VDD.t490 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.25
X253 VDD.t147 CLK.t8 w_55000_n73750# GND.t161 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X254 16to4_PriorityEncoder_v0p0p1_0.x22.Y 16to4_PriorityEncoder_v0p0p1_0.x22.A VDD.t451 VDD.t450 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X255 VV1.t8 VL.t4 GND.t52 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X256 w_55000_n62328# CLK.t9 frontAnalog_v0p0p1_11.x65.A.t1 VDD.t687 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X257 a_78243_n41309# 16to4_PriorityEncoder_v0p0p1_0.x5.x17.A a_78147_n41309# VDD.t410 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X258 OUT2.t117 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD.t1016 VDD.t1015 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X259 VDD.t1175 VDD.t1173 a_78649_n39527# VDD.t1174 sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X260 frontAnalog_v0p0p1_3.x63.X a_57123_n14879# GND.t93 GND.t92 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X261 OUT3.t52 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND.t321 GND.t320 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X262 VV10.t16 w_55000_n35950# error sky130_fd_pr__cap_var_lvt w=2 l=0.18
X263 S0.t0 R0.t5 a_55268_n84936# GND.t1228 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X264 a_53630_n68796# VV4.t16 w_55000_n67728# GND.t712 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X265 VDD.t1034 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t116 VDD.t1033 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X266 VV9.t3 VV8.t4 GND.t52 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X267 VDD.t316 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t119 VDD.t315 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X268 16to4_PriorityEncoder_v0p0p1_0.x3.x17.A a_77637_n50057# GND.t1306 GND.t1305 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.112 ps=1.04 w=0.65 l=0.15
X269 OUT0.t53 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND.t966 GND.t965 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X270 GND.t319 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t51 GND.t318 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X271 GND.t1192 frontAnalog_v0p0p1_9.x63.X frontAnalog_v0p0p1_9.RSfetsym_0.x1.Y GND.t1188 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X272 OUT3.t118 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD.t314 VDD.t313 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X273 16to4_PriorityEncoder_v0p0p1_0.x21.A 16to4_PriorityEncoder_v0p0p1_0.x2.X GND.t785 GND.t784 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X274 VIN.t4 w_55000_n8328# error sky130_fd_pr__cap_var_lvt w=2 l=0.18
X275 GND.t1224 16to4_PriorityEncoder_v0p0p1_0.x5.x21.B a_78183_n45737# GND.t1223 sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X276 VDD.t688 CLK.t10 w_55000_n30550# GND.t594 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X277 VDD.t124 frontAnalog_v0p0p1_4.x63.X I12.t2 VDD.t117 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.25
X278 w_55000_n19128# CLK.t11 frontAnalog_v0p0p1_4.x65.A.t1 VDD.t689 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X279 VDD.t642 16to4_PriorityEncoder_v0p0p1_0.x43.A 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD.t641 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X280 GND.t418 16to4_PriorityEncoder_v0p0p1_0.x42.A 16to4_PriorityEncoder_v0p0p1_0.x43.A GND.t417 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X281 GND.t1102 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t57 GND.t1101 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X282 a_78607_n53555# 16to4_PriorityEncoder_v0p0p1_0.x3.x20.X a_78525_n53555# VDD.t359 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X283 frontAnalog_v0p0p1_1.x65.A.t2 frontAnalog_v0p0p1_1.x63.A.t4 a_55268_n41736# GND.t1227 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X284 OUT2.t56 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND.t1100 GND.t1099 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X285 VDD.t495 frontAnalog_v0p0p1_11.x63.X frontAnalog_v0p0p1_11.RSfetsym_0.x1.Y VDD.t492 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X286 GND.t1514 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t56 GND.t1513 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X287 VV15.t5 VV14.t4 GND.t77 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X288 16to4_PriorityEncoder_v0p0p1_0.x3.x16.C I5.t8 GND.t747 GND.t746 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X289 OUT0.t117 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD.t906 VDD.t905 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X290 OUT3.t117 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD.t312 VDD.t311 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X291 GND.t101 frontAnalog_v0p0p1_10.x65.X frontAnalog_v0p0p1_10.RSfetsym_0.x2.Y GND.t100 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X292 VIN.t5 w_55000_n78528# error sky130_fd_pr__cap_var_lvt w=2 l=0.18
X293 OUT1.t55 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND.t1512 GND.t1511 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X294 frontAnalog_v0p0p1_4.RSfetsym_0.x1.Y frontAnalog_v0p0p1_4.x63.X VDD.t123 VDD.t119 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X295 VDD.t153 16to4_PriorityEncoder_v0p0p1_0.x1.A a_82988_n47995# VDD.t152 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X296 GND.t57 frontAnalog_v0p0p1_2.x63.X frontAnalog_v0p0p1_2.RSfetsym_0.x1.Y GND.t53 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X297 16to4_PriorityEncoder_v0p0p1_0.x21.A 16to4_PriorityEncoder_v0p0p1_0.x2.X VDD.t736 VDD.t735 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X298 a_77687_n44779# VDD.t1503 a_77605_n44779# GND.t678 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.109 ps=1.36 w=0.42 l=0.15
X299 a_77723_n42017# VDD.t1504 a_77637_n42017# GND.t696 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X300 VDD.t1244 16to4_PriorityEncoder_v0p0p1_0.x3.EI a_78649_n47567# VDD.t1243 sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X301 GND.t1098 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t55 GND.t1097 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X302 OUT2.t54 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND.t1096 GND.t1095 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X303 S1.t1 CLK.t12 R1.t1 VDD.t690 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X304 OUT2.t115 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD.t1032 VDD.t1031 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X305 16to4_PriorityEncoder_v0p0p1_0.x43.Y 16to4_PriorityEncoder_v0p0p1_0.x43.A VDD.t640 VDD.t639 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X306 frontAnalog_v0p0p1_8.x63.X a_57123_n47279# VDD.t1317 VDD.t1316 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X307 GND.t572 frontAnalog_v0p0p1_3.x65.X frontAnalog_v0p0p1_3.RSfetsym_0.x2.Y GND.t571 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X308 VIN.t6 w_55000_n35328# error sky130_fd_pr__cap_var_lvt w=2 l=0.18
X309 GND.t382 frontAnalog_v0p0p1_13.x63.X frontAnalog_v0p0p1_13.RSfetsym_0.x1.Y GND.t379 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X310 16to4_PriorityEncoder_v0p0p1_0.x43.Y 16to4_PriorityEncoder_v0p0p1_0.x43.A GND.t649 GND.t648 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X311 OUT1.t54 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND.t1510 GND.t1509 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X312 VDD.t1030 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t114 VDD.t1029 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X313 VDD.t310 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t116 VDD.t309 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X314 GND.t1336 16to4_PriorityEncoder_v0p0p1_0.x3.x21.B a_78183_n53777# GND.t1335 sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X315 a_53630_n74196# frontAnalog_v0p0p1_10.IB.t6 GND.t388 GND.t36 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X316 w_55000_n84550# VIN.t7 a_53630_n84996# GND.t1239 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X317 GND.t609 S1.t4 a_57123_n78159# GND.t608 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X318 OUT2.t53 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND.t1094 GND.t1093 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X319 VDD.t92 frontAnalog_v0p0p1_5.x65.A.t4 a_57123_n24159# VDD.t91 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X320 GND.t808 frontAnalog_v0p0p1_4.x63.A.t5 a_57123_n20279# GND.t807 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X321 R1.t2 S1.t5 a_55268_n79536# GND.t610 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X322 GND.t211 frontAnalog_v0p0p1_15.x65.X frontAnalog_v0p0p1_15.RSfetsym_0.x2.Y GND.t210 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X323 VDD.t1452 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t121 VDD.t1451 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X324 VDD.t543 frontAnalog_v0p0p1_3.x65.X frontAnalog_v0p0p1_3.RSfetsym_0.x2.Y VDD.t538 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X325 GND.t317 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t50 GND.t316 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X326 I1.t4 frontAnalog_v0p0p1_14.RSfetsym_0.QN.t5 VDD.t1066 VDD.t1065 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.3
X327 frontAnalog_v0p0p1_10.RSfetsym_0.x2.Y frontAnalog_v0p0p1_10.x65.X VDD.t84 VDD.t78 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X328 GND.t964 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t52 GND.t963 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X329 GND.t1561 16to4_PriorityEncoder_v0p0p1_0.x36.A 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND.t1560 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X330 w_55000_n19750# VIN.t8 a_53630_n20196# GND.t743 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X331 VDD.t1493 16to4_PriorityEncoder_v0p0p1_0.x36.A 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD.t1492 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X332 OUT3.t49 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND.t315 GND.t314 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X333 a_77881_n43295# 16to4_PriorityEncoder_v0p0p1_0.x5.x16.C a_77775_n43295# GND.t703 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X334 VDD.t1028 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t113 VDD.t1027 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X335 VDD.t308 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t115 VDD.t307 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X336 VV2.t15 VV1.t15 GND.t24 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X337 GND.t559 16to4_PriorityEncoder_v0p0p1_0.x29.A 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND.t558 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X338 VV2.t16 w_55000_n79150# error sky130_fd_pr__cap_var_lvt w=2 l=0.18
X339 w_55000_n41350# VIN.t9 a_53630_n41796# GND.t162 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X340 GND.t48 frontAnalog_v0p0p1_0.x65.X frontAnalog_v0p0p1_0.RSfetsym_0.x2.Y GND.t47 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X341 frontAnalog_v0p0p1_11.RSfetsym_0.x2.Y frontAnalog_v0p0p1_11.x65.X GND.t769 GND.t768 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X342 a_77723_n50057# 16to4_PriorityEncoder_v0p0p1_0.x3.EI a_77637_n50057# GND.t1304 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X343 GND.t679 16to4_PriorityEncoder_v0p0p1_0.x5.x19.D a_77881_n44779# GND.t678 sky130_fd_pr__nfet_01v8 ad=0.196 pd=1.33 as=0.0693 ps=0.75 w=0.42 l=0.15
X344 frontAnalog_v0p0p1_7.x63.A.t2 frontAnalog_v0p0p1_7.x65.A.t6 a_55268_n36336# GND.t1367 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X345 VV1.t6 VL.t2 GND.t202 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X346 VV11.t12 VV10.t10 GND.t106 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X347 I0.t4 frontAnalog_v0p0p1_15.RSfetsym_0.x2.Y GND.t520 GND.t519 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.25
X348 OUT1.t53 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND.t1508 GND.t1507 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X349 a_77775_n44527# I9.t5 a_77687_n44527# GND.t528 sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
X350 I9.t3 frontAnalog_v0p0p1_7.RSfetsym_0.QN.t5 VDD.t600 VDD.t504 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.3
X351 a_59578_n8370# frontAnalog_v0p0p1_0.x65.X frontAnalog_v0p0p1_0.RSfetsym_0.QN.t2 GND.t46 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.315 ps=2.72 w=1 l=0.15
X352 GND.t1092 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t52 GND.t1091 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X353 VDD.t1026 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t112 VDD.t1025 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X354 a_78147_n41309# 16to4_PriorityEncoder_v0p0p1_0.x5.x22.A a_78065_n41309# VDD.t410 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X355 VDD.t904 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t116 VDD.t903 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X356 OUT1.t52 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND.t1506 GND.t1505 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X357 OUT3.t48 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND.t313 GND.t312 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X358 I1.t2 frontAnalog_v0p0p1_14.x63.X VDD.t352 VDD.t349 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.25
X359 VV9.t12 VV8.t13 GND.t202 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X360 16to4_PriorityEncoder_v0p0p1_0.x36.Y 16to4_PriorityEncoder_v0p0p1_0.x36.A GND.t1559 GND.t1558 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X361 16to4_PriorityEncoder_v0p0p1_0.x36.Y 16to4_PriorityEncoder_v0p0p1_0.x36.A VDD.t1491 VDD.t1490 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X362 GND.t1504 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t51 GND.t1503 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X363 frontAnalog_v0p0p1_12.RSfetsym_0.x1.Y frontAnalog_v0p0p1_12.x63.X GND.t133 GND.t129 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X364 a_59577_n62883# frontAnalog_v0p0p1_11.x63.X I4.t1 GND.t511 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X365 I8.t4 frontAnalog_v0p0p1_1.RSfetsym_0.x2.Y GND.t757 GND.t526 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.25
X366 GND.t962 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t51 GND.t961 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X367 16to4_PriorityEncoder_v0p0p1_0.x3.x15.X a_77605_n51335# GND.t739 GND.t738 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.196 ps=1.33 w=0.65 l=0.15
X368 16to4_PriorityEncoder_v0p0p1_0.x43.Y 16to4_PriorityEncoder_v0p0p1_0.x43.A GND.t647 GND.t646 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X369 OUT0.t50 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND.t960 GND.t959 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X370 VDD.t691 CLK.t13 w_55000_n56928# GND.t732 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X371 GND.t1502 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t50 GND.t1501 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X372 a_53630_n47196# frontAnalog_v0p0p1_10.IB.t7 GND.t389 GND.t36 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X373 I9.t1 frontAnalog_v0p0p1_7.x63.X VDD.t553 VDD.t550 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.25
X374 OUT1.t120 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD.t1450 VDD.t1449 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X375 frontAnalog_v0p0p1_15.RSfetsym_0.x1.Y frontAnalog_v0p0p1_15.x63.X VDD.t487 VDD.t480 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X376 VDD.t1274 frontAnalog_v0p0p1_9.x65.X frontAnalog_v0p0p1_9.RSfetsym_0.x2.Y VDD.t1270 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X377 VDD.t1138 frontAnalog_v0p0p1_1.x63.A.t5 frontAnalog_v0p0p1_1.x65.A.t3 VDD.t1088 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X378 OUT2.t111 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD.t1024 VDD.t1023 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X379 frontAnalog_v0p0p1_6.RSfetsym_0.x1.Y frontAnalog_v0p0p1_6.x63.X GND.t616 GND.t612 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X380 frontAnalog_v0p0p1_13.RSfetsym_0.x2.Y frontAnalog_v0p0p1_13.x65.X GND.t1207 GND.t1206 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X381 16to4_PriorityEncoder_v0p0p1_0.x5.x14.A a_77637_n40777# VDD.t1131 VDD.t1130 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.167 ps=1.39 w=1 l=0.15
X382 VDD.t1448 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t119 VDD.t1447 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X383 16to4_PriorityEncoder_v0p0p1_0.x34.A a_82906_n43855# VDD.t1058 VDD.t1057 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.146 ps=1.34 w=1 l=0.15
X384 frontAnalog_v0p0p1_14.RSfetsym_0.QN.t1 I1.t5 VDD.t1215 VDD.t1065 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.3
X385 frontAnalog_v0p0p1_10.x65.X a_57123_n56559# GND.t76 GND.t75 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X386 GND.t19 I4.t6 a_59578_n62370# GND.t18 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X387 GND.t1235 frontAnalog_v0p0p1_9.RSfetsym_0.QN.t6 a_59577_n52083# GND.t1234 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X388 GND.t311 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t47 GND.t310 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X389 VV6.t3 VV5.t3 GND.t106 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X390 16to4_PriorityEncoder_v0p0p1_0.x5.x4.A VDD.t1505 GND.t698 GND.t697 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X391 a_77775_n52567# I1.t6 a_77687_n52567# GND.t153 sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
X392 VV10.t13 VV9.t11 GND.t24 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X393 a_16719_n13117.t20 a_16599_n13205.t7 a_16541_n13117.t5 GND.t721 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X394 VDD.t902 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t115 VDD.t901 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X395 VDD.t1078 16to4_PriorityEncoder_v0p0p1_0.x28.A 16to4_PriorityEncoder_v0p0p1_0.x29.A VDD.t1077 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X396 VDD.t692 CLK.t14 w_55000_n13728# GND.t597 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X397 OUT3.t46 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND.t309 GND.t308 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X398 VV3.t15 VV2.t14 GND.t123 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X399 OUT0.t49 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND.t958 GND.t957 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X400 OUT2.t51 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND.t1090 GND.t1089 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X401 VV14.t6 VV13.t5 GND.t106 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X402 VV13.t13 VV12.t14 GND.t24 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X403 16to4_PriorityEncoder_v0p0p1_0.x36.A 16to4_PriorityEncoder_v0p0p1_0.x35.A GND.t86 GND.t85 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X404 VDD.t306 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t114 VDD.t305 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X405 OUT0.t114 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD.t900 VDD.t899 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X406 GND.t557 16to4_PriorityEncoder_v0p0p1_0.x29.A 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND.t556 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X407 OUT2.t110 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD.t1022 VDD.t1021 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X408 frontAnalog_v0p0p1_1.RSfetsym_0.x1.Y frontAnalog_v0p0p1_1.x63.X VDD.t175 VDD.t168 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X409 frontAnalog_v0p0p1_14.RSfetsym_0.x2.Y frontAnalog_v0p0p1_14.x65.X VDD.t1128 VDD.t1123 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X410 GND.t307 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t45 GND.t306 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X411 GND.t645 16to4_PriorityEncoder_v0p0p1_0.x43.A 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND.t644 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X412 frontAnalog_v0p0p1_5.RSfetsym_0.x2.Y frontAnalog_v0p0p1_5.x65.X GND.t1379 GND.t1378 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X413 VDD.t586 frontAnalog_v0p0p1_13.x65.A.t4 a_57123_n67359# VDD.t585 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X414 frontAnalog_v0p0p1_14.RSfetsym_0.x1.Y frontAnalog_v0p0p1_14.x63.X GND.t358 GND.t353 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X415 VDD.t693 CLK.t15 w_55000_n14350# GND.t733 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X416 16to4_PriorityEncoder_v0p0p1_0.x5.x16.X a_77605_n43545# VDD.t797 VDD.t796 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.312 ps=1.68 w=1 l=0.15
X417 VDD.t83 frontAnalog_v0p0p1_10.x65.X frontAnalog_v0p0p1_10.RSfetsym_0.x2.Y VDD.t78 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X418 OUT1.t118 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD.t1446 VDD.t1445 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X419 VDD.t1444 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t117 VDD.t1443 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X420 frontAnalog_v0p0p1_7.RSfetsym_0.QN.t0 I9.t6 VDD.t505 VDD.t504 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.3
X421 frontAnalog_v0p0p1_3.x65.X a_57123_n13359# GND.t1362 GND.t92 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X422 GND.t658 R0.t6 a_57123_n85079# GND.t112 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X423 VV11.t3 VV10.t3 GND.t77 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X424 OUT3.t44 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND.t305 GND.t304 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X425 VDD.t140 I1.t7 a_77605_n52567# VDD.t139 sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X426 VV15.t3 VV14.t2 GND.t51 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X427 GND.t463 16to4_PriorityEncoder_v0p0p1_0.x22.A 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND.t462 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X428 OUT2.t109 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD.t1020 VDD.t1019 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X429 frontAnalog_v0p0p1_7.RSfetsym_0.x2.Y frontAnalog_v0p0p1_7.x65.X VDD.t1201 VDD.t1196 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X430 OUT0.t113 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD.t898 VDD.t897 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X431 GND.t1500 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t49 GND.t1499 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X432 frontAnalog_v0p0p1_7.RSfetsym_0.x1.Y frontAnalog_v0p0p1_7.x63.X GND.t582 GND.t577 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X433 VDD.t1018 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t108 VDD.t1017 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X434 16to4_PriorityEncoder_v0p0p1_0.x29.Y 16to4_PriorityEncoder_v0p0p1_0.x29.A GND.t555 GND.t554 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X435 OUT0.t48 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND.t956 GND.t955 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X436 16to4_PriorityEncoder_v0p0p1_0.x29.Y 16to4_PriorityEncoder_v0p0p1_0.x29.A VDD.t537 VDD.t536 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X437 GND.t758 frontAnalog_v0p0p1_1.x63.A.t6 a_57123_n41879# GND.t662 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X438 frontAnalog_v0p0p1_11.RSfetsym_0.QN.t3 frontAnalog_v0p0p1_11.x65.X VDD.t727 VDD.t723 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.25
X439 VDD.t460 I6.t6 a_77637_n50057# VDD.t459 sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X440 a_16719_n13117.t19 a_16599_n13205.t8 a_16541_n13117.t4 GND.t722 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X441 frontAnalog_v0p0p1_2.RSfetsym_0.x2.Y frontAnalog_v0p0p1_2.x65.X VDD.t1231 VDD.t1224 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X442 a_77723_n40777# VDD.t1506 a_77637_n40777# GND.t695 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X443 OUT0.t47 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND.t954 GND.t953 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X444 16to4_PriorityEncoder_v0p0p1_0.x3.EI 16to4_PriorityEncoder_v0p0p1_0.x5.EO VDD.t652 VDD.t651 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X445 frontAnalog_v0p0p1_8.RSfetsym_0.x1.Y frontAnalog_v0p0p1_8.x63.X VDD.t764 VDD.t759 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X446 GND.t303 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t43 GND.t302 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X447 GND.t952 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t46 GND.t951 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X448 GND.t1557 16to4_PriorityEncoder_v0p0p1_0.x36.A 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND.t1556 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X449 VDD.t449 16to4_PriorityEncoder_v0p0p1_0.x22.A 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD.t448 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X450 GND.t1177 I13.t8 a_77723_n41087# GND.t1176 sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X451 VIN.t10 w_55000_n19128# error sky130_fd_pr__cap_var_lvt w=2 l=0.18
X452 R0.t0 S0.t5 VDD.t98 VDD.t97 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X453 VDD.t36 frontAnalog_v0p0p1_0.x65.X frontAnalog_v0p0p1_0.RSfetsym_0.QN.t1 VDD.t29 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.25
X454 16to4_PriorityEncoder_v0p0p1_0.x3.x16.X a_77605_n51585# VDD.t1210 VDD.t1209 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.312 ps=1.68 w=1 l=0.15
X455 VDD.t1014 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t107 VDD.t1013 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X456 VDD.t638 16to4_PriorityEncoder_v0p0p1_0.x43.A 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD.t637 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X457 a_53630_n57996# frontAnalog_v0p0p1_10.IB.t8 GND.t1248 GND.t36 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X458 R1.t0 CLK.t16 w_55000_n79150# VDD.t386 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X459 OUT1.t116 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD.t1442 VDD.t1441 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X460 OUT0.t112 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD.t896 VDD.t895 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X461 VV6.t15 VV5.t13 GND.t77 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X462 GND.t950 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t45 GND.t949 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X463 VDD.t535 16to4_PriorityEncoder_v0p0p1_0.x29.A 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD.t534 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X464 GND.t1205 frontAnalog_v0p0p1_13.x65.X frontAnalog_v0p0p1_13.RSfetsym_0.x2.Y GND.t1204 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X465 16to4_PriorityEncoder_v0p0p1_0.x3.x19.D I6.t7 GND.t475 GND.t474 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X466 frontAnalog_v0p0p1_4.x65.A.t0 CLK.t17 frontAnalog_v0p0p1_4.x63.A.t2 VDD.t387 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X467 a_59578_n73170# frontAnalog_v0p0p1_12.x65.X frontAnalog_v0p0p1_12.RSfetsym_0.QN.t0 GND.t197 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.315 ps=2.72 w=1 l=0.15
X468 OUT0.t111 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD.t894 VDD.t893 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X469 VV16.t5 VV15.t8 GND.t33 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X470 a_77605_n52567# 16to4_PriorityEncoder_v0p0p1_0.x3.x19.C VDD.t610 VDD.t139 sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.109 ps=1.36 w=0.42 l=0.15
X471 GND.t301 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t42 GND.t300 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X472 VV14.t12 VV13.t14 GND.t77 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X473 frontAnalog_v0p0p1_1.x63.A.t1 frontAnalog_v0p0p1_1.x65.A.t5 VDD.t160 VDD.t159 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X474 VDD.t892 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t110 VDD.t891 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X475 OUT1.t48 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND.t1498 GND.t1497 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X476 OUT3.t41 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND.t299 GND.t298 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X477 frontAnalog_v0p0p1_8.x65.X a_57123_n45759# VDD.t1300 VDD.t1299 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X478 a_53630_n14796# frontAnalog_v0p0p1_10.IB.t9 GND.t1249 GND.t36 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X479 frontAnalog_v0p0p1_7.x63.A.t0 CLK.t18 w_55000_n35950# VDD.t179 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X480 16to4_PriorityEncoder_v0p0p1_0.x36.Y 16to4_PriorityEncoder_v0p0p1_0.x36.A VDD.t1489 VDD.t1488 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X481 GND.t1307 frontAnalog_v0p0p1_4.x65.A.t5 a_57123_n18759# GND.t807 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X482 frontAnalog_v0p0p1_10.RSfetsym_0.QN.t0 frontAnalog_v0p0p1_10.RSfetsym_0.x1.Y GND.t32 GND.t31 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.25
X483 GND.t17 16to4_PriorityEncoder_v0p0p1_0.x3.x17.A a_78065_n49349# GND.t16 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X484 GND.t361 frontAnalog_v0p0p1_2.x63.A.t6 a_57123_n4079# GND.t360 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X485 frontAnalog_v0p0p1_0.RSfetsym_0.x2.Y frontAnalog_v0p0p1_0.x65.X VDD.t35 VDD.t31 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X486 OUT3.t113 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD.t304 VDD.t303 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X487 GND.t1377 frontAnalog_v0p0p1_5.x65.X frontAnalog_v0p0p1_5.RSfetsym_0.x2.Y GND.t1376 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X488 GND.t357 frontAnalog_v0p0p1_14.x63.X frontAnalog_v0p0p1_14.RSfetsym_0.x1.Y GND.t353 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X489 VDD.t1440 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t115 VDD.t1439 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X490 VDD.t15 frontAnalog_v0p0p1_12.x63.A.t4 a_57123_n74279# VDD.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X491 I12.t3 frontAnalog_v0p0p1_4.RSfetsym_0.QN.t5 VDD.t681 VDD.t680 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.3
X492 GND.t461 16to4_PriorityEncoder_v0p0p1_0.x22.A 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND.t460 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X493 VDD.t122 frontAnalog_v0p0p1_4.x63.X frontAnalog_v0p0p1_4.RSfetsym_0.x1.Y VDD.t119 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X494 VDD.t890 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t109 VDD.t889 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X495 VDD.t388 CLK.t19 w_55000_n57550# GND.t399 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X496 VDD.t763 frontAnalog_v0p0p1_8.x63.X I7.t3 VDD.t757 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.25
X497 VDD.t1216 frontAnalog_v0p0p1_11.x63.A.t4 frontAnalog_v0p0p1_11.x65.A.t3 VDD.t668 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X498 w_55000_n46128# CLK.t20 frontAnalog_v0p0p1_8.x65.A.t0 VDD.t203 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X499 16to4_PriorityEncoder_v0p0p1_0.x43.Y 16to4_PriorityEncoder_v0p0p1_0.x43.A GND.t643 GND.t642 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X500 I14.t3 frontAnalog_v0p0p1_0.RSfetsym_0.x2.Y GND.t783 GND.t782 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.25
X501 OUT1.t47 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND.t1496 GND.t1495 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X502 VDD.t717 I15.t5 a_77639_n42341# VDD.t716 sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X503 VV13.t16 w_55000_n19750# error sky130_fd_pr__cap_var_lvt w=2 l=0.18
X504 a_16719_n13117.t18 a_16599_n13205.t9 a_16541_n13117.t3 GND.t723 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X505 frontAnalog_v0p0p1_13.x65.A.t1 frontAnalog_v0p0p1_13.x63.A.t5 a_55268_n68736# GND.t605 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X506 OUT2.t106 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD.t1012 VDD.t1011 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X507 GND.t1494 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t46 GND.t1493 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X508 OUT3.t112 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD.t302 VDD.t301 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X509 frontAnalog_v0p0p1_3.RSfetsym_0.QN.t4 frontAnalog_v0p0p1_3.RSfetsym_0.x1.Y GND.t1211 GND.t782 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.25
X510 VDD.t1438 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t114 VDD.t1437 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X511 GND.t581 frontAnalog_v0p0p1_7.x63.X frontAnalog_v0p0p1_7.RSfetsym_0.x1.Y GND.t577 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X512 VDD.t44 frontAnalog_v0p0p1_2.x63.X I15.t2 VDD.t37 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.25
X513 VDD.t775 frontAnalog_v0p0p1_6.x63.A.t4 a_57123_n31079# VDD.t774 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X514 VDD.t1487 16to4_PriorityEncoder_v0p0p1_0.x36.A 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD.t1486 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X515 a_53630_n74196# VV3.t16 w_55000_n73128# GND.t1170 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X516 VV5.t15 VV4.t15 GND.t52 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X517 VDD.t636 16to4_PriorityEncoder_v0p0p1_0.x43.A 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD.t635 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X518 VV12.t12 VV11.t13 GND.t122 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X519 GND.t948 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t44 GND.t947 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X520 VDD.t447 16to4_PriorityEncoder_v0p0p1_0.x22.A 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD.t446 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X521 OUT3.t40 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND.t297 GND.t296 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X522 VDD.t1208 16to4_PriorityEncoder_v0p0p1_0.x3.x19.D a_77605_n52567# VDD.t139 sky130_fd_pr__pfet_01v8_hvt ad=0.312 pd=1.68 as=0.0588 ps=0.7 w=0.42 l=0.15
X523 a_55268_n52536# CLK.t21 GND.t401 GND.t400 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X524 16to4_PriorityEncoder_v0p0p1_0.x22.Y 16to4_PriorityEncoder_v0p0p1_0.x22.A GND.t459 GND.t458 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X525 frontAnalog_v0p0p1_5.x65.A.t2 frontAnalog_v0p0p1_5.x63.A.t5 a_55268_n25536# GND.t419 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X526 GND.t641 16to4_PriorityEncoder_v0p0p1_0.x43.A 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND.t640 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X527 GND.t1088 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t50 GND.t1087 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X528 VDD.t762 frontAnalog_v0p0p1_8.x63.X frontAnalog_v0p0p1_8.RSfetsym_0.x1.Y VDD.t759 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X529 OUT3.t111 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD.t300 VDD.t299 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X530 VDD.t1436 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t113 VDD.t1435 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X531 GND.t800 frontAnalog_v0p0p1_7.RSfetsym_0.QN.t6 a_59577_n35883# GND.t799 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X532 a_53630_n30996# VV11.t16 w_55000_n29928# GND.t408 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X533 16to4_PriorityEncoder_v0p0p1_0.x36.Y 16to4_PriorityEncoder_v0p0p1_0.x36.A GND.t1555 GND.t1554 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X534 VDD.t298 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t110 VDD.t297 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X535 OUT1.t112 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD.t1434 VDD.t1433 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X536 VDD.t888 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t108 VDD.t887 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X537 a_55268_n9336# CLK.t22 GND.t403 GND.t402 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X538 GND.t767 frontAnalog_v0p0p1_11.x65.X frontAnalog_v0p0p1_11.RSfetsym_0.x2.Y GND.t766 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X539 VIN.t11 w_55000_n83928# error sky130_fd_pr__cap_var_lvt w=2 l=0.18
X540 frontAnalog_v0p0p1_5.RSfetsym_0.x1.Y frontAnalog_v0p0p1_5.x63.X VDD.t26 VDD.t19 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X541 VDD.t1064 I7.t5 a_77639_n50381# VDD.t1063 sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X542 16to4_PriorityEncoder_v0p0p1_0.x22.Y 16to4_PriorityEncoder_v0p0p1_0.x22.A VDD.t445 VDD.t444 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X543 VDD.t356 frontAnalog_v0p0p1_2.x63.A.t7 frontAnalog_v0p0p1_2.x65.A.t3 VDD.t355 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X544 VDD.t188 frontAnalog_v0p0p1_12.x65.X frontAnalog_v0p0p1_12.RSfetsym_0.QN.t2 VDD.t183 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.25
X545 16to4_PriorityEncoder_v0p0p1_0.x5.x21.B a_77605_n44527# GND.t118 GND.t117 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.196 ps=1.33 w=0.65 l=0.15
X546 OUT1.t45 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND.t1492 GND.t1491 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X547 16to4_PriorityEncoder_v0p0p1_0.x29.Y 16to4_PriorityEncoder_v0p0p1_0.x29.A VDD.t533 VDD.t532 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X548 frontAnalog_v0p0p1_2.x65.A.t1 CLK.t23 frontAnalog_v0p0p1_2.x63.A.t2 VDD.t417 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X549 VV11.t1 VV10.t1 GND.t51 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X550 VDD.t296 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t109 VDD.t295 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X551 OUT2.t105 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD.t1010 VDD.t1009 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X552 GND.t1490 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t44 GND.t1489 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X553 VV16.t14 VV15.t13 GND.t78 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X554 S0.t2 CLK.t24 R0.t2 VDD.t418 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X555 frontAnalog_v0p0p1_9.x63.X a_57123_n52679# VDD.t1183 VDD.t1182 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X556 OUT0.t43 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND.t946 GND.t945 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X557 w_55000_n68350# VIN.t12 a_53630_n68796# GND.t712 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X558 OUT2.t49 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND.t1086 GND.t1085 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X559 GND.t141 I10.t6 a_77605_n39305# GND.t140 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X560 GND.t132 frontAnalog_v0p0p1_12.x63.X frontAnalog_v0p0p1_12.RSfetsym_0.x1.Y GND.t129 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X561 VIN.t13 w_55000_n40728# error sky130_fd_pr__cap_var_lvt w=2 l=0.18
X562 VDD.t34 frontAnalog_v0p0p1_0.x65.X frontAnalog_v0p0p1_0.RSfetsym_0.x2.Y VDD.t31 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X563 VDD.t138 16to4_PriorityEncoder_v0p0p1_0.x5.x4.A a_78313_n39305# VDD.t137 sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X564 VDD.t1223 I12.t5 a_77855_n40069# VDD.t1222 sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X565 VV1.t1 VL.t1 GND.t24 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X566 GND.t113 S0.t6 a_57123_n83559# GND.t112 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X567 16to4_PriorityEncoder_v0p0p1_0.x3.x18.C I2.t6 GND.t345 GND.t344 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X568 a_77723_n49127# 16to4_PriorityEncoder_v0p0p1_0.x3.EI a_77637_n49127# GND.t1302 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X569 VDD.t294 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t108 VDD.t293 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X570 GND.t553 16to4_PriorityEncoder_v0p0p1_0.x29.A 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND.t552 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X571 R0.t1 S0.t7 a_55268_n84936# GND.t114 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X572 16to4_PriorityEncoder_v0p0p1_0.x3.A2 a_78065_n49349# VDD.t46 VDD.t45 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.148 ps=1.34 w=1 l=0.15
X573 I0.t0 frontAnalog_v0p0p1_15.RSfetsym_0.QN.t5 VDD.t108 VDD.t107 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.3
X574 VV9.t10 VV8.t10 GND.t24 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X575 frontAnalog_v0p0p1_1.x65.A.t0 CLK.t25 frontAnalog_v0p0p1_1.x63.A.t3 VDD.t419 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X576 frontAnalog_v0p0p1_11.RSfetsym_0.x2.Y frontAnalog_v0p0p1_11.x65.X VDD.t726 VDD.t720 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X577 VDD.t486 frontAnalog_v0p0p1_15.x63.X frontAnalog_v0p0p1_15.RSfetsym_0.x1.Y VDD.t480 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X578 GND.t1488 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t43 GND.t1487 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X579 OUT3.t107 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD.t292 VDD.t291 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X580 frontAnalog_v0p0p1_2.RSfetsym_0.x1.Y frontAnalog_v0p0p1_2.x63.X VDD.t43 VDD.t39 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X581 w_55000_n25150# VIN.t14 a_53630_n25596# GND.t606 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X582 GND.t615 frontAnalog_v0p0p1_6.x63.X frontAnalog_v0p0p1_6.RSfetsym_0.x1.Y GND.t612 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X583 OUT0.t42 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND.t944 GND.t943 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X584 frontAnalog_v0p0p1_8.RSfetsym_0.x2.Y frontAnalog_v0p0p1_8.x65.X GND.t1399 GND.t1398 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X585 OUT0.t107 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD.t886 VDD.t885 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X586 a_78065_n49349# 16to4_PriorityEncoder_v0p0p1_0.x3.x22.A GND.t1533 GND.t1532 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X587 frontAnalog_v0p0p1_11.x63.X a_57123_n63479# GND.t505 GND.t504 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X588 a_53630_n3996# VV16.t16 w_55000_n2928# GND.t1169 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X589 GND.t942 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t41 GND.t941 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X590 I3.t0 frontAnalog_v0p0p1_13.RSfetsym_0.x2.Y GND.t188 GND.t187 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.25
X591 VV1.t17 w_55000_n84550# error sky130_fd_pr__cap_var_lvt w=2 l=0.18
X592 a_78065_n41309# 16to4_PriorityEncoder_v0p0p1_0.x5.x11.X GND.t1569 GND.t1568 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X593 OUT1.t111 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD.t1432 VDD.t1431 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X594 GND.t663 frontAnalog_v0p0p1_1.x65.A.t6 a_57123_n40359# GND.t662 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X595 16to4_PriorityEncoder_v0p0p1_0.x3.x21.B a_77605_n52567# GND.t169 GND.t168 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.196 ps=1.33 w=0.65 l=0.15
X596 OUT3.t39 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND.t295 GND.t294 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X597 OUT2.t48 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND.t1084 GND.t1083 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X598 a_82988_n43855# 16to4_PriorityEncoder_v0p0p1_0.x3.A2 a_82906_n43855# VDD.t1255 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X599 GND.t1082 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t47 GND.t1081 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X600 16to4_PriorityEncoder_v0p0p1_0.x28.A 16to4_PriorityEncoder_v0p0p1_0.x1.X VDD.t664 VDD.t663 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X601 frontAnalog_v0p0p1_1.x63.A.t0 frontAnalog_v0p0p1_1.x65.A.t7 a_55268_n41736# GND.t664 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X602 GND.t1486 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t42 GND.t1485 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X603 VV6.t2 VV5.t2 GND.t51 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X604 I8.t3 frontAnalog_v0p0p1_1.RSfetsym_0.QN.t5 VDD.t601 VDD.t4 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.3
X605 GND.t293 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t38 GND.t292 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X606 VDD.t174 frontAnalog_v0p0p1_1.x63.X frontAnalog_v0p0p1_1.RSfetsym_0.x1.Y VDD.t168 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X607 GND.t1080 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t46 GND.t1079 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X608 VDD.t1127 frontAnalog_v0p0p1_14.x65.X frontAnalog_v0p0p1_14.RSfetsym_0.x2.Y VDD.t1123 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X609 OUT3.t106 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD.t290 VDD.t289 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X610 16to4_PriorityEncoder_v0p0p1_0.x29.Y 16to4_PriorityEncoder_v0p0p1_0.x29.A GND.t551 GND.t550 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X611 frontAnalog_v0p0p1_10.RSfetsym_0.x1.Y frontAnalog_v0p0p1_10.x63.X GND.t846 GND.t842 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X612 a_59577_n46683# frontAnalog_v0p0p1_8.x63.X I7.t1 GND.t813 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X613 VV14.t1 VV13.t0 GND.t51 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X614 a_59578_n56970# frontAnalog_v0p0p1_10.x65.X frontAnalog_v0p0p1_10.RSfetsym_0.QN.t1 GND.t99 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.315 ps=2.72 w=1 l=0.15
X615 VV5.t6 VV4.t5 GND.t202 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X616 GND.t855 I2.t7 a_77605_n47345# GND.t154 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X617 16to4_PriorityEncoder_v0p0p1_0.x3.x4.A 16to4_PriorityEncoder_v0p0p1_0.x3.EI VDD.t1242 VDD.t1241 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X618 OUT0.t106 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD.t884 VDD.t883 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X619 VDD.t100 16to4_PriorityEncoder_v0p0p1_0.x3.x4.A a_78313_n47345# VDD.t99 sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X620 VDD.t288 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t105 VDD.t287 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X621 I11.t4 frontAnalog_v0p0p1_5.RSfetsym_0.x2.Y GND.t852 GND.t851 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.25
X622 VV9.t17 w_55000_n41350# error sky130_fd_pr__cap_var_lvt w=2 l=0.18
X623 GND.t1137 frontAnalog_v0p0p1_14.RSfetsym_0.QN.t6 a_59577_n79083# GND.t1136 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X624 GND.t176 16to4_PriorityEncoder_v0p0p1_0.x5.x15.X a_78349_n43045# GND.t175 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X625 VDD.t882 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t105 VDD.t881 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X626 16to4_PriorityEncoder_v0p0p1_0.x3.x21.B a_77605_n52567# VDD.t156 VDD.t155 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.312 ps=1.68 w=1 l=0.15
X627 GND.t291 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t37 GND.t290 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X628 VDD.t1200 frontAnalog_v0p0p1_7.x65.X frontAnalog_v0p0p1_7.RSfetsym_0.x2.Y VDD.t1196 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X629 frontAnalog_v0p0p1_13.RSfetsym_0.x1.Y frontAnalog_v0p0p1_13.x63.X VDD.t379 VDD.t372 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X630 a_77775_n43295# 16to4_PriorityEncoder_v0p0p1_0.x5.x19.C a_77687_n43295# GND.t703 sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
X631 OUT2.t45 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND.t1078 GND.t1077 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X632 GND.t1076 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t44 GND.t1075 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X633 frontAnalog_v0p0p1_3.RSfetsym_0.x1.Y frontAnalog_v0p0p1_3.x63.X GND.t486 GND.t482 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X634 OUT1.t41 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND.t1484 GND.t1483 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X635 VDD.t634 16to4_PriorityEncoder_v0p0p1_0.x43.A 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD.t633 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X636 a_59578_n13770# frontAnalog_v0p0p1_3.x65.X frontAnalog_v0p0p1_3.RSfetsym_0.QN.t3 GND.t570 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.315 ps=2.72 w=1 l=0.15
X637 a_53630_n52596# frontAnalog_v0p0p1_10.IB.t10 GND.t1250 GND.t36 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X638 I8.t2 frontAnalog_v0p0p1_1.x63.X VDD.t173 VDD.t170 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.25
X639 16to4_PriorityEncoder_v0p0p1_0.x1.X a_82906_n47995# GND.t1369 GND.t1368 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1 ps=0.985 w=0.65 l=0.15
X640 16to4_PriorityEncoder_v0p0p1_0.x5.x17.A a_77637_n42017# VDD.t346 VDD.t345 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.167 ps=1.39 w=1 l=0.15
X641 VFS.t6 VV16.t11 GND.t709 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X642 VDD.t597 frontAnalog_v0p0p1_8.x63.A.t4 frontAnalog_v0p0p1_8.x65.A.t2 VDD.t596 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X643 GND.t1310 I7.t6 a_59578_n46170# GND.t1309 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X644 16to4_PriorityEncoder_v0p0p1_0.x3.EI 16to4_PriorityEncoder_v0p0p1_0.x5.EO GND.t667 GND.t666 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X645 OUT0.t40 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND.t940 GND.t939 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X646 frontAnalog_v0p0p1_2.RSfetsym_0.QN.t0 frontAnalog_v0p0p1_2.RSfetsym_0.x1.Y GND.t72 GND.t71 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.25
X647 VV4.t12 VV3.t12 GND.t33 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X648 VDD.t1230 frontAnalog_v0p0p1_2.x65.X frontAnalog_v0p0p1_2.RSfetsym_0.x2.Y VDD.t1224 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X649 GND.t362 frontAnalog_v0p0p1_2.x65.A.t5 a_57123_n2559# GND.t360 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X650 frontAnalog_v0p0p1_15.RSfetsym_0.QN.t4 I0.t6 VDD.t1068 VDD.t107 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.3
X651 VV8.t14 VV7.t15 GND.t52 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X652 GND.t289 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t36 GND.t288 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X653 frontAnalog_v0p0p1_11.x65.X a_57123_n61959# GND.t760 GND.t504 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X654 GND.t938 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t39 GND.t937 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X655 OUT1.t40 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND.t1482 GND.t1481 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X656 a_77605_n43295# 16to4_PriorityEncoder_v0p0p1_0.x5.x16.C VDD.t767 VDD.t766 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X657 VDD.t106 frontAnalog_v0p0p1_3.x63.A.t5 a_57123_n14879# VDD.t105 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X658 OUT3.t35 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND.t287 GND.t286 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X659 VDD.t286 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t104 VDD.t285 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X660 GND.t1180 I12.t6 a_77605_n40069# GND.t90 sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X661 frontAnalog_v0p0p1_4.RSfetsym_0.QN.t4 I12.t7 VDD.t1094 VDD.t680 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.3
X662 VDD.t1220 frontAnalog_v0p0p1_12.x65.A.t4 a_57123_n72759# VDD.t1219 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X663 GND.t1312 frontAnalog_v0p0p1_13.x63.A.t6 a_57123_n68879# GND.t848 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X664 VDD.t1008 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t104 VDD.t1007 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X665 16to4_PriorityEncoder_v0p0p1_0.x43.Y 16to4_PriorityEncoder_v0p0p1_0.x43.A VDD.t632 VDD.t631 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X666 VDD.t1430 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t110 VDD.t1429 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X667 VDD.t725 frontAnalog_v0p0p1_11.x65.X frontAnalog_v0p0p1_11.RSfetsym_0.x2.Y VDD.t720 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X668 VDD.t42 frontAnalog_v0p0p1_2.x63.X frontAnalog_v0p0p1_2.RSfetsym_0.x1.Y VDD.t39 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X669 GND.t457 16to4_PriorityEncoder_v0p0p1_0.x22.A 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND.t456 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X670 frontAnalog_v0p0p1_1.RSfetsym_0.QN.t4 I8.t5 VDD.t5 VDD.t4 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.3
X671 OUT0.t104 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD.t880 VDD.t879 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X672 a_77605_n39305# I11.t5 GND.t148 GND.t140 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X673 GND.t936 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t38 GND.t935 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X674 frontAnalog_v0p0p1_4.RSfetsym_0.x2.Y frontAnalog_v0p0p1_4.x65.X VDD.t479 VDD.t474 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X675 VDD.t878 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t103 VDD.t877 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X676 OUT1.t39 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND.t1480 GND.t1479 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X677 frontAnalog_v0p0p1_4.RSfetsym_0.x1.Y frontAnalog_v0p0p1_4.x63.X GND.t139 GND.t134 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X678 OUT3.t34 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND.t285 GND.t284 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X679 a_77855_n40069# I13.t9 a_77783_n40069# VDD.t1093 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X680 VV2.t3 VV1.t2 GND.t106 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X681 OUT2.t43 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND.t1074 GND.t1073 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X682 VDD.t284 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t103 VDD.t283 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X683 a_16719_n13117.t17 a_16599_n13205.t10 a_16541_n13117.t2 GND.t724 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X684 GND.t1478 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t38 GND.t1477 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X685 GND.t421 frontAnalog_v0p0p1_5.x63.A.t6 a_57123_n25679# GND.t420 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X686 frontAnalog_v0p0p1_8.RSfetsym_0.QN.t4 frontAnalog_v0p0p1_8.x65.X VDD.t1335 VDD.t1331 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.25
X687 frontAnalog_v0p0p1_1.RSfetsym_0.x1.Y frontAnalog_v0p0p1_1.x63.X GND.t181 GND.t177 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X688 OUT3.t102 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD.t282 VDD.t281 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X689 GND.t660 I14.t5 a_77723_n42017# GND.t659 sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X690 frontAnalog_v0p0p1_2.x63.A.t0 frontAnalog_v0p0p1_2.x65.A.t6 a_55268_n3936# GND.t363 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X691 GND.t934 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t37 GND.t933 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X692 VDD.t443 16to4_PriorityEncoder_v0p0p1_0.x22.A 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD.t442 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X693 VDD.t502 I8.t6 a_77855_n39305# VDD.t501 sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X694 OUT3.t33 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND.t283 GND.t282 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X695 16to4_PriorityEncoder_v0p0p1_0.x22.Y 16to4_PriorityEncoder_v0p0p1_0.x22.A GND.t455 GND.t454 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X696 VDD.t1006 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t103 VDD.t1005 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X697 VDD.t876 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t102 VDD.t875 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X698 a_77605_n51335# 16to4_PriorityEncoder_v0p0p1_0.x3.x16.C VDD.t337 VDD.t336 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X699 frontAnalog_v0p0p1_13.x63.A.t2 frontAnalog_v0p0p1_13.x65.A.t5 VDD.t587 VDD.t570 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X700 a_77881_n52819# 16to4_PriorityEncoder_v0p0p1_0.x3.x19.C a_77775_n52819# GND.t185 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X701 frontAnalog_v0p0p1_2.RSfetsym_0.QN.t4 frontAnalog_v0p0p1_2.x65.X VDD.t1229 VDD.t1227 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.25
X702 GND.t639 16to4_PriorityEncoder_v0p0p1_0.x43.A 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND.t638 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X703 frontAnalog_v0p0p1_9.RSfetsym_0.x1.Y frontAnalog_v0p0p1_9.x63.X VDD.t1102 VDD.t1097 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X704 GND.t1476 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t37 GND.t1475 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X705 GND.t21 I4.t7 a_77605_n48109# GND.t20 sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X706 OUT2.t102 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD.t1004 VDD.t1003 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X707 OUT3.t101 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD.t280 VDD.t279 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X708 VDD.t1428 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t109 VDD.t1427 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X709 OUT1.t108 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD.t1426 VDD.t1425 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X710 VDD.t542 frontAnalog_v0p0p1_3.x65.X frontAnalog_v0p0p1_3.RSfetsym_0.QN.t1 VDD.t541 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.25
X711 VDD.t874 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t101 VDD.t873 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X712 I0.t3 frontAnalog_v0p0p1_15.x63.X VDD.t485 VDD.t482 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.25
X713 a_77605_n47345# I3.t5 GND.t1195 GND.t154 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X714 OUT3.t32 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND.t281 GND.t280 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X715 frontAnalog_v0p0p1_5.x63.A.t0 frontAnalog_v0p0p1_5.x65.A.t5 VDD.t94 VDD.t93 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X716 OUT0.t36 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND.t932 GND.t931 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X717 a_59577_n3483# frontAnalog_v0p0p1_2.x63.X I15.t0 GND.t56 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X718 VV12.t13 VV11.t14 GND.t59 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X719 16to4_PriorityEncoder_v0p0p1_0.x2.X a_82906_n51645# GND.t1226 GND.t1225 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1 ps=0.985 w=0.65 l=0.15
X720 16to4_PriorityEncoder_v0p0p1_0.x22.Y 16to4_PriorityEncoder_v0p0p1_0.x22.A VDD.t441 VDD.t440 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X721 w_55000_n2928# CLK.t26 frontAnalog_v0p0p1_2.x65.A.t0 VDD.t420 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X722 frontAnalog_v0p0p1_6.x65.X a_57123_n29559# VDD.t1106 VDD.t1105 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X723 GND.t279 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t31 GND.t278 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X724 frontAnalog_v0p0p1_4.x63.A.t3 CLK.t27 w_55000_n19750# VDD.t421 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X725 VDD.t1002 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t101 VDD.t1001 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X726 OUT2.t100 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD.t1000 VDD.t999 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X727 16to4_PriorityEncoder_v0p0p1_0.x29.Y 16to4_PriorityEncoder_v0p0p1_0.x29.A GND.t549 GND.t548 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X728 GND.t477 I6.t8 a_77723_n50057# GND.t476 sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X729 frontAnalog_v0p0p1_9.x65.X a_57123_n51159# VDD.t1188 VDD.t1187 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X730 VV4.t9 VV3.t9 GND.t78 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X731 frontAnalog_v0p0p1_8.x63.X a_57123_n47279# GND.t1381 GND.t1364 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X732 VDD.t566 frontAnalog_v0p0p1_10.x63.A.t5 a_57123_n58079# VDD.t565 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X733 OUT1.t107 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD.t1424 VDD.t1423 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X734 VV10.t0 VV9.t0 GND.t106 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X735 VDD.t422 CLK.t28 w_55000_n62328# GND.t399 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X736 OUT0.t35 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND.t930 GND.t929 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X737 frontAnalog_v0p0p1_11.RSfetsym_0.QN.t1 frontAnalog_v0p0p1_11.RSfetsym_0.x1.Y GND.t718 GND.t170 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.25
X738 16to4_PriorityEncoder_v0p0p1_0.x5.x16.C I13.t10 GND.t1179 GND.t1178 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X739 a_78349_n51085# 16to4_PriorityEncoder_v0p0p1_0.x3.x16.X GND.t215 GND.t14 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X740 VDD.t1070 I0.t7 a_77855_n47345# VDD.t1069 sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X741 VV3.t2 VV2.t1 GND.t122 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X742 a_77687_n43545# I11.t6 a_77605_n43545# GND.t699 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.109 ps=1.36 w=0.42 l=0.15
X743 VV13.t1 VV12.t0 GND.t106 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X744 a_53630_n9396# frontAnalog_v0p0p1_10.IB.t11 GND.t1251 GND.t384 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X745 frontAnalog_v0p0p1_12.RSfetsym_0.x2.Y frontAnalog_v0p0p1_12.x65.X GND.t196 GND.t195 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X746 VDD.t748 I11.t7 a_77605_n44779# VDD.t747 sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X747 VV8.t2 VV7.t4 GND.t202 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X748 OUT2.t99 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD.t998 VDD.t997 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X749 VDD.t25 frontAnalog_v0p0p1_5.x63.X frontAnalog_v0p0p1_5.RSfetsym_0.x1.Y VDD.t19 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X750 VV2.t5 VV1.t3 GND.t77 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X751 OUT0.t100 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD.t872 VDD.t871 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X752 VDD.t1325 16to4_PriorityEncoder_v0p0p1_0.x5.x17.A a_78599_n43045# VDD.t1324 sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X753 VDD.t1101 frontAnalog_v0p0p1_9.x63.X I6.t2 VDD.t1100 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.25
X754 VDD.t423 CLK.t29 w_55000_n62950# GND.t435 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X755 GND.t277 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t30 GND.t276 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X756 16to4_PriorityEncoder_v0p0p1_0.x2.X a_82906_n51645# VDD.t1135 VDD.t1134 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.146 ps=1.34 w=1 l=0.15
X757 w_55000_n51528# CLK.t30 frontAnalog_v0p0p1_9.x65.A.t3 VDD.t556 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X758 OUT1.t36 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND.t1474 GND.t1473 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X759 VDD.t1485 16to4_PriorityEncoder_v0p0p1_0.x36.A 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD.t1484 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X760 GND.t138 frontAnalog_v0p0p1_4.x63.X frontAnalog_v0p0p1_4.RSfetsym_0.x1.Y GND.t134 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X761 16to4_PriorityEncoder_v0p0p1_0.x3.x19.C I4.t8 GND.t23 GND.t22 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X762 frontAnalog_v0p0p1_12.x65.A.t0 frontAnalog_v0p0p1_12.x63.A.t5 a_55268_n74136# GND.t13 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X763 a_53630_n57996# VV6.t16 w_55000_n56928# GND.t1282 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X764 GND.t547 16to4_PriorityEncoder_v0p0p1_0.x29.A 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND.t546 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X765 VDD.t531 16to4_PriorityEncoder_v0p0p1_0.x29.A 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD.t530 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X766 OUT0.t34 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND.t928 GND.t927 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X767 frontAnalog_v0p0p1_15.RSfetsym_0.x2.Y frontAnalog_v0p0p1_15.x65.X VDD.t198 VDD.t192 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X768 OUT0.t99 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD.t870 VDD.t869 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X769 GND.t180 frontAnalog_v0p0p1_1.x63.X frontAnalog_v0p0p1_1.RSfetsym_0.x1.Y GND.t177 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X770 frontAnalog_v0p0p1_0.x63.X a_57123_n9479# VDD.t684 VDD.t683 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X771 frontAnalog_v0p0p1_6.RSfetsym_0.x2.Y frontAnalog_v0p0p1_6.x65.X GND.t10 GND.t9 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X772 a_55268_n36336# CLK.t31 GND.t586 GND.t585 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X773 frontAnalog_v0p0p1_15.RSfetsym_0.x1.Y frontAnalog_v0p0p1_15.x63.X GND.t501 GND.t497 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X774 GND.t637 16to4_PriorityEncoder_v0p0p1_0.x43.A 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND.t636 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X775 GND.t926 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t33 GND.t925 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X776 VDD.t557 CLK.t32 w_55000_n19750# GND.t587 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X777 VFS.t0 VV16.t3 GND.t432 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X778 OUT1.t106 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD.t1422 VDD.t1421 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X779 OUT3.t29 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND.t275 GND.t274 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X780 VDD.t996 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t98 VDD.t995 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X781 GND.t513 frontAnalog_v0p0p1_0.RSfetsym_0.QN.t5 a_59577_n8883# GND.t512 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X782 OUT1.t105 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD.t1420 VDD.t1419 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X783 a_53630_n14796# VV14.t16 w_55000_n13728# GND.t740 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X784 GND.t711 frontAnalog_v0p0p1_4.RSfetsym_0.QN.t6 a_59577_n19683# GND.t710 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X785 GND.t143 I10.t7 a_59578_n29970# GND.t142 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X786 16to4_PriorityEncoder_v0p0p1_0.x36.Y 16to4_PriorityEncoder_v0p0p1_0.x36.A VDD.t1483 VDD.t1482 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X787 OUT3.t100 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD.t278 VDD.t277 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X788 VDD.t1099 frontAnalog_v0p0p1_9.x63.X frontAnalog_v0p0p1_9.RSfetsym_0.x1.Y VDD.t1097 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X789 VDD.t1418 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t104 VDD.t1417 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X790 frontAnalog_v0p0p1_1.RSfetsym_0.x2.Y frontAnalog_v0p0p1_1.x65.X VDD.t711 VDD.t704 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X791 frontAnalog_v0p0p1_14.x63.X a_57123_n79679# VDD.t1267 VDD.t1266 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X792 a_77687_n51585# I3.t6 a_77605_n51585# GND.t174 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.109 ps=1.36 w=0.42 l=0.15
X793 OUT0.t98 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD.t868 VDD.t867 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X794 a_78735_n39527# 16to4_PriorityEncoder_v0p0p1_0.x5.EO a_78649_n39527# GND.t665 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X795 GND.t1397 frontAnalog_v0p0p1_8.x65.X frontAnalog_v0p0p1_8.RSfetsym_0.x2.Y GND.t1396 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X796 16to4_PriorityEncoder_v0p0p1_0.x5.x11.X a_77637_n41087# VDD.t53 VDD.t52 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.167 ps=1.39 w=1 l=0.15
X797 VDD.t276 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t99 VDD.t275 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X798 VIN.t15 w_55000_n67728# error sky130_fd_pr__cap_var_lvt w=2 l=0.18
X799 GND.t700 VDD.t1507 a_77881_n43545# GND.t699 sky130_fd_pr__nfet_01v8 ad=0.196 pd=1.33 as=0.0693 ps=0.75 w=0.42 l=0.15
X800 GND.t924 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t32 GND.t923 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X801 VDD.t164 I3.t7 a_77605_n52819# VDD.t163 sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X802 a_77605_n44779# VDD.t1171 VDD.t1172 VDD.t731 sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.109 ps=1.36 w=0.42 l=0.15
X803 VDD.t18 16to4_PriorityEncoder_v0p0p1_0.x3.x17.A a_78599_n51085# VDD.t17 sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X804 GND.t84 16to4_PriorityEncoder_v0p0p1_0.x35.A 16to4_PriorityEncoder_v0p0p1_0.x36.A GND.t83 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X805 VDD.t866 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t97 VDD.t865 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X806 VDD.t82 frontAnalog_v0p0p1_10.x65.X frontAnalog_v0p0p1_10.RSfetsym_0.QN.t2 VDD.t81 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.25
X807 OUT3.t28 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND.t273 GND.t272 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X808 a_77855_n39305# I9.t7 a_77783_n39305# VDD.t777 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X809 a_78097_n45737# VDD.t1168 VDD.t1170 VDD.t1169 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X810 VDD.t398 16to4_PriorityEncoder_v0p0p1_0.x42.A 16to4_PriorityEncoder_v0p0p1_0.x43.A VDD.t397 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X811 VDD.t1416 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t103 VDD.t1415 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X812 GND.t271 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t27 GND.t270 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X813 VV10.t11 VV9.t9 GND.t77 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X814 OUT2.t42 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND.t1072 GND.t1071 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X815 frontAnalog_v0p0p1_13.x65.A.t2 CLK.t33 frontAnalog_v0p0p1_13.x63.A.t0 VDD.t558 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X816 OUT1.t35 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND.t1472 GND.t1471 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X817 frontAnalog_v0p0p1_7.x63.X a_57123_n36479# VDD.t361 VDD.t360 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X818 GND.t845 frontAnalog_v0p0p1_10.x63.X frontAnalog_v0p0p1_10.RSfetsym_0.x1.Y GND.t842 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X819 VIN.t16 w_55000_n24528# error sky130_fd_pr__cap_var_lvt w=2 l=0.18
X820 VV13.t9 VV12.t9 GND.t77 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X821 a_53630_n3996# frontAnalog_v0p0p1_10.IB.t12 GND.t1252 GND.t384 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X822 16to4_PriorityEncoder_v0p0p1_0.x22.Y 16to4_PriorityEncoder_v0p0p1_0.x22.A GND.t453 GND.t452 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X823 a_53630_n63396# frontAnalog_v0p0p1_10.IB.t13 GND.t37 GND.t36 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X824 VDD.t864 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t96 VDD.t863 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X825 R0.t3 CLK.t34 w_55000_n84550# VDD.t559 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X826 GND.t849 frontAnalog_v0p0p1_13.x65.A.t6 a_57123_n67359# GND.t848 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X827 OUT2.t97 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD.t994 VDD.t993 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X828 frontAnalog_v0p0p1_13.x63.A.t3 frontAnalog_v0p0p1_13.x65.A.t7 a_55268_n68736# GND.t850 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X829 GND.t194 frontAnalog_v0p0p1_12.x65.X frontAnalog_v0p0p1_12.RSfetsym_0.x2.Y GND.t193 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X830 16to4_PriorityEncoder_v0p0p1_0.x36.A 16to4_PriorityEncoder_v0p0p1_0.x35.A VDD.t67 VDD.t66 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X831 VDD.t529 16to4_PriorityEncoder_v0p0p1_0.x29.A 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD.t528 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X832 frontAnalog_v0p0p1_5.x65.A.t1 CLK.t35 frontAnalog_v0p0p1_5.x63.A.t3 VDD.t560 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X833 I3.t4 frontAnalog_v0p0p1_13.RSfetsym_0.QN.t5 VDD.t1072 VDD.t165 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.3
X834 VDD.t378 frontAnalog_v0p0p1_13.x63.X frontAnalog_v0p0p1_13.RSfetsym_0.x1.Y VDD.t372 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X835 frontAnalog_v0p0p1_8.RSfetsym_0.x2.Y frontAnalog_v0p0p1_8.x65.X VDD.t1334 VDD.t1329 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X836 16to4_PriorityEncoder_v0p0p1_0.x5.x15.X a_77605_n43295# GND.t150 GND.t149 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.196 ps=1.33 w=0.65 l=0.15
X837 GND.t485 frontAnalog_v0p0p1_3.x63.X frontAnalog_v0p0p1_3.RSfetsym_0.x1.Y GND.t482 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X838 GND.t1181 I12.t8 a_77723_n40777# GND.t1176 sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X839 a_78735_n47567# 16to4_PriorityEncoder_v0p0p1_0.x3.EO a_78649_n47567# GND.t109 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X840 GND.t1303 16to4_PriorityEncoder_v0p0p1_0.x3.EI a_77881_n51585# GND.t174 sky130_fd_pr__nfet_01v8 ad=0.196 pd=1.33 as=0.0693 ps=0.75 w=0.42 l=0.15
X841 a_77605_n52819# 16to4_PriorityEncoder_v0p0p1_0.x3.EI VDD.t1240 VDD.t700 sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.109 ps=1.36 w=0.42 l=0.15
X842 VV5.t14 VV4.t14 GND.t24 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X843 16to4_PriorityEncoder_v0p0p1_0.x43.Y 16to4_PriorityEncoder_v0p0p1_0.x43.A VDD.t630 VDD.t629 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X844 VV4.t17 w_55000_n68350# error sky130_fd_pr__cap_var_lvt w=2 l=0.18
X845 OUT0.t31 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND.t922 GND.t921 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X846 VDD.t662 16to4_PriorityEncoder_v0p0p1_0.x5.x19.D a_77605_n44779# VDD.t661 sky130_fd_pr__pfet_01v8_hvt ad=0.312 pd=1.68 as=0.0588 ps=0.7 w=0.42 l=0.15
X847 GND.t433 frontAnalog_v0p0p1_5.x65.A.t6 a_57123_n24159# GND.t420 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X848 frontAnalog_v0p0p1_9.RSfetsym_0.x2.Y frontAnalog_v0p0p1_9.x65.X GND.t1333 GND.t1332 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X849 16to4_PriorityEncoder_v0p0p1_0.x22.Y 16to4_PriorityEncoder_v0p0p1_0.x22.A VDD.t439 VDD.t438 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X850 frontAnalog_v0p0p1_5.x63.A.t1 frontAnalog_v0p0p1_5.x65.A.t7 a_55268_n25536# GND.t434 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X851 a_78097_n53777# 16to4_PriorityEncoder_v0p0p1_0.x3.EI VDD.t1239 VDD.t1238 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X852 GND.t451 16to4_PriorityEncoder_v0p0p1_0.x22.A 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND.t450 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X853 a_77855_n47345# I1.t8 a_77783_n47345# VDD.t141 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X854 GND.t8 frontAnalog_v0p0p1_6.x65.X frontAnalog_v0p0p1_6.RSfetsym_0.x2.Y GND.t7 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X855 GND.t500 frontAnalog_v0p0p1_15.x63.X frontAnalog_v0p0p1_15.RSfetsym_0.x1.Y GND.t497 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X856 I11.t3 frontAnalog_v0p0p1_5.RSfetsym_0.QN.t5 VDD.t734 VDD.t733 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.3
X857 VDD.t1414 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t102 VDD.t1413 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X858 a_78599_n43045# 16to4_PriorityEncoder_v0p0p1_0.x5.x22.A a_78527_n43045# VDD.t409 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X859 OUT2.t41 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND.t1070 GND.t1069 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X860 VDD.t274 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t98 VDD.t273 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X861 16to4_PriorityEncoder_v0p0p1_0.x29.Y 16to4_PriorityEncoder_v0p0p1_0.x29.A VDD.t527 VDD.t526 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X862 16to4_PriorityEncoder_v0p0p1_0.x5.x15.X a_77605_n43295# VDD.t136 VDD.t135 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.312 ps=1.68 w=1 l=0.15
X863 I3.t3 frontAnalog_v0p0p1_13.x63.X VDD.t377 VDD.t374 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.25
X864 a_53630_n79596# frontAnalog_v0p0p1_10.IB.t14 GND.t38 GND.t36 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X865 VV15.t1 VV14.t0 GND.t33 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X866 OUT3.t97 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD.t272 VDD.t271 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X867 VV12.t17 w_55000_n25150# error sky130_fd_pr__cap_var_lvt w=2 l=0.18
X868 frontAnalog_v0p0p1_11.RSfetsym_0.x1.Y frontAnalog_v0p0p1_11.x63.X GND.t510 GND.t506 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X869 OUT0.t95 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD.t862 VDD.t861 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X870 I10.t4 frontAnalog_v0p0p1_6.RSfetsym_0.x2.Y GND.t1390 GND.t583 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.25
X871 GND.t125 frontAnalog_v0p0p1_15.RSfetsym_0.QN.t6 a_59577_n84483# GND.t124 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X872 VDD.t437 16to4_PriorityEncoder_v0p0p1_0.x22.A 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD.t436 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X873 VDD.t1481 16to4_PriorityEncoder_v0p0p1_0.x36.A 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD.t1480 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X874 VDD.t478 frontAnalog_v0p0p1_4.x65.X frontAnalog_v0p0p1_4.RSfetsym_0.x2.Y VDD.t474 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X875 16to4_PriorityEncoder_v0p0p1_0.x3.x14.A a_77637_n48817# GND.t1323 GND.t1322 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.112 ps=1.04 w=0.65 l=0.15
X876 OUT2.t40 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND.t1068 GND.t1067 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X877 VDD.t778 I9.t8 a_77605_n44527# VDD.t659 sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X878 I11.t2 frontAnalog_v0p0p1_5.x63.X VDD.t24 VDD.t21 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.25
X879 a_53630_n36396# frontAnalog_v0p0p1_10.IB.t15 GND.t39 GND.t36 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X880 16to4_PriorityEncoder_v0p0p1_0.x3.x2.X a_77605_n48109# GND.t796 GND.t795 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.102 ps=0.99 w=0.65 l=0.15
X881 frontAnalog_v0p0p1_12.RSfetsym_0.x1.Y frontAnalog_v0p0p1_12.x63.X VDD.t116 VDD.t109 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X882 VDD.t776 frontAnalog_v0p0p1_6.x63.A.t5 frontAnalog_v0p0p1_6.x65.A.t3 VDD.t144 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X883 OUT3.t96 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD.t270 VDD.t269 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X884 a_16541_n13117.t0 GND.t393 GND.t392 sky130_fd_pr__res_xhigh_po_5p73 l=85.8
X885 VV2.t6 VV1.t4 GND.t51 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X886 VDD.t1207 16to4_PriorityEncoder_v0p0p1_0.x3.x19.D a_77605_n52819# VDD.t1206 sky130_fd_pr__pfet_01v8_hvt ad=0.312 pd=1.68 as=0.0588 ps=0.7 w=0.42 l=0.15
X887 GND.t425 16to4_PriorityEncoder_v0p0p1_0.x5.x22.A a_78525_n45515# GND.t424 sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X888 frontAnalog_v0p0p1_13.RSfetsym_0.QN.t0 I3.t8 VDD.t166 VDD.t165 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.3
X889 GND.t479 I6.t9 a_59578_n51570# GND.t478 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X890 frontAnalog_v0p0p1_8.x65.X a_57123_n45759# GND.t1365 GND.t1364 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X891 GND.t618 frontAnalog_v0p0p1_1.RSfetsym_0.QN.t6 a_59577_n41283# GND.t617 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X892 OUT0.t30 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND.t920 GND.t919 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X893 16to4_PriorityEncoder_v0p0p1_0.x36.Y 16to4_PriorityEncoder_v0p0p1_0.x36.A GND.t1553 GND.t1552 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X894 a_78599_n51085# 16to4_PriorityEncoder_v0p0p1_0.x3.x22.A a_78527_n51085# VDD.t1467 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X895 OUT1.t101 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD.t1412 VDD.t1411 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X896 w_55000_n3550# VIN.t17 a_53630_n3996# GND.t1169 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X897 16to4_PriorityEncoder_v0p0p1_0.x3.x15.X a_77605_n51335# VDD.t697 VDD.t696 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.312 ps=1.68 w=1 l=0.15
X898 16to4_PriorityEncoder_v0p0p1_0.x43.Y 16to4_PriorityEncoder_v0p0p1_0.x43.A VDD.t628 VDD.t627 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X899 frontAnalog_v0p0p1_6.RSfetsym_0.x1.Y frontAnalog_v0p0p1_6.x63.X VDD.t595 VDD.t588 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X900 VDD.t679 frontAnalog_v0p0p1_10.x65.A.t4 a_57123_n56559# VDD.t678 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X901 VDD.t1117 16to4_PriorityEncoder_v0p0p1_0.x3.x14.A a_78315_n49349# VDD.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X902 frontAnalog_v0p0p1_0.RSfetsym_0.x1.Y frontAnalog_v0p0p1_0.x63.X VDD.t369 VDD.t362 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X903 frontAnalog_v0p0p1_3.RSfetsym_0.x2.Y frontAnalog_v0p0p1_3.x65.X GND.t569 GND.t568 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X904 frontAnalog_v0p0p1_13.RSfetsym_0.x1.Y frontAnalog_v0p0p1_13.x63.X GND.t381 GND.t379 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X905 VV7.t7 VV6.t8 GND.t52 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X906 GND.t1470 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t34 GND.t1469 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X907 VDD.t1333 frontAnalog_v0p0p1_8.x65.X frontAnalog_v0p0p1_8.RSfetsym_0.x2.Y VDD.t1329 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X908 GND.t1144 16to4_PriorityEncoder_v0p0p1_0.x5.x2.X a_78159_n39549# GND.t1143 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X909 frontAnalog_v0p0p1_5.RSfetsym_0.QN.t0 I11.t8 VDD.t749 VDD.t733 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.3
X910 VV1.t10 VL.t6 GND.t106 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X911 GND.t798 frontAnalog_v0p0p1_12.x63.A.t6 a_57123_n74279# GND.t797 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X912 OUT2.t39 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND.t1066 GND.t1065 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X913 VDD.t268 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t95 VDD.t267 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X914 16to4_PriorityEncoder_v0p0p1_0.x5.x19.D I14.t6 GND.t147 GND.t146 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X915 OUT0.t94 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD.t860 VDD.t859 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X916 OUT1.t100 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD.t1410 VDD.t1409 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X917 w_55000_n73750# VIN.t18 a_53630_n74196# GND.t1170 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X918 VV9.t6 VV8.t7 GND.t106 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X919 a_77605_n44527# 16to4_PriorityEncoder_v0p0p1_0.x5.x19.C VDD.t743 VDD.t659 sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.109 ps=1.36 w=0.42 l=0.15
X920 OUT2.t38 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND.t1064 GND.t1063 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X921 GND.t1062 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t37 GND.t1061 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X922 GND.t1551 16to4_PriorityEncoder_v0p0p1_0.x36.A 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND.t1550 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X923 frontAnalog_v0p0p1_14.RSfetsym_0.x1.Y frontAnalog_v0p0p1_14.x63.X VDD.t351 VDD.t347 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X924 OUT3.t94 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD.t266 VDD.t265 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X925 VDD.t675 frontAnalog_v0p0p1_3.x65.A.t4 a_57123_n13359# VDD.t674 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X926 frontAnalog_v0p0p1_5.RSfetsym_0.x2.Y frontAnalog_v0p0p1_5.x65.X VDD.t1312 VDD.t1306 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X927 VDD.t1408 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t99 VDD.t1407 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X928 frontAnalog_v0p0p1_5.RSfetsym_0.x1.Y frontAnalog_v0p0p1_5.x63.X GND.t28 GND.t26 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X929 frontAnalog_v0p0p1_6.RSfetsym_0.QN.t2 frontAnalog_v0p0p1_6.x65.X VDD.t11 VDD.t6 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.25
X930 VDD.t264 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t93 VDD.t263 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X931 VDD.t626 16to4_PriorityEncoder_v0p0p1_0.x43.A 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD.t625 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X932 GND.t1531 16to4_PriorityEncoder_v0p0p1_0.x3.x22.A a_78525_n53555# GND.t1530 sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X933 frontAnalog_v0p0p1_0.x65.X a_57123_n7959# VDD.t1140 VDD.t1139 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X934 GND.t1186 frontAnalog_v0p0p1_6.x63.A.t6 a_57123_n31079# GND.t430 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X935 frontAnalog_v0p0p1_9.RSfetsym_0.QN.t4 frontAnalog_v0p0p1_9.x65.X VDD.t1273 VDD.t1268 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.25
X936 VDD.t710 frontAnalog_v0p0p1_1.x65.X frontAnalog_v0p0p1_1.RSfetsym_0.QN.t3 VDD.t707 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.25
X937 16to4_PriorityEncoder_v0p0p1_0.x5.GS a_78649_n39527# GND.t35 GND.t34 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.112 ps=1.04 w=0.65 l=0.15
X938 GND.t1468 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t33 GND.t1467 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X939 VV10.t5 VV9.t5 GND.t51 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X940 frontAnalog_v0p0p1_7.RSfetsym_0.x1.Y frontAnalog_v0p0p1_7.x63.X VDD.t552 VDD.t548 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X941 VV15.t11 VV14.t13 GND.t78 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X942 VV3.t0 VV2.t0 GND.t59 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X943 OUT3.t92 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD.t262 VDD.t261 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X944 OUT1.t32 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND.t1466 GND.t1465 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X945 VDD.t992 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t96 VDD.t991 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X946 VV13.t8 VV12.t6 GND.t51 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X947 frontAnalog_v0p0p1_12.x63.A.t2 frontAnalog_v0p0p1_12.x65.A.t5 VDD.t1221 VDD.t670 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X948 I2.t3 frontAnalog_v0p0p1_12.RSfetsym_0.x2.Y GND.t201 GND.t200 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.25
X949 GND.t1060 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t36 GND.t1059 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X950 a_77605_n39305# I9.t9 GND.t827 GND.t140 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X951 frontAnalog_v0p0p1_14.x65.X a_57123_n78159# VDD.t1262 VDD.t1261 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X952 GND.t204 16to4_PriorityEncoder_v0p0p1_0.x3.x2.X a_78159_n47589# GND.t203 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X953 16to4_PriorityEncoder_v0p0p1_0.x3.x16.C I5.t9 VDD.t703 VDD.t702 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X954 16to4_PriorityEncoder_v0p0p1_0.x36.Y 16to4_PriorityEncoder_v0p0p1_0.x36.A VDD.t1479 VDD.t1478 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X955 a_77723_n48817# 16to4_PriorityEncoder_v0p0p1_0.x3.EI a_77637_n48817# GND.t1302 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X956 frontAnalog_v0p0p1_13.x63.A.t1 CLK.t36 w_55000_n68350# VDD.t561 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X957 a_82988_n51645# 16to4_PriorityEncoder_v0p0p1_0.x3.A0 a_82906_n51645# VDD.t154 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X958 VDD.t197 frontAnalog_v0p0p1_15.x65.X frontAnalog_v0p0p1_15.RSfetsym_0.x2.Y VDD.t192 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X959 GND.t1058 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t35 GND.t1057 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X960 GND.t1133 I5.t10 a_77723_n49127# GND.t0 sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X961 16to4_PriorityEncoder_v0p0p1_0.x5.GS a_78649_n39527# VDD.t28 VDD.t27 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.167 ps=1.39 w=1 l=0.15
X962 a_59578_n62370# frontAnalog_v0p0p1_11.x65.X frontAnalog_v0p0p1_11.RSfetsym_0.QN.t4 GND.t765 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.315 ps=2.72 w=1 l=0.15
X963 a_59577_n52083# frontAnalog_v0p0p1_9.x63.X I6.t1 GND.t1191 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X964 VV8.t11 VV7.t13 GND.t24 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X965 VDD.t350 frontAnalog_v0p0p1_14.x63.X I1.t1 VDD.t349 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.25
X966 16to4_PriorityEncoder_v0p0p1_0.x43.Y 16to4_PriorityEncoder_v0p0p1_0.x43.A GND.t635 GND.t634 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X967 frontAnalog_v0p0p1_6.x63.A.t0 frontAnalog_v0p0p1_6.x65.A.t4 VDD.t77 VDD.t76 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X968 GND.t1464 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t31 GND.t1463 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X969 OUT1.t30 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND.t1462 GND.t1461 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X970 VDD.t660 16to4_PriorityEncoder_v0p0p1_0.x5.x19.D a_77605_n44527# VDD.t659 sky130_fd_pr__pfet_01v8_hvt ad=0.312 pd=1.68 as=0.0588 ps=0.7 w=0.42 l=0.15
X971 VDD.t260 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t91 VDD.t259 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X972 w_55000_n78528# CLK.t37 S1.t0 VDD.t581 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X973 OUT1.t98 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD.t1406 VDD.t1405 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X974 16to4_PriorityEncoder_v0p0p1_0.x5.A2 a_78065_n41309# GND.t429 GND.t428 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.102 ps=0.99 w=0.65 l=0.15
X975 frontAnalog_v0p0p1_7.x65.X a_57123_n34959# VDD.t1260 VDD.t1259 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X976 frontAnalog_v0p0p1_5.x63.A.t2 CLK.t38 w_55000_n25150# VDD.t405 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X977 VV1.t0 VL.t0 GND.t77 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X978 VDD.t1184 CLK.t39 w_55000_n46128# GND.t1161 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X979 VDD.t1404 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t97 VDD.t1403 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X980 frontAnalog_v0p0p1_8.RSfetsym_0.QN.t0 frontAnalog_v0p0p1_8.RSfetsym_0.x1.Y GND.t527 GND.t526 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.25
X981 VDD.t709 frontAnalog_v0p0p1_1.x65.X frontAnalog_v0p0p1_1.RSfetsym_0.x2.Y VDD.t704 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X982 16to4_PriorityEncoder_v0p0p1_0.x3.GS a_78649_n47567# GND.t657 GND.t656 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.112 ps=1.04 w=0.65 l=0.15
X983 OUT2.t95 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD.t990 VDD.t989 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X984 GND.t567 frontAnalog_v0p0p1_3.x65.X frontAnalog_v0p0p1_3.RSfetsym_0.x2.Y GND.t566 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X985 GND.t269 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t26 GND.t268 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X986 frontAnalog_v0p0p1_10.RSfetsym_0.x2.Y frontAnalog_v0p0p1_10.x65.X GND.t98 GND.t97 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X987 GND.t380 frontAnalog_v0p0p1_13.x63.X frontAnalog_v0p0p1_13.RSfetsym_0.x1.Y GND.t379 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X988 VDD.t1218 frontAnalog_v0p0p1_11.x63.A.t5 a_57123_n63479# VDD.t1217 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X989 VV9.t15 VV8.t15 GND.t77 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X990 VV11.t6 VV10.t6 GND.t33 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X991 OUT1.t29 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND.t1460 GND.t1459 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X992 VDD.t1185 CLK.t40 w_55000_n46750# GND.t837 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X993 frontAnalog_v0p0p1_2.RSfetsym_0.x1.Y frontAnalog_v0p0p1_2.x63.X GND.t55 GND.t53 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X994 VDD.t551 frontAnalog_v0p0p1_7.x63.X I9.t0 VDD.t550 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.25
X995 a_77775_n52819# I3.t9 a_77687_n52819# GND.t185 sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
X996 OUT3.t25 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND.t267 GND.t266 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X997 w_55000_n35328# CLK.t41 frontAnalog_v0p0p1_7.x65.A.t2 VDD.t1186 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X998 GND.t918 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t29 GND.t917 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X999 VDD.t342 frontAnalog_v0p0p1_9.x63.A.t4 frontAnalog_v0p0p1_9.x65.A.t1 VDD.t145 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1000 VDD.t258 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t90 VDD.t257 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1001 frontAnalog_v0p0p1_2.RSfetsym_0.x2.Y frontAnalog_v0p0p1_2.x65.X GND.t1292 GND.t1291 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1002 16to4_PriorityEncoder_v0p0p1_0.x36.A 16to4_PriorityEncoder_v0p0p1_0.x35.A GND.t82 GND.t81 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1003 a_55268_n84936# CLK.t42 GND.t1256 GND.t1255 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1004 GND.t545 16to4_PriorityEncoder_v0p0p1_0.x29.A 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND.t544 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1005 VDD.t525 16to4_PriorityEncoder_v0p0p1_0.x29.A 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD.t524 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1006 a_77605_n47345# I1.t9 GND.t155 GND.t154 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1007 frontAnalog_v0p0p1_10.x65.A.t3 frontAnalog_v0p0p1_10.x63.A.t6 a_55268_n57936# GND.t590 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1008 OUT3.t89 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD.t256 VDD.t255 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1009 VDD.t1402 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t96 VDD.t1401 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1010 VDD.t348 frontAnalog_v0p0p1_14.x63.X frontAnalog_v0p0p1_14.RSfetsym_0.x1.Y VDD.t347 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1011 VV7.t8 VV6.t10 GND.t202 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1012 frontAnalog_v0p0p1_13.RSfetsym_0.x2.Y frontAnalog_v0p0p1_13.x65.X VDD.t1115 VDD.t1109 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1013 GND.t27 frontAnalog_v0p0p1_5.x63.X frontAnalog_v0p0p1_5.RSfetsym_0.x1.Y GND.t26 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1014 a_78315_n49349# 16to4_PriorityEncoder_v0p0p1_0.x3.x11.X a_78243_n49349# VDD.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X1015 VDD.t1119 frontAnalog_v0p0p1_4.x63.A.t6 a_57123_n20279# VDD.t1118 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1016 a_53630_n63396# VV5.t16 w_55000_n62328# GND.t671 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1017 16to4_PriorityEncoder_v0p0p1_0.x3.GS a_78649_n47567# VDD.t646 VDD.t645 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.167 ps=1.39 w=1 l=0.15
X1018 OUT3.t24 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND.t265 GND.t264 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1019 GND.t1056 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t34 GND.t1055 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1020 a_55268_n41736# CLK.t43 GND.t1258 GND.t1257 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1021 VIN.t19 w_55000_n2928# error sky130_fd_pr__cap_var_lvt w=2 l=0.18
X1022 OUT2.t94 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD.t988 VDD.t987 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1023 VDD.t858 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t93 VDD.t857 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1024 GND.t1458 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t28 GND.t1457 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1025 VDD.t986 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t93 VDD.t985 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1026 16to4_PriorityEncoder_v0p0p1_0.x43.Y 16to4_PriorityEncoder_v0p0p1_0.x43.A VDD.t624 VDD.t623 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1027 frontAnalog_v0p0p1_3.x65.A.t2 frontAnalog_v0p0p1_3.x63.A.t6 a_55268_n14736# GND.t119 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1028 VDD.t1400 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t95 VDD.t1399 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1029 VDD.t549 frontAnalog_v0p0p1_7.x63.X frontAnalog_v0p0p1_7.RSfetsym_0.x1.Y VDD.t548 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1030 16to4_PriorityEncoder_v0p0p1_0.x29.Y 16to4_PriorityEncoder_v0p0p1_0.x29.A GND.t543 GND.t542 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1031 VDD.t984 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t92 VDD.t983 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1032 16to4_PriorityEncoder_v0p0p1_0.x5.x18.C I10.t8 GND.t145 GND.t144 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1033 16to4_PriorityEncoder_v0p0p1_0.x29.Y 16to4_PriorityEncoder_v0p0p1_0.x29.A VDD.t523 VDD.t522 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1034 GND.t916 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t28 GND.t915 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1035 VV6.t9 VV5.t9 GND.t33 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1036 OUT3.t23 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND.t263 GND.t262 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1037 OUT0.t27 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND.t914 GND.t913 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1038 frontAnalog_v0p0p1_0.RSfetsym_0.x2.Y frontAnalog_v0p0p1_0.x65.X GND.t45 GND.t44 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1039 GND.t1331 frontAnalog_v0p0p1_9.x65.X frontAnalog_v0p0p1_9.RSfetsym_0.x2.Y GND.t1330 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1040 GND.t261 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t22 GND.t260 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1041 VIN.t20 w_55000_n73128# error sky130_fd_pr__cap_var_lvt w=2 l=0.18
X1042 VV14.t11 VV13.t12 GND.t33 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1043 OUT3.t88 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD.t254 VDD.t253 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1044 VDD.t724 frontAnalog_v0p0p1_11.x65.X frontAnalog_v0p0p1_11.RSfetsym_0.QN.t2 VDD.t723 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.25
X1045 VDD.t982 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t91 VDD.t981 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1046 OUT2.t90 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD.t980 VDD.t979 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1047 VDD.t622 16to4_PriorityEncoder_v0p0p1_0.x43.A 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD.t621 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1048 OUT1.t94 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD.t1398 VDD.t1397 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1049 16to4_PriorityEncoder_v0p0p1_0.x1.X a_82906_n47995# VDD.t1305 VDD.t1304 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.146 ps=1.34 w=1 l=0.15
X1050 a_16599_n13205.t3 a_16599_n13205.t2 GND.t728 GND.t727 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1051 VDD.t856 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t92 VDD.t855 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1052 frontAnalog_v0p0p1_12.x65.A.t2 CLK.t44 frontAnalog_v0p0p1_12.x63.A.t0 VDD.t572 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1053 GND.t912 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t26 GND.t911 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1054 OUT0.t25 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND.t910 GND.t909 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1055 frontAnalog_v0p0p1_1.x63.X a_57123_n41879# VDD.t339 VDD.t338 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1056 a_53630_n47196# frontAnalog_v0p0p1_10.IB.t16 GND.t40 GND.t36 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1057 w_55000_n57550# VIN.t21 a_53630_n57996# GND.t777 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1058 GND.t509 frontAnalog_v0p0p1_11.x63.X frontAnalog_v0p0p1_11.RSfetsym_0.x1.Y GND.t506 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1059 OUT0.t91 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD.t854 VDD.t853 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1060 16to4_PriorityEncoder_v0p0p1_0.x5.x4.A VDD.t1165 VDD.t1167 VDD.t1166 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1061 frontAnalog_v0p0p1_14.RSfetsym_0.x2.Y frontAnalog_v0p0p1_14.x65.X GND.t1221 GND.t1220 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1062 frontAnalog_v0p0p1_0.x63.A.t3 frontAnalog_v0p0p1_0.x65.A.t4 VDD.t149 VDD.t148 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1063 GND.t96 frontAnalog_v0p0p1_10.x65.X frontAnalog_v0p0p1_10.RSfetsym_0.x2.Y GND.t95 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1064 OUT1.t27 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND.t1456 GND.t1455 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1065 VV16.t17 w_55000_n3550# error sky130_fd_pr__cap_var_lvt w=2 l=0.18
X1066 16to4_PriorityEncoder_v0p0p1_0.x29.A 16to4_PriorityEncoder_v0p0p1_0.x28.A GND.t1157 GND.t1156 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1067 OUT1.t93 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD.t1396 VDD.t1395 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1068 GND.t54 frontAnalog_v0p0p1_2.x63.X frontAnalog_v0p0p1_2.RSfetsym_0.x1.Y GND.t53 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1069 GND.t1280 frontAnalog_v0p0p1_12.x65.A.t6 a_57123_n72759# GND.t797 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X1070 16to4_PriorityEncoder_v0p0p1_0.x5.x21.B a_77605_n44527# VDD.t102 VDD.t101 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.312 ps=1.68 w=1 l=0.15
X1071 OUT0.t24 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND.t908 GND.t907 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1072 a_16719_n13117.t16 a_16599_n13205.t11 a_16541_n13117.t20 GND.t725 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1073 VV11.t4 VV10.t4 GND.t78 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1074 frontAnalog_v0p0p1_6.x65.A.t1 CLK.t45 frontAnalog_v0p0p1_6.x63.A.t2 VDD.t573 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1075 I2.t4 frontAnalog_v0p0p1_12.RSfetsym_0.QN.t5 VDD.t1263 VDD.t793 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.3
X1076 VDD.t115 frontAnalog_v0p0p1_12.x63.X frontAnalog_v0p0p1_12.RSfetsym_0.x1.Y VDD.t109 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1077 frontAnalog_v0p0p1_9.RSfetsym_0.x2.Y frontAnalog_v0p0p1_9.x65.X VDD.t1272 VDD.t1270 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1078 w_55000_n14350# VIN.t22 a_53630_n14796# GND.t740 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1079 frontAnalog_v0p0p1_7.RSfetsym_0.x2.Y frontAnalog_v0p0p1_7.x65.X GND.t1268 GND.t1267 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1080 GND.t449 16to4_PriorityEncoder_v0p0p1_0.x22.A 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND.t448 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1081 VDD.t852 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t90 VDD.t851 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1082 OUT0.t89 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD.t850 VDD.t849 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1083 VDD.t1 I4.t9 a_77855_n48109# VDD.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X1084 VDD.t742 16to4_PriorityEncoder_v0p0p1_0.x5.x19.C a_77605_n43545# VDD.t741 sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X1085 frontAnalog_v0p0p1_9.x63.X a_57123_n52679# GND.t1254 GND.t1253 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1086 16to4_PriorityEncoder_v0p0p1_0.x43.Y 16to4_PriorityEncoder_v0p0p1_0.x43.A GND.t633 GND.t632 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1087 I5.t0 frontAnalog_v0p0p1_10.RSfetsym_0.x2.Y GND.t171 GND.t170 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.25
X1088 VV3.t17 w_55000_n73750# error sky130_fd_pr__cap_var_lvt w=2 l=0.18
X1089 OUT1.t92 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD.t1394 VDD.t1393 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1090 frontAnalog_v0p0p1_6.x63.A.t1 frontAnalog_v0p0p1_6.x65.A.t5 a_55268_n30936# GND.t94 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1091 OUT2.t89 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD.t978 VDD.t977 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1092 a_77687_n51335# I2.t8 a_77605_n51335# GND.t346 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.109 ps=1.36 w=0.42 l=0.15
X1093 VDD.t1392 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t91 VDD.t1391 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1094 I10.t0 frontAnalog_v0p0p1_6.RSfetsym_0.QN.t5 VDD.t503 VDD.t125 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.3
X1095 VDD.t594 frontAnalog_v0p0p1_6.x63.X frontAnalog_v0p0p1_6.RSfetsym_0.x1.Y VDD.t588 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1096 a_59578_n2970# frontAnalog_v0p0p1_2.x65.X frontAnalog_v0p0p1_2.RSfetsym_0.QN.t2 GND.t1290 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.315 ps=2.72 w=1 l=0.15
X1097 OUT0.t88 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD.t848 VDD.t847 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1098 VDD.t368 frontAnalog_v0p0p1_0.x63.X frontAnalog_v0p0p1_0.RSfetsym_0.x1.Y VDD.t362 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1099 frontAnalog_v0p0p1_8.RSfetsym_0.x1.Y frontAnalog_v0p0p1_8.x63.X GND.t812 GND.t809 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1100 GND.t906 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t23 GND.t905 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1101 a_78065_n49349# 16to4_PriorityEncoder_v0p0p1_0.x3.x11.X GND.t789 GND.t788 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1102 a_59577_n35883# frontAnalog_v0p0p1_7.x63.X I9.t2 GND.t580 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1103 a_53630_n84996# frontAnalog_v0p0p1_10.IB.t17 GND.t41 GND.t36 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1104 VDD.t435 16to4_PriorityEncoder_v0p0p1_0.x22.A 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD.t434 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1105 a_77637_n42017# VDD.t1162 VDD.t1164 VDD.t1163 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X1106 I13.t4 frontAnalog_v0p0p1_3.RSfetsym_0.x2.Y GND.t1346 GND.t654 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.25
X1107 VV11.t17 w_55000_n30550# error sky130_fd_pr__cap_var_lvt w=2 l=0.18
X1108 frontAnalog_v0p0p1_0.x63.A.t1 CLK.t46 w_55000_n8950# VDD.t574 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1109 GND.t1146 frontAnalog_v0p0p1_13.RSfetsym_0.QN.t6 a_59577_n68283# GND.t1145 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1110 16to4_PriorityEncoder_v0p0p1_0.x22.Y 16to4_PriorityEncoder_v0p0p1_0.x22.A GND.t447 GND.t446 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1111 GND.t1233 I1.t10 a_59578_n78570# GND.t1232 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1112 GND.t541 16to4_PriorityEncoder_v0p0p1_0.x29.A 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND.t540 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1113 I14.t2 frontAnalog_v0p0p1_0.x63.X VDD.t367 VDD.t365 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.25
X1114 VV1.t13 VL.t7 GND.t51 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1115 GND.t43 frontAnalog_v0p0p1_0.x65.X frontAnalog_v0p0p1_0.RSfetsym_0.x2.Y GND.t42 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1116 VDD.t575 CLK.t47 w_55000_n29928# GND.t595 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1117 a_16719_n13117.t15 a_16599_n13205.t12 a_16541_n13117.t19 GND.t726 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1118 OUT3.t87 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD.t252 VDD.t251 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1119 VDD.t1390 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t90 VDD.t1389 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1120 VDD.t1311 frontAnalog_v0p0p1_5.x65.X frontAnalog_v0p0p1_5.RSfetsym_0.x2.Y VDD.t1306 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1121 frontAnalog_v0p0p1_10.RSfetsym_0.x1.Y frontAnalog_v0p0p1_10.x63.X VDD.t788 VDD.t783 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1122 VV6.t6 VV5.t7 GND.t78 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1123 OUT2.t33 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND.t1054 GND.t1053 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1124 VDD.t250 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t86 VDD.t249 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1125 VV9.t8 VV8.t8 GND.t51 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1126 a_53630_n41796# frontAnalog_v0p0p1_10.IB.t18 GND.t1124 GND.t36 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1127 16to4_PriorityEncoder_v0p0p1_0.x3.x11.X a_77637_n49127# GND.t1337 GND.t1322 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.112 ps=1.04 w=0.65 l=0.15
X1128 I14.t4 frontAnalog_v0p0p1_0.RSfetsym_0.QN.t6 VDD.t498 VDD.t129 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.3
X1129 VDD.t609 16to4_PriorityEncoder_v0p0p1_0.x3.x19.C a_77605_n51585# VDD.t176 sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X1130 a_77605_n43545# I11.t9 VDD.t1136 VDD.t741 sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.109 ps=1.36 w=0.42 l=0.15
X1131 VV14.t10 VV13.t11 GND.t78 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1132 VDD.t846 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t87 VDD.t845 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1133 GND.t1052 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t32 GND.t1051 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1134 GND.t781 frontAnalog_v0p0p1_5.RSfetsym_0.QN.t6 a_59577_n25083# GND.t780 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1135 frontAnalog_v0p0p1_6.x65.X a_57123_n29559# GND.t1194 GND.t719 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1136 16to4_PriorityEncoder_v0p0p1_0.x3.x19.D I6.t10 VDD.t1257 VDD.t1256 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1137 GND.t829 I9.t10 a_59578_n35370# GND.t828 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1138 16to4_PriorityEncoder_v0p0p1_0.x5.x2.X a_77605_n40069# VDD.t390 VDD.t389 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.148 ps=1.34 w=1 l=0.15
X1139 a_77605_n52567# 16to4_PriorityEncoder_v0p0p1_0.x3.x18.C VDD.t461 VDD.t139 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X1140 16to4_PriorityEncoder_v0p0p1_0.x22.Y 16to4_PriorityEncoder_v0p0p1_0.x22.A VDD.t433 VDD.t432 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1141 frontAnalog_v0p0p1_15.x63.X a_57123_n85079# VDD.t1501 VDD.t1500 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1142 frontAnalog_v0p0p1_3.RSfetsym_0.x1.Y frontAnalog_v0p0p1_3.x63.X VDD.t471 VDD.t464 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1143 VDD.t248 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t85 VDD.t247 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1144 16to4_PriorityEncoder_v0p0p1_0.x29.Y 16to4_PriorityEncoder_v0p0p1_0.x29.A VDD.t521 VDD.t520 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1145 GND.t1301 16to4_PriorityEncoder_v0p0p1_0.x3.EI a_77881_n51335# GND.t346 sky130_fd_pr__nfet_01v8 ad=0.196 pd=1.33 as=0.0693 ps=0.75 w=0.42 l=0.15
X1146 16to4_PriorityEncoder_v0p0p1_0.x3.x17.A a_77637_n50057# VDD.t1251 VDD.t1250 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.167 ps=1.39 w=1 l=0.15
X1147 a_77881_n44779# 16to4_PriorityEncoder_v0p0p1_0.x5.x19.C a_77775_n44779# GND.t678 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X1148 16to4_PriorityEncoder_v0p0p1_0.x3.x20.X a_77605_n53805# GND.t1383 GND.t1382 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X1149 VV12.t10 VV11.t8 GND.t709 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1150 OUT0.t22 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND.t904 GND.t903 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1151 VDD.t1150 frontAnalog_v0p0p1_11.x65.A.t4 a_57123_n61959# VDD.t1149 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1152 16to4_PriorityEncoder_v0p0p1_0.x22.A 16to4_PriorityEncoder_v0p0p1_0.x21.A GND.t1353 GND.t1352 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1153 GND.t592 frontAnalog_v0p0p1_10.x63.A.t7 a_57123_n58079# GND.t591 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X1154 frontAnalog_v0p0p1_14.RSfetsym_0.QN.t4 frontAnalog_v0p0p1_14.x65.X VDD.t1126 VDD.t1121 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.25
X1155 VDD.t1271 frontAnalog_v0p0p1_9.x65.X frontAnalog_v0p0p1_9.RSfetsym_0.x2.Y VDD.t1270 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1156 a_77783_n40069# I14.t7 a_77687_n40069# VDD.t128 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X1157 VDD.t246 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t84 VDD.t245 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1158 VDD.t576 CLK.t48 w_55000_n8328# GND.t596 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1159 OUT1.t89 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD.t1388 VDD.t1387 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1160 VV5.t8 VV4.t7 GND.t106 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1161 GND.t1050 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t31 GND.t1049 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1162 OUT3.t83 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD.t244 VDD.t243 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1163 a_77605_n51585# I3.t10 VDD.t177 VDD.t176 sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.109 ps=1.36 w=0.42 l=0.15
X1164 VDD.t519 16to4_PriorityEncoder_v0p0p1_0.x29.A 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD.t518 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1165 GND.t121 frontAnalog_v0p0p1_3.x63.A.t7 a_57123_n14879# GND.t120 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X1166 VDD.t577 CLK.t49 w_55000_n8950# GND.t597 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1167 frontAnalog_v0p0p1_7.RSfetsym_0.QN.t4 frontAnalog_v0p0p1_7.x65.X VDD.t1199 VDD.t1194 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.25
X1168 frontAnalog_v0p0p1_12.x63.A.t3 frontAnalog_v0p0p1_12.x65.A.t7 a_55268_n74136# GND.t1281 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1169 OUT0.t86 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD.t844 VDD.t843 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1170 VDD.t1161 VDD.t1160 a_77605_n43545# VDD.t741 sky130_fd_pr__pfet_01v8_hvt ad=0.312 pd=1.68 as=0.0588 ps=0.7 w=0.42 l=0.15
X1171 16to4_PriorityEncoder_v0p0p1_0.x22.A 16to4_PriorityEncoder_v0p0p1_0.x21.A VDD.t1294 VDD.t1293 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1172 VDD.t1133 16to4_PriorityEncoder_v0p0p1_0.x5.x21.B a_78097_n45737# VDD.t1132 sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X1173 frontAnalog_v0p0p1_4.RSfetsym_0.x1.Y frontAnalog_v0p0p1_4.x63.X VDD.t121 VDD.t119 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1174 a_59577_n79083# frontAnalog_v0p0p1_14.x63.X I1.t0 GND.t356 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1175 a_77855_n48109# I5.t11 a_77783_n48109# VDD.t1060 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X1176 a_78349_n43045# 16to4_PriorityEncoder_v0p0p1_0.x5.x16.X GND.t858 GND.t175 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X1177 GND.t1048 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t30 GND.t1047 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1178 a_77605_n45765# 16to4_PriorityEncoder_v0p0p1_0.x5.x19.D VDD.t658 VDD.t657 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X1179 GND.t1454 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t26 GND.t1453 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1180 frontAnalog_v0p0p1_0.RSfetsym_0.QN.t3 I14.t8 VDD.t130 VDD.t129 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.3
X1181 frontAnalog_v0p0p1_10.x63.A.t1 frontAnalog_v0p0p1_10.x65.A.t5 VDD.t694 VDD.t562 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1182 GND.t1289 frontAnalog_v0p0p1_2.x65.X frontAnalog_v0p0p1_2.RSfetsym_0.x2.Y GND.t1288 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1183 a_55268_n3936# CLK.t50 GND.t599 GND.t598 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1184 frontAnalog_v0p0p1_1.RSfetsym_0.x1.Y frontAnalog_v0p0p1_1.x63.X VDD.t172 VDD.t168 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1185 OUT3.t82 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD.t242 VDD.t241 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1186 a_53630_n30996# frontAnalog_v0p0p1_10.IB.t19 GND.t1125 GND.t36 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1187 16to4_PriorityEncoder_v0p0p1_0.x29.Y 16to4_PriorityEncoder_v0p0p1_0.x29.A GND.t539 GND.t538 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1188 GND.t445 16to4_PriorityEncoder_v0p0p1_0.x22.A 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND.t444 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1189 OUT3.t21 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND.t259 GND.t258 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1190 16to4_PriorityEncoder_v0p0p1_0.x5.x19.C I12.t9 GND.t803 GND.t802 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1191 VDD.t1114 frontAnalog_v0p0p1_13.x65.X frontAnalog_v0p0p1_13.RSfetsym_0.x2.Y VDD.t1109 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1192 a_59578_n46170# frontAnalog_v0p0p1_8.x65.X frontAnalog_v0p0p1_8.RSfetsym_0.QN.t2 GND.t1395 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.315 ps=2.72 w=1 l=0.15
X1193 VDD.t65 16to4_PriorityEncoder_v0p0p1_0.x35.A 16to4_PriorityEncoder_v0p0p1_0.x36.A VDD.t64 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1194 I2.t2 frontAnalog_v0p0p1_12.x63.X VDD.t114 VDD.t111 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.25
X1195 frontAnalog_v0p0p1_3.x63.A.t2 frontAnalog_v0p0p1_3.x65.A.t5 VDD.t677 VDD.t676 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1196 VDD.t768 R1.t6 S1.t3 VDD.t386 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1197 OUT3.t81 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD.t240 VDD.t239 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1198 frontAnalog_v0p0p1_4.x65.X a_57123_n18759# VDD.t96 VDD.t95 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1199 OUT2.t29 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND.t1046 GND.t1045 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1200 OUT2.t88 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD.t976 VDD.t975 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1201 VDD.t620 16to4_PriorityEncoder_v0p0p1_0.x43.A 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD.t619 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1202 OUT1.t88 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD.t1386 VDD.t1385 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1203 frontAnalog_v0p0p1_6.RSfetsym_0.QN.t3 frontAnalog_v0p0p1_6.RSfetsym_0.x1.Y GND.t1259 GND.t851 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.25
X1204 VDD.t1237 16to4_PriorityEncoder_v0p0p1_0.x3.EI a_77605_n51585# VDD.t176 sky130_fd_pr__pfet_01v8_hvt ad=0.312 pd=1.68 as=0.0588 ps=0.7 w=0.42 l=0.15
X1205 16to4_PriorityEncoder_v0p0p1_0.x3.A1 a_78349_n51085# GND.t1342 GND.t738 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.102 ps=0.99 w=0.65 l=0.15
X1206 VV7.t12 VV6.t12 GND.t24 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1207 VDD.t431 16to4_PriorityEncoder_v0p0p1_0.x22.A 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD.t430 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1208 OUT1.t25 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND.t1452 GND.t1451 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1209 VDD.t599 frontAnalog_v0p0p1_8.x63.A.t5 a_57123_n47279# VDD.t598 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1210 VDD.t1277 16to4_PriorityEncoder_v0p0p1_0.x3.x21.B a_78097_n53777# VDD.t1276 sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X1211 VDD.t780 CLK.t51 w_55000_n51528# GND.t837 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1212 I10.t2 frontAnalog_v0p0p1_6.x63.X VDD.t593 VDD.t590 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.25
X1213 VDD.t180 frontAnalog_v0p0p1_7.x63.A.t5 frontAnalog_v0p0p1_7.x65.A.t0 VDD.t179 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1214 GND.t257 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t20 GND.t256 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1215 a_77605_n53805# 16to4_PriorityEncoder_v0p0p1_0.x3.x19.D VDD.t1205 VDD.t1204 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X1216 frontAnalog_v0p0p1_11.RSfetsym_0.x2.Y frontAnalog_v0p0p1_11.x65.X GND.t764 GND.t763 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1217 a_55268_n68736# CLK.t52 GND.t839 GND.t838 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1218 OUT3.t80 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD.t238 VDD.t237 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1219 VV16.t1 VV15.t2 GND.t52 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1220 VDD.t781 CLK.t53 w_55000_n52150# GND.t732 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1221 VV5.t5 VV4.t4 GND.t77 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1222 16to4_PriorityEncoder_v0p0p1_0.x3.x18.C I2.t9 VDD.t792 VDD.t791 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1223 VDD.t171 frontAnalog_v0p0p1_1.x63.X I8.t1 VDD.t170 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.25
X1224 OUT3.t19 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND.t255 GND.t254 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1225 frontAnalog_v0p0p1_12.RSfetsym_0.QN.t4 I2.t10 VDD.t794 VDD.t793 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.3
X1226 a_77759_n53805# 16to4_PriorityEncoder_v0p0p1_0.x3.x19.D a_77687_n53805# GND.t1275 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X1227 frontAnalog_v0p0p1_9.x65.X a_57123_n51159# GND.t1260 GND.t1253 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1228 w_55000_n40728# CLK.t54 frontAnalog_v0p0p1_1.x65.A.t1 VDD.t159 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1229 VDD.t236 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t79 VDD.t235 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1230 I15.t4 frontAnalog_v0p0p1_2.RSfetsym_0.x2.Y GND.t1121 GND.t374 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.25
X1231 GND.t1343 I14.t9 a_77605_n40069# GND.t90 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X1232 GND.t253 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t18 GND.t252 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1233 frontAnalog_v0p0p1_11.x65.A.t2 frontAnalog_v0p0p1_11.x63.A.t6 a_55268_n63336# GND.t602 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1234 a_53630_n47196# VV8.t16 w_55000_n46128# GND.t673 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1235 a_78349_n51085# 16to4_PriorityEncoder_v0p0p1_0.x3.x22.A GND.t1529 GND.t14 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1236 GND.t1345 I14.t10 a_59578_n8370# GND.t1344 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1237 frontAnalog_v0p0p1_12.RSfetsym_0.x2.Y frontAnalog_v0p0p1_12.x65.X VDD.t187 VDD.t185 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1238 a_77637_n41087# VDD.t1158 VDD.t1159 VDD.t72 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X1239 a_55268_n25536# CLK.t55 GND.t841 GND.t840 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1240 frontAnalog_v0p0p1_12.RSfetsym_0.x1.Y frontAnalog_v0p0p1_12.x63.X GND.t131 GND.t129 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1241 a_78243_n49349# 16to4_PriorityEncoder_v0p0p1_0.x3.x17.A a_78147_n49349# VDD.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X1242 GND.t1219 frontAnalog_v0p0p1_14.x65.X frontAnalog_v0p0p1_14.RSfetsym_0.x2.Y GND.t1218 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1243 OUT1.t24 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND.t1450 GND.t1449 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1244 a_82988_n47995# 16to4_PriorityEncoder_v0p0p1_0.x3.A1 a_82906_n47995# VDD.t47 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X1245 GND.t1448 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t23 GND.t1447 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1246 a_77687_n40069# I15.t6 a_77605_n40069# VDD.t752 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X1247 VDD.t120 frontAnalog_v0p0p1_4.x63.X frontAnalog_v0p0p1_4.RSfetsym_0.x1.Y VDD.t119 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1248 VDD.t234 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t78 VDD.t233 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1249 frontAnalog_v0p0p1_0.x65.A.t3 frontAnalog_v0p0p1_0.x63.A.t4 a_55268_n9336# GND.t661 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1250 GND.t1446 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t22 GND.t1445 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1251 OUT2.t87 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD.t974 VDD.t973 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1252 a_77687_n44527# 16to4_PriorityEncoder_v0p0p1_0.x5.x19.C a_77605_n44527# GND.t528 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.109 ps=1.36 w=0.42 l=0.15
X1253 GND.t407 16to4_PriorityEncoder_v0p0p1_0.x5.A2 a_82906_n43855# GND.t406 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X1254 VDD.t169 frontAnalog_v0p0p1_1.x63.X frontAnalog_v0p0p1_1.RSfetsym_0.x1.Y VDD.t168 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1255 frontAnalog_v0p0p1_15.RSfetsym_0.x1.Y frontAnalog_v0p0p1_15.x63.X VDD.t484 VDD.t480 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1256 VDD.t648 frontAnalog_v0p0p1_0.x63.A.t5 a_57123_n9479# VDD.t647 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1257 frontAnalog_v0p0p1_6.RSfetsym_0.x2.Y frontAnalog_v0p0p1_6.x65.X VDD.t10 VDD.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1258 GND.t902 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t21 GND.t901 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1259 frontAnalog_v0p0p1_13.x63.X a_57123_n68879# VDD.t88 VDD.t87 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1260 frontAnalog_v0p0p1_6.RSfetsym_0.x1.Y frontAnalog_v0p0p1_6.x63.X GND.t614 GND.t612 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1261 GND.t1266 frontAnalog_v0p0p1_7.x65.X frontAnalog_v0p0p1_7.RSfetsym_0.x2.Y GND.t1265 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1262 VV12.t7 VV11.t5 GND.t432 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1263 a_77783_n39305# I10.t9 a_77687_n39305# VDD.t127 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X1264 VIN.t23 w_55000_n56928# error sky130_fd_pr__cap_var_lvt w=2 l=0.18
X1265 16to4_PriorityEncoder_v0p0p1_0.x22.Y 16to4_PriorityEncoder_v0p0p1_0.x22.A GND.t443 GND.t442 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1266 VDD.t618 16to4_PriorityEncoder_v0p0p1_0.x43.A 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD.t617 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1267 frontAnalog_v0p0p1_0.x63.X a_57123_n9479# GND.t717 GND.t716 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1268 VDD.t1332 frontAnalog_v0p0p1_8.x65.X frontAnalog_v0p0p1_8.RSfetsym_0.QN.t3 VDD.t1331 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.25
X1269 GND.t1316 I6.t11 a_77605_n48109# GND.t20 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X1270 OUT1.t21 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND.t1444 GND.t1443 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1271 GND.t1442 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t20 GND.t1441 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1272 OUT2.t86 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD.t972 VDD.t971 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1273 OUT3.t77 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD.t232 VDD.t231 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1274 frontAnalog_v0p0p1_10.x65.A.t0 CLK.t56 frontAnalog_v0p0p1_10.x63.A.t2 VDD.t782 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1275 frontAnalog_v0p0p1_5.x63.X a_57123_n25679# VDD.t715 VDD.t714 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1276 frontAnalog_v0p0p1_14.RSfetsym_0.x2.Y frontAnalog_v0p0p1_14.x65.X VDD.t1125 VDD.t1123 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1277 GND.t811 frontAnalog_v0p0p1_8.x63.X frontAnalog_v0p0p1_8.RSfetsym_0.x1.Y GND.t809 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1278 VV8.t6 VV7.t9 GND.t106 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1279 VIN.t24 w_55000_n13728# error sky130_fd_pr__cap_var_lvt w=2 l=0.18
X1280 R1.t3 S1.t6 VDD.t582 VDD.t581 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1281 VDD.t842 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t85 VDD.t841 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1282 VDD.t1228 frontAnalog_v0p0p1_2.x65.X frontAnalog_v0p0p1_2.RSfetsym_0.QN.t3 VDD.t1227 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.25
X1283 frontAnalog_v0p0p1_0.RSfetsym_0.x1.Y frontAnalog_v0p0p1_0.x63.X GND.t371 GND.t369 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1284 frontAnalog_v0p0p1_15.x65.X a_57123_n83559# VDD.t772 VDD.t771 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1285 GND.t1044 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t28 GND.t1043 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1286 frontAnalog_v0p0p1_14.x63.X a_57123_n79679# GND.t1324 GND.t1318 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1287 a_53630_n52596# frontAnalog_v0p0p1_10.IB.t20 GND.t1126 GND.t36 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1288 16to4_PriorityEncoder_v0p0p1_0.x36.Y 16to4_PriorityEncoder_v0p0p1_0.x36.A VDD.t1477 VDD.t1476 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1289 frontAnalog_v0p0p1_12.x63.A.t1 CLK.t57 w_55000_n73750# VDD.t750 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1290 16to4_PriorityEncoder_v0p0p1_0.x22.Y 16to4_PriorityEncoder_v0p0p1_0.x22.A VDD.t429 VDD.t428 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1291 GND.t251 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t17 GND.t250 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1292 VV2.t9 VV1.t11 GND.t33 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1293 GND.t734 frontAnalog_v0p0p1_10.x65.A.t6 a_57123_n56559# GND.t591 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X1294 OUT0.t20 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND.t900 GND.t899 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1295 a_77687_n52567# 16to4_PriorityEncoder_v0p0p1_0.x3.x19.C a_77605_n52567# GND.t153 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.109 ps=1.36 w=0.42 l=0.15
X1296 OUT3.t76 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD.t230 VDD.t229 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1297 frontAnalog_v0p0p1_10.x63.A.t0 frontAnalog_v0p0p1_10.x65.A.t7 a_55268_n57936# GND.t735 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1298 GND.t762 frontAnalog_v0p0p1_11.x65.X frontAnalog_v0p0p1_11.RSfetsym_0.x2.Y GND.t761 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1299 GND.t677 16to4_PriorityEncoder_v0p0p1_0.x5.x19.D a_77881_n44527# GND.t528 sky130_fd_pr__nfet_01v8 ad=0.196 pd=1.33 as=0.0693 ps=0.75 w=0.42 l=0.15
X1300 frontAnalog_v0p0p1_3.x65.A.t1 CLK.t58 frontAnalog_v0p0p1_3.x63.A.t0 VDD.t567 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1301 I5.t4 frontAnalog_v0p0p1_10.RSfetsym_0.QN.t5 VDD.t1129 VDD.t1061 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.3
X1302 frontAnalog_v0p0p1_7.RSfetsym_0.x2.Y frontAnalog_v0p0p1_7.x65.X VDD.t1198 VDD.t1196 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1303 VDD.t787 frontAnalog_v0p0p1_10.x63.X frontAnalog_v0p0p1_10.RSfetsym_0.x1.Y VDD.t783 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1304 VDD.t228 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t75 VDD.t227 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1305 VDD.t483 frontAnalog_v0p0p1_15.x63.X I0.t2 VDD.t482 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.25
X1306 VDD.t1384 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t87 VDD.t1383 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1307 frontAnalog_v0p0p1_4.RSfetsym_0.x2.Y frontAnalog_v0p0p1_4.x65.X GND.t492 GND.t491 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1308 w_55000_n83928# CLK.t59 S0.t3 VDD.t97 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1309 16to4_PriorityEncoder_v0p0p1_0.x5.x2.X a_77605_n40069# GND.t405 GND.t404 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.102 ps=0.99 w=0.65 l=0.15
X1310 a_77783_n47345# I2.t11 a_77687_n47345# VDD.t795 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X1311 frontAnalog_v0p0p1_1.x65.X a_57123_n40359# VDD.t1280 VDD.t1279 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1312 a_16719_n13117.t14 a_16599_n13205.t13 a_16541_n13117.t18 GND.t1356 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1313 frontAnalog_v0p0p1_7.x63.X a_57123_n36479# GND.t367 GND.t366 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1314 VV6.t17 w_55000_n57550# error sky130_fd_pr__cap_var_lvt w=2 l=0.18
X1315 OUT2.t85 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD.t970 VDD.t969 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1316 GND.t693 frontAnalog_v0p0p1_3.x65.A.t6 a_57123_n13359# GND.t120 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X1317 a_78527_n43045# 16to4_PriorityEncoder_v0p0p1_0.x5.x15.X a_78431_n43045# VDD.t167 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X1318 frontAnalog_v0p0p1_9.RSfetsym_0.QN.t0 frontAnalog_v0p0p1_9.RSfetsym_0.x1.Y GND.t822 GND.t821 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.25
X1319 frontAnalog_v0p0p1_2.RSfetsym_0.x2.Y frontAnalog_v0p0p1_2.x65.X VDD.t1226 VDD.t1224 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1320 VV16.t13 VV15.t10 GND.t202 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1321 frontAnalog_v0p0p1_3.x63.A.t3 frontAnalog_v0p0p1_3.x65.A.t7 a_55268_n14736# GND.t694 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1322 GND.t130 frontAnalog_v0p0p1_12.x63.X frontAnalog_v0p0p1_12.RSfetsym_0.x1.Y GND.t129 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1323 OUT1.t19 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND.t1440 GND.t1439 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1324 OUT2.t84 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD.t968 VDD.t967 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1325 VDD.t966 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t83 VDD.t965 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1326 VDD.t1475 16to4_PriorityEncoder_v0p0p1_0.x36.A 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD.t1474 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1327 OUT0.t84 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD.t840 VDD.t839 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1328 GND.t1 I4.t10 a_77723_n48817# GND.t0 sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X1329 I13.t0 frontAnalog_v0p0p1_3.RSfetsym_0.QN.t5 VDD.t416 VDD.t70 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.3
X1330 frontAnalog_v0p0p1_0.x65.X a_57123_n7959# GND.t1231 GND.t716 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1331 VDD.t470 frontAnalog_v0p0p1_3.x63.X frontAnalog_v0p0p1_3.RSfetsym_0.x1.Y VDD.t464 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1332 a_59577_n19683# frontAnalog_v0p0p1_4.x63.X I12.t0 GND.t137 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1333 OUT0.t19 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND.t898 GND.t897 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1334 a_59578_n29970# frontAnalog_v0p0p1_6.x65.X frontAnalog_v0p0p1_6.RSfetsym_0.QN.t0 GND.t6 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.315 ps=2.72 w=1 l=0.15
X1335 a_53630_n68796# frontAnalog_v0p0p1_10.IB.t21 GND.t1127 GND.t36 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1336 GND.t896 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t18 GND.t895 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1337 a_77605_n40069# I15.t7 GND.t801 GND.t90 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X1338 VV14.t17 w_55000_n14350# error sky130_fd_pr__cap_var_lvt w=2 l=0.18
X1339 GND.t894 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t17 GND.t893 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1340 frontAnalog_v0p0p1_9.RSfetsym_0.x1.Y frontAnalog_v0p0p1_9.x63.X GND.t1190 GND.t1188 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1341 a_16719_n13117.t13 a_16599_n13205.t14 a_16541_n13117.t17 GND.t1357 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1342 a_77637_n40777# VDD.t1155 VDD.t1157 VDD.t1156 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X1343 VDD.t481 frontAnalog_v0p0p1_15.x63.X frontAnalog_v0p0p1_15.RSfetsym_0.x1.Y VDD.t480 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1344 VDD.t1382 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t86 VDD.t1381 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1345 GND.t613 frontAnalog_v0p0p1_6.x63.X frontAnalog_v0p0p1_6.RSfetsym_0.x1.Y GND.t612 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1346 16to4_PriorityEncoder_v0p0p1_0.x43.A 16to4_PriorityEncoder_v0p0p1_0.x42.A GND.t416 GND.t415 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1347 GND.t1321 frontAnalog_v0p0p1_12.RSfetsym_0.QN.t6 a_59577_n73683# GND.t1320 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1348 OUT2.t27 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND.t1042 GND.t1041 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1349 GND.t1142 I0.t8 a_59578_n83970# GND.t1141 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1350 a_78147_n49349# 16to4_PriorityEncoder_v0p0p1_0.x3.x22.A a_78065_n49349# VDD.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X1351 GND.t1274 16to4_PriorityEncoder_v0p0p1_0.x3.x19.D a_77881_n52567# GND.t153 sky130_fd_pr__nfet_01v8 ad=0.196 pd=1.33 as=0.0693 ps=0.75 w=0.42 l=0.15
X1352 OUT1.t85 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD.t1380 VDD.t1379 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1353 16to4_PriorityEncoder_v0p0p1_0.x5.x19.X a_77605_n44779# GND.t1385 GND.t1384 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.196 ps=1.33 w=0.65 l=0.15
X1354 GND.t1040 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t26 GND.t1039 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1355 a_82906_n43855# 16to4_PriorityEncoder_v0p0p1_0.x3.A2 GND.t1315 GND.t1314 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1356 VDD.t964 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t82 VDD.t963 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1357 a_78313_n39305# 16to4_PriorityEncoder_v0p0p1_0.x5.x1.X a_78241_n39305# VDD.t578 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X1358 VV8.t0 VV7.t3 GND.t77 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1359 VV10.t2 VV9.t1 GND.t33 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1360 I13.t3 frontAnalog_v0p0p1_3.x63.X VDD.t469 VDD.t466 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.25
X1361 a_53630_n25596# frontAnalog_v0p0p1_10.IB.t22 GND.t1128 GND.t36 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1362 a_16719_n13117.t12 a_16599_n13205.t15 a_16541_n13117.t16 GND.t1358 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1363 VDD.t1120 frontAnalog_v0p0p1_4.x63.A.t7 frontAnalog_v0p0p1_4.x65.A.t3 VDD.t421 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1364 frontAnalog_v0p0p1_11.RSfetsym_0.x1.Y frontAnalog_v0p0p1_11.x63.X VDD.t494 VDD.t492 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1365 OUT0.t83 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD.t838 VDD.t837 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1366 GND.t805 I12.t10 a_59578_n19170# GND.t804 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1367 VV3.t8 VV2.t8 GND.t709 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1368 VDD.t836 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t82 VDD.t835 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1369 VV13.t15 VV12.t15 GND.t33 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1370 OUT0.t16 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND.t892 GND.t891 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1371 GND.t890 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t15 GND.t889 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1372 VV5.t1 VV4.t2 GND.t51 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1373 VDD.t1124 frontAnalog_v0p0p1_14.x65.X frontAnalog_v0p0p1_14.RSfetsym_0.x2.Y VDD.t1123 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1374 a_78527_n51085# 16to4_PriorityEncoder_v0p0p1_0.x3.x15.X a_78431_n51085# VDD.t1281 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X1375 GND.t80 16to4_PriorityEncoder_v0p0p1_0.x35.A 16to4_PriorityEncoder_v0p0p1_0.x36.A GND.t79 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1376 VDD.t962 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t81 VDD.t961 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1377 VDD.t834 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t81 VDD.t833 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1378 16to4_PriorityEncoder_v0p0p1_0.x3.A0 a_78525_n53555# GND.t1199 GND.t1198 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.102 ps=0.99 w=0.65 l=0.15
X1379 GND.t525 frontAnalog_v0p0p1_6.RSfetsym_0.QN.t6 a_59577_n30483# GND.t524 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1380 frontAnalog_v0p0p1_10.RSfetsym_0.QN.t4 I5.t12 VDD.t1062 VDD.t1061 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.3
X1381 frontAnalog_v0p0p1_7.x65.X a_57123_n34959# GND.t1317 GND.t366 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1382 GND.t522 I8.t7 a_59578_n40770# GND.t521 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1383 frontAnalog_v0p0p1_10.IB.t0 a_16719_n13117.t24 VDD.t1286 VDD.t1285 sky130_fd_pr__pfet_01v8_lvt ad=5.51 pd=38.6 as=5.51 ps=38.6 w=19 l=1
X1384 a_77687_n39305# I11.t10 a_77605_n39305# VDD.t1137 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X1385 VDD.t1378 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t84 VDD.t1377 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1386 OUT1.t83 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD.t1376 VDD.t1375 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1387 OUT2.t25 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND.t1038 GND.t1037 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1388 GND.t1036 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t24 GND.t1035 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1389 16to4_PriorityEncoder_v0p0p1_0.x3.x14.A a_77637_n48817# VDD.t1265 VDD.t1264 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.167 ps=1.39 w=1 l=0.15
X1390 a_77605_n48109# I7.t7 GND.t1311 GND.t20 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X1391 VDD.t202 frontAnalog_v0p0p1_8.x65.A.t4 a_57123_n45759# VDD.t201 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1392 VDD.t1197 frontAnalog_v0p0p1_7.x65.X frontAnalog_v0p0p1_7.RSfetsym_0.x2.Y VDD.t1196 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1393 16to4_PriorityEncoder_v0p0p1_0.x5.x16.C I13.t11 VDD.t69 VDD.t68 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1394 VV2.t13 VV1.t14 GND.t78 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1395 VFS.t5 VV16.t10 GND.t422 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1396 frontAnalog_v0p0p1_3.RSfetsym_0.QN.t0 I13.t12 VDD.t71 VDD.t70 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.3
X1397 OUT0.t80 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD.t832 VDD.t831 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1398 VDD.t830 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t79 VDD.t829 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1399 GND.t702 VDD.t1508 a_78735_n39527# GND.t701 sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X1400 VDD.t1288 a_16719_n13117.t25 a_16599_n13205.t1 VDD.t1287 sky130_fd_pr__pfet_01v8_lvt ad=5.51 pd=38.6 as=5.51 ps=38.6 w=19 l=1
X1401 OUT1.t82 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD.t1374 VDD.t1373 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1402 VV4.t0 VV3.t1 GND.t52 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1403 16to4_PriorityEncoder_v0p0p1_0.x3.x19.X a_77605_n52819# GND.t391 GND.t390 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.196 ps=1.33 w=0.65 l=0.15
X1404 16to4_PriorityEncoder_v0p0p1_0.x36.A 16to4_PriorityEncoder_v0p0p1_0.x35.A VDD.t63 VDD.t62 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1405 VDD.t517 16to4_PriorityEncoder_v0p0p1_0.x29.A 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD.t516 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1406 16to4_PriorityEncoder_v0p0p1_0.x3.x21.X a_78097_n53777# GND.t173 GND.t172 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.112 ps=1.04 w=0.65 l=0.15
X1407 w_55000_n62950# VIN.t25 a_53630_n63396# GND.t671 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1408 frontAnalog_v0p0p1_15.RSfetsym_0.x2.Y frontAnalog_v0p0p1_15.x65.X GND.t209 GND.t208 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1409 a_78313_n47345# 16to4_PriorityEncoder_v0p0p1_0.x3.x1.X a_78241_n47345# VDD.t682 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X1410 16to4_PriorityEncoder_v0p0p1_0.x36.Y 16to4_PriorityEncoder_v0p0p1_0.x36.A GND.t1549 GND.t1548 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1411 VDD.t1225 frontAnalog_v0p0p1_2.x65.X frontAnalog_v0p0p1_2.RSfetsym_0.x2.Y VDD.t1224 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1412 frontAnalog_v0p0p1_13.RSfetsym_0.x1.Y frontAnalog_v0p0p1_13.x63.X VDD.t376 VDD.t372 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1413 16to4_PriorityEncoder_v0p0p1_0.x3.x19.C I4.t11 VDD.t3 VDD.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1414 frontAnalog_v0p0p1_4.RSfetsym_0.QN.t2 frontAnalog_v0p0p1_4.x65.X VDD.t477 VDD.t472 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.25
X1415 frontAnalog_v0p0p1_3.RSfetsym_0.x1.Y frontAnalog_v0p0p1_3.x63.X GND.t484 GND.t482 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1416 VFS.t7 VV16.t12 GND.t214 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1417 OUT0.t14 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND.t888 GND.t887 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1418 a_77687_n47345# I3.t11 a_77605_n47345# VDD.t178 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X1419 VDD.t960 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t80 VDD.t959 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1420 VDD.t1372 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t81 VDD.t1371 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1421 frontAnalog_v0p0p1_1.RSfetsym_0.x2.Y frontAnalog_v0p0p1_1.x65.X GND.t752 GND.t751 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1422 frontAnalog_v0p0p1_5.RSfetsym_0.x1.Y frontAnalog_v0p0p1_5.x63.X VDD.t23 VDD.t19 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1423 a_59577_n84483# frontAnalog_v0p0p1_15.x63.X I0.t1 GND.t499 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1424 a_77775_n44779# I11.t11 a_77687_n44779# GND.t678 sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
X1425 OUT2.t23 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND.t1034 GND.t1033 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1426 I4.t0 frontAnalog_v0p0p1_11.RSfetsym_0.x2.Y GND.t157 GND.t156 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.25
X1427 16to4_PriorityEncoder_v0p0p1_0.x29.Y 16to4_PriorityEncoder_v0p0p1_0.x29.A VDD.t515 VDD.t514 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1428 frontAnalog_v0p0p1_11.x63.A.t3 frontAnalog_v0p0p1_11.x65.A.t5 VDD.t1151 VDD.t687 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1429 VDD.t151 frontAnalog_v0p0p1_0.x65.A.t5 a_57123_n7959# VDD.t150 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1430 GND.t1547 16to4_PriorityEncoder_v0p0p1_0.x36.A 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND.t1546 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1431 GND.t1300 16to4_PriorityEncoder_v0p0p1_0.x3.EI a_78735_n47567# GND.t1299 sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X1432 VDD.t568 CLK.t60 w_55000_n78528# GND.t161 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1433 OUT0.t78 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD.t828 VDD.t827 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1434 I5.t2 frontAnalog_v0p0p1_10.x63.X VDD.t786 VDD.t785 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.25
X1435 GND.t1155 16to4_PriorityEncoder_v0p0p1_0.x28.A 16to4_PriorityEncoder_v0p0p1_0.x29.A GND.t1154 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1436 a_77605_n44779# 16to4_PriorityEncoder_v0p0p1_0.x5.x19.C VDD.t740 VDD.t739 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X1437 VDD.t186 frontAnalog_v0p0p1_12.x65.X frontAnalog_v0p0p1_12.RSfetsym_0.x2.Y VDD.t185 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1438 GND.t1298 16to4_PriorityEncoder_v0p0p1_0.x3.EI a_77759_n53805# GND.t1297 sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X1439 a_59577_n41283# frontAnalog_v0p0p1_1.x63.X I8.t0 GND.t179 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1440 VV10.t7 VV9.t7 GND.t78 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1441 a_59578_n51570# frontAnalog_v0p0p1_9.x65.X frontAnalog_v0p0p1_9.RSfetsym_0.QN.t2 GND.t1329 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.315 ps=2.72 w=1 l=0.15
X1442 VDD.t375 frontAnalog_v0p0p1_13.x63.X I3.t2 VDD.t374 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.25
X1443 VDD.t569 CLK.t61 w_55000_n79150# GND.t593 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1444 frontAnalog_v0p0p1_4.x63.A.t1 frontAnalog_v0p0p1_4.x65.A.t6 VDD.t1252 VDD.t689 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1445 I12.t4 frontAnalog_v0p0p1_4.RSfetsym_0.x2.Y GND.t1197 GND.t1196 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.25
X1446 w_55000_n67728# CLK.t62 frontAnalog_v0p0p1_13.x65.A.t3 VDD.t570 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1447 VDD.t604 R0.t7 S0.t1 VDD.t559 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1448 OUT1.t18 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND.t1438 GND.t1437 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1449 frontAnalog_v0p0p1_14.x65.X a_57123_n78159# GND.t1319 GND.t1318 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1450 VV13.t4 VV12.t4 GND.t78 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1451 frontAnalog_v0p0p1_5.x65.X a_57123_n24159# VDD.t463 VDD.t462 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1452 frontAnalog_v0p0p1_4.x63.X a_57123_n20279# GND.t514 GND.t110 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1453 GND.t1032 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t22 GND.t1031 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1454 frontAnalog_v0p0p1_3.x63.A.t1 CLK.t63 w_55000_n14350# VDD.t103 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1455 VDD.t571 CLK.t64 w_55000_n35328# GND.t594 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1456 GND.t471 16to4_PriorityEncoder_v0p0p1_0.x5.x19.X a_78525_n45515# GND.t470 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X1457 frontAnalog_v0p0p1_7.RSfetsym_0.QN.t1 frontAnalog_v0p0p1_7.RSfetsym_0.x1.Y GND.t584 GND.t583 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.25
X1458 VDD.t9 frontAnalog_v0p0p1_6.x65.X frontAnalog_v0p0p1_6.RSfetsym_0.x2.Y VDD.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1459 frontAnalog_v0p0p1_8.RSfetsym_0.x2.Y frontAnalog_v0p0p1_8.x65.X GND.t1394 GND.t1393 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1460 VDD.t344 frontAnalog_v0p0p1_9.x63.A.t5 a_57123_n52679# VDD.t343 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1461 VDD.t22 frontAnalog_v0p0p1_5.x63.X I11.t1 VDD.t21 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.25
X1462 VDD.t1086 CLK.t65 w_55000_n35950# GND.t1158 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1463 OUT1.t80 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD.t1370 VDD.t1369 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1464 16to4_PriorityEncoder_v0p0p1_0.x29.A 16to4_PriorityEncoder_v0p0p1_0.x28.A VDD.t1076 VDD.t1075 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1465 w_55000_n24528# CLK.t66 frontAnalog_v0p0p1_5.x65.A.t0 VDD.t93 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1466 GND.t249 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t16 GND.t248 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1467 a_16719_n13117.t1 a_16719_n13117.t0 VDD.t1056 VDD.t1055 sky130_fd_pr__pfet_01v8_lvt ad=5.51 pd=38.6 as=5.51 ps=38.6 w=19 l=1
X1468 a_53630_n3996# frontAnalog_v0p0p1_10.IB.t23 GND.t790 GND.t384 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1469 GND.t1030 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t21 GND.t1029 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1470 a_55268_n74136# CLK.t67 GND.t1165 GND.t1164 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1471 16to4_PriorityEncoder_v0p0p1_0.x43.Y 16to4_PriorityEncoder_v0p0p1_0.x43.A VDD.t616 VDD.t615 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1472 frontAnalog_v0p0p1_8.x65.A.t3 frontAnalog_v0p0p1_8.x63.A.t6 a_55268_n47136# GND.t1338 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1473 VDD.t1284 I14.t11 a_77637_n42017# VDD.t1163 sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X1474 16to4_PriorityEncoder_v0p0p1_0.x5.EO a_78159_n39549# GND.t689 GND.t688 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.102 ps=0.99 w=0.65 l=0.15
X1475 VDD.t373 frontAnalog_v0p0p1_13.x63.X frontAnalog_v0p0p1_13.RSfetsym_0.x1.Y VDD.t372 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1476 a_77605_n52819# 16to4_PriorityEncoder_v0p0p1_0.x3.x19.C VDD.t608 VDD.t607 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X1477 GND.t483 frontAnalog_v0p0p1_3.x63.X frontAnalog_v0p0p1_3.RSfetsym_0.x1.Y GND.t482 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1478 frontAnalog_v0p0p1_10.RSfetsym_0.x2.Y frontAnalog_v0p0p1_10.x65.X VDD.t80 VDD.t78 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1479 VFS.t2 VV16.t6 GND.t394 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1480 frontAnalog_v0p0p1_10.RSfetsym_0.x1.Y frontAnalog_v0p0p1_10.x63.X GND.t844 GND.t842 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1481 a_53630_n52596# VV7.t17 w_55000_n51528# GND.t1148 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1482 a_16719_n13117.t11 a_16599_n13205.t16 a_16541_n13117.t15 GND.t1359 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1483 VV3.t13 VV2.t12 GND.t432 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1484 VDD.t226 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t74 VDD.t225 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1485 VV4.t13 VV3.t14 GND.t202 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1486 GND.t370 frontAnalog_v0p0p1_0.x63.X frontAnalog_v0p0p1_0.RSfetsym_0.x1.Y GND.t369 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1487 VV8.t3 VV7.t5 GND.t51 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1488 a_55268_n30936# CLK.t68 GND.t1167 GND.t1166 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1489 GND.t604 frontAnalog_v0p0p1_11.x63.A.t7 a_57123_n63479# GND.t603 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X1490 frontAnalog_v0p0p1_15.RSfetsym_0.QN.t0 frontAnalog_v0p0p1_15.x65.X VDD.t196 VDD.t195 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.25
X1491 GND.t1028 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t20 GND.t1027 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1492 OUT3.t73 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD.t224 VDD.t223 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1493 OUT1.t17 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND.t1436 GND.t1435 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1494 OUT2.t19 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND.t1026 GND.t1025 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1495 VDD.t20 frontAnalog_v0p0p1_5.x63.X frontAnalog_v0p0p1_5.RSfetsym_0.x1.Y VDD.t19 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1496 GND.t105 16to4_PriorityEncoder_v0p0p1_0.x3.x19.X a_78525_n53555# GND.t104 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X1497 frontAnalog_v0p0p1_3.RSfetsym_0.x2.Y frontAnalog_v0p0p1_3.x65.X VDD.t540 VDD.t538 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1498 16to4_PriorityEncoder_v0p0p1_0.x5.EO a_78159_n39549# VDD.t673 VDD.t672 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.148 ps=1.34 w=1 l=0.15
X1499 GND.t490 frontAnalog_v0p0p1_4.x65.X frontAnalog_v0p0p1_4.RSfetsym_0.x2.Y GND.t489 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1500 a_78159_n39549# 16to4_PriorityEncoder_v0p0p1_0.x5.x1.X GND.t601 GND.t600 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1501 OUT3.t72 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD.t222 VDD.t221 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1502 a_53630_n79596# frontAnalog_v0p0p1_10.IB.t24 GND.t791 GND.t36 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1503 frontAnalog_v0p0p1_1.RSfetsym_0.QN.t2 frontAnalog_v0p0p1_1.x65.X VDD.t708 VDD.t707 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.25
X1504 VDD.t7 frontAnalog_v0p0p1_6.x65.X frontAnalog_v0p0p1_6.RSfetsym_0.QN.t1 VDD.t6 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.25
X1505 VDD.t513 16to4_PriorityEncoder_v0p0p1_0.x29.A 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD.t512 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1506 OUT3.t15 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND.t247 GND.t246 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1507 16to4_PriorityEncoder_v0p0p1_0.x36.Y 16to4_PriorityEncoder_v0p0p1_0.x36.A GND.t1545 GND.t1544 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1508 16to4_PriorityEncoder_v0p0p1_0.x5.x22.A a_77639_n42341# GND.t350 GND.t349 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.112 ps=1.04 w=0.65 l=0.15
X1509 OUT1.t16 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND.t1434 GND.t1433 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1510 GND.t1351 16to4_PriorityEncoder_v0p0p1_0.x21.A 16to4_PriorityEncoder_v0p0p1_0.x22.A GND.t1350 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1511 VDD.t1269 frontAnalog_v0p0p1_9.x65.X frontAnalog_v0p0p1_9.RSfetsym_0.QN.t3 VDD.t1268 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.25
X1512 16to4_PriorityEncoder_v0p0p1_0.x3.EO a_78159_n47589# GND.t1245 GND.t1244 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.102 ps=0.99 w=0.65 l=0.15
X1513 OUT2.t79 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD.t958 VDD.t957 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1514 VV1.t7 VL.t3 GND.t33 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1515 a_77687_n43295# I10.t10 a_77605_n43295# GND.t703 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.109 ps=1.36 w=0.42 l=0.15
X1516 VDD.t956 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t78 VDD.t955 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1517 frontAnalog_v0p0p1_11.x65.A.t0 CLK.t69 frontAnalog_v0p0p1_11.x63.A.t1 VDD.t1087 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1518 frontAnalog_v0p0p1_13.x65.X a_57123_n67359# VDD.t1203 VDD.t1202 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1519 a_53630_n36396# frontAnalog_v0p0p1_10.IB.t25 GND.t792 GND.t36 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1520 OUT0.t13 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND.t886 GND.t885 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1521 OUT3.t71 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD.t220 VDD.t219 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1522 frontAnalog_v0p0p1_10.x63.A.t3 CLK.t70 w_55000_n57550# VDD.t563 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1523 GND.t1189 frontAnalog_v0p0p1_9.x63.X frontAnalog_v0p0p1_9.RSfetsym_0.x1.Y GND.t1188 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1524 16to4_PriorityEncoder_v0p0p1_0.x29.Y 16to4_PriorityEncoder_v0p0p1_0.x29.A GND.t537 GND.t536 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1525 VV9.t2 VV8.t1 GND.t33 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1526 frontAnalog_v0p0p1_14.RSfetsym_0.QN.t0 frontAnalog_v0p0p1_14.RSfetsym_0.x1.Y GND.t359 GND.t200 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.25
X1527 OUT3.t14 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND.t245 GND.t244 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1528 VDD.t218 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t70 VDD.t217 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1529 VV16.t0 VV15.t0 GND.t24 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1530 frontAnalog_v0p0p1_15.x63.X a_57123_n85079# GND.t1567 GND.t823 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1531 GND.t1392 frontAnalog_v0p0p1_8.x65.X frontAnalog_v0p0p1_8.RSfetsym_0.x2.Y GND.t1391 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1532 VV7.t10 VV6.t11 GND.t106 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1533 GND.t243 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t13 GND.t242 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1534 frontAnalog_v0p0p1_4.RSfetsym_0.x2.Y frontAnalog_v0p0p1_4.x65.X VDD.t476 VDD.t474 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1535 GND.t1117 frontAnalog_v0p0p1_11.x65.A.t6 a_57123_n61959# GND.t603 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X1536 VDD.t1292 16to4_PriorityEncoder_v0p0p1_0.x21.A 16to4_PriorityEncoder_v0p0p1_0.x22.A VDD.t1291 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1537 a_16719_n13117.t10 a_16599_n13205.t17 a_16541_n13117.t14 GND.t1360 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1538 16to4_PriorityEncoder_v0p0p1_0.x3.EO a_78159_n47589# VDD.t1148 VDD.t1147 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.148 ps=1.34 w=1 l=0.15
X1539 a_78159_n47589# 16to4_PriorityEncoder_v0p0p1_0.x3.x1.X GND.t715 GND.t714 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1540 VDD.t493 frontAnalog_v0p0p1_11.x63.X frontAnalog_v0p0p1_11.RSfetsym_0.x1.Y VDD.t492 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1541 frontAnalog_v0p0p1_1.RSfetsym_0.x2.Y frontAnalog_v0p0p1_1.x65.X VDD.t706 VDD.t704 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1542 OUT2.t18 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND.t1024 GND.t1023 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1543 frontAnalog_v0p0p1_5.RSfetsym_0.x2.Y frontAnalog_v0p0p1_5.x65.X GND.t1375 GND.t1374 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1544 frontAnalog_v0p0p1_14.RSfetsym_0.x1.Y frontAnalog_v0p0p1_14.x63.X GND.t355 GND.t353 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1545 OUT1.t15 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND.t1432 GND.t1431 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1546 a_78525_n45515# 16to4_PriorityEncoder_v0p0p1_0.x5.x20.X GND.t771 GND.t770 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X1547 OUT0.t77 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD.t826 VDD.t825 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1548 16to4_PriorityEncoder_v0p0p1_0.x5.x19.D I14.t12 VDD.t1315 VDD.t1314 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1549 16to4_PriorityEncoder_v0p0p1_0.x35.A 16to4_PriorityEncoder_v0p0p1_0.x34.A GND.t67 GND.t66 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1550 16to4_PriorityEncoder_v0p0p1_0.x3.x22.A a_77639_n50381# GND.t398 GND.t397 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.112 ps=1.04 w=0.65 l=0.15
X1551 frontAnalog_v0p0p1_1.x63.X a_57123_n41879# GND.t348 GND.t347 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1552 GND.t843 frontAnalog_v0p0p1_10.x63.X frontAnalog_v0p0p1_10.RSfetsym_0.x1.Y GND.t842 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1553 VV5.t17 w_55000_n62950# error sky130_fd_pr__cap_var_lvt w=2 l=0.18
X1554 OUT1.t14 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND.t1430 GND.t1429 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1555 GND.t1428 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t13 GND.t1427 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1556 GND.t535 16to4_PriorityEncoder_v0p0p1_0.x29.A 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND.t534 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1557 a_77605_n44527# 16to4_PriorityEncoder_v0p0p1_0.x5.x18.C VDD.t1328 VDD.t659 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X1558 VDD.t954 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t77 VDD.t953 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1559 a_77881_n43545# 16to4_PriorityEncoder_v0p0p1_0.x5.x16.C a_77775_n43545# GND.t699 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X1560 GND.t704 VDD.t1509 a_77881_n43295# GND.t703 sky130_fd_pr__nfet_01v8 ad=0.196 pd=1.33 as=0.0693 ps=0.75 w=0.42 l=0.15
X1561 a_77725_n42341# VDD.t1510 a_77639_n42341# GND.t705 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X1562 OUT3.t12 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND.t241 GND.t240 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1563 frontAnalog_v0p0p1_7.RSfetsym_0.x1.Y frontAnalog_v0p0p1_7.x63.X GND.t579 GND.t577 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1564 OUT0.t12 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND.t884 GND.t883 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1565 16to4_PriorityEncoder_v0p0p1_0.x5.x20.X a_77605_n45765# GND.t377 GND.t376 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X1566 VDD.t408 16to4_PriorityEncoder_v0p0p1_0.x5.x22.A a_78775_n45515# VDD.t407 sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X1567 GND.t239 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t11 GND.t238 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1568 GND.t3 frontAnalog_v0p0p1_10.RSfetsym_0.QN.t6 a_59577_n57483# GND.t2 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1569 GND.t1116 I3.t12 a_59578_n67770# GND.t1115 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1570 VDD.t952 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t76 VDD.t951 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1571 16to4_PriorityEncoder_v0p0p1_0.x43.Y 16to4_PriorityEncoder_v0p0p1_0.x43.A VDD.t614 VDD.t613 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1572 VDD.t1368 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t79 VDD.t1367 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1573 a_16719_n13117.t9 a_16599_n13205.t18 a_16541_n13117.t13 GND.t1361 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1574 16to4_PriorityEncoder_v0p0p1_0.x43.Y 16to4_PriorityEncoder_v0p0p1_0.x43.A GND.t631 GND.t630 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1575 frontAnalog_v0p0p1_2.x63.X a_57123_n4079# VDD.t1096 VDD.t1095 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1576 GND.t1426 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t12 GND.t1425 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1577 GND.t207 frontAnalog_v0p0p1_15.x65.X frontAnalog_v0p0p1_15.RSfetsym_0.x2.Y GND.t206 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1578 16to4_PriorityEncoder_v0p0p1_0.x29.Y 16to4_PriorityEncoder_v0p0p1_0.x29.A VDD.t511 VDD.t510 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1579 frontAnalog_v0p0p1_8.RSfetsym_0.x1.Y frontAnalog_v0p0p1_8.x63.X VDD.t761 VDD.t759 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1580 VV15.t7 VV14.t7 GND.t52 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1581 a_53630_n30996# frontAnalog_v0p0p1_10.IB.t26 GND.t793 GND.t36 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1582 a_78241_n39305# 16to4_PriorityEncoder_v0p0p1_0.x5.x2.X a_78159_n39549# VDD.t1071 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X1583 OUT0.t11 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND.t882 GND.t881 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1584 GND.t826 frontAnalog_v0p0p1_2.RSfetsym_0.QN.t5 a_59577_n3483# GND.t825 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1585 a_78525_n53555# 16to4_PriorityEncoder_v0p0p1_0.x3.x20.X GND.t365 GND.t364 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X1586 OUT0.t76 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD.t824 VDD.t823 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1587 GND.t1424 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t11 GND.t1423 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1588 16to4_PriorityEncoder_v0p0p1_0.x5.x20.X a_77605_n45765# VDD.t371 VDD.t370 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X1589 GND.t190 frontAnalog_v0p0p1_3.RSfetsym_0.QN.t6 a_59577_n14283# GND.t189 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1590 frontAnalog_v0p0p1_4.x65.X a_57123_n18759# GND.t111 GND.t110 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1591 GND.t816 I11.t12 a_59578_n24570# GND.t815 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1592 GND.t237 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t10 GND.t236 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1593 VV7.t0 VV6.t0 GND.t77 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1594 a_77605_n40069# I13.t13 GND.t91 GND.t90 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1595 a_16719_n13117.t8 a_16599_n13205.t19 a_16541_n13117.t12 GND.t832 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1596 frontAnalog_v0p0p1_12.x63.X a_57123_n74279# VDD.t1190 VDD.t1189 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1597 VV1.t9 VL.t5 GND.t78 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1598 a_77881_n51585# 16to4_PriorityEncoder_v0p0p1_0.x3.x16.C a_77775_n51585# GND.t174 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X1599 16to4_PriorityEncoder_v0p0p1_0.x5.A2 a_78065_n41309# VDD.t411 VDD.t52 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.148 ps=1.34 w=1 l=0.15
X1600 GND.t750 frontAnalog_v0p0p1_1.x65.X frontAnalog_v0p0p1_1.RSfetsym_0.x2.Y GND.t749 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1601 VIN.t26 w_55000_n62328# error sky130_fd_pr__cap_var_lvt w=2 l=0.18
X1602 OUT2.t75 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD.t950 VDD.t949 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1603 GND.t15 16to4_PriorityEncoder_v0p0p1_0.x3.x17.A a_78349_n51085# GND.t14 sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X1604 VDD.t413 frontAnalog_v0p0p1_6.x65.A.t6 a_57123_n29559# VDD.t412 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1605 16to4_PriorityEncoder_v0p0p1_0.x22.Y 16to4_PriorityEncoder_v0p0p1_0.x22.A GND.t441 GND.t440 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1606 16to4_PriorityEncoder_v0p0p1_0.x3.x2.X a_77605_n48109# VDD.t746 VDD.t745 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.148 ps=1.34 w=1 l=0.15
X1607 GND.t1022 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t17 GND.t1021 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1608 a_77725_n50381# 16to4_PriorityEncoder_v0p0p1_0.x3.EI a_77639_n50381# GND.t1296 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X1609 VDD.t73 I13.t14 a_77637_n41087# VDD.t72 sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X1610 VDD.t475 frontAnalog_v0p0p1_4.x65.X frontAnalog_v0p0p1_4.RSfetsym_0.x2.Y VDD.t474 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1611 OUT1.t78 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD.t1366 VDD.t1365 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1612 VV9.t4 VV8.t5 GND.t78 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1613 VDD.t1466 16to4_PriorityEncoder_v0p0p1_0.x3.x22.A a_78775_n53555# VDD.t1465 sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X1614 OUT0.t75 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD.t822 VDD.t821 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1615 VDD.t1192 frontAnalog_v0p0p1_9.x65.A.t6 a_57123_n51159# VDD.t1191 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1616 GND.t1339 frontAnalog_v0p0p1_8.x63.A.t7 a_57123_n47279# GND.t1172 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X1617 VDD.t705 frontAnalog_v0p0p1_1.x65.X frontAnalog_v0p0p1_1.RSfetsym_0.x2.Y VDD.t704 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1618 frontAnalog_v0p0p1_0.RSfetsym_0.x2.Y frontAnalog_v0p0p1_0.x65.X VDD.t33 VDD.t31 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1619 frontAnalog_v0p0p1_6.x63.X a_57123_n31079# VDD.t686 VDD.t685 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1620 frontAnalog_v0p0p1_15.RSfetsym_0.x2.Y frontAnalog_v0p0p1_15.x65.X VDD.t194 VDD.t192 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1621 16to4_PriorityEncoder_v0p0p1_0.x42.A 16to4_PriorityEncoder_v0p0p1_0.x5.GS GND.t411 GND.t410 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1622 16to4_PriorityEncoder_v0p0p1_0.x29.A 16to4_PriorityEncoder_v0p0p1_0.x28.A GND.t1153 GND.t1152 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1623 w_55000_n46750# VIN.t27 a_53630_n47196# GND.t673 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1624 frontAnalog_v0p0p1_13.RSfetsym_0.x2.Y frontAnalog_v0p0p1_13.x65.X GND.t1203 GND.t1202 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1625 OUT0.t10 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND.t880 GND.t879 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1626 16to4_PriorityEncoder_v0p0p1_0.x22.Y 16to4_PriorityEncoder_v0p0p1_0.x22.A VDD.t427 VDD.t426 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1627 a_78241_n47345# 16to4_PriorityEncoder_v0p0p1_0.x3.x2.X a_78159_n47589# VDD.t191 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X1628 frontAnalog_v0p0p1_5.RSfetsym_0.QN.t2 frontAnalog_v0p0p1_5.x65.X VDD.t1310 VDD.t1309 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.25
X1629 frontAnalog_v0p0p1_11.x63.A.t2 frontAnalog_v0p0p1_11.x65.A.t7 a_55268_n63336# GND.t1118 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1630 OUT0.t9 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND.t878 GND.t877 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1631 GND.t876 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t8 GND.t875 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1632 GND.t439 16to4_PriorityEncoder_v0p0p1_0.x22.A 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND.t438 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1633 16to4_PriorityEncoder_v0p0p1_0.x3.x20.X a_77605_n53805# VDD.t1319 VDD.t1318 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X1634 a_77783_n48109# I6.t12 a_77687_n48109# VDD.t1258 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X1635 16to4_PriorityEncoder_v0p0p1_0.x1.A a_78349_n43045# GND.t1389 GND.t149 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.102 ps=0.99 w=0.65 l=0.15
X1636 I4.t4 frontAnalog_v0p0p1_11.RSfetsym_0.QN.t5 VDD.t1146 VDD.t414 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.3
X1637 a_77605_n48109# I5.t13 GND.t1134 GND.t20 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1638 GND.t1422 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t10 GND.t1421 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1639 GND.t787 16to4_PriorityEncoder_v0p0p1_0.x5.x14.A a_78065_n41309# GND.t786 sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X1640 VDD.t1364 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t77 VDD.t1363 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1641 OUT1.t76 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD.t1362 VDD.t1361 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1642 a_59577_n68283# frontAnalog_v0p0p1_13.x63.X I3.t1 GND.t378 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1643 a_59578_n78570# frontAnalog_v0p0p1_14.x65.X frontAnalog_v0p0p1_14.RSfetsym_0.QN.t2 GND.t1217 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.315 ps=2.72 w=1 l=0.15
X1644 GND.t1020 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t16 GND.t1019 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1645 VDD.t1360 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t75 VDD.t1359 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1646 I7.t4 frontAnalog_v0p0p1_8.RSfetsym_0.x2.Y GND.t1400 GND.t821 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.25
X1647 frontAnalog_v0p0p1_8.x63.A.t3 frontAnalog_v0p0p1_8.x65.A.t5 VDD.t204 VDD.t203 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1648 16to4_PriorityEncoder_v0p0p1_0.x5.x18.C I10.t11 VDD.t1212 VDD.t1211 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1649 OUT0.t74 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD.t820 VDD.t819 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1650 OUT2.t15 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND.t1018 GND.t1017 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1651 frontAnalog_v0p0p1_4.x63.A.t0 frontAnalog_v0p0p1_4.x65.A.t7 a_55268_n20136# GND.t1308 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1652 a_77759_n45765# 16to4_PriorityEncoder_v0p0p1_0.x5.x19.D a_77687_n45765# GND.t676 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X1653 VDD.t392 16to4_PriorityEncoder_v0p0p1_0.x5.A2 a_82988_n43855# VDD.t391 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X1654 frontAnalog_v0p0p1_1.x63.A.t2 CLK.t71 w_55000_n41350# VDD.t1088 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1655 OUT0.t73 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD.t818 VDD.t817 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1656 VDD.t816 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t72 VDD.t815 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1657 VDD.t425 16to4_PriorityEncoder_v0p0p1_0.x22.A 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD.t424 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1658 VDD.t79 frontAnalog_v0p0p1_10.x65.X frontAnalog_v0p0p1_10.RSfetsym_0.x2.Y VDD.t78 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1659 a_78649_n39527# 16to4_PriorityEncoder_v0p0p1_0.x5.EO VDD.t650 VDD.t649 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X1660 GND.t874 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t7 GND.t873 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1661 16to4_PriorityEncoder_v0p0p1_0.x1.A a_78349_n43045# VDD.t1327 VDD.t1326 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.148 ps=1.34 w=1 l=0.15
X1662 VDD.t770 R1.t7 a_57123_n79679# VDD.t769 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1663 a_78349_n43045# 16to4_PriorityEncoder_v0p0p1_0.x5.x22.A GND.t423 GND.t175 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1664 a_59577_n25083# frontAnalog_v0p0p1_5.x63.X I11.t0 GND.t25 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1665 a_59578_n35370# frontAnalog_v0p0p1_7.x65.X frontAnalog_v0p0p1_7.RSfetsym_0.QN.t2 GND.t1264 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.315 ps=2.72 w=1 l=0.15
X1666 VDD.t1081 CLK.t72 w_55000_n83928# GND.t593 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1667 I4.t2 frontAnalog_v0p0p1_11.x63.X VDD.t491 VDD.t490 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.25
X1668 a_53630_n74196# frontAnalog_v0p0p1_10.IB.t27 GND.t794 GND.t36 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1669 a_78775_n45515# 16to4_PriorityEncoder_v0p0p1_0.x5.x21.X a_78703_n45515# VDD.t1059 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X1670 VDD.t1254 frontAnalog_v0p0p1_13.x63.A.t7 frontAnalog_v0p0p1_13.x65.A.t0 VDD.t561 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1671 VDD.t1358 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t74 VDD.t1357 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1672 OUT1.t73 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD.t1356 VDD.t1355 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1673 GND.t872 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t6 GND.t871 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1674 OUT3.t9 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND.t235 GND.t234 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1675 OUT2.t14 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND.t1016 GND.t1015 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1676 VDD.t1082 CLK.t73 w_55000_n19128# GND.t733 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1677 frontAnalog_v0p0p1_15.x65.X a_57123_n83559# GND.t824 GND.t823 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1678 frontAnalog_v0p0p1_4.RSfetsym_0.QN.t3 frontAnalog_v0p0p1_4.RSfetsym_0.x1.Y GND.t655 GND.t654 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.25
X1679 16to4_PriorityEncoder_v0p0p1_0.x43.A 16to4_PriorityEncoder_v0p0p1_0.x42.A GND.t414 GND.t410 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1680 VDD.t539 frontAnalog_v0p0p1_3.x65.X frontAnalog_v0p0p1_3.RSfetsym_0.x2.Y VDD.t538 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1681 VV15.t12 VV14.t14 GND.t202 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1682 OUT3.t69 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD.t216 VDD.t215 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1683 VDD.t366 frontAnalog_v0p0p1_0.x63.X I14.t1 VDD.t365 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.25
X1684 VDD.t182 frontAnalog_v0p0p1_7.x63.A.t6 a_57123_n36479# VDD.t181 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1685 a_53630_n79596# VV2.t17 w_55000_n78528# GND.t854 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1686 VDD.t1083 CLK.t74 w_55000_n40728# GND.t1158 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1687 I12.t1 frontAnalog_v0p0p1_4.x63.X VDD.t118 VDD.t117 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.25
X1688 VFS.t1 VV16.t4 GND.t123 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1689 VDD.t948 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t74 VDD.t947 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1690 VDD.t814 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t71 VDD.t813 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1691 a_77687_n53805# I5.t14 a_77605_n53805# GND.t1135 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X1692 VDD.t406 frontAnalog_v0p0p1_5.x63.A.t7 frontAnalog_v0p0p1_5.x65.A.t3 VDD.t405 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1693 VV4.t10 VV3.t10 GND.t24 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1694 frontAnalog_v0p0p1_9.RSfetsym_0.x2.Y frontAnalog_v0p0p1_9.x65.X GND.t1328 GND.t1327 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1695 a_55268_n57936# CLK.t75 GND.t1160 GND.t1159 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1696 VDD.t193 frontAnalog_v0p0p1_15.x65.X frontAnalog_v0p0p1_15.RSfetsym_0.x2.Y VDD.t192 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1697 VDD.t1084 CLK.t76 w_55000_n41350# GND.t1161 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1698 frontAnalog_v0p0p1_6.x65.A.t2 frontAnalog_v0p0p1_6.x63.A.t7 a_55268_n30936# GND.t1187 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1699 frontAnalog_v0p0p1_11.RSfetsym_0.QN.t0 I4.t12 VDD.t415 VDD.t414 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.3
X1700 VDD.t812 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t70 VDD.t811 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1701 GND.t1543 16to4_PriorityEncoder_v0p0p1_0.x36.A 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND.t1542 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1702 frontAnalog_v0p0p1_1.x65.X a_57123_n40359# GND.t1340 GND.t347 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1703 VDD.t756 I12.t11 a_77637_n40777# VDD.t755 sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X1704 16to4_PriorityEncoder_v0p0p1_0.x22.A 16to4_PriorityEncoder_v0p0p1_0.x21.A GND.t1349 GND.t1348 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1705 a_78649_n47567# 16to4_PriorityEncoder_v0p0p1_0.x3.EO VDD.t90 VDD.t89 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X1706 a_53630_n36396# VV10.t17 w_55000_n35328# GND.t127 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1707 16to4_PriorityEncoder_v0p0p1_0.x3.A1 a_78349_n51085# VDD.t1283 VDD.t1282 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.148 ps=1.34 w=1 l=0.15
X1708 GND.t413 16to4_PriorityEncoder_v0p0p1_0.x42.A 16to4_PriorityEncoder_v0p0p1_0.x43.A GND.t412 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1709 OUT2.t13 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND.t1014 GND.t1013 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1710 16to4_PriorityEncoder_v0p0p1_0.x3.x22.A a_77639_n50381# VDD.t385 VDD.t384 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.167 ps=1.39 w=1 l=0.15
X1711 a_78775_n53555# 16to4_PriorityEncoder_v0p0p1_0.x3.x21.X a_78703_n53555# VDD.t695 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X1712 frontAnalog_v0p0p1_11.RSfetsym_0.x2.Y frontAnalog_v0p0p1_11.x65.X VDD.t722 VDD.t720 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1713 frontAnalog_v0p0p1_2.RSfetsym_0.x1.Y frontAnalog_v0p0p1_2.x63.X VDD.t41 VDD.t39 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1714 VV11.t9 VV10.t8 GND.t52 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1715 a_55268_n14736# CLK.t77 GND.t1163 GND.t1162 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1716 frontAnalog_v0p0p1_11.RSfetsym_0.x1.Y frontAnalog_v0p0p1_11.x63.X GND.t508 GND.t506 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1717 frontAnalog_v0p0p1_13.RSfetsym_0.QN.t2 frontAnalog_v0p0p1_13.x65.X VDD.t1113 VDD.t1112 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.25
X1718 OUT2.t12 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND.t1012 GND.t1011 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1719 VDD.t214 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t68 VDD.t213 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1720 OUT1.t72 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD.t1354 VDD.t1353 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1721 GND.t233 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t8 GND.t232 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1722 GND.t1010 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t11 GND.t1009 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1723 VDD.t1122 frontAnalog_v0p0p1_14.x65.X frontAnalog_v0p0p1_14.RSfetsym_0.QN.t3 VDD.t1121 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.25
X1724 OUT3.t67 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD.t212 VDD.t211 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1725 GND.t870 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t5 GND.t869 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1726 a_77637_n49127# 16to4_PriorityEncoder_v0p0p1_0.x3.EI VDD.t1236 VDD.t698 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X1727 frontAnalog_v0p0p1_0.x65.A.t1 CLK.t78 frontAnalog_v0p0p1_0.x63.A.t0 VDD.t1085 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1728 VV7.t2 VV6.t5 GND.t51 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1729 VDD.t210 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t66 VDD.t209 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1730 16to4_PriorityEncoder_v0p0p1_0.x22.A 16to4_PriorityEncoder_v0p0p1_0.x21.A VDD.t1290 VDD.t1289 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1731 frontAnalog_v0p0p1_12.RSfetsym_0.x1.Y frontAnalog_v0p0p1_12.x63.X VDD.t113 VDD.t109 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1732 GND.t1373 frontAnalog_v0p0p1_5.x65.X frontAnalog_v0p0p1_5.RSfetsym_0.x2.Y GND.t1372 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1733 a_77687_n48109# I7.t8 a_77605_n48109# VDD.t1253 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X1734 GND.t354 frontAnalog_v0p0p1_14.x63.X frontAnalog_v0p0p1_14.RSfetsym_0.x1.Y GND.t353 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1735 VIN.t28 w_55000_n46128# error sky130_fd_pr__cap_var_lvt w=2 l=0.18
X1736 GND.t1008 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t10 GND.t1007 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1737 OUT2.t73 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD.t946 VDD.t945 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1738 frontAnalog_v0p0p1_2.x65.X a_57123_n2559# VDD.t383 VDD.t382 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1739 a_16719_n13117.t7 a_16599_n13205.t20 a_16541_n13117.t11 GND.t833 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1740 a_53630_n84996# frontAnalog_v0p0p1_10.IB.t28 GND.t529 GND.t36 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1741 VDD.t1195 frontAnalog_v0p0p1_7.x65.X frontAnalog_v0p0p1_7.RSfetsym_0.QN.t3 VDD.t1194 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.25
X1742 a_16719_n13117.t6 a_16599_n13205.t21 a_16541_n13117.t10 GND.t834 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1743 OUT1.t9 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND.t1420 GND.t1419 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1744 VDD.t944 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t72 VDD.t943 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1745 VDD.t810 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t69 VDD.t809 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1746 16to4_PriorityEncoder_v0p0p1_0.x3.x11.X a_77637_n49127# VDD.t1278 VDD.t45 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.167 ps=1.39 w=1 l=0.15
X1747 frontAnalog_v0p0p1_6.RSfetsym_0.x1.Y frontAnalog_v0p0p1_6.x63.X VDD.t592 VDD.t588 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1748 GND.t1418 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t8 GND.t1417 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1749 frontAnalog_v0p0p1_8.x65.A.t1 CLK.t79 frontAnalog_v0p0p1_8.x63.A.t0 VDD.t667 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1750 a_77605_n43545# 16to4_PriorityEncoder_v0p0p1_0.x5.x16.C VDD.t765 VDD.t741 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X1751 frontAnalog_v0p0p1_3.x63.X a_57123_n14879# VDD.t75 VDD.t74 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1752 frontAnalog_v0p0p1_13.RSfetsym_0.x2.Y frontAnalog_v0p0p1_13.x65.X VDD.t1111 VDD.t1109 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1753 frontAnalog_v0p0p1_0.RSfetsym_0.x1.Y frontAnalog_v0p0p1_0.x63.X VDD.t364 VDD.t362 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1754 a_53630_n20196# frontAnalog_v0p0p1_10.IB.t29 GND.t530 GND.t36 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1755 w_55000_n30550# VIN.t29 a_53630_n30996# GND.t408 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1756 GND.t578 frontAnalog_v0p0p1_7.x63.X frontAnalog_v0p0p1_7.RSfetsym_0.x1.Y GND.t577 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1757 VV6.t14 VV5.t12 GND.t52 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1758 VDD.t61 16to4_PriorityEncoder_v0p0p1_0.x35.A 16to4_PriorityEncoder_v0p0p1_0.x36.A VDD.t60 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1759 GND.t231 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t7 GND.t230 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1760 GND.t621 frontAnalog_v0p0p1_0.x63.A.t6 a_57123_n9479# GND.t87 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X1761 frontAnalog_v0p0p1_12.x65.X a_57123_n72759# VDD.t603 VDD.t602 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1762 frontAnalog_v0p0p1_13.x63.X a_57123_n68879# GND.t108 GND.t107 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1763 GND.t1541 16to4_PriorityEncoder_v0p0p1_0.x36.A 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND.t1540 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1764 a_53630_n9396# VV15.t17 w_55000_n8328# GND.t818 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1765 a_53630_n41796# frontAnalog_v0p0p1_10.IB.t30 GND.t531 GND.t36 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1766 frontAnalog_v0p0p1_11.x63.A.t0 CLK.t80 w_55000_n62950# VDD.t668 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1767 16to4_PriorityEncoder_v0p0p1_0.x5.x1.X a_77605_n39305# GND.t74 GND.t73 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.102 ps=0.99 w=0.65 l=0.15
X1768 VV14.t8 VV13.t7 GND.t52 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1769 GND.t1173 frontAnalog_v0p0p1_8.x65.A.t6 a_57123_n45759# GND.t1172 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X1770 VV5.t10 VV4.t11 GND.t33 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1771 OUT3.t6 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND.t229 GND.t228 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1772 frontAnalog_v0p0p1_15.RSfetsym_0.QN.t3 frontAnalog_v0p0p1_15.RSfetsym_0.x1.Y GND.t1371 GND.t436 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.25
X1773 OUT2.t71 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD.t942 VDD.t941 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1774 VDD.t940 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t70 VDD.t939 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1775 GND.t1326 frontAnalog_v0p0p1_9.x65.X frontAnalog_v0p0p1_9.RSfetsym_0.x2.Y GND.t1325 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1776 GND.t629 16to4_PriorityEncoder_v0p0p1_0.x43.A 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND.t628 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1777 I7.t0 frontAnalog_v0p0p1_8.RSfetsym_0.QN.t6 VDD.t666 VDD.t665 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.3
X1778 frontAnalog_v0p0p1_5.RSfetsym_0.x2.Y frontAnalog_v0p0p1_5.x65.X VDD.t1308 VDD.t1306 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1779 VDD.t669 CLK.t81 w_55000_n84550# GND.t684 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1780 VDD.t760 frontAnalog_v0p0p1_8.x63.X frontAnalog_v0p0p1_8.RSfetsym_0.x1.Y VDD.t759 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1781 VDD.t112 frontAnalog_v0p0p1_12.x63.X I2.t1 VDD.t111 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.25
X1782 w_55000_n73128# CLK.t82 frontAnalog_v0p0p1_12.x65.A.t3 VDD.t670 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1783 frontAnalog_v0p0p1_5.x63.X a_57123_n25679# GND.t759 GND.t480 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1784 GND.t1130 frontAnalog_v0p0p1_10.IB.t1 frontAnalog_v0p0p1_10.IB.t2 GND.t1129 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1785 VV8.t17 w_55000_n46750# error sky130_fd_pr__cap_var_lvt w=2 l=0.18
X1786 GND.t1006 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t9 GND.t1005 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1787 frontAnalog_v0p0p1_1.RSfetsym_0.QN.t0 frontAnalog_v0p0p1_1.RSfetsym_0.x1.Y GND.t184 GND.t183 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.25
X1788 16to4_PriorityEncoder_v0p0p1_0.x5.x1.X a_77605_n39305# VDD.t57 VDD.t56 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.148 ps=1.34 w=1 l=0.15
X1789 OUT3.t5 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND.t227 GND.t226 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1790 16to4_PriorityEncoder_v0p0p1_0.x2.A a_78525_n45515# GND.t773 GND.t772 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.102 ps=0.99 w=0.65 l=0.15
X1791 16to4_PriorityEncoder_v0p0p1_0.x36.Y 16to4_PriorityEncoder_v0p0p1_0.x36.A GND.t1539 GND.t1538 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1792 VDD.t208 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t65 VDD.t207 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1793 GND.t507 frontAnalog_v0p0p1_11.x63.X frontAnalog_v0p0p1_11.RSfetsym_0.x1.Y GND.t506 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1794 GND.t1416 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t7 GND.t1415 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1795 16to4_PriorityEncoder_v0p0p1_0.x36.Y 16to4_PriorityEncoder_v0p0p1_0.x36.A VDD.t1473 VDD.t1472 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1796 VDD.t591 frontAnalog_v0p0p1_6.x63.X I10.t1 VDD.t590 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.25
X1797 a_77605_n51585# 16to4_PriorityEncoder_v0p0p1_0.x3.x16.C VDD.t335 VDD.t176 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X1798 w_55000_n29928# CLK.t83 frontAnalog_v0p0p1_6.x65.A.t0 VDD.t76 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1799 frontAnalog_v0p0p1_4.RSfetsym_0.x1.Y frontAnalog_v0p0p1_4.x63.X GND.t136 GND.t134 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1800 a_53630_n57996# frontAnalog_v0p0p1_10.IB.t31 GND.t532 GND.t36 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1801 a_55268_n79536# CLK.t84 GND.t686 GND.t685 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1802 frontAnalog_v0p0p1_9.x65.A.t0 frontAnalog_v0p0p1_9.x63.A.t6 a_55268_n52536# GND.t1240 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1803 16to4_PriorityEncoder_v0p0p1_0.x43.Y 16to4_PriorityEncoder_v0p0p1_0.x43.A GND.t627 GND.t626 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1804 16to4_PriorityEncoder_v0p0p1_0.x3.x1.X a_77605_n47345# GND.t669 GND.t668 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.102 ps=0.99 w=0.65 l=0.15
X1805 VV11.t15 VV10.t12 GND.t202 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1806 VDD.t110 frontAnalog_v0p0p1_12.x63.X frontAnalog_v0p0p1_12.RSfetsym_0.x1.Y VDD.t109 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1807 GND.t1414 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t6 GND.t1413 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1808 frontAnalog_v0p0p1_0.RSfetsym_0.QN.t4 frontAnalog_v0p0p1_0.RSfetsym_0.x1.Y GND.t375 GND.t374 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.25
X1809 VDD.t32 frontAnalog_v0p0p1_0.x65.X frontAnalog_v0p0p1_0.RSfetsym_0.x2.Y VDD.t31 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1810 16to4_PriorityEncoder_v0p0p1_0.x3.x16.X a_77605_n51585# GND.t1277 GND.t1276 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.196 ps=1.33 w=0.65 l=0.15
X1811 GND.t225 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t4 GND.t224 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1812 GND.t88 frontAnalog_v0p0p1_0.x65.A.t6 a_57123_n7959# GND.t87 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X1813 GND.t1243 frontAnalog_v0p0p1_11.RSfetsym_0.QN.t6 a_59577_n62883# GND.t1242 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1814 GND.t1201 frontAnalog_v0p0p1_13.x65.X frontAnalog_v0p0p1_13.RSfetsym_0.x2.Y GND.t1200 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1815 16to4_PriorityEncoder_v0p0p1_0.x2.A a_78525_n45515# VDD.t730 VDD.t729 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.148 ps=1.34 w=1 l=0.15
X1816 OUT2.t69 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD.t938 VDD.t937 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1817 a_78525_n45515# 16to4_PriorityEncoder_v0p0p1_0.x5.x21.X GND.t1132 GND.t1131 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1818 VDD.t611 frontAnalog_v0p0p1_0.x63.A.t7 frontAnalog_v0p0p1_0.x65.A.t2 VDD.t574 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1819 16to4_PriorityEncoder_v0p0p1_0.x5.x21.X a_78097_n45737# GND.t65 GND.t64 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.112 ps=1.04 w=0.65 l=0.15
X1820 VDD.t1471 16to4_PriorityEncoder_v0p0p1_0.x36.A 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD.t1470 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1821 a_53630_n14796# frontAnalog_v0p0p1_10.IB.t32 GND.t533 GND.t36 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1822 a_77637_n48817# 16to4_PriorityEncoder_v0p0p1_0.x3.EI VDD.t1235 VDD.t1234 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X1823 16to4_PriorityEncoder_v0p0p1_0.x5.x19.C I12.t12 VDD.t1323 VDD.t1322 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1824 frontAnalog_v0p0p1_9.RSfetsym_0.x1.Y frontAnalog_v0p0p1_9.x63.X VDD.t1098 VDD.t1097 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1825 VDD.t584 S1.t7 a_57123_n78159# VDD.t583 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1826 VDD.t1074 16to4_PriorityEncoder_v0p0p1_0.x28.A 16to4_PriorityEncoder_v0p0p1_0.x29.A VDD.t1073 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1827 VDD.t589 frontAnalog_v0p0p1_6.x63.X frontAnalog_v0p0p1_6.RSfetsym_0.x1.Y VDD.t588 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1828 OUT0.t4 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND.t868 GND.t867 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1829 OUT2.t8 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND.t1004 GND.t1003 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1830 I15.t3 frontAnalog_v0p0p1_2.RSfetsym_0.QN.t6 VDD.t773 VDD.t753 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.3
X1831 VDD.t1110 frontAnalog_v0p0p1_13.x65.X frontAnalog_v0p0p1_13.RSfetsym_0.x2.Y VDD.t1109 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1832 VDD.t363 frontAnalog_v0p0p1_0.x63.X frontAnalog_v0p0p1_0.RSfetsym_0.x1.Y VDD.t362 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1833 frontAnalog_v0p0p1_10.x63.X a_57123_n58079# VDD.t656 VDD.t655 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1834 16to4_PriorityEncoder_v0p0p1_0.x3.x1.X a_77605_n47345# VDD.t654 VDD.t653 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.148 ps=1.34 w=1 l=0.15
X1835 GND.t223 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t3 GND.t222 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1836 GND.t866 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t3 GND.t865 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1837 OUT1.t5 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND.t1412 GND.t1411 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1838 a_77775_n43545# 16to4_PriorityEncoder_v0p0p1_0.x5.x19.C a_77687_n43545# GND.t699 sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
X1839 16to4_PriorityEncoder_v0p0p1_0.x43.A 16to4_PriorityEncoder_v0p0p1_0.x42.A VDD.t396 VDD.t395 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1840 OUT1.t71 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD.t1352 VDD.t1351 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1841 frontAnalog_v0p0p1_2.RSfetsym_0.x2.Y frontAnalog_v0p0p1_2.x65.X GND.t1287 GND.t1286 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1842 VDD.t936 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t68 VDD.t935 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1843 VDD.t1154 VDD.t1152 a_77605_n45765# VDD.t1153 sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X1844 16to4_PriorityEncoder_v0p0p1_0.x5.x21.X a_78097_n45737# VDD.t49 VDD.t48 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.167 ps=1.39 w=1 l=0.15
X1845 VDD.t1303 frontAnalog_v0p0p1_7.x65.A.t7 a_57123_n34959# VDD.t1302 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1846 VDD.t1307 frontAnalog_v0p0p1_5.x65.X frontAnalog_v0p0p1_5.RSfetsym_0.x2.Y VDD.t1306 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1847 VV16.t15 VV15.t15 GND.t106 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1848 VV6.t4 VV5.t4 GND.t202 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1849 VV5.t0 VV4.t1 GND.t78 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1850 OUT2.t7 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND.t1002 GND.t1001 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1851 OUT0.t68 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD.t808 VDD.t807 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1852 16to4_PriorityEncoder_v0p0p1_0.x3.A0 a_78525_n53555# VDD.t1108 VDD.t1107 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.148 ps=1.34 w=1 l=0.15
X1853 GND.t1000 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t6 GND.t999 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1854 a_78431_n43045# 16to4_PriorityEncoder_v0p0p1_0.x5.x16.X a_78349_n43045# VDD.t798 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X1855 VV14.t9 VV13.t10 GND.t202 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1856 GND.t707 VDD.t1511 a_77759_n45765# GND.t706 sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X1857 VDD.t934 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t67 VDD.t933 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1858 a_78525_n53555# 16to4_PriorityEncoder_v0p0p1_0.x3.x21.X GND.t737 GND.t736 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1859 VDD.t806 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t67 VDD.t805 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1860 a_77687_n52819# 16to4_PriorityEncoder_v0p0p1_0.x3.EI a_77605_n52819# GND.t185 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.109 ps=1.36 w=0.42 l=0.15
X1861 w_55000_n52150# VIN.t30 a_53630_n52596# GND.t1148 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1862 frontAnalog_v0p0p1_12.RSfetsym_0.x2.Y frontAnalog_v0p0p1_12.x65.X GND.t192 GND.t191 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1863 frontAnalog_v0p0p1_0.RSfetsym_0.QN.t0 frontAnalog_v0p0p1_0.x65.X VDD.t30 VDD.t29 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.25
X1864 GND.t152 16to4_PriorityEncoder_v0p0p1_0.x5.x4.A a_78159_n39549# GND.t151 sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X1865 frontAnalog_v0p0p1_2.x63.A.t3 frontAnalog_v0p0p1_2.x65.A.t7 VDD.t612 VDD.t420 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1866 VDD.t671 CLK.t85 w_55000_n2928# GND.t687 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1867 frontAnalog_v0p0p1_8.x63.A.t2 frontAnalog_v0p0p1_8.x65.A.t7 a_55268_n47136# GND.t1174 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1868 VV12.t11 VV11.t11 GND.t422 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1869 GND.t864 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t2 GND.t863 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1870 a_77775_n51585# 16to4_PriorityEncoder_v0p0p1_0.x3.x19.C a_77687_n51585# GND.t174 sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
X1871 16to4_PriorityEncoder_v0p0p1_0.x5.x14.A a_77637_n40777# GND.t1222 GND.t68 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.112 ps=1.04 w=0.65 l=0.15
X1872 VDD.t932 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t66 VDD.t931 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1873 frontAnalog_v0p0p1_6.RSfetsym_0.x2.Y frontAnalog_v0p0p1_6.x65.X GND.t5 GND.t4 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1874 frontAnalog_v0p0p1_15.RSfetsym_0.x1.Y frontAnalog_v0p0p1_15.x63.X GND.t498 GND.t497 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1875 OUT1.t70 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD.t1350 VDD.t1349 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1876 a_59577_n8883# frontAnalog_v0p0p1_0.x63.X I14.t0 GND.t368 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1877 frontAnalog_v0p0p1_3.RSfetsym_0.x1.Y frontAnalog_v0p0p1_3.x63.X VDD.t468 VDD.t464 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1878 w_55000_n8328# CLK.t86 frontAnalog_v0p0p1_0.x65.A.t0 VDD.t148 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1879 a_59577_n73683# frontAnalog_v0p0p1_12.x63.X I2.t0 GND.t128 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1880 a_59578_n83970# frontAnalog_v0p0p1_15.x65.X frontAnalog_v0p0p1_15.RSfetsym_0.QN.t2 GND.t205 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.315 ps=2.72 w=1 l=0.15
X1881 VDD.t1233 16to4_PriorityEncoder_v0p0p1_0.x3.EI a_77605_n53805# VDD.t1232 sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X1882 16to4_PriorityEncoder_v0p0p1_0.x3.x21.X a_78097_n53777# VDD.t162 VDD.t161 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.167 ps=1.39 w=1 l=0.15
X1883 OUT2.t65 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD.t930 VDD.t929 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1884 I6.t4 frontAnalog_v0p0p1_9.RSfetsym_0.x2.Y GND.t1334 GND.t31 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.25
X1885 GND.t165 16to4_PriorityEncoder_v0p0p1_0.x1.A a_82906_n47995# GND.t164 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X1886 frontAnalog_v0p0p1_2.RSfetsym_0.QN.t1 I15.t8 VDD.t754 VDD.t753 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.3
X1887 GND.t862 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t1 GND.t861 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1888 VV12.t3 VV11.t2 GND.t214 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1889 VV8.t12 VV7.t14 GND.t33 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1890 VV15.t4 VV14.t3 GND.t24 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1891 GND.t221 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t2 GND.t220 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1892 a_78183_n45737# VDD.t1512 a_78097_n45737# GND.t708 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X1893 VDD.t1089 CLK.t87 w_55000_n67728# GND.t435 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1894 a_59578_n19170# frontAnalog_v0p0p1_4.x65.X frontAnalog_v0p0p1_4.RSfetsym_0.QN.t0 GND.t488 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.315 ps=2.72 w=1 l=0.15
X1895 VDD.t804 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t66 VDD.t803 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1896 a_77881_n51335# 16to4_PriorityEncoder_v0p0p1_0.x3.x16.C a_77775_n51335# GND.t346 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X1897 I7.t2 frontAnalog_v0p0p1_8.x63.X VDD.t758 VDD.t757 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.25
X1898 VDD.t721 frontAnalog_v0p0p1_11.x65.X frontAnalog_v0p0p1_11.RSfetsym_0.x2.Y VDD.t720 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1899 a_78431_n51085# 16to4_PriorityEncoder_v0p0p1_0.x3.x16.X a_78349_n51085# VDD.t200 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X1900 VDD.t40 frontAnalog_v0p0p1_2.x63.X frontAnalog_v0p0p1_2.RSfetsym_0.x1.Y VDD.t39 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1901 OUT2.t5 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND.t998 GND.t997 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1902 frontAnalog_v0p0p1_1.RSfetsym_0.x1.Y frontAnalog_v0p0p1_1.x63.X GND.t178 GND.t177 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1903 frontAnalog_v0p0p1_14.RSfetsym_0.x2.Y frontAnalog_v0p0p1_14.x65.X GND.t1216 GND.t1215 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1904 OUT1.t69 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD.t1348 VDD.t1347 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1905 16to4_PriorityEncoder_v0p0p1_0.x36.Y 16to4_PriorityEncoder_v0p0p1_0.x36.A VDD.t1469 VDD.t1468 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1906 a_59577_n30483# frontAnalog_v0p0p1_6.x63.X I10.t3 GND.t611 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1907 a_59578_n40770# frontAnalog_v0p0p1_1.x65.X frontAnalog_v0p0p1_1.RSfetsym_0.QN.t1 GND.t748 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.315 ps=2.72 w=1 l=0.15
X1908 VDD.t1090 CLK.t88 w_55000_n68350# GND.t160 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1909 GND.t1273 16to4_PriorityEncoder_v0p0p1_0.x3.x19.D a_77881_n52819# GND.t185 sky130_fd_pr__nfet_01v8 ad=0.196 pd=1.33 as=0.0693 ps=0.75 w=0.42 l=0.15
X1910 VDD.t744 16to4_PriorityEncoder_v0p0p1_0.x5.x14.A a_78315_n41309# VDD.t410 sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X1911 GND.t116 16to4_PriorityEncoder_v0p0p1_0.x3.x4.A a_78159_n47589# GND.t115 sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X1912 GND.t996 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t4 GND.t995 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1913 VDD.t751 frontAnalog_v0p0p1_12.x63.A.t7 frontAnalog_v0p0p1_12.x65.A.t1 VDD.t750 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1914 frontAnalog_v0p0p1_2.x63.A.t1 CLK.t89 w_55000_n3550# VDD.t355 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1915 frontAnalog_v0p0p1_13.x65.X a_57123_n67359# GND.t1272 GND.t107 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1916 GND.t1184 I2.t12 a_59578_n73170# GND.t1183 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1917 VV16.t2 VV15.t6 GND.t77 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1918 VDD.t802 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t65 VDD.t801 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1919 I15.t1 frontAnalog_v0p0p1_2.x63.X VDD.t38 VDD.t37 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.25
X1920 GND.t1285 frontAnalog_v0p0p1_2.x65.X frontAnalog_v0p0p1_2.RSfetsym_0.x2.Y GND.t1284 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1921 VDD.t1091 CLK.t90 w_55000_n24528# GND.t587 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1922 OUT0.t0 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND.t860 GND.t859 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1923 GND.t1410 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t4 GND.t1409 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1924 16to4_PriorityEncoder_v0p0p1_0.x29.Y 16to4_PriorityEncoder_v0p0p1_0.x29.A VDD.t509 VDD.t508 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1925 frontAnalog_v0p0p1_7.RSfetsym_0.x2.Y frontAnalog_v0p0p1_7.x65.X GND.t1263 GND.t1262 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1926 VDD.t713 frontAnalog_v0p0p1_1.x63.A.t7 a_57123_n41879# VDD.t712 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1927 GND.t1537 16to4_PriorityEncoder_v0p0p1_0.x36.A 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND.t1536 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1928 VDD.t467 frontAnalog_v0p0p1_3.x63.X I13.t2 VDD.t466 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.25
X1929 VDD.t1092 CLK.t91 w_55000_n25150# GND.t595 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1930 16to4_PriorityEncoder_v0p0p1_0.x3.A2 a_78065_n49349# GND.t61 GND.t60 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.102 ps=0.99 w=0.65 l=0.15
X1931 w_55000_n13728# CLK.t92 frontAnalog_v0p0p1_3.x65.A.t0 VDD.t676 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1932 frontAnalog_v0p0p1_8.RSfetsym_0.QN.t1 I7.t9 VDD.t1067 VDD.t665 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.3
X1933 GND.t994 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t3 GND.t993 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1934 frontAnalog_v0p0p1_5.x65.X a_57123_n24159# GND.t481 GND.t480 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1935 GND.t516 I15.t9 a_77725_n42341# GND.t515 sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X1936 frontAnalog_v0p0p1_7.x65.A.t1 frontAnalog_v0p0p1_7.x63.A.t7 a_55268_n36336# GND.t186 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1937 a_53630_n20196# VV13.t17 w_55000_n19128# GND.t743 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1938 a_78183_n53777# 16to4_PriorityEncoder_v0p0p1_0.x3.EI a_78097_n53777# GND.t1295 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X1939 OUT2.t64 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD.t928 VDD.t927 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1940 OUT0.t64 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD.t800 VDD.t799 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1941 frontAnalog_v0p0p1_8.RSfetsym_0.x2.Y frontAnalog_v0p0p1_8.x65.X VDD.t1330 VDD.t1329 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1942 OUT1.t68 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD.t1346 VDD.t1345 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1943 frontAnalog_v0p0p1_8.RSfetsym_0.x1.Y frontAnalog_v0p0p1_8.x63.X GND.t810 GND.t809 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1944 16to4_PriorityEncoder_v0p0p1_0.x35.A 16to4_PriorityEncoder_v0p0p1_0.x34.A VDD.t51 VDD.t50 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1945 GND.t625 16to4_PriorityEncoder_v0p0p1_0.x43.A 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND.t624 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1946 GND.t992 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t2 GND.t991 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1947 VDD.t738 16to4_PriorityEncoder_v0p0p1_0.x5.x19.C a_77605_n43295# VDD.t737 sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X1948 frontAnalog_v0p0p1_0.x63.A.t2 frontAnalog_v0p0p1_0.x65.A.t7 a_55268_n9336# GND.t89 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1949 OUT1.t67 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD.t1344 VDD.t1343 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1950 VDD.t1342 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t66 VDD.t1341 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1951 VDD.t507 16to4_PriorityEncoder_v0p0p1_0.x29.A 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD.t506 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1952 GND.t518 I15.t10 a_59578_n2970# GND.t517 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1953 GND.t1241 frontAnalog_v0p0p1_9.x63.A.t7 a_57123_n52679# GND.t690 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X1954 a_55268_n20136# CLK.t93 GND.t831 GND.t830 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1955 frontAnalog_v0p0p1_12.RSfetsym_0.QN.t1 frontAnalog_v0p0p1_12.x65.X VDD.t184 VDD.t183 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.25
X1956 16to4_PriorityEncoder_v0p0p1_0.x36.Y 16to4_PriorityEncoder_v0p0p1_0.x36.A GND.t1535 GND.t1534 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1957 a_16719_n13117.t5 a_16599_n13205.t22 a_16541_n13117.t9 GND.t835 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1958 VDD.t206 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t64 VDD.t205 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1959 16to4_PriorityEncoder_v0p0p1_0.x3.x4.A 16to4_PriorityEncoder_v0p0p1_0.x3.EI GND.t1294 GND.t1293 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1960 VDD.t465 frontAnalog_v0p0p1_3.x63.X frontAnalog_v0p0p1_3.RSfetsym_0.x1.Y VDD.t464 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1961 frontAnalog_v0p0p1_10.RSfetsym_0.x1.Y frontAnalog_v0p0p1_10.x63.X VDD.t784 VDD.t783 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1962 VV12.t8 VV11.t7 GND.t394 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1963 VIN.t31 w_55000_n29928# error sky130_fd_pr__cap_var_lvt w=2 l=0.18
X1964 GND.t576 16to4_PriorityEncoder_v0p0p1_0.x2.A a_82906_n51645# GND.t575 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X1965 OUT1.t3 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND.t1408 GND.t1407 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1966 VDD.t779 CLK.t94 w_55000_n3550# GND.t596 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1967 VDD.t473 frontAnalog_v0p0p1_4.x65.X frontAnalog_v0p0p1_4.RSfetsym_0.QN.t1 VDD.t472 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.25
X1968 a_53630_n68796# frontAnalog_v0p0p1_10.IB.t33 GND.t472 GND.t36 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1969 OUT3.t1 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND.t219 GND.t218 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1970 VV8.t9 VV7.t11 GND.t78 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1971 OUT2.t1 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND.t990 GND.t989 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1972 GND.t1139 I7.t10 a_77725_n50381# GND.t1138 sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X1973 GND.t1406 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t2 GND.t1405 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1974 a_82906_n47995# 16to4_PriorityEncoder_v0p0p1_0.x3.A1 GND.t63 GND.t62 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1975 VDD.t1340 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t65 VDD.t1339 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1976 16to4_PriorityEncoder_v0p0p1_0.x34.A a_82906_n43855# GND.t1120 GND.t1119 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1 ps=0.985 w=0.65 l=0.15
X1977 frontAnalog_v0p0p1_2.x63.X a_57123_n4079# GND.t1185 GND.t395 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1978 GND.t1214 frontAnalog_v0p0p1_14.x65.X frontAnalog_v0p0p1_14.RSfetsym_0.x2.Y GND.t1213 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1979 GND.t1387 16to4_PriorityEncoder_v0p0p1_0.x5.x17.A a_78065_n41309# GND.t1386 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X1980 GND.t523 I8.t8 a_77605_n39305# GND.t140 sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X1981 GND.t135 frontAnalog_v0p0p1_4.x63.X frontAnalog_v0p0p1_4.RSfetsym_0.x1.Y GND.t134 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1982 frontAnalog_v0p0p1_9.x63.A.t3 frontAnalog_v0p0p1_9.x65.A.t7 VDD.t1193 VDD.t556 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1983 GND.t1151 16to4_PriorityEncoder_v0p0p1_0.x28.A 16to4_PriorityEncoder_v0p0p1_0.x29.A GND.t1150 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1984 VDD.t1338 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t64 VDD.t1337 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1985 frontAnalog_v0p0p1_10.x65.X a_57123_n56559# VDD.t59 VDD.t58 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1986 OUT3.t0 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND.t217 GND.t216 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1987 VDD.t606 16to4_PriorityEncoder_v0p0p1_0.x3.x19.C a_77605_n51335# VDD.t605 sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X1988 a_53630_n25596# frontAnalog_v0p0p1_10.IB.t34 GND.t473 GND.t36 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1989 OUT2.t0 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND.t988 GND.t987 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1990 a_77605_n43295# I10.t12 VDD.t1214 VDD.t1213 sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.109 ps=1.36 w=0.42 l=0.15
X1991 frontAnalog_v0p0p1_8.x63.A.t1 CLK.t95 w_55000_n46750# VDD.t596 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1992 GND.t431 frontAnalog_v0p0p1_6.x65.A.t7 a_57123_n29559# GND.t430 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X1993 VDD.t547 16to4_PriorityEncoder_v0p0p1_0.x2.A a_82988_n51645# VDD.t546 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X1994 a_16719_n13117.t4 a_16599_n13205.t23 a_16541_n13117.t8 GND.t836 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1995 frontAnalog_v0p0p1_13.RSfetsym_0.QN.t4 frontAnalog_v0p0p1_13.RSfetsym_0.x1.Y GND.t1212 GND.t156 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.25
X1996 GND.t623 16to4_PriorityEncoder_v0p0p1_0.x43.A 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND.t622 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1997 frontAnalog_v0p0p1_12.x63.X a_57123_n74279# GND.t1261 GND.t619 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1998 OUT1.t1 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND.t1404 GND.t1403 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1999 GND.t1402 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t0 GND.t1401 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
R0 GND.n6877 GND.n6876 5.63094e+06
R1 GND.n6798 GND 2.276e+06
R2 GND.n6798 GND 2.00869e+06
R3 GND GND.n5220 334900
R4 GND.n6874 GND 334900
R5 GND.n4916 GND.n4915 273240
R6 GND GND.n6794 271091
R7 GND.n4915 GND 271091
R8 GND.n5220 GND.n5177 215600
R9 GND.n6875 GND.n6874 215600
R10 GND GND.n7429 122896
R11 GND.n1329 GND.n1328 98120
R12 GND.n3587 GND.n3586 25854
R13 GND.n3558 GND.n3557 23278.5
R14 GND.n497 GND.n495 20340.7
R15 GND.n192 GND.n190 20340.7
R16 GND.n1478 GND.n1477 20340.7
R17 GND.n4200 GND.n4198 20340.7
R18 GND.n3394 GND.n3392 20340.7
R19 GND.n3237 GND.n3235 20340.7
R20 GND.n2940 GND.n2938 20340.7
R21 GND.n2615 GND.n2613 20340.7
R22 GND.n2291 GND.n2289 20340.7
R23 GND.n2129 GND.n2127 20340.7
R24 GND.n1261 GND.n1259 20340.7
R25 GND.n344 GND.n342 20340.7
R26 GND.n7427 GND.n7426 20340.7
R27 GND.n7429 GND.n7428 20223.1
R28 GND.n1980 GND.n1525 20169.3
R29 GND GND.n1982 13209.6
R30 GND.n495 GND 13209.6
R31 GND.n190 GND 13209.6
R32 GND.n1525 GND 13209.6
R33 GND.n1477 GND 13209.6
R34 GND.n4198 GND 13209.6
R35 GND.n3392 GND 13209.6
R36 GND.n3235 GND 13209.6
R37 GND.n2938 GND 13209.6
R38 GND.n2613 GND 13209.6
R39 GND.n2289 GND 13209.6
R40 GND.n2127 GND 13209.6
R41 GND.n1259 GND 13209.6
R42 GND.n342 GND 13209.6
R43 GND.n7426 GND 13209.6
R44 GND.n1982 GND.n1981 12525.6
R45 GND.n6795 GND.t397 10105.3
R46 GND.n4918 GND.t349 10105.3
R47 GND.n87 GND.n86 8769.23
R48 GND.t777 GND.n981 6847.68
R49 GND.n6796 GND.t60 5863.39
R50 GND.n4919 GND.t428 5863.39
R51 GND.n3562 GND.n3558 4921.69
R52 GND.n3591 GND.n3587 4780.92
R53 GND.n6735 GND 4548.57
R54 GND.n4149 GND.n4146 4526.39
R55 GND.n4145 GND.n4138 4526.07
R56 GND.n4157 GND.n4150 4525.74
R57 GND.n4128 GND.n4125 4519.41
R58 GND.n3609 GND.n3604 4519.41
R59 GND.n3609 GND.n3605 4519.41
R60 GND.n3603 GND.n3600 4519.41
R61 GND.n3599 GND.n3596 4519.41
R62 GND.n3595 GND.n3592 4519.41
R63 GND.n4130 GND.n4124 4519.41
R64 GND.n4137 GND.n4123 4519.41
R65 GND.n3585 GND.n3582 4519.41
R66 GND.n4122 GND.n4113 4519.41
R67 GND.n3581 GND.n3579 4519.41
R68 GND.n3578 GND.n3574 4519.41
R69 GND.n3578 GND.n3575 4519.41
R70 GND.n4112 GND.n4111 4519.41
R71 GND.n4110 GND.n4102 4519.41
R72 GND.n4110 GND.n4103 4519.41
R73 GND.n3573 GND.n3570 4519.41
R74 GND.n4101 GND.n4098 4519.41
R75 GND.n3565 GND.n3563 4519.41
R76 GND.n3562 GND.n3556 4519.41
R77 GND.n4092 GND.n4079 4519.41
R78 GND.n4085 GND.n4084 4519.41
R79 GND.n3555 GND.n3550 4519.41
R80 GND.n3555 GND.n3551 4519.41
R81 GND.n4078 GND.n4074 4377.09
R82 GND.n3624 GND.n3539 3876.26
R83 GND.n3682 GND.n3670 3876.26
R84 GND.n6876 GND.t34 3455.76
R85 GND.t236 GND.n4577 3428.59
R86 GND.n6874 GND.n6873 3003.29
R87 GND.n4976 GND.n4275 2817.54
R88 GND.n6735 GND.n5490 2744.41
R89 GND.n4917 GND.n4916 2744.41
R90 GND.n6797 GND.t656 2656.51
R91 GND.n1980 GND.n1540 2549.93
R92 GND.n6801 GND.n6800 2243.42
R93 GND.n6799 GND.n4426 1899.15
R94 GND.n7713 GND.n7712 1773
R95 GND.n666 GND.n665 1773
R96 GND.n6381 GND.n6380 1773
R97 GND.n6217 GND.n6216 1773
R98 GND.n6053 GND.n6052 1773
R99 GND.n5867 GND.n5866 1773
R100 GND.n5345 GND.n5344 1773
R101 GND.n5384 GND.n5383 1773
R102 GND.n4808 GND.n4807 1773
R103 GND.n7115 GND.n7114 1773
R104 GND.n2787 GND.n2786 1773
R105 GND.n2462 GND.n2461 1773
R106 GND.n6978 GND.n6977 1773
R107 GND.n1813 GND.n1812 1773
R108 GND.n1717 GND.n1716 1773
R109 GND.n1955 GND.n1954 1773
R110 GND.n6799 GND.n6798 1742.45
R111 GND.n6797 GND.n6796 1566.95
R112 GND.n6796 GND.n6795 1560.68
R113 GND.n4918 GND.n4917 1548.15
R114 GND.n4917 GND.n4426 1548.15
R115 GND.t208 GND.n7583 1465.31
R116 GND.n7658 GND.n7655 1390.42
R117 GND.n614 GND.n611 1390.42
R118 GND.n6326 GND.n6323 1390.42
R119 GND.n6162 GND.n6159 1390.42
R120 GND.n5995 GND.n5992 1390.42
R121 GND.n5812 GND.n5809 1390.42
R122 GND.n5290 GND.n5287 1390.42
R123 GND.n4849 GND.n4846 1390.42
R124 GND.n7156 GND.n7153 1390.42
R125 GND.n3056 GND.n3053 1390.42
R126 GND.n2732 GND.n2729 1390.42
R127 GND.n2407 GND.n2404 1390.42
R128 GND.n6923 GND.n6920 1390.42
R129 GND.n1758 GND.n1755 1390.42
R130 GND.n1567 GND.n1564 1390.42
R131 GND.n1549 GND.n1546 1390.42
R132 GND.n7715 GND.n7713 1384.79
R133 GND.n668 GND.n666 1384.79
R134 GND.n6383 GND.n6381 1384.79
R135 GND.n6219 GND.n6217 1384.79
R136 GND.n6055 GND.n6053 1384.79
R137 GND.n5869 GND.n5867 1384.79
R138 GND.n5347 GND.n5345 1384.79
R139 GND.n5386 GND.n5384 1384.79
R140 GND.n4810 GND.n4808 1384.79
R141 GND.n7117 GND.n7115 1384.79
R142 GND.n2789 GND.n2787 1384.79
R143 GND.n2464 GND.n2462 1384.79
R144 GND.n6980 GND.n6978 1384.79
R145 GND.n1815 GND.n1813 1384.79
R146 GND.n1719 GND.n1717 1384.79
R147 GND.n1957 GND.n1955 1384.79
R148 GND.n4920 GND.n4919 1309.97
R149 GND.t772 GND.n6799 1269.38
R150 GND.n7478 GND.n7477 1266.06
R151 GND GND.t1322 1255.01
R152 GND GND.t68 1255.01
R153 GND.n3847 GND.n3841 1176.21
R154 GND.n3822 GND.n3817 1176.21
R155 GND.n3807 GND.n3802 1176.21
R156 GND.n3792 GND.n3787 1176.21
R157 GND.n3777 GND.n3772 1176.21
R158 GND.n3758 GND.n3753 1176.21
R159 GND.n3743 GND.n3738 1176.21
R160 GND.n3728 GND.n3723 1176.21
R161 GND.n3713 GND.n3708 1176.21
R162 GND.n4032 GND.n3657 1176.21
R163 GND.n4025 GND.n4015 1176.21
R164 GND.n4010 GND.n4009 1176.21
R165 GND.n3995 GND.n3994 1176.21
R166 GND.n3980 GND.n3979 1176.21
R167 GND.n3965 GND.n3964 1176.21
R168 GND.n3948 GND.n3947 1176.21
R169 GND.n3933 GND.n3932 1176.21
R170 GND.n3918 GND.n3917 1176.21
R171 GND.n3903 GND.n3902 1176.21
R172 GND.n3888 GND.n3887 1176.21
R173 GND.n3867 GND.n3866 1176.21
R174 GND.n3849 GND.n3848 1176.21
R175 GND.n3824 GND.n3823 1176.21
R176 GND.n3809 GND.n3808 1176.21
R177 GND.n3794 GND.n3793 1176.21
R178 GND.n3779 GND.n3778 1176.21
R179 GND.n3760 GND.n3759 1176.21
R180 GND.n3745 GND.n3744 1176.21
R181 GND.n3730 GND.n3729 1176.21
R182 GND.n3715 GND.n3714 1176.21
R183 GND.n4033 GND.n3653 1176.21
R184 GND.n4024 GND.n4019 1176.21
R185 GND.n4008 GND.n4003 1176.21
R186 GND.n3993 GND.n3988 1176.21
R187 GND.n3978 GND.n3973 1176.21
R188 GND.n3963 GND.n3958 1176.21
R189 GND.n3946 GND.n3941 1176.21
R190 GND.n3931 GND.n3926 1176.21
R191 GND.n3916 GND.n3911 1176.21
R192 GND.n3901 GND.n3896 1176.21
R193 GND.n3886 GND.n3879 1176.21
R194 GND.n3865 GND.n3859 1176.21
R195 GND.n7483 GND.n7476 1153.03
R196 GND.n2071 GND.n2068 1153.03
R197 GND.n403 GND.n400 1153.03
R198 GND.n560 GND.n557 1153.03
R199 GND.n251 GND.n248 1153.03
R200 GND.n99 GND.n96 1153.03
R201 GND.n1432 GND.n1429 1153.03
R202 GND.n4259 GND.n4256 1153.03
R203 GND.n3456 GND.n3453 1153.03
R204 GND.n3298 GND.n3295 1153.03
R205 GND.n3002 GND.n2999 1153.03
R206 GND.n2678 GND.n2675 1153.03
R207 GND.n2353 GND.n2350 1153.03
R208 GND.n2195 GND.n2192 1153.03
R209 GND.n1312 GND.n1309 1153.03
R210 GND.n829 GND.n826 1153.03
R211 GND.t1198 GND.n6560 1137.9
R212 GND GND.t666 1129.73
R213 GND.n1038 GND.n1035 1077.71
R214 GND.n1034 GND.n1029 1077.71
R215 GND.n1034 GND.n1030 1077.71
R216 GND.n7449 GND.n7446 1077.71
R217 GND.n7451 GND.n7444 1077.71
R218 GND.n1349 GND.n1345 1077.71
R219 GND.n2036 GND.n2028 1077.71
R220 GND.n2038 GND.n2026 1077.71
R221 GND.n1344 GND.n1340 1077.71
R222 GND.n1344 GND.n1341 1077.71
R223 GND.n1023 GND.n1020 1077.71
R224 GND.n1019 GND.n1014 1077.71
R225 GND.n1019 GND.n1015 1077.71
R226 GND.n529 GND.n526 1077.71
R227 GND.n531 GND.n524 1077.71
R228 GND.n1003 GND.n999 1077.71
R229 GND.n998 GND.n994 1077.71
R230 GND.n998 GND.n995 1077.71
R231 GND.n224 GND.n221 1077.71
R232 GND.n226 GND.n219 1077.71
R233 GND.n993 GND.n988 1077.71
R234 GND.n987 GND.n979 1077.71
R235 GND.n987 GND.n980 1077.71
R236 GND.n60 GND.n59 1077.71
R237 GND.n65 GND.n64 1077.71
R238 GND.n978 GND.n974 1077.71
R239 GND.n978 GND.n975 1077.71
R240 GND.n973 GND.n969 1077.71
R241 GND.n1398 GND.n1395 1077.71
R242 GND.n1400 GND.n1393 1077.71
R243 GND.n968 GND.n965 1077.71
R244 GND.n964 GND.n959 1077.71
R245 GND.n964 GND.n960 1077.71
R246 GND.n4232 GND.n4229 1077.71
R247 GND.n4234 GND.n4227 1077.71
R248 GND.n958 GND.n954 1077.71
R249 GND.n953 GND.n949 1077.71
R250 GND.n953 GND.n950 1077.71
R251 GND.n3426 GND.n3423 1077.71
R252 GND.n3428 GND.n3421 1077.71
R253 GND.n948 GND.n944 1077.71
R254 GND.n948 GND.n945 1077.71
R255 GND.n943 GND.n939 1077.71
R256 GND.n3269 GND.n3266 1077.71
R257 GND.n3271 GND.n3264 1077.71
R258 GND.n938 GND.n935 1077.71
R259 GND.n934 GND.n929 1077.71
R260 GND.n934 GND.n930 1077.71
R261 GND.n2972 GND.n2969 1077.71
R262 GND.n2974 GND.n2967 1077.71
R263 GND.n928 GND.n924 1077.71
R264 GND.n928 GND.n925 1077.71
R265 GND.n923 GND.n919 1077.71
R266 GND.n2647 GND.n2644 1077.71
R267 GND.n2649 GND.n2642 1077.71
R268 GND.n918 GND.n913 1077.71
R269 GND.n918 GND.n914 1077.71
R270 GND.n912 GND.n909 1077.71
R271 GND.n2323 GND.n2320 1077.71
R272 GND.n2325 GND.n2318 1077.71
R273 GND.n908 GND.n904 1077.71
R274 GND.n908 GND.n905 1077.71
R275 GND.n903 GND.n899 1077.71
R276 GND.n2161 GND.n2158 1077.71
R277 GND.n2163 GND.n2156 1077.71
R278 GND.n1334 GND.n1330 1077.71
R279 GND.n1339 GND.n1335 1077.71
R280 GND.n1339 GND.n1336 1077.71
R281 GND.n1293 GND.n1290 1077.71
R282 GND.n1295 GND.n1288 1077.71
R283 GND.n1009 GND.n1004 1077.71
R284 GND.n1009 GND.n1005 1077.71
R285 GND.n376 GND.n373 1077.71
R286 GND.n378 GND.n371 1077.71
R287 GND.n1013 GND.n1010 1077.71
R288 GND.n801 GND.n798 1077.71
R289 GND.n1028 GND.n1024 1077.71
R290 GND.n1028 GND.n1025 1077.71
R291 GND.n803 GND.n796 1077.71
R292 GND.n1043 GND.n1039 1077.71
R293 GND GND.t497 1058.96
R294 GND GND.t353 1058.96
R295 GND GND.t129 1058.96
R296 GND GND.t379 1058.96
R297 GND GND.t506 1058.96
R298 GND GND.t842 1058.96
R299 GND GND.t1188 1058.96
R300 GND GND.t809 1058.96
R301 GND GND.t177 1058.96
R302 GND GND.t577 1058.96
R303 GND GND.t612 1058.96
R304 GND GND.t26 1058.96
R305 GND GND.t134 1058.96
R306 GND GND.t482 1058.96
R307 GND GND.t369 1058.96
R308 GND GND.t53 1058.96
R309 GND.n7451 GND.n7443 1054.53
R310 GND.n2038 GND.n2025 1054.53
R311 GND.n531 GND.n523 1054.53
R312 GND.n226 GND.n218 1054.53
R313 GND.n65 GND.n63 1054.53
R314 GND.n1400 GND.n1392 1054.53
R315 GND.n4234 GND.n4226 1054.53
R316 GND.n3428 GND.n3420 1054.53
R317 GND.n3271 GND.n3263 1054.53
R318 GND.n2974 GND.n2966 1054.53
R319 GND.n2649 GND.n2641 1054.53
R320 GND.n2325 GND.n2317 1054.53
R321 GND.n2163 GND.n2155 1054.53
R322 GND.n1295 GND.n1287 1054.53
R323 GND.n378 GND.n370 1054.53
R324 GND.n803 GND.n795 1054.53
R325 GND.n4915 GND.n4914 940.789
R326 GND.t1244 GND 917.571
R327 GND GND.t688 917.571
R328 GND.n7700 GND.n7696 915.471
R329 GND.n7723 GND.n7722 915.471
R330 GND.n7553 GND.n7552 915.471
R331 GND.n653 GND.n649 915.471
R332 GND.n676 GND.n675 915.471
R333 GND.n7684 GND.n7683 915.471
R334 GND.n6365 GND.n6361 915.471
R335 GND.n6391 GND.n6390 915.471
R336 GND.n637 GND.n636 915.471
R337 GND.n6201 GND.n6197 915.471
R338 GND.n6227 GND.n6226 915.471
R339 GND.n6349 GND.n6348 915.471
R340 GND.n6037 GND.n6033 915.471
R341 GND.n6063 GND.n6062 915.471
R342 GND.n6185 GND.n6184 915.471
R343 GND.n5854 GND.n5850 915.471
R344 GND.n5877 GND.n5876 915.471
R345 GND.n6021 GND.n6020 915.471
R346 GND.n5332 GND.n5328 915.471
R347 GND.n5355 GND.n5354 915.471
R348 GND.n5838 GND.n5837 915.471
R349 GND.n4891 GND.n4887 915.471
R350 GND.n5394 GND.n5393 915.471
R351 GND.n5316 GND.n5315 915.471
R352 GND.n7198 GND.n7194 915.471
R353 GND.n4818 GND.n4817 915.471
R354 GND.n4875 GND.n4874 915.471
R355 GND.n3098 GND.n3094 915.471
R356 GND.n7125 GND.n7124 915.471
R357 GND.n7182 GND.n7181 915.471
R358 GND.n2774 GND.n2770 915.471
R359 GND.n2797 GND.n2796 915.471
R360 GND.n3082 GND.n3081 915.471
R361 GND.n2449 GND.n2445 915.471
R362 GND.n2472 GND.n2471 915.471
R363 GND.n2758 GND.n2757 915.471
R364 GND.n6965 GND.n6961 915.471
R365 GND.n6988 GND.n6987 915.471
R366 GND.n2433 GND.n2432 915.471
R367 GND.n1800 GND.n1796 915.471
R368 GND.n1823 GND.n1822 915.471
R369 GND.n6949 GND.n6948 915.471
R370 GND.n1609 GND.n1605 915.471
R371 GND.n1727 GND.n1726 915.471
R372 GND.n1784 GND.n1783 915.471
R373 GND.n1545 GND.n1541 915.471
R374 GND.n1965 GND.n1964 915.471
R375 GND.n1593 GND.n1592 915.471
R376 GND.n7566 GND.n7563 841.244
R377 GND.n7702 GND.n7694 841.244
R378 GND.n655 GND.n647 841.244
R379 GND.n6367 GND.n6359 841.244
R380 GND.n6203 GND.n6195 841.244
R381 GND.n6039 GND.n6031 841.244
R382 GND.n5856 GND.n5848 841.244
R383 GND.n5334 GND.n5326 841.244
R384 GND.n4893 GND.n4885 841.244
R385 GND.n7200 GND.n7192 841.244
R386 GND.n3100 GND.n3092 841.244
R387 GND.n2776 GND.n2768 841.244
R388 GND.n2451 GND.n2443 841.244
R389 GND.n6967 GND.n6959 841.244
R390 GND.n1802 GND.n1794 841.244
R391 GND.n1611 GND.n1603 841.244
R392 GND.t1291 GND.n1891 808.275
R393 GND.t49 GND.n1848 808.275
R394 GND.n7043 GND.t573 808.275
R395 GND.t491 GND.n2497 808.275
R396 GND.t1374 GND.n2822 808.275
R397 GND.t4 GND.n3119 808.275
R398 GND.t1267 GND.n7219 808.275
R399 GND.t1322 GND.t0 806.792
R400 GND.t68 GND.t1176 806.792
R401 GND.n4071 GND.n4069 806.47
R402 GND GND.t154 784.713
R403 GND GND.t140 784.713
R404 GND.t1299 GND.t656 780.297
R405 GND.t34 GND.t701 780.297
R406 GND.n7815 GND.n7811 778.15
R407 GND.n7815 GND.n7812 778.15
R408 GND.n885 GND.n880 778.15
R409 GND.n885 GND.n881 778.15
R410 GND.n2060 GND.n2056 778.15
R411 GND.n2060 GND.n2059 778.15
R412 GND.n1663 GND.n1658 778.15
R413 GND.n1663 GND.n1659 778.15
R414 GND.n453 GND.n448 778.15
R415 GND.n453 GND.n449 778.15
R416 GND.n772 GND.n767 778.15
R417 GND.n772 GND.n768 778.15
R418 GND.n459 GND.n454 778.15
R419 GND.n459 GND.n455 778.15
R420 GND.n300 GND.n295 778.15
R421 GND.n300 GND.n296 778.15
R422 GND.n154 GND.n149 778.15
R423 GND.n154 GND.n150 778.15
R424 GND.n148 GND.n143 778.15
R425 GND.n148 GND.n144 778.15
R426 GND.n45 GND.n40 778.15
R427 GND.n45 GND.n41 778.15
R428 GND.n39 GND.n34 778.15
R429 GND.n39 GND.n35 778.15
R430 GND.n7301 GND.n7296 778.15
R431 GND.n7301 GND.n7297 778.15
R432 GND.n7295 GND.n7290 778.15
R433 GND.n7295 GND.n7291 778.15
R434 GND.n3511 GND.n3506 778.15
R435 GND.n3511 GND.n3507 778.15
R436 GND.n3505 GND.n3500 778.15
R437 GND.n3505 GND.n3501 778.15
R438 GND.n3353 GND.n3348 778.15
R439 GND.n3353 GND.n3349 778.15
R440 GND.n3347 GND.n3342 778.15
R441 GND.n3347 GND.n3343 778.15
R442 GND.n3196 GND.n3191 778.15
R443 GND.n3196 GND.n3192 778.15
R444 GND.n3190 GND.n3185 778.15
R445 GND.n3190 GND.n3186 778.15
R446 GND.n2899 GND.n2894 778.15
R447 GND.n2899 GND.n2895 778.15
R448 GND.n2893 GND.n2888 778.15
R449 GND.n2893 GND.n2889 778.15
R450 GND.n2574 GND.n2569 778.15
R451 GND.n2574 GND.n2570 778.15
R452 GND.n2568 GND.n2563 778.15
R453 GND.n2568 GND.n2564 778.15
R454 GND.n2250 GND.n2245 778.15
R455 GND.n2250 GND.n2246 778.15
R456 GND.n2244 GND.n2239 778.15
R457 GND.n2244 GND.n2240 778.15
R458 GND.n1225 GND.n1220 778.15
R459 GND.n1225 GND.n1221 778.15
R460 GND.n1219 GND.n1214 778.15
R461 GND.n1219 GND.n1215 778.15
R462 GND.n1677 GND.n1664 778.15
R463 GND.n1677 GND.n1665 778.15
R464 GND.n306 GND.n301 778.15
R465 GND.n306 GND.n302 778.15
R466 GND.n879 GND.n874 778.15
R467 GND.n879 GND.n875 778.15
R468 GND.n778 GND.n773 778.15
R469 GND.n778 GND.n774 778.15
R470 GND.t1305 GND.t1138 777.333
R471 GND.t515 GND.t351 777.333
R472 GND.t1302 GND 754.5
R473 GND.t695 GND 754.5
R474 GND.t60 GND.t1209 732.088
R475 GND.t428 GND.t786 732.088
R476 GND GND.t109 729.721
R477 GND.t665 GND 729.721
R478 GND.t1304 GND 726
R479 GND GND.t696 726
R480 GND.t16 GND.t1532 717.149
R481 GND.t1386 GND.t426 717.149
R482 GND.t115 GND.t1244 708.047
R483 GND.t688 GND.t151 708.047
R484 GND.t102 GND.n6088 706.715
R485 GND.t768 GND.n6252 706.715
R486 GND.t191 GND.n701 706.715
R487 GND.t1220 GND.n7748 706.715
R488 GND.t64 GND 654.159
R489 GND.n4976 GND 654.054
R490 GND.t1209 GND.t788 627.505
R491 GND.t788 GND.t16 627.505
R492 GND.t0 GND.t1302 627.505
R493 GND.t786 GND.t1568 627.505
R494 GND.t1568 GND.t1386 627.505
R495 GND.t1176 GND.t695 627.505
R496 GND.t109 GND.t1299 606.898
R497 GND.t714 GND.t115 606.898
R498 GND.t203 GND.t714 606.898
R499 GND.t701 GND.t665 606.898
R500 GND.t151 GND.t600 606.898
R501 GND.t600 GND.t1143 606.898
R502 GND.t476 GND.t1296 601.333
R503 GND.t705 GND.t659 601.333
R504 GND.t1202 GND.n6561 565.158
R505 GND.n4913 GND.t751 550.154
R506 GND GND.t20 546.497
R507 GND GND.t90 546.497
R508 GND.n7700 GND.n7697 521.471
R509 GND.n653 GND.n650 521.471
R510 GND.n6365 GND.n6362 521.471
R511 GND.n6201 GND.n6198 521.471
R512 GND.n6037 GND.n6034 521.471
R513 GND.n5854 GND.n5851 521.471
R514 GND.n5332 GND.n5329 521.471
R515 GND.n4891 GND.n4888 521.471
R516 GND.n7198 GND.n7195 521.471
R517 GND.n3098 GND.n3095 521.471
R518 GND.n2774 GND.n2771 521.471
R519 GND.n2449 GND.n2446 521.471
R520 GND.n6965 GND.n6962 521.471
R521 GND.n1800 GND.n1797 521.471
R522 GND.n1609 GND.n1606 521.471
R523 GND.n1545 GND.n1542 521.471
R524 GND.n7748 GND.n7747 515.509
R525 GND.n701 GND.n700 515.509
R526 GND.n6416 GND.n6415 515.509
R527 GND.n6252 GND.n6251 515.509
R528 GND.n6088 GND.n6087 515.509
R529 GND.n4912 GND.n4911 515.509
R530 GND.n7219 GND.n7218 515.509
R531 GND.n3119 GND.n3118 515.509
R532 GND.n2822 GND.n2821 515.509
R533 GND.n2497 GND.n2496 515.509
R534 GND.n7043 GND.n6878 515.509
R535 GND.n1848 GND.n1847 515.509
R536 GND.n1891 GND.n1890 515.509
R537 GND GND.t412 513.333
R538 GND.t706 GND.t376 498.408
R539 GND.n7660 GND 484.329
R540 GND.n616 GND 484.329
R541 GND.n6328 GND 484.329
R542 GND.n6164 GND 484.329
R543 GND.n5997 GND 484.329
R544 GND.n5814 GND 484.329
R545 GND.n5292 GND 484.329
R546 GND.n4851 GND 484.329
R547 GND.n7158 GND 484.329
R548 GND.n3058 GND 484.329
R549 GND.n2734 GND 484.329
R550 GND.n2409 GND 484.329
R551 GND.n6925 GND 484.329
R552 GND.n1760 GND 484.329
R553 GND.n1569 GND 484.329
R554 GND.n1551 GND 484.329
R555 GND.n7487 GND.n7486 480.913
R556 GND.n2077 GND.n2067 480.913
R557 GND.n409 GND.n399 480.913
R558 GND.n564 GND.n563 480.913
R559 GND.n255 GND.n254 480.913
R560 GND.n103 GND.n102 480.913
R561 GND.n1436 GND.n1435 480.913
R562 GND.n4263 GND.n4262 480.913
R563 GND.n3460 GND.n3459 480.913
R564 GND.n3302 GND.n3301 480.913
R565 GND.n3006 GND.n3005 480.913
R566 GND.n2682 GND.n2681 480.913
R567 GND.n2357 GND.n2356 480.913
R568 GND.n2199 GND.n2198 480.913
R569 GND.n1318 GND.n1308 480.913
R570 GND.n835 GND.n825 480.913
R571 GND.t376 GND 478.938
R572 GND.t1532 GND 478.099
R573 GND.t426 GND 478.099
R574 GND.n7566 GND.n7564 473.865
R575 GND.n7702 GND.n7695 473.865
R576 GND.n655 GND.n648 473.865
R577 GND.n6367 GND.n6360 473.865
R578 GND.n6203 GND.n6196 473.865
R579 GND.n6039 GND.n6032 473.865
R580 GND.n5856 GND.n5849 473.865
R581 GND.n5334 GND.n5327 473.865
R582 GND.n4893 GND.n4886 473.865
R583 GND.n7200 GND.n7193 473.865
R584 GND.n3100 GND.n3093 473.865
R585 GND.n2776 GND.n2769 473.865
R586 GND.n2451 GND.n2444 473.865
R587 GND.n6967 GND.n6960 473.865
R588 GND.n1802 GND.n1795 473.865
R589 GND.n1611 GND.n1604 473.865
R590 GND.n4919 GND.n4275 445.014
R591 GND.t1225 GND 426.178
R592 GND.t1223 GND.t64 420.531
R593 GND.n5177 GND 420.382
R594 GND.n6875 GND 420.382
R595 GND.n5177 GND.t203 419.048
R596 GND.t1143 GND.n6875 419.048
R597 GND.t823 GND.n7363 405.955
R598 GND GND.t708 393.274
R599 GND.t424 GND.t772 381.594
R600 GND.t770 GND.t470 373.805
R601 GND.n7045 GND.n6877 367.533
R602 GND GND.t346 339.942
R603 GND GND.t703 339.942
R604 GND.n7450 GND.n7445 331.909
R605 GND.n530 GND.n525 331.909
R606 GND.n377 GND.n372 331.909
R607 GND.n225 GND.n220 331.909
R608 GND.n4233 GND.n4228 331.909
R609 GND.n3270 GND.n3265 331.909
R610 GND.n2648 GND.n2643 331.909
R611 GND.n2162 GND.n2157 331.909
R612 GND.n1294 GND.n1289 331.909
R613 GND.n2324 GND.n2319 331.909
R614 GND.n2973 GND.n2968 331.909
R615 GND.n3427 GND.n3422 331.909
R616 GND.n1399 GND.n1394 331.909
R617 GND.n2037 GND.n2027 331.909
R618 GND.n802 GND.n797 331.909
R619 GND.n192 GND.n191 328.866
R620 GND.n1491 GND.n1490 328.866
R621 GND.n1980 GND.n1478 328.866
R622 GND.n4200 GND.n4199 328.866
R623 GND.n3394 GND.n3393 328.866
R624 GND.n3237 GND.n3236 328.866
R625 GND.n2940 GND.n2939 328.866
R626 GND.n2615 GND.n2614 328.866
R627 GND.n2291 GND.n2290 328.866
R628 GND.n2129 GND.n2128 328.866
R629 GND.n1261 GND.n1260 328.866
R630 GND.n1998 GND.n1997 328.866
R631 GND.n497 GND.n496 328.866
R632 GND.n344 GND.n343 328.866
R633 GND.n7428 GND.n7427 328.866
R634 GND.t1131 GND.t424 327.08
R635 GND.t470 GND.t1131 327.08
R636 GND.t708 GND.t1223 327.08
R637 GND.t630 GND.t640 324.212
R638 GND.t652 GND.t642 324.212
R639 GND.t632 GND.t652 324.212
R640 GND.t638 GND.t632 324.212
R641 GND.t648 GND.t638 324.212
R642 GND.t644 GND.t648 324.212
R643 GND.t626 GND.t636 324.212
R644 GND.t622 GND.t634 324.212
R645 GND.t412 GND.t415 324.212
R646 GND.t415 GND.t417 324.212
R647 GND.t417 GND.t410 324.212
R648 GND.t875 GND 308.692
R649 GND GND.t863 308.692
R650 GND GND.t941 308.692
R651 GND.t450 GND 308.692
R652 GND GND.t1350 306.387
R653 GND.t784 GND.n6734 304.084
R654 GND.t634 GND 301.053
R655 GND.n6800 GND 299.824
R656 GND.n3554 GND.n3552 293.647
R657 GND.n3554 GND.n3553 293.647
R658 GND.n3561 GND.n3559 293.647
R659 GND.n3561 GND.n3560 293.647
R660 GND.n3568 GND.n3566 293.647
R661 GND.n3568 GND.n3567 293.647
R662 GND.n3572 GND.n3571 293.647
R663 GND.n3577 GND.n3576 293.647
R664 GND.n3584 GND.n3583 293.647
R665 GND.n3590 GND.n3588 293.647
R666 GND.n3590 GND.n3589 293.647
R667 GND.n3594 GND.n3593 293.647
R668 GND.n3598 GND.n3597 293.647
R669 GND.n3602 GND.n3601 293.647
R670 GND.n3608 GND.n3606 293.647
R671 GND.n3608 GND.n3607 293.647
R672 GND.n92 GND.n91 290.183
R673 GND.n4978 GND.t646 285.615
R674 GND.n100 GND.n87 285.455
R675 GND.t676 GND.t706 280.354
R676 GND.t1175 GND.t676 280.354
R677 GND.n5015 GND.t628 270.175
R678 GND.n6757 GND.n6755 267.089
R679 GND GND.t153 266.514
R680 GND GND.t528 266.514
R681 GND GND.t1368 263.26
R682 GND.n4913 GND.n4912 258.123
R683 GND GND.t1175 253.097
R684 GND.n4920 GND.n4918 250.713
R685 GND GND.t770 249.204
R686 GND GND.t784 244.189
R687 GND GND.t174 230.905
R688 GND GND.t699 230.905
R689 GND.t1119 GND 227.501
R690 GND.t575 GND.t1225 223.457
R691 GND GND.t166 216.544
R692 GND.t1425 GND.n5509 214.877
R693 GND.n6757 GND.n6756 213.671
R694 GND.n6798 GND.n6797 213.106
R695 GND.n4977 GND 211.114
R696 GND.n991 GND.n990 209.695
R697 GND.n984 GND.n983 209.695
R698 GND.n7481 GND.n7480 203.294
R699 GND.n4275 GND.t644 196.843
R700 GND.n7459 GND.n7458 195.531
R701 GND.n2046 GND.n2045 195.531
R702 GND.n386 GND.n385 195.531
R703 GND.n539 GND.n538 195.531
R704 GND.n234 GND.n233 195.531
R705 GND.n1408 GND.n1407 195.531
R706 GND.n4242 GND.n4241 195.531
R707 GND.n3436 GND.n3435 195.531
R708 GND.n3279 GND.n3278 195.531
R709 GND.n2982 GND.n2981 195.531
R710 GND.n2657 GND.n2656 195.531
R711 GND.n2333 GND.n2332 195.531
R712 GND.n2171 GND.n2170 195.531
R713 GND.n1303 GND.n1302 195.531
R714 GND.n811 GND.n810 195.531
R715 GND.n6710 GND.t1349 193.933
R716 GND.n1929 GND.t54 193.933
R717 GND.n1894 GND.t1285 193.933
R718 GND.n1696 GND.t372 193.933
R719 GND.n1851 GND.t43 193.933
R720 GND.n6904 GND.t483 193.933
R721 GND.n6879 GND.t567 193.933
R722 GND.n2372 GND.t138 193.933
R723 GND.n2500 GND.t494 193.933
R724 GND.n2697 GND.t27 193.933
R725 GND.n2825 GND.t1377 193.933
R726 GND.n3021 GND.t613 193.933
R727 GND.n3122 GND.t8 193.933
R728 GND.n7094 GND.t581 193.933
R729 GND.n7222 GND.t1270 193.933
R730 GND.n4789 GND.t180 193.933
R731 GND.n4754 GND.t754 193.933
R732 GND.n5271 GND.t814 193.933
R733 GND.n5246 GND.t1392 193.933
R734 GND.n5793 GND.t1192 193.933
R735 GND.n5922 GND.t1326 193.933
R736 GND.n5960 GND.t843 193.933
R737 GND.n6091 GND.t96 193.933
R738 GND.n6127 GND.t507 193.933
R739 GND.n6255 GND.t762 193.933
R740 GND.n6291 GND.t380 193.933
R741 GND.n6564 GND.t1205 193.933
R742 GND.n579 GND.t130 193.933
R743 GND.n704 GND.t194 193.933
R744 GND.n7622 GND.t357 193.933
R745 GND.n7751 GND.t1214 193.933
R746 GND.n7502 GND.t500 193.933
R747 GND.n7586 GND.t211 193.933
R748 GND.n4950 GND.t414 193.933
R749 GND.n5741 GND.t1153 193.933
R750 GND.n5152 GND.t82 193.933
R751 GND.n5765 GND.t680 193.532
R752 GND.t899 GND.t873 193.508
R753 GND.t985 GND.t899 193.508
R754 GND.t877 GND.t985 193.508
R755 GND.t869 GND.t877 193.508
R756 GND.t891 GND.t869 193.508
R757 GND.t859 GND.t917 193.508
R758 GND.t895 GND.t859 193.508
R759 GND.t965 GND.t895 193.508
R760 GND.t861 GND.t965 193.508
R761 GND.t885 GND.t861 193.508
R762 GND.t949 GND.t885 193.508
R763 GND.t979 GND.t949 193.508
R764 GND.t911 GND.t979 193.508
R765 GND.t955 GND.t911 193.508
R766 GND.t943 GND.t875 193.508
R767 GND.t969 GND.t943 193.508
R768 GND.t867 GND.t969 193.508
R769 GND.t923 GND.t957 193.508
R770 GND.t957 GND.t889 193.508
R771 GND.t889 GND.t927 193.508
R772 GND.t927 GND.t961 193.508
R773 GND.t961 GND.t897 193.508
R774 GND.t897 GND.t977 193.508
R775 GND.t977 GND.t909 193.508
R776 GND.t909 GND.t935 193.508
R777 GND.t935 GND.t983 193.508
R778 GND.t983 GND.t915 193.508
R779 GND.t915 GND.t939 193.508
R780 GND.t863 GND.t921 193.508
R781 GND.t921 GND.t951 193.508
R782 GND.t951 GND.t887 193.508
R783 GND.t887 GND.t973 193.508
R784 GND.t947 GND.t883 193.508
R785 GND.t975 GND.t947 193.508
R786 GND.t905 GND.t975 193.508
R787 GND.t931 GND.t905 193.508
R788 GND.t963 GND.t907 193.508
R789 GND.t907 GND.t933 193.508
R790 GND.t933 GND.t879 193.508
R791 GND.t879 GND.t901 193.508
R792 GND.t901 GND.t919 193.508
R793 GND.t941 GND.t967 193.508
R794 GND.t967 GND.t865 193.508
R795 GND.t865 GND.t945 193.508
R796 GND.t903 GND.t971 193.508
R797 GND.t925 GND.t903 193.508
R798 GND.t959 GND.t925 193.508
R799 GND.t893 GND.t959 193.508
R800 GND.t929 GND.t893 193.508
R801 GND.t871 GND.t929 193.508
R802 GND.t953 GND.t871 193.508
R803 GND.t981 GND.t953 193.508
R804 GND.t913 GND.t981 193.508
R805 GND.t937 GND.t913 193.508
R806 GND.t881 GND.t937 193.508
R807 GND.t464 GND.t450 193.508
R808 GND.t444 GND.t464 193.508
R809 GND.t452 GND.t462 193.508
R810 GND.t462 GND.t458 193.508
R811 GND.t458 GND.t466 193.508
R812 GND.t466 GND.t446 193.508
R813 GND.t446 GND.t460 193.508
R814 GND.t460 GND.t468 193.508
R815 GND.t468 GND.t448 193.508
R816 GND.t448 GND.t454 193.508
R817 GND.t454 GND.t438 193.508
R818 GND.t438 GND.t442 193.508
R819 GND.t442 GND.t456 193.508
R820 GND.t456 GND.t440 193.508
R821 GND.t1350 GND.t1352 193.508
R822 GND.t1352 GND.t1354 193.508
R823 GND.t1354 GND.t1348 193.508
R824 GND.t166 GND.t575 193.508
R825 GND.n6700 GND.t1351 192.982
R826 GND.n1922 GND.t58 192.982
R827 GND.n1908 GND.t1292 192.982
R828 GND.n1689 GND.t371 192.982
R829 GND.n1865 GND.t50 192.982
R830 GND.n6897 GND.t486 192.982
R831 GND.n6886 GND.t574 192.982
R832 GND.n2365 GND.t136 192.982
R833 GND.n2514 GND.t492 192.982
R834 GND.n2690 GND.t30 192.982
R835 GND.n2839 GND.t1375 192.982
R836 GND.n3014 GND.t616 192.982
R837 GND.n3136 GND.t5 192.982
R838 GND.n7087 GND.t579 192.982
R839 GND.n7236 GND.t1268 192.982
R840 GND.n4782 GND.t178 192.982
R841 GND.n4768 GND.t752 192.982
R842 GND.n5264 GND.t812 192.982
R843 GND.n5253 GND.t1399 192.982
R844 GND.n5786 GND.t1190 192.982
R845 GND.n5936 GND.t1333 192.982
R846 GND.n5953 GND.t846 192.982
R847 GND.n6105 GND.t103 192.982
R848 GND.n6120 GND.t510 192.982
R849 GND.n6269 GND.t769 192.982
R850 GND.n6284 GND.t383 192.982
R851 GND.n6578 GND.t1203 192.982
R852 GND.n572 GND.t133 192.982
R853 GND.n718 GND.t192 192.982
R854 GND.n7615 GND.t355 192.982
R855 GND.n7765 GND.t1221 192.982
R856 GND.n7495 GND.t498 192.982
R857 GND.n7600 GND.t209 192.982
R858 GND.n4949 GND.t413 192.982
R859 GND.n5731 GND.t1155 192.982
R860 GND.n5142 GND.t84 192.982
R861 GND.t1427 GND 190.686
R862 GND GND.t1415 190.686
R863 GND.t1493 GND 190.686
R864 GND GND.t546 190.686
R865 GND GND.t1154 189.263
R866 GND.n7802 GND.n7799 185.779
R867 GND.t1059 GND.n4446 185.69
R868 GND.t360 GND 185.418
R869 GND GND.t797 185.418
R870 GND GND.t603 185.418
R871 GND GND.t591 185.418
R872 GND GND.t690 185.418
R873 GND GND.t1172 185.418
R874 GND GND.t662 185.418
R875 GND GND.t1278 185.418
R876 GND GND.t430 185.418
R877 GND GND.t420 185.418
R878 GND GND.t807 185.418
R879 GND GND.t120 185.418
R880 GND GND.t87 185.418
R881 GND GND.t848 185.418
R882 GND GND.t608 185.418
R883 GND.t112 GND 185.418
R884 GND.n5177 GND 182.167
R885 GND.n6875 GND 182.167
R886 GND GND.t185 181.03
R887 GND GND.t678 181.03
R888 GND GND.t955 179.686
R889 GND.t939 GND 179.686
R890 GND.t919 GND 179.686
R891 GND.t971 GND.n6657 179.686
R892 GND GND.t881 179.686
R893 GND.t440 GND 179.686
R894 GND.n5490 GND 176.386
R895 GND.n4916 GND 176.386
R896 GND.t1348 GND 172.775
R897 GND.n1267 GND.n1266 171.047
R898 GND.n2135 GND.n2134 171.047
R899 GND.n2297 GND.n2296 171.047
R900 GND.n2621 GND.n2620 171.047
R901 GND.n2946 GND.n2945 171.047
R902 GND.n3243 GND.n3242 171.047
R903 GND.n3400 GND.n3399 171.047
R904 GND.n4206 GND.n4205 171.047
R905 GND.n1449 GND.n1448 171.047
R906 GND.n1497 GND.n1496 171.047
R907 GND.n198 GND.n197 171.047
R908 GND.n2005 GND.n2003 171.047
R909 GND.n350 GND.n349 171.047
R910 GND.n503 GND.n502 171.047
R911 GND.n7398 GND.n7386 171.047
R912 GND GND.t1061 164.786
R913 GND.t1049 GND 164.786
R914 GND GND.t999 164.786
R915 GND.t1562 GND 164.786
R916 GND GND.t83 163.555
R917 GND.t66 GND.n5176 162.326
R918 GND.n3847 GND.n3840 162.236
R919 GND.t883 GND.n6559 161.257
R920 GND.t1332 GND.n5918 159.185
R921 GND.n6713 GND.t167 154.006
R922 GND.n5744 GND.t63 154.006
R923 GND.n5155 GND.t1315 154.006
R924 GND.n7470 GND.n7465 153.601
R925 GND.n7470 GND.n7469 153.601
R926 GND.n2064 GND.n2048 153.601
R927 GND.n2064 GND.n2063 153.601
R928 GND.n396 GND.n391 153.601
R929 GND.n551 GND.n545 153.601
R930 GND.n551 GND.n550 153.601
R931 GND.n242 GND.n240 153.601
R932 GND.n242 GND.n241 153.601
R933 GND.n81 GND.n76 153.601
R934 GND.n81 GND.n80 153.601
R935 GND.n1423 GND.n1414 153.601
R936 GND.n1423 GND.n1422 153.601
R937 GND.n4250 GND.n4244 153.601
R938 GND.n4250 GND.n4249 153.601
R939 GND.n3447 GND.n3441 153.601
R940 GND.n3447 GND.n3446 153.601
R941 GND.n3289 GND.n3284 153.601
R942 GND.n3289 GND.n3288 153.601
R943 GND.n2993 GND.n2988 153.601
R944 GND.n2993 GND.n2992 153.601
R945 GND.n2669 GND.n2663 153.601
R946 GND.n2669 GND.n2668 153.601
R947 GND.n2344 GND.n2338 153.601
R948 GND.n2344 GND.n2343 153.601
R949 GND.n2186 GND.n2176 153.601
R950 GND.n2186 GND.n2185 153.601
R951 GND.n396 GND.n395 153.601
R952 GND.n822 GND.n817 153.601
R953 GND.n822 GND.n821 153.601
R954 GND.t680 GND 150.841
R955 GND.n5468 GND.t365 150.465
R956 GND.n4399 GND.t771 150.465
R957 GND.n6776 GND.t215 150.465
R958 GND.n5233 GND.t1533 150.465
R959 GND.n5180 GND.t1311 150.465
R960 GND.n5213 GND.t1195 150.465
R961 GND.n4354 GND.t858 150.465
R962 GND.n4325 GND.t427 150.465
R963 GND.n4277 GND.t801 150.465
R964 GND.n4310 GND.t148 150.465
R965 GND.t222 GND 149.645
R966 GND GND.t252 149.645
R967 GND.t270 GND 149.645
R968 GND GND.t624 149.645
R969 GND.n1266 GND.n1261 148.436
R970 GND.n2134 GND.n2129 148.436
R971 GND.n2296 GND.n2291 148.436
R972 GND.n2620 GND.n2615 148.436
R973 GND.n2945 GND.n2940 148.436
R974 GND.n3242 GND.n3237 148.436
R975 GND.n3399 GND.n3394 148.436
R976 GND.n4205 GND.n4200 148.436
R977 GND.n1496 GND.n1491 148.436
R978 GND.n197 GND.n192 148.436
R979 GND.n2003 GND.n1998 148.436
R980 GND.n349 GND.n344 148.436
R981 GND.n502 GND.n497 148.436
R982 GND.n7427 GND.n7386 148.436
R983 GND.n6561 GND.n6416 141.556
R984 GND.n5435 GND.t1398 140.822
R985 GND.n6735 GND 138.286
R986 GND.n4426 GND 138.286
R987 GND.t1368 GND.t164 138.035
R988 GND.n2034 GND.n2033 137.827
R989 GND.n6794 GND.n6793 137.55
R990 GND.t62 GND 133.766
R991 GND.n3547 GND.n3540 131.194
R992 GND GND.t66 130.352
R993 GND.n6658 GND.t452 129.006
R994 GND.n6876 GND.n4275 128.821
R995 GND.n4920 GND.t630 127.368
R996 GND.n4275 GND.t626 127.368
R997 GND.n6472 GND.t891 124.398
R998 GND.n6473 GND.t923 124.398
R999 GND.n2016 GND.t395 123.612
R1000 GND.n514 GND.t619 123.612
R1001 GND.n209 GND.t504 123.612
R1002 GND.n1508 GND.t75 123.612
R1003 GND.n1460 GND.t1253 123.612
R1004 GND.n4217 GND.t1364 123.612
R1005 GND.n3411 GND.t347 123.612
R1006 GND.n3254 GND.t366 123.612
R1007 GND.n2957 GND.t719 123.612
R1008 GND.n2632 GND.t480 123.612
R1009 GND.n2308 GND.t110 123.612
R1010 GND.n2146 GND.t92 123.612
R1011 GND.n1278 GND.t716 123.612
R1012 GND.n361 GND.t107 123.612
R1013 GND.n7409 GND.t1318 123.612
R1014 GND.n7364 GND.t823 123.612
R1015 GND.n2053 GND.n2052 123.472
R1016 GND.n1938 GND.n1937 121.112
R1017 GND.n1905 GND.n1904 121.112
R1018 GND.n1705 GND.n1704 121.112
R1019 GND.n1862 GND.n1861 121.112
R1020 GND.n6913 GND.n6912 121.112
R1021 GND.n6883 GND.n6882 121.112
R1022 GND.n2381 GND.n2380 121.112
R1023 GND.n2511 GND.n2510 121.112
R1024 GND.n2706 GND.n2705 121.112
R1025 GND.n2836 GND.n2835 121.112
R1026 GND.n3030 GND.n3029 121.112
R1027 GND.n3133 GND.n3132 121.112
R1028 GND.n7103 GND.n7102 121.112
R1029 GND.n7233 GND.n7232 121.112
R1030 GND.n4798 GND.n4797 121.112
R1031 GND.n4765 GND.n4764 121.112
R1032 GND.n5280 GND.n5279 121.112
R1033 GND.n5250 GND.n5249 121.112
R1034 GND.n5802 GND.n5801 121.112
R1035 GND.n5933 GND.n5932 121.112
R1036 GND.n5969 GND.n5968 121.112
R1037 GND.n6102 GND.n6101 121.112
R1038 GND.n6136 GND.n6135 121.112
R1039 GND.n6266 GND.n6265 121.112
R1040 GND.n6300 GND.n6299 121.112
R1041 GND.n6575 GND.n6574 121.112
R1042 GND.n588 GND.n587 121.112
R1043 GND.n715 GND.n714 121.112
R1044 GND.n7631 GND.n7630 121.112
R1045 GND.n7762 GND.n7761 121.112
R1046 GND.n7511 GND.n7510 121.112
R1047 GND.n7597 GND.n7596 121.112
R1048 GND.n1983 GND.t360 120.669
R1049 GND.t797 GND.n494 120.669
R1050 GND.t603 GND.n189 120.669
R1051 GND.t591 GND.n1524 120.669
R1052 GND.t690 GND.n1476 120.669
R1053 GND.t1172 GND.n4197 120.669
R1054 GND.t662 GND.n3391 120.669
R1055 GND.t1278 GND.n3234 120.669
R1056 GND.t430 GND.n2937 120.669
R1057 GND.t420 GND.n2612 120.669
R1058 GND.t807 GND.n2288 120.669
R1059 GND.t120 GND.n2126 120.669
R1060 GND.t87 GND.n1258 120.669
R1061 GND.t848 GND.n341 120.669
R1062 GND.t608 GND.n7425 120.669
R1063 GND.n7430 GND.t112 120.669
R1064 GND.t1451 GND.t1425 119.534
R1065 GND.t1409 GND.t1451 119.534
R1066 GND.t1429 GND.t1409 119.534
R1067 GND.t1421 GND.t1429 119.534
R1068 GND.t1443 GND.t1421 119.534
R1069 GND.t1411 GND.t1469 119.534
R1070 GND.t1447 GND.t1411 119.534
R1071 GND.t1517 GND.t1447 119.534
R1072 GND.t1413 GND.t1517 119.534
R1073 GND.t1437 GND.t1413 119.534
R1074 GND.t1501 GND.t1437 119.534
R1075 GND.t1403 GND.t1501 119.534
R1076 GND.t1463 GND.t1403 119.534
R1077 GND.t1507 GND.t1463 119.534
R1078 GND.t1495 GND.t1427 119.534
R1079 GND.t1521 GND.t1495 119.534
R1080 GND.t1419 GND.t1521 119.534
R1081 GND.t1475 GND.t1509 119.534
R1082 GND.t1509 GND.t1441 119.534
R1083 GND.t1441 GND.t1479 119.534
R1084 GND.t1479 GND.t1513 119.534
R1085 GND.t1513 GND.t1449 119.534
R1086 GND.t1449 GND.t1401 119.534
R1087 GND.t1401 GND.t1461 119.534
R1088 GND.t1461 GND.t1487 119.534
R1089 GND.t1487 GND.t1407 119.534
R1090 GND.t1407 GND.t1467 119.534
R1091 GND.t1467 GND.t1491 119.534
R1092 GND.t1415 GND.t1473 119.534
R1093 GND.t1473 GND.t1503 119.534
R1094 GND.t1503 GND.t1439 119.534
R1095 GND.t1439 GND.t1525 119.534
R1096 GND.t1499 GND.t1435 119.534
R1097 GND.t1527 GND.t1499 119.534
R1098 GND.t1457 GND.t1527 119.534
R1099 GND.t1483 GND.t1457 119.534
R1100 GND.t1515 GND.t1483 119.534
R1101 GND.t1459 GND.t1515 119.534
R1102 GND.t1485 GND.t1459 119.534
R1103 GND.t1431 GND.t1485 119.534
R1104 GND.t1453 GND.t1431 119.534
R1105 GND.t1471 GND.t1453 119.534
R1106 GND.t1519 GND.t1493 119.534
R1107 GND.t1417 GND.t1519 119.534
R1108 GND.t1497 GND.t1417 119.534
R1109 GND.t1523 GND.t1455 119.534
R1110 GND.t1455 GND.t1477 119.534
R1111 GND.t1477 GND.t1511 119.534
R1112 GND.t1511 GND.t1445 119.534
R1113 GND.t1445 GND.t1481 119.534
R1114 GND.t1481 GND.t1423 119.534
R1115 GND.t1423 GND.t1505 119.534
R1116 GND.t1505 GND.t1405 119.534
R1117 GND.t1405 GND.t1465 119.534
R1118 GND.t1465 GND.t1489 119.534
R1119 GND.t1489 GND.t1433 119.534
R1120 GND.t546 GND.t560 119.534
R1121 GND.t560 GND.t540 119.534
R1122 GND.t548 GND.t558 119.534
R1123 GND.t558 GND.t554 119.534
R1124 GND.t554 GND.t562 119.534
R1125 GND.t562 GND.t542 119.534
R1126 GND.t542 GND.t556 119.534
R1127 GND.t556 GND.t564 119.534
R1128 GND.t564 GND.t544 119.534
R1129 GND.t544 GND.t550 119.534
R1130 GND.t550 GND.t534 119.534
R1131 GND.t534 GND.t538 119.534
R1132 GND.t538 GND.t552 119.534
R1133 GND.t552 GND.t536 119.534
R1134 GND.t1154 GND.t1156 119.534
R1135 GND.t1156 GND.t1150 119.534
R1136 GND.t1150 GND.t1152 119.534
R1137 GND.t164 GND.t62 119.534
R1138 GND.t406 GND.t1119 119.285
R1139 GND.t154 GND.t668 119.109
R1140 GND.t20 GND.t795 119.109
R1141 GND.t140 GND.t73 119.109
R1142 GND.t90 GND.t404 119.109
R1143 GND.n6718 GND.n6717 118.1
R1144 GND.n5749 GND.n5748 118.1
R1145 GND.n5160 GND.n5159 118.1
R1146 GND.n5191 GND.n5190 117.984
R1147 GND.n4288 GND.n4287 117.984
R1148 GND.n6421 GND.t874 117.626
R1149 GND.n5512 GND.t1426 117.626
R1150 GND.n4437 GND.t1060 117.626
R1151 GND.n4580 GND.t237 117.007
R1152 GND.n5767 GND.t1523 116.689
R1153 GND.n3837 GND.n3836 116.329
R1154 GND.n5488 GND.n5487 116.052
R1155 GND.n4419 GND.n4418 116.052
R1156 GND GND.t1314 115.596
R1157 GND.n7538 GND.n7537 115.201
R1158 GND.n7669 GND.n7668 115.201
R1159 GND.n6376 GND.n6375 115.201
R1160 GND.n6212 GND.n6211 115.201
R1161 GND.n6048 GND.n6047 115.201
R1162 GND.n6006 GND.n6005 115.201
R1163 GND.n5823 GND.n5822 115.201
R1164 GND.n5301 GND.n5300 115.201
R1165 GND.n4860 GND.n4859 115.201
R1166 GND.n7167 GND.n7166 115.201
R1167 GND.n3067 GND.n3066 115.201
R1168 GND.n2743 GND.n2742 115.201
R1169 GND.n2418 GND.n2417 115.201
R1170 GND.n6934 GND.n6933 115.201
R1171 GND.n1769 GND.n1768 115.201
R1172 GND.n1578 GND.n1577 115.201
R1173 GND.n6705 GND.n6704 114.713
R1174 GND.n5492 GND.n5491 114.713
R1175 GND.n6665 GND.n6664 114.713
R1176 GND.n6671 GND.n6670 114.713
R1177 GND.n6675 GND.n6674 114.713
R1178 GND.n6681 GND.n6680 114.713
R1179 GND.n6687 GND.n6686 114.713
R1180 GND.n6693 GND.n6692 114.713
R1181 GND.n6608 GND.n6607 114.713
R1182 GND.n6652 GND.n6651 114.713
R1183 GND.n6645 GND.n6644 114.713
R1184 GND.n6641 GND.n6640 114.713
R1185 GND.n6635 GND.n6634 114.713
R1186 GND.n6629 GND.n6628 114.713
R1187 GND.n6623 GND.n6622 114.713
R1188 GND.n6518 GND.n6517 114.713
R1189 GND.n6525 GND.n6524 114.713
R1190 GND.n6551 GND.n6550 114.713
R1191 GND.n6547 GND.n6546 114.713
R1192 GND.n6541 GND.n6540 114.713
R1193 GND.n6535 GND.n6534 114.713
R1194 GND.n6529 GND.n6528 114.713
R1195 GND.n6434 GND.n6433 114.713
R1196 GND.n6477 GND.n6476 114.713
R1197 GND.n6484 GND.n6483 114.713
R1198 GND.n6488 GND.n6487 114.713
R1199 GND.n6494 GND.n6493 114.713
R1200 GND.n6500 GND.n6499 114.713
R1201 GND.n6506 GND.n6505 114.713
R1202 GND.n6420 GND.n6419 114.713
R1203 GND.n6425 GND.n6424 114.713
R1204 GND.n6467 GND.n6466 114.713
R1205 GND.n6462 GND.n6461 114.713
R1206 GND.n6456 GND.n6455 114.713
R1207 GND.n6450 GND.n6449 114.713
R1208 GND.n6444 GND.n6443 114.713
R1209 GND.n4966 GND.n4965 114.713
R1210 GND.n4653 GND.n4652 114.713
R1211 GND.n4647 GND.n4646 114.713
R1212 GND.n4641 GND.n4640 114.713
R1213 GND.n4637 GND.n4636 114.713
R1214 GND.n4610 GND.n4609 114.713
R1215 GND.n4672 GND.n4671 114.713
R1216 GND.n4678 GND.n4677 114.713
R1217 GND.n4690 GND.n4689 114.713
R1218 GND.n4696 GND.n4695 114.713
R1219 GND.n4703 GND.n4702 114.713
R1220 GND.n4744 GND.n4743 114.713
R1221 GND.n4737 GND.n4736 114.713
R1222 GND.n4731 GND.n4730 114.713
R1223 GND.n4725 GND.n4724 114.713
R1224 GND.n4715 GND.n4714 114.713
R1225 GND.n4709 GND.n4708 114.713
R1226 GND.n4925 GND.n4924 114.713
R1227 GND.n4930 GND.n4929 114.713
R1228 GND.n4937 GND.n4936 114.713
R1229 GND.n4943 GND.n4942 114.713
R1230 GND.n5033 GND.n5032 114.713
R1231 GND.n5022 GND.n5021 114.713
R1232 GND.n5012 GND.n5011 114.713
R1233 GND.n5005 GND.n5004 114.713
R1234 GND.n5001 GND.n5000 114.713
R1235 GND.n4995 GND.n4994 114.713
R1236 GND.n4989 GND.n4988 114.713
R1237 GND.n4982 GND.n4981 114.713
R1238 GND.n4583 GND.n4582 114.713
R1239 GND.n4591 GND.n4590 114.713
R1240 GND.n4597 GND.n4596 114.713
R1241 GND.n4601 GND.n4600 114.713
R1242 GND.n4614 GND.n4613 114.713
R1243 GND.n4620 GND.n4619 114.713
R1244 GND.n4626 GND.n4625 114.713
R1245 GND.n5736 GND.n5735 114.713
R1246 GND.n5688 GND.n5687 114.713
R1247 GND.n5696 GND.n5695 114.713
R1248 GND.n5702 GND.n5701 114.713
R1249 GND.n5706 GND.n5705 114.713
R1250 GND.n5712 GND.n5711 114.713
R1251 GND.n5718 GND.n5717 114.713
R1252 GND.n5724 GND.n5723 114.713
R1253 GND.n5774 GND.n5773 114.713
R1254 GND.n5504 GND.n5503 114.713
R1255 GND.n5653 GND.n5652 114.713
R1256 GND.n5657 GND.n5656 114.713
R1257 GND.n5663 GND.n5662 114.713
R1258 GND.n5669 GND.n5668 114.713
R1259 GND.n5675 GND.n5674 114.713
R1260 GND.n5610 GND.n5609 114.713
R1261 GND.n5617 GND.n5616 114.713
R1262 GND.n5639 GND.n5638 114.713
R1263 GND.n5635 GND.n5634 114.713
R1264 GND.n5629 GND.n5628 114.713
R1265 GND.n5623 GND.n5622 114.713
R1266 GND.n5498 GND.n5497 114.713
R1267 GND.n5526 GND.n5525 114.713
R1268 GND.n5569 GND.n5568 114.713
R1269 GND.n5576 GND.n5575 114.713
R1270 GND.n5580 GND.n5579 114.713
R1271 GND.n5586 GND.n5585 114.713
R1272 GND.n5592 GND.n5591 114.713
R1273 GND.n5598 GND.n5597 114.713
R1274 GND.n5511 GND.n5510 114.713
R1275 GND.n5516 GND.n5515 114.713
R1276 GND.n5559 GND.n5558 114.713
R1277 GND.n5554 GND.n5553 114.713
R1278 GND.n5548 GND.n5547 114.713
R1279 GND.n5542 GND.n5541 114.713
R1280 GND.n5536 GND.n5535 114.713
R1281 GND.n5147 GND.n5146 114.713
R1282 GND.n4428 GND.n4427 114.713
R1283 GND.n5107 GND.n5106 114.713
R1284 GND.n5113 GND.n5112 114.713
R1285 GND.n5117 GND.n5116 114.713
R1286 GND.n5123 GND.n5122 114.713
R1287 GND.n5129 GND.n5128 114.713
R1288 GND.n5135 GND.n5134 114.713
R1289 GND.n5050 GND.n5049 114.713
R1290 GND.n5094 GND.n5093 114.713
R1291 GND.n5087 GND.n5086 114.713
R1292 GND.n5083 GND.n5082 114.713
R1293 GND.n5077 GND.n5076 114.713
R1294 GND.n5071 GND.n5070 114.713
R1295 GND.n5065 GND.n5064 114.713
R1296 GND.n4498 GND.n4497 114.713
R1297 GND.n4432 GND.n4431 114.713
R1298 GND.n4550 GND.n4549 114.713
R1299 GND.n4554 GND.n4553 114.713
R1300 GND.n4560 GND.n4559 114.713
R1301 GND.n4566 GND.n4565 114.713
R1302 GND.n4572 GND.n4571 114.713
R1303 GND.n4486 GND.n4485 114.713
R1304 GND.n4537 GND.n4536 114.713
R1305 GND.n4530 GND.n4529 114.713
R1306 GND.n4526 GND.n4525 114.713
R1307 GND.n4520 GND.n4519 114.713
R1308 GND.n4514 GND.n4513 114.713
R1309 GND.n4508 GND.n4507 114.713
R1310 GND.n4436 GND.n4435 114.713
R1311 GND.n4441 GND.n4440 114.713
R1312 GND.n4451 GND.n4450 114.713
R1313 GND.n4456 GND.n4455 114.713
R1314 GND.n4462 GND.n4461 114.713
R1315 GND.n4468 GND.n4467 114.713
R1316 GND.n4474 GND.n4473 114.713
R1317 GND.n6615 GND.t451 113.734
R1318 GND.n6603 GND.t942 113.734
R1319 GND.n6513 GND.t864 113.734
R1320 GND.n6431 GND.t876 113.734
R1321 GND.n4659 GND.t223 113.734
R1322 GND.n4685 GND.t253 113.734
R1323 GND.n4707 GND.t271 113.734
R1324 GND.n4947 GND.t625 113.734
R1325 GND.n5682 GND.t547 113.734
R1326 GND.n5502 GND.t1494 113.734
R1327 GND.n5605 GND.t1416 113.734
R1328 GND.n5523 GND.t1428 113.734
R1329 GND.n5057 GND.t1563 113.734
R1330 GND.n5045 GND.t1000 113.734
R1331 GND.n4493 GND.t1050 113.734
R1332 GND.n4481 GND.t1062 113.734
R1333 GND.n6560 GND.t931 112.88
R1334 GND.n5480 GND.n5479 111.957
R1335 GND.n4411 GND.n4410 111.957
R1336 GND.n5449 GND.n5448 111.957
R1337 GND.n5451 GND.n5450 111.957
R1338 GND.n5235 GND.n5234 111.957
R1339 GND.n5240 GND.n5225 111.957
R1340 GND.n6854 GND.n6853 111.957
R1341 GND.n6856 GND.n6855 111.957
R1342 GND.n4327 GND.n4326 111.957
R1343 GND.n4332 GND.n4317 111.957
R1344 GND.n6712 GND.t785 111.924
R1345 GND.n4955 GND.t411 111.924
R1346 GND.n4952 GND.t667 111.924
R1347 GND.n5743 GND.t681 111.924
R1348 GND.n6806 GND.t1294 111.924
R1349 GND.n6807 GND.t475 111.924
R1350 GND.n6808 GND.t747 111.924
R1351 GND.n6809 GND.t23 111.924
R1352 GND.n6810 GND.t345 111.924
R1353 GND.n7051 GND.t698 111.924
R1354 GND.n7052 GND.t147 111.924
R1355 GND.n7053 GND.t1179 111.924
R1356 GND.n7054 GND.t803 111.924
R1357 GND.n7055 GND.t145 111.924
R1358 GND.n5154 GND.t67 111.924
R1359 GND.n6699 GND.t441 111.296
R1360 GND.n6614 GND.t882 111.296
R1361 GND.n6602 GND.t920 111.296
R1362 GND.n6512 GND.t940 111.296
R1363 GND.n6430 GND.t956 111.296
R1364 GND.n4660 GND.t295 111.296
R1365 GND.n4683 GND.t219 111.296
R1366 GND.n4706 GND.t217 111.296
R1367 GND.n4946 GND.t241 111.296
R1368 GND.n4948 GND.t635 111.296
R1369 GND.n5730 GND.t537 111.296
R1370 GND.n5681 GND.t1434 111.296
R1371 GND.n5501 GND.t1472 111.296
R1372 GND.n5604 GND.t1492 111.296
R1373 GND.n5522 GND.t1508 111.296
R1374 GND.n5141 GND.t1553 111.296
R1375 GND.n5056 GND.t1068 111.296
R1376 GND.n5044 GND.t1106 111.296
R1377 GND.n4492 GND.t998 111.296
R1378 GND.n4480 GND.t1014 111.296
R1379 GND GND.t1507 110.996
R1380 GND.t1491 GND 110.996
R1381 GND GND.t1471 110.996
R1382 GND.t1433 GND 110.996
R1383 GND.t536 GND 110.996
R1384 GND.n5220 GND.n5219 110.841
R1385 GND.n7360 GND.n7359 109.394
R1386 GND.n2013 GND.n2012 109.394
R1387 GND.n511 GND.n510 109.394
R1388 GND.n206 GND.n205 109.394
R1389 GND.n1505 GND.n1504 109.394
R1390 GND.n1457 GND.n1456 109.394
R1391 GND.n4214 GND.n4213 109.394
R1392 GND.n3408 GND.n3407 109.394
R1393 GND.n3251 GND.n3250 109.394
R1394 GND.n2954 GND.n2953 109.394
R1395 GND.n2629 GND.n2628 109.394
R1396 GND.n2305 GND.n2304 109.394
R1397 GND.n2143 GND.n2142 109.394
R1398 GND.n1275 GND.n1274 109.394
R1399 GND.n358 GND.n357 109.394
R1400 GND.n7406 GND.n7405 109.394
R1401 GND.n5470 GND.n5469 109.359
R1402 GND.n4401 GND.n4400 109.359
R1403 GND.n6773 GND.n6772 109.314
R1404 GND.n5230 GND.n5229 109.314
R1405 GND.n4351 GND.n4350 109.314
R1406 GND.n4322 GND.n4321 109.314
R1407 GND.n6742 GND.t1274 108.505
R1408 GND.n6739 GND.t1273 108.505
R1409 GND.n6769 GND.t1303 108.505
R1410 GND.n6766 GND.t1301 108.505
R1411 GND.n4381 GND.t677 108.505
R1412 GND.n4378 GND.t679 108.505
R1413 GND.n4347 GND.t700 108.505
R1414 GND.n4344 GND.t704 108.505
R1415 GND.n5472 GND.n5471 108.016
R1416 GND.n4403 GND.n4402 108.016
R1417 GND.n6774 GND.n6771 108.016
R1418 GND.n5228 GND.n5227 108.016
R1419 GND.n5207 GND.n5206 108.016
R1420 GND.n5211 GND.n5181 108.016
R1421 GND.n5187 GND.n5186 108.016
R1422 GND.n4352 GND.n4349 108.016
R1423 GND.n4320 GND.n4319 108.016
R1424 GND.n4304 GND.n4303 108.016
R1425 GND.n4308 GND.n4278 108.016
R1426 GND.n4284 GND.n4283 108.016
R1427 GND.n7374 GND.n7373 107.24
R1428 GND.n1370 GND.n1369 107.24
R1429 GND.n327 GND.n326 107.24
R1430 GND.n480 GND.n479 107.24
R1431 GND.n175 GND.n174 107.24
R1432 GND.n1484 GND.n1483 107.24
R1433 GND.n1383 GND.n1382 107.24
R1434 GND.n4183 GND.n4182 107.24
R1435 GND.n3377 GND.n3376 107.24
R1436 GND.n3220 GND.n3219 107.24
R1437 GND.n2923 GND.n2922 107.24
R1438 GND.n2598 GND.n2597 107.24
R1439 GND.n2274 GND.n2273 107.24
R1440 GND.n2112 GND.n2111 107.24
R1441 GND.n1244 GND.n1243 107.24
R1442 GND.n7392 GND.n7391 107.24
R1443 GND.t1152 GND 106.728
R1444 GND.n5204 GND.n5203 105.975
R1445 GND.n5184 GND.n5183 105.975
R1446 GND.n5194 GND.n5189 105.975
R1447 GND.n4301 GND.n4300 105.975
R1448 GND.n4281 GND.n4280 105.975
R1449 GND.n4291 GND.n4286 105.975
R1450 GND.t1435 GND.n5647 105.305
R1451 GND.n4914 GND.t1293 103.51
R1452 GND.t1085 GND.t1059 103.299
R1453 GND.t1043 GND.t1085 103.299
R1454 GND.t1063 GND.t1043 103.299
R1455 GND.t1055 GND.t1063 103.299
R1456 GND.t1077 GND.t1055 103.299
R1457 GND.t1103 GND.t1045 103.299
R1458 GND.t1045 GND.t1081 103.299
R1459 GND.t1081 GND.t1023 103.299
R1460 GND.t1023 GND.t1047 103.299
R1461 GND.t1047 GND.t1071 103.299
R1462 GND.t1071 GND.t1007 103.299
R1463 GND.t1007 GND.t1037 103.299
R1464 GND.t1037 GND.t1097 103.299
R1465 GND.t1097 GND.t1013 103.299
R1466 GND.t1061 GND.t1001 103.299
R1467 GND.t1001 GND.t1027 103.299
R1468 GND.t1027 GND.t1053 103.299
R1469 GND.t1015 GND.t1109 103.299
R1470 GND.t1075 GND.t1015 103.299
R1471 GND.t1113 GND.t1075 103.299
R1472 GND.t1019 GND.t1113 103.299
R1473 GND.t1083 GND.t1019 103.299
R1474 GND.t1035 GND.t1083 103.299
R1475 GND.t1095 GND.t1035 103.299
R1476 GND.t993 GND.t1095 103.299
R1477 GND.t1041 GND.t993 103.299
R1478 GND.t1101 GND.t1041 103.299
R1479 GND.t997 GND.t1101 103.299
R1480 GND.t1107 GND.t1049 103.299
R1481 GND.t1009 GND.t1107 103.299
R1482 GND.t1073 GND.t1009 103.299
R1483 GND.t1031 GND.t1073 103.299
R1484 GND.t1069 GND.t1005 103.299
R1485 GND.t1005 GND.t1033 103.299
R1486 GND.t1033 GND.t1091 103.299
R1487 GND.t1091 GND.t989 103.299
R1488 GND.t989 GND.t1021 103.299
R1489 GND.t1021 GND.t1093 103.299
R1490 GND.t1093 GND.t991 103.299
R1491 GND.t991 GND.t1065 103.299
R1492 GND.t1065 GND.t1087 103.299
R1493 GND.t1087 GND.t1105 103.299
R1494 GND.t999 GND.t1025 103.299
R1495 GND.t1025 GND.t1051 103.299
R1496 GND.t1051 GND.t1003 103.299
R1497 GND.t1089 GND.t1029 103.299
R1498 GND.t1111 GND.t1089 103.299
R1499 GND.t1017 GND.t1111 103.299
R1500 GND.t1079 GND.t1017 103.299
R1501 GND.t987 GND.t1079 103.299
R1502 GND.t1057 GND.t987 103.299
R1503 GND.t1011 GND.t1057 103.299
R1504 GND.t1039 GND.t1011 103.299
R1505 GND.t1099 GND.t1039 103.299
R1506 GND.t995 GND.t1099 103.299
R1507 GND.t1067 GND.t995 103.299
R1508 GND.t1544 GND.t1562 103.299
R1509 GND.t1556 GND.t1544 103.299
R1510 GND.t1564 GND.t1542 103.299
R1511 GND.t1542 GND.t1538 103.299
R1512 GND.t1538 GND.t1546 103.299
R1513 GND.t1546 GND.t1558 103.299
R1514 GND.t1558 GND.t1540 103.299
R1515 GND.t1540 GND.t1548 103.299
R1516 GND.t1548 GND.t1560 103.299
R1517 GND.t1560 GND.t1534 103.299
R1518 GND.t1534 GND.t1550 103.299
R1519 GND.t1550 GND.t1554 103.299
R1520 GND.t1554 GND.t1536 103.299
R1521 GND.t1536 GND.t1552 103.299
R1522 GND.t83 GND.t85 103.299
R1523 GND.t85 GND.t79 103.299
R1524 GND.t79 GND.t81 103.299
R1525 GND.t1314 GND.t406 103.299
R1526 GND.n1992 GND.n1991 101.948
R1527 GND.n5487 GND.t1298 101.43
R1528 GND.n4418 GND.t707 101.43
R1529 GND.n7793 GND.n7786 100.894
R1530 GND.n854 GND.n845 100.894
R1531 GND.n747 GND.n738 100.894
R1532 GND.n428 GND.n419 100.894
R1533 GND.n1638 GND.n1629 100.894
R1534 GND.n275 GND.n266 100.894
R1535 GND.n123 GND.n114 100.894
R1536 GND.n14 GND.n5 100.894
R1537 GND.n7270 GND.n7261 100.894
R1538 GND.n3480 GND.n3471 100.894
R1539 GND.n3322 GND.n3313 100.894
R1540 GND.n3165 GND.n3156 100.894
R1541 GND.n2868 GND.n2859 100.894
R1542 GND.n2543 GND.n2534 100.894
R1543 GND.n2219 GND.n2210 100.894
R1544 GND.n1194 GND.n1185 100.894
R1545 GND.n1980 GND.n1526 100.692
R1546 GND GND.t474 98.3051
R1547 GND GND.t746 98.3051
R1548 GND GND.t344 98.3051
R1549 GND GND.t22 97.1486
R1550 GND.t1013 GND 95.92
R1551 GND GND.t997 95.92
R1552 GND.t1105 GND 95.92
R1553 GND.t1029 GND.n5099 95.92
R1554 GND GND.t1067 95.92
R1555 GND.t1552 GND 95.92
R1556 GND.t254 GND.t236 93.8076
R1557 GND.t326 GND.t226 93.8076
R1558 GND.t226 GND.t276 93.8076
R1559 GND.t276 GND.t312 93.8076
R1560 GND.t312 GND.t230 93.8076
R1561 GND.t230 GND.t280 93.8076
R1562 GND.t280 GND.t316 93.8076
R1563 GND.t338 GND.t304 93.8076
R1564 GND.t234 GND.t338 93.8076
R1565 GND.t310 GND.t234 93.8076
R1566 GND.t342 GND.t310 93.8076
R1567 GND.t268 GND.t342 93.8076
R1568 GND.t272 GND.t222 93.8076
R1569 GND.t306 GND.t272 93.8076
R1570 GND.t258 GND.t306 93.8076
R1571 GND.t220 GND.t258 93.8076
R1572 GND.t244 GND.t220 93.8076
R1573 GND.t300 GND.t244 93.8076
R1574 GND.t332 GND.t300 93.8076
R1575 GND.t232 GND.t332 93.8076
R1576 GND.t284 GND.t232 93.8076
R1577 GND.t336 GND.t284 93.8076
R1578 GND.t262 GND.t288 93.8076
R1579 GND.t288 GND.t320 93.8076
R1580 GND.t320 GND.t256 93.8076
R1581 GND.t256 GND.t218 93.8076
R1582 GND.t252 GND.t324 93.8076
R1583 GND.t324 GND.t238 93.8076
R1584 GND.t238 GND.t296 93.8076
R1585 GND.t296 GND.t328 93.8076
R1586 GND.t328 GND.t228 93.8076
R1587 GND.t228 GND.t278 93.8076
R1588 GND.t250 GND.t314 93.8076
R1589 GND.t282 GND.t250 93.8076
R1590 GND.t248 GND.t282 93.8076
R1591 GND.t308 GND.t248 93.8076
R1592 GND.t340 GND.t308 93.8076
R1593 GND.t266 GND.t340 93.8076
R1594 GND.t292 GND.t266 93.8076
R1595 GND.t216 GND.t292 93.8076
R1596 GND.t322 GND.t270 93.8076
R1597 GND.t224 GND.t322 93.8076
R1598 GND.t274 GND.t224 93.8076
R1599 GND.t242 GND.t274 93.8076
R1600 GND.t298 GND.t242 93.8076
R1601 GND.t330 GND.t246 93.8076
R1602 GND.t246 GND.t302 93.8076
R1603 GND.t302 GND.t334 93.8076
R1604 GND.t334 GND.t260 93.8076
R1605 GND.t260 GND.t286 93.8076
R1606 GND.t286 GND.t318 93.8076
R1607 GND.t318 GND.t264 93.8076
R1608 GND.t264 GND.t290 93.8076
R1609 GND.t290 GND.t240 93.8076
R1610 GND.t81 GND 92.2308
R1611 GND.t1255 GND.t114 91.9116
R1612 GND.n7808 GND.n7805 91.8593
R1613 GND.n871 GND.n868 91.8593
R1614 GND.n764 GND.n761 91.8593
R1615 GND.n445 GND.n442 91.8593
R1616 GND.n1655 GND.n1652 91.8593
R1617 GND.n292 GND.n289 91.8593
R1618 GND.n140 GND.n137 91.8593
R1619 GND.n31 GND.n28 91.8593
R1620 GND.n7287 GND.n7284 91.8593
R1621 GND.n3497 GND.n3494 91.8593
R1622 GND.n3339 GND.n3336 91.8593
R1623 GND.n3182 GND.n3179 91.8593
R1624 GND.n2885 GND.n2882 91.8593
R1625 GND.n2560 GND.n2557 91.8593
R1626 GND.n2236 GND.n2233 91.8593
R1627 GND.n1211 GND.n1208 91.8593
R1628 GND.n7562 GND.n7561 90.3534
R1629 GND.n7693 GND.n7692 90.3534
R1630 GND.n646 GND.n645 90.3534
R1631 GND.n6358 GND.n6357 90.3534
R1632 GND.n6194 GND.n6193 90.3534
R1633 GND.n6030 GND.n6029 90.3534
R1634 GND.n5847 GND.n5846 90.3534
R1635 GND.n5325 GND.n5324 90.3534
R1636 GND.n4884 GND.n4883 90.3534
R1637 GND.n7191 GND.n7190 90.3534
R1638 GND.n3091 GND.n3090 90.3534
R1639 GND.n2767 GND.n2766 90.3534
R1640 GND.n2442 GND.n2441 90.3534
R1641 GND.n6958 GND.n6957 90.3534
R1642 GND.n1793 GND.n1792 90.3534
R1643 GND.n1602 GND.n1601 90.3534
R1644 GND.n1548 GND.n1547 90.3427
R1645 GND.n1566 GND.n1565 90.3427
R1646 GND.n1757 GND.n1756 90.3427
R1647 GND.n6922 GND.n6921 90.3427
R1648 GND.n2406 GND.n2405 90.3427
R1649 GND.n2731 GND.n2730 90.3427
R1650 GND.n3055 GND.n3054 90.3427
R1651 GND.n7155 GND.n7154 90.3427
R1652 GND.n4848 GND.n4847 90.3427
R1653 GND.n5289 GND.n5288 90.3427
R1654 GND.n5811 GND.n5810 90.3427
R1655 GND.n5994 GND.n5993 90.3427
R1656 GND.n6161 GND.n6160 90.3427
R1657 GND.n6325 GND.n6324 90.3427
R1658 GND.n613 GND.n612 90.3427
R1659 GND.n7657 GND.n7656 90.3427
R1660 GND.n6734 GND 87.5398
R1661 GND.n4664 GND.t268 87.1071
R1662 GND GND.t294 87.1071
R1663 GND.t218 GND 87.1071
R1664 GND GND.t216 87.1071
R1665 GND.t240 GND 87.1071
R1666 GND.n1558 GND.n1557 86.1558
R1667 GND.n1747 GND.n1746 86.1558
R1668 GND.n7019 GND.n7018 86.1558
R1669 GND.n2396 GND.n2395 86.1558
R1670 GND.n2721 GND.n2720 86.1558
R1671 GND.n3045 GND.n3044 86.1558
R1672 GND.n7145 GND.n7144 86.1558
R1673 GND.n4838 GND.n4837 86.1558
R1674 GND.n5414 GND.n5413 86.1558
R1675 GND.n5909 GND.n5908 86.1558
R1676 GND.n5984 GND.n5983 86.1558
R1677 GND.n6151 GND.n6150 86.1558
R1678 GND.n6315 GND.n6314 86.1558
R1679 GND.n603 GND.n602 86.1558
R1680 GND.n7646 GND.n7645 86.1558
R1681 GND.n7526 GND.n7525 86.1558
R1682 GND.n7581 GND.n7580 86.1558
R1683 GND.n7745 GND.n7744 86.1558
R1684 GND.n698 GND.n697 86.1558
R1685 GND.n6413 GND.n6412 86.1558
R1686 GND.n6249 GND.n6248 86.1558
R1687 GND.n6085 GND.n6084 86.1558
R1688 GND.n5899 GND.n5898 86.1558
R1689 GND.n5377 GND.n5376 86.1558
R1690 GND.n4909 GND.n4908 86.1558
R1691 GND.n7216 GND.n7215 86.1558
R1692 GND.n3116 GND.n3115 86.1558
R1693 GND.n2819 GND.n2818 86.1558
R1694 GND.n2494 GND.n2493 86.1558
R1695 GND.n7009 GND.n7008 86.1558
R1696 GND.n1845 GND.n1844 86.1558
R1697 GND.n1888 GND.n1887 86.1558
R1698 GND.n4543 GND.t1069 86.0821
R1699 GND.n5766 GND.t548 85.3821
R1700 GND.n1203 GND.n1200 83.5572
R1701 GND.n2228 GND.n2225 83.5572
R1702 GND.n2552 GND.n2549 83.5572
R1703 GND.n2877 GND.n2874 83.5572
R1704 GND.n3174 GND.n3171 83.5572
R1705 GND.n3331 GND.n3328 83.5572
R1706 GND.n3489 GND.n3486 83.5572
R1707 GND.n7279 GND.n7276 83.5572
R1708 GND.n23 GND.n20 83.5572
R1709 GND.n132 GND.n129 83.5572
R1710 GND.n284 GND.n281 83.5572
R1711 GND.n1647 GND.n1644 83.5572
R1712 GND.n437 GND.n434 83.5572
R1713 GND.n756 GND.n753 83.5572
R1714 GND.n863 GND.n860 83.5572
R1715 GND.n5565 GND.t1475 82.5361
R1716 GND.n2135 GND.n2106 81.2313
R1717 GND.n2621 GND.n2592 81.2313
R1718 GND.n3243 GND.n3214 81.2313
R1719 GND.n4206 GND.n4177 81.2313
R1720 GND.n198 GND.n169 81.2313
R1721 GND.n503 GND.n474 81.2313
R1722 GND.n6560 GND.t963 80.6288
R1723 GND.n4665 GND.t262 80.4066
R1724 GND.n1980 GND.n1529 79.3342
R1725 GND.n7788 GND.n7787 78.6829
R1726 GND.n2033 GND.n2032 78.6829
R1727 GND.n7482 GND.n7481 74.9181
R1728 GND.n2070 GND.n2069 74.9181
R1729 GND.n402 GND.n401 74.9181
R1730 GND.n559 GND.n558 74.9181
R1731 GND.n250 GND.n249 74.9181
R1732 GND.n98 GND.n97 74.9181
R1733 GND.n1431 GND.n1430 74.9181
R1734 GND.n4258 GND.n4257 74.9181
R1735 GND.n3455 GND.n3454 74.9181
R1736 GND.n3297 GND.n3296 74.9181
R1737 GND.n3001 GND.n3000 74.9181
R1738 GND.n2677 GND.n2676 74.9181
R1739 GND.n2352 GND.n2351 74.9181
R1740 GND.n2194 GND.n2193 74.9181
R1741 GND.n1311 GND.n1310 74.9181
R1742 GND.n828 GND.n827 74.9181
R1743 GND.t174 GND.t1276 73.7614
R1744 GND.t699 GND.t856 73.7614
R1745 GND.n5479 GND.t1336 72.8576
R1746 GND.n4410 GND.t1224 72.8576
R1747 GND.n5448 GND.t1139 72.8576
R1748 GND.n5450 GND.t477 72.8576
R1749 GND.n5234 GND.t1133 72.8576
R1750 GND.n5225 GND.t1 72.8576
R1751 GND.n5190 GND.t1300 72.8576
R1752 GND.n6853 GND.t516 72.8576
R1753 GND.n6855 GND.t660 72.8576
R1754 GND.n4326 GND.t1177 72.8576
R1755 GND.n4317 GND.t1181 72.8576
R1756 GND.n4287 GND.t702 72.8576
R1757 GND.t77 GND.t123 72.82
R1758 GND.t24 GND.t59 72.82
R1759 GND.t122 GND.t33 72.82
R1760 GND.t214 GND.t106 72.82
R1761 GND.t394 GND.t78 72.82
R1762 GND.n5177 GND 72.2501
R1763 GND.n6875 GND 72.2501
R1764 GND.t436 GND.n7661 71.7802
R1765 GND.t200 GND.n617 71.7802
R1766 GND.t187 GND.n6329 71.7802
R1767 GND.t156 GND.n6165 71.7802
R1768 GND.t170 GND.n5998 71.7802
R1769 GND.t31 GND.n5815 71.7802
R1770 GND.t821 GND.n5293 71.7802
R1771 GND.t526 GND.n4852 71.7802
R1772 GND.t183 GND.n7159 71.7802
R1773 GND.t583 GND.n3059 71.7802
R1774 GND.t851 GND.n2735 71.7802
R1775 GND.t1196 GND.n2410 71.7802
R1776 GND.t654 GND.n6926 71.7802
R1777 GND.t782 GND.n1761 71.7802
R1778 GND.t374 GND.n1570 71.7802
R1779 GND.n5564 GND.t1443 71.1519
R1780 GND.n7452 GND.n7442 70.024
R1781 GND.n7448 GND.n7447 70.024
R1782 GND.n1033 GND.n1031 70.024
R1783 GND.n1033 GND.n1032 70.024
R1784 GND.n1037 GND.n1036 70.024
R1785 GND.n1343 GND.n1342 70.024
R1786 GND.n1348 GND.n1346 70.024
R1787 GND.n1348 GND.n1347 70.024
R1788 GND.n2035 GND.n2034 70.024
R1789 GND.n2039 GND.n2024 70.024
R1790 GND.n1012 GND.n1011 70.024
R1791 GND.n1022 GND.n1021 70.024
R1792 GND.n1018 GND.n1016 70.024
R1793 GND.n1018 GND.n1017 70.024
R1794 GND.n528 GND.n527 70.024
R1795 GND.n532 GND.n522 70.024
R1796 GND.n227 GND.n217 70.024
R1797 GND.n223 GND.n222 70.024
R1798 GND.n997 GND.n996 70.024
R1799 GND.n1002 GND.n1000 70.024
R1800 GND.n1002 GND.n1001 70.024
R1801 GND.n992 GND.n991 70.024
R1802 GND.n986 GND.n984 70.024
R1803 GND.n986 GND.n985 70.024
R1804 GND.n61 GND.n58 70.024
R1805 GND.n66 GND.n62 70.024
R1806 GND.n977 GND.n976 70.024
R1807 GND.n972 GND.n970 70.024
R1808 GND.n972 GND.n971 70.024
R1809 GND.n1397 GND.n1396 70.024
R1810 GND.n1401 GND.n1391 70.024
R1811 GND.n4235 GND.n4225 70.024
R1812 GND.n4231 GND.n4230 70.024
R1813 GND.n963 GND.n961 70.024
R1814 GND.n963 GND.n962 70.024
R1815 GND.n967 GND.n966 70.024
R1816 GND.n957 GND.n955 70.024
R1817 GND.n957 GND.n956 70.024
R1818 GND.n952 GND.n951 70.024
R1819 GND.n3425 GND.n3424 70.024
R1820 GND.n3429 GND.n3419 70.024
R1821 GND.n3272 GND.n3262 70.024
R1822 GND.n3268 GND.n3267 70.024
R1823 GND.n942 GND.n940 70.024
R1824 GND.n942 GND.n941 70.024
R1825 GND.n947 GND.n946 70.024
R1826 GND.n937 GND.n936 70.024
R1827 GND.n933 GND.n931 70.024
R1828 GND.n933 GND.n932 70.024
R1829 GND.n2971 GND.n2970 70.024
R1830 GND.n2975 GND.n2965 70.024
R1831 GND.n2650 GND.n2640 70.024
R1832 GND.n2646 GND.n2645 70.024
R1833 GND.n922 GND.n920 70.024
R1834 GND.n922 GND.n921 70.024
R1835 GND.n927 GND.n926 70.024
R1836 GND.n917 GND.n915 70.024
R1837 GND.n917 GND.n916 70.024
R1838 GND.n911 GND.n910 70.024
R1839 GND.n2322 GND.n2321 70.024
R1840 GND.n2326 GND.n2316 70.024
R1841 GND.n2164 GND.n2154 70.024
R1842 GND.n2160 GND.n2159 70.024
R1843 GND.n902 GND.n900 70.024
R1844 GND.n902 GND.n901 70.024
R1845 GND.n907 GND.n906 70.024
R1846 GND.n1296 GND.n1286 70.024
R1847 GND.n1292 GND.n1291 70.024
R1848 GND.n1338 GND.n1337 70.024
R1849 GND.n1333 GND.n1331 70.024
R1850 GND.n1333 GND.n1332 70.024
R1851 GND.n1008 GND.n1006 70.024
R1852 GND.n1008 GND.n1007 70.024
R1853 GND.n375 GND.n374 70.024
R1854 GND.n379 GND.n369 70.024
R1855 GND.n1042 GND.n1040 70.024
R1856 GND.n1042 GND.n1041 70.024
R1857 GND.n1027 GND.n1026 70.024
R1858 GND.n800 GND.n799 70.024
R1859 GND.n804 GND.n794 70.024
R1860 GND.t917 GND.n6472 69.1104
R1861 GND.n6473 GND.t867 69.1104
R1862 GND.n5100 GND.t1564 68.8658
R1863 GND.n5436 GND.n5435 68.1084
R1864 GND.n6743 GND.n6742 67.973
R1865 GND.n6740 GND.n6739 67.973
R1866 GND.n6780 GND.n6769 67.973
R1867 GND.n6767 GND.n6766 67.973
R1868 GND.n4382 GND.n4381 67.973
R1869 GND.n4379 GND.n4378 67.973
R1870 GND.n4358 GND.n4347 67.973
R1871 GND.n4345 GND.n4344 67.973
R1872 GND.n2063 GND.n2062 67.5205
R1873 GND.n1674 GND.n1673 67.5205
R1874 GND.n4578 GND.t254 67.0056
R1875 GND.n4447 GND.t1077 66.4063
R1876 GND.t1109 GND.n4542 66.4063
R1877 GND.n4921 GND.t298 64.7721
R1878 GND.n6658 GND.t444 64.5031
R1879 GND.n1981 GND.n1980 64.3169
R1880 GND.t1293 GND 61.2963
R1881 GND.t474 GND 61.2963
R1882 GND.t746 GND 61.2963
R1883 GND.t22 GND 61.2963
R1884 GND.t344 GND 61.2963
R1885 GND.n1544 GND.n1543 59.4829
R1886 GND.n1608 GND.n1607 59.4829
R1887 GND.n1799 GND.n1798 59.4829
R1888 GND.n6964 GND.n6963 59.4829
R1889 GND.n2448 GND.n2447 59.4829
R1890 GND.n2773 GND.n2772 59.4829
R1891 GND.n3097 GND.n3096 59.4829
R1892 GND.n7197 GND.n7196 59.4829
R1893 GND.n4890 GND.n4889 59.4829
R1894 GND.n5331 GND.n5330 59.4829
R1895 GND.n5853 GND.n5852 59.4829
R1896 GND.n6036 GND.n6035 59.4829
R1897 GND.n6200 GND.n6199 59.4829
R1898 GND.n6364 GND.n6363 59.4829
R1899 GND.n652 GND.n651 59.4829
R1900 GND.n7699 GND.n7698 59.4829
R1901 GND.n67 GND.n61 57.977
R1902 GND.t153 GND.t168 57.8291
R1903 GND.t185 GND.t390 57.8291
R1904 GND.t528 GND.t117 57.8291
R1905 GND.t678 GND.t1384 57.8291
R1906 GND.n7459 GND.n7452 57.224
R1907 GND.n2046 GND.n2039 57.224
R1908 GND.n539 GND.n532 57.224
R1909 GND.n234 GND.n227 57.224
R1910 GND.n67 GND.n66 57.224
R1911 GND.n1408 GND.n1401 57.224
R1912 GND.n4242 GND.n4235 57.224
R1913 GND.n3436 GND.n3429 57.224
R1914 GND.n3279 GND.n3272 57.224
R1915 GND.n2982 GND.n2975 57.224
R1916 GND.n2657 GND.n2650 57.224
R1917 GND.n2333 GND.n2326 57.224
R1918 GND.n2171 GND.n2164 57.224
R1919 GND.n1303 GND.n1296 57.224
R1920 GND.n386 GND.n379 57.224
R1921 GND.n811 GND.n804 57.224
R1922 GND.t624 GND.n4920 56.9548
R1923 GND.n6717 GND.t576 55.7148
R1924 GND.n5748 GND.t165 55.7148
R1925 GND.n5159 GND.t407 55.7148
R1926 GND.n2030 GND.n2029 54.813
R1927 GND.n7567 GND.n7562 54.66
R1928 GND.n7703 GND.n7693 54.66
R1929 GND.n656 GND.n646 54.66
R1930 GND.n6368 GND.n6358 54.66
R1931 GND.n6204 GND.n6194 54.66
R1932 GND.n6040 GND.n6030 54.66
R1933 GND.n5857 GND.n5847 54.66
R1934 GND.n5335 GND.n5325 54.66
R1935 GND.n4894 GND.n4884 54.66
R1936 GND.n7201 GND.n7191 54.66
R1937 GND.n3101 GND.n3091 54.66
R1938 GND.n2777 GND.n2767 54.66
R1939 GND.n2452 GND.n2442 54.66
R1940 GND.n6968 GND.n6958 54.66
R1941 GND.n1803 GND.n1793 54.66
R1942 GND.n1612 GND.n1602 54.66
R1943 GND.t14 GND.t738 54.5194
R1944 GND.n5490 GND 54.5194
R1945 GND.t175 GND.t149 54.5194
R1946 GND.n4916 GND 54.5194
R1947 GND.n5015 GND.t650 54.0356
R1948 GND.t314 GND.n4749 53.6046
R1949 GND.t384 GND.n1350 52.9309
R1950 GND.n2093 GND.t384 52.9309
R1951 GND.n5469 GND.t1531 52.8576
R1952 GND.n4400 GND.t425 52.8576
R1953 GND.n6772 GND.t15 52.8576
R1954 GND.n5229 GND.t1210 52.8576
R1955 GND.n5203 GND.t21 52.8576
R1956 GND.n5183 GND.t1140 52.8576
R1957 GND.n5189 GND.t116 52.8576
R1958 GND.n4350 GND.t1388 52.8576
R1959 GND.n4321 GND.t787 52.8576
R1960 GND.n4300 GND.t1180 52.8576
R1961 GND.n4280 GND.t523 52.8576
R1962 GND.n4286 GND.t152 52.8576
R1963 GND.n1980 GND.n1527 51.4154
R1964 GND.n1980 GND.n1528 51.4154
R1965 GND.n1980 GND.n1530 51.4154
R1966 GND.n1980 GND.n1531 51.4154
R1967 GND.n1980 GND.n1532 51.4154
R1968 GND.n1980 GND.n1533 51.4154
R1969 GND.n1980 GND.n1534 51.4154
R1970 GND.n1980 GND.n1535 51.4154
R1971 GND.n1980 GND.n1536 51.4154
R1972 GND.n1980 GND.n1537 51.4154
R1973 GND.n1980 GND.n1538 51.4154
R1974 GND.n1980 GND.n1539 51.4154
R1975 GND.n7814 GND.n7813 50.5605
R1976 GND.n884 GND.n882 50.5605
R1977 GND.n884 GND.n883 50.5605
R1978 GND.n1662 GND.n1660 50.5605
R1979 GND.n1662 GND.n1661 50.5605
R1980 GND.n2062 GND.n2061 50.5605
R1981 GND.n452 GND.n450 50.5605
R1982 GND.n452 GND.n451 50.5605
R1983 GND.n771 GND.n769 50.5605
R1984 GND.n771 GND.n770 50.5605
R1985 GND.n458 GND.n456 50.5605
R1986 GND.n458 GND.n457 50.5605
R1987 GND.n299 GND.n297 50.5605
R1988 GND.n299 GND.n298 50.5605
R1989 GND.n153 GND.n151 50.5605
R1990 GND.n153 GND.n152 50.5605
R1991 GND.n147 GND.n145 50.5605
R1992 GND.n147 GND.n146 50.5605
R1993 GND.n44 GND.n42 50.5605
R1994 GND.n44 GND.n43 50.5605
R1995 GND.n38 GND.n36 50.5605
R1996 GND.n38 GND.n37 50.5605
R1997 GND.n7300 GND.n7298 50.5605
R1998 GND.n7300 GND.n7299 50.5605
R1999 GND.n7294 GND.n7292 50.5605
R2000 GND.n7294 GND.n7293 50.5605
R2001 GND.n3510 GND.n3508 50.5605
R2002 GND.n3510 GND.n3509 50.5605
R2003 GND.n3504 GND.n3502 50.5605
R2004 GND.n3504 GND.n3503 50.5605
R2005 GND.n3352 GND.n3350 50.5605
R2006 GND.n3352 GND.n3351 50.5605
R2007 GND.n3346 GND.n3344 50.5605
R2008 GND.n3346 GND.n3345 50.5605
R2009 GND.n3195 GND.n3193 50.5605
R2010 GND.n3195 GND.n3194 50.5605
R2011 GND.n3189 GND.n3187 50.5605
R2012 GND.n3189 GND.n3188 50.5605
R2013 GND.n2898 GND.n2896 50.5605
R2014 GND.n2898 GND.n2897 50.5605
R2015 GND.n2892 GND.n2890 50.5605
R2016 GND.n2892 GND.n2891 50.5605
R2017 GND.n2573 GND.n2571 50.5605
R2018 GND.n2573 GND.n2572 50.5605
R2019 GND.n2567 GND.n2565 50.5605
R2020 GND.n2567 GND.n2566 50.5605
R2021 GND.n2249 GND.n2247 50.5605
R2022 GND.n2249 GND.n2248 50.5605
R2023 GND.n2243 GND.n2241 50.5605
R2024 GND.n2243 GND.n2242 50.5605
R2025 GND.n1224 GND.n1222 50.5605
R2026 GND.n1224 GND.n1223 50.5605
R2027 GND.n1218 GND.n1216 50.5605
R2028 GND.n1218 GND.n1217 50.5605
R2029 GND.n1676 GND.n1674 50.5605
R2030 GND.n1676 GND.n1675 50.5605
R2031 GND.n305 GND.n303 50.5605
R2032 GND.n305 GND.n304 50.5605
R2033 GND.n878 GND.n876 50.5605
R2034 GND.n878 GND.n877 50.5605
R2035 GND.n777 GND.n775 50.5605
R2036 GND.n777 GND.n776 50.5605
R2037 GND.n1979 GND.t517 50.1906
R2038 GND.t1469 GND.n5564 48.3834
R2039 GND GND.n5765 48.3834
R2040 GND.n6735 GND 47.7719
R2041 GND.n4426 GND 47.7719
R2042 GND.n3623 GND.t432 47.3332
R2043 GND.n3684 GND.n3683 47.2744
R2044 GND.n5176 GND 46.7305
R2045 GND.n7367 GND.n7358 46.2978
R2046 GND.n517 GND.n509 46.2978
R2047 GND.n212 GND.n204 46.2978
R2048 GND.n1511 GND.n1503 46.2978
R2049 GND.n1463 GND.n1455 46.2978
R2050 GND.n4220 GND.n4212 46.2978
R2051 GND.n3414 GND.n3406 46.2978
R2052 GND.n3257 GND.n3249 46.2978
R2053 GND.n2960 GND.n2952 46.2978
R2054 GND.n2635 GND.n2627 46.2978
R2055 GND.n2311 GND.n2303 46.2978
R2056 GND.n2149 GND.n2141 46.2978
R2057 GND.n1281 GND.n1273 46.2978
R2058 GND.n2019 GND.n2011 46.2978
R2059 GND.n364 GND.n356 46.2978
R2060 GND.n7412 GND.n7404 46.2978
R2061 GND.n1892 GND 46.1266
R2062 GND.n1849 GND 46.1266
R2063 GND GND.n7042 46.1266
R2064 GND.n2498 GND 46.1266
R2065 GND.n2823 GND 46.1266
R2066 GND.n3120 GND 46.1266
R2067 GND.n7220 GND 46.1266
R2068 GND.n4752 GND 46.1266
R2069 GND GND.n5434 46.1266
R2070 GND.t684 GND.n7355 43.8159
R2071 GND.t71 GND.n1551 43.4986
R2072 GND GND.n4913 43.3696
R2073 GND.n1996 GND.n1995 42.8187
R2074 GND.n7437 GND.n7436 42.8174
R2075 GND.n320 GND.n319 42.8174
R2076 GND.n473 GND.n472 42.8174
R2077 GND.n168 GND.n167 42.8174
R2078 GND.n1514 GND.n1513 42.8174
R2079 GND.n1466 GND.n1465 42.8174
R2080 GND.n4176 GND.n4175 42.8174
R2081 GND.n3370 GND.n3369 42.8174
R2082 GND.n3213 GND.n3212 42.8174
R2083 GND.n2916 GND.n2915 42.8174
R2084 GND.n2591 GND.n2590 42.8174
R2085 GND.n2267 GND.n2266 42.8174
R2086 GND.n2105 GND.n2104 42.8174
R2087 GND.n1237 GND.n1236 42.8174
R2088 GND.n7415 GND.n7414 42.8174
R2089 GND.n7045 GND.t697 42.5398
R2090 GND.n6089 GND 40.3307
R2091 GND.n6253 GND 40.3307
R2092 GND.n6562 GND 40.3307
R2093 GND.n702 GND 40.3307
R2094 GND.n7749 GND 40.3307
R2095 GND.n7584 GND 40.3307
R2096 GND.n4749 GND.t278 40.2035
R2097 GND.t422 GND.n3610 40.1687
R2098 GND.n4129 GND.t202 40.1687
R2099 GND.n7460 GND.n7441 39.6805
R2100 GND.n2047 GND.n2023 39.6805
R2101 GND.n540 GND.n521 39.6805
R2102 GND.n235 GND.n216 39.6805
R2103 GND.n1409 GND.n1390 39.6805
R2104 GND.n4243 GND.n4224 39.6805
R2105 GND.n3437 GND.n3418 39.6805
R2106 GND.n3280 GND.n3261 39.6805
R2107 GND.n2983 GND.n2964 39.6805
R2108 GND.n2658 GND.n2639 39.6805
R2109 GND.n2334 GND.n2315 39.6805
R2110 GND.n2172 GND.n2153 39.6805
R2111 GND.n1304 GND.n1285 39.6805
R2112 GND.n387 GND.n368 39.6805
R2113 GND.n812 GND.n793 39.6805
R2114 GND.n4961 GND.n4951 39.2858
R2115 GND.n6753 GND.n6752 39.2858
R2116 GND.n6790 GND.n6789 39.2858
R2117 GND.n5455 GND.n5445 39.2858
R2118 GND.n5459 GND.n5458 39.2858
R2119 GND.n5245 GND.n5244 39.2858
R2120 GND.n4392 GND.n4391 39.2858
R2121 GND.n4368 GND.n4367 39.2858
R2122 GND.n6860 GND.n6850 39.2858
R2123 GND.n6864 GND.n6863 39.2858
R2124 GND.n4337 GND.n4336 39.2858
R2125 GND.n6749 GND.n6736 38.7881
R2126 GND.n6786 GND.n6763 38.7881
R2127 GND.n5241 GND.n5222 38.7881
R2128 GND.n4388 GND.n4375 38.7881
R2129 GND.n4364 GND.n4341 38.7881
R2130 GND.n4333 GND.n4314 38.7881
R2131 GND.n6742 GND.t169 38.7697
R2132 GND.n6739 GND.t391 38.7697
R2133 GND.n6769 GND.t1277 38.7697
R2134 GND.n6766 GND.t739 38.7697
R2135 GND.n4381 GND.t118 38.7697
R2136 GND.n4378 GND.t1385 38.7697
R2137 GND.n4347 GND.t857 38.7697
R2138 GND.n4344 GND.t150 38.7697
R2139 GND.n5193 GND.n5191 38.7523
R2140 GND.n4290 GND.n4288 38.7523
R2141 GND.n4978 GND.t622 38.597
R2142 GND.n5471 GND.t737 38.5719
R2143 GND.n5471 GND.t105 38.5719
R2144 GND.n4402 GND.t1132 38.5719
R2145 GND.n4402 GND.t471 38.5719
R2146 GND.n6771 GND.t1529 38.5719
R2147 GND.n6771 GND.t1341 38.5719
R2148 GND.n5227 GND.t789 38.5719
R2149 GND.n5227 GND.t17 38.5719
R2150 GND.n5206 GND.t1134 38.5719
R2151 GND.n5206 GND.t1316 38.5719
R2152 GND.n5181 GND.t155 38.5719
R2153 GND.n5181 GND.t855 38.5719
R2154 GND.n5186 GND.t715 38.5719
R2155 GND.n5186 GND.t204 38.5719
R2156 GND.n4349 GND.t423 38.5719
R2157 GND.n4349 GND.t176 38.5719
R2158 GND.n4319 GND.t1569 38.5719
R2159 GND.n4319 GND.t1387 38.5719
R2160 GND.n4303 GND.t91 38.5719
R2161 GND.n4303 GND.t1343 38.5719
R2162 GND.n4278 GND.t827 38.5719
R2163 GND.n4278 GND.t141 38.5719
R2164 GND.n4283 GND.t601 38.5719
R2165 GND.n4283 GND.t1144 38.5719
R2166 GND.n7791 GND.n7790 37.1561
R2167 GND.n5565 GND.t1419 36.9992
R2168 GND.n4447 GND.t1103 36.8926
R2169 GND.n4542 GND.t1053 36.8926
R2170 GND.t51 GND.n3617 36.469
R2171 GND.t402 GND.t119 36.3723
R2172 GND.t1162 GND.t806 36.3723
R2173 GND.t830 GND.t419 36.3723
R2174 GND.t840 GND.t1187 36.3723
R2175 GND.t1166 GND.t186 36.3723
R2176 GND.t585 GND.t1227 36.3723
R2177 GND.t1257 GND.t1338 36.3723
R2178 GND.t158 GND.t1240 36.3723
R2179 GND.t400 GND.t590 36.3723
R2180 GND.t1159 GND.t602 36.3723
R2181 GND.t588 GND.t605 36.3723
R2182 GND.t598 GND.t661 36.3723
R2183 GND.t838 GND.t13 36.3723
R2184 GND.t1164 GND.t819 36.3723
R2185 GND.t685 GND.t1228 36.3723
R2186 GND.n350 GND.n321 35.6515
R2187 GND.n1449 GND.n1443 35.6515
R2188 GND.n3400 GND.n3371 35.6515
R2189 GND.n2946 GND.n2917 35.6515
R2190 GND.n2297 GND.n2268 35.6515
R2191 GND.n1267 GND.n1238 35.6515
R2192 GND.n1497 GND.n1489 35.6515
R2193 GND.n2005 GND.n2004 35.6515
R2194 GND.n7398 GND.n7397 35.6515
R2195 GND.n6725 GND.n6724 34.6358
R2196 GND.n5478 GND.n5477 34.6358
R2197 GND.n5481 GND.n5466 34.6358
R2198 GND.n5485 GND.n5466 34.6358
R2199 GND.n5486 GND.n5485 34.6358
R2200 GND.n4409 GND.n4408 34.6358
R2201 GND.n4412 GND.n4397 34.6358
R2202 GND.n4416 GND.n4397 34.6358
R2203 GND.n4417 GND.n4416 34.6358
R2204 GND.n5756 GND.n5755 34.6358
R2205 GND.n6745 GND.n6744 34.6358
R2206 GND.n6744 GND.n6737 34.6358
R2207 GND.n6752 GND.n6737 34.6358
R2208 GND.n6748 GND.n6747 34.6358
R2209 GND.n6749 GND.n6748 34.6358
R2210 GND.n6782 GND.n6781 34.6358
R2211 GND.n6781 GND.n6764 34.6358
R2212 GND.n6789 GND.n6764 34.6358
R2213 GND.n6785 GND.n6784 34.6358
R2214 GND.n6786 GND.n6785 34.6358
R2215 GND.n5455 GND.n5454 34.6358
R2216 GND.n5458 GND.n5446 34.6358
R2217 GND.n5244 GND.n5223 34.6358
R2218 GND.n5237 GND.n5236 34.6358
R2219 GND.n5200 GND.n5199 34.6358
R2220 GND.n6834 GND.n6833 34.6358
R2221 GND.n6828 GND.n6827 34.6358
R2222 GND.n6816 GND.n6815 34.6358
R2223 GND.n4384 GND.n4383 34.6358
R2224 GND.n4383 GND.n4376 34.6358
R2225 GND.n4391 GND.n4376 34.6358
R2226 GND.n4387 GND.n4386 34.6358
R2227 GND.n4388 GND.n4387 34.6358
R2228 GND.n4360 GND.n4359 34.6358
R2229 GND.n4359 GND.n4342 34.6358
R2230 GND.n4367 GND.n4342 34.6358
R2231 GND.n4363 GND.n4362 34.6358
R2232 GND.n4364 GND.n4363 34.6358
R2233 GND.n6860 GND.n6859 34.6358
R2234 GND.n6863 GND.n6851 34.6358
R2235 GND.n4336 GND.n4315 34.6358
R2236 GND.n4329 GND.n4328 34.6358
R2237 GND.n4297 GND.n4296 34.6358
R2238 GND.n7079 GND.n7078 34.6358
R2239 GND.n7073 GND.n7072 34.6358
R2240 GND.n7061 GND.n7060 34.6358
R2241 GND.n5167 GND.n5166 34.6358
R2242 GND.n5100 GND.t1556 34.4331
R2243 GND.t540 GND.n5766 34.1532
R2244 GND.n6822 GND.n6821 33.8829
R2245 GND.n7067 GND.n7066 33.8829
R2246 GND.n7359 GND.t1567 33.462
R2247 GND.n7359 GND.t658 33.462
R2248 GND.n7373 GND.t824 33.462
R2249 GND.n7373 GND.t113 33.462
R2250 GND.n1369 GND.t396 33.462
R2251 GND.n1369 GND.t362 33.462
R2252 GND.n2012 GND.t1185 33.462
R2253 GND.n2012 GND.t361 33.462
R2254 GND.n326 GND.t1272 33.462
R2255 GND.n326 GND.t849 33.462
R2256 GND.n479 GND.t620 33.462
R2257 GND.n479 GND.t1280 33.462
R2258 GND.n510 GND.t1261 33.462
R2259 GND.n510 GND.t798 33.462
R2260 GND.n174 GND.t760 33.462
R2261 GND.n174 GND.t1117 33.462
R2262 GND.n205 GND.t505 33.462
R2263 GND.n205 GND.t604 33.462
R2264 GND.n1483 GND.t76 33.462
R2265 GND.n1483 GND.t734 33.462
R2266 GND.n1504 GND.t675 33.462
R2267 GND.n1504 GND.t592 33.462
R2268 GND.n1382 GND.t1260 33.462
R2269 GND.n1382 GND.t691 33.462
R2270 GND.n1456 GND.t1254 33.462
R2271 GND.n1456 GND.t1241 33.462
R2272 GND.n4182 GND.t1365 33.462
R2273 GND.n4182 GND.t1173 33.462
R2274 GND.n4213 GND.t1381 33.462
R2275 GND.n4213 GND.t1339 33.462
R2276 GND.n3376 GND.t1340 33.462
R2277 GND.n3376 GND.t663 33.462
R2278 GND.n3407 GND.t348 33.462
R2279 GND.n3407 GND.t758 33.462
R2280 GND.n3219 GND.t1317 33.462
R2281 GND.n3219 GND.t1366 33.462
R2282 GND.n3250 GND.t367 33.462
R2283 GND.n3250 GND.t1279 33.462
R2284 GND.n2922 GND.t1194 33.462
R2285 GND.n2922 GND.t431 33.462
R2286 GND.n2953 GND.t720 33.462
R2287 GND.n2953 GND.t1186 33.462
R2288 GND.n2597 GND.t481 33.462
R2289 GND.n2597 GND.t433 33.462
R2290 GND.n2628 GND.t759 33.462
R2291 GND.n2628 GND.t421 33.462
R2292 GND.n2273 GND.t111 33.462
R2293 GND.n2273 GND.t1307 33.462
R2294 GND.n2304 GND.t514 33.462
R2295 GND.n2304 GND.t808 33.462
R2296 GND.n2111 GND.t1362 33.462
R2297 GND.n2111 GND.t693 33.462
R2298 GND.n2142 GND.t93 33.462
R2299 GND.n2142 GND.t121 33.462
R2300 GND.n1243 GND.t1231 33.462
R2301 GND.n1243 GND.t88 33.462
R2302 GND.n1274 GND.t717 33.462
R2303 GND.n1274 GND.t621 33.462
R2304 GND.n357 GND.t108 33.462
R2305 GND.n357 GND.t1312 33.462
R2306 GND.n7391 GND.t1319 33.462
R2307 GND.n7391 GND.t609 33.462
R2308 GND.n7405 GND.t1324 33.462
R2309 GND.n7405 GND.t820 33.462
R2310 GND.n6559 GND.t973 32.2518
R2311 GND.n6780 GND.n6779 32.1329
R2312 GND.n4358 GND.n4357 32.1329
R2313 GND.n1980 GND.n1979 31.7876
R2314 GND.n7568 GND.n7567 30.7897
R2315 GND.n7704 GND.n7703 30.7897
R2316 GND.n657 GND.n656 30.7897
R2317 GND.n6369 GND.n6368 30.7897
R2318 GND.n6205 GND.n6204 30.7897
R2319 GND.n6041 GND.n6040 30.7897
R2320 GND.n5858 GND.n5857 30.7897
R2321 GND.n5336 GND.n5335 30.7897
R2322 GND.n4895 GND.n4894 30.7897
R2323 GND.n7202 GND.n7201 30.7897
R2324 GND.n3102 GND.n3101 30.7897
R2325 GND.n2778 GND.n2777 30.7897
R2326 GND.n2453 GND.n2452 30.7897
R2327 GND.n6969 GND.n6968 30.7897
R2328 GND.n1804 GND.n1803 30.7897
R2329 GND.n1613 GND.n1612 30.7897
R2330 GND.n7660 GND.n7654 30.5561
R2331 GND.n4921 GND.t330 29.036
R2332 GND.n7044 GND.n7043 29.0202
R2333 GND.n7798 GND.n7793 28.9511
R2334 GND.n859 GND.n854 28.9511
R2335 GND.n752 GND.n747 28.9511
R2336 GND.n433 GND.n428 28.9511
R2337 GND.n1643 GND.n1638 28.9511
R2338 GND.n280 GND.n275 28.9511
R2339 GND.n128 GND.n123 28.9511
R2340 GND.n19 GND.n14 28.9511
R2341 GND.n7275 GND.n7270 28.9511
R2342 GND.n3485 GND.n3480 28.9511
R2343 GND.n3327 GND.n3322 28.9511
R2344 GND.n3170 GND.n3165 28.9511
R2345 GND.n2873 GND.n2868 28.9511
R2346 GND.n2548 GND.n2543 28.9511
R2347 GND.n2224 GND.n2219 28.9511
R2348 GND.n1199 GND.n1194 28.9511
R2349 GND.n7660 GND.n7659 28.8988
R2350 GND.n616 GND.n615 28.8988
R2351 GND.n6328 GND.n6327 28.8988
R2352 GND.n6164 GND.n6163 28.8988
R2353 GND.n5997 GND.n5996 28.8988
R2354 GND.n5814 GND.n5813 28.8988
R2355 GND.n5292 GND.n5291 28.8988
R2356 GND.n4851 GND.n4850 28.8988
R2357 GND.n7158 GND.n7157 28.8988
R2358 GND.n3058 GND.n3057 28.8988
R2359 GND.n2734 GND.n2733 28.8988
R2360 GND.n2409 GND.n2408 28.8988
R2361 GND.n6925 GND.n6924 28.8988
R2362 GND.n1760 GND.n1759 28.8988
R2363 GND.n1569 GND.n1568 28.8988
R2364 GND.n7557 GND.n7556 28.8193
R2365 GND.n7688 GND.n7687 28.8193
R2366 GND.n641 GND.n640 28.8193
R2367 GND.n6353 GND.n6352 28.8193
R2368 GND.n6189 GND.n6188 28.8193
R2369 GND.n6025 GND.n6024 28.8193
R2370 GND.n5842 GND.n5841 28.8193
R2371 GND.n5320 GND.n5319 28.8193
R2372 GND.n4879 GND.n4878 28.8193
R2373 GND.n7186 GND.n7185 28.8193
R2374 GND.n3086 GND.n3085 28.8193
R2375 GND.n2762 GND.n2761 28.8193
R2376 GND.n2437 GND.n2436 28.8193
R2377 GND.n6953 GND.n6952 28.8193
R2378 GND.n1788 GND.n1787 28.8193
R2379 GND.n1597 GND.n1596 28.8193
R2380 GND.n6615 GND.n6614 27.8593
R2381 GND.n6603 GND.n6602 27.8593
R2382 GND.n6513 GND.n6512 27.8593
R2383 GND.n6431 GND.n6430 27.8593
R2384 GND.n4660 GND.n4659 27.8593
R2385 GND.n4707 GND.n4706 27.8593
R2386 GND.n4947 GND.n4946 27.8593
R2387 GND.n5682 GND.n5681 27.8593
R2388 GND.n5502 GND.n5501 27.8593
R2389 GND.n5605 GND.n5604 27.8593
R2390 GND.n5523 GND.n5522 27.8593
R2391 GND.n5057 GND.n5056 27.8593
R2392 GND.n5045 GND.n5044 27.8593
R2393 GND.n4493 GND.n4492 27.8593
R2394 GND.n4481 GND.n4480 27.8593
R2395 GND.n5469 GND.t1199 27.5691
R2396 GND.n4400 GND.t773 27.5691
R2397 GND.n6772 GND.t1342 27.5691
R2398 GND.n5229 GND.t61 27.5691
R2399 GND.n5203 GND.t796 27.5691
R2400 GND.n5183 GND.t669 27.5691
R2401 GND.n5189 GND.t1245 27.5691
R2402 GND.n4350 GND.t1389 27.5691
R2403 GND.n4321 GND.t429 27.5691
R2404 GND.n4300 GND.t405 27.5691
R2405 GND.n4280 GND.t74 27.5691
R2406 GND.n4286 GND.t689 27.5691
R2407 GND.n4959 GND.n4950 27.1064
R2408 GND.n5919 GND 26.9763
R2409 GND.n4047 GND.t1130 26.8697
R2410 GND.n6717 GND.t1226 26.8576
R2411 GND.n5748 GND.t1369 26.8576
R2412 GND.n5159 GND.t1120 26.8576
R2413 GND.n4578 GND.t326 26.8025
R2414 GND.n1971 GND.n1970 26.7111
R2415 GND.n1733 GND.n1732 26.7111
R2416 GND.n1829 GND.n1828 26.7111
R2417 GND.n6994 GND.n6993 26.7111
R2418 GND.n2478 GND.n2477 26.7111
R2419 GND.n2803 GND.n2802 26.7111
R2420 GND.n7131 GND.n7130 26.7111
R2421 GND.n4824 GND.n4823 26.7111
R2422 GND.n5400 GND.n5399 26.7111
R2423 GND.n5361 GND.n5360 26.7111
R2424 GND.n5883 GND.n5882 26.7111
R2425 GND.n6069 GND.n6068 26.7111
R2426 GND.n6233 GND.n6232 26.7111
R2427 GND.n6397 GND.n6396 26.7111
R2428 GND.n682 GND.n681 26.7111
R2429 GND.n7729 GND.n7728 26.7111
R2430 GND.t410 GND.n4977 26.1036
R2431 GND.n5487 GND.t1383 25.9346
R2432 GND.n4418 GND.t377 25.9346
R2433 GND.t1284 GND.t1286 25.66
R2434 GND.t1286 GND.t1288 25.66
R2435 GND.t1288 GND.t1291 25.66
R2436 GND.t42 GND.t44 25.66
R2437 GND.t44 GND.t47 25.66
R2438 GND.t47 GND.t49 25.66
R2439 GND.t568 GND.t566 25.66
R2440 GND.t571 GND.t568 25.66
R2441 GND.t573 GND.t571 25.66
R2442 GND.t493 GND.t495 25.66
R2443 GND.t495 GND.t489 25.66
R2444 GND.t489 GND.t491 25.66
R2445 GND.t1376 GND.t1378 25.66
R2446 GND.t1378 GND.t1372 25.66
R2447 GND.t1372 GND.t1374 25.66
R2448 GND.t7 GND.t9 25.66
R2449 GND.t9 GND.t11 25.66
R2450 GND.t11 GND.t4 25.66
R2451 GND.t1269 GND.t1262 25.66
R2452 GND.t1262 GND.t1265 25.66
R2453 GND.t1265 GND.t1267 25.66
R2454 GND.t753 GND.t755 25.66
R2455 GND.t755 GND.t749 25.66
R2456 GND.t749 GND.t751 25.66
R2457 GND.t1393 GND.t1391 25.66
R2458 GND.t1396 GND.t1393 25.66
R2459 GND.t1398 GND.t1396 25.66
R2460 GND.n3623 GND.t52 25.4873
R2461 GND.n7818 GND.n7808 25.0358
R2462 GND.n890 GND.n871 25.0358
R2463 GND.n783 GND.n764 25.0358
R2464 GND.n464 GND.n445 25.0358
R2465 GND.n1682 GND.n1655 25.0358
R2466 GND.n311 GND.n292 25.0358
R2467 GND.n159 GND.n140 25.0358
R2468 GND.n50 GND.n31 25.0358
R2469 GND.n7306 GND.n7287 25.0358
R2470 GND.n3516 GND.n3497 25.0358
R2471 GND.n3358 GND.n3339 25.0358
R2472 GND.n3201 GND.n3182 25.0358
R2473 GND.n2904 GND.n2885 25.0358
R2474 GND.n2579 GND.n2560 25.0358
R2475 GND.n2255 GND.n2236 25.0358
R2476 GND.n1230 GND.n1211 25.0358
R2477 GND.n6704 GND.t1353 24.9236
R2478 GND.n6704 GND.t1355 24.9236
R2479 GND.n5491 GND.t465 24.9236
R2480 GND.n5491 GND.t445 24.9236
R2481 GND.n6664 GND.t453 24.9236
R2482 GND.n6664 GND.t463 24.9236
R2483 GND.n6670 GND.t459 24.9236
R2484 GND.n6670 GND.t467 24.9236
R2485 GND.n6674 GND.t447 24.9236
R2486 GND.n6674 GND.t461 24.9236
R2487 GND.n6680 GND.t469 24.9236
R2488 GND.n6680 GND.t449 24.9236
R2489 GND.n6686 GND.t455 24.9236
R2490 GND.n6686 GND.t439 24.9236
R2491 GND.n6692 GND.t443 24.9236
R2492 GND.n6692 GND.t457 24.9236
R2493 GND.n6607 GND.t968 24.9236
R2494 GND.n6607 GND.t866 24.9236
R2495 GND.n6651 GND.t946 24.9236
R2496 GND.n6651 GND.t972 24.9236
R2497 GND.n6644 GND.t904 24.9236
R2498 GND.n6644 GND.t926 24.9236
R2499 GND.n6640 GND.t960 24.9236
R2500 GND.n6640 GND.t894 24.9236
R2501 GND.n6634 GND.t930 24.9236
R2502 GND.n6634 GND.t872 24.9236
R2503 GND.n6628 GND.t954 24.9236
R2504 GND.n6628 GND.t982 24.9236
R2505 GND.n6622 GND.t914 24.9236
R2506 GND.n6622 GND.t938 24.9236
R2507 GND.n6517 GND.t922 24.9236
R2508 GND.n6517 GND.t952 24.9236
R2509 GND.n6524 GND.t888 24.9236
R2510 GND.n6524 GND.t974 24.9236
R2511 GND.n6550 GND.t884 24.9236
R2512 GND.n6550 GND.t948 24.9236
R2513 GND.n6546 GND.t976 24.9236
R2514 GND.n6546 GND.t906 24.9236
R2515 GND.n6540 GND.t932 24.9236
R2516 GND.n6540 GND.t964 24.9236
R2517 GND.n6534 GND.t908 24.9236
R2518 GND.n6534 GND.t934 24.9236
R2519 GND.n6528 GND.t880 24.9236
R2520 GND.n6528 GND.t902 24.9236
R2521 GND.n6433 GND.t944 24.9236
R2522 GND.n6433 GND.t970 24.9236
R2523 GND.n6476 GND.t868 24.9236
R2524 GND.n6476 GND.t924 24.9236
R2525 GND.n6483 GND.t958 24.9236
R2526 GND.n6483 GND.t890 24.9236
R2527 GND.n6487 GND.t928 24.9236
R2528 GND.n6487 GND.t962 24.9236
R2529 GND.n6493 GND.t898 24.9236
R2530 GND.n6493 GND.t978 24.9236
R2531 GND.n6499 GND.t910 24.9236
R2532 GND.n6499 GND.t936 24.9236
R2533 GND.n6505 GND.t984 24.9236
R2534 GND.n6505 GND.t916 24.9236
R2535 GND.n6419 GND.t900 24.9236
R2536 GND.n6419 GND.t986 24.9236
R2537 GND.n6424 GND.t878 24.9236
R2538 GND.n6424 GND.t870 24.9236
R2539 GND.n6466 GND.t892 24.9236
R2540 GND.n6466 GND.t918 24.9236
R2541 GND.n6461 GND.t860 24.9236
R2542 GND.n6461 GND.t896 24.9236
R2543 GND.n6455 GND.t966 24.9236
R2544 GND.n6455 GND.t862 24.9236
R2545 GND.n6449 GND.t886 24.9236
R2546 GND.n6449 GND.t950 24.9236
R2547 GND.n6443 GND.t980 24.9236
R2548 GND.n6443 GND.t912 24.9236
R2549 GND.n1937 GND.t55 24.9236
R2550 GND.n1937 GND.t57 24.9236
R2551 GND.n1904 GND.t1287 24.9236
R2552 GND.n1904 GND.t1289 24.9236
R2553 GND.n1704 GND.t373 24.9236
R2554 GND.n1704 GND.t370 24.9236
R2555 GND.n1861 GND.t45 24.9236
R2556 GND.n1861 GND.t48 24.9236
R2557 GND.n6912 GND.t484 24.9236
R2558 GND.n6912 GND.t485 24.9236
R2559 GND.n6882 GND.t569 24.9236
R2560 GND.n6882 GND.t572 24.9236
R2561 GND.n2380 GND.t139 24.9236
R2562 GND.n2380 GND.t135 24.9236
R2563 GND.n2510 GND.t496 24.9236
R2564 GND.n2510 GND.t490 24.9236
R2565 GND.n2705 GND.t28 24.9236
R2566 GND.n2705 GND.t29 24.9236
R2567 GND.n2835 GND.t1379 24.9236
R2568 GND.n2835 GND.t1373 24.9236
R2569 GND.n3029 GND.t614 24.9236
R2570 GND.n3029 GND.t615 24.9236
R2571 GND.n3132 GND.t10 24.9236
R2572 GND.n3132 GND.t12 24.9236
R2573 GND.n7102 GND.t582 24.9236
R2574 GND.n7102 GND.t578 24.9236
R2575 GND.n7232 GND.t1263 24.9236
R2576 GND.n7232 GND.t1266 24.9236
R2577 GND.n4797 GND.t181 24.9236
R2578 GND.n4797 GND.t182 24.9236
R2579 GND.n4764 GND.t756 24.9236
R2580 GND.n4764 GND.t750 24.9236
R2581 GND.n5279 GND.t810 24.9236
R2582 GND.n5279 GND.t811 24.9236
R2583 GND.n5249 GND.t1394 24.9236
R2584 GND.n5249 GND.t1397 24.9236
R2585 GND.n5801 GND.t1193 24.9236
R2586 GND.n5801 GND.t1189 24.9236
R2587 GND.n5932 GND.t1328 24.9236
R2588 GND.n5932 GND.t1331 24.9236
R2589 GND.n5968 GND.t844 24.9236
R2590 GND.n5968 GND.t845 24.9236
R2591 GND.n6101 GND.t98 24.9236
R2592 GND.n6101 GND.t101 24.9236
R2593 GND.n6135 GND.t508 24.9236
R2594 GND.n6135 GND.t509 24.9236
R2595 GND.n6265 GND.t764 24.9236
R2596 GND.n6265 GND.t767 24.9236
R2597 GND.n6299 GND.t381 24.9236
R2598 GND.n6299 GND.t382 24.9236
R2599 GND.n6574 GND.t1207 24.9236
R2600 GND.n6574 GND.t1201 24.9236
R2601 GND.n587 GND.t131 24.9236
R2602 GND.n587 GND.t132 24.9236
R2603 GND.n714 GND.t196 24.9236
R2604 GND.n714 GND.t199 24.9236
R2605 GND.n7630 GND.t358 24.9236
R2606 GND.n7630 GND.t354 24.9236
R2607 GND.n7761 GND.t1216 24.9236
R2608 GND.n7761 GND.t1219 24.9236
R2609 GND.n7510 GND.t501 24.9236
R2610 GND.n7510 GND.t502 24.9236
R2611 GND.n7596 GND.t213 24.9236
R2612 GND.n7596 GND.t207 24.9236
R2613 GND.n4965 GND.t416 24.9236
R2614 GND.n4965 GND.t418 24.9236
R2615 GND.n4652 GND.t273 24.9236
R2616 GND.n4652 GND.t307 24.9236
R2617 GND.n4646 GND.t259 24.9236
R2618 GND.n4646 GND.t221 24.9236
R2619 GND.n4640 GND.t245 24.9236
R2620 GND.n4640 GND.t301 24.9236
R2621 GND.n4636 GND.t333 24.9236
R2622 GND.n4636 GND.t233 24.9236
R2623 GND.n4609 GND.t285 24.9236
R2624 GND.n4609 GND.t337 24.9236
R2625 GND.n4671 GND.t263 24.9236
R2626 GND.n4671 GND.t289 24.9236
R2627 GND.n4677 GND.t321 24.9236
R2628 GND.n4677 GND.t257 24.9236
R2629 GND.n4689 GND.t325 24.9236
R2630 GND.n4689 GND.t239 24.9236
R2631 GND.n4695 GND.t297 24.9236
R2632 GND.n4695 GND.t329 24.9236
R2633 GND.n4702 GND.t229 24.9236
R2634 GND.n4702 GND.t279 24.9236
R2635 GND.n4743 GND.t315 24.9236
R2636 GND.n4743 GND.t251 24.9236
R2637 GND.n4736 GND.t283 24.9236
R2638 GND.n4736 GND.t249 24.9236
R2639 GND.n4730 GND.t309 24.9236
R2640 GND.n4730 GND.t341 24.9236
R2641 GND.n4724 GND.t267 24.9236
R2642 GND.n4724 GND.t293 24.9236
R2643 GND.n4714 GND.t323 24.9236
R2644 GND.n4714 GND.t225 24.9236
R2645 GND.n4708 GND.t275 24.9236
R2646 GND.n4708 GND.t243 24.9236
R2647 GND.n4924 GND.t299 24.9236
R2648 GND.n4924 GND.t331 24.9236
R2649 GND.n4929 GND.t247 24.9236
R2650 GND.n4929 GND.t303 24.9236
R2651 GND.n4936 GND.t335 24.9236
R2652 GND.n4936 GND.t261 24.9236
R2653 GND.n4942 GND.t287 24.9236
R2654 GND.n4942 GND.t319 24.9236
R2655 GND.n5032 GND.t265 24.9236
R2656 GND.n5032 GND.t291 24.9236
R2657 GND.n5021 GND.t631 24.9236
R2658 GND.n5021 GND.t641 24.9236
R2659 GND.n5011 GND.t651 24.9236
R2660 GND.n5011 GND.t629 24.9236
R2661 GND.n5004 GND.t643 24.9236
R2662 GND.n5004 GND.t653 24.9236
R2663 GND.n5000 GND.t633 24.9236
R2664 GND.n5000 GND.t639 24.9236
R2665 GND.n4994 GND.t649 24.9236
R2666 GND.n4994 GND.t645 24.9236
R2667 GND.n4988 GND.t627 24.9236
R2668 GND.n4988 GND.t637 24.9236
R2669 GND.n4981 GND.t647 24.9236
R2670 GND.n4981 GND.t623 24.9236
R2671 GND.n4582 GND.t255 24.9236
R2672 GND.n4582 GND.t327 24.9236
R2673 GND.n4590 GND.t227 24.9236
R2674 GND.n4590 GND.t277 24.9236
R2675 GND.n4596 GND.t313 24.9236
R2676 GND.n4596 GND.t231 24.9236
R2677 GND.n4600 GND.t281 24.9236
R2678 GND.n4600 GND.t317 24.9236
R2679 GND.n4613 GND.t305 24.9236
R2680 GND.n4613 GND.t339 24.9236
R2681 GND.n4619 GND.t235 24.9236
R2682 GND.n4619 GND.t311 24.9236
R2683 GND.n4625 GND.t343 24.9236
R2684 GND.n4625 GND.t269 24.9236
R2685 GND.n5735 GND.t1157 24.9236
R2686 GND.n5735 GND.t1151 24.9236
R2687 GND.n5687 GND.t561 24.9236
R2688 GND.n5687 GND.t541 24.9236
R2689 GND.n5695 GND.t549 24.9236
R2690 GND.n5695 GND.t559 24.9236
R2691 GND.n5701 GND.t555 24.9236
R2692 GND.n5701 GND.t563 24.9236
R2693 GND.n5705 GND.t543 24.9236
R2694 GND.n5705 GND.t557 24.9236
R2695 GND.n5711 GND.t565 24.9236
R2696 GND.n5711 GND.t545 24.9236
R2697 GND.n5717 GND.t551 24.9236
R2698 GND.n5717 GND.t535 24.9236
R2699 GND.n5723 GND.t539 24.9236
R2700 GND.n5723 GND.t553 24.9236
R2701 GND.n5773 GND.t1520 24.9236
R2702 GND.n5773 GND.t1418 24.9236
R2703 GND.n5503 GND.t1498 24.9236
R2704 GND.n5503 GND.t1524 24.9236
R2705 GND.n5652 GND.t1456 24.9236
R2706 GND.n5652 GND.t1478 24.9236
R2707 GND.n5656 GND.t1512 24.9236
R2708 GND.n5656 GND.t1446 24.9236
R2709 GND.n5662 GND.t1482 24.9236
R2710 GND.n5662 GND.t1424 24.9236
R2711 GND.n5668 GND.t1506 24.9236
R2712 GND.n5668 GND.t1406 24.9236
R2713 GND.n5674 GND.t1466 24.9236
R2714 GND.n5674 GND.t1490 24.9236
R2715 GND.n5609 GND.t1474 24.9236
R2716 GND.n5609 GND.t1504 24.9236
R2717 GND.n5616 GND.t1440 24.9236
R2718 GND.n5616 GND.t1526 24.9236
R2719 GND.n5638 GND.t1436 24.9236
R2720 GND.n5638 GND.t1500 24.9236
R2721 GND.n5634 GND.t1528 24.9236
R2722 GND.n5634 GND.t1458 24.9236
R2723 GND.n5628 GND.t1484 24.9236
R2724 GND.n5628 GND.t1516 24.9236
R2725 GND.n5622 GND.t1460 24.9236
R2726 GND.n5622 GND.t1486 24.9236
R2727 GND.n5497 GND.t1432 24.9236
R2728 GND.n5497 GND.t1454 24.9236
R2729 GND.n5525 GND.t1496 24.9236
R2730 GND.n5525 GND.t1522 24.9236
R2731 GND.n5568 GND.t1420 24.9236
R2732 GND.n5568 GND.t1476 24.9236
R2733 GND.n5575 GND.t1510 24.9236
R2734 GND.n5575 GND.t1442 24.9236
R2735 GND.n5579 GND.t1480 24.9236
R2736 GND.n5579 GND.t1514 24.9236
R2737 GND.n5585 GND.t1450 24.9236
R2738 GND.n5585 GND.t1402 24.9236
R2739 GND.n5591 GND.t1462 24.9236
R2740 GND.n5591 GND.t1488 24.9236
R2741 GND.n5597 GND.t1408 24.9236
R2742 GND.n5597 GND.t1468 24.9236
R2743 GND.n5510 GND.t1452 24.9236
R2744 GND.n5510 GND.t1410 24.9236
R2745 GND.n5515 GND.t1430 24.9236
R2746 GND.n5515 GND.t1422 24.9236
R2747 GND.n5558 GND.t1444 24.9236
R2748 GND.n5558 GND.t1470 24.9236
R2749 GND.n5553 GND.t1412 24.9236
R2750 GND.n5553 GND.t1448 24.9236
R2751 GND.n5547 GND.t1518 24.9236
R2752 GND.n5547 GND.t1414 24.9236
R2753 GND.n5541 GND.t1438 24.9236
R2754 GND.n5541 GND.t1502 24.9236
R2755 GND.n5535 GND.t1404 24.9236
R2756 GND.n5535 GND.t1464 24.9236
R2757 GND.n5146 GND.t86 24.9236
R2758 GND.n5146 GND.t80 24.9236
R2759 GND.n4427 GND.t1545 24.9236
R2760 GND.n4427 GND.t1557 24.9236
R2761 GND.n5106 GND.t1565 24.9236
R2762 GND.n5106 GND.t1543 24.9236
R2763 GND.n5112 GND.t1539 24.9236
R2764 GND.n5112 GND.t1547 24.9236
R2765 GND.n5116 GND.t1559 24.9236
R2766 GND.n5116 GND.t1541 24.9236
R2767 GND.n5122 GND.t1549 24.9236
R2768 GND.n5122 GND.t1561 24.9236
R2769 GND.n5128 GND.t1535 24.9236
R2770 GND.n5128 GND.t1551 24.9236
R2771 GND.n5134 GND.t1555 24.9236
R2772 GND.n5134 GND.t1537 24.9236
R2773 GND.n5049 GND.t1026 24.9236
R2774 GND.n5049 GND.t1052 24.9236
R2775 GND.n5093 GND.t1004 24.9236
R2776 GND.n5093 GND.t1030 24.9236
R2777 GND.n5086 GND.t1090 24.9236
R2778 GND.n5086 GND.t1112 24.9236
R2779 GND.n5082 GND.t1018 24.9236
R2780 GND.n5082 GND.t1080 24.9236
R2781 GND.n5076 GND.t988 24.9236
R2782 GND.n5076 GND.t1058 24.9236
R2783 GND.n5070 GND.t1012 24.9236
R2784 GND.n5070 GND.t1040 24.9236
R2785 GND.n5064 GND.t1100 24.9236
R2786 GND.n5064 GND.t996 24.9236
R2787 GND.n4497 GND.t1108 24.9236
R2788 GND.n4497 GND.t1010 24.9236
R2789 GND.n4431 GND.t1074 24.9236
R2790 GND.n4431 GND.t1032 24.9236
R2791 GND.n4549 GND.t1070 24.9236
R2792 GND.n4549 GND.t1006 24.9236
R2793 GND.n4553 GND.t1034 24.9236
R2794 GND.n4553 GND.t1092 24.9236
R2795 GND.n4559 GND.t990 24.9236
R2796 GND.n4559 GND.t1022 24.9236
R2797 GND.n4565 GND.t1094 24.9236
R2798 GND.n4565 GND.t992 24.9236
R2799 GND.n4571 GND.t1066 24.9236
R2800 GND.n4571 GND.t1088 24.9236
R2801 GND.n4485 GND.t1002 24.9236
R2802 GND.n4485 GND.t1028 24.9236
R2803 GND.n4536 GND.t1054 24.9236
R2804 GND.n4536 GND.t1110 24.9236
R2805 GND.n4529 GND.t1016 24.9236
R2806 GND.n4529 GND.t1076 24.9236
R2807 GND.n4525 GND.t1114 24.9236
R2808 GND.n4525 GND.t1020 24.9236
R2809 GND.n4519 GND.t1084 24.9236
R2810 GND.n4519 GND.t1036 24.9236
R2811 GND.n4513 GND.t1096 24.9236
R2812 GND.n4513 GND.t994 24.9236
R2813 GND.n4507 GND.t1042 24.9236
R2814 GND.n4507 GND.t1102 24.9236
R2815 GND.n4435 GND.t1086 24.9236
R2816 GND.n4435 GND.t1044 24.9236
R2817 GND.n4440 GND.t1064 24.9236
R2818 GND.n4440 GND.t1056 24.9236
R2819 GND.n4450 GND.t1078 24.9236
R2820 GND.n4450 GND.t1104 24.9236
R2821 GND.n4455 GND.t1046 24.9236
R2822 GND.n4455 GND.t1082 24.9236
R2823 GND.n4461 GND.t1024 24.9236
R2824 GND.n4461 GND.t1048 24.9236
R2825 GND.n4467 GND.t1072 24.9236
R2826 GND.n4467 GND.t1008 24.9236
R2827 GND.n4473 GND.t1038 24.9236
R2828 GND.n4473 GND.t1098 24.9236
R2829 GND.n6700 GND.n6699 24.4711
R2830 GND.n5477 GND.n5468 24.4711
R2831 GND.n4408 GND.n4399 24.4711
R2832 GND.n4949 GND.n4948 24.4711
R2833 GND.n5731 GND.n5730 24.4711
R2834 GND.n5237 GND.n5233 24.4711
R2835 GND.n5194 GND.n5193 24.4711
R2836 GND.n4329 GND.n4325 24.4711
R2837 GND.n4291 GND.n4290 24.4711
R2838 GND.n5142 GND.n5141 24.4711
R2839 GND.t596 GND.n2006 23.9028
R2840 GND.t597 GND.n1268 23.9028
R2841 GND.t587 GND.n2298 23.9028
R2842 GND.t594 GND.n2947 23.9028
R2843 GND.t1161 GND.n3401 23.9028
R2844 GND.t732 GND.n1450 23.9028
R2845 GND.t399 GND.n1498 23.9028
R2846 GND.t160 GND.n351 23.9028
R2847 GND.t593 GND.n7399 23.9028
R2848 GND.n5200 GND.n5184 23.7181
R2849 GND.n4297 GND.n4281 23.7181
R2850 GND.n7460 GND.n7459 23.4245
R2851 GND.n2047 GND.n2046 23.4245
R2852 GND.n540 GND.n539 23.4245
R2853 GND.n235 GND.n234 23.4245
R2854 GND.n68 GND.n67 23.4245
R2855 GND.n1409 GND.n1408 23.4245
R2856 GND.n4243 GND.n4242 23.4245
R2857 GND.n3437 GND.n3436 23.4245
R2858 GND.n3280 GND.n3279 23.4245
R2859 GND.n2983 GND.n2982 23.4245
R2860 GND.n2658 GND.n2657 23.4245
R2861 GND.n2334 GND.n2333 23.4245
R2862 GND.n2172 GND.n2171 23.4245
R2863 GND.n1304 GND.n1303 23.4245
R2864 GND.n387 GND.n386 23.4245
R2865 GND.n812 GND.n811 23.4245
R2866 GND.n5473 GND.n5472 22.9652
R2867 GND.n4404 GND.n4403 22.9652
R2868 GND.n6775 GND.n6774 22.9652
R2869 GND.n5232 GND.n5228 22.9652
R2870 GND.n5207 GND.n5205 22.9652
R2871 GND.n5212 GND.n5211 22.9652
R2872 GND.n4353 GND.n4352 22.9652
R2873 GND.n4324 GND.n4320 22.9652
R2874 GND.n4304 GND.n4302 22.9652
R2875 GND.n4309 GND.n4308 22.9652
R2876 GND.n7569 GND.n7568 22.9087
R2877 GND.n7705 GND.n7704 22.9087
R2878 GND.n658 GND.n657 22.9087
R2879 GND.n6370 GND.n6369 22.9087
R2880 GND.n6206 GND.n6205 22.9087
R2881 GND.n6042 GND.n6041 22.9087
R2882 GND.n5859 GND.n5858 22.9087
R2883 GND.n5337 GND.n5336 22.9087
R2884 GND.n4896 GND.n4895 22.9087
R2885 GND.n7203 GND.n7202 22.9087
R2886 GND.n3103 GND.n3102 22.9087
R2887 GND.n2779 GND.n2778 22.9087
R2888 GND.n2454 GND.n2453 22.9087
R2889 GND.n6970 GND.n6969 22.9087
R2890 GND.n1805 GND.n1804 22.9087
R2891 GND.n1614 GND.n1613 22.9087
R2892 GND.t733 GND.n2136 22.765
R2893 GND.t595 GND.n2622 22.765
R2894 GND.t1158 GND.n3244 22.765
R2895 GND.t837 GND.n4207 22.765
R2896 GND.t435 GND.n199 22.765
R2897 GND.t161 GND.n504 22.765
R2898 GND.n6049 GND.n6048 22.5323
R2899 GND.n6213 GND.n6212 22.5323
R2900 GND.n6377 GND.n6376 22.5323
R2901 GND.t1325 GND.t1327 22.4359
R2902 GND.t1327 GND.t1330 22.4359
R2903 GND.t1330 GND.t1332 22.4359
R2904 GND.t95 GND.t97 22.4359
R2905 GND.t97 GND.t100 22.4359
R2906 GND.t100 GND.t102 22.4359
R2907 GND.t761 GND.t763 22.4359
R2908 GND.t763 GND.t766 22.4359
R2909 GND.t766 GND.t768 22.4359
R2910 GND.t1204 GND.t1206 22.4359
R2911 GND.t1206 GND.t1200 22.4359
R2912 GND.t1200 GND.t1202 22.4359
R2913 GND.t193 GND.t195 22.4359
R2914 GND.t195 GND.t198 22.4359
R2915 GND.t198 GND.t191 22.4359
R2916 GND.t1213 GND.t1215 22.4359
R2917 GND.t1215 GND.t1218 22.4359
R2918 GND.t1218 GND.t1220 22.4359
R2919 GND.t210 GND.t212 22.4359
R2920 GND.t212 GND.t206 22.4359
R2921 GND.t206 GND.t208 22.4359
R2922 GND.n1579 GND.n1578 22.4086
R2923 GND.n1770 GND.n1769 22.4086
R2924 GND.n6935 GND.n6934 22.4086
R2925 GND.n2419 GND.n2418 22.4086
R2926 GND.n2744 GND.n2743 22.4086
R2927 GND.n3068 GND.n3067 22.4086
R2928 GND.n7168 GND.n7167 22.4086
R2929 GND.n4861 GND.n4860 22.4086
R2930 GND.n5302 GND.n5301 22.4086
R2931 GND.n5824 GND.n5823 22.4086
R2932 GND.n6007 GND.n6006 22.4086
R2933 GND.n7670 GND.n7669 22.4086
R2934 GND.n7539 GND.n7538 22.4086
R2935 GND.n5479 GND.t173 22.3257
R2936 GND.n4410 GND.t65 22.3257
R2937 GND.n5448 GND.t398 22.3257
R2938 GND.n5450 GND.t1306 22.3257
R2939 GND.n5234 GND.t1337 22.3257
R2940 GND.n5225 GND.t1323 22.3257
R2941 GND.n5190 GND.t657 22.3257
R2942 GND.n6853 GND.t350 22.3257
R2943 GND.n6855 GND.t352 22.3257
R2944 GND.n4326 GND.t69 22.3257
R2945 GND.n4317 GND.t1222 22.3257
R2946 GND.n4287 GND.t35 22.3257
R2947 GND.t172 GND 22.2656
R2948 GND.n5199 GND.n5187 22.2123
R2949 GND.n5195 GND.n5187 22.2123
R2950 GND.n4296 GND.n4284 22.2123
R2951 GND.n4292 GND.n4284 22.2123
R2952 GND.n1974 GND.n1973 22.0429
R2953 GND.n1736 GND.n1735 22.0429
R2954 GND.n1832 GND.n1831 22.0429
R2955 GND.n6997 GND.n6996 22.0429
R2956 GND.n2481 GND.n2480 22.0429
R2957 GND.n2806 GND.n2805 22.0429
R2958 GND.n7134 GND.n7133 22.0429
R2959 GND.n4827 GND.n4826 22.0429
R2960 GND.n5403 GND.n5402 22.0429
R2961 GND.n5364 GND.n5363 22.0429
R2962 GND.n5886 GND.n5885 22.0429
R2963 GND.n6072 GND.n6071 22.0429
R2964 GND.n6236 GND.n6235 22.0429
R2965 GND.n6400 GND.n6399 22.0429
R2966 GND.n685 GND.n684 22.0429
R2967 GND.n7732 GND.n7731 22.0429
R2968 GND.n1930 GND.n1929 21.8358
R2969 GND.n1697 GND.n1696 21.8358
R2970 GND.n6905 GND.n6904 21.8358
R2971 GND.n2373 GND.n2372 21.8358
R2972 GND.n2698 GND.n2697 21.8358
R2973 GND.n3022 GND.n3021 21.8358
R2974 GND.n7095 GND.n7094 21.8358
R2975 GND.n4790 GND.n4789 21.8358
R2976 GND.n5272 GND.n5271 21.8358
R2977 GND.n5794 GND.n5793 21.8358
R2978 GND.n5961 GND.n5960 21.8358
R2979 GND.n6128 GND.n6127 21.8358
R2980 GND.n6292 GND.n6291 21.8358
R2981 GND.n580 GND.n579 21.8358
R2982 GND.n7623 GND.n7622 21.8358
R2983 GND.n7503 GND.n7502 21.8358
R2984 GND.n5488 GND.n5486 21.4593
R2985 GND.n4419 GND.n4417 21.4593
R2986 GND.n6745 GND.n6743 21.4593
R2987 GND.n6747 GND.n6740 21.4593
R2988 GND.n6782 GND.n6780 21.4593
R2989 GND.n6784 GND.n6767 21.4593
R2990 GND.n5208 GND.n5207 21.4593
R2991 GND.n5211 GND.n5210 21.4593
R2992 GND.n4384 GND.n4382 21.4593
R2993 GND.n4386 GND.n4379 21.4593
R2994 GND.n4360 GND.n4358 21.4593
R2995 GND.n4362 GND.n4345 21.4593
R2996 GND.n4305 GND.n4304 21.4593
R2997 GND.n4308 GND.n4307 21.4593
R2998 GND.n6755 GND.n6735 21.3675
R2999 GND.n408 GND.n407 20.6255
R3000 GND.n1433 GND.n1428 20.6255
R3001 GND.n3457 GND.n3452 20.6255
R3002 GND.n3003 GND.n2998 20.6255
R3003 GND.n2354 GND.n2349 20.6255
R3004 GND.n1317 GND.n1316 20.6255
R3005 GND.n2196 GND.n2191 20.6255
R3006 GND.n2679 GND.n2674 20.6255
R3007 GND.n3299 GND.n3294 20.6255
R3008 GND.n4260 GND.n4255 20.6255
R3009 GND.n252 GND.n247 20.6255
R3010 GND.n2076 GND.n2075 20.6255
R3011 GND.n834 GND.n833 20.6255
R3012 GND.n561 GND.n556 20.6255
R3013 GND.n7484 GND.n7475 20.6255
R3014 GND.n1350 GND.n1329 20.0775
R3015 GND.n5473 GND.n5468 19.9534
R3016 GND.n4404 GND.n4399 19.9534
R3017 GND.n6776 GND.n6775 19.9534
R3018 GND.n5233 GND.n5232 19.9534
R3019 GND.n5205 GND.n5180 19.9534
R3020 GND.n5213 GND.n5212 19.9534
R3021 GND.n4354 GND.n4353 19.9534
R3022 GND.n4325 GND.n4324 19.9534
R3023 GND.n4302 GND.n4277 19.9534
R3024 GND.n4310 GND.n4309 19.9534
R3025 GND.n7803 GND.n7802 19.5561
R3026 GND.t346 GND.t14 19.2425
R3027 GND.t703 GND.t175 19.2425
R3028 GND.n1995 GND.n1994 19.2005
R3029 GND.n1943 GND.t518 17.475
R3030 GND.n1712 GND.t1345 17.475
R3031 GND.n7024 GND.t775 17.475
R3032 GND.n2388 GND.t805 17.475
R3033 GND.n2713 GND.t816 17.475
R3034 GND.n3037 GND.t143 17.475
R3035 GND.n7110 GND.t829 17.475
R3036 GND.n4803 GND.t522 17.475
R3037 GND.n5419 GND.t1310 17.475
R3038 GND.n5914 GND.t479 17.475
R3039 GND.n5976 GND.t745 17.475
R3040 GND.n6143 GND.t19 17.475
R3041 GND.n6307 GND.t1116 17.475
R3042 GND.n595 GND.t1184 17.475
R3043 GND.n7638 GND.t1233 17.475
R3044 GND.n7518 GND.t1142 17.475
R3045 GND.n7782 GND.t1256 17.4601
R3046 GND.n841 GND.t686 17.4601
R3047 GND.n734 GND.t1165 17.4601
R3048 GND.n415 GND.t839 17.4601
R3049 GND.n1625 GND.t599 17.4601
R3050 GND.n262 GND.t589 17.4601
R3051 GND.n110 GND.t1160 17.4601
R3052 GND.n1 GND.t401 17.4601
R3053 GND.n7257 GND.t159 17.4601
R3054 GND.n3467 GND.t1258 17.4601
R3055 GND.n3309 GND.t586 17.4601
R3056 GND.n3152 GND.t1167 17.4601
R3057 GND.n2855 GND.t841 17.4601
R3058 GND.n2530 GND.t831 17.4601
R3059 GND.n2206 GND.t1163 17.4601
R3060 GND.n1181 GND.t403 17.4601
R3061 GND.n1943 GND.t826 17.4528
R3062 GND.n1712 GND.t513 17.4528
R3063 GND.n7024 GND.t190 17.4528
R3064 GND.n2388 GND.t711 17.4528
R3065 GND.n2713 GND.t781 17.4528
R3066 GND.n3037 GND.t525 17.4528
R3067 GND.n7110 GND.t800 17.4528
R3068 GND.n4803 GND.t618 17.4528
R3069 GND.n5419 GND.t683 17.4528
R3070 GND.n5914 GND.t1235 17.4528
R3071 GND.n5976 GND.t3 17.4528
R3072 GND.n6143 GND.t1243 17.4528
R3073 GND.n6307 GND.t1146 17.4528
R3074 GND.n595 GND.t1321 17.4528
R3075 GND.n7638 GND.t1137 17.4528
R3076 GND.n7518 GND.t125 17.4528
R3077 GND.n1551 GND.n1550 17.2882
R3078 GND.n4543 GND.t1031 17.2168
R3079 GND GND.t146 17.1372
R3080 GND GND.t1178 17.1372
R3081 GND GND.t144 17.1372
R3082 GND.t1297 GND.t1382 16.9644
R3083 GND.n6676 GND.n6675 16.9417
R3084 GND.n6642 GND.n6641 16.9417
R3085 GND.n6548 GND.n6547 16.9417
R3086 GND.n6489 GND.n6488 16.9417
R3087 GND.n6463 GND.n6462 16.9417
R3088 GND.n4638 GND.n4637 16.9417
R3089 GND.n4745 GND.n4744 16.9417
R3090 GND.n4931 GND.n4930 16.9417
R3091 GND.n5002 GND.n5001 16.9417
R3092 GND.n4602 GND.n4601 16.9417
R3093 GND.n5707 GND.n5706 16.9417
R3094 GND.n5658 GND.n5657 16.9417
R3095 GND.n5636 GND.n5635 16.9417
R3096 GND.n5581 GND.n5580 16.9417
R3097 GND.n5555 GND.n5554 16.9417
R3098 GND.n5208 GND.n5204 16.9417
R3099 GND.n5210 GND.n5184 16.9417
R3100 GND.n4305 GND.n4301 16.9417
R3101 GND.n4307 GND.n4281 16.9417
R3102 GND.n5118 GND.n5117 16.9417
R3103 GND.n5084 GND.n5083 16.9417
R3104 GND.n4555 GND.n4554 16.9417
R3105 GND.n4527 GND.n4526 16.9417
R3106 GND.n4457 GND.n4456 16.9417
R3107 GND GND.t802 16.9356
R3108 GND.t1382 GND 16.3017
R3109 GND.n1895 GND.n1894 16.1887
R3110 GND.n1852 GND.n1851 16.1887
R3111 GND.n7039 GND.n6879 16.1887
R3112 GND.n2501 GND.n2500 16.1887
R3113 GND.n2826 GND.n2825 16.1887
R3114 GND.n3123 GND.n3122 16.1887
R3115 GND.n7223 GND.n7222 16.1887
R3116 GND.n4755 GND.n4754 16.1887
R3117 GND.n5431 GND.n5246 16.1887
R3118 GND.n5923 GND.n5922 16.1887
R3119 GND.n6092 GND.n6091 16.1887
R3120 GND.n6256 GND.n6255 16.1887
R3121 GND.n6565 GND.n6564 16.1887
R3122 GND.n705 GND.n704 16.1887
R3123 GND.n7752 GND.n7751 16.1887
R3124 GND.n7587 GND.n7586 16.1887
R3125 GND.n5195 GND.n5194 16.1887
R3126 GND.n4292 GND.n4291 16.1887
R3127 GND.n7463 GND.n7461 14.7755
R3128 GND.n7467 GND.n7466 14.7755
R3129 GND.n2054 GND.n2049 14.7755
R3130 GND.n1668 GND.n1667 14.7755
R3131 GND.n389 GND.n388 14.7755
R3132 GND.n543 GND.n541 14.7755
R3133 GND.n548 GND.n546 14.7755
R3134 GND.n238 GND.n236 14.7755
R3135 GND.n72 GND.n70 14.7755
R3136 GND.n74 GND.n69 14.7755
R3137 GND.n78 GND.n77 14.7755
R3138 GND.n1412 GND.n1410 14.7755
R3139 GND.n1420 GND.n1415 14.7755
R3140 GND.n1418 GND.n1416 14.7755
R3141 GND.n4247 GND.n4245 14.7755
R3142 GND.n3439 GND.n3438 14.7755
R3143 GND.n3444 GND.n3442 14.7755
R3144 GND.n3282 GND.n3281 14.7755
R3145 GND.n3286 GND.n3285 14.7755
R3146 GND.n2986 GND.n2984 14.7755
R3147 GND.n2990 GND.n2989 14.7755
R3148 GND.n2661 GND.n2659 14.7755
R3149 GND.n2666 GND.n2664 14.7755
R3150 GND.n2336 GND.n2335 14.7755
R3151 GND.n2341 GND.n2339 14.7755
R3152 GND.n2174 GND.n2173 14.7755
R3153 GND.n2183 GND.n2177 14.7755
R3154 GND.n2181 GND.n2178 14.7755
R3155 GND.n1671 GND.n1670 14.7755
R3156 GND.n393 GND.n392 14.7755
R3157 GND.n815 GND.n813 14.7755
R3158 GND.n819 GND.n818 14.7755
R3159 GND.t397 GND.t1305 14.6672
R3160 GND.t1138 GND.t476 14.6672
R3161 GND.t1296 GND.t1304 14.6672
R3162 GND.t351 GND.t349 14.6672
R3163 GND.t659 GND.t515 14.6672
R3164 GND.t696 GND.t705 14.6672
R3165 GND.n6733 GND.n6709 14.5711
R3166 GND.n5764 GND.n5740 14.5711
R3167 GND.n5175 GND.n5151 14.5711
R3168 GND.t687 GND.n1992 14.4569
R3169 GND.t1335 GND.t172 14.3138
R3170 GND.n5647 GND.t1525 14.2308
R3171 GND.n6657 GND.t945 13.8225
R3172 GND.n7816 GND.t1255 13.6894
R3173 GND.n5452 GND.n5449 13.5727
R3174 GND.n6857 GND.n6854 13.5727
R3175 GND.n5452 GND.n5451 13.5705
R3176 GND.n6857 GND.n6856 13.5705
R3177 GND.n5240 GND.n5239 13.5646
R3178 GND.n4332 GND.n4331 13.5646
R3179 GND.n3843 GND.n3842 13.4405
R3180 GND.n4665 GND.t336 13.4015
R3181 GND GND.t1295 13.386
R3182 GND.n5920 GND.n5919 13.3549
R3183 GND.t1530 GND.t1198 12.9885
R3184 GND.t364 GND.t104 12.7234
R3185 GND GND.t1284 12.5248
R3186 GND GND.t42 12.5248
R3187 GND.t566 GND 12.5248
R3188 GND GND.t493 12.5248
R3189 GND GND.t1376 12.5248
R3190 GND GND.t7 12.5248
R3191 GND GND.t1269 12.5248
R3192 GND GND.t753 12.5248
R3193 GND.t1391 GND 12.5248
R3194 GND.t36 GND.n1044 11.9218
R3195 GND.n7348 GND.t36 11.9218
R3196 GND.t1129 GND.n3656 11.9218
R3197 GND.t1358 GND.n4018 11.9218
R3198 GND.t722 GND.n4002 11.9218
R3199 GND.t836 GND.n3987 11.9218
R3200 GND.t726 GND.n3972 11.9218
R3201 GND.t833 GND.n3957 11.9218
R3202 GND.t1356 GND.n3940 11.9218
R3203 GND.t721 GND.n3925 11.9218
R3204 GND.t835 GND.n3910 11.9218
R3205 GND.t725 GND.n3895 11.9218
R3206 GND.t1359 GND.n3878 11.9218
R3207 GND.t727 GND.n3858 11.9218
R3208 GND.t723 GND.n3816 11.9218
R3209 GND.t832 GND.n3801 11.9218
R3210 GND.t729 GND.n3786 11.9218
R3211 GND.t1361 GND.n3771 11.9218
R3212 GND.t724 GND.n3752 11.9218
R3213 GND.t731 GND.n3737 11.9218
R3214 GND.t1357 GND.n3722 11.9218
R3215 GND.t834 GND.n3707 11.9218
R3216 GND.n6672 GND.n6671 11.6711
R3217 GND.n6646 GND.n6645 11.6711
R3218 GND.n6552 GND.n6551 11.6711
R3219 GND.n6485 GND.n6484 11.6711
R3220 GND.n6468 GND.n6467 11.6711
R3221 GND.n4642 GND.n4641 11.6711
R3222 GND.n4704 GND.n4703 11.6711
R3223 GND.n4926 GND.n4925 11.6711
R3224 GND.n5006 GND.n5005 11.6711
R3225 GND.n4598 GND.n4597 11.6711
R3226 GND.n5703 GND.n5702 11.6711
R3227 GND.n5654 GND.n5653 11.6711
R3228 GND.n5640 GND.n5639 11.6711
R3229 GND.n5577 GND.n5576 11.6711
R3230 GND.n5560 GND.n5559 11.6711
R3231 GND.n5114 GND.n5113 11.6711
R3232 GND.n5088 GND.n5087 11.6711
R3233 GND.n4551 GND.n4550 11.6711
R3234 GND.n4531 GND.n4530 11.6711
R3235 GND.n4452 GND.n4451 11.6711
R3236 GND.t730 GND.n3831 11.5107
R3237 GND.n4955 GND.n4954 11.427
R3238 GND.n4953 GND.n4952 11.427
R3239 GND.n6811 GND.n6810 11.427
R3240 GND.n7056 GND.n7055 11.427
R3241 GND.t736 GND.t1530 11.133
R3242 GND.t104 GND.t736 11.133
R3243 GND.t1295 GND.t1335 11.133
R3244 GND GND.t1325 10.9511
R3245 GND GND.t95 10.9511
R3246 GND GND.t761 10.9511
R3247 GND GND.t1204 10.9511
R3248 GND GND.t193 10.9511
R3249 GND GND.t1213 10.9511
R3250 GND GND.t210 10.9511
R3251 GND.n6682 GND.n6681 10.9181
R3252 GND.n6636 GND.n6635 10.9181
R3253 GND.n6542 GND.n6541 10.9181
R3254 GND.n6495 GND.n6494 10.9181
R3255 GND.n6457 GND.n6456 10.9181
R3256 GND.n4611 GND.n4610 10.9181
R3257 GND.n4738 GND.n4737 10.9181
R3258 GND.n4938 GND.n4937 10.9181
R3259 GND.n4996 GND.n4995 10.9181
R3260 GND.n4615 GND.n4614 10.9181
R3261 GND.n5713 GND.n5712 10.9181
R3262 GND.n5664 GND.n5663 10.9181
R3263 GND.n5630 GND.n5629 10.9181
R3264 GND.n5587 GND.n5586 10.9181
R3265 GND.n5549 GND.n5548 10.9181
R3266 GND.n5124 GND.n5123 10.9181
R3267 GND.n5078 GND.n5077 10.9181
R3268 GND.n4561 GND.n4560 10.9181
R3269 GND.n4521 GND.n4520 10.9181
R3270 GND.n4463 GND.n4462 10.9181
R3271 GND.t697 GND 10.6857
R3272 GND.t146 GND 10.6857
R3273 GND.t1178 GND 10.6857
R3274 GND.t802 GND 10.6857
R3275 GND.t144 GND 10.6857
R3276 GND.n4956 GND.n4955 10.5417
R3277 GND.n4163 GND.t392 10.3949
R3278 GND.n6561 GND 10.2053
R3279 GND.n1191 GND.n1188 9.8307
R3280 GND.t119 GND.t89 9.8307
R3281 GND.n1206 GND.n1203 9.8307
R3282 GND.n2216 GND.n2213 9.8307
R3283 GND.t806 GND.t694 9.8307
R3284 GND.n2231 GND.n2228 9.8307
R3285 GND.n2540 GND.n2537 9.8307
R3286 GND.t419 GND.t1308 9.8307
R3287 GND.n2555 GND.n2552 9.8307
R3288 GND.n2865 GND.n2862 9.8307
R3289 GND.t1187 GND.t434 9.8307
R3290 GND.n2880 GND.n2877 9.8307
R3291 GND.n3162 GND.n3159 9.8307
R3292 GND.t186 GND.t94 9.8307
R3293 GND.n3177 GND.n3174 9.8307
R3294 GND.n3319 GND.n3316 9.8307
R3295 GND.t1227 GND.t1367 9.8307
R3296 GND.n3334 GND.n3331 9.8307
R3297 GND.n3477 GND.n3474 9.8307
R3298 GND.t1338 GND.t664 9.8307
R3299 GND.n3492 GND.n3489 9.8307
R3300 GND.n7267 GND.n7264 9.8307
R3301 GND.t1240 GND.t1174 9.8307
R3302 GND.n7282 GND.n7279 9.8307
R3303 GND.n11 GND.n10 9.8307
R3304 GND.t590 GND.t692 9.8307
R3305 GND.n26 GND.n23 9.8307
R3306 GND.n120 GND.n117 9.8307
R3307 GND.t602 GND.t735 9.8307
R3308 GND.n135 GND.n132 9.8307
R3309 GND.n272 GND.n269 9.8307
R3310 GND.t605 GND.t1118 9.8307
R3311 GND.n287 GND.n284 9.8307
R3312 GND.n1635 GND.n1632 9.8307
R3313 GND.t661 GND.t363 9.8307
R3314 GND.n1650 GND.n1647 9.8307
R3315 GND.n425 GND.n422 9.8307
R3316 GND.t13 GND.t850 9.8307
R3317 GND.n440 GND.n437 9.8307
R3318 GND.n744 GND.n741 9.8307
R3319 GND.t819 GND.t1281 9.8307
R3320 GND.n759 GND.n756 9.8307
R3321 GND.n851 GND.n848 9.8307
R3322 GND.t1228 GND.t610 9.8307
R3323 GND.n866 GND.n863 9.8307
R3324 GND.t1275 GND.t1297 9.54267
R3325 GND.t1135 GND.t1275 9.54267
R3326 GND.n5480 GND.n5478 9.41227
R3327 GND.n4411 GND.n4409 9.41227
R3328 GND.n5236 GND.n5235 9.41227
R3329 GND.n4328 GND.n4327 9.41227
R3330 GND.n1925 GND.n1924 9.3005
R3331 GND.n1931 GND.n1930 9.3005
R3332 GND.n1933 GND.n1932 9.3005
R3333 GND.n1927 GND.n1926 9.3005
R3334 GND.n1911 GND.n1910 9.3005
R3335 GND.n1896 GND.n1895 9.3005
R3336 GND.n1559 GND.n1558 9.3005
R3337 GND.n1948 GND.n1947 9.3005
R3338 GND.n1975 GND.n1974 9.3005
R3339 GND.n1950 GND.n1949 9.3005
R3340 GND.n1972 GND.n1971 9.3005
R3341 GND.n1963 GND.n1962 9.3005
R3342 GND.n1961 GND.n1960 9.3005
R3343 GND.n1952 GND.n1951 9.3005
R3344 GND.n1692 GND.n1691 9.3005
R3345 GND.n1698 GND.n1697 9.3005
R3346 GND.n1700 GND.n1699 9.3005
R3347 GND.n1694 GND.n1693 9.3005
R3348 GND.n1868 GND.n1867 9.3005
R3349 GND.n1853 GND.n1852 9.3005
R3350 GND.n1748 GND.n1747 9.3005
R3351 GND.n1743 GND.n1742 9.3005
R3352 GND.n1737 GND.n1736 9.3005
R3353 GND.n1741 GND.n1740 9.3005
R3354 GND.n1734 GND.n1733 9.3005
R3355 GND.n1725 GND.n1724 9.3005
R3356 GND.n1723 GND.n1722 9.3005
R3357 GND.n1714 GND.n1713 9.3005
R3358 GND.n6900 GND.n6899 9.3005
R3359 GND.n6906 GND.n6905 9.3005
R3360 GND.n6908 GND.n6907 9.3005
R3361 GND.n6902 GND.n6901 9.3005
R3362 GND.n6889 GND.n6888 9.3005
R3363 GND.n7040 GND.n7039 9.3005
R3364 GND.n7020 GND.n7019 9.3005
R3365 GND.n7015 GND.n7014 9.3005
R3366 GND.n1833 GND.n1832 9.3005
R3367 GND.n7013 GND.n7012 9.3005
R3368 GND.n1830 GND.n1829 9.3005
R3369 GND.n1821 GND.n1820 9.3005
R3370 GND.n1819 GND.n1818 9.3005
R3371 GND.n1810 GND.n1809 9.3005
R3372 GND.n2368 GND.n2367 9.3005
R3373 GND.n2374 GND.n2373 9.3005
R3374 GND.n2376 GND.n2375 9.3005
R3375 GND.n2370 GND.n2369 9.3005
R3376 GND.n2517 GND.n2516 9.3005
R3377 GND.n2502 GND.n2501 9.3005
R3378 GND.n2397 GND.n2396 9.3005
R3379 GND.n2392 GND.n2391 9.3005
R3380 GND.n6998 GND.n6997 9.3005
R3381 GND.n2390 GND.n2389 9.3005
R3382 GND.n6995 GND.n6994 9.3005
R3383 GND.n6986 GND.n6985 9.3005
R3384 GND.n6984 GND.n6983 9.3005
R3385 GND.n6975 GND.n6974 9.3005
R3386 GND.n2693 GND.n2692 9.3005
R3387 GND.n2699 GND.n2698 9.3005
R3388 GND.n2701 GND.n2700 9.3005
R3389 GND.n2695 GND.n2694 9.3005
R3390 GND.n2842 GND.n2841 9.3005
R3391 GND.n2827 GND.n2826 9.3005
R3392 GND.n2722 GND.n2721 9.3005
R3393 GND.n2717 GND.n2716 9.3005
R3394 GND.n2482 GND.n2481 9.3005
R3395 GND.n2715 GND.n2714 9.3005
R3396 GND.n2479 GND.n2478 9.3005
R3397 GND.n2470 GND.n2469 9.3005
R3398 GND.n2468 GND.n2467 9.3005
R3399 GND.n2459 GND.n2458 9.3005
R3400 GND.n3017 GND.n3016 9.3005
R3401 GND.n3023 GND.n3022 9.3005
R3402 GND.n3025 GND.n3024 9.3005
R3403 GND.n3019 GND.n3018 9.3005
R3404 GND.n3139 GND.n3138 9.3005
R3405 GND.n3124 GND.n3123 9.3005
R3406 GND.n3046 GND.n3045 9.3005
R3407 GND.n3041 GND.n3040 9.3005
R3408 GND.n2807 GND.n2806 9.3005
R3409 GND.n3039 GND.n3038 9.3005
R3410 GND.n2804 GND.n2803 9.3005
R3411 GND.n2795 GND.n2794 9.3005
R3412 GND.n2793 GND.n2792 9.3005
R3413 GND.n2784 GND.n2783 9.3005
R3414 GND.n7090 GND.n7089 9.3005
R3415 GND.n7096 GND.n7095 9.3005
R3416 GND.n7098 GND.n7097 9.3005
R3417 GND.n7092 GND.n7091 9.3005
R3418 GND.n7239 GND.n7238 9.3005
R3419 GND.n7224 GND.n7223 9.3005
R3420 GND.n7146 GND.n7145 9.3005
R3421 GND.n7141 GND.n7140 9.3005
R3422 GND.n7135 GND.n7134 9.3005
R3423 GND.n7139 GND.n7138 9.3005
R3424 GND.n7132 GND.n7131 9.3005
R3425 GND.n7123 GND.n7122 9.3005
R3426 GND.n7121 GND.n7120 9.3005
R3427 GND.n7112 GND.n7111 9.3005
R3428 GND.n4785 GND.n4784 9.3005
R3429 GND.n4791 GND.n4790 9.3005
R3430 GND.n4793 GND.n4792 9.3005
R3431 GND.n4787 GND.n4786 9.3005
R3432 GND.n4771 GND.n4770 9.3005
R3433 GND.n4756 GND.n4755 9.3005
R3434 GND.n4839 GND.n4838 9.3005
R3435 GND.n4834 GND.n4833 9.3005
R3436 GND.n4828 GND.n4827 9.3005
R3437 GND.n4832 GND.n4831 9.3005
R3438 GND.n4825 GND.n4824 9.3005
R3439 GND.n4816 GND.n4815 9.3005
R3440 GND.n4814 GND.n4813 9.3005
R3441 GND.n4805 GND.n4804 9.3005
R3442 GND.n5267 GND.n5266 9.3005
R3443 GND.n5273 GND.n5272 9.3005
R3444 GND.n5275 GND.n5274 9.3005
R3445 GND.n5269 GND.n5268 9.3005
R3446 GND.n5256 GND.n5255 9.3005
R3447 GND.n5432 GND.n5431 9.3005
R3448 GND.n5415 GND.n5414 9.3005
R3449 GND.n5410 GND.n5409 9.3005
R3450 GND.n5404 GND.n5403 9.3005
R3451 GND.n5408 GND.n5407 9.3005
R3452 GND.n5401 GND.n5400 9.3005
R3453 GND.n5392 GND.n5391 9.3005
R3454 GND.n5390 GND.n5389 9.3005
R3455 GND.n5381 GND.n5380 9.3005
R3456 GND.n5789 GND.n5788 9.3005
R3457 GND.n5795 GND.n5794 9.3005
R3458 GND.n5797 GND.n5796 9.3005
R3459 GND.n5791 GND.n5790 9.3005
R3460 GND.n5939 GND.n5938 9.3005
R3461 GND.n5924 GND.n5923 9.3005
R3462 GND.n5910 GND.n5909 9.3005
R3463 GND.n5905 GND.n5904 9.3005
R3464 GND.n5365 GND.n5364 9.3005
R3465 GND.n5903 GND.n5902 9.3005
R3466 GND.n5362 GND.n5361 9.3005
R3467 GND.n5353 GND.n5352 9.3005
R3468 GND.n5351 GND.n5350 9.3005
R3469 GND.n5342 GND.n5341 9.3005
R3470 GND.n5956 GND.n5955 9.3005
R3471 GND.n5962 GND.n5961 9.3005
R3472 GND.n5964 GND.n5963 9.3005
R3473 GND.n5958 GND.n5957 9.3005
R3474 GND.n6108 GND.n6107 9.3005
R3475 GND.n6093 GND.n6092 9.3005
R3476 GND.n5985 GND.n5984 9.3005
R3477 GND.n5980 GND.n5979 9.3005
R3478 GND.n5887 GND.n5886 9.3005
R3479 GND.n5978 GND.n5977 9.3005
R3480 GND.n5884 GND.n5883 9.3005
R3481 GND.n5875 GND.n5874 9.3005
R3482 GND.n5873 GND.n5872 9.3005
R3483 GND.n5864 GND.n5863 9.3005
R3484 GND.n6123 GND.n6122 9.3005
R3485 GND.n6129 GND.n6128 9.3005
R3486 GND.n6131 GND.n6130 9.3005
R3487 GND.n6125 GND.n6124 9.3005
R3488 GND.n6272 GND.n6271 9.3005
R3489 GND.n6257 GND.n6256 9.3005
R3490 GND.n6152 GND.n6151 9.3005
R3491 GND.n6147 GND.n6146 9.3005
R3492 GND.n6073 GND.n6072 9.3005
R3493 GND.n6145 GND.n6144 9.3005
R3494 GND.n6070 GND.n6069 9.3005
R3495 GND.n6061 GND.n6060 9.3005
R3496 GND.n6059 GND.n6058 9.3005
R3497 GND.n6050 GND.n6049 9.3005
R3498 GND.n6287 GND.n6286 9.3005
R3499 GND.n6293 GND.n6292 9.3005
R3500 GND.n6295 GND.n6294 9.3005
R3501 GND.n6289 GND.n6288 9.3005
R3502 GND.n6581 GND.n6580 9.3005
R3503 GND.n6566 GND.n6565 9.3005
R3504 GND.n6316 GND.n6315 9.3005
R3505 GND.n6311 GND.n6310 9.3005
R3506 GND.n6237 GND.n6236 9.3005
R3507 GND.n6309 GND.n6308 9.3005
R3508 GND.n6234 GND.n6233 9.3005
R3509 GND.n6225 GND.n6224 9.3005
R3510 GND.n6223 GND.n6222 9.3005
R3511 GND.n6214 GND.n6213 9.3005
R3512 GND.n575 GND.n574 9.3005
R3513 GND.n581 GND.n580 9.3005
R3514 GND.n583 GND.n582 9.3005
R3515 GND.n577 GND.n576 9.3005
R3516 GND.n721 GND.n720 9.3005
R3517 GND.n706 GND.n705 9.3005
R3518 GND.n604 GND.n603 9.3005
R3519 GND.n599 GND.n598 9.3005
R3520 GND.n6401 GND.n6400 9.3005
R3521 GND.n597 GND.n596 9.3005
R3522 GND.n6398 GND.n6397 9.3005
R3523 GND.n6389 GND.n6388 9.3005
R3524 GND.n6387 GND.n6386 9.3005
R3525 GND.n6378 GND.n6377 9.3005
R3526 GND.n7618 GND.n7617 9.3005
R3527 GND.n7624 GND.n7623 9.3005
R3528 GND.n7626 GND.n7625 9.3005
R3529 GND.n7620 GND.n7619 9.3005
R3530 GND.n7768 GND.n7767 9.3005
R3531 GND.n7753 GND.n7752 9.3005
R3532 GND.n7647 GND.n7646 9.3005
R3533 GND.n7642 GND.n7641 9.3005
R3534 GND.n686 GND.n685 9.3005
R3535 GND.n7640 GND.n7639 9.3005
R3536 GND.n683 GND.n682 9.3005
R3537 GND.n674 GND.n673 9.3005
R3538 GND.n672 GND.n671 9.3005
R3539 GND.n663 GND.n662 9.3005
R3540 GND.n1437 GND.n1436 9.3005
R3541 GND.n3461 GND.n3460 9.3005
R3542 GND.n3007 GND.n3006 9.3005
R3543 GND.n2358 GND.n2357 9.3005
R3544 GND.n1319 GND.n1318 9.3005
R3545 GND.n1318 GND.n1317 9.3005
R3546 GND.n2200 GND.n2199 9.3005
R3547 GND.n2683 GND.n2682 9.3005
R3548 GND.n3303 GND.n3302 9.3005
R3549 GND.n4264 GND.n4263 9.3005
R3550 GND.n104 GND.n103 9.3005
R3551 GND.n256 GND.n255 9.3005
R3552 GND.n410 GND.n409 9.3005
R3553 GND.n409 GND.n408 9.3005
R3554 GND.n2078 GND.n2077 9.3005
R3555 GND.n2077 GND.n2076 9.3005
R3556 GND.n3767 GND.n3766 9.3005
R3557 GND.n3679 GND.n3678 9.3005
R3558 GND.n3650 GND.n3649 9.3005
R3559 GND.n3954 GND.n3953 9.3005
R3560 GND.n4044 GND.n4043 9.3005
R3561 GND.n836 GND.n835 9.3005
R3562 GND.n835 GND.n834 9.3005
R3563 GND.n565 GND.n564 9.3005
R3564 GND.n7488 GND.n7487 9.3005
R3565 GND.n7498 GND.n7497 9.3005
R3566 GND.n7504 GND.n7503 9.3005
R3567 GND.n7506 GND.n7505 9.3005
R3568 GND.n7500 GND.n7499 9.3005
R3569 GND.n7603 GND.n7602 9.3005
R3570 GND.n7588 GND.n7587 9.3005
R3571 GND.n7527 GND.n7526 9.3005
R3572 GND.n7522 GND.n7521 9.3005
R3573 GND.n7733 GND.n7732 9.3005
R3574 GND.n7520 GND.n7519 9.3005
R3575 GND.n7730 GND.n7729 9.3005
R3576 GND.n7721 GND.n7720 9.3005
R3577 GND.n7719 GND.n7718 9.3005
R3578 GND.n7710 GND.n7709 9.3005
R3579 GND.n7535 GND.n7534 9.3005
R3580 GND.n7580 GND.n7579 9.3005
R3581 GND.n7570 GND.n7569 9.3005
R3582 GND.n7549 GND.n7548 9.3005
R3583 GND.n7558 GND.n7557 9.3005
R3584 GND.n7540 GND.n7539 9.3005
R3585 GND.n7547 GND.n7546 9.3005
R3586 GND.n7666 GND.n7665 9.3005
R3587 GND.n7744 GND.n7743 9.3005
R3588 GND.n7706 GND.n7705 9.3005
R3589 GND.n7680 GND.n7679 9.3005
R3590 GND.n7689 GND.n7688 9.3005
R3591 GND.n7671 GND.n7670 9.3005
R3592 GND.n7678 GND.n7677 9.3005
R3593 GND.n622 GND.n621 9.3005
R3594 GND.n697 GND.n696 9.3005
R3595 GND.n659 GND.n658 9.3005
R3596 GND.n633 GND.n632 9.3005
R3597 GND.n642 GND.n641 9.3005
R3598 GND.n624 GND.n623 9.3005
R3599 GND.n631 GND.n630 9.3005
R3600 GND.n6334 GND.n6333 9.3005
R3601 GND.n6412 GND.n6411 9.3005
R3602 GND.n6371 GND.n6370 9.3005
R3603 GND.n6345 GND.n6344 9.3005
R3604 GND.n6354 GND.n6353 9.3005
R3605 GND.n6336 GND.n6335 9.3005
R3606 GND.n6343 GND.n6342 9.3005
R3607 GND.n6170 GND.n6169 9.3005
R3608 GND.n6248 GND.n6247 9.3005
R3609 GND.n6207 GND.n6206 9.3005
R3610 GND.n6181 GND.n6180 9.3005
R3611 GND.n6190 GND.n6189 9.3005
R3612 GND.n6172 GND.n6171 9.3005
R3613 GND.n6179 GND.n6178 9.3005
R3614 GND.n6003 GND.n6002 9.3005
R3615 GND.n6084 GND.n6083 9.3005
R3616 GND.n6043 GND.n6042 9.3005
R3617 GND.n6017 GND.n6016 9.3005
R3618 GND.n6026 GND.n6025 9.3005
R3619 GND.n6008 GND.n6007 9.3005
R3620 GND.n6015 GND.n6014 9.3005
R3621 GND.n5820 GND.n5819 9.3005
R3622 GND.n5900 GND.n5899 9.3005
R3623 GND.n5860 GND.n5859 9.3005
R3624 GND.n5834 GND.n5833 9.3005
R3625 GND.n5843 GND.n5842 9.3005
R3626 GND.n5825 GND.n5824 9.3005
R3627 GND.n5832 GND.n5831 9.3005
R3628 GND.n5298 GND.n5297 9.3005
R3629 GND.n5378 GND.n5377 9.3005
R3630 GND.n5338 GND.n5337 9.3005
R3631 GND.n5312 GND.n5311 9.3005
R3632 GND.n5321 GND.n5320 9.3005
R3633 GND.n5303 GND.n5302 9.3005
R3634 GND.n5310 GND.n5309 9.3005
R3635 GND.n4857 GND.n4856 9.3005
R3636 GND.n4908 GND.n4907 9.3005
R3637 GND.n4897 GND.n4896 9.3005
R3638 GND.n4871 GND.n4870 9.3005
R3639 GND.n4880 GND.n4879 9.3005
R3640 GND.n4862 GND.n4861 9.3005
R3641 GND.n4869 GND.n4868 9.3005
R3642 GND.n7164 GND.n7163 9.3005
R3643 GND.n7215 GND.n7214 9.3005
R3644 GND.n7204 GND.n7203 9.3005
R3645 GND.n7178 GND.n7177 9.3005
R3646 GND.n7187 GND.n7186 9.3005
R3647 GND.n7169 GND.n7168 9.3005
R3648 GND.n7176 GND.n7175 9.3005
R3649 GND.n3064 GND.n3063 9.3005
R3650 GND.n3115 GND.n3114 9.3005
R3651 GND.n3104 GND.n3103 9.3005
R3652 GND.n3078 GND.n3077 9.3005
R3653 GND.n3087 GND.n3086 9.3005
R3654 GND.n3069 GND.n3068 9.3005
R3655 GND.n3076 GND.n3075 9.3005
R3656 GND.n2740 GND.n2739 9.3005
R3657 GND.n2818 GND.n2817 9.3005
R3658 GND.n2780 GND.n2779 9.3005
R3659 GND.n2754 GND.n2753 9.3005
R3660 GND.n2763 GND.n2762 9.3005
R3661 GND.n2745 GND.n2744 9.3005
R3662 GND.n2752 GND.n2751 9.3005
R3663 GND.n2415 GND.n2414 9.3005
R3664 GND.n2493 GND.n2492 9.3005
R3665 GND.n2455 GND.n2454 9.3005
R3666 GND.n2429 GND.n2428 9.3005
R3667 GND.n2438 GND.n2437 9.3005
R3668 GND.n2420 GND.n2419 9.3005
R3669 GND.n2427 GND.n2426 9.3005
R3670 GND.n6931 GND.n6930 9.3005
R3671 GND.n7010 GND.n7009 9.3005
R3672 GND.n6971 GND.n6970 9.3005
R3673 GND.n6945 GND.n6944 9.3005
R3674 GND.n6954 GND.n6953 9.3005
R3675 GND.n6936 GND.n6935 9.3005
R3676 GND.n6943 GND.n6942 9.3005
R3677 GND.n1766 GND.n1765 9.3005
R3678 GND.n1844 GND.n1843 9.3005
R3679 GND.n1806 GND.n1805 9.3005
R3680 GND.n1780 GND.n1779 9.3005
R3681 GND.n1789 GND.n1788 9.3005
R3682 GND.n1771 GND.n1770 9.3005
R3683 GND.n1778 GND.n1777 9.3005
R3684 GND.n1575 GND.n1574 9.3005
R3685 GND.n1887 GND.n1886 9.3005
R3686 GND.n1615 GND.n1614 9.3005
R3687 GND.n1589 GND.n1588 9.3005
R3688 GND.n1598 GND.n1597 9.3005
R3689 GND.n1580 GND.n1579 9.3005
R3690 GND.n1587 GND.n1586 9.3005
R3691 GND.n7487 GND.n7485 9.1766
R3692 GND.n564 GND.n562 9.1766
R3693 GND.n255 GND.n253 9.1766
R3694 GND.n103 GND.n101 9.1766
R3695 GND.n1436 GND.n1434 9.1766
R3696 GND.n4263 GND.n4261 9.1766
R3697 GND.n3460 GND.n3458 9.1766
R3698 GND.n3302 GND.n3300 9.1766
R3699 GND.n3006 GND.n3004 9.1766
R3700 GND.n2682 GND.n2680 9.1766
R3701 GND.n2357 GND.n2355 9.1766
R3702 GND.n2199 GND.n2197 9.1766
R3703 GND.n1192 GND.n1191 8.84768
R3704 GND.n2217 GND.n2216 8.84768
R3705 GND.n2541 GND.n2540 8.84768
R3706 GND.n2866 GND.n2865 8.84768
R3707 GND.n3163 GND.n3162 8.84768
R3708 GND.n3320 GND.n3319 8.84768
R3709 GND.n3478 GND.n3477 8.84768
R3710 GND.n7268 GND.n7267 8.84768
R3711 GND.n12 GND.n11 8.84768
R3712 GND.n121 GND.n120 8.84768
R3713 GND.n273 GND.n272 8.84768
R3714 GND.n1636 GND.n1635 8.84768
R3715 GND.n426 GND.n425 8.84768
R3716 GND.n745 GND.n744 8.84768
R3717 GND.n852 GND.n851 8.84768
R3718 GND.n1560 GND.t72 8.70904
R3719 GND.n1749 GND.t375 8.70904
R3720 GND.n7021 GND.t1211 8.70904
R3721 GND.n2398 GND.t655 8.70904
R3722 GND.n2723 GND.t1247 8.70904
R3723 GND.n3047 GND.t1259 8.70904
R3724 GND.n7147 GND.t584 8.70904
R3725 GND.n4840 GND.t184 8.70904
R3726 GND.n5416 GND.t527 8.70904
R3727 GND.n5911 GND.t822 8.70904
R3728 GND.n5986 GND.t32 8.70904
R3729 GND.n6153 GND.t718 8.70904
R3730 GND.n6317 GND.t1212 8.70904
R3731 GND.n605 GND.t503 8.70904
R3732 GND.n7648 GND.t359 8.70904
R3733 GND.n7528 GND.t1371 8.70904
R3734 GND.n1573 GND.t1121 8.70236
R3735 GND.n1764 GND.t783 8.70236
R3736 GND.n6929 GND.t1346 8.70236
R3737 GND.n2413 GND.t1197 8.70236
R3738 GND.n2738 GND.t852 8.70236
R3739 GND.n3062 GND.t1390 8.70236
R3740 GND.n7162 GND.t674 8.70236
R3741 GND.n4855 GND.t757 8.70236
R3742 GND.n5296 GND.t1400 8.70236
R3743 GND.n5818 GND.t1334 8.70236
R3744 GND.n6001 GND.t171 8.70236
R3745 GND.n6168 GND.t157 8.70236
R3746 GND.n6332 GND.t188 8.70236
R3747 GND.n620 GND.t201 8.70236
R3748 GND.n7664 GND.t437 8.70236
R3749 GND.n7533 GND.t520 8.70236
R3750 GND GND.t1135 8.61496
R3751 GND GND.t364 8.48243
R3752 GND.t1141 GND.t124 8.20945
R3753 GND.t1232 GND.t1136 8.20945
R3754 GND.t1183 GND.t1320 8.20945
R3755 GND.t1115 GND.t1145 8.20945
R3756 GND.t18 GND.t1242 8.20945
R3757 GND.t744 GND.t2 8.20945
R3758 GND.t478 GND.t1234 8.20945
R3759 GND.t1309 GND.t682 8.20945
R3760 GND.t521 GND.t617 8.20945
R3761 GND.t828 GND.t799 8.20945
R3762 GND.t142 GND.t524 8.20945
R3763 GND.t815 GND.t780 8.20945
R3764 GND.t804 GND.t710 8.20945
R3765 GND.t774 GND.t189 8.20945
R3766 GND.t1344 GND.t512 8.20945
R3767 GND.t517 GND.t825 8.20945
R3768 GND.n7360 GND 8.05791
R3769 GND.n2013 GND 8.05791
R3770 GND.n511 GND 8.05791
R3771 GND.n206 GND 8.05791
R3772 GND.n1505 GND 8.05791
R3773 GND.n1457 GND 8.05791
R3774 GND.n4214 GND 8.05791
R3775 GND.n3408 GND 8.05791
R3776 GND.n3251 GND 8.05791
R3777 GND.n2954 GND 8.05791
R3778 GND.n2629 GND 8.05791
R3779 GND.n2305 GND 8.05791
R3780 GND.n2143 GND 8.05791
R3781 GND.n1275 GND 8.05791
R3782 GND.n358 GND 8.05791
R3783 GND.n7406 GND 8.05791
R3784 GND.t1246 GND.n3839 8.04588
R3785 GND.n7358 GND.n7357 7.90638
R3786 GND.n2011 GND.n2010 7.90638
R3787 GND.n356 GND.n355 7.90638
R3788 GND.n509 GND.n508 7.90638
R3789 GND.n204 GND.n203 7.90638
R3790 GND.n1503 GND.n1502 7.90638
R3791 GND.n1455 GND.n1454 7.90638
R3792 GND.n4212 GND.n4211 7.90638
R3793 GND.n3406 GND.n3405 7.90638
R3794 GND.n3249 GND.n3248 7.90638
R3795 GND.n2952 GND.n2951 7.90638
R3796 GND.n2627 GND.n2626 7.90638
R3797 GND.n2303 GND.n2302 7.90638
R3798 GND.n2141 GND.n2140 7.90638
R3799 GND.n1273 GND.n1272 7.90638
R3800 GND.n7404 GND.n7403 7.90638
R3801 GND GND.n7044 7.56079
R3802 GND.n5099 GND.t1003 7.37892
R3803 GND.n1228 GND.t402 6.88164
R3804 GND.n2253 GND.t1162 6.88164
R3805 GND.n2577 GND.t830 6.88164
R3806 GND.n2902 GND.t840 6.88164
R3807 GND.n3199 GND.t1166 6.88164
R3808 GND.n3356 GND.t585 6.88164
R3809 GND.n3514 GND.t1257 6.88164
R3810 GND.n7304 GND.t158 6.88164
R3811 GND.n48 GND.t400 6.88164
R3812 GND.n157 GND.t1159 6.88164
R3813 GND.n309 GND.t588 6.88164
R3814 GND.n1680 GND.t598 6.88164
R3815 GND.n462 GND.t838 6.88164
R3816 GND.n781 GND.t1164 6.88164
R3817 GND.n888 GND.t685 6.88164
R3818 GND.n6725 GND.n6712 6.77697
R3819 GND.n5756 GND.n5743 6.77697
R3820 GND.n6834 GND.n6806 6.77697
R3821 GND.n6828 GND.n6807 6.77697
R3822 GND.n6822 GND.n6808 6.77697
R3823 GND.n6816 GND.n6809 6.77697
R3824 GND.n7079 GND.n7051 6.77697
R3825 GND.n7073 GND.n7052 6.77697
R3826 GND.n7067 GND.n7053 6.77697
R3827 GND.n7061 GND.n7054 6.77697
R3828 GND.n5167 GND.n5154 6.77697
R3829 GND.t294 GND.n4664 6.70101
R3830 GND.n2065 GND.n2064 6.52989
R3831 GND.n397 GND.n396 6.52989
R3832 GND.n823 GND.n822 6.52989
R3833 GND.n7471 GND.n7470 6.5285
R3834 GND.n552 GND.n551 6.5285
R3835 GND.n243 GND.n242 6.5285
R3836 GND.n82 GND.n81 6.5285
R3837 GND.n1424 GND.n1423 6.5285
R3838 GND.n4251 GND.n4250 6.5285
R3839 GND.n3448 GND.n3447 6.5285
R3840 GND.n3290 GND.n3289 6.5285
R3841 GND.n2994 GND.n2993 6.5285
R3842 GND.n2670 GND.n2669 6.5285
R3843 GND.n2345 GND.n2344 6.5285
R3844 GND.n2187 GND.n2186 6.5285
R3845 GND.n1306 GND.n1305 6.5285
R3846 GND.n5481 GND.n5480 6.4005
R3847 GND.n4412 GND.n4411 6.4005
R3848 GND.n5454 GND.n5449 6.4005
R3849 GND.n5451 GND.n5446 6.4005
R3850 GND.n5235 GND.n5223 6.4005
R3851 GND.n5241 GND.n5240 6.4005
R3852 GND.n6859 GND.n6854 6.4005
R3853 GND.n6856 GND.n6851 6.4005
R3854 GND.n4327 GND.n4315 6.4005
R3855 GND.n4333 GND.n4332 6.4005
R3856 GND.n6714 GND.n6713 6.15638
R3857 GND.n5745 GND.n5744 6.15638
R3858 GND.n5156 GND.n5155 6.15638
R3859 GND.n6666 GND.n6665 5.64756
R3860 GND.n6653 GND.n6652 5.64756
R3861 GND.n6526 GND.n6525 5.64756
R3862 GND.n6478 GND.n6477 5.64756
R3863 GND.n6426 GND.n6425 5.64756
R3864 GND.n7378 GND 5.64756
R3865 GND.n1374 GND 5.64756
R3866 GND.n336 GND 5.64756
R3867 GND.n489 GND 5.64756
R3868 GND.n184 GND 5.64756
R3869 GND.n1519 GND 5.64756
R3870 GND.n1471 GND 5.64756
R3871 GND.n4192 GND 5.64756
R3872 GND.n3386 GND 5.64756
R3873 GND.n3229 GND 5.64756
R3874 GND.n2932 GND 5.64756
R3875 GND.n2607 GND 5.64756
R3876 GND.n2283 GND 5.64756
R3877 GND.n2121 GND 5.64756
R3878 GND.n1253 GND 5.64756
R3879 GND.n7420 GND 5.64756
R3880 GND.n4648 GND.n4647 5.64756
R3881 GND.n4697 GND.n4696 5.64756
R3882 GND.n4710 GND.n4709 5.64756
R3883 GND.n5013 GND.n5012 5.64756
R3884 GND.n4592 GND.n4591 5.64756
R3885 GND.n5697 GND.n5696 5.64756
R3886 GND.n5505 GND.n5504 5.64756
R3887 GND.n5618 GND.n5617 5.64756
R3888 GND.n5570 GND.n5569 5.64756
R3889 GND.n5517 GND.n5516 5.64756
R3890 GND.n5108 GND.n5107 5.64756
R3891 GND.n5095 GND.n5094 5.64756
R3892 GND.n4433 GND.n4432 5.64756
R3893 GND.n4538 GND.n4537 5.64756
R3894 GND.n4442 GND.n4441 5.64756
R3895 GND.n7712 GND.n7711 5.62907
R3896 GND.n665 GND.n664 5.62907
R3897 GND.n6380 GND.n6379 5.62907
R3898 GND.n6216 GND.n6215 5.62907
R3899 GND.n6052 GND.n6051 5.62907
R3900 GND.n5866 GND.n5865 5.62907
R3901 GND.n5344 GND.n5343 5.62907
R3902 GND.n5383 GND.n5382 5.62907
R3903 GND.n4807 GND.n4806 5.62907
R3904 GND.n7114 GND.n7113 5.62907
R3905 GND.n2786 GND.n2785 5.62907
R3906 GND.n2461 GND.n2460 5.62907
R3907 GND.n6977 GND.n6976 5.62907
R3908 GND.n1812 GND.n1811 5.62907
R3909 GND.n1716 GND.n1715 5.62907
R3910 GND.n1954 GND.n1953 5.62907
R3911 GND.n7818 GND.n7798 5.1205
R3912 GND.n890 GND.n859 5.1205
R3913 GND.n783 GND.n752 5.1205
R3914 GND.n464 GND.n433 5.1205
R3915 GND.n1682 GND.n1643 5.1205
R3916 GND.n311 GND.n280 5.1205
R3917 GND.n159 GND.n128 5.1205
R3918 GND.n50 GND.n19 5.1205
R3919 GND.n7306 GND.n7275 5.1205
R3920 GND.n3516 GND.n3485 5.1205
R3921 GND.n3358 GND.n3327 5.1205
R3922 GND.n3201 GND.n3170 5.1205
R3923 GND.n2904 GND.n2873 5.1205
R3924 GND.n2579 GND.n2548 5.1205
R3925 GND.n2255 GND.n2224 5.1205
R3926 GND.n1230 GND.n1199 5.1205
R3927 GND.n3764 GND.n3763 4.90717
R3928 GND.n6688 GND.n6687 4.89462
R3929 GND.n6630 GND.n6629 4.89462
R3930 GND.n6536 GND.n6535 4.89462
R3931 GND.n6501 GND.n6500 4.89462
R3932 GND.n6451 GND.n6450 4.89462
R3933 GND.n4673 GND.n4672 4.89462
R3934 GND.n4732 GND.n4731 4.89462
R3935 GND.n4944 GND.n4943 4.89462
R3936 GND.n4990 GND.n4989 4.89462
R3937 GND.n4621 GND.n4620 4.89462
R3938 GND.n5719 GND.n5718 4.89462
R3939 GND.n5670 GND.n5669 4.89462
R3940 GND.n5624 GND.n5623 4.89462
R3941 GND.n5593 GND.n5592 4.89462
R3942 GND.n5543 GND.n5542 4.89462
R3943 GND.n5130 GND.n5129 4.89462
R3944 GND.n5072 GND.n5071 4.89462
R3945 GND.n4567 GND.n4566 4.89462
R3946 GND.n4515 GND.n4514 4.89462
R3947 GND.n4469 GND.n4468 4.89462
R3948 GND.n3855 GND.t728 4.78444
R3949 GND.n1929 GND 4.66821
R3950 GND.n1696 GND 4.66821
R3951 GND.n6904 GND 4.66821
R3952 GND.n2372 GND 4.66821
R3953 GND.n2697 GND 4.66821
R3954 GND.n3021 GND 4.66821
R3955 GND.n7094 GND 4.66821
R3956 GND.n4789 GND 4.66821
R3957 GND.n5271 GND 4.66821
R3958 GND.n5793 GND 4.66821
R3959 GND.n5960 GND 4.66821
R3960 GND.n6127 GND 4.66821
R3961 GND.n6291 GND 4.66821
R3962 GND.n579 GND 4.66821
R3963 GND.n7622 GND 4.66821
R3964 GND.n7502 GND 4.66821
R3965 GND.n5475 GND.n5468 4.6505
R3966 GND.n5486 GND.n5465 4.6505
R3967 GND.n5485 GND.n5484 4.6505
R3968 GND.n5483 GND.n5466 4.6505
R3969 GND.n5482 GND.n5481 4.6505
R3970 GND.n5478 GND.n5467 4.6505
R3971 GND.n5477 GND.n5476 4.6505
R3972 GND.n5474 GND.n5473 4.6505
R3973 GND.n1923 GND.n1922 4.6505
R3974 GND.n1894 GND.n1893 4.6505
R3975 GND.n1909 GND.n1908 4.6505
R3976 GND.n1690 GND.n1689 4.6505
R3977 GND.n1851 GND.n1850 4.6505
R3978 GND.n1866 GND.n1865 4.6505
R3979 GND.n6898 GND.n6897 4.6505
R3980 GND.n7041 GND.n6879 4.6505
R3981 GND.n6887 GND.n6886 4.6505
R3982 GND.n2366 GND.n2365 4.6505
R3983 GND.n2500 GND.n2499 4.6505
R3984 GND.n2515 GND.n2514 4.6505
R3985 GND.n2691 GND.n2690 4.6505
R3986 GND.n2825 GND.n2824 4.6505
R3987 GND.n2840 GND.n2839 4.6505
R3988 GND.n3015 GND.n3014 4.6505
R3989 GND.n3122 GND.n3121 4.6505
R3990 GND.n3137 GND.n3136 4.6505
R3991 GND.n7088 GND.n7087 4.6505
R3992 GND.n7222 GND.n7221 4.6505
R3993 GND.n7237 GND.n7236 4.6505
R3994 GND.n4783 GND.n4782 4.6505
R3995 GND.n4754 GND.n4753 4.6505
R3996 GND.n4769 GND.n4768 4.6505
R3997 GND.n5265 GND.n5264 4.6505
R3998 GND.n5433 GND.n5246 4.6505
R3999 GND.n5254 GND.n5253 4.6505
R4000 GND.n5787 GND.n5786 4.6505
R4001 GND.n5922 GND.n5921 4.6505
R4002 GND.n5937 GND.n5936 4.6505
R4003 GND.n5954 GND.n5953 4.6505
R4004 GND.n6091 GND.n6090 4.6505
R4005 GND.n6106 GND.n6105 4.6505
R4006 GND.n6121 GND.n6120 4.6505
R4007 GND.n6255 GND.n6254 4.6505
R4008 GND.n6270 GND.n6269 4.6505
R4009 GND.n6285 GND.n6284 4.6505
R4010 GND.n6564 GND.n6563 4.6505
R4011 GND.n6579 GND.n6578 4.6505
R4012 GND.n573 GND.n572 4.6505
R4013 GND.n704 GND.n703 4.6505
R4014 GND.n719 GND.n718 4.6505
R4015 GND.n7616 GND.n7615 4.6505
R4016 GND.n7751 GND.n7750 4.6505
R4017 GND.n7766 GND.n7765 4.6505
R4018 GND.n7496 GND.n7495 4.6505
R4019 GND.n7586 GND.n7585 4.6505
R4020 GND.n7601 GND.n7600 4.6505
R4021 GND.n4406 GND.n4399 4.6505
R4022 GND.n4417 GND.n4396 4.6505
R4023 GND.n4416 GND.n4415 4.6505
R4024 GND.n4414 GND.n4397 4.6505
R4025 GND.n4413 GND.n4412 4.6505
R4026 GND.n4409 GND.n4398 4.6505
R4027 GND.n4408 GND.n4407 4.6505
R4028 GND.n4405 GND.n4404 4.6505
R4029 GND.n4958 GND.n4951 4.6505
R4030 GND.n4970 GND.n4949 4.6505
R4031 GND.n4962 GND.n4950 4.6505
R4032 GND.n4969 GND.n4968 4.6505
R4033 GND.n4967 GND.n4966 4.6505
R4034 GND.n4964 GND.n4963 4.6505
R4035 GND.n4960 GND.n4959 4.6505
R4036 GND.n4957 GND.n4956 4.6505
R4037 GND.n5028 GND.n4946 4.6505
R4038 GND.n5027 GND.n4947 4.6505
R4039 GND.n4972 GND.n4948 4.6505
R4040 GND.n5026 GND.n5025 4.6505
R4041 GND.n5024 GND.n5023 4.6505
R4042 GND.n5019 GND.n5018 4.6505
R4043 GND.n5014 GND.n5013 4.6505
R4044 GND.n5009 GND.n5008 4.6505
R4045 GND.n5007 GND.n5006 4.6505
R4046 GND.n5003 GND.n5002 4.6505
R4047 GND.n4999 GND.n4998 4.6505
R4048 GND.n4997 GND.n4996 4.6505
R4049 GND.n4993 GND.n4992 4.6505
R4050 GND.n4991 GND.n4990 4.6505
R4051 GND.n4987 GND.n4986 4.6505
R4052 GND.n4984 GND.n4983 4.6505
R4053 GND.n4975 GND.n4974 4.6505
R4054 GND.n4935 GND.n4934 4.6505
R4055 GND.n4939 GND.n4938 4.6505
R4056 GND.n4941 GND.n4940 4.6505
R4057 GND.n4945 GND.n4944 4.6505
R4058 GND.n5037 GND.n5036 4.6505
R4059 GND.n5035 GND.n5034 4.6505
R4060 GND.n5031 GND.n5030 4.6505
R4061 GND.n4659 GND.n4658 4.6505
R4062 GND.n4684 GND.n4683 4.6505
R4063 GND.n4686 GND.n4685 4.6505
R4064 GND.n4721 GND.n4706 4.6505
R4065 GND.n4720 GND.n4707 4.6505
R4066 GND.n4657 GND.n4656 4.6505
R4067 GND.n4655 GND.n4654 4.6505
R4068 GND.n4651 GND.n4650 4.6505
R4069 GND.n4649 GND.n4648 4.6505
R4070 GND.n4645 GND.n4644 4.6505
R4071 GND.n4643 GND.n4642 4.6505
R4072 GND.n4639 GND.n4638 4.6505
R4073 GND.n4635 GND.n4634 4.6505
R4074 GND.n4612 GND.n4611 4.6505
R4075 GND.n4669 GND.n4668 4.6505
R4076 GND.n4674 GND.n4673 4.6505
R4077 GND.n4676 GND.n4675 4.6505
R4078 GND.n4680 GND.n4679 4.6505
R4079 GND.n4682 GND.n4681 4.6505
R4080 GND.n4688 GND.n4687 4.6505
R4081 GND.n4692 GND.n4691 4.6505
R4082 GND.n4694 GND.n4693 4.6505
R4083 GND.n4698 GND.n4697 4.6505
R4084 GND.n4700 GND.n4699 4.6505
R4085 GND.n4705 GND.n4704 4.6505
R4086 GND.n4746 GND.n4745 4.6505
R4087 GND.n4741 GND.n4740 4.6505
R4088 GND.n4739 GND.n4738 4.6505
R4089 GND.n4735 GND.n4734 4.6505
R4090 GND.n4733 GND.n4732 4.6505
R4091 GND.n4729 GND.n4728 4.6505
R4092 GND.n4727 GND.n4726 4.6505
R4093 GND.n4723 GND.n4722 4.6505
R4094 GND.n4719 GND.n4718 4.6505
R4095 GND.n4717 GND.n4716 4.6505
R4096 GND.n4713 GND.n4712 4.6505
R4097 GND.n4711 GND.n4710 4.6505
R4098 GND.n4608 GND.n4607 4.6505
R4099 GND.n4927 GND.n4926 4.6505
R4100 GND.n4932 GND.n4931 4.6505
R4101 GND.n4661 GND.n4660 4.6505
R4102 GND.n4632 GND.n4631 4.6505
R4103 GND.n4585 GND.n4584 4.6505
R4104 GND.n4588 GND.n4587 4.6505
R4105 GND.n4593 GND.n4592 4.6505
R4106 GND.n4595 GND.n4594 4.6505
R4107 GND.n4599 GND.n4598 4.6505
R4108 GND.n4603 GND.n4602 4.6505
R4109 GND.n4605 GND.n4604 4.6505
R4110 GND.n4616 GND.n4615 4.6505
R4111 GND.n4618 GND.n4617 4.6505
R4112 GND.n4622 GND.n4621 4.6505
R4113 GND.n4624 GND.n4623 4.6505
R4114 GND.n4628 GND.n4627 4.6505
R4115 GND.n5532 GND.n5522 4.6505
R4116 GND.n5531 GND.n5523 4.6505
R4117 GND.n5604 GND.n5603 4.6505
R4118 GND.n5606 GND.n5605 4.6505
R4119 GND.n5780 GND.n5501 4.6505
R4120 GND.n5779 GND.n5502 4.6505
R4121 GND.n5681 GND.n5680 4.6505
R4122 GND.n5683 GND.n5682 4.6505
R4123 GND.n5730 GND.n5729 4.6505
R4124 GND.n5732 GND.n5731 4.6505
R4125 GND.n5742 GND.n5741 4.6505
R4126 GND.n5514 GND.n5513 4.6505
R4127 GND.n5518 GND.n5517 4.6505
R4128 GND.n5521 GND.n5520 4.6505
R4129 GND.n5561 GND.n5560 4.6505
R4130 GND.n5556 GND.n5555 4.6505
R4131 GND.n5552 GND.n5551 4.6505
R4132 GND.n5550 GND.n5549 4.6505
R4133 GND.n5546 GND.n5545 4.6505
R4134 GND.n5544 GND.n5543 4.6505
R4135 GND.n5540 GND.n5539 4.6505
R4136 GND.n5538 GND.n5537 4.6505
R4137 GND.n5534 GND.n5533 4.6505
R4138 GND.n5530 GND.n5529 4.6505
R4139 GND.n5528 GND.n5527 4.6505
R4140 GND.n5508 GND.n5507 4.6505
R4141 GND.n5571 GND.n5570 4.6505
R4142 GND.n5574 GND.n5573 4.6505
R4143 GND.n5578 GND.n5577 4.6505
R4144 GND.n5582 GND.n5581 4.6505
R4145 GND.n5584 GND.n5583 4.6505
R4146 GND.n5588 GND.n5587 4.6505
R4147 GND.n5590 GND.n5589 4.6505
R4148 GND.n5594 GND.n5593 4.6505
R4149 GND.n5596 GND.n5595 4.6505
R4150 GND.n5600 GND.n5599 4.6505
R4151 GND.n5602 GND.n5601 4.6505
R4152 GND.n5608 GND.n5607 4.6505
R4153 GND.n5612 GND.n5611 4.6505
R4154 GND.n5614 GND.n5613 4.6505
R4155 GND.n5619 GND.n5618 4.6505
R4156 GND.n5644 GND.n5643 4.6505
R4157 GND.n5641 GND.n5640 4.6505
R4158 GND.n5637 GND.n5636 4.6505
R4159 GND.n5633 GND.n5632 4.6505
R4160 GND.n5631 GND.n5630 4.6505
R4161 GND.n5627 GND.n5626 4.6505
R4162 GND.n5625 GND.n5624 4.6505
R4163 GND.n5621 GND.n5620 4.6505
R4164 GND.n5500 GND.n5499 4.6505
R4165 GND.n5782 GND.n5781 4.6505
R4166 GND.n5778 GND.n5777 4.6505
R4167 GND.n5776 GND.n5775 4.6505
R4168 GND.n5771 GND.n5770 4.6505
R4169 GND.n5506 GND.n5505 4.6505
R4170 GND.n5651 GND.n5650 4.6505
R4171 GND.n5655 GND.n5654 4.6505
R4172 GND.n5659 GND.n5658 4.6505
R4173 GND.n5661 GND.n5660 4.6505
R4174 GND.n5665 GND.n5664 4.6505
R4175 GND.n5667 GND.n5666 4.6505
R4176 GND.n5671 GND.n5670 4.6505
R4177 GND.n5673 GND.n5672 4.6505
R4178 GND.n5677 GND.n5676 4.6505
R4179 GND.n5679 GND.n5678 4.6505
R4180 GND.n5685 GND.n5684 4.6505
R4181 GND.n5690 GND.n5689 4.6505
R4182 GND.n5693 GND.n5692 4.6505
R4183 GND.n5698 GND.n5697 4.6505
R4184 GND.n5700 GND.n5699 4.6505
R4185 GND.n5704 GND.n5703 4.6505
R4186 GND.n5708 GND.n5707 4.6505
R4187 GND.n5710 GND.n5709 4.6505
R4188 GND.n5714 GND.n5713 4.6505
R4189 GND.n5716 GND.n5715 4.6505
R4190 GND.n5720 GND.n5719 4.6505
R4191 GND.n5722 GND.n5721 4.6505
R4192 GND.n5726 GND.n5725 4.6505
R4193 GND.n5728 GND.n5727 4.6505
R4194 GND.n5734 GND.n5733 4.6505
R4195 GND.n5737 GND.n5736 4.6505
R4196 GND.n5739 GND.n5738 4.6505
R4197 GND.n5762 GND.n5761 4.6505
R4198 GND.n5759 GND.n5758 4.6505
R4199 GND.n5757 GND.n5756 4.6505
R4200 GND.n5755 GND.n5754 4.6505
R4201 GND.n5753 GND.n5752 4.6505
R4202 GND.n5751 GND.n5750 4.6505
R4203 GND.n5747 GND.n5746 4.6505
R4204 GND.n6750 GND.n6749 4.6505
R4205 GND.n6748 GND.n6738 4.6505
R4206 GND.n6747 GND.n6746 4.6505
R4207 GND.n6746 GND.n6745 4.6505
R4208 GND.n6744 GND.n6738 4.6505
R4209 GND.n6750 GND.n6737 4.6505
R4210 GND.n6752 GND.n6751 4.6505
R4211 GND.n6775 GND.n6770 4.6505
R4212 GND.n6777 GND.n6776 4.6505
R4213 GND.n6784 GND.n6783 4.6505
R4214 GND.n6785 GND.n6765 4.6505
R4215 GND.n6787 GND.n6786 4.6505
R4216 GND.n6780 GND.n6768 4.6505
R4217 GND.n6783 GND.n6782 4.6505
R4218 GND.n6781 GND.n6765 4.6505
R4219 GND.n6787 GND.n6764 4.6505
R4220 GND.n6789 GND.n6788 4.6505
R4221 GND.n5447 GND.n5446 4.6505
R4222 GND.n5458 GND.n5457 4.6505
R4223 GND.n5454 GND.n5453 4.6505
R4224 GND.n5456 GND.n5455 4.6505
R4225 GND.n5242 GND.n5241 4.6505
R4226 GND.n5233 GND.n5226 4.6505
R4227 GND.n5232 GND.n5231 4.6505
R4228 GND.n5238 GND.n5237 4.6505
R4229 GND.n5236 GND.n5224 4.6505
R4230 GND.n5242 GND.n5223 4.6505
R4231 GND.n5244 GND.n5243 4.6505
R4232 GND.n5194 GND.n5188 4.6505
R4233 GND.n5197 GND.n5187 4.6505
R4234 GND.n5185 GND.n5184 4.6505
R4235 GND.n5211 GND.n5182 4.6505
R4236 GND.n5193 GND.n5192 4.6505
R4237 GND.n5196 GND.n5195 4.6505
R4238 GND.n5199 GND.n5198 4.6505
R4239 GND.n5201 GND.n5200 4.6505
R4240 GND.n5210 GND.n5209 4.6505
R4241 GND.n5212 GND.n5179 4.6505
R4242 GND.n5214 GND.n5213 4.6505
R4243 GND.n5207 GND.n5182 4.6505
R4244 GND.n5209 GND.n5208 4.6505
R4245 GND.n5205 GND.n5179 4.6505
R4246 GND.n5214 GND.n5180 4.6505
R4247 GND.n6813 GND.n6812 4.6505
R4248 GND.n6815 GND.n6814 4.6505
R4249 GND.n6817 GND.n6816 4.6505
R4250 GND.n6819 GND.n6818 4.6505
R4251 GND.n6821 GND.n6820 4.6505
R4252 GND.n6823 GND.n6822 4.6505
R4253 GND.n6825 GND.n6824 4.6505
R4254 GND.n6827 GND.n6826 4.6505
R4255 GND.n6829 GND.n6828 4.6505
R4256 GND.n6831 GND.n6830 4.6505
R4257 GND.n6833 GND.n6832 4.6505
R4258 GND.n6835 GND.n6834 4.6505
R4259 GND.n4389 GND.n4388 4.6505
R4260 GND.n4387 GND.n4377 4.6505
R4261 GND.n4386 GND.n4385 4.6505
R4262 GND.n4385 GND.n4384 4.6505
R4263 GND.n4383 GND.n4377 4.6505
R4264 GND.n4389 GND.n4376 4.6505
R4265 GND.n4391 GND.n4390 4.6505
R4266 GND.n4353 GND.n4348 4.6505
R4267 GND.n4355 GND.n4354 4.6505
R4268 GND.n4362 GND.n4361 4.6505
R4269 GND.n4363 GND.n4343 4.6505
R4270 GND.n4365 GND.n4364 4.6505
R4271 GND.n4358 GND.n4346 4.6505
R4272 GND.n4361 GND.n4360 4.6505
R4273 GND.n4359 GND.n4343 4.6505
R4274 GND.n4365 GND.n4342 4.6505
R4275 GND.n4367 GND.n4366 4.6505
R4276 GND.n6852 GND.n6851 4.6505
R4277 GND.n6863 GND.n6862 4.6505
R4278 GND.n6859 GND.n6858 4.6505
R4279 GND.n6861 GND.n6860 4.6505
R4280 GND.n4334 GND.n4333 4.6505
R4281 GND.n4325 GND.n4318 4.6505
R4282 GND.n4324 GND.n4323 4.6505
R4283 GND.n4330 GND.n4329 4.6505
R4284 GND.n4328 GND.n4316 4.6505
R4285 GND.n4334 GND.n4315 4.6505
R4286 GND.n4336 GND.n4335 4.6505
R4287 GND.n4291 GND.n4285 4.6505
R4288 GND.n4294 GND.n4284 4.6505
R4289 GND.n4282 GND.n4281 4.6505
R4290 GND.n4308 GND.n4279 4.6505
R4291 GND.n4290 GND.n4289 4.6505
R4292 GND.n4293 GND.n4292 4.6505
R4293 GND.n4296 GND.n4295 4.6505
R4294 GND.n4298 GND.n4297 4.6505
R4295 GND.n4307 GND.n4306 4.6505
R4296 GND.n4309 GND.n4276 4.6505
R4297 GND.n4311 GND.n4310 4.6505
R4298 GND.n4304 GND.n4279 4.6505
R4299 GND.n4306 GND.n4305 4.6505
R4300 GND.n4302 GND.n4276 4.6505
R4301 GND.n4311 GND.n4277 4.6505
R4302 GND.n7058 GND.n7057 4.6505
R4303 GND.n7060 GND.n7059 4.6505
R4304 GND.n7062 GND.n7061 4.6505
R4305 GND.n7064 GND.n7063 4.6505
R4306 GND.n7066 GND.n7065 4.6505
R4307 GND.n7068 GND.n7067 4.6505
R4308 GND.n7070 GND.n7069 4.6505
R4309 GND.n7072 GND.n7071 4.6505
R4310 GND.n7074 GND.n7073 4.6505
R4311 GND.n7076 GND.n7075 4.6505
R4312 GND.n7078 GND.n7077 4.6505
R4313 GND.n7080 GND.n7079 4.6505
R4314 GND.n4480 GND.n4479 4.6505
R4315 GND.n4482 GND.n4481 4.6505
R4316 GND.n4504 GND.n4492 4.6505
R4317 GND.n4503 GND.n4493 4.6505
R4318 GND.n5044 GND.n5043 4.6505
R4319 GND.n5046 GND.n5045 4.6505
R4320 GND.n5061 GND.n5056 4.6505
R4321 GND.n5060 GND.n5057 4.6505
R4322 GND.n5141 GND.n5140 4.6505
R4323 GND.n5143 GND.n5142 4.6505
R4324 GND.n5153 GND.n5152 4.6505
R4325 GND.n4439 GND.n4438 4.6505
R4326 GND.n4443 GND.n4442 4.6505
R4327 GND.n4445 GND.n4444 4.6505
R4328 GND.n4453 GND.n4452 4.6505
R4329 GND.n4458 GND.n4457 4.6505
R4330 GND.n4460 GND.n4459 4.6505
R4331 GND.n4464 GND.n4463 4.6505
R4332 GND.n4466 GND.n4465 4.6505
R4333 GND.n4470 GND.n4469 4.6505
R4334 GND.n4472 GND.n4471 4.6505
R4335 GND.n4476 GND.n4475 4.6505
R4336 GND.n4478 GND.n4477 4.6505
R4337 GND.n4484 GND.n4483 4.6505
R4338 GND.n4488 GND.n4487 4.6505
R4339 GND.n4491 GND.n4490 4.6505
R4340 GND.n4539 GND.n4538 4.6505
R4341 GND.n4534 GND.n4533 4.6505
R4342 GND.n4532 GND.n4531 4.6505
R4343 GND.n4528 GND.n4527 4.6505
R4344 GND.n4524 GND.n4523 4.6505
R4345 GND.n4522 GND.n4521 4.6505
R4346 GND.n4518 GND.n4517 4.6505
R4347 GND.n4516 GND.n4515 4.6505
R4348 GND.n4512 GND.n4511 4.6505
R4349 GND.n4510 GND.n4509 4.6505
R4350 GND.n4506 GND.n4505 4.6505
R4351 GND.n4502 GND.n4501 4.6505
R4352 GND.n4500 GND.n4499 4.6505
R4353 GND.n4496 GND.n4495 4.6505
R4354 GND.n4434 GND.n4433 4.6505
R4355 GND.n4547 GND.n4546 4.6505
R4356 GND.n4552 GND.n4551 4.6505
R4357 GND.n4556 GND.n4555 4.6505
R4358 GND.n4558 GND.n4557 4.6505
R4359 GND.n4562 GND.n4561 4.6505
R4360 GND.n4564 GND.n4563 4.6505
R4361 GND.n4568 GND.n4567 4.6505
R4362 GND.n4570 GND.n4569 4.6505
R4363 GND.n4574 GND.n4573 4.6505
R4364 GND.n4576 GND.n4575 4.6505
R4365 GND.n5048 GND.n5047 4.6505
R4366 GND.n5052 GND.n5051 4.6505
R4367 GND.n5055 GND.n5054 4.6505
R4368 GND.n5096 GND.n5095 4.6505
R4369 GND.n5091 GND.n5090 4.6505
R4370 GND.n5089 GND.n5088 4.6505
R4371 GND.n5085 GND.n5084 4.6505
R4372 GND.n5081 GND.n5080 4.6505
R4373 GND.n5079 GND.n5078 4.6505
R4374 GND.n5075 GND.n5074 4.6505
R4375 GND.n5073 GND.n5072 4.6505
R4376 GND.n5069 GND.n5068 4.6505
R4377 GND.n5067 GND.n5066 4.6505
R4378 GND.n5063 GND.n5062 4.6505
R4379 GND.n5059 GND.n5058 4.6505
R4380 GND.n4430 GND.n4429 4.6505
R4381 GND.n5104 GND.n5103 4.6505
R4382 GND.n5109 GND.n5108 4.6505
R4383 GND.n5111 GND.n5110 4.6505
R4384 GND.n5115 GND.n5114 4.6505
R4385 GND.n5119 GND.n5118 4.6505
R4386 GND.n5121 GND.n5120 4.6505
R4387 GND.n5125 GND.n5124 4.6505
R4388 GND.n5127 GND.n5126 4.6505
R4389 GND.n5131 GND.n5130 4.6505
R4390 GND.n5133 GND.n5132 4.6505
R4391 GND.n5137 GND.n5136 4.6505
R4392 GND.n5139 GND.n5138 4.6505
R4393 GND.n5145 GND.n5144 4.6505
R4394 GND.n5148 GND.n5147 4.6505
R4395 GND.n5150 GND.n5149 4.6505
R4396 GND.n5173 GND.n5172 4.6505
R4397 GND.n5170 GND.n5169 4.6505
R4398 GND.n5168 GND.n5167 4.6505
R4399 GND.n5166 GND.n5165 4.6505
R4400 GND.n5164 GND.n5163 4.6505
R4401 GND.n5162 GND.n5161 4.6505
R4402 GND.n5158 GND.n5157 4.6505
R4403 GND.n6440 GND.n6430 4.6505
R4404 GND.n6439 GND.n6431 4.6505
R4405 GND.n6512 GND.n6511 4.6505
R4406 GND.n6514 GND.n6513 4.6505
R4407 GND.n6602 GND.n6601 4.6505
R4408 GND.n6604 GND.n6603 4.6505
R4409 GND.n6619 GND.n6614 4.6505
R4410 GND.n6618 GND.n6615 4.6505
R4411 GND.n6699 GND.n6698 4.6505
R4412 GND.n6701 GND.n6700 4.6505
R4413 GND.n6711 GND.n6710 4.6505
R4414 GND.n6423 GND.n6422 4.6505
R4415 GND.n6427 GND.n6426 4.6505
R4416 GND.n6429 GND.n6428 4.6505
R4417 GND.n6469 GND.n6468 4.6505
R4418 GND.n6464 GND.n6463 4.6505
R4419 GND.n6460 GND.n6459 4.6505
R4420 GND.n6458 GND.n6457 4.6505
R4421 GND.n6454 GND.n6453 4.6505
R4422 GND.n6452 GND.n6451 4.6505
R4423 GND.n6448 GND.n6447 4.6505
R4424 GND.n6446 GND.n6445 4.6505
R4425 GND.n6442 GND.n6441 4.6505
R4426 GND.n6438 GND.n6437 4.6505
R4427 GND.n6436 GND.n6435 4.6505
R4428 GND.n6418 GND.n6417 4.6505
R4429 GND.n6479 GND.n6478 4.6505
R4430 GND.n6482 GND.n6481 4.6505
R4431 GND.n6486 GND.n6485 4.6505
R4432 GND.n6490 GND.n6489 4.6505
R4433 GND.n6492 GND.n6491 4.6505
R4434 GND.n6496 GND.n6495 4.6505
R4435 GND.n6498 GND.n6497 4.6505
R4436 GND.n6502 GND.n6501 4.6505
R4437 GND.n6504 GND.n6503 4.6505
R4438 GND.n6508 GND.n6507 4.6505
R4439 GND.n6510 GND.n6509 4.6505
R4440 GND.n6516 GND.n6515 4.6505
R4441 GND.n6520 GND.n6519 4.6505
R4442 GND.n6522 GND.n6521 4.6505
R4443 GND.n6527 GND.n6526 4.6505
R4444 GND.n6556 GND.n6555 4.6505
R4445 GND.n6553 GND.n6552 4.6505
R4446 GND.n6549 GND.n6548 4.6505
R4447 GND.n6545 GND.n6544 4.6505
R4448 GND.n6543 GND.n6542 4.6505
R4449 GND.n6539 GND.n6538 4.6505
R4450 GND.n6537 GND.n6536 4.6505
R4451 GND.n6533 GND.n6532 4.6505
R4452 GND.n6531 GND.n6530 4.6505
R4453 GND.n5496 GND.n5495 4.6505
R4454 GND.n6606 GND.n6605 4.6505
R4455 GND.n6610 GND.n6609 4.6505
R4456 GND.n6613 GND.n6612 4.6505
R4457 GND.n6654 GND.n6653 4.6505
R4458 GND.n6649 GND.n6648 4.6505
R4459 GND.n6647 GND.n6646 4.6505
R4460 GND.n6643 GND.n6642 4.6505
R4461 GND.n6639 GND.n6638 4.6505
R4462 GND.n6637 GND.n6636 4.6505
R4463 GND.n6633 GND.n6632 4.6505
R4464 GND.n6631 GND.n6630 4.6505
R4465 GND.n6627 GND.n6626 4.6505
R4466 GND.n6625 GND.n6624 4.6505
R4467 GND.n6621 GND.n6620 4.6505
R4468 GND.n6617 GND.n6616 4.6505
R4469 GND.n5494 GND.n5493 4.6505
R4470 GND.n6662 GND.n6661 4.6505
R4471 GND.n6667 GND.n6666 4.6505
R4472 GND.n6669 GND.n6668 4.6505
R4473 GND.n6673 GND.n6672 4.6505
R4474 GND.n6677 GND.n6676 4.6505
R4475 GND.n6679 GND.n6678 4.6505
R4476 GND.n6683 GND.n6682 4.6505
R4477 GND.n6685 GND.n6684 4.6505
R4478 GND.n6689 GND.n6688 4.6505
R4479 GND.n6691 GND.n6690 4.6505
R4480 GND.n6695 GND.n6694 4.6505
R4481 GND.n6697 GND.n6696 4.6505
R4482 GND.n6703 GND.n6702 4.6505
R4483 GND.n6706 GND.n6705 4.6505
R4484 GND.n6708 GND.n6707 4.6505
R4485 GND.n6731 GND.n6730 4.6505
R4486 GND.n6728 GND.n6727 4.6505
R4487 GND.n6726 GND.n6725 4.6505
R4488 GND.n6724 GND.n6723 4.6505
R4489 GND.n6722 GND.n6721 4.6505
R4490 GND.n6720 GND.n6719 4.6505
R4491 GND.n6716 GND.n6715 4.6505
R4492 GND.n4074 GND.n4073 4.52281
R4493 GND.n1044 GND.n898 4.52235
R4494 GND.n1935 GND.n1934 4.5005
R4495 GND.n1928 GND.n1921 4.5005
R4496 GND.n1900 GND.n1899 4.5005
R4497 GND.n1913 GND.n1907 4.5005
R4498 GND.n1702 GND.n1701 4.5005
R4499 GND.n1695 GND.n1688 4.5005
R4500 GND.n1857 GND.n1856 4.5005
R4501 GND.n1870 GND.n1864 4.5005
R4502 GND.n6910 GND.n6909 4.5005
R4503 GND.n6903 GND.n6896 4.5005
R4504 GND.n7037 GND.n6881 4.5005
R4505 GND.n6891 GND.n6885 4.5005
R4506 GND.n2378 GND.n2377 4.5005
R4507 GND.n2371 GND.n2364 4.5005
R4508 GND.n2506 GND.n2505 4.5005
R4509 GND.n2519 GND.n2513 4.5005
R4510 GND.n2703 GND.n2702 4.5005
R4511 GND.n2696 GND.n2689 4.5005
R4512 GND.n2831 GND.n2830 4.5005
R4513 GND.n2844 GND.n2838 4.5005
R4514 GND.n3027 GND.n3026 4.5005
R4515 GND.n3020 GND.n3013 4.5005
R4516 GND.n3128 GND.n3127 4.5005
R4517 GND.n3141 GND.n3135 4.5005
R4518 GND.n7100 GND.n7099 4.5005
R4519 GND.n7093 GND.n7086 4.5005
R4520 GND.n7228 GND.n7227 4.5005
R4521 GND.n7241 GND.n7235 4.5005
R4522 GND.n4795 GND.n4794 4.5005
R4523 GND.n4788 GND.n4781 4.5005
R4524 GND.n4760 GND.n4759 4.5005
R4525 GND.n4773 GND.n4767 4.5005
R4526 GND.n5277 GND.n5276 4.5005
R4527 GND.n5270 GND.n5263 4.5005
R4528 GND.n5429 GND.n5248 4.5005
R4529 GND.n5258 GND.n5252 4.5005
R4530 GND.n5799 GND.n5798 4.5005
R4531 GND.n5792 GND.n5785 4.5005
R4532 GND.n5928 GND.n5927 4.5005
R4533 GND.n5941 GND.n5935 4.5005
R4534 GND.n5966 GND.n5965 4.5005
R4535 GND.n5959 GND.n5952 4.5005
R4536 GND.n6097 GND.n6096 4.5005
R4537 GND.n6110 GND.n6104 4.5005
R4538 GND.n6133 GND.n6132 4.5005
R4539 GND.n6126 GND.n6119 4.5005
R4540 GND.n6261 GND.n6260 4.5005
R4541 GND.n6274 GND.n6268 4.5005
R4542 GND.n6297 GND.n6296 4.5005
R4543 GND.n6290 GND.n6283 4.5005
R4544 GND.n6570 GND.n6569 4.5005
R4545 GND.n6583 GND.n6577 4.5005
R4546 GND.n585 GND.n584 4.5005
R4547 GND.n578 GND.n571 4.5005
R4548 GND.n710 GND.n709 4.5005
R4549 GND.n723 GND.n717 4.5005
R4550 GND.n7628 GND.n7627 4.5005
R4551 GND.n7621 GND.n7614 4.5005
R4552 GND.n7757 GND.n7756 4.5005
R4553 GND.n7770 GND.n7764 4.5005
R4554 GND.n3855 GND.n3658 4.5005
R4555 GND.n3855 GND.n3854 4.5005
R4556 GND.n7508 GND.n7507 4.5005
R4557 GND.n7501 GND.n7494 4.5005
R4558 GND.n7592 GND.n7591 4.5005
R4559 GND.n7605 GND.n7599 4.5005
R4560 GND.n4049 GND.n4048 4.4805
R4561 GND.n4037 GND.n4036 4.4805
R4562 GND.n6421 GND.n6420 4.45136
R4563 GND.n5512 GND.n5511 4.45136
R4564 GND.n4437 GND.n4436 4.45136
R4565 GND.n1145 GND.t791 4.41708
R4566 GND.n7352 GND.t529 4.41708
R4567 GND.n2087 GND.t790 4.41708
R4568 GND.n1129 GND.t472 4.41708
R4569 GND.n1137 GND.t388 4.41708
R4570 GND.n1121 GND.t37 4.41708
R4571 GND.n1113 GND.t1248 4.41708
R4572 GND.n7314 GND.t1126 4.41708
R4573 GND.n4172 GND.t40 4.41708
R4574 GND.n3366 GND.t531 4.41708
R4575 GND.n3209 GND.t792 4.41708
R4576 GND.n2912 GND.t1125 4.41708
R4577 GND.n2587 GND.t473 4.41708
R4578 GND.n2263 GND.t530 4.41708
R4579 GND.n7342 GND.t1249 4.41708
R4580 GND.n2097 GND.t1251 4.41708
R4581 GND.n789 GND.t38 4.35136
R4582 GND.n7353 GND.t41 4.35136
R4583 GND.n2085 GND.t1252 4.35136
R4584 GND.n317 GND.t1127 4.35136
R4585 GND.n470 GND.t794 4.35136
R4586 GND.n165 GND.t386 4.35136
R4587 GND.n56 GND.t532 4.35136
R4588 GND.n7315 GND.t1250 4.35136
R4589 GND.n4173 GND.t389 4.35136
R4590 GND.n3367 GND.t1124 4.35136
R4591 GND.n3210 GND.t39 4.35136
R4592 GND.n2913 GND.t793 4.35136
R4593 GND.n2588 GND.t1128 4.35136
R4594 GND.n2264 GND.t387 4.35136
R4595 GND.n7340 GND.t533 4.35136
R4596 GND.n2098 GND.t385 4.35136
R4597 GND.n4977 GND.n4976 4.25025
R4598 GND.n5489 GND.n5488 4.06709
R4599 GND.n4420 GND.n4419 4.06709
R4600 GND.n6741 GND.n6740 4.06409
R4601 GND.n4380 GND.n4379 4.06409
R4602 GND.n6743 GND.n6741 4.0631
R4603 GND.n4382 GND.n4380 4.0631
R4604 GND.n6778 GND.n6767 4.05611
R4605 GND.n4356 GND.n4345 4.05611
R4606 GND.n5204 GND.n5202 3.98881
R4607 GND.n4301 GND.n4299 3.98881
R4608 GND.n2079 GND.n2078 3.9685
R4609 GND.n411 GND.n410 3.9685
R4610 GND.n837 GND.n836 3.9685
R4611 GND.n4046 GND.n4045 3.84205
R4612 GND.n6774 GND.n6773 3.80559
R4613 GND.n5230 GND.n5228 3.80559
R4614 GND.n4352 GND.n4351 3.80559
R4615 GND.n4322 GND.n4320 3.80559
R4616 GND.n5472 GND.n5470 3.80083
R4617 GND.n4403 GND.n4401 3.80083
R4618 GND.n3839 GND.n3834 3.7002
R4619 GND.n100 GND.n95 3.63686
R4620 GND.n3692 GND.n3659 3.38533
R4621 GND.n3677 GND.n3675 3.20453
R4622 GND.n1939 GND.n1938 3.03311
R4623 GND.n1915 GND.n1905 3.03311
R4624 GND.n1706 GND.n1705 3.03311
R4625 GND.n1872 GND.n1862 3.03311
R4626 GND.n6914 GND.n6913 3.03311
R4627 GND.n6893 GND.n6883 3.03311
R4628 GND.n2382 GND.n2381 3.03311
R4629 GND.n2521 GND.n2511 3.03311
R4630 GND.n2707 GND.n2706 3.03311
R4631 GND.n2846 GND.n2836 3.03311
R4632 GND.n3031 GND.n3030 3.03311
R4633 GND.n3143 GND.n3133 3.03311
R4634 GND.n7104 GND.n7103 3.03311
R4635 GND.n7243 GND.n7233 3.03311
R4636 GND.n4799 GND.n4798 3.03311
R4637 GND.n4775 GND.n4765 3.03311
R4638 GND.n5281 GND.n5280 3.03311
R4639 GND.n5260 GND.n5250 3.03311
R4640 GND.n5803 GND.n5802 3.03311
R4641 GND.n5943 GND.n5933 3.03311
R4642 GND.n5970 GND.n5969 3.03311
R4643 GND.n6112 GND.n6102 3.03311
R4644 GND.n6137 GND.n6136 3.03311
R4645 GND.n6276 GND.n6266 3.03311
R4646 GND.n6301 GND.n6300 3.03311
R4647 GND.n6585 GND.n6575 3.03311
R4648 GND.n589 GND.n588 3.03311
R4649 GND.n725 GND.n715 3.03311
R4650 GND.n7632 GND.n7631 3.03311
R4651 GND.n7772 GND.n7762 3.03311
R4652 GND.n7375 GND.n7374 3.03311
R4653 GND.n7379 GND.n7378 3.03311
R4654 GND.n1371 GND.n1370 3.03311
R4655 GND.n1375 GND.n1374 3.03311
R4656 GND.n328 GND.n327 3.03311
R4657 GND.n337 GND.n336 3.03311
R4658 GND.n481 GND.n480 3.03311
R4659 GND.n490 GND.n489 3.03311
R4660 GND.n176 GND.n175 3.03311
R4661 GND.n185 GND.n184 3.03311
R4662 GND.n1485 GND.n1484 3.03311
R4663 GND.n1520 GND.n1519 3.03311
R4664 GND.n1384 GND.n1383 3.03311
R4665 GND.n1472 GND.n1471 3.03311
R4666 GND.n4184 GND.n4183 3.03311
R4667 GND.n4193 GND.n4192 3.03311
R4668 GND.n3378 GND.n3377 3.03311
R4669 GND.n3387 GND.n3386 3.03311
R4670 GND.n3221 GND.n3220 3.03311
R4671 GND.n3230 GND.n3229 3.03311
R4672 GND.n2924 GND.n2923 3.03311
R4673 GND.n2933 GND.n2932 3.03311
R4674 GND.n2599 GND.n2598 3.03311
R4675 GND.n2608 GND.n2607 3.03311
R4676 GND.n2275 GND.n2274 3.03311
R4677 GND.n2284 GND.n2283 3.03311
R4678 GND.n2113 GND.n2112 3.03311
R4679 GND.n2122 GND.n2121 3.03311
R4680 GND.n1245 GND.n1244 3.03311
R4681 GND.n1254 GND.n1253 3.03311
R4682 GND.n7393 GND.n7392 3.03311
R4683 GND.n7421 GND.n7420 3.03311
R4684 GND.n7512 GND.n7511 3.03311
R4685 GND.n7607 GND.n7597 3.03311
R4686 GND.n7362 GND 3.0005
R4687 GND.n2015 GND 3.0005
R4688 GND.n513 GND 3.0005
R4689 GND.n208 GND 3.0005
R4690 GND.n1507 GND 3.0005
R4691 GND.n1459 GND 3.0005
R4692 GND.n4216 GND 3.0005
R4693 GND.n3410 GND 3.0005
R4694 GND.n3253 GND 3.0005
R4695 GND.n2956 GND 3.0005
R4696 GND.n2631 GND 3.0005
R4697 GND.n2307 GND 3.0005
R4698 GND.n2145 GND 3.0005
R4699 GND.n1277 GND 3.0005
R4700 GND.n360 GND 3.0005
R4701 GND.n7408 GND 3.0005
R4702 GND.n5767 GND.t1497 2.84655
R4703 GND.n2136 GND.n2135 2.5872
R4704 GND.n2622 GND.n2621 2.5872
R4705 GND.n3244 GND.n3243 2.5872
R4706 GND.n4207 GND.n4206 2.5872
R4707 GND.n199 GND.n198 2.5872
R4708 GND.n504 GND.n503 2.5872
R4709 GND.n1268 GND.n1267 2.56838
R4710 GND.n2298 GND.n2297 2.56838
R4711 GND.n2947 GND.n2946 2.56838
R4712 GND.n3401 GND.n3400 2.56838
R4713 GND.n1450 GND.n1449 2.56838
R4714 GND.n1498 GND.n1497 2.56838
R4715 GND.n2006 GND.n2005 2.56838
R4716 GND.n351 GND.n350 2.56838
R4717 GND.n7399 GND.n7398 2.56838
R4718 GND.n3642 GND.t1271 2.36824
R4719 GND.n3639 GND.t393 2.36824
R4720 GND.n6719 GND.n6718 2.25932
R4721 GND.n5750 GND.n5749 2.25932
R4722 GND.n5161 GND.n5160 2.25932
R4723 GND.n1211 GND.n1210 1.93119
R4724 GND.n1210 GND.n1209 1.93119
R4725 GND.n2236 GND.n2235 1.93119
R4726 GND.n2235 GND.n2234 1.93119
R4727 GND.n2560 GND.n2559 1.93119
R4728 GND.n2559 GND.n2558 1.93119
R4729 GND.n2885 GND.n2884 1.93119
R4730 GND.n2884 GND.n2883 1.93119
R4731 GND.n3182 GND.n3181 1.93119
R4732 GND.n3181 GND.n3180 1.93119
R4733 GND.n3339 GND.n3338 1.93119
R4734 GND.n3338 GND.n3337 1.93119
R4735 GND.n3497 GND.n3496 1.93119
R4736 GND.n3496 GND.n3495 1.93119
R4737 GND.n7287 GND.n7286 1.93119
R4738 GND.n7286 GND.n7285 1.93119
R4739 GND.n31 GND.n30 1.93119
R4740 GND.n30 GND.n29 1.93119
R4741 GND.n140 GND.n139 1.93119
R4742 GND.n139 GND.n138 1.93119
R4743 GND.n292 GND.n291 1.93119
R4744 GND.n291 GND.n290 1.93119
R4745 GND.n1655 GND.n1654 1.93119
R4746 GND.n1654 GND.n1653 1.93119
R4747 GND.n445 GND.n444 1.93119
R4748 GND.n444 GND.n443 1.93119
R4749 GND.n764 GND.n763 1.93119
R4750 GND.n763 GND.n762 1.93119
R4751 GND.n871 GND.n870 1.93119
R4752 GND.n870 GND.n869 1.93119
R4753 GND.n7808 GND.n7807 1.93119
R4754 GND.n7807 GND.n7806 1.93119
R4755 GND.n3677 GND.n3676 1.85757
R4756 GND.n95 GND.n92 1.81868
R4757 GND.n3636 GND.n3635 1.70717
R4758 GND.n7490 GND.n7489 1.64041
R4759 GND.n567 GND.n566 1.64041
R4760 GND.n258 GND.n257 1.64041
R4761 GND.n106 GND.n105 1.64041
R4762 GND.n1439 GND.n1438 1.64041
R4763 GND.n4266 GND.n4265 1.64041
R4764 GND.n3463 GND.n3462 1.64041
R4765 GND.n3305 GND.n3304 1.64041
R4766 GND.n3009 GND.n3008 1.64041
R4767 GND.n2685 GND.n2684 1.64041
R4768 GND.n2360 GND.n2359 1.64041
R4769 GND.n2202 GND.n2201 1.64041
R4770 GND.n1321 GND.n1320 1.64041
R4771 GND.n1438 GND.n1437 1.63319
R4772 GND.n3462 GND.n3461 1.63319
R4773 GND.n3008 GND.n3007 1.63319
R4774 GND.n2359 GND.n2358 1.63319
R4775 GND.n1320 GND.n1319 1.63319
R4776 GND.n2201 GND.n2200 1.63319
R4777 GND.n2684 GND.n2683 1.63319
R4778 GND.n3304 GND.n3303 1.63319
R4779 GND.n4265 GND.n4264 1.63319
R4780 GND.n105 GND.n104 1.63319
R4781 GND.n257 GND.n256 1.63319
R4782 GND.n566 GND.n565 1.63319
R4783 GND.n7489 GND.n7488 1.63319
R4784 GND.n3861 GND.n3860 1.49383
R4785 GND.n3691 GND.n3689 1.40675
R4786 GND.n3687 GND.n3666 1.40675
R4787 GND.n3674 GND.n3672 1.3822
R4788 GND.n3680 GND.n3679 1.3822
R4789 GND.n4065 GND.n4064 1.2805
R4790 GND.n4056 GND.n4055 1.2805
R4791 GND.n7823 GND.n7781 1.22123
R4792 GND.n7780 GND.n895 1.20741
R4793 GND.n788 GND.n733 1.20741
R4794 GND.n1881 GND.n1687 1.20741
R4795 GND.n5951 GND.n55 1.20741
R4796 GND.n7311 GND.n7256 1.20741
R4797 GND.n3206 GND.n3151 1.20741
R4798 GND.n2909 GND.n2854 1.20741
R4799 GND.n2584 GND.n2529 1.20741
R4800 GND.n7026 GND.n2260 1.20741
R4801 GND.n1879 GND.n1235 1.20741
R4802 GND.n6694 GND.n6693 1.12991
R4803 GND.n6624 GND.n6623 1.12991
R4804 GND.n6530 GND.n6529 1.12991
R4805 GND.n6507 GND.n6506 1.12991
R4806 GND.n6445 GND.n6444 1.12991
R4807 GND.n1907 GND.n1906 1.12991
R4808 GND.n1864 GND.n1863 1.12991
R4809 GND.n6885 GND.n6884 1.12991
R4810 GND.n2513 GND.n2512 1.12991
R4811 GND.n2838 GND.n2837 1.12991
R4812 GND.n3135 GND.n3134 1.12991
R4813 GND.n7235 GND.n7234 1.12991
R4814 GND.n4767 GND.n4766 1.12991
R4815 GND.n5252 GND.n5251 1.12991
R4816 GND.n5935 GND.n5934 1.12991
R4817 GND.n6104 GND.n6103 1.12991
R4818 GND.n6268 GND.n6267 1.12991
R4819 GND.n6577 GND.n6576 1.12991
R4820 GND.n717 GND.n716 1.12991
R4821 GND.n7764 GND.n7763 1.12991
R4822 GND.n7599 GND.n7598 1.12991
R4823 GND.n4679 GND.n4678 1.12991
R4824 GND.n4726 GND.n4725 1.12991
R4825 GND.n5034 GND.n5033 1.12991
R4826 GND.n4983 GND.n4982 1.12991
R4827 GND.n4627 GND.n4626 1.12991
R4828 GND.n5725 GND.n5724 1.12991
R4829 GND.n5676 GND.n5675 1.12991
R4830 GND.n5499 GND.n5498 1.12991
R4831 GND.n5599 GND.n5598 1.12991
R4832 GND.n5537 GND.n5536 1.12991
R4833 GND.n5136 GND.n5135 1.12991
R4834 GND.n5066 GND.n5065 1.12991
R4835 GND.n4573 GND.n4572 1.12991
R4836 GND.n4509 GND.n4508 1.12991
R4837 GND.n4475 GND.n4474 1.12991
R4838 GND.n7492 GND.n7491 1.10116
R4839 GND.n2081 GND.n2080 1.10116
R4840 GND.n569 GND.n568 1.10116
R4841 GND.n260 GND.n259 1.10116
R4842 GND.n108 GND.n107 1.10116
R4843 GND.n1441 GND.n1440 1.10116
R4844 GND.n4268 GND.n4267 1.10116
R4845 GND.n3465 GND.n3464 1.10116
R4846 GND.n3307 GND.n3306 1.10116
R4847 GND.n3011 GND.n3010 1.10116
R4848 GND.n2687 GND.n2686 1.10116
R4849 GND.n2362 GND.n2361 1.10116
R4850 GND.n2204 GND.n2203 1.10116
R4851 GND.n1323 GND.n1322 1.10116
R4852 GND.n413 GND.n412 1.10116
R4853 GND.n839 GND.n838 1.10116
R4854 GND.n7465 GND.n7464 0.9605
R4855 GND.n7469 GND.n7468 0.9605
R4856 GND.n2063 GND.n2055 0.9605
R4857 GND.n391 GND.n390 0.9605
R4858 GND.n545 GND.n544 0.9605
R4859 GND.n550 GND.n549 0.9605
R4860 GND.n240 GND.n239 0.9605
R4861 GND.n76 GND.n75 0.9605
R4862 GND.n80 GND.n79 0.9605
R4863 GND.n1414 GND.n1413 0.9605
R4864 GND.n1422 GND.n1421 0.9605
R4865 GND.n4249 GND.n4248 0.9605
R4866 GND.n3441 GND.n3440 0.9605
R4867 GND.n3446 GND.n3445 0.9605
R4868 GND.n3284 GND.n3283 0.9605
R4869 GND.n3288 GND.n3287 0.9605
R4870 GND.n2988 GND.n2987 0.9605
R4871 GND.n2992 GND.n2991 0.9605
R4872 GND.n2663 GND.n2662 0.9605
R4873 GND.n2668 GND.n2667 0.9605
R4874 GND.n2338 GND.n2337 0.9605
R4875 GND.n2343 GND.n2342 0.9605
R4876 GND.n2176 GND.n2175 0.9605
R4877 GND.n2185 GND.n2184 0.9605
R4878 GND.n2180 GND.n2179 0.9605
R4879 GND.n1673 GND.n1672 0.9605
R4880 GND.n395 GND.n394 0.9605
R4881 GND.n817 GND.n816 0.9605
R4882 GND.n821 GND.n820 0.9605
R4883 GND.n7661 GND.n7660 0.932703
R4884 GND.n7701 GND.t1141 0.932703
R4885 GND.n617 GND.n616 0.932703
R4886 GND.n654 GND.t1232 0.932703
R4887 GND.n6329 GND.n6328 0.932703
R4888 GND.n6366 GND.t1183 0.932703
R4889 GND.n6165 GND.n6164 0.932703
R4890 GND.n6202 GND.t1115 0.932703
R4891 GND.n5998 GND.n5997 0.932703
R4892 GND.n6038 GND.t18 0.932703
R4893 GND.n5815 GND.n5814 0.932703
R4894 GND.n5855 GND.t744 0.932703
R4895 GND.n5293 GND.n5292 0.932703
R4896 GND.n5333 GND.t478 0.932703
R4897 GND.n4852 GND.n4851 0.932703
R4898 GND.n4892 GND.t1309 0.932703
R4899 GND.n7159 GND.n7158 0.932703
R4900 GND.n7199 GND.t521 0.932703
R4901 GND.n3059 GND.n3058 0.932703
R4902 GND.n3099 GND.t828 0.932703
R4903 GND.n2735 GND.n2734 0.932703
R4904 GND.n2775 GND.t142 0.932703
R4905 GND.n2410 GND.n2409 0.932703
R4906 GND.n2450 GND.t815 0.932703
R4907 GND.n6926 GND.n6925 0.932703
R4908 GND.n6966 GND.t804 0.932703
R4909 GND.n1761 GND.n1760 0.932703
R4910 GND.n1801 GND.t774 0.932703
R4911 GND.n1570 GND.n1569 0.932703
R4912 GND.n1610 GND.t1344 0.932703
R4913 GND.n2092 GND.n2091 0.795683
R4914 GND.n7347 GND.n7346 0.795683
R4915 GND.n2091 GND.n2090 0.795337
R4916 GND.n1363 GND.n1362 0.795337
R4917 GND.n2093 GND.n1363 0.795337
R4918 GND.n7346 GND.n7345 0.795337
R4919 GND.n1180 GND.n1179 0.795337
R4920 GND.n7348 GND.n1180 0.795337
R4921 GND.n1178 GND.n1177 0.795337
R4922 GND.n7348 GND.n1178 0.795337
R4923 GND.n1176 GND.n1175 0.795337
R4924 GND.n7348 GND.n1176 0.795337
R4925 GND.n1174 GND.n1173 0.795337
R4926 GND.n7348 GND.n1174 0.795337
R4927 GND.n1172 GND.n1171 0.795337
R4928 GND.n7348 GND.n1172 0.795337
R4929 GND.n1170 GND.n1169 0.795337
R4930 GND.n7348 GND.n1170 0.795337
R4931 GND.n1168 GND.n1167 0.795337
R4932 GND.n7348 GND.n1168 0.795337
R4933 GND.n1166 GND.n1165 0.795337
R4934 GND.n7348 GND.n1166 0.795337
R4935 GND.n1164 GND.n1163 0.795337
R4936 GND.n7348 GND.n1164 0.795337
R4937 GND.n1162 GND.n1161 0.795337
R4938 GND.n7348 GND.n1162 0.795337
R4939 GND.n1160 GND.n1159 0.795337
R4940 GND.n7348 GND.n1160 0.795337
R4941 GND.n1156 GND.n1155 0.795337
R4942 GND.n7348 GND.n1156 0.795337
R4943 GND.n1158 GND.n1157 0.795337
R4944 GND.n7348 GND.n1158 0.795337
R4945 GND.n4581 GND.n4580 0.705542
R4946 GND.n3628 GND.n3626 0.6255
R4947 GND.n1882 GND 0.589529
R4948 GND.n3661 GND.n3660 0.549071
R4949 GND.n3647 GND.n3646 0.54612
R4950 GND.n1886 GND.n1624 0.533636
R4951 GND.n1843 GND.n1842 0.533636
R4952 GND.n7011 GND.n7010 0.533636
R4953 GND.n2492 GND.n2491 0.533636
R4954 GND.n2817 GND.n2816 0.533636
R4955 GND.n3114 GND.n3113 0.533636
R4956 GND.n7214 GND.n7213 0.533636
R4957 GND.n4907 GND.n4906 0.533636
R4958 GND.n5379 GND.n5378 0.533636
R4959 GND.n5901 GND.n5900 0.533636
R4960 GND.n6083 GND.n6082 0.533636
R4961 GND.n6247 GND.n6246 0.533636
R4962 GND.n6411 GND.n6410 0.533636
R4963 GND.n696 GND.n695 0.533636
R4964 GND.n7743 GND.n7742 0.533636
R4965 GND.n7579 GND.n7578 0.533636
R4966 GND.n5039 GND.n4606 0.53211
R4967 GND.n7824 GND.n7493 0.520438
R4968 GND.n2083 GND.n2082 0.520438
R4969 GND.n7830 GND.n570 0.520438
R4970 GND.n7836 GND.n261 0.520438
R4971 GND.n7839 GND.n109 0.520438
R4972 GND.n1442 GND.n0 0.520438
R4973 GND.n7319 GND.n4269 0.520438
R4974 GND.n7323 GND.n3466 0.520438
R4975 GND.n7326 GND.n3308 0.520438
R4976 GND.n7329 GND.n3012 0.520438
R4977 GND.n7332 GND.n2688 0.520438
R4978 GND.n7335 GND.n2363 0.520438
R4979 GND.n7338 GND.n2205 0.520438
R4980 GND.n2101 GND.n1324 0.520438
R4981 GND.n7833 GND.n414 0.520438
R4982 GND.n7827 GND.n840 0.520438
R4983 GND.n5042 GND.n5041 0.48654
R4984 GND.n5784 GND.n5783 0.479239
R4985 GND.n1194 GND.n1193 0.436742
R4986 GND.n1193 GND.n1192 0.436742
R4987 GND.n2219 GND.n2218 0.436742
R4988 GND.n2218 GND.n2217 0.436742
R4989 GND.n2543 GND.n2542 0.436742
R4990 GND.n2542 GND.n2541 0.436742
R4991 GND.n2868 GND.n2867 0.436742
R4992 GND.n2867 GND.n2866 0.436742
R4993 GND.n3165 GND.n3164 0.436742
R4994 GND.n3164 GND.n3163 0.436742
R4995 GND.n3322 GND.n3321 0.436742
R4996 GND.n3321 GND.n3320 0.436742
R4997 GND.n3480 GND.n3479 0.436742
R4998 GND.n3479 GND.n3478 0.436742
R4999 GND.n7270 GND.n7269 0.436742
R5000 GND.n7269 GND.n7268 0.436742
R5001 GND.n14 GND.n13 0.436742
R5002 GND.n13 GND.n12 0.436742
R5003 GND.n123 GND.n122 0.436742
R5004 GND.n122 GND.n121 0.436742
R5005 GND.n275 GND.n274 0.436742
R5006 GND.n274 GND.n273 0.436742
R5007 GND.n1638 GND.n1637 0.436742
R5008 GND.n1637 GND.n1636 0.436742
R5009 GND.n428 GND.n427 0.436742
R5010 GND.n427 GND.n426 0.436742
R5011 GND.n747 GND.n746 0.436742
R5012 GND.n746 GND.n745 0.436742
R5013 GND.n854 GND.n853 0.436742
R5014 GND.n853 GND.n852 0.436742
R5015 GND.n7793 GND.n7792 0.436742
R5016 GND.n7792 GND.n7791 0.436742
R5017 GND.n3632 GND.n3631 0.427167
R5018 GND.n3871 GND.n3870 0.427167
R5019 GND.n1560 GND.n1559 0.425574
R5020 GND.n1749 GND.n1748 0.425574
R5021 GND.n7021 GND.n7020 0.425574
R5022 GND.n2398 GND.n2397 0.425574
R5023 GND.n2723 GND.n2722 0.425574
R5024 GND.n3047 GND.n3046 0.425574
R5025 GND.n7147 GND.n7146 0.425574
R5026 GND.n4840 GND.n4839 0.425574
R5027 GND.n5416 GND.n5415 0.425574
R5028 GND.n5911 GND.n5910 0.425574
R5029 GND.n5986 GND.n5985 0.425574
R5030 GND.n6153 GND.n6152 0.425574
R5031 GND.n6317 GND.n6316 0.425574
R5032 GND.n605 GND.n604 0.425574
R5033 GND.n7648 GND.n7647 0.425574
R5034 GND.n7528 GND.n7527 0.425574
R5035 GND.n6759 GND.n6758 0.414845
R5036 GND.n6841 GND.n4422 0.414845
R5037 GND GND.n7823 0.383725
R5038 GND.n1615 GND.n1598 0.38056
R5039 GND.n1806 GND.n1789 0.38056
R5040 GND.n6971 GND.n6954 0.38056
R5041 GND.n2455 GND.n2438 0.38056
R5042 GND.n2780 GND.n2763 0.38056
R5043 GND.n3104 GND.n3087 0.38056
R5044 GND.n7204 GND.n7187 0.38056
R5045 GND.n4897 GND.n4880 0.38056
R5046 GND.n5338 GND.n5321 0.38056
R5047 GND.n5860 GND.n5843 0.38056
R5048 GND.n6043 GND.n6026 0.38056
R5049 GND.n6207 GND.n6190 0.38056
R5050 GND.n6371 GND.n6354 0.38056
R5051 GND.n659 GND.n642 0.38056
R5052 GND.n7706 GND.n7689 0.38056
R5053 GND.n7570 GND.n7558 0.38056
R5054 GND.n7826 GND.n895 0.378813
R5055 GND.n7829 GND.n788 0.378813
R5056 GND.n7832 GND.n469 0.378813
R5057 GND.n1687 GND.n1325 0.378813
R5058 GND.n7835 GND.n316 0.378813
R5059 GND.n7838 GND.n164 0.378813
R5060 GND.n7841 GND.n55 0.378813
R5061 GND.n7318 GND.n7311 0.378813
R5062 GND.n7322 GND.n3521 0.378813
R5063 GND.n7325 GND.n3363 0.378813
R5064 GND.n7328 GND.n3206 0.378813
R5065 GND.n7331 GND.n2909 0.378813
R5066 GND.n7334 GND.n2584 0.378813
R5067 GND.n7337 GND.n2260 0.378813
R5068 GND.n2102 GND.n1235 0.378813
R5069 GND.n1587 GND.n1585 0.377583
R5070 GND.n1778 GND.n1776 0.377583
R5071 GND.n6943 GND.n6941 0.377583
R5072 GND.n2427 GND.n2425 0.377583
R5073 GND.n2752 GND.n2750 0.377583
R5074 GND.n3076 GND.n3074 0.377583
R5075 GND.n7176 GND.n7174 0.377583
R5076 GND.n4869 GND.n4867 0.377583
R5077 GND.n5310 GND.n5308 0.377583
R5078 GND.n5832 GND.n5830 0.377583
R5079 GND.n6015 GND.n6013 0.377583
R5080 GND.n6179 GND.n6177 0.377583
R5081 GND.n6343 GND.n6341 0.377583
R5082 GND.n631 GND.n629 0.377583
R5083 GND.n7678 GND.n7676 0.377583
R5084 GND.n7547 GND.n7545 0.377583
R5085 GND.n5493 GND.n5492 0.376971
R5086 GND.n6609 GND.n6608 0.376971
R5087 GND.n6519 GND.n6518 0.376971
R5088 GND.n6435 GND.n6434 0.376971
R5089 GND.n1899 GND.n1898 0.376971
R5090 GND.n1856 GND.n1855 0.376971
R5091 GND.n6881 GND.n6880 0.376971
R5092 GND.n2505 GND.n2504 0.376971
R5093 GND.n2830 GND.n2829 0.376971
R5094 GND.n3127 GND.n3126 0.376971
R5095 GND.n7227 GND.n7226 0.376971
R5096 GND.n4759 GND.n4758 0.376971
R5097 GND.n5248 GND.n5247 0.376971
R5098 GND.n5927 GND.n5926 0.376971
R5099 GND.n6096 GND.n6095 0.376971
R5100 GND.n6260 GND.n6259 0.376971
R5101 GND.n6569 GND.n6568 0.376971
R5102 GND.n709 GND.n708 0.376971
R5103 GND.n7756 GND.n7755 0.376971
R5104 GND.n7591 GND.n7590 0.376971
R5105 GND.n4654 GND.n4653 0.376971
R5106 GND.n4691 GND.n4690 0.376971
R5107 GND.n4716 GND.n4715 0.376971
R5108 GND.n5023 GND.n5022 0.376971
R5109 GND.n4584 GND.n4583 0.376971
R5110 GND.n5689 GND.n5688 0.376971
R5111 GND.n5775 GND.n5774 0.376971
R5112 GND.n5611 GND.n5610 0.376971
R5113 GND.n5527 GND.n5526 0.376971
R5114 GND.n4429 GND.n4428 0.376971
R5115 GND.n5051 GND.n5050 0.376971
R5116 GND.n4499 GND.n4498 0.376971
R5117 GND.n4487 GND.n4486 0.376971
R5118 GND.n6760 GND.n5464 0.375505
R5119 GND.n6842 GND.n4395 0.375505
R5120 GND.n1583 GND.n1580 0.3755
R5121 GND.n1774 GND.n1771 0.3755
R5122 GND.n6939 GND.n6936 0.3755
R5123 GND.n2423 GND.n2420 0.3755
R5124 GND.n2748 GND.n2745 0.3755
R5125 GND.n3072 GND.n3069 0.3755
R5126 GND.n7172 GND.n7169 0.3755
R5127 GND.n4865 GND.n4862 0.3755
R5128 GND.n5306 GND.n5303 0.3755
R5129 GND.n5828 GND.n5825 0.3755
R5130 GND.n6011 GND.n6008 0.3755
R5131 GND.n6175 GND.n6172 0.3755
R5132 GND.n6339 GND.n6336 0.3755
R5133 GND.n627 GND.n624 0.3755
R5134 GND.n7674 GND.n7671 0.3755
R5135 GND.n7543 GND.n7540 0.3755
R5136 GND.n1961 GND.n1959 0.373417
R5137 GND.n1959 GND.n1952 0.373417
R5138 GND.n1723 GND.n1721 0.373417
R5139 GND.n1721 GND.n1714 0.373417
R5140 GND.n1819 GND.n1817 0.373417
R5141 GND.n1817 GND.n1810 0.373417
R5142 GND.n6984 GND.n6982 0.373417
R5143 GND.n6982 GND.n6975 0.373417
R5144 GND.n2468 GND.n2466 0.373417
R5145 GND.n2466 GND.n2459 0.373417
R5146 GND.n2793 GND.n2791 0.373417
R5147 GND.n2791 GND.n2784 0.373417
R5148 GND.n7121 GND.n7119 0.373417
R5149 GND.n7119 GND.n7112 0.373417
R5150 GND.n4814 GND.n4812 0.373417
R5151 GND.n4812 GND.n4805 0.373417
R5152 GND.n5390 GND.n5388 0.373417
R5153 GND.n5388 GND.n5381 0.373417
R5154 GND.n5351 GND.n5349 0.373417
R5155 GND.n5349 GND.n5342 0.373417
R5156 GND.n5873 GND.n5871 0.373417
R5157 GND.n5871 GND.n5864 0.373417
R5158 GND.n6059 GND.n6057 0.373417
R5159 GND.n6057 GND.n6050 0.373417
R5160 GND.n6223 GND.n6221 0.373417
R5161 GND.n6221 GND.n6214 0.373417
R5162 GND.n6387 GND.n6385 0.373417
R5163 GND.n6385 GND.n6378 0.373417
R5164 GND.n672 GND.n670 0.373417
R5165 GND.n670 GND.n663 0.373417
R5166 GND.n7719 GND.n7717 0.373417
R5167 GND.n7717 GND.n7710 0.373417
R5168 GND.n7537 GND.n7536 0.366214
R5169 GND.n7668 GND.n7667 0.366214
R5170 GND.n6375 GND.n6374 0.366214
R5171 GND.n6211 GND.n6210 0.366214
R5172 GND.n6047 GND.n6046 0.366214
R5173 GND.n6005 GND.n6004 0.366214
R5174 GND.n5822 GND.n5821 0.366214
R5175 GND.n5300 GND.n5299 0.366214
R5176 GND.n4859 GND.n4858 0.366214
R5177 GND.n7166 GND.n7165 0.366214
R5178 GND.n3066 GND.n3065 0.366214
R5179 GND.n2742 GND.n2741 0.366214
R5180 GND.n2417 GND.n2416 0.366214
R5181 GND.n6933 GND.n6932 0.366214
R5182 GND.n1768 GND.n1767 0.366214
R5183 GND.n1577 GND.n1576 0.366214
R5184 GND.n1623 GND.n1622 0.355857
R5185 GND.n1841 GND.n1840 0.355857
R5186 GND.n7006 GND.n7005 0.355857
R5187 GND.n2490 GND.n2489 0.355857
R5188 GND.n2815 GND.n2814 0.355857
R5189 GND.n3112 GND.n3111 0.355857
R5190 GND.n7212 GND.n7211 0.355857
R5191 GND.n4905 GND.n4904 0.355857
R5192 GND.n5373 GND.n5372 0.355857
R5193 GND.n5895 GND.n5894 0.355857
R5194 GND.n6081 GND.n6080 0.355857
R5195 GND.n6245 GND.n6244 0.355857
R5196 GND.n6409 GND.n6408 0.355857
R5197 GND.n694 GND.n693 0.355857
R5198 GND.n7741 GND.n7740 0.355857
R5199 GND.n7577 GND.n7576 0.355857
R5200 GND.n7362 GND 0.354667
R5201 GND.n2015 GND 0.354667
R5202 GND.n513 GND 0.354667
R5203 GND.n208 GND 0.354667
R5204 GND.n1507 GND 0.354667
R5205 GND.n1459 GND 0.354667
R5206 GND.n4216 GND 0.354667
R5207 GND.n3410 GND 0.354667
R5208 GND.n3253 GND 0.354667
R5209 GND.n2956 GND 0.354667
R5210 GND.n2631 GND 0.354667
R5211 GND.n2307 GND 0.354667
R5212 GND.n2145 GND 0.354667
R5213 GND.n1277 GND 0.354667
R5214 GND.n360 GND 0.354667
R5215 GND.n7408 GND 0.354667
R5216 GND.n6599 GND.n6598 0.353
R5217 GND.n4035 GND.n3652 0.352931
R5218 GND.n4022 GND.n4021 0.352931
R5219 GND.n4006 GND.n4005 0.352931
R5220 GND.n3991 GND.n3990 0.352931
R5221 GND.n3976 GND.n3975 0.352931
R5222 GND.n3961 GND.n3960 0.352931
R5223 GND.n3944 GND.n3943 0.352931
R5224 GND.n3929 GND.n3928 0.352931
R5225 GND.n3914 GND.n3913 0.352931
R5226 GND.n3899 GND.n3898 0.352931
R5227 GND.n3863 GND.n3862 0.352931
R5228 GND.n3845 GND.n3844 0.352931
R5229 GND.n3820 GND.n3819 0.352931
R5230 GND.n3805 GND.n3804 0.352931
R5231 GND.n3790 GND.n3789 0.352931
R5232 GND.n3775 GND.n3774 0.352931
R5233 GND.n3756 GND.n3755 0.352931
R5234 GND.n3741 GND.n3740 0.352931
R5235 GND.n3726 GND.n3725 0.352931
R5236 GND.n3711 GND.n3710 0.352931
R5237 GND.n3884 GND.n3883 0.347722
R5238 GND.n1946 GND.n1554 0.345738
R5239 GND.n6762 GND.n6761 0.33677
R5240 GND.n6843 GND.n4373 0.33677
R5241 GND.n5041 GND.n5040 0.336652
R5242 GND.n6837 GND 0.327423
R5243 GND.n7082 GND 0.327423
R5244 GND.n5438 GND.n5437 0.326891
R5245 GND.n6869 GND.n4339 0.326891
R5246 GND.n5217 GND.n4423 0.325812
R5247 GND.n6871 GND.n6870 0.325812
R5248 GND.n7367 GND.n7366 0.321569
R5249 GND.n7437 GND.n7435 0.321569
R5250 GND.n1996 GND.n1988 0.321569
R5251 GND.n2019 GND.n2018 0.321569
R5252 GND.n332 GND.n320 0.321569
R5253 GND.n517 GND.n516 0.321569
R5254 GND.n485 GND.n473 0.321569
R5255 GND.n212 GND.n211 0.321569
R5256 GND.n180 GND.n168 0.321569
R5257 GND.n1511 GND.n1510 0.321569
R5258 GND.n1515 GND.n1514 0.321569
R5259 GND.n1463 GND.n1462 0.321569
R5260 GND.n1467 GND.n1466 0.321569
R5261 GND.n4220 GND.n4219 0.321569
R5262 GND.n4188 GND.n4176 0.321569
R5263 GND.n3414 GND.n3413 0.321569
R5264 GND.n3382 GND.n3370 0.321569
R5265 GND.n3257 GND.n3256 0.321569
R5266 GND.n3225 GND.n3213 0.321569
R5267 GND.n2960 GND.n2959 0.321569
R5268 GND.n2928 GND.n2916 0.321569
R5269 GND.n2635 GND.n2634 0.321569
R5270 GND.n2603 GND.n2591 0.321569
R5271 GND.n2311 GND.n2310 0.321569
R5272 GND.n2279 GND.n2267 0.321569
R5273 GND.n2149 GND.n2148 0.321569
R5274 GND.n2117 GND.n2105 0.321569
R5275 GND.n1281 GND.n1280 0.321569
R5276 GND.n1249 GND.n1237 0.321569
R5277 GND.n364 GND.n363 0.321569
R5278 GND.n7416 GND.n7415 0.321569
R5279 GND.n7412 GND.n7411 0.321569
R5280 GND.n4059 GND.n4056 0.3205
R5281 GND.n5040 GND.n5039 0.31982
R5282 GND.n7493 GND.n7438 0.314812
R5283 GND.n2082 GND.n2020 0.314812
R5284 GND.n570 GND.n518 0.314812
R5285 GND.n261 GND.n213 0.314812
R5286 GND.n1512 GND.n109 0.314812
R5287 GND.n1464 GND.n1442 0.314812
R5288 GND.n4269 GND.n4221 0.314812
R5289 GND.n3466 GND.n3415 0.314812
R5290 GND.n3308 GND.n3258 0.314812
R5291 GND.n3012 GND.n2961 0.314812
R5292 GND.n2688 GND.n2636 0.314812
R5293 GND.n2363 GND.n2312 0.314812
R5294 GND.n2205 GND.n2150 0.314812
R5295 GND.n1324 GND.n1282 0.314812
R5296 GND.n414 GND.n365 0.314812
R5297 GND.n7413 GND.n840 0.314812
R5298 GND.n1975 GND.n1972 0.313
R5299 GND.n1737 GND.n1734 0.313
R5300 GND.n1833 GND.n1830 0.313
R5301 GND.n6998 GND.n6995 0.313
R5302 GND.n2482 GND.n2479 0.313
R5303 GND.n2807 GND.n2804 0.313
R5304 GND.n7135 GND.n7132 0.313
R5305 GND.n4828 GND.n4825 0.313
R5306 GND.n5404 GND.n5401 0.313
R5307 GND.n5365 GND.n5362 0.313
R5308 GND.n5887 GND.n5884 0.313
R5309 GND.n6073 GND.n6070 0.313
R5310 GND.n6237 GND.n6234 0.313
R5311 GND.n6401 GND.n6398 0.313
R5312 GND.n686 GND.n683 0.313
R5313 GND.n7733 GND.n7730 0.313
R5314 GND.n6599 GND.n5784 0.309146
R5315 GND.n4038 GND.n4035 0.302583
R5316 GND GND.n5489 0.295209
R5317 GND GND.n4420 0.295209
R5318 GND.n7362 GND.n7360 0.295052
R5319 GND.n2015 GND.n2013 0.295052
R5320 GND.n513 GND.n511 0.295052
R5321 GND.n208 GND.n206 0.295052
R5322 GND.n1507 GND.n1505 0.295052
R5323 GND.n1459 GND.n1457 0.295052
R5324 GND.n4216 GND.n4214 0.295052
R5325 GND.n3410 GND.n3408 0.295052
R5326 GND.n3253 GND.n3251 0.295052
R5327 GND.n2956 GND.n2954 0.295052
R5328 GND.n2631 GND.n2629 0.295052
R5329 GND.n2307 GND.n2305 0.295052
R5330 GND.n2145 GND.n2143 0.295052
R5331 GND.n1277 GND.n1275 0.295052
R5332 GND.n360 GND.n358 0.295052
R5333 GND.n7408 GND.n7406 0.295052
R5334 GND.n1575 GND.n1573 0.290381
R5335 GND.n1766 GND.n1764 0.290381
R5336 GND.n6931 GND.n6929 0.290381
R5337 GND.n2415 GND.n2413 0.290381
R5338 GND.n2740 GND.n2738 0.290381
R5339 GND.n3064 GND.n3062 0.290381
R5340 GND.n7164 GND.n7162 0.290381
R5341 GND.n4857 GND.n4855 0.290381
R5342 GND.n5298 GND.n5296 0.290381
R5343 GND.n5820 GND.n5818 0.290381
R5344 GND.n6003 GND.n6001 0.290381
R5345 GND.n6170 GND.n6168 0.290381
R5346 GND.n6334 GND.n6332 0.290381
R5347 GND.n622 GND.n620 0.290381
R5348 GND.n7666 GND.n7664 0.290381
R5349 GND.n7535 GND.n7533 0.290381
R5350 GND.n7252 GND.n7085 0.283189
R5351 GND.n5463 GND.n5462 0.280127
R5352 GND.n6868 GND.n6867 0.280127
R5353 GND.n3638 GND.n3637 0.270108
R5354 GND.n4072 GND.n4071 0.260982
R5355 GND.n4071 GND.n4070 0.2605
R5356 GND.n1589 GND.n1587 0.24425
R5357 GND.n1780 GND.n1778 0.24425
R5358 GND.n6945 GND.n6943 0.24425
R5359 GND.n2429 GND.n2427 0.24425
R5360 GND.n2754 GND.n2752 0.24425
R5361 GND.n3078 GND.n3076 0.24425
R5362 GND.n7178 GND.n7176 0.24425
R5363 GND.n4871 GND.n4869 0.24425
R5364 GND.n5312 GND.n5310 0.24425
R5365 GND.n5834 GND.n5832 0.24425
R5366 GND.n6017 GND.n6015 0.24425
R5367 GND.n6181 GND.n6179 0.24425
R5368 GND.n6345 GND.n6343 0.24425
R5369 GND.n633 GND.n631 0.24425
R5370 GND.n7680 GND.n7678 0.24425
R5371 GND.n7549 GND.n7547 0.24425
R5372 GND.n1945 GND.n1944 0.243155
R5373 GND.n1751 GND.n1750 0.243155
R5374 GND.n7023 GND.n7022 0.243155
R5375 GND.n2400 GND.n2399 0.243155
R5376 GND.n2725 GND.n2724 0.243155
R5377 GND.n3049 GND.n3048 0.243155
R5378 GND.n7149 GND.n7148 0.243155
R5379 GND.n4842 GND.n4841 0.243155
R5380 GND.n5418 GND.n5417 0.243155
R5381 GND.n5913 GND.n5912 0.243155
R5382 GND.n5988 GND.n5987 0.243155
R5383 GND.n6155 GND.n6154 0.243155
R5384 GND.n6319 GND.n6318 0.243155
R5385 GND.n607 GND.n606 0.243155
R5386 GND.n7650 GND.n7649 0.243155
R5387 GND.n7530 GND.n7529 0.243155
R5388 GND.n1963 GND.n1961 0.238893
R5389 GND.n1725 GND.n1723 0.238893
R5390 GND.n1821 GND.n1819 0.238893
R5391 GND.n6986 GND.n6984 0.238893
R5392 GND.n2470 GND.n2468 0.238893
R5393 GND.n2795 GND.n2793 0.238893
R5394 GND.n7123 GND.n7121 0.238893
R5395 GND.n4816 GND.n4814 0.238893
R5396 GND.n5392 GND.n5390 0.238893
R5397 GND.n5353 GND.n5351 0.238893
R5398 GND.n5875 GND.n5873 0.238893
R5399 GND.n6061 GND.n6059 0.238893
R5400 GND.n6225 GND.n6223 0.238893
R5401 GND.n6389 GND.n6387 0.238893
R5402 GND.n674 GND.n672 0.238893
R5403 GND.n7721 GND.n7719 0.238893
R5404 GND.n4933 GND 0.228789
R5405 GND.n5474 GND.n5470 0.226583
R5406 GND.n4405 GND.n4401 0.226583
R5407 GND.n1942 GND.n1920 0.224247
R5408 GND.n1877 GND.n1709 0.224247
R5409 GND.n7029 GND.n7025 0.224247
R5410 GND.n2526 GND.n2385 0.224247
R5411 GND.n2851 GND.n2710 0.224247
R5412 GND.n3148 GND.n3034 0.224247
R5413 GND.n7248 GND.n7107 0.224247
R5414 GND.n4802 GND.n4780 0.224247
R5415 GND.n5421 GND.n5420 0.224247
R5416 GND.n5948 GND.n5915 0.224247
R5417 GND.n6117 GND.n5973 0.224247
R5418 GND.n6281 GND.n6140 0.224247
R5419 GND.n6590 GND.n6304 0.224247
R5420 GND.n730 GND.n592 0.224247
R5421 GND.n7777 GND.n7635 0.224247
R5422 GND.n7612 GND.n7515 0.224247
R5423 GND.n4589 GND 0.209082
R5424 GND.n1950 GND.n1948 0.200996
R5425 GND.n1743 GND.n1741 0.200996
R5426 GND.n7015 GND.n7013 0.200996
R5427 GND.n2392 GND.n2390 0.200996
R5428 GND.n2717 GND.n2715 0.200996
R5429 GND.n3041 GND.n3039 0.200996
R5430 GND.n7141 GND.n7139 0.200996
R5431 GND.n4834 GND.n4832 0.200996
R5432 GND.n5410 GND.n5408 0.200996
R5433 GND.n5905 GND.n5903 0.200996
R5434 GND.n5980 GND.n5978 0.200996
R5435 GND.n6147 GND.n6145 0.200996
R5436 GND.n6311 GND.n6309 0.200996
R5437 GND.n599 GND.n597 0.200996
R5438 GND.n7642 GND.n7640 0.200996
R5439 GND.n7522 GND.n7520 0.200996
R5440 GND.n7431 GND.n7381 0.197423
R5441 GND.n1984 GND.n1377 0.197423
R5442 GND.n340 GND.n322 0.197423
R5443 GND.n493 GND.n475 0.197423
R5444 GND.n188 GND.n170 0.197423
R5445 GND.n1523 GND.n1479 0.197423
R5446 GND.n1475 GND.n1378 0.197423
R5447 GND.n4196 GND.n4178 0.197423
R5448 GND.n3390 GND.n3372 0.197423
R5449 GND.n3233 GND.n3215 0.197423
R5450 GND.n2936 GND.n2918 0.197423
R5451 GND.n2611 GND.n2593 0.197423
R5452 GND.n2287 GND.n2269 0.197423
R5453 GND.n2125 GND.n2107 0.197423
R5454 GND.n1257 GND.n1239 0.197423
R5455 GND.n7424 GND.n7387 0.197423
R5456 GND.n3640 GND.n3639 0.196239
R5457 GND.n3642 GND.n3641 0.190273
R5458 GND.n6773 GND.n6770 0.189094
R5459 GND.n5231 GND.n5230 0.189094
R5460 GND.n4351 GND.n4348 0.189094
R5461 GND.n4323 GND.n4322 0.189094
R5462 GND.n3647 GND.n3642 0.188284
R5463 GND.n4063 GND.n3650 0.181849
R5464 GND.n1624 GND.n1623 0.181736
R5465 GND.n1842 GND.n1841 0.181736
R5466 GND.n7011 GND.n7006 0.181736
R5467 GND.n2491 GND.n2490 0.181736
R5468 GND.n2816 GND.n2815 0.181736
R5469 GND.n3113 GND.n3112 0.181736
R5470 GND.n7213 GND.n7212 0.181736
R5471 GND.n4906 GND.n4905 0.181736
R5472 GND.n5379 GND.n5373 0.181736
R5473 GND.n5901 GND.n5895 0.181736
R5474 GND.n6082 GND.n6081 0.181736
R5475 GND.n6246 GND.n6245 0.181736
R5476 GND.n6410 GND.n6409 0.181736
R5477 GND.n695 GND.n694 0.181736
R5478 GND.n7742 GND.n7741 0.181736
R5479 GND.n7578 GND.n7577 0.181736
R5480 GND.n3639 GND.n3638 0.178057
R5481 GND.n1944 GND.n1624 0.17675
R5482 GND.n1842 GND.n1751 0.17675
R5483 GND.n7023 GND.n7011 0.17675
R5484 GND.n2491 GND.n2400 0.17675
R5485 GND.n2816 GND.n2725 0.17675
R5486 GND.n3113 GND.n3049 0.17675
R5487 GND.n7213 GND.n7149 0.17675
R5488 GND.n4906 GND.n4842 0.17675
R5489 GND.n5418 GND.n5379 0.17675
R5490 GND.n5913 GND.n5901 0.17675
R5491 GND.n6082 GND.n5988 0.17675
R5492 GND.n6246 GND.n6155 0.17675
R5493 GND.n6410 GND.n6319 0.17675
R5494 GND.n695 GND.n607 0.17675
R5495 GND.n7742 GND.n7650 0.17675
R5496 GND.n7578 GND.n7530 0.17675
R5497 GND.t730 GND.t1246 0.176676
R5498 GND.n3684 GND.n3669 0.176676
R5499 GND.n1591 GND.n1589 0.171333
R5500 GND.n1782 GND.n1780 0.171333
R5501 GND.n6947 GND.n6945 0.171333
R5502 GND.n2431 GND.n2429 0.171333
R5503 GND.n2756 GND.n2754 0.171333
R5504 GND.n3080 GND.n3078 0.171333
R5505 GND.n7180 GND.n7178 0.171333
R5506 GND.n4873 GND.n4871 0.171333
R5507 GND.n5314 GND.n5312 0.171333
R5508 GND.n5836 GND.n5834 0.171333
R5509 GND.n6019 GND.n6017 0.171333
R5510 GND.n6183 GND.n6181 0.171333
R5511 GND.n6347 GND.n6345 0.171333
R5512 GND.n635 GND.n633 0.171333
R5513 GND.n7682 GND.n7680 0.171333
R5514 GND.n7551 GND.n7549 0.171333
R5515 GND.n1598 GND.n1595 0.16925
R5516 GND.n1789 GND.n1786 0.16925
R5517 GND.n6954 GND.n6951 0.16925
R5518 GND.n2438 GND.n2435 0.16925
R5519 GND.n2763 GND.n2760 0.16925
R5520 GND.n3087 GND.n3084 0.16925
R5521 GND.n7187 GND.n7184 0.16925
R5522 GND.n4880 GND.n4877 0.16925
R5523 GND.n5321 GND.n5318 0.16925
R5524 GND.n5843 GND.n5840 0.16925
R5525 GND.n6026 GND.n6023 0.16925
R5526 GND.n6190 GND.n6187 0.16925
R5527 GND.n6354 GND.n6351 0.16925
R5528 GND.n642 GND.n639 0.16925
R5529 GND.n7689 GND.n7686 0.16925
R5530 GND.n7558 GND.n7555 0.16925
R5531 GND.n4272 GND 0.165163
R5532 GND.n1976 GND.n1950 0.164786
R5533 GND.n1976 GND.n1975 0.164786
R5534 GND.n1741 GND.n1739 0.164786
R5535 GND.n1739 GND.n1737 0.164786
R5536 GND.n1834 GND.n1833 0.164786
R5537 GND.n6999 GND.n6998 0.164786
R5538 GND.n2483 GND.n2482 0.164786
R5539 GND.n2808 GND.n2807 0.164786
R5540 GND.n7139 GND.n7137 0.164786
R5541 GND.n7137 GND.n7135 0.164786
R5542 GND.n4832 GND.n4830 0.164786
R5543 GND.n4830 GND.n4828 0.164786
R5544 GND.n5408 GND.n5406 0.164786
R5545 GND.n5406 GND.n5404 0.164786
R5546 GND.n5366 GND.n5365 0.164786
R5547 GND.n5888 GND.n5887 0.164786
R5548 GND.n6074 GND.n6073 0.164786
R5549 GND.n6238 GND.n6237 0.164786
R5550 GND.n6402 GND.n6401 0.164786
R5551 GND.n687 GND.n686 0.164786
R5552 GND.n7734 GND.n7733 0.164786
R5553 GND.n1617 GND.n1615 0.159429
R5554 GND.n1808 GND.n1806 0.159429
R5555 GND.n6973 GND.n6971 0.159429
R5556 GND.n2457 GND.n2455 0.159429
R5557 GND.n2782 GND.n2780 0.159429
R5558 GND.n3106 GND.n3104 0.159429
R5559 GND.n7206 GND.n7204 0.159429
R5560 GND.n4899 GND.n4897 0.159429
R5561 GND.n5340 GND.n5338 0.159429
R5562 GND.n5862 GND.n5860 0.159429
R5563 GND.n6045 GND.n6043 0.159429
R5564 GND.n6209 GND.n6207 0.159429
R5565 GND.n6373 GND.n6371 0.159429
R5566 GND.n661 GND.n659 0.159429
R5567 GND.n7708 GND.n7706 0.159429
R5568 GND.n7572 GND.n7570 0.159429
R5569 GND.n6837 GND.n6836 0.15606
R5570 GND.n7082 GND.n7081 0.15606
R5571 GND.n1972 GND.n1969 0.148714
R5572 GND.n1967 GND.n1963 0.148714
R5573 GND.n1734 GND.n1731 0.148714
R5574 GND.n1729 GND.n1725 0.148714
R5575 GND.n1830 GND.n1827 0.148714
R5576 GND.n1825 GND.n1821 0.148714
R5577 GND.n6995 GND.n6992 0.148714
R5578 GND.n6990 GND.n6986 0.148714
R5579 GND.n2479 GND.n2476 0.148714
R5580 GND.n2474 GND.n2470 0.148714
R5581 GND.n2804 GND.n2801 0.148714
R5582 GND.n2799 GND.n2795 0.148714
R5583 GND.n7132 GND.n7129 0.148714
R5584 GND.n7127 GND.n7123 0.148714
R5585 GND.n4825 GND.n4822 0.148714
R5586 GND.n4820 GND.n4816 0.148714
R5587 GND.n5401 GND.n5398 0.148714
R5588 GND.n5396 GND.n5392 0.148714
R5589 GND.n5362 GND.n5359 0.148714
R5590 GND.n5357 GND.n5353 0.148714
R5591 GND.n5884 GND.n5881 0.148714
R5592 GND.n5879 GND.n5875 0.148714
R5593 GND.n6070 GND.n6067 0.148714
R5594 GND.n6065 GND.n6061 0.148714
R5595 GND.n6234 GND.n6231 0.148714
R5596 GND.n6229 GND.n6225 0.148714
R5597 GND.n6398 GND.n6395 0.148714
R5598 GND.n6393 GND.n6389 0.148714
R5599 GND.n683 GND.n680 0.148714
R5600 GND.n678 GND.n674 0.148714
R5601 GND.n7730 GND.n7727 0.148714
R5602 GND.n7725 GND.n7721 0.148714
R5603 GND.n3648 GND.n3647 0.148287
R5604 GND.n790 GND.n789 0.142154
R5605 GND.n7354 GND.n7353 0.142154
R5606 GND.n2086 GND.n2085 0.142154
R5607 GND.n318 GND.n317 0.142154
R5608 GND.n471 GND.n470 0.142154
R5609 GND.n166 GND.n165 0.142154
R5610 GND.n57 GND.n56 0.142154
R5611 GND.n7316 GND.n7315 0.142154
R5612 GND.n4174 GND.n4173 0.142154
R5613 GND.n3368 GND.n3367 0.142154
R5614 GND.n3211 GND.n3210 0.142154
R5615 GND.n2914 GND.n2913 0.142154
R5616 GND.n2589 GND.n2588 0.142154
R5617 GND.n2265 GND.n2264 0.142154
R5618 GND.n7341 GND.n7340 0.142154
R5619 GND.n2099 GND.n2098 0.142154
R5620 GND.n4030 GND.n4029 0.141472
R5621 GND.n4029 GND.n4027 0.141472
R5622 GND.n4027 GND.n4014 0.141472
R5623 GND.n4014 GND.n4012 0.141472
R5624 GND.n4012 GND.n3999 0.141472
R5625 GND.n3999 GND.n3997 0.141472
R5626 GND.n3997 GND.n3984 0.141472
R5627 GND.n3984 GND.n3982 0.141472
R5628 GND.n3982 GND.n3969 0.141472
R5629 GND.n3969 GND.n3967 0.141472
R5630 GND.n3952 GND.n3950 0.141472
R5631 GND.n3950 GND.n3937 0.141472
R5632 GND.n3937 GND.n3935 0.141472
R5633 GND.n3935 GND.n3922 0.141472
R5634 GND.n3922 GND.n3920 0.141472
R5635 GND.n3920 GND.n3907 0.141472
R5636 GND.n3907 GND.n3905 0.141472
R5637 GND.n3905 GND.n3892 0.141472
R5638 GND.n3892 GND.n3890 0.141472
R5639 GND.n3872 GND.n3869 0.141472
R5640 GND.n3853 GND.n3851 0.141472
R5641 GND.n3851 GND.n3828 0.141472
R5642 GND.n3828 GND.n3826 0.141472
R5643 GND.n3826 GND.n3813 0.141472
R5644 GND.n3813 GND.n3811 0.141472
R5645 GND.n3811 GND.n3798 0.141472
R5646 GND.n3798 GND.n3796 0.141472
R5647 GND.n3796 GND.n3783 0.141472
R5648 GND.n3783 GND.n3781 0.141472
R5649 GND.n3765 GND.n3762 0.141472
R5650 GND.n3762 GND.n3749 0.141472
R5651 GND.n3749 GND.n3747 0.141472
R5652 GND.n3747 GND.n3734 0.141472
R5653 GND.n3734 GND.n3732 0.141472
R5654 GND.n3732 GND.n3719 0.141472
R5655 GND.n3719 GND.n3717 0.141472
R5656 GND.n3717 GND.n3704 0.141472
R5657 GND.n3704 GND.n3702 0.141472
R5658 GND.n91 GND.n90 0.140882
R5659 GND.n6838 GND 0.140869
R5660 GND.n7083 GND 0.140869
R5661 GND.n3890 GND.n3875 0.136611
R5662 GND.n6758 GND 0.134348
R5663 GND.n4422 GND 0.134348
R5664 GND.n3668 GND.n3667 0.134262
R5665 GND.n403 GND.n402 0.131784
R5666 GND.n1432 GND.n1431 0.131784
R5667 GND.n1433 GND.n1432 0.131784
R5668 GND.n3456 GND.n3455 0.131784
R5669 GND.n3457 GND.n3456 0.131784
R5670 GND.n3002 GND.n3001 0.131784
R5671 GND.n3003 GND.n3002 0.131784
R5672 GND.n2353 GND.n2352 0.131784
R5673 GND.n2354 GND.n2353 0.131784
R5674 GND.n1312 GND.n1311 0.131784
R5675 GND.n2195 GND.n2194 0.131784
R5676 GND.n2196 GND.n2195 0.131784
R5677 GND.n2678 GND.n2677 0.131784
R5678 GND.n2679 GND.n2678 0.131784
R5679 GND.n3298 GND.n3297 0.131784
R5680 GND.n3299 GND.n3298 0.131784
R5681 GND.n4259 GND.n4258 0.131784
R5682 GND.n4260 GND.n4259 0.131784
R5683 GND.n99 GND.n98 0.131784
R5684 GND.n100 GND.n99 0.131784
R5685 GND.n251 GND.n250 0.131784
R5686 GND.n252 GND.n251 0.131784
R5687 GND.n2071 GND.n2070 0.131784
R5688 GND.n829 GND.n828 0.131784
R5689 GND.n560 GND.n559 0.131784
R5690 GND.n561 GND.n560 0.131784
R5691 GND.n7483 GND.n7482 0.131784
R5692 GND.n7484 GND.n7483 0.131784
R5693 GND.n406 GND.n403 0.13084
R5694 GND.n1315 GND.n1312 0.13084
R5695 GND.n2074 GND.n2071 0.13084
R5696 GND.n832 GND.n829 0.13084
R5697 GND.n6836 GND.n6835 0.12814
R5698 GND.n7081 GND.n7080 0.12814
R5699 GND.n3679 GND.n3677 0.127732
R5700 GND.n405 GND.n404 0.126877
R5701 GND.n1427 GND.n1426 0.126877
R5702 GND.n3451 GND.n3450 0.126877
R5703 GND.n2997 GND.n2996 0.126877
R5704 GND.n2348 GND.n2347 0.126877
R5705 GND.n1314 GND.n1313 0.126877
R5706 GND.n2190 GND.n2189 0.126877
R5707 GND.n2673 GND.n2672 0.126877
R5708 GND.n3293 GND.n3292 0.126877
R5709 GND.n4254 GND.n4253 0.126877
R5710 GND.n85 GND.n84 0.126877
R5711 GND.n246 GND.n245 0.126877
R5712 GND.n2073 GND.n2072 0.126877
R5713 GND.n831 GND.n830 0.126877
R5714 GND.n555 GND.n554 0.126877
R5715 GND.n7474 GND.n7473 0.126877
R5716 GND.n2074 GND.n2073 0.125988
R5717 GND.n406 GND.n405 0.125988
R5718 GND.n1315 GND.n1314 0.125988
R5719 GND.n832 GND.n831 0.125988
R5720 GND.n1434 GND.n1427 0.125687
R5721 GND.n3458 GND.n3451 0.125687
R5722 GND.n3004 GND.n2997 0.125687
R5723 GND.n2355 GND.n2348 0.125687
R5724 GND.n2197 GND.n2190 0.125687
R5725 GND.n2680 GND.n2673 0.125687
R5726 GND.n3300 GND.n3293 0.125687
R5727 GND.n4261 GND.n4254 0.125687
R5728 GND.n101 GND.n85 0.125687
R5729 GND.n253 GND.n246 0.125687
R5730 GND.n562 GND.n555 0.125687
R5731 GND.n7485 GND.n7474 0.125687
R5732 GND.n3781 GND.n3768 0.1255
R5733 GND.n1883 GND.n1882 0.122252
R5734 GND.n1880 GND.n1878 0.122252
R5735 GND.n7028 GND.n7027 0.122252
R5736 GND.n2528 GND.n2527 0.122252
R5737 GND.n2853 GND.n2852 0.122252
R5738 GND.n3150 GND.n3149 0.122252
R5739 GND.n7250 GND.n7249 0.122252
R5740 GND.n7253 GND.n4271 0.122252
R5741 GND.n7255 GND.n4270 0.122252
R5742 GND.n5950 GND.n5949 0.122252
R5743 GND.n6597 GND.n6118 0.122252
R5744 GND.n6595 GND.n6282 0.122252
R5745 GND.n6593 GND.n6591 0.122252
R5746 GND.n732 GND.n731 0.122252
R5747 GND.n7779 GND.n7778 0.122252
R5748 GND.n7781 GND.n7613 0.122252
R5749 GND.n1893 GND.n1892 0.122064
R5750 GND.n1850 GND.n1849 0.122064
R5751 GND.n7042 GND.n7041 0.122064
R5752 GND.n2499 GND.n2498 0.122064
R5753 GND.n2824 GND.n2823 0.122064
R5754 GND.n3121 GND.n3120 0.122064
R5755 GND.n7221 GND.n7220 0.122064
R5756 GND.n4753 GND.n4752 0.122064
R5757 GND.n5434 GND.n5433 0.122064
R5758 GND.n6090 GND.n6089 0.122064
R5759 GND.n5921 GND.n5920 0.122064
R5760 GND.n6254 GND.n6253 0.122064
R5761 GND.n6563 GND.n6562 0.122064
R5762 GND.n703 GND.n702 0.122064
R5763 GND.n7750 GND.n7749 0.122064
R5764 GND.n7585 GND.n7584 0.122064
R5765 GND.n3648 GND.n2103 0.118
R5766 GND.n3610 GND.n3547 0.117951
R5767 GND.t52 GND.t422 0.117951
R5768 GND.t432 GND.t77 0.117951
R5769 GND.t123 GND.t24 0.117951
R5770 GND.t59 GND.t51 0.117951
R5771 GND.t33 GND.t709 0.117951
R5772 GND.t106 GND.t122 0.117951
R5773 GND.t78 GND.t214 0.117951
R5774 GND.t202 GND.t394 0.117951
R5775 GND.n3702 GND.n3696 0.117167
R5776 GND.n6832 GND.n6831 0.1155
R5777 GND.n6831 GND.n6829 0.1155
R5778 GND.n6826 GND.n6825 0.1155
R5779 GND.n6825 GND.n6823 0.1155
R5780 GND.n6820 GND.n6819 0.1155
R5781 GND.n6819 GND.n6817 0.1155
R5782 GND.n6814 GND.n6813 0.1155
R5783 GND.n6813 GND.n6811 0.1155
R5784 GND.n7077 GND.n7076 0.1155
R5785 GND.n7076 GND.n7074 0.1155
R5786 GND.n7071 GND.n7070 0.1155
R5787 GND.n7070 GND.n7068 0.1155
R5788 GND.n7065 GND.n7064 0.1155
R5789 GND.n7064 GND.n7062 0.1155
R5790 GND.n7059 GND.n7058 0.1155
R5791 GND.n7058 GND.n7056 0.1155
R5792 GND.n1946 GND.n1945 0.112135
R5793 GND.n1750 GND.n1744 0.112135
R5794 GND.n7022 GND.n7016 0.112135
R5795 GND.n2399 GND.n2393 0.112135
R5796 GND.n2724 GND.n2718 0.112135
R5797 GND.n3048 GND.n3042 0.112135
R5798 GND.n7148 GND.n7142 0.112135
R5799 GND.n4841 GND.n4835 0.112135
R5800 GND.n5417 GND.n5411 0.112135
R5801 GND.n5912 GND.n5906 0.112135
R5802 GND.n5987 GND.n5981 0.112135
R5803 GND.n6154 GND.n6148 0.112135
R5804 GND.n6318 GND.n6312 0.112135
R5805 GND.n606 GND.n600 0.112135
R5806 GND.n7649 GND.n7643 0.112135
R5807 GND.n7529 GND.n7523 0.112135
R5808 GND.n5489 GND.n5465 0.110055
R5809 GND.n4420 GND.n4396 0.110055
R5810 GND.n1213 GND.n1212 0.10956
R5811 GND.t89 GND.n1213 0.10956
R5812 GND.n1219 GND.n1218 0.10956
R5813 GND.t89 GND.n1219 0.10956
R5814 GND.n1208 GND.n1207 0.10956
R5815 GND.n1207 GND.n1206 0.10956
R5816 GND.n1185 GND.n1184 0.10956
R5817 GND.n1184 GND.n1183 0.10956
R5818 GND.n1227 GND.n1226 0.10956
R5819 GND.t119 GND.n1227 0.10956
R5820 GND.t119 GND.n1225 0.10956
R5821 GND.n1225 GND.n1224 0.10956
R5822 GND.n2238 GND.n2237 0.10956
R5823 GND.t694 GND.n2238 0.10956
R5824 GND.n2244 GND.n2243 0.10956
R5825 GND.t694 GND.n2244 0.10956
R5826 GND.n2233 GND.n2232 0.10956
R5827 GND.n2232 GND.n2231 0.10956
R5828 GND.n2210 GND.n2209 0.10956
R5829 GND.n2209 GND.n2208 0.10956
R5830 GND.n2252 GND.n2251 0.10956
R5831 GND.t806 GND.n2252 0.10956
R5832 GND.t806 GND.n2250 0.10956
R5833 GND.n2250 GND.n2249 0.10956
R5834 GND.n2562 GND.n2561 0.10956
R5835 GND.t1308 GND.n2562 0.10956
R5836 GND.n2568 GND.n2567 0.10956
R5837 GND.t1308 GND.n2568 0.10956
R5838 GND.n2557 GND.n2556 0.10956
R5839 GND.n2556 GND.n2555 0.10956
R5840 GND.n2534 GND.n2533 0.10956
R5841 GND.n2533 GND.n2532 0.10956
R5842 GND.n2576 GND.n2575 0.10956
R5843 GND.t419 GND.n2576 0.10956
R5844 GND.t419 GND.n2574 0.10956
R5845 GND.n2574 GND.n2573 0.10956
R5846 GND.n2887 GND.n2886 0.10956
R5847 GND.t434 GND.n2887 0.10956
R5848 GND.n2893 GND.n2892 0.10956
R5849 GND.t434 GND.n2893 0.10956
R5850 GND.n2882 GND.n2881 0.10956
R5851 GND.n2881 GND.n2880 0.10956
R5852 GND.n2859 GND.n2858 0.10956
R5853 GND.n2858 GND.n2857 0.10956
R5854 GND.n2901 GND.n2900 0.10956
R5855 GND.t1187 GND.n2901 0.10956
R5856 GND.t1187 GND.n2899 0.10956
R5857 GND.n2899 GND.n2898 0.10956
R5858 GND.n3184 GND.n3183 0.10956
R5859 GND.t94 GND.n3184 0.10956
R5860 GND.n3190 GND.n3189 0.10956
R5861 GND.t94 GND.n3190 0.10956
R5862 GND.n3179 GND.n3178 0.10956
R5863 GND.n3178 GND.n3177 0.10956
R5864 GND.n3156 GND.n3155 0.10956
R5865 GND.n3155 GND.n3154 0.10956
R5866 GND.n3198 GND.n3197 0.10956
R5867 GND.t186 GND.n3198 0.10956
R5868 GND.t186 GND.n3196 0.10956
R5869 GND.n3196 GND.n3195 0.10956
R5870 GND.n3341 GND.n3340 0.10956
R5871 GND.t1367 GND.n3341 0.10956
R5872 GND.n3347 GND.n3346 0.10956
R5873 GND.t1367 GND.n3347 0.10956
R5874 GND.n3336 GND.n3335 0.10956
R5875 GND.n3335 GND.n3334 0.10956
R5876 GND.n3313 GND.n3312 0.10956
R5877 GND.n3312 GND.n3311 0.10956
R5878 GND.n3355 GND.n3354 0.10956
R5879 GND.t1227 GND.n3355 0.10956
R5880 GND.t1227 GND.n3353 0.10956
R5881 GND.n3353 GND.n3352 0.10956
R5882 GND.n3499 GND.n3498 0.10956
R5883 GND.t664 GND.n3499 0.10956
R5884 GND.n3505 GND.n3504 0.10956
R5885 GND.t664 GND.n3505 0.10956
R5886 GND.n3494 GND.n3493 0.10956
R5887 GND.n3493 GND.n3492 0.10956
R5888 GND.n3471 GND.n3470 0.10956
R5889 GND.n3470 GND.n3469 0.10956
R5890 GND.n3513 GND.n3512 0.10956
R5891 GND.t1338 GND.n3513 0.10956
R5892 GND.t1338 GND.n3511 0.10956
R5893 GND.n3511 GND.n3510 0.10956
R5894 GND.n7289 GND.n7288 0.10956
R5895 GND.t1174 GND.n7289 0.10956
R5896 GND.n7295 GND.n7294 0.10956
R5897 GND.t1174 GND.n7295 0.10956
R5898 GND.n7284 GND.n7283 0.10956
R5899 GND.n7283 GND.n7282 0.10956
R5900 GND.n7261 GND.n7260 0.10956
R5901 GND.n7260 GND.n7259 0.10956
R5902 GND.n7303 GND.n7302 0.10956
R5903 GND.t1240 GND.n7303 0.10956
R5904 GND.t1240 GND.n7301 0.10956
R5905 GND.n7301 GND.n7300 0.10956
R5906 GND.n28 GND.n27 0.10956
R5907 GND.n27 GND.n26 0.10956
R5908 GND.n5 GND.n4 0.10956
R5909 GND.n4 GND.n3 0.10956
R5910 GND.n33 GND.n32 0.10956
R5911 GND.t692 GND.n33 0.10956
R5912 GND.n39 GND.n38 0.10956
R5913 GND.t692 GND.n39 0.10956
R5914 GND.n47 GND.n46 0.10956
R5915 GND.t590 GND.n47 0.10956
R5916 GND.t590 GND.n45 0.10956
R5917 GND.n45 GND.n44 0.10956
R5918 GND.n142 GND.n141 0.10956
R5919 GND.t735 GND.n142 0.10956
R5920 GND.n148 GND.n147 0.10956
R5921 GND.t735 GND.n148 0.10956
R5922 GND.n137 GND.n136 0.10956
R5923 GND.n136 GND.n135 0.10956
R5924 GND.n114 GND.n113 0.10956
R5925 GND.n113 GND.n112 0.10956
R5926 GND.n156 GND.n155 0.10956
R5927 GND.t602 GND.n156 0.10956
R5928 GND.t602 GND.n154 0.10956
R5929 GND.n154 GND.n153 0.10956
R5930 GND.n294 GND.n293 0.10956
R5931 GND.t1118 GND.n294 0.10956
R5932 GND.n300 GND.n299 0.10956
R5933 GND.t1118 GND.n300 0.10956
R5934 GND.n289 GND.n288 0.10956
R5935 GND.n288 GND.n287 0.10956
R5936 GND.n266 GND.n265 0.10956
R5937 GND.n265 GND.n264 0.10956
R5938 GND.n308 GND.n307 0.10956
R5939 GND.t605 GND.n308 0.10956
R5940 GND.t605 GND.n306 0.10956
R5941 GND.n306 GND.n305 0.10956
R5942 GND.n1657 GND.n1656 0.10956
R5943 GND.t363 GND.n1657 0.10956
R5944 GND.n1663 GND.n1662 0.10956
R5945 GND.t363 GND.n1663 0.10956
R5946 GND.n1652 GND.n1651 0.10956
R5947 GND.n1651 GND.n1650 0.10956
R5948 GND.n1629 GND.n1628 0.10956
R5949 GND.n1628 GND.n1627 0.10956
R5950 GND.n1679 GND.n1678 0.10956
R5951 GND.t661 GND.n1679 0.10956
R5952 GND.t661 GND.n1677 0.10956
R5953 GND.n1677 GND.n1676 0.10956
R5954 GND.n2060 GND.t70 0.10956
R5955 GND.n2058 GND.n2057 0.10956
R5956 GND.t70 GND.n2058 0.10956
R5957 GND.n2061 GND.n2060 0.10956
R5958 GND.n3830 GND.n3829 0.10956
R5959 GND.n3831 GND.n3830 0.10956
R5960 GND.n3838 GND.n3837 0.10956
R5961 GND.n3839 GND.n3838 0.10956
R5962 GND.n447 GND.n446 0.10956
R5963 GND.t850 GND.n447 0.10956
R5964 GND.n453 GND.n452 0.10956
R5965 GND.t850 GND.n453 0.10956
R5966 GND.n442 GND.n441 0.10956
R5967 GND.n441 GND.n440 0.10956
R5968 GND.n419 GND.n418 0.10956
R5969 GND.n418 GND.n417 0.10956
R5970 GND.n461 GND.n460 0.10956
R5971 GND.t13 GND.n461 0.10956
R5972 GND.t13 GND.n459 0.10956
R5973 GND.n459 GND.n458 0.10956
R5974 GND.n766 GND.n765 0.10956
R5975 GND.t1281 GND.n766 0.10956
R5976 GND.n772 GND.n771 0.10956
R5977 GND.t1281 GND.n772 0.10956
R5978 GND.n761 GND.n760 0.10956
R5979 GND.n760 GND.n759 0.10956
R5980 GND.n738 GND.n737 0.10956
R5981 GND.n737 GND.n736 0.10956
R5982 GND.n780 GND.n779 0.10956
R5983 GND.t819 GND.n780 0.10956
R5984 GND.t819 GND.n778 0.10956
R5985 GND.n778 GND.n777 0.10956
R5986 GND.n873 GND.n872 0.10956
R5987 GND.t610 GND.n873 0.10956
R5988 GND.n879 GND.n878 0.10956
R5989 GND.t610 GND.n879 0.10956
R5990 GND.n868 GND.n867 0.10956
R5991 GND.n867 GND.n866 0.10956
R5992 GND.n845 GND.n844 0.10956
R5993 GND.n844 GND.n843 0.10956
R5994 GND.n887 GND.n886 0.10956
R5995 GND.t1228 GND.n887 0.10956
R5996 GND.t1228 GND.n885 0.10956
R5997 GND.n885 GND.n884 0.10956
R5998 GND.n7810 GND.n7809 0.10956
R5999 GND.t114 GND.n7810 0.10956
R6000 GND.n7815 GND.n7814 0.10956
R6001 GND.t114 GND.n7815 0.10956
R6002 GND.n7805 GND.n7804 0.10956
R6003 GND.n7804 GND.n7803 0.10956
R6004 GND.n7786 GND.n7785 0.10956
R6005 GND.n7785 GND.n7784 0.10956
R6006 GND.n7567 GND.n7566 0.10956
R6007 GND.n7566 GND.n7565 0.10956
R6008 GND.n7700 GND.n7699 0.10956
R6009 GND.t1141 GND.n7700 0.10956
R6010 GND.n7703 GND.n7702 0.10956
R6011 GND.n7702 GND.n7701 0.10956
R6012 GND.n653 GND.n652 0.10956
R6013 GND.t1232 GND.n653 0.10956
R6014 GND.n656 GND.n655 0.10956
R6015 GND.n655 GND.n654 0.10956
R6016 GND.n6365 GND.n6364 0.10956
R6017 GND.t1183 GND.n6365 0.10956
R6018 GND.n6368 GND.n6367 0.10956
R6019 GND.n6367 GND.n6366 0.10956
R6020 GND.n6201 GND.n6200 0.10956
R6021 GND.t1115 GND.n6201 0.10956
R6022 GND.n6204 GND.n6203 0.10956
R6023 GND.n6203 GND.n6202 0.10956
R6024 GND.n6037 GND.n6036 0.10956
R6025 GND.t18 GND.n6037 0.10956
R6026 GND.n6040 GND.n6039 0.10956
R6027 GND.n6039 GND.n6038 0.10956
R6028 GND.n5854 GND.n5853 0.10956
R6029 GND.t744 GND.n5854 0.10956
R6030 GND.n5857 GND.n5856 0.10956
R6031 GND.n5856 GND.n5855 0.10956
R6032 GND.n5332 GND.n5331 0.10956
R6033 GND.t478 GND.n5332 0.10956
R6034 GND.n5335 GND.n5334 0.10956
R6035 GND.n5334 GND.n5333 0.10956
R6036 GND.n4891 GND.n4890 0.10956
R6037 GND.t1309 GND.n4891 0.10956
R6038 GND.n4894 GND.n4893 0.10956
R6039 GND.n4893 GND.n4892 0.10956
R6040 GND.n7198 GND.n7197 0.10956
R6041 GND.t521 GND.n7198 0.10956
R6042 GND.n7201 GND.n7200 0.10956
R6043 GND.n7200 GND.n7199 0.10956
R6044 GND.n3098 GND.n3097 0.10956
R6045 GND.t828 GND.n3098 0.10956
R6046 GND.n3101 GND.n3100 0.10956
R6047 GND.n3100 GND.n3099 0.10956
R6048 GND.n2774 GND.n2773 0.10956
R6049 GND.t142 GND.n2774 0.10956
R6050 GND.n2777 GND.n2776 0.10956
R6051 GND.n2776 GND.n2775 0.10956
R6052 GND.n2449 GND.n2448 0.10956
R6053 GND.t815 GND.n2449 0.10956
R6054 GND.n2452 GND.n2451 0.10956
R6055 GND.n2451 GND.n2450 0.10956
R6056 GND.n6965 GND.n6964 0.10956
R6057 GND.t804 GND.n6965 0.10956
R6058 GND.n6968 GND.n6967 0.10956
R6059 GND.n6967 GND.n6966 0.10956
R6060 GND.n1800 GND.n1799 0.10956
R6061 GND.t774 GND.n1800 0.10956
R6062 GND.n1803 GND.n1802 0.10956
R6063 GND.n1802 GND.n1801 0.10956
R6064 GND.n1609 GND.n1608 0.10956
R6065 GND.t1344 GND.n1609 0.10956
R6066 GND.n1612 GND.n1611 0.10956
R6067 GND.n1611 GND.n1610 0.10956
R6068 GND.n1545 GND.n1544 0.10956
R6069 GND.t517 GND.n1545 0.10956
R6070 GND.n1199 GND.n1198 0.104537
R6071 GND.n1198 GND.n1197 0.104537
R6072 GND.n2224 GND.n2223 0.104537
R6073 GND.n2223 GND.n2222 0.104537
R6074 GND.n2548 GND.n2547 0.104537
R6075 GND.n2547 GND.n2546 0.104537
R6076 GND.n2873 GND.n2872 0.104537
R6077 GND.n2872 GND.n2871 0.104537
R6078 GND.n3170 GND.n3169 0.104537
R6079 GND.n3169 GND.n3168 0.104537
R6080 GND.n3327 GND.n3326 0.104537
R6081 GND.n3326 GND.n3325 0.104537
R6082 GND.n3485 GND.n3484 0.104537
R6083 GND.n3484 GND.n3483 0.104537
R6084 GND.n7275 GND.n7274 0.104537
R6085 GND.n7274 GND.n7273 0.104537
R6086 GND.n19 GND.n18 0.104537
R6087 GND.n18 GND.n17 0.104537
R6088 GND.n128 GND.n127 0.104537
R6089 GND.n127 GND.n126 0.104537
R6090 GND.n280 GND.n279 0.104537
R6091 GND.n279 GND.n278 0.104537
R6092 GND.n1643 GND.n1642 0.104537
R6093 GND.n1642 GND.n1641 0.104537
R6094 GND.n433 GND.n432 0.104537
R6095 GND.n432 GND.n431 0.104537
R6096 GND.n752 GND.n751 0.104537
R6097 GND.n751 GND.n750 0.104537
R6098 GND.n859 GND.n858 0.104537
R6099 GND.n858 GND.n857 0.104537
R6100 GND.n7798 GND.n7797 0.104537
R6101 GND.n7797 GND.n7796 0.104537
R6102 GND.n4395 GND.n4374 0.102336
R6103 GND.n5918 GND.n5464 0.102336
R6104 GND.n1945 GND.n1560 0.102333
R6105 GND.n1750 GND.n1749 0.102333
R6106 GND.n7022 GND.n7021 0.102333
R6107 GND.n2399 GND.n2398 0.102333
R6108 GND.n2724 GND.n2723 0.102333
R6109 GND.n3048 GND.n3047 0.102333
R6110 GND.n7148 GND.n7147 0.102333
R6111 GND.n4841 GND.n4840 0.102333
R6112 GND.n5417 GND.n5416 0.102333
R6113 GND.n5912 GND.n5911 0.102333
R6114 GND.n5987 GND.n5986 0.102333
R6115 GND.n6154 GND.n6153 0.102333
R6116 GND.n6318 GND.n6317 0.102333
R6117 GND.n606 GND.n605 0.102333
R6118 GND.n7649 GND.n7648 0.102333
R6119 GND.n7529 GND.n7528 0.102333
R6120 GND.n6779 GND 0.101889
R6121 GND.n4357 GND 0.101889
R6122 GND GND.n3648 0.0991625
R6123 GND.n5475 GND.n5474 0.0963333
R6124 GND.n5476 GND.n5467 0.0963333
R6125 GND.n5482 GND.n5467 0.0963333
R6126 GND.n5483 GND.n5482 0.0963333
R6127 GND.n5484 GND.n5483 0.0963333
R6128 GND.n4406 GND.n4405 0.0963333
R6129 GND.n4407 GND.n4398 0.0963333
R6130 GND.n4413 GND.n4398 0.0963333
R6131 GND.n4414 GND.n4413 0.0963333
R6132 GND.n4415 GND.n4414 0.0963333
R6133 GND.n3836 GND.n3835 0.0944005
R6134 GND.n7582 GND.n7581 0.0944005
R6135 GND.n7583 GND.n7582 0.0944005
R6136 GND.n7525 GND.n7524 0.0944005
R6137 GND.n7746 GND.n7745 0.0944005
R6138 GND.n7747 GND.n7746 0.0944005
R6139 GND.n7645 GND.n7644 0.0944005
R6140 GND.n699 GND.n698 0.0944005
R6141 GND.n700 GND.n699 0.0944005
R6142 GND.n602 GND.n601 0.0944005
R6143 GND.n6414 GND.n6413 0.0944005
R6144 GND.n6415 GND.n6414 0.0944005
R6145 GND.n6314 GND.n6313 0.0944005
R6146 GND.n6250 GND.n6249 0.0944005
R6147 GND.n6251 GND.n6250 0.0944005
R6148 GND.n6150 GND.n6149 0.0944005
R6149 GND.n6086 GND.n6085 0.0944005
R6150 GND.n6087 GND.n6086 0.0944005
R6151 GND.n5983 GND.n5982 0.0944005
R6152 GND.n5898 GND.n5897 0.0944005
R6153 GND.n5897 GND.n5896 0.0944005
R6154 GND.n5908 GND.n5907 0.0944005
R6155 GND.n5376 GND.n5375 0.0944005
R6156 GND.n5375 GND.n5374 0.0944005
R6157 GND.n5413 GND.n5412 0.0944005
R6158 GND.n4910 GND.n4909 0.0944005
R6159 GND.n4911 GND.n4910 0.0944005
R6160 GND.n4837 GND.n4836 0.0944005
R6161 GND.n7217 GND.n7216 0.0944005
R6162 GND.n7218 GND.n7217 0.0944005
R6163 GND.n7144 GND.n7143 0.0944005
R6164 GND.n3117 GND.n3116 0.0944005
R6165 GND.n3118 GND.n3117 0.0944005
R6166 GND.n3044 GND.n3043 0.0944005
R6167 GND.n2820 GND.n2819 0.0944005
R6168 GND.n2821 GND.n2820 0.0944005
R6169 GND.n2720 GND.n2719 0.0944005
R6170 GND.n2495 GND.n2494 0.0944005
R6171 GND.n2496 GND.n2495 0.0944005
R6172 GND.n2395 GND.n2394 0.0944005
R6173 GND.n7008 GND.n7007 0.0944005
R6174 GND.n7007 GND.n6878 0.0944005
R6175 GND.n7018 GND.n7017 0.0944005
R6176 GND.n1846 GND.n1845 0.0944005
R6177 GND.n1847 GND.n1846 0.0944005
R6178 GND.n1746 GND.n1745 0.0944005
R6179 GND.n1889 GND.n1888 0.0944005
R6180 GND.n1890 GND.n1889 0.0944005
R6181 GND.n1557 GND.n1556 0.0944005
R6182 GND.n1556 GND.n1555 0.0944005
R6183 GND.n1925 GND.n1923 0.0921667
R6184 GND.n1692 GND.n1690 0.0921667
R6185 GND.n6900 GND.n6898 0.0921667
R6186 GND.n2368 GND.n2366 0.0921667
R6187 GND.n2693 GND.n2691 0.0921667
R6188 GND.n3017 GND.n3015 0.0921667
R6189 GND.n7090 GND.n7088 0.0921667
R6190 GND.n4785 GND.n4783 0.0921667
R6191 GND.n5267 GND.n5265 0.0921667
R6192 GND.n5789 GND.n5787 0.0921667
R6193 GND.n5956 GND.n5954 0.0921667
R6194 GND.n6123 GND.n6121 0.0921667
R6195 GND.n6287 GND.n6285 0.0921667
R6196 GND.n575 GND.n573 0.0921667
R6197 GND.n7618 GND.n7616 0.0921667
R6198 GND.n7498 GND.n7496 0.0921667
R6199 GND.n4040 GND.n4038 0.0920099
R6200 GND.n5514 GND.n5512 0.0894537
R6201 GND.n4439 GND.n4437 0.0894537
R6202 GND.n6423 GND.n6421 0.0894537
R6203 GND.n2084 GND 0.0891586
R6204 GND.n1911 GND.n1909 0.0891364
R6205 GND.n1868 GND.n1866 0.0891364
R6206 GND.n6889 GND.n6887 0.0891364
R6207 GND.n2517 GND.n2515 0.0891364
R6208 GND.n2842 GND.n2840 0.0891364
R6209 GND.n3139 GND.n3137 0.0891364
R6210 GND.n7239 GND.n7237 0.0891364
R6211 GND.n4771 GND.n4769 0.0891364
R6212 GND.n5256 GND.n5254 0.0891364
R6213 GND.n5939 GND.n5937 0.0891364
R6214 GND.n6108 GND.n6106 0.0891364
R6215 GND.n6272 GND.n6270 0.0891364
R6216 GND.n6581 GND.n6579 0.0891364
R6217 GND.n721 GND.n719 0.0891364
R6218 GND.n7768 GND.n7766 0.0891364
R6219 GND.n7603 GND.n7601 0.0891364
R6220 GND.n7438 GND.n7367 0.08745
R6221 GND.n2020 GND.n2019 0.08745
R6222 GND.n518 GND.n517 0.08745
R6223 GND.n213 GND.n212 0.08745
R6224 GND.n1512 GND.n1511 0.08745
R6225 GND.n1464 GND.n1463 0.08745
R6226 GND.n4221 GND.n4220 0.08745
R6227 GND.n3415 GND.n3414 0.08745
R6228 GND.n3258 GND.n3257 0.08745
R6229 GND.n2961 GND.n2960 0.08745
R6230 GND.n2636 GND.n2635 0.08745
R6231 GND.n2312 GND.n2311 0.08745
R6232 GND.n2150 GND.n2149 0.08745
R6233 GND.n1282 GND.n1281 0.08745
R6234 GND.n365 GND.n364 0.08745
R6235 GND.n7413 GND.n7412 0.08745
R6236 GND.n7438 GND.n7437 0.0868625
R6237 GND.n2020 GND.n1996 0.0868625
R6238 GND.n365 GND.n320 0.0868625
R6239 GND.n518 GND.n473 0.0868625
R6240 GND.n213 GND.n168 0.0868625
R6241 GND.n1514 GND.n1512 0.0868625
R6242 GND.n1466 GND.n1464 0.0868625
R6243 GND.n4221 GND.n4176 0.0868625
R6244 GND.n3415 GND.n3370 0.0868625
R6245 GND.n3258 GND.n3213 0.0868625
R6246 GND.n2961 GND.n2916 0.0868625
R6247 GND.n2636 GND.n2591 0.0868625
R6248 GND.n2312 GND.n2267 0.0868625
R6249 GND.n2150 GND.n2105 0.0868625
R6250 GND.n1282 GND.n1237 0.0868625
R6251 GND.n7415 GND.n7413 0.0868625
R6252 GND.n3666 GND.n3664 0.0853214
R6253 GND.n1920 GND.n1883 0.0845572
R6254 GND.n1878 GND.n1877 0.0845572
R6255 GND.n7029 GND.n7028 0.0845572
R6256 GND.n2527 GND.n2526 0.0845572
R6257 GND.n2852 GND.n2851 0.0845572
R6258 GND.n3149 GND.n3148 0.0845572
R6259 GND.n7249 GND.n7248 0.0845572
R6260 GND.n4780 GND.n4271 0.0845572
R6261 GND.n5421 GND.n4270 0.0845572
R6262 GND.n5949 GND.n5948 0.0845572
R6263 GND.n6118 GND.n6117 0.0845572
R6264 GND.n6282 GND.n6281 0.0845572
R6265 GND.n6591 GND.n6590 0.0845572
R6266 GND.n731 GND.n730 0.0845572
R6267 GND.n7778 GND.n7777 0.0845572
R6268 GND.n7613 GND.n7612 0.0845572
R6269 GND.n3967 GND.n3954 0.0838333
R6270 GND.n5437 GND 0.0824444
R6271 GND.n4339 GND 0.0824444
R6272 GND.n5040 GND.n4272 0.0795145
R6273 GND.n1931 GND 0.0775833
R6274 GND.n1698 GND 0.0775833
R6275 GND.n6906 GND 0.0775833
R6276 GND.n2374 GND 0.0775833
R6277 GND.n2699 GND 0.0775833
R6278 GND.n3023 GND 0.0775833
R6279 GND.n7096 GND 0.0775833
R6280 GND.n4791 GND 0.0775833
R6281 GND.n5273 GND 0.0775833
R6282 GND.n5795 GND 0.0775833
R6283 GND.n5962 GND 0.0775833
R6284 GND.n6129 GND 0.0775833
R6285 GND.n6293 GND 0.0775833
R6286 GND.n581 GND 0.0775833
R6287 GND.n7624 GND 0.0775833
R6288 GND.n7504 GND 0.0775833
R6289 GND.n6868 GND.n6843 0.0740087
R6290 GND.n6761 GND.n5463 0.0740087
R6291 GND.n6869 GND.n6868 0.0732412
R6292 GND.n5463 GND.n5438 0.0732412
R6293 GND.n6870 GND.n6869 0.0727407
R6294 GND.n5438 GND.n4423 0.0727407
R6295 GND.n3855 GND.n3853 0.0727222
R6296 GND.n6840 GND.n4423 0.0714246
R6297 GND.n6600 GND.n6599 0.0711855
R6298 GND.n6839 GND.n6805 0.0696598
R6299 GND.n7084 GND.n7050 0.0696598
R6300 GND.n6843 GND.n6842 0.0692593
R6301 GND.n6761 GND.n6760 0.0692593
R6302 GND.n3869 GND.n3855 0.06925
R6303 GND.n1896 GND 0.0675455
R6304 GND.n1853 GND 0.0675455
R6305 GND GND.n7040 0.0675455
R6306 GND.n2502 GND 0.0675455
R6307 GND.n2827 GND 0.0675455
R6308 GND.n3124 GND 0.0675455
R6309 GND.n7224 GND 0.0675455
R6310 GND.n4756 GND 0.0675455
R6311 GND GND.n5432 0.0675455
R6312 GND.n5924 GND 0.0675455
R6313 GND.n6093 GND 0.0675455
R6314 GND.n6257 GND 0.0675455
R6315 GND.n6566 GND 0.0675455
R6316 GND.n706 GND 0.0675455
R6317 GND.n7753 GND 0.0675455
R6318 GND.n7588 GND 0.0675455
R6319 GND.n7321 GND.n4169 0.0666615
R6320 GND.n6746 GND.n6741 0.0659695
R6321 GND.n4385 GND.n4380 0.0659695
R6322 GND.n4077 GND.n4076 0.0653227
R6323 GND.n4970 GND.n4969 0.0643889
R6324 GND.n4969 GND.n4967 0.0643889
R6325 GND.n4967 GND.n4964 0.0643889
R6326 GND.n4964 GND.n4962 0.0643889
R6327 GND.n6746 GND.n6738 0.0643889
R6328 GND.n6750 GND.n6738 0.0643889
R6329 GND.n6751 GND.n6750 0.0643889
R6330 GND.n6777 GND.n6770 0.0643889
R6331 GND.n6783 GND.n6768 0.0643889
R6332 GND.n6783 GND.n6765 0.0643889
R6333 GND.n6787 GND.n6765 0.0643889
R6334 GND.n6788 GND.n6787 0.0643889
R6335 GND.n5231 GND.n5226 0.0643889
R6336 GND.n5242 GND.n5224 0.0643889
R6337 GND.n5243 GND.n5242 0.0643889
R6338 GND.n4385 GND.n4377 0.0643889
R6339 GND.n4389 GND.n4377 0.0643889
R6340 GND.n4390 GND.n4389 0.0643889
R6341 GND.n4355 GND.n4348 0.0643889
R6342 GND.n4361 GND.n4346 0.0643889
R6343 GND.n4361 GND.n4343 0.0643889
R6344 GND.n4365 GND.n4343 0.0643889
R6345 GND.n4366 GND.n4365 0.0643889
R6346 GND.n4323 GND.n4318 0.0643889
R6347 GND.n4334 GND.n4316 0.0643889
R6348 GND.n4335 GND.n4334 0.0643889
R6349 GND.n7449 GND.n7448 0.0636886
R6350 GND.n7450 GND.n7449 0.0636886
R6351 GND.n7452 GND.n7451 0.0636886
R6352 GND.n7451 GND.n7450 0.0636886
R6353 GND.n529 GND.n528 0.0636886
R6354 GND.n530 GND.n529 0.0636886
R6355 GND.n532 GND.n531 0.0636886
R6356 GND.n531 GND.n530 0.0636886
R6357 GND.n224 GND.n223 0.0636886
R6358 GND.n225 GND.n224 0.0636886
R6359 GND.n227 GND.n226 0.0636886
R6360 GND.n226 GND.n225 0.0636886
R6361 GND.n4232 GND.n4231 0.0636886
R6362 GND.n4233 GND.n4232 0.0636886
R6363 GND.n4235 GND.n4234 0.0636886
R6364 GND.n4234 GND.n4233 0.0636886
R6365 GND.n3269 GND.n3268 0.0636886
R6366 GND.n3270 GND.n3269 0.0636886
R6367 GND.n3272 GND.n3271 0.0636886
R6368 GND.n3271 GND.n3270 0.0636886
R6369 GND.n2647 GND.n2646 0.0636886
R6370 GND.n2648 GND.n2647 0.0636886
R6371 GND.n2650 GND.n2649 0.0636886
R6372 GND.n2649 GND.n2648 0.0636886
R6373 GND.n2161 GND.n2160 0.0636886
R6374 GND.n2162 GND.n2161 0.0636886
R6375 GND.n2164 GND.n2163 0.0636886
R6376 GND.n2163 GND.n2162 0.0636886
R6377 GND.n1293 GND.n1292 0.0636886
R6378 GND.n1294 GND.n1293 0.0636886
R6379 GND.n1296 GND.n1295 0.0636886
R6380 GND.n1295 GND.n1294 0.0636886
R6381 GND.n1271 GND.t597 0.0636886
R6382 GND.n1272 GND.n1271 0.0636886
R6383 GND.n1270 GND.n1269 0.0636886
R6384 GND.t597 GND.n1270 0.0636886
R6385 GND.n2140 GND.n2139 0.0636886
R6386 GND.n2139 GND.t733 0.0636886
R6387 GND.t733 GND.n2138 0.0636886
R6388 GND.n2138 GND.n2137 0.0636886
R6389 GND.n2323 GND.n2322 0.0636886
R6390 GND.n2324 GND.n2323 0.0636886
R6391 GND.n2326 GND.n2325 0.0636886
R6392 GND.n2325 GND.n2324 0.0636886
R6393 GND.n2302 GND.n2301 0.0636886
R6394 GND.n2301 GND.t587 0.0636886
R6395 GND.t587 GND.n2300 0.0636886
R6396 GND.n2300 GND.n2299 0.0636886
R6397 GND.n2626 GND.n2625 0.0636886
R6398 GND.n2625 GND.t595 0.0636886
R6399 GND.t595 GND.n2624 0.0636886
R6400 GND.n2624 GND.n2623 0.0636886
R6401 GND.n2972 GND.n2971 0.0636886
R6402 GND.n2973 GND.n2972 0.0636886
R6403 GND.n2975 GND.n2974 0.0636886
R6404 GND.n2974 GND.n2973 0.0636886
R6405 GND.n2951 GND.n2950 0.0636886
R6406 GND.n2950 GND.t594 0.0636886
R6407 GND.t594 GND.n2949 0.0636886
R6408 GND.n2949 GND.n2948 0.0636886
R6409 GND.n3248 GND.n3247 0.0636886
R6410 GND.n3247 GND.t1158 0.0636886
R6411 GND.t1158 GND.n3246 0.0636886
R6412 GND.n3246 GND.n3245 0.0636886
R6413 GND.n3426 GND.n3425 0.0636886
R6414 GND.n3427 GND.n3426 0.0636886
R6415 GND.n3429 GND.n3428 0.0636886
R6416 GND.n3428 GND.n3427 0.0636886
R6417 GND.n3405 GND.n3404 0.0636886
R6418 GND.n3404 GND.t1161 0.0636886
R6419 GND.t1161 GND.n3403 0.0636886
R6420 GND.n3403 GND.n3402 0.0636886
R6421 GND.n4211 GND.n4210 0.0636886
R6422 GND.n4210 GND.t837 0.0636886
R6423 GND.t837 GND.n4209 0.0636886
R6424 GND.n4209 GND.n4208 0.0636886
R6425 GND.n1398 GND.n1397 0.0636886
R6426 GND.n1399 GND.n1398 0.0636886
R6427 GND.n1401 GND.n1400 0.0636886
R6428 GND.n1400 GND.n1399 0.0636886
R6429 GND.n1454 GND.n1453 0.0636886
R6430 GND.n1453 GND.t732 0.0636886
R6431 GND.n1452 GND.n1451 0.0636886
R6432 GND.t732 GND.n1452 0.0636886
R6433 GND.n61 GND.n60 0.0636886
R6434 GND.n66 GND.n65 0.0636886
R6435 GND.n1502 GND.n1501 0.0636886
R6436 GND.n1501 GND.t399 0.0636886
R6437 GND.t399 GND.n1500 0.0636886
R6438 GND.n1500 GND.n1499 0.0636886
R6439 GND.n203 GND.n202 0.0636886
R6440 GND.n202 GND.t435 0.0636886
R6441 GND.t435 GND.n201 0.0636886
R6442 GND.n201 GND.n200 0.0636886
R6443 GND.n376 GND.n375 0.0636886
R6444 GND.n377 GND.n376 0.0636886
R6445 GND.n379 GND.n378 0.0636886
R6446 GND.n378 GND.n377 0.0636886
R6447 GND.n2010 GND.n2009 0.0636886
R6448 GND.n2009 GND.t596 0.0636886
R6449 GND.t596 GND.n2008 0.0636886
R6450 GND.n2008 GND.n2007 0.0636886
R6451 GND.n1994 GND.n1993 0.0636886
R6452 GND.n1993 GND.t687 0.0636886
R6453 GND.n2036 GND.n2035 0.0636886
R6454 GND.n2037 GND.n2036 0.0636886
R6455 GND.n2039 GND.n2038 0.0636886
R6456 GND.n2038 GND.n2037 0.0636886
R6457 GND.n1349 GND.n1348 0.0636886
R6458 GND.n1350 GND.n1349 0.0636886
R6459 GND.n1344 GND.n1343 0.0636886
R6460 GND.n1350 GND.n1344 0.0636886
R6461 GND.n1354 GND.n1353 0.0636886
R6462 GND.t384 GND.n1354 0.0636886
R6463 GND.n1334 GND.n1333 0.0636886
R6464 GND.n1350 GND.n1334 0.0636886
R6465 GND.n1339 GND.n1338 0.0636886
R6466 GND.n1350 GND.n1339 0.0636886
R6467 GND.n1352 GND.n1351 0.0636886
R6468 GND.t384 GND.n1352 0.0636886
R6469 GND.n903 GND.n902 0.0636886
R6470 GND.n1044 GND.n903 0.0636886
R6471 GND.n908 GND.n907 0.0636886
R6472 GND.n1044 GND.n908 0.0636886
R6473 GND.n1072 GND.n1071 0.0636886
R6474 GND.t36 GND.n1072 0.0636886
R6475 GND.n918 GND.n917 0.0636886
R6476 GND.n1044 GND.n918 0.0636886
R6477 GND.n912 GND.n911 0.0636886
R6478 GND.n1044 GND.n912 0.0636886
R6479 GND.n1070 GND.n1069 0.0636886
R6480 GND.t36 GND.n1070 0.0636886
R6481 GND.n928 GND.n927 0.0636886
R6482 GND.n1044 GND.n928 0.0636886
R6483 GND.n923 GND.n922 0.0636886
R6484 GND.n1044 GND.n923 0.0636886
R6485 GND.n1068 GND.n1067 0.0636886
R6486 GND.t36 GND.n1068 0.0636886
R6487 GND.n938 GND.n937 0.0636886
R6488 GND.n1044 GND.n938 0.0636886
R6489 GND.n934 GND.n933 0.0636886
R6490 GND.n1044 GND.n934 0.0636886
R6491 GND.n1066 GND.n1065 0.0636886
R6492 GND.t36 GND.n1066 0.0636886
R6493 GND.n948 GND.n947 0.0636886
R6494 GND.n1044 GND.n948 0.0636886
R6495 GND.n943 GND.n942 0.0636886
R6496 GND.n1044 GND.n943 0.0636886
R6497 GND.n1064 GND.n1063 0.0636886
R6498 GND.t36 GND.n1064 0.0636886
R6499 GND.n958 GND.n957 0.0636886
R6500 GND.n1044 GND.n958 0.0636886
R6501 GND.n953 GND.n952 0.0636886
R6502 GND.n1044 GND.n953 0.0636886
R6503 GND.n1062 GND.n1061 0.0636886
R6504 GND.t36 GND.n1062 0.0636886
R6505 GND.n968 GND.n967 0.0636886
R6506 GND.n1044 GND.n968 0.0636886
R6507 GND.n964 GND.n963 0.0636886
R6508 GND.n1044 GND.n964 0.0636886
R6509 GND.n1060 GND.n1059 0.0636886
R6510 GND.t36 GND.n1060 0.0636886
R6511 GND.n973 GND.n972 0.0636886
R6512 GND.n1044 GND.n973 0.0636886
R6513 GND.n978 GND.n977 0.0636886
R6514 GND.n1044 GND.n978 0.0636886
R6515 GND.n1058 GND.n1057 0.0636886
R6516 GND.t36 GND.n1058 0.0636886
R6517 GND.n987 GND.n986 0.0636886
R6518 GND.n1044 GND.n987 0.0636886
R6519 GND.n993 GND.n992 0.0636886
R6520 GND.n1044 GND.n993 0.0636886
R6521 GND.n1056 GND.n1055 0.0636886
R6522 GND.t36 GND.n1056 0.0636886
R6523 GND.n1003 GND.n1002 0.0636886
R6524 GND.n1044 GND.n1003 0.0636886
R6525 GND.n998 GND.n997 0.0636886
R6526 GND.n1044 GND.n998 0.0636886
R6527 GND.n1054 GND.n1053 0.0636886
R6528 GND.t36 GND.n1054 0.0636886
R6529 GND.n1013 GND.n1012 0.0636886
R6530 GND.n1044 GND.n1013 0.0636886
R6531 GND.n1009 GND.n1008 0.0636886
R6532 GND.n1044 GND.n1009 0.0636886
R6533 GND.n1052 GND.n1051 0.0636886
R6534 GND.t36 GND.n1052 0.0636886
R6535 GND.n1023 GND.n1022 0.0636886
R6536 GND.n1044 GND.n1023 0.0636886
R6537 GND.n1019 GND.n1018 0.0636886
R6538 GND.n1044 GND.n1019 0.0636886
R6539 GND.n1050 GND.n1049 0.0636886
R6540 GND.t36 GND.n1050 0.0636886
R6541 GND.n1038 GND.n1037 0.0636886
R6542 GND.n1044 GND.n1038 0.0636886
R6543 GND.n1034 GND.n1033 0.0636886
R6544 GND.n1044 GND.n1034 0.0636886
R6545 GND.n1046 GND.n1045 0.0636886
R6546 GND.t36 GND.n1046 0.0636886
R6547 GND.n1043 GND.n1042 0.0636886
R6548 GND.n1044 GND.n1043 0.0636886
R6549 GND.n1048 GND.n1047 0.0636886
R6550 GND.t36 GND.n1048 0.0636886
R6551 GND.n1044 GND.n1028 0.0636886
R6552 GND.n1028 GND.n1027 0.0636886
R6553 GND.n355 GND.n354 0.0636886
R6554 GND.n354 GND.t160 0.0636886
R6555 GND.t160 GND.n353 0.0636886
R6556 GND.n353 GND.n352 0.0636886
R6557 GND.n508 GND.n507 0.0636886
R6558 GND.n507 GND.t161 0.0636886
R6559 GND.t161 GND.n506 0.0636886
R6560 GND.n506 GND.n505 0.0636886
R6561 GND.n801 GND.n800 0.0636886
R6562 GND.n802 GND.n801 0.0636886
R6563 GND.n804 GND.n803 0.0636886
R6564 GND.n803 GND.n802 0.0636886
R6565 GND.n7402 GND.t593 0.0636886
R6566 GND.n7403 GND.n7402 0.0636886
R6567 GND.n7401 GND.n7400 0.0636886
R6568 GND.t593 GND.n7401 0.0636886
R6569 GND.n7357 GND.n7356 0.0636886
R6570 GND.n7356 GND.t684 0.0636886
R6571 GND.n4394 GND.n4393 0.0636834
R6572 GND.n6755 GND.n6754 0.0636834
R6573 GND.n6842 GND 0.0628765
R6574 GND.n6760 GND 0.0628765
R6575 GND.n5192 GND.n5188 0.0610263
R6576 GND.n5196 GND.n5188 0.0610263
R6577 GND.n5197 GND.n5196 0.0610263
R6578 GND.n5198 GND.n5197 0.0610263
R6579 GND.n5209 GND.n5185 0.0610263
R6580 GND.n5209 GND.n5182 0.0610263
R6581 GND.n5182 GND.n5179 0.0610263
R6582 GND.n5214 GND.n5179 0.0610263
R6583 GND.n4289 GND.n4285 0.0610263
R6584 GND.n4293 GND.n4285 0.0610263
R6585 GND.n4294 GND.n4293 0.0610263
R6586 GND.n4295 GND.n4294 0.0610263
R6587 GND.n4306 GND.n4282 0.0610263
R6588 GND.n4306 GND.n4279 0.0610263
R6589 GND.n4279 GND.n4276 0.0610263
R6590 GND.n4311 GND.n4276 0.0610263
R6591 GND.n1883 GND 0.060284
R6592 GND.n1878 GND 0.060284
R6593 GND.n7028 GND 0.060284
R6594 GND.n2527 GND 0.060284
R6595 GND.n2852 GND 0.060284
R6596 GND.n3149 GND 0.060284
R6597 GND.n7249 GND 0.060284
R6598 GND.n4271 GND 0.060284
R6599 GND.n4270 GND 0.060284
R6600 GND.n5949 GND 0.060284
R6601 GND.n6118 GND 0.060284
R6602 GND.n6282 GND 0.060284
R6603 GND.n6591 GND 0.060284
R6604 GND.n731 GND 0.060284
R6605 GND.n7778 GND 0.060284
R6606 GND.n7613 GND 0.060284
R6607 GND.n6870 GND.n4272 0.0593951
R6608 GND.n4044 GND.n4042 0.0589677
R6609 GND.n7365 GND.n7364 0.0588369
R6610 GND.n2017 GND.n2016 0.0588344
R6611 GND.n515 GND.n514 0.0588344
R6612 GND.n210 GND.n209 0.0588344
R6613 GND.n1509 GND.n1508 0.0588344
R6614 GND.n1461 GND.n1460 0.0588344
R6615 GND.n4218 GND.n4217 0.0588344
R6616 GND.n3412 GND.n3411 0.0588344
R6617 GND.n3255 GND.n3254 0.0588344
R6618 GND.n2958 GND.n2957 0.0588344
R6619 GND.n2633 GND.n2632 0.0588344
R6620 GND.n2309 GND.n2308 0.0588344
R6621 GND.n2147 GND.n2146 0.0588344
R6622 GND.n1279 GND.n1278 0.0588344
R6623 GND.n362 GND.n361 0.0588344
R6624 GND.n7410 GND.n7409 0.0588344
R6625 GND.n1940 GND.n1928 0.0582982
R6626 GND.n1707 GND.n1695 0.0582982
R6627 GND.n6915 GND.n6903 0.0582982
R6628 GND.n2383 GND.n2371 0.0582982
R6629 GND.n2708 GND.n2696 0.0582982
R6630 GND.n3032 GND.n3020 0.0582982
R6631 GND.n7105 GND.n7093 0.0582982
R6632 GND.n4800 GND.n4788 0.0582982
R6633 GND.n5282 GND.n5270 0.0582982
R6634 GND.n5804 GND.n5792 0.0582982
R6635 GND.n5971 GND.n5959 0.0582982
R6636 GND.n6138 GND.n6126 0.0582982
R6637 GND.n6302 GND.n6290 0.0582982
R6638 GND.n590 GND.n578 0.0582982
R6639 GND.n7633 GND.n7621 0.0582982
R6640 GND.n7513 GND.n7501 0.0582982
R6641 GND.n3954 GND.n3952 0.0581389
R6642 GND.n5453 GND.n5452 0.0580634
R6643 GND.n6858 GND.n6857 0.0580634
R6644 GND.n6753 GND.n6736 0.0580441
R6645 GND.n6790 GND.n6763 0.0580441
R6646 GND.n5239 GND.n5238 0.0580441
R6647 GND.n5245 GND.n5222 0.0580441
R6648 GND.n4392 GND.n4375 0.0580441
R6649 GND.n4368 GND.n4341 0.0580441
R6650 GND.n4331 GND.n4330 0.0580441
R6651 GND.n4337 GND.n4314 0.0580441
R6652 GND.n6832 GND 0.058
R6653 GND.n6826 GND 0.058
R6654 GND.n6814 GND 0.058
R6655 GND.n7077 GND 0.058
R6656 GND.n7071 GND 0.058
R6657 GND.n7059 GND 0.058
R6658 GND.n3637 GND.n3634 0.0570476
R6659 GND.n1902 GND.n1901 0.05675
R6660 GND.n1859 GND.n1858 0.05675
R6661 GND.n7035 GND.n7034 0.05675
R6662 GND.n2508 GND.n2507 0.05675
R6663 GND.n2833 GND.n2832 0.05675
R6664 GND.n3130 GND.n3129 0.05675
R6665 GND.n7230 GND.n7229 0.05675
R6666 GND.n4762 GND.n4761 0.05675
R6667 GND.n5427 GND.n5426 0.05675
R6668 GND.n5930 GND.n5929 0.05675
R6669 GND.n6099 GND.n6098 0.05675
R6670 GND.n6263 GND.n6262 0.05675
R6671 GND.n6572 GND.n6571 0.05675
R6672 GND.n712 GND.n711 0.05675
R6673 GND.n7759 GND.n7758 0.05675
R6674 GND.n7594 GND.n7593 0.05675
R6675 GND.n5456 GND.n5447 0.05675
R6676 GND.n5457 GND.n5445 0.05675
R6677 GND.n6861 GND.n6852 0.05675
R6678 GND.n6862 GND.n6850 0.05675
R6679 GND.n6779 GND.n6778 0.0567153
R6680 GND.n4357 GND.n4356 0.0567153
R6681 GND.n6839 GND.n6838 0.0558279
R6682 GND.n7084 GND.n7083 0.0558279
R6683 GND.n6820 GND 0.0555
R6684 GND.n7065 GND 0.0555
R6685 GND.n3692 GND.n3691 0.0540714
R6686 GND.n1915 GND.n1914 0.0532741
R6687 GND.n1872 GND.n1871 0.0532741
R6688 GND.n6893 GND.n6892 0.0532741
R6689 GND.n2521 GND.n2520 0.0532741
R6690 GND.n2846 GND.n2845 0.0532741
R6691 GND.n3143 GND.n3142 0.0532741
R6692 GND.n7243 GND.n7242 0.0532741
R6693 GND.n4775 GND.n4774 0.0532741
R6694 GND.n5260 GND.n5259 0.0532741
R6695 GND.n5943 GND.n5942 0.0532741
R6696 GND.n6112 GND.n6111 0.0532741
R6697 GND.n6276 GND.n6275 0.0532741
R6698 GND.n6585 GND.n6584 0.0532741
R6699 GND.n725 GND.n724 0.0532741
R6700 GND.n7772 GND.n7771 0.0532741
R6701 GND.n7607 GND.n7606 0.0532741
R6702 GND.n3633 GND.n3630 0.0530794
R6703 GND.n5202 GND.n5201 0.052907
R6704 GND.n4299 GND.n4298 0.052907
R6705 GND.n1359 GND.n1356 0.0528195
R6706 GND.n1077 GND.n1074 0.0528195
R6707 GND.n1909 GND 0.0527727
R6708 GND.n1866 GND 0.0527727
R6709 GND.n6887 GND 0.0527727
R6710 GND.n2515 GND 0.0527727
R6711 GND.n2840 GND 0.0527727
R6712 GND.n3137 GND 0.0527727
R6713 GND.n7237 GND 0.0527727
R6714 GND.n4769 GND 0.0527727
R6715 GND.n5254 GND 0.0527727
R6716 GND.n5937 GND 0.0527727
R6717 GND.n6106 GND 0.0527727
R6718 GND.n6270 GND 0.0527727
R6719 GND.n6579 GND 0.0527727
R6720 GND.n719 GND 0.0527727
R6721 GND.n7766 GND 0.0527727
R6722 GND.n7601 GND 0.0527727
R6723 GND.n1187 GND.n1186 0.0525185
R6724 GND.n1188 GND.n1187 0.0525185
R6725 GND.n1202 GND.n1201 0.0525185
R6726 GND.n1203 GND.n1202 0.0525185
R6727 GND.n1196 GND.n1195 0.0525185
R6728 GND.n1197 GND.n1196 0.0525185
R6729 GND.n1190 GND.n1189 0.0525185
R6730 GND.n1191 GND.n1190 0.0525185
R6731 GND.n1205 GND.n1204 0.0525185
R6732 GND.n1206 GND.n1205 0.0525185
R6733 GND.n2212 GND.n2211 0.0525185
R6734 GND.n2213 GND.n2212 0.0525185
R6735 GND.n2227 GND.n2226 0.0525185
R6736 GND.n2228 GND.n2227 0.0525185
R6737 GND.n2221 GND.n2220 0.0525185
R6738 GND.n2222 GND.n2221 0.0525185
R6739 GND.n2215 GND.n2214 0.0525185
R6740 GND.n2216 GND.n2215 0.0525185
R6741 GND.n2230 GND.n2229 0.0525185
R6742 GND.n2231 GND.n2230 0.0525185
R6743 GND.n2536 GND.n2535 0.0525185
R6744 GND.n2537 GND.n2536 0.0525185
R6745 GND.n2551 GND.n2550 0.0525185
R6746 GND.n2552 GND.n2551 0.0525185
R6747 GND.n2545 GND.n2544 0.0525185
R6748 GND.n2546 GND.n2545 0.0525185
R6749 GND.n2539 GND.n2538 0.0525185
R6750 GND.n2540 GND.n2539 0.0525185
R6751 GND.n2554 GND.n2553 0.0525185
R6752 GND.n2555 GND.n2554 0.0525185
R6753 GND.n2861 GND.n2860 0.0525185
R6754 GND.n2862 GND.n2861 0.0525185
R6755 GND.n2876 GND.n2875 0.0525185
R6756 GND.n2877 GND.n2876 0.0525185
R6757 GND.n2870 GND.n2869 0.0525185
R6758 GND.n2871 GND.n2870 0.0525185
R6759 GND.n2864 GND.n2863 0.0525185
R6760 GND.n2865 GND.n2864 0.0525185
R6761 GND.n2879 GND.n2878 0.0525185
R6762 GND.n2880 GND.n2879 0.0525185
R6763 GND.n3158 GND.n3157 0.0525185
R6764 GND.n3159 GND.n3158 0.0525185
R6765 GND.n3173 GND.n3172 0.0525185
R6766 GND.n3174 GND.n3173 0.0525185
R6767 GND.n3167 GND.n3166 0.0525185
R6768 GND.n3168 GND.n3167 0.0525185
R6769 GND.n3161 GND.n3160 0.0525185
R6770 GND.n3162 GND.n3161 0.0525185
R6771 GND.n3176 GND.n3175 0.0525185
R6772 GND.n3177 GND.n3176 0.0525185
R6773 GND.n3315 GND.n3314 0.0525185
R6774 GND.n3316 GND.n3315 0.0525185
R6775 GND.n3330 GND.n3329 0.0525185
R6776 GND.n3331 GND.n3330 0.0525185
R6777 GND.n3324 GND.n3323 0.0525185
R6778 GND.n3325 GND.n3324 0.0525185
R6779 GND.n3318 GND.n3317 0.0525185
R6780 GND.n3319 GND.n3318 0.0525185
R6781 GND.n3333 GND.n3332 0.0525185
R6782 GND.n3334 GND.n3333 0.0525185
R6783 GND.n3473 GND.n3472 0.0525185
R6784 GND.n3474 GND.n3473 0.0525185
R6785 GND.n3488 GND.n3487 0.0525185
R6786 GND.n3489 GND.n3488 0.0525185
R6787 GND.n3482 GND.n3481 0.0525185
R6788 GND.n3483 GND.n3482 0.0525185
R6789 GND.n3476 GND.n3475 0.0525185
R6790 GND.n3477 GND.n3476 0.0525185
R6791 GND.n3491 GND.n3490 0.0525185
R6792 GND.n3492 GND.n3491 0.0525185
R6793 GND.n7263 GND.n7262 0.0525185
R6794 GND.n7264 GND.n7263 0.0525185
R6795 GND.n7278 GND.n7277 0.0525185
R6796 GND.n7279 GND.n7278 0.0525185
R6797 GND.n7272 GND.n7271 0.0525185
R6798 GND.n7273 GND.n7272 0.0525185
R6799 GND.n7266 GND.n7265 0.0525185
R6800 GND.n7267 GND.n7266 0.0525185
R6801 GND.n7281 GND.n7280 0.0525185
R6802 GND.n7282 GND.n7281 0.0525185
R6803 GND.n16 GND.n15 0.0525185
R6804 GND.n17 GND.n16 0.0525185
R6805 GND.n9 GND.n8 0.0525185
R6806 GND.n10 GND.n9 0.0525185
R6807 GND.n22 GND.n21 0.0525185
R6808 GND.n23 GND.n22 0.0525185
R6809 GND.n7 GND.n6 0.0525185
R6810 GND.n11 GND.n7 0.0525185
R6811 GND.n25 GND.n24 0.0525185
R6812 GND.n26 GND.n25 0.0525185
R6813 GND.n116 GND.n115 0.0525185
R6814 GND.n117 GND.n116 0.0525185
R6815 GND.n131 GND.n130 0.0525185
R6816 GND.n132 GND.n131 0.0525185
R6817 GND.n125 GND.n124 0.0525185
R6818 GND.n126 GND.n125 0.0525185
R6819 GND.n119 GND.n118 0.0525185
R6820 GND.n120 GND.n119 0.0525185
R6821 GND.n134 GND.n133 0.0525185
R6822 GND.n135 GND.n134 0.0525185
R6823 GND.n268 GND.n267 0.0525185
R6824 GND.n269 GND.n268 0.0525185
R6825 GND.n283 GND.n282 0.0525185
R6826 GND.n284 GND.n283 0.0525185
R6827 GND.n277 GND.n276 0.0525185
R6828 GND.n278 GND.n277 0.0525185
R6829 GND.n271 GND.n270 0.0525185
R6830 GND.n272 GND.n271 0.0525185
R6831 GND.n286 GND.n285 0.0525185
R6832 GND.n287 GND.n286 0.0525185
R6833 GND.n1631 GND.n1630 0.0525185
R6834 GND.n1632 GND.n1631 0.0525185
R6835 GND.n1646 GND.n1645 0.0525185
R6836 GND.n1647 GND.n1646 0.0525185
R6837 GND.n1640 GND.n1639 0.0525185
R6838 GND.n1641 GND.n1640 0.0525185
R6839 GND.n1634 GND.n1633 0.0525185
R6840 GND.n1635 GND.n1634 0.0525185
R6841 GND.n1649 GND.n1648 0.0525185
R6842 GND.n1650 GND.n1649 0.0525185
R6843 GND.n2051 GND.n2050 0.0525185
R6844 GND.n2052 GND.n2051 0.0525185
R6845 GND.n2032 GND.n2031 0.0525185
R6846 GND.n2031 GND.n2030 0.0525185
R6847 GND.n421 GND.n420 0.0525185
R6848 GND.n422 GND.n421 0.0525185
R6849 GND.n436 GND.n435 0.0525185
R6850 GND.n437 GND.n436 0.0525185
R6851 GND.n430 GND.n429 0.0525185
R6852 GND.n431 GND.n430 0.0525185
R6853 GND.n424 GND.n423 0.0525185
R6854 GND.n425 GND.n424 0.0525185
R6855 GND.n439 GND.n438 0.0525185
R6856 GND.n440 GND.n439 0.0525185
R6857 GND.n740 GND.n739 0.0525185
R6858 GND.n741 GND.n740 0.0525185
R6859 GND.n755 GND.n754 0.0525185
R6860 GND.n756 GND.n755 0.0525185
R6861 GND.n749 GND.n748 0.0525185
R6862 GND.n750 GND.n749 0.0525185
R6863 GND.n743 GND.n742 0.0525185
R6864 GND.n744 GND.n743 0.0525185
R6865 GND.n758 GND.n757 0.0525185
R6866 GND.n759 GND.n758 0.0525185
R6867 GND.n847 GND.n846 0.0525185
R6868 GND.n848 GND.n847 0.0525185
R6869 GND.n862 GND.n861 0.0525185
R6870 GND.n863 GND.n862 0.0525185
R6871 GND.n856 GND.n855 0.0525185
R6872 GND.n857 GND.n856 0.0525185
R6873 GND.n850 GND.n849 0.0525185
R6874 GND.n851 GND.n850 0.0525185
R6875 GND.n865 GND.n864 0.0525185
R6876 GND.n866 GND.n865 0.0525185
R6877 GND.n7789 GND.n7788 0.0525185
R6878 GND.n7790 GND.n7789 0.0525185
R6879 GND.n7801 GND.n7800 0.0525185
R6880 GND.n7802 GND.n7801 0.0525185
R6881 GND.n7795 GND.n7794 0.0525185
R6882 GND.n7796 GND.n7795 0.0525185
R6883 GND.n1356 GND.n1355 0.0523204
R6884 GND.n1361 GND.n1360 0.0523204
R6885 GND.n2093 GND.n1361 0.0523204
R6886 GND.n1074 GND.n1073 0.0523204
R6887 GND.n1082 GND.n1081 0.0523204
R6888 GND.n7348 GND.n1082 0.0523204
R6889 GND.n1087 GND.n1086 0.0523204
R6890 GND.n7348 GND.n1087 0.0523204
R6891 GND.n1092 GND.n1091 0.0523204
R6892 GND.n7348 GND.n1092 0.0523204
R6893 GND.n1097 GND.n1096 0.0523204
R6894 GND.n7348 GND.n1097 0.0523204
R6895 GND.n1102 GND.n1101 0.0523204
R6896 GND.n7348 GND.n1102 0.0523204
R6897 GND.n1107 GND.n1106 0.0523204
R6898 GND.n7348 GND.n1107 0.0523204
R6899 GND.n1112 GND.n1111 0.0523204
R6900 GND.n7348 GND.n1112 0.0523204
R6901 GND.n1120 GND.n1119 0.0523204
R6902 GND.n7348 GND.n1120 0.0523204
R6903 GND.n1128 GND.n1127 0.0523204
R6904 GND.n7348 GND.n1128 0.0523204
R6905 GND.n1136 GND.n1135 0.0523204
R6906 GND.n7348 GND.n1136 0.0523204
R6907 GND.n1144 GND.n1143 0.0523204
R6908 GND.n7348 GND.n1144 0.0523204
R6909 GND.n1154 GND.n1153 0.0523204
R6910 GND.n7348 GND.n1154 0.0523204
R6911 GND.n1152 GND.n1151 0.0523204
R6912 GND.n7348 GND.n1152 0.0523204
R6913 GND.n1903 GND.n1900 0.0516364
R6914 GND.n1860 GND.n1857 0.0516364
R6915 GND.n7037 GND.n7036 0.0516364
R6916 GND.n2509 GND.n2506 0.0516364
R6917 GND.n2834 GND.n2831 0.0516364
R6918 GND.n3131 GND.n3128 0.0516364
R6919 GND.n7231 GND.n7228 0.0516364
R6920 GND.n4763 GND.n4760 0.0516364
R6921 GND.n5429 GND.n5428 0.0516364
R6922 GND.n5931 GND.n5928 0.0516364
R6923 GND.n6100 GND.n6097 0.0516364
R6924 GND.n6264 GND.n6261 0.0516364
R6925 GND.n6573 GND.n6570 0.0516364
R6926 GND.n713 GND.n710 0.0516364
R6927 GND.n7760 GND.n7757 0.0516364
R6928 GND.n7595 GND.n7592 0.0516364
R6929 GND.n6841 GND.n6840 0.0500734
R6930 GND.n1944 GND.n1943 0.0494583
R6931 GND.n1751 GND.n1712 0.0494583
R6932 GND.n7024 GND.n7023 0.0494583
R6933 GND.n2400 GND.n2388 0.0494583
R6934 GND.n2725 GND.n2713 0.0494583
R6935 GND.n3049 GND.n3037 0.0494583
R6936 GND.n7149 GND.n7110 0.0494583
R6937 GND.n4842 GND.n4803 0.0494583
R6938 GND.n5419 GND.n5418 0.0494583
R6939 GND.n5914 GND.n5913 0.0494583
R6940 GND.n5988 GND.n5976 0.0494583
R6941 GND.n6155 GND.n6143 0.0494583
R6942 GND.n6319 GND.n6307 0.0494583
R6943 GND.n607 GND.n595 0.0494583
R6944 GND.n7650 GND.n7638 0.0494583
R6945 GND.n7530 GND.n7518 0.0494583
R6946 GND.n1916 GND.n1903 0.0493636
R6947 GND.n1873 GND.n1860 0.0493636
R6948 GND.n7036 GND.n7033 0.0493636
R6949 GND.n2522 GND.n2509 0.0493636
R6950 GND.n2847 GND.n2834 0.0493636
R6951 GND.n3144 GND.n3131 0.0493636
R6952 GND.n7244 GND.n7231 0.0493636
R6953 GND.n4776 GND.n4763 0.0493636
R6954 GND.n5428 GND.n5425 0.0493636
R6955 GND.n5944 GND.n5931 0.0493636
R6956 GND.n6113 GND.n6100 0.0493636
R6957 GND.n6277 GND.n6264 0.0493636
R6958 GND.n6586 GND.n6573 0.0493636
R6959 GND.n726 GND.n713 0.0493636
R6960 GND.n7773 GND.n7760 0.0493636
R6961 GND.n7608 GND.n7595 0.0493636
R6962 GND GND.n5191 0.0490201
R6963 GND GND.n4288 0.0490201
R6964 GND.n5476 GND 0.0484167
R6965 GND GND.n5465 0.0484167
R6966 GND.n1923 GND 0.0484167
R6967 GND.n1690 GND 0.0484167
R6968 GND.n6898 GND 0.0484167
R6969 GND.n2366 GND 0.0484167
R6970 GND.n2691 GND 0.0484167
R6971 GND.n3015 GND 0.0484167
R6972 GND.n7088 GND 0.0484167
R6973 GND.n4783 GND 0.0484167
R6974 GND.n5265 GND 0.0484167
R6975 GND.n5787 GND 0.0484167
R6976 GND.n5954 GND 0.0484167
R6977 GND.n6121 GND 0.0484167
R6978 GND.n6285 GND 0.0484167
R6979 GND.n573 GND 0.0484167
R6980 GND.n7616 GND 0.0484167
R6981 GND.n7496 GND 0.0484167
R6982 GND.n4407 GND 0.0484167
R6983 GND GND.n4396 0.0484167
R6984 GND.n1914 GND.n1913 0.0483725
R6985 GND.n1871 GND.n1870 0.0483725
R6986 GND.n6892 GND.n6891 0.0483725
R6987 GND.n2520 GND.n2519 0.0483725
R6988 GND.n2845 GND.n2844 0.0483725
R6989 GND.n3142 GND.n3141 0.0483725
R6990 GND.n7242 GND.n7241 0.0483725
R6991 GND.n4774 GND.n4773 0.0483725
R6992 GND.n5259 GND.n5258 0.0483725
R6993 GND.n5942 GND.n5941 0.0483725
R6994 GND.n6111 GND.n6110 0.0483725
R6995 GND.n6275 GND.n6274 0.0483725
R6996 GND.n6584 GND.n6583 0.0483725
R6997 GND.n724 GND.n723 0.0483725
R6998 GND.n7771 GND.n7770 0.0483725
R6999 GND.n7606 GND.n7605 0.0483725
R7000 GND.n3646 GND.n3644 0.048348
R7001 GND.n1145 GND.n790 0.0483051
R7002 GND.n7354 GND.n7352 0.0483051
R7003 GND.n2087 GND.n2086 0.0483051
R7004 GND.n1129 GND.n318 0.0483051
R7005 GND.n1137 GND.n471 0.0483051
R7006 GND.n1121 GND.n166 0.0483051
R7007 GND.n7316 GND.n7314 0.0483051
R7008 GND.n4174 GND.n4172 0.0483051
R7009 GND.n3368 GND.n3366 0.0483051
R7010 GND.n3211 GND.n3209 0.0483051
R7011 GND.n2914 GND.n2912 0.0483051
R7012 GND.n2589 GND.n2587 0.0483051
R7013 GND.n2265 GND.n2263 0.0483051
R7014 GND.n7342 GND.n7341 0.0483051
R7015 GND.n2099 GND.n2097 0.0483051
R7016 GND.n1939 GND.n1936 0.0464802
R7017 GND.n1706 GND.n1703 0.0464802
R7018 GND.n6914 GND.n6911 0.0464802
R7019 GND.n2382 GND.n2379 0.0464802
R7020 GND.n2707 GND.n2704 0.0464802
R7021 GND.n3031 GND.n3028 0.0464802
R7022 GND.n7104 GND.n7101 0.0464802
R7023 GND.n4799 GND.n4796 0.0464802
R7024 GND.n5281 GND.n5278 0.0464802
R7025 GND.n5803 GND.n5800 0.0464802
R7026 GND.n5970 GND.n5967 0.0464802
R7027 GND.n6137 GND.n6134 0.0464802
R7028 GND.n6301 GND.n6298 0.0464802
R7029 GND.n589 GND.n586 0.0464802
R7030 GND.n7632 GND.n7629 0.0464802
R7031 GND.n7512 GND.n7509 0.0464802
R7032 GND.n6791 GND 0.04425
R7033 GND.n4369 GND 0.04425
R7034 GND.n7561 GND.n7560 0.0425017
R7035 GND.n7560 GND.n7559 0.0425017
R7036 GND.n7658 GND.n7657 0.0425017
R7037 GND.n7659 GND.n7658 0.0425017
R7038 GND.n7692 GND.n7691 0.0425017
R7039 GND.n7691 GND.n7690 0.0425017
R7040 GND.n614 GND.n613 0.0425017
R7041 GND.n615 GND.n614 0.0425017
R7042 GND.n645 GND.n644 0.0425017
R7043 GND.n644 GND.n643 0.0425017
R7044 GND.n6326 GND.n6325 0.0425017
R7045 GND.n6327 GND.n6326 0.0425017
R7046 GND.n6357 GND.n6356 0.0425017
R7047 GND.n6356 GND.n6355 0.0425017
R7048 GND.n6162 GND.n6161 0.0425017
R7049 GND.n6163 GND.n6162 0.0425017
R7050 GND.n6193 GND.n6192 0.0425017
R7051 GND.n6192 GND.n6191 0.0425017
R7052 GND.n5995 GND.n5994 0.0425017
R7053 GND.n5996 GND.n5995 0.0425017
R7054 GND.n6029 GND.n6028 0.0425017
R7055 GND.n6028 GND.n6027 0.0425017
R7056 GND.n5812 GND.n5811 0.0425017
R7057 GND.n5813 GND.n5812 0.0425017
R7058 GND.n5846 GND.n5845 0.0425017
R7059 GND.n5845 GND.n5844 0.0425017
R7060 GND.n5290 GND.n5289 0.0425017
R7061 GND.n5291 GND.n5290 0.0425017
R7062 GND.n5324 GND.n5323 0.0425017
R7063 GND.n5323 GND.n5322 0.0425017
R7064 GND.n4849 GND.n4848 0.0425017
R7065 GND.n4850 GND.n4849 0.0425017
R7066 GND.n4883 GND.n4882 0.0425017
R7067 GND.n4882 GND.n4881 0.0425017
R7068 GND.n7156 GND.n7155 0.0425017
R7069 GND.n7157 GND.n7156 0.0425017
R7070 GND.n7190 GND.n7189 0.0425017
R7071 GND.n7189 GND.n7188 0.0425017
R7072 GND.n3056 GND.n3055 0.0425017
R7073 GND.n3057 GND.n3056 0.0425017
R7074 GND.n3090 GND.n3089 0.0425017
R7075 GND.n3089 GND.n3088 0.0425017
R7076 GND.n2732 GND.n2731 0.0425017
R7077 GND.n2733 GND.n2732 0.0425017
R7078 GND.n2766 GND.n2765 0.0425017
R7079 GND.n2765 GND.n2764 0.0425017
R7080 GND.n2407 GND.n2406 0.0425017
R7081 GND.n2408 GND.n2407 0.0425017
R7082 GND.n2441 GND.n2440 0.0425017
R7083 GND.n2440 GND.n2439 0.0425017
R7084 GND.n6923 GND.n6922 0.0425017
R7085 GND.n6924 GND.n6923 0.0425017
R7086 GND.n6957 GND.n6956 0.0425017
R7087 GND.n6956 GND.n6955 0.0425017
R7088 GND.n1758 GND.n1757 0.0425017
R7089 GND.n1759 GND.n1758 0.0425017
R7090 GND.n1792 GND.n1791 0.0425017
R7091 GND.n1791 GND.n1790 0.0425017
R7092 GND.n1567 GND.n1566 0.0425017
R7093 GND.n1568 GND.n1567 0.0425017
R7094 GND.n1601 GND.n1600 0.0425017
R7095 GND.n1600 GND.n1599 0.0425017
R7096 GND.n1549 GND.n1548 0.0425017
R7097 GND.n1550 GND.n1549 0.0425017
R7098 GND.n7369 GND.n7368 0.0415714
R7099 GND.n1365 GND.n1364 0.0415714
R7100 GND.n330 GND.n329 0.0415714
R7101 GND.n483 GND.n482 0.0415714
R7102 GND.n178 GND.n177 0.0415714
R7103 GND.n1487 GND.n1486 0.0415714
R7104 GND.n1386 GND.n1385 0.0415714
R7105 GND.n4186 GND.n4185 0.0415714
R7106 GND.n3380 GND.n3379 0.0415714
R7107 GND.n3223 GND.n3222 0.0415714
R7108 GND.n2926 GND.n2925 0.0415714
R7109 GND.n2601 GND.n2600 0.0415714
R7110 GND.n2277 GND.n2276 0.0415714
R7111 GND.n2115 GND.n2114 0.0415714
R7112 GND.n1247 GND.n1246 0.0415714
R7113 GND.n7395 GND.n7394 0.0415714
R7114 GND.n7435 GND.n7434 0.0406786
R7115 GND.n1988 GND.n1987 0.0406786
R7116 GND.n332 GND.n331 0.0406786
R7117 GND.n485 GND.n484 0.0406786
R7118 GND.n180 GND.n179 0.0406786
R7119 GND.n1515 GND.n1488 0.0406786
R7120 GND.n1467 GND.n1387 0.0406786
R7121 GND.n4188 GND.n4187 0.0406786
R7122 GND.n3382 GND.n3381 0.0406786
R7123 GND.n3225 GND.n3224 0.0406786
R7124 GND.n2928 GND.n2927 0.0406786
R7125 GND.n2603 GND.n2602 0.0406786
R7126 GND.n2279 GND.n2278 0.0406786
R7127 GND.n2117 GND.n2116 0.0406786
R7128 GND.n1249 GND.n1248 0.0406786
R7129 GND.n7416 GND.n7396 0.0406786
R7130 GND.n4160 GND.n4159 0.0390862
R7131 GND.n789 GND 0.0386944
R7132 GND.n7353 GND 0.0386944
R7133 GND.n2085 GND 0.0386944
R7134 GND.n317 GND 0.0386944
R7135 GND.n470 GND 0.0386944
R7136 GND.n165 GND 0.0386944
R7137 GND.n56 GND 0.0386944
R7138 GND.n7315 GND 0.0386944
R7139 GND.n4173 GND 0.0386944
R7140 GND.n3367 GND 0.0386944
R7141 GND.n3210 GND 0.0386944
R7142 GND.n2913 GND 0.0386944
R7143 GND.n2588 GND 0.0386944
R7144 GND.n2264 GND 0.0386944
R7145 GND.n7340 GND 0.0386944
R7146 GND.n2098 GND 0.0386944
R7147 GND.n3641 GND.n3628 0.0381984
R7148 GND.n4042 GND.n4040 0.0367903
R7149 GND.n6754 GND.n5464 0.0356562
R7150 GND.n4395 GND.n4394 0.0356562
R7151 GND.n5215 GND 0.0353684
R7152 GND.n4312 GND 0.0353684
R7153 GND.n4958 GND.n4957 0.0352222
R7154 GND.n1948 GND.n1946 0.0345278
R7155 GND.n1744 GND.n1743 0.0345278
R7156 GND.n7016 GND.n7015 0.0345278
R7157 GND.n2393 GND.n2392 0.0345278
R7158 GND.n2718 GND.n2717 0.0345278
R7159 GND.n3042 GND.n3041 0.0345278
R7160 GND.n7142 GND.n7141 0.0345278
R7161 GND.n4835 GND.n4834 0.0345278
R7162 GND.n5411 GND.n5410 0.0345278
R7163 GND.n5906 GND.n5905 0.0345278
R7164 GND.n5981 GND.n5980 0.0345278
R7165 GND.n6148 GND.n6147 0.0345278
R7166 GND.n6312 GND.n6311 0.0345278
R7167 GND.n600 GND.n599 0.0345278
R7168 GND.n7643 GND.n7642 0.0345278
R7169 GND.n7523 GND.n7522 0.0345278
R7170 GND.n3664 GND.n3663 0.0339821
R7171 GND.n1943 GND.n1942 0.0337917
R7172 GND.n1712 GND.n1709 0.0337917
R7173 GND.n7025 GND.n7024 0.0337917
R7174 GND.n2388 GND.n2385 0.0337917
R7175 GND.n2713 GND.n2710 0.0337917
R7176 GND.n3037 GND.n3034 0.0337917
R7177 GND.n7110 GND.n7107 0.0337917
R7178 GND.n4803 GND.n4802 0.0337917
R7179 GND.n5420 GND.n5419 0.0337917
R7180 GND.n5915 GND.n5914 0.0337917
R7181 GND.n5976 GND.n5973 0.0337917
R7182 GND.n6143 GND.n6140 0.0337917
R7183 GND.n6307 GND.n6304 0.0337917
R7184 GND.n595 GND.n592 0.0337917
R7185 GND.n7638 GND.n7635 0.0337917
R7186 GND.n7518 GND.n7515 0.0337917
R7187 GND.n5460 GND 0.033625
R7188 GND.n6865 GND 0.033625
R7189 GND.n1936 GND.n1935 0.0335935
R7190 GND.n1703 GND.n1702 0.0335935
R7191 GND.n6911 GND.n6910 0.0335935
R7192 GND.n2379 GND.n2378 0.0335935
R7193 GND.n2704 GND.n2703 0.0335935
R7194 GND.n3028 GND.n3027 0.0335935
R7195 GND.n7101 GND.n7100 0.0335935
R7196 GND.n4796 GND.n4795 0.0335935
R7197 GND.n5278 GND.n5277 0.0335935
R7198 GND.n5800 GND.n5799 0.0335935
R7199 GND.n5967 GND.n5966 0.0335935
R7200 GND.n6134 GND.n6133 0.0335935
R7201 GND.n6298 GND.n6297 0.0335935
R7202 GND.n586 GND.n585 0.0335935
R7203 GND.n7629 GND.n7628 0.0335935
R7204 GND.n7509 GND.n7508 0.0335935
R7205 GND GND.n4970 0.0324444
R7206 GND GND.n4960 0.0324444
R7207 GND.n5238 GND 0.0324444
R7208 GND.n4330 GND 0.0324444
R7209 GND.n3680 GND.n3674 0.03175
R7210 GND.n6792 GND.n6791 0.03175
R7211 GND.n4370 GND.n4369 0.03175
R7212 GND.n5027 GND.n5026 0.0307632
R7213 GND.n5026 GND.n5024 0.0307632
R7214 GND.n5009 GND.n5007 0.0307632
R7215 GND.n5007 GND.n5003 0.0307632
R7216 GND.n5003 GND.n4999 0.0307632
R7217 GND.n4999 GND.n4997 0.0307632
R7218 GND.n4997 GND.n4993 0.0307632
R7219 GND.n4993 GND.n4991 0.0307632
R7220 GND.n4991 GND.n4987 0.0307632
R7221 GND.n4658 GND.n4657 0.0307632
R7222 GND.n4657 GND.n4655 0.0307632
R7223 GND.n4655 GND.n4651 0.0307632
R7224 GND.n4651 GND.n4649 0.0307632
R7225 GND.n4649 GND.n4645 0.0307632
R7226 GND.n4645 GND.n4643 0.0307632
R7227 GND.n4643 GND.n4639 0.0307632
R7228 GND.n4639 GND.n4635 0.0307632
R7229 GND.n4635 GND.n4612 0.0307632
R7230 GND.n4676 GND.n4674 0.0307632
R7231 GND.n4680 GND.n4676 0.0307632
R7232 GND.n4682 GND.n4680 0.0307632
R7233 GND.n4684 GND.n4682 0.0307632
R7234 GND.n4688 GND.n4686 0.0307632
R7235 GND.n4692 GND.n4688 0.0307632
R7236 GND.n4694 GND.n4692 0.0307632
R7237 GND.n4698 GND.n4694 0.0307632
R7238 GND.n4700 GND.n4698 0.0307632
R7239 GND.n4741 GND.n4739 0.0307632
R7240 GND.n4739 GND.n4735 0.0307632
R7241 GND.n4735 GND.n4733 0.0307632
R7242 GND.n4733 GND.n4729 0.0307632
R7243 GND.n4729 GND.n4727 0.0307632
R7244 GND.n4727 GND.n4723 0.0307632
R7245 GND.n4723 GND.n4721 0.0307632
R7246 GND.n4720 GND.n4719 0.0307632
R7247 GND.n4719 GND.n4717 0.0307632
R7248 GND.n4717 GND.n4713 0.0307632
R7249 GND.n4713 GND.n4711 0.0307632
R7250 GND.n4711 GND.n4608 0.0307632
R7251 GND.n5192 GND 0.0307632
R7252 GND.n5201 GND 0.0307632
R7253 GND.n4289 GND 0.0307632
R7254 GND.n4298 GND 0.0307632
R7255 GND.n5216 GND.n5215 0.0301053
R7256 GND.n4313 GND.n4312 0.0301053
R7257 GND.n3650 GND 0.0300162
R7258 GND.n4960 GND.n4958 0.0296667
R7259 GND.n4957 GND.n4953 0.0296667
R7260 GND.n7783 GND.n7782 0.0296391
R7261 GND.n842 GND.n841 0.0296391
R7262 GND.n735 GND.n734 0.0296391
R7263 GND.n416 GND.n415 0.0296391
R7264 GND.n1626 GND.n1625 0.0296391
R7265 GND.n263 GND.n262 0.0296391
R7266 GND.n111 GND.n110 0.0296391
R7267 GND.n2 GND.n1 0.0296391
R7268 GND.n7258 GND.n7257 0.0296391
R7269 GND.n3468 GND.n3467 0.0296391
R7270 GND.n3310 GND.n3309 0.0296391
R7271 GND.n3153 GND.n3152 0.0296391
R7272 GND.n2856 GND.n2855 0.0296391
R7273 GND.n2531 GND.n2530 0.0296391
R7274 GND.n2207 GND.n2206 0.0296391
R7275 GND.n1182 GND.n1181 0.0296391
R7276 GND.n4933 GND.n4932 0.0294474
R7277 GND.n5461 GND.n5460 0.028625
R7278 GND.n5462 GND.n5461 0.028625
R7279 GND.n6866 GND.n6865 0.028625
R7280 GND.n6867 GND.n6866 0.028625
R7281 GND.n4973 GND.n4972 0.0284605
R7282 GND.n4667 GND.n4612 0.0282663
R7283 GND.n6754 GND 0.0268889
R7284 GND.n4394 GND 0.0268889
R7285 GND.n4923 GND.n4608 0.0262926
R7286 GND.n5024 GND.n5020 0.0238553
R7287 GND.n4701 GND.n4700 0.0231974
R7288 GND.n4662 GND.n4661 0.0225395
R7289 GND.n4742 GND.n4741 0.0225395
R7290 GND.n5010 GND.n5009 0.0218816
R7291 GND.n6835 GND 0.02175
R7292 GND.n6829 GND 0.02175
R7293 GND.n6823 GND 0.02175
R7294 GND.n6817 GND 0.02175
R7295 GND.n6811 GND 0.02175
R7296 GND.n7080 GND 0.02175
R7297 GND.n7074 GND 0.02175
R7298 GND.n7068 GND 0.02175
R7299 GND.n7062 GND 0.02175
R7300 GND.n7056 GND 0.02175
R7301 GND.n4980 GND.n4975 0.0212237
R7302 GND.n6805 GND.n6804 0.0209918
R7303 GND.n7050 GND.n7049 0.0209918
R7304 GND.n7372 GND.n7371 0.0208901
R7305 GND.n7375 GND.n7372 0.0208901
R7306 GND.n7380 GND.n7379 0.0208901
R7307 GND.n1368 GND.n1367 0.0208901
R7308 GND.n1371 GND.n1368 0.0208901
R7309 GND.n1376 GND.n1375 0.0208901
R7310 GND.n325 GND.n324 0.0208901
R7311 GND.n328 GND.n325 0.0208901
R7312 GND.n338 GND.n337 0.0208901
R7313 GND.n478 GND.n477 0.0208901
R7314 GND.n481 GND.n478 0.0208901
R7315 GND.n491 GND.n490 0.0208901
R7316 GND.n173 GND.n172 0.0208901
R7317 GND.n176 GND.n173 0.0208901
R7318 GND.n186 GND.n185 0.0208901
R7319 GND.n1482 GND.n1481 0.0208901
R7320 GND.n1485 GND.n1482 0.0208901
R7321 GND.n1521 GND.n1520 0.0208901
R7322 GND.n1381 GND.n1380 0.0208901
R7323 GND.n1384 GND.n1381 0.0208901
R7324 GND.n1473 GND.n1472 0.0208901
R7325 GND.n4181 GND.n4180 0.0208901
R7326 GND.n4184 GND.n4181 0.0208901
R7327 GND.n4194 GND.n4193 0.0208901
R7328 GND.n3375 GND.n3374 0.0208901
R7329 GND.n3378 GND.n3375 0.0208901
R7330 GND.n3388 GND.n3387 0.0208901
R7331 GND.n3218 GND.n3217 0.0208901
R7332 GND.n3221 GND.n3218 0.0208901
R7333 GND.n3231 GND.n3230 0.0208901
R7334 GND.n2921 GND.n2920 0.0208901
R7335 GND.n2924 GND.n2921 0.0208901
R7336 GND.n2934 GND.n2933 0.0208901
R7337 GND.n2596 GND.n2595 0.0208901
R7338 GND.n2599 GND.n2596 0.0208901
R7339 GND.n2609 GND.n2608 0.0208901
R7340 GND.n2272 GND.n2271 0.0208901
R7341 GND.n2275 GND.n2272 0.0208901
R7342 GND.n2285 GND.n2284 0.0208901
R7343 GND.n2110 GND.n2109 0.0208901
R7344 GND.n2113 GND.n2110 0.0208901
R7345 GND.n2123 GND.n2122 0.0208901
R7346 GND.n1242 GND.n1241 0.0208901
R7347 GND.n1245 GND.n1242 0.0208901
R7348 GND.n1255 GND.n1254 0.0208901
R7349 GND.n7390 GND.n7389 0.0208901
R7350 GND.n7393 GND.n7390 0.0208901
R7351 GND.n7422 GND.n7421 0.0208901
R7352 GND.n6596 GND.n6595 0.020607
R7353 GND.n6594 GND.n6593 0.020607
R7354 GND.n7781 GND.n7780 0.020607
R7355 GND.n4670 GND.n4669 0.0205658
R7356 GND.n1881 GND.n1880 0.0203417
R7357 GND.n7255 GND.n7254 0.0203417
R7358 GND.n4072 GND.n4068 0.0202922
R7359 GND.n7365 GND.n7362 0.0200011
R7360 GND.n2017 GND.n2015 0.0200011
R7361 GND.n515 GND.n513 0.0200011
R7362 GND.n210 GND.n208 0.0200011
R7363 GND.n1509 GND.n1507 0.0200011
R7364 GND.n1461 GND.n1459 0.0200011
R7365 GND.n4218 GND.n4216 0.0200011
R7366 GND.n3412 GND.n3410 0.0200011
R7367 GND.n3255 GND.n3253 0.0200011
R7368 GND.n2958 GND.n2956 0.0200011
R7369 GND.n2633 GND.n2631 0.0200011
R7370 GND.n2309 GND.n2307 0.0200011
R7371 GND.n2147 GND.n2145 0.0200011
R7372 GND.n1279 GND.n1277 0.0200011
R7373 GND.n362 GND.n360 0.0200011
R7374 GND.n7410 GND.n7408 0.0200011
R7375 GND.n1893 GND 0.0198182
R7376 GND.n1850 GND 0.0198182
R7377 GND.n7041 GND 0.0198182
R7378 GND.n2499 GND 0.0198182
R7379 GND.n2824 GND 0.0198182
R7380 GND.n3121 GND 0.0198182
R7381 GND.n7221 GND 0.0198182
R7382 GND.n4753 GND 0.0198182
R7383 GND.n5433 GND 0.0198182
R7384 GND.n5921 GND 0.0198182
R7385 GND.n6090 GND 0.0198182
R7386 GND.n6254 GND 0.0198182
R7387 GND.n6563 GND 0.0198182
R7388 GND.n703 GND 0.0198182
R7389 GND.n7750 GND 0.0198182
R7390 GND.n7585 GND 0.0198182
R7391 GND.n4068 GND.n4067 0.0197936
R7392 GND.n7432 GND.n7380 0.0195603
R7393 GND.n1985 GND.n1376 0.0195603
R7394 GND.n339 GND.n338 0.0195603
R7395 GND.n492 GND.n491 0.0195603
R7396 GND.n187 GND.n186 0.0195603
R7397 GND.n1522 GND.n1521 0.0195603
R7398 GND.n1474 GND.n1473 0.0195603
R7399 GND.n4195 GND.n4194 0.0195603
R7400 GND.n3389 GND.n3388 0.0195603
R7401 GND.n3232 GND.n3231 0.0195603
R7402 GND.n2935 GND.n2934 0.0195603
R7403 GND.n2610 GND.n2609 0.0195603
R7404 GND.n2286 GND.n2285 0.0195603
R7405 GND.n2124 GND.n2123 0.0195603
R7406 GND.n1256 GND.n1255 0.0195603
R7407 GND.n7423 GND.n7422 0.0195603
R7408 GND.n7253 GND.n7252 0.0191946
R7409 GND.n1897 GND.n1896 0.0186818
R7410 GND.n1854 GND.n1853 0.0186818
R7411 GND.n7040 GND.n7038 0.0186818
R7412 GND.n2503 GND.n2502 0.0186818
R7413 GND.n2828 GND.n2827 0.0186818
R7414 GND.n3125 GND.n3124 0.0186818
R7415 GND.n7225 GND.n7224 0.0186818
R7416 GND.n4757 GND.n4756 0.0186818
R7417 GND.n5432 GND.n5430 0.0186818
R7418 GND.n5925 GND.n5924 0.0186818
R7419 GND.n6094 GND.n6093 0.0186818
R7420 GND.n6258 GND.n6257 0.0186818
R7421 GND.n6567 GND.n6566 0.0186818
R7422 GND.n707 GND.n706 0.0186818
R7423 GND.n7754 GND.n7753 0.0186818
R7424 GND.n7589 GND.n7588 0.0186818
R7425 GND.n4928 GND.n4927 0.0185921
R7426 GND.n3641 GND.n3633 0.0183571
R7427 GND.n5484 GND 0.0182083
R7428 GND.n4415 GND 0.0182083
R7429 GND.n4062 GND.n4061 0.0179743
R7430 GND GND.n4961 0.0178611
R7431 GND.n7472 GND.n7471 0.0176904
R7432 GND.n553 GND.n552 0.0176904
R7433 GND.n244 GND.n243 0.0176904
R7434 GND.n83 GND.n82 0.0176904
R7435 GND.n1425 GND.n1424 0.0176904
R7436 GND.n4252 GND.n4251 0.0176904
R7437 GND.n3449 GND.n3448 0.0176904
R7438 GND.n3291 GND.n3290 0.0176904
R7439 GND.n2995 GND.n2994 0.0176904
R7440 GND.n2671 GND.n2670 0.0176904
R7441 GND.n2346 GND.n2345 0.0176904
R7442 GND.n2188 GND.n2187 0.0176904
R7443 GND.n1307 GND.n1306 0.0176904
R7444 GND.n4987 GND.n4985 0.0172763
R7445 GND.n824 GND.n823 0.0172687
R7446 GND.n2066 GND.n2065 0.0172687
R7447 GND.n398 GND.n397 0.0172687
R7448 GND GND.n5475 0.0171667
R7449 GND.n1935 GND.n1933 0.0171667
R7450 GND.n1702 GND.n1700 0.0171667
R7451 GND.n6910 GND.n6908 0.0171667
R7452 GND.n2378 GND.n2376 0.0171667
R7453 GND.n2703 GND.n2701 0.0171667
R7454 GND.n3027 GND.n3025 0.0171667
R7455 GND.n7100 GND.n7098 0.0171667
R7456 GND.n4795 GND.n4793 0.0171667
R7457 GND.n5277 GND.n5275 0.0171667
R7458 GND.n5799 GND.n5797 0.0171667
R7459 GND.n5966 GND.n5964 0.0171667
R7460 GND.n6133 GND.n6131 0.0171667
R7461 GND.n6297 GND.n6295 0.0171667
R7462 GND.n585 GND.n583 0.0171667
R7463 GND.n7628 GND.n7626 0.0171667
R7464 GND.n7508 GND.n7506 0.0171667
R7465 GND GND.n4406 0.0171667
R7466 GND.n4939 GND.n4935 0.0171667
R7467 GND.n4941 GND.n4939 0.0171667
R7468 GND.n4945 GND.n4941 0.0171667
R7469 GND.n5037 GND.n5035 0.0171667
R7470 GND.n5035 GND.n5031 0.0171667
R7471 GND.n3637 GND.n3636 0.0167601
R7472 GND.n5019 GND.n5017 0.0166184
R7473 GND.n1912 GND.n1911 0.0164091
R7474 GND.n1869 GND.n1868 0.0164091
R7475 GND.n6890 GND.n6889 0.0164091
R7476 GND.n2518 GND.n2517 0.0164091
R7477 GND.n2843 GND.n2842 0.0164091
R7478 GND.n3140 GND.n3139 0.0164091
R7479 GND.n7240 GND.n7239 0.0164091
R7480 GND.n4772 GND.n4771 0.0164091
R7481 GND.n5257 GND.n5256 0.0164091
R7482 GND.n5940 GND.n5939 0.0164091
R7483 GND.n6109 GND.n6108 0.0164091
R7484 GND.n6273 GND.n6272 0.0164091
R7485 GND.n6582 GND.n6581 0.0164091
R7486 GND.n722 GND.n721 0.0164091
R7487 GND.n7769 GND.n7768 0.0164091
R7488 GND.n7604 GND.n7603 0.0164091
R7489 GND.n3689 GND.n3687 0.016125
R7490 GND.n4747 GND.n4705 0.0159605
R7491 GND.n4630 GND 0.0158101
R7492 GND.n5031 GND.n5029 0.0157174
R7493 GND GND.n5027 0.0156316
R7494 GND.n4658 GND 0.0156316
R7495 GND.n4686 GND 0.0156316
R7496 GND GND.n4720 0.0156316
R7497 GND.n4747 GND.n4746 0.0153026
R7498 GND.n7822 GND.n7821 0.0152059
R7499 GND.n894 GND.n893 0.0152059
R7500 GND.n787 GND.n786 0.0152059
R7501 GND.n468 GND.n467 0.0152059
R7502 GND.n1686 GND.n1685 0.0152059
R7503 GND.n315 GND.n314 0.0152059
R7504 GND.n163 GND.n162 0.0152059
R7505 GND.n54 GND.n53 0.0152059
R7506 GND.n7310 GND.n7309 0.0152059
R7507 GND.n3520 GND.n3519 0.0152059
R7508 GND.n3362 GND.n3361 0.0152059
R7509 GND.n3205 GND.n3204 0.0152059
R7510 GND.n2908 GND.n2907 0.0152059
R7511 GND.n2583 GND.n2582 0.0152059
R7512 GND.n2259 GND.n2258 0.0152059
R7513 GND.n1234 GND.n1233 0.0152059
R7514 GND.n7458 GND.n7457 0.015169
R7515 GND.n7457 GND.t1239 0.015169
R7516 GND.n7456 GND.n7455 0.015169
R7517 GND.t1239 GND.n7456 0.015169
R7518 GND.n7454 GND.n7453 0.015169
R7519 GND.t1239 GND.n7454 0.015169
R7520 GND.n538 GND.n537 0.015169
R7521 GND.n537 GND.t1170 0.015169
R7522 GND.n536 GND.n535 0.015169
R7523 GND.t1170 GND.n536 0.015169
R7524 GND.n534 GND.n533 0.015169
R7525 GND.t1170 GND.n534 0.015169
R7526 GND.n233 GND.n232 0.015169
R7527 GND.n232 GND.t671 0.015169
R7528 GND.n231 GND.n230 0.015169
R7529 GND.t671 GND.n231 0.015169
R7530 GND.n229 GND.n228 0.015169
R7531 GND.t671 GND.n229 0.015169
R7532 GND.n4241 GND.n4240 0.015169
R7533 GND.n4240 GND.t673 0.015169
R7534 GND.n4239 GND.n4238 0.015169
R7535 GND.t673 GND.n4239 0.015169
R7536 GND.n4237 GND.n4236 0.015169
R7537 GND.t673 GND.n4237 0.015169
R7538 GND.n3278 GND.n3277 0.015169
R7539 GND.n3277 GND.t127 0.015169
R7540 GND.n3276 GND.n3275 0.015169
R7541 GND.t127 GND.n3276 0.015169
R7542 GND.n3274 GND.n3273 0.015169
R7543 GND.t127 GND.n3274 0.015169
R7544 GND.n2656 GND.n2655 0.015169
R7545 GND.n2655 GND.t606 0.015169
R7546 GND.n2654 GND.n2653 0.015169
R7547 GND.t606 GND.n2654 0.015169
R7548 GND.n2652 GND.n2651 0.015169
R7549 GND.t606 GND.n2652 0.015169
R7550 GND.n2170 GND.n2169 0.015169
R7551 GND.n2169 GND.t740 0.015169
R7552 GND.n2168 GND.n2167 0.015169
R7553 GND.t740 GND.n2168 0.015169
R7554 GND.n2166 GND.n2165 0.015169
R7555 GND.t740 GND.n2166 0.015169
R7556 GND.n1302 GND.n1301 0.015169
R7557 GND.n1301 GND.t818 0.015169
R7558 GND.n1300 GND.n1299 0.015169
R7559 GND.t818 GND.n1300 0.015169
R7560 GND.n1298 GND.n1297 0.015169
R7561 GND.t818 GND.n1298 0.015169
R7562 GND.n1265 GND.n1264 0.015169
R7563 GND.n1266 GND.n1265 0.015169
R7564 GND.n2181 GND.n2180 0.015169
R7565 GND.n2182 GND.n2181 0.015169
R7566 GND.n2184 GND.n2183 0.015169
R7567 GND.n2183 GND.n2182 0.015169
R7568 GND.n1263 GND.n1262 0.015169
R7569 GND.n1266 GND.n1263 0.015169
R7570 GND.n2133 GND.n2132 0.015169
R7571 GND.n2134 GND.n2133 0.015169
R7572 GND.n2175 GND.n2174 0.015169
R7573 GND.n2342 GND.n2341 0.015169
R7574 GND.n2341 GND.n2340 0.015169
R7575 GND.n2131 GND.n2130 0.015169
R7576 GND.n2134 GND.n2131 0.015169
R7577 GND.n2332 GND.n2331 0.015169
R7578 GND.n2331 GND.t743 0.015169
R7579 GND.n2330 GND.n2329 0.015169
R7580 GND.t743 GND.n2330 0.015169
R7581 GND.n2328 GND.n2327 0.015169
R7582 GND.t743 GND.n2328 0.015169
R7583 GND.n2295 GND.n2294 0.015169
R7584 GND.n2296 GND.n2295 0.015169
R7585 GND.n2337 GND.n2336 0.015169
R7586 GND.n2667 GND.n2666 0.015169
R7587 GND.n2666 GND.n2665 0.015169
R7588 GND.n2293 GND.n2292 0.015169
R7589 GND.n2296 GND.n2293 0.015169
R7590 GND.n2619 GND.n2618 0.015169
R7591 GND.n2620 GND.n2619 0.015169
R7592 GND.n2662 GND.n2661 0.015169
R7593 GND.n2661 GND.n2660 0.015169
R7594 GND.n2991 GND.n2990 0.015169
R7595 GND.n2617 GND.n2616 0.015169
R7596 GND.n2620 GND.n2617 0.015169
R7597 GND.n2981 GND.n2980 0.015169
R7598 GND.n2980 GND.t408 0.015169
R7599 GND.n2979 GND.n2978 0.015169
R7600 GND.t408 GND.n2979 0.015169
R7601 GND.n2977 GND.n2976 0.015169
R7602 GND.t408 GND.n2977 0.015169
R7603 GND.n2944 GND.n2943 0.015169
R7604 GND.n2945 GND.n2944 0.015169
R7605 GND.n2987 GND.n2986 0.015169
R7606 GND.n2986 GND.n2985 0.015169
R7607 GND.n3287 GND.n3286 0.015169
R7608 GND.n2942 GND.n2941 0.015169
R7609 GND.n2945 GND.n2942 0.015169
R7610 GND.n3241 GND.n3240 0.015169
R7611 GND.n3242 GND.n3241 0.015169
R7612 GND.n3283 GND.n3282 0.015169
R7613 GND.n3445 GND.n3444 0.015169
R7614 GND.n3444 GND.n3443 0.015169
R7615 GND.n3239 GND.n3238 0.015169
R7616 GND.n3242 GND.n3239 0.015169
R7617 GND.n3435 GND.n3434 0.015169
R7618 GND.n3434 GND.t162 0.015169
R7619 GND.n3433 GND.n3432 0.015169
R7620 GND.t162 GND.n3433 0.015169
R7621 GND.n3431 GND.n3430 0.015169
R7622 GND.t162 GND.n3431 0.015169
R7623 GND.n3398 GND.n3397 0.015169
R7624 GND.n3399 GND.n3398 0.015169
R7625 GND.n3440 GND.n3439 0.015169
R7626 GND.n4248 GND.n4247 0.015169
R7627 GND.n4247 GND.n4246 0.015169
R7628 GND.n3396 GND.n3395 0.015169
R7629 GND.n3399 GND.n3396 0.015169
R7630 GND.n4204 GND.n4203 0.015169
R7631 GND.n4205 GND.n4204 0.015169
R7632 GND.n1418 GND.n1417 0.015169
R7633 GND.n1419 GND.n1418 0.015169
R7634 GND.n1421 GND.n1420 0.015169
R7635 GND.n1420 GND.n1419 0.015169
R7636 GND.n4202 GND.n4201 0.015169
R7637 GND.n4205 GND.n4202 0.015169
R7638 GND.n1407 GND.n1406 0.015169
R7639 GND.n1406 GND.t1148 0.015169
R7640 GND.n1405 GND.n1404 0.015169
R7641 GND.t1148 GND.n1405 0.015169
R7642 GND.n1403 GND.n1402 0.015169
R7643 GND.t1148 GND.n1403 0.015169
R7644 GND.n1447 GND.n1446 0.015169
R7645 GND.n1448 GND.n1447 0.015169
R7646 GND.n1413 GND.n1412 0.015169
R7647 GND.n1412 GND.n1411 0.015169
R7648 GND.n79 GND.n78 0.015169
R7649 GND.n1445 GND.n1444 0.015169
R7650 GND.n1448 GND.n1445 0.015169
R7651 GND.n983 GND.n982 0.015169
R7652 GND.n982 GND.t777 0.015169
R7653 GND.n94 GND.n93 0.015169
R7654 GND.n95 GND.n94 0.015169
R7655 GND.n990 GND.n989 0.015169
R7656 GND.n989 GND.t1282 0.015169
R7657 GND.n1495 GND.n1494 0.015169
R7658 GND.n1496 GND.n1495 0.015169
R7659 GND.n75 GND.n74 0.015169
R7660 GND.n74 GND.n73 0.015169
R7661 GND.n72 GND.n71 0.015169
R7662 GND.n73 GND.n72 0.015169
R7663 GND.n1493 GND.n1492 0.015169
R7664 GND.n1496 GND.n1493 0.015169
R7665 GND.n196 GND.n195 0.015169
R7666 GND.n197 GND.n196 0.015169
R7667 GND.n239 GND.n238 0.015169
R7668 GND.n238 GND.n237 0.015169
R7669 GND.n194 GND.n193 0.015169
R7670 GND.n197 GND.n194 0.015169
R7671 GND.n394 GND.n393 0.015169
R7672 GND.n385 GND.n384 0.015169
R7673 GND.n384 GND.t712 0.015169
R7674 GND.n381 GND.n380 0.015169
R7675 GND.t712 GND.n381 0.015169
R7676 GND.n383 GND.n382 0.015169
R7677 GND.t712 GND.n383 0.015169
R7678 GND.n1668 GND.n1666 0.015169
R7679 GND.n1669 GND.n1668 0.015169
R7680 GND.n1672 GND.n1671 0.015169
R7681 GND.n1671 GND.n1669 0.015169
R7682 GND.n2000 GND.n1999 0.015169
R7683 GND.n2003 GND.n2000 0.015169
R7684 GND.n2002 GND.n2001 0.015169
R7685 GND.n2003 GND.n2002 0.015169
R7686 GND.n2055 GND.n2054 0.015169
R7687 GND.n2054 GND.n2053 0.015169
R7688 GND.n1990 GND.n1989 0.015169
R7689 GND.n1991 GND.n1990 0.015169
R7690 GND.n2043 GND.n2042 0.015169
R7691 GND.t1169 GND.n2043 0.015169
R7692 GND.n2044 GND.t1169 0.015169
R7693 GND.n2045 GND.n2044 0.015169
R7694 GND.n2041 GND.n2040 0.015169
R7695 GND.t1169 GND.n2041 0.015169
R7696 GND.n3706 GND.n3705 0.015169
R7697 GND.n3707 GND.n3706 0.015169
R7698 GND.n3721 GND.n3720 0.015169
R7699 GND.n3722 GND.n3721 0.015169
R7700 GND.n3736 GND.n3735 0.015169
R7701 GND.n3737 GND.n3736 0.015169
R7702 GND.n3751 GND.n3750 0.015169
R7703 GND.n3752 GND.n3751 0.015169
R7704 GND.n3770 GND.n3769 0.015169
R7705 GND.n3771 GND.n3770 0.015169
R7706 GND.n3785 GND.n3784 0.015169
R7707 GND.n3786 GND.n3785 0.015169
R7708 GND.n3800 GND.n3799 0.015169
R7709 GND.n3801 GND.n3800 0.015169
R7710 GND.n3815 GND.n3814 0.015169
R7711 GND.n3816 GND.n3815 0.015169
R7712 GND.n3833 GND.n3832 0.015169
R7713 GND.n3834 GND.n3833 0.015169
R7714 GND.n3857 GND.n3856 0.015169
R7715 GND.n3858 GND.n3857 0.015169
R7716 GND.n3877 GND.n3876 0.015169
R7717 GND.n3878 GND.n3877 0.015169
R7718 GND.n3894 GND.n3893 0.015169
R7719 GND.n3895 GND.n3894 0.015169
R7720 GND.n3909 GND.n3908 0.015169
R7721 GND.n3910 GND.n3909 0.015169
R7722 GND.n3924 GND.n3923 0.015169
R7723 GND.n3925 GND.n3924 0.015169
R7724 GND.n3939 GND.n3938 0.015169
R7725 GND.n3940 GND.n3939 0.015169
R7726 GND.n3956 GND.n3955 0.015169
R7727 GND.n3957 GND.n3956 0.015169
R7728 GND.n3971 GND.n3970 0.015169
R7729 GND.n3972 GND.n3971 0.015169
R7730 GND.n3986 GND.n3985 0.015169
R7731 GND.n3987 GND.n3986 0.015169
R7732 GND.n4001 GND.n4000 0.015169
R7733 GND.n4002 GND.n4001 0.015169
R7734 GND.n3669 GND.n3668 0.015169
R7735 GND.n4017 GND.n4016 0.015169
R7736 GND.n4018 GND.n4017 0.015169
R7737 GND.n3655 GND.n3654 0.015169
R7738 GND.n3656 GND.n3655 0.015169
R7739 GND.n348 GND.n347 0.015169
R7740 GND.n349 GND.n348 0.015169
R7741 GND.n390 GND.n389 0.015169
R7742 GND.n549 GND.n548 0.015169
R7743 GND.n548 GND.n547 0.015169
R7744 GND.n346 GND.n345 0.015169
R7745 GND.n349 GND.n346 0.015169
R7746 GND.n501 GND.n500 0.015169
R7747 GND.n502 GND.n501 0.015169
R7748 GND.n544 GND.n543 0.015169
R7749 GND.n543 GND.n542 0.015169
R7750 GND.n820 GND.n819 0.015169
R7751 GND.n499 GND.n498 0.015169
R7752 GND.n502 GND.n499 0.015169
R7753 GND.n810 GND.n809 0.015169
R7754 GND.n809 GND.t854 0.015169
R7755 GND.n808 GND.n807 0.015169
R7756 GND.t854 GND.n808 0.015169
R7757 GND.n806 GND.n805 0.015169
R7758 GND.t854 GND.n806 0.015169
R7759 GND.n7385 GND.n7384 0.015169
R7760 GND.n7386 GND.n7385 0.015169
R7761 GND.n816 GND.n815 0.015169
R7762 GND.n815 GND.n814 0.015169
R7763 GND.n7468 GND.n7467 0.015169
R7764 GND.n7383 GND.n7382 0.015169
R7765 GND.n7386 GND.n7383 0.015169
R7766 GND.n7480 GND.n7479 0.015169
R7767 GND.n7479 GND.n7478 0.015169
R7768 GND.n7464 GND.n7463 0.015169
R7769 GND.n7463 GND.n7462 0.015169
R7770 GND.n2094 GND.n1327 0.014943
R7771 GND.n1080 GND.n1079 0.014943
R7772 GND.n1085 GND.n1084 0.014943
R7773 GND.n1090 GND.n1089 0.014943
R7774 GND.n1095 GND.n1094 0.014943
R7775 GND.n1100 GND.n1099 0.014943
R7776 GND.n1105 GND.n1104 0.014943
R7777 GND.n1110 GND.n1109 0.014943
R7778 GND.n1118 GND.n1117 0.014943
R7779 GND.n1126 GND.n1125 0.014943
R7780 GND.n1134 GND.n1133 0.014943
R7781 GND.n1142 GND.n1141 0.014943
R7782 GND.n7349 GND.n897 0.014943
R7783 GND.n1150 GND.n1149 0.014943
R7784 GND.n1359 GND.n1358 0.014943
R7785 GND.n1077 GND.n1076 0.014943
R7786 GND.n5017 GND.n5014 0.0146447
R7787 GND.n4588 GND.n4586 0.0146077
R7788 GND.n1358 GND.n1357 0.0144432
R7789 GND.n1327 GND.n1326 0.0144432
R7790 GND.n1076 GND.n1075 0.0144432
R7791 GND.n1079 GND.n1078 0.0144432
R7792 GND.n1084 GND.n1083 0.0144432
R7793 GND.n1089 GND.n1088 0.0144432
R7794 GND.n1094 GND.n1093 0.0144432
R7795 GND.n1099 GND.n1098 0.0144432
R7796 GND.n1104 GND.n1103 0.0144432
R7797 GND.n1109 GND.n1108 0.0144432
R7798 GND.n1117 GND.n1116 0.0144432
R7799 GND.n1125 GND.n1124 0.0144432
R7800 GND.n1133 GND.n1132 0.0144432
R7801 GND.n1141 GND.n1140 0.0144432
R7802 GND.n897 GND.n896 0.0144432
R7803 GND.n1149 GND.n1148 0.0144432
R7804 GND.n3620 GND.n3619 0.0143889
R7805 GND.n6597 GND.n6596 0.0143235
R7806 GND.n6595 GND.n6594 0.0143235
R7807 GND.n6593 GND.n6592 0.0143235
R7808 GND.n733 GND.n732 0.0143235
R7809 GND.n7780 GND.n7779 0.0143235
R7810 GND.n1882 GND.n1881 0.0141412
R7811 GND.n1880 GND.n1879 0.0141412
R7812 GND.n7027 GND.n7026 0.0141412
R7813 GND.n2529 GND.n2528 0.0141412
R7814 GND.n2854 GND.n2853 0.0141412
R7815 GND.n3151 GND.n3150 0.0141412
R7816 GND.n7251 GND.n7250 0.0141412
R7817 GND.n7254 GND.n7253 0.0141412
R7818 GND.n7256 GND.n7255 0.0141412
R7819 GND.n5951 GND.n5950 0.0141412
R7820 GND.n1928 GND.n1927 0.0140417
R7821 GND.n1695 GND.n1694 0.0140417
R7822 GND.n6903 GND.n6902 0.0140417
R7823 GND.n2371 GND.n2370 0.0140417
R7824 GND.n2696 GND.n2695 0.0140417
R7825 GND.n3020 GND.n3019 0.0140417
R7826 GND.n7093 GND.n7092 0.0140417
R7827 GND.n4788 GND.n4787 0.0140417
R7828 GND.n5270 GND.n5269 0.0140417
R7829 GND.n5792 GND.n5791 0.0140417
R7830 GND.n5959 GND.n5958 0.0140417
R7831 GND.n6126 GND.n6125 0.0140417
R7832 GND.n6290 GND.n6289 0.0140417
R7833 GND.n578 GND.n577 0.0140417
R7834 GND.n7621 GND.n7620 0.0140417
R7835 GND.n7501 GND.n7500 0.0140417
R7836 GND.n4985 GND.n4984 0.0139868
R7837 GND.n7377 GND.n7376 0.0138596
R7838 GND.n1373 GND.n1372 0.0138596
R7839 GND.n335 GND.n334 0.0138596
R7840 GND.n488 GND.n487 0.0138596
R7841 GND.n183 GND.n182 0.0138596
R7842 GND.n1518 GND.n1517 0.0138596
R7843 GND.n1470 GND.n1469 0.0138596
R7844 GND.n4191 GND.n4190 0.0138596
R7845 GND.n3385 GND.n3384 0.0138596
R7846 GND.n3228 GND.n3227 0.0138596
R7847 GND.n2931 GND.n2930 0.0138596
R7848 GND.n2606 GND.n2605 0.0138596
R7849 GND.n2282 GND.n2281 0.0138596
R7850 GND.n2120 GND.n2119 0.0138596
R7851 GND.n1252 GND.n1251 0.0138596
R7852 GND.n7419 GND.n7418 0.0138596
R7853 GND.n5518 GND.n5514 0.012734
R7854 GND.n5556 GND.n5552 0.012734
R7855 GND.n5552 GND.n5550 0.012734
R7856 GND.n5550 GND.n5546 0.012734
R7857 GND.n5546 GND.n5544 0.012734
R7858 GND.n5544 GND.n5540 0.012734
R7859 GND.n5540 GND.n5538 0.012734
R7860 GND.n5538 GND.n5534 0.012734
R7861 GND.n5534 GND.n5532 0.012734
R7862 GND.n5531 GND.n5530 0.012734
R7863 GND.n5530 GND.n5528 0.012734
R7864 GND.n5578 GND.n5574 0.012734
R7865 GND.n5582 GND.n5578 0.012734
R7866 GND.n5584 GND.n5582 0.012734
R7867 GND.n5588 GND.n5584 0.012734
R7868 GND.n5590 GND.n5588 0.012734
R7869 GND.n5594 GND.n5590 0.012734
R7870 GND.n5596 GND.n5594 0.012734
R7871 GND.n5600 GND.n5596 0.012734
R7872 GND.n5602 GND.n5600 0.012734
R7873 GND.n5603 GND.n5602 0.012734
R7874 GND.n5608 GND.n5606 0.012734
R7875 GND.n5612 GND.n5608 0.012734
R7876 GND.n5614 GND.n5612 0.012734
R7877 GND.n5641 GND.n5637 0.012734
R7878 GND.n5637 GND.n5633 0.012734
R7879 GND.n5633 GND.n5631 0.012734
R7880 GND.n5631 GND.n5627 0.012734
R7881 GND.n5627 GND.n5625 0.012734
R7882 GND.n5625 GND.n5621 0.012734
R7883 GND.n5621 GND.n5500 0.012734
R7884 GND.n5782 GND.n5780 0.012734
R7885 GND.n5779 GND.n5778 0.012734
R7886 GND.n5778 GND.n5776 0.012734
R7887 GND.n5655 GND.n5651 0.012734
R7888 GND.n5659 GND.n5655 0.012734
R7889 GND.n5661 GND.n5659 0.012734
R7890 GND.n5665 GND.n5661 0.012734
R7891 GND.n5667 GND.n5665 0.012734
R7892 GND.n5671 GND.n5667 0.012734
R7893 GND.n5673 GND.n5671 0.012734
R7894 GND.n5677 GND.n5673 0.012734
R7895 GND.n5679 GND.n5677 0.012734
R7896 GND.n5680 GND.n5679 0.012734
R7897 GND.n5685 GND.n5683 0.012734
R7898 GND.n5700 GND.n5698 0.012734
R7899 GND.n5704 GND.n5700 0.012734
R7900 GND.n5708 GND.n5704 0.012734
R7901 GND.n5710 GND.n5708 0.012734
R7902 GND.n5714 GND.n5710 0.012734
R7903 GND.n5716 GND.n5714 0.012734
R7904 GND.n5720 GND.n5716 0.012734
R7905 GND.n5722 GND.n5720 0.012734
R7906 GND.n5726 GND.n5722 0.012734
R7907 GND.n5728 GND.n5726 0.012734
R7908 GND.n5729 GND.n5728 0.012734
R7909 GND.n5734 GND.n5732 0.012734
R7910 GND.n5737 GND.n5734 0.012734
R7911 GND.n5739 GND.n5737 0.012734
R7912 GND.n5759 GND.n5757 0.012734
R7913 GND.n5754 GND.n5753 0.012734
R7914 GND.n5753 GND.n5751 0.012734
R7915 GND.n5751 GND.n5747 0.012734
R7916 GND.n5747 GND.n5745 0.012734
R7917 GND.n4443 GND.n4439 0.012734
R7918 GND.n4445 GND.n4443 0.012734
R7919 GND.n4460 GND.n4458 0.012734
R7920 GND.n4464 GND.n4460 0.012734
R7921 GND.n4466 GND.n4464 0.012734
R7922 GND.n4470 GND.n4466 0.012734
R7923 GND.n4472 GND.n4470 0.012734
R7924 GND.n4476 GND.n4472 0.012734
R7925 GND.n4478 GND.n4476 0.012734
R7926 GND.n4479 GND.n4478 0.012734
R7927 GND.n4484 GND.n4482 0.012734
R7928 GND.n4488 GND.n4484 0.012734
R7929 GND.n4534 GND.n4532 0.012734
R7930 GND.n4532 GND.n4528 0.012734
R7931 GND.n4528 GND.n4524 0.012734
R7932 GND.n4524 GND.n4522 0.012734
R7933 GND.n4522 GND.n4518 0.012734
R7934 GND.n4518 GND.n4516 0.012734
R7935 GND.n4516 GND.n4512 0.012734
R7936 GND.n4512 GND.n4510 0.012734
R7937 GND.n4510 GND.n4506 0.012734
R7938 GND.n4506 GND.n4504 0.012734
R7939 GND.n4503 GND.n4502 0.012734
R7940 GND.n4502 GND.n4500 0.012734
R7941 GND.n4500 GND.n4496 0.012734
R7942 GND.n4556 GND.n4552 0.012734
R7943 GND.n4558 GND.n4556 0.012734
R7944 GND.n4562 GND.n4558 0.012734
R7945 GND.n4564 GND.n4562 0.012734
R7946 GND.n4568 GND.n4564 0.012734
R7947 GND.n4570 GND.n4568 0.012734
R7948 GND.n4574 GND.n4570 0.012734
R7949 GND.n4576 GND.n4574 0.012734
R7950 GND.n5048 GND.n5046 0.012734
R7951 GND.n5052 GND.n5048 0.012734
R7952 GND.n5091 GND.n5089 0.012734
R7953 GND.n5089 GND.n5085 0.012734
R7954 GND.n5085 GND.n5081 0.012734
R7955 GND.n5081 GND.n5079 0.012734
R7956 GND.n5079 GND.n5075 0.012734
R7957 GND.n5075 GND.n5073 0.012734
R7958 GND.n5073 GND.n5069 0.012734
R7959 GND.n5069 GND.n5067 0.012734
R7960 GND.n5067 GND.n5063 0.012734
R7961 GND.n5063 GND.n5061 0.012734
R7962 GND.n5060 GND.n5059 0.012734
R7963 GND.n5059 GND.n4430 0.012734
R7964 GND.n5111 GND.n5109 0.012734
R7965 GND.n5115 GND.n5111 0.012734
R7966 GND.n5119 GND.n5115 0.012734
R7967 GND.n5121 GND.n5119 0.012734
R7968 GND.n5125 GND.n5121 0.012734
R7969 GND.n5127 GND.n5125 0.012734
R7970 GND.n5131 GND.n5127 0.012734
R7971 GND.n5133 GND.n5131 0.012734
R7972 GND.n5137 GND.n5133 0.012734
R7973 GND.n5139 GND.n5137 0.012734
R7974 GND.n5140 GND.n5139 0.012734
R7975 GND.n5145 GND.n5143 0.012734
R7976 GND.n5148 GND.n5145 0.012734
R7977 GND.n5150 GND.n5148 0.012734
R7978 GND.n5170 GND.n5168 0.012734
R7979 GND.n5165 GND.n5164 0.012734
R7980 GND.n5164 GND.n5162 0.012734
R7981 GND.n5162 GND.n5158 0.012734
R7982 GND.n5158 GND.n5156 0.012734
R7983 GND.n6427 GND.n6423 0.012734
R7984 GND.n6429 GND.n6427 0.012734
R7985 GND.n6464 GND.n6460 0.012734
R7986 GND.n6460 GND.n6458 0.012734
R7987 GND.n6458 GND.n6454 0.012734
R7988 GND.n6454 GND.n6452 0.012734
R7989 GND.n6452 GND.n6448 0.012734
R7990 GND.n6448 GND.n6446 0.012734
R7991 GND.n6446 GND.n6442 0.012734
R7992 GND.n6442 GND.n6440 0.012734
R7993 GND.n6439 GND.n6438 0.012734
R7994 GND.n6438 GND.n6436 0.012734
R7995 GND.n6486 GND.n6482 0.012734
R7996 GND.n6490 GND.n6486 0.012734
R7997 GND.n6492 GND.n6490 0.012734
R7998 GND.n6496 GND.n6492 0.012734
R7999 GND.n6498 GND.n6496 0.012734
R8000 GND.n6502 GND.n6498 0.012734
R8001 GND.n6504 GND.n6502 0.012734
R8002 GND.n6508 GND.n6504 0.012734
R8003 GND.n6510 GND.n6508 0.012734
R8004 GND.n6511 GND.n6510 0.012734
R8005 GND.n6516 GND.n6514 0.012734
R8006 GND.n6520 GND.n6516 0.012734
R8007 GND.n6522 GND.n6520 0.012734
R8008 GND.n6553 GND.n6549 0.012734
R8009 GND.n6549 GND.n6545 0.012734
R8010 GND.n6545 GND.n6543 0.012734
R8011 GND.n6543 GND.n6539 0.012734
R8012 GND.n6539 GND.n6537 0.012734
R8013 GND.n6537 GND.n6533 0.012734
R8014 GND.n6533 GND.n6531 0.012734
R8015 GND.n6531 GND.n5496 0.012734
R8016 GND.n6606 GND.n6604 0.012734
R8017 GND.n6610 GND.n6606 0.012734
R8018 GND.n6649 GND.n6647 0.012734
R8019 GND.n6647 GND.n6643 0.012734
R8020 GND.n6643 GND.n6639 0.012734
R8021 GND.n6639 GND.n6637 0.012734
R8022 GND.n6637 GND.n6633 0.012734
R8023 GND.n6633 GND.n6631 0.012734
R8024 GND.n6631 GND.n6627 0.012734
R8025 GND.n6627 GND.n6625 0.012734
R8026 GND.n6625 GND.n6621 0.012734
R8027 GND.n6621 GND.n6619 0.012734
R8028 GND.n6618 GND.n6617 0.012734
R8029 GND.n6617 GND.n5494 0.012734
R8030 GND.n6669 GND.n6667 0.012734
R8031 GND.n6673 GND.n6669 0.012734
R8032 GND.n6677 GND.n6673 0.012734
R8033 GND.n6679 GND.n6677 0.012734
R8034 GND.n6683 GND.n6679 0.012734
R8035 GND.n6685 GND.n6683 0.012734
R8036 GND.n6689 GND.n6685 0.012734
R8037 GND.n6691 GND.n6689 0.012734
R8038 GND.n6695 GND.n6691 0.012734
R8039 GND.n6697 GND.n6695 0.012734
R8040 GND.n6698 GND.n6697 0.012734
R8041 GND.n6703 GND.n6701 0.012734
R8042 GND.n6706 GND.n6703 0.012734
R8043 GND.n6708 GND.n6706 0.012734
R8044 GND.n6728 GND.n6726 0.012734
R8045 GND.n6723 GND.n6722 0.012734
R8046 GND.n6722 GND.n6720 0.012734
R8047 GND.n6720 GND.n6716 0.012734
R8048 GND.n6716 GND.n6714 0.012734
R8049 GND.n4932 GND.n4928 0.0126711
R8050 GND.n5519 GND.n5518 0.0126011
R8051 GND.n5043 GND.n5042 0.0126011
R8052 GND.n6601 GND.n6600 0.0126011
R8053 GND.n5198 GND 0.0123421
R8054 GND.n4295 GND 0.0123421
R8055 GND.n5783 GND.n5500 0.0123351
R8056 GND.n5686 GND.n5685 0.0123351
R8057 GND.n4962 GND 0.0123056
R8058 GND GND.n4953 0.0123056
R8059 GND.n4954 GND 0.0123056
R8060 GND GND.n6753 0.0123056
R8061 GND GND.n6790 0.0123056
R8062 GND GND.n5245 0.0123056
R8063 GND GND.n4392 0.0123056
R8064 GND GND.n4368 0.0123056
R8065 GND GND.n4337 0.0123056
R8066 GND.n7362 GND.n7361 0.0120741
R8067 GND.n2015 GND.n2014 0.0120741
R8068 GND.n513 GND.n512 0.0120741
R8069 GND.n208 GND.n207 0.0120741
R8070 GND.n1507 GND.n1506 0.0120741
R8071 GND.n1459 GND.n1458 0.0120741
R8072 GND.n4216 GND.n4215 0.0120741
R8073 GND.n3410 GND.n3409 0.0120741
R8074 GND.n3253 GND.n3252 0.0120741
R8075 GND.n2956 GND.n2955 0.0120741
R8076 GND.n2631 GND.n2630 0.0120741
R8077 GND.n2307 GND.n2306 0.0120741
R8078 GND.n2145 GND.n2144 0.0120741
R8079 GND.n1277 GND.n1276 0.0120741
R8080 GND.n360 GND.n359 0.0120741
R8081 GND.n7408 GND.n7407 0.0120741
R8082 GND.n4489 GND.n4488 0.0120691
R8083 GND.n6436 GND.n6432 0.0120691
R8084 GND.n5038 GND.n5037 0.0117319
R8085 GND GND.n6777 0.0116111
R8086 GND.n5226 GND 0.0116111
R8087 GND GND.n4355 0.0116111
R8088 GND.n4318 GND 0.0116111
R8089 GND.n6598 GND.n5951 0.0115679
R8090 GND.n5528 GND.n5524 0.0115372
R8091 GND.n2100 GND.n1325 0.0114919
R8092 GND.n7337 GND.n7336 0.0114919
R8093 GND.n7334 GND.n7333 0.0114919
R8094 GND.n7331 GND.n7330 0.0114919
R8095 GND.n7328 GND.n7327 0.0114919
R8096 GND.n7325 GND.n7324 0.0114919
R8097 GND.n7318 GND.n7317 0.0114919
R8098 GND.n7841 GND.n7840 0.0114919
R8099 GND.n7838 GND.n7837 0.0114919
R8100 GND.n7835 GND.n7834 0.0114919
R8101 GND.n7832 GND.n7831 0.0114919
R8102 GND.n7829 GND.n7828 0.0114919
R8103 GND.n7826 GND.n7825 0.0114919
R8104 GND.n1623 GND.n1575 0.0112143
R8105 GND.n1841 GND.n1766 0.0112143
R8106 GND.n7006 GND.n6931 0.0112143
R8107 GND.n2490 GND.n2415 0.0112143
R8108 GND.n2815 GND.n2740 0.0112143
R8109 GND.n3112 GND.n3064 0.0112143
R8110 GND.n7212 GND.n7164 0.0112143
R8111 GND.n4905 GND.n4857 0.0112143
R8112 GND.n5373 GND.n5298 0.0112143
R8113 GND.n5895 GND.n5820 0.0112143
R8114 GND.n6081 GND.n6003 0.0112143
R8115 GND.n6245 GND.n6170 0.0112143
R8116 GND.n6409 GND.n6334 0.0112143
R8117 GND.n694 GND.n622 0.0112143
R8118 GND.n7741 GND.n7666 0.0112143
R8119 GND.n7577 GND.n7535 0.0112143
R8120 GND.n7361 GND 0.0111481
R8121 GND.n2014 GND 0.0111481
R8122 GND.n512 GND 0.0111481
R8123 GND.n207 GND 0.0111481
R8124 GND.n1506 GND 0.0111481
R8125 GND.n1458 GND 0.0111481
R8126 GND.n4215 GND 0.0111481
R8127 GND.n3409 GND 0.0111481
R8128 GND.n3252 GND 0.0111481
R8129 GND.n2955 GND 0.0111481
R8130 GND.n2630 GND 0.0111481
R8131 GND.n2306 GND 0.0111481
R8132 GND.n2144 GND 0.0111481
R8133 GND.n1276 GND 0.0111481
R8134 GND.n359 GND 0.0111481
R8135 GND.n7407 GND 0.0111481
R8136 GND GND.n5214 0.0110263
R8137 GND GND.n4311 0.0110263
R8138 GND.n3696 GND.n3694 0.0109167
R8139 GND.n5642 GND.n5641 0.0107394
R8140 GND.n5651 GND.n5649 0.0107394
R8141 GND.n5151 GND.n5150 0.0107394
R8142 GND.n6709 GND.n6708 0.0107394
R8143 GND.n4449 GND.n4445 0.0107015
R8144 GND.n6470 GND.n6429 0.0107015
R8145 GND.n4674 GND.n4670 0.0106974
R8146 GND.n5102 GND.n4430 0.0104355
R8147 GND.n6660 GND.n5494 0.0104355
R8148 GND.n3768 GND.n3767 0.0102222
R8149 GND.n5740 GND.n5739 0.0102074
R8150 GND.n4552 GND.n4548 0.0102074
R8151 GND.n5092 GND.n5091 0.0102074
R8152 GND.n6554 GND.n6553 0.0102074
R8153 GND.n6650 GND.n6649 0.0102074
R8154 GND.n3546 GND.n3545 0.0101468
R8155 GND.n3547 GND.n3546 0.0101468
R8156 GND.n3609 GND.n3608 0.0101468
R8157 GND.n3610 GND.n3609 0.0101468
R8158 GND.n3603 GND.n3602 0.0101468
R8159 GND.n3610 GND.n3603 0.0101468
R8160 GND.n3599 GND.n3598 0.0101468
R8161 GND.n3610 GND.n3599 0.0101468
R8162 GND.n3595 GND.n3594 0.0101468
R8163 GND.n3610 GND.n3595 0.0101468
R8164 GND.n3544 GND.n3543 0.0101468
R8165 GND.n3547 GND.n3544 0.0101468
R8166 GND.n3591 GND.n3590 0.0101468
R8167 GND.n3610 GND.n3591 0.0101468
R8168 GND.n3585 GND.n3584 0.0101468
R8169 GND.n3610 GND.n3585 0.0101468
R8170 GND.n3581 GND.n3580 0.0101468
R8171 GND.n3610 GND.n3581 0.0101468
R8172 GND.n3578 GND.n3577 0.0101468
R8173 GND.n3610 GND.n3578 0.0101468
R8174 GND.n3573 GND.n3572 0.0101468
R8175 GND.n3610 GND.n3573 0.0101468
R8176 GND.n3569 GND.n3568 0.0101468
R8177 GND.n3610 GND.n3569 0.0101468
R8178 GND.n3565 GND.n3564 0.0101468
R8179 GND.n3610 GND.n3565 0.0101468
R8180 GND.n3562 GND.n3561 0.0101468
R8181 GND.n3610 GND.n3562 0.0101468
R8182 GND.n3542 GND.n3541 0.0101468
R8183 GND.n3547 GND.n3542 0.0101468
R8184 GND.n3555 GND.n3554 0.0101468
R8185 GND.n3610 GND.n3555 0.0101468
R8186 GND.n3549 GND.n3548 0.0101468
R8187 GND.n3610 GND.n3549 0.0101468
R8188 GND.n4984 GND.n4980 0.0100395
R8189 GND.n4585 GND.n4581 0.0100149
R8190 GND GND.n5459 0.009875
R8191 GND GND.n6864 0.009875
R8192 GND.n5562 GND.n5521 0.00967553
R8193 GND.n3696 GND.n3695 0.00959091
R8194 GND.n5202 GND.n5185 0.00950855
R8195 GND.n4299 GND.n4282 0.00950855
R8196 GND.n4595 GND.n4593 0.00941473
R8197 GND.n4599 GND.n4595 0.00941473
R8198 GND.n4603 GND.n4599 0.00941473
R8199 GND.n4605 GND.n4603 0.00941473
R8200 GND.n4618 GND.n4616 0.00941473
R8201 GND.n4622 GND.n4618 0.00941473
R8202 GND.n4624 GND.n4622 0.00941473
R8203 GND.n4628 GND.n4624 0.00941473
R8204 GND.n5691 GND.n5690 0.00940957
R8205 GND.n5014 GND.n5010 0.00938158
R8206 GND.n6598 GND.n6597 0.00932473
R8207 GND.n4540 GND.n4491 0.00914362
R8208 GND.n6475 GND.n6418 0.00914362
R8209 GND.n6778 GND.n6768 0.00906279
R8210 GND.n4356 GND.n4346 0.00906279
R8211 GND.n4087 GND.n4083 0.00904142
R8212 GND.n4155 GND.n4154 0.00898517
R8213 GND.n4143 GND.n4142 0.00898517
R8214 GND.n4095 GND.n4094 0.00898517
R8215 GND.n4090 GND.n4089 0.00898517
R8216 GND.n4089 GND.n4087 0.00898517
R8217 GND.n4143 GND.n4140 0.00897458
R8218 GND.n4155 GND.n4152 0.00896398
R8219 GND.n4134 GND.n4132 0.00896398
R8220 GND.n4135 GND.n4134 0.00896398
R8221 GND.n4166 GND.n3523 0.00896398
R8222 GND.n4119 GND.n4117 0.00896398
R8223 GND.n4108 GND.n4107 0.00896398
R8224 GND.n4090 GND.n4081 0.00896398
R8225 GND.n4108 GND.n4105 0.0089428
R8226 GND.n5760 GND.n5759 0.00887766
R8227 GND.n4496 GND.n4494 0.00887766
R8228 GND.n5053 GND.n5052 0.00887766
R8229 GND.n6523 GND.n6522 0.00887766
R8230 GND.n6611 GND.n6610 0.00887766
R8231 GND.n7321 GND.n7320 0.00878716
R8232 GND.n4662 GND.n4632 0.00872368
R8233 GND.n4746 GND.n4742 0.00872368
R8234 GND.n5567 GND.n5508 0.0086117
R8235 GND.n4052 GND.n4044 0.00856452
R8236 GND.n5615 GND.n5614 0.00834574
R8237 GND.n5776 GND.n5772 0.00834574
R8238 GND.n5171 GND.n5170 0.00834574
R8239 GND.n6729 GND.n6728 0.00834574
R8240 GND GND.n4119 0.00822246
R8241 GND GND.n4971 0.00806579
R8242 GND.n4705 GND.n4701 0.00806579
R8243 GND.n7379 GND.n7377 0.00783909
R8244 GND.n1375 GND.n1373 0.00783909
R8245 GND.n337 GND.n335 0.00783909
R8246 GND.n490 GND.n488 0.00783909
R8247 GND.n185 GND.n183 0.00783909
R8248 GND.n1520 GND.n1518 0.00783909
R8249 GND.n1472 GND.n1470 0.00783909
R8250 GND.n4193 GND.n4191 0.00783909
R8251 GND.n3387 GND.n3385 0.00783909
R8252 GND.n3230 GND.n3228 0.00783909
R8253 GND.n2933 GND.n2931 0.00783909
R8254 GND.n2608 GND.n2606 0.00783909
R8255 GND.n2284 GND.n2282 0.00783909
R8256 GND.n2122 GND.n2120 0.00783909
R8257 GND.n1254 GND.n1252 0.00783909
R8258 GND.n7421 GND.n7419 0.00783909
R8259 GND.n5645 GND.n5644 0.00781383
R8260 GND.n5769 GND.n5506 0.00781383
R8261 GND.n3646 GND.n3645 0.00779984
R8262 GND.n6751 GND.n6736 0.00775202
R8263 GND.n6788 GND.n6763 0.00775202
R8264 GND.n5239 GND.n5224 0.00775202
R8265 GND.n5243 GND.n5222 0.00775202
R8266 GND.n4390 GND.n4375 0.00775202
R8267 GND.n4366 GND.n4341 0.00775202
R8268 GND.n4331 GND.n4316 0.00775202
R8269 GND.n4335 GND.n4314 0.00775202
R8270 GND.n4050 GND.n4049 0.00769258
R8271 GND.n4038 GND.n4037 0.00769258
R8272 GND.n5574 GND.n5572 0.00754787
R8273 GND.n3534 GND.n3533 0.00744444
R8274 GND.n3626 GND.n3538 0.00744444
R8275 GND.n5020 GND.n5019 0.00740789
R8276 GND.n7371 GND.n7370 0.00739975
R8277 GND.n1367 GND.n1366 0.00739975
R8278 GND.n324 GND.n323 0.00739975
R8279 GND.n477 GND.n476 0.00739975
R8280 GND.n172 GND.n171 0.00739975
R8281 GND.n1481 GND.n1480 0.00739975
R8282 GND.n1380 GND.n1379 0.00739975
R8283 GND.n4180 GND.n4179 0.00739975
R8284 GND.n3374 GND.n3373 0.00739975
R8285 GND.n3217 GND.n3216 0.00739975
R8286 GND.n2920 GND.n2919 0.00739975
R8287 GND.n2595 GND.n2594 0.00739975
R8288 GND.n2271 GND.n2270 0.00739975
R8289 GND.n2109 GND.n2108 0.00739975
R8290 GND.n1241 GND.n1240 0.00739975
R8291 GND.n7389 GND.n7388 0.00739975
R8292 GND.n3633 GND.n3632 0.00738379
R8293 GND.n4454 GND.n4453 0.00728191
R8294 GND.n4547 GND.n4545 0.00728191
R8295 GND.n5097 GND.n5096 0.00728191
R8296 GND.n6469 GND.n6465 0.00728191
R8297 GND.n6557 GND.n6556 0.00728191
R8298 GND.n6655 GND.n6654 0.00728191
R8299 GND.n3663 GND.n3662 0.00719643
R8300 GND.n4632 GND.n4630 0.00707895
R8301 GND.n4535 GND.n4534 0.00701596
R8302 GND.n5105 GND.n5104 0.00701596
R8303 GND.n6482 GND.n6480 0.00701596
R8304 GND.n6663 GND.n6662 0.00701596
R8305 GND.n3767 GND.n3765 0.00675
R8306 GND.n5561 GND.n5557 0.00675
R8307 GND.n5698 GND.n5694 0.00675
R8308 GND.n3694 GND.n3693 0.0066794
R8309 GND.n3662 GND.n3661 0.0066794
R8310 GND.n7339 GND.n2103 0.00666458
R8311 GND GND.n5531 0.00661702
R8312 GND.n5606 GND 0.00661702
R8313 GND GND.n5779 0.00661702
R8314 GND.n5683 GND 0.00661702
R8315 GND.n5732 GND 0.00661702
R8316 GND.n5754 GND 0.00661702
R8317 GND.n4482 GND 0.00661702
R8318 GND GND.n4503 0.00661702
R8319 GND.n5046 GND 0.00661702
R8320 GND GND.n5060 0.00661702
R8321 GND.n5143 GND 0.00661702
R8322 GND.n5165 GND 0.00661702
R8323 GND GND.n6439 0.00661702
R8324 GND.n6514 GND 0.00661702
R8325 GND.n6604 GND 0.00661702
R8326 GND GND.n6618 0.00661702
R8327 GND.n6701 GND 0.00661702
R8328 GND.n6723 GND 0.00661702
R8329 GND.n5557 GND.n5556 0.00648404
R8330 GND.n5694 GND.n5693 0.00648404
R8331 GND.n4589 GND.n4588 0.00647015
R8332 GND.n4593 GND.n4589 0.00631395
R8333 GND.n4539 GND.n4535 0.00621809
R8334 GND.n5109 GND.n5105 0.00621809
R8335 GND.n6480 GND.n6479 0.00621809
R8336 GND.n6667 GND.n6663 0.00621809
R8337 GND.n5028 GND 0.00609211
R8338 GND.n4972 GND 0.00609211
R8339 GND GND.n4684 0.00609211
R8340 GND.n4721 GND 0.00609211
R8341 GND.n3694 GND.n3692 0.00605556
R8342 GND.n5763 GND.n5762 0.00595213
R8343 GND.n4458 GND.n4454 0.00595213
R8344 GND.n4545 GND.n4434 0.00595213
R8345 GND.n5097 GND.n5055 0.00595213
R8346 GND.n6465 GND.n6464 0.00595213
R8347 GND.n6557 GND.n6527 0.00595213
R8348 GND.n6655 GND.n6613 0.00595213
R8349 GND.n5038 GND.n4945 0.00593478
R8350 GND.n4927 GND.n4923 0.00593421
R8351 GND.n1969 GND.n1967 0.00585714
R8352 GND.n1731 GND.n1729 0.00585714
R8353 GND.n1827 GND.n1825 0.00585714
R8354 GND.n6992 GND.n6990 0.00585714
R8355 GND.n2476 GND.n2474 0.00585714
R8356 GND.n2801 GND.n2799 0.00585714
R8357 GND.n7129 GND.n7127 0.00585714
R8358 GND.n4822 GND.n4820 0.00585714
R8359 GND.n5398 GND.n5396 0.00585714
R8360 GND.n5359 GND.n5357 0.00585714
R8361 GND.n5881 GND.n5879 0.00585714
R8362 GND.n6067 GND.n6065 0.00585714
R8363 GND.n6231 GND.n6229 0.00585714
R8364 GND.n6395 GND.n6393 0.00585714
R8365 GND.n680 GND.n678 0.00585714
R8366 GND.n7727 GND.n7725 0.00585714
R8367 GND.n4169 GND.n4166 0.00571186
R8368 GND.n3883 GND.n3881 0.00570833
R8369 GND.n5572 GND.n5571 0.00568617
R8370 GND.n5645 GND.n5619 0.00542021
R8371 GND.n5771 GND.n5769 0.00542021
R8372 GND.n5174 GND.n5173 0.00542021
R8373 GND.n6732 GND.n6731 0.00542021
R8374 GND GND.n1325 0.00541226
R8375 GND.n2102 GND 0.00541226
R8376 GND GND.n7337 0.00541226
R8377 GND GND.n7334 0.00541226
R8378 GND GND.n7331 0.00541226
R8379 GND GND.n7328 0.00541226
R8380 GND GND.n7325 0.00541226
R8381 GND GND.n7322 0.00541226
R8382 GND GND.n7318 0.00541226
R8383 GND GND.n7841 0.00541226
R8384 GND GND.n7838 0.00541226
R8385 GND GND.n7835 0.00541226
R8386 GND GND.n7832 0.00541226
R8387 GND GND.n7829 0.00541226
R8388 GND GND.n7826 0.00541226
R8389 GND.n4616 GND.n4606 0.00534496
R8390 GND.n2103 GND.n2102 0.00532736
R8391 GND GND.n4633 0.00510526
R8392 GND.n838 GND.n824 0.00507317
R8393 GND.n7491 GND.n7472 0.00507317
R8394 GND.n2080 GND.n2066 0.00507317
R8395 GND.n412 GND.n398 0.00507317
R8396 GND.n568 GND.n553 0.00507317
R8397 GND.n259 GND.n244 0.00507317
R8398 GND.n107 GND.n83 0.00507317
R8399 GND.n1440 GND.n1425 0.00507317
R8400 GND.n4267 GND.n4252 0.00507317
R8401 GND.n3464 GND.n3449 0.00507317
R8402 GND.n3306 GND.n3291 0.00507317
R8403 GND.n3010 GND.n2995 0.00507317
R8404 GND.n2686 GND.n2671 0.00507317
R8405 GND.n2361 GND.n2346 0.00507317
R8406 GND.n2203 GND.n2188 0.00507317
R8407 GND.n1322 GND.n1307 0.00507317
R8408 GND.n4629 GND.n4628 0.00505426
R8409 GND.n5029 GND 0.00502899
R8410 GND.n7085 GND.n4272 0.00498679
R8411 GND.n5619 GND.n5615 0.0048883
R8412 GND.n5772 GND.n5771 0.0048883
R8413 GND.n5173 GND.n5171 0.0048883
R8414 GND.n6731 GND.n6729 0.0048883
R8415 GND.n3641 GND.n3640 0.00476136
R8416 GND.n1927 GND.n1925 0.00466667
R8417 GND.n1585 GND.n1583 0.00466667
R8418 GND.n1694 GND.n1692 0.00466667
R8419 GND.n1776 GND.n1774 0.00466667
R8420 GND.n6902 GND.n6900 0.00466667
R8421 GND.n6941 GND.n6939 0.00466667
R8422 GND.n2370 GND.n2368 0.00466667
R8423 GND.n2425 GND.n2423 0.00466667
R8424 GND.n2695 GND.n2693 0.00466667
R8425 GND.n2750 GND.n2748 0.00466667
R8426 GND.n3019 GND.n3017 0.00466667
R8427 GND.n3074 GND.n3072 0.00466667
R8428 GND.n7092 GND.n7090 0.00466667
R8429 GND.n7174 GND.n7172 0.00466667
R8430 GND.n4787 GND.n4785 0.00466667
R8431 GND.n4867 GND.n4865 0.00466667
R8432 GND.n5269 GND.n5267 0.00466667
R8433 GND.n5308 GND.n5306 0.00466667
R8434 GND.n5791 GND.n5789 0.00466667
R8435 GND.n5830 GND.n5828 0.00466667
R8436 GND.n5958 GND.n5956 0.00466667
R8437 GND.n6013 GND.n6011 0.00466667
R8438 GND.n6125 GND.n6123 0.00466667
R8439 GND.n6177 GND.n6175 0.00466667
R8440 GND.n6289 GND.n6287 0.00466667
R8441 GND.n6341 GND.n6339 0.00466667
R8442 GND.n577 GND.n575 0.00466667
R8443 GND.n629 GND.n627 0.00466667
R8444 GND.n7620 GND.n7618 0.00466667
R8445 GND.n7676 GND.n7674 0.00466667
R8446 GND.n7500 GND.n7498 0.00466667
R8447 GND.n7545 GND.n7543 0.00466667
R8448 GND.n4971 GND 0.00466667
R8449 GND.n5571 GND.n5567 0.00462234
R8450 GND.n4606 GND.n4605 0.00456977
R8451 GND.n6759 GND 0.00456173
R8452 GND.n4586 GND.n4585 0.00454478
R8453 GND.n3704 GND.n3703 0.00438796
R8454 GND.n3719 GND.n3718 0.00438796
R8455 GND.n3734 GND.n3733 0.00438796
R8456 GND.n3749 GND.n3748 0.00438796
R8457 GND.n3765 GND.n3764 0.00438796
R8458 GND.n3783 GND.n3782 0.00438796
R8459 GND.n3798 GND.n3797 0.00438796
R8460 GND.n3813 GND.n3812 0.00438796
R8461 GND.n3828 GND.n3827 0.00438796
R8462 GND.n3853 GND.n3852 0.00438796
R8463 GND.n3872 GND.n3871 0.00438796
R8464 GND.n3892 GND.n3891 0.00438796
R8465 GND.n3907 GND.n3906 0.00438796
R8466 GND.n3922 GND.n3921 0.00438796
R8467 GND.n3937 GND.n3936 0.00438796
R8468 GND.n3952 GND.n3951 0.00438796
R8469 GND.n3969 GND.n3968 0.00438796
R8470 GND.n3984 GND.n3983 0.00438796
R8471 GND.n3999 GND.n3998 0.00438796
R8472 GND.n4014 GND.n4013 0.00438796
R8473 GND.n4029 GND.n4028 0.00438796
R8474 GND.n3652 GND.n3651 0.00438796
R8475 GND.n4021 GND.n4020 0.00438796
R8476 GND.n4005 GND.n4004 0.00438796
R8477 GND.n3990 GND.n3989 0.00438796
R8478 GND.n3975 GND.n3974 0.00438796
R8479 GND.n3960 GND.n3959 0.00438796
R8480 GND.n3943 GND.n3942 0.00438796
R8481 GND.n3928 GND.n3927 0.00438796
R8482 GND.n3913 GND.n3912 0.00438796
R8483 GND.n3898 GND.n3897 0.00438796
R8484 GND.n3881 GND.n3880 0.00438796
R8485 GND.n3862 GND.n3861 0.00438796
R8486 GND.n3844 GND.n3843 0.00438796
R8487 GND.n3819 GND.n3818 0.00438796
R8488 GND.n3804 GND.n3803 0.00438796
R8489 GND.n3789 GND.n3788 0.00438796
R8490 GND.n3774 GND.n3773 0.00438796
R8491 GND.n3755 GND.n3754 0.00438796
R8492 GND.n3740 GND.n3739 0.00438796
R8493 GND.n3725 GND.n3724 0.00438796
R8494 GND.n3710 GND.n3709 0.00438796
R8495 GND.n5762 GND.n5760 0.00435638
R8496 GND.n4494 GND.n4434 0.00435638
R8497 GND.n5055 GND.n5053 0.00435638
R8498 GND.n6527 GND.n6523 0.00435638
R8499 GND.n6613 GND.n6611 0.00435638
R8500 GND.n1917 GND.n1885 0.00425
R8501 GND.n1874 GND.n1711 0.00425
R8502 GND.n7032 GND.n6895 0.00425
R8503 GND.n2523 GND.n2387 0.00425
R8504 GND.n2848 GND.n2712 0.00425
R8505 GND.n3145 GND.n3036 0.00425
R8506 GND.n7245 GND.n7109 0.00425
R8507 GND.n4777 GND.n4751 0.00425
R8508 GND.n5424 GND.n5262 0.00425
R8509 GND.n5945 GND.n5917 0.00425
R8510 GND.n6114 GND.n5975 0.00425
R8511 GND.n6278 GND.n6142 0.00425
R8512 GND.n6587 GND.n6306 0.00425
R8513 GND.n727 GND.n594 0.00425
R8514 GND.n7774 GND.n7637 0.00425
R8515 GND.n7609 GND.n7517 0.00425
R8516 GND.n1230 GND.n1229 0.00420666
R8517 GND.n1229 GND.n1228 0.00420666
R8518 GND.n2255 GND.n2254 0.00420666
R8519 GND.n2254 GND.n2253 0.00420666
R8520 GND.n2579 GND.n2578 0.00420666
R8521 GND.n2578 GND.n2577 0.00420666
R8522 GND.n2904 GND.n2903 0.00420666
R8523 GND.n2903 GND.n2902 0.00420666
R8524 GND.n3201 GND.n3200 0.00420666
R8525 GND.n3200 GND.n3199 0.00420666
R8526 GND.n3358 GND.n3357 0.00420666
R8527 GND.n3357 GND.n3356 0.00420666
R8528 GND.n3516 GND.n3515 0.00420666
R8529 GND.n3515 GND.n3514 0.00420666
R8530 GND.n7306 GND.n7305 0.00420666
R8531 GND.n7305 GND.n7304 0.00420666
R8532 GND.n50 GND.n49 0.00420666
R8533 GND.n49 GND.n48 0.00420666
R8534 GND.n159 GND.n158 0.00420666
R8535 GND.n158 GND.n157 0.00420666
R8536 GND.n311 GND.n310 0.00420666
R8537 GND.n310 GND.n309 0.00420666
R8538 GND.n1682 GND.n1681 0.00420666
R8539 GND.n1681 GND.n1680 0.00420666
R8540 GND.n464 GND.n463 0.00420666
R8541 GND.n463 GND.n462 0.00420666
R8542 GND.n783 GND.n782 0.00420666
R8543 GND.n782 GND.n781 0.00420666
R8544 GND.n890 GND.n889 0.00420666
R8545 GND.n889 GND.n888 0.00420666
R8546 GND.n7818 GND.n7817 0.00420666
R8547 GND.n7817 GND.n7816 0.00420666
R8548 GND.n4540 GND.n4539 0.00409043
R8549 GND.n6479 GND.n6475 0.00409043
R8550 GND.n3875 GND.n3873 0.00397222
R8551 GND.n7725 GND.n7724 0.00396756
R8552 GND.n7555 GND.n7554 0.00396756
R8553 GND.n678 GND.n677 0.00396756
R8554 GND.n7686 GND.n7685 0.00396756
R8555 GND.n6393 GND.n6392 0.00396756
R8556 GND.n639 GND.n638 0.00396756
R8557 GND.n6229 GND.n6228 0.00396756
R8558 GND.n6351 GND.n6350 0.00396756
R8559 GND.n6065 GND.n6064 0.00396756
R8560 GND.n6187 GND.n6186 0.00396756
R8561 GND.n5879 GND.n5878 0.00396756
R8562 GND.n6023 GND.n6022 0.00396756
R8563 GND.n5357 GND.n5356 0.00396756
R8564 GND.n5840 GND.n5839 0.00396756
R8565 GND.n5396 GND.n5395 0.00396756
R8566 GND.n5318 GND.n5317 0.00396756
R8567 GND.n4820 GND.n4819 0.00396756
R8568 GND.n4877 GND.n4876 0.00396756
R8569 GND.n7127 GND.n7126 0.00396756
R8570 GND.n7184 GND.n7183 0.00396756
R8571 GND.n2799 GND.n2798 0.00396756
R8572 GND.n3084 GND.n3083 0.00396756
R8573 GND.n2474 GND.n2473 0.00396756
R8574 GND.n2760 GND.n2759 0.00396756
R8575 GND.n6990 GND.n6989 0.00396756
R8576 GND.n2435 GND.n2434 0.00396756
R8577 GND.n1825 GND.n1824 0.00396756
R8578 GND.n6951 GND.n6950 0.00396756
R8579 GND.n1729 GND.n1728 0.00396756
R8580 GND.n1786 GND.n1785 0.00396756
R8581 GND.n1967 GND.n1966 0.00396756
R8582 GND.n1595 GND.n1594 0.00396756
R8583 GND.n4669 GND.n4667 0.00396053
R8584 GND.n1920 GND.n1919 0.00395031
R8585 GND.n1877 GND.n1876 0.00395031
R8586 GND.n7030 GND.n7029 0.00395031
R8587 GND.n2526 GND.n2525 0.00395031
R8588 GND.n2851 GND.n2850 0.00395031
R8589 GND.n3148 GND.n3147 0.00395031
R8590 GND.n7248 GND.n7247 0.00395031
R8591 GND.n4780 GND.n4779 0.00395031
R8592 GND.n5422 GND.n5421 0.00395031
R8593 GND.n5948 GND.n5947 0.00395031
R8594 GND.n6117 GND.n6116 0.00395031
R8595 GND.n6281 GND.n6280 0.00395031
R8596 GND.n6590 GND.n6589 0.00395031
R8597 GND.n730 GND.n729 0.00395031
R8598 GND.n7777 GND.n7776 0.00395031
R8599 GND.n7612 GND.n7611 0.00395031
R8600 GND.n7724 GND.n7723 0.0039133
R8601 GND.n7723 GND.t205 0.0039133
R8602 GND.n7554 GND.n7553 0.0039133
R8603 GND.n7553 GND.t499 0.0039133
R8604 GND.n677 GND.n676 0.0039133
R8605 GND.n676 GND.t1217 0.0039133
R8606 GND.n7685 GND.n7684 0.0039133
R8607 GND.n7684 GND.t356 0.0039133
R8608 GND.n6392 GND.n6391 0.0039133
R8609 GND.n6391 GND.t197 0.0039133
R8610 GND.n638 GND.n637 0.0039133
R8611 GND.n637 GND.t128 0.0039133
R8612 GND.n6228 GND.n6227 0.0039133
R8613 GND.n6227 GND.t1208 0.0039133
R8614 GND.n6350 GND.n6349 0.0039133
R8615 GND.n6349 GND.t378 0.0039133
R8616 GND.n6064 GND.n6063 0.0039133
R8617 GND.n6063 GND.t765 0.0039133
R8618 GND.n6186 GND.n6185 0.0039133
R8619 GND.n6185 GND.t511 0.0039133
R8620 GND.n5878 GND.n5877 0.0039133
R8621 GND.n5877 GND.t99 0.0039133
R8622 GND.n6022 GND.n6021 0.0039133
R8623 GND.n6021 GND.t847 0.0039133
R8624 GND.n5356 GND.n5355 0.0039133
R8625 GND.n5355 GND.t1329 0.0039133
R8626 GND.n5839 GND.n5838 0.0039133
R8627 GND.n5838 GND.t1191 0.0039133
R8628 GND.n5395 GND.n5394 0.0039133
R8629 GND.n5394 GND.t1395 0.0039133
R8630 GND.n5317 GND.n5316 0.0039133
R8631 GND.n5316 GND.t813 0.0039133
R8632 GND.n4819 GND.n4818 0.0039133
R8633 GND.n4818 GND.t748 0.0039133
R8634 GND.n4876 GND.n4875 0.0039133
R8635 GND.n4875 GND.t179 0.0039133
R8636 GND.n7126 GND.n7125 0.0039133
R8637 GND.n7125 GND.t1264 0.0039133
R8638 GND.n7183 GND.n7182 0.0039133
R8639 GND.n7182 GND.t580 0.0039133
R8640 GND.n2798 GND.n2797 0.0039133
R8641 GND.n2797 GND.t6 0.0039133
R8642 GND.n3083 GND.n3082 0.0039133
R8643 GND.n3082 GND.t611 0.0039133
R8644 GND.n2473 GND.n2472 0.0039133
R8645 GND.n2472 GND.t1380 0.0039133
R8646 GND.n2759 GND.n2758 0.0039133
R8647 GND.n2758 GND.t25 0.0039133
R8648 GND.n6989 GND.n6988 0.0039133
R8649 GND.n6988 GND.t488 0.0039133
R8650 GND.n2434 GND.n2433 0.0039133
R8651 GND.n2433 GND.t137 0.0039133
R8652 GND.n1824 GND.n1823 0.0039133
R8653 GND.n1823 GND.t570 0.0039133
R8654 GND.n6950 GND.n6949 0.0039133
R8655 GND.n6949 GND.t487 0.0039133
R8656 GND.n1728 GND.n1727 0.0039133
R8657 GND.n1727 GND.t46 0.0039133
R8658 GND.n1785 GND.n1784 0.0039133
R8659 GND.n1784 GND.t368 0.0039133
R8660 GND.n1966 GND.n1965 0.0039133
R8661 GND.n1965 GND.t1290 0.0039133
R8662 GND.n1594 GND.n1593 0.0039133
R8663 GND.n1593 GND.t56 0.0039133
R8664 GND.n1916 GND.n1915 0.00390909
R8665 GND.n1913 GND.n1912 0.00390909
R8666 GND.n1873 GND.n1872 0.00390909
R8667 GND.n1870 GND.n1869 0.00390909
R8668 GND.n7033 GND.n6893 0.00390909
R8669 GND.n6891 GND.n6890 0.00390909
R8670 GND.n2522 GND.n2521 0.00390909
R8671 GND.n2519 GND.n2518 0.00390909
R8672 GND.n2847 GND.n2846 0.00390909
R8673 GND.n2844 GND.n2843 0.00390909
R8674 GND.n3144 GND.n3143 0.00390909
R8675 GND.n3141 GND.n3140 0.00390909
R8676 GND.n7244 GND.n7243 0.00390909
R8677 GND.n7241 GND.n7240 0.00390909
R8678 GND.n4776 GND.n4775 0.00390909
R8679 GND.n4773 GND.n4772 0.00390909
R8680 GND.n5425 GND.n5260 0.00390909
R8681 GND.n5258 GND.n5257 0.00390909
R8682 GND.n5944 GND.n5943 0.00390909
R8683 GND.n5941 GND.n5940 0.00390909
R8684 GND.n6113 GND.n6112 0.00390909
R8685 GND.n6110 GND.n6109 0.00390909
R8686 GND.n6277 GND.n6276 0.00390909
R8687 GND.n6274 GND.n6273 0.00390909
R8688 GND.n6586 GND.n6585 0.00390909
R8689 GND.n6583 GND.n6582 0.00390909
R8690 GND.n726 GND.n725 0.00390909
R8691 GND.n723 GND.n722 0.00390909
R8692 GND.n7773 GND.n7772 0.00390909
R8693 GND.n7770 GND.n7769 0.00390909
R8694 GND.n7608 GND.n7607 0.00390909
R8695 GND.n7605 GND.n7604 0.00390909
R8696 GND.n5693 GND.n5691 0.00382447
R8697 GND.n5104 GND.n5102 0.00379255
R8698 GND.n6662 GND.n6660 0.00379255
R8699 GND.n4169 GND.n4168 0.00377331
R8700 GND.n5562 GND.n5561 0.00355851
R8701 GND.n4453 GND.n4449 0.0035266
R8702 GND.n6470 GND.n6469 0.0035266
R8703 GND.n7576 GND.n7575 0.0034846
R8704 GND.n7740 GND.n7739 0.0034846
R8705 GND.n693 GND.n692 0.0034846
R8706 GND.n6408 GND.n6407 0.0034846
R8707 GND.n6244 GND.n6243 0.0034846
R8708 GND.n6080 GND.n6079 0.0034846
R8709 GND.n5894 GND.n5893 0.0034846
R8710 GND.n5372 GND.n5371 0.0034846
R8711 GND.n4904 GND.n4903 0.0034846
R8712 GND.n7211 GND.n7210 0.0034846
R8713 GND.n3111 GND.n3110 0.0034846
R8714 GND.n2814 GND.n2813 0.0034846
R8715 GND.n2489 GND.n2488 0.0034846
R8716 GND.n7005 GND.n7004 0.0034846
R8717 GND.n1840 GND.n1839 0.0034846
R8718 GND.n1622 GND.n1621 0.0034846
R8719 GND.n7575 GND.n7574 0.00343883
R8720 GND.n7574 GND.n7573 0.00343883
R8721 GND.n7736 GND.n7735 0.00343883
R8722 GND.n7737 GND.n7736 0.00343883
R8723 GND.n7739 GND.n7738 0.00343883
R8724 GND.n7738 GND.n7737 0.00343883
R8725 GND.n689 GND.n688 0.00343883
R8726 GND.n690 GND.n689 0.00343883
R8727 GND.n692 GND.n691 0.00343883
R8728 GND.n691 GND.n690 0.00343883
R8729 GND.n6404 GND.n6403 0.00343883
R8730 GND.n6405 GND.n6404 0.00343883
R8731 GND.n6407 GND.n6406 0.00343883
R8732 GND.n6406 GND.n6405 0.00343883
R8733 GND.n6240 GND.n6239 0.00343883
R8734 GND.n6241 GND.n6240 0.00343883
R8735 GND.n6243 GND.n6242 0.00343883
R8736 GND.n6242 GND.n6241 0.00343883
R8737 GND.n6076 GND.n6075 0.00343883
R8738 GND.n6077 GND.n6076 0.00343883
R8739 GND.n6079 GND.n6078 0.00343883
R8740 GND.n6078 GND.n6077 0.00343883
R8741 GND.n5890 GND.n5889 0.00343883
R8742 GND.n5891 GND.n5890 0.00343883
R8743 GND.n5893 GND.n5892 0.00343883
R8744 GND.n5892 GND.n5891 0.00343883
R8745 GND.n5368 GND.n5367 0.00343883
R8746 GND.n5369 GND.n5368 0.00343883
R8747 GND.n5371 GND.n5370 0.00343883
R8748 GND.n5370 GND.n5369 0.00343883
R8749 GND.n4901 GND.n4900 0.00343883
R8750 GND.n4903 GND.n4902 0.00343883
R8751 GND.n4902 GND.n4901 0.00343883
R8752 GND.n7208 GND.n7207 0.00343883
R8753 GND.n7210 GND.n7209 0.00343883
R8754 GND.n7209 GND.n7208 0.00343883
R8755 GND.n3108 GND.n3107 0.00343883
R8756 GND.n3110 GND.n3109 0.00343883
R8757 GND.n3109 GND.n3108 0.00343883
R8758 GND.n2810 GND.n2809 0.00343883
R8759 GND.n2811 GND.n2810 0.00343883
R8760 GND.n2813 GND.n2812 0.00343883
R8761 GND.n2812 GND.n2811 0.00343883
R8762 GND.n2485 GND.n2484 0.00343883
R8763 GND.n2486 GND.n2485 0.00343883
R8764 GND.n2488 GND.n2487 0.00343883
R8765 GND.n2487 GND.n2486 0.00343883
R8766 GND.n7001 GND.n7000 0.00343883
R8767 GND.n7002 GND.n7001 0.00343883
R8768 GND.n7004 GND.n7003 0.00343883
R8769 GND.n7003 GND.n7002 0.00343883
R8770 GND.n1836 GND.n1835 0.00343883
R8771 GND.n1837 GND.n1836 0.00343883
R8772 GND.n1839 GND.n1838 0.00343883
R8773 GND.n1838 GND.n1837 0.00343883
R8774 GND.n1619 GND.n1618 0.00343883
R8775 GND.n1621 GND.n1620 0.00343883
R8776 GND.n1620 GND.n1619 0.00343883
R8777 GND.n1978 GND.n1977 0.00343883
R8778 GND.n1979 GND.n1978 0.00343883
R8779 GND GND.n6841 0.00340123
R8780 GND GND.n6759 0.00340123
R8781 GND.n4961 GND 0.00327778
R8782 GND.n4954 GND 0.00327778
R8783 GND.n7322 GND.n7321 0.00320477
R8784 GND.n5029 GND.n5028 0.00313158
R8785 GND.n1940 GND.n1939 0.00308428
R8786 GND.n1707 GND.n1706 0.00308428
R8787 GND.n6915 GND.n6914 0.00308428
R8788 GND.n2383 GND.n2382 0.00308428
R8789 GND.n2708 GND.n2707 0.00308428
R8790 GND.n3032 GND.n3031 0.00308428
R8791 GND.n7105 GND.n7104 0.00308428
R8792 GND.n4800 GND.n4799 0.00308428
R8793 GND.n5282 GND.n5281 0.00308428
R8794 GND.n5804 GND.n5803 0.00308428
R8795 GND.n5971 GND.n5970 0.00308428
R8796 GND.n6138 GND.n6137 0.00308428
R8797 GND.n6302 GND.n6301 0.00308428
R8798 GND.n590 GND.n589 0.00308428
R8799 GND.n7633 GND.n7632 0.00308428
R8800 GND.n7513 GND.n7512 0.00308428
R8801 GND.n4425 GND.n4424 0.00307458
R8802 GND.n5742 GND.n5740 0.0030266
R8803 GND.n4548 GND.n4547 0.0030266
R8804 GND.n5096 GND.n5092 0.0030266
R8805 GND.n6556 GND.n6554 0.0030266
R8806 GND.n6654 GND.n6650 0.0030266
R8807 GND.n1885 GND.n1884 0.003
R8808 GND.n1711 GND.n1710 0.003
R8809 GND.n6895 GND.n6894 0.003
R8810 GND.n2387 GND.n2386 0.003
R8811 GND.n2712 GND.n2711 0.003
R8812 GND.n3036 GND.n3035 0.003
R8813 GND.n7109 GND.n7108 0.003
R8814 GND.n4751 GND.n4750 0.003
R8815 GND.n5262 GND.n5261 0.003
R8816 GND.n5917 GND.n5916 0.003
R8817 GND.n5975 GND.n5974 0.003
R8818 GND.n6142 GND.n6141 0.003
R8819 GND.n6306 GND.n6305 0.003
R8820 GND.n594 GND.n593 0.003
R8821 GND.n7637 GND.n7636 0.003
R8822 GND.n7517 GND.n7516 0.003
R8823 GND.n3698 GND.n3697 0.00299232
R8824 GND.n4630 GND.n4629 0.00292248
R8825 GND.n6838 GND.n6837 0.00290385
R8826 GND.n7083 GND.n7082 0.00290385
R8827 GND.n4975 GND.n4973 0.00280263
R8828 GND.n5444 GND.n5441 0.00277946
R8829 GND.n6849 GND.n6846 0.00277946
R8830 GND.n5532 GND 0.00276064
R8831 GND.n5603 GND 0.00276064
R8832 GND.n5780 GND 0.00276064
R8833 GND.n5680 GND 0.00276064
R8834 GND.n5729 GND 0.00276064
R8835 GND GND.n5742 0.00276064
R8836 GND.n5757 GND 0.00276064
R8837 GND.n5745 GND 0.00276064
R8838 GND.n4479 GND 0.00276064
R8839 GND.n4504 GND 0.00276064
R8840 GND.n5043 GND 0.00276064
R8841 GND.n5061 GND 0.00276064
R8842 GND.n5140 GND 0.00276064
R8843 GND GND.n5153 0.00276064
R8844 GND.n5168 GND 0.00276064
R8845 GND.n5156 GND 0.00276064
R8846 GND.n6440 GND 0.00276064
R8847 GND.n6511 GND 0.00276064
R8848 GND.n6601 GND 0.00276064
R8849 GND.n6619 GND 0.00276064
R8850 GND.n6698 GND 0.00276064
R8851 GND GND.n6711 0.00276064
R8852 GND.n6726 GND 0.00276064
R8853 GND.n6714 GND 0.00276064
R8854 GND.n1434 GND.n1433 0.00266776
R8855 GND.n3458 GND.n3457 0.00266776
R8856 GND.n3004 GND.n3003 0.00266776
R8857 GND.n2355 GND.n2354 0.00266776
R8858 GND.n2197 GND.n2196 0.00266776
R8859 GND.n2680 GND.n2679 0.00266776
R8860 GND.n3300 GND.n3299 0.00266776
R8861 GND.n4261 GND.n4260 0.00266776
R8862 GND.n101 GND.n100 0.00266776
R8863 GND.n253 GND.n252 0.00266776
R8864 GND.n562 GND.n561 0.00266776
R8865 GND.n7485 GND.n7484 0.00266776
R8866 GND.n1595 GND.n1591 0.00258333
R8867 GND.n1786 GND.n1782 0.00258333
R8868 GND.n6951 GND.n6947 0.00258333
R8869 GND.n2435 GND.n2431 0.00258333
R8870 GND.n2760 GND.n2756 0.00258333
R8871 GND.n3084 GND.n3080 0.00258333
R8872 GND.n7184 GND.n7180 0.00258333
R8873 GND.n4877 GND.n4873 0.00258333
R8874 GND.n5318 GND.n5314 0.00258333
R8875 GND.n5840 GND.n5836 0.00258333
R8876 GND.n6023 GND.n6019 0.00258333
R8877 GND.n6187 GND.n6183 0.00258333
R8878 GND.n6351 GND.n6347 0.00258333
R8879 GND.n639 GND.n635 0.00258333
R8880 GND.n7686 GND.n7682 0.00258333
R8881 GND.n7555 GND.n7551 0.00258333
R8882 GND.n4061 GND.n4060 0.00253688
R8883 GND.n4052 GND.n4051 0.00253688
R8884 GND.n4035 GND.n4034 0.00250907
R8885 GND.n4023 GND.n4022 0.00250907
R8886 GND.n4007 GND.n4006 0.00250907
R8887 GND.n3992 GND.n3991 0.00250907
R8888 GND.n3977 GND.n3976 0.00250907
R8889 GND.n3962 GND.n3961 0.00250907
R8890 GND.n3945 GND.n3944 0.00250907
R8891 GND.n3930 GND.n3929 0.00250907
R8892 GND.n3915 GND.n3914 0.00250907
R8893 GND.n3900 GND.n3899 0.00250907
R8894 GND.n3885 GND.n3884 0.00250907
R8895 GND.n3864 GND.n3863 0.00250907
R8896 GND.n3846 GND.n3845 0.00250907
R8897 GND.n3821 GND.n3820 0.00250907
R8898 GND.n3806 GND.n3805 0.00250907
R8899 GND.n3791 GND.n3790 0.00250907
R8900 GND.n3776 GND.n3775 0.00250907
R8901 GND.n3757 GND.n3756 0.00250907
R8902 GND.n3742 GND.n3741 0.00250907
R8903 GND.n3727 GND.n3726 0.00250907
R8904 GND.n3712 GND.n3711 0.00250907
R8905 GND.n3702 GND.n3701 0.00250907
R8906 GND.n3717 GND.n3716 0.00250907
R8907 GND.n3732 GND.n3731 0.00250907
R8908 GND.n3747 GND.n3746 0.00250907
R8909 GND.n3762 GND.n3761 0.00250907
R8910 GND.n3781 GND.n3780 0.00250907
R8911 GND.n3796 GND.n3795 0.00250907
R8912 GND.n3811 GND.n3810 0.00250907
R8913 GND.n3826 GND.n3825 0.00250907
R8914 GND.n3851 GND.n3850 0.00250907
R8915 GND.n3869 GND.n3868 0.00250907
R8916 GND.n3890 GND.n3889 0.00250907
R8917 GND.n3905 GND.n3904 0.00250907
R8918 GND.n3920 GND.n3919 0.00250907
R8919 GND.n3935 GND.n3934 0.00250907
R8920 GND.n3950 GND.n3949 0.00250907
R8921 GND.n3967 GND.n3966 0.00250907
R8922 GND.n3982 GND.n3981 0.00250907
R8923 GND.n3997 GND.n3996 0.00250907
R8924 GND.n4012 GND.n4011 0.00250907
R8925 GND.n4027 GND.n4026 0.00250907
R8926 GND.n4031 GND.n4030 0.00250907
R8927 GND.n5644 GND.n5642 0.00249468
R8928 GND.n5649 GND.n5506 0.00249468
R8929 GND.n5153 GND.n5151 0.00249468
R8930 GND.n6711 GND.n6709 0.00249468
R8931 GND.n3700 GND.t1360 0.00247763
R8932 GND.n3715 GND.t834 0.00247763
R8933 GND.n3730 GND.t1357 0.00247763
R8934 GND.n3745 GND.t731 0.00247763
R8935 GND.n3760 GND.t724 0.00247763
R8936 GND.n3779 GND.t1361 0.00247763
R8937 GND.n3794 GND.t729 0.00247763
R8938 GND.n3809 GND.t832 0.00247763
R8939 GND.n3824 GND.t723 0.00247763
R8940 GND.n3849 GND.t730 0.00247763
R8941 GND.n3867 GND.t727 0.00247763
R8942 GND.n3888 GND.t1359 0.00247763
R8943 GND.n3903 GND.t725 0.00247763
R8944 GND.n3918 GND.t835 0.00247763
R8945 GND.n3933 GND.t721 0.00247763
R8946 GND.n3948 GND.t1356 0.00247763
R8947 GND.n3965 GND.t833 0.00247763
R8948 GND.n3980 GND.t726 0.00247763
R8949 GND.n3995 GND.t836 0.00247763
R8950 GND.n4010 GND.t722 0.00247763
R8951 GND.n4008 GND.n4007 0.00247763
R8952 GND.t722 GND.n4008 0.00247763
R8953 GND.n3993 GND.n3992 0.00247763
R8954 GND.t836 GND.n3993 0.00247763
R8955 GND.n3978 GND.n3977 0.00247763
R8956 GND.t726 GND.n3978 0.00247763
R8957 GND.n3963 GND.n3962 0.00247763
R8958 GND.t833 GND.n3963 0.00247763
R8959 GND.n3946 GND.n3945 0.00247763
R8960 GND.t1356 GND.n3946 0.00247763
R8961 GND.n3931 GND.n3930 0.00247763
R8962 GND.t721 GND.n3931 0.00247763
R8963 GND.n3916 GND.n3915 0.00247763
R8964 GND.t835 GND.n3916 0.00247763
R8965 GND.n3901 GND.n3900 0.00247763
R8966 GND.t725 GND.n3901 0.00247763
R8967 GND.n3886 GND.n3885 0.00247763
R8968 GND.t1359 GND.n3886 0.00247763
R8969 GND.n3865 GND.n3864 0.00247763
R8970 GND.t727 GND.n3865 0.00247763
R8971 GND.n3847 GND.n3846 0.00247763
R8972 GND.t730 GND.n3847 0.00247763
R8973 GND.n3822 GND.n3821 0.00247763
R8974 GND.t723 GND.n3822 0.00247763
R8975 GND.n3807 GND.n3806 0.00247763
R8976 GND.t832 GND.n3807 0.00247763
R8977 GND.n3792 GND.n3791 0.00247763
R8978 GND.t729 GND.n3792 0.00247763
R8979 GND.n3777 GND.n3776 0.00247763
R8980 GND.t1361 GND.n3777 0.00247763
R8981 GND.n3758 GND.n3757 0.00247763
R8982 GND.t724 GND.n3758 0.00247763
R8983 GND.n3743 GND.n3742 0.00247763
R8984 GND.t731 GND.n3743 0.00247763
R8985 GND.n3728 GND.n3727 0.00247763
R8986 GND.t1357 GND.n3728 0.00247763
R8987 GND.n3713 GND.n3712 0.00247763
R8988 GND.t834 GND.n3713 0.00247763
R8989 GND.n3699 GND.n3698 0.00247763
R8990 GND.t1360 GND.n3699 0.00247763
R8991 GND.n3701 GND.n3700 0.00247763
R8992 GND.n3716 GND.n3715 0.00247763
R8993 GND.n3731 GND.n3730 0.00247763
R8994 GND.n3746 GND.n3745 0.00247763
R8995 GND.n3761 GND.n3760 0.00247763
R8996 GND.n3780 GND.n3779 0.00247763
R8997 GND.n3795 GND.n3794 0.00247763
R8998 GND.n3810 GND.n3809 0.00247763
R8999 GND.n3825 GND.n3824 0.00247763
R9000 GND.n3850 GND.n3849 0.00247763
R9001 GND.n3868 GND.n3867 0.00247763
R9002 GND.n3889 GND.n3888 0.00247763
R9003 GND.n3904 GND.n3903 0.00247763
R9004 GND.n3919 GND.n3918 0.00247763
R9005 GND.n3934 GND.n3933 0.00247763
R9006 GND.n3949 GND.n3948 0.00247763
R9007 GND.n3966 GND.n3965 0.00247763
R9008 GND.n3981 GND.n3980 0.00247763
R9009 GND.n3996 GND.n3995 0.00247763
R9010 GND.n4011 GND.n4010 0.00247763
R9011 GND.n4026 GND.n4025 0.00247763
R9012 GND.n4025 GND.t1358 0.00247763
R9013 GND.n4024 GND.n4023 0.00247763
R9014 GND.t1358 GND.n4024 0.00247763
R9015 GND.n4034 GND.n4033 0.00247763
R9016 GND.n4033 GND.t1129 0.00247763
R9017 GND.t1129 GND.n4032 0.00247763
R9018 GND.n4032 GND.n4031 0.00247763
R9019 GND.n4971 GND 0.00247368
R9020 GND.n1919 GND.n1918 0.00245833
R9021 GND.n1876 GND.n1875 0.00245833
R9022 GND.n7031 GND.n7030 0.00245833
R9023 GND.n2525 GND.n2524 0.00245833
R9024 GND.n2850 GND.n2849 0.00245833
R9025 GND.n3147 GND.n3146 0.00245833
R9026 GND.n7247 GND.n7246 0.00245833
R9027 GND.n4779 GND.n4778 0.00245833
R9028 GND.n5423 GND.n5422 0.00245833
R9029 GND.n5947 GND.n5946 0.00245833
R9030 GND.n6116 GND.n6115 0.00245833
R9031 GND.n6280 GND.n6279 0.00245833
R9032 GND.n6589 GND.n6588 0.00245833
R9033 GND.n729 GND.n728 0.00245833
R9034 GND.n7776 GND.n7775 0.00245833
R9035 GND.n7611 GND.n7610 0.00245833
R9036 GND.n1622 GND.n1617 0.00228571
R9037 GND.n1840 GND.n1808 0.00228571
R9038 GND.n7005 GND.n6973 0.00228571
R9039 GND.n2489 GND.n2457 0.00228571
R9040 GND.n2814 GND.n2782 0.00228571
R9041 GND.n3111 GND.n3106 0.00228571
R9042 GND.n7211 GND.n7206 0.00228571
R9043 GND.n4904 GND.n4899 0.00228571
R9044 GND.n5372 GND.n5340 0.00228571
R9045 GND.n5894 GND.n5862 0.00228571
R9046 GND.n6080 GND.n6045 0.00228571
R9047 GND.n6244 GND.n6209 0.00228571
R9048 GND.n6408 GND.n6373 0.00228571
R9049 GND.n693 GND.n661 0.00228571
R9050 GND.n7740 GND.n7708 0.00228571
R9051 GND.n7576 GND.n7572 0.00228571
R9052 GND.n7376 GND 0.00217027
R9053 GND.n1372 GND 0.00217027
R9054 GND.n334 GND 0.00217027
R9055 GND.n487 GND 0.00217027
R9056 GND.n182 GND 0.00217027
R9057 GND.n1517 GND 0.00217027
R9058 GND.n1469 GND 0.00217027
R9059 GND.n4190 GND 0.00217027
R9060 GND.n3384 GND 0.00217027
R9061 GND.n3227 GND 0.00217027
R9062 GND.n2930 GND 0.00217027
R9063 GND.n2605 GND 0.00217027
R9064 GND.n2281 GND 0.00217027
R9065 GND.n2119 GND 0.00217027
R9066 GND.n1251 GND 0.00217027
R9067 GND.n7418 GND 0.00217027
R9068 GND.n6849 GND.n6848 0.00193331
R9069 GND.n5444 GND.n5443 0.00193331
R9070 GND.n3873 GND.n3872 0.00188889
R9071 GND.n3614 GND.n3613 0.00186977
R9072 GND.n3617 GND.n3614 0.00186977
R9073 GND.n3616 GND.n3615 0.00186977
R9074 GND.n3617 GND.n3616 0.00186977
R9075 GND.n3612 GND.n3611 0.00186977
R9076 GND.n3617 GND.n3612 0.00186977
R9077 GND.n7543 GND.n7542 0.00183506
R9078 GND.n7674 GND.n7673 0.00183506
R9079 GND.n627 GND.n626 0.00183506
R9080 GND.n6339 GND.n6338 0.00183506
R9081 GND.n6175 GND.n6174 0.00183506
R9082 GND.n6011 GND.n6010 0.00183506
R9083 GND.n5828 GND.n5827 0.00183506
R9084 GND.n5306 GND.n5305 0.00183506
R9085 GND.n4865 GND.n4864 0.00183506
R9086 GND.n7172 GND.n7171 0.00183506
R9087 GND.n3072 GND.n3071 0.00183506
R9088 GND.n2748 GND.n2747 0.00183506
R9089 GND.n2423 GND.n2422 0.00183506
R9090 GND.n6939 GND.n6938 0.00183506
R9091 GND.n1774 GND.n1773 0.00183506
R9092 GND.n1583 GND.n1582 0.00183506
R9093 GND.n7542 GND.n7541 0.00181454
R9094 GND.n7716 GND.n7715 0.00181454
R9095 GND.n7715 GND.n7714 0.00181454
R9096 GND.n7673 GND.n7672 0.00181454
R9097 GND.n669 GND.n668 0.00181454
R9098 GND.n668 GND.n667 0.00181454
R9099 GND.n626 GND.n625 0.00181454
R9100 GND.n6384 GND.n6383 0.00181454
R9101 GND.n6383 GND.n6382 0.00181454
R9102 GND.n6338 GND.n6337 0.00181454
R9103 GND.n6220 GND.n6219 0.00181454
R9104 GND.n6219 GND.n6218 0.00181454
R9105 GND.n6174 GND.n6173 0.00181454
R9106 GND.n6056 GND.n6055 0.00181454
R9107 GND.n6055 GND.n6054 0.00181454
R9108 GND.n6010 GND.n6009 0.00181454
R9109 GND.n5870 GND.n5869 0.00181454
R9110 GND.n5869 GND.n5868 0.00181454
R9111 GND.n5827 GND.n5826 0.00181454
R9112 GND.n5348 GND.n5347 0.00181454
R9113 GND.n5347 GND.n5346 0.00181454
R9114 GND.n5305 GND.n5304 0.00181454
R9115 GND.n5387 GND.n5386 0.00181454
R9116 GND.n5386 GND.n5385 0.00181454
R9117 GND.n4864 GND.n4863 0.00181454
R9118 GND.n4811 GND.n4810 0.00181454
R9119 GND.n4810 GND.n4809 0.00181454
R9120 GND.n7171 GND.n7170 0.00181454
R9121 GND.n7118 GND.n7117 0.00181454
R9122 GND.n7117 GND.n7116 0.00181454
R9123 GND.n3071 GND.n3070 0.00181454
R9124 GND.n2790 GND.n2789 0.00181454
R9125 GND.n2789 GND.n2788 0.00181454
R9126 GND.n2747 GND.n2746 0.00181454
R9127 GND.n2465 GND.n2464 0.00181454
R9128 GND.n2464 GND.n2463 0.00181454
R9129 GND.n2422 GND.n2421 0.00181454
R9130 GND.n6981 GND.n6980 0.00181454
R9131 GND.n6980 GND.n6979 0.00181454
R9132 GND.n6938 GND.n6937 0.00181454
R9133 GND.n1816 GND.n1815 0.00181454
R9134 GND.n1815 GND.n1814 0.00181454
R9135 GND.n1773 GND.n1772 0.00181454
R9136 GND.n1720 GND.n1719 0.00181454
R9137 GND.n1719 GND.n1718 0.00181454
R9138 GND.n1582 GND.n1581 0.00181454
R9139 GND.n1958 GND.n1957 0.00181454
R9140 GND.n1957 GND.n1956 0.00181454
R9141 GND.n5453 GND.n5447 0.00175
R9142 GND.n5457 GND.n5456 0.00175
R9143 GND.n5459 GND.n5445 0.00175
R9144 GND.n6858 GND.n6852 0.00175
R9145 GND.n6862 GND.n6861 0.00175
R9146 GND.n6864 GND.n6850 0.00175
R9147 GND.n7820 GND.n7783 0.00174202
R9148 GND.n892 GND.n842 0.00174202
R9149 GND.n785 GND.n735 0.00174202
R9150 GND.n466 GND.n416 0.00174202
R9151 GND.n1684 GND.n1626 0.00174202
R9152 GND.n313 GND.n263 0.00174202
R9153 GND.n161 GND.n111 0.00174202
R9154 GND.n52 GND.n2 0.00174202
R9155 GND.n7308 GND.n7258 0.00174202
R9156 GND.n3518 GND.n3468 0.00174202
R9157 GND.n3360 GND.n3310 0.00174202
R9158 GND.n3203 GND.n3153 0.00174202
R9159 GND.n2906 GND.n2856 0.00174202
R9160 GND.n2581 GND.n2531 0.00174202
R9161 GND.n2257 GND.n2207 0.00174202
R9162 GND.n1232 GND.n1182 0.00174202
R9163 GND.n3529 GND.n3528 0.00172549
R9164 GND.n408 GND.n406 0.001708
R9165 GND.n1317 GND.n1315 0.001708
R9166 GND.n2076 GND.n2074 0.001708
R9167 GND.n834 GND.n832 0.001708
R9168 GND.n5524 GND.n5508 0.00169681
R9169 GND.n5174 GND 0.00169681
R9170 GND.n6732 GND 0.00169681
R9171 GND.n4120 GND.n4115 0.00166525
R9172 GND.n7252 GND.n7251 0.0016471
R9173 GND.n1900 GND.n1897 0.00163636
R9174 GND.n1857 GND.n1854 0.00163636
R9175 GND.n7038 GND.n7037 0.00163636
R9176 GND.n2506 GND.n2503 0.00163636
R9177 GND.n2831 GND.n2828 0.00163636
R9178 GND.n3128 GND.n3125 0.00163636
R9179 GND.n7228 GND.n7225 0.00163636
R9180 GND.n4760 GND.n4757 0.00163636
R9181 GND.n5430 GND.n5429 0.00163636
R9182 GND.n5928 GND.n5925 0.00163636
R9183 GND.n6097 GND.n6094 0.00163636
R9184 GND.n6261 GND.n6258 0.00163636
R9185 GND.n6570 GND.n6567 0.00163636
R9186 GND.n710 GND.n707 0.00163636
R9187 GND.n7757 GND.n7754 0.00163636
R9188 GND.n7592 GND.n7589 0.00163636
R9189 GND.n1933 GND.n1931 0.00154167
R9190 GND.n1700 GND.n1698 0.00154167
R9191 GND.n6908 GND.n6906 0.00154167
R9192 GND.n2376 GND.n2374 0.00154167
R9193 GND.n2701 GND.n2699 0.00154167
R9194 GND.n3025 GND.n3023 0.00154167
R9195 GND.n7098 GND.n7096 0.00154167
R9196 GND.n4793 GND.n4791 0.00154167
R9197 GND.n5275 GND.n5273 0.00154167
R9198 GND.n5797 GND.n5795 0.00154167
R9199 GND.n5964 GND.n5962 0.00154167
R9200 GND.n6131 GND.n6129 0.00154167
R9201 GND.n6295 GND.n6293 0.00154167
R9202 GND.n583 GND.n581 0.00154167
R9203 GND.n7626 GND.n7624 0.00154167
R9204 GND.n7506 GND.n7504 0.00154167
R9205 GND.n7491 GND.n7490 0.00150729
R9206 GND.n568 GND.n567 0.00150729
R9207 GND.n259 GND.n258 0.00150729
R9208 GND.n107 GND.n106 0.00150729
R9209 GND.n1440 GND.n1439 0.00150729
R9210 GND.n4267 GND.n4266 0.00150729
R9211 GND.n3464 GND.n3463 0.00150729
R9212 GND.n3306 GND.n3305 0.00150729
R9213 GND.n3010 GND.n3009 0.00150729
R9214 GND.n2686 GND.n2685 0.00150729
R9215 GND.n2361 GND.n2360 0.00150729
R9216 GND.n2203 GND.n2202 0.00150729
R9217 GND.n1322 GND.n1321 0.00150729
R9218 GND.n7085 GND.n7084 0.00150166
R9219 GND.n6840 GND.n6839 0.00150121
R9220 GND.n4661 GND.n4633 0.00148684
R9221 GND.n7435 GND.n7369 0.00139286
R9222 GND.n1988 GND.n1365 0.00139286
R9223 GND.n332 GND.n330 0.00139286
R9224 GND.n485 GND.n483 0.00139286
R9225 GND.n180 GND.n178 0.00139286
R9226 GND.n1515 GND.n1487 0.00139286
R9227 GND.n1467 GND.n1386 0.00139286
R9228 GND.n4188 GND.n4186 0.00139286
R9229 GND.n3382 GND.n3380 0.00139286
R9230 GND.n3225 GND.n3223 0.00139286
R9231 GND.n2928 GND.n2926 0.00139286
R9232 GND.n2603 GND.n2601 0.00139286
R9233 GND.n2279 GND.n2277 0.00139286
R9234 GND.n2117 GND.n2115 0.00139286
R9235 GND.n1249 GND.n1247 0.00139286
R9236 GND.n7416 GND.n7395 0.00139286
R9237 GND.n7433 GND.n7432 0.00138653
R9238 GND.n1986 GND.n1985 0.00138653
R9239 GND.n339 GND.n333 0.00138653
R9240 GND.n492 GND.n486 0.00138653
R9241 GND.n187 GND.n181 0.00138653
R9242 GND.n1522 GND.n1516 0.00138653
R9243 GND.n1474 GND.n1468 0.00138653
R9244 GND.n4195 GND.n4189 0.00138653
R9245 GND.n3389 GND.n3383 0.00138653
R9246 GND.n3232 GND.n3226 0.00138653
R9247 GND.n2935 GND.n2929 0.00138653
R9248 GND.n2610 GND.n2604 0.00138653
R9249 GND.n2286 GND.n2280 0.00138653
R9250 GND.n2124 GND.n2118 0.00138653
R9251 GND.n1256 GND.n1250 0.00138653
R9252 GND.n7423 GND.n7417 0.00138653
R9253 GND.n7350 GND.n7349 0.00132676
R9254 GND.n1142 GND.n1139 0.00132676
R9255 GND.n1126 GND.n1123 0.00132676
R9256 GND.n1118 GND.n1115 0.00132676
R9257 GND.n7312 GND.n1110 0.00132676
R9258 GND.n4170 GND.n1105 0.00132676
R9259 GND.n3364 GND.n1100 0.00132676
R9260 GND.n3207 GND.n1095 0.00132676
R9261 GND.n2910 GND.n1090 0.00132676
R9262 GND.n2585 GND.n1085 0.00132676
R9263 GND.n2261 GND.n1080 0.00132676
R9264 GND.n2095 GND.n2094 0.00132676
R9265 GND.n1134 GND.n1131 0.00132676
R9266 GND.n1150 GND.n1147 0.00132676
R9267 GND.n2092 GND.n2089 0.0013267
R9268 GND.n7347 GND.n7344 0.0013267
R9269 GND.n7531 GND.t519 0.00131092
R9270 GND.n7532 GND.n7531 0.00131092
R9271 GND.n7653 GND.n7652 0.00131092
R9272 GND.t436 GND.n7653 0.00131092
R9273 GND.n7662 GND.t436 0.00131092
R9274 GND.n7663 GND.n7662 0.00131092
R9275 GND.n610 GND.n609 0.00131092
R9276 GND.t200 GND.n610 0.00131092
R9277 GND.n618 GND.t200 0.00131092
R9278 GND.n619 GND.n618 0.00131092
R9279 GND.n6322 GND.n6321 0.00131092
R9280 GND.t187 GND.n6322 0.00131092
R9281 GND.n6330 GND.t187 0.00131092
R9282 GND.n6331 GND.n6330 0.00131092
R9283 GND.n6158 GND.n6157 0.00131092
R9284 GND.t156 GND.n6158 0.00131092
R9285 GND.n6166 GND.t156 0.00131092
R9286 GND.n6167 GND.n6166 0.00131092
R9287 GND.n5991 GND.n5990 0.00131092
R9288 GND.t170 GND.n5991 0.00131092
R9289 GND.n5999 GND.t170 0.00131092
R9290 GND.n6000 GND.n5999 0.00131092
R9291 GND.n5808 GND.n5807 0.00131092
R9292 GND.t31 GND.n5808 0.00131092
R9293 GND.n5816 GND.t31 0.00131092
R9294 GND.n5817 GND.n5816 0.00131092
R9295 GND.n5286 GND.n5285 0.00131092
R9296 GND.t821 GND.n5286 0.00131092
R9297 GND.n5294 GND.t821 0.00131092
R9298 GND.n5295 GND.n5294 0.00131092
R9299 GND.n4845 GND.n4844 0.00131092
R9300 GND.t526 GND.n4845 0.00131092
R9301 GND.n4853 GND.t526 0.00131092
R9302 GND.n4854 GND.n4853 0.00131092
R9303 GND.n7152 GND.n7151 0.00131092
R9304 GND.t183 GND.n7152 0.00131092
R9305 GND.n7160 GND.t183 0.00131092
R9306 GND.n7161 GND.n7160 0.00131092
R9307 GND.n3052 GND.n3051 0.00131092
R9308 GND.t583 GND.n3052 0.00131092
R9309 GND.n3060 GND.t583 0.00131092
R9310 GND.n3061 GND.n3060 0.00131092
R9311 GND.n2728 GND.n2727 0.00131092
R9312 GND.t851 GND.n2728 0.00131092
R9313 GND.n2736 GND.t851 0.00131092
R9314 GND.n2737 GND.n2736 0.00131092
R9315 GND.n2403 GND.n2402 0.00131092
R9316 GND.t1196 GND.n2403 0.00131092
R9317 GND.n2411 GND.t1196 0.00131092
R9318 GND.n2412 GND.n2411 0.00131092
R9319 GND.n6919 GND.n6918 0.00131092
R9320 GND.t654 GND.n6919 0.00131092
R9321 GND.n6927 GND.t654 0.00131092
R9322 GND.n6928 GND.n6927 0.00131092
R9323 GND.n1754 GND.n1753 0.00131092
R9324 GND.t782 GND.n1754 0.00131092
R9325 GND.n1762 GND.t782 0.00131092
R9326 GND.n1763 GND.n1762 0.00131092
R9327 GND.n1563 GND.n1562 0.00131092
R9328 GND.t374 GND.n1563 0.00131092
R9329 GND.n1571 GND.t374 0.00131092
R9330 GND.n1572 GND.n1571 0.00131092
R9331 GND.n1553 GND.n1552 0.00131092
R9332 GND.n1552 GND.t71 0.00131092
R9333 GND.n4051 GND.n4050 0.00125043
R9334 GND.n4120 GND 0.00124153
R9335 GND.n4935 GND.n4933 0.00122464
R9336 GND.n5763 GND 0.00116489
R9337 GND.n4491 GND.n4489 0.00116489
R9338 GND.n6432 GND.n6418 0.00116489
R9339 GND.n7047 GND.n7046 0.00115206
R9340 GND.n7046 GND.n4274 0.00115206
R9341 GND.n4063 GND.n4062 0.00114322
R9342 GND.n6802 GND.n6801 0.00109111
R9343 GND.n5461 GND.n5444 0.00108327
R9344 GND.n6866 GND.n6849 0.00108327
R9345 GND.n6803 GND.n6802 0.00107707
R9346 GND.n7048 GND.n7047 0.00107707
R9347 GND.n4422 GND.n4421 0.00107231
R9348 GND.n6758 GND.n6757 0.00107231
R9349 GND.n7366 GND.n7365 0.00103916
R9350 GND.n2018 GND.n2017 0.00103916
R9351 GND.n516 GND.n515 0.00103916
R9352 GND.n211 GND.n210 0.00103916
R9353 GND.n1510 GND.n1509 0.00103916
R9354 GND.n1462 GND.n1461 0.00103916
R9355 GND.n4219 GND.n4218 0.00103916
R9356 GND.n3413 GND.n3412 0.00103916
R9357 GND.n3256 GND.n3255 0.00103916
R9358 GND.n2959 GND.n2958 0.00103916
R9359 GND.n2634 GND.n2633 0.00103916
R9360 GND.n2310 GND.n2309 0.00103916
R9361 GND.n2148 GND.n2147 0.00103916
R9362 GND.n1280 GND.n1279 0.00103916
R9363 GND.n363 GND.n362 0.00103916
R9364 GND.n7411 GND.n7410 0.00103916
R9365 GND.n4050 GND.n4047 0.00103602
R9366 GND.n7493 GND.n7492 0.00101312
R9367 GND.n2082 GND.n2081 0.00101312
R9368 GND.n570 GND.n569 0.00101312
R9369 GND.n261 GND.n260 0.00101312
R9370 GND.n109 GND.n108 0.00101312
R9371 GND.n1442 GND.n1441 0.00101312
R9372 GND.n4269 GND.n4268 0.00101312
R9373 GND.n3466 GND.n3465 0.00101312
R9374 GND.n3308 GND.n3307 0.00101312
R9375 GND.n3012 GND.n3011 0.00101312
R9376 GND.n2688 GND.n2687 0.00101312
R9377 GND.n2363 GND.n2362 0.00101312
R9378 GND.n2205 GND.n2204 0.00101312
R9379 GND.n1324 GND.n1323 0.00101312
R9380 GND.n414 GND.n413 0.00101312
R9381 GND.n840 GND.n839 0.00101312
R9382 GND.n7492 GND.n7460 0.00100714
R9383 GND.n2081 GND.n2047 0.00100714
R9384 GND.n569 GND.n540 0.00100714
R9385 GND.n260 GND.n235 0.00100714
R9386 GND.n108 GND.n68 0.00100714
R9387 GND.n1441 GND.n1409 0.00100714
R9388 GND.n4268 GND.n4243 0.00100714
R9389 GND.n3465 GND.n3437 0.00100714
R9390 GND.n3307 GND.n3280 0.00100714
R9391 GND.n3011 GND.n2983 0.00100714
R9392 GND.n2687 GND.n2658 0.00100714
R9393 GND.n2362 GND.n2334 0.00100714
R9394 GND.n2204 GND.n2172 0.00100714
R9395 GND.n1323 GND.n1304 0.00100714
R9396 GND.n413 GND.n387 0.00100714
R9397 GND.n839 GND.n812 0.00100714
R9398 GND.n4076 GND.n4075 0.00100417
R9399 GND.n7819 GND.n7818 0.001004
R9400 GND.n891 GND.n890 0.001004
R9401 GND.n784 GND.n783 0.001004
R9402 GND.n465 GND.n464 0.001004
R9403 GND.n1683 GND.n1682 0.001004
R9404 GND.n312 GND.n311 0.001004
R9405 GND.n160 GND.n159 0.001004
R9406 GND.n51 GND.n50 0.001004
R9407 GND.n7307 GND.n7306 0.001004
R9408 GND.n3517 GND.n3516 0.001004
R9409 GND.n3359 GND.n3358 0.001004
R9410 GND.n3202 GND.n3201 0.001004
R9411 GND.n2905 GND.n2904 0.001004
R9412 GND.n2580 GND.n2579 0.001004
R9413 GND.n2256 GND.n2255 0.001004
R9414 GND.n1231 GND.n1230 0.001004
R9415 GND.n4127 GND.n4126 0.00100271
R9416 GND.n6762 GND.n5221 0.00100171
R9417 GND.n5218 GND.n5217 0.00100171
R9418 GND.n4373 GND.n4372 0.00100171
R9419 GND.n6872 GND.n6871 0.00100171
R9420 GND.n6792 GND.n6762 0.00100166
R9421 GND.n5217 GND.n5216 0.00100166
R9422 GND.n4373 GND.n4370 0.00100166
R9423 GND.n6871 GND.n4313 0.00100166
R9424 GND.n4163 GND.n4072 0.00100126
R9425 GND.n6660 GND.n6659 0.00100097
R9426 GND.n4449 GND.n4448 0.00100097
R9427 GND.n5102 GND.n5101 0.00100097
R9428 GND.n6471 GND.n6470 0.00100097
R9429 GND.n4586 GND.n4579 0.00100097
R9430 GND.n4667 GND.n4666 0.00100097
R9431 GND.n4923 GND.n4922 0.00100097
R9432 GND.n1941 GND.n1940 0.00100095
R9433 GND.n1708 GND.n1707 0.00100095
R9434 GND.n6916 GND.n6915 0.00100095
R9435 GND.n2384 GND.n2383 0.00100095
R9436 GND.n2709 GND.n2708 0.00100095
R9437 GND.n3033 GND.n3032 0.00100095
R9438 GND.n7106 GND.n7105 0.00100095
R9439 GND.n4801 GND.n4800 0.00100095
R9440 GND.n5283 GND.n5282 0.00100095
R9441 GND.n5805 GND.n5804 0.00100095
R9442 GND.n5972 GND.n5971 0.00100095
R9443 GND.n6139 GND.n6138 0.00100095
R9444 GND.n6303 GND.n6302 0.00100095
R9445 GND.n591 GND.n590 0.00100095
R9446 GND.n7634 GND.n7633 0.00100095
R9447 GND.n7514 GND.n7513 0.00100095
R9448 GND.n6804 GND.n4425 0.00100086
R9449 GND.n7049 GND.n4273 0.00100086
R9450 GND.n2093 GND.n1359 0.00100018
R9451 GND.n7348 GND.n1077 0.00100018
R9452 GND.n7049 GND.n7048 0.00100017
R9453 GND.n6804 GND.n6803 0.00100017
R9454 GND.n2093 GND.n2092 0.00100006
R9455 GND.n7348 GND.n7347 0.00100006
R9456 GND.n4052 GND.n4046 0.00100003
R9457 GND.n7820 GND.n7819 0.00100001
R9458 GND.n892 GND.n891 0.00100001
R9459 GND.n785 GND.n784 0.00100001
R9460 GND.n466 GND.n465 0.00100001
R9461 GND.n1684 GND.n1683 0.00100001
R9462 GND.n313 GND.n312 0.00100001
R9463 GND.n161 GND.n160 0.00100001
R9464 GND.n52 GND.n51 0.00100001
R9465 GND.n7308 GND.n7307 0.00100001
R9466 GND.n3518 GND.n3517 0.00100001
R9467 GND.n3360 GND.n3359 0.00100001
R9468 GND.n3203 GND.n3202 0.00100001
R9469 GND.n2906 GND.n2905 0.00100001
R9470 GND.n2581 GND.n2580 0.00100001
R9471 GND.n2257 GND.n2256 0.00100001
R9472 GND.n1232 GND.n1231 0.00100001
R9473 GND.n2094 GND.n2093 0.001
R9474 GND.n7348 GND.n1080 0.001
R9475 GND.n7348 GND.n1085 0.001
R9476 GND.n7348 GND.n1090 0.001
R9477 GND.n7348 GND.n1095 0.001
R9478 GND.n7348 GND.n1100 0.001
R9479 GND.n7348 GND.n1105 0.001
R9480 GND.n7348 GND.n1110 0.001
R9481 GND.n7348 GND.n1118 0.001
R9482 GND.n7348 GND.n1126 0.001
R9483 GND.n7348 GND.n1134 0.001
R9484 GND.n7348 GND.n1142 0.001
R9485 GND.n7349 GND.n7348 0.001
R9486 GND.n7348 GND.n1150 0.001
R9487 GND.n5437 GND.n5436 0.001
R9488 GND.n7046 GND.n7045 0.001
R9489 GND.n4339 GND.n4338 0.001
R9490 GND.n4060 GND.n4059 0.000966399
R9491 GND.n4059 GND.n4058 0.000959101
R9492 GND.n4058 GND.n4057 0.000959101
R9493 GND.n7433 GND.n7375 0.000943262
R9494 GND.n1986 GND.n1371 0.000943262
R9495 GND.n333 GND.n328 0.000943262
R9496 GND.n486 GND.n481 0.000943262
R9497 GND.n181 GND.n176 0.000943262
R9498 GND.n1516 GND.n1485 0.000943262
R9499 GND.n1468 GND.n1384 0.000943262
R9500 GND.n4189 GND.n4184 0.000943262
R9501 GND.n3383 GND.n3378 0.000943262
R9502 GND.n3226 GND.n3221 0.000943262
R9503 GND.n2929 GND.n2924 0.000943262
R9504 GND.n2604 GND.n2599 0.000943262
R9505 GND.n2280 GND.n2275 0.000943262
R9506 GND.n2118 GND.n2113 0.000943262
R9507 GND.n1250 GND.n1245 0.000943262
R9508 GND.n7417 GND.n7393 0.000943262
R9509 GND.n5783 GND.n5782 0.000898936
R9510 GND.n5690 GND.n5686 0.000898936
R9511 GND.n3681 GND.n3680 0.000864406
R9512 GND.n3687 GND.n3686 0.000864406
R9513 GND.n3682 GND.n3681 0.000858717
R9514 GND.n3684 GND.n3682 0.000858717
R9515 GND.n3686 GND.n3685 0.000858717
R9516 GND.n3685 GND.n3684 0.000858717
R9517 GND.n3625 GND.n3624 0.000858717
R9518 GND.n3624 GND.n3623 0.000858717
R9519 GND.n3622 GND.n3621 0.000858717
R9520 GND.n3623 GND.n3622 0.000858717
R9521 GND.n4078 GND.n4077 0.000840211
R9522 GND.n4163 GND.n4078 0.000840211
R9523 GND.n2089 GND.n2088 0.000826763
R9524 GND.n2096 GND.n2095 0.000826763
R9525 GND.n7344 GND.n7343 0.000826763
R9526 GND.n2262 GND.n2261 0.000826763
R9527 GND.n2586 GND.n2585 0.000826763
R9528 GND.n2911 GND.n2910 0.000826763
R9529 GND.n3208 GND.n3207 0.000826763
R9530 GND.n3365 GND.n3364 0.000826763
R9531 GND.n4171 GND.n4170 0.000826763
R9532 GND.n7313 GND.n7312 0.000826763
R9533 GND.n1115 GND.n1114 0.000826763
R9534 GND.n1123 GND.n1122 0.000826763
R9535 GND.n1131 GND.n1130 0.000826763
R9536 GND.n1139 GND.n1138 0.000826763
R9537 GND.n7351 GND.n7350 0.000826763
R9538 GND.n1147 GND.n1146 0.000826763
R9539 GND.n2083 GND 0.000803226
R9540 GND GND.n2101 0.000803226
R9541 GND.n7338 GND 0.000803226
R9542 GND.n7335 GND 0.000803226
R9543 GND.n7332 GND 0.000803226
R9544 GND.n7329 GND 0.000803226
R9545 GND.n7326 GND 0.000803226
R9546 GND.n7323 GND 0.000803226
R9547 GND.n7319 GND 0.000803226
R9548 GND GND.n0 0.000803226
R9549 GND.n7839 GND 0.000803226
R9550 GND.n7836 GND 0.000803226
R9551 GND.n7833 GND 0.000803226
R9552 GND.n7830 GND 0.000803226
R9553 GND.n7827 GND 0.000803226
R9554 GND.n7824 GND 0.000803226
R9555 GND.n4128 GND.n4127 0.000801918
R9556 GND.n4129 GND.n4128 0.000801918
R9557 GND.n4162 GND.n4161 0.000801918
R9558 GND.n4163 GND.n4162 0.000801918
R9559 GND.n4157 GND.n4156 0.000801918
R9560 GND.n4163 GND.n4157 0.000801918
R9561 GND.n4149 GND.n4148 0.000801918
R9562 GND.n4163 GND.n4149 0.000801918
R9563 GND.n4145 GND.n4144 0.000801918
R9564 GND.n4163 GND.n4145 0.000801918
R9565 GND.n4131 GND.n4130 0.000801918
R9566 GND.n4130 GND.n4129 0.000801918
R9567 GND.n4137 GND.n4136 0.000801918
R9568 GND.n4163 GND.n4137 0.000801918
R9569 GND.n4165 GND.n4164 0.000801918
R9570 GND.n4164 GND.n4163 0.000801918
R9571 GND.n4122 GND.n4121 0.000801918
R9572 GND.n4163 GND.n4122 0.000801918
R9573 GND.n4116 GND.n4112 0.000801918
R9574 GND.n4163 GND.n4112 0.000801918
R9575 GND.n4110 GND.n4109 0.000801918
R9576 GND.n4163 GND.n4110 0.000801918
R9577 GND.n4101 GND.n4100 0.000801918
R9578 GND.n4163 GND.n4101 0.000801918
R9579 GND.n4097 GND.n4096 0.000801918
R9580 GND.n4163 GND.n4097 0.000801918
R9581 GND.n4092 GND.n4091 0.000801918
R9582 GND.n4163 GND.n4092 0.000801918
R9583 GND.n4086 GND.n4085 0.000801918
R9584 GND.n3526 GND.n3525 0.000801918
R9585 GND.n4163 GND.n3526 0.000801918
R9586 GND.n7441 GND.n7440 0.000756235
R9587 GND.n7440 GND.n7439 0.000756235
R9588 GND.n521 GND.n520 0.000756235
R9589 GND.n520 GND.n519 0.000756235
R9590 GND.n216 GND.n215 0.000756235
R9591 GND.n215 GND.n214 0.000756235
R9592 GND.n1390 GND.n1389 0.000756235
R9593 GND.n1389 GND.n1388 0.000756235
R9594 GND.n4224 GND.n4223 0.000756235
R9595 GND.n4223 GND.n4222 0.000756235
R9596 GND.n3418 GND.n3417 0.000756235
R9597 GND.n3417 GND.n3416 0.000756235
R9598 GND.n3261 GND.n3260 0.000756235
R9599 GND.n3260 GND.n3259 0.000756235
R9600 GND.n2964 GND.n2963 0.000756235
R9601 GND.n2963 GND.n2962 0.000756235
R9602 GND.n2639 GND.n2638 0.000756235
R9603 GND.n2638 GND.n2637 0.000756235
R9604 GND.n2315 GND.n2314 0.000756235
R9605 GND.n2314 GND.n2313 0.000756235
R9606 GND.n2153 GND.n2152 0.000756235
R9607 GND.n2152 GND.n2151 0.000756235
R9608 GND.n1285 GND.n1284 0.000756235
R9609 GND.n1284 GND.n1283 0.000756235
R9610 GND.n89 GND.n88 0.000756235
R9611 GND.n92 GND.n89 0.000756235
R9612 GND.n368 GND.n367 0.000756235
R9613 GND.n367 GND.n366 0.000756235
R9614 GND.n2023 GND.n2022 0.000756235
R9615 GND.n2022 GND.n2021 0.000756235
R9616 GND.n793 GND.n792 0.000756235
R9617 GND.n792 GND.n791 0.000756235
R9618 GND.n4060 GND.n4054 0.000714408
R9619 GND.n2084 GND.n2083 0.000666774
R9620 GND.n2101 GND.n2100 0.000666774
R9621 GND.n7339 GND.n7338 0.000666774
R9622 GND.n7336 GND.n7335 0.000666774
R9623 GND.n7333 GND.n7332 0.000666774
R9624 GND.n7330 GND.n7329 0.000666774
R9625 GND.n7327 GND.n7326 0.000666774
R9626 GND.n7324 GND.n7323 0.000666774
R9627 GND.n7320 GND.n7319 0.000666774
R9628 GND.n7317 GND.n0 0.000666774
R9629 GND.n7840 GND.n7839 0.000666774
R9630 GND.n7837 GND.n7836 0.000666774
R9631 GND.n7834 GND.n7833 0.000666774
R9632 GND.n7831 GND.n7830 0.000666774
R9633 GND.n7828 GND.n7827 0.000666774
R9634 GND.n7825 GND.n7824 0.000666774
R9635 GND.n5521 GND.n5519 0.000632979
R9636 GND.n5042 GND.n4576 0.000632979
R9637 GND.n6600 GND.n5496 0.000632979
R9638 GND.n4054 GND.n4052 0.000607204
R9639 GND.n4040 GND.n4039 0.000567786
R9640 GND.n4370 GND.n4340 0.000560793
R9641 GND.n5216 GND.n5178 0.000560793
R9642 GND.n6793 GND.n6792 0.000560793
R9643 GND.n6873 GND.n6872 0.000557763
R9644 GND.n4372 GND.n4371 0.000557763
R9645 GND.n5219 GND.n5218 0.000557763
R9646 GND.n5919 GND.n5221 0.000557763
R9647 GND.n3666 GND.n3665 0.000557678
R9648 GND.n1903 GND.n1902 0.000544755
R9649 GND.n1860 GND.n1859 0.000544755
R9650 GND.n7036 GND.n7035 0.000544755
R9651 GND.n2509 GND.n2508 0.000544755
R9652 GND.n2834 GND.n2833 0.000544755
R9653 GND.n3131 GND.n3130 0.000544755
R9654 GND.n7231 GND.n7230 0.000544755
R9655 GND.n4763 GND.n4762 0.000544755
R9656 GND.n5428 GND.n5427 0.000544755
R9657 GND.n5931 GND.n5930 0.000544755
R9658 GND.n6100 GND.n6099 0.000544755
R9659 GND.n6264 GND.n6263 0.000544755
R9660 GND.n6573 GND.n6572 0.000544755
R9661 GND.n713 GND.n712 0.000544755
R9662 GND.n7760 GND.n7759 0.000544755
R9663 GND.n7595 GND.n7594 0.000544755
R9664 GND.n3672 GND.n3671 0.000538452
R9665 GND.n3628 GND.n3627 0.000537082
R9666 GND.n7551 GND.n7550 0.000530553
R9667 GND.n7682 GND.n7681 0.000530553
R9668 GND.n635 GND.n634 0.000530553
R9669 GND.n6347 GND.n6346 0.000530553
R9670 GND.n6183 GND.n6182 0.000530553
R9671 GND.n6019 GND.n6018 0.000530553
R9672 GND.n5836 GND.n5835 0.000530553
R9673 GND.n5314 GND.n5313 0.000530553
R9674 GND.n4873 GND.n4872 0.000530553
R9675 GND.n7180 GND.n7179 0.000530553
R9676 GND.n3080 GND.n3079 0.000530553
R9677 GND.n2756 GND.n2755 0.000530553
R9678 GND.n2431 GND.n2430 0.000530553
R9679 GND.n6947 GND.n6946 0.000530553
R9680 GND.n1782 GND.n1781 0.000530553
R9681 GND.n1591 GND.n1590 0.000530553
R9682 GND.n6846 GND.n6845 0.000528881
R9683 GND.n6845 GND.n6844 0.000528881
R9684 GND.n6848 GND.n6847 0.000528881
R9685 GND.n5441 GND.n5440 0.000528881
R9686 GND.n5440 GND.n5439 0.000528881
R9687 GND.n5443 GND.n5442 0.000528881
R9688 GND.n7572 GND.n7571 0.00052846
R9689 GND.n7708 GND.n7707 0.00052846
R9690 GND.n661 GND.n660 0.00052846
R9691 GND.n6373 GND.n6372 0.00052846
R9692 GND.n6209 GND.n6208 0.00052846
R9693 GND.n6045 GND.n6044 0.00052846
R9694 GND.n5862 GND.n5861 0.00052846
R9695 GND.n5340 GND.n5339 0.00052846
R9696 GND.n4899 GND.n4898 0.00052846
R9697 GND.n7206 GND.n7205 0.00052846
R9698 GND.n3106 GND.n3105 0.00052846
R9699 GND.n2782 GND.n2781 0.00052846
R9700 GND.n2457 GND.n2456 0.00052846
R9701 GND.n6973 GND.n6972 0.00052846
R9702 GND.n1808 GND.n1807 0.00052846
R9703 GND.n1617 GND.n1616 0.00052846
R9704 GND.n1969 GND.n1968 0.00052846
R9705 GND.n1731 GND.n1730 0.00052846
R9706 GND.n1827 GND.n1826 0.00052846
R9707 GND.n6992 GND.n6991 0.00052846
R9708 GND.n2476 GND.n2475 0.00052846
R9709 GND.n2801 GND.n2800 0.00052846
R9710 GND.n7129 GND.n7128 0.00052846
R9711 GND.n4822 GND.n4821 0.00052846
R9712 GND.n5398 GND.n5397 0.00052846
R9713 GND.n5359 GND.n5358 0.00052846
R9714 GND.n5881 GND.n5880 0.00052846
R9715 GND.n6067 GND.n6066 0.00052846
R9716 GND.n6231 GND.n6230 0.00052846
R9717 GND.n6395 GND.n6394 0.00052846
R9718 GND.n680 GND.n679 0.00052846
R9719 GND.n7727 GND.n7726 0.00052846
R9720 GND.n3691 GND.n3690 0.000526656
R9721 GND.n7735 GND.n7734 0.0005264
R9722 GND.n688 GND.n687 0.0005264
R9723 GND.n6403 GND.n6402 0.0005264
R9724 GND.n6239 GND.n6238 0.0005264
R9725 GND.n6075 GND.n6074 0.0005264
R9726 GND.n5889 GND.n5888 0.0005264
R9727 GND.n5367 GND.n5366 0.0005264
R9728 GND.n5406 GND.n5405 0.0005264
R9729 GND.n4830 GND.n4829 0.0005264
R9730 GND.n7137 GND.n7136 0.0005264
R9731 GND.n2809 GND.n2808 0.0005264
R9732 GND.n2484 GND.n2483 0.0005264
R9733 GND.n7000 GND.n6999 0.0005264
R9734 GND.n1835 GND.n1834 0.0005264
R9735 GND.n1739 GND.n1738 0.0005264
R9736 GND.n1977 GND.n1976 0.0005264
R9737 GND.n4042 GND.n4041 0.000525991
R9738 GND.n3630 GND.n3629 0.000524722
R9739 GND.n3535 GND.n3534 0.000523819
R9740 GND.n4065 GND.n4063 0.000523819
R9741 GND.n3530 GND.n3529 0.000523819
R9742 GND.t392 GND.n3536 0.000523446
R9743 GND.n4066 GND.n4065 0.000523446
R9744 GND.t392 GND.n4066 0.000523446
R9745 GND.n3536 GND.n3535 0.000523446
R9746 GND.n3531 GND.n3530 0.000523446
R9747 GND.t392 GND.n3531 0.000523446
R9748 GND.n3644 GND.n3643 0.000517138
R9749 GND.n7717 GND.n7716 0.000512627
R9750 GND.n670 GND.n669 0.000512627
R9751 GND.n6385 GND.n6384 0.000512627
R9752 GND.n6221 GND.n6220 0.000512627
R9753 GND.n6057 GND.n6056 0.000512627
R9754 GND.n5871 GND.n5870 0.000512627
R9755 GND.n5349 GND.n5348 0.000512627
R9756 GND.n5388 GND.n5387 0.000512627
R9757 GND.n4812 GND.n4811 0.000512627
R9758 GND.n7119 GND.n7118 0.000512627
R9759 GND.n2791 GND.n2790 0.000512627
R9760 GND.n2466 GND.n2465 0.000512627
R9761 GND.n6982 GND.n6981 0.000512627
R9762 GND.n1817 GND.n1816 0.000512627
R9763 GND.n1721 GND.n1720 0.000512627
R9764 GND.n1959 GND.n1958 0.000512627
R9765 GND.n7545 GND.n7544 0.000512369
R9766 GND.n7676 GND.n7675 0.000512369
R9767 GND.n629 GND.n628 0.000512369
R9768 GND.n6341 GND.n6340 0.000512369
R9769 GND.n6177 GND.n6176 0.000512369
R9770 GND.n6013 GND.n6012 0.000512369
R9771 GND.n5830 GND.n5829 0.000512369
R9772 GND.n5308 GND.n5307 0.000512369
R9773 GND.n4867 GND.n4866 0.000512369
R9774 GND.n7174 GND.n7173 0.000512369
R9775 GND.n3074 GND.n3073 0.000512369
R9776 GND.n2750 GND.n2749 0.000512369
R9777 GND.n2425 GND.n2424 0.000512369
R9778 GND.n6941 GND.n6940 0.000512369
R9779 GND.n1776 GND.n1775 0.000512369
R9780 GND.n1585 GND.n1584 0.000512369
R9781 GND.n4091 GND.n4090 0.000508571
R9782 GND.n4096 GND.n4095 0.000508571
R9783 GND.n4100 GND.n4099 0.000508571
R9784 GND.n4109 GND.n4108 0.000508571
R9785 GND.n4117 GND.n4116 0.000508571
R9786 GND.n4121 GND.n4120 0.000508571
R9787 GND.n4166 GND.n4165 0.000508571
R9788 GND.n4136 GND.n4135 0.000508571
R9789 GND.n4144 GND.n4143 0.000508571
R9790 GND.n4148 GND.n4147 0.000508571
R9791 GND.n4156 GND.n4155 0.000508571
R9792 GND.n4161 GND.n4160 0.000508571
R9793 GND.n3525 GND.n3524 0.000508571
R9794 GND.n7652 GND.n7651 0.000507826
R9795 GND.n609 GND.n608 0.000507826
R9796 GND.n6321 GND.n6320 0.000507826
R9797 GND.n6157 GND.n6156 0.000507826
R9798 GND.n5990 GND.n5989 0.000507826
R9799 GND.n5807 GND.n5806 0.000507826
R9800 GND.n5285 GND.n5284 0.000507826
R9801 GND.n4844 GND.n4843 0.000507826
R9802 GND.n7151 GND.n7150 0.000507826
R9803 GND.n3051 GND.n3050 0.000507826
R9804 GND.n2727 GND.n2726 0.000507826
R9805 GND.n2402 GND.n2401 0.000507826
R9806 GND.n6918 GND.n6917 0.000507826
R9807 GND.n1753 GND.n1752 0.000507826
R9808 GND.n1562 GND.n1561 0.000507826
R9809 GND.n1554 GND.n1553 0.000507826
R9810 GND.n7533 GND.n7532 0.000507826
R9811 GND.n7664 GND.n7663 0.000507826
R9812 GND.n620 GND.n619 0.000507826
R9813 GND.n6332 GND.n6331 0.000507826
R9814 GND.n6168 GND.n6167 0.000507826
R9815 GND.n6001 GND.n6000 0.000507826
R9816 GND.n5818 GND.n5817 0.000507826
R9817 GND.n5296 GND.n5295 0.000507826
R9818 GND.n4855 GND.n4854 0.000507826
R9819 GND.n7162 GND.n7161 0.000507826
R9820 GND.n3062 GND.n3061 0.000507826
R9821 GND.n2738 GND.n2737 0.000507826
R9822 GND.n2413 GND.n2412 0.000507826
R9823 GND.n6929 GND.n6928 0.000507826
R9824 GND.n1764 GND.n1763 0.000507826
R9825 GND.n1573 GND.n1572 0.000507826
R9826 GND.n2080 GND.n2079 0.000507291
R9827 GND.n412 GND.n411 0.000507291
R9828 GND.n838 GND.n837 0.000507291
R9829 GND.n4448 GND.n4447 0.000506774
R9830 GND.n4542 GND.n4541 0.000506774
R9831 GND.n5101 GND.n5100 0.000506774
R9832 GND.n5176 GND.n5175 0.000506774
R9833 GND.n5099 GND.n5098 0.000506774
R9834 GND.n4544 GND.n4543 0.000506774
R9835 GND.n5564 GND.n5563 0.000506774
R9836 GND.n5566 GND.n5565 0.000506774
R9837 GND.n5766 GND.n5648 0.000506774
R9838 GND.n5765 GND.n5764 0.000506774
R9839 GND.n5768 GND.n5767 0.000506774
R9840 GND.n5647 GND.n5646 0.000506774
R9841 GND.n4666 GND.n4665 0.000506774
R9842 GND.n4922 GND.n4921 0.000506774
R9843 GND.n4579 GND.n4578 0.000506774
R9844 GND.n4664 GND.n4663 0.000506774
R9845 GND.n4749 GND.n4748 0.000506774
R9846 GND.n4979 GND.n4978 0.000506774
R9847 GND.n5016 GND.n5015 0.000506774
R9848 GND.n6474 GND.n6473 0.000506774
R9849 GND.n6659 GND.n6658 0.000506774
R9850 GND.n6734 GND.n6733 0.000506774
R9851 GND.n6657 GND.n6656 0.000506774
R9852 GND.n6559 GND.n6558 0.000506774
R9853 GND.n6472 GND.n6471 0.000506774
R9854 GND.n1984 GND.n1983 0.000505544
R9855 GND.n494 GND.n493 0.000505544
R9856 GND.n189 GND.n188 0.000505544
R9857 GND.n1524 GND.n1523 0.000505544
R9858 GND.n1476 GND.n1475 0.000505544
R9859 GND.n4197 GND.n4196 0.000505544
R9860 GND.n3391 GND.n3390 0.000505544
R9861 GND.n3234 GND.n3233 0.000505544
R9862 GND.n2937 GND.n2936 0.000505544
R9863 GND.n2612 GND.n2611 0.000505544
R9864 GND.n2288 GND.n2287 0.000505544
R9865 GND.n2126 GND.n2125 0.000505544
R9866 GND.n1258 GND.n1257 0.000505544
R9867 GND.n341 GND.n340 0.000505544
R9868 GND.n7425 GND.n7424 0.000505544
R9869 GND.n7431 GND.n7430 0.000505544
R9870 GND.n1942 GND.n1941 0.000504863
R9871 GND.n1709 GND.n1708 0.000504863
R9872 GND.n7025 GND.n6916 0.000504863
R9873 GND.n2385 GND.n2384 0.000504863
R9874 GND.n2710 GND.n2709 0.000504863
R9875 GND.n3034 GND.n3033 0.000504863
R9876 GND.n7107 GND.n7106 0.000504863
R9877 GND.n4802 GND.n4801 0.000504863
R9878 GND.n5420 GND.n5283 0.000504863
R9879 GND.n5915 GND.n5805 0.000504863
R9880 GND.n5973 GND.n5972 0.000504863
R9881 GND.n6140 GND.n6139 0.000504863
R9882 GND.n6304 GND.n6303 0.000504863
R9883 GND.n592 GND.n591 0.000504863
R9884 GND.n7635 GND.n7634 0.000504863
R9885 GND.n7515 GND.n7514 0.000504863
R9886 GND.n4105 GND.n4104 0.000504378
R9887 GND.n4087 GND.n4086 0.000504346
R9888 GND.n4132 GND.n4131 0.000504346
R9889 GND.n4159 GND.n4158 0.00050424
R9890 GND.n4152 GND.n4151 0.00050424
R9891 GND.n4134 GND.n4133 0.00050424
R9892 GND.n3523 GND.n3522 0.00050424
R9893 GND.n4119 GND.n4118 0.00050424
R9894 GND.n4107 GND.n4106 0.00050424
R9895 GND.n4081 GND.n4080 0.00050424
R9896 GND.n4083 GND.n4082 0.00050424
R9897 GND.n4140 GND.n4139 0.000504176
R9898 GND.n4154 GND.n4153 0.000504112
R9899 GND.n4142 GND.n4141 0.000504112
R9900 GND.n4168 GND.n4167 0.000504112
R9901 GND.n4094 GND.n4093 0.000504112
R9902 GND.n4089 GND.n4088 0.000504112
R9903 GND.n7821 GND.n7820 0.000504005
R9904 GND.n893 GND.n892 0.000504005
R9905 GND.n786 GND.n785 0.000504005
R9906 GND.n467 GND.n466 0.000504005
R9907 GND.n1685 GND.n1684 0.000504005
R9908 GND.n314 GND.n313 0.000504005
R9909 GND.n162 GND.n161 0.000504005
R9910 GND.n53 GND.n52 0.000504005
R9911 GND.n7309 GND.n7308 0.000504005
R9912 GND.n3519 GND.n3518 0.000504005
R9913 GND.n3361 GND.n3360 0.000504005
R9914 GND.n3204 GND.n3203 0.000504005
R9915 GND.n2907 GND.n2906 0.000504005
R9916 GND.n2582 GND.n2581 0.000504005
R9917 GND.n2258 GND.n2257 0.000504005
R9918 GND.n1233 GND.n1232 0.000504005
R9919 GND.n4054 GND.n4053 0.00050212
R9920 GND.n895 GND.n894 0.000501449
R9921 GND.n788 GND.n787 0.000501449
R9922 GND.n469 GND.n468 0.000501449
R9923 GND.n1687 GND.n1686 0.000501449
R9924 GND.n316 GND.n315 0.000501449
R9925 GND.n164 GND.n163 0.000501449
R9926 GND.n55 GND.n54 0.000501449
R9927 GND.n7311 GND.n7310 0.000501449
R9928 GND.n3521 GND.n3520 0.000501449
R9929 GND.n3363 GND.n3362 0.000501449
R9930 GND.n3206 GND.n3205 0.000501449
R9931 GND.n2909 GND.n2908 0.000501449
R9932 GND.n2584 GND.n2583 0.000501449
R9933 GND.n2260 GND.n2259 0.000501449
R9934 GND.n1235 GND.n1234 0.000501449
R9935 GND.n7823 GND.n7822 0.000501449
R9936 GND.n1918 GND.n1917 0.000501292
R9937 GND.n1917 GND.n1916 0.000501292
R9938 GND.n1875 GND.n1874 0.000501292
R9939 GND.n1874 GND.n1873 0.000501292
R9940 GND.n7032 GND.n7031 0.000501292
R9941 GND.n7033 GND.n7032 0.000501292
R9942 GND.n2524 GND.n2523 0.000501292
R9943 GND.n2523 GND.n2522 0.000501292
R9944 GND.n2849 GND.n2848 0.000501292
R9945 GND.n2848 GND.n2847 0.000501292
R9946 GND.n3146 GND.n3145 0.000501292
R9947 GND.n3145 GND.n3144 0.000501292
R9948 GND.n7246 GND.n7245 0.000501292
R9949 GND.n7245 GND.n7244 0.000501292
R9950 GND.n4778 GND.n4777 0.000501292
R9951 GND.n4777 GND.n4776 0.000501292
R9952 GND.n5424 GND.n5423 0.000501292
R9953 GND.n5425 GND.n5424 0.000501292
R9954 GND.n5946 GND.n5945 0.000501292
R9955 GND.n5945 GND.n5944 0.000501292
R9956 GND.n6115 GND.n6114 0.000501292
R9957 GND.n6114 GND.n6113 0.000501292
R9958 GND.n6279 GND.n6278 0.000501292
R9959 GND.n6278 GND.n6277 0.000501292
R9960 GND.n6588 GND.n6587 0.000501292
R9961 GND.n6587 GND.n6586 0.000501292
R9962 GND.n728 GND.n727 0.000501292
R9963 GND.n727 GND.n726 0.000501292
R9964 GND.n7775 GND.n7774 0.000501292
R9965 GND.n7774 GND.n7773 0.000501292
R9966 GND.n7610 GND.n7609 0.000501292
R9967 GND.n7609 GND.n7608 0.000501292
R9968 GND.n3626 GND.n3625 0.00050117
R9969 GND.n3621 GND.n3620 0.00050117
R9970 GND.n4541 GND.n4540 0.00050097
R9971 GND.n5175 GND.n5174 0.00050097
R9972 GND.n5098 GND.n5097 0.00050097
R9973 GND.n4545 GND.n4544 0.00050097
R9974 GND.n5563 GND.n5562 0.00050097
R9975 GND.n5567 GND.n5566 0.00050097
R9976 GND.n5691 GND.n5648 0.00050097
R9977 GND.n5764 GND.n5763 0.00050097
R9978 GND.n5769 GND.n5768 0.00050097
R9979 GND.n5646 GND.n5645 0.00050097
R9980 GND.n4748 GND.n4747 0.00050097
R9981 GND.n4980 GND.n4979 0.00050097
R9982 GND.n5017 GND.n5016 0.00050097
R9983 GND.n6475 GND.n6474 0.00050097
R9984 GND.n6733 GND.n6732 0.00050097
R9985 GND.n6656 GND.n6655 0.00050097
R9986 GND.n6558 GND.n6557 0.00050097
R9987 GND.n4663 GND.n4662 0.00050097
R9988 GND.n1985 GND.n1984 0.000500915
R9989 GND.n493 GND.n492 0.000500915
R9990 GND.n188 GND.n187 0.000500915
R9991 GND.n1523 GND.n1522 0.000500915
R9992 GND.n1475 GND.n1474 0.000500915
R9993 GND.n4196 GND.n4195 0.000500915
R9994 GND.n3390 GND.n3389 0.000500915
R9995 GND.n3233 GND.n3232 0.000500915
R9996 GND.n2936 GND.n2935 0.000500915
R9997 GND.n2611 GND.n2610 0.000500915
R9998 GND.n2287 GND.n2286 0.000500915
R9999 GND.n2125 GND.n2124 0.000500915
R10000 GND.n1257 GND.n1256 0.000500915
R10001 GND.n340 GND.n339 0.000500915
R10002 GND.n7424 GND.n7423 0.000500915
R10003 GND.n7432 GND.n7431 0.000500915
R10004 GND.n3674 GND.n3673 0.000500552
R10005 GND.n3689 GND.n3688 0.000500539
R10006 GND.n7352 GND.n7351 0.000500526
R10007 GND.n2088 GND.n2087 0.000500526
R10008 GND.n1138 GND.n1137 0.000500526
R10009 GND.n1122 GND.n1121 0.000500526
R10010 GND.n1114 GND.n1113 0.000500526
R10011 GND.n7314 GND.n7313 0.000500526
R10012 GND.n4172 GND.n4171 0.000500526
R10013 GND.n3366 GND.n3365 0.000500526
R10014 GND.n3209 GND.n3208 0.000500526
R10015 GND.n2912 GND.n2911 0.000500526
R10016 GND.n2587 GND.n2586 0.000500526
R10017 GND.n2263 GND.n2262 0.000500526
R10018 GND.n7343 GND.n7342 0.000500526
R10019 GND.n2097 GND.n2096 0.000500526
R10020 GND.n1130 GND.n1129 0.000500526
R10021 GND.n1146 GND.n1145 0.000500526
R10022 GND.n3619 GND.n3618 0.000500355
R10023 GND.n3538 GND.n3537 0.000500347
R10024 GND.n7435 GND.n7433 0.000500286
R10025 GND.n1988 GND.n1986 0.000500286
R10026 GND.n333 GND.n332 0.000500286
R10027 GND.n486 GND.n485 0.000500286
R10028 GND.n181 GND.n180 0.000500286
R10029 GND.n1516 GND.n1515 0.000500286
R10030 GND.n1468 GND.n1467 0.000500286
R10031 GND.n4189 GND.n4188 0.000500286
R10032 GND.n3383 GND.n3382 0.000500286
R10033 GND.n3226 GND.n3225 0.000500286
R10034 GND.n2929 GND.n2928 0.000500286
R10035 GND.n2604 GND.n2603 0.000500286
R10036 GND.n2280 GND.n2279 0.000500286
R10037 GND.n2118 GND.n2117 0.000500286
R10038 GND.n1250 GND.n1249 0.000500286
R10039 GND.n7417 GND.n7416 0.000500286
R10040 GND.n3875 GND.n3874 0.000500199
R10041 GND.n5039 GND.n5038 0.00050016
R10042 GND.n3883 GND.n3882 0.000500107
R10043 GND.n2086 GND.n2084 0.000500059
R10044 GND.n2100 GND.n2099 0.000500059
R10045 GND.n7341 GND.n7339 0.000500059
R10046 GND.n7336 GND.n2265 0.000500059
R10047 GND.n7333 GND.n2589 0.000500059
R10048 GND.n7330 GND.n2914 0.000500059
R10049 GND.n7327 GND.n3211 0.000500059
R10050 GND.n7840 GND.n57 0.000500059
R10051 GND.n7317 GND.n7316 0.000500059
R10052 GND.n7324 GND.n3368 0.000500059
R10053 GND.n7320 GND.n4174 0.000500059
R10054 GND.n7837 GND.n166 0.000500059
R10055 GND.n7834 GND.n318 0.000500059
R10056 GND.n7831 GND.n471 0.000500059
R10057 GND.n7828 GND.n790 0.000500059
R10058 GND.n7825 GND.n7354 0.000500059
R10059 GND.n3533 GND.n3532 0.000500053
R10060 GND.n3528 GND.n3527 0.000500023
R10061 GND.n4115 GND.n4114 0.00050002
R10062 VDD.n1970 VDD.n1931 8089.41
R10063 VDD.n1951 VDD.n1949 8089.41
R10064 VDD.n1954 VDD.n1948 6801.18
R10065 VDD.n1913 VDD.n1895 2565.88
R10066 VDD.n1913 VDD.n1896 2565.88
R10067 VDD.n1878 VDD.n1823 2565.88
R10068 VDD.n1859 VDD.n1848 2565.88
R10069 VDD.n1864 VDD.n1848 2565.88
R10070 VDD.n2180 VDD.n2169 2565.88
R10071 VDD.n2185 VDD.n2169 2565.88
R10072 VDD.n2199 VDD.n2144 2565.88
R10073 VDD.n2234 VDD.n2216 2565.88
R10074 VDD.n2234 VDD.n2217 2565.88
R10075 VDD.n2438 VDD.n2427 2565.88
R10076 VDD.n2443 VDD.n2427 2565.88
R10077 VDD.n2457 VDD.n2402 2565.88
R10078 VDD.n2492 VDD.n2474 2565.88
R10079 VDD.n2492 VDD.n2475 2565.88
R10080 VDD.n2696 VDD.n2685 2565.88
R10081 VDD.n2701 VDD.n2685 2565.88
R10082 VDD.n2715 VDD.n2660 2565.88
R10083 VDD.n2750 VDD.n2732 2565.88
R10084 VDD.n2750 VDD.n2733 2565.88
R10085 VDD.n2954 VDD.n2943 2565.88
R10086 VDD.n2959 VDD.n2943 2565.88
R10087 VDD.n2973 VDD.n2918 2565.88
R10088 VDD.n3008 VDD.n2990 2565.88
R10089 VDD.n3008 VDD.n2991 2565.88
R10090 VDD.n3212 VDD.n3201 2565.88
R10091 VDD.n3217 VDD.n3201 2565.88
R10092 VDD.n3231 VDD.n3176 2565.88
R10093 VDD.n3266 VDD.n3248 2565.88
R10094 VDD.n3266 VDD.n3249 2565.88
R10095 VDD.n3470 VDD.n3459 2565.88
R10096 VDD.n3475 VDD.n3459 2565.88
R10097 VDD.n3489 VDD.n3434 2565.88
R10098 VDD.n3524 VDD.n3506 2565.88
R10099 VDD.n3524 VDD.n3507 2565.88
R10100 VDD.n5797 VDD.n5786 2565.88
R10101 VDD.n5802 VDD.n5786 2565.88
R10102 VDD.n5816 VDD.n5761 2565.88
R10103 VDD.n5851 VDD.n5833 2565.88
R10104 VDD.n5851 VDD.n5834 2565.88
R10105 VDD.n5543 VDD.n5532 2565.88
R10106 VDD.n5548 VDD.n5532 2565.88
R10107 VDD.n5562 VDD.n5507 2565.88
R10108 VDD.n5597 VDD.n5579 2565.88
R10109 VDD.n5597 VDD.n5580 2565.88
R10110 VDD.n3728 VDD.n3717 2565.88
R10111 VDD.n3733 VDD.n3717 2565.88
R10112 VDD.n3747 VDD.n3692 2565.88
R10113 VDD.n3782 VDD.n3764 2565.88
R10114 VDD.n3782 VDD.n3765 2565.88
R10115 VDD.n3986 VDD.n3975 2565.88
R10116 VDD.n3991 VDD.n3975 2565.88
R10117 VDD.n4005 VDD.n3950 2565.88
R10118 VDD.n4040 VDD.n4022 2565.88
R10119 VDD.n4040 VDD.n4023 2565.88
R10120 VDD.n4244 VDD.n4233 2565.88
R10121 VDD.n4249 VDD.n4233 2565.88
R10122 VDD.n4263 VDD.n4208 2565.88
R10123 VDD.n4298 VDD.n4280 2565.88
R10124 VDD.n4298 VDD.n4281 2565.88
R10125 VDD.n4502 VDD.n4491 2565.88
R10126 VDD.n4507 VDD.n4491 2565.88
R10127 VDD.n4521 VDD.n4466 2565.88
R10128 VDD.n4556 VDD.n4538 2565.88
R10129 VDD.n4556 VDD.n4539 2565.88
R10130 VDD.n4760 VDD.n4749 2565.88
R10131 VDD.n4765 VDD.n4749 2565.88
R10132 VDD.n4779 VDD.n4724 2565.88
R10133 VDD.n4814 VDD.n4796 2565.88
R10134 VDD.n4814 VDD.n4797 2565.88
R10135 VDD.n5075 VDD.n5057 2565.88
R10136 VDD.n5075 VDD.n5058 2565.88
R10137 VDD.n5040 VDD.n4985 2565.88
R10138 VDD.n5021 VDD.n5010 2565.88
R10139 VDD.n5026 VDD.n5010 2565.88
R10140 VDD.n5337 VDD.n5319 2565.88
R10141 VDD.n5337 VDD.n5320 2565.88
R10142 VDD.n5302 VDD.n5247 2565.88
R10143 VDD.n5283 VDD.n5272 2565.88
R10144 VDD.n5288 VDD.n5272 2565.88
R10145 VDD.n1744 VDD.n1713 2082.55
R10146 VDD.n2093 VDD.n2062 2082.55
R10147 VDD.n2323 VDD.n2292 2082.55
R10148 VDD.n2581 VDD.n2550 2082.55
R10149 VDD.n2839 VDD.n2808 2082.55
R10150 VDD.n3097 VDD.n3066 2082.55
R10151 VDD.n3355 VDD.n3324 2082.55
R10152 VDD.n5685 VDD.n5654 2082.55
R10153 VDD.n5431 VDD.n5400 2082.55
R10154 VDD.n3613 VDD.n3582 2082.55
R10155 VDD.n3871 VDD.n3840 2082.55
R10156 VDD.n4129 VDD.n4098 2082.55
R10157 VDD.n4387 VDD.n4356 2082.55
R10158 VDD.n4645 VDD.n4614 2082.55
R10159 VDD.n4903 VDD.n4872 2082.55
R10160 VDD.n5195 VDD.n5164 2082.55
R10161 VDD.n1694 VDD.n1674 2080.64
R10162 VDD.n2043 VDD.n2023 2080.64
R10163 VDD.n2273 VDD.n2253 2080.64
R10164 VDD.n2531 VDD.n2511 2080.64
R10165 VDD.n2789 VDD.n2769 2080.64
R10166 VDD.n3047 VDD.n3027 2080.64
R10167 VDD.n3305 VDD.n3285 2080.64
R10168 VDD.n5635 VDD.n5615 2080.64
R10169 VDD.n5381 VDD.n5361 2080.64
R10170 VDD.n3563 VDD.n3543 2080.64
R10171 VDD.n3821 VDD.n3801 2080.64
R10172 VDD.n4079 VDD.n4059 2080.64
R10173 VDD.n4337 VDD.n4317 2080.64
R10174 VDD.n4595 VDD.n4575 2080.64
R10175 VDD.n4853 VDD.n4833 2080.64
R10176 VDD.n5145 VDD.n5125 2080.64
R10177 VDD.n1742 VDD.n1712 2015.29
R10178 VDD.n1698 VDD.n1678 2015.29
R10179 VDD.n2091 VDD.n2061 2015.29
R10180 VDD.n2047 VDD.n2027 2015.29
R10181 VDD.n2321 VDD.n2291 2015.29
R10182 VDD.n2277 VDD.n2257 2015.29
R10183 VDD.n2579 VDD.n2549 2015.29
R10184 VDD.n2535 VDD.n2515 2015.29
R10185 VDD.n2837 VDD.n2807 2015.29
R10186 VDD.n2793 VDD.n2773 2015.29
R10187 VDD.n3095 VDD.n3065 2015.29
R10188 VDD.n3051 VDD.n3031 2015.29
R10189 VDD.n3353 VDD.n3323 2015.29
R10190 VDD.n3309 VDD.n3289 2015.29
R10191 VDD.n5683 VDD.n5653 2015.29
R10192 VDD.n5639 VDD.n5619 2015.29
R10193 VDD.n5429 VDD.n5399 2015.29
R10194 VDD.n5385 VDD.n5365 2015.29
R10195 VDD.n3611 VDD.n3581 2015.29
R10196 VDD.n3567 VDD.n3547 2015.29
R10197 VDD.n3869 VDD.n3839 2015.29
R10198 VDD.n3825 VDD.n3805 2015.29
R10199 VDD.n4127 VDD.n4097 2015.29
R10200 VDD.n4083 VDD.n4063 2015.29
R10201 VDD.n4385 VDD.n4355 2015.29
R10202 VDD.n4341 VDD.n4321 2015.29
R10203 VDD.n4643 VDD.n4613 2015.29
R10204 VDD.n4599 VDD.n4579 2015.29
R10205 VDD.n4901 VDD.n4871 2015.29
R10206 VDD.n4857 VDD.n4837 2015.29
R10207 VDD.n5193 VDD.n5163 2015.29
R10208 VDD.n5149 VDD.n5129 2015.29
R10209 VDD.n1904 VDD.n1894 1997.65
R10210 VDD.n1899 VDD.n1894 1997.65
R10211 VDD.n1868 VDD.n1850 1997.65
R10212 VDD.n1868 VDD.n1851 1997.65
R10213 VDD.n2189 VDD.n2171 1997.65
R10214 VDD.n2189 VDD.n2172 1997.65
R10215 VDD.n2225 VDD.n2215 1997.65
R10216 VDD.n2220 VDD.n2215 1997.65
R10217 VDD.n2447 VDD.n2429 1997.65
R10218 VDD.n2447 VDD.n2430 1997.65
R10219 VDD.n2483 VDD.n2473 1997.65
R10220 VDD.n2478 VDD.n2473 1997.65
R10221 VDD.n2705 VDD.n2687 1997.65
R10222 VDD.n2705 VDD.n2688 1997.65
R10223 VDD.n2741 VDD.n2731 1997.65
R10224 VDD.n2736 VDD.n2731 1997.65
R10225 VDD.n2963 VDD.n2945 1997.65
R10226 VDD.n2963 VDD.n2946 1997.65
R10227 VDD.n2999 VDD.n2989 1997.65
R10228 VDD.n2994 VDD.n2989 1997.65
R10229 VDD.n3221 VDD.n3203 1997.65
R10230 VDD.n3221 VDD.n3204 1997.65
R10231 VDD.n3257 VDD.n3247 1997.65
R10232 VDD.n3252 VDD.n3247 1997.65
R10233 VDD.n3479 VDD.n3461 1997.65
R10234 VDD.n3479 VDD.n3462 1997.65
R10235 VDD.n3515 VDD.n3505 1997.65
R10236 VDD.n3510 VDD.n3505 1997.65
R10237 VDD.n5806 VDD.n5788 1997.65
R10238 VDD.n5806 VDD.n5789 1997.65
R10239 VDD.n5842 VDD.n5832 1997.65
R10240 VDD.n5837 VDD.n5832 1997.65
R10241 VDD.n5552 VDD.n5534 1997.65
R10242 VDD.n5552 VDD.n5535 1997.65
R10243 VDD.n5588 VDD.n5578 1997.65
R10244 VDD.n5583 VDD.n5578 1997.65
R10245 VDD.n3737 VDD.n3719 1997.65
R10246 VDD.n3737 VDD.n3720 1997.65
R10247 VDD.n3773 VDD.n3763 1997.65
R10248 VDD.n3768 VDD.n3763 1997.65
R10249 VDD.n3995 VDD.n3977 1997.65
R10250 VDD.n3995 VDD.n3978 1997.65
R10251 VDD.n4031 VDD.n4021 1997.65
R10252 VDD.n4026 VDD.n4021 1997.65
R10253 VDD.n4253 VDD.n4235 1997.65
R10254 VDD.n4253 VDD.n4236 1997.65
R10255 VDD.n4289 VDD.n4279 1997.65
R10256 VDD.n4284 VDD.n4279 1997.65
R10257 VDD.n4511 VDD.n4493 1997.65
R10258 VDD.n4511 VDD.n4494 1997.65
R10259 VDD.n4547 VDD.n4537 1997.65
R10260 VDD.n4542 VDD.n4537 1997.65
R10261 VDD.n4769 VDD.n4751 1997.65
R10262 VDD.n4769 VDD.n4752 1997.65
R10263 VDD.n4805 VDD.n4795 1997.65
R10264 VDD.n4800 VDD.n4795 1997.65
R10265 VDD.n5066 VDD.n5056 1997.65
R10266 VDD.n5061 VDD.n5056 1997.65
R10267 VDD.n5030 VDD.n5012 1997.65
R10268 VDD.n5030 VDD.n5013 1997.65
R10269 VDD.n5328 VDD.n5318 1997.65
R10270 VDD.n5323 VDD.n5318 1997.65
R10271 VDD.n5292 VDD.n5274 1997.65
R10272 VDD.n5292 VDD.n5275 1997.65
R10273 VDD.n1878 VDD.n1819 1814.12
R10274 VDD.n2199 VDD.n2140 1814.12
R10275 VDD.n2457 VDD.n2398 1814.12
R10276 VDD.n2715 VDD.n2656 1814.12
R10277 VDD.n2973 VDD.n2914 1814.12
R10278 VDD.n3231 VDD.n3172 1814.12
R10279 VDD.n3489 VDD.n3430 1814.12
R10280 VDD.n5816 VDD.n5757 1814.12
R10281 VDD.n5562 VDD.n5503 1814.12
R10282 VDD.n3747 VDD.n3688 1814.12
R10283 VDD.n4005 VDD.n3946 1814.12
R10284 VDD.n4263 VDD.n4204 1814.12
R10285 VDD.n4521 VDD.n4462 1814.12
R10286 VDD.n4779 VDD.n4720 1814.12
R10287 VDD.n5040 VDD.n4981 1814.12
R10288 VDD.n5302 VDD.n5243 1814.12
R10289 VDD.n1881 VDD.n1880 1598.82
R10290 VDD.n2202 VDD.n2201 1598.82
R10291 VDD.n2460 VDD.n2459 1598.82
R10292 VDD.n2718 VDD.n2717 1598.82
R10293 VDD.n2976 VDD.n2975 1598.82
R10294 VDD.n3234 VDD.n3233 1598.82
R10295 VDD.n3492 VDD.n3491 1598.82
R10296 VDD.n5819 VDD.n5818 1598.82
R10297 VDD.n5565 VDD.n5564 1598.82
R10298 VDD.n3750 VDD.n3749 1598.82
R10299 VDD.n4008 VDD.n4007 1598.82
R10300 VDD.n4266 VDD.n4265 1598.82
R10301 VDD.n4524 VDD.n4523 1598.82
R10302 VDD.n4782 VDD.n4781 1598.82
R10303 VDD.n5043 VDD.n5042 1598.82
R10304 VDD.n5305 VDD.n5304 1598.82
R10305 VDD.n1698 VDD.n1697 1514.12
R10306 VDD.n2047 VDD.n2046 1514.12
R10307 VDD.n2277 VDD.n2276 1514.12
R10308 VDD.n2535 VDD.n2534 1514.12
R10309 VDD.n2793 VDD.n2792 1514.12
R10310 VDD.n3051 VDD.n3050 1514.12
R10311 VDD.n3309 VDD.n3308 1514.12
R10312 VDD.n5639 VDD.n5638 1514.12
R10313 VDD.n5385 VDD.n5384 1514.12
R10314 VDD.n3567 VDD.n3566 1514.12
R10315 VDD.n3825 VDD.n3824 1514.12
R10316 VDD.n4083 VDD.n4082 1514.12
R10317 VDD.n4341 VDD.n4340 1514.12
R10318 VDD.n4599 VDD.n4598 1514.12
R10319 VDD.n4857 VDD.n4856 1514.12
R10320 VDD.n5149 VDD.n5148 1514.12
R10321 VDD.n1856 VDD.n1844 1440
R10322 VDD.n1869 VDD.n1846 1440
R10323 VDD.n2177 VDD.n2165 1440
R10324 VDD.n2190 VDD.n2167 1440
R10325 VDD.n2435 VDD.n2423 1440
R10326 VDD.n2448 VDD.n2425 1440
R10327 VDD.n2693 VDD.n2681 1440
R10328 VDD.n2706 VDD.n2683 1440
R10329 VDD.n2951 VDD.n2939 1440
R10330 VDD.n2964 VDD.n2941 1440
R10331 VDD.n3209 VDD.n3197 1440
R10332 VDD.n3222 VDD.n3199 1440
R10333 VDD.n3467 VDD.n3455 1440
R10334 VDD.n3480 VDD.n3457 1440
R10335 VDD.n5794 VDD.n5782 1440
R10336 VDD.n5807 VDD.n5784 1440
R10337 VDD.n5540 VDD.n5528 1440
R10338 VDD.n5553 VDD.n5530 1440
R10339 VDD.n3725 VDD.n3713 1440
R10340 VDD.n3738 VDD.n3715 1440
R10341 VDD.n3983 VDD.n3971 1440
R10342 VDD.n3996 VDD.n3973 1440
R10343 VDD.n4241 VDD.n4229 1440
R10344 VDD.n4254 VDD.n4231 1440
R10345 VDD.n4499 VDD.n4487 1440
R10346 VDD.n4512 VDD.n4489 1440
R10347 VDD.n4757 VDD.n4745 1440
R10348 VDD.n4770 VDD.n4747 1440
R10349 VDD.n5018 VDD.n5006 1440
R10350 VDD.n5031 VDD.n5008 1440
R10351 VDD.n5280 VDD.n5268 1440
R10352 VDD.n5293 VDD.n5270 1440
R10353 VDD.n1915 VDD.n1890 1422.35
R10354 VDD.n1900 VDD.n1891 1422.35
R10355 VDD.n2236 VDD.n2211 1422.35
R10356 VDD.n2221 VDD.n2212 1422.35
R10357 VDD.n2494 VDD.n2469 1422.35
R10358 VDD.n2479 VDD.n2470 1422.35
R10359 VDD.n2752 VDD.n2727 1422.35
R10360 VDD.n2737 VDD.n2728 1422.35
R10361 VDD.n3010 VDD.n2985 1422.35
R10362 VDD.n2995 VDD.n2986 1422.35
R10363 VDD.n3268 VDD.n3243 1422.35
R10364 VDD.n3253 VDD.n3244 1422.35
R10365 VDD.n3526 VDD.n3501 1422.35
R10366 VDD.n3511 VDD.n3502 1422.35
R10367 VDD.n5853 VDD.n5828 1422.35
R10368 VDD.n5838 VDD.n5829 1422.35
R10369 VDD.n5599 VDD.n5574 1422.35
R10370 VDD.n5584 VDD.n5575 1422.35
R10371 VDD.n3784 VDD.n3759 1422.35
R10372 VDD.n3769 VDD.n3760 1422.35
R10373 VDD.n4042 VDD.n4017 1422.35
R10374 VDD.n4027 VDD.n4018 1422.35
R10375 VDD.n4300 VDD.n4275 1422.35
R10376 VDD.n4285 VDD.n4276 1422.35
R10377 VDD.n4558 VDD.n4533 1422.35
R10378 VDD.n4543 VDD.n4534 1422.35
R10379 VDD.n4816 VDD.n4791 1422.35
R10380 VDD.n4801 VDD.n4792 1422.35
R10381 VDD.n5077 VDD.n5052 1422.35
R10382 VDD.n5062 VDD.n5053 1422.35
R10383 VDD.n5339 VDD.n5314 1422.35
R10384 VDD.n5324 VDD.n5315 1422.35
R10385 VDD.n1174 VDD 1319.65
R10386 VDD.n1240 VDD 1319.65
R10387 VDD.n1713 VDD.n1676 1231.76
R10388 VDD.n2062 VDD.n2025 1231.76
R10389 VDD.n2292 VDD.n2255 1231.76
R10390 VDD.n2550 VDD.n2513 1231.76
R10391 VDD.n2808 VDD.n2771 1231.76
R10392 VDD.n3066 VDD.n3029 1231.76
R10393 VDD.n3324 VDD.n3287 1231.76
R10394 VDD.n5654 VDD.n5617 1231.76
R10395 VDD.n5400 VDD.n5363 1231.76
R10396 VDD.n3582 VDD.n3545 1231.76
R10397 VDD.n3840 VDD.n3803 1231.76
R10398 VDD.n4098 VDD.n4061 1231.76
R10399 VDD.n4356 VDD.n4319 1231.76
R10400 VDD.n4614 VDD.n4577 1231.76
R10401 VDD.n4872 VDD.n4835 1231.76
R10402 VDD.n5164 VDD.n5127 1231.76
R10403 VDD.n1765 VDD.n1674 1228.24
R10404 VDD.n2114 VDD.n2023 1228.24
R10405 VDD.n2344 VDD.n2253 1228.24
R10406 VDD.n2602 VDD.n2511 1228.24
R10407 VDD.n2860 VDD.n2769 1228.24
R10408 VDD.n3118 VDD.n3027 1228.24
R10409 VDD.n3376 VDD.n3285 1228.24
R10410 VDD.n5706 VDD.n5615 1228.24
R10411 VDD.n5452 VDD.n5361 1228.24
R10412 VDD.n3634 VDD.n3543 1228.24
R10413 VDD.n3892 VDD.n3801 1228.24
R10414 VDD.n4150 VDD.n4059 1228.24
R10415 VDD.n4408 VDD.n4317 1228.24
R10416 VDD.n4666 VDD.n4575 1228.24
R10417 VDD.n4924 VDD.n4833 1228.24
R10418 VDD.n5216 VDD.n5125 1228.24
R10419 VDD.n1765 VDD.n1675 1224.71
R10420 VDD.n1676 VDD.n1675 1224.71
R10421 VDD.n2114 VDD.n2024 1224.71
R10422 VDD.n2025 VDD.n2024 1224.71
R10423 VDD.n2344 VDD.n2254 1224.71
R10424 VDD.n2255 VDD.n2254 1224.71
R10425 VDD.n2602 VDD.n2512 1224.71
R10426 VDD.n2513 VDD.n2512 1224.71
R10427 VDD.n2860 VDD.n2770 1224.71
R10428 VDD.n2771 VDD.n2770 1224.71
R10429 VDD.n3118 VDD.n3028 1224.71
R10430 VDD.n3029 VDD.n3028 1224.71
R10431 VDD.n3376 VDD.n3286 1224.71
R10432 VDD.n3287 VDD.n3286 1224.71
R10433 VDD.n5706 VDD.n5616 1224.71
R10434 VDD.n5617 VDD.n5616 1224.71
R10435 VDD.n5452 VDD.n5362 1224.71
R10436 VDD.n5363 VDD.n5362 1224.71
R10437 VDD.n3634 VDD.n3544 1224.71
R10438 VDD.n3545 VDD.n3544 1224.71
R10439 VDD.n3892 VDD.n3802 1224.71
R10440 VDD.n3803 VDD.n3802 1224.71
R10441 VDD.n4150 VDD.n4060 1224.71
R10442 VDD.n4061 VDD.n4060 1224.71
R10443 VDD.n4408 VDD.n4318 1224.71
R10444 VDD.n4319 VDD.n4318 1224.71
R10445 VDD.n4666 VDD.n4576 1224.71
R10446 VDD.n4577 VDD.n4576 1224.71
R10447 VDD.n4924 VDD.n4834 1224.71
R10448 VDD.n4835 VDD.n4834 1224.71
R10449 VDD.n5216 VDD.n5126 1224.71
R10450 VDD.n5127 VDD.n5126 1224.71
R10451 VDD.n1718 VDD.n1675 1153.33
R10452 VDD.n2067 VDD.n2024 1153.33
R10453 VDD.n2297 VDD.n2254 1153.33
R10454 VDD.n2555 VDD.n2512 1153.33
R10455 VDD.n2813 VDD.n2770 1153.33
R10456 VDD.n3071 VDD.n3028 1153.33
R10457 VDD.n3329 VDD.n3286 1153.33
R10458 VDD.n5659 VDD.n5616 1153.33
R10459 VDD.n5405 VDD.n5362 1153.33
R10460 VDD.n3587 VDD.n3544 1153.33
R10461 VDD.n3845 VDD.n3802 1153.33
R10462 VDD.n4103 VDD.n4060 1153.33
R10463 VDD.n4361 VDD.n4318 1153.33
R10464 VDD.n4619 VDD.n4576 1153.33
R10465 VDD.n4877 VDD.n4834 1153.33
R10466 VDD.n5169 VDD.n5126 1153.33
R10467 VDD.n1902 VDD.n1900 1143.53
R10468 VDD.n2223 VDD.n2221 1143.53
R10469 VDD.n2481 VDD.n2479 1143.53
R10470 VDD.n2739 VDD.n2737 1143.53
R10471 VDD.n2997 VDD.n2995 1143.53
R10472 VDD.n3255 VDD.n3253 1143.53
R10473 VDD.n3513 VDD.n3511 1143.53
R10474 VDD.n5840 VDD.n5838 1143.53
R10475 VDD.n5586 VDD.n5584 1143.53
R10476 VDD.n3771 VDD.n3769 1143.53
R10477 VDD.n4029 VDD.n4027 1143.53
R10478 VDD.n4287 VDD.n4285 1143.53
R10479 VDD.n4545 VDD.n4543 1143.53
R10480 VDD.n4803 VDD.n4801 1143.53
R10481 VDD.n5064 VDD.n5062 1143.53
R10482 VDD.n5326 VDD.n5324 1143.53
R10483 VDD.n1862 VDD.n1846 1125.88
R10484 VDD.n2183 VDD.n2167 1125.88
R10485 VDD.n2441 VDD.n2425 1125.88
R10486 VDD.n2699 VDD.n2683 1125.88
R10487 VDD.n2957 VDD.n2941 1125.88
R10488 VDD.n3215 VDD.n3199 1125.88
R10489 VDD.n3473 VDD.n3457 1125.88
R10490 VDD.n5800 VDD.n5784 1125.88
R10491 VDD.n5546 VDD.n5530 1125.88
R10492 VDD.n3731 VDD.n3715 1125.88
R10493 VDD.n3989 VDD.n3973 1125.88
R10494 VDD.n4247 VDD.n4231 1125.88
R10495 VDD.n4505 VDD.n4489 1125.88
R10496 VDD.n4763 VDD.n4747 1125.88
R10497 VDD.n5024 VDD.n5008 1125.88
R10498 VDD.n5286 VDD.n5270 1125.88
R10499 VDD.n1756 VDD.n1718 1072.94
R10500 VDD.n2105 VDD.n2067 1072.94
R10501 VDD.n2335 VDD.n2297 1072.94
R10502 VDD.n2593 VDD.n2555 1072.94
R10503 VDD.n2851 VDD.n2813 1072.94
R10504 VDD.n3109 VDD.n3071 1072.94
R10505 VDD.n3367 VDD.n3329 1072.94
R10506 VDD.n5697 VDD.n5659 1072.94
R10507 VDD.n5443 VDD.n5405 1072.94
R10508 VDD.n3625 VDD.n3587 1072.94
R10509 VDD.n3883 VDD.n3845 1072.94
R10510 VDD.n4141 VDD.n4103 1072.94
R10511 VDD.n4399 VDD.n4361 1072.94
R10512 VDD.n4657 VDD.n4619 1072.94
R10513 VDD.n4915 VDD.n4877 1072.94
R10514 VDD.n5207 VDD.n5169 1072.94
R10515 VDD.n1718 VDD.n1670 1069.41
R10516 VDD.n2067 VDD.n2019 1069.41
R10517 VDD.n2297 VDD.n2249 1069.41
R10518 VDD.n2555 VDD.n2507 1069.41
R10519 VDD.n2813 VDD.n2765 1069.41
R10520 VDD.n3071 VDD.n3023 1069.41
R10521 VDD.n3329 VDD.n3281 1069.41
R10522 VDD.n5659 VDD.n5611 1069.41
R10523 VDD.n5405 VDD.n5357 1069.41
R10524 VDD.n3587 VDD.n3539 1069.41
R10525 VDD.n3845 VDD.n3797 1069.41
R10526 VDD.n4103 VDD.n4055 1069.41
R10527 VDD.n4361 VDD.n4313 1069.41
R10528 VDD.n4619 VDD.n4571 1069.41
R10529 VDD.n4877 VDD.n4829 1069.41
R10530 VDD.n5169 VDD.n5121 1069.41
R10531 VDD.n1906 VDD.n1890 1051.76
R10532 VDD.n1856 VDD.n1855 1051.76
R10533 VDD.n2177 VDD.n2176 1051.76
R10534 VDD.n2227 VDD.n2211 1051.76
R10535 VDD.n2435 VDD.n2434 1051.76
R10536 VDD.n2485 VDD.n2469 1051.76
R10537 VDD.n2693 VDD.n2692 1051.76
R10538 VDD.n2743 VDD.n2727 1051.76
R10539 VDD.n2951 VDD.n2950 1051.76
R10540 VDD.n3001 VDD.n2985 1051.76
R10541 VDD.n3209 VDD.n3208 1051.76
R10542 VDD.n3259 VDD.n3243 1051.76
R10543 VDD.n3467 VDD.n3466 1051.76
R10544 VDD.n3517 VDD.n3501 1051.76
R10545 VDD.n5794 VDD.n5793 1051.76
R10546 VDD.n5844 VDD.n5828 1051.76
R10547 VDD.n5540 VDD.n5539 1051.76
R10548 VDD.n5590 VDD.n5574 1051.76
R10549 VDD.n3725 VDD.n3724 1051.76
R10550 VDD.n3775 VDD.n3759 1051.76
R10551 VDD.n3983 VDD.n3982 1051.76
R10552 VDD.n4033 VDD.n4017 1051.76
R10553 VDD.n4241 VDD.n4240 1051.76
R10554 VDD.n4291 VDD.n4275 1051.76
R10555 VDD.n4499 VDD.n4498 1051.76
R10556 VDD.n4549 VDD.n4533 1051.76
R10557 VDD.n4757 VDD.n4756 1051.76
R10558 VDD.n4807 VDD.n4791 1051.76
R10559 VDD.n5068 VDD.n5052 1051.76
R10560 VDD.n5018 VDD.n5017 1051.76
R10561 VDD.n5330 VDD.n5314 1051.76
R10562 VDD.n5280 VDD.n5279 1051.76
R10563 VDD.n1960 VDD.n1942 862.871
R10564 VDD.n1950 VDD.n1942 862.871
R10565 VDD.n1971 VDD.n1930 862.871
R10566 VDD.n1967 VDD.n1930 862.871
R10567 VDD.n1759 VDD.n1758 861.178
R10568 VDD.n2108 VDD.n2107 861.178
R10569 VDD.n2338 VDD.n2337 861.178
R10570 VDD.n2596 VDD.n2595 861.178
R10571 VDD.n2854 VDD.n2853 861.178
R10572 VDD.n3112 VDD.n3111 861.178
R10573 VDD.n3370 VDD.n3369 861.178
R10574 VDD.n5700 VDD.n5699 861.178
R10575 VDD.n5446 VDD.n5445 861.178
R10576 VDD.n3628 VDD.n3627 861.178
R10577 VDD.n3886 VDD.n3885 861.178
R10578 VDD.n4144 VDD.n4143 861.178
R10579 VDD.n4402 VDD.n4401 861.178
R10580 VDD.n4660 VDD.n4659 861.178
R10581 VDD.n4918 VDD.n4917 861.178
R10582 VDD.n5210 VDD.n5209 861.178
R10583 VDD.n1962 VDD.n1961 857.648
R10584 VDD.n1963 VDD.n1962 857.648
R10585 VDD.n1963 VDD.n1928 857.648
R10586 VDD.n1970 VDD.n1928 857.648
R10587 VDD.n1951 VDD.n1938 857.648
R10588 VDD.n1964 VDD.n1938 857.648
R10589 VDD.n1964 VDD.n1932 857.648
R10590 VDD.n1968 VDD.n1932 857.648
R10591 VDD.n1883 VDD.n1819 751.765
R10592 VDD.n2204 VDD.n2140 751.765
R10593 VDD.n2462 VDD.n2398 751.765
R10594 VDD.n2720 VDD.n2656 751.765
R10595 VDD.n2978 VDD.n2914 751.765
R10596 VDD.n3236 VDD.n3172 751.765
R10597 VDD.n3494 VDD.n3430 751.765
R10598 VDD.n5821 VDD.n5757 751.765
R10599 VDD.n5567 VDD.n5503 751.765
R10600 VDD.n3752 VDD.n3688 751.765
R10601 VDD.n4010 VDD.n3946 751.765
R10602 VDD.n4268 VDD.n4204 751.765
R10603 VDD.n4526 VDD.n4462 751.765
R10604 VDD.n4784 VDD.n4720 751.765
R10605 VDD.n5045 VDD.n4981 751.765
R10606 VDD.n5307 VDD.n5243 751.765
R10607 VDD.n1714 VDD.n1712 723.529
R10608 VDD.n2063 VDD.n2061 723.529
R10609 VDD.n2293 VDD.n2291 723.529
R10610 VDD.n2551 VDD.n2549 723.529
R10611 VDD.n2809 VDD.n2807 723.529
R10612 VDD.n3067 VDD.n3065 723.529
R10613 VDD.n3325 VDD.n3323 723.529
R10614 VDD.n5655 VDD.n5653 723.529
R10615 VDD.n5401 VDD.n5399 723.529
R10616 VDD.n3583 VDD.n3581 723.529
R10617 VDD.n3841 VDD.n3839 723.529
R10618 VDD.n4099 VDD.n4097 723.529
R10619 VDD.n4357 VDD.n4355 723.529
R10620 VDD.n4615 VDD.n4613 723.529
R10621 VDD.n4873 VDD.n4871 723.529
R10622 VDD.n5165 VDD.n5163 723.529
R10623 VDD.n1680 VDD.n1678 720
R10624 VDD.n2029 VDD.n2027 720
R10625 VDD.n2259 VDD.n2257 720
R10626 VDD.n2517 VDD.n2515 720
R10627 VDD.n2775 VDD.n2773 720
R10628 VDD.n3033 VDD.n3031 720
R10629 VDD.n3291 VDD.n3289 720
R10630 VDD.n5621 VDD.n5619 720
R10631 VDD.n5367 VDD.n5365 720
R10632 VDD.n3549 VDD.n3547 720
R10633 VDD.n3807 VDD.n3805 720
R10634 VDD.n4065 VDD.n4063 720
R10635 VDD.n4323 VDD.n4321 720
R10636 VDD.n4581 VDD.n4579 720
R10637 VDD.n4839 VDD.n4837 720
R10638 VDD.n5131 VDD.n5129 720
R10639 VDD.n1695 VDD.t1227 632.183
R10640 VDD.n2044 VDD.t29 632.183
R10641 VDD.n2274 VDD.t541 632.183
R10642 VDD.n2532 VDD.t472 632.183
R10643 VDD.n2790 VDD.t1309 632.183
R10644 VDD.n3048 VDD.t6 632.183
R10645 VDD.n3306 VDD.t1194 632.183
R10646 VDD.n5636 VDD.t707 632.183
R10647 VDD.n5382 VDD.t1331 632.183
R10648 VDD.n3564 VDD.t1268 632.183
R10649 VDD.n3822 VDD.t81 632.183
R10650 VDD.n4080 VDD.t723 632.183
R10651 VDD.n4338 VDD.t1112 632.183
R10652 VDD.n4596 VDD.t183 632.183
R10653 VDD.n4854 VDD.t1121 632.183
R10654 VDD.n5146 VDD.t195 632.183
R10655 VDD.n1677 VDD.n1674 593.144
R10656 VDD.n1680 VDD.n1677 593.144
R10657 VDD.n2026 VDD.n2023 593.144
R10658 VDD.n2029 VDD.n2026 593.144
R10659 VDD.n2256 VDD.n2253 593.144
R10660 VDD.n2259 VDD.n2256 593.144
R10661 VDD.n2514 VDD.n2511 593.144
R10662 VDD.n2517 VDD.n2514 593.144
R10663 VDD.n2772 VDD.n2769 593.144
R10664 VDD.n2775 VDD.n2772 593.144
R10665 VDD.n3030 VDD.n3027 593.144
R10666 VDD.n3033 VDD.n3030 593.144
R10667 VDD.n3288 VDD.n3285 593.144
R10668 VDD.n3291 VDD.n3288 593.144
R10669 VDD.n5618 VDD.n5615 593.144
R10670 VDD.n5621 VDD.n5618 593.144
R10671 VDD.n5364 VDD.n5361 593.144
R10672 VDD.n5367 VDD.n5364 593.144
R10673 VDD.n3546 VDD.n3543 593.144
R10674 VDD.n3549 VDD.n3546 593.144
R10675 VDD.n3804 VDD.n3801 593.144
R10676 VDD.n3807 VDD.n3804 593.144
R10677 VDD.n4062 VDD.n4059 593.144
R10678 VDD.n4065 VDD.n4062 593.144
R10679 VDD.n4320 VDD.n4317 593.144
R10680 VDD.n4323 VDD.n4320 593.144
R10681 VDD.n4578 VDD.n4575 593.144
R10682 VDD.n4581 VDD.n4578 593.144
R10683 VDD.n4836 VDD.n4833 593.144
R10684 VDD.n4839 VDD.n4836 593.144
R10685 VDD.n5128 VDD.n5125 593.144
R10686 VDD.n5131 VDD.n5128 593.144
R10687 VDD.n1795 VDD.t41 584.644
R10688 VDD.n1781 VDD.t1231 584.644
R10689 VDD.n2003 VDD.t369 584.644
R10690 VDD.n1989 VDD.t33 584.644
R10691 VDD.n2374 VDD.t471 584.644
R10692 VDD.n2360 VDD.t540 584.644
R10693 VDD.n2632 VDD.t123 584.644
R10694 VDD.n2618 VDD.t479 584.644
R10695 VDD.n2890 VDD.t26 584.644
R10696 VDD.n2876 VDD.t1312 584.644
R10697 VDD.n3148 VDD.t595 584.644
R10698 VDD.n3134 VDD.t10 584.644
R10699 VDD.n3406 VDD.t555 584.644
R10700 VDD.n3392 VDD.t1201 584.644
R10701 VDD.n5736 VDD.t175 584.644
R10702 VDD.n5722 VDD.t711 584.644
R10703 VDD.n5482 VDD.t761 584.644
R10704 VDD.n5468 VDD.t1330 584.644
R10705 VDD.n3664 VDD.t1098 584.644
R10706 VDD.n3650 VDD.t1275 584.644
R10707 VDD.n3922 VDD.t788 584.644
R10708 VDD.n3908 VDD.t80 584.644
R10709 VDD.n4180 VDD.t494 584.644
R10710 VDD.n4166 VDD.t722 584.644
R10711 VDD.n4438 VDD.t379 584.644
R10712 VDD.n4424 VDD.t1115 584.644
R10713 VDD.n4696 VDD.t116 584.644
R10714 VDD.n4682 VDD.t187 584.644
R10715 VDD.n4955 VDD.t354 584.644
R10716 VDD.n4941 VDD.t1128 584.644
R10717 VDD.n5105 VDD.t487 584.644
R10718 VDD.n5091 VDD.t198 584.644
R10719 VDD.n840 VDD.t1292 584.644
R10720 VDD.n45 VDD.t65 584.644
R10721 VDD.n439 VDD.t1074 584.644
R10722 VDD.n1348 VDD.t400 584.644
R10723 VDD.n1763 VDD.n1713 576.668
R10724 VDD.n1763 VDD.n1714 576.668
R10725 VDD.n2112 VDD.n2062 576.668
R10726 VDD.n2112 VDD.n2063 576.668
R10727 VDD.n2342 VDD.n2292 576.668
R10728 VDD.n2342 VDD.n2293 576.668
R10729 VDD.n2600 VDD.n2550 576.668
R10730 VDD.n2600 VDD.n2551 576.668
R10731 VDD.n2858 VDD.n2808 576.668
R10732 VDD.n2858 VDD.n2809 576.668
R10733 VDD.n3116 VDD.n3066 576.668
R10734 VDD.n3116 VDD.n3067 576.668
R10735 VDD.n3374 VDD.n3324 576.668
R10736 VDD.n3374 VDD.n3325 576.668
R10737 VDD.n5704 VDD.n5654 576.668
R10738 VDD.n5704 VDD.n5655 576.668
R10739 VDD.n5450 VDD.n5400 576.668
R10740 VDD.n5450 VDD.n5401 576.668
R10741 VDD.n3632 VDD.n3582 576.668
R10742 VDD.n3632 VDD.n3583 576.668
R10743 VDD.n3890 VDD.n3840 576.668
R10744 VDD.n3890 VDD.n3841 576.668
R10745 VDD.n4148 VDD.n4098 576.668
R10746 VDD.n4148 VDD.n4099 576.668
R10747 VDD.n4406 VDD.n4356 576.668
R10748 VDD.n4406 VDD.n4357 576.668
R10749 VDD.n4664 VDD.n4614 576.668
R10750 VDD.n4664 VDD.n4615 576.668
R10751 VDD.n4922 VDD.n4872 576.668
R10752 VDD.n4922 VDD.n4873 576.668
R10753 VDD.n5214 VDD.n5164 576.668
R10754 VDD.n5214 VDD.n5165 576.668
R10755 VDD.n1906 VDD.n1904 568.236
R10756 VDD.n1899 VDD.n1896 568.236
R10757 VDD.n1902 VDD.n1899 568.236
R10758 VDD.n1904 VDD.n1895 568.236
R10759 VDD.n1859 VDD.n1850 568.236
R10760 VDD.n1862 VDD.n1851 568.236
R10761 VDD.n1864 VDD.n1851 568.236
R10762 VDD.n1855 VDD.n1850 568.236
R10763 VDD.n2180 VDD.n2171 568.236
R10764 VDD.n2183 VDD.n2172 568.236
R10765 VDD.n2185 VDD.n2172 568.236
R10766 VDD.n2176 VDD.n2171 568.236
R10767 VDD.n2227 VDD.n2225 568.236
R10768 VDD.n2220 VDD.n2217 568.236
R10769 VDD.n2223 VDD.n2220 568.236
R10770 VDD.n2225 VDD.n2216 568.236
R10771 VDD.n2438 VDD.n2429 568.236
R10772 VDD.n2441 VDD.n2430 568.236
R10773 VDD.n2443 VDD.n2430 568.236
R10774 VDD.n2434 VDD.n2429 568.236
R10775 VDD.n2485 VDD.n2483 568.236
R10776 VDD.n2478 VDD.n2475 568.236
R10777 VDD.n2481 VDD.n2478 568.236
R10778 VDD.n2483 VDD.n2474 568.236
R10779 VDD.n2696 VDD.n2687 568.236
R10780 VDD.n2699 VDD.n2688 568.236
R10781 VDD.n2701 VDD.n2688 568.236
R10782 VDD.n2692 VDD.n2687 568.236
R10783 VDD.n2743 VDD.n2741 568.236
R10784 VDD.n2736 VDD.n2733 568.236
R10785 VDD.n2739 VDD.n2736 568.236
R10786 VDD.n2741 VDD.n2732 568.236
R10787 VDD.n2954 VDD.n2945 568.236
R10788 VDD.n2957 VDD.n2946 568.236
R10789 VDD.n2959 VDD.n2946 568.236
R10790 VDD.n2950 VDD.n2945 568.236
R10791 VDD.n3001 VDD.n2999 568.236
R10792 VDD.n2994 VDD.n2991 568.236
R10793 VDD.n2997 VDD.n2994 568.236
R10794 VDD.n2999 VDD.n2990 568.236
R10795 VDD.n3212 VDD.n3203 568.236
R10796 VDD.n3215 VDD.n3204 568.236
R10797 VDD.n3217 VDD.n3204 568.236
R10798 VDD.n3208 VDD.n3203 568.236
R10799 VDD.n3259 VDD.n3257 568.236
R10800 VDD.n3252 VDD.n3249 568.236
R10801 VDD.n3255 VDD.n3252 568.236
R10802 VDD.n3257 VDD.n3248 568.236
R10803 VDD.n3470 VDD.n3461 568.236
R10804 VDD.n3473 VDD.n3462 568.236
R10805 VDD.n3475 VDD.n3462 568.236
R10806 VDD.n3466 VDD.n3461 568.236
R10807 VDD.n3517 VDD.n3515 568.236
R10808 VDD.n3510 VDD.n3507 568.236
R10809 VDD.n3513 VDD.n3510 568.236
R10810 VDD.n3515 VDD.n3506 568.236
R10811 VDD.n5797 VDD.n5788 568.236
R10812 VDD.n5800 VDD.n5789 568.236
R10813 VDD.n5802 VDD.n5789 568.236
R10814 VDD.n5793 VDD.n5788 568.236
R10815 VDD.n5844 VDD.n5842 568.236
R10816 VDD.n5837 VDD.n5834 568.236
R10817 VDD.n5840 VDD.n5837 568.236
R10818 VDD.n5842 VDD.n5833 568.236
R10819 VDD.n5543 VDD.n5534 568.236
R10820 VDD.n5546 VDD.n5535 568.236
R10821 VDD.n5548 VDD.n5535 568.236
R10822 VDD.n5539 VDD.n5534 568.236
R10823 VDD.n5590 VDD.n5588 568.236
R10824 VDD.n5583 VDD.n5580 568.236
R10825 VDD.n5586 VDD.n5583 568.236
R10826 VDD.n5588 VDD.n5579 568.236
R10827 VDD.n3728 VDD.n3719 568.236
R10828 VDD.n3731 VDD.n3720 568.236
R10829 VDD.n3733 VDD.n3720 568.236
R10830 VDD.n3724 VDD.n3719 568.236
R10831 VDD.n3775 VDD.n3773 568.236
R10832 VDD.n3768 VDD.n3765 568.236
R10833 VDD.n3771 VDD.n3768 568.236
R10834 VDD.n3773 VDD.n3764 568.236
R10835 VDD.n3986 VDD.n3977 568.236
R10836 VDD.n3989 VDD.n3978 568.236
R10837 VDD.n3991 VDD.n3978 568.236
R10838 VDD.n3982 VDD.n3977 568.236
R10839 VDD.n4033 VDD.n4031 568.236
R10840 VDD.n4026 VDD.n4023 568.236
R10841 VDD.n4029 VDD.n4026 568.236
R10842 VDD.n4031 VDD.n4022 568.236
R10843 VDD.n4244 VDD.n4235 568.236
R10844 VDD.n4247 VDD.n4236 568.236
R10845 VDD.n4249 VDD.n4236 568.236
R10846 VDD.n4240 VDD.n4235 568.236
R10847 VDD.n4291 VDD.n4289 568.236
R10848 VDD.n4284 VDD.n4281 568.236
R10849 VDD.n4287 VDD.n4284 568.236
R10850 VDD.n4289 VDD.n4280 568.236
R10851 VDD.n4502 VDD.n4493 568.236
R10852 VDD.n4505 VDD.n4494 568.236
R10853 VDD.n4507 VDD.n4494 568.236
R10854 VDD.n4498 VDD.n4493 568.236
R10855 VDD.n4549 VDD.n4547 568.236
R10856 VDD.n4542 VDD.n4539 568.236
R10857 VDD.n4545 VDD.n4542 568.236
R10858 VDD.n4547 VDD.n4538 568.236
R10859 VDD.n4760 VDD.n4751 568.236
R10860 VDD.n4763 VDD.n4752 568.236
R10861 VDD.n4765 VDD.n4752 568.236
R10862 VDD.n4756 VDD.n4751 568.236
R10863 VDD.n4807 VDD.n4805 568.236
R10864 VDD.n4800 VDD.n4797 568.236
R10865 VDD.n4803 VDD.n4800 568.236
R10866 VDD.n4805 VDD.n4796 568.236
R10867 VDD.n5068 VDD.n5066 568.236
R10868 VDD.n5061 VDD.n5058 568.236
R10869 VDD.n5064 VDD.n5061 568.236
R10870 VDD.n5066 VDD.n5057 568.236
R10871 VDD.n5021 VDD.n5012 568.236
R10872 VDD.n5024 VDD.n5013 568.236
R10873 VDD.n5026 VDD.n5013 568.236
R10874 VDD.n5017 VDD.n5012 568.236
R10875 VDD.n5330 VDD.n5328 568.236
R10876 VDD.n5323 VDD.n5320 568.236
R10877 VDD.n5326 VDD.n5323 568.236
R10878 VDD.n5328 VDD.n5319 568.236
R10879 VDD.n5283 VDD.n5274 568.236
R10880 VDD.n5286 VDD.n5275 568.236
R10881 VDD.n5288 VDD.n5275 568.236
R10882 VDD.n5279 VDD.n5274 568.236
R10883 VDD.n1174 VDD.t1241 533.735
R10884 VDD.n1240 VDD.t1166 533.735
R10885 VDD.n1744 VDD.n1743 481.226
R10886 VDD.n2093 VDD.n2092 481.226
R10887 VDD.n2323 VDD.n2322 481.226
R10888 VDD.n2581 VDD.n2580 481.226
R10889 VDD.n2839 VDD.n2838 481.226
R10890 VDD.n3097 VDD.n3096 481.226
R10891 VDD.n3355 VDD.n3354 481.226
R10892 VDD.n5685 VDD.n5684 481.226
R10893 VDD.n5431 VDD.n5430 481.226
R10894 VDD.n3613 VDD.n3612 481.226
R10895 VDD.n3871 VDD.n3870 481.226
R10896 VDD.n4129 VDD.n4128 481.226
R10897 VDD.n4387 VDD.n4386 481.226
R10898 VDD.n4645 VDD.n4644 481.226
R10899 VDD.n4903 VDD.n4902 481.226
R10900 VDD.n5195 VDD.n5194 481.226
R10901 VDD.n1857 VDD.n1847 473.839
R10902 VDD.t355 VDD.n1849 473.839
R10903 VDD.n2178 VDD.n2168 473.839
R10904 VDD.t574 VDD.n2170 473.839
R10905 VDD.n2436 VDD.n2426 473.839
R10906 VDD.t103 VDD.n2428 473.839
R10907 VDD.n2694 VDD.n2684 473.839
R10908 VDD.t421 VDD.n2686 473.839
R10909 VDD.n2952 VDD.n2942 473.839
R10910 VDD.t405 VDD.n2944 473.839
R10911 VDD.n3210 VDD.n3200 473.839
R10912 VDD.t144 VDD.n3202 473.839
R10913 VDD.n3468 VDD.n3458 473.839
R10914 VDD.t179 VDD.n3460 473.839
R10915 VDD.n5795 VDD.n5785 473.839
R10916 VDD.t1088 VDD.n5787 473.839
R10917 VDD.n5541 VDD.n5531 473.839
R10918 VDD.t596 VDD.n5533 473.839
R10919 VDD.n3726 VDD.n3716 473.839
R10920 VDD.t145 VDD.n3718 473.839
R10921 VDD.n3984 VDD.n3974 473.839
R10922 VDD.t563 VDD.n3976 473.839
R10923 VDD.n4242 VDD.n4232 473.839
R10924 VDD.t668 VDD.n4234 473.839
R10925 VDD.n4500 VDD.n4490 473.839
R10926 VDD.t561 VDD.n4492 473.839
R10927 VDD.n4758 VDD.n4748 473.839
R10928 VDD.t750 VDD.n4750 473.839
R10929 VDD.n5019 VDD.n5009 473.839
R10930 VDD.t386 VDD.n5011 473.839
R10931 VDD.n5281 VDD.n5271 473.839
R10932 VDD.t559 VDD.n5273 473.839
R10933 VDD.n1914 VDD.n1892 468.033
R10934 VDD.t420 VDD.n1893 468.033
R10935 VDD.n2235 VDD.n2213 468.033
R10936 VDD.t148 VDD.n2214 468.033
R10937 VDD.n2493 VDD.n2471 468.033
R10938 VDD.t676 VDD.n2472 468.033
R10939 VDD.n2751 VDD.n2729 468.033
R10940 VDD.t689 VDD.n2730 468.033
R10941 VDD.n3009 VDD.n2987 468.033
R10942 VDD.t93 VDD.n2988 468.033
R10943 VDD.n3267 VDD.n3245 468.033
R10944 VDD.t76 VDD.n3246 468.033
R10945 VDD.n3525 VDD.n3503 468.033
R10946 VDD.t1186 VDD.n3504 468.033
R10947 VDD.n5852 VDD.n5830 468.033
R10948 VDD.t159 VDD.n5831 468.033
R10949 VDD.n5598 VDD.n5576 468.033
R10950 VDD.t203 VDD.n5577 468.033
R10951 VDD.n3783 VDD.n3761 468.033
R10952 VDD.t556 VDD.n3762 468.033
R10953 VDD.n4041 VDD.n4019 468.033
R10954 VDD.t562 VDD.n4020 468.033
R10955 VDD.n4299 VDD.n4277 468.033
R10956 VDD.t687 VDD.n4278 468.033
R10957 VDD.n4557 VDD.n4535 468.033
R10958 VDD.t570 VDD.n4536 468.033
R10959 VDD.n4815 VDD.n4793 468.033
R10960 VDD.t670 VDD.n4794 468.033
R10961 VDD.n5076 VDD.n5054 468.033
R10962 VDD.t581 VDD.n5055 468.033
R10963 VDD.n5338 VDD.n5316 468.033
R10964 VDD.t97 VDD.n5317 468.033
R10965 VDD.n1933 VDD.n1925 459.009
R10966 VDD.n1935 VDD.n1932 437.647
R10967 VDD.n1974 VDD.n1928 430.589
R10968 VDD.n1962 VDD.n1940 430.589
R10969 VDD.n800 VDD.n799 425.228
R10970 VDD.n398 VDD.n397 425.228
R10971 VDD VDD.t651 421.082
R10972 VDD.n1948 VDD.n1938 420
R10973 VDD.n724 VDD.t745 396.079
R10974 VDD.n1565 VDD.t389 396.079
R10975 VDD.n9 VDD.t1246 382.793
R10976 VDD.n782 VDD.t1239 382.793
R10977 VDD.n729 VDD.t1249 382.793
R10978 VDD.n728 VDD.t1236 382.793
R10979 VDD.n710 VDD.t1235 382.793
R10980 VDD.n380 VDD.t1170 382.793
R10981 VDD.n326 VDD.t1178 382.793
R10982 VDD.n1570 VDD.t1164 382.793
R10983 VDD.n1569 VDD.t1159 382.793
R10984 VDD.n1551 VDD.t1157 382.793
R10985 VDD.n1122 VDD.t90 382.793
R10986 VDD.n1188 VDD.t650 382.793
R10987 VDD VDD.t1256 374.711
R10988 VDD VDD.t702 374.711
R10989 VDD VDD.t791 374.711
R10990 VDD VDD.t1314 374.711
R10991 VDD VDD.t68 374.711
R10992 VDD VDD.t1211 374.711
R10993 VDD.n1709 VDD.n1680 370.589
R10994 VDD.n1759 VDD.n1714 370.589
R10995 VDD.n2058 VDD.n2029 370.589
R10996 VDD.n2108 VDD.n2063 370.589
R10997 VDD.n2288 VDD.n2259 370.589
R10998 VDD.n2338 VDD.n2293 370.589
R10999 VDD.n2546 VDD.n2517 370.589
R11000 VDD.n2596 VDD.n2551 370.589
R11001 VDD.n2804 VDD.n2775 370.589
R11002 VDD.n2854 VDD.n2809 370.589
R11003 VDD.n3062 VDD.n3033 370.589
R11004 VDD.n3112 VDD.n3067 370.589
R11005 VDD.n3320 VDD.n3291 370.589
R11006 VDD.n3370 VDD.n3325 370.589
R11007 VDD.n5650 VDD.n5621 370.589
R11008 VDD.n5700 VDD.n5655 370.589
R11009 VDD.n5396 VDD.n5367 370.589
R11010 VDD.n5446 VDD.n5401 370.589
R11011 VDD.n3578 VDD.n3549 370.589
R11012 VDD.n3628 VDD.n3583 370.589
R11013 VDD.n3836 VDD.n3807 370.589
R11014 VDD.n3886 VDD.n3841 370.589
R11015 VDD.n4094 VDD.n4065 370.589
R11016 VDD.n4144 VDD.n4099 370.589
R11017 VDD.n4352 VDD.n4323 370.589
R11018 VDD.n4402 VDD.n4357 370.589
R11019 VDD.n4610 VDD.n4581 370.589
R11020 VDD.n4660 VDD.n4615 370.589
R11021 VDD.n4868 VDD.n4839 370.589
R11022 VDD.n4918 VDD.n4873 370.589
R11023 VDD.n5160 VDD.n5131 370.589
R11024 VDD.n5210 VDD.n5165 370.589
R11025 VDD.n12 VDD.t334 370.341
R11026 VDD.n790 VDD.t1240 370.341
R11027 VDD.n762 VDD.t177 370.341
R11028 VDD.n763 VDD.t610 370.341
R11029 VDD.n388 VDD.t1172 370.341
R11030 VDD.n359 VDD.t1136 370.341
R11031 VDD.n360 VDD.t743 370.341
R11032 VDD.n329 VDD.t1214 370.341
R11033 VDD VDD.t2 370.303
R11034 VDD VDD.t1322 370.303
R11035 VDD.t753 VDD.t1227 333.365
R11036 VDD.t753 VDD.t37 333.365
R11037 VDD.t129 VDD.t29 333.365
R11038 VDD.t129 VDD.t365 333.365
R11039 VDD.t70 VDD.t541 333.365
R11040 VDD.t70 VDD.t466 333.365
R11041 VDD.t680 VDD.t472 333.365
R11042 VDD.t680 VDD.t117 333.365
R11043 VDD.t733 VDD.t1309 333.365
R11044 VDD.t733 VDD.t21 333.365
R11045 VDD.t125 VDD.t6 333.365
R11046 VDD.t125 VDD.t590 333.365
R11047 VDD.t504 VDD.t1194 333.365
R11048 VDD.t504 VDD.t550 333.365
R11049 VDD.t4 VDD.t707 333.365
R11050 VDD.t4 VDD.t170 333.365
R11051 VDD.t665 VDD.t1331 333.365
R11052 VDD.t665 VDD.t757 333.365
R11053 VDD.t1141 VDD.t1268 333.365
R11054 VDD.t1141 VDD.t1100 333.365
R11055 VDD.t1061 VDD.t81 333.365
R11056 VDD.t1061 VDD.t785 333.365
R11057 VDD.t414 VDD.t723 333.365
R11058 VDD.t414 VDD.t490 333.365
R11059 VDD.t165 VDD.t1112 333.365
R11060 VDD.t165 VDD.t374 333.365
R11061 VDD.t793 VDD.t183 333.365
R11062 VDD.t793 VDD.t111 333.365
R11063 VDD.t1065 VDD.t1121 333.365
R11064 VDD.t1065 VDD.t349 333.365
R11065 VDD.t107 VDD.t195 333.365
R11066 VDD.t107 VDD.t482 333.365
R11067 VDD VDD.t696 331.981
R11068 VDD VDD.t135 331.981
R11069 VDD.n1634 VDD.t1179 330.12
R11070 VDD.n1635 VDD.t1160 330.002
R11071 VDD.n1541 VDD 323.514
R11072 VDD.n1643 VDD.t1171 323.342
R11073 VDD.n34 VDD.t1282 321.801
R11074 VDD.n351 VDD.t1326 321.801
R11075 VDD.n793 VDD.n792 318.678
R11076 VDD.n391 VDD.n390 318.678
R11077 VDD.n828 VDD.t1107 318.108
R11078 VDD.n426 VDD.t729 318.108
R11079 VDD VDD.t1134 313.839
R11080 VDD VDD.t1057 313.839
R11081 VDD VDD.t1304 313.839
R11082 VDD.n8 VDD.n7 307.24
R11083 VDD.n789 VDD.n788 307.24
R11084 VDD.n759 VDD.n758 307.24
R11085 VDD.n761 VDD.n760 307.24
R11086 VDD.n387 VDD.n386 307.24
R11087 VDD.n356 VDD.n355 307.24
R11088 VDD.n358 VDD.n357 307.24
R11089 VDD.n325 VDD.n324 307.24
R11090 VDD.t753 VDD.n1678 298.82
R11091 VDD.t753 VDD.n1712 298.82
R11092 VDD.t129 VDD.n2027 298.82
R11093 VDD.t129 VDD.n2061 298.82
R11094 VDD.t70 VDD.n2257 298.82
R11095 VDD.t70 VDD.n2291 298.82
R11096 VDD.t680 VDD.n2515 298.82
R11097 VDD.t680 VDD.n2549 298.82
R11098 VDD.t733 VDD.n2773 298.82
R11099 VDD.t733 VDD.n2807 298.82
R11100 VDD.t125 VDD.n3031 298.82
R11101 VDD.t125 VDD.n3065 298.82
R11102 VDD.t504 VDD.n3289 298.82
R11103 VDD.t504 VDD.n3323 298.82
R11104 VDD.t4 VDD.n5619 298.82
R11105 VDD.t4 VDD.n5653 298.82
R11106 VDD.t665 VDD.n5365 298.82
R11107 VDD.t665 VDD.n5399 298.82
R11108 VDD.t1141 VDD.n3547 298.82
R11109 VDD.t1141 VDD.n3581 298.82
R11110 VDD.t1061 VDD.n3805 298.82
R11111 VDD.t1061 VDD.n3839 298.82
R11112 VDD.t414 VDD.n4063 298.82
R11113 VDD.t414 VDD.n4097 298.82
R11114 VDD.t165 VDD.n4321 298.82
R11115 VDD.t165 VDD.n4355 298.82
R11116 VDD.t793 VDD.n4579 298.82
R11117 VDD.t793 VDD.n4613 298.82
R11118 VDD.t1065 VDD.n4837 298.82
R11119 VDD.t1065 VDD.n4871 298.82
R11120 VDD.t107 VDD.n5129 298.82
R11121 VDD.t107 VDD.n5163 298.82
R11122 VDD.n1912 VDD.n1897 273.695
R11123 VDD.n1912 VDD.n1911 273.695
R11124 VDD.n1877 VDD.n1824 273.695
R11125 VDD.n1824 VDD.n1822 273.695
R11126 VDD.n1861 VDD.n1860 273.695
R11127 VDD.n1865 VDD.n1861 273.695
R11128 VDD.n2182 VDD.n2181 273.695
R11129 VDD.n2186 VDD.n2182 273.695
R11130 VDD.n2198 VDD.n2145 273.695
R11131 VDD.n2145 VDD.n2143 273.695
R11132 VDD.n2233 VDD.n2218 273.695
R11133 VDD.n2233 VDD.n2232 273.695
R11134 VDD.n2440 VDD.n2439 273.695
R11135 VDD.n2444 VDD.n2440 273.695
R11136 VDD.n2456 VDD.n2403 273.695
R11137 VDD.n2403 VDD.n2401 273.695
R11138 VDD.n2491 VDD.n2476 273.695
R11139 VDD.n2491 VDD.n2490 273.695
R11140 VDD.n2698 VDD.n2697 273.695
R11141 VDD.n2702 VDD.n2698 273.695
R11142 VDD.n2714 VDD.n2661 273.695
R11143 VDD.n2661 VDD.n2659 273.695
R11144 VDD.n2749 VDD.n2734 273.695
R11145 VDD.n2749 VDD.n2748 273.695
R11146 VDD.n2956 VDD.n2955 273.695
R11147 VDD.n2960 VDD.n2956 273.695
R11148 VDD.n2972 VDD.n2919 273.695
R11149 VDD.n2919 VDD.n2917 273.695
R11150 VDD.n3007 VDD.n2992 273.695
R11151 VDD.n3007 VDD.n3006 273.695
R11152 VDD.n3214 VDD.n3213 273.695
R11153 VDD.n3218 VDD.n3214 273.695
R11154 VDD.n3230 VDD.n3177 273.695
R11155 VDD.n3177 VDD.n3175 273.695
R11156 VDD.n3265 VDD.n3250 273.695
R11157 VDD.n3265 VDD.n3264 273.695
R11158 VDD.n3472 VDD.n3471 273.695
R11159 VDD.n3476 VDD.n3472 273.695
R11160 VDD.n3488 VDD.n3435 273.695
R11161 VDD.n3435 VDD.n3433 273.695
R11162 VDD.n3523 VDD.n3508 273.695
R11163 VDD.n3523 VDD.n3522 273.695
R11164 VDD.n5799 VDD.n5798 273.695
R11165 VDD.n5803 VDD.n5799 273.695
R11166 VDD.n5815 VDD.n5762 273.695
R11167 VDD.n5762 VDD.n5760 273.695
R11168 VDD.n5850 VDD.n5835 273.695
R11169 VDD.n5850 VDD.n5849 273.695
R11170 VDD.n5545 VDD.n5544 273.695
R11171 VDD.n5549 VDD.n5545 273.695
R11172 VDD.n5561 VDD.n5508 273.695
R11173 VDD.n5508 VDD.n5506 273.695
R11174 VDD.n5596 VDD.n5581 273.695
R11175 VDD.n5596 VDD.n5595 273.695
R11176 VDD.n3730 VDD.n3729 273.695
R11177 VDD.n3734 VDD.n3730 273.695
R11178 VDD.n3746 VDD.n3693 273.695
R11179 VDD.n3693 VDD.n3691 273.695
R11180 VDD.n3781 VDD.n3766 273.695
R11181 VDD.n3781 VDD.n3780 273.695
R11182 VDD.n3988 VDD.n3987 273.695
R11183 VDD.n3992 VDD.n3988 273.695
R11184 VDD.n4004 VDD.n3951 273.695
R11185 VDD.n3951 VDD.n3949 273.695
R11186 VDD.n4039 VDD.n4024 273.695
R11187 VDD.n4039 VDD.n4038 273.695
R11188 VDD.n4246 VDD.n4245 273.695
R11189 VDD.n4250 VDD.n4246 273.695
R11190 VDD.n4262 VDD.n4209 273.695
R11191 VDD.n4209 VDD.n4207 273.695
R11192 VDD.n4297 VDD.n4282 273.695
R11193 VDD.n4297 VDD.n4296 273.695
R11194 VDD.n4504 VDD.n4503 273.695
R11195 VDD.n4508 VDD.n4504 273.695
R11196 VDD.n4520 VDD.n4467 273.695
R11197 VDD.n4467 VDD.n4465 273.695
R11198 VDD.n4555 VDD.n4540 273.695
R11199 VDD.n4555 VDD.n4554 273.695
R11200 VDD.n4762 VDD.n4761 273.695
R11201 VDD.n4766 VDD.n4762 273.695
R11202 VDD.n4778 VDD.n4725 273.695
R11203 VDD.n4725 VDD.n4723 273.695
R11204 VDD.n4813 VDD.n4798 273.695
R11205 VDD.n4813 VDD.n4812 273.695
R11206 VDD.n5074 VDD.n5059 273.695
R11207 VDD.n5074 VDD.n5073 273.695
R11208 VDD.n5039 VDD.n4986 273.695
R11209 VDD.n4986 VDD.n4984 273.695
R11210 VDD.n5023 VDD.n5022 273.695
R11211 VDD.n5027 VDD.n5023 273.695
R11212 VDD.n5336 VDD.n5321 273.695
R11213 VDD.n5336 VDD.n5335 273.695
R11214 VDD.n5301 VDD.n5248 273.695
R11215 VDD.n5248 VDD.n5246 273.695
R11216 VDD.n5285 VDD.n5284 273.695
R11217 VDD.n5289 VDD.n5285 273.695
R11218 VDD.n1616 VDD.t1173 260.435
R11219 VDD.n1624 VDD.t1155 256.07
R11220 VDD.n1627 VDD.t1158 256.07
R11221 VDD.n1629 VDD.t1162 256.07
R11222 VDD.n1632 VDD.t1176 256.07
R11223 VDD.n1649 VDD.t1168 251.637
R11224 VDD.t696 VDD.t1247 246.023
R11225 VDD.t135 VDD.t1180 246.023
R11226 VDD VDD.t161 241.819
R11227 VDD VDD.t48 241.819
R11228 VDD.t1241 VDD 233.643
R11229 VDD.t1256 VDD 233.643
R11230 VDD.t702 VDD 233.643
R11231 VDD.t2 VDD 233.643
R11232 VDD.t791 VDD 233.643
R11233 VDD.t1166 VDD 233.643
R11234 VDD.t1314 VDD 233.643
R11235 VDD.t68 VDD 233.643
R11236 VDD.t1322 VDD 233.643
R11237 VDD.t1211 VDD 233.643
R11238 VDD.n1605 VDD.t1165 229.433
R11239 VDD.t815 VDD 227.321
R11240 VDD VDD.t803 227.321
R11241 VDD.t881 VDD 227.321
R11242 VDD.t436 VDD 227.321
R11243 VDD.t965 VDD 227.321
R11244 VDD VDD.t953 227.321
R11245 VDD.t1033 VDD 227.321
R11246 VDD.t1486 VDD 227.321
R11247 VDD.t1341 VDD 227.321
R11248 VDD VDD.t1457 227.321
R11249 VDD.t1407 VDD 227.321
R11250 VDD.t518 VDD 227.321
R11251 VDD.t1291 VDD 225.625
R11252 VDD.t64 VDD 225.625
R11253 VDD.t1073 VDD 225.625
R11254 VDD.n1909 VDD.n1908 213.083
R11255 VDD.n1910 VDD.n1909 213.083
R11256 VDD.n1867 VDD.n1852 213.083
R11257 VDD.n1867 VDD.n1866 213.083
R11258 VDD.n2188 VDD.n2173 213.083
R11259 VDD.n2188 VDD.n2187 213.083
R11260 VDD.n2230 VDD.n2229 213.083
R11261 VDD.n2231 VDD.n2230 213.083
R11262 VDD.n2446 VDD.n2431 213.083
R11263 VDD.n2446 VDD.n2445 213.083
R11264 VDD.n2488 VDD.n2487 213.083
R11265 VDD.n2489 VDD.n2488 213.083
R11266 VDD.n2704 VDD.n2689 213.083
R11267 VDD.n2704 VDD.n2703 213.083
R11268 VDD.n2746 VDD.n2745 213.083
R11269 VDD.n2747 VDD.n2746 213.083
R11270 VDD.n2962 VDD.n2947 213.083
R11271 VDD.n2962 VDD.n2961 213.083
R11272 VDD.n3004 VDD.n3003 213.083
R11273 VDD.n3005 VDD.n3004 213.083
R11274 VDD.n3220 VDD.n3205 213.083
R11275 VDD.n3220 VDD.n3219 213.083
R11276 VDD.n3262 VDD.n3261 213.083
R11277 VDD.n3263 VDD.n3262 213.083
R11278 VDD.n3478 VDD.n3463 213.083
R11279 VDD.n3478 VDD.n3477 213.083
R11280 VDD.n3520 VDD.n3519 213.083
R11281 VDD.n3521 VDD.n3520 213.083
R11282 VDD.n5805 VDD.n5790 213.083
R11283 VDD.n5805 VDD.n5804 213.083
R11284 VDD.n5847 VDD.n5846 213.083
R11285 VDD.n5848 VDD.n5847 213.083
R11286 VDD.n5551 VDD.n5536 213.083
R11287 VDD.n5551 VDD.n5550 213.083
R11288 VDD.n5593 VDD.n5592 213.083
R11289 VDD.n5594 VDD.n5593 213.083
R11290 VDD.n3736 VDD.n3721 213.083
R11291 VDD.n3736 VDD.n3735 213.083
R11292 VDD.n3778 VDD.n3777 213.083
R11293 VDD.n3779 VDD.n3778 213.083
R11294 VDD.n3994 VDD.n3979 213.083
R11295 VDD.n3994 VDD.n3993 213.083
R11296 VDD.n4036 VDD.n4035 213.083
R11297 VDD.n4037 VDD.n4036 213.083
R11298 VDD.n4252 VDD.n4237 213.083
R11299 VDD.n4252 VDD.n4251 213.083
R11300 VDD.n4294 VDD.n4293 213.083
R11301 VDD.n4295 VDD.n4294 213.083
R11302 VDD.n4510 VDD.n4495 213.083
R11303 VDD.n4510 VDD.n4509 213.083
R11304 VDD.n4552 VDD.n4551 213.083
R11305 VDD.n4553 VDD.n4552 213.083
R11306 VDD.n4768 VDD.n4753 213.083
R11307 VDD.n4768 VDD.n4767 213.083
R11308 VDD.n4810 VDD.n4809 213.083
R11309 VDD.n4811 VDD.n4810 213.083
R11310 VDD.n5071 VDD.n5070 213.083
R11311 VDD.n5072 VDD.n5071 213.083
R11312 VDD.n5029 VDD.n5014 213.083
R11313 VDD.n5029 VDD.n5028 213.083
R11314 VDD.n5333 VDD.n5332 213.083
R11315 VDD.n5334 VDD.n5333 213.083
R11316 VDD.n5291 VDD.n5276 213.083
R11317 VDD.n5291 VDD.n5290 213.083
R11318 VDD.n848 VDD.t814 204.903
R11319 VDD.n53 VDD.t964 204.903
R11320 VDD.n447 VDD.t1340 204.903
R11321 VDD.n1249 VDD.t322 204.9
R11322 VDD.n1634 VDD.t1509 201.587
R11323 VDD.n859 VDD.t816 201.012
R11324 VDD.n938 VDD.t804 201.012
R11325 VDD.n834 VDD.t882 201.012
R11326 VDD.n837 VDD.t437 201.012
R11327 VDD.n64 VDD.t966 201.012
R11328 VDD.n143 VDD.t954 201.012
R11329 VDD.n39 VDD.t1034 201.012
R11330 VDD.n42 VDD.t1487 201.012
R11331 VDD.n458 VDD.t1342 201.012
R11332 VDD.n537 VDD.t1458 201.012
R11333 VDD.n433 VDD.t1408 201.012
R11334 VDD.n436 VDD.t519 201.012
R11335 VDD.n1313 VDD.t228 201.012
R11336 VDD.n1342 VDD.t638 201.012
R11337 VDD.n1263 VDD.t210 201.012
R11338 VDD.n1260 VDD.t308 201.012
R11339 VDD.n1635 VDD.t1507 200.782
R11340 VDD.n1643 VDD.t1503 194.809
R11341 VDD.n1901 VDD.n1893 189.304
R11342 VDD.n2222 VDD.n2214 189.304
R11343 VDD.n2480 VDD.n2472 189.304
R11344 VDD.n2738 VDD.n2730 189.304
R11345 VDD.n2996 VDD.n2988 189.304
R11346 VDD.n3254 VDD.n3246 189.304
R11347 VDD.n3512 VDD.n3504 189.304
R11348 VDD.n5839 VDD.n5831 189.304
R11349 VDD.n5585 VDD.n5577 189.304
R11350 VDD.n3770 VDD.n3762 189.304
R11351 VDD.n4028 VDD.n4020 189.304
R11352 VDD.n4286 VDD.n4278 189.304
R11353 VDD.n4544 VDD.n4536 189.304
R11354 VDD.n4802 VDD.n4794 189.304
R11355 VDD.n5063 VDD.n5055 189.304
R11356 VDD.n5325 VDD.n5317 189.304
R11357 VDD.n1954 VDD.n1939 185
R11358 VDD.n1900 VDD.n1898 185
R11359 VDD.n1900 VDD.n1893 185
R11360 VDD.n1890 VDD.n1888 185
R11361 VDD.n1892 VDD.n1890 185
R11362 VDD.n1697 VDD.n1682 185
R11363 VDD.n2046 VDD.n2031 185
R11364 VDD.n2221 VDD.n2219 185
R11365 VDD.n2221 VDD.n2214 185
R11366 VDD.n2211 VDD.n2209 185
R11367 VDD.n2213 VDD.n2211 185
R11368 VDD.n2276 VDD.n2261 185
R11369 VDD.n2479 VDD.n2477 185
R11370 VDD.n2479 VDD.n2472 185
R11371 VDD.n2469 VDD.n2467 185
R11372 VDD.n2471 VDD.n2469 185
R11373 VDD.n2534 VDD.n2519 185
R11374 VDD.n2737 VDD.n2735 185
R11375 VDD.n2737 VDD.n2730 185
R11376 VDD.n2727 VDD.n2725 185
R11377 VDD.n2729 VDD.n2727 185
R11378 VDD.n2792 VDD.n2777 185
R11379 VDD.n2995 VDD.n2993 185
R11380 VDD.n2995 VDD.n2988 185
R11381 VDD.n2985 VDD.n2983 185
R11382 VDD.n2987 VDD.n2985 185
R11383 VDD.n3050 VDD.n3035 185
R11384 VDD.n3253 VDD.n3251 185
R11385 VDD.n3253 VDD.n3246 185
R11386 VDD.n3243 VDD.n3241 185
R11387 VDD.n3245 VDD.n3243 185
R11388 VDD.n3308 VDD.n3293 185
R11389 VDD.n3511 VDD.n3509 185
R11390 VDD.n3511 VDD.n3504 185
R11391 VDD.n3501 VDD.n3499 185
R11392 VDD.n3503 VDD.n3501 185
R11393 VDD.n5638 VDD.n5623 185
R11394 VDD.n5838 VDD.n5836 185
R11395 VDD.n5838 VDD.n5831 185
R11396 VDD.n5828 VDD.n5826 185
R11397 VDD.n5830 VDD.n5828 185
R11398 VDD.n5384 VDD.n5369 185
R11399 VDD.n5584 VDD.n5582 185
R11400 VDD.n5584 VDD.n5577 185
R11401 VDD.n5574 VDD.n5572 185
R11402 VDD.n5576 VDD.n5574 185
R11403 VDD.n3566 VDD.n3551 185
R11404 VDD.n3769 VDD.n3767 185
R11405 VDD.n3769 VDD.n3762 185
R11406 VDD.n3759 VDD.n3757 185
R11407 VDD.n3761 VDD.n3759 185
R11408 VDD.n3824 VDD.n3809 185
R11409 VDD.n4027 VDD.n4025 185
R11410 VDD.n4027 VDD.n4020 185
R11411 VDD.n4017 VDD.n4015 185
R11412 VDD.n4019 VDD.n4017 185
R11413 VDD.n4082 VDD.n4067 185
R11414 VDD.n4285 VDD.n4283 185
R11415 VDD.n4285 VDD.n4278 185
R11416 VDD.n4275 VDD.n4273 185
R11417 VDD.n4277 VDD.n4275 185
R11418 VDD.n4340 VDD.n4325 185
R11419 VDD.n4543 VDD.n4541 185
R11420 VDD.n4543 VDD.n4536 185
R11421 VDD.n4533 VDD.n4531 185
R11422 VDD.n4535 VDD.n4533 185
R11423 VDD.n4598 VDD.n4583 185
R11424 VDD.n4801 VDD.n4799 185
R11425 VDD.n4801 VDD.n4794 185
R11426 VDD.n4791 VDD.n4789 185
R11427 VDD.n4793 VDD.n4791 185
R11428 VDD.n4856 VDD.n4841 185
R11429 VDD.n5062 VDD.n5060 185
R11430 VDD.n5062 VDD.n5055 185
R11431 VDD.n5052 VDD.n5050 185
R11432 VDD.n5054 VDD.n5052 185
R11433 VDD.n5148 VDD.n5133 185
R11434 VDD.n5324 VDD.n5322 185
R11435 VDD.n5324 VDD.n5317 185
R11436 VDD.n5314 VDD.n5312 185
R11437 VDD.n5316 VDD.n5314 185
R11438 VDD.n1863 VDD.n1849 183.496
R11439 VDD.n2184 VDD.n2170 183.496
R11440 VDD.n2442 VDD.n2428 183.496
R11441 VDD.n2700 VDD.n2686 183.496
R11442 VDD.n2958 VDD.n2944 183.496
R11443 VDD.n3216 VDD.n3202 183.496
R11444 VDD.n3474 VDD.n3460 183.496
R11445 VDD.n5801 VDD.n5787 183.496
R11446 VDD.n5547 VDD.n5533 183.496
R11447 VDD.n3732 VDD.n3718 183.496
R11448 VDD.n3990 VDD.n3976 183.496
R11449 VDD.n4248 VDD.n4234 183.496
R11450 VDD.n4506 VDD.n4492 183.496
R11451 VDD.n4764 VDD.n4750 183.496
R11452 VDD.n5025 VDD.n5011 183.496
R11453 VDD.n5287 VDD.n5273 183.496
R11454 VDD.n1124 VDD.n1123 183.363
R11455 VDD.n1190 VDD.n1189 183.363
R11456 VDD.n1793 VDD.n1792 180.994
R11457 VDD.n1790 VDD.n1788 180.994
R11458 VDD.n2001 VDD.n2000 180.994
R11459 VDD.n1998 VDD.n1996 180.994
R11460 VDD.n2372 VDD.n2371 180.994
R11461 VDD.n2369 VDD.n2367 180.994
R11462 VDD.n2630 VDD.n2629 180.994
R11463 VDD.n2627 VDD.n2625 180.994
R11464 VDD.n2888 VDD.n2887 180.994
R11465 VDD.n2885 VDD.n2883 180.994
R11466 VDD.n3146 VDD.n3145 180.994
R11467 VDD.n3143 VDD.n3141 180.994
R11468 VDD.n3404 VDD.n3403 180.994
R11469 VDD.n3401 VDD.n3399 180.994
R11470 VDD.n5734 VDD.n5733 180.994
R11471 VDD.n5731 VDD.n5729 180.994
R11472 VDD.n5480 VDD.n5479 180.994
R11473 VDD.n5477 VDD.n5475 180.994
R11474 VDD.n3662 VDD.n3661 180.994
R11475 VDD.n3659 VDD.n3657 180.994
R11476 VDD.n3920 VDD.n3919 180.994
R11477 VDD.n3917 VDD.n3915 180.994
R11478 VDD.n4178 VDD.n4177 180.994
R11479 VDD.n4175 VDD.n4173 180.994
R11480 VDD.n4436 VDD.n4435 180.994
R11481 VDD.n4433 VDD.n4431 180.994
R11482 VDD.n4694 VDD.n4693 180.994
R11483 VDD.n4691 VDD.n4689 180.994
R11484 VDD.n4953 VDD.n4952 180.994
R11485 VDD.n4950 VDD.n4948 180.994
R11486 VDD.n5103 VDD.n5102 180.994
R11487 VDD.n5100 VDD.n5098 180.994
R11488 VDD.t735 VDD 179.821
R11489 VDD.t154 VDD 179.821
R11490 VDD.t50 VDD 179.821
R11491 VDD.t1255 VDD 179.821
R11492 VDD.n582 VDD.t663 179.821
R11493 VDD.t663 VDD 179.821
R11494 VDD.t47 VDD 179.821
R11495 VDD.n19 VDD.n5 179.131
R11496 VDD.n812 VDD.n811 179.131
R11497 VDD.n740 VDD.n739 179.131
R11498 VDD.n736 VDD.n735 179.131
R11499 VDD.n719 VDD.n718 179.131
R11500 VDD.n410 VDD.n409 179.131
R11501 VDD.n336 VDD.n322 179.131
R11502 VDD.n1581 VDD.n1580 179.131
R11503 VDD.n1577 VDD.n1576 179.131
R11504 VDD.n1560 VDD.n1559 179.131
R11505 VDD.t1224 VDD.n1803 174.632
R11506 VDD.t31 VDD.n2011 174.632
R11507 VDD.t538 VDD.n2382 174.632
R11508 VDD.t474 VDD.n2640 174.632
R11509 VDD.t1306 VDD.n2898 174.632
R11510 VDD.t8 VDD.n3156 174.632
R11511 VDD.t1196 VDD.n3414 174.632
R11512 VDD.t704 VDD.n5744 174.632
R11513 VDD.t1329 VDD.n5490 174.632
R11514 VDD.t1270 VDD.n3672 174.632
R11515 VDD.t78 VDD.n3930 174.632
R11516 VDD.t720 VDD.n4188 174.632
R11517 VDD.t1109 VDD.n4446 174.632
R11518 VDD.t185 VDD.n4704 174.632
R11519 VDD.t1123 VDD.n4963 174.632
R11520 VDD.t192 VDD.n5113 174.632
R11521 VDD.t1147 VDD 174.602
R11522 VDD.t672 VDD 174.602
R11523 VDD.n1010 VDD.n1009 174.595
R11524 VDD.n873 VDD.n872 174.595
R11525 VDD.n879 VDD.n878 174.595
R11526 VDD.n885 VDD.n884 174.595
R11527 VDD.n891 VDD.n890 174.595
R11528 VDD.n896 VDD.n895 174.595
R11529 VDD.n852 VDD.n851 174.595
R11530 VDD.n847 VDD.n846 174.595
R11531 VDD.n931 VDD.n930 174.595
R11532 VDD.n925 VDD.n924 174.595
R11533 VDD.n919 VDD.n918 174.595
R11534 VDD.n913 VDD.n912 174.595
R11535 VDD.n909 VDD.n908 174.595
R11536 VDD.n843 VDD.n842 174.595
R11537 VDD.n863 VDD.n862 174.595
R11538 VDD.n956 VDD.n955 174.595
R11539 VDD.n962 VDD.n961 174.595
R11540 VDD.n968 VDD.n967 174.595
R11541 VDD.n974 VDD.n973 174.595
R11542 VDD.n979 VDD.n978 174.595
R11543 VDD.n949 VDD.n948 174.595
R11544 VDD.n943 VDD.n942 174.595
R11545 VDD.n1066 VDD.n1065 174.595
R11546 VDD.n1072 VDD.n1071 174.595
R11547 VDD.n1078 VDD.n1077 174.595
R11548 VDD.n1084 VDD.n1083 174.595
R11549 VDD.n1088 VDD.n1087 174.595
R11550 VDD.n1095 VDD.n1094 174.595
R11551 VDD.n1103 VDD.n1102 174.595
R11552 VDD.n1019 VDD.n1018 174.595
R11553 VDD.n1025 VDD.n1024 174.595
R11554 VDD.n1031 VDD.n1030 174.595
R11555 VDD.n1037 VDD.n1036 174.595
R11556 VDD.n1041 VDD.n1040 174.595
R11557 VDD.n1047 VDD.n1046 174.595
R11558 VDD.n1055 VDD.n1054 174.595
R11559 VDD.n215 VDD.n214 174.595
R11560 VDD.n78 VDD.n77 174.595
R11561 VDD.n84 VDD.n83 174.595
R11562 VDD.n90 VDD.n89 174.595
R11563 VDD.n96 VDD.n95 174.595
R11564 VDD.n101 VDD.n100 174.595
R11565 VDD.n57 VDD.n56 174.595
R11566 VDD.n52 VDD.n51 174.595
R11567 VDD.n136 VDD.n135 174.595
R11568 VDD.n130 VDD.n129 174.595
R11569 VDD.n124 VDD.n123 174.595
R11570 VDD.n118 VDD.n117 174.595
R11571 VDD.n114 VDD.n113 174.595
R11572 VDD.n48 VDD.n47 174.595
R11573 VDD.n68 VDD.n67 174.595
R11574 VDD.n161 VDD.n160 174.595
R11575 VDD.n167 VDD.n166 174.595
R11576 VDD.n173 VDD.n172 174.595
R11577 VDD.n179 VDD.n178 174.595
R11578 VDD.n184 VDD.n183 174.595
R11579 VDD.n154 VDD.n153 174.595
R11580 VDD.n148 VDD.n147 174.595
R11581 VDD.n271 VDD.n270 174.595
R11582 VDD.n277 VDD.n276 174.595
R11583 VDD.n283 VDD.n282 174.595
R11584 VDD.n289 VDD.n288 174.595
R11585 VDD.n293 VDD.n292 174.595
R11586 VDD.n300 VDD.n299 174.595
R11587 VDD.n308 VDD.n307 174.595
R11588 VDD.n224 VDD.n223 174.595
R11589 VDD.n230 VDD.n229 174.595
R11590 VDD.n236 VDD.n235 174.595
R11591 VDD.n242 VDD.n241 174.595
R11592 VDD.n246 VDD.n245 174.595
R11593 VDD.n252 VDD.n251 174.595
R11594 VDD.n260 VDD.n259 174.595
R11595 VDD.n605 VDD.n604 174.595
R11596 VDD.n472 VDD.n471 174.595
R11597 VDD.n478 VDD.n477 174.595
R11598 VDD.n484 VDD.n483 174.595
R11599 VDD.n490 VDD.n489 174.595
R11600 VDD.n495 VDD.n494 174.595
R11601 VDD.n451 VDD.n450 174.595
R11602 VDD.n446 VDD.n445 174.595
R11603 VDD.n530 VDD.n529 174.595
R11604 VDD.n524 VDD.n523 174.595
R11605 VDD.n518 VDD.n517 174.595
R11606 VDD.n512 VDD.n511 174.595
R11607 VDD.n508 VDD.n507 174.595
R11608 VDD.n442 VDD.n441 174.595
R11609 VDD.n462 VDD.n461 174.595
R11610 VDD.n429 VDD.n428 174.595
R11611 VDD.n557 VDD.n556 174.595
R11612 VDD.n563 VDD.n562 174.595
R11613 VDD.n569 VDD.n568 174.595
R11614 VDD.n574 VDD.n573 174.595
R11615 VDD.n548 VDD.n547 174.595
R11616 VDD.n542 VDD.n541 174.595
R11617 VDD.n661 VDD.n660 174.595
R11618 VDD.n667 VDD.n666 174.595
R11619 VDD.n673 VDD.n672 174.595
R11620 VDD.n679 VDD.n678 174.595
R11621 VDD.n683 VDD.n682 174.595
R11622 VDD.n690 VDD.n689 174.595
R11623 VDD.n698 VDD.n697 174.595
R11624 VDD.n614 VDD.n613 174.595
R11625 VDD.n620 VDD.n619 174.595
R11626 VDD.n626 VDD.n625 174.595
R11627 VDD.n632 VDD.n631 174.595
R11628 VDD.n636 VDD.n635 174.595
R11629 VDD.n642 VDD.n641 174.595
R11630 VDD.n650 VDD.n649 174.595
R11631 VDD.n1353 VDD.n1352 174.595
R11632 VDD.n1335 VDD.n1334 174.595
R11633 VDD.n1329 VDD.n1328 174.595
R11634 VDD.n1322 VDD.n1321 174.595
R11635 VDD.n1435 VDD.n1434 174.595
R11636 VDD.n1439 VDD.n1438 174.595
R11637 VDD.n1445 VDD.n1444 174.595
R11638 VDD.n1451 VDD.n1450 174.595
R11639 VDD.n1379 VDD.n1378 174.595
R11640 VDD.n1385 VDD.n1384 174.595
R11641 VDD.n1391 VDD.n1390 174.595
R11642 VDD.n1403 VDD.n1402 174.595
R11643 VDD.n1408 VDD.n1407 174.595
R11644 VDD.n1414 VDD.n1413 174.595
R11645 VDD.n1420 VDD.n1419 174.595
R11646 VDD.n1306 VDD.n1305 174.595
R11647 VDD.n1299 VDD.n1298 174.595
R11648 VDD.n1293 VDD.n1292 174.595
R11649 VDD.n1268 VDD.n1267 174.595
R11650 VDD.n1272 VDD.n1271 174.595
R11651 VDD.n1278 VDD.n1277 174.595
R11652 VDD.n1265 VDD.n1264 174.595
R11653 VDD.n1465 VDD.n1464 174.595
R11654 VDD.n1471 VDD.n1470 174.595
R11655 VDD.n1477 VDD.n1476 174.595
R11656 VDD.n1483 VDD.n1482 174.595
R11657 VDD.n1487 VDD.n1486 174.595
R11658 VDD.n1493 VDD.n1492 174.595
R11659 VDD.n1499 VDD.n1498 174.595
R11660 VDD.n1515 VDD.n1514 174.595
R11661 VDD.n1521 VDD.n1520 174.595
R11662 VDD.n1257 VDD.n1256 174.595
R11663 VDD.n1531 VDD.n1530 174.595
R11664 VDD.n1535 VDD.n1534 174.595
R11665 VDD.n1253 VDD.n1252 174.595
R11666 VDD.n1248 VDD.n1247 174.595
R11667 VDD VDD.t209 174.385
R11668 VDD VDD.t227 174.385
R11669 VDD VDD.t399 173.083
R11670 VDD.n987 VDD.t735 173.036
R11671 VDD.n192 VDD.t50 173.036
R11672 VDD.n1822 VDD.n1820 170.542
R11673 VDD.n2143 VDD.n2141 170.542
R11674 VDD.n2401 VDD.n2399 170.542
R11675 VDD.n2659 VDD.n2657 170.542
R11676 VDD.n2917 VDD.n2915 170.542
R11677 VDD.n3175 VDD.n3173 170.542
R11678 VDD.n3433 VDD.n3431 170.542
R11679 VDD.n5760 VDD.n5758 170.542
R11680 VDD.n5506 VDD.n5504 170.542
R11681 VDD.n3691 VDD.n3689 170.542
R11682 VDD.n3949 VDD.n3947 170.542
R11683 VDD.n4207 VDD.n4205 170.542
R11684 VDD.n4465 VDD.n4463 170.542
R11685 VDD.n4723 VDD.n4721 170.542
R11686 VDD.n4984 VDD.n4982 170.542
R11687 VDD.n5246 VDD.n5244 170.542
R11688 VDD.t653 VDD 170.478
R11689 VDD.t56 VDD 170.478
R11690 VDD VDD.n1428 169.179
R11691 VDD.n32 VDD.n31 169.107
R11692 VDD.n826 VDD.n825 169.107
R11693 VDD.n753 VDD.n752 169.107
R11694 VDD.n722 VDD.n721 169.107
R11695 VDD.n424 VDD.n423 169.107
R11696 VDD.n349 VDD.n348 169.107
R11697 VDD.n1594 VDD.n1593 169.107
R11698 VDD.n1563 VDD.n1562 169.107
R11699 VDD.n1136 VDD.n1117 169.107
R11700 VDD.n1129 VDD.n1120 169.107
R11701 VDD.n1202 VDD.n1183 169.107
R11702 VDD.n1195 VDD.n1186 169.107
R11703 VDD.n990 VDD.n989 169.017
R11704 VDD.n195 VDD.n194 169.017
R11705 VDD.n585 VDD.n584 169.017
R11706 VDD.n1645 VDD.t1152 168.561
R11707 VDD.n1689 VDD.n1673 167.234
R11708 VDD.n2038 VDD.n2022 167.234
R11709 VDD.n2268 VDD.n2252 167.234
R11710 VDD.n2526 VDD.n2510 167.234
R11711 VDD.n2784 VDD.n2768 167.234
R11712 VDD.n3042 VDD.n3026 167.234
R11713 VDD.n3300 VDD.n3284 167.234
R11714 VDD.n5630 VDD.n5614 167.234
R11715 VDD.n5376 VDD.n5360 167.234
R11716 VDD.n3558 VDD.n3542 167.234
R11717 VDD.n3816 VDD.n3800 167.234
R11718 VDD.n4074 VDD.n4058 167.234
R11719 VDD.n4332 VDD.n4316 167.234
R11720 VDD.n4590 VDD.n4574 167.234
R11721 VDD.n4848 VDD.n4832 167.234
R11722 VDD.n5140 VDD.n5124 167.234
R11723 VDD.n1746 VDD.n1715 166.812
R11724 VDD.n2095 VDD.n2064 166.812
R11725 VDD.n2325 VDD.n2294 166.812
R11726 VDD.n2583 VDD.n2552 166.812
R11727 VDD.n2841 VDD.n2810 166.812
R11728 VDD.n3099 VDD.n3068 166.812
R11729 VDD.n3357 VDD.n3326 166.812
R11730 VDD.n5687 VDD.n5656 166.812
R11731 VDD.n5433 VDD.n5402 166.812
R11732 VDD.n3615 VDD.n3584 166.812
R11733 VDD.n3873 VDD.n3842 166.812
R11734 VDD.n4131 VDD.n4100 166.812
R11735 VDD.n4389 VDD.n4358 166.812
R11736 VDD.n4647 VDD.n4616 166.812
R11737 VDD.n4905 VDD.n4874 166.812
R11738 VDD.n5197 VDD.n5166 166.812
R11739 VDD.n1645 VDD.t1511 166.328
R11740 VDD.n1834 VDD.n1830 165.767
R11741 VDD.n1814 VDD.n1813 165.767
R11742 VDD.n2135 VDD.n2134 165.767
R11743 VDD.n2155 VDD.n2151 165.767
R11744 VDD.n2393 VDD.n2392 165.767
R11745 VDD.n2413 VDD.n2409 165.767
R11746 VDD.n2651 VDD.n2650 165.767
R11747 VDD.n2671 VDD.n2667 165.767
R11748 VDD.n2909 VDD.n2908 165.767
R11749 VDD.n2929 VDD.n2925 165.767
R11750 VDD.n3167 VDD.n3166 165.767
R11751 VDD.n3187 VDD.n3183 165.767
R11752 VDD.n3425 VDD.n3424 165.767
R11753 VDD.n3445 VDD.n3441 165.767
R11754 VDD.n5752 VDD.n5751 165.767
R11755 VDD.n5772 VDD.n5768 165.767
R11756 VDD.n5498 VDD.n5497 165.767
R11757 VDD.n5518 VDD.n5514 165.767
R11758 VDD.n3683 VDD.n3682 165.767
R11759 VDD.n3703 VDD.n3699 165.767
R11760 VDD.n3941 VDD.n3940 165.767
R11761 VDD.n3961 VDD.n3957 165.767
R11762 VDD.n4199 VDD.n4198 165.767
R11763 VDD.n4219 VDD.n4215 165.767
R11764 VDD.n4457 VDD.n4456 165.767
R11765 VDD.n4477 VDD.n4473 165.767
R11766 VDD.n4715 VDD.n4714 165.767
R11767 VDD.n4735 VDD.n4731 165.767
R11768 VDD.n4996 VDD.n4992 165.767
R11769 VDD.n4976 VDD.n4975 165.767
R11770 VDD.n5258 VDD.n5254 165.767
R11771 VDD.n5238 VDD.n5237 165.767
R11772 VDD.t1134 VDD.t546 164.554
R11773 VDD.t1057 VDD.t391 164.554
R11774 VDD.t1304 VDD.t152 164.554
R11775 VDD.n24 VDD.n1 164.215
R11776 VDD.n805 VDD.n785 164.215
R11777 VDD.n757 VDD.n756 164.215
R11778 VDD.n777 VDD.n776 164.215
R11779 VDD.n403 VDD.n383 164.215
R11780 VDD.n354 VDD.n353 164.215
R11781 VDD.n374 VDD.n373 164.215
R11782 VDD.n341 VDD.n318 164.215
R11783 VDD.n1699 VDD.n1682 161.506
R11784 VDD.n2048 VDD.n2031 161.506
R11785 VDD.n2278 VDD.n2261 161.506
R11786 VDD.n2536 VDD.n2519 161.506
R11787 VDD.n2794 VDD.n2777 161.506
R11788 VDD.n3052 VDD.n3035 161.506
R11789 VDD.n3310 VDD.n3293 161.506
R11790 VDD.n5640 VDD.n5623 161.506
R11791 VDD.n5386 VDD.n5369 161.506
R11792 VDD.n3568 VDD.n3551 161.506
R11793 VDD.n3826 VDD.n3809 161.506
R11794 VDD.n4084 VDD.n4067 161.506
R11795 VDD.n4342 VDD.n4325 161.506
R11796 VDD.n4600 VDD.n4583 161.506
R11797 VDD.n4858 VDD.n4841 161.506
R11798 VDD.n5150 VDD.n5133 161.506
R11799 VDD.n1741 VDD.n1728 159.143
R11800 VDD.n2090 VDD.n2077 159.143
R11801 VDD.n2320 VDD.n2307 159.143
R11802 VDD.n2578 VDD.n2565 159.143
R11803 VDD.n2836 VDD.n2823 159.143
R11804 VDD.n3094 VDD.n3081 159.143
R11805 VDD.n3352 VDD.n3339 159.143
R11806 VDD.n5682 VDD.n5669 159.143
R11807 VDD.n5428 VDD.n5415 159.143
R11808 VDD.n3610 VDD.n3597 159.143
R11809 VDD.n3868 VDD.n3855 159.143
R11810 VDD.n4126 VDD.n4113 159.143
R11811 VDD.n4384 VDD.n4371 159.143
R11812 VDD.n4642 VDD.n4629 159.143
R11813 VDD.n4900 VDD.n4887 159.143
R11814 VDD.n5192 VDD.n5179 159.143
R11815 VDD.n1905 VDD.n1892 159.108
R11816 VDD.n1858 VDD.n1857 159.108
R11817 VDD.n2179 VDD.n2178 159.108
R11818 VDD.n2226 VDD.n2213 159.108
R11819 VDD.n2437 VDD.n2436 159.108
R11820 VDD.n2484 VDD.n2471 159.108
R11821 VDD.n2695 VDD.n2694 159.108
R11822 VDD.n2742 VDD.n2729 159.108
R11823 VDD.n2953 VDD.n2952 159.108
R11824 VDD.n3000 VDD.n2987 159.108
R11825 VDD.n3211 VDD.n3210 159.108
R11826 VDD.n3258 VDD.n3245 159.108
R11827 VDD.n3469 VDD.n3468 159.108
R11828 VDD.n3516 VDD.n3503 159.108
R11829 VDD.n5796 VDD.n5795 159.108
R11830 VDD.n5843 VDD.n5830 159.108
R11831 VDD.n5542 VDD.n5541 159.108
R11832 VDD.n5589 VDD.n5576 159.108
R11833 VDD.n3727 VDD.n3726 159.108
R11834 VDD.n3774 VDD.n3761 159.108
R11835 VDD.n3985 VDD.n3984 159.108
R11836 VDD.n4032 VDD.n4019 159.108
R11837 VDD.n4243 VDD.n4242 159.108
R11838 VDD.n4290 VDD.n4277 159.108
R11839 VDD.n4501 VDD.n4500 159.108
R11840 VDD.n4548 VDD.n4535 159.108
R11841 VDD.n4759 VDD.n4758 159.108
R11842 VDD.n4806 VDD.n4793 159.108
R11843 VDD.n5067 VDD.n5054 159.108
R11844 VDD.n5020 VDD.n5019 159.108
R11845 VDD.n5329 VDD.n5316 159.108
R11846 VDD.n5282 VDD.n5281 159.108
R11847 VDD.n1605 VDD.t1505 158.886
R11848 VDD.n1700 VDD.n1699 158.776
R11849 VDD.n2049 VDD.n2048 158.776
R11850 VDD.n2279 VDD.n2278 158.776
R11851 VDD.n2537 VDD.n2536 158.776
R11852 VDD.n2795 VDD.n2794 158.776
R11853 VDD.n3053 VDD.n3052 158.776
R11854 VDD.n3311 VDD.n3310 158.776
R11855 VDD.n5641 VDD.n5640 158.776
R11856 VDD.n5387 VDD.n5386 158.776
R11857 VDD.n3569 VDD.n3568 158.776
R11858 VDD.n3827 VDD.n3826 158.776
R11859 VDD.n4085 VDD.n4084 158.776
R11860 VDD.n4343 VDD.n4342 158.776
R11861 VDD.n4601 VDD.n4600 158.776
R11862 VDD.n4859 VDD.n4858 158.776
R11863 VDD.n5151 VDD.n5150 158.776
R11864 VDD.n858 VDD.t896 158.117
R11865 VDD.n937 VDD.t880 158.117
R11866 VDD.n833 VDD.t860 158.117
R11867 VDD.n836 VDD.t822 158.117
R11868 VDD.n839 VDD.t427 158.117
R11869 VDD.n63 VDD.t1046 158.117
R11870 VDD.n142 VDD.t1032 158.117
R11871 VDD.n38 VDD.t1010 158.117
R11872 VDD.n41 VDD.t972 158.117
R11873 VDD.n44 VDD.t1477 158.117
R11874 VDD.n457 VDD.t1422 158.117
R11875 VDD.n536 VDD.t1406 158.117
R11876 VDD.n432 VDD.t1386 158.117
R11877 VDD.n435 VDD.t1348 158.117
R11878 VDD.n438 VDD.t509 158.117
R11879 VDD.n1341 VDD.t326 158.117
R11880 VDD.n1347 VDD.t616 158.117
R11881 VDD.n1312 VDD.t302 158.117
R11882 VDD.n1262 VDD.t304 158.117
R11883 VDD.n1259 VDD.t252 158.117
R11884 VDD.n988 VDD.t736 158.06
R11885 VDD.n193 VDD.t51 158.06
R11886 VDD.n583 VDD.t664 158.06
R11887 VDD.n1362 VDD.t394 158.06
R11888 VDD.n1143 VDD.t792 158.06
R11889 VDD.n1142 VDD.t3 158.06
R11890 VDD.n1141 VDD.t703 158.06
R11891 VDD.n1140 VDD.t1257 158.06
R11892 VDD.n1139 VDD.t1242 158.06
R11893 VDD.n1542 VDD.t652 158.06
R11894 VDD.n1209 VDD.t1212 158.06
R11895 VDD.n1208 VDD.t1323 158.06
R11896 VDD.n1207 VDD.t69 158.06
R11897 VDD.n1206 VDD.t1315 158.06
R11898 VDD.n1205 VDD.t1167 158.06
R11899 VDD.n1616 VDD.t1508 156.403
R11900 VDD.t161 VDD.t1276 155.456
R11901 VDD.t48 VDD.t1132 155.456
R11902 VDD.n1679 VDD.n1670 155.294
R11903 VDD.n2028 VDD.n2019 155.294
R11904 VDD.n2258 VDD.n2249 155.294
R11905 VDD.n2516 VDD.n2507 155.294
R11906 VDD.n2774 VDD.n2765 155.294
R11907 VDD.n3032 VDD.n3023 155.294
R11908 VDD.n3290 VDD.n3281 155.294
R11909 VDD.n5620 VDD.n5611 155.294
R11910 VDD.n5366 VDD.n5357 155.294
R11911 VDD.n3548 VDD.n3539 155.294
R11912 VDD.n3806 VDD.n3797 155.294
R11913 VDD.n4064 VDD.n4055 155.294
R11914 VDD.n4322 VDD.n4313 155.294
R11915 VDD.n4580 VDD.n4571 155.294
R11916 VDD.n4838 VDD.n4829 155.294
R11917 VDD.n5130 VDD.n5121 155.294
R11918 VDD.n1507 VDD.t307 153.562
R11919 VDD VDD.t1206 151.137
R11920 VDD VDD.t661 151.137
R11921 VDD.n1784 VDD.t42 151.123
R11922 VDD.n1786 VDD.t1225 151.123
R11923 VDD.n1992 VDD.t363 151.123
R11924 VDD.n1994 VDD.t34 151.123
R11925 VDD.n2363 VDD.t465 151.123
R11926 VDD.n2365 VDD.t543 151.123
R11927 VDD.n2621 VDD.t120 151.123
R11928 VDD.n2623 VDD.t475 151.123
R11929 VDD.n2879 VDD.t20 151.123
R11930 VDD.n2881 VDD.t1307 151.123
R11931 VDD.n3137 VDD.t589 151.123
R11932 VDD.n3139 VDD.t12 151.123
R11933 VDD.n3395 VDD.t549 151.123
R11934 VDD.n3397 VDD.t1197 151.123
R11935 VDD.n5725 VDD.t169 151.123
R11936 VDD.n5727 VDD.t705 151.123
R11937 VDD.n5471 VDD.t762 151.123
R11938 VDD.n5473 VDD.t1333 151.123
R11939 VDD.n3653 VDD.t1099 151.123
R11940 VDD.n3655 VDD.t1271 151.123
R11941 VDD.n3911 VDD.t789 151.123
R11942 VDD.n3913 VDD.t83 151.123
R11943 VDD.n4169 VDD.t495 151.123
R11944 VDD.n4171 VDD.t725 151.123
R11945 VDD.n4427 VDD.t373 151.123
R11946 VDD.n4429 VDD.t1110 151.123
R11947 VDD.n4685 VDD.t110 151.123
R11948 VDD.n4687 VDD.t189 151.123
R11949 VDD.n4944 VDD.t348 151.123
R11950 VDD.n4946 VDD.t1124 151.123
R11951 VDD.n5094 VDD.t481 151.123
R11952 VDD.n5096 VDD.t193 151.123
R11953 VDD.n841 VDD.t1290 151.123
R11954 VDD.n46 VDD.t63 151.123
R11955 VDD.n440 VDD.t1080 151.123
R11956 VDD.n1357 VDD.t402 151.123
R11957 VDD.n1624 VDD.t1506 150.03
R11958 VDD.n1627 VDD.t1502 150.03
R11959 VDD.n1629 VDD.t1504 150.03
R11960 VDD.n1632 VDD.t1510 150.03
R11961 VDD.t1243 VDD.t645 148.481
R11962 VDD.t1174 VDD.t27 148.481
R11963 VDD.n1802 VDD.t39 146.691
R11964 VDD.n2010 VDD.t362 146.691
R11965 VDD.n2381 VDD.t464 146.691
R11966 VDD.n2639 VDD.t119 146.691
R11967 VDD.n2897 VDD.t19 146.691
R11968 VDD.n3155 VDD.t588 146.691
R11969 VDD.n3413 VDD.t548 146.691
R11970 VDD.n5743 VDD.t168 146.691
R11971 VDD.n5489 VDD.t759 146.691
R11972 VDD.n3671 VDD.t1097 146.691
R11973 VDD.n3929 VDD.t783 146.691
R11974 VDD.n4187 VDD.t492 146.691
R11975 VDD.n4445 VDD.t372 146.691
R11976 VDD.n4703 VDD.t109 146.691
R11977 VDD.n4962 VDD.t347 146.691
R11978 VDD.n5112 VDD.t480 146.691
R11979 VDD.t1282 VDD.t17 145.243
R11980 VDD.t1326 VDD.t1324 145.243
R11981 VDD.n1647 VDD.t1512 145.043
R11982 VDD.n1741 VDD.n1740 143.435
R11983 VDD.n2090 VDD.n2089 143.435
R11984 VDD.n2320 VDD.n2319 143.435
R11985 VDD.n2578 VDD.n2577 143.435
R11986 VDD.n2836 VDD.n2835 143.435
R11987 VDD.n3094 VDD.n3093 143.435
R11988 VDD.n3352 VDD.n3351 143.435
R11989 VDD.n5682 VDD.n5681 143.435
R11990 VDD.n5428 VDD.n5427 143.435
R11991 VDD.n3610 VDD.n3609 143.435
R11992 VDD.n3868 VDD.n3867 143.435
R11993 VDD.n4126 VDD.n4125 143.435
R11994 VDD.n4384 VDD.n4383 143.435
R11995 VDD.n4642 VDD.n4641 143.435
R11996 VDD.n4900 VDD.n4899 143.435
R11997 VDD.n5192 VDD.n5191 143.435
R11998 VDD.t745 VDD.t0 143.232
R11999 VDD.t389 VDD.t1222 143.232
R12000 VDD.t839 VDD.t813 142.5
R12001 VDD.t925 VDD.t839 142.5
R12002 VDD.t817 VDD.t925 142.5
R12003 VDD.t809 VDD.t817 142.5
R12004 VDD.t831 VDD.t809 142.5
R12005 VDD.t799 VDD.t857 142.5
R12006 VDD.t835 VDD.t799 142.5
R12007 VDD.t905 VDD.t835 142.5
R12008 VDD.t801 VDD.t905 142.5
R12009 VDD.t825 VDD.t801 142.5
R12010 VDD.t889 VDD.t825 142.5
R12011 VDD.t919 VDD.t889 142.5
R12012 VDD.t851 VDD.t919 142.5
R12013 VDD.t895 VDD.t851 142.5
R12014 VDD.t883 VDD.t815 142.5
R12015 VDD.t909 VDD.t883 142.5
R12016 VDD.t807 VDD.t909 142.5
R12017 VDD.t863 VDD.t807 142.5
R12018 VDD.t897 VDD.t829 142.5
R12019 VDD.t829 VDD.t867 142.5
R12020 VDD.t867 VDD.t901 142.5
R12021 VDD.t901 VDD.t837 142.5
R12022 VDD.t837 VDD.t917 142.5
R12023 VDD.t917 VDD.t849 142.5
R12024 VDD.t849 VDD.t875 142.5
R12025 VDD.t875 VDD.t923 142.5
R12026 VDD.t923 VDD.t855 142.5
R12027 VDD.t855 VDD.t879 142.5
R12028 VDD.t803 VDD.t861 142.5
R12029 VDD.t861 VDD.t891 142.5
R12030 VDD.t891 VDD.t827 142.5
R12031 VDD.t827 VDD.t913 142.5
R12032 VDD.t913 VDD.t823 142.5
R12033 VDD.t915 VDD.t887 142.5
R12034 VDD.t845 VDD.t915 142.5
R12035 VDD.t871 VDD.t845 142.5
R12036 VDD.t903 VDD.t871 142.5
R12037 VDD.t847 VDD.t903 142.5
R12038 VDD.t873 VDD.t847 142.5
R12039 VDD.t819 VDD.t873 142.5
R12040 VDD.t841 VDD.t819 142.5
R12041 VDD.t859 VDD.t841 142.5
R12042 VDD.t907 VDD.t881 142.5
R12043 VDD.t805 VDD.t907 142.5
R12044 VDD.t885 VDD.t805 142.5
R12045 VDD.t843 VDD.t911 142.5
R12046 VDD.t865 VDD.t843 142.5
R12047 VDD.t899 VDD.t865 142.5
R12048 VDD.t833 VDD.t899 142.5
R12049 VDD.t869 VDD.t833 142.5
R12050 VDD.t811 VDD.t869 142.5
R12051 VDD.t893 VDD.t811 142.5
R12052 VDD.t921 VDD.t893 142.5
R12053 VDD.t853 VDD.t921 142.5
R12054 VDD.t877 VDD.t853 142.5
R12055 VDD.t821 VDD.t877 142.5
R12056 VDD.t450 VDD.t436 142.5
R12057 VDD.t438 VDD.t430 142.5
R12058 VDD.t448 VDD.t438 142.5
R12059 VDD.t444 VDD.t448 142.5
R12060 VDD.t452 VDD.t444 142.5
R12061 VDD.t432 VDD.t452 142.5
R12062 VDD.t446 VDD.t432 142.5
R12063 VDD.t454 VDD.t446 142.5
R12064 VDD.t434 VDD.t454 142.5
R12065 VDD.t440 VDD.t434 142.5
R12066 VDD.t424 VDD.t440 142.5
R12067 VDD.t428 VDD.t424 142.5
R12068 VDD.t442 VDD.t428 142.5
R12069 VDD.t426 VDD.t442 142.5
R12070 VDD.t1293 VDD.t1291 142.5
R12071 VDD.t1295 VDD.t1293 142.5
R12072 VDD.t1289 VDD.t1295 142.5
R12073 VDD.t989 VDD.t963 142.5
R12074 VDD.t947 VDD.t989 142.5
R12075 VDD.t967 VDD.t947 142.5
R12076 VDD.t959 VDD.t967 142.5
R12077 VDD.t979 VDD.t959 142.5
R12078 VDD.t949 VDD.t1007 142.5
R12079 VDD.t985 VDD.t949 142.5
R12080 VDD.t927 VDD.t985 142.5
R12081 VDD.t951 VDD.t927 142.5
R12082 VDD.t975 VDD.t951 142.5
R12083 VDD.t1039 VDD.t975 142.5
R12084 VDD.t941 VDD.t1039 142.5
R12085 VDD.t1001 VDD.t941 142.5
R12086 VDD.t1045 VDD.t1001 142.5
R12087 VDD.t1015 VDD.t965 142.5
R12088 VDD.t931 VDD.t1015 142.5
R12089 VDD.t957 VDD.t931 142.5
R12090 VDD.t1013 VDD.t957 142.5
R12091 VDD.t1047 VDD.t981 142.5
R12092 VDD.t981 VDD.t1019 142.5
R12093 VDD.t1019 VDD.t1051 142.5
R12094 VDD.t1051 VDD.t987 142.5
R12095 VDD.t987 VDD.t939 142.5
R12096 VDD.t939 VDD.t999 142.5
R12097 VDD.t999 VDD.t1027 142.5
R12098 VDD.t1027 VDD.t945 142.5
R12099 VDD.t945 VDD.t1005 142.5
R12100 VDD.t1005 VDD.t1031 142.5
R12101 VDD.t953 VDD.t1011 142.5
R12102 VDD.t1011 VDD.t1041 142.5
R12103 VDD.t1041 VDD.t977 142.5
R12104 VDD.t977 VDD.t935 142.5
R12105 VDD.t935 VDD.t973 142.5
R12106 VDD.t937 VDD.t1037 142.5
R12107 VDD.t995 VDD.t937 142.5
R12108 VDD.t1023 VDD.t995 142.5
R12109 VDD.t1053 VDD.t1023 142.5
R12110 VDD.t997 VDD.t1053 142.5
R12111 VDD.t1025 VDD.t997 142.5
R12112 VDD.t969 VDD.t1025 142.5
R12113 VDD.t991 VDD.t969 142.5
R12114 VDD.t1009 VDD.t991 142.5
R12115 VDD.t929 VDD.t1033 142.5
R12116 VDD.t955 VDD.t929 142.5
R12117 VDD.t1035 VDD.t955 142.5
R12118 VDD.t993 VDD.t933 142.5
R12119 VDD.t1017 VDD.t993 142.5
R12120 VDD.t1049 VDD.t1017 142.5
R12121 VDD.t983 VDD.t1049 142.5
R12122 VDD.t1021 VDD.t983 142.5
R12123 VDD.t961 VDD.t1021 142.5
R12124 VDD.t1043 VDD.t961 142.5
R12125 VDD.t943 VDD.t1043 142.5
R12126 VDD.t1003 VDD.t943 142.5
R12127 VDD.t1029 VDD.t1003 142.5
R12128 VDD.t971 VDD.t1029 142.5
R12129 VDD.t1468 VDD.t1486 142.5
R12130 VDD.t1488 VDD.t1480 142.5
R12131 VDD.t1498 VDD.t1488 142.5
R12132 VDD.t1494 VDD.t1498 142.5
R12133 VDD.t1470 VDD.t1494 142.5
R12134 VDD.t1482 VDD.t1470 142.5
R12135 VDD.t1496 VDD.t1482 142.5
R12136 VDD.t1472 VDD.t1496 142.5
R12137 VDD.t1484 VDD.t1472 142.5
R12138 VDD.t1490 VDD.t1484 142.5
R12139 VDD.t1474 VDD.t1490 142.5
R12140 VDD.t1478 VDD.t1474 142.5
R12141 VDD.t1492 VDD.t1478 142.5
R12142 VDD.t1476 VDD.t1492 142.5
R12143 VDD.t66 VDD.t64 142.5
R12144 VDD.t60 VDD.t66 142.5
R12145 VDD.t62 VDD.t60 142.5
R12146 VDD.t1365 VDD.t1339 142.5
R12147 VDD.t1451 VDD.t1365 142.5
R12148 VDD.t1343 VDD.t1451 142.5
R12149 VDD.t1463 VDD.t1343 142.5
R12150 VDD.t1355 VDD.t1463 142.5
R12151 VDD.t1453 VDD.t1383 142.5
R12152 VDD.t1363 VDD.t1453 142.5
R12153 VDD.t1431 VDD.t1363 142.5
R12154 VDD.t1455 VDD.t1431 142.5
R12155 VDD.t1351 VDD.t1455 142.5
R12156 VDD.t1415 VDD.t1351 142.5
R12157 VDD.t1445 VDD.t1415 142.5
R12158 VDD.t1377 VDD.t1445 142.5
R12159 VDD.t1421 VDD.t1377 142.5
R12160 VDD.t1409 VDD.t1341 142.5
R12161 VDD.t1435 VDD.t1409 142.5
R12162 VDD.t1461 VDD.t1435 142.5
R12163 VDD.t1389 VDD.t1461 142.5
R12164 VDD.t1423 VDD.t1357 142.5
R12165 VDD.t1357 VDD.t1393 142.5
R12166 VDD.t1393 VDD.t1427 142.5
R12167 VDD.t1427 VDD.t1361 142.5
R12168 VDD.t1361 VDD.t1443 142.5
R12169 VDD.t1443 VDD.t1375 142.5
R12170 VDD.t1375 VDD.t1401 142.5
R12171 VDD.t1401 VDD.t1449 142.5
R12172 VDD.t1449 VDD.t1381 142.5
R12173 VDD.t1381 VDD.t1405 142.5
R12174 VDD.t1457 VDD.t1387 142.5
R12175 VDD.t1387 VDD.t1417 142.5
R12176 VDD.t1417 VDD.t1353 142.5
R12177 VDD.t1353 VDD.t1439 142.5
R12178 VDD.t1439 VDD.t1349 142.5
R12179 VDD.t1441 VDD.t1413 142.5
R12180 VDD.t1371 VDD.t1441 142.5
R12181 VDD.t1397 VDD.t1371 142.5
R12182 VDD.t1429 VDD.t1397 142.5
R12183 VDD.t1373 VDD.t1429 142.5
R12184 VDD.t1399 VDD.t1373 142.5
R12185 VDD.t1345 VDD.t1399 142.5
R12186 VDD.t1367 VDD.t1345 142.5
R12187 VDD.t1385 VDD.t1367 142.5
R12188 VDD.t1433 VDD.t1407 142.5
R12189 VDD.t1459 VDD.t1433 142.5
R12190 VDD.t1411 VDD.t1459 142.5
R12191 VDD.t1369 VDD.t1437 142.5
R12192 VDD.t1391 VDD.t1369 142.5
R12193 VDD.t1425 VDD.t1391 142.5
R12194 VDD.t1359 VDD.t1425 142.5
R12195 VDD.t1395 VDD.t1359 142.5
R12196 VDD.t1337 VDD.t1395 142.5
R12197 VDD.t1419 VDD.t1337 142.5
R12198 VDD.t1447 VDD.t1419 142.5
R12199 VDD.t1379 VDD.t1447 142.5
R12200 VDD.t1403 VDD.t1379 142.5
R12201 VDD.t1347 VDD.t1403 142.5
R12202 VDD.t532 VDD.t518 142.5
R12203 VDD.t520 VDD.t512 142.5
R12204 VDD.t530 VDD.t520 142.5
R12205 VDD.t526 VDD.t530 142.5
R12206 VDD.t534 VDD.t526 142.5
R12207 VDD.t514 VDD.t534 142.5
R12208 VDD.t528 VDD.t514 142.5
R12209 VDD.t536 VDD.t528 142.5
R12210 VDD.t516 VDD.t536 142.5
R12211 VDD.t522 VDD.t516 142.5
R12212 VDD.t506 VDD.t522 142.5
R12213 VDD.t510 VDD.t506 142.5
R12214 VDD.t524 VDD.t510 142.5
R12215 VDD.t508 VDD.t524 142.5
R12216 VDD.t1075 VDD.t1073 142.5
R12217 VDD.t1077 VDD.t1075 142.5
R12218 VDD.t1079 VDD.t1077 142.5
R12219 VDD.t17 VDD.t1467 142.279
R12220 VDD.t1281 VDD.t200 142.279
R12221 VDD.t1324 VDD.t409 142.279
R12222 VDD.t167 VDD.t798 142.279
R12223 VDD.t1107 VDD.t1465 141.061
R12224 VDD.t729 VDD.t407 141.061
R12225 VDD.n986 VDD.t450 139.107
R12226 VDD.n191 VDD.t1468 139.107
R12227 VDD.t1437 VDD.n580 139.107
R12228 VDD VDD.t89 138.857
R12229 VDD VDD.t649 138.857
R12230 VDD.t1465 VDD.t695 138.183
R12231 VDD.t86 VDD.t359 138.183
R12232 VDD.t407 VDD.t1059 138.183
R12233 VDD.t456 VDD.t728 138.183
R12234 VDD.t393 VDD 137.946
R12235 VDD.t417 VDD.n1821 136.591
R12236 VDD.t1085 VDD.n2142 136.591
R12237 VDD.t567 VDD.n2400 136.591
R12238 VDD.t387 VDD.n2658 136.591
R12239 VDD.t560 VDD.n2916 136.591
R12240 VDD.t573 VDD.n3174 136.591
R12241 VDD.t143 VDD.n3432 136.591
R12242 VDD.t419 VDD.n5759 136.591
R12243 VDD.t667 VDD.n5505 136.591
R12244 VDD.t142 VDD.n3690 136.591
R12245 VDD.t782 VDD.n3948 136.591
R12246 VDD.t1087 VDD.n4206 136.591
R12247 VDD.t558 VDD.n4464 136.591
R12248 VDD.t572 VDD.n4722 136.591
R12249 VDD.t690 VDD.n4983 136.591
R12250 VDD.t418 VDD.n5245 136.591
R12251 VDD.n1697 VDD.n1696 135.117
R12252 VDD.n2046 VDD.n2045 135.117
R12253 VDD.n2276 VDD.n2275 135.117
R12254 VDD.n2534 VDD.n2533 135.117
R12255 VDD.n2792 VDD.n2791 135.117
R12256 VDD.n3050 VDD.n3049 135.117
R12257 VDD.n3308 VDD.n3307 135.117
R12258 VDD.n5638 VDD.n5637 135.117
R12259 VDD.n5384 VDD.n5383 135.117
R12260 VDD.n3566 VDD.n3565 135.117
R12261 VDD.n3824 VDD.n3823 135.117
R12262 VDD.n4082 VDD.n4081 135.117
R12263 VDD.n4340 VDD.n4339 135.117
R12264 VDD.n4598 VDD.n4597 135.117
R12265 VDD.n4856 VDD.n4855 135.117
R12266 VDD.n5148 VDD.n5147 135.117
R12267 VDD.t99 VDD.t1147 134.732
R12268 VDD.t1069 VDD.t653 134.732
R12269 VDD.t137 VDD.t672 134.732
R12270 VDD.t501 VDD.t56 134.732
R12271 VDD.n1371 VDD.t393 132.74
R12272 VDD VDD.t895 132.321
R12273 VDD.t879 VDD 132.321
R12274 VDD VDD.t859 132.321
R12275 VDD.t911 VDD.n985 132.321
R12276 VDD VDD.t821 132.321
R12277 VDD VDD.t426 132.321
R12278 VDD VDD.t1045 132.321
R12279 VDD.t1031 VDD 132.321
R12280 VDD VDD.t1009 132.321
R12281 VDD.t933 VDD.n190 132.321
R12282 VDD VDD.t971 132.321
R12283 VDD VDD.t1476 132.321
R12284 VDD VDD.t1421 132.321
R12285 VDD.t1405 VDD 132.321
R12286 VDD VDD.t1385 132.321
R12287 VDD VDD.t1347 132.321
R12288 VDD.n581 VDD.t532 132.321
R12289 VDD VDD.t508 132.321
R12290 VDD.t682 VDD.t99 131.983
R12291 VDD.t141 VDD.t1069 131.983
R12292 VDD.t178 VDD.t795 131.983
R12293 VDD.t578 VDD.t137 131.983
R12294 VDD.t777 VDD.t501 131.983
R12295 VDD.t1137 VDD.t127 131.983
R12296 VDD.n1715 VDD.n1672 131.388
R12297 VDD.n2064 VDD.n2021 131.388
R12298 VDD.n2294 VDD.n2251 131.388
R12299 VDD.n2552 VDD.n2509 131.388
R12300 VDD.n2810 VDD.n2767 131.388
R12301 VDD.n3068 VDD.n3025 131.388
R12302 VDD.n3326 VDD.n3283 131.388
R12303 VDD.n5656 VDD.n5613 131.388
R12304 VDD.n5402 VDD.n5359 131.388
R12305 VDD.n3584 VDD.n3541 131.388
R12306 VDD.n3842 VDD.n3799 131.388
R12307 VDD.n4100 VDD.n4057 131.388
R12308 VDD.n4358 VDD.n4315 131.388
R12309 VDD.n4616 VDD.n4573 131.388
R12310 VDD.n4874 VDD.n4831 131.388
R12311 VDD.n5166 VDD.n5123 131.388
R12312 VDD.n1766 VDD.n1673 131.012
R12313 VDD.n2115 VDD.n2022 131.012
R12314 VDD.n2345 VDD.n2252 131.012
R12315 VDD.n2603 VDD.n2510 131.012
R12316 VDD.n2861 VDD.n2768 131.012
R12317 VDD.n3119 VDD.n3026 131.012
R12318 VDD.n3377 VDD.n3284 131.012
R12319 VDD.n5707 VDD.n5614 131.012
R12320 VDD.n5453 VDD.n5360 131.012
R12321 VDD.n3635 VDD.n3542 131.012
R12322 VDD.n3893 VDD.n3800 131.012
R12323 VDD.n4151 VDD.n4058 131.012
R12324 VDD.n4409 VDD.n4316 131.012
R12325 VDD.n4667 VDD.n4574 131.012
R12326 VDD.n4925 VDD.n4832 131.012
R12327 VDD.n5217 VDD.n5124 131.012
R12328 VDD.n1767 VDD.n1672 130.636
R12329 VDD.n1767 VDD.n1766 130.636
R12330 VDD.n2116 VDD.n2021 130.636
R12331 VDD.n2116 VDD.n2115 130.636
R12332 VDD.n2346 VDD.n2251 130.636
R12333 VDD.n2346 VDD.n2345 130.636
R12334 VDD.n2604 VDD.n2509 130.636
R12335 VDD.n2604 VDD.n2603 130.636
R12336 VDD.n2862 VDD.n2767 130.636
R12337 VDD.n2862 VDD.n2861 130.636
R12338 VDD.n3120 VDD.n3025 130.636
R12339 VDD.n3120 VDD.n3119 130.636
R12340 VDD.n3378 VDD.n3283 130.636
R12341 VDD.n3378 VDD.n3377 130.636
R12342 VDD.n5708 VDD.n5613 130.636
R12343 VDD.n5708 VDD.n5707 130.636
R12344 VDD.n5454 VDD.n5359 130.636
R12345 VDD.n5454 VDD.n5453 130.636
R12346 VDD.n3636 VDD.n3541 130.636
R12347 VDD.n3636 VDD.n3635 130.636
R12348 VDD.n3894 VDD.n3799 130.636
R12349 VDD.n3894 VDD.n3893 130.636
R12350 VDD.n4152 VDD.n4057 130.636
R12351 VDD.n4152 VDD.n4151 130.636
R12352 VDD.n4410 VDD.n4315 130.636
R12353 VDD.n4410 VDD.n4409 130.636
R12354 VDD.n4668 VDD.n4573 130.636
R12355 VDD.n4668 VDD.n4667 130.636
R12356 VDD.n4926 VDD.n4831 130.636
R12357 VDD.n4926 VDD.n4925 130.636
R12358 VDD.n5218 VDD.n5123 130.636
R12359 VDD.n5218 VDD.n5217 130.636
R12360 VDD.n1879 VDD.n1823 129.691
R12361 VDD.n2200 VDD.n2144 129.691
R12362 VDD.n2458 VDD.n2402 129.691
R12363 VDD.n2716 VDD.n2660 129.691
R12364 VDD.n2974 VDD.n2918 129.691
R12365 VDD.n3232 VDD.n3176 129.691
R12366 VDD.n3490 VDD.n3434 129.691
R12367 VDD.n5817 VDD.n5761 129.691
R12368 VDD.n5563 VDD.n5507 129.691
R12369 VDD.n3748 VDD.n3692 129.691
R12370 VDD.n4006 VDD.n3950 129.691
R12371 VDD.n4264 VDD.n4208 129.691
R12372 VDD.n4522 VDD.n4466 129.691
R12373 VDD.n4780 VDD.n4724 129.691
R12374 VDD.n5041 VDD.n4985 129.691
R12375 VDD.n5303 VDD.n5247 129.691
R12376 VDD VDD.t698 129.228
R12377 VDD VDD.t72 129.228
R12378 VDD VDD.t1289 127.233
R12379 VDD VDD.t62 127.233
R12380 VDD VDD.t1079 127.233
R12381 VDD.t357 VDD 126.02
R12382 VDD.t150 VDD 126.02
R12383 VDD.t674 VDD 126.02
R12384 VDD.t1144 VDD 126.02
R12385 VDD.t91 VDD 126.02
R12386 VDD.t412 VDD 126.02
R12387 VDD.t1302 VDD 126.02
R12388 VDD.t157 VDD 126.02
R12389 VDD.t201 VDD 126.02
R12390 VDD.t1191 VDD 126.02
R12391 VDD.t678 VDD 126.02
R12392 VDD.t1149 VDD 126.02
R12393 VDD.t585 VDD 126.02
R12394 VDD.t1219 VDD 126.02
R12395 VDD.t583 VDD 126.02
R12396 VDD.t133 VDD 126.02
R12397 VDD.t546 VDD.t154 122.144
R12398 VDD.t391 VDD.t1255 122.144
R12399 VDD.t152 VDD.t47 122.144
R12400 VDD.n1903 VDD.n1898 121.977
R12401 VDD.n2224 VDD.n2219 121.977
R12402 VDD.n2482 VDD.n2477 121.977
R12403 VDD.n2740 VDD.n2735 121.977
R12404 VDD.n2998 VDD.n2993 121.977
R12405 VDD.n3256 VDD.n3251 121.977
R12406 VDD.n3514 VDD.n3509 121.977
R12407 VDD.n5841 VDD.n5836 121.977
R12408 VDD.n5587 VDD.n5582 121.977
R12409 VDD.n3772 VDD.n3767 121.977
R12410 VDD.n4030 VDD.n4025 121.977
R12411 VDD.n4288 VDD.n4283 121.977
R12412 VDD.n4546 VDD.n4541 121.977
R12413 VDD.n4804 VDD.n4799 121.977
R12414 VDD.n5065 VDD.n5060 121.977
R12415 VDD.n5327 VDD.n5322 121.977
R12416 VDD.t336 VDD.t1063 121.529
R12417 VDD.t766 VDD.t716 121.529
R12418 VDD.n1764 VDD.t753 121.114
R12419 VDD.t753 VDD.n1711 121.114
R12420 VDD.n2113 VDD.t129 121.114
R12421 VDD.t129 VDD.n2060 121.114
R12422 VDD.n2343 VDD.t70 121.114
R12423 VDD.t70 VDD.n2290 121.114
R12424 VDD.n2601 VDD.t680 121.114
R12425 VDD.t680 VDD.n2548 121.114
R12426 VDD.n2859 VDD.t733 121.114
R12427 VDD.t733 VDD.n2806 121.114
R12428 VDD.n3117 VDD.t125 121.114
R12429 VDD.t125 VDD.n3064 121.114
R12430 VDD.n3375 VDD.t504 121.114
R12431 VDD.t504 VDD.n3322 121.114
R12432 VDD.n5705 VDD.t4 121.114
R12433 VDD.t4 VDD.n5652 121.114
R12434 VDD.n5451 VDD.t665 121.114
R12435 VDD.t665 VDD.n5398 121.114
R12436 VDD.n3633 VDD.t1141 121.114
R12437 VDD.t1141 VDD.n3580 121.114
R12438 VDD.n3891 VDD.t1061 121.114
R12439 VDD.t1061 VDD.n3838 121.114
R12440 VDD.n4149 VDD.t414 121.114
R12441 VDD.t414 VDD.n4096 121.114
R12442 VDD.n4407 VDD.t165 121.114
R12443 VDD.t165 VDD.n4354 121.114
R12444 VDD.n4665 VDD.t793 121.114
R12445 VDD.t793 VDD.n4612 121.114
R12446 VDD.n4923 VDD.t1065 121.114
R12447 VDD.t1065 VDD.n4870 121.114
R12448 VDD.n5215 VDD.t107 121.114
R12449 VDD.t107 VDD.n5162 121.114
R12450 VDD.t1276 VDD.t1238 120.909
R12451 VDD.t1204 VDD.t700 120.909
R12452 VDD.t1132 VDD.t1169 120.909
R12453 VDD.t657 VDD.t731 120.909
R12454 VDD.n1853 VDD.n1845 120.094
R12455 VDD.n2174 VDD.n2166 120.094
R12456 VDD.n2432 VDD.n2424 120.094
R12457 VDD.n2690 VDD.n2682 120.094
R12458 VDD.n2948 VDD.n2940 120.094
R12459 VDD.n3206 VDD.n3198 120.094
R12460 VDD.n3464 VDD.n3456 120.094
R12461 VDD.n5791 VDD.n5783 120.094
R12462 VDD.n5537 VDD.n5529 120.094
R12463 VDD.n3722 VDD.n3714 120.094
R12464 VDD.n3980 VDD.n3972 120.094
R12465 VDD.n4238 VDD.n4230 120.094
R12466 VDD.n4496 VDD.n4488 120.094
R12467 VDD.n4754 VDD.n4746 120.094
R12468 VDD.n5015 VDD.n5007 120.094
R12469 VDD.n5277 VDD.n5269 120.094
R12470 VDD.n1 VDD.t1248 117.451
R12471 VDD.n785 VDD.t1207 117.451
R12472 VDD.n756 VDD.t1237 117.451
R12473 VDD.n776 VDD.t1208 117.451
R12474 VDD.n383 VDD.t662 117.451
R12475 VDD.n353 VDD.t1161 117.451
R12476 VDD.n373 VDD.t660 117.451
R12477 VDD.n318 VDD.t1181 117.451
R12478 VDD.n5 VDD.t1064 116.322
R12479 VDD.n811 VDD.t1277 116.322
R12480 VDD.n739 VDD.t460 116.322
R12481 VDD.n735 VDD.t699 116.322
R12482 VDD.n718 VDD.t458 116.322
R12483 VDD.n409 VDD.t1133 116.322
R12484 VDD.n322 VDD.t717 116.322
R12485 VDD.n1580 VDD.t1284 116.322
R12486 VDD.n1576 VDD.t73 116.322
R12487 VDD.n1559 VDD.t756 116.322
R12488 VDD.n1123 VDD.t1244 116.322
R12489 VDD.n1189 VDD.t1175 116.322
R12490 VDD.n1768 VDD.n1767 116.267
R12491 VDD.n2117 VDD.n2116 116.267
R12492 VDD.n2347 VDD.n2346 116.267
R12493 VDD.n2605 VDD.n2604 116.267
R12494 VDD.n2863 VDD.n2862 116.267
R12495 VDD.n3121 VDD.n3120 116.267
R12496 VDD.n3379 VDD.n3378 116.267
R12497 VDD.n5709 VDD.n5708 116.267
R12498 VDD.n5455 VDD.n5454 116.267
R12499 VDD.n3637 VDD.n3636 116.267
R12500 VDD.n3895 VDD.n3894 116.267
R12501 VDD.n4153 VDD.n4152 116.267
R12502 VDD.n4411 VDD.n4410 116.267
R12503 VDD.n4669 VDD.n4668 116.267
R12504 VDD.n4927 VDD.n4926 116.267
R12505 VDD.n5219 VDD.n5218 116.267
R12506 VDD.t89 VDD.t1243 115.486
R12507 VDD.t649 VDD.t1174 115.486
R12508 VDD.n987 VDD 115.358
R12509 VDD.n192 VDD 115.358
R12510 VDD.t1413 VDD.n579 115.358
R12511 VDD.n1907 VDD.n1888 112.189
R12512 VDD.n1854 VDD.n1843 112.189
R12513 VDD.n2175 VDD.n2164 112.189
R12514 VDD.n2228 VDD.n2209 112.189
R12515 VDD.n2433 VDD.n2422 112.189
R12516 VDD.n2486 VDD.n2467 112.189
R12517 VDD.n2691 VDD.n2680 112.189
R12518 VDD.n2744 VDD.n2725 112.189
R12519 VDD.n2949 VDD.n2938 112.189
R12520 VDD.n3002 VDD.n2983 112.189
R12521 VDD.n3207 VDD.n3196 112.189
R12522 VDD.n3260 VDD.n3241 112.189
R12523 VDD.n3465 VDD.n3454 112.189
R12524 VDD.n3518 VDD.n3499 112.189
R12525 VDD.n5792 VDD.n5781 112.189
R12526 VDD.n5845 VDD.n5826 112.189
R12527 VDD.n5538 VDD.n5527 112.189
R12528 VDD.n5591 VDD.n5572 112.189
R12529 VDD.n3723 VDD.n3712 112.189
R12530 VDD.n3776 VDD.n3757 112.189
R12531 VDD.n3981 VDD.n3970 112.189
R12532 VDD.n4034 VDD.n4015 112.189
R12533 VDD.n4239 VDD.n4228 112.189
R12534 VDD.n4292 VDD.n4273 112.189
R12535 VDD.n4497 VDD.n4486 112.189
R12536 VDD.n4550 VDD.n4531 112.189
R12537 VDD.n4755 VDD.n4744 112.189
R12538 VDD.n4808 VDD.n4789 112.189
R12539 VDD.n5069 VDD.n5050 112.189
R12540 VDD.n5016 VDD.n5005 112.189
R12541 VDD.n5331 VDD.n5312 112.189
R12542 VDD.n5278 VDD.n5267 112.189
R12543 VDD.t1232 VDD.t163 110.834
R12544 VDD.t1153 VDD.t747 110.834
R12545 VDD.t211 VDD.t321 109.316
R12546 VDD.t283 VDD.t211 109.316
R12547 VDD.t311 VDD.t283 109.316
R12548 VDD.t233 VDD.t311 109.316
R12549 VDD.t269 VDD.t233 109.316
R12550 VDD.t315 VDD.t269 109.316
R12551 VDD.t237 VDD.t315 109.316
R12552 VDD.t273 VDD.t237 109.316
R12553 VDD.t261 VDD.t273 109.316
R12554 VDD.t295 VDD.t261 109.316
R12555 VDD.t319 VDD.t295 109.316
R12556 VDD.t267 VDD.t319 109.316
R12557 VDD.t299 VDD.t267 109.316
R12558 VDD.t225 VDD.t299 109.316
R12559 VDD.t251 VDD.t225 109.316
R12560 VDD.t307 VDD.t229 109.316
R12561 VDD.t229 VDD.t263 109.316
R12562 VDD.t263 VDD.t215 109.316
R12563 VDD.t215 VDD.t305 109.316
R12564 VDD.t305 VDD.t329 109.316
R12565 VDD.t329 VDD.t257 109.316
R12566 VDD.t257 VDD.t289 109.316
R12567 VDD.t241 VDD.t317 109.316
R12568 VDD.t293 VDD.t241 109.316
R12569 VDD.t219 VDD.t293 109.316
R12570 VDD.t245 VDD.t219 109.316
R12571 VDD.t277 VDD.t245 109.316
R12572 VDD.t213 VDD.t277 109.316
R12573 VDD.t303 VDD.t213 109.316
R12574 VDD.t209 VDD.t281 109.316
R12575 VDD.t223 VDD.t249 109.316
R12576 VDD.t249 VDD.t301 109.316
R12577 VDD.t279 VDD.t309 109.316
R12578 VDD.t309 VDD.t231 109.316
R12579 VDD.t231 VDD.t327 109.316
R12580 VDD.t287 VDD.t255 109.316
R12581 VDD.t331 VDD.t287 109.316
R12582 VDD.t259 VDD.t331 109.316
R12583 VDD.t291 VDD.t217 109.316
R12584 VDD.t217 VDD.t243 109.316
R12585 VDD.t243 VDD.t275 109.316
R12586 VDD.t275 VDD.t221 109.316
R12587 VDD.t221 VDD.t247 109.316
R12588 VDD.t247 VDD.t325 109.316
R12589 VDD.t637 VDD.t643 109.316
R12590 VDD.t643 VDD.t621 109.316
R12591 VDD.t621 VDD.t631 109.316
R12592 VDD.t623 VDD.t641 109.316
R12593 VDD.t633 VDD.t623 109.316
R12594 VDD.t613 VDD.t633 109.316
R12595 VDD.t619 VDD.t629 109.316
R12596 VDD.t629 VDD.t625 109.316
R12597 VDD.t625 VDD.t639 109.316
R12598 VDD.t627 VDD.t617 109.316
R12599 VDD.t635 VDD.t627 109.316
R12600 VDD.t399 VDD.t395 109.316
R12601 VDD.t395 VDD.t397 109.316
R12602 VDD.t397 VDD.t401 109.316
R12603 VDD.t887 VDD.n984 108.572
R12604 VDD.t1037 VDD.n189 108.572
R12605 VDD.n582 VDD 108.572
R12606 VDD.t1467 VDD.t1281 106.709
R12607 VDD.t409 VDD.t167 106.709
R12608 VDD.t695 VDD.t86 103.636
R12609 VDD.t1059 VDD.t456 103.636
R12610 VDD.n1769 VDD.n1768 102.721
R12611 VDD.n1755 VDD.n1671 102.721
R12612 VDD.n2118 VDD.n2117 102.721
R12613 VDD.n2104 VDD.n2020 102.721
R12614 VDD.n2348 VDD.n2347 102.721
R12615 VDD.n2334 VDD.n2250 102.721
R12616 VDD.n2606 VDD.n2605 102.721
R12617 VDD.n2592 VDD.n2508 102.721
R12618 VDD.n2864 VDD.n2863 102.721
R12619 VDD.n2850 VDD.n2766 102.721
R12620 VDD.n3122 VDD.n3121 102.721
R12621 VDD.n3108 VDD.n3024 102.721
R12622 VDD.n3380 VDD.n3379 102.721
R12623 VDD.n3366 VDD.n3282 102.721
R12624 VDD.n5710 VDD.n5709 102.721
R12625 VDD.n5696 VDD.n5612 102.721
R12626 VDD.n5456 VDD.n5455 102.721
R12627 VDD.n5442 VDD.n5358 102.721
R12628 VDD.n3638 VDD.n3637 102.721
R12629 VDD.n3624 VDD.n3540 102.721
R12630 VDD.n3896 VDD.n3895 102.721
R12631 VDD.n3882 VDD.n3798 102.721
R12632 VDD.n4154 VDD.n4153 102.721
R12633 VDD.n4140 VDD.n4056 102.721
R12634 VDD.n4412 VDD.n4411 102.721
R12635 VDD.n4398 VDD.n4314 102.721
R12636 VDD.n4670 VDD.n4669 102.721
R12637 VDD.n4656 VDD.n4572 102.721
R12638 VDD.n4928 VDD.n4927 102.721
R12639 VDD.n4914 VDD.n4830 102.721
R12640 VDD.n5220 VDD.n5219 102.721
R12641 VDD.n5206 VDD.n5122 102.721
R12642 VDD VDD.t251 101.507
R12643 VDD.t301 VDD 101.507
R12644 VDD.t325 VDD 101.507
R12645 VDD.t615 VDD 101.507
R12646 VDD.t54 VDD 99.5973
R12647 VDD.t647 VDD 99.5973
R12648 VDD.t105 VDD 99.5973
R12649 VDD.t1118 VDD 99.5973
R12650 VDD.t403 VDD 99.5973
R12651 VDD.t774 VDD 99.5973
R12652 VDD.t181 VDD 99.5973
R12653 VDD.t712 VDD 99.5973
R12654 VDD.t598 VDD 99.5973
R12655 VDD.t343 VDD 99.5973
R12656 VDD.t565 VDD 99.5973
R12657 VDD.t1217 VDD 99.5973
R12658 VDD.t579 VDD 99.5973
R12659 VDD.t14 VDD 99.5973
R12660 VDD.t769 VDD 99.5973
R12661 VDD.t131 VDD 99.5973
R12662 VDD VDD.t459 99.5409
R12663 VDD VDD.t1163 99.5409
R12664 VDD.t191 VDD.t682 98.9875
R12665 VDD.t795 VDD.t141 98.9875
R12666 VDD.t1071 VDD.t578 98.9875
R12667 VDD.t127 VDD.t777 98.9875
R12668 VDD.n1429 VDD.t259 98.9046
R12669 VDD.t1318 VDD.t607 97.8793
R12670 VDD.t370 VDD.t739 97.8793
R12671 VDD.t401 VDD 97.6032
R12672 VDD.n31 VDD.t18 96.1553
R12673 VDD.n989 VDD.t547 96.1553
R12674 VDD.n825 VDD.t1466 96.1553
R12675 VDD.n752 VDD.t1117 96.1553
R12676 VDD.n721 VDD.t1 96.1553
R12677 VDD.n423 VDD.t408 96.1553
R12678 VDD.n348 VDD.t1325 96.1553
R12679 VDD.n1593 VDD.t744 96.1553
R12680 VDD.n1562 VDD.t1223 96.1553
R12681 VDD.n1117 VDD.t1070 96.1553
R12682 VDD.n1120 VDD.t100 96.1553
R12683 VDD.n194 VDD.t392 96.1553
R12684 VDD.n584 VDD.t153 96.1553
R12685 VDD.n1183 VDD.t502 96.1553
R12686 VDD.n1186 VDD.t138 96.1553
R12687 VDD.n902 VDD.t863 95.0005
R12688 VDD.n107 VDD.t1013 95.0005
R12689 VDD.t200 VDD 94.8523
R12690 VDD.t798 VDD 94.8523
R12691 VDD.n799 VDD.t1233 93.81
R12692 VDD.n397 VDD.t1154 93.81
R12693 VDD.t700 VDD 93.5611
R12694 VDD.t731 VDD 93.5611
R12695 VDD.t1253 VDD 93.539
R12696 VDD.t752 VDD 93.539
R12697 VDD VDD.t191 93.4882
R12698 VDD VDD.t1071 93.4882
R12699 VDD.t333 VDD 93.3702
R12700 VDD.t1213 VDD 93.3702
R12701 VDD.n1733 VDD.n1730 92.5005
R12702 VDD.n2082 VDD.n2079 92.5005
R12703 VDD.n2312 VDD.n2309 92.5005
R12704 VDD.n2570 VDD.n2567 92.5005
R12705 VDD.n2828 VDD.n2825 92.5005
R12706 VDD.n3086 VDD.n3083 92.5005
R12707 VDD.n3344 VDD.n3341 92.5005
R12708 VDD.n5674 VDD.n5671 92.5005
R12709 VDD.n5420 VDD.n5417 92.5005
R12710 VDD.n3602 VDD.n3599 92.5005
R12711 VDD.n3860 VDD.n3857 92.5005
R12712 VDD.n4118 VDD.n4115 92.5005
R12713 VDD.n4376 VDD.n4373 92.5005
R12714 VDD.n4634 VDD.n4631 92.5005
R12715 VDD.n4892 VDD.n4889 92.5005
R12716 VDD.n5184 VDD.n5181 92.5005
R12717 VDD.t359 VDD 92.1217
R12718 VDD.t728 VDD 92.1217
R12719 VDD.t605 VDD.t1245 91.8882
R12720 VDD.t737 VDD.t1177 91.8882
R12721 VDD.n1915 VDD.n1891 91.7652
R12722 VDD.n2236 VDD.n2212 91.7652
R12723 VDD.n2494 VDD.n2470 91.7652
R12724 VDD.n2752 VDD.n2728 91.7652
R12725 VDD.n3010 VDD.n2986 91.7652
R12726 VDD.n3268 VDD.n3244 91.7652
R12727 VDD.n3526 VDD.n3502 91.7652
R12728 VDD.n5853 VDD.n5829 91.7652
R12729 VDD.n5599 VDD.n5575 91.7652
R12730 VDD.n3784 VDD.n3760 91.7652
R12731 VDD.n4042 VDD.n4018 91.7652
R12732 VDD.n4300 VDD.n4276 91.7652
R12733 VDD.n4558 VDD.n4534 91.7652
R12734 VDD.n4816 VDD.n4792 91.7652
R12735 VDD.n5077 VDD.n5053 91.7652
R12736 VDD.n5339 VDD.n5315 91.7652
R12737 VDD.t1383 VDD.n500 91.6076
R12738 VDD.n1960 VDD.n1959 91.4829
R12739 VDD.n1959 VDD.n1929 91.4829
R12740 VDD.n1972 VDD.n1929 91.4829
R12741 VDD.n1972 VDD.n1971 91.4829
R12742 VDD.n1950 VDD.n1937 91.4829
R12743 VDD.n1965 VDD.n1937 91.4829
R12744 VDD.n1966 VDD.n1965 91.4829
R12745 VDD.n1967 VDD.n1966 91.4829
R12746 VDD.n1884 VDD.n1820 91.343
R12747 VDD.n2205 VDD.n2141 91.343
R12748 VDD.n2463 VDD.n2399 91.343
R12749 VDD.n2721 VDD.n2657 91.343
R12750 VDD.n2979 VDD.n2915 91.343
R12751 VDD.n3237 VDD.n3173 91.343
R12752 VDD.n3495 VDD.n3431 91.343
R12753 VDD.n5822 VDD.n5758 91.343
R12754 VDD.n5568 VDD.n5504 91.343
R12755 VDD.n3753 VDD.n3689 91.343
R12756 VDD.n4011 VDD.n3947 91.343
R12757 VDD.n4269 VDD.n4205 91.343
R12758 VDD.n4527 VDD.n4463 91.343
R12759 VDD.n4785 VDD.n4721 91.343
R12760 VDD.n5046 VDD.n4982 91.343
R12761 VDD.n5308 VDD.n5244 91.343
R12762 VDD.n1372 VDD.t635 91.0964
R12763 VDD.n1827 VDD.t357 89.1694
R12764 VDD.n2148 VDD.t150 89.1694
R12765 VDD.n2406 VDD.t674 89.1694
R12766 VDD.n2664 VDD.t1144 89.1694
R12767 VDD.n2922 VDD.t91 89.1694
R12768 VDD.n3180 VDD.t412 89.1694
R12769 VDD.n3438 VDD.t1302 89.1694
R12770 VDD.n5765 VDD.t157 89.1694
R12771 VDD.n5511 VDD.t201 89.1694
R12772 VDD.n3696 VDD.t1191 89.1694
R12773 VDD.n3954 VDD.t678 89.1694
R12774 VDD.n4212 VDD.t1149 89.1694
R12775 VDD.n4470 VDD.t585 89.1694
R12776 VDD.n4728 VDD.t1219 89.1694
R12777 VDD.n4989 VDD.t583 89.1694
R12778 VDD.n5251 VDD.t133 89.1694
R12779 VDD.t1247 VDD.t384 88.9241
R12780 VDD.t1180 VDD.t340 88.9241
R12781 VDD VDD.n1371 88.4936
R12782 VDD.n501 VDD.t1389 88.2148
R12783 VDD VDD.t178 87.9889
R12784 VDD VDD.t1137 87.9889
R12785 VDD.t380 VDD 87.8035
R12786 VDD.t1320 VDD 87.8035
R12787 VDD.t1264 VDD.t1060 87.6928
R12788 VDD.t1258 VDD.t1234 87.6928
R12789 VDD.t1130 VDD.t1093 87.6928
R12790 VDD.t128 VDD.t1156 87.6928
R12791 VDD.n7 VDD.t337 86.7743
R12792 VDD.n7 VDD.t606 86.7743
R12793 VDD.n788 VDD.t608 86.7743
R12794 VDD.n788 VDD.t164 86.7743
R12795 VDD.n758 VDD.t335 86.7743
R12796 VDD.n758 VDD.t609 86.7743
R12797 VDD.n760 VDD.t461 86.7743
R12798 VDD.n760 VDD.t140 86.7743
R12799 VDD.n386 VDD.t740 86.7743
R12800 VDD.n386 VDD.t748 86.7743
R12801 VDD.n355 VDD.t765 86.7743
R12802 VDD.n355 VDD.t742 86.7743
R12803 VDD.n357 VDD.t1328 86.7743
R12804 VDD.n357 VDD.t778 86.7743
R12805 VDD.n324 VDD.t767 86.7743
R12806 VDD.n324 VDD.t738 86.7743
R12807 VDD.t857 VDD.n901 84.8219
R12808 VDD.t1007 VDD.n106 84.8219
R12809 VDD.n755 VDD.n725 83.3098
R12810 VDD.n1596 VDD.n1566 83.3098
R12811 VDD.n1827 VDD.t382 81.2688
R12812 VDD.n2148 VDD.t1139 81.2688
R12813 VDD.n2406 VDD.t1297 81.2688
R12814 VDD.n2664 VDD.t95 81.2688
R12815 VDD.n2922 VDD.t462 81.2688
R12816 VDD.n3180 VDD.t1105 81.2688
R12817 VDD.n3438 VDD.t1259 81.2688
R12818 VDD.n5765 VDD.t1279 81.2688
R12819 VDD.n5511 VDD.t1299 81.2688
R12820 VDD.n3696 VDD.t1187 81.2688
R12821 VDD.n3954 VDD.t58 81.2688
R12822 VDD.n4212 VDD.t718 81.2688
R12823 VDD.n4470 VDD.t1202 81.2688
R12824 VDD.n4728 VDD.t602 81.2688
R12825 VDD.n4989 VDD.t1261 81.2688
R12826 VDD.n5251 VDD.t771 81.2688
R12827 VDD.n1457 VDD.t303 80.6854
R12828 VDD.n1760 VDD.n1717 80.5087
R12829 VDD.n2109 VDD.n2066 80.5087
R12830 VDD.n2339 VDD.n2296 80.5087
R12831 VDD.n2597 VDD.n2554 80.5087
R12832 VDD.n2855 VDD.n2812 80.5087
R12833 VDD.n3113 VDD.n3070 80.5087
R12834 VDD.n3371 VDD.n3328 80.5087
R12835 VDD.n5701 VDD.n5658 80.5087
R12836 VDD.n5447 VDD.n5404 80.5087
R12837 VDD.n3629 VDD.n3586 80.5087
R12838 VDD.n3887 VDD.n3844 80.5087
R12839 VDD.n4145 VDD.n4102 80.5087
R12840 VDD.n4403 VDD.n4360 80.5087
R12841 VDD.n4661 VDD.n4618 80.5087
R12842 VDD.n4919 VDD.n4876 80.5087
R12843 VDD.n5211 VDD.n5168 80.5087
R12844 VDD.n1708 VDD.n1669 80.2452
R12845 VDD.n2057 VDD.n2018 80.2452
R12846 VDD.n2287 VDD.n2248 80.2452
R12847 VDD.n2545 VDD.n2506 80.2452
R12848 VDD.n2803 VDD.n2764 80.2452
R12849 VDD.n3061 VDD.n3022 80.2452
R12850 VDD.n3319 VDD.n3280 80.2452
R12851 VDD.n5649 VDD.n5610 80.2452
R12852 VDD.n5395 VDD.n5356 80.2452
R12853 VDD.n3577 VDD.n3538 80.2452
R12854 VDD.n3835 VDD.n3796 80.2452
R12855 VDD.n4093 VDD.n4054 80.2452
R12856 VDD.n4351 VDD.n4312 80.2452
R12857 VDD.n4609 VDD.n4570 80.2452
R12858 VDD.n4867 VDD.n4828 80.2452
R12859 VDD.n5159 VDD.n5120 80.2452
R12860 VDD VDD.n1643 79.5475
R12861 VDD.t281 VDD.t323 78.5727
R12862 VDD VDD.n1634 78.5148
R12863 VDD.n1633 VDD.n1632 77.1383
R12864 VDD.n1870 VDD.n1845 76.5328
R12865 VDD.n2191 VDD.n2166 76.5328
R12866 VDD.n2449 VDD.n2424 76.5328
R12867 VDD.n2707 VDD.n2682 76.5328
R12868 VDD.n2965 VDD.n2940 76.5328
R12869 VDD.n3223 VDD.n3198 76.5328
R12870 VDD.n3481 VDD.n3456 76.5328
R12871 VDD.n5808 VDD.n5783 76.5328
R12872 VDD.n5554 VDD.n5529 76.5328
R12873 VDD.n3739 VDD.n3714 76.5328
R12874 VDD.n3997 VDD.n3972 76.5328
R12875 VDD.n4255 VDD.n4230 76.5328
R12876 VDD.n4513 VDD.n4488 76.5328
R12877 VDD.n4771 VDD.n4746 76.5328
R12878 VDD.n5032 VDD.n5007 76.5328
R12879 VDD.n5294 VDD.n5269 76.5328
R12880 VDD.n1625 VDD.n1624 76.0005
R12881 VDD.n1628 VDD.n1627 76.0005
R12882 VDD.n1630 VDD.n1629 76.0005
R12883 VDD.n1397 VDD.t613 75.48
R12884 VDD.n1869 VDD.n1844 74.1181
R12885 VDD.n2190 VDD.n2165 74.1181
R12886 VDD.n2448 VDD.n2423 74.1181
R12887 VDD.n2706 VDD.n2681 74.1181
R12888 VDD.n2964 VDD.n2939 74.1181
R12889 VDD.n3222 VDD.n3197 74.1181
R12890 VDD.n3480 VDD.n3455 74.1181
R12891 VDD.n5807 VDD.n5782 74.1181
R12892 VDD.n5553 VDD.n5528 74.1181
R12893 VDD.n3738 VDD.n3713 74.1181
R12894 VDD.n3996 VDD.n3971 74.1181
R12895 VDD.n4254 VDD.n4229 74.1181
R12896 VDD.n4512 VDD.n4487 74.1181
R12897 VDD.n4770 VDD.n4745 74.1181
R12898 VDD.n5031 VDD.n5006 74.1181
R12899 VDD.n5293 VDD.n5268 74.1181
R12900 VDD.n1871 VDD.n1843 71.6136
R12901 VDD.n2192 VDD.n2164 71.6136
R12902 VDD.n2450 VDD.n2422 71.6136
R12903 VDD.n2708 VDD.n2680 71.6136
R12904 VDD.n2966 VDD.n2938 71.6136
R12905 VDD.n3224 VDD.n3196 71.6136
R12906 VDD.n3482 VDD.n3454 71.6136
R12907 VDD.n5809 VDD.n5781 71.6136
R12908 VDD.n5555 VDD.n5527 71.6136
R12909 VDD.n3740 VDD.n3712 71.6136
R12910 VDD.n3998 VDD.n3970 71.6136
R12911 VDD.n4256 VDD.n4228 71.6136
R12912 VDD.n4514 VDD.n4486 71.6136
R12913 VDD.n4772 VDD.n4744 71.6136
R12914 VDD.n5033 VDD.n5005 71.6136
R12915 VDD.n5295 VDD.n5267 71.6136
R12916 VDD.n1809 VDD.t54 70.4844
R12917 VDD.n2130 VDD.t647 70.4844
R12918 VDD.n2388 VDD.t105 70.4844
R12919 VDD.n2646 VDD.t1118 70.4844
R12920 VDD.n2904 VDD.t403 70.4844
R12921 VDD.n3162 VDD.t774 70.4844
R12922 VDD.n3420 VDD.t181 70.4844
R12923 VDD.n5747 VDD.t712 70.4844
R12924 VDD.n5493 VDD.t598 70.4844
R12925 VDD.n3678 VDD.t343 70.4844
R12926 VDD.n3936 VDD.t565 70.4844
R12927 VDD.n4194 VDD.t1217 70.4844
R12928 VDD.n4452 VDD.t579 70.4844
R12929 VDD.n4710 VDD.t14 70.4844
R12930 VDD.n4971 VDD.t769 70.4844
R12931 VDD.n5233 VDD.t131 70.4844
R12932 VDD.t1060 VDD.t457 70.1543
R12933 VDD.t1093 VDD.t755 70.1543
R12934 VDD.n1877 VDD.n1876 66.2808
R12935 VDD.n2198 VDD.n2197 66.2808
R12936 VDD.n2456 VDD.n2455 66.2808
R12937 VDD.n2714 VDD.n2713 66.2808
R12938 VDD.n2972 VDD.n2971 66.2808
R12939 VDD.n3230 VDD.n3229 66.2808
R12940 VDD.n3488 VDD.n3487 66.2808
R12941 VDD.n5815 VDD.n5814 66.2808
R12942 VDD.n5561 VDD.n5560 66.2808
R12943 VDD.n3746 VDD.n3745 66.2808
R12944 VDD.n4004 VDD.n4003 66.2808
R12945 VDD.n4262 VDD.n4261 66.2808
R12946 VDD.n4520 VDD.n4519 66.2808
R12947 VDD.n4778 VDD.n4777 66.2808
R12948 VDD.n5039 VDD.n5038 66.2808
R12949 VDD.n5301 VDD.n5300 66.2808
R12950 VDD.n1898 VDD.n1889 65.0929
R12951 VDD.n2219 VDD.n2210 65.0929
R12952 VDD.n2477 VDD.n2468 65.0929
R12953 VDD.n2735 VDD.n2726 65.0929
R12954 VDD.n2993 VDD.n2984 65.0929
R12955 VDD.n3251 VDD.n3242 65.0929
R12956 VDD.n3509 VDD.n3500 65.0929
R12957 VDD.n5836 VDD.n5827 65.0929
R12958 VDD.n5582 VDD.n5573 65.0929
R12959 VDD.n3767 VDD.n3758 65.0929
R12960 VDD.n4025 VDD.n4016 65.0929
R12961 VDD.n4283 VDD.n4274 65.0929
R12962 VDD.n4541 VDD.n4532 65.0929
R12963 VDD.n4799 VDD.n4790 65.0929
R12964 VDD.n5060 VDD.n5051 65.0929
R12965 VDD.n5322 VDD.n5313 65.0929
R12966 VDD.n1809 VDD.t1095 64.3553
R12967 VDD.n2130 VDD.t683 64.3553
R12968 VDD.n2388 VDD.t74 64.3553
R12969 VDD.n2646 VDD.t499 64.3553
R12970 VDD.n2904 VDD.t714 64.3553
R12971 VDD.n3162 VDD.t685 64.3553
R12972 VDD.n3420 VDD.t360 64.3553
R12973 VDD.n5747 VDD.t338 64.3553
R12974 VDD.n5493 VDD.t1316 64.3553
R12975 VDD.n3678 VDD.t1182 64.3553
R12976 VDD.n3936 VDD.t655 64.3553
R12977 VDD.n4194 VDD.t488 64.3553
R12978 VDD.n4452 VDD.t87 64.3553
R12979 VDD.n4710 VDD.t1189 64.3553
R12980 VDD.n4971 VDD.t1266 64.3553
R12981 VDD.n5233 VDD.t1500 64.3553
R12982 VDD.n792 VDD.t1205 63.3219
R12983 VDD.n792 VDD.t701 63.3219
R12984 VDD.n390 VDD.t658 63.3219
R12985 VDD.n390 VDD.t732 63.3219
R12986 VDD.n1706 VDD.n1673 63.2691
R12987 VDD.n1707 VDD.n1706 63.2691
R12988 VDD.n2055 VDD.n2022 63.2691
R12989 VDD.n2056 VDD.n2055 63.2691
R12990 VDD.n2285 VDD.n2252 63.2691
R12991 VDD.n2286 VDD.n2285 63.2691
R12992 VDD.n2543 VDD.n2510 63.2691
R12993 VDD.n2544 VDD.n2543 63.2691
R12994 VDD.n2801 VDD.n2768 63.2691
R12995 VDD.n2802 VDD.n2801 63.2691
R12996 VDD.n3059 VDD.n3026 63.2691
R12997 VDD.n3060 VDD.n3059 63.2691
R12998 VDD.n3317 VDD.n3284 63.2691
R12999 VDD.n3318 VDD.n3317 63.2691
R13000 VDD.n5647 VDD.n5614 63.2691
R13001 VDD.n5648 VDD.n5647 63.2691
R13002 VDD.n5393 VDD.n5360 63.2691
R13003 VDD.n5394 VDD.n5393 63.2691
R13004 VDD.n3575 VDD.n3542 63.2691
R13005 VDD.n3576 VDD.n3575 63.2691
R13006 VDD.n3833 VDD.n3800 63.2691
R13007 VDD.n3834 VDD.n3833 63.2691
R13008 VDD.n4091 VDD.n4058 63.2691
R13009 VDD.n4092 VDD.n4091 63.2691
R13010 VDD.n4349 VDD.n4316 63.2691
R13011 VDD.n4350 VDD.n4349 63.2691
R13012 VDD.n4607 VDD.n4574 63.2691
R13013 VDD.n4608 VDD.n4607 63.2691
R13014 VDD.n4865 VDD.n4832 63.2691
R13015 VDD.n4866 VDD.n4865 63.2691
R13016 VDD.n5157 VDD.n5124 63.2691
R13017 VDD.n5158 VDD.n5157 63.2691
R13018 VDD.n1762 VDD.n1715 61.5116
R13019 VDD.n1762 VDD.n1761 61.5116
R13020 VDD.n2111 VDD.n2064 61.5116
R13021 VDD.n2111 VDD.n2110 61.5116
R13022 VDD.n2341 VDD.n2294 61.5116
R13023 VDD.n2341 VDD.n2340 61.5116
R13024 VDD.n2599 VDD.n2552 61.5116
R13025 VDD.n2599 VDD.n2598 61.5116
R13026 VDD.n2857 VDD.n2810 61.5116
R13027 VDD.n2857 VDD.n2856 61.5116
R13028 VDD.n3115 VDD.n3068 61.5116
R13029 VDD.n3115 VDD.n3114 61.5116
R13030 VDD.n3373 VDD.n3326 61.5116
R13031 VDD.n3373 VDD.n3372 61.5116
R13032 VDD.n5703 VDD.n5656 61.5116
R13033 VDD.n5703 VDD.n5702 61.5116
R13034 VDD.n5449 VDD.n5402 61.5116
R13035 VDD.n5449 VDD.n5448 61.5116
R13036 VDD.n3631 VDD.n3584 61.5116
R13037 VDD.n3631 VDD.n3630 61.5116
R13038 VDD.n3889 VDD.n3842 61.5116
R13039 VDD.n3889 VDD.n3888 61.5116
R13040 VDD.n4147 VDD.n4100 61.5116
R13041 VDD.n4147 VDD.n4146 61.5116
R13042 VDD.n4405 VDD.n4358 61.5116
R13043 VDD.n4405 VDD.n4404 61.5116
R13044 VDD.n4663 VDD.n4616 61.5116
R13045 VDD.n4663 VDD.n4662 61.5116
R13046 VDD.n4921 VDD.n4874 61.5116
R13047 VDD.n4921 VDD.n4920 61.5116
R13048 VDD.n5213 VDD.n5166 61.5116
R13049 VDD.n5213 VDD.n5212 61.5116
R13050 VDD.n1908 VDD.n1897 60.6123
R13051 VDD.n1911 VDD.n1910 60.6123
R13052 VDD.n1910 VDD.n1903 60.6123
R13053 VDD.n1908 VDD.n1907 60.6123
R13054 VDD.n1860 VDD.n1852 60.6123
R13055 VDD.n1866 VDD.n1853 60.6123
R13056 VDD.n1866 VDD.n1865 60.6123
R13057 VDD.n1854 VDD.n1852 60.6123
R13058 VDD.n2181 VDD.n2173 60.6123
R13059 VDD.n2187 VDD.n2174 60.6123
R13060 VDD.n2187 VDD.n2186 60.6123
R13061 VDD.n2175 VDD.n2173 60.6123
R13062 VDD.n2229 VDD.n2218 60.6123
R13063 VDD.n2232 VDD.n2231 60.6123
R13064 VDD.n2231 VDD.n2224 60.6123
R13065 VDD.n2229 VDD.n2228 60.6123
R13066 VDD.n2439 VDD.n2431 60.6123
R13067 VDD.n2445 VDD.n2432 60.6123
R13068 VDD.n2445 VDD.n2444 60.6123
R13069 VDD.n2433 VDD.n2431 60.6123
R13070 VDD.n2487 VDD.n2476 60.6123
R13071 VDD.n2490 VDD.n2489 60.6123
R13072 VDD.n2489 VDD.n2482 60.6123
R13073 VDD.n2487 VDD.n2486 60.6123
R13074 VDD.n2697 VDD.n2689 60.6123
R13075 VDD.n2703 VDD.n2690 60.6123
R13076 VDD.n2703 VDD.n2702 60.6123
R13077 VDD.n2691 VDD.n2689 60.6123
R13078 VDD.n2745 VDD.n2734 60.6123
R13079 VDD.n2748 VDD.n2747 60.6123
R13080 VDD.n2747 VDD.n2740 60.6123
R13081 VDD.n2745 VDD.n2744 60.6123
R13082 VDD.n2955 VDD.n2947 60.6123
R13083 VDD.n2961 VDD.n2948 60.6123
R13084 VDD.n2961 VDD.n2960 60.6123
R13085 VDD.n2949 VDD.n2947 60.6123
R13086 VDD.n3003 VDD.n2992 60.6123
R13087 VDD.n3006 VDD.n3005 60.6123
R13088 VDD.n3005 VDD.n2998 60.6123
R13089 VDD.n3003 VDD.n3002 60.6123
R13090 VDD.n3213 VDD.n3205 60.6123
R13091 VDD.n3219 VDD.n3206 60.6123
R13092 VDD.n3219 VDD.n3218 60.6123
R13093 VDD.n3207 VDD.n3205 60.6123
R13094 VDD.n3261 VDD.n3250 60.6123
R13095 VDD.n3264 VDD.n3263 60.6123
R13096 VDD.n3263 VDD.n3256 60.6123
R13097 VDD.n3261 VDD.n3260 60.6123
R13098 VDD.n3471 VDD.n3463 60.6123
R13099 VDD.n3477 VDD.n3464 60.6123
R13100 VDD.n3477 VDD.n3476 60.6123
R13101 VDD.n3465 VDD.n3463 60.6123
R13102 VDD.n3519 VDD.n3508 60.6123
R13103 VDD.n3522 VDD.n3521 60.6123
R13104 VDD.n3521 VDD.n3514 60.6123
R13105 VDD.n3519 VDD.n3518 60.6123
R13106 VDD.n5798 VDD.n5790 60.6123
R13107 VDD.n5804 VDD.n5791 60.6123
R13108 VDD.n5804 VDD.n5803 60.6123
R13109 VDD.n5792 VDD.n5790 60.6123
R13110 VDD.n5846 VDD.n5835 60.6123
R13111 VDD.n5849 VDD.n5848 60.6123
R13112 VDD.n5848 VDD.n5841 60.6123
R13113 VDD.n5846 VDD.n5845 60.6123
R13114 VDD.n5544 VDD.n5536 60.6123
R13115 VDD.n5550 VDD.n5537 60.6123
R13116 VDD.n5550 VDD.n5549 60.6123
R13117 VDD.n5538 VDD.n5536 60.6123
R13118 VDD.n5592 VDD.n5581 60.6123
R13119 VDD.n5595 VDD.n5594 60.6123
R13120 VDD.n5594 VDD.n5587 60.6123
R13121 VDD.n5592 VDD.n5591 60.6123
R13122 VDD.n3729 VDD.n3721 60.6123
R13123 VDD.n3735 VDD.n3722 60.6123
R13124 VDD.n3735 VDD.n3734 60.6123
R13125 VDD.n3723 VDD.n3721 60.6123
R13126 VDD.n3777 VDD.n3766 60.6123
R13127 VDD.n3780 VDD.n3779 60.6123
R13128 VDD.n3779 VDD.n3772 60.6123
R13129 VDD.n3777 VDD.n3776 60.6123
R13130 VDD.n3987 VDD.n3979 60.6123
R13131 VDD.n3993 VDD.n3980 60.6123
R13132 VDD.n3993 VDD.n3992 60.6123
R13133 VDD.n3981 VDD.n3979 60.6123
R13134 VDD.n4035 VDD.n4024 60.6123
R13135 VDD.n4038 VDD.n4037 60.6123
R13136 VDD.n4037 VDD.n4030 60.6123
R13137 VDD.n4035 VDD.n4034 60.6123
R13138 VDD.n4245 VDD.n4237 60.6123
R13139 VDD.n4251 VDD.n4238 60.6123
R13140 VDD.n4251 VDD.n4250 60.6123
R13141 VDD.n4239 VDD.n4237 60.6123
R13142 VDD.n4293 VDD.n4282 60.6123
R13143 VDD.n4296 VDD.n4295 60.6123
R13144 VDD.n4295 VDD.n4288 60.6123
R13145 VDD.n4293 VDD.n4292 60.6123
R13146 VDD.n4503 VDD.n4495 60.6123
R13147 VDD.n4509 VDD.n4496 60.6123
R13148 VDD.n4509 VDD.n4508 60.6123
R13149 VDD.n4497 VDD.n4495 60.6123
R13150 VDD.n4551 VDD.n4540 60.6123
R13151 VDD.n4554 VDD.n4553 60.6123
R13152 VDD.n4553 VDD.n4546 60.6123
R13153 VDD.n4551 VDD.n4550 60.6123
R13154 VDD.n4761 VDD.n4753 60.6123
R13155 VDD.n4767 VDD.n4754 60.6123
R13156 VDD.n4767 VDD.n4766 60.6123
R13157 VDD.n4755 VDD.n4753 60.6123
R13158 VDD.n4809 VDD.n4798 60.6123
R13159 VDD.n4812 VDD.n4811 60.6123
R13160 VDD.n4811 VDD.n4804 60.6123
R13161 VDD.n4809 VDD.n4808 60.6123
R13162 VDD.n5070 VDD.n5059 60.6123
R13163 VDD.n5073 VDD.n5072 60.6123
R13164 VDD.n5072 VDD.n5065 60.6123
R13165 VDD.n5070 VDD.n5069 60.6123
R13166 VDD.n5022 VDD.n5014 60.6123
R13167 VDD.n5028 VDD.n5015 60.6123
R13168 VDD.n5028 VDD.n5027 60.6123
R13169 VDD.n5016 VDD.n5014 60.6123
R13170 VDD.n5332 VDD.n5321 60.6123
R13171 VDD.n5335 VDD.n5334 60.6123
R13172 VDD.n5334 VDD.n5327 60.6123
R13173 VDD.n5332 VDD.n5331 60.6123
R13174 VDD.n5284 VDD.n5276 60.6123
R13175 VDD.n5290 VDD.n5277 60.6123
R13176 VDD.n5290 VDD.n5289 60.6123
R13177 VDD.n5278 VDD.n5276 60.6123
R13178 VDD.n1456 VDD.t279 59.8635
R13179 VDD.n1916 VDD.n1888 58.0325
R13180 VDD.n2237 VDD.n2209 58.0325
R13181 VDD.n2495 VDD.n2467 58.0325
R13182 VDD.n2753 VDD.n2725 58.0325
R13183 VDD.n3011 VDD.n2983 58.0325
R13184 VDD.n3269 VDD.n3241 58.0325
R13185 VDD.n3527 VDD.n3499 58.0325
R13186 VDD.n5854 VDD.n5826 58.0325
R13187 VDD.n5600 VDD.n5572 58.0325
R13188 VDD.n3785 VDD.n3757 58.0325
R13189 VDD.n4043 VDD.n4015 58.0325
R13190 VDD.n4301 VDD.n4273 58.0325
R13191 VDD.n4559 VDD.n4531 58.0325
R13192 VDD.n4817 VDD.n4789 58.0325
R13193 VDD.n5078 VDD.n5050 58.0325
R13194 VDD.n5340 VDD.n5312 58.0325
R13195 VDD.n901 VDD.t831 57.6791
R13196 VDD.n106 VDD.t979 57.6791
R13197 VDD.t1238 VDD.t380 57.5763
R13198 VDD.t1169 VDD.t1320 57.5763
R13199 VDD VDD.t176 57.5434
R13200 VDD VDD.t741 57.5434
R13201 VDD.t1245 VDD.t333 56.3188
R13202 VDD.t1177 VDD.t1213 56.3188
R13203 VDD.n1732 VDD.n1731 55.4672
R13204 VDD.n1733 VDD.n1729 55.4672
R13205 VDD.n2081 VDD.n2080 55.4672
R13206 VDD.n2082 VDD.n2078 55.4672
R13207 VDD.n2311 VDD.n2310 55.4672
R13208 VDD.n2312 VDD.n2308 55.4672
R13209 VDD.n2569 VDD.n2568 55.4672
R13210 VDD.n2570 VDD.n2566 55.4672
R13211 VDD.n2827 VDD.n2826 55.4672
R13212 VDD.n2828 VDD.n2824 55.4672
R13213 VDD.n3085 VDD.n3084 55.4672
R13214 VDD.n3086 VDD.n3082 55.4672
R13215 VDD.n3343 VDD.n3342 55.4672
R13216 VDD.n3344 VDD.n3340 55.4672
R13217 VDD.n5673 VDD.n5672 55.4672
R13218 VDD.n5674 VDD.n5670 55.4672
R13219 VDD.n5419 VDD.n5418 55.4672
R13220 VDD.n5420 VDD.n5416 55.4672
R13221 VDD.n3601 VDD.n3600 55.4672
R13222 VDD.n3602 VDD.n3598 55.4672
R13223 VDD.n3859 VDD.n3858 55.4672
R13224 VDD.n3860 VDD.n3856 55.4672
R13225 VDD.n4117 VDD.n4116 55.4672
R13226 VDD.n4118 VDD.n4114 55.4672
R13227 VDD.n4375 VDD.n4374 55.4672
R13228 VDD.n4376 VDD.n4372 55.4672
R13229 VDD.n4633 VDD.n4632 55.4672
R13230 VDD.n4634 VDD.n4630 55.4672
R13231 VDD.n4891 VDD.n4890 55.4672
R13232 VDD.n4892 VDD.n4888 55.4672
R13233 VDD.n5183 VDD.n5182 55.4672
R13234 VDD.n5184 VDD.n5180 55.4672
R13235 VDD.n1803 VDD 54.4858
R13236 VDD.n2011 VDD 54.4858
R13237 VDD.n2382 VDD 54.4858
R13238 VDD.n2640 VDD 54.4858
R13239 VDD.n2898 VDD 54.4858
R13240 VDD.n3156 VDD 54.4858
R13241 VDD.n3414 VDD 54.4858
R13242 VDD.n5744 VDD 54.4858
R13243 VDD.n5490 VDD 54.4858
R13244 VDD.n3672 VDD 54.4858
R13245 VDD.n3930 VDD 54.4858
R13246 VDD.n4188 VDD 54.4858
R13247 VDD.n4446 VDD 54.4858
R13248 VDD.n4704 VDD 54.4858
R13249 VDD.n4963 VDD 54.4858
R13250 VDD.n5113 VDD 54.4858
R13251 VDD.t1055 VDD.n1927 54.472
R13252 VDD.t1287 VDD.n1927 54.472
R13253 VDD.n501 VDD.t1423 54.2862
R13254 VDD.n1953 VDD.t1285 54.2478
R13255 VDD.n1949 VDD.n1941 54.1098
R13256 VDD.n1969 VDD.n1931 54.1091
R13257 VDD.t0 VDD.t1264 52.6159
R13258 VDD.t1234 VDD.t1253 52.6159
R13259 VDD.t1222 VDD.t1130 52.6159
R13260 VDD.t1156 VDD.t752 52.6159
R13261 VDD.n500 VDD.t1355 50.8934
R13262 VDD.t1055 VDD.n1939 50.8854
R13263 VDD.t45 VDD.t16 50.6439
R13264 VDD.t52 VDD.t410 50.6439
R13265 VDD.n1876 VDD.n1818 50.1034
R13266 VDD.n2197 VDD.n2139 50.1034
R13267 VDD.n2455 VDD.n2397 50.1034
R13268 VDD.n2713 VDD.n2655 50.1034
R13269 VDD.n2971 VDD.n2913 50.1034
R13270 VDD.n3229 VDD.n3171 50.1034
R13271 VDD.n3487 VDD.n3429 50.1034
R13272 VDD.n5814 VDD.n5756 50.1034
R13273 VDD.n5560 VDD.n5502 50.1034
R13274 VDD.n3745 VDD.n3687 50.1034
R13275 VDD.n4003 VDD.n3945 50.1034
R13276 VDD.n4261 VDD.n4203 50.1034
R13277 VDD.n4519 VDD.n4461 50.1034
R13278 VDD.n4777 VDD.n4719 50.1034
R13279 VDD.n5038 VDD.n4980 50.1034
R13280 VDD.n5300 VDD.n5242 50.1034
R13281 VDD.t227 VDD.n1456 49.4526
R13282 VDD.t323 VDD.t253 49.2598
R13283 VDD.t253 VDD.t285 49.2598
R13284 VDD.t285 VDD.t313 49.2598
R13285 VDD.t313 VDD.t235 49.2598
R13286 VDD.t235 VDD.t271 49.2598
R13287 VDD.t271 VDD.t207 49.2598
R13288 VDD.t207 VDD.t239 49.2598
R13289 VDD.t239 VDD.t205 49.2598
R13290 VDD.t205 VDD.t265 49.2598
R13291 VDD.t265 VDD.t297 49.2598
R13292 VDD.t39 VDD.n1801 49.1183
R13293 VDD.t362 VDD.n2009 49.1183
R13294 VDD.t464 VDD.n2380 49.1183
R13295 VDD.t119 VDD.n2638 49.1183
R13296 VDD.t19 VDD.n2896 49.1183
R13297 VDD.t588 VDD.n3154 49.1183
R13298 VDD.t548 VDD.n3412 49.1183
R13299 VDD.t168 VDD.n5742 49.1183
R13300 VDD.t759 VDD.n5488 49.1183
R13301 VDD.t1097 VDD.n3670 49.1183
R13302 VDD.t783 VDD.n3928 49.1183
R13303 VDD.t492 VDD.n4186 49.1183
R13304 VDD.t372 VDD.n4444 49.1183
R13305 VDD.t109 VDD.n4702 49.1183
R13306 VDD.t347 VDD.n4961 49.1183
R13307 VDD.t480 VDD.n5111 49.1183
R13308 VDD.t297 VDD.t223 47.9846
R13309 VDD.n902 VDD.t897 47.5005
R13310 VDD.n107 VDD.t1047 47.5005
R13311 VDD.n1700 VDD.n1681 47.0405
R13312 VDD.n2049 VDD.n2030 47.0405
R13313 VDD.n2279 VDD.n2260 47.0405
R13314 VDD.n2537 VDD.n2518 47.0405
R13315 VDD.n2795 VDD.n2776 47.0405
R13316 VDD.n3053 VDD.n3034 47.0405
R13317 VDD.n3311 VDD.n3292 47.0405
R13318 VDD.n5641 VDD.n5622 47.0405
R13319 VDD.n5387 VDD.n5368 47.0405
R13320 VDD.n3569 VDD.n3550 47.0405
R13321 VDD.n3827 VDD.n3808 47.0405
R13322 VDD.n4085 VDD.n4066 47.0405
R13323 VDD.n4343 VDD.n4324 47.0405
R13324 VDD.n4601 VDD.n4582 47.0405
R13325 VDD.n4859 VDD.n4840 47.0405
R13326 VDD.n5151 VDD.n5132 47.0405
R13327 VDD.n1966 VDD.n1936 46.6829
R13328 VDD.n1973 VDD.n1972 45.9299
R13329 VDD.n1959 VDD.n1958 45.9299
R13330 VDD.n1705 VDD.n1704 45.7605
R13331 VDD.n1689 VDD.n1685 45.7605
R13332 VDD.n2054 VDD.n2053 45.7605
R13333 VDD.n2038 VDD.n2034 45.7605
R13334 VDD.n2284 VDD.n2283 45.7605
R13335 VDD.n2268 VDD.n2264 45.7605
R13336 VDD.n2542 VDD.n2541 45.7605
R13337 VDD.n2526 VDD.n2522 45.7605
R13338 VDD.n2800 VDD.n2799 45.7605
R13339 VDD.n2784 VDD.n2780 45.7605
R13340 VDD.n3058 VDD.n3057 45.7605
R13341 VDD.n3042 VDD.n3038 45.7605
R13342 VDD.n3316 VDD.n3315 45.7605
R13343 VDD.n3300 VDD.n3296 45.7605
R13344 VDD.n5646 VDD.n5645 45.7605
R13345 VDD.n5630 VDD.n5626 45.7605
R13346 VDD.n5392 VDD.n5391 45.7605
R13347 VDD.n5376 VDD.n5372 45.7605
R13348 VDD.n3574 VDD.n3573 45.7605
R13349 VDD.n3558 VDD.n3554 45.7605
R13350 VDD.n3832 VDD.n3831 45.7605
R13351 VDD.n3816 VDD.n3812 45.7605
R13352 VDD.n4090 VDD.n4089 45.7605
R13353 VDD.n4074 VDD.n4070 45.7605
R13354 VDD.n4348 VDD.n4347 45.7605
R13355 VDD.n4332 VDD.n4328 45.7605
R13356 VDD.n4606 VDD.n4605 45.7605
R13357 VDD.n4590 VDD.n4586 45.7605
R13358 VDD.n4864 VDD.n4863 45.7605
R13359 VDD.n4848 VDD.n4844 45.7605
R13360 VDD.n5156 VDD.n5155 45.7605
R13361 VDD.n5140 VDD.n5136 45.7605
R13362 VDD.n1684 VDD.n1682 45.4405
R13363 VDD.n2033 VDD.n2031 45.4405
R13364 VDD.n2263 VDD.n2261 45.4405
R13365 VDD.n2521 VDD.n2519 45.4405
R13366 VDD.n2779 VDD.n2777 45.4405
R13367 VDD.n3037 VDD.n3035 45.4405
R13368 VDD.n3295 VDD.n3293 45.4405
R13369 VDD.n5625 VDD.n5623 45.4405
R13370 VDD.n5371 VDD.n5369 45.4405
R13371 VDD.n3553 VDD.n3551 45.4405
R13372 VDD.n3811 VDD.n3809 45.4405
R13373 VDD.n4069 VDD.n4067 45.4405
R13374 VDD.n4327 VDD.n4325 45.4405
R13375 VDD.n4585 VDD.n4583 45.4405
R13376 VDD.n4843 VDD.n4841 45.4405
R13377 VDD.n5135 VDD.n5133 45.4405
R13378 VDD.n1947 VDD.n1937 44.8005
R13379 VDD.n725 VDD 43.6586
R13380 VDD.n1566 VDD 43.6586
R13381 VDD.n1 VDD.t697 42.3555
R13382 VDD.n785 VDD.t381 42.3555
R13383 VDD.n756 VDD.t1210 42.3555
R13384 VDD.n776 VDD.t156 42.3555
R13385 VDD.n383 VDD.t1321 42.3555
R13386 VDD.n353 VDD.t797 42.3555
R13387 VDD.n373 VDD.t102 42.3555
R13388 VDD.n318 VDD.t136 42.3555
R13389 VDD.n1947 VDD.n1946 41.323
R13390 VDD.n1936 VDD.n1933 41.2617
R13391 VDD.n1708 VDD.n1707 39.5299
R13392 VDD.n1761 VDD.n1760 39.5299
R13393 VDD.n2057 VDD.n2056 39.5299
R13394 VDD.n2110 VDD.n2109 39.5299
R13395 VDD.n2287 VDD.n2286 39.5299
R13396 VDD.n2340 VDD.n2339 39.5299
R13397 VDD.n2545 VDD.n2544 39.5299
R13398 VDD.n2598 VDD.n2597 39.5299
R13399 VDD.n2803 VDD.n2802 39.5299
R13400 VDD.n2856 VDD.n2855 39.5299
R13401 VDD.n3061 VDD.n3060 39.5299
R13402 VDD.n3114 VDD.n3113 39.5299
R13403 VDD.n3319 VDD.n3318 39.5299
R13404 VDD.n3372 VDD.n3371 39.5299
R13405 VDD.n5649 VDD.n5648 39.5299
R13406 VDD.n5702 VDD.n5701 39.5299
R13407 VDD.n5395 VDD.n5394 39.5299
R13408 VDD.n5448 VDD.n5447 39.5299
R13409 VDD.n3577 VDD.n3576 39.5299
R13410 VDD.n3630 VDD.n3629 39.5299
R13411 VDD.n3835 VDD.n3834 39.5299
R13412 VDD.n3888 VDD.n3887 39.5299
R13413 VDD.n4093 VDD.n4092 39.5299
R13414 VDD.n4146 VDD.n4145 39.5299
R13415 VDD.n4351 VDD.n4350 39.5299
R13416 VDD.n4404 VDD.n4403 39.5299
R13417 VDD.n4609 VDD.n4608 39.5299
R13418 VDD.n4662 VDD.n4661 39.5299
R13419 VDD.n4867 VDD.n4866 39.5299
R13420 VDD.n4920 VDD.n4919 39.5299
R13421 VDD.n5159 VDD.n5158 39.5299
R13422 VDD.n5212 VDD.n5211 39.5299
R13423 VDD.n20 VDD.n3 39.2858
R13424 VDD.n337 VDD.n320 39.2858
R13425 VDD VDD.t139 39.0862
R13426 VDD VDD.t659 39.0862
R13427 VDD.n1885 VDD.n1884 38.9491
R13428 VDD.n2206 VDD.n2205 38.9491
R13429 VDD.n2464 VDD.n2463 38.9491
R13430 VDD.n2722 VDD.n2721 38.9491
R13431 VDD.n2980 VDD.n2979 38.9491
R13432 VDD.n3238 VDD.n3237 38.9491
R13433 VDD.n3496 VDD.n3495 38.9491
R13434 VDD.n5823 VDD.n5822 38.9491
R13435 VDD.n5569 VDD.n5568 38.9491
R13436 VDD.n3754 VDD.n3753 38.9491
R13437 VDD.n4012 VDD.n4011 38.9491
R13438 VDD.n4270 VDD.n4269 38.9491
R13439 VDD.n4528 VDD.n4527 38.9491
R13440 VDD.n4786 VDD.n4785 38.9491
R13441 VDD.n5047 VDD.n5046 38.9491
R13442 VDD.n5309 VDD.n5308 38.9491
R13443 VDD.t607 VDD.t1232 38.8641
R13444 VDD.t739 VDD.t1153 38.8641
R13445 VDD.t384 VDD.t336 38.534
R13446 VDD.t340 VDD.t766 38.534
R13447 VDD.n1746 VDD.n1745 37.3765
R13448 VDD.n1728 VDD.n1725 37.3765
R13449 VDD.n2095 VDD.n2094 37.3765
R13450 VDD.n2077 VDD.n2074 37.3765
R13451 VDD.n2325 VDD.n2324 37.3765
R13452 VDD.n2307 VDD.n2304 37.3765
R13453 VDD.n2583 VDD.n2582 37.3765
R13454 VDD.n2565 VDD.n2562 37.3765
R13455 VDD.n2841 VDD.n2840 37.3765
R13456 VDD.n2823 VDD.n2820 37.3765
R13457 VDD.n3099 VDD.n3098 37.3765
R13458 VDD.n3081 VDD.n3078 37.3765
R13459 VDD.n3357 VDD.n3356 37.3765
R13460 VDD.n3339 VDD.n3336 37.3765
R13461 VDD.n5687 VDD.n5686 37.3765
R13462 VDD.n5669 VDD.n5666 37.3765
R13463 VDD.n5433 VDD.n5432 37.3765
R13464 VDD.n5415 VDD.n5412 37.3765
R13465 VDD.n3615 VDD.n3614 37.3765
R13466 VDD.n3597 VDD.n3594 37.3765
R13467 VDD.n3873 VDD.n3872 37.3765
R13468 VDD.n3855 VDD.n3852 37.3765
R13469 VDD.n4131 VDD.n4130 37.3765
R13470 VDD.n4113 VDD.n4110 37.3765
R13471 VDD.n4389 VDD.n4388 37.3765
R13472 VDD.n4371 VDD.n4368 37.3765
R13473 VDD.n4647 VDD.n4646 37.3765
R13474 VDD.n4629 VDD.n4626 37.3765
R13475 VDD.n4905 VDD.n4904 37.3765
R13476 VDD.n4887 VDD.n4884 37.3765
R13477 VDD.n5197 VDD.n5196 37.3765
R13478 VDD.n5179 VDD.n5176 37.3765
R13479 VDD.n1830 VDD.t383 36.1587
R13480 VDD.n1830 VDD.t358 36.1587
R13481 VDD.n1813 VDD.t1096 36.1587
R13482 VDD.n1813 VDD.t55 36.1587
R13483 VDD.n2134 VDD.t684 36.1587
R13484 VDD.n2134 VDD.t648 36.1587
R13485 VDD.n2151 VDD.t1140 36.1587
R13486 VDD.n2151 VDD.t151 36.1587
R13487 VDD.n2392 VDD.t75 36.1587
R13488 VDD.n2392 VDD.t106 36.1587
R13489 VDD.n2409 VDD.t1298 36.1587
R13490 VDD.n2409 VDD.t675 36.1587
R13491 VDD.n2650 VDD.t500 36.1587
R13492 VDD.n2650 VDD.t1119 36.1587
R13493 VDD.n2667 VDD.t96 36.1587
R13494 VDD.n2667 VDD.t1145 36.1587
R13495 VDD.n2908 VDD.t715 36.1587
R13496 VDD.n2908 VDD.t404 36.1587
R13497 VDD.n2925 VDD.t463 36.1587
R13498 VDD.n2925 VDD.t92 36.1587
R13499 VDD.n3166 VDD.t686 36.1587
R13500 VDD.n3166 VDD.t775 36.1587
R13501 VDD.n3183 VDD.t1106 36.1587
R13502 VDD.n3183 VDD.t413 36.1587
R13503 VDD.n3424 VDD.t361 36.1587
R13504 VDD.n3424 VDD.t182 36.1587
R13505 VDD.n3441 VDD.t1260 36.1587
R13506 VDD.n3441 VDD.t1303 36.1587
R13507 VDD.n5751 VDD.t339 36.1587
R13508 VDD.n5751 VDD.t713 36.1587
R13509 VDD.n5768 VDD.t1280 36.1587
R13510 VDD.n5768 VDD.t158 36.1587
R13511 VDD.n5497 VDD.t1317 36.1587
R13512 VDD.n5497 VDD.t599 36.1587
R13513 VDD.n5514 VDD.t1300 36.1587
R13514 VDD.n5514 VDD.t202 36.1587
R13515 VDD.n3682 VDD.t1183 36.1587
R13516 VDD.n3682 VDD.t344 36.1587
R13517 VDD.n3699 VDD.t1188 36.1587
R13518 VDD.n3699 VDD.t1192 36.1587
R13519 VDD.n3940 VDD.t656 36.1587
R13520 VDD.n3940 VDD.t566 36.1587
R13521 VDD.n3957 VDD.t59 36.1587
R13522 VDD.n3957 VDD.t679 36.1587
R13523 VDD.n4198 VDD.t489 36.1587
R13524 VDD.n4198 VDD.t1218 36.1587
R13525 VDD.n4215 VDD.t719 36.1587
R13526 VDD.n4215 VDD.t1150 36.1587
R13527 VDD.n4456 VDD.t88 36.1587
R13528 VDD.n4456 VDD.t580 36.1587
R13529 VDD.n4473 VDD.t1203 36.1587
R13530 VDD.n4473 VDD.t586 36.1587
R13531 VDD.n4714 VDD.t1190 36.1587
R13532 VDD.n4714 VDD.t15 36.1587
R13533 VDD.n4731 VDD.t603 36.1587
R13534 VDD.n4731 VDD.t1220 36.1587
R13535 VDD.n4992 VDD.t1262 36.1587
R13536 VDD.n4992 VDD.t584 36.1587
R13537 VDD.n4975 VDD.t1267 36.1587
R13538 VDD.n4975 VDD.t770 36.1587
R13539 VDD.n5254 VDD.t772 36.1587
R13540 VDD.n5254 VDD.t134 36.1587
R13541 VDD.n5237 VDD.t1501 36.1587
R13542 VDD.n5237 VDD.t132 36.1587
R13543 VDD.t457 VDD.t1258 35.0774
R13544 VDD.t755 VDD.t128 35.0774
R13545 VDD VDD.n1802 34.927
R13546 VDD VDD.n2010 34.927
R13547 VDD VDD.n2381 34.927
R13548 VDD VDD.n2639 34.927
R13549 VDD VDD.n2897 34.927
R13550 VDD VDD.n3155 34.927
R13551 VDD VDD.n3413 34.927
R13552 VDD VDD.n5743 34.927
R13553 VDD VDD.n5489 34.927
R13554 VDD VDD.n3671 34.927
R13555 VDD VDD.n3929 34.927
R13556 VDD VDD.n4187 34.927
R13557 VDD VDD.n4445 34.927
R13558 VDD VDD.n4703 34.927
R13559 VDD VDD.n4962 34.927
R13560 VDD VDD.n5112 34.927
R13561 VDD.n23 VDD.n2 34.6358
R13562 VDD.n18 VDD.n6 34.6358
R13563 VDD.n996 VDD.n995 34.6358
R13564 VDD.n817 VDD.n816 34.6358
R13565 VDD.n744 VDD.n743 34.6358
R13566 VDD.n415 VDD.n414 34.6358
R13567 VDD.n340 VDD.n319 34.6358
R13568 VDD.n335 VDD.n323 34.6358
R13569 VDD.n1585 VDD.n1584 34.6358
R13570 VDD.n1149 VDD.n1148 34.6358
R13571 VDD.n1161 VDD.n1160 34.6358
R13572 VDD.n1167 VDD.n1166 34.6358
R13573 VDD.n1130 VDD.n1118 34.6358
R13574 VDD.n1134 VDD.n1118 34.6358
R13575 VDD.n1135 VDD.n1134 34.6358
R13576 VDD.n1128 VDD.n1121 34.6358
R13577 VDD.n201 VDD.n200 34.6358
R13578 VDD.n591 VDD.n590 34.6358
R13579 VDD.n1215 VDD.n1214 34.6358
R13580 VDD.n1227 VDD.n1226 34.6358
R13581 VDD.n1233 VDD.n1232 34.6358
R13582 VDD.n1196 VDD.n1184 34.6358
R13583 VDD.n1200 VDD.n1184 34.6358
R13584 VDD.n1201 VDD.n1200 34.6358
R13585 VDD.n1194 VDD.n1187 34.6358
R13586 VDD.n984 VDD.t823 33.9291
R13587 VDD.n189 VDD.t973 33.9291
R13588 VDD.n1155 VDD.n1154 33.8829
R13589 VDD.n1221 VDD.n1220 33.8829
R13590 VDD.n1958 VDD.n1957 33.8422
R13591 VDD.n1397 VDD.t619 33.8361
R13592 VDD.n1973 VDD.n1923 33.6292
R13593 VDD.t1063 VDD.t605 32.6058
R13594 VDD.t716 VDD.t737 32.6058
R13595 VDD.t176 VDD.t1209 31.4862
R13596 VDD.t139 VDD.t155 31.4862
R13597 VDD.t741 VDD.t796 31.4862
R13598 VDD.t659 VDD.t101 31.4862
R13599 VDD.n1914 VDD.t420 30.1961
R13600 VDD.n2235 VDD.t148 30.1961
R13601 VDD.n2493 VDD.t676 30.1961
R13602 VDD.n2751 VDD.t689 30.1961
R13603 VDD.n3009 VDD.t93 30.1961
R13604 VDD.n3267 VDD.t76 30.1961
R13605 VDD.n3525 VDD.t1186 30.1961
R13606 VDD.n5852 VDD.t159 30.1961
R13607 VDD.n5598 VDD.t203 30.1961
R13608 VDD.n3783 VDD.t556 30.1961
R13609 VDD.n4041 VDD.t562 30.1961
R13610 VDD.n4299 VDD.t687 30.1961
R13611 VDD.n4557 VDD.t570 30.1961
R13612 VDD.n4815 VDD.t670 30.1961
R13613 VDD.n5076 VDD.t581 30.1961
R13614 VDD.n5338 VDD.t97 30.1961
R13615 VDD.n859 VDD.n858 29.3652
R13616 VDD.n938 VDD.n937 29.3652
R13617 VDD.n834 VDD.n833 29.3652
R13618 VDD.n837 VDD.n836 29.3652
R13619 VDD.n64 VDD.n63 29.3652
R13620 VDD.n143 VDD.n142 29.3652
R13621 VDD.n39 VDD.n38 29.3652
R13622 VDD.n42 VDD.n41 29.3652
R13623 VDD.n458 VDD.n457 29.3652
R13624 VDD.n537 VDD.n536 29.3652
R13625 VDD.n433 VDD.n432 29.3652
R13626 VDD.n436 VDD.n435 29.3652
R13627 VDD.n1313 VDD.n1312 29.3652
R13628 VDD.n1342 VDD.n1341 29.3652
R13629 VDD.n840 VDD.n839 28.9887
R13630 VDD.n45 VDD.n44 28.9887
R13631 VDD.n439 VDD.n438 28.9887
R13632 VDD.n1348 VDD.n1347 28.9887
R13633 VDD.n5 VDD.t385 28.4628
R13634 VDD.n811 VDD.t162 28.4628
R13635 VDD.n739 VDD.t1251 28.4628
R13636 VDD.n735 VDD.t1278 28.4628
R13637 VDD.n718 VDD.t1265 28.4628
R13638 VDD.n409 VDD.t49 28.4628
R13639 VDD.n322 VDD.t341 28.4628
R13640 VDD.n1580 VDD.t346 28.4628
R13641 VDD.n1576 VDD.t53 28.4628
R13642 VDD.n1559 VDD.t1131 28.4628
R13643 VDD.n1123 VDD.t646 28.4628
R13644 VDD.n1189 VDD.t28 28.4628
R13645 VDD.n1793 VDD.n1782 28.2358
R13646 VDD.n1794 VDD.n1793 28.2358
R13647 VDD.n1790 VDD.n1787 28.2358
R13648 VDD.n1790 VDD.n1789 28.2358
R13649 VDD.n2001 VDD.n1990 28.2358
R13650 VDD.n2002 VDD.n2001 28.2358
R13651 VDD.n1998 VDD.n1995 28.2358
R13652 VDD.n1998 VDD.n1997 28.2358
R13653 VDD.n2372 VDD.n2361 28.2358
R13654 VDD.n2373 VDD.n2372 28.2358
R13655 VDD.n2369 VDD.n2366 28.2358
R13656 VDD.n2369 VDD.n2368 28.2358
R13657 VDD.n2630 VDD.n2619 28.2358
R13658 VDD.n2631 VDD.n2630 28.2358
R13659 VDD.n2627 VDD.n2624 28.2358
R13660 VDD.n2627 VDD.n2626 28.2358
R13661 VDD.n2888 VDD.n2877 28.2358
R13662 VDD.n2889 VDD.n2888 28.2358
R13663 VDD.n2885 VDD.n2882 28.2358
R13664 VDD.n2885 VDD.n2884 28.2358
R13665 VDD.n3146 VDD.n3135 28.2358
R13666 VDD.n3147 VDD.n3146 28.2358
R13667 VDD.n3143 VDD.n3140 28.2358
R13668 VDD.n3143 VDD.n3142 28.2358
R13669 VDD.n3404 VDD.n3393 28.2358
R13670 VDD.n3405 VDD.n3404 28.2358
R13671 VDD.n3401 VDD.n3398 28.2358
R13672 VDD.n3401 VDD.n3400 28.2358
R13673 VDD.n5734 VDD.n5723 28.2358
R13674 VDD.n5735 VDD.n5734 28.2358
R13675 VDD.n5731 VDD.n5728 28.2358
R13676 VDD.n5731 VDD.n5730 28.2358
R13677 VDD.n5480 VDD.n5469 28.2358
R13678 VDD.n5481 VDD.n5480 28.2358
R13679 VDD.n5477 VDD.n5474 28.2358
R13680 VDD.n5477 VDD.n5476 28.2358
R13681 VDD.n3662 VDD.n3651 28.2358
R13682 VDD.n3663 VDD.n3662 28.2358
R13683 VDD.n3659 VDD.n3656 28.2358
R13684 VDD.n3659 VDD.n3658 28.2358
R13685 VDD.n3920 VDD.n3909 28.2358
R13686 VDD.n3921 VDD.n3920 28.2358
R13687 VDD.n3917 VDD.n3914 28.2358
R13688 VDD.n3917 VDD.n3916 28.2358
R13689 VDD.n4178 VDD.n4167 28.2358
R13690 VDD.n4179 VDD.n4178 28.2358
R13691 VDD.n4175 VDD.n4172 28.2358
R13692 VDD.n4175 VDD.n4174 28.2358
R13693 VDD.n4436 VDD.n4425 28.2358
R13694 VDD.n4437 VDD.n4436 28.2358
R13695 VDD.n4433 VDD.n4430 28.2358
R13696 VDD.n4433 VDD.n4432 28.2358
R13697 VDD.n4694 VDD.n4683 28.2358
R13698 VDD.n4695 VDD.n4694 28.2358
R13699 VDD.n4691 VDD.n4688 28.2358
R13700 VDD.n4691 VDD.n4690 28.2358
R13701 VDD.n4953 VDD.n4942 28.2358
R13702 VDD.n4954 VDD.n4953 28.2358
R13703 VDD.n4950 VDD.n4947 28.2358
R13704 VDD.n4950 VDD.n4949 28.2358
R13705 VDD.n5103 VDD.n5092 28.2358
R13706 VDD.n5104 VDD.n5103 28.2358
R13707 VDD.n5100 VDD.n5097 28.2358
R13708 VDD.n5100 VDD.n5099 28.2358
R13709 VDD.n13 VDD.n8 28.2358
R13710 VDD.n330 VDD.n325 28.2358
R13711 VDD.n780 VDD 28.2291
R13712 VDD.n377 VDD 28.2291
R13713 VDD.n579 VDD.t1349 27.1434
R13714 VDD.n799 VDD.t1319 26.9729
R13715 VDD.n397 VDD.t371 26.9729
R13716 VDD.n1835 VDD.n1834 26.8623
R13717 VDD.n2156 VDD.n2155 26.8623
R13718 VDD.n2414 VDD.n2413 26.8623
R13719 VDD.n2672 VDD.n2671 26.8623
R13720 VDD.n2930 VDD.n2929 26.8623
R13721 VDD.n3188 VDD.n3187 26.8623
R13722 VDD.n3446 VDD.n3445 26.8623
R13723 VDD.n5773 VDD.n5772 26.8623
R13724 VDD.n5519 VDD.n5518 26.8623
R13725 VDD.n3704 VDD.n3703 26.8623
R13726 VDD.n3962 VDD.n3961 26.8623
R13727 VDD.n4220 VDD.n4219 26.8623
R13728 VDD.n4478 VDD.n4477 26.8623
R13729 VDD.n4736 VDD.n4735 26.8623
R13730 VDD.n4997 VDD.n4996 26.8623
R13731 VDD.n5259 VDD.n5258 26.8623
R13732 VDD.n1656 VDD 26.615
R13733 VDD.n31 VDD.t1283 26.5955
R13734 VDD.n825 VDD.t1108 26.5955
R13735 VDD.n752 VDD.t46 26.5955
R13736 VDD.n721 VDD.t746 26.5955
R13737 VDD.n423 VDD.t730 26.5955
R13738 VDD.n348 VDD.t1327 26.5955
R13739 VDD.n1593 VDD.t411 26.5955
R13740 VDD.n1562 VDD.t390 26.5955
R13741 VDD.n1117 VDD.t654 26.5955
R13742 VDD.n1120 VDD.t1148 26.5955
R13743 VDD.n1183 VDD.t57 26.5955
R13744 VDD.n1186 VDD.t673 26.5955
R13745 VDD.n1792 VDD.t43 26.5955
R13746 VDD.n1792 VDD.t40 26.5955
R13747 VDD.n1788 VDD.t1226 26.5955
R13748 VDD.n1788 VDD.t1230 26.5955
R13749 VDD.n2000 VDD.t364 26.5955
R13750 VDD.n2000 VDD.t368 26.5955
R13751 VDD.n1996 VDD.t35 26.5955
R13752 VDD.n1996 VDD.t32 26.5955
R13753 VDD.n2371 VDD.t468 26.5955
R13754 VDD.n2371 VDD.t470 26.5955
R13755 VDD.n2367 VDD.t544 26.5955
R13756 VDD.n2367 VDD.t539 26.5955
R13757 VDD.n2629 VDD.t121 26.5955
R13758 VDD.n2629 VDD.t122 26.5955
R13759 VDD.n2625 VDD.t476 26.5955
R13760 VDD.n2625 VDD.t478 26.5955
R13761 VDD.n2887 VDD.t23 26.5955
R13762 VDD.n2887 VDD.t25 26.5955
R13763 VDD.n2883 VDD.t1308 26.5955
R13764 VDD.n2883 VDD.t1311 26.5955
R13765 VDD.n3145 VDD.t592 26.5955
R13766 VDD.n3145 VDD.t594 26.5955
R13767 VDD.n3141 VDD.t13 26.5955
R13768 VDD.n3141 VDD.t9 26.5955
R13769 VDD.n3403 VDD.t552 26.5955
R13770 VDD.n3403 VDD.t554 26.5955
R13771 VDD.n3399 VDD.t1198 26.5955
R13772 VDD.n3399 VDD.t1200 26.5955
R13773 VDD.n5733 VDD.t172 26.5955
R13774 VDD.n5733 VDD.t174 26.5955
R13775 VDD.n5729 VDD.t706 26.5955
R13776 VDD.n5729 VDD.t709 26.5955
R13777 VDD.n5479 VDD.t764 26.5955
R13778 VDD.n5479 VDD.t760 26.5955
R13779 VDD.n5475 VDD.t1334 26.5955
R13780 VDD.n5475 VDD.t1336 26.5955
R13781 VDD.n3661 VDD.t1102 26.5955
R13782 VDD.n3661 VDD.t1104 26.5955
R13783 VDD.n3657 VDD.t1272 26.5955
R13784 VDD.n3657 VDD.t1274 26.5955
R13785 VDD.n3919 VDD.t784 26.5955
R13786 VDD.n3919 VDD.t787 26.5955
R13787 VDD.n3915 VDD.t84 26.5955
R13788 VDD.n3915 VDD.t79 26.5955
R13789 VDD.n4177 VDD.t497 26.5955
R13790 VDD.n4177 VDD.t493 26.5955
R13791 VDD.n4173 VDD.t726 26.5955
R13792 VDD.n4173 VDD.t721 26.5955
R13793 VDD.n4435 VDD.t376 26.5955
R13794 VDD.n4435 VDD.t378 26.5955
R13795 VDD.n4431 VDD.t1111 26.5955
R13796 VDD.n4431 VDD.t1114 26.5955
R13797 VDD.n4693 VDD.t113 26.5955
R13798 VDD.n4693 VDD.t115 26.5955
R13799 VDD.n4689 VDD.t190 26.5955
R13800 VDD.n4689 VDD.t186 26.5955
R13801 VDD.n4952 VDD.t351 26.5955
R13802 VDD.n4952 VDD.t353 26.5955
R13803 VDD.n4948 VDD.t1125 26.5955
R13804 VDD.n4948 VDD.t1127 26.5955
R13805 VDD.n5102 VDD.t484 26.5955
R13806 VDD.n5102 VDD.t486 26.5955
R13807 VDD.n5098 VDD.t194 26.5955
R13808 VDD.n5098 VDD.t197 26.5955
R13809 VDD.n1009 VDD.t1294 26.5955
R13810 VDD.n1009 VDD.t1296 26.5955
R13811 VDD.n872 VDD.t920 26.5955
R13812 VDD.n872 VDD.t852 26.5955
R13813 VDD.n878 VDD.t826 26.5955
R13814 VDD.n878 VDD.t890 26.5955
R13815 VDD.n884 VDD.t906 26.5955
R13816 VDD.n884 VDD.t802 26.5955
R13817 VDD.n890 VDD.t800 26.5955
R13818 VDD.n890 VDD.t836 26.5955
R13819 VDD.n895 VDD.t832 26.5955
R13820 VDD.n895 VDD.t858 26.5955
R13821 VDD.n851 VDD.t818 26.5955
R13822 VDD.n851 VDD.t810 26.5955
R13823 VDD.n846 VDD.t840 26.5955
R13824 VDD.n846 VDD.t926 26.5955
R13825 VDD.n930 VDD.t924 26.5955
R13826 VDD.n930 VDD.t856 26.5955
R13827 VDD.n924 VDD.t850 26.5955
R13828 VDD.n924 VDD.t876 26.5955
R13829 VDD.n918 VDD.t838 26.5955
R13830 VDD.n918 VDD.t918 26.5955
R13831 VDD.n912 VDD.t868 26.5955
R13832 VDD.n912 VDD.t902 26.5955
R13833 VDD.n908 VDD.t898 26.5955
R13834 VDD.n908 VDD.t830 26.5955
R13835 VDD.n842 VDD.t808 26.5955
R13836 VDD.n842 VDD.t864 26.5955
R13837 VDD.n862 VDD.t884 26.5955
R13838 VDD.n862 VDD.t910 26.5955
R13839 VDD.n955 VDD.t820 26.5955
R13840 VDD.n955 VDD.t842 26.5955
R13841 VDD.n961 VDD.t848 26.5955
R13842 VDD.n961 VDD.t874 26.5955
R13843 VDD.n967 VDD.t872 26.5955
R13844 VDD.n967 VDD.t904 26.5955
R13845 VDD.n973 VDD.t916 26.5955
R13846 VDD.n973 VDD.t846 26.5955
R13847 VDD.n978 VDD.t824 26.5955
R13848 VDD.n978 VDD.t888 26.5955
R13849 VDD.n948 VDD.t828 26.5955
R13850 VDD.n948 VDD.t914 26.5955
R13851 VDD.n942 VDD.t862 26.5955
R13852 VDD.n942 VDD.t892 26.5955
R13853 VDD.n1065 VDD.t854 26.5955
R13854 VDD.n1065 VDD.t878 26.5955
R13855 VDD.n1071 VDD.t894 26.5955
R13856 VDD.n1071 VDD.t922 26.5955
R13857 VDD.n1077 VDD.t870 26.5955
R13858 VDD.n1077 VDD.t812 26.5955
R13859 VDD.n1083 VDD.t900 26.5955
R13860 VDD.n1083 VDD.t834 26.5955
R13861 VDD.n1087 VDD.t844 26.5955
R13862 VDD.n1087 VDD.t866 26.5955
R13863 VDD.n1094 VDD.t886 26.5955
R13864 VDD.n1094 VDD.t912 26.5955
R13865 VDD.n1102 VDD.t908 26.5955
R13866 VDD.n1102 VDD.t806 26.5955
R13867 VDD.n1018 VDD.t429 26.5955
R13868 VDD.n1018 VDD.t443 26.5955
R13869 VDD.n1024 VDD.t441 26.5955
R13870 VDD.n1024 VDD.t425 26.5955
R13871 VDD.n1030 VDD.t455 26.5955
R13872 VDD.n1030 VDD.t435 26.5955
R13873 VDD.n1036 VDD.t433 26.5955
R13874 VDD.n1036 VDD.t447 26.5955
R13875 VDD.n1040 VDD.t445 26.5955
R13876 VDD.n1040 VDD.t453 26.5955
R13877 VDD.n1046 VDD.t439 26.5955
R13878 VDD.n1046 VDD.t449 26.5955
R13879 VDD.n1054 VDD.t451 26.5955
R13880 VDD.n1054 VDD.t431 26.5955
R13881 VDD.n214 VDD.t67 26.5955
R13882 VDD.n214 VDD.t61 26.5955
R13883 VDD.n77 VDD.t942 26.5955
R13884 VDD.n77 VDD.t1002 26.5955
R13885 VDD.n83 VDD.t976 26.5955
R13886 VDD.n83 VDD.t1040 26.5955
R13887 VDD.n89 VDD.t928 26.5955
R13888 VDD.n89 VDD.t952 26.5955
R13889 VDD.n95 VDD.t950 26.5955
R13890 VDD.n95 VDD.t986 26.5955
R13891 VDD.n100 VDD.t980 26.5955
R13892 VDD.n100 VDD.t1008 26.5955
R13893 VDD.n56 VDD.t968 26.5955
R13894 VDD.n56 VDD.t960 26.5955
R13895 VDD.n51 VDD.t990 26.5955
R13896 VDD.n51 VDD.t948 26.5955
R13897 VDD.n135 VDD.t946 26.5955
R13898 VDD.n135 VDD.t1006 26.5955
R13899 VDD.n129 VDD.t1000 26.5955
R13900 VDD.n129 VDD.t1028 26.5955
R13901 VDD.n123 VDD.t988 26.5955
R13902 VDD.n123 VDD.t940 26.5955
R13903 VDD.n117 VDD.t1020 26.5955
R13904 VDD.n117 VDD.t1052 26.5955
R13905 VDD.n113 VDD.t1048 26.5955
R13906 VDD.n113 VDD.t982 26.5955
R13907 VDD.n47 VDD.t958 26.5955
R13908 VDD.n47 VDD.t1014 26.5955
R13909 VDD.n67 VDD.t1016 26.5955
R13910 VDD.n67 VDD.t932 26.5955
R13911 VDD.n160 VDD.t970 26.5955
R13912 VDD.n160 VDD.t992 26.5955
R13913 VDD.n166 VDD.t998 26.5955
R13914 VDD.n166 VDD.t1026 26.5955
R13915 VDD.n172 VDD.t1024 26.5955
R13916 VDD.n172 VDD.t1054 26.5955
R13917 VDD.n178 VDD.t938 26.5955
R13918 VDD.n178 VDD.t996 26.5955
R13919 VDD.n183 VDD.t974 26.5955
R13920 VDD.n183 VDD.t1038 26.5955
R13921 VDD.n153 VDD.t978 26.5955
R13922 VDD.n153 VDD.t936 26.5955
R13923 VDD.n147 VDD.t1012 26.5955
R13924 VDD.n147 VDD.t1042 26.5955
R13925 VDD.n270 VDD.t1004 26.5955
R13926 VDD.n270 VDD.t1030 26.5955
R13927 VDD.n276 VDD.t1044 26.5955
R13928 VDD.n276 VDD.t944 26.5955
R13929 VDD.n282 VDD.t1022 26.5955
R13930 VDD.n282 VDD.t962 26.5955
R13931 VDD.n288 VDD.t1050 26.5955
R13932 VDD.n288 VDD.t984 26.5955
R13933 VDD.n292 VDD.t994 26.5955
R13934 VDD.n292 VDD.t1018 26.5955
R13935 VDD.n299 VDD.t1036 26.5955
R13936 VDD.n299 VDD.t934 26.5955
R13937 VDD.n307 VDD.t930 26.5955
R13938 VDD.n307 VDD.t956 26.5955
R13939 VDD.n223 VDD.t1479 26.5955
R13940 VDD.n223 VDD.t1493 26.5955
R13941 VDD.n229 VDD.t1491 26.5955
R13942 VDD.n229 VDD.t1475 26.5955
R13943 VDD.n235 VDD.t1473 26.5955
R13944 VDD.n235 VDD.t1485 26.5955
R13945 VDD.n241 VDD.t1483 26.5955
R13946 VDD.n241 VDD.t1497 26.5955
R13947 VDD.n245 VDD.t1495 26.5955
R13948 VDD.n245 VDD.t1471 26.5955
R13949 VDD.n251 VDD.t1489 26.5955
R13950 VDD.n251 VDD.t1499 26.5955
R13951 VDD.n259 VDD.t1469 26.5955
R13952 VDD.n259 VDD.t1481 26.5955
R13953 VDD.n604 VDD.t1076 26.5955
R13954 VDD.n604 VDD.t1078 26.5955
R13955 VDD.n471 VDD.t1446 26.5955
R13956 VDD.n471 VDD.t1378 26.5955
R13957 VDD.n477 VDD.t1352 26.5955
R13958 VDD.n477 VDD.t1416 26.5955
R13959 VDD.n483 VDD.t1432 26.5955
R13960 VDD.n483 VDD.t1456 26.5955
R13961 VDD.n489 VDD.t1454 26.5955
R13962 VDD.n489 VDD.t1364 26.5955
R13963 VDD.n494 VDD.t1356 26.5955
R13964 VDD.n494 VDD.t1384 26.5955
R13965 VDD.n450 VDD.t1344 26.5955
R13966 VDD.n450 VDD.t1464 26.5955
R13967 VDD.n445 VDD.t1366 26.5955
R13968 VDD.n445 VDD.t1452 26.5955
R13969 VDD.n529 VDD.t1450 26.5955
R13970 VDD.n529 VDD.t1382 26.5955
R13971 VDD.n523 VDD.t1376 26.5955
R13972 VDD.n523 VDD.t1402 26.5955
R13973 VDD.n517 VDD.t1362 26.5955
R13974 VDD.n517 VDD.t1444 26.5955
R13975 VDD.n511 VDD.t1394 26.5955
R13976 VDD.n511 VDD.t1428 26.5955
R13977 VDD.n507 VDD.t1424 26.5955
R13978 VDD.n507 VDD.t1358 26.5955
R13979 VDD.n441 VDD.t1462 26.5955
R13980 VDD.n441 VDD.t1390 26.5955
R13981 VDD.n461 VDD.t1410 26.5955
R13982 VDD.n461 VDD.t1436 26.5955
R13983 VDD.n428 VDD.t1346 26.5955
R13984 VDD.n428 VDD.t1368 26.5955
R13985 VDD.n556 VDD.t1374 26.5955
R13986 VDD.n556 VDD.t1400 26.5955
R13987 VDD.n562 VDD.t1398 26.5955
R13988 VDD.n562 VDD.t1430 26.5955
R13989 VDD.n568 VDD.t1442 26.5955
R13990 VDD.n568 VDD.t1372 26.5955
R13991 VDD.n573 VDD.t1350 26.5955
R13992 VDD.n573 VDD.t1414 26.5955
R13993 VDD.n547 VDD.t1354 26.5955
R13994 VDD.n547 VDD.t1440 26.5955
R13995 VDD.n541 VDD.t1388 26.5955
R13996 VDD.n541 VDD.t1418 26.5955
R13997 VDD.n660 VDD.t1380 26.5955
R13998 VDD.n660 VDD.t1404 26.5955
R13999 VDD.n666 VDD.t1420 26.5955
R14000 VDD.n666 VDD.t1448 26.5955
R14001 VDD.n672 VDD.t1396 26.5955
R14002 VDD.n672 VDD.t1338 26.5955
R14003 VDD.n678 VDD.t1426 26.5955
R14004 VDD.n678 VDD.t1360 26.5955
R14005 VDD.n682 VDD.t1370 26.5955
R14006 VDD.n682 VDD.t1392 26.5955
R14007 VDD.n689 VDD.t1412 26.5955
R14008 VDD.n689 VDD.t1438 26.5955
R14009 VDD.n697 VDD.t1434 26.5955
R14010 VDD.n697 VDD.t1460 26.5955
R14011 VDD.n613 VDD.t511 26.5955
R14012 VDD.n613 VDD.t525 26.5955
R14013 VDD.n619 VDD.t523 26.5955
R14014 VDD.n619 VDD.t507 26.5955
R14015 VDD.n625 VDD.t537 26.5955
R14016 VDD.n625 VDD.t517 26.5955
R14017 VDD.n631 VDD.t515 26.5955
R14018 VDD.n631 VDD.t529 26.5955
R14019 VDD.n635 VDD.t527 26.5955
R14020 VDD.n635 VDD.t535 26.5955
R14021 VDD.n641 VDD.t521 26.5955
R14022 VDD.n641 VDD.t531 26.5955
R14023 VDD.n649 VDD.t533 26.5955
R14024 VDD.n649 VDD.t513 26.5955
R14025 VDD.n1352 VDD.t396 26.5955
R14026 VDD.n1352 VDD.t398 26.5955
R14027 VDD.n1334 VDD.t222 26.5955
R14028 VDD.n1334 VDD.t248 26.5955
R14029 VDD.n1328 VDD.t244 26.5955
R14030 VDD.n1328 VDD.t276 26.5955
R14031 VDD.n1321 VDD.t292 26.5955
R14032 VDD.n1321 VDD.t218 26.5955
R14033 VDD.n1434 VDD.t332 26.5955
R14034 VDD.n1434 VDD.t260 26.5955
R14035 VDD.n1438 VDD.t256 26.5955
R14036 VDD.n1438 VDD.t288 26.5955
R14037 VDD.n1444 VDD.t232 26.5955
R14038 VDD.n1444 VDD.t328 26.5955
R14039 VDD.n1450 VDD.t280 26.5955
R14040 VDD.n1450 VDD.t310 26.5955
R14041 VDD.n1378 VDD.t628 26.5955
R14042 VDD.n1378 VDD.t636 26.5955
R14043 VDD.n1384 VDD.t640 26.5955
R14044 VDD.n1384 VDD.t618 26.5955
R14045 VDD.n1390 VDD.t630 26.5955
R14046 VDD.n1390 VDD.t626 26.5955
R14047 VDD.n1402 VDD.t614 26.5955
R14048 VDD.n1402 VDD.t620 26.5955
R14049 VDD.n1407 VDD.t624 26.5955
R14050 VDD.n1407 VDD.t634 26.5955
R14051 VDD.n1413 VDD.t632 26.5955
R14052 VDD.n1413 VDD.t642 26.5955
R14053 VDD.n1419 VDD.t644 26.5955
R14054 VDD.n1419 VDD.t622 26.5955
R14055 VDD.n1305 VDD.t224 26.5955
R14056 VDD.n1305 VDD.t250 26.5955
R14057 VDD.n1298 VDD.t266 26.5955
R14058 VDD.n1298 VDD.t298 26.5955
R14059 VDD.n1292 VDD.t240 26.5955
R14060 VDD.n1292 VDD.t206 26.5955
R14061 VDD.n1267 VDD.t272 26.5955
R14062 VDD.n1267 VDD.t208 26.5955
R14063 VDD.n1271 VDD.t314 26.5955
R14064 VDD.n1271 VDD.t236 26.5955
R14065 VDD.n1277 VDD.t254 26.5955
R14066 VDD.n1277 VDD.t286 26.5955
R14067 VDD.n1264 VDD.t282 26.5955
R14068 VDD.n1264 VDD.t324 26.5955
R14069 VDD.n1464 VDD.t278 26.5955
R14070 VDD.n1464 VDD.t214 26.5955
R14071 VDD.n1470 VDD.t220 26.5955
R14072 VDD.n1470 VDD.t246 26.5955
R14073 VDD.n1476 VDD.t242 26.5955
R14074 VDD.n1476 VDD.t294 26.5955
R14075 VDD.n1482 VDD.t290 26.5955
R14076 VDD.n1482 VDD.t318 26.5955
R14077 VDD.n1486 VDD.t330 26.5955
R14078 VDD.n1486 VDD.t258 26.5955
R14079 VDD.n1492 VDD.t216 26.5955
R14080 VDD.n1492 VDD.t306 26.5955
R14081 VDD.n1498 VDD.t230 26.5955
R14082 VDD.n1498 VDD.t264 26.5955
R14083 VDD.n1514 VDD.t300 26.5955
R14084 VDD.n1514 VDD.t226 26.5955
R14085 VDD.n1520 VDD.t320 26.5955
R14086 VDD.n1520 VDD.t268 26.5955
R14087 VDD.n1256 VDD.t262 26.5955
R14088 VDD.n1256 VDD.t296 26.5955
R14089 VDD.n1530 VDD.t238 26.5955
R14090 VDD.n1530 VDD.t274 26.5955
R14091 VDD.n1534 VDD.t270 26.5955
R14092 VDD.n1534 VDD.t316 26.5955
R14093 VDD.n1252 VDD.t312 26.5955
R14094 VDD.n1252 VDD.t234 26.5955
R14095 VDD.n1247 VDD.t212 26.5955
R14096 VDD.n1247 VDD.t284 26.5955
R14097 VDD.n1129 VDD.n1128 25.977
R14098 VDD.n1195 VDD.n1194 25.977
R14099 VDD.t1206 VDD.t1318 25.9096
R14100 VDD.t661 VDD.t370 25.9096
R14101 VDD.n989 VDD.t1135 25.6105
R14102 VDD.n194 VDD.t1058 25.6105
R14103 VDD.n584 VDD.t1305 25.6105
R14104 VDD.n1136 VDD.n1135 25.224
R14105 VDD.n1202 VDD.n1201 25.224
R14106 VDD.t355 VDD.n1847 24.3893
R14107 VDD.t574 VDD.n2168 24.3893
R14108 VDD.t103 VDD.n2426 24.3893
R14109 VDD.t421 VDD.n2684 24.3893
R14110 VDD.t405 VDD.n2942 24.3893
R14111 VDD.t144 VDD.n3200 24.3893
R14112 VDD.t179 VDD.n3458 24.3893
R14113 VDD.t1088 VDD.n5785 24.3893
R14114 VDD.t596 VDD.n5531 24.3893
R14115 VDD.t145 VDD.n3716 24.3893
R14116 VDD.t563 VDD.n3974 24.3893
R14117 VDD.t668 VDD.n4232 24.3893
R14118 VDD.t561 VDD.n4490 24.3893
R14119 VDD.t750 VDD.n4748 24.3893
R14120 VDD.t386 VDD.n5009 24.3893
R14121 VDD.t559 VDD.n5271 24.3893
R14122 VDD.t163 VDD.t1204 23.0308
R14123 VDD.t747 VDD.t657 23.0308
R14124 VDD.n725 VDD 22.7027
R14125 VDD.n1566 VDD 22.7027
R14126 VDD.n1660 VDD.n1626 22.5125
R14127 VDD.n1834 VDD.n1833 22.2123
R14128 VDD.n1814 VDD.n1812 22.2123
R14129 VDD.n1784 VDD.n1782 22.2123
R14130 VDD.n1795 VDD.n1794 22.2123
R14131 VDD.n1787 VDD.n1786 22.2123
R14132 VDD.n1789 VDD.n1781 22.2123
R14133 VDD.n2135 VDD.n2133 22.2123
R14134 VDD.n2155 VDD.n2154 22.2123
R14135 VDD.n1992 VDD.n1990 22.2123
R14136 VDD.n2003 VDD.n2002 22.2123
R14137 VDD.n1995 VDD.n1994 22.2123
R14138 VDD.n1997 VDD.n1989 22.2123
R14139 VDD.n2393 VDD.n2391 22.2123
R14140 VDD.n2413 VDD.n2412 22.2123
R14141 VDD.n2363 VDD.n2361 22.2123
R14142 VDD.n2374 VDD.n2373 22.2123
R14143 VDD.n2366 VDD.n2365 22.2123
R14144 VDD.n2368 VDD.n2360 22.2123
R14145 VDD.n2651 VDD.n2649 22.2123
R14146 VDD.n2671 VDD.n2670 22.2123
R14147 VDD.n2621 VDD.n2619 22.2123
R14148 VDD.n2632 VDD.n2631 22.2123
R14149 VDD.n2624 VDD.n2623 22.2123
R14150 VDD.n2626 VDD.n2618 22.2123
R14151 VDD.n2909 VDD.n2907 22.2123
R14152 VDD.n2929 VDD.n2928 22.2123
R14153 VDD.n2879 VDD.n2877 22.2123
R14154 VDD.n2890 VDD.n2889 22.2123
R14155 VDD.n2882 VDD.n2881 22.2123
R14156 VDD.n2884 VDD.n2876 22.2123
R14157 VDD.n3167 VDD.n3165 22.2123
R14158 VDD.n3187 VDD.n3186 22.2123
R14159 VDD.n3137 VDD.n3135 22.2123
R14160 VDD.n3148 VDD.n3147 22.2123
R14161 VDD.n3140 VDD.n3139 22.2123
R14162 VDD.n3142 VDD.n3134 22.2123
R14163 VDD.n3425 VDD.n3423 22.2123
R14164 VDD.n3445 VDD.n3444 22.2123
R14165 VDD.n3395 VDD.n3393 22.2123
R14166 VDD.n3406 VDD.n3405 22.2123
R14167 VDD.n3398 VDD.n3397 22.2123
R14168 VDD.n3400 VDD.n3392 22.2123
R14169 VDD.n5752 VDD.n5750 22.2123
R14170 VDD.n5772 VDD.n5771 22.2123
R14171 VDD.n5725 VDD.n5723 22.2123
R14172 VDD.n5736 VDD.n5735 22.2123
R14173 VDD.n5728 VDD.n5727 22.2123
R14174 VDD.n5730 VDD.n5722 22.2123
R14175 VDD.n5498 VDD.n5496 22.2123
R14176 VDD.n5518 VDD.n5517 22.2123
R14177 VDD.n5471 VDD.n5469 22.2123
R14178 VDD.n5482 VDD.n5481 22.2123
R14179 VDD.n5474 VDD.n5473 22.2123
R14180 VDD.n5476 VDD.n5468 22.2123
R14181 VDD.n3683 VDD.n3681 22.2123
R14182 VDD.n3703 VDD.n3702 22.2123
R14183 VDD.n3653 VDD.n3651 22.2123
R14184 VDD.n3664 VDD.n3663 22.2123
R14185 VDD.n3656 VDD.n3655 22.2123
R14186 VDD.n3658 VDD.n3650 22.2123
R14187 VDD.n3941 VDD.n3939 22.2123
R14188 VDD.n3961 VDD.n3960 22.2123
R14189 VDD.n3911 VDD.n3909 22.2123
R14190 VDD.n3922 VDD.n3921 22.2123
R14191 VDD.n3914 VDD.n3913 22.2123
R14192 VDD.n3916 VDD.n3908 22.2123
R14193 VDD.n4199 VDD.n4197 22.2123
R14194 VDD.n4219 VDD.n4218 22.2123
R14195 VDD.n4169 VDD.n4167 22.2123
R14196 VDD.n4180 VDD.n4179 22.2123
R14197 VDD.n4172 VDD.n4171 22.2123
R14198 VDD.n4174 VDD.n4166 22.2123
R14199 VDD.n4457 VDD.n4455 22.2123
R14200 VDD.n4477 VDD.n4476 22.2123
R14201 VDD.n4427 VDD.n4425 22.2123
R14202 VDD.n4438 VDD.n4437 22.2123
R14203 VDD.n4430 VDD.n4429 22.2123
R14204 VDD.n4432 VDD.n4424 22.2123
R14205 VDD.n4715 VDD.n4713 22.2123
R14206 VDD.n4735 VDD.n4734 22.2123
R14207 VDD.n4685 VDD.n4683 22.2123
R14208 VDD.n4696 VDD.n4695 22.2123
R14209 VDD.n4688 VDD.n4687 22.2123
R14210 VDD.n4690 VDD.n4682 22.2123
R14211 VDD.n4944 VDD.n4942 22.2123
R14212 VDD.n4955 VDD.n4954 22.2123
R14213 VDD.n4947 VDD.n4946 22.2123
R14214 VDD.n4949 VDD.n4941 22.2123
R14215 VDD.n4996 VDD.n4995 22.2123
R14216 VDD.n4976 VDD.n4974 22.2123
R14217 VDD.n5094 VDD.n5092 22.2123
R14218 VDD.n5105 VDD.n5104 22.2123
R14219 VDD.n5097 VDD.n5096 22.2123
R14220 VDD.n5099 VDD.n5091 22.2123
R14221 VDD.n5258 VDD.n5257 22.2123
R14222 VDD.n5238 VDD.n5236 22.2123
R14223 VDD.n1130 VDD.n1129 22.2123
R14224 VDD.n1196 VDD.n1195 22.2123
R14225 VDD.n1804 VDD.t1224 20.9587
R14226 VDD.n2012 VDD.t31 20.9587
R14227 VDD.n2383 VDD.t538 20.9587
R14228 VDD.n2641 VDD.t474 20.9587
R14229 VDD.n2899 VDD.t1306 20.9587
R14230 VDD.n3157 VDD.t8 20.9587
R14231 VDD.n3415 VDD.t1196 20.9587
R14232 VDD.n5745 VDD.t704 20.9587
R14233 VDD.n5491 VDD.t1329 20.9587
R14234 VDD.n3673 VDD.t1270 20.9587
R14235 VDD.n3931 VDD.t78 20.9587
R14236 VDD.n4189 VDD.t720 20.9587
R14237 VDD.n4447 VDD.t1109 20.9587
R14238 VDD.n4705 VDD.t185 20.9587
R14239 VDD.n4964 VDD.t1123 20.9587
R14240 VDD.n5114 VDD.t192 20.9587
R14241 VDD.n1507 VDD 20.8224
R14242 VDD.n1457 VDD 20.8224
R14243 VDD.n1707 VDD.n1705 20.5934
R14244 VDD.n2056 VDD.n2054 20.5934
R14245 VDD.n2286 VDD.n2284 20.5934
R14246 VDD.n2544 VDD.n2542 20.5934
R14247 VDD.n2802 VDD.n2800 20.5934
R14248 VDD.n3060 VDD.n3058 20.5934
R14249 VDD.n3318 VDD.n3316 20.5934
R14250 VDD.n5648 VDD.n5646 20.5934
R14251 VDD.n5394 VDD.n5392 20.5934
R14252 VDD.n3576 VDD.n3574 20.5934
R14253 VDD.n3834 VDD.n3832 20.5934
R14254 VDD.n4092 VDD.n4090 20.5934
R14255 VDD.n4350 VDD.n4348 20.5934
R14256 VDD.n4608 VDD.n4606 20.5934
R14257 VDD.n4866 VDD.n4864 20.5934
R14258 VDD.n5158 VDD.n5156 20.5934
R14259 VDD.n13 VDD.n12 19.9534
R14260 VDD.n330 VDD.n329 19.9534
R14261 VDD.n1840 VDD.n1839 18.6543
R14262 VDD.n2161 VDD.n2160 18.6543
R14263 VDD.n2419 VDD.n2418 18.6543
R14264 VDD.n2677 VDD.n2676 18.6543
R14265 VDD.n2935 VDD.n2934 18.6543
R14266 VDD.n3193 VDD.n3192 18.6543
R14267 VDD.n3451 VDD.n3450 18.6543
R14268 VDD.n5778 VDD.n5777 18.6543
R14269 VDD.n5524 VDD.n5523 18.6543
R14270 VDD.n3709 VDD.n3708 18.6543
R14271 VDD.n3967 VDD.n3966 18.6543
R14272 VDD.n4225 VDD.n4224 18.6543
R14273 VDD.n4483 VDD.n4482 18.6543
R14274 VDD.n4741 VDD.n4740 18.6543
R14275 VDD.n5002 VDD.n5001 18.6543
R14276 VDD.n5264 VDD.n5263 18.6543
R14277 VDD.n1372 VDD.t615 18.2197
R14278 VDD.n1654 VDD 17.4176
R14279 VDD.n1761 VDD.n1716 17.109
R14280 VDD.n2110 VDD.n2065 17.109
R14281 VDD.n2340 VDD.n2295 17.109
R14282 VDD.n2598 VDD.n2553 17.109
R14283 VDD.n2856 VDD.n2811 17.109
R14284 VDD.n3114 VDD.n3069 17.109
R14285 VDD.n3372 VDD.n3327 17.109
R14286 VDD.n5702 VDD.n5657 17.109
R14287 VDD.n5448 VDD.n5403 17.109
R14288 VDD.n3630 VDD.n3585 17.109
R14289 VDD.n3888 VDD.n3843 17.109
R14290 VDD.n4146 VDD.n4101 17.109
R14291 VDD.n4404 VDD.n4359 17.109
R14292 VDD.n4662 VDD.n4617 17.109
R14293 VDD.n4920 VDD.n4875 17.109
R14294 VDD.n5212 VDD.n5167 17.109
R14295 VDD.n24 VDD.n23 16.9417
R14296 VDD.n892 VDD.n891 16.9417
R14297 VDD.n914 VDD.n913 16.9417
R14298 VDD.n975 VDD.n974 16.9417
R14299 VDD.n1085 VDD.n1084 16.9417
R14300 VDD.n1038 VDD.n1037 16.9417
R14301 VDD.n805 VDD.n804 16.9417
R14302 VDD.n403 VDD.n402 16.9417
R14303 VDD.n341 VDD.n340 16.9417
R14304 VDD.n97 VDD.n96 16.9417
R14305 VDD.n119 VDD.n118 16.9417
R14306 VDD.n180 VDD.n179 16.9417
R14307 VDD.n290 VDD.n289 16.9417
R14308 VDD.n243 VDD.n242 16.9417
R14309 VDD.n491 VDD.n490 16.9417
R14310 VDD.n513 VDD.n512 16.9417
R14311 VDD.n570 VDD.n569 16.9417
R14312 VDD.n680 VDD.n679 16.9417
R14313 VDD.n633 VDD.n632 16.9417
R14314 VDD.n1436 VDD.n1435 16.9417
R14315 VDD.n1404 VDD.n1403 16.9417
R14316 VDD.n1269 VDD.n1268 16.9417
R14317 VDD.n1484 VDD.n1483 16.9417
R14318 VDD.n1532 VDD.n1531 16.9417
R14319 VDD.n8 VDD.n2 16.1887
R14320 VDD.n325 VDD.n319 16.1887
R14321 VDD.n1005 VDD.n1004 14.5711
R14322 VDD.n210 VDD.n209 14.5711
R14323 VDD.n600 VDD.n599 14.5711
R14324 VDD.n1659 VDD 14.551
R14325 VDD.n1686 VDD.t1228 14.2962
R14326 VDD.n2035 VDD.t36 14.2962
R14327 VDD.n2265 VDD.t542 14.2962
R14328 VDD.n2523 VDD.t473 14.2962
R14329 VDD.n2781 VDD.t1313 14.2962
R14330 VDD.n3039 VDD.t7 14.2962
R14331 VDD.n3297 VDD.t1195 14.2962
R14332 VDD.n5627 VDD.t710 14.2962
R14333 VDD.n5373 VDD.t1332 14.2962
R14334 VDD.n3555 VDD.t1269 14.2962
R14335 VDD.n3813 VDD.t82 14.2962
R14336 VDD.n4071 VDD.t724 14.2962
R14337 VDD.n4329 VDD.t1116 14.2962
R14338 VDD.n4587 VDD.t188 14.2962
R14339 VDD.n4845 VDD.t1122 14.2962
R14340 VDD.n5137 VDD.t199 14.2962
R14341 VDD.n1666 VDD.t1229 14.2955
R14342 VDD.n2015 VDD.t30 14.2955
R14343 VDD.n2245 VDD.t545 14.2955
R14344 VDD.n2503 VDD.t477 14.2955
R14345 VDD.n2761 VDD.t1310 14.2955
R14346 VDD.n3019 VDD.t11 14.2955
R14347 VDD.n3277 VDD.t1199 14.2955
R14348 VDD.n5607 VDD.t708 14.2955
R14349 VDD.n5353 VDD.t1335 14.2955
R14350 VDD.n3535 VDD.t1273 14.2955
R14351 VDD.n3793 VDD.t85 14.2955
R14352 VDD.n4051 VDD.t727 14.2955
R14353 VDD.n4309 VDD.t1113 14.2955
R14354 VDD.n4567 VDD.t184 14.2955
R14355 VDD.n4825 VDD.t1126 14.2955
R14356 VDD.n5117 VDD.t196 14.2955
R14357 VDD.n1749 VDD.t44 14.2865
R14358 VDD.n2098 VDD.t366 14.2865
R14359 VDD.n2328 VDD.t467 14.2865
R14360 VDD.n2586 VDD.t124 14.2865
R14361 VDD.n2844 VDD.t22 14.2865
R14362 VDD.n3102 VDD.t591 14.2865
R14363 VDD.n3360 VDD.t551 14.2865
R14364 VDD.n5690 VDD.t171 14.2865
R14365 VDD.n5436 VDD.t763 14.2865
R14366 VDD.n3618 VDD.t1101 14.2865
R14367 VDD.n3876 VDD.t790 14.2865
R14368 VDD.n4134 VDD.t496 14.2865
R14369 VDD.n4392 VDD.t375 14.2865
R14370 VDD.n4650 VDD.t112 14.2865
R14371 VDD.n4908 VDD.t350 14.2865
R14372 VDD.n5200 VDD.t483 14.2865
R14373 VDD.n1737 VDD.t38 14.2864
R14374 VDD.n2086 VDD.t367 14.2864
R14375 VDD.n2316 VDD.t469 14.2864
R14376 VDD.n2574 VDD.t118 14.2864
R14377 VDD.n2832 VDD.t24 14.2864
R14378 VDD.n3090 VDD.t593 14.2864
R14379 VDD.n3348 VDD.t553 14.2864
R14380 VDD.n5678 VDD.t173 14.2864
R14381 VDD.n5424 VDD.t758 14.2864
R14382 VDD.n3606 VDD.t1103 14.2864
R14383 VDD.n3864 VDD.t786 14.2864
R14384 VDD.n4122 VDD.t491 14.2864
R14385 VDD.n4380 VDD.t377 14.2864
R14386 VDD.n4638 VDD.t114 14.2864
R14387 VDD.n4896 VDD.t352 14.2864
R14388 VDD.n5188 VDD.t485 14.2864
R14389 VDD.n1771 VDD.t754 14.2849
R14390 VDD.n1753 VDD.t773 14.2849
R14391 VDD.n2120 VDD.t130 14.2849
R14392 VDD.n2102 VDD.t498 14.2849
R14393 VDD.n2350 VDD.t71 14.2849
R14394 VDD.n2332 VDD.t416 14.2849
R14395 VDD.n2608 VDD.t1094 14.2849
R14396 VDD.n2590 VDD.t681 14.2849
R14397 VDD.n2866 VDD.t749 14.2849
R14398 VDD.n2848 VDD.t734 14.2849
R14399 VDD.n3124 VDD.t126 14.2849
R14400 VDD.n3106 VDD.t503 14.2849
R14401 VDD.n3382 VDD.t505 14.2849
R14402 VDD.n3364 VDD.t600 14.2849
R14403 VDD.n5712 VDD.t5 14.2849
R14404 VDD.n5694 VDD.t601 14.2849
R14405 VDD.n5458 VDD.t1067 14.2849
R14406 VDD.n5440 VDD.t666 14.2849
R14407 VDD.n3640 VDD.t1142 14.2849
R14408 VDD.n3622 VDD.t1143 14.2849
R14409 VDD.n3898 VDD.t1062 14.2849
R14410 VDD.n3880 VDD.t1129 14.2849
R14411 VDD.n4156 VDD.t415 14.2849
R14412 VDD.n4138 VDD.t1146 14.2849
R14413 VDD.n4414 VDD.t166 14.2849
R14414 VDD.n4396 VDD.t1072 14.2849
R14415 VDD.n4672 VDD.t794 14.2849
R14416 VDD.n4654 VDD.t1263 14.2849
R14417 VDD.n4930 VDD.t1215 14.2849
R14418 VDD.n4912 VDD.t1066 14.2849
R14419 VDD.n5222 VDD.t1068 14.2849
R14420 VDD.n5204 VDD.t108 14.2849
R14421 VDD.n1620 VDD.n1619 14.1868
R14422 VDD.n1769 VDD.n1669 14.0805
R14423 VDD.n2118 VDD.n2018 14.0805
R14424 VDD.n2348 VDD.n2248 14.0805
R14425 VDD.n2606 VDD.n2506 14.0805
R14426 VDD.n2864 VDD.n2764 14.0805
R14427 VDD.n3122 VDD.n3022 14.0805
R14428 VDD.n3380 VDD.n3280 14.0805
R14429 VDD.n5710 VDD.n5610 14.0805
R14430 VDD.n5456 VDD.n5356 14.0805
R14431 VDD.n3638 VDD.n3538 14.0805
R14432 VDD.n3896 VDD.n3796 14.0805
R14433 VDD.n4154 VDD.n4054 14.0805
R14434 VDD.n4412 VDD.n4312 14.0805
R14435 VDD.n4670 VDD.n4570 14.0805
R14436 VDD.n4928 VDD.n4828 14.0805
R14437 VDD.n5220 VDD.n5120 14.0805
R14438 VDD.t698 VDD.t45 13.9711
R14439 VDD.t459 VDD.t1250 13.9711
R14440 VDD.t72 VDD.t52 13.9711
R14441 VDD.t1163 VDD.t345 13.9711
R14442 VDD.n1755 VDD.n1717 13.7605
R14443 VDD.n2104 VDD.n2066 13.7605
R14444 VDD.n2334 VDD.n2296 13.7605
R14445 VDD.n2592 VDD.n2554 13.7605
R14446 VDD.n2850 VDD.n2812 13.7605
R14447 VDD.n3108 VDD.n3070 13.7605
R14448 VDD.n3366 VDD.n3328 13.7605
R14449 VDD.n5696 VDD.n5658 13.7605
R14450 VDD.n5442 VDD.n5404 13.7605
R14451 VDD.n3624 VDD.n3586 13.7605
R14452 VDD.n3882 VDD.n3844 13.7605
R14453 VDD.n4140 VDD.n4102 13.7605
R14454 VDD.n4398 VDD.n4360 13.7605
R14455 VDD.n4656 VDD.n4618 13.7605
R14456 VDD.n4914 VDD.n4876 13.7605
R14457 VDD.n5206 VDD.n5168 13.7605
R14458 VDD.n1658 VDD.n1631 13.4428
R14459 VDD.n1657 VDD 13.4235
R14460 VDD.n1124 VDD.n1122 13.3488
R14461 VDD.n1190 VDD.n1188 13.3488
R14462 VDD.n1144 VDD.n1143 12.9329
R14463 VDD.n1543 VDD.n1542 12.9329
R14464 VDD.n1363 VDD.n1362 12.9329
R14465 VDD.n1210 VDD.n1209 12.9329
R14466 VDD.n897 VDD.n896 11.6711
R14467 VDD.n910 VDD.n909 11.6711
R14468 VDD.n980 VDD.n979 11.6711
R14469 VDD.n1089 VDD.n1088 11.6711
R14470 VDD.n1042 VDD.n1041 11.6711
R14471 VDD.n102 VDD.n101 11.6711
R14472 VDD.n115 VDD.n114 11.6711
R14473 VDD.n185 VDD.n184 11.6711
R14474 VDD.n294 VDD.n293 11.6711
R14475 VDD.n247 VDD.n246 11.6711
R14476 VDD.n496 VDD.n495 11.6711
R14477 VDD.n509 VDD.n508 11.6711
R14478 VDD.n575 VDD.n574 11.6711
R14479 VDD.n684 VDD.n683 11.6711
R14480 VDD.n637 VDD.n636 11.6711
R14481 VDD.n1440 VDD.n1439 11.6711
R14482 VDD.n1409 VDD.n1408 11.6711
R14483 VDD.n1273 VDD.n1272 11.6711
R14484 VDD.n1488 VDD.n1487 11.6711
R14485 VDD.n1536 VDD.n1535 11.6711
R14486 VDD.n886 VDD.n885 10.9181
R14487 VDD.n920 VDD.n919 10.9181
R14488 VDD.n969 VDD.n968 10.9181
R14489 VDD.n1079 VDD.n1078 10.9181
R14490 VDD.n1032 VDD.n1031 10.9181
R14491 VDD.n91 VDD.n90 10.9181
R14492 VDD.n125 VDD.n124 10.9181
R14493 VDD.n174 VDD.n173 10.9181
R14494 VDD.n284 VDD.n283 10.9181
R14495 VDD.n237 VDD.n236 10.9181
R14496 VDD.n485 VDD.n484 10.9181
R14497 VDD.n519 VDD.n518 10.9181
R14498 VDD.n564 VDD.n563 10.9181
R14499 VDD.n674 VDD.n673 10.9181
R14500 VDD.n627 VDD.n626 10.9181
R14501 VDD.n1323 VDD.n1322 10.9181
R14502 VDD.n1392 VDD.n1391 10.9181
R14503 VDD.n1294 VDD.n1293 10.9181
R14504 VDD.n1478 VDD.n1477 10.9181
R14505 VDD.n1258 VDD.n1257 10.9181
R14506 VDD.n1957 VDD.n1956 10.8802
R14507 VDD.n780 VDD 10.8576
R14508 VDD.n377 VDD 10.8576
R14509 VDD.n1955 VDD.n1954 10.5887
R14510 VDD.n1429 VDD.t291 10.4115
R14511 VDD.n985 VDD.t885 10.1791
R14512 VDD.n190 VDD.t1035 10.1791
R14513 VDD.t512 VDD.n581 10.1791
R14514 VDD.n1617 VDD 9.58775
R14515 VDD.n9 VDD.n6 9.41227
R14516 VDD.n326 VDD.n323 9.41227
R14517 VDD.n1954 VDD.n1953 9.3005
R14518 VDD.n1916 VDD.n1915 9.3005
R14519 VDD.n1915 VDD.n1914 9.3005
R14520 VDD.n1828 VDD.n1826 9.3005
R14521 VDD.n1747 VDD.n1746 9.3005
R14522 VDD.n1728 VDD.n1727 9.3005
R14523 VDD.n1731 VDD.n1722 9.3005
R14524 VDD.n1705 VDD.n1667 9.3005
R14525 VDD.n1690 VDD.n1689 9.3005
R14526 VDD.n2096 VDD.n2095 9.3005
R14527 VDD.n2077 VDD.n2076 9.3005
R14528 VDD.n2080 VDD.n2071 9.3005
R14529 VDD.n2054 VDD.n2016 9.3005
R14530 VDD.n2039 VDD.n2038 9.3005
R14531 VDD.n2237 VDD.n2236 9.3005
R14532 VDD.n2236 VDD.n2235 9.3005
R14533 VDD.n2149 VDD.n2147 9.3005
R14534 VDD.n2326 VDD.n2325 9.3005
R14535 VDD.n2307 VDD.n2306 9.3005
R14536 VDD.n2310 VDD.n2301 9.3005
R14537 VDD.n2284 VDD.n2246 9.3005
R14538 VDD.n2269 VDD.n2268 9.3005
R14539 VDD.n2495 VDD.n2494 9.3005
R14540 VDD.n2494 VDD.n2493 9.3005
R14541 VDD.n2407 VDD.n2405 9.3005
R14542 VDD.n2584 VDD.n2583 9.3005
R14543 VDD.n2565 VDD.n2564 9.3005
R14544 VDD.n2568 VDD.n2559 9.3005
R14545 VDD.n2542 VDD.n2504 9.3005
R14546 VDD.n2527 VDD.n2526 9.3005
R14547 VDD.n2753 VDD.n2752 9.3005
R14548 VDD.n2752 VDD.n2751 9.3005
R14549 VDD.n2665 VDD.n2663 9.3005
R14550 VDD.n2842 VDD.n2841 9.3005
R14551 VDD.n2823 VDD.n2822 9.3005
R14552 VDD.n2826 VDD.n2817 9.3005
R14553 VDD.n2800 VDD.n2762 9.3005
R14554 VDD.n2785 VDD.n2784 9.3005
R14555 VDD.n3011 VDD.n3010 9.3005
R14556 VDD.n3010 VDD.n3009 9.3005
R14557 VDD.n2923 VDD.n2921 9.3005
R14558 VDD.n3100 VDD.n3099 9.3005
R14559 VDD.n3081 VDD.n3080 9.3005
R14560 VDD.n3084 VDD.n3075 9.3005
R14561 VDD.n3058 VDD.n3020 9.3005
R14562 VDD.n3043 VDD.n3042 9.3005
R14563 VDD.n3269 VDD.n3268 9.3005
R14564 VDD.n3268 VDD.n3267 9.3005
R14565 VDD.n3181 VDD.n3179 9.3005
R14566 VDD.n3358 VDD.n3357 9.3005
R14567 VDD.n3339 VDD.n3338 9.3005
R14568 VDD.n3342 VDD.n3333 9.3005
R14569 VDD.n3316 VDD.n3278 9.3005
R14570 VDD.n3301 VDD.n3300 9.3005
R14571 VDD.n3527 VDD.n3526 9.3005
R14572 VDD.n3526 VDD.n3525 9.3005
R14573 VDD.n3439 VDD.n3437 9.3005
R14574 VDD.n5688 VDD.n5687 9.3005
R14575 VDD.n5669 VDD.n5668 9.3005
R14576 VDD.n5672 VDD.n5663 9.3005
R14577 VDD.n5646 VDD.n5608 9.3005
R14578 VDD.n5631 VDD.n5630 9.3005
R14579 VDD.n5854 VDD.n5853 9.3005
R14580 VDD.n5853 VDD.n5852 9.3005
R14581 VDD.n5766 VDD.n5764 9.3005
R14582 VDD.n5434 VDD.n5433 9.3005
R14583 VDD.n5415 VDD.n5414 9.3005
R14584 VDD.n5418 VDD.n5409 9.3005
R14585 VDD.n5392 VDD.n5354 9.3005
R14586 VDD.n5377 VDD.n5376 9.3005
R14587 VDD.n5600 VDD.n5599 9.3005
R14588 VDD.n5599 VDD.n5598 9.3005
R14589 VDD.n5512 VDD.n5510 9.3005
R14590 VDD.n3616 VDD.n3615 9.3005
R14591 VDD.n3597 VDD.n3596 9.3005
R14592 VDD.n3600 VDD.n3591 9.3005
R14593 VDD.n3574 VDD.n3536 9.3005
R14594 VDD.n3559 VDD.n3558 9.3005
R14595 VDD.n3785 VDD.n3784 9.3005
R14596 VDD.n3784 VDD.n3783 9.3005
R14597 VDD.n3697 VDD.n3695 9.3005
R14598 VDD.n3874 VDD.n3873 9.3005
R14599 VDD.n3855 VDD.n3854 9.3005
R14600 VDD.n3858 VDD.n3849 9.3005
R14601 VDD.n3832 VDD.n3794 9.3005
R14602 VDD.n3817 VDD.n3816 9.3005
R14603 VDD.n4043 VDD.n4042 9.3005
R14604 VDD.n4042 VDD.n4041 9.3005
R14605 VDD.n3955 VDD.n3953 9.3005
R14606 VDD.n4132 VDD.n4131 9.3005
R14607 VDD.n4113 VDD.n4112 9.3005
R14608 VDD.n4116 VDD.n4107 9.3005
R14609 VDD.n4090 VDD.n4052 9.3005
R14610 VDD.n4075 VDD.n4074 9.3005
R14611 VDD.n4301 VDD.n4300 9.3005
R14612 VDD.n4300 VDD.n4299 9.3005
R14613 VDD.n4213 VDD.n4211 9.3005
R14614 VDD.n4390 VDD.n4389 9.3005
R14615 VDD.n4371 VDD.n4370 9.3005
R14616 VDD.n4374 VDD.n4365 9.3005
R14617 VDD.n4348 VDD.n4310 9.3005
R14618 VDD.n4333 VDD.n4332 9.3005
R14619 VDD.n4559 VDD.n4558 9.3005
R14620 VDD.n4558 VDD.n4557 9.3005
R14621 VDD.n4471 VDD.n4469 9.3005
R14622 VDD.n4648 VDD.n4647 9.3005
R14623 VDD.n4629 VDD.n4628 9.3005
R14624 VDD.n4632 VDD.n4623 9.3005
R14625 VDD.n4606 VDD.n4568 9.3005
R14626 VDD.n4591 VDD.n4590 9.3005
R14627 VDD.n4817 VDD.n4816 9.3005
R14628 VDD.n4816 VDD.n4815 9.3005
R14629 VDD.n4729 VDD.n4727 9.3005
R14630 VDD.n4906 VDD.n4905 9.3005
R14631 VDD.n4887 VDD.n4886 9.3005
R14632 VDD.n4890 VDD.n4881 9.3005
R14633 VDD.n4864 VDD.n4826 9.3005
R14634 VDD.n4849 VDD.n4848 9.3005
R14635 VDD.n5078 VDD.n5077 9.3005
R14636 VDD.n5077 VDD.n5076 9.3005
R14637 VDD.n4990 VDD.n4988 9.3005
R14638 VDD.n5198 VDD.n5197 9.3005
R14639 VDD.n5179 VDD.n5178 9.3005
R14640 VDD.n5182 VDD.n5173 9.3005
R14641 VDD.n5156 VDD.n5118 9.3005
R14642 VDD.n5141 VDD.n5140 9.3005
R14643 VDD.n5340 VDD.n5339 9.3005
R14644 VDD.n5339 VDD.n5338 9.3005
R14645 VDD.n5252 VDD.n5250 9.3005
R14646 VDD.n1618 VDD.n1617 9.3005
R14647 VDD VDD.n1628 9.22489
R14648 VDD.n1646 VDD.n1645 9.0245
R14649 VDD.n1734 VDD.n1733 8.88939
R14650 VDD.n2083 VDD.n2082 8.88939
R14651 VDD.n2313 VDD.n2312 8.88939
R14652 VDD.n2571 VDD.n2570 8.88939
R14653 VDD.n2829 VDD.n2828 8.88939
R14654 VDD.n3087 VDD.n3086 8.88939
R14655 VDD.n3345 VDD.n3344 8.88939
R14656 VDD.n5675 VDD.n5674 8.88939
R14657 VDD.n5421 VDD.n5420 8.88939
R14658 VDD.n3603 VDD.n3602 8.88939
R14659 VDD.n3861 VDD.n3860 8.88939
R14660 VDD.n4119 VDD.n4118 8.88939
R14661 VDD.n4377 VDD.n4376 8.88939
R14662 VDD.n4635 VDD.n4634 8.88939
R14663 VDD.n4893 VDD.n4892 8.88939
R14664 VDD.n5185 VDD.n5184 8.88939
R14665 VDD.n1954 VDD.n1943 8.85536
R14666 VDD.n10 VDD.n9 8.79168
R14667 VDD.n730 VDD.n729 8.79168
R14668 VDD.n730 VDD.n728 8.79168
R14669 VDD.n711 VDD.n710 8.79168
R14670 VDD.n327 VDD.n326 8.79168
R14671 VDD.n1571 VDD.n1570 8.79168
R14672 VDD.n1571 VDD.n1569 8.79168
R14673 VDD.n1552 VDD.n1551 8.79168
R14674 VDD.n1652 VDD.n1649 8.76429
R14675 VDD.n5083 VDD.n4935 8.39231
R14676 VDD.n996 VDD.n988 8.28285
R14677 VDD.n1149 VDD.n1142 8.28285
R14678 VDD.n1155 VDD.n1141 8.28285
R14679 VDD.n1161 VDD.n1140 8.28285
R14680 VDD.n1167 VDD.n1139 8.28285
R14681 VDD.n201 VDD.n193 8.28285
R14682 VDD.n591 VDD.n583 8.28285
R14683 VDD.n1215 VDD.n1208 8.28285
R14684 VDD.n1221 VDD.n1207 8.28285
R14685 VDD.n1227 VDD.n1206 8.28285
R14686 VDD.n1233 VDD.n1205 8.28285
R14687 VDD.n1977 VDD.n1923 7.681
R14688 VDD.n1628 VDD 7.6805
R14689 VDD.n1618 VDD.n1616 7.60183
R14690 VDD.n741 VDD.n740 7.54105
R14691 VDD.n720 VDD.n719 7.54105
R14692 VDD.n1582 VDD.n1581 7.54105
R14693 VDD.n1561 VDD.n1560 7.54105
R14694 VDD.n1885 VDD.n1818 7.49764
R14695 VDD.n2206 VDD.n2139 7.49764
R14696 VDD.n2464 VDD.n2397 7.49764
R14697 VDD.n2722 VDD.n2655 7.49764
R14698 VDD.n2980 VDD.n2913 7.49764
R14699 VDD.n3238 VDD.n3171 7.49764
R14700 VDD.n3496 VDD.n3429 7.49764
R14701 VDD.n5823 VDD.n5756 7.49764
R14702 VDD.n5569 VDD.n5502 7.49764
R14703 VDD.n3754 VDD.n3687 7.49764
R14704 VDD.n4012 VDD.n3945 7.49764
R14705 VDD.n4270 VDD.n4203 7.49764
R14706 VDD.n4528 VDD.n4461 7.49764
R14707 VDD.n4786 VDD.n4719 7.49764
R14708 VDD.n5047 VDD.n4980 7.49764
R14709 VDD.n5309 VDD.n5242 7.49764
R14710 VDD.n1606 VDD.n1605 7.39078
R14711 VDD.n1636 VDD.n1635 7.27155
R14712 VDD.n1917 VDD.t612 7.15136
R14713 VDD.n2238 VDD.t149 7.15136
R14714 VDD.n2496 VDD.t677 7.15136
R14715 VDD.n2754 VDD.t1252 7.15136
R14716 VDD.n3012 VDD.t94 7.15136
R14717 VDD.n3270 VDD.t77 7.15136
R14718 VDD.n3528 VDD.t1301 7.15136
R14719 VDD.n5855 VDD.t160 7.15136
R14720 VDD.n5601 VDD.t204 7.15136
R14721 VDD.n3786 VDD.t1193 7.15136
R14722 VDD.n4044 VDD.t694 7.15136
R14723 VDD.n4302 VDD.t1151 7.15136
R14724 VDD.n4560 VDD.t587 7.15136
R14725 VDD.n4818 VDD.t1221 7.15136
R14726 VDD.n5079 VDD.t582 7.15136
R14727 VDD.n5341 VDD.t98 7.15136
R14728 VDD.n1872 VDD.t356 7.14897
R14729 VDD.n2193 VDD.t611 7.14897
R14730 VDD.n2451 VDD.t104 7.14897
R14731 VDD.n2709 VDD.t1120 7.14897
R14732 VDD.n2967 VDD.t406 7.14897
R14733 VDD.n3225 VDD.t776 7.14897
R14734 VDD.n3483 VDD.t180 7.14897
R14735 VDD.n5810 VDD.t1138 7.14897
R14736 VDD.n5556 VDD.t597 7.14897
R14737 VDD.n3741 VDD.t342 7.14897
R14738 VDD.n3999 VDD.t564 7.14897
R14739 VDD.n4257 VDD.t1216 7.14897
R14740 VDD.n4515 VDD.t1254 7.14897
R14741 VDD.n4773 VDD.t751 7.14897
R14742 VDD.n5034 VDD.t768 7.14897
R14743 VDD.n5296 VDD.t604 7.14897
R14744 VDD.n1976 VDD.n1926 7.05932
R14745 VDD.n1625 VDD 6.73734
R14746 VDD.n1833 VDD 6.4005
R14747 VDD.n1812 VDD 6.4005
R14748 VDD.n2133 VDD 6.4005
R14749 VDD.n2154 VDD 6.4005
R14750 VDD.n2391 VDD 6.4005
R14751 VDD.n2412 VDD 6.4005
R14752 VDD.n2649 VDD 6.4005
R14753 VDD.n2670 VDD 6.4005
R14754 VDD.n2907 VDD 6.4005
R14755 VDD.n2928 VDD 6.4005
R14756 VDD.n3165 VDD 6.4005
R14757 VDD.n3186 VDD 6.4005
R14758 VDD.n3423 VDD 6.4005
R14759 VDD.n3444 VDD 6.4005
R14760 VDD.n5750 VDD 6.4005
R14761 VDD.n5771 VDD 6.4005
R14762 VDD.n5496 VDD 6.4005
R14763 VDD.n5517 VDD 6.4005
R14764 VDD.n3681 VDD 6.4005
R14765 VDD.n3702 VDD 6.4005
R14766 VDD.n3939 VDD 6.4005
R14767 VDD.n3960 VDD 6.4005
R14768 VDD.n4197 VDD 6.4005
R14769 VDD.n4218 VDD 6.4005
R14770 VDD.n4455 VDD 6.4005
R14771 VDD.n4476 VDD 6.4005
R14772 VDD.n4713 VDD 6.4005
R14773 VDD.n4734 VDD 6.4005
R14774 VDD.n4995 VDD 6.4005
R14775 VDD.n4974 VDD 6.4005
R14776 VDD.n5257 VDD 6.4005
R14777 VDD.n5236 VDD 6.4005
R14778 VDD.n19 VDD.n18 6.4005
R14779 VDD.n336 VDD.n335 6.4005
R14780 VDD.n1646 VDD.n1644 6.23487
R14781 VDD.n1652 VDD 5.65631
R14782 VDD.n1631 VDD 5.65631
R14783 VDD.n853 VDD.n852 5.64756
R14784 VDD.n844 VDD.n843 5.64756
R14785 VDD.n950 VDD.n949 5.64756
R14786 VDD.n1096 VDD.n1095 5.64756
R14787 VDD.n1048 VDD.n1047 5.64756
R14788 VDD.n58 VDD.n57 5.64756
R14789 VDD.n49 VDD.n48 5.64756
R14790 VDD.n155 VDD.n154 5.64756
R14791 VDD.n301 VDD.n300 5.64756
R14792 VDD.n253 VDD.n252 5.64756
R14793 VDD.n452 VDD.n451 5.64756
R14794 VDD.n443 VDD.n442 5.64756
R14795 VDD.n549 VDD.n548 5.64756
R14796 VDD.n691 VDD.n690 5.64756
R14797 VDD.n643 VDD.n642 5.64756
R14798 VDD.n1446 VDD.n1445 5.64756
R14799 VDD.n1415 VDD.n1414 5.64756
R14800 VDD.n1279 VDD.n1278 5.64756
R14801 VDD.n1494 VDD.n1493 5.64756
R14802 VDD.n1254 VDD.n1253 5.64756
R14803 VDD.n2128 VDD.n2013 5.34133
R14804 VDD.n1626 VDD 5.31371
R14805 VDD.n1360 VDD.n1359 5.27114
R14806 VDD.n1505 VDD.n1504 5.27114
R14807 VDD.n1288 VDD.n1287 5.27114
R14808 VDD.n1428 VDD.t637 5.20598
R14809 VDD.n1653 VDD.n1652 4.99699
R14810 VDD.n1648 VDD.n1647 4.98671
R14811 VDD.n880 VDD.n879 4.89462
R14812 VDD.n926 VDD.n925 4.89462
R14813 VDD.n963 VDD.n962 4.89462
R14814 VDD.n1073 VDD.n1072 4.89462
R14815 VDD.n1026 VDD.n1025 4.89462
R14816 VDD.n85 VDD.n84 4.89462
R14817 VDD.n131 VDD.n130 4.89462
R14818 VDD.n168 VDD.n167 4.89462
R14819 VDD.n278 VDD.n277 4.89462
R14820 VDD.n231 VDD.n230 4.89462
R14821 VDD.n479 VDD.n478 4.89462
R14822 VDD.n525 VDD.n524 4.89462
R14823 VDD.n558 VDD.n557 4.89462
R14824 VDD.n668 VDD.n667 4.89462
R14825 VDD.n621 VDD.n620 4.89462
R14826 VDD.n1330 VDD.n1329 4.89462
R14827 VDD.n1386 VDD.n1385 4.89462
R14828 VDD.n1300 VDD.n1299 4.89462
R14829 VDD.n1472 VDD.n1471 4.89462
R14830 VDD.n1522 VDD.n1521 4.89462
R14831 VDD.n1618 VDD 4.8645
R14832 VDD.n1833 VDD.n1832 4.6505
R14833 VDD.n1834 VDD.n1829 4.6505
R14834 VDD.n1812 VDD.n1811 4.6505
R14835 VDD.n1796 VDD.n1781 4.6505
R14836 VDD.n1796 VDD.n1795 4.6505
R14837 VDD.n1791 VDD.n1790 4.6505
R14838 VDD.n1793 VDD.n1791 4.6505
R14839 VDD.n1789 VDD.n1780 4.6505
R14840 VDD.n1787 VDD.n1783 4.6505
R14841 VDD.n1786 VDD.n1785 4.6505
R14842 VDD.n1794 VDD.n1780 4.6505
R14843 VDD.n1783 VDD.n1782 4.6505
R14844 VDD.n1785 VDD.n1784 4.6505
R14845 VDD.n2133 VDD.n2132 4.6505
R14846 VDD.n2154 VDD.n2153 4.6505
R14847 VDD.n2155 VDD.n2150 4.6505
R14848 VDD.n2004 VDD.n1989 4.6505
R14849 VDD.n2004 VDD.n2003 4.6505
R14850 VDD.n1999 VDD.n1998 4.6505
R14851 VDD.n2001 VDD.n1999 4.6505
R14852 VDD.n1997 VDD.n1988 4.6505
R14853 VDD.n1995 VDD.n1991 4.6505
R14854 VDD.n1994 VDD.n1993 4.6505
R14855 VDD.n2002 VDD.n1988 4.6505
R14856 VDD.n1991 VDD.n1990 4.6505
R14857 VDD.n1993 VDD.n1992 4.6505
R14858 VDD.n2391 VDD.n2390 4.6505
R14859 VDD.n2412 VDD.n2411 4.6505
R14860 VDD.n2413 VDD.n2408 4.6505
R14861 VDD.n2375 VDD.n2360 4.6505
R14862 VDD.n2375 VDD.n2374 4.6505
R14863 VDD.n2370 VDD.n2369 4.6505
R14864 VDD.n2372 VDD.n2370 4.6505
R14865 VDD.n2368 VDD.n2359 4.6505
R14866 VDD.n2366 VDD.n2362 4.6505
R14867 VDD.n2365 VDD.n2364 4.6505
R14868 VDD.n2373 VDD.n2359 4.6505
R14869 VDD.n2362 VDD.n2361 4.6505
R14870 VDD.n2364 VDD.n2363 4.6505
R14871 VDD.n2649 VDD.n2648 4.6505
R14872 VDD.n2670 VDD.n2669 4.6505
R14873 VDD.n2671 VDD.n2666 4.6505
R14874 VDD.n2633 VDD.n2618 4.6505
R14875 VDD.n2633 VDD.n2632 4.6505
R14876 VDD.n2628 VDD.n2627 4.6505
R14877 VDD.n2630 VDD.n2628 4.6505
R14878 VDD.n2626 VDD.n2617 4.6505
R14879 VDD.n2624 VDD.n2620 4.6505
R14880 VDD.n2623 VDD.n2622 4.6505
R14881 VDD.n2631 VDD.n2617 4.6505
R14882 VDD.n2620 VDD.n2619 4.6505
R14883 VDD.n2622 VDD.n2621 4.6505
R14884 VDD.n2907 VDD.n2906 4.6505
R14885 VDD.n2928 VDD.n2927 4.6505
R14886 VDD.n2929 VDD.n2924 4.6505
R14887 VDD.n2891 VDD.n2876 4.6505
R14888 VDD.n2891 VDD.n2890 4.6505
R14889 VDD.n2886 VDD.n2885 4.6505
R14890 VDD.n2888 VDD.n2886 4.6505
R14891 VDD.n2884 VDD.n2875 4.6505
R14892 VDD.n2882 VDD.n2878 4.6505
R14893 VDD.n2881 VDD.n2880 4.6505
R14894 VDD.n2889 VDD.n2875 4.6505
R14895 VDD.n2878 VDD.n2877 4.6505
R14896 VDD.n2880 VDD.n2879 4.6505
R14897 VDD.n3165 VDD.n3164 4.6505
R14898 VDD.n3186 VDD.n3185 4.6505
R14899 VDD.n3187 VDD.n3182 4.6505
R14900 VDD.n3149 VDD.n3134 4.6505
R14901 VDD.n3149 VDD.n3148 4.6505
R14902 VDD.n3144 VDD.n3143 4.6505
R14903 VDD.n3146 VDD.n3144 4.6505
R14904 VDD.n3142 VDD.n3133 4.6505
R14905 VDD.n3140 VDD.n3136 4.6505
R14906 VDD.n3139 VDD.n3138 4.6505
R14907 VDD.n3147 VDD.n3133 4.6505
R14908 VDD.n3136 VDD.n3135 4.6505
R14909 VDD.n3138 VDD.n3137 4.6505
R14910 VDD.n3423 VDD.n3422 4.6505
R14911 VDD.n3444 VDD.n3443 4.6505
R14912 VDD.n3445 VDD.n3440 4.6505
R14913 VDD.n3407 VDD.n3392 4.6505
R14914 VDD.n3407 VDD.n3406 4.6505
R14915 VDD.n3402 VDD.n3401 4.6505
R14916 VDD.n3404 VDD.n3402 4.6505
R14917 VDD.n3400 VDD.n3391 4.6505
R14918 VDD.n3398 VDD.n3394 4.6505
R14919 VDD.n3397 VDD.n3396 4.6505
R14920 VDD.n3405 VDD.n3391 4.6505
R14921 VDD.n3394 VDD.n3393 4.6505
R14922 VDD.n3396 VDD.n3395 4.6505
R14923 VDD.n5750 VDD.n5749 4.6505
R14924 VDD.n5771 VDD.n5770 4.6505
R14925 VDD.n5772 VDD.n5767 4.6505
R14926 VDD.n5737 VDD.n5722 4.6505
R14927 VDD.n5737 VDD.n5736 4.6505
R14928 VDD.n5732 VDD.n5731 4.6505
R14929 VDD.n5734 VDD.n5732 4.6505
R14930 VDD.n5730 VDD.n5721 4.6505
R14931 VDD.n5728 VDD.n5724 4.6505
R14932 VDD.n5727 VDD.n5726 4.6505
R14933 VDD.n5735 VDD.n5721 4.6505
R14934 VDD.n5724 VDD.n5723 4.6505
R14935 VDD.n5726 VDD.n5725 4.6505
R14936 VDD.n5496 VDD.n5495 4.6505
R14937 VDD.n5517 VDD.n5516 4.6505
R14938 VDD.n5518 VDD.n5513 4.6505
R14939 VDD.n5483 VDD.n5468 4.6505
R14940 VDD.n5483 VDD.n5482 4.6505
R14941 VDD.n5478 VDD.n5477 4.6505
R14942 VDD.n5480 VDD.n5478 4.6505
R14943 VDD.n5476 VDD.n5467 4.6505
R14944 VDD.n5474 VDD.n5470 4.6505
R14945 VDD.n5473 VDD.n5472 4.6505
R14946 VDD.n5481 VDD.n5467 4.6505
R14947 VDD.n5470 VDD.n5469 4.6505
R14948 VDD.n5472 VDD.n5471 4.6505
R14949 VDD.n3681 VDD.n3680 4.6505
R14950 VDD.n3702 VDD.n3701 4.6505
R14951 VDD.n3703 VDD.n3698 4.6505
R14952 VDD.n3665 VDD.n3650 4.6505
R14953 VDD.n3665 VDD.n3664 4.6505
R14954 VDD.n3660 VDD.n3659 4.6505
R14955 VDD.n3662 VDD.n3660 4.6505
R14956 VDD.n3658 VDD.n3649 4.6505
R14957 VDD.n3656 VDD.n3652 4.6505
R14958 VDD.n3655 VDD.n3654 4.6505
R14959 VDD.n3663 VDD.n3649 4.6505
R14960 VDD.n3652 VDD.n3651 4.6505
R14961 VDD.n3654 VDD.n3653 4.6505
R14962 VDD.n3939 VDD.n3938 4.6505
R14963 VDD.n3960 VDD.n3959 4.6505
R14964 VDD.n3961 VDD.n3956 4.6505
R14965 VDD.n3923 VDD.n3908 4.6505
R14966 VDD.n3923 VDD.n3922 4.6505
R14967 VDD.n3918 VDD.n3917 4.6505
R14968 VDD.n3920 VDD.n3918 4.6505
R14969 VDD.n3916 VDD.n3907 4.6505
R14970 VDD.n3914 VDD.n3910 4.6505
R14971 VDD.n3913 VDD.n3912 4.6505
R14972 VDD.n3921 VDD.n3907 4.6505
R14973 VDD.n3910 VDD.n3909 4.6505
R14974 VDD.n3912 VDD.n3911 4.6505
R14975 VDD.n4197 VDD.n4196 4.6505
R14976 VDD.n4218 VDD.n4217 4.6505
R14977 VDD.n4219 VDD.n4214 4.6505
R14978 VDD.n4181 VDD.n4166 4.6505
R14979 VDD.n4181 VDD.n4180 4.6505
R14980 VDD.n4176 VDD.n4175 4.6505
R14981 VDD.n4178 VDD.n4176 4.6505
R14982 VDD.n4174 VDD.n4165 4.6505
R14983 VDD.n4172 VDD.n4168 4.6505
R14984 VDD.n4171 VDD.n4170 4.6505
R14985 VDD.n4179 VDD.n4165 4.6505
R14986 VDD.n4168 VDD.n4167 4.6505
R14987 VDD.n4170 VDD.n4169 4.6505
R14988 VDD.n4455 VDD.n4454 4.6505
R14989 VDD.n4476 VDD.n4475 4.6505
R14990 VDD.n4477 VDD.n4472 4.6505
R14991 VDD.n4439 VDD.n4424 4.6505
R14992 VDD.n4439 VDD.n4438 4.6505
R14993 VDD.n4434 VDD.n4433 4.6505
R14994 VDD.n4436 VDD.n4434 4.6505
R14995 VDD.n4432 VDD.n4423 4.6505
R14996 VDD.n4430 VDD.n4426 4.6505
R14997 VDD.n4429 VDD.n4428 4.6505
R14998 VDD.n4437 VDD.n4423 4.6505
R14999 VDD.n4426 VDD.n4425 4.6505
R15000 VDD.n4428 VDD.n4427 4.6505
R15001 VDD.n4713 VDD.n4712 4.6505
R15002 VDD.n4734 VDD.n4733 4.6505
R15003 VDD.n4735 VDD.n4730 4.6505
R15004 VDD.n4697 VDD.n4682 4.6505
R15005 VDD.n4697 VDD.n4696 4.6505
R15006 VDD.n4692 VDD.n4691 4.6505
R15007 VDD.n4694 VDD.n4692 4.6505
R15008 VDD.n4690 VDD.n4681 4.6505
R15009 VDD.n4688 VDD.n4684 4.6505
R15010 VDD.n4687 VDD.n4686 4.6505
R15011 VDD.n4695 VDD.n4681 4.6505
R15012 VDD.n4684 VDD.n4683 4.6505
R15013 VDD.n4686 VDD.n4685 4.6505
R15014 VDD.n4956 VDD.n4941 4.6505
R15015 VDD.n4956 VDD.n4955 4.6505
R15016 VDD.n4951 VDD.n4950 4.6505
R15017 VDD.n4953 VDD.n4951 4.6505
R15018 VDD.n4949 VDD.n4940 4.6505
R15019 VDD.n4947 VDD.n4943 4.6505
R15020 VDD.n4946 VDD.n4945 4.6505
R15021 VDD.n4954 VDD.n4940 4.6505
R15022 VDD.n4943 VDD.n4942 4.6505
R15023 VDD.n4945 VDD.n4944 4.6505
R15024 VDD.n4995 VDD.n4994 4.6505
R15025 VDD.n4996 VDD.n4991 4.6505
R15026 VDD.n4974 VDD.n4973 4.6505
R15027 VDD.n5106 VDD.n5091 4.6505
R15028 VDD.n5106 VDD.n5105 4.6505
R15029 VDD.n5101 VDD.n5100 4.6505
R15030 VDD.n5103 VDD.n5101 4.6505
R15031 VDD.n5099 VDD.n5090 4.6505
R15032 VDD.n5097 VDD.n5093 4.6505
R15033 VDD.n5096 VDD.n5095 4.6505
R15034 VDD.n5104 VDD.n5090 4.6505
R15035 VDD.n5093 VDD.n5092 4.6505
R15036 VDD.n5095 VDD.n5094 4.6505
R15037 VDD.n5257 VDD.n5256 4.6505
R15038 VDD.n5258 VDD.n5253 4.6505
R15039 VDD.n5236 VDD.n5235 4.6505
R15040 VDD.n12 VDD.n11 4.6505
R15041 VDD.n14 VDD.n13 4.6505
R15042 VDD.n16 VDD.n8 4.6505
R15043 VDD.n4 VDD.n2 4.6505
R15044 VDD.n23 VDD.n22 4.6505
R15045 VDD.n15 VDD.n6 4.6505
R15046 VDD.n18 VDD.n17 4.6505
R15047 VDD.n21 VDD.n20 4.6505
R15048 VDD.n30 VDD.n29 4.6505
R15049 VDD.n1006 VDD.n841 4.6505
R15050 VDD.n1014 VDD.n840 4.6505
R15051 VDD.n1015 VDD.n839 4.6505
R15052 VDD.n1061 VDD.n837 4.6505
R15053 VDD.n1062 VDD.n836 4.6505
R15054 VDD.n1108 VDD.n834 4.6505
R15055 VDD.n1109 VDD.n833 4.6505
R15056 VDD.n939 VDD.n938 4.6505
R15057 VDD.n937 VDD.n936 4.6505
R15058 VDD.n868 VDD.n859 4.6505
R15059 VDD.n869 VDD.n858 4.6505
R15060 VDD.n993 VDD.n992 4.6505
R15061 VDD.n995 VDD.n994 4.6505
R15062 VDD.n997 VDD.n996 4.6505
R15063 VDD.n999 VDD.n998 4.6505
R15064 VDD.n1002 VDD.n1001 4.6505
R15065 VDD.n1008 VDD.n1007 4.6505
R15066 VDD.n1011 VDD.n1010 4.6505
R15067 VDD.n1013 VDD.n1012 4.6505
R15068 VDD.n1017 VDD.n1016 4.6505
R15069 VDD.n1021 VDD.n1020 4.6505
R15070 VDD.n1023 VDD.n1022 4.6505
R15071 VDD.n1027 VDD.n1026 4.6505
R15072 VDD.n1029 VDD.n1028 4.6505
R15073 VDD.n1033 VDD.n1032 4.6505
R15074 VDD.n1035 VDD.n1034 4.6505
R15075 VDD.n1039 VDD.n1038 4.6505
R15076 VDD.n1043 VDD.n1042 4.6505
R15077 VDD.n1045 VDD.n1044 4.6505
R15078 VDD.n1049 VDD.n1048 4.6505
R15079 VDD.n1052 VDD.n1051 4.6505
R15080 VDD.n1057 VDD.n1056 4.6505
R15081 VDD.n1060 VDD.n1059 4.6505
R15082 VDD.n1064 VDD.n1063 4.6505
R15083 VDD.n1068 VDD.n1067 4.6505
R15084 VDD.n1070 VDD.n1069 4.6505
R15085 VDD.n1074 VDD.n1073 4.6505
R15086 VDD.n1076 VDD.n1075 4.6505
R15087 VDD.n1080 VDD.n1079 4.6505
R15088 VDD.n1082 VDD.n1081 4.6505
R15089 VDD.n1086 VDD.n1085 4.6505
R15090 VDD.n1090 VDD.n1089 4.6505
R15091 VDD.n1092 VDD.n1091 4.6505
R15092 VDD.n1097 VDD.n1096 4.6505
R15093 VDD.n1100 VDD.n1099 4.6505
R15094 VDD.n1105 VDD.n1104 4.6505
R15095 VDD.n1107 VDD.n1106 4.6505
R15096 VDD.n832 VDD.n831 4.6505
R15097 VDD.n958 VDD.n957 4.6505
R15098 VDD.n960 VDD.n959 4.6505
R15099 VDD.n964 VDD.n963 4.6505
R15100 VDD.n966 VDD.n965 4.6505
R15101 VDD.n970 VDD.n969 4.6505
R15102 VDD.n972 VDD.n971 4.6505
R15103 VDD.n976 VDD.n975 4.6505
R15104 VDD.n981 VDD.n980 4.6505
R15105 VDD.n954 VDD.n953 4.6505
R15106 VDD.n951 VDD.n950 4.6505
R15107 VDD.n947 VDD.n946 4.6505
R15108 VDD.n945 VDD.n944 4.6505
R15109 VDD.n941 VDD.n940 4.6505
R15110 VDD.n935 VDD.n934 4.6505
R15111 VDD.n933 VDD.n932 4.6505
R15112 VDD.n929 VDD.n928 4.6505
R15113 VDD.n927 VDD.n926 4.6505
R15114 VDD.n923 VDD.n922 4.6505
R15115 VDD.n921 VDD.n920 4.6505
R15116 VDD.n917 VDD.n916 4.6505
R15117 VDD.n915 VDD.n914 4.6505
R15118 VDD.n911 VDD.n910 4.6505
R15119 VDD.n906 VDD.n905 4.6505
R15120 VDD.n845 VDD.n844 4.6505
R15121 VDD.n861 VDD.n860 4.6505
R15122 VDD.n865 VDD.n864 4.6505
R15123 VDD.n867 VDD.n866 4.6505
R15124 VDD.n871 VDD.n870 4.6505
R15125 VDD.n875 VDD.n874 4.6505
R15126 VDD.n877 VDD.n876 4.6505
R15127 VDD.n881 VDD.n880 4.6505
R15128 VDD.n883 VDD.n882 4.6505
R15129 VDD.n887 VDD.n886 4.6505
R15130 VDD.n889 VDD.n888 4.6505
R15131 VDD.n893 VDD.n892 4.6505
R15132 VDD.n898 VDD.n897 4.6505
R15133 VDD.n857 VDD.n856 4.6505
R15134 VDD.n854 VDD.n853 4.6505
R15135 VDD.n850 VDD.n849 4.6505
R15136 VDD.n791 VDD.n790 4.6505
R15137 VDD.n797 VDD.n789 4.6505
R15138 VDD.n797 VDD.n787 4.6505
R15139 VDD.n796 VDD.n795 4.6505
R15140 VDD.n802 VDD.n800 4.6505
R15141 VDD.n803 VDD.n786 4.6505
R15142 VDD.n784 VDD.n783 4.6505
R15143 VDD.n808 VDD.n807 4.6505
R15144 VDD.n810 VDD.n809 4.6505
R15145 VDD.n814 VDD.n813 4.6505
R15146 VDD.n816 VDD.n815 4.6505
R15147 VDD.n818 VDD.n817 4.6505
R15148 VDD.n820 VDD.n819 4.6505
R15149 VDD.n822 VDD.n821 4.6505
R15150 VDD.n824 VDD.n823 4.6505
R15151 VDD.n802 VDD.n801 4.6505
R15152 VDD.n804 VDD.n803 4.6505
R15153 VDD.n764 VDD.n763 4.6505
R15154 VDD.n768 VDD.n761 4.6505
R15155 VDD.n767 VDD.n765 4.6505
R15156 VDD.n771 VDD.n769 4.6505
R15157 VDD.n774 VDD.n772 4.6505
R15158 VDD.n764 VDD.n762 4.6505
R15159 VDD.n767 VDD.n766 4.6505
R15160 VDD.n768 VDD.n759 4.6505
R15161 VDD.n771 VDD.n770 4.6505
R15162 VDD.n774 VDD.n773 4.6505
R15163 VDD.n775 VDD.n757 4.6505
R15164 VDD.n732 VDD.n727 4.6505
R15165 VDD.n734 VDD.n726 4.6505
R15166 VDD.n732 VDD.n731 4.6505
R15167 VDD.n734 VDD.n733 4.6505
R15168 VDD.n738 VDD.n737 4.6505
R15169 VDD.n743 VDD.n742 4.6505
R15170 VDD.n745 VDD.n744 4.6505
R15171 VDD.n747 VDD.n746 4.6505
R15172 VDD.n749 VDD.n748 4.6505
R15173 VDD.n751 VDD.n750 4.6505
R15174 VDD.n713 VDD.n709 4.6505
R15175 VDD.n715 VDD.n708 4.6505
R15176 VDD.n715 VDD.n714 4.6505
R15177 VDD.n717 VDD.n716 4.6505
R15178 VDD.n389 VDD.n388 4.6505
R15179 VDD.n395 VDD.n387 4.6505
R15180 VDD.n395 VDD.n385 4.6505
R15181 VDD.n394 VDD.n393 4.6505
R15182 VDD.n400 VDD.n398 4.6505
R15183 VDD.n401 VDD.n384 4.6505
R15184 VDD.n382 VDD.n381 4.6505
R15185 VDD.n406 VDD.n405 4.6505
R15186 VDD.n408 VDD.n407 4.6505
R15187 VDD.n412 VDD.n411 4.6505
R15188 VDD.n414 VDD.n413 4.6505
R15189 VDD.n416 VDD.n415 4.6505
R15190 VDD.n418 VDD.n417 4.6505
R15191 VDD.n420 VDD.n419 4.6505
R15192 VDD.n422 VDD.n421 4.6505
R15193 VDD.n400 VDD.n399 4.6505
R15194 VDD.n402 VDD.n401 4.6505
R15195 VDD.n361 VDD.n360 4.6505
R15196 VDD.n365 VDD.n358 4.6505
R15197 VDD.n364 VDD.n362 4.6505
R15198 VDD.n368 VDD.n366 4.6505
R15199 VDD.n371 VDD.n369 4.6505
R15200 VDD.n361 VDD.n359 4.6505
R15201 VDD.n364 VDD.n363 4.6505
R15202 VDD.n365 VDD.n356 4.6505
R15203 VDD.n368 VDD.n367 4.6505
R15204 VDD.n371 VDD.n370 4.6505
R15205 VDD.n372 VDD.n354 4.6505
R15206 VDD.n329 VDD.n328 4.6505
R15207 VDD.n331 VDD.n330 4.6505
R15208 VDD.n333 VDD.n325 4.6505
R15209 VDD.n321 VDD.n319 4.6505
R15210 VDD.n340 VDD.n339 4.6505
R15211 VDD.n332 VDD.n323 4.6505
R15212 VDD.n335 VDD.n334 4.6505
R15213 VDD.n338 VDD.n337 4.6505
R15214 VDD.n347 VDD.n346 4.6505
R15215 VDD.n1573 VDD.n1568 4.6505
R15216 VDD.n1575 VDD.n1567 4.6505
R15217 VDD.n1573 VDD.n1572 4.6505
R15218 VDD.n1575 VDD.n1574 4.6505
R15219 VDD.n1579 VDD.n1578 4.6505
R15220 VDD.n1584 VDD.n1583 4.6505
R15221 VDD.n1586 VDD.n1585 4.6505
R15222 VDD.n1588 VDD.n1587 4.6505
R15223 VDD.n1590 VDD.n1589 4.6505
R15224 VDD.n1592 VDD.n1591 4.6505
R15225 VDD.n1554 VDD.n1550 4.6505
R15226 VDD.n1556 VDD.n1549 4.6505
R15227 VDD.n1556 VDD.n1555 4.6505
R15228 VDD.n1558 VDD.n1557 4.6505
R15229 VDD.n1168 VDD.n1167 4.6505
R15230 VDD.n1166 VDD.n1165 4.6505
R15231 VDD.n1164 VDD.n1163 4.6505
R15232 VDD.n1162 VDD.n1161 4.6505
R15233 VDD.n1160 VDD.n1159 4.6505
R15234 VDD.n1158 VDD.n1157 4.6505
R15235 VDD.n1156 VDD.n1155 4.6505
R15236 VDD.n1154 VDD.n1153 4.6505
R15237 VDD.n1152 VDD.n1151 4.6505
R15238 VDD.n1150 VDD.n1149 4.6505
R15239 VDD.n1148 VDD.n1147 4.6505
R15240 VDD.n1146 VDD.n1145 4.6505
R15241 VDD.n1125 VDD.n1121 4.6505
R15242 VDD.n1129 VDD.n1119 4.6505
R15243 VDD.n1135 VDD.n1116 4.6505
R15244 VDD.n1134 VDD.n1133 4.6505
R15245 VDD.n1132 VDD.n1118 4.6505
R15246 VDD.n1131 VDD.n1130 4.6505
R15247 VDD.n1128 VDD.n1127 4.6505
R15248 VDD.n1546 VDD.n1545 4.6505
R15249 VDD.n211 VDD.n46 4.6505
R15250 VDD.n219 VDD.n45 4.6505
R15251 VDD.n220 VDD.n44 4.6505
R15252 VDD.n266 VDD.n42 4.6505
R15253 VDD.n267 VDD.n41 4.6505
R15254 VDD.n313 VDD.n39 4.6505
R15255 VDD.n314 VDD.n38 4.6505
R15256 VDD.n144 VDD.n143 4.6505
R15257 VDD.n142 VDD.n141 4.6505
R15258 VDD.n73 VDD.n64 4.6505
R15259 VDD.n74 VDD.n63 4.6505
R15260 VDD.n198 VDD.n197 4.6505
R15261 VDD.n200 VDD.n199 4.6505
R15262 VDD.n202 VDD.n201 4.6505
R15263 VDD.n204 VDD.n203 4.6505
R15264 VDD.n207 VDD.n206 4.6505
R15265 VDD.n213 VDD.n212 4.6505
R15266 VDD.n216 VDD.n215 4.6505
R15267 VDD.n218 VDD.n217 4.6505
R15268 VDD.n222 VDD.n221 4.6505
R15269 VDD.n226 VDD.n225 4.6505
R15270 VDD.n228 VDD.n227 4.6505
R15271 VDD.n232 VDD.n231 4.6505
R15272 VDD.n234 VDD.n233 4.6505
R15273 VDD.n238 VDD.n237 4.6505
R15274 VDD.n240 VDD.n239 4.6505
R15275 VDD.n244 VDD.n243 4.6505
R15276 VDD.n248 VDD.n247 4.6505
R15277 VDD.n250 VDD.n249 4.6505
R15278 VDD.n254 VDD.n253 4.6505
R15279 VDD.n257 VDD.n256 4.6505
R15280 VDD.n262 VDD.n261 4.6505
R15281 VDD.n265 VDD.n264 4.6505
R15282 VDD.n269 VDD.n268 4.6505
R15283 VDD.n273 VDD.n272 4.6505
R15284 VDD.n275 VDD.n274 4.6505
R15285 VDD.n279 VDD.n278 4.6505
R15286 VDD.n281 VDD.n280 4.6505
R15287 VDD.n285 VDD.n284 4.6505
R15288 VDD.n287 VDD.n286 4.6505
R15289 VDD.n291 VDD.n290 4.6505
R15290 VDD.n295 VDD.n294 4.6505
R15291 VDD.n297 VDD.n296 4.6505
R15292 VDD.n302 VDD.n301 4.6505
R15293 VDD.n305 VDD.n304 4.6505
R15294 VDD.n310 VDD.n309 4.6505
R15295 VDD.n312 VDD.n311 4.6505
R15296 VDD.n37 VDD.n36 4.6505
R15297 VDD.n163 VDD.n162 4.6505
R15298 VDD.n165 VDD.n164 4.6505
R15299 VDD.n169 VDD.n168 4.6505
R15300 VDD.n171 VDD.n170 4.6505
R15301 VDD.n175 VDD.n174 4.6505
R15302 VDD.n177 VDD.n176 4.6505
R15303 VDD.n181 VDD.n180 4.6505
R15304 VDD.n186 VDD.n185 4.6505
R15305 VDD.n159 VDD.n158 4.6505
R15306 VDD.n156 VDD.n155 4.6505
R15307 VDD.n152 VDD.n151 4.6505
R15308 VDD.n150 VDD.n149 4.6505
R15309 VDD.n146 VDD.n145 4.6505
R15310 VDD.n140 VDD.n139 4.6505
R15311 VDD.n138 VDD.n137 4.6505
R15312 VDD.n134 VDD.n133 4.6505
R15313 VDD.n132 VDD.n131 4.6505
R15314 VDD.n128 VDD.n127 4.6505
R15315 VDD.n126 VDD.n125 4.6505
R15316 VDD.n122 VDD.n121 4.6505
R15317 VDD.n120 VDD.n119 4.6505
R15318 VDD.n116 VDD.n115 4.6505
R15319 VDD.n111 VDD.n110 4.6505
R15320 VDD.n50 VDD.n49 4.6505
R15321 VDD.n66 VDD.n65 4.6505
R15322 VDD.n70 VDD.n69 4.6505
R15323 VDD.n72 VDD.n71 4.6505
R15324 VDD.n76 VDD.n75 4.6505
R15325 VDD.n80 VDD.n79 4.6505
R15326 VDD.n82 VDD.n81 4.6505
R15327 VDD.n86 VDD.n85 4.6505
R15328 VDD.n88 VDD.n87 4.6505
R15329 VDD.n92 VDD.n91 4.6505
R15330 VDD.n94 VDD.n93 4.6505
R15331 VDD.n98 VDD.n97 4.6505
R15332 VDD.n103 VDD.n102 4.6505
R15333 VDD.n62 VDD.n61 4.6505
R15334 VDD.n59 VDD.n58 4.6505
R15335 VDD.n55 VDD.n54 4.6505
R15336 VDD.n601 VDD.n440 4.6505
R15337 VDD.n609 VDD.n439 4.6505
R15338 VDD.n610 VDD.n438 4.6505
R15339 VDD.n656 VDD.n436 4.6505
R15340 VDD.n657 VDD.n435 4.6505
R15341 VDD.n703 VDD.n433 4.6505
R15342 VDD.n704 VDD.n432 4.6505
R15343 VDD.n538 VDD.n537 4.6505
R15344 VDD.n536 VDD.n535 4.6505
R15345 VDD.n467 VDD.n458 4.6505
R15346 VDD.n468 VDD.n457 4.6505
R15347 VDD.n588 VDD.n587 4.6505
R15348 VDD.n590 VDD.n589 4.6505
R15349 VDD.n592 VDD.n591 4.6505
R15350 VDD.n594 VDD.n593 4.6505
R15351 VDD.n597 VDD.n596 4.6505
R15352 VDD.n603 VDD.n602 4.6505
R15353 VDD.n606 VDD.n605 4.6505
R15354 VDD.n608 VDD.n607 4.6505
R15355 VDD.n612 VDD.n611 4.6505
R15356 VDD.n616 VDD.n615 4.6505
R15357 VDD.n618 VDD.n617 4.6505
R15358 VDD.n622 VDD.n621 4.6505
R15359 VDD.n624 VDD.n623 4.6505
R15360 VDD.n628 VDD.n627 4.6505
R15361 VDD.n630 VDD.n629 4.6505
R15362 VDD.n634 VDD.n633 4.6505
R15363 VDD.n638 VDD.n637 4.6505
R15364 VDD.n640 VDD.n639 4.6505
R15365 VDD.n644 VDD.n643 4.6505
R15366 VDD.n647 VDD.n646 4.6505
R15367 VDD.n652 VDD.n651 4.6505
R15368 VDD.n655 VDD.n654 4.6505
R15369 VDD.n659 VDD.n658 4.6505
R15370 VDD.n663 VDD.n662 4.6505
R15371 VDD.n665 VDD.n664 4.6505
R15372 VDD.n669 VDD.n668 4.6505
R15373 VDD.n671 VDD.n670 4.6505
R15374 VDD.n675 VDD.n674 4.6505
R15375 VDD.n677 VDD.n676 4.6505
R15376 VDD.n681 VDD.n680 4.6505
R15377 VDD.n685 VDD.n684 4.6505
R15378 VDD.n687 VDD.n686 4.6505
R15379 VDD.n692 VDD.n691 4.6505
R15380 VDD.n695 VDD.n694 4.6505
R15381 VDD.n700 VDD.n699 4.6505
R15382 VDD.n702 VDD.n701 4.6505
R15383 VDD.n706 VDD.n705 4.6505
R15384 VDD.n431 VDD.n430 4.6505
R15385 VDD.n555 VDD.n554 4.6505
R15386 VDD.n559 VDD.n558 4.6505
R15387 VDD.n561 VDD.n560 4.6505
R15388 VDD.n565 VDD.n564 4.6505
R15389 VDD.n567 VDD.n566 4.6505
R15390 VDD.n571 VDD.n570 4.6505
R15391 VDD.n576 VDD.n575 4.6505
R15392 VDD.n553 VDD.n552 4.6505
R15393 VDD.n550 VDD.n549 4.6505
R15394 VDD.n546 VDD.n545 4.6505
R15395 VDD.n544 VDD.n543 4.6505
R15396 VDD.n540 VDD.n539 4.6505
R15397 VDD.n534 VDD.n533 4.6505
R15398 VDD.n532 VDD.n531 4.6505
R15399 VDD.n528 VDD.n527 4.6505
R15400 VDD.n526 VDD.n525 4.6505
R15401 VDD.n522 VDD.n521 4.6505
R15402 VDD.n520 VDD.n519 4.6505
R15403 VDD.n516 VDD.n515 4.6505
R15404 VDD.n514 VDD.n513 4.6505
R15405 VDD.n510 VDD.n509 4.6505
R15406 VDD.n505 VDD.n504 4.6505
R15407 VDD.n444 VDD.n443 4.6505
R15408 VDD.n460 VDD.n459 4.6505
R15409 VDD.n464 VDD.n463 4.6505
R15410 VDD.n466 VDD.n465 4.6505
R15411 VDD.n470 VDD.n469 4.6505
R15412 VDD.n474 VDD.n473 4.6505
R15413 VDD.n476 VDD.n475 4.6505
R15414 VDD.n480 VDD.n479 4.6505
R15415 VDD.n482 VDD.n481 4.6505
R15416 VDD.n486 VDD.n485 4.6505
R15417 VDD.n488 VDD.n487 4.6505
R15418 VDD.n492 VDD.n491 4.6505
R15419 VDD.n497 VDD.n496 4.6505
R15420 VDD.n456 VDD.n455 4.6505
R15421 VDD.n453 VDD.n452 4.6505
R15422 VDD.n449 VDD.n448 4.6505
R15423 VDD.n1358 VDD.n1357 4.6505
R15424 VDD.n1349 VDD.n1348 4.6505
R15425 VDD.n1347 VDD.n1346 4.6505
R15426 VDD.n1343 VDD.n1342 4.6505
R15427 VDD.n1341 VDD.n1340 4.6505
R15428 VDD.n1314 VDD.n1313 4.6505
R15429 VDD.n1365 VDD.n1364 4.6505
R15430 VDD.n1368 VDD.n1367 4.6505
R15431 VDD.n1356 VDD.n1355 4.6505
R15432 VDD.n1354 VDD.n1353 4.6505
R15433 VDD.n1351 VDD.n1350 4.6505
R15434 VDD.n1376 VDD.n1375 4.6505
R15435 VDD.n1381 VDD.n1380 4.6505
R15436 VDD.n1383 VDD.n1382 4.6505
R15437 VDD.n1387 VDD.n1386 4.6505
R15438 VDD.n1389 VDD.n1388 4.6505
R15439 VDD.n1393 VDD.n1392 4.6505
R15440 VDD.n1396 VDD.n1395 4.6505
R15441 VDD.n1405 VDD.n1404 4.6505
R15442 VDD.n1410 VDD.n1409 4.6505
R15443 VDD.n1412 VDD.n1411 4.6505
R15444 VDD.n1416 VDD.n1415 4.6505
R15445 VDD.n1418 VDD.n1417 4.6505
R15446 VDD.n1422 VDD.n1421 4.6505
R15447 VDD.n1425 VDD.n1424 4.6505
R15448 VDD.n1339 VDD.n1338 4.6505
R15449 VDD.n1337 VDD.n1336 4.6505
R15450 VDD.n1333 VDD.n1332 4.6505
R15451 VDD.n1331 VDD.n1330 4.6505
R15452 VDD.n1327 VDD.n1326 4.6505
R15453 VDD.n1324 VDD.n1323 4.6505
R15454 VDD.n1433 VDD.n1432 4.6505
R15455 VDD.n1437 VDD.n1436 4.6505
R15456 VDD.n1441 VDD.n1440 4.6505
R15457 VDD.n1443 VDD.n1442 4.6505
R15458 VDD.n1447 VDD.n1446 4.6505
R15459 VDD.n1449 VDD.n1448 4.6505
R15460 VDD.n1453 VDD.n1452 4.6505
R15461 VDD.n1317 VDD.n1316 4.6505
R15462 VDD.n1312 VDD.n1311 4.6505
R15463 VDD.n1310 VDD.n1309 4.6505
R15464 VDD.n1308 VDD.n1307 4.6505
R15465 VDD.n1527 VDD.n1258 4.6505
R15466 VDD.n1529 VDD.n1528 4.6505
R15467 VDD.n1533 VDD.n1532 4.6505
R15468 VDD.n1537 VDD.n1536 4.6505
R15469 VDD.n1539 VDD.n1538 4.6505
R15470 VDD.n1255 VDD.n1254 4.6505
R15471 VDD.n1251 VDD.n1250 4.6505
R15472 VDD.n1286 VDD.n1263 4.6505
R15473 VDD.n1460 VDD.n1262 4.6505
R15474 VDD.n1261 VDD.n1260 4.6505
R15475 VDD.n1510 VDD.n1259 4.6505
R15476 VDD.n1283 VDD.n1266 4.6505
R15477 VDD.n1285 VDD.n1284 4.6505
R15478 VDD.n1463 VDD.n1462 4.6505
R15479 VDD.n1467 VDD.n1466 4.6505
R15480 VDD.n1469 VDD.n1468 4.6505
R15481 VDD.n1473 VDD.n1472 4.6505
R15482 VDD.n1475 VDD.n1474 4.6505
R15483 VDD.n1479 VDD.n1478 4.6505
R15484 VDD.n1481 VDD.n1480 4.6505
R15485 VDD.n1485 VDD.n1484 4.6505
R15486 VDD.n1489 VDD.n1488 4.6505
R15487 VDD.n1491 VDD.n1490 4.6505
R15488 VDD.n1495 VDD.n1494 4.6505
R15489 VDD.n1497 VDD.n1496 4.6505
R15490 VDD.n1501 VDD.n1500 4.6505
R15491 VDD.n1503 VDD.n1502 4.6505
R15492 VDD.n1513 VDD.n1512 4.6505
R15493 VDD.n1517 VDD.n1516 4.6505
R15494 VDD.n1519 VDD.n1518 4.6505
R15495 VDD.n1523 VDD.n1522 4.6505
R15496 VDD.n1525 VDD.n1524 4.6505
R15497 VDD.n1303 VDD.n1302 4.6505
R15498 VDD.n1301 VDD.n1300 4.6505
R15499 VDD.n1297 VDD.n1296 4.6505
R15500 VDD.n1295 VDD.n1294 4.6505
R15501 VDD.n1291 VDD.n1290 4.6505
R15502 VDD.n1270 VDD.n1269 4.6505
R15503 VDD.n1274 VDD.n1273 4.6505
R15504 VDD.n1276 VDD.n1275 4.6505
R15505 VDD.n1280 VDD.n1279 4.6505
R15506 VDD.n1282 VDD.n1281 4.6505
R15507 VDD.n1234 VDD.n1233 4.6505
R15508 VDD.n1232 VDD.n1231 4.6505
R15509 VDD.n1230 VDD.n1229 4.6505
R15510 VDD.n1228 VDD.n1227 4.6505
R15511 VDD.n1226 VDD.n1225 4.6505
R15512 VDD.n1224 VDD.n1223 4.6505
R15513 VDD.n1222 VDD.n1221 4.6505
R15514 VDD.n1220 VDD.n1219 4.6505
R15515 VDD.n1218 VDD.n1217 4.6505
R15516 VDD.n1216 VDD.n1215 4.6505
R15517 VDD.n1214 VDD.n1213 4.6505
R15518 VDD.n1212 VDD.n1211 4.6505
R15519 VDD.n1191 VDD.n1187 4.6505
R15520 VDD.n1195 VDD.n1185 4.6505
R15521 VDD.n1201 VDD.n1182 4.6505
R15522 VDD.n1200 VDD.n1199 4.6505
R15523 VDD.n1198 VDD.n1184 4.6505
R15524 VDD.n1197 VDD.n1196 4.6505
R15525 VDD.n1194 VDD.n1193 4.6505
R15526 VDD.n1653 VDD.n1646 4.61128
R15527 VDD.n1946 VDD.n1943 4.58799
R15528 VDD.n1751 VDD.n1721 4.5005
R15529 VDD.n1751 VDD.n1716 4.5005
R15530 VDD.n1751 VDD.n1750 4.5005
R15531 VDD.n1777 VDD.n1776 4.5005
R15532 VDD.n1800 VDD.n1779 4.5005
R15533 VDD.n1800 VDD.n1799 4.5005
R15534 VDD.n1797 VDD.n1779 4.5005
R15535 VDD.n2100 VDD.n2070 4.5005
R15536 VDD.n2100 VDD.n2065 4.5005
R15537 VDD.n2100 VDD.n2099 4.5005
R15538 VDD.n1985 VDD.n1984 4.5005
R15539 VDD.n2008 VDD.n1987 4.5005
R15540 VDD.n2008 VDD.n2007 4.5005
R15541 VDD.n2005 VDD.n1987 4.5005
R15542 VDD.n2330 VDD.n2300 4.5005
R15543 VDD.n2330 VDD.n2295 4.5005
R15544 VDD.n2330 VDD.n2329 4.5005
R15545 VDD.n2356 VDD.n2355 4.5005
R15546 VDD.n2379 VDD.n2358 4.5005
R15547 VDD.n2379 VDD.n2378 4.5005
R15548 VDD.n2376 VDD.n2358 4.5005
R15549 VDD.n2588 VDD.n2558 4.5005
R15550 VDD.n2588 VDD.n2553 4.5005
R15551 VDD.n2588 VDD.n2587 4.5005
R15552 VDD.n2614 VDD.n2613 4.5005
R15553 VDD.n2637 VDD.n2616 4.5005
R15554 VDD.n2637 VDD.n2636 4.5005
R15555 VDD.n2634 VDD.n2616 4.5005
R15556 VDD.n2846 VDD.n2816 4.5005
R15557 VDD.n2846 VDD.n2811 4.5005
R15558 VDD.n2846 VDD.n2845 4.5005
R15559 VDD.n2872 VDD.n2871 4.5005
R15560 VDD.n2895 VDD.n2874 4.5005
R15561 VDD.n2895 VDD.n2894 4.5005
R15562 VDD.n2892 VDD.n2874 4.5005
R15563 VDD.n3104 VDD.n3074 4.5005
R15564 VDD.n3104 VDD.n3069 4.5005
R15565 VDD.n3104 VDD.n3103 4.5005
R15566 VDD.n3130 VDD.n3129 4.5005
R15567 VDD.n3153 VDD.n3132 4.5005
R15568 VDD.n3153 VDD.n3152 4.5005
R15569 VDD.n3150 VDD.n3132 4.5005
R15570 VDD.n3362 VDD.n3332 4.5005
R15571 VDD.n3362 VDD.n3327 4.5005
R15572 VDD.n3362 VDD.n3361 4.5005
R15573 VDD.n3388 VDD.n3387 4.5005
R15574 VDD.n3411 VDD.n3390 4.5005
R15575 VDD.n3411 VDD.n3410 4.5005
R15576 VDD.n3408 VDD.n3390 4.5005
R15577 VDD.n5692 VDD.n5662 4.5005
R15578 VDD.n5692 VDD.n5657 4.5005
R15579 VDD.n5692 VDD.n5691 4.5005
R15580 VDD.n5718 VDD.n5717 4.5005
R15581 VDD.n5741 VDD.n5720 4.5005
R15582 VDD.n5741 VDD.n5740 4.5005
R15583 VDD.n5738 VDD.n5720 4.5005
R15584 VDD.n5438 VDD.n5408 4.5005
R15585 VDD.n5438 VDD.n5403 4.5005
R15586 VDD.n5438 VDD.n5437 4.5005
R15587 VDD.n5464 VDD.n5463 4.5005
R15588 VDD.n5487 VDD.n5466 4.5005
R15589 VDD.n5487 VDD.n5486 4.5005
R15590 VDD.n5484 VDD.n5466 4.5005
R15591 VDD.n3620 VDD.n3590 4.5005
R15592 VDD.n3620 VDD.n3585 4.5005
R15593 VDD.n3620 VDD.n3619 4.5005
R15594 VDD.n3646 VDD.n3645 4.5005
R15595 VDD.n3669 VDD.n3648 4.5005
R15596 VDD.n3669 VDD.n3668 4.5005
R15597 VDD.n3666 VDD.n3648 4.5005
R15598 VDD.n3878 VDD.n3848 4.5005
R15599 VDD.n3878 VDD.n3843 4.5005
R15600 VDD.n3878 VDD.n3877 4.5005
R15601 VDD.n3904 VDD.n3903 4.5005
R15602 VDD.n3927 VDD.n3906 4.5005
R15603 VDD.n3927 VDD.n3926 4.5005
R15604 VDD.n3924 VDD.n3906 4.5005
R15605 VDD.n4136 VDD.n4106 4.5005
R15606 VDD.n4136 VDD.n4101 4.5005
R15607 VDD.n4136 VDD.n4135 4.5005
R15608 VDD.n4162 VDD.n4161 4.5005
R15609 VDD.n4185 VDD.n4164 4.5005
R15610 VDD.n4185 VDD.n4184 4.5005
R15611 VDD.n4182 VDD.n4164 4.5005
R15612 VDD.n4394 VDD.n4364 4.5005
R15613 VDD.n4394 VDD.n4359 4.5005
R15614 VDD.n4394 VDD.n4393 4.5005
R15615 VDD.n4420 VDD.n4419 4.5005
R15616 VDD.n4443 VDD.n4422 4.5005
R15617 VDD.n4443 VDD.n4442 4.5005
R15618 VDD.n4440 VDD.n4422 4.5005
R15619 VDD.n4652 VDD.n4622 4.5005
R15620 VDD.n4652 VDD.n4617 4.5005
R15621 VDD.n4652 VDD.n4651 4.5005
R15622 VDD.n4678 VDD.n4677 4.5005
R15623 VDD.n4701 VDD.n4680 4.5005
R15624 VDD.n4701 VDD.n4700 4.5005
R15625 VDD.n4698 VDD.n4680 4.5005
R15626 VDD.n4910 VDD.n4880 4.5005
R15627 VDD.n4910 VDD.n4875 4.5005
R15628 VDD.n4910 VDD.n4909 4.5005
R15629 VDD.n4937 VDD.n4936 4.5005
R15630 VDD.n4960 VDD.n4939 4.5005
R15631 VDD.n4960 VDD.n4959 4.5005
R15632 VDD.n4957 VDD.n4939 4.5005
R15633 VDD.n5202 VDD.n5172 4.5005
R15634 VDD.n5202 VDD.n5167 4.5005
R15635 VDD.n5202 VDD.n5201 4.5005
R15636 VDD.n5087 VDD.n5086 4.5005
R15637 VDD.n5110 VDD.n5089 4.5005
R15638 VDD.n5110 VDD.n5109 4.5005
R15639 VDD.n5107 VDD.n5089 4.5005
R15640 VDD.n1249 VDD.n1248 4.45149
R15641 VDD.n848 VDD.n847 4.4514
R15642 VDD.n53 VDD.n52 4.4514
R15643 VDD.n447 VDD.n446 4.4514
R15644 VDD.n1649 VDD.n1648 4.43268
R15645 VDD.n1887 VDD.t779 4.35136
R15646 VDD.n1874 VDD.t671 4.35136
R15647 VDD.n2195 VDD.t576 4.35136
R15648 VDD.n2208 VDD.t577 4.35136
R15649 VDD.n2453 VDD.t692 4.35136
R15650 VDD.n2466 VDD.t693 4.35136
R15651 VDD.n2711 VDD.t1082 4.35136
R15652 VDD.n2724 VDD.t557 4.35136
R15653 VDD.n2969 VDD.t1091 4.35136
R15654 VDD.n2982 VDD.t1092 4.35136
R15655 VDD.n3227 VDD.t575 4.35136
R15656 VDD.n3240 VDD.t688 4.35136
R15657 VDD.n3485 VDD.t571 4.35136
R15658 VDD.n3498 VDD.t1086 4.35136
R15659 VDD.n5812 VDD.t1083 4.35136
R15660 VDD.n5825 VDD.t1084 4.35136
R15661 VDD.n5558 VDD.t1184 4.35136
R15662 VDD.n5571 VDD.t1185 4.35136
R15663 VDD.n3743 VDD.t780 4.35136
R15664 VDD.n3756 VDD.t781 4.35136
R15665 VDD.n4001 VDD.t691 4.35136
R15666 VDD.n4014 VDD.t388 4.35136
R15667 VDD.n4259 VDD.t422 4.35136
R15668 VDD.n4272 VDD.t423 4.35136
R15669 VDD.n4517 VDD.t1089 4.35136
R15670 VDD.n4530 VDD.t1090 4.35136
R15671 VDD.n4775 VDD.t146 4.35136
R15672 VDD.n4788 VDD.t147 4.35136
R15673 VDD.n5049 VDD.t569 4.35136
R15674 VDD.n5036 VDD.t568 4.35136
R15675 VDD.n5311 VDD.t669 4.35136
R15676 VDD.n5298 VDD.t1081 4.35136
R15677 VDD.n1633 VDD 4.26717
R15678 VDD.n991 VDD.n990 4.14756
R15679 VDD.n196 VDD.n195 4.14756
R15680 VDD.n586 VDD.n585 4.14756
R15681 VDD.n783 VDD.n782 4.14168
R15682 VDD.n381 VDD.n380 4.14168
R15683 VDD.n1122 VDD.n1121 4.14168
R15684 VDD.n1188 VDD.n1187 4.14168
R15685 VDD.n806 VDD.n805 4.05611
R15686 VDD.n404 VDD.n403 4.05611
R15687 VDD.n25 VDD.n24 4.05569
R15688 VDD.n778 VDD.n777 4.05569
R15689 VDD.n375 VDD.n374 4.05569
R15690 VDD.n342 VDD.n341 4.05569
R15691 VDD.n1626 VDD.n1625 4.04261
R15692 VDD.n827 VDD.n826 4.01726
R15693 VDD.n754 VDD.n753 4.01726
R15694 VDD.n723 VDD.n722 4.01726
R15695 VDD.n425 VDD.n424 4.01726
R15696 VDD.n1595 VDD.n1594 4.01726
R15697 VDD.n1564 VDD.n1563 4.01726
R15698 VDD.n33 VDD.n32 4.01682
R15699 VDD.n350 VDD.n349 4.01682
R15700 VDD.n1815 VDD.n1814 3.96837
R15701 VDD.n2136 VDD.n2135 3.96837
R15702 VDD.n2394 VDD.n2393 3.96837
R15703 VDD.n2652 VDD.n2651 3.96837
R15704 VDD.n2910 VDD.n2909 3.96837
R15705 VDD.n3168 VDD.n3167 3.96837
R15706 VDD.n3426 VDD.n3425 3.96837
R15707 VDD.n5753 VDD.n5752 3.96837
R15708 VDD.n5499 VDD.n5498 3.96837
R15709 VDD.n3684 VDD.n3683 3.96837
R15710 VDD.n3942 VDD.n3941 3.96837
R15711 VDD.n4200 VDD.n4199 3.96837
R15712 VDD.n4458 VDD.n4457 3.96837
R15713 VDD.n4716 VDD.n4715 3.96837
R15714 VDD.n4977 VDD.n4976 3.96837
R15715 VDD.n5239 VDD.n5238 3.96837
R15716 VDD.n1137 VDD.n1136 3.96556
R15717 VDD.n1203 VDD.n1202 3.96556
R15718 VDD.n1638 VDD.n1637 3.88621
R15719 VDD.n1952 VDD.n1939 3.5871
R15720 VDD.n1694 VDD.n1683 3.52991
R15721 VDD.n2043 VDD.n2032 3.52991
R15722 VDD.n2273 VDD.n2262 3.52991
R15723 VDD.n2531 VDD.n2520 3.52991
R15724 VDD.n2789 VDD.n2778 3.52991
R15725 VDD.n3047 VDD.n3036 3.52991
R15726 VDD.n3305 VDD.n3294 3.52991
R15727 VDD.n5635 VDD.n5624 3.52991
R15728 VDD.n5381 VDD.n5370 3.52991
R15729 VDD.n3563 VDD.n3552 3.52991
R15730 VDD.n3821 VDD.n3810 3.52991
R15731 VDD.n4079 VDD.n4068 3.52991
R15732 VDD.n4337 VDD.n4326 3.52991
R15733 VDD.n4595 VDD.n4584 3.52991
R15734 VDD.n4853 VDD.n4842 3.52991
R15735 VDD.n5145 VDD.n5134 3.52991
R15736 VDD.n1608 VDD.n1607 3.46717
R15737 VDD.t430 VDD.n986 3.39336
R15738 VDD.t1480 VDD.n191 3.39336
R15739 VDD.n580 VDD.t1411 3.39336
R15740 VDD.n20 VDD.n19 3.38874
R15741 VDD.n813 VDD.n812 3.38874
R15742 VDD.n737 VDD.n736 3.38874
R15743 VDD.n411 VDD.n410 3.38874
R15744 VDD.n337 VDD.n336 3.38874
R15745 VDD.n1578 VDD.n1577 3.38874
R15746 VDD.n1980 VDD.n1922 3.1102
R15747 VDD.n1980 VDD.n1979 3.08146
R15748 VDD.n1701 VDD.n1700 3.03311
R15749 VDD.n2050 VDD.n2049 3.03311
R15750 VDD.n2280 VDD.n2279 3.03311
R15751 VDD.n2538 VDD.n2537 3.03311
R15752 VDD.n2796 VDD.n2795 3.03311
R15753 VDD.n3054 VDD.n3053 3.03311
R15754 VDD.n3312 VDD.n3311 3.03311
R15755 VDD.n5642 VDD.n5641 3.03311
R15756 VDD.n5388 VDD.n5387 3.03311
R15757 VDD.n3570 VDD.n3569 3.03311
R15758 VDD.n3828 VDD.n3827 3.03311
R15759 VDD.n4086 VDD.n4085 3.03311
R15760 VDD.n4344 VDD.n4343 3.03311
R15761 VDD.n4602 VDD.n4601 3.03311
R15762 VDD.n4860 VDD.n4859 3.03311
R15763 VDD.n5152 VDD.n5151 3.03311
R15764 VDD.n1609 VDD.n1608 3.03311
R15765 VDD VDD.n1622 3.02091
R15766 VDD.n1831 VDD 3.0005
R15767 VDD.n2152 VDD 3.0005
R15768 VDD.n2410 VDD 3.0005
R15769 VDD.n2668 VDD 3.0005
R15770 VDD.n2926 VDD 3.0005
R15771 VDD.n3184 VDD 3.0005
R15772 VDD.n3442 VDD 3.0005
R15773 VDD.n5769 VDD 3.0005
R15774 VDD.n5515 VDD 3.0005
R15775 VDD.n3700 VDD 3.0005
R15776 VDD.n3958 VDD 3.0005
R15777 VDD.n4216 VDD 3.0005
R15778 VDD.n4474 VDD 3.0005
R15779 VDD.n4732 VDD 3.0005
R15780 VDD.n4993 VDD 3.0005
R15781 VDD.n5255 VDD 3.0005
R15782 VDD.n1871 VDD.n1870 2.98717
R15783 VDD.n2192 VDD.n2191 2.98717
R15784 VDD.n2450 VDD.n2449 2.98717
R15785 VDD.n2708 VDD.n2707 2.98717
R15786 VDD.n2966 VDD.n2965 2.98717
R15787 VDD.n3224 VDD.n3223 2.98717
R15788 VDD.n3482 VDD.n3481 2.98717
R15789 VDD.n5809 VDD.n5808 2.98717
R15790 VDD.n5555 VDD.n5554 2.98717
R15791 VDD.n3740 VDD.n3739 2.98717
R15792 VDD.n3998 VDD.n3997 2.98717
R15793 VDD.n4256 VDD.n4255 2.98717
R15794 VDD.n4514 VDD.n4513 2.98717
R15795 VDD.n4772 VDD.n4771 2.98717
R15796 VDD.n5033 VDD.n5032 2.98717
R15797 VDD.n5295 VDD.n5294 2.98717
R15798 VDD.n4934 VDD.n4823 2.94072
R15799 VDD.n5345 VDD.n5344 2.81521
R15800 VDD.n1916 VDD.n1889 2.72837
R15801 VDD.n2237 VDD.n2210 2.72837
R15802 VDD.n2495 VDD.n2468 2.72837
R15803 VDD.n2753 VDD.n2726 2.72837
R15804 VDD.n3011 VDD.n2984 2.72837
R15805 VDD.n3269 VDD.n3242 2.72837
R15806 VDD.n3527 VDD.n3500 2.72837
R15807 VDD.n5854 VDD.n5827 2.72837
R15808 VDD.n5600 VDD.n5573 2.72837
R15809 VDD.n3785 VDD.n3758 2.72837
R15810 VDD.n4043 VDD.n4016 2.72837
R15811 VDD.n4301 VDD.n4274 2.72837
R15812 VDD.n4559 VDD.n4532 2.72837
R15813 VDD.n4817 VDD.n4790 2.72837
R15814 VDD.n5078 VDD.n5051 2.72837
R15815 VDD.n5340 VDD.n5313 2.72837
R15816 VDD.n794 VDD.n793 2.30978
R15817 VDD.n392 VDD.n391 2.30978
R15818 VDD.n1622 VDD.n1614 2.251
R15819 VDD.n1778 VDD.n1777 2.2278
R15820 VDD.n1986 VDD.n1985 2.2278
R15821 VDD.n2357 VDD.n2356 2.2278
R15822 VDD.n2615 VDD.n2614 2.2278
R15823 VDD.n2873 VDD.n2872 2.2278
R15824 VDD.n3131 VDD.n3130 2.2278
R15825 VDD.n3389 VDD.n3388 2.2278
R15826 VDD.n5719 VDD.n5718 2.2278
R15827 VDD.n5465 VDD.n5464 2.2278
R15828 VDD.n3647 VDD.n3646 2.2278
R15829 VDD.n3905 VDD.n3904 2.2278
R15830 VDD.n4163 VDD.n4162 2.2278
R15831 VDD.n4421 VDD.n4420 2.2278
R15832 VDD.n4679 VDD.n4678 2.2278
R15833 VDD.n4938 VDD.n4937 2.2278
R15834 VDD.n5088 VDD.n5087 2.2278
R15835 VDD VDD.n1633 2.13383
R15836 VDD.n1644 VDD 2.11184
R15837 VDD.n5345 VDD.n5085 1.85789
R15838 VDD.n1655 VDD.n1642 1.59861
R15839 VDD.n1630 VDD 1.53093
R15840 VDD.n1981 VDD 1.52828
R15841 VDD.n1772 VDD.n1771 1.51475
R15842 VDD.n2121 VDD.n2120 1.51475
R15843 VDD.n2351 VDD.n2350 1.51475
R15844 VDD.n2609 VDD.n2608 1.51475
R15845 VDD.n2867 VDD.n2866 1.51475
R15846 VDD.n3125 VDD.n3124 1.51475
R15847 VDD.n3383 VDD.n3382 1.51475
R15848 VDD.n5713 VDD.n5712 1.51475
R15849 VDD.n5459 VDD.n5458 1.51475
R15850 VDD.n3641 VDD.n3640 1.51475
R15851 VDD.n3899 VDD.n3898 1.51475
R15852 VDD.n4157 VDD.n4156 1.51475
R15853 VDD.n4415 VDD.n4414 1.51475
R15854 VDD.n4673 VDD.n4672 1.51475
R15855 VDD.n4931 VDD.n4930 1.51475
R15856 VDD.n5223 VDD.n5222 1.51475
R15857 VDD.n1945 VDD.t1286 1.50409
R15858 VDD.n1924 VDD.t1056 1.50409
R15859 VDD.n1924 VDD.t1288 1.50409
R15860 VDD.n1918 VDD.n1917 1.49778
R15861 VDD.n2239 VDD.n2238 1.49778
R15862 VDD.n2497 VDD.n2496 1.49778
R15863 VDD.n2755 VDD.n2754 1.49778
R15864 VDD.n3013 VDD.n3012 1.49778
R15865 VDD.n3271 VDD.n3270 1.49778
R15866 VDD.n3529 VDD.n3528 1.49778
R15867 VDD.n5856 VDD.n5855 1.49778
R15868 VDD.n5602 VDD.n5601 1.49778
R15869 VDD.n3787 VDD.n3786 1.49778
R15870 VDD.n4045 VDD.n4044 1.49778
R15871 VDD.n4303 VDD.n4302 1.49778
R15872 VDD.n4561 VDD.n4560 1.49778
R15873 VDD.n4819 VDD.n4818 1.49778
R15874 VDD.n5080 VDD.n5079 1.49778
R15875 VDD.n5342 VDD.n5341 1.49778
R15876 VDD.n2013 VDD.n2012 1.47642
R15877 VDD.n1661 VDD.n1660 1.43354
R15878 VDD.n1740 VDD.n1729 1.42272
R15879 VDD.n2089 VDD.n2078 1.42272
R15880 VDD.n2319 VDD.n2308 1.42272
R15881 VDD.n2577 VDD.n2566 1.42272
R15882 VDD.n2835 VDD.n2824 1.42272
R15883 VDD.n3093 VDD.n3082 1.42272
R15884 VDD.n3351 VDD.n3340 1.42272
R15885 VDD.n5681 VDD.n5670 1.42272
R15886 VDD.n5427 VDD.n5416 1.42272
R15887 VDD.n3609 VDD.n3598 1.42272
R15888 VDD.n3867 VDD.n3856 1.42272
R15889 VDD.n4125 VDD.n4114 1.42272
R15890 VDD.n4383 VDD.n4372 1.42272
R15891 VDD.n4641 VDD.n4630 1.42272
R15892 VDD.n4899 VDD.n4888 1.42272
R15893 VDD.n5191 VDD.n5180 1.42272
R15894 VDD.n1663 VDD.n1662 1.39179
R15895 VDD.n1887 VDD.n1886 1.25748
R15896 VDD.n2208 VDD.n2207 1.25748
R15897 VDD.n2466 VDD.n2465 1.25748
R15898 VDD.n2724 VDD.n2723 1.25748
R15899 VDD.n2982 VDD.n2981 1.25748
R15900 VDD.n3240 VDD.n3239 1.25748
R15901 VDD.n3498 VDD.n3497 1.25748
R15902 VDD.n5825 VDD.n5824 1.25748
R15903 VDD.n5571 VDD.n5570 1.25748
R15904 VDD.n3756 VDD.n3755 1.25748
R15905 VDD.n4014 VDD.n4013 1.25748
R15906 VDD.n4272 VDD.n4271 1.25748
R15907 VDD.n4530 VDD.n4529 1.25748
R15908 VDD.n4788 VDD.n4787 1.25748
R15909 VDD.n5049 VDD.n5048 1.25748
R15910 VDD.n5311 VDD.n5310 1.25748
R15911 VDD.n1651 VDD.n1650 1.25267
R15912 VDD.n1655 VDD.n1654 1.21925
R15913 VDD.n874 VDD.n873 1.12991
R15914 VDD.n932 VDD.n931 1.12991
R15915 VDD.n957 VDD.n956 1.12991
R15916 VDD.n1067 VDD.n1066 1.12991
R15917 VDD.n1020 VDD.n1019 1.12991
R15918 VDD.n79 VDD.n78 1.12991
R15919 VDD.n137 VDD.n136 1.12991
R15920 VDD.n162 VDD.n161 1.12991
R15921 VDD.n272 VDD.n271 1.12991
R15922 VDD.n225 VDD.n224 1.12991
R15923 VDD.n473 VDD.n472 1.12991
R15924 VDD.n531 VDD.n530 1.12991
R15925 VDD.n430 VDD.n429 1.12991
R15926 VDD.n662 VDD.n661 1.12991
R15927 VDD.n615 VDD.n614 1.12991
R15928 VDD.n1336 VDD.n1335 1.12991
R15929 VDD.n1380 VDD.n1379 1.12991
R15930 VDD.n1307 VDD.n1306 1.12991
R15931 VDD.n1466 VDD.n1465 1.12991
R15932 VDD.n1516 VDD.n1515 1.12991
R15933 VDD.n1652 VDD.n1651 1.11354
R15934 VDD.n1631 VDD.n1630 1.11354
R15935 VDD.n1623 VDD.n1613 1.10388
R15936 VDD.n1731 VDD.n1716 1.06717
R15937 VDD.n2080 VDD.n2065 1.06717
R15938 VDD.n2310 VDD.n2295 1.06717
R15939 VDD.n2568 VDD.n2553 1.06717
R15940 VDD.n2826 VDD.n2811 1.06717
R15941 VDD.n3084 VDD.n3069 1.06717
R15942 VDD.n3342 VDD.n3327 1.06717
R15943 VDD.n5672 VDD.n5657 1.06717
R15944 VDD.n5418 VDD.n5403 1.06717
R15945 VDD.n3600 VDD.n3585 1.06717
R15946 VDD.n3858 VDD.n3843 1.06717
R15947 VDD.n4116 VDD.n4101 1.06717
R15948 VDD.n4374 VDD.n4359 1.06717
R15949 VDD.n4632 VDD.n4617 1.06717
R15950 VDD.n4890 VDD.n4875 1.06717
R15951 VDD.n5182 VDD.n5167 1.06717
R15952 VDD.n1608 VDD.n1606 1.06717
R15953 VDD.n1607 VDD 1.06717
R15954 VDD.n1873 VDD.n1872 1.00783
R15955 VDD.n2194 VDD.n2193 1.00687
R15956 VDD.n2452 VDD.n2451 1.00687
R15957 VDD.n2710 VDD.n2709 1.00687
R15958 VDD.n2968 VDD.n2967 1.00687
R15959 VDD.n3226 VDD.n3225 1.00687
R15960 VDD.n3484 VDD.n3483 1.00687
R15961 VDD.n5811 VDD.n5810 1.00687
R15962 VDD.n5557 VDD.n5556 1.00687
R15963 VDD.n3742 VDD.n3741 1.00687
R15964 VDD.n4000 VDD.n3999 1.00687
R15965 VDD.n4258 VDD.n4257 1.00687
R15966 VDD.n4516 VDD.n4515 1.00687
R15967 VDD.n4774 VDD.n4773 1.00687
R15968 VDD.n5035 VDD.n5034 1.00687
R15969 VDD.n5297 VDD.n5296 1.00687
R15970 VDD.n1644 VDD 0.970197
R15971 VDD.n1704 VDD.n1681 0.9605
R15972 VDD.n2053 VDD.n2030 0.9605
R15973 VDD.n2283 VDD.n2260 0.9605
R15974 VDD.n2541 VDD.n2518 0.9605
R15975 VDD.n2799 VDD.n2776 0.9605
R15976 VDD.n3057 VDD.n3034 0.9605
R15977 VDD.n3315 VDD.n3292 0.9605
R15978 VDD.n5645 VDD.n5622 0.9605
R15979 VDD.n5391 VDD.n5368 0.9605
R15980 VDD.n3573 VDD.n3550 0.9605
R15981 VDD.n3831 VDD.n3808 0.9605
R15982 VDD.n4089 VDD.n4066 0.9605
R15983 VDD.n4347 VDD.n4324 0.9605
R15984 VDD.n4605 VDD.n4582 0.9605
R15985 VDD.n4863 VDD.n4840 0.9605
R15986 VDD.n5155 VDD.n5132 0.9605
R15987 VDD.n1603 VDD.n1245 0.939577
R15988 VDD.n5866 VDD.n1982 0.885753
R15989 VDD.n1662 VDD.n1661 0.87764
R15990 VDD.n1113 VDD.n724 0.826983
R15991 VDD.n1598 VDD.n1565 0.826983
R15992 VDD.n1933 VDD.n1924 0.800961
R15993 VDD.n5868 VDD 0.78236
R15994 VDD.n1619 VDD.n1618 0.7685
R15995 VDD.n1956 VDD.n1943 0.738962
R15996 VDD.n1638 VDD.n1636 0.686214
R15997 VDD.n1657 VDD.n1656 0.683536
R15998 VDD.n1663 VDD.n1603 0.673542
R15999 VDD.n1693 VDD.n1685 0.6405
R16000 VDD.n2042 VDD.n2034 0.6405
R16001 VDD.n2272 VDD.n2264 0.6405
R16002 VDD.n2530 VDD.n2522 0.6405
R16003 VDD.n2788 VDD.n2780 0.6405
R16004 VDD.n3046 VDD.n3038 0.6405
R16005 VDD.n3304 VDD.n3296 0.6405
R16006 VDD.n5634 VDD.n5626 0.6405
R16007 VDD.n5380 VDD.n5372 0.6405
R16008 VDD.n3562 VDD.n3554 0.6405
R16009 VDD.n3820 VDD.n3812 0.6405
R16010 VDD.n4078 VDD.n4070 0.6405
R16011 VDD.n4336 VDD.n4328 0.6405
R16012 VDD.n4594 VDD.n4586 0.6405
R16013 VDD.n4852 VDD.n4844 0.6405
R16014 VDD.n5144 VDD.n5136 0.6405
R16015 VDD.n1688 VDD.n1687 0.590778
R16016 VDD.n2037 VDD.n2036 0.590778
R16017 VDD.n2267 VDD.n2266 0.590778
R16018 VDD.n2525 VDD.n2524 0.590778
R16019 VDD.n2783 VDD.n2782 0.590778
R16020 VDD.n3041 VDD.n3040 0.590778
R16021 VDD.n3299 VDD.n3298 0.590778
R16022 VDD.n5629 VDD.n5628 0.590778
R16023 VDD.n5375 VDD.n5374 0.590778
R16024 VDD.n3557 VDD.n3556 0.590778
R16025 VDD.n3815 VDD.n3814 0.590778
R16026 VDD.n4073 VDD.n4072 0.590778
R16027 VDD.n4331 VDD.n4330 0.590778
R16028 VDD.n4589 VDD.n4588 0.590778
R16029 VDD.n4847 VDD.n4846 0.590778
R16030 VDD.n5139 VDD.n5138 0.590778
R16031 VDD.n5746 VDD.n5745 0.588569
R16032 VDD.n5492 VDD.n5491 0.588569
R16033 VDD.n1805 VDD.n1804 0.580785
R16034 VDD.n2384 VDD.n2383 0.580785
R16035 VDD.n2642 VDD.n2641 0.580785
R16036 VDD.n2900 VDD.n2899 0.580785
R16037 VDD.n3158 VDD.n3157 0.580785
R16038 VDD.n3416 VDD.n3415 0.580785
R16039 VDD.n3674 VDD.n3673 0.580785
R16040 VDD.n3932 VDD.n3931 0.580785
R16041 VDD.n4190 VDD.n4189 0.580785
R16042 VDD.n4448 VDD.n4447 0.580785
R16043 VDD.n4706 VDD.n4705 0.580785
R16044 VDD.n4965 VDD.n4964 0.577251
R16045 VDD.n5115 VDD.n5114 0.577251
R16046 VDD.n1658 VDD.n1657 0.571929
R16047 VDD.n1660 VDD.n1659 0.558536
R16048 VDD.n1112 VDD.n755 0.557954
R16049 VDD.n1597 VDD.n1596 0.557954
R16050 VDD.n1659 VDD.n1658 0.549607
R16051 VDD.n1748 VDD.n1723 0.514389
R16052 VDD.n2097 VDD.n2072 0.514389
R16053 VDD.n2327 VDD.n2302 0.514389
R16054 VDD.n2585 VDD.n2560 0.514389
R16055 VDD.n2843 VDD.n2818 0.514389
R16056 VDD.n3101 VDD.n3076 0.514389
R16057 VDD.n3359 VDD.n3334 0.514389
R16058 VDD.n5689 VDD.n5664 0.514389
R16059 VDD.n5435 VDD.n5410 0.514389
R16060 VDD.n3617 VDD.n3592 0.514389
R16061 VDD.n3875 VDD.n3850 0.514389
R16062 VDD.n4133 VDD.n4108 0.514389
R16063 VDD.n4391 VDD.n4366 0.514389
R16064 VDD.n4649 VDD.n4624 0.514389
R16065 VDD.n4907 VDD.n4882 0.514389
R16066 VDD.n5199 VDD.n5174 0.514389
R16067 VDD.n1977 VDD.n1925 0.5125
R16068 VDD.n1839 VDD.n1826 0.492808
R16069 VDD.n2160 VDD.n2147 0.492808
R16070 VDD.n2418 VDD.n2405 0.492808
R16071 VDD.n2676 VDD.n2663 0.492808
R16072 VDD.n2934 VDD.n2921 0.492808
R16073 VDD.n3192 VDD.n3179 0.492808
R16074 VDD.n3450 VDD.n3437 0.492808
R16075 VDD.n5777 VDD.n5764 0.492808
R16076 VDD.n5523 VDD.n5510 0.492808
R16077 VDD.n3708 VDD.n3695 0.492808
R16078 VDD.n3966 VDD.n3953 0.492808
R16079 VDD.n4224 VDD.n4211 0.492808
R16080 VDD.n4482 VDD.n4469 0.492808
R16081 VDD.n4740 VDD.n4727 0.492808
R16082 VDD.n5001 VDD.n4988 0.492808
R16083 VDD.n5263 VDD.n5250 0.492808
R16084 VDD.n26 VDD 0.476404
R16085 VDD.n343 VDD 0.476404
R16086 VDD.n1686 VDD.n1665 0.471224
R16087 VDD.n2035 VDD.n2014 0.471224
R16088 VDD.n2265 VDD.n2244 0.471224
R16089 VDD.n2523 VDD.n2502 0.471224
R16090 VDD.n2781 VDD.n2760 0.471224
R16091 VDD.n3039 VDD.n3018 0.471224
R16092 VDD.n3297 VDD.n3276 0.471224
R16093 VDD.n5627 VDD.n5606 0.471224
R16094 VDD.n5373 VDD.n5352 0.471224
R16095 VDD.n3555 VDD.n3534 0.471224
R16096 VDD.n3813 VDD.n3792 0.471224
R16097 VDD.n4071 VDD.n4050 0.471224
R16098 VDD.n4329 VDD.n4308 0.471224
R16099 VDD.n4587 VDD.n4566 0.471224
R16100 VDD.n4845 VDD.n4824 0.471224
R16101 VDD.n5137 VDD.n5116 0.471224
R16102 VDD.n1773 VDD.n1666 0.467504
R16103 VDD.n2122 VDD.n2015 0.467504
R16104 VDD.n2352 VDD.n2245 0.467504
R16105 VDD.n2610 VDD.n2503 0.467504
R16106 VDD.n2868 VDD.n2761 0.467504
R16107 VDD.n3126 VDD.n3019 0.467504
R16108 VDD.n3384 VDD.n3277 0.467504
R16109 VDD.n5714 VDD.n5607 0.467504
R16110 VDD.n5460 VDD.n5353 0.467504
R16111 VDD.n3642 VDD.n3535 0.467504
R16112 VDD.n3900 VDD.n3793 0.467504
R16113 VDD.n4158 VDD.n4051 0.467504
R16114 VDD.n4416 VDD.n4309 0.467504
R16115 VDD.n4674 VDD.n4567 0.467504
R16116 VDD.n4932 VDD.n4825 0.467504
R16117 VDD.n5224 VDD.n5117 0.467504
R16118 VDD.n1654 VDD.n1653 0.464786
R16119 VDD.n1637 VDD 0.457643
R16120 VDD.n1661 VDD.n1623 0.424377
R16121 VDD.n1810 VDD 0.411214
R16122 VDD.n2131 VDD 0.411214
R16123 VDD.n2389 VDD 0.411214
R16124 VDD.n2647 VDD 0.411214
R16125 VDD.n2905 VDD 0.411214
R16126 VDD.n3163 VDD 0.411214
R16127 VDD.n3421 VDD 0.411214
R16128 VDD.n5748 VDD 0.411214
R16129 VDD.n5494 VDD 0.411214
R16130 VDD.n3679 VDD 0.411214
R16131 VDD.n3937 VDD 0.411214
R16132 VDD.n4195 VDD 0.411214
R16133 VDD.n4453 VDD 0.411214
R16134 VDD.n4711 VDD 0.411214
R16135 VDD.n4972 VDD 0.411214
R16136 VDD.n5234 VDD 0.411214
R16137 VDD.n1753 VDD.n1752 0.410606
R16138 VDD.n2102 VDD.n2101 0.410606
R16139 VDD.n2332 VDD.n2331 0.410606
R16140 VDD.n2590 VDD.n2589 0.410606
R16141 VDD.n2848 VDD.n2847 0.410606
R16142 VDD.n3106 VDD.n3105 0.410606
R16143 VDD.n3364 VDD.n3363 0.410606
R16144 VDD.n5694 VDD.n5693 0.410606
R16145 VDD.n5440 VDD.n5439 0.410606
R16146 VDD.n3622 VDD.n3621 0.410606
R16147 VDD.n3880 VDD.n3879 0.410606
R16148 VDD.n4138 VDD.n4137 0.410606
R16149 VDD.n4396 VDD.n4395 0.410606
R16150 VDD.n4654 VDD.n4653 0.410606
R16151 VDD.n4912 VDD.n4911 0.410606
R16152 VDD.n5204 VDD.n5203 0.410606
R16153 VDD.n1921 VDD.n1920 0.409102
R16154 VDD.n2242 VDD.n2241 0.409102
R16155 VDD.n2500 VDD.n2499 0.409102
R16156 VDD.n2758 VDD.n2757 0.409102
R16157 VDD.n3016 VDD.n3015 0.409102
R16158 VDD.n3274 VDD.n3273 0.409102
R16159 VDD.n3532 VDD.n3531 0.409102
R16160 VDD.n3790 VDD.n3789 0.409102
R16161 VDD.n4048 VDD.n4047 0.409102
R16162 VDD.n4306 VDD.n4305 0.409102
R16163 VDD.n4564 VDD.n4563 0.409102
R16164 VDD.n4822 VDD.n4821 0.409102
R16165 VDD VDD.n26 0.403703
R16166 VDD VDD.n343 0.403703
R16167 VDD.n4970 VDD.n4969 0.403161
R16168 VDD.n5228 VDD.n5227 0.403161
R16169 VDD.n5232 VDD.n5231 0.403161
R16170 VDD.n1738 VDD.n1737 0.399706
R16171 VDD.n2087 VDD.n2086 0.399706
R16172 VDD.n2317 VDD.n2316 0.399706
R16173 VDD.n2575 VDD.n2574 0.399706
R16174 VDD.n2833 VDD.n2832 0.399706
R16175 VDD.n3091 VDD.n3090 0.399706
R16176 VDD.n3349 VDD.n3348 0.399706
R16177 VDD.n5679 VDD.n5678 0.399706
R16178 VDD.n5425 VDD.n5424 0.399706
R16179 VDD.n3607 VDD.n3606 0.399706
R16180 VDD.n3865 VDD.n3864 0.399706
R16181 VDD.n4123 VDD.n4122 0.399706
R16182 VDD.n4381 VDD.n4380 0.399706
R16183 VDD.n4639 VDD.n4638 0.399706
R16184 VDD.n4897 VDD.n4896 0.399706
R16185 VDD.n5189 VDD.n5188 0.399706
R16186 VDD.n830 VDD.n781 0.399037
R16187 VDD.n379 VDD.n378 0.399037
R16188 VDD.n1749 VDD.n1748 0.398914
R16189 VDD.n2098 VDD.n2097 0.398914
R16190 VDD.n2328 VDD.n2327 0.398914
R16191 VDD.n2586 VDD.n2585 0.398914
R16192 VDD.n2844 VDD.n2843 0.398914
R16193 VDD.n3102 VDD.n3101 0.398914
R16194 VDD.n3360 VDD.n3359 0.398914
R16195 VDD.n5690 VDD.n5689 0.398914
R16196 VDD.n5436 VDD.n5435 0.398914
R16197 VDD.n3618 VDD.n3617 0.398914
R16198 VDD.n3876 VDD.n3875 0.398914
R16199 VDD.n4134 VDD.n4133 0.398914
R16200 VDD.n4392 VDD.n4391 0.398914
R16201 VDD.n4650 VDD.n4649 0.398914
R16202 VDD.n4908 VDD.n4907 0.398914
R16203 VDD.n5200 VDD.n5199 0.398914
R16204 VDD.n1737 VDD.n1723 0.398403
R16205 VDD.n2086 VDD.n2072 0.398403
R16206 VDD.n2316 VDD.n2302 0.398403
R16207 VDD.n2574 VDD.n2560 0.398403
R16208 VDD.n2832 VDD.n2818 0.398403
R16209 VDD.n3090 VDD.n3076 0.398403
R16210 VDD.n3348 VDD.n3334 0.398403
R16211 VDD.n5678 VDD.n5664 0.398403
R16212 VDD.n5424 VDD.n5410 0.398403
R16213 VDD.n3606 VDD.n3592 0.398403
R16214 VDD.n3864 VDD.n3850 0.398403
R16215 VDD.n4122 VDD.n4108 0.398403
R16216 VDD.n4380 VDD.n4366 0.398403
R16217 VDD.n4638 VDD.n4624 0.398403
R16218 VDD.n4896 VDD.n4882 0.398403
R16219 VDD.n5188 VDD.n5174 0.398403
R16220 VDD.n1656 VDD.n1655 0.384429
R16221 VDD.n1807 VDD.n1806 0.3805
R16222 VDD.n2127 VDD.n2126 0.3805
R16223 VDD.n2386 VDD.n2385 0.3805
R16224 VDD.n2644 VDD.n2643 0.3805
R16225 VDD.n2902 VDD.n2901 0.3805
R16226 VDD.n3160 VDD.n3159 0.3805
R16227 VDD.n3418 VDD.n3417 0.3805
R16228 VDD.n3676 VDD.n3675 0.3805
R16229 VDD.n3934 VDD.n3933 0.3805
R16230 VDD.n4192 VDD.n4191 0.3805
R16231 VDD.n4450 VDD.n4449 0.3805
R16232 VDD.n4708 VDD.n4707 0.3805
R16233 VDD.n864 VDD.n863 0.376971
R16234 VDD.n944 VDD.n943 0.376971
R16235 VDD.n1104 VDD.n1103 0.376971
R16236 VDD.n1056 VDD.n1055 0.376971
R16237 VDD.n69 VDD.n68 0.376971
R16238 VDD.n149 VDD.n148 0.376971
R16239 VDD.n309 VDD.n308 0.376971
R16240 VDD.n261 VDD.n260 0.376971
R16241 VDD.n463 VDD.n462 0.376971
R16242 VDD.n543 VDD.n542 0.376971
R16243 VDD.n699 VDD.n698 0.376971
R16244 VDD.n651 VDD.n650 0.376971
R16245 VDD.n1452 VDD.n1451 0.376971
R16246 VDD.n1421 VDD.n1420 0.376971
R16247 VDD.n1266 VDD.n1265 0.376971
R16248 VDD.n1500 VDD.n1499 0.376971
R16249 VDD.n1687 VDD.n1686 0.368458
R16250 VDD.n2036 VDD.n2035 0.368458
R16251 VDD.n2266 VDD.n2265 0.368458
R16252 VDD.n2524 VDD.n2523 0.368458
R16253 VDD.n2782 VDD.n2781 0.368458
R16254 VDD.n3040 VDD.n3039 0.368458
R16255 VDD.n3298 VDD.n3297 0.368458
R16256 VDD.n5628 VDD.n5627 0.368458
R16257 VDD.n5374 VDD.n5373 0.368458
R16258 VDD.n3556 VDD.n3555 0.368458
R16259 VDD.n3814 VDD.n3813 0.368458
R16260 VDD.n4072 VDD.n4071 0.368458
R16261 VDD.n4330 VDD.n4329 0.368458
R16262 VDD.n4588 VDD.n4587 0.368458
R16263 VDD.n4846 VDD.n4845 0.368458
R16264 VDD.n5138 VDD.n5137 0.368458
R16265 VDD.n1688 VDD.n1666 0.361663
R16266 VDD.n2037 VDD.n2015 0.361663
R16267 VDD.n2267 VDD.n2245 0.361663
R16268 VDD.n2525 VDD.n2503 0.361663
R16269 VDD.n2783 VDD.n2761 0.361663
R16270 VDD.n3041 VDD.n3019 0.361663
R16271 VDD.n3299 VDD.n3277 0.361663
R16272 VDD.n5629 VDD.n5607 0.361663
R16273 VDD.n5375 VDD.n5353 0.361663
R16274 VDD.n3557 VDD.n3535 0.361663
R16275 VDD.n3815 VDD.n3793 0.361663
R16276 VDD.n4073 VDD.n4051 0.361663
R16277 VDD.n4331 VDD.n4309 0.361663
R16278 VDD.n4589 VDD.n4567 0.361663
R16279 VDD.n4847 VDD.n4825 0.361663
R16280 VDD.n5139 VDD.n5117 0.361663
R16281 VDD.n1750 VDD.n1749 0.357683
R16282 VDD.n2099 VDD.n2098 0.357683
R16283 VDD.n2329 VDD.n2328 0.357683
R16284 VDD.n2587 VDD.n2586 0.357683
R16285 VDD.n2845 VDD.n2844 0.357683
R16286 VDD.n3103 VDD.n3102 0.357683
R16287 VDD.n3361 VDD.n3360 0.357683
R16288 VDD.n5691 VDD.n5690 0.357683
R16289 VDD.n5437 VDD.n5436 0.357683
R16290 VDD.n3619 VDD.n3618 0.357683
R16291 VDD.n3877 VDD.n3876 0.357683
R16292 VDD.n4135 VDD.n4134 0.357683
R16293 VDD.n4393 VDD.n4392 0.357683
R16294 VDD.n4651 VDD.n4650 0.357683
R16295 VDD.n4909 VDD.n4908 0.357683
R16296 VDD.n5201 VDD.n5200 0.357683
R16297 VDD.n1734 VDD.n1732 0.356056
R16298 VDD.n2083 VDD.n2081 0.356056
R16299 VDD.n2313 VDD.n2311 0.356056
R16300 VDD.n2571 VDD.n2569 0.356056
R16301 VDD.n2829 VDD.n2827 0.356056
R16302 VDD.n3087 VDD.n3085 0.356056
R16303 VDD.n3345 VDD.n3343 0.356056
R16304 VDD.n5675 VDD.n5673 0.356056
R16305 VDD.n5421 VDD.n5419 0.356056
R16306 VDD.n3603 VDD.n3601 0.356056
R16307 VDD.n3861 VDD.n3859 0.356056
R16308 VDD.n4119 VDD.n4117 0.356056
R16309 VDD.n4377 VDD.n4375 0.356056
R16310 VDD.n4635 VDD.n4633 0.356056
R16311 VDD.n4893 VDD.n4891 0.356056
R16312 VDD.n5185 VDD.n5183 0.356056
R16313 VDD.n35 VDD.n34 0.35558
R16314 VDD.n352 VDD.n351 0.35558
R16315 VDD.n1836 VDD 0.355332
R16316 VDD.n2157 VDD 0.355332
R16317 VDD.n2415 VDD 0.355332
R16318 VDD.n2673 VDD 0.355332
R16319 VDD.n2931 VDD 0.355332
R16320 VDD.n3189 VDD 0.355332
R16321 VDD.n3447 VDD 0.355332
R16322 VDD.n5774 VDD 0.355332
R16323 VDD.n5520 VDD 0.355332
R16324 VDD.n3705 VDD 0.355332
R16325 VDD.n3963 VDD 0.355332
R16326 VDD.n4221 VDD 0.355332
R16327 VDD.n4479 VDD 0.355332
R16328 VDD.n4737 VDD 0.355332
R16329 VDD.n4998 VDD 0.355332
R16330 VDD.n5260 VDD 0.355332
R16331 VDD.n1918 VDD.n1887 0.349136
R16332 VDD.n2239 VDD.n2208 0.349136
R16333 VDD.n2497 VDD.n2466 0.349136
R16334 VDD.n2755 VDD.n2724 0.349136
R16335 VDD.n3013 VDD.n2982 0.349136
R16336 VDD.n3271 VDD.n3240 0.349136
R16337 VDD.n3529 VDD.n3498 0.349136
R16338 VDD.n5856 VDD.n5825 0.349136
R16339 VDD.n5602 VDD.n5571 0.349136
R16340 VDD.n3787 VDD.n3756 0.349136
R16341 VDD.n4045 VDD.n4014 0.349136
R16342 VDD.n4303 VDD.n4272 0.349136
R16343 VDD.n4561 VDD.n4530 0.349136
R16344 VDD.n4819 VDD.n4788 0.349136
R16345 VDD.n5080 VDD.n5049 0.349136
R16346 VDD.n5342 VDD.n5311 0.349136
R16347 VDD.n0 VDD 0.340206
R16348 VDD.n317 VDD 0.340206
R16349 VDD.n1692 VDD.n1687 0.340142
R16350 VDD.n2041 VDD.n2036 0.340142
R16351 VDD.n2271 VDD.n2266 0.340142
R16352 VDD.n2529 VDD.n2524 0.340142
R16353 VDD.n2787 VDD.n2782 0.340142
R16354 VDD.n3045 VDD.n3040 0.340142
R16355 VDD.n3303 VDD.n3298 0.340142
R16356 VDD.n5633 VDD.n5628 0.340142
R16357 VDD.n5379 VDD.n5374 0.340142
R16358 VDD.n3561 VDD.n3556 0.340142
R16359 VDD.n3819 VDD.n3814 0.340142
R16360 VDD.n4077 VDD.n4072 0.340142
R16361 VDD.n4335 VDD.n4330 0.340142
R16362 VDD.n4593 VDD.n4588 0.340142
R16363 VDD.n4851 VDD.n4846 0.340142
R16364 VDD.n5143 VDD.n5138 0.340142
R16365 VDD.n1283 VDD 0.330819
R16366 VDD VDD.n5870 0.330551
R16367 VDD.n1768 VDD.n1671 0.3205
R16368 VDD.n1693 VDD.n1684 0.3205
R16369 VDD.n2117 VDD.n2020 0.3205
R16370 VDD.n2042 VDD.n2033 0.3205
R16371 VDD.n2347 VDD.n2250 0.3205
R16372 VDD.n2272 VDD.n2263 0.3205
R16373 VDD.n2605 VDD.n2508 0.3205
R16374 VDD.n2530 VDD.n2521 0.3205
R16375 VDD.n2863 VDD.n2766 0.3205
R16376 VDD.n2788 VDD.n2779 0.3205
R16377 VDD.n3121 VDD.n3024 0.3205
R16378 VDD.n3046 VDD.n3037 0.3205
R16379 VDD.n3379 VDD.n3282 0.3205
R16380 VDD.n3304 VDD.n3295 0.3205
R16381 VDD.n5709 VDD.n5612 0.3205
R16382 VDD.n5634 VDD.n5625 0.3205
R16383 VDD.n5455 VDD.n5358 0.3205
R16384 VDD.n5380 VDD.n5371 0.3205
R16385 VDD.n3637 VDD.n3540 0.3205
R16386 VDD.n3562 VDD.n3553 0.3205
R16387 VDD.n3895 VDD.n3798 0.3205
R16388 VDD.n3820 VDD.n3811 0.3205
R16389 VDD.n4153 VDD.n4056 0.3205
R16390 VDD.n4078 VDD.n4069 0.3205
R16391 VDD.n4411 VDD.n4314 0.3205
R16392 VDD.n4336 VDD.n4327 0.3205
R16393 VDD.n4669 VDD.n4572 0.3205
R16394 VDD.n4594 VDD.n4585 0.3205
R16395 VDD.n4927 VDD.n4830 0.3205
R16396 VDD.n4852 VDD.n4843 0.3205
R16397 VDD.n5219 VDD.n5122 0.3205
R16398 VDD.n5144 VDD.n5135 0.3205
R16399 VDD.n1919 VDD.n1918 0.314572
R16400 VDD.n2240 VDD.n2239 0.314572
R16401 VDD.n2498 VDD.n2497 0.314572
R16402 VDD.n2756 VDD.n2755 0.314572
R16403 VDD.n3014 VDD.n3013 0.314572
R16404 VDD.n3272 VDD.n3271 0.314572
R16405 VDD.n3530 VDD.n3529 0.314572
R16406 VDD.n5857 VDD.n5856 0.314572
R16407 VDD.n5603 VDD.n5602 0.314572
R16408 VDD.n3788 VDD.n3787 0.314572
R16409 VDD.n4046 VDD.n4045 0.314572
R16410 VDD.n4304 VDD.n4303 0.314572
R16411 VDD.n4562 VDD.n4561 0.314572
R16412 VDD.n4820 VDD.n4819 0.314572
R16413 VDD.n5081 VDD.n5080 0.314572
R16414 VDD.n5343 VDD.n5342 0.314572
R16415 VDD.n1874 VDD.n1873 0.311403
R16416 VDD.n2195 VDD.n2194 0.311403
R16417 VDD.n2453 VDD.n2452 0.311403
R16418 VDD.n2711 VDD.n2710 0.311403
R16419 VDD.n2969 VDD.n2968 0.311403
R16420 VDD.n3227 VDD.n3226 0.311403
R16421 VDD.n3485 VDD.n3484 0.311403
R16422 VDD.n5812 VDD.n5811 0.311403
R16423 VDD.n5558 VDD.n5557 0.311403
R16424 VDD.n3743 VDD.n3742 0.311403
R16425 VDD.n4001 VDD.n4000 0.311403
R16426 VDD.n4259 VDD.n4258 0.311403
R16427 VDD.n4517 VDD.n4516 0.311403
R16428 VDD.n4775 VDD.n4774 0.311403
R16429 VDD.n5036 VDD.n5035 0.311403
R16430 VDD.n5298 VDD.n5297 0.311403
R16431 VDD.n1691 VDD.n1690 0.296036
R16432 VDD.n2040 VDD.n2039 0.296036
R16433 VDD.n2270 VDD.n2269 0.296036
R16434 VDD.n2528 VDD.n2527 0.296036
R16435 VDD.n2786 VDD.n2785 0.296036
R16436 VDD.n3044 VDD.n3043 0.296036
R16437 VDD.n3302 VDD.n3301 0.296036
R16438 VDD.n5632 VDD.n5631 0.296036
R16439 VDD.n5378 VDD.n5377 0.296036
R16440 VDD.n3560 VDD.n3559 0.296036
R16441 VDD.n3818 VDD.n3817 0.296036
R16442 VDD.n4076 VDD.n4075 0.296036
R16443 VDD.n4334 VDD.n4333 0.296036
R16444 VDD.n4592 VDD.n4591 0.296036
R16445 VDD.n4850 VDD.n4849 0.296036
R16446 VDD.n5142 VDD.n5141 0.296036
R16447 VDD.n1650 VDD 0.278761
R16448 VDD.n5083 VDD.n4823 0.27093
R16449 VDD.n5869 VDD.n1181 0.261949
R16450 VDD.n1747 VDD.n1724 0.261214
R16451 VDD.n1727 VDD.n1726 0.261214
R16452 VDD.n2096 VDD.n2073 0.261214
R16453 VDD.n2076 VDD.n2075 0.261214
R16454 VDD.n2326 VDD.n2303 0.261214
R16455 VDD.n2306 VDD.n2305 0.261214
R16456 VDD.n2584 VDD.n2561 0.261214
R16457 VDD.n2564 VDD.n2563 0.261214
R16458 VDD.n2842 VDD.n2819 0.261214
R16459 VDD.n2822 VDD.n2821 0.261214
R16460 VDD.n3100 VDD.n3077 0.261214
R16461 VDD.n3080 VDD.n3079 0.261214
R16462 VDD.n3358 VDD.n3335 0.261214
R16463 VDD.n3338 VDD.n3337 0.261214
R16464 VDD.n5688 VDD.n5665 0.261214
R16465 VDD.n5668 VDD.n5667 0.261214
R16466 VDD.n5434 VDD.n5411 0.261214
R16467 VDD.n5414 VDD.n5413 0.261214
R16468 VDD.n3616 VDD.n3593 0.261214
R16469 VDD.n3596 VDD.n3595 0.261214
R16470 VDD.n3874 VDD.n3851 0.261214
R16471 VDD.n3854 VDD.n3853 0.261214
R16472 VDD.n4132 VDD.n4109 0.261214
R16473 VDD.n4112 VDD.n4111 0.261214
R16474 VDD.n4390 VDD.n4367 0.261214
R16475 VDD.n4370 VDD.n4369 0.261214
R16476 VDD.n4648 VDD.n4625 0.261214
R16477 VDD.n4628 VDD.n4627 0.261214
R16478 VDD.n4906 VDD.n4883 0.261214
R16479 VDD.n4886 VDD.n4885 0.261214
R16480 VDD.n5198 VDD.n5175 0.261214
R16481 VDD.n5178 VDD.n5177 0.261214
R16482 VDD.n1745 VDD.n1725 0.2565
R16483 VDD.n2094 VDD.n2074 0.2565
R16484 VDD.n2324 VDD.n2304 0.2565
R16485 VDD.n2582 VDD.n2562 0.2565
R16486 VDD.n2840 VDD.n2820 0.2565
R16487 VDD.n3098 VDD.n3078 0.2565
R16488 VDD.n3356 VDD.n3336 0.2565
R16489 VDD.n5686 VDD.n5666 0.2565
R16490 VDD.n5432 VDD.n5412 0.2565
R16491 VDD.n3614 VDD.n3594 0.2565
R16492 VDD.n3872 VDD.n3852 0.2565
R16493 VDD.n4130 VDD.n4110 0.2565
R16494 VDD.n4388 VDD.n4368 0.2565
R16495 VDD.n4646 VDD.n4626 0.2565
R16496 VDD.n4904 VDD.n4884 0.2565
R16497 VDD.n5196 VDD.n5176 0.2565
R16498 VDD.n1736 VDD.n1735 0.251889
R16499 VDD.n2085 VDD.n2084 0.251889
R16500 VDD.n2315 VDD.n2314 0.251889
R16501 VDD.n2573 VDD.n2572 0.251889
R16502 VDD.n2831 VDD.n2830 0.251889
R16503 VDD.n3089 VDD.n3088 0.251889
R16504 VDD.n3347 VDD.n3346 0.251889
R16505 VDD.n5677 VDD.n5676 0.251889
R16506 VDD.n5423 VDD.n5422 0.251889
R16507 VDD.n3605 VDD.n3604 0.251889
R16508 VDD.n3863 VDD.n3862 0.251889
R16509 VDD.n4121 VDD.n4120 0.251889
R16510 VDD.n4379 VDD.n4378 0.251889
R16511 VDD.n4637 VDD.n4636 0.251889
R16512 VDD.n4895 VDD.n4894 0.251889
R16513 VDD.n5187 VDD.n5186 0.251889
R16514 VDD.n1754 VDD.n1719 0.248103
R16515 VDD.n2103 VDD.n2068 0.248103
R16516 VDD.n2333 VDD.n2298 0.248103
R16517 VDD.n2591 VDD.n2556 0.248103
R16518 VDD.n2849 VDD.n2814 0.248103
R16519 VDD.n3107 VDD.n3072 0.248103
R16520 VDD.n3365 VDD.n3330 0.248103
R16521 VDD.n5695 VDD.n5660 0.248103
R16522 VDD.n5441 VDD.n5406 0.248103
R16523 VDD.n3623 VDD.n3588 0.248103
R16524 VDD.n3881 VDD.n3846 0.248103
R16525 VDD.n4139 VDD.n4104 0.248103
R16526 VDD.n4397 VDD.n4362 0.248103
R16527 VDD.n4655 VDD.n4620 0.248103
R16528 VDD.n4913 VDD.n4878 0.248103
R16529 VDD.n5205 VDD.n5170 0.248103
R16530 VDD.n1770 VDD.n1668 0.247868
R16531 VDD.n2119 VDD.n2017 0.247868
R16532 VDD.n2349 VDD.n2247 0.247868
R16533 VDD.n2607 VDD.n2505 0.247868
R16534 VDD.n2865 VDD.n2763 0.247868
R16535 VDD.n3123 VDD.n3021 0.247868
R16536 VDD.n3381 VDD.n3279 0.247868
R16537 VDD.n5711 VDD.n5609 0.247868
R16538 VDD.n5457 VDD.n5355 0.247868
R16539 VDD.n3639 VDD.n3537 0.247868
R16540 VDD.n3897 VDD.n3795 0.247868
R16541 VDD.n4155 VDD.n4053 0.247868
R16542 VDD.n4413 VDD.n4311 0.247868
R16543 VDD.n4671 VDD.n4569 0.247868
R16544 VDD.n4929 VDD.n4827 0.247868
R16545 VDD.n5221 VDD.n5119 0.247868
R16546 VDD.n1125 VDD.n1124 0.240091
R16547 VDD.n1191 VDD.n1190 0.240091
R16548 VDD.n1738 VDD.n1721 0.232755
R16549 VDD.n2087 VDD.n2070 0.232755
R16550 VDD.n2317 VDD.n2300 0.232755
R16551 VDD.n2575 VDD.n2558 0.232755
R16552 VDD.n2833 VDD.n2816 0.232755
R16553 VDD.n3091 VDD.n3074 0.232755
R16554 VDD.n3349 VDD.n3332 0.232755
R16555 VDD.n5679 VDD.n5662 0.232755
R16556 VDD.n5425 VDD.n5408 0.232755
R16557 VDD.n3607 VDD.n3590 0.232755
R16558 VDD.n3865 VDD.n3848 0.232755
R16559 VDD.n4123 VDD.n4106 0.232755
R16560 VDD.n4381 VDD.n4364 0.232755
R16561 VDD.n4639 VDD.n4622 0.232755
R16562 VDD.n4897 VDD.n4880 0.232755
R16563 VDD.n5189 VDD.n5172 0.232755
R16564 VDD.n1953 VDD.n1952 0.224662
R16565 VDD.n1730 VDD.n1722 0.217167
R16566 VDD.n2079 VDD.n2071 0.217167
R16567 VDD.n2309 VDD.n2301 0.217167
R16568 VDD.n2567 VDD.n2559 0.217167
R16569 VDD.n2825 VDD.n2817 0.217167
R16570 VDD.n3083 VDD.n3075 0.217167
R16571 VDD.n3341 VDD.n3333 0.217167
R16572 VDD.n5671 VDD.n5663 0.217167
R16573 VDD.n5417 VDD.n5409 0.217167
R16574 VDD.n3599 VDD.n3591 0.217167
R16575 VDD.n3857 VDD.n3849 0.217167
R16576 VDD.n4115 VDD.n4107 0.217167
R16577 VDD.n4373 VDD.n4365 0.217167
R16578 VDD.n4631 VDD.n4623 0.217167
R16579 VDD.n4889 VDD.n4881 0.217167
R16580 VDD.n5181 VDD.n5173 0.217167
R16581 VDD.n829 VDD.n828 0.212557
R16582 VDD.n427 VDD.n426 0.212557
R16583 VDD.n724 VDD.n723 0.211096
R16584 VDD.n1565 VDD.n1564 0.211096
R16585 VDD.n798 VDD 0.210222
R16586 VDD.n396 VDD 0.210222
R16587 VDD.n1702 VDD.n1701 0.204667
R16588 VDD.n2051 VDD.n2050 0.204667
R16589 VDD.n2281 VDD.n2280 0.204667
R16590 VDD.n2539 VDD.n2538 0.204667
R16591 VDD.n2797 VDD.n2796 0.204667
R16592 VDD.n3055 VDD.n3054 0.204667
R16593 VDD.n3313 VDD.n3312 0.204667
R16594 VDD.n5643 VDD.n5642 0.204667
R16595 VDD.n5389 VDD.n5388 0.204667
R16596 VDD.n3571 VDD.n3570 0.204667
R16597 VDD.n3829 VDD.n3828 0.204667
R16598 VDD.n4087 VDD.n4086 0.204667
R16599 VDD.n4345 VDD.n4344 0.204667
R16600 VDD.n4603 VDD.n4602 0.204667
R16601 VDD.n4861 VDD.n4860 0.204667
R16602 VDD.n5153 VDD.n5152 0.204667
R16603 VDD.n1662 VDD 0.2005
R16604 VDD.n1703 VDD.n1667 0.199111
R16605 VDD.n2052 VDD.n2016 0.199111
R16606 VDD.n2282 VDD.n2246 0.199111
R16607 VDD.n2540 VDD.n2504 0.199111
R16608 VDD.n2798 VDD.n2762 0.199111
R16609 VDD.n3056 VDD.n3020 0.199111
R16610 VDD.n3314 VDD.n3278 0.199111
R16611 VDD.n5644 VDD.n5608 0.199111
R16612 VDD.n5390 VDD.n5354 0.199111
R16613 VDD.n3572 VDD.n3536 0.199111
R16614 VDD.n3830 VDD.n3794 0.199111
R16615 VDD.n4088 VDD.n4052 0.199111
R16616 VDD.n4346 VDD.n4310 0.199111
R16617 VDD.n4604 VDD.n4568 0.199111
R16618 VDD.n4862 VDD.n4826 0.199111
R16619 VDD.n5154 VDD.n5118 0.199111
R16620 VDD.n28 VDD 0.196824
R16621 VDD.n345 VDD 0.196824
R16622 VDD.n1816 VDD.n1815 0.192557
R16623 VDD.n2137 VDD.n2136 0.192557
R16624 VDD.n2395 VDD.n2394 0.192557
R16625 VDD.n2653 VDD.n2652 0.192557
R16626 VDD.n2911 VDD.n2910 0.192557
R16627 VDD.n3169 VDD.n3168 0.192557
R16628 VDD.n3427 VDD.n3426 0.192557
R16629 VDD.n5754 VDD.n5753 0.192557
R16630 VDD.n5500 VDD.n5499 0.192557
R16631 VDD.n3685 VDD.n3684 0.192557
R16632 VDD.n3943 VDD.n3942 0.192557
R16633 VDD.n4201 VDD.n4200 0.192557
R16634 VDD.n4459 VDD.n4458 0.192557
R16635 VDD.n4717 VDD.n4716 0.192557
R16636 VDD.n4978 VDD.n4977 0.192557
R16637 VDD.n5240 VDD.n5239 0.192557
R16638 VDD.n1811 VDD.n1810 0.192167
R16639 VDD.n2132 VDD.n2131 0.192167
R16640 VDD.n2390 VDD.n2389 0.192167
R16641 VDD.n2648 VDD.n2647 0.192167
R16642 VDD.n2906 VDD.n2905 0.192167
R16643 VDD.n3164 VDD.n3163 0.192167
R16644 VDD.n3422 VDD.n3421 0.192167
R16645 VDD.n5749 VDD.n5748 0.192167
R16646 VDD.n5495 VDD.n5494 0.192167
R16647 VDD.n3680 VDD.n3679 0.192167
R16648 VDD.n3938 VDD.n3937 0.192167
R16649 VDD.n4196 VDD.n4195 0.192167
R16650 VDD.n4454 VDD.n4453 0.192167
R16651 VDD.n4712 VDD.n4711 0.192167
R16652 VDD.n4973 VDD.n4972 0.192167
R16653 VDD.n5235 VDD.n5234 0.192167
R16654 VDD.n5870 VDD.n1180 0.189
R16655 VDD.n34 VDD.n33 0.183651
R16656 VDD.n351 VDD.n350 0.183651
R16657 VDD.n1804 VDD.n1776 0.180841
R16658 VDD.n2012 VDD.n1984 0.180841
R16659 VDD.n2383 VDD.n2355 0.180841
R16660 VDD.n2641 VDD.n2613 0.180841
R16661 VDD.n2899 VDD.n2871 0.180841
R16662 VDD.n3157 VDD.n3129 0.180841
R16663 VDD.n3415 VDD.n3387 0.180841
R16664 VDD.n5745 VDD.n5717 0.180841
R16665 VDD.n5491 VDD.n5463 0.180841
R16666 VDD.n3673 VDD.n3645 0.180841
R16667 VDD.n3931 VDD.n3903 0.180841
R16668 VDD.n4189 VDD.n4161 0.180841
R16669 VDD.n4447 VDD.n4419 0.180841
R16670 VDD.n4705 VDD.n4677 0.180841
R16671 VDD.n4964 VDD.n4936 0.180841
R16672 VDD.n5114 VDD.n5086 0.180841
R16673 VDD.n828 VDD.n827 0.175873
R16674 VDD.n426 VDD.n425 0.175873
R16675 VDD.n1599 VDD.n1548 0.168948
R16676 VDD.n1760 VDD.n1759 0.164944
R16677 VDD.n1759 VDD.n1711 0.164944
R16678 VDD.n2109 VDD.n2108 0.164944
R16679 VDD.n2108 VDD.n2060 0.164944
R16680 VDD.n2339 VDD.n2338 0.164944
R16681 VDD.n2338 VDD.n2290 0.164944
R16682 VDD.n2597 VDD.n2596 0.164944
R16683 VDD.n2596 VDD.n2548 0.164944
R16684 VDD.n2855 VDD.n2854 0.164944
R16685 VDD.n2854 VDD.n2806 0.164944
R16686 VDD.n3113 VDD.n3112 0.164944
R16687 VDD.n3112 VDD.n3064 0.164944
R16688 VDD.n3371 VDD.n3370 0.164944
R16689 VDD.n3370 VDD.n3322 0.164944
R16690 VDD.n5701 VDD.n5700 0.164944
R16691 VDD.n5700 VDD.n5652 0.164944
R16692 VDD.n5447 VDD.n5446 0.164944
R16693 VDD.n5446 VDD.n5398 0.164944
R16694 VDD.n3629 VDD.n3628 0.164944
R16695 VDD.n3628 VDD.n3580 0.164944
R16696 VDD.n3887 VDD.n3886 0.164944
R16697 VDD.n3886 VDD.n3838 0.164944
R16698 VDD.n4145 VDD.n4144 0.164944
R16699 VDD.n4144 VDD.n4096 0.164944
R16700 VDD.n4403 VDD.n4402 0.164944
R16701 VDD.n4402 VDD.n4354 0.164944
R16702 VDD.n4661 VDD.n4660 0.164944
R16703 VDD.n4660 VDD.n4612 0.164944
R16704 VDD.n4919 VDD.n4918 0.164944
R16705 VDD.n4918 VDD.n4870 0.164944
R16706 VDD.n5211 VDD.n5210 0.164944
R16707 VDD.n5210 VDD.n5162 0.164944
R16708 VDD.n1710 VDD.n1709 0.159358
R16709 VDD.n2059 VDD.n2058 0.159358
R16710 VDD.n2289 VDD.n2288 0.159358
R16711 VDD.n2547 VDD.n2546 0.159358
R16712 VDD.n2805 VDD.n2804 0.159358
R16713 VDD.n3063 VDD.n3062 0.159358
R16714 VDD.n3321 VDD.n3320 0.159358
R16715 VDD.n5651 VDD.n5650 0.159358
R16716 VDD.n5397 VDD.n5396 0.159358
R16717 VDD.n3579 VDD.n3578 0.159358
R16718 VDD.n3837 VDD.n3836 0.159358
R16719 VDD.n4095 VDD.n4094 0.159358
R16720 VDD.n4353 VDD.n4352 0.159358
R16721 VDD.n4611 VDD.n4610 0.159358
R16722 VDD.n4869 VDD.n4868 0.159358
R16723 VDD.n5161 VDD.n5160 0.159358
R16724 VDD.n1709 VDD.n1708 0.15889
R16725 VDD.n2058 VDD.n2057 0.15889
R16726 VDD.n2288 VDD.n2287 0.15889
R16727 VDD.n2546 VDD.n2545 0.15889
R16728 VDD.n2804 VDD.n2803 0.15889
R16729 VDD.n3062 VDD.n3061 0.15889
R16730 VDD.n3320 VDD.n3319 0.15889
R16731 VDD.n5650 VDD.n5649 0.15889
R16732 VDD.n5396 VDD.n5395 0.15889
R16733 VDD.n3578 VDD.n3577 0.15889
R16734 VDD.n3836 VDD.n3835 0.15889
R16735 VDD.n4094 VDD.n4093 0.15889
R16736 VDD.n4352 VDD.n4351 0.15889
R16737 VDD.n4610 VDD.n4609 0.15889
R16738 VDD.n4868 VDD.n4867 0.15889
R16739 VDD.n5160 VDD.n5159 0.15889
R16740 VDD.n755 VDD.n754 0.155541
R16741 VDD.n1596 VDD.n1595 0.155541
R16742 VDD.n27 VDD 0.145087
R16743 VDD.n344 VDD 0.145087
R16744 VDD VDD.n1137 0.137071
R16745 VDD VDD.n1203 0.137071
R16746 VDD.n5868 VDD.n1663 0.134625
R16747 VDD.n1169 VDD.n1168 0.128415
R16748 VDD.n1235 VDD.n1234 0.128415
R16749 VDD.n781 VDD.n779 0.120987
R16750 VDD.n378 VDD.n376 0.120987
R16751 VDD.n1170 VDD.n1169 0.119283
R16752 VDD.n1236 VDD.n1235 0.119283
R16753 VDD.n1774 VDD.n1773 0.117306
R16754 VDD.n2123 VDD.n2122 0.117306
R16755 VDD.n2353 VDD.n2352 0.117306
R16756 VDD.n2611 VDD.n2610 0.117306
R16757 VDD.n2869 VDD.n2868 0.117306
R16758 VDD.n3127 VDD.n3126 0.117306
R16759 VDD.n3385 VDD.n3384 0.117306
R16760 VDD.n5715 VDD.n5714 0.117306
R16761 VDD.n5461 VDD.n5460 0.117306
R16762 VDD.n3643 VDD.n3642 0.117306
R16763 VDD.n3901 VDD.n3900 0.117306
R16764 VDD.n4159 VDD.n4158 0.117306
R16765 VDD.n4417 VDD.n4416 0.117306
R16766 VDD.n4675 VDD.n4674 0.117306
R16767 VDD.n4933 VDD.n4932 0.117306
R16768 VDD.n5225 VDD.n5224 0.117306
R16769 VDD.n1111 VDD.n1110 0.116581
R16770 VDD.n1165 VDD.n1164 0.1155
R16771 VDD.n1164 VDD.n1162 0.1155
R16772 VDD.n1159 VDD.n1158 0.1155
R16773 VDD.n1158 VDD.n1156 0.1155
R16774 VDD.n1153 VDD.n1152 0.1155
R16775 VDD.n1152 VDD.n1150 0.1155
R16776 VDD.n1147 VDD.n1146 0.1155
R16777 VDD.n1146 VDD.n1144 0.1155
R16778 VDD.n1231 VDD.n1230 0.1155
R16779 VDD.n1230 VDD.n1228 0.1155
R16780 VDD.n1225 VDD.n1224 0.1155
R16781 VDD.n1224 VDD.n1222 0.1155
R16782 VDD.n1219 VDD.n1218 0.1155
R16783 VDD.n1218 VDD.n1216 0.1155
R16784 VDD.n1213 VDD.n1212 0.1155
R16785 VDD.n1212 VDD.n1210 0.1155
R16786 VDD.n5858 VDD.n5746 0.109623
R16787 VDD.n5604 VDD.n5492 0.109623
R16788 VDD.n1179 VDD 0.109094
R16789 VDD.n1245 VDD 0.109094
R16790 VDD.n1179 VDD.n1178 0.107922
R16791 VDD.n1245 VDD.n1244 0.107922
R16792 VDD.n1948 VDD.n1947 0.107375
R16793 VDD.n1952 VDD.n1948 0.107375
R16794 VDD.n1856 VDD.n1843 0.104784
R16795 VDD.n1857 VDD.n1856 0.104784
R16796 VDD.n2177 VDD.n2164 0.104784
R16797 VDD.n2178 VDD.n2177 0.104784
R16798 VDD.n2435 VDD.n2422 0.104784
R16799 VDD.n2436 VDD.n2435 0.104784
R16800 VDD.n2693 VDD.n2680 0.104784
R16801 VDD.n2694 VDD.n2693 0.104784
R16802 VDD.n2951 VDD.n2938 0.104784
R16803 VDD.n2952 VDD.n2951 0.104784
R16804 VDD.n3209 VDD.n3196 0.104784
R16805 VDD.n3210 VDD.n3209 0.104784
R16806 VDD.n3467 VDD.n3454 0.104784
R16807 VDD.n3468 VDD.n3467 0.104784
R16808 VDD.n5794 VDD.n5781 0.104784
R16809 VDD.n5795 VDD.n5794 0.104784
R16810 VDD.n5540 VDD.n5527 0.104784
R16811 VDD.n5541 VDD.n5540 0.104784
R16812 VDD.n3725 VDD.n3712 0.104784
R16813 VDD.n3726 VDD.n3725 0.104784
R16814 VDD.n3983 VDD.n3970 0.104784
R16815 VDD.n3984 VDD.n3983 0.104784
R16816 VDD.n4241 VDD.n4228 0.104784
R16817 VDD.n4242 VDD.n4241 0.104784
R16818 VDD.n4499 VDD.n4486 0.104784
R16819 VDD.n4500 VDD.n4499 0.104784
R16820 VDD.n4757 VDD.n4744 0.104784
R16821 VDD.n4758 VDD.n4757 0.104784
R16822 VDD.n5018 VDD.n5005 0.104784
R16823 VDD.n5019 VDD.n5018 0.104784
R16824 VDD.n5280 VDD.n5267 0.104784
R16825 VDD.n5281 VDD.n5280 0.104784
R16826 VDD.n1114 VDD.n707 0.102139
R16827 VDD.n1975 VDD.n1974 0.100461
R16828 VDD.n1944 VDD.n1940 0.100461
R16829 VDD.n1974 VDD.n1973 0.0999624
R16830 VDD.n1958 VDD.n1940 0.0999624
R16831 VDD.n1873 VDD.n1842 0.0972991
R16832 VDD.n2194 VDD.n2163 0.0972991
R16833 VDD.n2452 VDD.n2421 0.0972991
R16834 VDD.n2710 VDD.n2679 0.0972991
R16835 VDD.n2968 VDD.n2937 0.0972991
R16836 VDD.n3226 VDD.n3195 0.0972991
R16837 VDD.n3484 VDD.n3453 0.0972991
R16838 VDD.n5811 VDD.n5780 0.0972991
R16839 VDD.n5557 VDD.n5526 0.0972991
R16840 VDD.n3742 VDD.n3711 0.0972991
R16841 VDD.n4000 VDD.n3969 0.0972991
R16842 VDD.n4258 VDD.n4227 0.0972991
R16843 VDD.n4516 VDD.n4485 0.0972991
R16844 VDD.n4774 VDD.n4743 0.0972991
R16845 VDD.n5035 VDD.n5004 0.0972991
R16846 VDD.n5297 VDD.n5266 0.0972991
R16847 VDD.n1811 VDD 0.0963333
R16848 VDD.n2132 VDD 0.0963333
R16849 VDD.n2390 VDD 0.0963333
R16850 VDD.n2648 VDD 0.0963333
R16851 VDD.n2906 VDD 0.0963333
R16852 VDD.n3164 VDD 0.0963333
R16853 VDD.n3422 VDD 0.0963333
R16854 VDD.n5749 VDD 0.0963333
R16855 VDD.n5495 VDD 0.0963333
R16856 VDD.n3680 VDD 0.0963333
R16857 VDD.n3938 VDD 0.0963333
R16858 VDD.n4196 VDD 0.0963333
R16859 VDD.n4454 VDD 0.0963333
R16860 VDD.n4712 VDD 0.0963333
R16861 VDD.n4973 VDD 0.0963333
R16862 VDD.n5235 VDD 0.0963333
R16863 VDD.n1935 VDD.n1934 0.0960166
R16864 VDD.n1936 VDD.n1935 0.095518
R16865 VDD.n1170 VDD 0.0950313
R16866 VDD.n1236 VDD 0.0950313
R16867 VDD.n1841 VDD 0.0948131
R16868 VDD.n2162 VDD 0.0948131
R16869 VDD.n2420 VDD 0.0948131
R16870 VDD.n2678 VDD 0.0948131
R16871 VDD.n2936 VDD 0.0948131
R16872 VDD.n3194 VDD 0.0948131
R16873 VDD.n3452 VDD 0.0948131
R16874 VDD.n5779 VDD 0.0948131
R16875 VDD.n5525 VDD 0.0948131
R16876 VDD.n3710 VDD 0.0948131
R16877 VDD.n3968 VDD 0.0948131
R16878 VDD.n4226 VDD 0.0948131
R16879 VDD.n4484 VDD 0.0948131
R16880 VDD.n4742 VDD 0.0948131
R16881 VDD.n5003 VDD 0.0948131
R16882 VDD.n5265 VDD 0.0948131
R16883 VDD.n1875 VDD.n1817 0.0945934
R16884 VDD.n2196 VDD.n2138 0.0945934
R16885 VDD.n2454 VDD.n2396 0.0945934
R16886 VDD.n2712 VDD.n2654 0.0945934
R16887 VDD.n2970 VDD.n2912 0.0945934
R16888 VDD.n3228 VDD.n3170 0.0945934
R16889 VDD.n3486 VDD.n3428 0.0945934
R16890 VDD.n5813 VDD.n5755 0.0945934
R16891 VDD.n5559 VDD.n5501 0.0945934
R16892 VDD.n3744 VDD.n3686 0.0945934
R16893 VDD.n4002 VDD.n3944 0.0945934
R16894 VDD.n4260 VDD.n4202 0.0945934
R16895 VDD.n4518 VDD.n4460 0.0945934
R16896 VDD.n4776 VDD.n4718 0.0945934
R16897 VDD.n5037 VDD.n4979 0.0945934
R16898 VDD.n5299 VDD.n5241 0.0945934
R16899 VDD.n1836 VDD 0.0902606
R16900 VDD.n2157 VDD 0.0902606
R16901 VDD.n2415 VDD 0.0902606
R16902 VDD.n2673 VDD 0.0902606
R16903 VDD.n2931 VDD 0.0902606
R16904 VDD.n3189 VDD 0.0902606
R16905 VDD.n3447 VDD 0.0902606
R16906 VDD.n5774 VDD 0.0902606
R16907 VDD.n5520 VDD 0.0902606
R16908 VDD.n3705 VDD 0.0902606
R16909 VDD.n3963 VDD 0.0902606
R16910 VDD.n4221 VDD 0.0902606
R16911 VDD.n4479 VDD 0.0902606
R16912 VDD.n4737 VDD 0.0902606
R16913 VDD.n4998 VDD 0.0902606
R16914 VDD.n5260 VDD 0.0902606
R16915 VDD.n1111 VDD 0.0900726
R16916 VDD.n850 VDD.n848 0.0892839
R16917 VDD.n55 VDD.n53 0.0892839
R16918 VDD.n449 VDD.n447 0.0892839
R16919 VDD.n1251 VDD.n1249 0.088354
R16920 VDD.n1797 VDD.n1778 0.0864543
R16921 VDD.n1800 VDD.n1778 0.0864543
R16922 VDD.n2005 VDD.n1986 0.0864543
R16923 VDD.n2008 VDD.n1986 0.0864543
R16924 VDD.n2376 VDD.n2357 0.0864543
R16925 VDD.n2379 VDD.n2357 0.0864543
R16926 VDD.n2634 VDD.n2615 0.0864543
R16927 VDD.n2637 VDD.n2615 0.0864543
R16928 VDD.n2892 VDD.n2873 0.0864543
R16929 VDD.n2895 VDD.n2873 0.0864543
R16930 VDD.n3150 VDD.n3131 0.0864543
R16931 VDD.n3153 VDD.n3131 0.0864543
R16932 VDD.n3408 VDD.n3389 0.0864543
R16933 VDD.n3411 VDD.n3389 0.0864543
R16934 VDD.n5738 VDD.n5719 0.0864543
R16935 VDD.n5741 VDD.n5719 0.0864543
R16936 VDD.n5484 VDD.n5465 0.0864543
R16937 VDD.n5487 VDD.n5465 0.0864543
R16938 VDD.n3666 VDD.n3647 0.0864543
R16939 VDD.n3669 VDD.n3647 0.0864543
R16940 VDD.n3924 VDD.n3905 0.0864543
R16941 VDD.n3927 VDD.n3905 0.0864543
R16942 VDD.n4182 VDD.n4163 0.0864543
R16943 VDD.n4185 VDD.n4163 0.0864543
R16944 VDD.n4440 VDD.n4421 0.0864543
R16945 VDD.n4443 VDD.n4421 0.0864543
R16946 VDD.n4698 VDD.n4679 0.0864543
R16947 VDD.n4701 VDD.n4679 0.0864543
R16948 VDD.n4957 VDD.n4938 0.0864543
R16949 VDD.n4960 VDD.n4938 0.0864543
R16950 VDD.n5107 VDD.n5088 0.0864543
R16951 VDD.n5110 VDD.n5088 0.0864543
R16952 VDD.n5869 VDD.n5868 0.0862917
R16953 VDD.n1774 VDD.n1665 0.0855148
R16954 VDD.n2123 VDD.n2014 0.0855148
R16955 VDD.n2353 VDD.n2244 0.0855148
R16956 VDD.n2611 VDD.n2502 0.0855148
R16957 VDD.n2869 VDD.n2760 0.0855148
R16958 VDD.n3127 VDD.n3018 0.0855148
R16959 VDD.n3385 VDD.n3276 0.0855148
R16960 VDD.n5715 VDD.n5606 0.0855148
R16961 VDD.n5461 VDD.n5352 0.0855148
R16962 VDD.n3643 VDD.n3534 0.0855148
R16963 VDD.n3901 VDD.n3792 0.0855148
R16964 VDD.n4159 VDD.n4050 0.0855148
R16965 VDD.n4417 VDD.n4308 0.0855148
R16966 VDD.n4675 VDD.n4566 0.0855148
R16967 VDD.n4933 VDD.n4824 0.0855148
R16968 VDD.n5225 VDD.n5116 0.0855148
R16969 VDD.n26 VDD.n25 0.0849867
R16970 VDD.n343 VDD.n342 0.0849867
R16971 VDD.n1832 VDD.n1825 0.0832206
R16972 VDD.n2153 VDD.n2146 0.0832206
R16973 VDD.n2411 VDD.n2404 0.0832206
R16974 VDD.n2669 VDD.n2662 0.0832206
R16975 VDD.n2927 VDD.n2920 0.0832206
R16976 VDD.n3185 VDD.n3178 0.0832206
R16977 VDD.n3443 VDD.n3436 0.0832206
R16978 VDD.n5770 VDD.n5763 0.0832206
R16979 VDD.n5516 VDD.n5509 0.0832206
R16980 VDD.n3701 VDD.n3694 0.0832206
R16981 VDD.n3959 VDD.n3952 0.0832206
R16982 VDD.n4217 VDD.n4210 0.0832206
R16983 VDD.n4475 VDD.n4468 0.0832206
R16984 VDD.n4733 VDD.n4726 0.0832206
R16985 VDD.n4994 VDD.n4987 0.0832206
R16986 VDD.n5256 VDD.n5249 0.0832206
R16987 VDD.n316 VDD.n315 0.082109
R16988 VDD.n1727 VDD.n1723 0.07913
R16989 VDD.n2076 VDD.n2072 0.07913
R16990 VDD.n2306 VDD.n2302 0.07913
R16991 VDD.n2564 VDD.n2560 0.07913
R16992 VDD.n2822 VDD.n2818 0.07913
R16993 VDD.n3080 VDD.n3076 0.07913
R16994 VDD.n3338 VDD.n3334 0.07913
R16995 VDD.n5668 VDD.n5664 0.07913
R16996 VDD.n5414 VDD.n5410 0.07913
R16997 VDD.n3596 VDD.n3592 0.07913
R16998 VDD.n3854 VDD.n3850 0.07913
R16999 VDD.n4112 VDD.n4108 0.07913
R17000 VDD.n4370 VDD.n4366 0.07913
R17001 VDD.n4628 VDD.n4624 0.07913
R17002 VDD.n4886 VDD.n4882 0.07913
R17003 VDD.n5178 VDD.n5174 0.07913
R17004 VDD.n1835 VDD.n1828 0.078625
R17005 VDD.n2156 VDD.n2149 0.078625
R17006 VDD.n2414 VDD.n2407 0.078625
R17007 VDD.n2672 VDD.n2665 0.078625
R17008 VDD.n2930 VDD.n2923 0.078625
R17009 VDD.n3188 VDD.n3181 0.078625
R17010 VDD.n3446 VDD.n3439 0.078625
R17011 VDD.n5773 VDD.n5766 0.078625
R17012 VDD.n5519 VDD.n5512 0.078625
R17013 VDD.n3704 VDD.n3697 0.078625
R17014 VDD.n3962 VDD.n3955 0.078625
R17015 VDD.n4220 VDD.n4213 0.078625
R17016 VDD.n4478 VDD.n4471 0.078625
R17017 VDD.n4736 VDD.n4729 0.078625
R17018 VDD.n4997 VDD.n4990 0.078625
R17019 VDD.n5259 VDD.n5252 0.078625
R17020 VDD.n33 VDD.n30 0.0777407
R17021 VDD.n350 VDD.n347 0.0777407
R17022 VDD.n1748 VDD.n1747 0.0773443
R17023 VDD.n2097 VDD.n2096 0.0773443
R17024 VDD.n2327 VDD.n2326 0.0773443
R17025 VDD.n2585 VDD.n2584 0.0773443
R17026 VDD.n2843 VDD.n2842 0.0773443
R17027 VDD.n3101 VDD.n3100 0.0773443
R17028 VDD.n3359 VDD.n3358 0.0773443
R17029 VDD.n5689 VDD.n5688 0.0773443
R17030 VDD.n5435 VDD.n5434 0.0773443
R17031 VDD.n3617 VDD.n3616 0.0773443
R17032 VDD.n3875 VDD.n3874 0.0773443
R17033 VDD.n4133 VDD.n4132 0.0773443
R17034 VDD.n4391 VDD.n4390 0.0773443
R17035 VDD.n4649 VDD.n4648 0.0773443
R17036 VDD.n4907 VDD.n4906 0.0773443
R17037 VDD.n5199 VDD.n5198 0.0773443
R17038 VDD.n1690 VDD.n1688 0.0755586
R17039 VDD.n2039 VDD.n2037 0.0755586
R17040 VDD.n2269 VDD.n2267 0.0755586
R17041 VDD.n2527 VDD.n2525 0.0755586
R17042 VDD.n2785 VDD.n2783 0.0755586
R17043 VDD.n3043 VDD.n3041 0.0755586
R17044 VDD.n3301 VDD.n3299 0.0755586
R17045 VDD.n5631 VDD.n5629 0.0755586
R17046 VDD.n5377 VDD.n5375 0.0755586
R17047 VDD.n3559 VDD.n3557 0.0755586
R17048 VDD.n3817 VDD.n3815 0.0755586
R17049 VDD.n4075 VDD.n4073 0.0755586
R17050 VDD.n4333 VDD.n4331 0.0755586
R17051 VDD.n4591 VDD.n4589 0.0755586
R17052 VDD.n4849 VDD.n4847 0.0755586
R17053 VDD.n5141 VDD.n5139 0.0755586
R17054 VDD.n827 VDD.n824 0.0734782
R17055 VDD.n754 VDD.n751 0.0734782
R17056 VDD.n425 VDD.n422 0.0734782
R17057 VDD.n1595 VDD.n1592 0.0734782
R17058 VDD.n1842 VDD.n1841 0.0710611
R17059 VDD.n2163 VDD.n2162 0.0710611
R17060 VDD.n2421 VDD.n2420 0.0710611
R17061 VDD.n2679 VDD.n2678 0.0710611
R17062 VDD.n2937 VDD.n2936 0.0710611
R17063 VDD.n3195 VDD.n3194 0.0710611
R17064 VDD.n3453 VDD.n3452 0.0710611
R17065 VDD.n5780 VDD.n5779 0.0710611
R17066 VDD.n5526 VDD.n5525 0.0710611
R17067 VDD.n3711 VDD.n3710 0.0710611
R17068 VDD.n3969 VDD.n3968 0.0710611
R17069 VDD.n4227 VDD.n4226 0.0710611
R17070 VDD.n4485 VDD.n4484 0.0710611
R17071 VDD.n4743 VDD.n4742 0.0710611
R17072 VDD.n5004 VDD.n5003 0.0710611
R17073 VDD.n5266 VDD.n5265 0.0710611
R17074 VDD.n1919 VDD.n1816 0.0705353
R17075 VDD.n2240 VDD.n2137 0.0705353
R17076 VDD.n2498 VDD.n2395 0.0705353
R17077 VDD.n2756 VDD.n2653 0.0705353
R17078 VDD.n3014 VDD.n2911 0.0705353
R17079 VDD.n3272 VDD.n3169 0.0705353
R17080 VDD.n3530 VDD.n3427 0.0705353
R17081 VDD.n5857 VDD.n5754 0.0705353
R17082 VDD.n5603 VDD.n5500 0.0705353
R17083 VDD.n3788 VDD.n3685 0.0705353
R17084 VDD.n4046 VDD.n3943 0.0705353
R17085 VDD.n4304 VDD.n4201 0.0705353
R17086 VDD.n4562 VDD.n4459 0.0705353
R17087 VDD.n4820 VDD.n4717 0.0705353
R17088 VDD.n5081 VDD.n4978 0.0705353
R17089 VDD.n5343 VDD.n5240 0.0705353
R17090 VDD.n1846 VDD.n1845 0.0694784
R17091 VDD.n1849 VDD.n1846 0.0694784
R17092 VDD.n2167 VDD.n2166 0.0694784
R17093 VDD.n2170 VDD.n2167 0.0694784
R17094 VDD.n2425 VDD.n2424 0.0694784
R17095 VDD.n2428 VDD.n2425 0.0694784
R17096 VDD.n2683 VDD.n2682 0.0694784
R17097 VDD.n2686 VDD.n2683 0.0694784
R17098 VDD.n2941 VDD.n2940 0.0694784
R17099 VDD.n2944 VDD.n2941 0.0694784
R17100 VDD.n3199 VDD.n3198 0.0694784
R17101 VDD.n3202 VDD.n3199 0.0694784
R17102 VDD.n3457 VDD.n3456 0.0694784
R17103 VDD.n3460 VDD.n3457 0.0694784
R17104 VDD.n5784 VDD.n5783 0.0694784
R17105 VDD.n5787 VDD.n5784 0.0694784
R17106 VDD.n5530 VDD.n5529 0.0694784
R17107 VDD.n5533 VDD.n5530 0.0694784
R17108 VDD.n3715 VDD.n3714 0.0694784
R17109 VDD.n3718 VDD.n3715 0.0694784
R17110 VDD.n3973 VDD.n3972 0.0694784
R17111 VDD.n3976 VDD.n3973 0.0694784
R17112 VDD.n4231 VDD.n4230 0.0694784
R17113 VDD.n4234 VDD.n4231 0.0694784
R17114 VDD.n4489 VDD.n4488 0.0694784
R17115 VDD.n4492 VDD.n4489 0.0694784
R17116 VDD.n4747 VDD.n4746 0.0694784
R17117 VDD.n4750 VDD.n4747 0.0694784
R17118 VDD.n5008 VDD.n5007 0.0694784
R17119 VDD.n5011 VDD.n5008 0.0694784
R17120 VDD.n5270 VDD.n5269 0.0694784
R17121 VDD.n5273 VDD.n5270 0.0694784
R17122 VDD.n775 VDD.n774 0.0681471
R17123 VDD.n774 VDD.n771 0.0681471
R17124 VDD.n771 VDD.n768 0.0681471
R17125 VDD.n768 VDD.n767 0.0681471
R17126 VDD.n767 VDD.n764 0.0681471
R17127 VDD.n372 VDD.n371 0.0681471
R17128 VDD.n371 VDD.n368 0.0681471
R17129 VDD.n368 VDD.n365 0.0681471
R17130 VDD.n365 VDD.n364 0.0681471
R17131 VDD.n364 VDD.n361 0.0681471
R17132 VDD.n723 VDD.n720 0.0671334
R17133 VDD.n1564 VDD.n1561 0.0671334
R17134 VDD.n22 VDD.n21 0.065907
R17135 VDD.n17 VDD.n4 0.065907
R17136 VDD.n16 VDD.n15 0.065907
R17137 VDD.n14 VDD.n10 0.065907
R17138 VDD.n339 VDD.n338 0.065907
R17139 VDD.n334 VDD.n321 0.065907
R17140 VDD.n333 VDD.n332 0.065907
R17141 VDD.n331 VDD.n327 0.065907
R17142 VDD.n797 VDD.n796 0.0658409
R17143 VDD.n395 VDD.n394 0.0658409
R17144 VDD.n5746 VDD 0.0644514
R17145 VDD.n5492 VDD 0.0644514
R17146 VDD.n1791 VDD.n1783 0.0643889
R17147 VDD.n1791 VDD.n1780 0.0643889
R17148 VDD.n1796 VDD.n1780 0.0643889
R17149 VDD.n1999 VDD.n1991 0.0643889
R17150 VDD.n1999 VDD.n1988 0.0643889
R17151 VDD.n2004 VDD.n1988 0.0643889
R17152 VDD.n2370 VDD.n2362 0.0643889
R17153 VDD.n2370 VDD.n2359 0.0643889
R17154 VDD.n2375 VDD.n2359 0.0643889
R17155 VDD.n2628 VDD.n2620 0.0643889
R17156 VDD.n2628 VDD.n2617 0.0643889
R17157 VDD.n2633 VDD.n2617 0.0643889
R17158 VDD.n2886 VDD.n2878 0.0643889
R17159 VDD.n2886 VDD.n2875 0.0643889
R17160 VDD.n2891 VDD.n2875 0.0643889
R17161 VDD.n3144 VDD.n3136 0.0643889
R17162 VDD.n3144 VDD.n3133 0.0643889
R17163 VDD.n3149 VDD.n3133 0.0643889
R17164 VDD.n3402 VDD.n3394 0.0643889
R17165 VDD.n3402 VDD.n3391 0.0643889
R17166 VDD.n3407 VDD.n3391 0.0643889
R17167 VDD.n5732 VDD.n5724 0.0643889
R17168 VDD.n5732 VDD.n5721 0.0643889
R17169 VDD.n5737 VDD.n5721 0.0643889
R17170 VDD.n5478 VDD.n5470 0.0643889
R17171 VDD.n5478 VDD.n5467 0.0643889
R17172 VDD.n5483 VDD.n5467 0.0643889
R17173 VDD.n3660 VDD.n3652 0.0643889
R17174 VDD.n3660 VDD.n3649 0.0643889
R17175 VDD.n3665 VDD.n3649 0.0643889
R17176 VDD.n3918 VDD.n3910 0.0643889
R17177 VDD.n3918 VDD.n3907 0.0643889
R17178 VDD.n3923 VDD.n3907 0.0643889
R17179 VDD.n4176 VDD.n4168 0.0643889
R17180 VDD.n4176 VDD.n4165 0.0643889
R17181 VDD.n4181 VDD.n4165 0.0643889
R17182 VDD.n4434 VDD.n4426 0.0643889
R17183 VDD.n4434 VDD.n4423 0.0643889
R17184 VDD.n4439 VDD.n4423 0.0643889
R17185 VDD.n4692 VDD.n4684 0.0643889
R17186 VDD.n4692 VDD.n4681 0.0643889
R17187 VDD.n4697 VDD.n4681 0.0643889
R17188 VDD.n4951 VDD.n4943 0.0643889
R17189 VDD.n4951 VDD.n4940 0.0643889
R17190 VDD.n4956 VDD.n4940 0.0643889
R17191 VDD.n5101 VDD.n5093 0.0643889
R17192 VDD.n5101 VDD.n5090 0.0643889
R17193 VDD.n5106 VDD.n5090 0.0643889
R17194 VDD.n824 VDD.n822 0.0643889
R17195 VDD.n822 VDD.n820 0.0643889
R17196 VDD.n820 VDD.n818 0.0643889
R17197 VDD.n815 VDD.n814 0.0643889
R17198 VDD.n814 VDD.n810 0.0643889
R17199 VDD.n810 VDD.n808 0.0643889
R17200 VDD.n803 VDD.n802 0.0643889
R17201 VDD.n751 VDD.n749 0.0643889
R17202 VDD.n749 VDD.n747 0.0643889
R17203 VDD.n747 VDD.n745 0.0643889
R17204 VDD.n738 VDD.n734 0.0643889
R17205 VDD.n734 VDD.n732 0.0643889
R17206 VDD.n732 VDD.n730 0.0643889
R17207 VDD.n717 VDD.n715 0.0643889
R17208 VDD.n715 VDD.n713 0.0643889
R17209 VDD.n422 VDD.n420 0.0643889
R17210 VDD.n420 VDD.n418 0.0643889
R17211 VDD.n418 VDD.n416 0.0643889
R17212 VDD.n413 VDD.n412 0.0643889
R17213 VDD.n412 VDD.n408 0.0643889
R17214 VDD.n408 VDD.n406 0.0643889
R17215 VDD.n401 VDD.n400 0.0643889
R17216 VDD.n1592 VDD.n1590 0.0643889
R17217 VDD.n1590 VDD.n1588 0.0643889
R17218 VDD.n1588 VDD.n1586 0.0643889
R17219 VDD.n1579 VDD.n1575 0.0643889
R17220 VDD.n1575 VDD.n1573 0.0643889
R17221 VDD.n1573 VDD.n1571 0.0643889
R17222 VDD.n1558 VDD.n1556 0.0643889
R17223 VDD.n1556 VDD.n1554 0.0643889
R17224 VDD.n1526 VDD 0.0639804
R17225 VDD.n1806 VDD 0.0630006
R17226 VDD.n2126 VDD 0.0630006
R17227 VDD.n2385 VDD 0.0630006
R17228 VDD.n2643 VDD 0.0630006
R17229 VDD.n2901 VDD 0.0630006
R17230 VDD.n3159 VDD 0.0630006
R17231 VDD.n3417 VDD 0.0630006
R17232 VDD.n3675 VDD 0.0630006
R17233 VDD.n3933 VDD 0.0630006
R17234 VDD.n4191 VDD 0.0630006
R17235 VDD.n4449 VDD 0.0630006
R17236 VDD.n4707 VDD 0.0630006
R17237 VDD.n4966 VDD 0.0630006
R17238 VDD.n5228 VDD 0.0630006
R17239 VDD.n1623 VDD 0.0604792
R17240 VDD.n779 VDD.n778 0.0599867
R17241 VDD.n376 VDD.n375 0.0599867
R17242 VDD.n1772 VDD.n1667 0.0588333
R17243 VDD.n2121 VDD.n2016 0.0588333
R17244 VDD.n2351 VDD.n2246 0.0588333
R17245 VDD.n2609 VDD.n2504 0.0588333
R17246 VDD.n2867 VDD.n2762 0.0588333
R17247 VDD.n3125 VDD.n3020 0.0588333
R17248 VDD.n3383 VDD.n3278 0.0588333
R17249 VDD.n5713 VDD.n5608 0.0588333
R17250 VDD.n5459 VDD.n5354 0.0588333
R17251 VDD.n3641 VDD.n3536 0.0588333
R17252 VDD.n3899 VDD.n3794 0.0588333
R17253 VDD.n4157 VDD.n4052 0.0588333
R17254 VDD.n4415 VDD.n4310 0.0588333
R17255 VDD.n4673 VDD.n4568 0.0588333
R17256 VDD.n4931 VDD.n4826 0.0588333
R17257 VDD.n5223 VDD.n5118 0.0588333
R17258 VDD.n712 VDD.n711 0.0587674
R17259 VDD.n1553 VDD.n1552 0.0587674
R17260 VDD.n742 VDD.n741 0.0580441
R17261 VDD.n1583 VDD.n1582 0.0580441
R17262 VDD.n1165 VDD 0.058
R17263 VDD.n1159 VDD 0.058
R17264 VDD.n1147 VDD 0.058
R17265 VDD.n1231 VDD 0.058
R17266 VDD.n1225 VDD 0.058
R17267 VDD.n1213 VDD 0.058
R17268 VDD.n808 VDD.n806 0.0567153
R17269 VDD.n406 VDD.n404 0.0567153
R17270 VDD.n5870 VDD.n5869 0.0560833
R17271 VDD.n1153 VDD 0.0555
R17272 VDD.n1219 VDD 0.0555
R17273 VDD VDD.n1783 0.0525833
R17274 VDD VDD.n1991 0.0525833
R17275 VDD VDD.n2362 0.0525833
R17276 VDD VDD.n2620 0.0525833
R17277 VDD VDD.n2878 0.0525833
R17278 VDD VDD.n3136 0.0525833
R17279 VDD VDD.n3394 0.0525833
R17280 VDD VDD.n5724 0.0525833
R17281 VDD VDD.n5470 0.0525833
R17282 VDD VDD.n3652 0.0525833
R17283 VDD VDD.n3910 0.0525833
R17284 VDD VDD.n4168 0.0525833
R17285 VDD VDD.n4426 0.0525833
R17286 VDD VDD.n4684 0.0525833
R17287 VDD VDD.n4943 0.0525833
R17288 VDD VDD.n5093 0.0525833
R17289 VDD.n798 VDD.n797 0.0516364
R17290 VDD.n396 VDD.n395 0.0516364
R17291 VDD VDD.n5867 0.0470704
R17292 VDD.n1799 VDD 0.0470278
R17293 VDD.n2007 VDD 0.0470278
R17294 VDD.n2378 VDD 0.0470278
R17295 VDD.n2636 VDD 0.0470278
R17296 VDD.n2894 VDD 0.0470278
R17297 VDD.n3152 VDD 0.0470278
R17298 VDD.n3410 VDD 0.0470278
R17299 VDD.n5740 VDD 0.0470278
R17300 VDD.n5486 VDD 0.0470278
R17301 VDD.n3668 VDD 0.0470278
R17302 VDD.n3926 VDD 0.0470278
R17303 VDD.n4184 VDD 0.0470278
R17304 VDD.n4442 VDD 0.0470278
R17305 VDD.n4700 VDD 0.0470278
R17306 VDD.n4959 VDD 0.0470278
R17307 VDD.n5109 VDD 0.0470278
R17308 VDD.n5083 VDD.n5082 0.0460643
R17309 VDD.n5346 VDD.n5345 0.0438717
R17310 VDD.n5226 VDD.n5084 0.0438548
R17311 VDD.n25 VDD.n0 0.0418891
R17312 VDD.n342 VDD.n317 0.0418891
R17313 VDD.n1832 VDD.n1831 0.0409412
R17314 VDD.n2153 VDD.n2152 0.0409412
R17315 VDD.n2411 VDD.n2410 0.0409412
R17316 VDD.n2669 VDD.n2668 0.0409412
R17317 VDD.n2927 VDD.n2926 0.0409412
R17318 VDD.n3185 VDD.n3184 0.0409412
R17319 VDD.n3443 VDD.n3442 0.0409412
R17320 VDD.n5770 VDD.n5769 0.0409412
R17321 VDD.n5516 VDD.n5515 0.0409412
R17322 VDD.n3701 VDD.n3700 0.0409412
R17323 VDD.n3959 VDD.n3958 0.0409412
R17324 VDD.n4217 VDD.n4216 0.0409412
R17325 VDD.n4475 VDD.n4474 0.0409412
R17326 VDD.n4733 VDD.n4732 0.0409412
R17327 VDD.n4994 VDD.n4993 0.0409412
R17328 VDD.n5256 VDD.n5255 0.0409412
R17329 VDD.n30 VDD.n28 0.0409412
R17330 VDD.n347 VDD.n345 0.0409412
R17331 VDD.n5716 VDD.n5715 0.0399318
R17332 VDD.n5462 VDD.n5461 0.0399318
R17333 VDD.n1137 VDD.n1116 0.03976
R17334 VDD.n1203 VDD.n1182 0.03976
R17335 VDD.n1797 VDD.n1776 0.0395625
R17336 VDD.n2005 VDD.n1984 0.0395625
R17337 VDD.n2376 VDD.n2355 0.0395625
R17338 VDD.n2634 VDD.n2613 0.0395625
R17339 VDD.n2892 VDD.n2871 0.0395625
R17340 VDD.n3150 VDD.n3129 0.0395625
R17341 VDD.n3408 VDD.n3387 0.0395625
R17342 VDD.n5738 VDD.n5717 0.0395625
R17343 VDD.n5484 VDD.n5463 0.0395625
R17344 VDD.n3666 VDD.n3645 0.0395625
R17345 VDD.n3924 VDD.n3903 0.0395625
R17346 VDD.n4182 VDD.n4161 0.0395625
R17347 VDD.n4440 VDD.n4419 0.0395625
R17348 VDD.n4698 VDD.n4677 0.0395625
R17349 VDD.n4957 VDD.n4936 0.0395625
R17350 VDD.n5107 VDD.n5086 0.0395625
R17351 VDD.n5082 VDD.n4970 0.0394687
R17352 VDD.n1114 VDD 0.0390887
R17353 VDD.n1171 VDD.n1170 0.0376094
R17354 VDD.n1237 VDD.n1236 0.0376094
R17355 VDD.n1836 VDD.n1835 0.0372647
R17356 VDD.n2157 VDD.n2156 0.0372647
R17357 VDD.n2415 VDD.n2414 0.0372647
R17358 VDD.n2673 VDD.n2672 0.0372647
R17359 VDD.n2931 VDD.n2930 0.0372647
R17360 VDD.n3189 VDD.n3188 0.0372647
R17361 VDD.n3447 VDD.n3446 0.0372647
R17362 VDD.n5774 VDD.n5773 0.0372647
R17363 VDD.n5520 VDD.n5519 0.0372647
R17364 VDD.n3705 VDD.n3704 0.0372647
R17365 VDD.n3963 VDD.n3962 0.0372647
R17366 VDD.n4221 VDD.n4220 0.0372647
R17367 VDD.n4479 VDD.n4478 0.0372647
R17368 VDD.n4737 VDD.n4736 0.0372647
R17369 VDD.n4998 VDD.n4997 0.0372647
R17370 VDD.n5260 VDD.n5259 0.0372647
R17371 VDD.n28 VDD.n27 0.0371297
R17372 VDD.n345 VDD.n344 0.0371297
R17373 VDD.n1701 VDD.n1665 0.0364409
R17374 VDD.n2050 VDD.n2014 0.0364409
R17375 VDD.n2280 VDD.n2244 0.0364409
R17376 VDD.n2538 VDD.n2502 0.0364409
R17377 VDD.n2796 VDD.n2760 0.0364409
R17378 VDD.n3054 VDD.n3018 0.0364409
R17379 VDD.n3312 VDD.n3276 0.0364409
R17380 VDD.n5642 VDD.n5606 0.0364409
R17381 VDD.n5388 VDD.n5352 0.0364409
R17382 VDD.n3570 VDD.n3534 0.0364409
R17383 VDD.n3828 VDD.n3792 0.0364409
R17384 VDD.n4086 VDD.n4050 0.0364409
R17385 VDD.n4344 VDD.n4308 0.0364409
R17386 VDD.n4602 VDD.n4566 0.0364409
R17387 VDD.n4860 VDD.n4824 0.0364409
R17388 VDD.n5152 VDD.n5116 0.0364409
R17389 VDD.n1837 VDD.n1836 0.0361152
R17390 VDD.n2158 VDD.n2157 0.0361152
R17391 VDD.n2416 VDD.n2415 0.0361152
R17392 VDD.n2674 VDD.n2673 0.0361152
R17393 VDD.n2932 VDD.n2931 0.0361152
R17394 VDD.n3190 VDD.n3189 0.0361152
R17395 VDD.n3448 VDD.n3447 0.0361152
R17396 VDD.n5775 VDD.n5774 0.0361152
R17397 VDD.n5521 VDD.n5520 0.0361152
R17398 VDD.n3706 VDD.n3705 0.0361152
R17399 VDD.n3964 VDD.n3963 0.0361152
R17400 VDD.n4222 VDD.n4221 0.0361152
R17401 VDD.n4480 VDD.n4479 0.0361152
R17402 VDD.n4738 VDD.n4737 0.0361152
R17403 VDD.n4999 VDD.n4998 0.0361152
R17404 VDD.n5261 VDD.n5260 0.0361152
R17405 VDD.n1752 VDD.n1751 0.0357224
R17406 VDD.n2101 VDD.n2100 0.0357224
R17407 VDD.n2331 VDD.n2330 0.0357224
R17408 VDD.n2589 VDD.n2588 0.0357224
R17409 VDD.n2847 VDD.n2846 0.0357224
R17410 VDD.n3105 VDD.n3104 0.0357224
R17411 VDD.n3363 VDD.n3362 0.0357224
R17412 VDD.n5693 VDD.n5692 0.0357224
R17413 VDD.n5439 VDD.n5438 0.0357224
R17414 VDD.n3621 VDD.n3620 0.0357224
R17415 VDD.n3879 VDD.n3878 0.0357224
R17416 VDD.n4137 VDD.n4136 0.0357224
R17417 VDD.n4395 VDD.n4394 0.0357224
R17418 VDD.n4653 VDD.n4652 0.0357224
R17419 VDD.n4911 VDD.n4910 0.0357224
R17420 VDD.n5203 VDD.n5202 0.0357224
R17421 VDD.n1684 VDD.n1683 0.034445
R17422 VDD.n2033 VDD.n2032 0.034445
R17423 VDD.n2263 VDD.n2262 0.034445
R17424 VDD.n2521 VDD.n2520 0.034445
R17425 VDD.n2779 VDD.n2778 0.034445
R17426 VDD.n3037 VDD.n3036 0.034445
R17427 VDD.n3295 VDD.n3294 0.034445
R17428 VDD.n5625 VDD.n5624 0.034445
R17429 VDD.n5371 VDD.n5370 0.034445
R17430 VDD.n3553 VDD.n3552 0.034445
R17431 VDD.n3811 VDD.n3810 0.034445
R17432 VDD.n4069 VDD.n4068 0.034445
R17433 VDD.n4327 VDD.n4326 0.034445
R17434 VDD.n4585 VDD.n4584 0.034445
R17435 VDD.n4843 VDD.n4842 0.034445
R17436 VDD.n5135 VDD.n5134 0.034445
R17437 VDD.n3 VDD.n0 0.0339302
R17438 VDD.n320 VDD.n317 0.0339302
R17439 VDD.n1127 VDD.n1119 0.033737
R17440 VDD.n1131 VDD.n1119 0.033737
R17441 VDD.n1132 VDD.n1131 0.033737
R17442 VDD.n1133 VDD.n1132 0.033737
R17443 VDD.n1193 VDD.n1185 0.033737
R17444 VDD.n1197 VDD.n1185 0.033737
R17445 VDD.n1198 VDD.n1197 0.033737
R17446 VDD.n1199 VDD.n1198 0.033737
R17447 VDD.n796 VDD.n794 0.0334425
R17448 VDD.n794 VDD.n791 0.0334425
R17449 VDD.n394 VDD.n392 0.0334425
R17450 VDD.n392 VDD.n389 0.0334425
R17451 VDD.n1548 VDD.n1547 0.0333707
R17452 VDD.n1180 VDD.n1115 0.0325611
R17453 VDD VDD.n1796 0.0324444
R17454 VDD VDD.n2004 0.0324444
R17455 VDD VDD.n2375 0.0324444
R17456 VDD VDD.n2633 0.0324444
R17457 VDD VDD.n2891 0.0324444
R17458 VDD VDD.n3149 0.0324444
R17459 VDD VDD.n3407 0.0324444
R17460 VDD VDD.n5737 0.0324444
R17461 VDD VDD.n5483 0.0324444
R17462 VDD VDD.n3665 0.0324444
R17463 VDD VDD.n3923 0.0324444
R17464 VDD VDD.n4181 0.0324444
R17465 VDD VDD.n4439 0.0324444
R17466 VDD VDD.n4697 0.0324444
R17467 VDD VDD.n4956 0.0324444
R17468 VDD VDD.n5106 0.0324444
R17469 VDD.n815 VDD 0.0324444
R17470 VDD.n803 VDD 0.0324444
R17471 VDD.n742 VDD 0.0324444
R17472 VDD.n413 VDD 0.0324444
R17473 VDD.n401 VDD 0.0324444
R17474 VDD.n1583 VDD 0.0324444
R17475 VDD.n5867 VDD.n1921 0.0317545
R17476 VDD.n5865 VDD.n2242 0.0317545
R17477 VDD.n5864 VDD.n2500 0.0317545
R17478 VDD.n5863 VDD.n2758 0.0317545
R17479 VDD.n5862 VDD.n3016 0.0317545
R17480 VDD.n5861 VDD.n3274 0.0317545
R17481 VDD.n5860 VDD.n3532 0.0317545
R17482 VDD.n5351 VDD.n3790 0.0317545
R17483 VDD.n5350 VDD.n4048 0.0317545
R17484 VDD.n5349 VDD.n4306 0.0317545
R17485 VDD.n5348 VDD.n4564 0.0317545
R17486 VDD.n5347 VDD.n4822 0.0317545
R17487 VDD.n1640 VDD.n1639 0.0308571
R17488 VDD.n5344 VDD.n5232 0.0302768
R17489 VDD.n427 VDD.n379 0.0299677
R17490 VDD.n1115 VDD.n427 0.0299677
R17491 VDD.n830 VDD.n829 0.0299677
R17492 VDD.n1771 VDD.n1770 0.0294474
R17493 VDD.n2120 VDD.n2119 0.0294474
R17494 VDD.n2350 VDD.n2349 0.0294474
R17495 VDD.n2608 VDD.n2607 0.0294474
R17496 VDD.n2866 VDD.n2865 0.0294474
R17497 VDD.n3124 VDD.n3123 0.0294474
R17498 VDD.n3382 VDD.n3381 0.0294474
R17499 VDD.n5712 VDD.n5711 0.0294474
R17500 VDD.n5458 VDD.n5457 0.0294474
R17501 VDD.n3640 VDD.n3639 0.0294474
R17502 VDD.n3898 VDD.n3897 0.0294474
R17503 VDD.n4156 VDD.n4155 0.0294474
R17504 VDD.n4414 VDD.n4413 0.0294474
R17505 VDD.n4672 VDD.n4671 0.0294474
R17506 VDD.n4930 VDD.n4929 0.0294474
R17507 VDD.n5222 VDD.n5221 0.0294474
R17508 VDD.n1598 VDD.n1597 0.0292661
R17509 VDD.n1113 VDD.n1112 0.0292661
R17510 VDD.n379 VDD.n352 0.0290323
R17511 VDD.n1754 VDD.n1753 0.0287895
R17512 VDD.n2103 VDD.n2102 0.0287895
R17513 VDD.n2333 VDD.n2332 0.0287895
R17514 VDD.n2591 VDD.n2590 0.0287895
R17515 VDD.n2849 VDD.n2848 0.0287895
R17516 VDD.n3107 VDD.n3106 0.0287895
R17517 VDD.n3365 VDD.n3364 0.0287895
R17518 VDD.n5695 VDD.n5694 0.0287895
R17519 VDD.n5441 VDD.n5440 0.0287895
R17520 VDD.n3623 VDD.n3622 0.0287895
R17521 VDD.n3881 VDD.n3880 0.0287895
R17522 VDD.n4139 VDD.n4138 0.0287895
R17523 VDD.n4397 VDD.n4396 0.0287895
R17524 VDD.n4655 VDD.n4654 0.0287895
R17525 VDD.n4913 VDD.n4912 0.0287895
R17526 VDD.n5205 VDD.n5204 0.0287895
R17527 VDD.n1750 VDD.n1720 0.0282778
R17528 VDD.n2099 VDD.n2069 0.0282778
R17529 VDD.n2329 VDD.n2299 0.0282778
R17530 VDD.n2587 VDD.n2557 0.0282778
R17531 VDD.n2845 VDD.n2815 0.0282778
R17532 VDD.n3103 VDD.n3073 0.0282778
R17533 VDD.n3361 VDD.n3331 0.0282778
R17534 VDD.n5691 VDD.n5661 0.0282778
R17535 VDD.n5437 VDD.n5407 0.0282778
R17536 VDD.n3619 VDD.n3589 0.0282778
R17537 VDD.n3877 VDD.n3847 0.0282778
R17538 VDD.n4135 VDD.n4105 0.0282778
R17539 VDD.n4393 VDD.n4363 0.0282778
R17540 VDD.n4651 VDD.n4621 0.0282778
R17541 VDD.n4909 VDD.n4879 0.0282778
R17542 VDD.n5201 VDD.n5171 0.0282778
R17543 VDD.t753 VDD.n1763 0.0282694
R17544 VDD.n1763 VDD.n1762 0.0282694
R17545 VDD.t753 VDD.n1677 0.0282694
R17546 VDD.n1706 VDD.n1677 0.0282694
R17547 VDD.t129 VDD.n2112 0.0282694
R17548 VDD.n2112 VDD.n2111 0.0282694
R17549 VDD.t129 VDD.n2026 0.0282694
R17550 VDD.n2055 VDD.n2026 0.0282694
R17551 VDD.t70 VDD.n2342 0.0282694
R17552 VDD.n2342 VDD.n2341 0.0282694
R17553 VDD.t70 VDD.n2256 0.0282694
R17554 VDD.n2285 VDD.n2256 0.0282694
R17555 VDD.t680 VDD.n2600 0.0282694
R17556 VDD.n2600 VDD.n2599 0.0282694
R17557 VDD.t680 VDD.n2514 0.0282694
R17558 VDD.n2543 VDD.n2514 0.0282694
R17559 VDD.t733 VDD.n2858 0.0282694
R17560 VDD.n2858 VDD.n2857 0.0282694
R17561 VDD.t733 VDD.n2772 0.0282694
R17562 VDD.n2801 VDD.n2772 0.0282694
R17563 VDD.t125 VDD.n3116 0.0282694
R17564 VDD.n3116 VDD.n3115 0.0282694
R17565 VDD.t125 VDD.n3030 0.0282694
R17566 VDD.n3059 VDD.n3030 0.0282694
R17567 VDD.t504 VDD.n3374 0.0282694
R17568 VDD.n3374 VDD.n3373 0.0282694
R17569 VDD.t504 VDD.n3288 0.0282694
R17570 VDD.n3317 VDD.n3288 0.0282694
R17571 VDD.t4 VDD.n5704 0.0282694
R17572 VDD.n5704 VDD.n5703 0.0282694
R17573 VDD.t4 VDD.n5618 0.0282694
R17574 VDD.n5647 VDD.n5618 0.0282694
R17575 VDD.t665 VDD.n5450 0.0282694
R17576 VDD.n5450 VDD.n5449 0.0282694
R17577 VDD.t665 VDD.n5364 0.0282694
R17578 VDD.n5393 VDD.n5364 0.0282694
R17579 VDD.t1141 VDD.n3632 0.0282694
R17580 VDD.n3632 VDD.n3631 0.0282694
R17581 VDD.t1141 VDD.n3546 0.0282694
R17582 VDD.n3575 VDD.n3546 0.0282694
R17583 VDD.t1061 VDD.n3890 0.0282694
R17584 VDD.n3890 VDD.n3889 0.0282694
R17585 VDD.t1061 VDD.n3804 0.0282694
R17586 VDD.n3833 VDD.n3804 0.0282694
R17587 VDD.t414 VDD.n4148 0.0282694
R17588 VDD.n4148 VDD.n4147 0.0282694
R17589 VDD.t414 VDD.n4062 0.0282694
R17590 VDD.n4091 VDD.n4062 0.0282694
R17591 VDD.t165 VDD.n4406 0.0282694
R17592 VDD.n4406 VDD.n4405 0.0282694
R17593 VDD.t165 VDD.n4320 0.0282694
R17594 VDD.n4349 VDD.n4320 0.0282694
R17595 VDD.t793 VDD.n4664 0.0282694
R17596 VDD.n4664 VDD.n4663 0.0282694
R17597 VDD.t793 VDD.n4578 0.0282694
R17598 VDD.n4607 VDD.n4578 0.0282694
R17599 VDD.t1065 VDD.n4922 0.0282694
R17600 VDD.n4922 VDD.n4921 0.0282694
R17601 VDD.t1065 VDD.n4836 0.0282694
R17602 VDD.n4865 VDD.n4836 0.0282694
R17603 VDD.t107 VDD.n5214 0.0282694
R17604 VDD.n5214 VDD.n5213 0.0282694
R17605 VDD.t107 VDD.n5128 0.0282694
R17606 VDD.n5157 VDD.n5128 0.0282694
R17607 VDD.n991 VDD 0.0279106
R17608 VDD.n196 VDD 0.0279106
R17609 VDD.n586 VDD 0.0279106
R17610 VDD.n5346 VDD.n5083 0.0269368
R17611 VDD.n1897 VDD.n1895 0.0265784
R17612 VDD.n1905 VDD.n1895 0.0265784
R17613 VDD.n1911 VDD.n1896 0.0265784
R17614 VDD.n1901 VDD.n1896 0.0265784
R17615 VDD.n1903 VDD.n1902 0.0265784
R17616 VDD.n1902 VDD.n1901 0.0265784
R17617 VDD.n1907 VDD.n1906 0.0265784
R17618 VDD.n1906 VDD.n1905 0.0265784
R17619 VDD.n1878 VDD.n1877 0.0265784
R17620 VDD.t417 VDD.n1878 0.0265784
R17621 VDD.n1880 VDD.n1822 0.0265784
R17622 VDD.n1860 VDD.n1859 0.0265784
R17623 VDD.n1859 VDD.n1858 0.0265784
R17624 VDD.n1862 VDD.n1853 0.0265784
R17625 VDD.n1863 VDD.n1862 0.0265784
R17626 VDD.n1865 VDD.n1864 0.0265784
R17627 VDD.n1864 VDD.n1863 0.0265784
R17628 VDD.n1858 VDD.n1855 0.0265784
R17629 VDD.n1855 VDD.n1854 0.0265784
R17630 VDD.n2181 VDD.n2180 0.0265784
R17631 VDD.n2180 VDD.n2179 0.0265784
R17632 VDD.n2183 VDD.n2174 0.0265784
R17633 VDD.n2184 VDD.n2183 0.0265784
R17634 VDD.n2186 VDD.n2185 0.0265784
R17635 VDD.n2185 VDD.n2184 0.0265784
R17636 VDD.n2179 VDD.n2176 0.0265784
R17637 VDD.n2176 VDD.n2175 0.0265784
R17638 VDD.n2199 VDD.n2198 0.0265784
R17639 VDD.t1085 VDD.n2199 0.0265784
R17640 VDD.n2201 VDD.n2143 0.0265784
R17641 VDD.n2218 VDD.n2216 0.0265784
R17642 VDD.n2226 VDD.n2216 0.0265784
R17643 VDD.n2232 VDD.n2217 0.0265784
R17644 VDD.n2222 VDD.n2217 0.0265784
R17645 VDD.n2224 VDD.n2223 0.0265784
R17646 VDD.n2223 VDD.n2222 0.0265784
R17647 VDD.n2228 VDD.n2227 0.0265784
R17648 VDD.n2227 VDD.n2226 0.0265784
R17649 VDD.n2439 VDD.n2438 0.0265784
R17650 VDD.n2438 VDD.n2437 0.0265784
R17651 VDD.n2441 VDD.n2432 0.0265784
R17652 VDD.n2442 VDD.n2441 0.0265784
R17653 VDD.n2444 VDD.n2443 0.0265784
R17654 VDD.n2443 VDD.n2442 0.0265784
R17655 VDD.n2437 VDD.n2434 0.0265784
R17656 VDD.n2434 VDD.n2433 0.0265784
R17657 VDD.n2457 VDD.n2456 0.0265784
R17658 VDD.t567 VDD.n2457 0.0265784
R17659 VDD.n2459 VDD.n2401 0.0265784
R17660 VDD.n2476 VDD.n2474 0.0265784
R17661 VDD.n2484 VDD.n2474 0.0265784
R17662 VDD.n2490 VDD.n2475 0.0265784
R17663 VDD.n2480 VDD.n2475 0.0265784
R17664 VDD.n2482 VDD.n2481 0.0265784
R17665 VDD.n2481 VDD.n2480 0.0265784
R17666 VDD.n2486 VDD.n2485 0.0265784
R17667 VDD.n2485 VDD.n2484 0.0265784
R17668 VDD.n2697 VDD.n2696 0.0265784
R17669 VDD.n2696 VDD.n2695 0.0265784
R17670 VDD.n2699 VDD.n2690 0.0265784
R17671 VDD.n2700 VDD.n2699 0.0265784
R17672 VDD.n2702 VDD.n2701 0.0265784
R17673 VDD.n2701 VDD.n2700 0.0265784
R17674 VDD.n2695 VDD.n2692 0.0265784
R17675 VDD.n2692 VDD.n2691 0.0265784
R17676 VDD.n2715 VDD.n2714 0.0265784
R17677 VDD.t387 VDD.n2715 0.0265784
R17678 VDD.n2717 VDD.n2659 0.0265784
R17679 VDD.n2734 VDD.n2732 0.0265784
R17680 VDD.n2742 VDD.n2732 0.0265784
R17681 VDD.n2748 VDD.n2733 0.0265784
R17682 VDD.n2738 VDD.n2733 0.0265784
R17683 VDD.n2740 VDD.n2739 0.0265784
R17684 VDD.n2739 VDD.n2738 0.0265784
R17685 VDD.n2744 VDD.n2743 0.0265784
R17686 VDD.n2743 VDD.n2742 0.0265784
R17687 VDD.n2955 VDD.n2954 0.0265784
R17688 VDD.n2954 VDD.n2953 0.0265784
R17689 VDD.n2957 VDD.n2948 0.0265784
R17690 VDD.n2958 VDD.n2957 0.0265784
R17691 VDD.n2960 VDD.n2959 0.0265784
R17692 VDD.n2959 VDD.n2958 0.0265784
R17693 VDD.n2953 VDD.n2950 0.0265784
R17694 VDD.n2950 VDD.n2949 0.0265784
R17695 VDD.n2973 VDD.n2972 0.0265784
R17696 VDD.t560 VDD.n2973 0.0265784
R17697 VDD.n2975 VDD.n2917 0.0265784
R17698 VDD.n2992 VDD.n2990 0.0265784
R17699 VDD.n3000 VDD.n2990 0.0265784
R17700 VDD.n3006 VDD.n2991 0.0265784
R17701 VDD.n2996 VDD.n2991 0.0265784
R17702 VDD.n2998 VDD.n2997 0.0265784
R17703 VDD.n2997 VDD.n2996 0.0265784
R17704 VDD.n3002 VDD.n3001 0.0265784
R17705 VDD.n3001 VDD.n3000 0.0265784
R17706 VDD.n3213 VDD.n3212 0.0265784
R17707 VDD.n3212 VDD.n3211 0.0265784
R17708 VDD.n3215 VDD.n3206 0.0265784
R17709 VDD.n3216 VDD.n3215 0.0265784
R17710 VDD.n3218 VDD.n3217 0.0265784
R17711 VDD.n3217 VDD.n3216 0.0265784
R17712 VDD.n3211 VDD.n3208 0.0265784
R17713 VDD.n3208 VDD.n3207 0.0265784
R17714 VDD.n3231 VDD.n3230 0.0265784
R17715 VDD.t573 VDD.n3231 0.0265784
R17716 VDD.n3233 VDD.n3175 0.0265784
R17717 VDD.n3250 VDD.n3248 0.0265784
R17718 VDD.n3258 VDD.n3248 0.0265784
R17719 VDD.n3264 VDD.n3249 0.0265784
R17720 VDD.n3254 VDD.n3249 0.0265784
R17721 VDD.n3256 VDD.n3255 0.0265784
R17722 VDD.n3255 VDD.n3254 0.0265784
R17723 VDD.n3260 VDD.n3259 0.0265784
R17724 VDD.n3259 VDD.n3258 0.0265784
R17725 VDD.n3471 VDD.n3470 0.0265784
R17726 VDD.n3470 VDD.n3469 0.0265784
R17727 VDD.n3473 VDD.n3464 0.0265784
R17728 VDD.n3474 VDD.n3473 0.0265784
R17729 VDD.n3476 VDD.n3475 0.0265784
R17730 VDD.n3475 VDD.n3474 0.0265784
R17731 VDD.n3469 VDD.n3466 0.0265784
R17732 VDD.n3466 VDD.n3465 0.0265784
R17733 VDD.n3489 VDD.n3488 0.0265784
R17734 VDD.t143 VDD.n3489 0.0265784
R17735 VDD.n3491 VDD.n3433 0.0265784
R17736 VDD.n3508 VDD.n3506 0.0265784
R17737 VDD.n3516 VDD.n3506 0.0265784
R17738 VDD.n3522 VDD.n3507 0.0265784
R17739 VDD.n3512 VDD.n3507 0.0265784
R17740 VDD.n3514 VDD.n3513 0.0265784
R17741 VDD.n3513 VDD.n3512 0.0265784
R17742 VDD.n3518 VDD.n3517 0.0265784
R17743 VDD.n3517 VDD.n3516 0.0265784
R17744 VDD.n5798 VDD.n5797 0.0265784
R17745 VDD.n5797 VDD.n5796 0.0265784
R17746 VDD.n5800 VDD.n5791 0.0265784
R17747 VDD.n5801 VDD.n5800 0.0265784
R17748 VDD.n5803 VDD.n5802 0.0265784
R17749 VDD.n5802 VDD.n5801 0.0265784
R17750 VDD.n5796 VDD.n5793 0.0265784
R17751 VDD.n5793 VDD.n5792 0.0265784
R17752 VDD.n5816 VDD.n5815 0.0265784
R17753 VDD.t419 VDD.n5816 0.0265784
R17754 VDD.n5818 VDD.n5760 0.0265784
R17755 VDD.n5835 VDD.n5833 0.0265784
R17756 VDD.n5843 VDD.n5833 0.0265784
R17757 VDD.n5849 VDD.n5834 0.0265784
R17758 VDD.n5839 VDD.n5834 0.0265784
R17759 VDD.n5841 VDD.n5840 0.0265784
R17760 VDD.n5840 VDD.n5839 0.0265784
R17761 VDD.n5845 VDD.n5844 0.0265784
R17762 VDD.n5844 VDD.n5843 0.0265784
R17763 VDD.n5544 VDD.n5543 0.0265784
R17764 VDD.n5543 VDD.n5542 0.0265784
R17765 VDD.n5546 VDD.n5537 0.0265784
R17766 VDD.n5547 VDD.n5546 0.0265784
R17767 VDD.n5549 VDD.n5548 0.0265784
R17768 VDD.n5548 VDD.n5547 0.0265784
R17769 VDD.n5542 VDD.n5539 0.0265784
R17770 VDD.n5539 VDD.n5538 0.0265784
R17771 VDD.n5562 VDD.n5561 0.0265784
R17772 VDD.t667 VDD.n5562 0.0265784
R17773 VDD.n5564 VDD.n5506 0.0265784
R17774 VDD.n5581 VDD.n5579 0.0265784
R17775 VDD.n5589 VDD.n5579 0.0265784
R17776 VDD.n5595 VDD.n5580 0.0265784
R17777 VDD.n5585 VDD.n5580 0.0265784
R17778 VDD.n5587 VDD.n5586 0.0265784
R17779 VDD.n5586 VDD.n5585 0.0265784
R17780 VDD.n5591 VDD.n5590 0.0265784
R17781 VDD.n5590 VDD.n5589 0.0265784
R17782 VDD.n3729 VDD.n3728 0.0265784
R17783 VDD.n3728 VDD.n3727 0.0265784
R17784 VDD.n3731 VDD.n3722 0.0265784
R17785 VDD.n3732 VDD.n3731 0.0265784
R17786 VDD.n3734 VDD.n3733 0.0265784
R17787 VDD.n3733 VDD.n3732 0.0265784
R17788 VDD.n3727 VDD.n3724 0.0265784
R17789 VDD.n3724 VDD.n3723 0.0265784
R17790 VDD.n3747 VDD.n3746 0.0265784
R17791 VDD.t142 VDD.n3747 0.0265784
R17792 VDD.n3749 VDD.n3691 0.0265784
R17793 VDD.n3766 VDD.n3764 0.0265784
R17794 VDD.n3774 VDD.n3764 0.0265784
R17795 VDD.n3780 VDD.n3765 0.0265784
R17796 VDD.n3770 VDD.n3765 0.0265784
R17797 VDD.n3772 VDD.n3771 0.0265784
R17798 VDD.n3771 VDD.n3770 0.0265784
R17799 VDD.n3776 VDD.n3775 0.0265784
R17800 VDD.n3775 VDD.n3774 0.0265784
R17801 VDD.n3987 VDD.n3986 0.0265784
R17802 VDD.n3986 VDD.n3985 0.0265784
R17803 VDD.n3989 VDD.n3980 0.0265784
R17804 VDD.n3990 VDD.n3989 0.0265784
R17805 VDD.n3992 VDD.n3991 0.0265784
R17806 VDD.n3991 VDD.n3990 0.0265784
R17807 VDD.n3985 VDD.n3982 0.0265784
R17808 VDD.n3982 VDD.n3981 0.0265784
R17809 VDD.n4005 VDD.n4004 0.0265784
R17810 VDD.t782 VDD.n4005 0.0265784
R17811 VDD.n4007 VDD.n3949 0.0265784
R17812 VDD.n4024 VDD.n4022 0.0265784
R17813 VDD.n4032 VDD.n4022 0.0265784
R17814 VDD.n4038 VDD.n4023 0.0265784
R17815 VDD.n4028 VDD.n4023 0.0265784
R17816 VDD.n4030 VDD.n4029 0.0265784
R17817 VDD.n4029 VDD.n4028 0.0265784
R17818 VDD.n4034 VDD.n4033 0.0265784
R17819 VDD.n4033 VDD.n4032 0.0265784
R17820 VDD.n4245 VDD.n4244 0.0265784
R17821 VDD.n4244 VDD.n4243 0.0265784
R17822 VDD.n4247 VDD.n4238 0.0265784
R17823 VDD.n4248 VDD.n4247 0.0265784
R17824 VDD.n4250 VDD.n4249 0.0265784
R17825 VDD.n4249 VDD.n4248 0.0265784
R17826 VDD.n4243 VDD.n4240 0.0265784
R17827 VDD.n4240 VDD.n4239 0.0265784
R17828 VDD.n4263 VDD.n4262 0.0265784
R17829 VDD.t1087 VDD.n4263 0.0265784
R17830 VDD.n4265 VDD.n4207 0.0265784
R17831 VDD.n4282 VDD.n4280 0.0265784
R17832 VDD.n4290 VDD.n4280 0.0265784
R17833 VDD.n4296 VDD.n4281 0.0265784
R17834 VDD.n4286 VDD.n4281 0.0265784
R17835 VDD.n4288 VDD.n4287 0.0265784
R17836 VDD.n4287 VDD.n4286 0.0265784
R17837 VDD.n4292 VDD.n4291 0.0265784
R17838 VDD.n4291 VDD.n4290 0.0265784
R17839 VDD.n4503 VDD.n4502 0.0265784
R17840 VDD.n4502 VDD.n4501 0.0265784
R17841 VDD.n4505 VDD.n4496 0.0265784
R17842 VDD.n4506 VDD.n4505 0.0265784
R17843 VDD.n4508 VDD.n4507 0.0265784
R17844 VDD.n4507 VDD.n4506 0.0265784
R17845 VDD.n4501 VDD.n4498 0.0265784
R17846 VDD.n4498 VDD.n4497 0.0265784
R17847 VDD.n4521 VDD.n4520 0.0265784
R17848 VDD.t558 VDD.n4521 0.0265784
R17849 VDD.n4523 VDD.n4465 0.0265784
R17850 VDD.n4540 VDD.n4538 0.0265784
R17851 VDD.n4548 VDD.n4538 0.0265784
R17852 VDD.n4554 VDD.n4539 0.0265784
R17853 VDD.n4544 VDD.n4539 0.0265784
R17854 VDD.n4546 VDD.n4545 0.0265784
R17855 VDD.n4545 VDD.n4544 0.0265784
R17856 VDD.n4550 VDD.n4549 0.0265784
R17857 VDD.n4549 VDD.n4548 0.0265784
R17858 VDD.n4761 VDD.n4760 0.0265784
R17859 VDD.n4760 VDD.n4759 0.0265784
R17860 VDD.n4763 VDD.n4754 0.0265784
R17861 VDD.n4764 VDD.n4763 0.0265784
R17862 VDD.n4766 VDD.n4765 0.0265784
R17863 VDD.n4765 VDD.n4764 0.0265784
R17864 VDD.n4759 VDD.n4756 0.0265784
R17865 VDD.n4756 VDD.n4755 0.0265784
R17866 VDD.n4779 VDD.n4778 0.0265784
R17867 VDD.t572 VDD.n4779 0.0265784
R17868 VDD.n4781 VDD.n4723 0.0265784
R17869 VDD.n4798 VDD.n4796 0.0265784
R17870 VDD.n4806 VDD.n4796 0.0265784
R17871 VDD.n4812 VDD.n4797 0.0265784
R17872 VDD.n4802 VDD.n4797 0.0265784
R17873 VDD.n4804 VDD.n4803 0.0265784
R17874 VDD.n4803 VDD.n4802 0.0265784
R17875 VDD.n4808 VDD.n4807 0.0265784
R17876 VDD.n4807 VDD.n4806 0.0265784
R17877 VDD.n5059 VDD.n5057 0.0265784
R17878 VDD.n5067 VDD.n5057 0.0265784
R17879 VDD.n5073 VDD.n5058 0.0265784
R17880 VDD.n5063 VDD.n5058 0.0265784
R17881 VDD.n5065 VDD.n5064 0.0265784
R17882 VDD.n5064 VDD.n5063 0.0265784
R17883 VDD.n5069 VDD.n5068 0.0265784
R17884 VDD.n5068 VDD.n5067 0.0265784
R17885 VDD.n5040 VDD.n5039 0.0265784
R17886 VDD.t690 VDD.n5040 0.0265784
R17887 VDD.n5042 VDD.n4984 0.0265784
R17888 VDD.n5022 VDD.n5021 0.0265784
R17889 VDD.n5021 VDD.n5020 0.0265784
R17890 VDD.n5024 VDD.n5015 0.0265784
R17891 VDD.n5025 VDD.n5024 0.0265784
R17892 VDD.n5027 VDD.n5026 0.0265784
R17893 VDD.n5026 VDD.n5025 0.0265784
R17894 VDD.n5020 VDD.n5017 0.0265784
R17895 VDD.n5017 VDD.n5016 0.0265784
R17896 VDD.n5321 VDD.n5319 0.0265784
R17897 VDD.n5329 VDD.n5319 0.0265784
R17898 VDD.n5335 VDD.n5320 0.0265784
R17899 VDD.n5325 VDD.n5320 0.0265784
R17900 VDD.n5327 VDD.n5326 0.0265784
R17901 VDD.n5326 VDD.n5325 0.0265784
R17902 VDD.n5331 VDD.n5330 0.0265784
R17903 VDD.n5330 VDD.n5329 0.0265784
R17904 VDD.n5302 VDD.n5301 0.0265784
R17905 VDD.t418 VDD.n5302 0.0265784
R17906 VDD.n5304 VDD.n5246 0.0265784
R17907 VDD.n5284 VDD.n5283 0.0265784
R17908 VDD.n5283 VDD.n5282 0.0265784
R17909 VDD.n5286 VDD.n5277 0.0265784
R17910 VDD.n5287 VDD.n5286 0.0265784
R17911 VDD.n5289 VDD.n5288 0.0265784
R17912 VDD.n5288 VDD.n5287 0.0265784
R17913 VDD.n5282 VDD.n5279 0.0265784
R17914 VDD.n5279 VDD.n5278 0.0265784
R17915 VDD.n5859 VDD.n5858 0.0261294
R17916 VDD.n5605 VDD.n5604 0.0261294
R17917 VDD.n1840 VDD.n1825 0.0261194
R17918 VDD.n2161 VDD.n2146 0.0261194
R17919 VDD.n2419 VDD.n2404 0.0261194
R17920 VDD.n2677 VDD.n2662 0.0261194
R17921 VDD.n2935 VDD.n2920 0.0261194
R17922 VDD.n3193 VDD.n3178 0.0261194
R17923 VDD.n3451 VDD.n3436 0.0261194
R17924 VDD.n5778 VDD.n5763 0.0261194
R17925 VDD.n5524 VDD.n5509 0.0261194
R17926 VDD.n3709 VDD.n3694 0.0261194
R17927 VDD.n3967 VDD.n3952 0.0261194
R17928 VDD.n4225 VDD.n4210 0.0261194
R17929 VDD.n4483 VDD.n4468 0.0261194
R17930 VDD.n4741 VDD.n4726 0.0261194
R17931 VDD.n5002 VDD.n4987 0.0261194
R17932 VDD.n5264 VDD.n5249 0.0261194
R17933 VDD.n1304 VDD 0.0260435
R17934 VDD.n1945 VDD.n1922 0.0258165
R17935 VDD.n1696 VDD.n1683 0.0257918
R17936 VDD.n2045 VDD.n2032 0.0257918
R17937 VDD.n2275 VDD.n2262 0.0257918
R17938 VDD.n2533 VDD.n2520 0.0257918
R17939 VDD.n2791 VDD.n2778 0.0257918
R17940 VDD.n3049 VDD.n3036 0.0257918
R17941 VDD.n3307 VDD.n3294 0.0257918
R17942 VDD.n5637 VDD.n5624 0.0257918
R17943 VDD.n5383 VDD.n5370 0.0257918
R17944 VDD.n3565 VDD.n3552 0.0257918
R17945 VDD.n3823 VDD.n3810 0.0257918
R17946 VDD.n4081 VDD.n4068 0.0257918
R17947 VDD.n4339 VDD.n4326 0.0257918
R17948 VDD.n4597 VDD.n4584 0.0257918
R17949 VDD.n4855 VDD.n4842 0.0257918
R17950 VDD.n5147 VDD.n5134 0.0257918
R17951 VDD.n1880 VDD.n1879 0.02576
R17952 VDD.n2201 VDD.n2200 0.02576
R17953 VDD.n2459 VDD.n2458 0.02576
R17954 VDD.n2717 VDD.n2716 0.02576
R17955 VDD.n2975 VDD.n2974 0.02576
R17956 VDD.n3233 VDD.n3232 0.02576
R17957 VDD.n3491 VDD.n3490 0.02576
R17958 VDD.n5818 VDD.n5817 0.02576
R17959 VDD.n5564 VDD.n5563 0.02576
R17960 VDD.n3749 VDD.n3748 0.02576
R17961 VDD.n4007 VDD.n4006 0.02576
R17962 VDD.n4265 VDD.n4264 0.02576
R17963 VDD.n4523 VDD.n4522 0.02576
R17964 VDD.n4781 VDD.n4780 0.02576
R17965 VDD.n5042 VDD.n5041 0.02576
R17966 VDD.n5304 VDD.n5303 0.02576
R17967 VDD.n1315 VDD.n1314 0.0254026
R17968 VDD.n1310 VDD.n1308 0.0249681
R17969 VDD.n1311 VDD.n1310 0.0249681
R17970 VDD.n1453 VDD.n1449 0.0249681
R17971 VDD.n1449 VDD.n1447 0.0249681
R17972 VDD.n1447 VDD.n1443 0.0249681
R17973 VDD.n1443 VDD.n1441 0.0249681
R17974 VDD.n1441 VDD.n1437 0.0249681
R17975 VDD.n1437 VDD.n1433 0.0249681
R17976 VDD.n1331 VDD.n1327 0.0249681
R17977 VDD.n1333 VDD.n1331 0.0249681
R17978 VDD.n1337 VDD.n1333 0.0249681
R17979 VDD.n1339 VDD.n1337 0.0249681
R17980 VDD.n1340 VDD.n1339 0.0249681
R17981 VDD.n1422 VDD.n1418 0.0249681
R17982 VDD.n1418 VDD.n1416 0.0249681
R17983 VDD.n1416 VDD.n1412 0.0249681
R17984 VDD.n1412 VDD.n1410 0.0249681
R17985 VDD.n1393 VDD.n1389 0.0249681
R17986 VDD.n1389 VDD.n1387 0.0249681
R17987 VDD.n1387 VDD.n1383 0.0249681
R17988 VDD.n1383 VDD.n1381 0.0249681
R17989 VDD.n1351 VDD.n1349 0.0249681
R17990 VDD.n1354 VDD.n1351 0.0249681
R17991 VDD.n1356 VDD.n1354 0.0249681
R17992 VDD.n1358 VDD.n1356 0.0249681
R17993 VDD.n1365 VDD.n1363 0.0249681
R17994 VDD.n1525 VDD.n1523 0.0249681
R17995 VDD.n1523 VDD.n1519 0.0249681
R17996 VDD.n1519 VDD.n1517 0.0249681
R17997 VDD.n1517 VDD.n1513 0.0249681
R17998 VDD.n1503 VDD.n1501 0.0249681
R17999 VDD.n1501 VDD.n1497 0.0249681
R18000 VDD.n1497 VDD.n1495 0.0249681
R18001 VDD.n1495 VDD.n1491 0.0249681
R18002 VDD.n1491 VDD.n1489 0.0249681
R18003 VDD.n1489 VDD.n1485 0.0249681
R18004 VDD.n1485 VDD.n1481 0.0249681
R18005 VDD.n1481 VDD.n1479 0.0249681
R18006 VDD.n1479 VDD.n1475 0.0249681
R18007 VDD.n1475 VDD.n1473 0.0249681
R18008 VDD.n1473 VDD.n1469 0.0249681
R18009 VDD.n1469 VDD.n1467 0.0249681
R18010 VDD.n1467 VDD.n1463 0.0249681
R18011 VDD.n1286 VDD.n1285 0.0249681
R18012 VDD.n1285 VDD.n1283 0.0249681
R18013 VDD.n1546 VDD.n1544 0.0243281
R18014 VDD.n1454 VDD.n1453 0.0241145
R18015 VDD.n5345 VDD.n5084 0.0238663
R18016 VDD.n5858 VDD.n5857 0.0228694
R18017 VDD.n5604 VDD.n5603 0.0228694
R18018 VDD.n1882 VDD.n1881 0.0228205
R18019 VDD.n2203 VDD.n2202 0.0228205
R18020 VDD.n2461 VDD.n2460 0.0228205
R18021 VDD.n2719 VDD.n2718 0.0228205
R18022 VDD.n2977 VDD.n2976 0.0228205
R18023 VDD.n3235 VDD.n3234 0.0228205
R18024 VDD.n3493 VDD.n3492 0.0228205
R18025 VDD.n5820 VDD.n5819 0.0228205
R18026 VDD.n5566 VDD.n5565 0.0228205
R18027 VDD.n3751 VDD.n3750 0.0228205
R18028 VDD.n4009 VDD.n4008 0.0228205
R18029 VDD.n4267 VDD.n4266 0.0228205
R18030 VDD.n4525 VDD.n4524 0.0228205
R18031 VDD.n4783 VDD.n4782 0.0228205
R18032 VDD.n5044 VDD.n5043 0.0228205
R18033 VDD.n5306 VDD.n5305 0.0228205
R18034 VDD.n1881 VDD.n1820 0.0223212
R18035 VDD.n2202 VDD.n2141 0.0223212
R18036 VDD.n2460 VDD.n2399 0.0223212
R18037 VDD.n2718 VDD.n2657 0.0223212
R18038 VDD.n2976 VDD.n2915 0.0223212
R18039 VDD.n3234 VDD.n3173 0.0223212
R18040 VDD.n3492 VDD.n3431 0.0223212
R18041 VDD.n5819 VDD.n5758 0.0223212
R18042 VDD.n5565 VDD.n5504 0.0223212
R18043 VDD.n3750 VDD.n3689 0.0223212
R18044 VDD.n4008 VDD.n3947 0.0223212
R18045 VDD.n4266 VDD.n4205 0.0223212
R18046 VDD.n4524 VDD.n4463 0.0223212
R18047 VDD.n4782 VDD.n4721 0.0223212
R18048 VDD.n5043 VDD.n4982 0.0223212
R18049 VDD.n5305 VDD.n5244 0.0223212
R18050 VDD.n1374 VDD.n1346 0.0218724
R18051 VDD.n1168 VDD 0.02175
R18052 VDD.n1162 VDD 0.02175
R18053 VDD.n1156 VDD 0.02175
R18054 VDD.n1150 VDD 0.02175
R18055 VDD.n1144 VDD 0.02175
R18056 VDD.n1234 VDD 0.02175
R18057 VDD.n1228 VDD 0.02175
R18058 VDD.n1222 VDD 0.02175
R18059 VDD.n1216 VDD 0.02175
R18060 VDD.n1210 VDD 0.02175
R18061 VDD.n1600 VDD 0.0213145
R18062 VDD.n1410 VDD.n1406 0.0212447
R18063 VDD.n1504 VDD.n1503 0.0207128
R18064 VDD.n1622 VDD.n1621 0.0205312
R18065 VDD.n1433 VDD.n1431 0.0198592
R18066 VDD.n1461 VDD.n1460 0.0188511
R18067 VDD.n5226 VDD.n5225 0.0185136
R18068 VDD.n1946 VDD.n1945 0.0183679
R18069 VDD.n1799 VDD.n1798 0.0182941
R18070 VDD.n2007 VDD.n2006 0.0182941
R18071 VDD.n2378 VDD.n2377 0.0182941
R18072 VDD.n2636 VDD.n2635 0.0182941
R18073 VDD.n2894 VDD.n2893 0.0182941
R18074 VDD.n3152 VDD.n3151 0.0182941
R18075 VDD.n3410 VDD.n3409 0.0182941
R18076 VDD.n5740 VDD.n5739 0.0182941
R18077 VDD.n5486 VDD.n5485 0.0182941
R18078 VDD.n3668 VDD.n3667 0.0182941
R18079 VDD.n3926 VDD.n3925 0.0182941
R18080 VDD.n4184 VDD.n4183 0.0182941
R18081 VDD.n4442 VDD.n4441 0.0182941
R18082 VDD.n4700 VDD.n4699 0.0182941
R18083 VDD.n4959 VDD.n4958 0.0182941
R18084 VDD.n5109 VDD.n5108 0.0182941
R18085 VDD.n1779 VDD.n1777 0.0178611
R18086 VDD.n1987 VDD.n1985 0.0178611
R18087 VDD.n2358 VDD.n2356 0.0178611
R18088 VDD.n2616 VDD.n2614 0.0178611
R18089 VDD.n2874 VDD.n2872 0.0178611
R18090 VDD.n3132 VDD.n3130 0.0178611
R18091 VDD.n3390 VDD.n3388 0.0178611
R18092 VDD.n5720 VDD.n5718 0.0178611
R18093 VDD.n5466 VDD.n5464 0.0178611
R18094 VDD.n3648 VDD.n3646 0.0178611
R18095 VDD.n3906 VDD.n3904 0.0178611
R18096 VDD.n4164 VDD.n4162 0.0178611
R18097 VDD.n4422 VDD.n4420 0.0178611
R18098 VDD.n4680 VDD.n4678 0.0178611
R18099 VDD.n4939 VDD.n4937 0.0178611
R18100 VDD.n5089 VDD.n5087 0.0178611
R18101 VDD.n1808 VDD.n1807 0.0177731
R18102 VDD.n2387 VDD.n2386 0.0177731
R18103 VDD.n2645 VDD.n2644 0.0177731
R18104 VDD.n2903 VDD.n2902 0.0177731
R18105 VDD.n3161 VDD.n3160 0.0177731
R18106 VDD.n3419 VDD.n3418 0.0177731
R18107 VDD.n3677 VDD.n3676 0.0177731
R18108 VDD.n3935 VDD.n3934 0.0177731
R18109 VDD.n4193 VDD.n4192 0.0177731
R18110 VDD.n4451 VDD.n4450 0.0177731
R18111 VDD.n4709 VDD.n4708 0.0177731
R18112 VDD.n1368 VDD.n1366 0.0172553
R18113 VDD.n5859 VDD.n5605 0.0171851
R18114 VDD.n1127 VDD 0.0171185
R18115 VDD VDD.n1116 0.0171185
R18116 VDD.n1193 VDD 0.0171185
R18117 VDD VDD.n1182 0.0171185
R18118 VDD.n1758 VDD.n1757 0.0168386
R18119 VDD.n2107 VDD.n2106 0.0168386
R18120 VDD.n2337 VDD.n2336 0.0168386
R18121 VDD.n2595 VDD.n2594 0.0168386
R18122 VDD.n2853 VDD.n2852 0.0168386
R18123 VDD.n3111 VDD.n3110 0.0168386
R18124 VDD.n3369 VDD.n3368 0.0168386
R18125 VDD.n5699 VDD.n5698 0.0168386
R18126 VDD.n5445 VDD.n5444 0.0168386
R18127 VDD.n3627 VDD.n3626 0.0168386
R18128 VDD.n3885 VDD.n3884 0.0168386
R18129 VDD.n4143 VDD.n4142 0.0168386
R18130 VDD.n4401 VDD.n4400 0.0168386
R18131 VDD.n4659 VDD.n4658 0.0168386
R18132 VDD.n4917 VDD.n4916 0.0168386
R18133 VDD.n5209 VDD.n5208 0.0168386
R18134 VDD.n1710 VDD.n1679 0.0168372
R18135 VDD.n2059 VDD.n2028 0.0168372
R18136 VDD.n2289 VDD.n2258 0.0168372
R18137 VDD.n2547 VDD.n2516 0.0168372
R18138 VDD.n2805 VDD.n2774 0.0168372
R18139 VDD.n3063 VDD.n3032 0.0168372
R18140 VDD.n3321 VDD.n3290 0.0168372
R18141 VDD.n5651 VDD.n5620 0.0168372
R18142 VDD.n5397 VDD.n5366 0.0168372
R18143 VDD.n3579 VDD.n3548 0.0168372
R18144 VDD.n3837 VDD.n3806 0.0168372
R18145 VDD.n4095 VDD.n4064 0.0168372
R18146 VDD.n4353 VDD.n4322 0.0168372
R18147 VDD.n4611 VDD.n4580 0.0168372
R18148 VDD.n4869 VDD.n4838 0.0168372
R18149 VDD.n5161 VDD.n5130 0.0168372
R18150 VDD.n1178 VDD.n1177 0.0165987
R18151 VDD.n1244 VDD.n1243 0.0165987
R18152 VDD.n5860 VDD.n5859 0.0164899
R18153 VDD.n1679 VDD.n1669 0.0163404
R18154 VDD.n1758 VDD.n1717 0.0163404
R18155 VDD.n2028 VDD.n2018 0.0163404
R18156 VDD.n2107 VDD.n2066 0.0163404
R18157 VDD.n2258 VDD.n2248 0.0163404
R18158 VDD.n2337 VDD.n2296 0.0163404
R18159 VDD.n2516 VDD.n2506 0.0163404
R18160 VDD.n2595 VDD.n2554 0.0163404
R18161 VDD.n2774 VDD.n2764 0.0163404
R18162 VDD.n2853 VDD.n2812 0.0163404
R18163 VDD.n3032 VDD.n3022 0.0163404
R18164 VDD.n3111 VDD.n3070 0.0163404
R18165 VDD.n3290 VDD.n3280 0.0163404
R18166 VDD.n3369 VDD.n3328 0.0163404
R18167 VDD.n5620 VDD.n5610 0.0163404
R18168 VDD.n5699 VDD.n5658 0.0163404
R18169 VDD.n5366 VDD.n5356 0.0163404
R18170 VDD.n5445 VDD.n5404 0.0163404
R18171 VDD.n3548 VDD.n3538 0.0163404
R18172 VDD.n3627 VDD.n3586 0.0163404
R18173 VDD.n3806 VDD.n3796 0.0163404
R18174 VDD.n3885 VDD.n3844 0.0163404
R18175 VDD.n4064 VDD.n4054 0.0163404
R18176 VDD.n4143 VDD.n4102 0.0163404
R18177 VDD.n4322 VDD.n4312 0.0163404
R18178 VDD.n4401 VDD.n4360 0.0163404
R18179 VDD.n4580 VDD.n4570 0.0163404
R18180 VDD.n4659 VDD.n4618 0.0163404
R18181 VDD.n4838 VDD.n4828 0.0163404
R18182 VDD.n4917 VDD.n4876 0.0163404
R18183 VDD.n5130 VDD.n5120 0.0163404
R18184 VDD.n5209 VDD.n5168 0.0163404
R18185 VDD.n1423 VDD.n1422 0.0161915
R18186 VDD.n1172 VDD.n1171 0.016125
R18187 VDD.n1238 VDD.n1237 0.016125
R18188 VDD.n5605 VDD.n5351 0.0161096
R18189 VDD.n1961 VDD.n1941 0.0154506
R18190 VDD.n1969 VDD.n1968 0.015449
R18191 VDD.n5865 VDD.n5864 0.0154143
R18192 VDD.n5864 VDD.n5863 0.0154143
R18193 VDD.n5863 VDD.n5862 0.0154143
R18194 VDD.n5862 VDD.n5861 0.0154143
R18195 VDD.n5861 VDD.n5860 0.0154143
R18196 VDD.n5351 VDD.n5350 0.0154143
R18197 VDD.n5350 VDD.n5349 0.0154143
R18198 VDD.n5349 VDD.n5348 0.0154143
R18199 VDD.n5348 VDD.n5347 0.0154143
R18200 VDD.n5347 VDD.n5346 0.0154143
R18201 VDD.n1405 VDD.n1401 0.0153936
R18202 VDD.n1513 VDD.n1511 0.0151277
R18203 VDD.n1971 VDD.n1970 0.0150463
R18204 VDD.n1970 VDD.t1287 0.0150463
R18205 VDD.n1963 VDD.n1929 0.0150463
R18206 VDD.t1055 VDD.n1963 0.0150463
R18207 VDD.n1961 VDD.n1960 0.0150463
R18208 VDD.n1964 VDD.t1055 0.0150463
R18209 VDD.n1968 VDD.n1967 0.0150463
R18210 VDD.n1965 VDD.n1964 0.0150463
R18211 VDD.t1285 VDD.n1951 0.0150463
R18212 VDD.n1951 VDD.n1950 0.0150463
R18213 VDD.n1111 VDD.n830 0.015
R18214 VDD.n1839 VDD.n1827 0.0149834
R18215 VDD.n2160 VDD.n2148 0.0149834
R18216 VDD.n2418 VDD.n2406 0.0149834
R18217 VDD.n2676 VDD.n2664 0.0149834
R18218 VDD.n2934 VDD.n2922 0.0149834
R18219 VDD.n3192 VDD.n3180 0.0149834
R18220 VDD.n3450 VDD.n3438 0.0149834
R18221 VDD.n5777 VDD.n5765 0.0149834
R18222 VDD.n5523 VDD.n5511 0.0149834
R18223 VDD.n3708 VDD.n3696 0.0149834
R18224 VDD.n3966 VDD.n3954 0.0149834
R18225 VDD.n4224 VDD.n4212 0.0149834
R18226 VDD.n4482 VDD.n4470 0.0149834
R18227 VDD.n4740 VDD.n4728 0.0149834
R18228 VDD.n5001 VDD.n4989 0.0149834
R18229 VDD.n5263 VDD.n5251 0.0149834
R18230 VDD.n1325 VDD.n1324 0.0148617
R18231 VDD.n5867 VDD.n5866 0.0147238
R18232 VDD.n993 VDD.n991 0.0146339
R18233 VDD.n198 VDD.n196 0.0146339
R18234 VDD.n588 VDD.n586 0.0146339
R18235 VDD.n1394 VDD.n1393 0.0145957
R18236 VDD.n1377 VDD.n1376 0.0145957
R18237 VDD.n1886 VDD.n1817 0.0145797
R18238 VDD.n2207 VDD.n2138 0.0145797
R18239 VDD.n2465 VDD.n2396 0.0145797
R18240 VDD.n2723 VDD.n2654 0.0145797
R18241 VDD.n2981 VDD.n2912 0.0145797
R18242 VDD.n3239 VDD.n3170 0.0145797
R18243 VDD.n3497 VDD.n3428 0.0145797
R18244 VDD.n5824 VDD.n5755 0.0145797
R18245 VDD.n5570 VDD.n5501 0.0145797
R18246 VDD.n3755 VDD.n3686 0.0145797
R18247 VDD.n4013 VDD.n3944 0.0145797
R18248 VDD.n4271 VDD.n4202 0.0145797
R18249 VDD.n4529 VDD.n4460 0.0145797
R18250 VDD.n4787 VDD.n4718 0.0145797
R18251 VDD.n5048 VDD.n4979 0.0145797
R18252 VDD.n5310 VDD.n5241 0.0145797
R18253 VDD.n1721 VDD.n1720 0.0143889
R18254 VDD.n2070 VDD.n2069 0.0143889
R18255 VDD.n2300 VDD.n2299 0.0143889
R18256 VDD.n2558 VDD.n2557 0.0143889
R18257 VDD.n2816 VDD.n2815 0.0143889
R18258 VDD.n3074 VDD.n3073 0.0143889
R18259 VDD.n3332 VDD.n3331 0.0143889
R18260 VDD.n5662 VDD.n5661 0.0143889
R18261 VDD.n5408 VDD.n5407 0.0143889
R18262 VDD.n3590 VDD.n3589 0.0143889
R18263 VDD.n3848 VDD.n3847 0.0143889
R18264 VDD.n4106 VDD.n4105 0.0143889
R18265 VDD.n4364 VDD.n4363 0.0143889
R18266 VDD.n4622 VDD.n4621 0.0143889
R18267 VDD.n4880 VDD.n4879 0.0143889
R18268 VDD.n5172 VDD.n5171 0.0143889
R18269 VDD.n802 VDD.n798 0.0143889
R18270 VDD.n400 VDD.n396 0.0143889
R18271 VDD.n1308 VDD.n1304 0.0143298
R18272 VDD.n352 VDD.n316 0.0142984
R18273 VDD.n5858 VDD.n5716 0.0142906
R18274 VDD.n5604 VDD.n5462 0.0142906
R18275 VDD.n1979 VDD.n1978 0.0138929
R18276 VDD.n1345 VDD.n1343 0.0137979
R18277 VDD VDD.n1840 0.0131689
R18278 VDD VDD.n2161 0.0131689
R18279 VDD VDD.n2419 0.0131689
R18280 VDD VDD.n2677 0.0131689
R18281 VDD VDD.n2935 0.0131689
R18282 VDD VDD.n3193 0.0131689
R18283 VDD VDD.n3451 0.0131689
R18284 VDD VDD.n5778 0.0131689
R18285 VDD VDD.n5524 0.0131689
R18286 VDD VDD.n3709 0.0131689
R18287 VDD VDD.n3967 0.0131689
R18288 VDD VDD.n4225 0.0131689
R18289 VDD VDD.n4483 0.0131689
R18290 VDD VDD.n4741 0.0131689
R18291 VDD VDD.n5002 0.0131689
R18292 VDD VDD.n5264 0.0131689
R18293 VDD.n764 VDD 0.013
R18294 VDD.n361 VDD 0.013
R18295 VDD.n1314 VDD 0.012734
R18296 VDD.n1349 VDD 0.012734
R18297 VDD.n1261 VDD 0.012734
R18298 VDD.n1544 VDD.n1543 0.0126094
R18299 VDD.n854 VDD.n850 0.0126053
R18300 VDD.n893 VDD.n889 0.0126053
R18301 VDD.n889 VDD.n887 0.0126053
R18302 VDD.n887 VDD.n883 0.0126053
R18303 VDD.n883 VDD.n881 0.0126053
R18304 VDD.n881 VDD.n877 0.0126053
R18305 VDD.n877 VDD.n875 0.0126053
R18306 VDD.n875 VDD.n871 0.0126053
R18307 VDD.n871 VDD.n869 0.0126053
R18308 VDD.n868 VDD.n867 0.0126053
R18309 VDD.n867 VDD.n865 0.0126053
R18310 VDD.n865 VDD.n861 0.0126053
R18311 VDD.n861 VDD.n845 0.0126053
R18312 VDD.n915 VDD.n911 0.0126053
R18313 VDD.n917 VDD.n915 0.0126053
R18314 VDD.n921 VDD.n917 0.0126053
R18315 VDD.n923 VDD.n921 0.0126053
R18316 VDD.n927 VDD.n923 0.0126053
R18317 VDD.n929 VDD.n927 0.0126053
R18318 VDD.n933 VDD.n929 0.0126053
R18319 VDD.n935 VDD.n933 0.0126053
R18320 VDD.n936 VDD.n935 0.0126053
R18321 VDD.n941 VDD.n939 0.0126053
R18322 VDD.n945 VDD.n941 0.0126053
R18323 VDD.n947 VDD.n945 0.0126053
R18324 VDD.n951 VDD.n947 0.0126053
R18325 VDD.n976 VDD.n972 0.0126053
R18326 VDD.n972 VDD.n970 0.0126053
R18327 VDD.n970 VDD.n966 0.0126053
R18328 VDD.n966 VDD.n964 0.0126053
R18329 VDD.n964 VDD.n960 0.0126053
R18330 VDD.n960 VDD.n958 0.0126053
R18331 VDD.n958 VDD.n832 0.0126053
R18332 VDD.n1108 VDD.n1107 0.0126053
R18333 VDD.n1107 VDD.n1105 0.0126053
R18334 VDD.n1092 VDD.n1090 0.0126053
R18335 VDD.n1090 VDD.n1086 0.0126053
R18336 VDD.n1086 VDD.n1082 0.0126053
R18337 VDD.n1082 VDD.n1080 0.0126053
R18338 VDD.n1080 VDD.n1076 0.0126053
R18339 VDD.n1076 VDD.n1074 0.0126053
R18340 VDD.n1074 VDD.n1070 0.0126053
R18341 VDD.n1070 VDD.n1068 0.0126053
R18342 VDD.n1068 VDD.n1064 0.0126053
R18343 VDD.n1064 VDD.n1062 0.0126053
R18344 VDD.n1061 VDD.n1060 0.0126053
R18345 VDD.n1049 VDD.n1045 0.0126053
R18346 VDD.n1045 VDD.n1043 0.0126053
R18347 VDD.n1043 VDD.n1039 0.0126053
R18348 VDD.n1039 VDD.n1035 0.0126053
R18349 VDD.n1035 VDD.n1033 0.0126053
R18350 VDD.n1033 VDD.n1029 0.0126053
R18351 VDD.n1029 VDD.n1027 0.0126053
R18352 VDD.n1027 VDD.n1023 0.0126053
R18353 VDD.n1023 VDD.n1021 0.0126053
R18354 VDD.n1021 VDD.n1017 0.0126053
R18355 VDD.n1017 VDD.n1015 0.0126053
R18356 VDD.n1014 VDD.n1013 0.0126053
R18357 VDD.n1013 VDD.n1011 0.0126053
R18358 VDD.n1011 VDD.n1008 0.0126053
R18359 VDD.n1008 VDD.n1006 0.0126053
R18360 VDD.n999 VDD.n997 0.0126053
R18361 VDD.n994 VDD.n993 0.0126053
R18362 VDD.n59 VDD.n55 0.0126053
R18363 VDD.n98 VDD.n94 0.0126053
R18364 VDD.n94 VDD.n92 0.0126053
R18365 VDD.n92 VDD.n88 0.0126053
R18366 VDD.n88 VDD.n86 0.0126053
R18367 VDD.n86 VDD.n82 0.0126053
R18368 VDD.n82 VDD.n80 0.0126053
R18369 VDD.n80 VDD.n76 0.0126053
R18370 VDD.n76 VDD.n74 0.0126053
R18371 VDD.n73 VDD.n72 0.0126053
R18372 VDD.n72 VDD.n70 0.0126053
R18373 VDD.n70 VDD.n66 0.0126053
R18374 VDD.n66 VDD.n50 0.0126053
R18375 VDD.n120 VDD.n116 0.0126053
R18376 VDD.n122 VDD.n120 0.0126053
R18377 VDD.n126 VDD.n122 0.0126053
R18378 VDD.n128 VDD.n126 0.0126053
R18379 VDD.n132 VDD.n128 0.0126053
R18380 VDD.n134 VDD.n132 0.0126053
R18381 VDD.n138 VDD.n134 0.0126053
R18382 VDD.n140 VDD.n138 0.0126053
R18383 VDD.n141 VDD.n140 0.0126053
R18384 VDD.n146 VDD.n144 0.0126053
R18385 VDD.n150 VDD.n146 0.0126053
R18386 VDD.n152 VDD.n150 0.0126053
R18387 VDD.n156 VDD.n152 0.0126053
R18388 VDD.n181 VDD.n177 0.0126053
R18389 VDD.n177 VDD.n175 0.0126053
R18390 VDD.n175 VDD.n171 0.0126053
R18391 VDD.n171 VDD.n169 0.0126053
R18392 VDD.n169 VDD.n165 0.0126053
R18393 VDD.n165 VDD.n163 0.0126053
R18394 VDD.n163 VDD.n37 0.0126053
R18395 VDD.n313 VDD.n312 0.0126053
R18396 VDD.n312 VDD.n310 0.0126053
R18397 VDD.n297 VDD.n295 0.0126053
R18398 VDD.n295 VDD.n291 0.0126053
R18399 VDD.n291 VDD.n287 0.0126053
R18400 VDD.n287 VDD.n285 0.0126053
R18401 VDD.n285 VDD.n281 0.0126053
R18402 VDD.n281 VDD.n279 0.0126053
R18403 VDD.n279 VDD.n275 0.0126053
R18404 VDD.n275 VDD.n273 0.0126053
R18405 VDD.n273 VDD.n269 0.0126053
R18406 VDD.n269 VDD.n267 0.0126053
R18407 VDD.n266 VDD.n265 0.0126053
R18408 VDD.n254 VDD.n250 0.0126053
R18409 VDD.n250 VDD.n248 0.0126053
R18410 VDD.n248 VDD.n244 0.0126053
R18411 VDD.n244 VDD.n240 0.0126053
R18412 VDD.n240 VDD.n238 0.0126053
R18413 VDD.n238 VDD.n234 0.0126053
R18414 VDD.n234 VDD.n232 0.0126053
R18415 VDD.n232 VDD.n228 0.0126053
R18416 VDD.n228 VDD.n226 0.0126053
R18417 VDD.n226 VDD.n222 0.0126053
R18418 VDD.n222 VDD.n220 0.0126053
R18419 VDD.n219 VDD.n218 0.0126053
R18420 VDD.n218 VDD.n216 0.0126053
R18421 VDD.n216 VDD.n213 0.0126053
R18422 VDD.n213 VDD.n211 0.0126053
R18423 VDD.n204 VDD.n202 0.0126053
R18424 VDD.n199 VDD.n198 0.0126053
R18425 VDD.n453 VDD.n449 0.0126053
R18426 VDD.n492 VDD.n488 0.0126053
R18427 VDD.n488 VDD.n486 0.0126053
R18428 VDD.n486 VDD.n482 0.0126053
R18429 VDD.n482 VDD.n480 0.0126053
R18430 VDD.n480 VDD.n476 0.0126053
R18431 VDD.n476 VDD.n474 0.0126053
R18432 VDD.n474 VDD.n470 0.0126053
R18433 VDD.n470 VDD.n468 0.0126053
R18434 VDD.n467 VDD.n466 0.0126053
R18435 VDD.n466 VDD.n464 0.0126053
R18436 VDD.n464 VDD.n460 0.0126053
R18437 VDD.n460 VDD.n444 0.0126053
R18438 VDD.n514 VDD.n510 0.0126053
R18439 VDD.n516 VDD.n514 0.0126053
R18440 VDD.n520 VDD.n516 0.0126053
R18441 VDD.n522 VDD.n520 0.0126053
R18442 VDD.n526 VDD.n522 0.0126053
R18443 VDD.n528 VDD.n526 0.0126053
R18444 VDD.n532 VDD.n528 0.0126053
R18445 VDD.n534 VDD.n532 0.0126053
R18446 VDD.n535 VDD.n534 0.0126053
R18447 VDD.n540 VDD.n538 0.0126053
R18448 VDD.n544 VDD.n540 0.0126053
R18449 VDD.n546 VDD.n544 0.0126053
R18450 VDD.n550 VDD.n546 0.0126053
R18451 VDD.n571 VDD.n567 0.0126053
R18452 VDD.n567 VDD.n565 0.0126053
R18453 VDD.n565 VDD.n561 0.0126053
R18454 VDD.n561 VDD.n559 0.0126053
R18455 VDD.n559 VDD.n555 0.0126053
R18456 VDD.n555 VDD.n431 0.0126053
R18457 VDD.n706 VDD.n704 0.0126053
R18458 VDD.n703 VDD.n702 0.0126053
R18459 VDD.n702 VDD.n700 0.0126053
R18460 VDD.n687 VDD.n685 0.0126053
R18461 VDD.n685 VDD.n681 0.0126053
R18462 VDD.n681 VDD.n677 0.0126053
R18463 VDD.n677 VDD.n675 0.0126053
R18464 VDD.n675 VDD.n671 0.0126053
R18465 VDD.n671 VDD.n669 0.0126053
R18466 VDD.n669 VDD.n665 0.0126053
R18467 VDD.n665 VDD.n663 0.0126053
R18468 VDD.n663 VDD.n659 0.0126053
R18469 VDD.n659 VDD.n657 0.0126053
R18470 VDD.n656 VDD.n655 0.0126053
R18471 VDD.n644 VDD.n640 0.0126053
R18472 VDD.n640 VDD.n638 0.0126053
R18473 VDD.n638 VDD.n634 0.0126053
R18474 VDD.n634 VDD.n630 0.0126053
R18475 VDD.n630 VDD.n628 0.0126053
R18476 VDD.n628 VDD.n624 0.0126053
R18477 VDD.n624 VDD.n622 0.0126053
R18478 VDD.n622 VDD.n618 0.0126053
R18479 VDD.n618 VDD.n616 0.0126053
R18480 VDD.n616 VDD.n612 0.0126053
R18481 VDD.n612 VDD.n610 0.0126053
R18482 VDD.n609 VDD.n608 0.0126053
R18483 VDD.n608 VDD.n606 0.0126053
R18484 VDD.n606 VDD.n603 0.0126053
R18485 VDD.n603 VDD.n601 0.0126053
R18486 VDD.n594 VDD.n592 0.0126053
R18487 VDD.n589 VDD.n588 0.0126053
R18488 VDD.n791 VDD 0.0125739
R18489 VDD.n389 VDD 0.0125739
R18490 VDD.n1611 VDD.n1609 0.0125192
R18491 VDD.n1110 VDD.n1109 0.0124737
R18492 VDD.n315 VDD.n314 0.0124737
R18493 VDD.n1785 VDD 0.0123056
R18494 VDD.n1993 VDD 0.0123056
R18495 VDD.n2364 VDD 0.0123056
R18496 VDD.n2622 VDD 0.0123056
R18497 VDD.n2880 VDD 0.0123056
R18498 VDD.n3138 VDD 0.0123056
R18499 VDD.n3396 VDD 0.0123056
R18500 VDD.n5726 VDD 0.0123056
R18501 VDD.n5472 VDD 0.0123056
R18502 VDD.n3654 VDD 0.0123056
R18503 VDD.n3912 VDD 0.0123056
R18504 VDD.n4170 VDD 0.0123056
R18505 VDD.n4428 VDD 0.0123056
R18506 VDD.n4686 VDD 0.0123056
R18507 VDD.n4945 VDD 0.0123056
R18508 VDD.n5095 VDD 0.0123056
R18509 VDD VDD.n784 0.0123056
R18510 VDD.n730 VDD 0.0123056
R18511 VDD VDD.n382 0.0123056
R18512 VDD.n1571 VDD 0.0123056
R18513 VDD.n707 VDD.n431 0.0122105
R18514 VDD.n4967 VDD.n4935 0.0121683
R18515 VDD.n904 VDD.n845 0.0119152
R18516 VDD.n109 VDD.n50 0.0119152
R18517 VDD.n1842 VDD 0.0118881
R18518 VDD.n2163 VDD 0.0118881
R18519 VDD.n2421 VDD 0.0118881
R18520 VDD.n2679 VDD 0.0118881
R18521 VDD.n2937 VDD 0.0118881
R18522 VDD.n3195 VDD 0.0118881
R18523 VDD.n3453 VDD 0.0118881
R18524 VDD.n5780 VDD 0.0118881
R18525 VDD.n5526 VDD 0.0118881
R18526 VDD.n3711 VDD 0.0118881
R18527 VDD.n3969 VDD 0.0118881
R18528 VDD.n4227 VDD 0.0118881
R18529 VDD.n4485 VDD 0.0118881
R18530 VDD.n4743 VDD 0.0118881
R18531 VDD.n5004 VDD 0.0118881
R18532 VDD.n5266 VDD 0.0118881
R18533 VDD.n1255 VDD.n1251 0.0117745
R18534 VDD.n1539 VDD.n1537 0.0117745
R18535 VDD.n1537 VDD.n1533 0.0117745
R18536 VDD.n1533 VDD.n1529 0.0117745
R18537 VDD.n1529 VDD.n1527 0.0117745
R18538 VDD.n1613 VDD.n1611 0.0117367
R18539 VDD.n818 VDD 0.0116111
R18540 VDD.n745 VDD 0.0116111
R18541 VDD.n711 VDD 0.0116111
R18542 VDD.n416 VDD 0.0116111
R18543 VDD.n1586 VDD 0.0116111
R18544 VDD.n1552 VDD 0.0116111
R18545 VDD.n11 VDD 0.0114012
R18546 VDD.n328 VDD 0.0114012
R18547 VDD.n503 VDD.n444 0.0113889
R18548 VDD.n1875 VDD.n1874 0.0111456
R18549 VDD.n2196 VDD.n2195 0.0111456
R18550 VDD.n2454 VDD.n2453 0.0111456
R18551 VDD.n2712 VDD.n2711 0.0111456
R18552 VDD.n2970 VDD.n2969 0.0111456
R18553 VDD.n3228 VDD.n3227 0.0111456
R18554 VDD.n3486 VDD.n3485 0.0111456
R18555 VDD.n5813 VDD.n5812 0.0111456
R18556 VDD.n5559 VDD.n5558 0.0111456
R18557 VDD.n3744 VDD.n3743 0.0111456
R18558 VDD.n4002 VDD.n4001 0.0111456
R18559 VDD.n4260 VDD.n4259 0.0111456
R18560 VDD.n4518 VDD.n4517 0.0111456
R18561 VDD.n4776 VDD.n4775 0.0111456
R18562 VDD.n5037 VDD.n5036 0.0111456
R18563 VDD.n5299 VDD.n5298 0.0111456
R18564 VDD.n572 VDD.n571 0.0108947
R18565 VDD.n1396 VDD.n1394 0.0108723
R18566 VDD.n1381 VDD.n1377 0.0108723
R18567 VDD.n1957 VDD.n1922 0.0108144
R18568 VDD.n688 VDD.n687 0.0106316
R18569 VDD.n645 VDD.n644 0.0106316
R18570 VDD.n1327 VDD.n1325 0.0106064
R18571 VDD.n855 VDD.n854 0.0103684
R18572 VDD.n977 VDD.n976 0.0103684
R18573 VDD.n60 VDD.n59 0.0103684
R18574 VDD.n182 VDD.n181 0.0103684
R18575 VDD.n1426 VDD.n1425 0.0103404
R18576 VDD.n1511 VDD.n1510 0.0103404
R18577 VDD.n1527 VDD.n1526 0.0103039
R18578 VDD.n1696 VDD.n1695 0.0101514
R18579 VDD.n2045 VDD.n2044 0.0101514
R18580 VDD.n2275 VDD.n2274 0.0101514
R18581 VDD.n2533 VDD.n2532 0.0101514
R18582 VDD.n2791 VDD.n2790 0.0101514
R18583 VDD.n3049 VDD.n3048 0.0101514
R18584 VDD.n3307 VDD.n3306 0.0101514
R18585 VDD.n5637 VDD.n5636 0.0101514
R18586 VDD.n5383 VDD.n5382 0.0101514
R18587 VDD.n3565 VDD.n3564 0.0101514
R18588 VDD.n3823 VDD.n3822 0.0101514
R18589 VDD.n4081 VDD.n4080 0.0101514
R18590 VDD.n4339 VDD.n4338 0.0101514
R18591 VDD.n4597 VDD.n4596 0.0101514
R18592 VDD.n4855 VDD.n4854 0.0101514
R18593 VDD.n5147 VDD.n5146 0.0101514
R18594 VDD.n1093 VDD.n1092 0.0101053
R18595 VDD.n1050 VDD.n1049 0.0101053
R18596 VDD.n298 VDD.n297 0.0101053
R18597 VDD.n255 VDD.n254 0.0101053
R18598 VDD.n1883 VDD.n1882 0.0101
R18599 VDD.n2204 VDD.n2203 0.0101
R18600 VDD.n2462 VDD.n2461 0.0101
R18601 VDD.n2720 VDD.n2719 0.0101
R18602 VDD.n2978 VDD.n2977 0.0101
R18603 VDD.n3236 VDD.n3235 0.0101
R18604 VDD.n3494 VDD.n3493 0.0101
R18605 VDD.n5821 VDD.n5820 0.0101
R18606 VDD.n5567 VDD.n5566 0.0101
R18607 VDD.n3752 VDD.n3751 0.0101
R18608 VDD.n4010 VDD.n4009 0.0101
R18609 VDD.n4268 VDD.n4267 0.0101
R18610 VDD.n4526 VDD.n4525 0.0101
R18611 VDD.n4784 VDD.n4783 0.0101
R18612 VDD.n5045 VDD.n5044 0.0101
R18613 VDD.n5307 VDD.n5306 0.0101
R18614 VDD.n1597 VDD.n1181 0.00985484
R18615 VDD.n454 VDD.n453 0.00984211
R18616 VDD.n2129 VDD.n2128 0.00977468
R18617 VDD.n1884 VDD.n1883 0.0096003
R18618 VDD.n1870 VDD.n1869 0.0096003
R18619 VDD.n1869 VDD.t355 0.0096003
R18620 VDD.n2191 VDD.n2190 0.0096003
R18621 VDD.n2190 VDD.t574 0.0096003
R18622 VDD.n2205 VDD.n2204 0.0096003
R18623 VDD.n2449 VDD.n2448 0.0096003
R18624 VDD.n2448 VDD.t103 0.0096003
R18625 VDD.n2463 VDD.n2462 0.0096003
R18626 VDD.n2707 VDD.n2706 0.0096003
R18627 VDD.n2706 VDD.t421 0.0096003
R18628 VDD.n2721 VDD.n2720 0.0096003
R18629 VDD.n2965 VDD.n2964 0.0096003
R18630 VDD.n2964 VDD.t405 0.0096003
R18631 VDD.n2979 VDD.n2978 0.0096003
R18632 VDD.n3223 VDD.n3222 0.0096003
R18633 VDD.n3222 VDD.t144 0.0096003
R18634 VDD.n3237 VDD.n3236 0.0096003
R18635 VDD.n3481 VDD.n3480 0.0096003
R18636 VDD.n3480 VDD.t179 0.0096003
R18637 VDD.n3495 VDD.n3494 0.0096003
R18638 VDD.n5808 VDD.n5807 0.0096003
R18639 VDD.n5807 VDD.t1088 0.0096003
R18640 VDD.n5822 VDD.n5821 0.0096003
R18641 VDD.n5554 VDD.n5553 0.0096003
R18642 VDD.n5553 VDD.t596 0.0096003
R18643 VDD.n5568 VDD.n5567 0.0096003
R18644 VDD.n3739 VDD.n3738 0.0096003
R18645 VDD.n3738 VDD.t145 0.0096003
R18646 VDD.n3753 VDD.n3752 0.0096003
R18647 VDD.n3997 VDD.n3996 0.0096003
R18648 VDD.n3996 VDD.t563 0.0096003
R18649 VDD.n4011 VDD.n4010 0.0096003
R18650 VDD.n4255 VDD.n4254 0.0096003
R18651 VDD.n4254 VDD.t668 0.0096003
R18652 VDD.n4269 VDD.n4268 0.0096003
R18653 VDD.n4513 VDD.n4512 0.0096003
R18654 VDD.n4512 VDD.t561 0.0096003
R18655 VDD.n4527 VDD.n4526 0.0096003
R18656 VDD.n4771 VDD.n4770 0.0096003
R18657 VDD.n4770 VDD.t750 0.0096003
R18658 VDD.n4785 VDD.n4784 0.0096003
R18659 VDD.n5046 VDD.n5045 0.0096003
R18660 VDD.n5032 VDD.n5031 0.0096003
R18661 VDD.n5031 VDD.t386 0.0096003
R18662 VDD.n5308 VDD.n5307 0.0096003
R18663 VDD.n5294 VDD.n5293 0.0096003
R18664 VDD.n5293 VDD.t559 0.0096003
R18665 VDD.t420 VDD.n1891 0.00959985
R18666 VDD.n1891 VDD.n1889 0.00959985
R18667 VDD.t148 VDD.n2212 0.00959985
R18668 VDD.n2212 VDD.n2210 0.00959985
R18669 VDD.t676 VDD.n2470 0.00959985
R18670 VDD.n2470 VDD.n2468 0.00959985
R18671 VDD.t689 VDD.n2728 0.00959985
R18672 VDD.n2728 VDD.n2726 0.00959985
R18673 VDD.t93 VDD.n2986 0.00959985
R18674 VDD.n2986 VDD.n2984 0.00959985
R18675 VDD.t76 VDD.n3244 0.00959985
R18676 VDD.n3244 VDD.n3242 0.00959985
R18677 VDD.t1186 VDD.n3502 0.00959985
R18678 VDD.n3502 VDD.n3500 0.00959985
R18679 VDD.t159 VDD.n5829 0.00959985
R18680 VDD.n5829 VDD.n5827 0.00959985
R18681 VDD.t203 VDD.n5575 0.00959985
R18682 VDD.n5575 VDD.n5573 0.00959985
R18683 VDD.t556 VDD.n3760 0.00959985
R18684 VDD.n3760 VDD.n3758 0.00959985
R18685 VDD.t562 VDD.n4018 0.00959985
R18686 VDD.n4018 VDD.n4016 0.00959985
R18687 VDD.t687 VDD.n4276 0.00959985
R18688 VDD.n4276 VDD.n4274 0.00959985
R18689 VDD.t570 VDD.n4534 0.00959985
R18690 VDD.n4534 VDD.n4532 0.00959985
R18691 VDD.t670 VDD.n4792 0.00959985
R18692 VDD.n4792 VDD.n4790 0.00959985
R18693 VDD.t581 VDD.n5053 0.00959985
R18694 VDD.n5053 VDD.n5051 0.00959985
R18695 VDD.t97 VDD.n5315 0.00959985
R18696 VDD.n5315 VDD.n5313 0.00959985
R18697 VDD.n1361 VDD 0.00954255
R18698 VDD.n778 VDD.n775 0.0095362
R18699 VDD.n375 VDD.n372 0.0095362
R18700 VDD.n1425 VDD.n1423 0.0092766
R18701 VDD.n806 VDD.n784 0.00906279
R18702 VDD.n404 VDD.n382 0.00906279
R18703 VDD.n493 VDD.n492 0.00905263
R18704 VDD.n1283 VDD.n1282 0.00883333
R18705 VDD.n1282 VDD.n1280 0.00883333
R18706 VDD.n1280 VDD.n1276 0.00883333
R18707 VDD.n1276 VDD.n1274 0.00883333
R18708 VDD.n1274 VDD.n1270 0.00883333
R18709 VDD.n1295 VDD.n1291 0.00883333
R18710 VDD.n1297 VDD.n1295 0.00883333
R18711 VDD.n1301 VDD.n1297 0.00883333
R18712 VDD.n1303 VDD.n1301 0.00883333
R18713 VDD.n1105 VDD.n1101 0.00878947
R18714 VDD.n1060 VDD.n1058 0.00878947
R18715 VDD.n1002 VDD.n1000 0.00878947
R18716 VDD.n310 VDD.n306 0.00878947
R18717 VDD.n265 VDD.n263 0.00878947
R18718 VDD.n207 VDD.n205 0.00878947
R18719 VDD.n1399 VDD.n1396 0.00874468
R18720 VDD.n894 VDD.n893 0.00852632
R18721 VDD.n907 VDD.n906 0.00852632
R18722 VDD.n952 VDD.n951 0.00852632
R18723 VDD.n99 VDD.n98 0.00852632
R18724 VDD.n112 VDD.n111 0.00852632
R18725 VDD.n157 VDD.n156 0.00852632
R18726 VDD.n2128 VDD.n2127 0.00849839
R18727 VDD.n1287 VDD 0.00847872
R18728 VDD.n1742 VDD.n1741 0.0084202
R18729 VDD.n1699 VDD.n1698 0.0084202
R18730 VDD.n1698 VDD.t1227 0.0084202
R18731 VDD.n1676 VDD.n1672 0.0084202
R18732 VDD.n1764 VDD.n1676 0.0084202
R18733 VDD.n1766 VDD.n1765 0.0084202
R18734 VDD.n1765 VDD.n1764 0.0084202
R18735 VDD.n2091 VDD.n2090 0.0084202
R18736 VDD.n2048 VDD.n2047 0.0084202
R18737 VDD.n2047 VDD.t29 0.0084202
R18738 VDD.n2025 VDD.n2021 0.0084202
R18739 VDD.n2113 VDD.n2025 0.0084202
R18740 VDD.n2115 VDD.n2114 0.0084202
R18741 VDD.n2114 VDD.n2113 0.0084202
R18742 VDD.n2321 VDD.n2320 0.0084202
R18743 VDD.n2278 VDD.n2277 0.0084202
R18744 VDD.n2277 VDD.t541 0.0084202
R18745 VDD.n2255 VDD.n2251 0.0084202
R18746 VDD.n2343 VDD.n2255 0.0084202
R18747 VDD.n2345 VDD.n2344 0.0084202
R18748 VDD.n2344 VDD.n2343 0.0084202
R18749 VDD.n2579 VDD.n2578 0.0084202
R18750 VDD.n2536 VDD.n2535 0.0084202
R18751 VDD.n2535 VDD.t472 0.0084202
R18752 VDD.n2513 VDD.n2509 0.0084202
R18753 VDD.n2601 VDD.n2513 0.0084202
R18754 VDD.n2603 VDD.n2602 0.0084202
R18755 VDD.n2602 VDD.n2601 0.0084202
R18756 VDD.n2837 VDD.n2836 0.0084202
R18757 VDD.n2794 VDD.n2793 0.0084202
R18758 VDD.n2793 VDD.t1309 0.0084202
R18759 VDD.n2771 VDD.n2767 0.0084202
R18760 VDD.n2859 VDD.n2771 0.0084202
R18761 VDD.n2861 VDD.n2860 0.0084202
R18762 VDD.n2860 VDD.n2859 0.0084202
R18763 VDD.n3095 VDD.n3094 0.0084202
R18764 VDD.n3052 VDD.n3051 0.0084202
R18765 VDD.n3051 VDD.t6 0.0084202
R18766 VDD.n3029 VDD.n3025 0.0084202
R18767 VDD.n3117 VDD.n3029 0.0084202
R18768 VDD.n3119 VDD.n3118 0.0084202
R18769 VDD.n3118 VDD.n3117 0.0084202
R18770 VDD.n3353 VDD.n3352 0.0084202
R18771 VDD.n3310 VDD.n3309 0.0084202
R18772 VDD.n3309 VDD.t1194 0.0084202
R18773 VDD.n3287 VDD.n3283 0.0084202
R18774 VDD.n3375 VDD.n3287 0.0084202
R18775 VDD.n3377 VDD.n3376 0.0084202
R18776 VDD.n3376 VDD.n3375 0.0084202
R18777 VDD.n5683 VDD.n5682 0.0084202
R18778 VDD.n5640 VDD.n5639 0.0084202
R18779 VDD.n5639 VDD.t707 0.0084202
R18780 VDD.n5617 VDD.n5613 0.0084202
R18781 VDD.n5705 VDD.n5617 0.0084202
R18782 VDD.n5707 VDD.n5706 0.0084202
R18783 VDD.n5706 VDD.n5705 0.0084202
R18784 VDD.n5429 VDD.n5428 0.0084202
R18785 VDD.n5386 VDD.n5385 0.0084202
R18786 VDD.n5385 VDD.t1331 0.0084202
R18787 VDD.n5363 VDD.n5359 0.0084202
R18788 VDD.n5451 VDD.n5363 0.0084202
R18789 VDD.n5453 VDD.n5452 0.0084202
R18790 VDD.n5452 VDD.n5451 0.0084202
R18791 VDD.n3611 VDD.n3610 0.0084202
R18792 VDD.n3568 VDD.n3567 0.0084202
R18793 VDD.n3567 VDD.t1268 0.0084202
R18794 VDD.n3545 VDD.n3541 0.0084202
R18795 VDD.n3633 VDD.n3545 0.0084202
R18796 VDD.n3635 VDD.n3634 0.0084202
R18797 VDD.n3634 VDD.n3633 0.0084202
R18798 VDD.n3869 VDD.n3868 0.0084202
R18799 VDD.n3826 VDD.n3825 0.0084202
R18800 VDD.n3825 VDD.t81 0.0084202
R18801 VDD.n3803 VDD.n3799 0.0084202
R18802 VDD.n3891 VDD.n3803 0.0084202
R18803 VDD.n3893 VDD.n3892 0.0084202
R18804 VDD.n3892 VDD.n3891 0.0084202
R18805 VDD.n4127 VDD.n4126 0.0084202
R18806 VDD.n4084 VDD.n4083 0.0084202
R18807 VDD.n4083 VDD.t723 0.0084202
R18808 VDD.n4061 VDD.n4057 0.0084202
R18809 VDD.n4149 VDD.n4061 0.0084202
R18810 VDD.n4151 VDD.n4150 0.0084202
R18811 VDD.n4150 VDD.n4149 0.0084202
R18812 VDD.n4385 VDD.n4384 0.0084202
R18813 VDD.n4342 VDD.n4341 0.0084202
R18814 VDD.n4341 VDD.t1112 0.0084202
R18815 VDD.n4319 VDD.n4315 0.0084202
R18816 VDD.n4407 VDD.n4319 0.0084202
R18817 VDD.n4409 VDD.n4408 0.0084202
R18818 VDD.n4408 VDD.n4407 0.0084202
R18819 VDD.n4643 VDD.n4642 0.0084202
R18820 VDD.n4600 VDD.n4599 0.0084202
R18821 VDD.n4599 VDD.t183 0.0084202
R18822 VDD.n4577 VDD.n4573 0.0084202
R18823 VDD.n4665 VDD.n4577 0.0084202
R18824 VDD.n4667 VDD.n4666 0.0084202
R18825 VDD.n4666 VDD.n4665 0.0084202
R18826 VDD.n4901 VDD.n4900 0.0084202
R18827 VDD.n4858 VDD.n4857 0.0084202
R18828 VDD.n4857 VDD.t1121 0.0084202
R18829 VDD.n4835 VDD.n4831 0.0084202
R18830 VDD.n4923 VDD.n4835 0.0084202
R18831 VDD.n4925 VDD.n4924 0.0084202
R18832 VDD.n4924 VDD.n4923 0.0084202
R18833 VDD.n5193 VDD.n5192 0.0084202
R18834 VDD.n5150 VDD.n5149 0.0084202
R18835 VDD.n5149 VDD.t195 0.0084202
R18836 VDD.n5127 VDD.n5123 0.0084202
R18837 VDD.n5215 VDD.n5127 0.0084202
R18838 VDD.n5217 VDD.n5216 0.0084202
R18839 VDD.n5216 VDD.n5215 0.0084202
R18840 VDD.n1615 VDD.n1614 0.0083125
R18841 VDD.n700 VDD.n696 0.00826316
R18842 VDD.n655 VDD.n653 0.00826316
R18843 VDD.n597 VDD.n595 0.00826316
R18844 VDD.n1366 VDD.n1365 0.00821277
R18845 VDD.n5227 VDD.n5226 0.00811918
R18846 VDD.n713 VDD.n712 0.00802802
R18847 VDD.n1554 VDD.n1553 0.00802802
R18848 VDD.n506 VDD.n505 0.008
R18849 VDD.n551 VDD.n550 0.008
R18850 VDD.n577 VDD.n576 0.008
R18851 VDD.n741 VDD.n738 0.00775202
R18852 VDD.n720 VDD.n717 0.00775202
R18853 VDD.n1582 VDD.n1579 0.00775202
R18854 VDD.n1561 VDD.n1558 0.00775202
R18855 VDD.n693 VDD.n692 0.00773684
R18856 VDD.n648 VDD.n647 0.00773684
R18857 VDD.n899 VDD.n857 0.00747368
R18858 VDD.n982 VDD.n981 0.00747368
R18859 VDD.n104 VDD.n62 0.00747368
R18860 VDD.n187 VDD.n186 0.00747368
R18861 VDD VDD.n1320 0.00741489
R18862 VDD.n1098 VDD.n1097 0.00721053
R18863 VDD.n1053 VDD.n1052 0.00721053
R18864 VDD.n303 VDD.n302 0.00721053
R18865 VDD.n258 VDD.n257 0.00721053
R18866 VDD.n1543 VDD 0.00714063
R18867 VDD.n1743 VDD.n1742 0.00702894
R18868 VDD.n2092 VDD.n2091 0.00702894
R18869 VDD.n2322 VDD.n2321 0.00702894
R18870 VDD.n2580 VDD.n2579 0.00702894
R18871 VDD.n2838 VDD.n2837 0.00702894
R18872 VDD.n3096 VDD.n3095 0.00702894
R18873 VDD.n3354 VDD.n3353 0.00702894
R18874 VDD.n5684 VDD.n5683 0.00702894
R18875 VDD.n5430 VDD.n5429 0.00702894
R18876 VDD.n3612 VDD.n3611 0.00702894
R18877 VDD.n3870 VDD.n3869 0.00702894
R18878 VDD.n4128 VDD.n4127 0.00702894
R18879 VDD.n4386 VDD.n4385 0.00702894
R18880 VDD.n4644 VDD.n4643 0.00702894
R18881 VDD.n4902 VDD.n4901 0.00702894
R18882 VDD.n5194 VDD.n5193 0.00702894
R18883 VDD.n1291 VDD.n1246 0.00702174
R18884 VDD.n1133 VDD 0.00700289
R18885 VDD.n1199 VDD 0.00700289
R18886 VDD.n498 VDD.n456 0.00694737
R18887 VDD.n1829 VDD.n1828 0.00693382
R18888 VDD.n2150 VDD.n2149 0.00693382
R18889 VDD.n2408 VDD.n2407 0.00693382
R18890 VDD.n2666 VDD.n2665 0.00693382
R18891 VDD.n2924 VDD.n2923 0.00693382
R18892 VDD.n3182 VDD.n3181 0.00693382
R18893 VDD.n3440 VDD.n3439 0.00693382
R18894 VDD.n5767 VDD.n5766 0.00693382
R18895 VDD.n5513 VDD.n5512 0.00693382
R18896 VDD.n3698 VDD.n3697 0.00693382
R18897 VDD.n3956 VDD.n3955 0.00693382
R18898 VDD.n4214 VDD.n4213 0.00693382
R18899 VDD.n4472 VDD.n4471 0.00693382
R18900 VDD.n4730 VDD.n4729 0.00693382
R18901 VDD.n4991 VDD.n4990 0.00693382
R18902 VDD.n5253 VDD.n5252 0.00693382
R18903 VDD.n1126 VDD 0.00675
R18904 VDD.n1192 VDD 0.00675
R18905 VDD.n1540 VDD.n1255 0.00662745
R18906 VDD.n1463 VDD.n1461 0.00661702
R18907 VDD VDD.n868 0.00655263
R18908 VDD.n939 VDD 0.00655263
R18909 VDD VDD.n1108 0.00655263
R18910 VDD VDD.n1061 0.00655263
R18911 VDD VDD.n1014 0.00655263
R18912 VDD.n994 VDD 0.00655263
R18913 VDD VDD.n73 0.00655263
R18914 VDD.n144 VDD 0.00655263
R18915 VDD VDD.n313 0.00655263
R18916 VDD VDD.n266 0.00655263
R18917 VDD VDD.n219 0.00655263
R18918 VDD.n199 VDD 0.00655263
R18919 VDD VDD.n467 0.00655263
R18920 VDD.n538 VDD 0.00655263
R18921 VDD VDD.n703 0.00655263
R18922 VDD VDD.n656 0.00655263
R18923 VDD VDD.n609 0.00655263
R18924 VDD.n589 VDD 0.00655263
R18925 VDD.n1111 VDD.n35 0.00638056
R18926 VDD.n498 VDD.n497 0.00615789
R18927 VDD VDD.n1125 0.00609211
R18928 VDD VDD.n1191 0.00609211
R18929 VDD.n1739 VDD.n1736 0.00605556
R18930 VDD.n2088 VDD.n2085 0.00605556
R18931 VDD.n2318 VDD.n2315 0.00605556
R18932 VDD.n2576 VDD.n2573 0.00605556
R18933 VDD.n2834 VDD.n2831 0.00605556
R18934 VDD.n3092 VDD.n3089 0.00605556
R18935 VDD.n3350 VDD.n3347 0.00605556
R18936 VDD.n5680 VDD.n5677 0.00605556
R18937 VDD.n5426 VDD.n5423 0.00605556
R18938 VDD.n3608 VDD.n3605 0.00605556
R18939 VDD.n3866 VDD.n3863 0.00605556
R18940 VDD.n4124 VDD.n4121 0.00605556
R18941 VDD.n4382 VDD.n4379 0.00605556
R18942 VDD.n4640 VDD.n4637 0.00605556
R18943 VDD.n4898 VDD.n4895 0.00605556
R18944 VDD.n5190 VDD.n5187 0.00605556
R18945 VDD.n4935 VDD.n4934 0.00602323
R18946 VDD.n1100 VDD.n1098 0.00589474
R18947 VDD.n1057 VDD.n1053 0.00589474
R18948 VDD.n305 VDD.n303 0.00589474
R18949 VDD.n262 VDD.n258 0.00589474
R18950 VDD.n1343 VDD.n1320 0.00581915
R18951 VDD.n1982 VDD.n1981 0.00573228
R18952 VDD.n1982 VDD.n1980 0.00573228
R18953 VDD.n1540 VDD.n1539 0.00564706
R18954 VDD.n899 VDD.n898 0.00563158
R18955 VDD.n982 VDD.n954 0.00563158
R18956 VDD.n1003 VDD 0.00563158
R18957 VDD.n104 VDD.n103 0.00563158
R18958 VDD.n187 VDD.n159 0.00563158
R18959 VDD.n208 VDD 0.00563158
R18960 VDD.n1376 VDD.n1374 0.00552129
R18961 VDD.n1603 VDD.n1602 0.00542857
R18962 VDD.n695 VDD.n693 0.00536842
R18963 VDD.n652 VDD.n648 0.00536842
R18964 VDD.n1617 VDD.n1615 0.0051875
R18965 VDD.n510 VDD.n506 0.00510526
R18966 VDD.n553 VDD.n551 0.00510526
R18967 VDD.n577 VDD.n553 0.00510526
R18968 VDD.n598 VDD 0.00510526
R18969 VDD.n1913 VDD.n1912 0.00505015
R18970 VDD.t420 VDD.n1913 0.00505015
R18971 VDD.t420 VDD.n1894 0.00505015
R18972 VDD.n1909 VDD.n1894 0.00505015
R18973 VDD.n1824 VDD.n1823 0.00505015
R18974 VDD.n1861 VDD.n1848 0.00505015
R18975 VDD.t355 VDD.n1848 0.00505015
R18976 VDD.n1868 VDD.n1867 0.00505015
R18977 VDD.t355 VDD.n1868 0.00505015
R18978 VDD.n2182 VDD.n2169 0.00505015
R18979 VDD.t574 VDD.n2169 0.00505015
R18980 VDD.n2189 VDD.n2188 0.00505015
R18981 VDD.t574 VDD.n2189 0.00505015
R18982 VDD.n2145 VDD.n2144 0.00505015
R18983 VDD.n2234 VDD.n2233 0.00505015
R18984 VDD.t148 VDD.n2234 0.00505015
R18985 VDD.t148 VDD.n2215 0.00505015
R18986 VDD.n2230 VDD.n2215 0.00505015
R18987 VDD.n2440 VDD.n2427 0.00505015
R18988 VDD.t103 VDD.n2427 0.00505015
R18989 VDD.n2447 VDD.n2446 0.00505015
R18990 VDD.t103 VDD.n2447 0.00505015
R18991 VDD.n2403 VDD.n2402 0.00505015
R18992 VDD.n2492 VDD.n2491 0.00505015
R18993 VDD.t676 VDD.n2492 0.00505015
R18994 VDD.t676 VDD.n2473 0.00505015
R18995 VDD.n2488 VDD.n2473 0.00505015
R18996 VDD.n2698 VDD.n2685 0.00505015
R18997 VDD.t421 VDD.n2685 0.00505015
R18998 VDD.n2705 VDD.n2704 0.00505015
R18999 VDD.t421 VDD.n2705 0.00505015
R19000 VDD.n2661 VDD.n2660 0.00505015
R19001 VDD.n2750 VDD.n2749 0.00505015
R19002 VDD.t689 VDD.n2750 0.00505015
R19003 VDD.t689 VDD.n2731 0.00505015
R19004 VDD.n2746 VDD.n2731 0.00505015
R19005 VDD.n2956 VDD.n2943 0.00505015
R19006 VDD.t405 VDD.n2943 0.00505015
R19007 VDD.n2963 VDD.n2962 0.00505015
R19008 VDD.t405 VDD.n2963 0.00505015
R19009 VDD.n2919 VDD.n2918 0.00505015
R19010 VDD.n3008 VDD.n3007 0.00505015
R19011 VDD.t93 VDD.n3008 0.00505015
R19012 VDD.t93 VDD.n2989 0.00505015
R19013 VDD.n3004 VDD.n2989 0.00505015
R19014 VDD.n3214 VDD.n3201 0.00505015
R19015 VDD.t144 VDD.n3201 0.00505015
R19016 VDD.n3221 VDD.n3220 0.00505015
R19017 VDD.t144 VDD.n3221 0.00505015
R19018 VDD.n3177 VDD.n3176 0.00505015
R19019 VDD.n3266 VDD.n3265 0.00505015
R19020 VDD.t76 VDD.n3266 0.00505015
R19021 VDD.t76 VDD.n3247 0.00505015
R19022 VDD.n3262 VDD.n3247 0.00505015
R19023 VDD.n3472 VDD.n3459 0.00505015
R19024 VDD.t179 VDD.n3459 0.00505015
R19025 VDD.n3479 VDD.n3478 0.00505015
R19026 VDD.t179 VDD.n3479 0.00505015
R19027 VDD.n3435 VDD.n3434 0.00505015
R19028 VDD.n3524 VDD.n3523 0.00505015
R19029 VDD.t1186 VDD.n3524 0.00505015
R19030 VDD.t1186 VDD.n3505 0.00505015
R19031 VDD.n3520 VDD.n3505 0.00505015
R19032 VDD.n5799 VDD.n5786 0.00505015
R19033 VDD.t1088 VDD.n5786 0.00505015
R19034 VDD.n5806 VDD.n5805 0.00505015
R19035 VDD.t1088 VDD.n5806 0.00505015
R19036 VDD.n5762 VDD.n5761 0.00505015
R19037 VDD.n5851 VDD.n5850 0.00505015
R19038 VDD.t159 VDD.n5851 0.00505015
R19039 VDD.t159 VDD.n5832 0.00505015
R19040 VDD.n5847 VDD.n5832 0.00505015
R19041 VDD.n5545 VDD.n5532 0.00505015
R19042 VDD.t596 VDD.n5532 0.00505015
R19043 VDD.n5552 VDD.n5551 0.00505015
R19044 VDD.t596 VDD.n5552 0.00505015
R19045 VDD.n5508 VDD.n5507 0.00505015
R19046 VDD.n5597 VDD.n5596 0.00505015
R19047 VDD.t203 VDD.n5597 0.00505015
R19048 VDD.t203 VDD.n5578 0.00505015
R19049 VDD.n5593 VDD.n5578 0.00505015
R19050 VDD.n3730 VDD.n3717 0.00505015
R19051 VDD.t145 VDD.n3717 0.00505015
R19052 VDD.n3737 VDD.n3736 0.00505015
R19053 VDD.t145 VDD.n3737 0.00505015
R19054 VDD.n3693 VDD.n3692 0.00505015
R19055 VDD.n3782 VDD.n3781 0.00505015
R19056 VDD.t556 VDD.n3782 0.00505015
R19057 VDD.t556 VDD.n3763 0.00505015
R19058 VDD.n3778 VDD.n3763 0.00505015
R19059 VDD.n3988 VDD.n3975 0.00505015
R19060 VDD.t563 VDD.n3975 0.00505015
R19061 VDD.n3995 VDD.n3994 0.00505015
R19062 VDD.t563 VDD.n3995 0.00505015
R19063 VDD.n3951 VDD.n3950 0.00505015
R19064 VDD.n4040 VDD.n4039 0.00505015
R19065 VDD.t562 VDD.n4040 0.00505015
R19066 VDD.t562 VDD.n4021 0.00505015
R19067 VDD.n4036 VDD.n4021 0.00505015
R19068 VDD.n4246 VDD.n4233 0.00505015
R19069 VDD.t668 VDD.n4233 0.00505015
R19070 VDD.n4253 VDD.n4252 0.00505015
R19071 VDD.t668 VDD.n4253 0.00505015
R19072 VDD.n4209 VDD.n4208 0.00505015
R19073 VDD.n4298 VDD.n4297 0.00505015
R19074 VDD.t687 VDD.n4298 0.00505015
R19075 VDD.t687 VDD.n4279 0.00505015
R19076 VDD.n4294 VDD.n4279 0.00505015
R19077 VDD.n4504 VDD.n4491 0.00505015
R19078 VDD.t561 VDD.n4491 0.00505015
R19079 VDD.n4511 VDD.n4510 0.00505015
R19080 VDD.t561 VDD.n4511 0.00505015
R19081 VDD.n4467 VDD.n4466 0.00505015
R19082 VDD.n4556 VDD.n4555 0.00505015
R19083 VDD.t570 VDD.n4556 0.00505015
R19084 VDD.t570 VDD.n4537 0.00505015
R19085 VDD.n4552 VDD.n4537 0.00505015
R19086 VDD.n4762 VDD.n4749 0.00505015
R19087 VDD.t750 VDD.n4749 0.00505015
R19088 VDD.n4769 VDD.n4768 0.00505015
R19089 VDD.t750 VDD.n4769 0.00505015
R19090 VDD.n4725 VDD.n4724 0.00505015
R19091 VDD.n4814 VDD.n4813 0.00505015
R19092 VDD.t670 VDD.n4814 0.00505015
R19093 VDD.t670 VDD.n4795 0.00505015
R19094 VDD.n4810 VDD.n4795 0.00505015
R19095 VDD.n5075 VDD.n5074 0.00505015
R19096 VDD.t581 VDD.n5075 0.00505015
R19097 VDD.t581 VDD.n5056 0.00505015
R19098 VDD.n5071 VDD.n5056 0.00505015
R19099 VDD.n4986 VDD.n4985 0.00505015
R19100 VDD.n5023 VDD.n5010 0.00505015
R19101 VDD.t386 VDD.n5010 0.00505015
R19102 VDD.n5030 VDD.n5029 0.00505015
R19103 VDD.t386 VDD.n5030 0.00505015
R19104 VDD.n5337 VDD.n5336 0.00505015
R19105 VDD.t97 VDD.n5337 0.00505015
R19106 VDD.t97 VDD.n5318 0.00505015
R19107 VDD.n5333 VDD.n5318 0.00505015
R19108 VDD.n5248 VDD.n5247 0.00505015
R19109 VDD.n5285 VDD.n5272 0.00505015
R19110 VDD.t559 VDD.n5272 0.00505015
R19111 VDD.n5292 VDD.n5291 0.00505015
R19112 VDD.t559 VDD.n5292 0.00505015
R19113 VDD.n1311 VDD 0.00502128
R19114 VDD.n1340 VDD 0.00502128
R19115 VDD VDD.n1346 0.00502128
R19116 VDD.n1363 VDD 0.00502128
R19117 VDD.n1510 VDD 0.00502128
R19118 VDD.n696 VDD.n695 0.00484211
R19119 VDD.n653 VDD.n652 0.00484211
R19120 VDD.n595 VDD.n594 0.00484211
R19121 VDD.n1324 VDD.n1319 0.00475532
R19122 VDD VDD.n1509 0.00475532
R19123 VDD.n1504 VDD.n1261 0.00475532
R19124 VDD.n1287 VDD.n1286 0.00475532
R19125 VDD.n1751 VDD.n1722 0.00466667
R19126 VDD.n1703 VDD.n1702 0.00466667
R19127 VDD.n1692 VDD.n1691 0.00466667
R19128 VDD.n2100 VDD.n2071 0.00466667
R19129 VDD.n2052 VDD.n2051 0.00466667
R19130 VDD.n2041 VDD.n2040 0.00466667
R19131 VDD.n2330 VDD.n2301 0.00466667
R19132 VDD.n2282 VDD.n2281 0.00466667
R19133 VDD.n2271 VDD.n2270 0.00466667
R19134 VDD.n2588 VDD.n2559 0.00466667
R19135 VDD.n2540 VDD.n2539 0.00466667
R19136 VDD.n2529 VDD.n2528 0.00466667
R19137 VDD.n2846 VDD.n2817 0.00466667
R19138 VDD.n2798 VDD.n2797 0.00466667
R19139 VDD.n2787 VDD.n2786 0.00466667
R19140 VDD.n3104 VDD.n3075 0.00466667
R19141 VDD.n3056 VDD.n3055 0.00466667
R19142 VDD.n3045 VDD.n3044 0.00466667
R19143 VDD.n3362 VDD.n3333 0.00466667
R19144 VDD.n3314 VDD.n3313 0.00466667
R19145 VDD.n3303 VDD.n3302 0.00466667
R19146 VDD.n5692 VDD.n5663 0.00466667
R19147 VDD.n5644 VDD.n5643 0.00466667
R19148 VDD.n5633 VDD.n5632 0.00466667
R19149 VDD.n5438 VDD.n5409 0.00466667
R19150 VDD.n5390 VDD.n5389 0.00466667
R19151 VDD.n5379 VDD.n5378 0.00466667
R19152 VDD.n3620 VDD.n3591 0.00466667
R19153 VDD.n3572 VDD.n3571 0.00466667
R19154 VDD.n3561 VDD.n3560 0.00466667
R19155 VDD.n3878 VDD.n3849 0.00466667
R19156 VDD.n3830 VDD.n3829 0.00466667
R19157 VDD.n3819 VDD.n3818 0.00466667
R19158 VDD.n4136 VDD.n4107 0.00466667
R19159 VDD.n4088 VDD.n4087 0.00466667
R19160 VDD.n4077 VDD.n4076 0.00466667
R19161 VDD.n4394 VDD.n4365 0.00466667
R19162 VDD.n4346 VDD.n4345 0.00466667
R19163 VDD.n4335 VDD.n4334 0.00466667
R19164 VDD.n4652 VDD.n4623 0.00466667
R19165 VDD.n4604 VDD.n4603 0.00466667
R19166 VDD.n4593 VDD.n4592 0.00466667
R19167 VDD.n4910 VDD.n4881 0.00466667
R19168 VDD.n4862 VDD.n4861 0.00466667
R19169 VDD.n4851 VDD.n4850 0.00466667
R19170 VDD.n5202 VDD.n5173 0.00466667
R19171 VDD.n5154 VDD.n5153 0.00466667
R19172 VDD.n5143 VDD.n5142 0.00466667
R19173 VDD VDD.n35 0.00460833
R19174 VDD.n898 VDD.n894 0.00457895
R19175 VDD.n911 VDD.n907 0.00457895
R19176 VDD.n954 VDD.n952 0.00457895
R19177 VDD.n103 VDD.n99 0.00457895
R19178 VDD.n116 VDD.n112 0.00457895
R19179 VDD.n159 VDD.n157 0.00457895
R19180 VDD.n1547 VDD.n1546 0.00451563
R19181 VDD.n1101 VDD.n1100 0.00431579
R19182 VDD.n1058 VDD.n1057 0.00431579
R19183 VDD.n1000 VDD.n999 0.00431579
R19184 VDD.n306 VDD.n305 0.00431579
R19185 VDD.n263 VDD.n262 0.00431579
R19186 VDD.n205 VDD.n204 0.00431579
R19187 VDD.n1406 VDD.n1405 0.0042234
R19188 VDD.n1304 VDD.n1303 0.00412319
R19189 VDD VDD.n1126 0.00411272
R19190 VDD VDD.n1192 0.00411272
R19191 VDD.n1611 VDD.n1610 0.00410577
R19192 VDD.n497 VDD.n493 0.00405263
R19193 VDD.n829 VDD 0.00400806
R19194 VDD.n2125 VDD.n2013 0.00390318
R19195 VDD.n1126 VDD 0.00378947
R19196 VDD.n1192 VDD 0.00378947
R19197 VDD.n1526 VDD.n1525 0.00369149
R19198 VDD.n1816 VDD.n1809 0.00364862
R19199 VDD.n2137 VDD.n2130 0.00364862
R19200 VDD.n2395 VDD.n2388 0.00364862
R19201 VDD.n2653 VDD.n2646 0.00364862
R19202 VDD.n2911 VDD.n2904 0.00364862
R19203 VDD.n3169 VDD.n3162 0.00364862
R19204 VDD.n3427 VDD.n3420 0.00364862
R19205 VDD.n5754 VDD.n5747 0.00364862
R19206 VDD.n5500 VDD.n5493 0.00364862
R19207 VDD.n3685 VDD.n3678 0.00364862
R19208 VDD.n3943 VDD.n3936 0.00364862
R19209 VDD.n4201 VDD.n4194 0.00364862
R19210 VDD.n4459 VDD.n4452 0.00364862
R19211 VDD.n4717 VDD.n4710 0.00364862
R19212 VDD.n4978 VDD.n4971 0.00364862
R19213 VDD.n5240 VDD.n5233 0.00364862
R19214 VDD.n1289 VDD 0.00342553
R19215 VDD.n1609 VDD.n1604 0.00339649
R19216 VDD VDD.n1113 0.00330645
R19217 VDD.n456 VDD.n454 0.00326316
R19218 VDD.n1934 VDD.n1926 0.00317113
R19219 VDD.n1955 VDD.n1944 0.00317113
R19220 VDD.n1359 VDD.n1358 0.00315957
R19221 VDD.n1600 VDD 0.00304286
R19222 VDD.n1097 VDD.n1093 0.003
R19223 VDD.n1052 VDD.n1050 0.003
R19224 VDD.n302 VDD.n298 0.003
R19225 VDD.n257 VDD.n255 0.003
R19226 VDD.n1743 VDD.t37 0.00289124
R19227 VDD.n2092 VDD.t365 0.00289124
R19228 VDD.n2322 VDD.t466 0.00289124
R19229 VDD.n2580 VDD.t117 0.00289124
R19230 VDD.n2838 VDD.t21 0.00289124
R19231 VDD.n3096 VDD.t590 0.00289124
R19232 VDD.n3354 VDD.t550 0.00289124
R19233 VDD.n5684 VDD.t170 0.00289124
R19234 VDD.n5430 VDD.t757 0.00289124
R19235 VDD.n3612 VDD.t1100 0.00289124
R19236 VDD.n3870 VDD.t785 0.00289124
R19237 VDD.n4128 VDD.t490 0.00289124
R19238 VDD.n4386 VDD.t374 0.00289124
R19239 VDD.n4644 VDD.t111 0.00289124
R19240 VDD.n4902 VDD.t349 0.00289124
R19241 VDD.n5194 VDD.t482 0.00289124
R19242 VDD.n857 VDD.n855 0.00273684
R19243 VDD.n869 VDD 0.00273684
R19244 VDD.n936 VDD 0.00273684
R19245 VDD.n981 VDD.n977 0.00273684
R19246 VDD.n1109 VDD 0.00273684
R19247 VDD.n1062 VDD 0.00273684
R19248 VDD.n1015 VDD 0.00273684
R19249 VDD.n997 VDD 0.00273684
R19250 VDD.n62 VDD.n60 0.00273684
R19251 VDD.n74 VDD 0.00273684
R19252 VDD.n141 VDD 0.00273684
R19253 VDD.n186 VDD.n182 0.00273684
R19254 VDD.n314 VDD 0.00273684
R19255 VDD.n267 VDD 0.00273684
R19256 VDD.n220 VDD 0.00273684
R19257 VDD.n202 VDD 0.00273684
R19258 VDD.n468 VDD 0.00273684
R19259 VDD.n535 VDD 0.00273684
R19260 VDD.n704 VDD 0.00273684
R19261 VDD.n657 VDD 0.00273684
R19262 VDD.n610 VDD 0.00273684
R19263 VDD.n592 VDD 0.00273684
R19264 VDD.n505 VDD.n503 0.00271053
R19265 VDD.n1926 VDD.n1925 0.00267116
R19266 VDD.n1956 VDD.n1955 0.00267116
R19267 VDD.n4934 VDD.n4933 0.0026624
R19268 VDD.n1506 VDD 0.00262766
R19269 VDD.n1006 VDD.n1005 0.00247368
R19270 VDD.n211 VDD.n210 0.00247368
R19271 VDD.n692 VDD.n688 0.00247368
R19272 VDD.n647 VDD.n645 0.00247368
R19273 VDD.n1838 VDD.n1837 0.00240766
R19274 VDD.n2159 VDD.n2158 0.00240766
R19275 VDD.n2417 VDD.n2416 0.00240766
R19276 VDD.n2675 VDD.n2674 0.00240766
R19277 VDD.n2933 VDD.n2932 0.00240766
R19278 VDD.n3191 VDD.n3190 0.00240766
R19279 VDD.n3449 VDD.n3448 0.00240766
R19280 VDD.n5776 VDD.n5775 0.00240766
R19281 VDD.n5522 VDD.n5521 0.00240766
R19282 VDD.n3707 VDD.n3706 0.00240766
R19283 VDD.n3965 VDD.n3964 0.00240766
R19284 VDD.n4223 VDD.n4222 0.00240766
R19285 VDD.n4481 VDD.n4480 0.00240766
R19286 VDD.n4739 VDD.n4738 0.00240766
R19287 VDD.n5000 VDD.n4999 0.00240766
R19288 VDD.n5262 VDD.n5261 0.00240766
R19289 VDD.n1601 VDD.n1600 0.00237143
R19290 VDD.n1359 VDD 0.0023617
R19291 VDD.n1369 VDD.n1368 0.0023617
R19292 VDD.n1829 VDD.n1825 0.00233824
R19293 VDD.n1831 VDD 0.00233824
R19294 VDD.n2150 VDD.n2146 0.00233824
R19295 VDD.n2152 VDD 0.00233824
R19296 VDD.n2408 VDD.n2404 0.00233824
R19297 VDD.n2410 VDD 0.00233824
R19298 VDD.n2666 VDD.n2662 0.00233824
R19299 VDD.n2668 VDD 0.00233824
R19300 VDD.n2924 VDD.n2920 0.00233824
R19301 VDD.n2926 VDD 0.00233824
R19302 VDD.n3182 VDD.n3178 0.00233824
R19303 VDD.n3184 VDD 0.00233824
R19304 VDD.n3440 VDD.n3436 0.00233824
R19305 VDD.n3442 VDD 0.00233824
R19306 VDD.n5767 VDD.n5763 0.00233824
R19307 VDD.n5769 VDD 0.00233824
R19308 VDD.n5513 VDD.n5509 0.00233824
R19309 VDD.n5515 VDD 0.00233824
R19310 VDD.n3698 VDD.n3694 0.00233824
R19311 VDD.n3700 VDD 0.00233824
R19312 VDD.n3956 VDD.n3952 0.00233824
R19313 VDD.n3958 VDD 0.00233824
R19314 VDD.n4214 VDD.n4210 0.00233824
R19315 VDD.n4216 VDD 0.00233824
R19316 VDD.n4472 VDD.n4468 0.00233824
R19317 VDD.n4474 VDD 0.00233824
R19318 VDD.n4730 VDD.n4726 0.00233824
R19319 VDD.n4732 VDD 0.00233824
R19320 VDD.n4991 VDD.n4987 0.00233824
R19321 VDD.n4993 VDD 0.00233824
R19322 VDD.n5253 VDD.n5249 0.00233824
R19323 VDD.n5255 VDD 0.00233824
R19324 VDD.n1454 VDD.n1317 0.00232979
R19325 VDD.n1431 VDD.n1319 0.00232979
R19326 VDD.n1879 VDD.t417 0.00231811
R19327 VDD.n2200 VDD.t1085 0.00231811
R19328 VDD.n2458 VDD.t567 0.00231811
R19329 VDD.n2716 VDD.t387 0.00231811
R19330 VDD.n2974 VDD.t560 0.00231811
R19331 VDD.n3232 VDD.t573 0.00231811
R19332 VDD.n3490 VDD.t143 0.00231811
R19333 VDD.n5817 VDD.t419 0.00231811
R19334 VDD.n5563 VDD.t667 0.00231811
R19335 VDD.n3748 VDD.t142 0.00231811
R19336 VDD.n4006 VDD.t782 0.00231811
R19337 VDD.n4264 VDD.t1087 0.00231811
R19338 VDD.n4522 VDD.t558 0.00231811
R19339 VDD.n4780 VDD.t572 0.00231811
R19340 VDD.n5041 VDD.t690 0.00231811
R19341 VDD.n5303 VDD.t418 0.00231811
R19342 VDD.n1270 VDD.n1246 0.00231159
R19343 VDD.n1726 VDD.n1724 0.00228571
R19344 VDD.n2075 VDD.n2073 0.00228571
R19345 VDD.n2305 VDD.n2303 0.00228571
R19346 VDD.n2563 VDD.n2561 0.00228571
R19347 VDD.n2821 VDD.n2819 0.00228571
R19348 VDD.n3079 VDD.n3077 0.00228571
R19349 VDD.n3337 VDD.n3335 0.00228571
R19350 VDD.n5667 VDD.n5665 0.00228571
R19351 VDD.n5413 VDD.n5411 0.00228571
R19352 VDD.n3595 VDD.n3593 0.00228571
R19353 VDD.n3853 VDD.n3851 0.00228571
R19354 VDD.n4111 VDD.n4109 0.00228571
R19355 VDD.n4369 VDD.n4367 0.00228571
R19356 VDD.n4627 VDD.n4625 0.00228571
R19357 VDD.n4885 VDD.n4883 0.00228571
R19358 VDD.n5177 VDD.n5175 0.00228571
R19359 VDD.n1694 VDD.n1693 0.00221302
R19360 VDD.n1695 VDD.n1694 0.00221302
R19361 VDD.n2043 VDD.n2042 0.00221302
R19362 VDD.n2044 VDD.n2043 0.00221302
R19363 VDD.n2273 VDD.n2272 0.00221302
R19364 VDD.n2274 VDD.n2273 0.00221302
R19365 VDD.n2531 VDD.n2530 0.00221302
R19366 VDD.n2532 VDD.n2531 0.00221302
R19367 VDD.n2789 VDD.n2788 0.00221302
R19368 VDD.n2790 VDD.n2789 0.00221302
R19369 VDD.n3047 VDD.n3046 0.00221302
R19370 VDD.n3048 VDD.n3047 0.00221302
R19371 VDD.n3305 VDD.n3304 0.00221302
R19372 VDD.n3306 VDD.n3305 0.00221302
R19373 VDD.n5635 VDD.n5634 0.00221302
R19374 VDD.n5636 VDD.n5635 0.00221302
R19375 VDD.n5381 VDD.n5380 0.00221302
R19376 VDD.n5382 VDD.n5381 0.00221302
R19377 VDD.n3563 VDD.n3562 0.00221302
R19378 VDD.n3564 VDD.n3563 0.00221302
R19379 VDD.n3821 VDD.n3820 0.00221302
R19380 VDD.n3822 VDD.n3821 0.00221302
R19381 VDD.n4079 VDD.n4078 0.00221302
R19382 VDD.n4080 VDD.n4079 0.00221302
R19383 VDD.n4337 VDD.n4336 0.00221302
R19384 VDD.n4338 VDD.n4337 0.00221302
R19385 VDD.n4595 VDD.n4594 0.00221302
R19386 VDD.n4596 VDD.n4595 0.00221302
R19387 VDD.n4853 VDD.n4852 0.00221302
R19388 VDD.n4854 VDD.n4853 0.00221302
R19389 VDD.n5145 VDD.n5144 0.00221302
R19390 VDD.n5146 VDD.n5145 0.00221302
R19391 VDD.n1693 VDD.n1692 0.00221271
R19392 VDD.n2042 VDD.n2041 0.00221271
R19393 VDD.n2272 VDD.n2271 0.00221271
R19394 VDD.n2530 VDD.n2529 0.00221271
R19395 VDD.n2788 VDD.n2787 0.00221271
R19396 VDD.n3046 VDD.n3045 0.00221271
R19397 VDD.n3304 VDD.n3303 0.00221271
R19398 VDD.n5634 VDD.n5633 0.00221271
R19399 VDD.n5380 VDD.n5379 0.00221271
R19400 VDD.n3562 VDD.n3561 0.00221271
R19401 VDD.n3820 VDD.n3819 0.00221271
R19402 VDD.n4078 VDD.n4077 0.00221271
R19403 VDD.n4336 VDD.n4335 0.00221271
R19404 VDD.n4594 VDD.n4593 0.00221271
R19405 VDD.n4852 VDD.n4851 0.00221271
R19406 VDD.n5144 VDD.n5143 0.00221271
R19407 VDD.n576 VDD.n572 0.00221053
R19408 VDD.n1732 VDD.n1730 0.00220611
R19409 VDD.n2081 VDD.n2079 0.00220611
R19410 VDD.n2311 VDD.n2309 0.00220611
R19411 VDD.n2569 VDD.n2567 0.00220611
R19412 VDD.n2827 VDD.n2825 0.00220611
R19413 VDD.n3085 VDD.n3083 0.00220611
R19414 VDD.n3343 VDD.n3341 0.00220611
R19415 VDD.n5673 VDD.n5671 0.00220611
R19416 VDD.n5419 VDD.n5417 0.00220611
R19417 VDD.n3601 VDD.n3599 0.00220611
R19418 VDD.n3859 VDD.n3857 0.00220611
R19419 VDD.n4117 VDD.n4115 0.00220611
R19420 VDD.n4375 VDD.n4373 0.00220611
R19421 VDD.n4633 VDD.n4631 0.00220611
R19422 VDD.n4891 VDD.n4889 0.00220611
R19423 VDD.n5183 VDD.n5181 0.00220611
R19424 VDD.n1702 VDD.n1681 0.0022058
R19425 VDD.n2051 VDD.n2030 0.0022058
R19426 VDD.n2281 VDD.n2260 0.0022058
R19427 VDD.n2539 VDD.n2518 0.0022058
R19428 VDD.n2797 VDD.n2776 0.0022058
R19429 VDD.n3055 VDD.n3034 0.0022058
R19430 VDD.n3313 VDD.n3292 0.0022058
R19431 VDD.n5643 VDD.n5622 0.0022058
R19432 VDD.n5389 VDD.n5368 0.0022058
R19433 VDD.n3571 VDD.n3550 0.0022058
R19434 VDD.n3829 VDD.n3808 0.0022058
R19435 VDD.n4087 VDD.n4066 0.0022058
R19436 VDD.n4345 VDD.n4324 0.0022058
R19437 VDD.n4603 VDD.n4582 0.0022058
R19438 VDD.n4861 VDD.n4840 0.0022058
R19439 VDD.n5153 VDD.n5132 0.0022058
R19440 VDD.n1745 VDD.n1724 0.0022058
R19441 VDD.n2094 VDD.n2073 0.0022058
R19442 VDD.n2324 VDD.n2303 0.0022058
R19443 VDD.n2582 VDD.n2561 0.0022058
R19444 VDD.n2840 VDD.n2819 0.0022058
R19445 VDD.n3098 VDD.n3077 0.0022058
R19446 VDD.n3356 VDD.n3335 0.0022058
R19447 VDD.n5686 VDD.n5665 0.0022058
R19448 VDD.n5432 VDD.n5411 0.0022058
R19449 VDD.n3614 VDD.n3593 0.0022058
R19450 VDD.n3872 VDD.n3851 0.0022058
R19451 VDD.n4130 VDD.n4109 0.0022058
R19452 VDD.n4388 VDD.n4367 0.0022058
R19453 VDD.n4646 VDD.n4625 0.0022058
R19454 VDD.n4904 VDD.n4883 0.0022058
R19455 VDD.n5196 VDD.n5175 0.0022058
R19456 VDD.n906 VDD.n904 0.00218421
R19457 VDD.n111 VDD.n109 0.00218421
R19458 VDD.n1745 VDD.n1744 0.00212475
R19459 VDD.n1681 VDD.n1678 0.00212475
R19460 VDD.n1732 VDD.n1712 0.00212475
R19461 VDD.n2094 VDD.n2093 0.00212475
R19462 VDD.n2030 VDD.n2027 0.00212475
R19463 VDD.n2081 VDD.n2061 0.00212475
R19464 VDD.n2324 VDD.n2323 0.00212475
R19465 VDD.n2260 VDD.n2257 0.00212475
R19466 VDD.n2311 VDD.n2291 0.00212475
R19467 VDD.n2582 VDD.n2581 0.00212475
R19468 VDD.n2518 VDD.n2515 0.00212475
R19469 VDD.n2569 VDD.n2549 0.00212475
R19470 VDD.n2840 VDD.n2839 0.00212475
R19471 VDD.n2776 VDD.n2773 0.00212475
R19472 VDD.n2827 VDD.n2807 0.00212475
R19473 VDD.n3098 VDD.n3097 0.00212475
R19474 VDD.n3034 VDD.n3031 0.00212475
R19475 VDD.n3085 VDD.n3065 0.00212475
R19476 VDD.n3356 VDD.n3355 0.00212475
R19477 VDD.n3292 VDD.n3289 0.00212475
R19478 VDD.n3343 VDD.n3323 0.00212475
R19479 VDD.n5686 VDD.n5685 0.00212475
R19480 VDD.n5622 VDD.n5619 0.00212475
R19481 VDD.n5673 VDD.n5653 0.00212475
R19482 VDD.n5432 VDD.n5431 0.00212475
R19483 VDD.n5368 VDD.n5365 0.00212475
R19484 VDD.n5419 VDD.n5399 0.00212475
R19485 VDD.n3614 VDD.n3613 0.00212475
R19486 VDD.n3550 VDD.n3547 0.00212475
R19487 VDD.n3601 VDD.n3581 0.00212475
R19488 VDD.n3872 VDD.n3871 0.00212475
R19489 VDD.n3808 VDD.n3805 0.00212475
R19490 VDD.n3859 VDD.n3839 0.00212475
R19491 VDD.n4130 VDD.n4129 0.00212475
R19492 VDD.n4066 VDD.n4063 0.00212475
R19493 VDD.n4117 VDD.n4097 0.00212475
R19494 VDD.n4388 VDD.n4387 0.00212475
R19495 VDD.n4324 VDD.n4321 0.00212475
R19496 VDD.n4375 VDD.n4355 0.00212475
R19497 VDD.n4646 VDD.n4645 0.00212475
R19498 VDD.n4582 VDD.n4579 0.00212475
R19499 VDD.n4633 VDD.n4613 0.00212475
R19500 VDD.n4904 VDD.n4903 0.00212475
R19501 VDD.n4840 VDD.n4837 0.00212475
R19502 VDD.n4891 VDD.n4871 0.00212475
R19503 VDD.n5196 VDD.n5195 0.00212475
R19504 VDD.n5132 VDD.n5129 0.00212475
R19505 VDD.n5183 VDD.n5163 0.00212475
R19506 VDD.n5229 VDD.n5085 0.00202384
R19507 VDD VDD.n1599 0.00202016
R19508 VDD.n22 VDD.n3 0.00195349
R19509 VDD.n21 VDD.n4 0.00195349
R19510 VDD.n17 VDD.n16 0.00195349
R19511 VDD.n15 VDD.n14 0.00195349
R19512 VDD.n11 VDD.n10 0.00195349
R19513 VDD.n339 VDD.n320 0.00195349
R19514 VDD.n338 VDD.n321 0.00195349
R19515 VDD.n334 VDD.n333 0.00195349
R19516 VDD.n332 VDD.n331 0.00195349
R19517 VDD.n328 VDD.n327 0.00195349
R19518 VDD.n601 VDD.n600 0.00194737
R19519 VDD.n598 VDD.n597 0.00194737
R19520 VDD.n1757 VDD.n1756 0.00194704
R19521 VDD.n2106 VDD.n2105 0.00194704
R19522 VDD.n2336 VDD.n2335 0.00194704
R19523 VDD.n2594 VDD.n2593 0.00194704
R19524 VDD.n2852 VDD.n2851 0.00194704
R19525 VDD.n3110 VDD.n3109 0.00194704
R19526 VDD.n3368 VDD.n3367 0.00194704
R19527 VDD.n5698 VDD.n5697 0.00194704
R19528 VDD.n5444 VDD.n5443 0.00194704
R19529 VDD.n3626 VDD.n3625 0.00194704
R19530 VDD.n3884 VDD.n3883 0.00194704
R19531 VDD.n4142 VDD.n4141 0.00194704
R19532 VDD.n4400 VDD.n4399 0.00194704
R19533 VDD.n4658 VDD.n4657 0.00194704
R19534 VDD.n4916 VDD.n4915 0.00194704
R19535 VDD.n5208 VDD.n5207 0.00194704
R19536 VDD.n1112 VDD.n1111 0.00190323
R19537 VDD.n1735 VDD.n1730 0.00188889
R19538 VDD.n2084 VDD.n2079 0.00188889
R19539 VDD.n2314 VDD.n2309 0.00188889
R19540 VDD.n2572 VDD.n2567 0.00188889
R19541 VDD.n2830 VDD.n2825 0.00188889
R19542 VDD.n3088 VDD.n3083 0.00188889
R19543 VDD.n3346 VDD.n3341 0.00188889
R19544 VDD.n5676 VDD.n5671 0.00188889
R19545 VDD.n5422 VDD.n5417 0.00188889
R19546 VDD.n3604 VDD.n3599 0.00188889
R19547 VDD.n3862 VDD.n3857 0.00188889
R19548 VDD.n4120 VDD.n4115 0.00188889
R19549 VDD.n4378 VDD.n4373 0.00188889
R19550 VDD.n4636 VDD.n4631 0.00188889
R19551 VDD.n4894 VDD.n4889 0.00188889
R19552 VDD.n5186 VDD.n5181 0.00188889
R19553 VDD.n1426 VDD.n1345 0.00182979
R19554 VDD.n1401 VDD.n1399 0.00182979
R19555 VDD.n1369 VDD.n1361 0.00182979
R19556 VDD.n1509 VDD.n1506 0.00182979
R19557 VDD.n1459 VDD.n1289 0.00182979
R19558 VDD.n1599 VDD.n1598 0.00178629
R19559 VDD.n1803 VDD.n1777 0.00175592
R19560 VDD.n1802 VDD.n1777 0.00175592
R19561 VDD.n2011 VDD.n1985 0.00175592
R19562 VDD.n2010 VDD.n1985 0.00175592
R19563 VDD.n2382 VDD.n2356 0.00175592
R19564 VDD.n2381 VDD.n2356 0.00175592
R19565 VDD.n2640 VDD.n2614 0.00175592
R19566 VDD.n2639 VDD.n2614 0.00175592
R19567 VDD.n2898 VDD.n2872 0.00175592
R19568 VDD.n2897 VDD.n2872 0.00175592
R19569 VDD.n3156 VDD.n3130 0.00175592
R19570 VDD.n3155 VDD.n3130 0.00175592
R19571 VDD.n3414 VDD.n3388 0.00175592
R19572 VDD.n3413 VDD.n3388 0.00175592
R19573 VDD.n5744 VDD.n5718 0.00175592
R19574 VDD.n5743 VDD.n5718 0.00175592
R19575 VDD.n5490 VDD.n5464 0.00175592
R19576 VDD.n5489 VDD.n5464 0.00175592
R19577 VDD.n3672 VDD.n3646 0.00175592
R19578 VDD.n3671 VDD.n3646 0.00175592
R19579 VDD.n3930 VDD.n3904 0.00175592
R19580 VDD.n3929 VDD.n3904 0.00175592
R19581 VDD.n4188 VDD.n4162 0.00175592
R19582 VDD.n4187 VDD.n4162 0.00175592
R19583 VDD.n4446 VDD.n4420 0.00175592
R19584 VDD.n4445 VDD.n4420 0.00175592
R19585 VDD.n4704 VDD.n4678 0.00175592
R19586 VDD.n4703 VDD.n4678 0.00175592
R19587 VDD.n4963 VDD.n4937 0.00175592
R19588 VDD.n4962 VDD.n4937 0.00175592
R19589 VDD.n5113 VDD.n5087 0.00175592
R19590 VDD.n5112 VDD.n5087 0.00175592
R19591 VDD.n4968 VDD.n4965 0.00169131
R19592 VDD.n1838 VDD.n1825 0.00162613
R19593 VDD.n2159 VDD.n2146 0.00162613
R19594 VDD.n2417 VDD.n2404 0.00162613
R19595 VDD.n2675 VDD.n2662 0.00162613
R19596 VDD.n2933 VDD.n2920 0.00162613
R19597 VDD.n3191 VDD.n3178 0.00162613
R19598 VDD.n3449 VDD.n3436 0.00162613
R19599 VDD.n5776 VDD.n5763 0.00162613
R19600 VDD.n5522 VDD.n5509 0.00162613
R19601 VDD.n3707 VDD.n3694 0.00162613
R19602 VDD.n3965 VDD.n3952 0.00162613
R19603 VDD.n4223 VDD.n4210 0.00162613
R19604 VDD.n4481 VDD.n4468 0.00162613
R19605 VDD.n4739 VDD.n4726 0.00162613
R19606 VDD.n5000 VDD.n4987 0.00162613
R19607 VDD.n5262 VDD.n5249 0.00162613
R19608 VDD.n1921 VDD.n1664 0.00162258
R19609 VDD.n2242 VDD.n1983 0.00162258
R19610 VDD.n2500 VDD.n2243 0.00162258
R19611 VDD.n2758 VDD.n2501 0.00162258
R19612 VDD.n3016 VDD.n2759 0.00162258
R19613 VDD.n3274 VDD.n3017 0.00162258
R19614 VDD.n3532 VDD.n3275 0.00162258
R19615 VDD.n3790 VDD.n3533 0.00162258
R19616 VDD.n4048 VDD.n3791 0.00162258
R19617 VDD.n4306 VDD.n4049 0.00162258
R19618 VDD.n4564 VDD.n4307 0.00162258
R19619 VDD.n4822 VDD.n4565 0.00162258
R19620 VDD.n1815 VDD.n1810 0.00161113
R19621 VDD.n2136 VDD.n2131 0.00161113
R19622 VDD.n2394 VDD.n2389 0.00161113
R19623 VDD.n2652 VDD.n2647 0.00161113
R19624 VDD.n2910 VDD.n2905 0.00161113
R19625 VDD.n3168 VDD.n3163 0.00161113
R19626 VDD.n3426 VDD.n3421 0.00161113
R19627 VDD.n5753 VDD.n5748 0.00161113
R19628 VDD.n5499 VDD.n5494 0.00161113
R19629 VDD.n3684 VDD.n3679 0.00161113
R19630 VDD.n3942 VDD.n3937 0.00161113
R19631 VDD.n4200 VDD.n4195 0.00161113
R19632 VDD.n4458 VDD.n4453 0.00161113
R19633 VDD.n4716 VDD.n4711 0.00161113
R19634 VDD.n4977 VDD.n4972 0.00161113
R19635 VDD.n5239 VDD.n5234 0.00161113
R19636 VDD.n1808 VDD.n1664 0.00160808
R19637 VDD.n2129 VDD.n1983 0.00160808
R19638 VDD.n2387 VDD.n2243 0.00160808
R19639 VDD.n2645 VDD.n2501 0.00160808
R19640 VDD.n2903 VDD.n2759 0.00160808
R19641 VDD.n3161 VDD.n3017 0.00160808
R19642 VDD.n3419 VDD.n3275 0.00160808
R19643 VDD.n3677 VDD.n3533 0.00160808
R19644 VDD.n3935 VDD.n3791 0.00160808
R19645 VDD.n4193 VDD.n4049 0.00160808
R19646 VDD.n4451 VDD.n4307 0.00160808
R19647 VDD.n4709 VDD.n4565 0.00160808
R19648 VDD.n4970 VDD.n4965 0.00160622
R19649 VDD.n5230 VDD.n5115 0.00159967
R19650 VDD.n1949 VDD.n1942 0.00158558
R19651 VDD.n1931 VDD.n1930 0.00158558
R19652 VDD.n1807 VDD.n1775 0.00157581
R19653 VDD.n2127 VDD.n2124 0.00157581
R19654 VDD.n2386 VDD.n2354 0.00157581
R19655 VDD.n2644 VDD.n2612 0.00157581
R19656 VDD.n2902 VDD.n2870 0.00157581
R19657 VDD.n3160 VDD.n3128 0.00157581
R19658 VDD.n3418 VDD.n3386 0.00157581
R19659 VDD.n3676 VDD.n3644 0.00157581
R19660 VDD.n3934 VDD.n3902 0.00157581
R19661 VDD.n4192 VDD.n4160 0.00157581
R19662 VDD.n4450 VDD.n4418 0.00157581
R19663 VDD.n4708 VDD.n4676 0.00157581
R19664 VDD.n5232 VDD.n5115 0.00152113
R19665 VDD.n1801 VDD.n1800 0.00151809
R19666 VDD.n2009 VDD.n2008 0.00151809
R19667 VDD.n2380 VDD.n2379 0.00151809
R19668 VDD.n2638 VDD.n2637 0.00151809
R19669 VDD.n2896 VDD.n2895 0.00151809
R19670 VDD.n3154 VDD.n3153 0.00151809
R19671 VDD.n3412 VDD.n3411 0.00151809
R19672 VDD.n5742 VDD.n5741 0.00151809
R19673 VDD.n5488 VDD.n5487 0.00151809
R19674 VDD.n3670 VDD.n3669 0.00151809
R19675 VDD.n3928 VDD.n3927 0.00151809
R19676 VDD.n4186 VDD.n4185 0.00151809
R19677 VDD.n4444 VDD.n4443 0.00151809
R19678 VDD.n4702 VDD.n4701 0.00151809
R19679 VDD.n4961 VDD.n4960 0.00151809
R19680 VDD.n5111 VDD.n5110 0.00151809
R19681 VDD.n1801 VDD.n1777 0.00149567
R19682 VDD.n2009 VDD.n1985 0.00149567
R19683 VDD.n2380 VDD.n2356 0.00149567
R19684 VDD.n2638 VDD.n2614 0.00149567
R19685 VDD.n2896 VDD.n2872 0.00149567
R19686 VDD.n3154 VDD.n3130 0.00149567
R19687 VDD.n3412 VDD.n3388 0.00149567
R19688 VDD.n5742 VDD.n5718 0.00149567
R19689 VDD.n5488 VDD.n5464 0.00149567
R19690 VDD.n3670 VDD.n3646 0.00149567
R19691 VDD.n3928 VDD.n3904 0.00149567
R19692 VDD.n4186 VDD.n4162 0.00149567
R19693 VDD.n4444 VDD.n4420 0.00149567
R19694 VDD.n4702 VDD.n4678 0.00149567
R19695 VDD.n4961 VDD.n4937 0.00149567
R19696 VDD.n5111 VDD.n5087 0.00149567
R19697 VDD.n1917 VDD.n1916 0.00148913
R19698 VDD.n2238 VDD.n2237 0.00148913
R19699 VDD.n2496 VDD.n2495 0.00148913
R19700 VDD.n2754 VDD.n2753 0.00148913
R19701 VDD.n3012 VDD.n3011 0.00148913
R19702 VDD.n3270 VDD.n3269 0.00148913
R19703 VDD.n3528 VDD.n3527 0.00148913
R19704 VDD.n5855 VDD.n5854 0.00148913
R19705 VDD.n5601 VDD.n5600 0.00148913
R19706 VDD.n3786 VDD.n3785 0.00148913
R19707 VDD.n4044 VDD.n4043 0.00148913
R19708 VDD.n4302 VDD.n4301 0.00148913
R19709 VDD.n4560 VDD.n4559 0.00148913
R19710 VDD.n4818 VDD.n4817 0.00148913
R19711 VDD.n5079 VDD.n5078 0.00148913
R19712 VDD.n5341 VDD.n5340 0.00148913
R19713 VDD.n1602 VDD.n1601 0.00147143
R19714 VDD.n1806 VDD.n1805 0.00147065
R19715 VDD.n2126 VDD.n2125 0.00147065
R19716 VDD.n2385 VDD.n2384 0.00147065
R19717 VDD.n2643 VDD.n2642 0.00147065
R19718 VDD.n2901 VDD.n2900 0.00147065
R19719 VDD.n3159 VDD.n3158 0.00147065
R19720 VDD.n3417 VDD.n3416 0.00147065
R19721 VDD.n3675 VDD.n3674 0.00147065
R19722 VDD.n3933 VDD.n3932 0.00147065
R19723 VDD.n4191 VDD.n4190 0.00147065
R19724 VDD.n4449 VDD.n4448 0.00147065
R19725 VDD.n4707 VDD.n4706 0.00147065
R19726 VDD.n1769 VDD.n1670 0.00145131
R19727 VDD.n1711 VDD.n1670 0.00145131
R19728 VDD.n2118 VDD.n2019 0.00145131
R19729 VDD.n2060 VDD.n2019 0.00145131
R19730 VDD.n2348 VDD.n2249 0.00145131
R19731 VDD.n2290 VDD.n2249 0.00145131
R19732 VDD.n2606 VDD.n2507 0.00145131
R19733 VDD.n2548 VDD.n2507 0.00145131
R19734 VDD.n2864 VDD.n2765 0.00145131
R19735 VDD.n2806 VDD.n2765 0.00145131
R19736 VDD.n3122 VDD.n3023 0.00145131
R19737 VDD.n3064 VDD.n3023 0.00145131
R19738 VDD.n3380 VDD.n3281 0.00145131
R19739 VDD.n3322 VDD.n3281 0.00145131
R19740 VDD.n5710 VDD.n5611 0.00145131
R19741 VDD.n5652 VDD.n5611 0.00145131
R19742 VDD.n5456 VDD.n5357 0.00145131
R19743 VDD.n5398 VDD.n5357 0.00145131
R19744 VDD.n3638 VDD.n3539 0.00145131
R19745 VDD.n3580 VDD.n3539 0.00145131
R19746 VDD.n3896 VDD.n3797 0.00145131
R19747 VDD.n3838 VDD.n3797 0.00145131
R19748 VDD.n4154 VDD.n4055 0.00145131
R19749 VDD.n4096 VDD.n4055 0.00145131
R19750 VDD.n4412 VDD.n4313 0.00145131
R19751 VDD.n4354 VDD.n4313 0.00145131
R19752 VDD.n4670 VDD.n4571 0.00145131
R19753 VDD.n4612 VDD.n4571 0.00145131
R19754 VDD.n4928 VDD.n4829 0.00145131
R19755 VDD.n4870 VDD.n4829 0.00145131
R19756 VDD.n5220 VDD.n5121 0.00145131
R19757 VDD.n5162 VDD.n5121 0.00145131
R19758 VDD.n1770 VDD.n1769 0.00145112
R19759 VDD.n2119 VDD.n2118 0.00145112
R19760 VDD.n2349 VDD.n2348 0.00145112
R19761 VDD.n2607 VDD.n2606 0.00145112
R19762 VDD.n2865 VDD.n2864 0.00145112
R19763 VDD.n3123 VDD.n3122 0.00145112
R19764 VDD.n3381 VDD.n3380 0.00145112
R19765 VDD.n5711 VDD.n5710 0.00145112
R19766 VDD.n5457 VDD.n5456 0.00145112
R19767 VDD.n3639 VDD.n3638 0.00145112
R19768 VDD.n3897 VDD.n3896 0.00145112
R19769 VDD.n4155 VDD.n4154 0.00145112
R19770 VDD.n4413 VDD.n4412 0.00145112
R19771 VDD.n4671 VDD.n4670 0.00145112
R19772 VDD.n4929 VDD.n4928 0.00145112
R19773 VDD.n5221 VDD.n5220 0.00145112
R19774 VDD.n1756 VDD.n1755 0.00144714
R19775 VDD.n2105 VDD.n2104 0.00144714
R19776 VDD.n2335 VDD.n2334 0.00144714
R19777 VDD.n2593 VDD.n2592 0.00144714
R19778 VDD.n2851 VDD.n2850 0.00144714
R19779 VDD.n3109 VDD.n3108 0.00144714
R19780 VDD.n3367 VDD.n3366 0.00144714
R19781 VDD.n5697 VDD.n5696 0.00144714
R19782 VDD.n5443 VDD.n5442 0.00144714
R19783 VDD.n3625 VDD.n3624 0.00144714
R19784 VDD.n3883 VDD.n3882 0.00144714
R19785 VDD.n4141 VDD.n4140 0.00144714
R19786 VDD.n4399 VDD.n4398 0.00144714
R19787 VDD.n4657 VDD.n4656 0.00144714
R19788 VDD.n4915 VDD.n4914 0.00144714
R19789 VDD.n5207 VDD.n5206 0.00144714
R19790 VDD.n1755 VDD.n1754 0.00144695
R19791 VDD.n2104 VDD.n2103 0.00144695
R19792 VDD.n2334 VDD.n2333 0.00144695
R19793 VDD.n2592 VDD.n2591 0.00144695
R19794 VDD.n2850 VDD.n2849 0.00144695
R19795 VDD.n3108 VDD.n3107 0.00144695
R19796 VDD.n3366 VDD.n3365 0.00144695
R19797 VDD.n5696 VDD.n5695 0.00144695
R19798 VDD.n5442 VDD.n5441 0.00144695
R19799 VDD.n3624 VDD.n3623 0.00144695
R19800 VDD.n3882 VDD.n3881 0.00144695
R19801 VDD.n4140 VDD.n4139 0.00144695
R19802 VDD.n4398 VDD.n4397 0.00144695
R19803 VDD.n4656 VDD.n4655 0.00144695
R19804 VDD.n4914 VDD.n4913 0.00144695
R19805 VDD.n5206 VDD.n5205 0.00144695
R19806 VDD.n1115 VDD.n1114 0.00143548
R19807 VDD.n1003 VDD.n1002 0.00142105
R19808 VDD.n208 VDD.n207 0.00142105
R19809 VDD.n1978 VDD.n1924 0.00139286
R19810 VDD.n1719 VDD.n1668 0.00139286
R19811 VDD.n2068 VDD.n2017 0.00139286
R19812 VDD.n2298 VDD.n2247 0.00139286
R19813 VDD.n2556 VDD.n2505 0.00139286
R19814 VDD.n2814 VDD.n2763 0.00139286
R19815 VDD.n3072 VDD.n3021 0.00139286
R19816 VDD.n3330 VDD.n3279 0.00139286
R19817 VDD.n5660 VDD.n5609 0.00139286
R19818 VDD.n5406 VDD.n5355 0.00139286
R19819 VDD.n3588 VDD.n3537 0.00139286
R19820 VDD.n3846 VDD.n3795 0.00139286
R19821 VDD.n4104 VDD.n4053 0.00139286
R19822 VDD.n4362 VDD.n4311 0.00139286
R19823 VDD.n4620 VDD.n4569 0.00139286
R19824 VDD.n4878 VDD.n4827 0.00139286
R19825 VDD.n5170 VDD.n5119 0.00139286
R19826 VDD.t1285 VDD.n1941 0.00134143
R19827 VDD.n4969 VDD.n4966 0.00133929
R19828 VDD.n5231 VDD.n5228 0.00133929
R19829 VDD.n1885 VDD.n1819 0.00133663
R19830 VDD.n1821 VDD.n1819 0.00133663
R19831 VDD.n2206 VDD.n2140 0.00133663
R19832 VDD.n2142 VDD.n2140 0.00133663
R19833 VDD.n2464 VDD.n2398 0.00133663
R19834 VDD.n2400 VDD.n2398 0.00133663
R19835 VDD.n2722 VDD.n2656 0.00133663
R19836 VDD.n2658 VDD.n2656 0.00133663
R19837 VDD.n2980 VDD.n2914 0.00133663
R19838 VDD.n2916 VDD.n2914 0.00133663
R19839 VDD.n3238 VDD.n3172 0.00133663
R19840 VDD.n3174 VDD.n3172 0.00133663
R19841 VDD.n3496 VDD.n3430 0.00133663
R19842 VDD.n3432 VDD.n3430 0.00133663
R19843 VDD.n5823 VDD.n5757 0.00133663
R19844 VDD.n5759 VDD.n5757 0.00133663
R19845 VDD.n5569 VDD.n5503 0.00133663
R19846 VDD.n5505 VDD.n5503 0.00133663
R19847 VDD.n3754 VDD.n3688 0.00133663
R19848 VDD.n3690 VDD.n3688 0.00133663
R19849 VDD.n4012 VDD.n3946 0.00133663
R19850 VDD.n3948 VDD.n3946 0.00133663
R19851 VDD.n4270 VDD.n4204 0.00133663
R19852 VDD.n4206 VDD.n4204 0.00133663
R19853 VDD.n4528 VDD.n4462 0.00133663
R19854 VDD.n4464 VDD.n4462 0.00133663
R19855 VDD.n4786 VDD.n4720 0.00133663
R19856 VDD.n4722 VDD.n4720 0.00133663
R19857 VDD.n5047 VDD.n4981 0.00133663
R19858 VDD.n4983 VDD.n4981 0.00133663
R19859 VDD.n5309 VDD.n5243 0.00133663
R19860 VDD.n5245 VDD.n5243 0.00133663
R19861 VDD.n1981 VDD 0.00130357
R19862 VDD.n600 VDD 0.00128947
R19863 VDD.n1805 VDD.n1775 0.00120516
R19864 VDD.n2125 VDD.n2124 0.00120516
R19865 VDD.n2384 VDD.n2354 0.00120516
R19866 VDD.n2642 VDD.n2612 0.00120516
R19867 VDD.n2900 VDD.n2870 0.00120516
R19868 VDD.n3158 VDD.n3128 0.00120516
R19869 VDD.n3416 VDD.n3386 0.00120516
R19870 VDD.n3674 VDD.n3644 0.00120516
R19871 VDD.n3932 VDD.n3902 0.00120516
R19872 VDD.n4190 VDD.n4160 0.00120516
R19873 VDD.n4448 VDD.n4418 0.00120516
R19874 VDD.n4706 VDD.n4676 0.00120516
R19875 VDD.n5866 VDD.n5865 0.00119048
R19876 VDD.n1172 VDD.n1138 0.00116652
R19877 VDD.n1238 VDD.n1204 0.00116652
R19878 VDD.n5344 VDD.n5343 0.00115375
R19879 VDD.n5082 VDD.n5081 0.00115374
R19880 VDD.n1176 VDD.n1175 0.00114708
R19881 VDD.n1175 VDD.n1173 0.00114708
R19882 VDD.n1242 VDD.n1241 0.00114708
R19883 VDD.n1241 VDD.n1239 0.00114708
R19884 VDD.n1871 VDD.n1844 0.00114565
R19885 VDD.n1847 VDD.n1844 0.00114565
R19886 VDD.n2192 VDD.n2165 0.00114565
R19887 VDD.n2168 VDD.n2165 0.00114565
R19888 VDD.n2450 VDD.n2423 0.00114565
R19889 VDD.n2426 VDD.n2423 0.00114565
R19890 VDD.n2708 VDD.n2681 0.00114565
R19891 VDD.n2684 VDD.n2681 0.00114565
R19892 VDD.n2966 VDD.n2939 0.00114565
R19893 VDD.n2942 VDD.n2939 0.00114565
R19894 VDD.n3224 VDD.n3197 0.00114565
R19895 VDD.n3200 VDD.n3197 0.00114565
R19896 VDD.n3482 VDD.n3455 0.00114565
R19897 VDD.n3458 VDD.n3455 0.00114565
R19898 VDD.n5809 VDD.n5782 0.00114565
R19899 VDD.n5785 VDD.n5782 0.00114565
R19900 VDD.n5555 VDD.n5528 0.00114565
R19901 VDD.n5531 VDD.n5528 0.00114565
R19902 VDD.n3740 VDD.n3713 0.00114565
R19903 VDD.n3716 VDD.n3713 0.00114565
R19904 VDD.n3998 VDD.n3971 0.00114565
R19905 VDD.n3974 VDD.n3971 0.00114565
R19906 VDD.n4256 VDD.n4229 0.00114565
R19907 VDD.n4232 VDD.n4229 0.00114565
R19908 VDD.n4514 VDD.n4487 0.00114565
R19909 VDD.n4490 VDD.n4487 0.00114565
R19910 VDD.n4772 VDD.n4745 0.00114565
R19911 VDD.n4748 VDD.n4745 0.00114565
R19912 VDD.n5033 VDD.n5006 0.00114565
R19913 VDD.n5009 VDD.n5006 0.00114565
R19914 VDD.n5295 VDD.n5268 0.00114565
R19915 VDD.n5271 VDD.n5268 0.00114565
R19916 VDD.n1739 VDD.n1738 0.00113805
R19917 VDD.n2088 VDD.n2087 0.00113805
R19918 VDD.n2318 VDD.n2317 0.00113805
R19919 VDD.n2576 VDD.n2575 0.00113805
R19920 VDD.n2834 VDD.n2833 0.00113805
R19921 VDD.n3092 VDD.n3091 0.00113805
R19922 VDD.n3350 VDD.n3349 0.00113805
R19923 VDD.n5680 VDD.n5679 0.00113805
R19924 VDD.n5426 VDD.n5425 0.00113805
R19925 VDD.n3608 VDD.n3607 0.00113805
R19926 VDD.n3866 VDD.n3865 0.00113805
R19927 VDD.n4124 VDD.n4123 0.00113805
R19928 VDD.n4382 VDD.n4381 0.00113805
R19929 VDD.n4640 VDD.n4639 0.00113805
R19930 VDD.n4898 VDD.n4897 0.00113805
R19931 VDD.n5190 VDD.n5189 0.00113805
R19932 VDD.n1621 VDD.n1620 0.00111657
R19933 VDD.n1976 VDD.n1975 0.00111635
R19934 VDD.t1287 VDD.n1969 0.0010973
R19935 VDD.n5227 VDD.n5085 0.00109697
R19936 VDD.n1798 VDD.n1797 0.00108642
R19937 VDD.n2006 VDD.n2005 0.00108642
R19938 VDD.n2377 VDD.n2376 0.00108642
R19939 VDD.n2635 VDD.n2634 0.00108642
R19940 VDD.n2893 VDD.n2892 0.00108642
R19941 VDD.n3151 VDD.n3150 0.00108642
R19942 VDD.n3409 VDD.n3408 0.00108642
R19943 VDD.n5739 VDD.n5738 0.00108642
R19944 VDD.n5485 VDD.n5484 0.00108642
R19945 VDD.n3667 VDD.n3666 0.00108642
R19946 VDD.n3925 VDD.n3924 0.00108642
R19947 VDD.n4183 VDD.n4182 0.00108642
R19948 VDD.n4441 VDD.n4440 0.00108642
R19949 VDD.n4699 VDD.n4698 0.00108642
R19950 VDD.n4958 VDD.n4957 0.00108642
R19951 VDD.n5108 VDD.n5107 0.00108642
R19952 VDD.n4968 VDD.n4967 0.00108509
R19953 VDD.n1177 VDD.n1176 0.00107711
R19954 VDD.n1243 VDD.n1242 0.00107711
R19955 VDD.n1642 VDD.n1641 0.00107006
R19956 VDD.n1613 VDD.n1612 0.00106596
R19957 VDD.n1752 VDD.n1720 0.00105202
R19958 VDD.n2101 VDD.n2069 0.00105202
R19959 VDD.n2331 VDD.n2299 0.00105202
R19960 VDD.n2589 VDD.n2557 0.00105202
R19961 VDD.n2847 VDD.n2815 0.00105202
R19962 VDD.n3105 VDD.n3073 0.00105202
R19963 VDD.n3363 VDD.n3331 0.00105202
R19964 VDD.n5693 VDD.n5661 0.00105202
R19965 VDD.n5439 VDD.n5407 0.00105202
R19966 VDD.n3621 VDD.n3589 0.00105202
R19967 VDD.n3879 VDD.n3847 0.00105202
R19968 VDD.n4137 VDD.n4105 0.00105202
R19969 VDD.n4395 VDD.n4363 0.00105202
R19970 VDD.n4653 VDD.n4621 0.00105202
R19971 VDD.n4911 VDD.n4879 0.00105202
R19972 VDD.n5203 VDD.n5171 0.00105202
R19973 VDD.n1431 VDD.n1430 0.00100344
R19974 VDD.n1455 VDD.n1454 0.00100344
R19975 VDD.n1374 VDD.n1373 0.00100342
R19976 VDD.n1711 VDD.n1710 0.00100293
R19977 VDD.n2060 VDD.n2059 0.00100293
R19978 VDD.n2290 VDD.n2289 0.00100293
R19979 VDD.n2548 VDD.n2547 0.00100293
R19980 VDD.n2806 VDD.n2805 0.00100293
R19981 VDD.n3064 VDD.n3063 0.00100293
R19982 VDD.n3322 VDD.n3321 0.00100293
R19983 VDD.n5652 VDD.n5651 0.00100293
R19984 VDD.n5398 VDD.n5397 0.00100293
R19985 VDD.n3580 VDD.n3579 0.00100293
R19986 VDD.n3838 VDD.n3837 0.00100293
R19987 VDD.n4096 VDD.n4095 0.00100293
R19988 VDD.n4354 VDD.n4353 0.00100293
R19989 VDD.n4612 VDD.n4611 0.00100293
R19990 VDD.n4870 VDD.n4869 0.00100293
R19991 VDD.n5162 VDD.n5161 0.00100293
R19992 VDD.n781 VDD.n780 0.00100258
R19993 VDD.n378 VDD.n377 0.00100258
R19994 VDD.n1837 VDD.n1826 0.00100132
R19995 VDD.n2158 VDD.n2147 0.00100132
R19996 VDD.n2416 VDD.n2405 0.00100132
R19997 VDD.n2674 VDD.n2663 0.00100132
R19998 VDD.n2932 VDD.n2921 0.00100132
R19999 VDD.n3190 VDD.n3179 0.00100132
R20000 VDD.n3448 VDD.n3437 0.00100132
R20001 VDD.n5775 VDD.n5764 0.00100132
R20002 VDD.n5521 VDD.n5510 0.00100132
R20003 VDD.n3706 VDD.n3695 0.00100132
R20004 VDD.n3964 VDD.n3953 0.00100132
R20005 VDD.n4222 VDD.n4211 0.00100132
R20006 VDD.n4480 VDD.n4469 0.00100132
R20007 VDD.n4738 VDD.n4727 0.00100132
R20008 VDD.n4999 VDD.n4988 0.00100132
R20009 VDD.n5261 VDD.n5250 0.00100132
R20010 VDD.n904 VDD.n903 0.00100097
R20011 VDD.n109 VDD.n108 0.00100097
R20012 VDD.n503 VDD.n502 0.00100097
R20013 VDD.n1547 VDD.n1541 0.00100097
R20014 VDD.n1620 VDD.n1614 0.00100057
R20015 VDD.n1798 VDD.n1777 0.00100033
R20016 VDD.n2006 VDD.n1985 0.00100033
R20017 VDD.n2377 VDD.n2356 0.00100033
R20018 VDD.n2635 VDD.n2614 0.00100033
R20019 VDD.n2893 VDD.n2872 0.00100033
R20020 VDD.n3151 VDD.n3130 0.00100033
R20021 VDD.n3409 VDD.n3388 0.00100033
R20022 VDD.n5739 VDD.n5718 0.00100033
R20023 VDD.n5485 VDD.n5464 0.00100033
R20024 VDD.n3667 VDD.n3646 0.00100033
R20025 VDD.n3925 VDD.n3904 0.00100033
R20026 VDD.n4183 VDD.n4162 0.00100033
R20027 VDD.n4441 VDD.n4420 0.00100033
R20028 VDD.n4699 VDD.n4678 0.00100033
R20029 VDD.n4958 VDD.n4937 0.00100033
R20030 VDD.n5108 VDD.n5087 0.00100033
R20031 VDD.n1882 VDD.n1821 0.00100021
R20032 VDD.n2203 VDD.n2142 0.00100021
R20033 VDD.n2461 VDD.n2400 0.00100021
R20034 VDD.n2719 VDD.n2658 0.00100021
R20035 VDD.n2977 VDD.n2916 0.00100021
R20036 VDD.n3235 VDD.n3174 0.00100021
R20037 VDD.n3493 VDD.n3432 0.00100021
R20038 VDD.n5820 VDD.n5759 0.00100021
R20039 VDD.n5566 VDD.n5505 0.00100021
R20040 VDD.n3751 VDD.n3690 0.00100021
R20041 VDD.n4009 VDD.n3948 0.00100021
R20042 VDD.n4267 VDD.n4206 0.00100021
R20043 VDD.n4525 VDD.n4464 0.00100021
R20044 VDD.n4783 VDD.n4722 0.00100021
R20045 VDD.n5044 VDD.n4983 0.00100021
R20046 VDD.n5306 VDD.n5245 0.00100021
R20047 VDD.n1177 VDD.n1172 0.00100013
R20048 VDD.n1243 VDD.n1238 0.00100013
R20049 VDD.n1757 VDD.n1711 0.0010001
R20050 VDD.n2106 VDD.n2060 0.0010001
R20051 VDD.n2336 VDD.n2290 0.0010001
R20052 VDD.n2594 VDD.n2548 0.0010001
R20053 VDD.n2852 VDD.n2806 0.0010001
R20054 VDD.n3110 VDD.n3064 0.0010001
R20055 VDD.n3368 VDD.n3322 0.0010001
R20056 VDD.n5698 VDD.n5652 0.0010001
R20057 VDD.n5444 VDD.n5398 0.0010001
R20058 VDD.n3626 VDD.n3580 0.0010001
R20059 VDD.n3884 VDD.n3838 0.0010001
R20060 VDD.n4142 VDD.n4096 0.0010001
R20061 VDD.n4400 VDD.n4354 0.0010001
R20062 VDD.n4658 VDD.n4612 0.0010001
R20063 VDD.n4916 VDD.n4870 0.0010001
R20064 VDD.n5208 VDD.n5162 0.0010001
R20065 VDD.n4967 VDD.n4966 0.00100008
R20066 VDD.n1641 VDD.n1640 0.00100008
R20067 VDD.n1952 VDD.n1944 0.00100003
R20068 VDD.n1934 VDD.n1927 0.00100003
R20069 VDD.n1920 VDD.n1808 0.00100002
R20070 VDD.n2241 VDD.n2129 0.00100002
R20071 VDD.n2499 VDD.n2387 0.00100002
R20072 VDD.n2757 VDD.n2645 0.00100002
R20073 VDD.n3015 VDD.n2903 0.00100002
R20074 VDD.n3273 VDD.n3161 0.00100002
R20075 VDD.n3531 VDD.n3419 0.00100002
R20076 VDD.n3789 VDD.n3677 0.00100002
R20077 VDD.n4047 VDD.n3935 0.00100002
R20078 VDD.n4305 VDD.n4193 0.00100002
R20079 VDD.n4563 VDD.n4451 0.00100002
R20080 VDD.n4821 VDD.n4709 0.00100002
R20081 VDD.n1317 VDD.n1315 0.001
R20082 VDD.n1975 VDD.n1927 0.001
R20083 VDD.n1979 VDD.n1923 0.001
R20084 VDD.n1175 VDD.n1174 0.001
R20085 VDD.n1241 VDD.n1240 0.001
R20086 VDD.n707 VDD.n706 0.000894737
R20087 VDD.n1640 VDD.n1638 0.000834423
R20088 VDD.n1460 VDD.n1459 0.000765957
R20089 VDD.n1005 VDD 0.000763158
R20090 VDD.n210 VDD 0.000763158
R20091 VDD.n1110 VDD.n832 0.000631579
R20092 VDD.n315 VDD.n37 0.000631579
R20093 VDD.n1621 VDD.n1615 0.000625544
R20094 VDD.n1619 VDD.n1615 0.000625542
R20095 VDD.n1977 VDD.n1976 0.00061635
R20096 VDD.n1978 VDD.n1977 0.000616347
R20097 VDD.n1736 VDD.n1729 0.000594432
R20098 VDD.n2085 VDD.n2078 0.000594432
R20099 VDD.n2315 VDD.n2308 0.000594432
R20100 VDD.n2573 VDD.n2566 0.000594432
R20101 VDD.n2831 VDD.n2824 0.000594432
R20102 VDD.n3089 VDD.n3082 0.000594432
R20103 VDD.n3347 VDD.n3340 0.000594432
R20104 VDD.n5677 VDD.n5670 0.000594432
R20105 VDD.n5423 VDD.n5416 0.000594432
R20106 VDD.n3605 VDD.n3598 0.000594432
R20107 VDD.n3863 VDD.n3856 0.000594432
R20108 VDD.n4121 VDD.n4114 0.000594432
R20109 VDD.n4379 VDD.n4372 0.000594432
R20110 VDD.n4637 VDD.n4630 0.000594432
R20111 VDD.n4895 VDD.n4888 0.000594432
R20112 VDD.n5187 VDD.n5180 0.000594432
R20113 VDD.n4969 VDD.n4968 0.000578904
R20114 VDD.n5231 VDD.n5230 0.000578904
R20115 VDD.n5230 VDD.n5229 0.000578548
R20116 VDD.n1773 VDD.n1772 0.000558569
R20117 VDD.n2122 VDD.n2121 0.000558569
R20118 VDD.n2352 VDD.n2351 0.000558569
R20119 VDD.n2610 VDD.n2609 0.000558569
R20120 VDD.n2868 VDD.n2867 0.000558569
R20121 VDD.n3126 VDD.n3125 0.000558569
R20122 VDD.n3384 VDD.n3383 0.000558569
R20123 VDD.n5714 VDD.n5713 0.000558569
R20124 VDD.n5460 VDD.n5459 0.000558569
R20125 VDD.n3642 VDD.n3641 0.000558569
R20126 VDD.n3900 VDD.n3899 0.000558569
R20127 VDD.n4158 VDD.n4157 0.000558569
R20128 VDD.n4416 VDD.n4415 0.000558569
R20129 VDD.n4674 VDD.n4673 0.000558569
R20130 VDD.n4932 VDD.n4931 0.000558569
R20131 VDD.n5224 VDD.n5223 0.000558569
R20132 VDD.n1740 VDD.n1739 0.000555817
R20133 VDD.n2089 VDD.n2088 0.000555817
R20134 VDD.n2319 VDD.n2318 0.000555817
R20135 VDD.n2577 VDD.n2576 0.000555817
R20136 VDD.n2835 VDD.n2834 0.000555817
R20137 VDD.n3093 VDD.n3092 0.000555817
R20138 VDD.n3351 VDD.n3350 0.000555817
R20139 VDD.n5681 VDD.n5680 0.000555817
R20140 VDD.n5427 VDD.n5426 0.000555817
R20141 VDD.n3609 VDD.n3608 0.000555817
R20142 VDD.n3867 VDD.n3866 0.000555817
R20143 VDD.n4125 VDD.n4124 0.000555817
R20144 VDD.n4383 VDD.n4382 0.000555817
R20145 VDD.n4641 VDD.n4640 0.000555817
R20146 VDD.n4899 VDD.n4898 0.000555817
R20147 VDD.n5191 VDD.n5190 0.000555817
R20148 VDD.n1768 VDD.n1668 0.000534058
R20149 VDD.n2117 VDD.n2017 0.000534058
R20150 VDD.n2347 VDD.n2247 0.000534058
R20151 VDD.n2605 VDD.n2505 0.000534058
R20152 VDD.n2863 VDD.n2763 0.000534058
R20153 VDD.n3121 VDD.n3021 0.000534058
R20154 VDD.n3379 VDD.n3279 0.000534058
R20155 VDD.n5709 VDD.n5609 0.000534058
R20156 VDD.n5455 VDD.n5355 0.000534058
R20157 VDD.n3637 VDD.n3537 0.000534058
R20158 VDD.n3895 VDD.n3795 0.000534058
R20159 VDD.n4153 VDD.n4053 0.000534058
R20160 VDD.n4411 VDD.n4311 0.000534058
R20161 VDD.n4669 VDD.n4569 0.000534058
R20162 VDD.n4927 VDD.n4827 0.000534058
R20163 VDD.n5219 VDD.n5119 0.000534058
R20164 VDD.n1886 VDD.n1885 0.000523376
R20165 VDD.n2207 VDD.n2206 0.000523376
R20166 VDD.n2465 VDD.n2464 0.000523376
R20167 VDD.n2723 VDD.n2722 0.000523376
R20168 VDD.n2981 VDD.n2980 0.000523376
R20169 VDD.n3239 VDD.n3238 0.000523376
R20170 VDD.n3497 VDD.n3496 0.000523376
R20171 VDD.n5824 VDD.n5823 0.000523376
R20172 VDD.n5570 VDD.n5569 0.000523376
R20173 VDD.n3755 VDD.n3754 0.000523376
R20174 VDD.n4013 VDD.n4012 0.000523376
R20175 VDD.n4271 VDD.n4270 0.000523376
R20176 VDD.n4529 VDD.n4528 0.000523376
R20177 VDD.n4787 VDD.n4786 0.000523376
R20178 VDD.n5048 VDD.n5047 0.000523376
R20179 VDD.n5310 VDD.n5309 0.000523376
R20180 VDD.n1704 VDD.n1703 0.000516232
R20181 VDD.n1691 VDD.n1685 0.000516232
R20182 VDD.n2053 VDD.n2052 0.000516232
R20183 VDD.n2040 VDD.n2034 0.000516232
R20184 VDD.n2283 VDD.n2282 0.000516232
R20185 VDD.n2270 VDD.n2264 0.000516232
R20186 VDD.n2541 VDD.n2540 0.000516232
R20187 VDD.n2528 VDD.n2522 0.000516232
R20188 VDD.n2799 VDD.n2798 0.000516232
R20189 VDD.n2786 VDD.n2780 0.000516232
R20190 VDD.n3057 VDD.n3056 0.000516232
R20191 VDD.n3044 VDD.n3038 0.000516232
R20192 VDD.n3315 VDD.n3314 0.000516232
R20193 VDD.n3302 VDD.n3296 0.000516232
R20194 VDD.n5645 VDD.n5644 0.000516232
R20195 VDD.n5632 VDD.n5626 0.000516232
R20196 VDD.n5391 VDD.n5390 0.000516232
R20197 VDD.n5378 VDD.n5372 0.000516232
R20198 VDD.n3573 VDD.n3572 0.000516232
R20199 VDD.n3560 VDD.n3554 0.000516232
R20200 VDD.n3831 VDD.n3830 0.000516232
R20201 VDD.n3818 VDD.n3812 0.000516232
R20202 VDD.n4089 VDD.n4088 0.000516232
R20203 VDD.n4076 VDD.n4070 0.000516232
R20204 VDD.n4347 VDD.n4346 0.000516232
R20205 VDD.n4334 VDD.n4328 0.000516232
R20206 VDD.n4605 VDD.n4604 0.000516232
R20207 VDD.n4592 VDD.n4586 0.000516232
R20208 VDD.n4863 VDD.n4862 0.000516232
R20209 VDD.n4850 VDD.n4844 0.000516232
R20210 VDD.n5155 VDD.n5154 0.000516232
R20211 VDD.n5142 VDD.n5136 0.000516232
R20212 VDD.n1735 VDD.n1734 0.000515622
R20213 VDD.n2084 VDD.n2083 0.000515622
R20214 VDD.n2314 VDD.n2313 0.000515622
R20215 VDD.n2572 VDD.n2571 0.000515622
R20216 VDD.n2830 VDD.n2829 0.000515622
R20217 VDD.n3088 VDD.n3087 0.000515622
R20218 VDD.n3346 VDD.n3345 0.000515622
R20219 VDD.n5676 VDD.n5675 0.000515622
R20220 VDD.n5422 VDD.n5421 0.000515622
R20221 VDD.n3604 VDD.n3603 0.000515622
R20222 VDD.n3862 VDD.n3861 0.000515622
R20223 VDD.n4120 VDD.n4119 0.000515622
R20224 VDD.n4378 VDD.n4377 0.000515622
R20225 VDD.n4636 VDD.n4635 0.000515622
R20226 VDD.n4894 VDD.n4893 0.000515622
R20227 VDD.n5186 VDD.n5185 0.000515622
R20228 VDD.n1876 VDD.n1875 0.000514451
R20229 VDD.n2197 VDD.n2196 0.000514451
R20230 VDD.n2455 VDD.n2454 0.000514451
R20231 VDD.n2713 VDD.n2712 0.000514451
R20232 VDD.n2971 VDD.n2970 0.000514451
R20233 VDD.n3229 VDD.n3228 0.000514451
R20234 VDD.n3487 VDD.n3486 0.000514451
R20235 VDD.n5814 VDD.n5813 0.000514451
R20236 VDD.n5560 VDD.n5559 0.000514451
R20237 VDD.n3745 VDD.n3744 0.000514451
R20238 VDD.n4003 VDD.n4002 0.000514451
R20239 VDD.n4261 VDD.n4260 0.000514451
R20240 VDD.n4519 VDD.n4518 0.000514451
R20241 VDD.n4777 VDD.n4776 0.000514451
R20242 VDD.n5038 VDD.n5037 0.000514451
R20243 VDD.n5300 VDD.n5299 0.000514451
R20244 VDD.n986 VDD.n838 0.000506553
R20245 VDD.n985 VDD.n835 0.000506553
R20246 VDD.n984 VDD.n983 0.000506553
R20247 VDD.n903 VDD.n902 0.000506553
R20248 VDD.n901 VDD.n900 0.000506553
R20249 VDD.n1004 VDD.n987 0.000506553
R20250 VDD.n191 VDD.n43 0.000506553
R20251 VDD.n190 VDD.n40 0.000506553
R20252 VDD.n189 VDD.n188 0.000506553
R20253 VDD.n108 VDD.n107 0.000506553
R20254 VDD.n106 VDD.n105 0.000506553
R20255 VDD.n209 VDD.n192 0.000506553
R20256 VDD.n581 VDD.n437 0.000506553
R20257 VDD.n580 VDD.n434 0.000506553
R20258 VDD.n579 VDD.n578 0.000506553
R20259 VDD.n502 VDD.n501 0.000506553
R20260 VDD.n500 VDD.n499 0.000506553
R20261 VDD.n599 VDD.n582 0.000506553
R20262 VDD.n1458 VDD.n1457 0.000506553
R20263 VDD.n1508 VDD.n1507 0.000506553
R20264 VDD.n1456 VDD.n1455 0.000506553
R20265 VDD.n1430 VDD.n1429 0.000506553
R20266 VDD.n1398 VDD.n1397 0.000506553
R20267 VDD.n1373 VDD.n1372 0.000506553
R20268 VDD.n1371 VDD.n1370 0.000506553
R20269 VDD.n1428 VDD.n1427 0.000506553
R20270 VDD.n1726 VDD.n1725 0.000505865
R20271 VDD.n2075 VDD.n2074 0.000505865
R20272 VDD.n2305 VDD.n2304 0.000505865
R20273 VDD.n2563 VDD.n2562 0.000505865
R20274 VDD.n2821 VDD.n2820 0.000505865
R20275 VDD.n3079 VDD.n3078 0.000505865
R20276 VDD.n3337 VDD.n3336 0.000505865
R20277 VDD.n5667 VDD.n5666 0.000505865
R20278 VDD.n5413 VDD.n5412 0.000505865
R20279 VDD.n3595 VDD.n3594 0.000505865
R20280 VDD.n3853 VDD.n3852 0.000505865
R20281 VDD.n4111 VDD.n4110 0.000505865
R20282 VDD.n4369 VDD.n4368 0.000505865
R20283 VDD.n4627 VDD.n4626 0.000505865
R20284 VDD.n4885 VDD.n4884 0.000505865
R20285 VDD.n5177 VDD.n5176 0.000505865
R20286 VDD.n1839 VDD.n1838 0.000504381
R20287 VDD.n2160 VDD.n2159 0.000504381
R20288 VDD.n2418 VDD.n2417 0.000504381
R20289 VDD.n2676 VDD.n2675 0.000504381
R20290 VDD.n2934 VDD.n2933 0.000504381
R20291 VDD.n3192 VDD.n3191 0.000504381
R20292 VDD.n3450 VDD.n3449 0.000504381
R20293 VDD.n5777 VDD.n5776 0.000504381
R20294 VDD.n5523 VDD.n5522 0.000504381
R20295 VDD.n3708 VDD.n3707 0.000504381
R20296 VDD.n3966 VDD.n3965 0.000504381
R20297 VDD.n4224 VDD.n4223 0.000504381
R20298 VDD.n4482 VDD.n4481 0.000504381
R20299 VDD.n4740 VDD.n4739 0.000504381
R20300 VDD.n5001 VDD.n5000 0.000504381
R20301 VDD.n5263 VDD.n5262 0.000504381
R20302 VDD.n1719 VDD.n1671 0.000503792
R20303 VDD.n2068 VDD.n2020 0.000503792
R20304 VDD.n2298 VDD.n2250 0.000503792
R20305 VDD.n2556 VDD.n2508 0.000503792
R20306 VDD.n2814 VDD.n2766 0.000503792
R20307 VDD.n3072 VDD.n3024 0.000503792
R20308 VDD.n3330 VDD.n3282 0.000503792
R20309 VDD.n5660 VDD.n5612 0.000503792
R20310 VDD.n5406 VDD.n5358 0.000503792
R20311 VDD.n3588 VDD.n3540 0.000503792
R20312 VDD.n3846 VDD.n3798 0.000503792
R20313 VDD.n4104 VDD.n4056 0.000503792
R20314 VDD.n4362 VDD.n4314 0.000503792
R20315 VDD.n4620 VDD.n4572 0.000503792
R20316 VDD.n4878 VDD.n4830 0.000503792
R20317 VDD.n5170 VDD.n5122 0.000503792
R20318 VDD.n1427 VDD.n1426 0.000503441
R20319 VDD.n1399 VDD.n1398 0.000503441
R20320 VDD.n1370 VDD.n1369 0.000503441
R20321 VDD.n1459 VDD.n1458 0.000503441
R20322 VDD.n1509 VDD.n1508 0.000503441
R20323 VDD.n1345 VDD.n1344 0.000501258
R20324 VDD.n1319 VDD.n1318 0.000501258
R20325 VDD.n1401 VDD.n1400 0.000501258
R20326 VDD.n1361 VDD.n1360 0.000501258
R20327 VDD.n1289 VDD.n1288 0.000501258
R20328 VDD.n1506 VDD.n1505 0.000501258
R20329 VDD.n1818 VDD.n1817 0.000501164
R20330 VDD.n2139 VDD.n2138 0.000501164
R20331 VDD.n2397 VDD.n2396 0.000501164
R20332 VDD.n2655 VDD.n2654 0.000501164
R20333 VDD.n2913 VDD.n2912 0.000501164
R20334 VDD.n3171 VDD.n3170 0.000501164
R20335 VDD.n3429 VDD.n3428 0.000501164
R20336 VDD.n5756 VDD.n5755 0.000501164
R20337 VDD.n5502 VDD.n5501 0.000501164
R20338 VDD.n3687 VDD.n3686 0.000501164
R20339 VDD.n3945 VDD.n3944 0.000501164
R20340 VDD.n4203 VDD.n4202 0.000501164
R20341 VDD.n4461 VDD.n4460 0.000501164
R20342 VDD.n4719 VDD.n4718 0.000501164
R20343 VDD.n4980 VDD.n4979 0.000501164
R20344 VDD.n5242 VDD.n5241 0.000501164
R20345 VDD.n1053 VDD.n838 0.00050097
R20346 VDD.n1098 VDD.n835 0.00050097
R20347 VDD.n983 VDD.n982 0.00050097
R20348 VDD.n900 VDD.n899 0.00050097
R20349 VDD.n258 VDD.n43 0.00050097
R20350 VDD.n303 VDD.n40 0.00050097
R20351 VDD.n188 VDD.n187 0.00050097
R20352 VDD.n105 VDD.n104 0.00050097
R20353 VDD.n648 VDD.n437 0.00050097
R20354 VDD.n693 VDD.n434 0.00050097
R20355 VDD.n578 VDD.n577 0.00050097
R20356 VDD.n499 VDD.n498 0.00050097
R20357 VDD.n1004 VDD.n1003 0.00050097
R20358 VDD.n209 VDD.n208 0.00050097
R20359 VDD.n599 VDD.n598 0.00050097
R20360 VDD.n2193 VDD.n2192 0.000500414
R20361 VDD.n2451 VDD.n2450 0.000500414
R20362 VDD.n2709 VDD.n2708 0.000500414
R20363 VDD.n2967 VDD.n2966 0.000500414
R20364 VDD.n3225 VDD.n3224 0.000500414
R20365 VDD.n3483 VDD.n3482 0.000500414
R20366 VDD.n5810 VDD.n5809 0.000500414
R20367 VDD.n5556 VDD.n5555 0.000500414
R20368 VDD.n3741 VDD.n3740 0.000500414
R20369 VDD.n3999 VDD.n3998 0.000500414
R20370 VDD.n4257 VDD.n4256 0.000500414
R20371 VDD.n4515 VDD.n4514 0.000500414
R20372 VDD.n4773 VDD.n4772 0.000500414
R20373 VDD.n5034 VDD.n5033 0.000500414
R20374 VDD.n5296 VDD.n5295 0.000500414
R20375 VDD.n1872 VDD.n1871 0.000500414
R20376 VDD.n1180 VDD.n1179 0.000500259
R20377 VDD.n1920 VDD.n1919 0.000500184
R20378 VDD.n2241 VDD.n2240 0.000500184
R20379 VDD.n2499 VDD.n2498 0.000500184
R20380 VDD.n2757 VDD.n2756 0.000500184
R20381 VDD.n3015 VDD.n3014 0.000500184
R20382 VDD.n3273 VDD.n3272 0.000500184
R20383 VDD.n3531 VDD.n3530 0.000500184
R20384 VDD.n3789 VDD.n3788 0.000500184
R20385 VDD.n4047 VDD.n4046 0.000500184
R20386 VDD.n4305 VDD.n4304 0.000500184
R20387 VDD.n4563 VDD.n4562 0.000500184
R20388 VDD.n4821 VDD.n4820 0.000500184
R20389 VDD.n1775 VDD.n1774 0.000500121
R20390 VDD.n2124 VDD.n2123 0.000500121
R20391 VDD.n2354 VDD.n2353 0.000500121
R20392 VDD.n2612 VDD.n2611 0.000500121
R20393 VDD.n2870 VDD.n2869 0.000500121
R20394 VDD.n3128 VDD.n3127 0.000500121
R20395 VDD.n3386 VDD.n3385 0.000500121
R20396 VDD.n3644 VDD.n3643 0.000500121
R20397 VDD.n3902 VDD.n3901 0.000500121
R20398 VDD.n4160 VDD.n4159 0.000500121
R20399 VDD.n4418 VDD.n4417 0.000500121
R20400 VDD.n4676 VDD.n4675 0.000500121
R20401 VDD.n2162 VDD.n1983 0.000500117
R20402 VDD.n2420 VDD.n2243 0.000500117
R20403 VDD.n2678 VDD.n2501 0.000500117
R20404 VDD.n2936 VDD.n2759 0.000500117
R20405 VDD.n3194 VDD.n3017 0.000500117
R20406 VDD.n3452 VDD.n3275 0.000500117
R20407 VDD.n5779 VDD.n5716 0.000500117
R20408 VDD.n5525 VDD.n5462 0.000500117
R20409 VDD.n3710 VDD.n3533 0.000500117
R20410 VDD.n3968 VDD.n3791 0.000500117
R20411 VDD.n4226 VDD.n4049 0.000500117
R20412 VDD.n4484 VDD.n4307 0.000500117
R20413 VDD.n4742 VDD.n4565 0.000500117
R20414 VDD.n1841 VDD.n1664 0.000500117
R20415 VDD.n5003 VDD.n4823 0.000500117
R20416 VDD.n5265 VDD.n5084 0.000500117
R20417 VDD.n5229 VDD.n5228 0.000500084
R20418 VDD.n1602 VDD.n1246 0.000500071
R20419 VDD.n1601 VDD.n1540 0.000500071
R20420 OUT3.n142 OUT3.n140 145.809
R20421 OUT3.n91 OUT3.n89 145.809
R20422 OUT3.n53 OUT3.n51 145.809
R20423 OUT3.n7 OUT3.n5 145.809
R20424 OUT3.n91 OUT3.n90 107.409
R20425 OUT3.n93 OUT3.n92 107.409
R20426 OUT3.n95 OUT3.n94 107.409
R20427 OUT3.n97 OUT3.n96 107.409
R20428 OUT3.n99 OUT3.n98 107.409
R20429 OUT3.n101 OUT3.n100 107.409
R20430 OUT3.n53 OUT3.n52 107.409
R20431 OUT3.n55 OUT3.n54 107.409
R20432 OUT3.n57 OUT3.n56 107.409
R20433 OUT3.n59 OUT3.n58 107.409
R20434 OUT3.n61 OUT3.n60 107.409
R20435 OUT3.n63 OUT3.n62 107.409
R20436 OUT3.n7 OUT3.n6 107.409
R20437 OUT3.n9 OUT3.n8 107.409
R20438 OUT3.n11 OUT3.n10 107.409
R20439 OUT3.n13 OUT3.n12 107.409
R20440 OUT3.n15 OUT3.n14 107.409
R20441 OUT3.n17 OUT3.n16 107.409
R20442 OUT3.n142 OUT3.n141 107.407
R20443 OUT3.n144 OUT3.n143 107.407
R20444 OUT3.n146 OUT3.n145 107.407
R20445 OUT3.n148 OUT3.n147 107.407
R20446 OUT3.n150 OUT3.n149 107.407
R20447 OUT3.n152 OUT3.n151 107.407
R20448 OUT3.n160 OUT3.n158 87.1779
R20449 OUT3.n114 OUT3.n112 87.1779
R20450 OUT3.n72 OUT3.n70 87.1779
R20451 OUT3.n26 OUT3.n24 87.1779
R20452 OUT3.n160 OUT3.n159 52.82
R20453 OUT3.n162 OUT3.n161 52.82
R20454 OUT3.n164 OUT3.n163 52.82
R20455 OUT3.n166 OUT3.n165 52.82
R20456 OUT3.n168 OUT3.n167 52.82
R20457 OUT3.n170 OUT3.n169 52.82
R20458 OUT3.n114 OUT3.n113 52.82
R20459 OUT3.n116 OUT3.n115 52.82
R20460 OUT3.n118 OUT3.n117 52.82
R20461 OUT3.n120 OUT3.n119 52.82
R20462 OUT3.n122 OUT3.n121 52.82
R20463 OUT3.n124 OUT3.n123 52.82
R20464 OUT3.n72 OUT3.n71 52.82
R20465 OUT3.n74 OUT3.n73 52.82
R20466 OUT3.n76 OUT3.n75 52.82
R20467 OUT3.n78 OUT3.n77 52.82
R20468 OUT3.n80 OUT3.n79 52.82
R20469 OUT3.n82 OUT3.n81 52.82
R20470 OUT3.n26 OUT3.n25 52.82
R20471 OUT3.n28 OUT3.n27 52.82
R20472 OUT3.n30 OUT3.n29 52.82
R20473 OUT3.n32 OUT3.n31 52.82
R20474 OUT3.n34 OUT3.n33 52.82
R20475 OUT3.n36 OUT3.n35 52.82
R20476 OUT3.n144 OUT3.n142 38.4005
R20477 OUT3.n146 OUT3.n144 38.4005
R20478 OUT3.n148 OUT3.n146 38.4005
R20479 OUT3.n150 OUT3.n148 38.4005
R20480 OUT3.n152 OUT3.n150 38.4005
R20481 OUT3.n153 OUT3.n152 38.4005
R20482 OUT3.n93 OUT3.n91 38.4005
R20483 OUT3.n95 OUT3.n93 38.4005
R20484 OUT3.n97 OUT3.n95 38.4005
R20485 OUT3.n99 OUT3.n97 38.4005
R20486 OUT3.n101 OUT3.n99 38.4005
R20487 OUT3.n102 OUT3.n101 38.4005
R20488 OUT3.n55 OUT3.n53 38.4005
R20489 OUT3.n57 OUT3.n55 38.4005
R20490 OUT3.n59 OUT3.n57 38.4005
R20491 OUT3.n61 OUT3.n59 38.4005
R20492 OUT3.n63 OUT3.n61 38.4005
R20493 OUT3.n64 OUT3.n63 38.4005
R20494 OUT3.n9 OUT3.n7 38.4005
R20495 OUT3.n11 OUT3.n9 38.4005
R20496 OUT3.n13 OUT3.n11 38.4005
R20497 OUT3.n15 OUT3.n13 38.4005
R20498 OUT3.n17 OUT3.n15 38.4005
R20499 OUT3.n18 OUT3.n17 38.4005
R20500 OUT3.n162 OUT3.n160 34.3584
R20501 OUT3.n164 OUT3.n162 34.3584
R20502 OUT3.n166 OUT3.n164 34.3584
R20503 OUT3.n168 OUT3.n166 34.3584
R20504 OUT3.n170 OUT3.n168 34.3584
R20505 OUT3.n174 OUT3.n170 34.3584
R20506 OUT3.n116 OUT3.n114 34.3584
R20507 OUT3.n118 OUT3.n116 34.3584
R20508 OUT3.n120 OUT3.n118 34.3584
R20509 OUT3.n122 OUT3.n120 34.3584
R20510 OUT3.n124 OUT3.n122 34.3584
R20511 OUT3.n129 OUT3.n124 34.3584
R20512 OUT3.n74 OUT3.n72 34.3584
R20513 OUT3.n76 OUT3.n74 34.3584
R20514 OUT3.n78 OUT3.n76 34.3584
R20515 OUT3.n80 OUT3.n78 34.3584
R20516 OUT3.n82 OUT3.n80 34.3584
R20517 OUT3.n83 OUT3.n82 34.3584
R20518 OUT3.n28 OUT3.n26 34.3584
R20519 OUT3.n30 OUT3.n28 34.3584
R20520 OUT3.n32 OUT3.n30 34.3584
R20521 OUT3.n34 OUT3.n32 34.3584
R20522 OUT3.n36 OUT3.n34 34.3584
R20523 OUT3.n40 OUT3.n36 34.3584
R20524 OUT3.n135 OUT3.t75 26.5955
R20525 OUT3.n135 OUT3.t101 26.5955
R20526 OUT3.n140 OUT3.t85 26.5955
R20527 OUT3.n140 OUT3.t124 26.5955
R20528 OUT3.n141 OUT3.t99 26.5955
R20529 OUT3.n141 OUT3.t72 26.5955
R20530 OUT3.n143 OUT3.t70 26.5955
R20531 OUT3.n143 OUT3.t83 26.5955
R20532 OUT3.n145 OUT3.t91 26.5955
R20533 OUT3.n145 OUT3.t107 26.5955
R20534 OUT3.n147 OUT3.t105 26.5955
R20535 OUT3.n147 OUT3.t127 26.5955
R20536 OUT3.n149 OUT3.t125 26.5955
R20537 OUT3.n149 OUT3.t89 26.5955
R20538 OUT3.n151 OUT3.t116 26.5955
R20539 OUT3.n151 OUT3.t77 26.5955
R20540 OUT3.n89 OUT3.t86 26.5955
R20541 OUT3.n89 OUT3.t112 26.5955
R20542 OUT3.n90 OUT3.t110 26.5955
R20543 OUT3.n90 OUT3.t73 26.5955
R20544 OUT3.n92 OUT3.t64 26.5955
R20545 OUT3.n92 OUT3.t94 26.5955
R20546 OUT3.n94 OUT3.t65 26.5955
R20547 OUT3.n94 OUT3.t81 26.5955
R20548 OUT3.n96 OUT3.t79 26.5955
R20549 OUT3.n96 OUT3.t97 26.5955
R20550 OUT3.n98 OUT3.t104 26.5955
R20551 OUT3.n98 OUT3.t118 26.5955
R20552 OUT3.n100 OUT3.t123 26.5955
R20553 OUT3.n100 OUT3.t88 26.5955
R20554 OUT3.n51 OUT3.t68 26.5955
R20555 OUT3.n51 OUT3.t113 26.5955
R20556 OUT3.n52 OUT3.t84 26.5955
R20557 OUT3.n52 OUT3.t100 26.5955
R20558 OUT3.n54 OUT3.t108 26.5955
R20559 OUT3.n54 OUT3.t71 26.5955
R20560 OUT3.n56 OUT3.t120 26.5955
R20561 OUT3.n56 OUT3.t82 26.5955
R20562 OUT3.n58 OUT3.t90 26.5955
R20563 OUT3.n58 OUT3.t106 26.5955
R20564 OUT3.n60 OUT3.t114 26.5955
R20565 OUT3.n60 OUT3.t126 26.5955
R20566 OUT3.n62 OUT3.t93 26.5955
R20567 OUT3.n62 OUT3.t69 26.5955
R20568 OUT3.n1 OUT3.t122 26.5955
R20569 OUT3.n1 OUT3.t67 26.5955
R20570 OUT3.n5 OUT3.t74 26.5955
R20571 OUT3.n5 OUT3.t87 26.5955
R20572 OUT3.n6 OUT3.t95 26.5955
R20573 OUT3.n6 OUT3.t111 26.5955
R20574 OUT3.n8 OUT3.t109 26.5955
R20575 OUT3.n8 OUT3.t121 26.5955
R20576 OUT3.n10 OUT3.t98 26.5955
R20577 OUT3.n10 OUT3.t92 26.5955
R20578 OUT3.n12 OUT3.t119 26.5955
R20579 OUT3.n12 OUT3.t80 26.5955
R20580 OUT3.n14 OUT3.t78 26.5955
R20581 OUT3.n14 OUT3.t96 26.5955
R20582 OUT3.n16 OUT3.t103 26.5955
R20583 OUT3.n16 OUT3.t117 26.5955
R20584 OUT3.n46 OUT3.t115 25.6105
R20585 OUT3.n171 OUT3.t27 24.9236
R20586 OUT3.n171 OUT3.t53 24.9236
R20587 OUT3.n158 OUT3.t37 24.9236
R20588 OUT3.n158 OUT3.t12 24.9236
R20589 OUT3.n159 OUT3.t51 24.9236
R20590 OUT3.n159 OUT3.t24 24.9236
R20591 OUT3.n161 OUT3.t22 24.9236
R20592 OUT3.n161 OUT3.t35 24.9236
R20593 OUT3.n163 OUT3.t43 24.9236
R20594 OUT3.n163 OUT3.t59 24.9236
R20595 OUT3.n165 OUT3.t57 24.9236
R20596 OUT3.n165 OUT3.t15 24.9236
R20597 OUT3.n167 OUT3.t13 24.9236
R20598 OUT3.n167 OUT3.t41 24.9236
R20599 OUT3.n169 OUT3.t4 24.9236
R20600 OUT3.n169 OUT3.t29 24.9236
R20601 OUT3.n112 OUT3.t38 24.9236
R20602 OUT3.n112 OUT3.t0 24.9236
R20603 OUT3.n113 OUT3.t62 24.9236
R20604 OUT3.n113 OUT3.t25 24.9236
R20605 OUT3.n115 OUT3.t16 24.9236
R20606 OUT3.n115 OUT3.t46 24.9236
R20607 OUT3.n117 OUT3.t17 24.9236
R20608 OUT3.n117 OUT3.t33 24.9236
R20609 OUT3.n119 OUT3.t31 24.9236
R20610 OUT3.n119 OUT3.t49 24.9236
R20611 OUT3.n121 OUT3.t56 24.9236
R20612 OUT3.n121 OUT3.t6 24.9236
R20613 OUT3.n123 OUT3.t11 24.9236
R20614 OUT3.n123 OUT3.t40 24.9236
R20615 OUT3.n70 OUT3.t20 24.9236
R20616 OUT3.n70 OUT3.t1 24.9236
R20617 OUT3.n71 OUT3.t36 24.9236
R20618 OUT3.n71 OUT3.t52 24.9236
R20619 OUT3.n73 OUT3.t60 24.9236
R20620 OUT3.n73 OUT3.t23 24.9236
R20621 OUT3.n75 OUT3.t8 24.9236
R20622 OUT3.n75 OUT3.t34 24.9236
R20623 OUT3.n77 OUT3.t42 24.9236
R20624 OUT3.n77 OUT3.t58 24.9236
R20625 OUT3.n79 OUT3.t2 24.9236
R20626 OUT3.n79 OUT3.t14 24.9236
R20627 OUT3.n81 OUT3.t45 24.9236
R20628 OUT3.n81 OUT3.t21 24.9236
R20629 OUT3.n37 OUT3.t10 24.9236
R20630 OUT3.n37 OUT3.t19 24.9236
R20631 OUT3.n24 OUT3.t26 24.9236
R20632 OUT3.n24 OUT3.t39 24.9236
R20633 OUT3.n25 OUT3.t47 24.9236
R20634 OUT3.n25 OUT3.t63 24.9236
R20635 OUT3.n27 OUT3.t61 24.9236
R20636 OUT3.n27 OUT3.t9 24.9236
R20637 OUT3.n29 OUT3.t50 24.9236
R20638 OUT3.n29 OUT3.t44 24.9236
R20639 OUT3.n31 OUT3.t7 24.9236
R20640 OUT3.n31 OUT3.t32 24.9236
R20641 OUT3.n33 OUT3.t30 24.9236
R20642 OUT3.n33 OUT3.t48 24.9236
R20643 OUT3.n35 OUT3.t55 24.9236
R20644 OUT3.n35 OUT3.t5 24.9236
R20645 OUT3.n68 OUT3.t3 24.7196
R20646 OUT3.n105 OUT3.t66 24.6255
R20647 OUT3.n68 OUT3.t28 23.9564
R20648 OUT3.n127 OUT3.t18 23.1655
R20649 OUT3.n103 OUT3.t102 19.1164
R20650 OUT3.n126 OUT3.n125 13.8467
R20651 OUT3 OUT3.n174 11.4429
R20652 OUT3 OUT3.n129 11.4429
R20653 OUT3 OUT3.n83 11.4429
R20654 OUT3 OUT3.n40 11.4429
R20655 OUT3.n125 OUT3.t54 11.0774
R20656 OUT3.n47 OUT3.t76 10.8355
R20657 OUT3.n106 OUT3.n105 9.3005
R20658 OUT3.n110 OUT3.n109 9.3005
R20659 OUT3.n128 OUT3.n127 8.77252
R20660 OUT3.n136 OUT3.n135 8.76605
R20661 OUT3.n2 OUT3.n1 8.76605
R20662 OUT3.n50 OUT3.n49 8.70762
R20663 OUT3.n49 OUT3.n48 8.69892
R20664 OUT3.n172 OUT3.n171 7.87147
R20665 OUT3.n38 OUT3.n37 7.87147
R20666 OUT3.n48 OUT3.n47 7.77627
R20667 OUT3.n104 OUT3.n103 7.29637
R20668 OUT3.n69 OUT3.n68 6.88889
R20669 OUT3.n85 OUT3.n69 4.758
R20670 OUT3.n128 OUT3.n111 4.6505
R20671 OUT3.n107 OUT3.n106 4.6505
R20672 OUT3.n39 OUT3.n23 4.6505
R20673 OUT3.n20 OUT3.n19 4.6505
R20674 OUT3.n3 OUT3.n2 4.26717
R20675 OUT3.n175 OUT3 3.10353
R20676 OUT3.n130 OUT3 3.10353
R20677 OUT3.n84 OUT3 3.10353
R20678 OUT3.n41 OUT3 3.10353
R20679 OUT3.n173 OUT3.n157 3.1005
R20680 OUT3.n137 OUT3.n136 3.1005
R20681 OUT3.n155 OUT3.n154 3.1005
R20682 OUT3.n66 OUT3.n65 2.75
R20683 OUT3.n154 OUT3.n153 2.71565
R20684 OUT3.n106 OUT3.n102 2.71565
R20685 OUT3.n65 OUT3.n64 2.71565
R20686 OUT3.n19 OUT3.n18 2.71565
R20687 OUT3.n66 OUT3.n50 2.69896
R20688 OUT3.n105 OUT3.n104 1.9705
R20689 OUT3.n174 OUT3 1.74595
R20690 OUT3 OUT3.n173 1.74595
R20691 OUT3.n129 OUT3 1.74595
R20692 OUT3 OUT3.n128 1.74595
R20693 OUT3.n83 OUT3 1.74595
R20694 OUT3.n40 OUT3 1.74595
R20695 OUT3 OUT3.n39 1.74595
R20696 OUT3.n127 OUT3.n126 1.74224
R20697 OUT3.n181 OUT3.n180 0.810582
R20698 OUT3 OUT3.n183 0.597838
R20699 OUT3.n183 OUT3.n182 0.531962
R20700 OUT3.n182 OUT3.n181 0.531962
R20701 OUT3.n182 OUT3.n86 0.475506
R20702 OUT3 OUT3.n69 0.388379
R20703 OUT3.n173 OUT3.n172 0.300854
R20704 OUT3.n39 OUT3.n38 0.300854
R20705 OUT3.n183 OUT3.n45 0.275505
R20706 OUT3.n181 OUT3.n134 0.263005
R20707 OUT3.n180 OUT3.n179 0.1755
R20708 OUT3.n134 OUT3.n133 0.1755
R20709 OUT3.n45 OUT3.n44 0.1755
R20710 OUT3.n176 OUT3.n157 0.11675
R20711 OUT3.n131 OUT3.n111 0.11675
R20712 OUT3.n42 OUT3.n23 0.11675
R20713 OUT3.n132 OUT3.n107 0.10425
R20714 OUT3.n178 OUT3.n155 0.09175
R20715 OUT3.n43 OUT3.n20 0.09175
R20716 OUT3.n86 OUT3.n66 0.0855244
R20717 OUT3.n49 OUT3.n46 0.0578287
R20718 OUT3.n86 OUT3.n85 0.0505
R20719 OUT3.n155 OUT3.n139 0.04425
R20720 OUT3.n20 OUT3.n4 0.04425
R20721 OUT3.n107 OUT3.n88 0.043
R20722 OUT3.n111 OUT3.n110 0.03175
R20723 OUT3.n139 OUT3.n137 0.028
R20724 OUT3.n4 OUT3.n0 0.028
R20725 OUT3.n178 OUT3.n176 0.0255
R20726 OUT3.n157 OUT3.n156 0.0255
R20727 OUT3.n43 OUT3.n42 0.0255
R20728 OUT3.n23 OUT3.n22 0.0255
R20729 OUT3.n132 OUT3.n131 0.013
R20730 OUT3.n88 OUT3.n87 0.00450862
R20731 OUT3.n139 OUT3.n138 0.0025557
R20732 OUT3.n4 OUT3.n3 0.0025557
R20733 OUT3.n176 OUT3.n175 0.00053521
R20734 OUT3.n131 OUT3.n130 0.00053521
R20735 OUT3.n85 OUT3.n84 0.00053521
R20736 OUT3.n42 OUT3.n41 0.00053521
R20737 OUT3.n178 OUT3.n177 0.00050852
R20738 OUT3.n132 OUT3.n108 0.00050852
R20739 OUT3.n86 OUT3.n67 0.00050852
R20740 OUT3.n43 OUT3.n21 0.00050852
R20741 OUT3.n179 OUT3.n178 0.000500999
R20742 OUT3.n133 OUT3.n132 0.000500999
R20743 OUT3.n44 OUT3.n43 0.000500999
R20744 R0.n0 R0.t4 260.322
R20745 R0.n5 R0.t5 233.888
R20746 R0.n0 R0.t6 175.169
R20747 R0.n4 R0.t7 159.725
R20748 R0.n6 R0.t1 17.4109
R20749 R0.n1 R0.n0 9.75129
R20750 R0.n6 R0.t0 9.6037
R20751 R0.n2 R0 9.3005
R20752 R0.n8 R0.t2 8.40929
R20753 R0.n4 R0.t3 8.06629
R20754 R0 R0.n1 3.11453
R20755 R0.n5 R0.n4 1.73501
R20756 R0.n7 R0.n5 0.99025
R20757 R0.n8 R0.n7 0.853186
R20758 R0 R0.n9 0.315016
R20759 R0.n3 R0 0.310984
R20760 R0.n3 R0.n2 0.195812
R20761 R0.n8 R0 0.109296
R20762 R0 R0.n3 0.0776605
R20763 R0.n2 R0.n1 0.0292043
R20764 R0.n9 R0.n8 0.0120741
R20765 R0.n9 R0 0.00654839
R20766 R0.n9 R0 0.00281481
R20767 R0.n7 R0.n6 0.000500726
R20768 OUT0.n122 OUT0.n120 145.809
R20769 OUT0.n65 OUT0.n63 145.809
R20770 OUT0.n25 OUT0.n23 145.809
R20771 OUT0.n102 OUT0.n100 145.808
R20772 OUT0.n65 OUT0.n64 107.409
R20773 OUT0.n67 OUT0.n66 107.409
R20774 OUT0.n69 OUT0.n68 107.409
R20775 OUT0.n71 OUT0.n70 107.409
R20776 OUT0.n73 OUT0.n72 107.409
R20777 OUT0.n75 OUT0.n74 107.409
R20778 OUT0.n25 OUT0.n24 107.409
R20779 OUT0.n27 OUT0.n26 107.409
R20780 OUT0.n29 OUT0.n28 107.409
R20781 OUT0.n31 OUT0.n30 107.409
R20782 OUT0.n33 OUT0.n32 107.409
R20783 OUT0.n35 OUT0.n34 107.409
R20784 OUT0.n122 OUT0.n121 107.407
R20785 OUT0.n124 OUT0.n123 107.407
R20786 OUT0.n126 OUT0.n125 107.407
R20787 OUT0.n128 OUT0.n127 107.407
R20788 OUT0.n130 OUT0.n129 107.407
R20789 OUT0.n132 OUT0.n131 107.407
R20790 OUT0.n102 OUT0.n101 107.407
R20791 OUT0.n104 OUT0.n103 107.407
R20792 OUT0.n106 OUT0.n105 107.407
R20793 OUT0.n108 OUT0.n107 107.407
R20794 OUT0.n110 OUT0.n109 107.407
R20795 OUT0.n112 OUT0.n111 107.407
R20796 OUT0.n138 OUT0.n136 87.1779
R20797 OUT0.n83 OUT0.n81 87.1779
R20798 OUT0.n44 OUT0.n42 87.1779
R20799 OUT0.n4 OUT0.n2 87.1779
R20800 OUT0.n54 OUT0.n53 52.82
R20801 OUT0.n14 OUT0.n13 52.82
R20802 OUT0.n138 OUT0.n137 52.82
R20803 OUT0.n140 OUT0.n139 52.82
R20804 OUT0.n142 OUT0.n141 52.82
R20805 OUT0.n144 OUT0.n143 52.82
R20806 OUT0.n146 OUT0.n145 52.82
R20807 OUT0.n148 OUT0.n147 52.82
R20808 OUT0.n83 OUT0.n82 52.82
R20809 OUT0.n85 OUT0.n84 52.82
R20810 OUT0.n87 OUT0.n86 52.82
R20811 OUT0.n89 OUT0.n88 52.82
R20812 OUT0.n91 OUT0.n90 52.82
R20813 OUT0.n93 OUT0.n92 52.82
R20814 OUT0.n44 OUT0.n43 52.82
R20815 OUT0.n46 OUT0.n45 52.82
R20816 OUT0.n48 OUT0.n47 52.82
R20817 OUT0.n50 OUT0.n49 52.82
R20818 OUT0.n52 OUT0.n51 52.82
R20819 OUT0.n4 OUT0.n3 52.82
R20820 OUT0.n6 OUT0.n5 52.82
R20821 OUT0.n8 OUT0.n7 52.82
R20822 OUT0.n10 OUT0.n9 52.82
R20823 OUT0.n12 OUT0.n11 52.82
R20824 OUT0 OUT0.n149 51.0745
R20825 OUT0 OUT0.n94 51.0745
R20826 OUT0.n124 OUT0.n122 38.4005
R20827 OUT0.n126 OUT0.n124 38.4005
R20828 OUT0.n128 OUT0.n126 38.4005
R20829 OUT0.n130 OUT0.n128 38.4005
R20830 OUT0.n132 OUT0.n130 38.4005
R20831 OUT0.n133 OUT0.n132 38.4005
R20832 OUT0.n104 OUT0.n102 38.4005
R20833 OUT0.n106 OUT0.n104 38.4005
R20834 OUT0.n108 OUT0.n106 38.4005
R20835 OUT0.n110 OUT0.n108 38.4005
R20836 OUT0.n112 OUT0.n110 38.4005
R20837 OUT0.n113 OUT0.n112 38.4005
R20838 OUT0.n67 OUT0.n65 38.4005
R20839 OUT0.n69 OUT0.n67 38.4005
R20840 OUT0.n71 OUT0.n69 38.4005
R20841 OUT0.n73 OUT0.n71 38.4005
R20842 OUT0.n75 OUT0.n73 38.4005
R20843 OUT0.n76 OUT0.n75 38.4005
R20844 OUT0.n27 OUT0.n25 38.4005
R20845 OUT0.n29 OUT0.n27 38.4005
R20846 OUT0.n31 OUT0.n29 38.4005
R20847 OUT0.n33 OUT0.n31 38.4005
R20848 OUT0.n35 OUT0.n33 38.4005
R20849 OUT0.n36 OUT0.n35 38.4005
R20850 OUT0.n140 OUT0.n138 34.3584
R20851 OUT0.n142 OUT0.n140 34.3584
R20852 OUT0.n144 OUT0.n142 34.3584
R20853 OUT0.n146 OUT0.n144 34.3584
R20854 OUT0.n148 OUT0.n146 34.3584
R20855 OUT0.n150 OUT0.n148 34.3584
R20856 OUT0.n85 OUT0.n83 34.3584
R20857 OUT0.n87 OUT0.n85 34.3584
R20858 OUT0.n89 OUT0.n87 34.3584
R20859 OUT0.n91 OUT0.n89 34.3584
R20860 OUT0.n93 OUT0.n91 34.3584
R20861 OUT0.n95 OUT0.n93 34.3584
R20862 OUT0.n46 OUT0.n44 34.3584
R20863 OUT0.n48 OUT0.n46 34.3584
R20864 OUT0.n50 OUT0.n48 34.3584
R20865 OUT0.n52 OUT0.n50 34.3584
R20866 OUT0.n54 OUT0.n52 34.3584
R20867 OUT0.n58 OUT0.n54 34.3584
R20868 OUT0.n6 OUT0.n4 34.3584
R20869 OUT0.n8 OUT0.n6 34.3584
R20870 OUT0.n10 OUT0.n8 34.3584
R20871 OUT0.n12 OUT0.n10 34.3584
R20872 OUT0.n14 OUT0.n12 34.3584
R20873 OUT0.n18 OUT0.n14 34.3584
R20874 OUT0.n118 OUT0.t105 26.5955
R20875 OUT0.n118 OUT0.t118 26.5955
R20876 OUT0.n120 OUT0.t103 26.5955
R20877 OUT0.n120 OUT0.t75 26.5955
R20878 OUT0.n121 OUT0.t125 26.5955
R20879 OUT0.n121 OUT0.t91 26.5955
R20880 OUT0.n123 OUT0.t70 26.5955
R20881 OUT0.n123 OUT0.t111 26.5955
R20882 OUT0.n125 OUT0.t81 26.5955
R20883 OUT0.n125 OUT0.t99 26.5955
R20884 OUT0.n127 OUT0.t97 26.5955
R20885 OUT0.n127 OUT0.t114 26.5955
R20886 OUT0.n129 OUT0.t120 26.5955
R20887 OUT0.n129 OUT0.t86 26.5955
R20888 OUT0.n131 OUT0.t67 26.5955
R20889 OUT0.n131 OUT0.t107 26.5955
R20890 OUT0.n99 OUT0.t66 26.5955
R20891 OUT0.n99 OUT0.t95 26.5955
R20892 OUT0.n100 OUT0.t85 26.5955
R20893 OUT0.n100 OUT0.t94 26.5955
R20894 OUT0.n101 OUT0.t101 26.5955
R20895 OUT0.n101 OUT0.t74 26.5955
R20896 OUT0.n103 OUT0.t116 26.5955
R20897 OUT0.n103 OUT0.t88 26.5955
R20898 OUT0.n105 OUT0.t87 26.5955
R20899 OUT0.n105 OUT0.t100 26.5955
R20900 OUT0.n107 OUT0.t108 26.5955
R20901 OUT0.n107 OUT0.t122 26.5955
R20902 OUT0.n109 OUT0.t121 26.5955
R20903 OUT0.n109 OUT0.t76 26.5955
R20904 OUT0.n111 OUT0.t110 26.5955
R20905 OUT0.n111 OUT0.t78 26.5955
R20906 OUT0.n62 OUT0.t72 26.5955
R20907 OUT0.n62 OUT0.t106 26.5955
R20908 OUT0.n63 OUT0.t92 26.5955
R20909 OUT0.n63 OUT0.t104 26.5955
R20910 OUT0.n64 OUT0.t102 26.5955
R20911 OUT0.n64 OUT0.t126 26.5955
R20912 OUT0.n66 OUT0.t123 26.5955
R20913 OUT0.n66 OUT0.t89 26.5955
R20914 OUT0.n68 OUT0.t115 26.5955
R20915 OUT0.n68 OUT0.t83 26.5955
R20916 OUT0.n70 OUT0.t79 26.5955
R20917 OUT0.n70 OUT0.t98 26.5955
R20918 OUT0.n72 OUT0.t96 26.5955
R20919 OUT0.n72 OUT0.t113 26.5955
R20920 OUT0.n74 OUT0.t119 26.5955
R20921 OUT0.n74 OUT0.t68 26.5955
R20922 OUT0.n22 OUT0.t71 26.5955
R20923 OUT0.n22 OUT0.t84 26.5955
R20924 OUT0.n23 OUT0.t90 26.5955
R20925 OUT0.n23 OUT0.t112 26.5955
R20926 OUT0.n24 OUT0.t109 26.5955
R20927 OUT0.n24 OUT0.t124 26.5955
R20928 OUT0.n26 OUT0.t65 26.5955
R20929 OUT0.n26 OUT0.t77 26.5955
R20930 OUT0.n28 OUT0.t82 26.5955
R20931 OUT0.n28 OUT0.t117 26.5955
R20932 OUT0.n30 OUT0.t93 26.5955
R20933 OUT0.n30 OUT0.t64 26.5955
R20934 OUT0.n32 OUT0.t69 26.5955
R20935 OUT0.n32 OUT0.t80 26.5955
R20936 OUT0.n34 OUT0.t127 26.5955
R20937 OUT0.n34 OUT0.t73 26.5955
R20938 OUT0.n149 OUT0.t41 24.9236
R20939 OUT0.n149 OUT0.t54 24.9236
R20940 OUT0.n136 OUT0.t39 24.9236
R20941 OUT0.n136 OUT0.t11 24.9236
R20942 OUT0.n137 OUT0.t61 24.9236
R20943 OUT0.n137 OUT0.t27 24.9236
R20944 OUT0.n139 OUT0.t6 24.9236
R20945 OUT0.n139 OUT0.t47 24.9236
R20946 OUT0.n141 OUT0.t17 24.9236
R20947 OUT0.n141 OUT0.t35 24.9236
R20948 OUT0.n143 OUT0.t33 24.9236
R20949 OUT0.n143 OUT0.t50 24.9236
R20950 OUT0.n145 OUT0.t56 24.9236
R20951 OUT0.n145 OUT0.t22 24.9236
R20952 OUT0.n147 OUT0.t3 24.9236
R20953 OUT0.n147 OUT0.t43 24.9236
R20954 OUT0.n94 OUT0.t2 24.9236
R20955 OUT0.n94 OUT0.t31 24.9236
R20956 OUT0.n81 OUT0.t21 24.9236
R20957 OUT0.n81 OUT0.t30 24.9236
R20958 OUT0.n82 OUT0.t37 24.9236
R20959 OUT0.n82 OUT0.t10 24.9236
R20960 OUT0.n84 OUT0.t52 24.9236
R20961 OUT0.n84 OUT0.t24 24.9236
R20962 OUT0.n86 OUT0.t23 24.9236
R20963 OUT0.n86 OUT0.t36 24.9236
R20964 OUT0.n88 OUT0.t44 24.9236
R20965 OUT0.n88 OUT0.t58 24.9236
R20966 OUT0.n90 OUT0.t57 24.9236
R20967 OUT0.n90 OUT0.t12 24.9236
R20968 OUT0.n92 OUT0.t46 24.9236
R20969 OUT0.n92 OUT0.t14 24.9236
R20970 OUT0.n55 OUT0.t8 24.9236
R20971 OUT0.n55 OUT0.t42 24.9236
R20972 OUT0.n42 OUT0.t28 24.9236
R20973 OUT0.n42 OUT0.t40 24.9236
R20974 OUT0.n43 OUT0.t38 24.9236
R20975 OUT0.n43 OUT0.t62 24.9236
R20976 OUT0.n45 OUT0.t59 24.9236
R20977 OUT0.n45 OUT0.t25 24.9236
R20978 OUT0.n47 OUT0.t51 24.9236
R20979 OUT0.n47 OUT0.t19 24.9236
R20980 OUT0.n49 OUT0.t15 24.9236
R20981 OUT0.n49 OUT0.t34 24.9236
R20982 OUT0.n51 OUT0.t32 24.9236
R20983 OUT0.n51 OUT0.t49 24.9236
R20984 OUT0.n53 OUT0.t55 24.9236
R20985 OUT0.n53 OUT0.t4 24.9236
R20986 OUT0.n15 OUT0.t7 24.9236
R20987 OUT0.n15 OUT0.t20 24.9236
R20988 OUT0.n2 OUT0.t26 24.9236
R20989 OUT0.n2 OUT0.t48 24.9236
R20990 OUT0.n3 OUT0.t45 24.9236
R20991 OUT0.n3 OUT0.t60 24.9236
R20992 OUT0.n5 OUT0.t1 24.9236
R20993 OUT0.n5 OUT0.t13 24.9236
R20994 OUT0.n7 OUT0.t18 24.9236
R20995 OUT0.n7 OUT0.t53 24.9236
R20996 OUT0.n9 OUT0.t29 24.9236
R20997 OUT0.n9 OUT0.t0 24.9236
R20998 OUT0.n11 OUT0.t5 24.9236
R20999 OUT0.n11 OUT0.t16 24.9236
R21000 OUT0.n13 OUT0.t63 24.9236
R21001 OUT0.n13 OUT0.t9 24.9236
R21002 OUT0 OUT0.n150 11.4429
R21003 OUT0 OUT0.n95 11.4429
R21004 OUT0 OUT0.n58 11.4429
R21005 OUT0 OUT0.n18 11.4429
R21006 OUT0.n77 OUT0.n62 8.55118
R21007 OUT0.n37 OUT0.n22 8.55118
R21008 OUT0.n114 OUT0.n99 8.55117
R21009 OUT0.n119 OUT0.n118 8.47293
R21010 OUT0.n56 OUT0.n55 7.80093
R21011 OUT0.n16 OUT0.n15 7.80093
R21012 OUT0.n78 OUT0.n77 3.20954
R21013 OUT0.n38 OUT0.n37 3.20953
R21014 OUT0.n115 OUT0.n114 3.20289
R21015 OUT0.n151 OUT0 3.10353
R21016 OUT0.n96 OUT0 3.10353
R21017 OUT0.n59 OUT0 3.10353
R21018 OUT0.n19 OUT0 3.10353
R21019 OUT0.n135 OUT0.n134 3.1005
R21020 OUT0.n57 OUT0.n41 3.1005
R21021 OUT0.n17 OUT0.n1 3.1005
R21022 OUT0.n134 OUT0.n133 2.71565
R21023 OUT0.n114 OUT0.n113 2.13383
R21024 OUT0.n77 OUT0.n76 2.13383
R21025 OUT0.n37 OUT0.n36 2.13383
R21026 OUT0.n150 OUT0 1.74595
R21027 OUT0.n95 OUT0 1.74595
R21028 OUT0.n58 OUT0.n57 1.16414
R21029 OUT0.n18 OUT0.n17 1.16414
R21030 OUT0.n157 OUT0.n156 1.07337
R21031 OUT0.n158 OUT0.n157 0.69375
R21032 OUT0.n159 OUT0.n158 0.68905
R21033 OUT0.n56 OUT0 0.488972
R21034 OUT0.n16 OUT0 0.488972
R21035 OUT0.n158 OUT0.n79 0.414635
R21036 OUT0.n157 OUT0.n116 0.382465
R21037 OUT0.n159 OUT0.n39 0.368576
R21038 OUT0 OUT0.n159 0.281623
R21039 OUT0.n134 OUT0.n119 0.196887
R21040 OUT0.n79 OUT0.n78 0.157252
R21041 OUT0.n39 OUT0.n38 0.139891
R21042 OUT0.n156 OUT0.n155 0.139389
R21043 OUT0.n116 OUT0.n115 0.132946
R21044 OUT0.n60 OUT0.n41 0.113
R21045 OUT0.n20 OUT0.n1 0.113
R21046 OUT0.n154 OUT0.n135 0.101889
R21047 OUT0.n57 OUT0.n56 0.0893205
R21048 OUT0.n17 OUT0.n16 0.0893205
R21049 OUT0.n154 OUT0.n152 0.0282778
R21050 OUT0.n135 OUT0.n117 0.0268889
R21051 OUT0.n98 OUT0.n97 0.0213333
R21052 OUT0.n61 OUT0.n60 0.0143889
R21053 OUT0.n21 OUT0.n20 0.0143889
R21054 OUT0.n115 OUT0.n98 0.00100004
R21055 OUT0.n38 OUT0.n21 0.00100004
R21056 OUT0.n78 OUT0.n61 0.00100004
R21057 OUT0.n152 OUT0.n151 0.000513335
R21058 OUT0.n97 OUT0.n96 0.000513335
R21059 OUT0.n60 OUT0.n59 0.000513218
R21060 OUT0.n20 OUT0.n19 0.000513218
R21061 OUT0.n98 OUT0.n80 0.00050517
R21062 OUT0.n154 OUT0.n153 0.000504838
R21063 OUT0.n61 OUT0.n40 0.000504838
R21064 OUT0.n21 OUT0.n0 0.000504838
R21065 OUT0.n155 OUT0.n154 0.000501713
R21066 I5.t11 I5.t13 618.109
R21067 I5.n12 I5.t6 259.74
R21068 I5 I5.t11 253.56
R21069 I5.n3 I5.t9 228.899
R21070 I5.n18 I5.t7 180.286
R21071 I5.n3 I5.t8 159.411
R21072 I5.n12 I5.t10 157.083
R21073 I5.n20 I5.n19 152
R21074 I5.n26 I5.t5 117.314
R21075 I5.n20 I5.t14 111.091
R21076 I5.n26 I5.t12 110.853
R21077 I5.n18 I5.n17 74.4551
R21078 I5.n24 I5 37.6855
R21079 I5.n28 I5.t1 17.6181
R21080 I5.n29 I5.t4 14.2865
R21081 I5.n31 I5.t3 14.283
R21082 I5.n31 I5.t2 14.283
R21083 I5.n6 I5.n2 9.3005
R21084 I5.n6 I5.n5 9.3005
R21085 I5.n21 I5.n20 9.3005
R21086 I5.n14 I5 9.3005
R21087 I5.n33 I5.t0 8.77744
R21088 I5.n22 I5.n21 7.80966
R21089 I5.n13 I5.n12 7.57248
R21090 I5.n5 I5.n3 7.36978
R21091 I5.n20 I5.n18 6.53562
R21092 I5 I5.n13 4.8645
R21093 I5.n14 I5.n10 4.50988
R21094 I5.n4 I5.n2 3.46717
R21095 I5 I5.n34 3.14231
R21096 I5.n4 I5.n1 3.03286
R21097 I5.n19 I5.n17 2.32777
R21098 I5.n8 I5.n0 2.26553
R21099 I5.n7 I5.n1 2.26468
R21100 I5.n16 I5.n15 2.251
R21101 I5.n22 I5.n16 2.19001
R21102 I5.n19 I5 1.4966
R21103 I5.n23 I5.n9 1.36032
R21104 I5.n33 I5.n32 1.20426
R21105 I5.n23 I5.n22 1.07639
R21106 I5.n5 I5.n4 1.06717
R21107 I5.n2 I5 1.06717
R21108 I5.n9 I5.n8 0.71595
R21109 I5.n35 I5 0.588
R21110 I5 I5.n25 0.577033
R21111 I5.n21 I5.n17 0.499201
R21112 I5 I5.n35 0.441125
R21113 I5.n25 I5.n24 0.435179
R21114 I5.n34 I5.n33 0.32511
R21115 I5.n29 I5.n28 0.314673
R21116 I5.n30 I5.n29 0.299251
R21117 I5.n9 I5 0.221483
R21118 I5.n25 I5 0.20675
R21119 I5.n27 I5.n26 0.159555
R21120 I5.n32 I5.n31 0.106617
R21121 I5.n30 I5.n27 0.0796167
R21122 I5.n32 I5.n30 0.0480595
R21123 I5.n34 I5 0.046937
R21124 I5.n15 I5.n14 0.0301875
R21125 I5.n16 I5.n10 0.0205312
R21126 I5.n35 I5 0.0161667
R21127 I5.n35 I5 0.01225
R21128 I5.n6 I5.n0 0.00618182
R21129 I5.n1 I5.n0 0.00555107
R21130 I5.n7 I5.n6 0.00530477
R21131 I5.n11 I5.n10 0.00210765
R21132 I5.n13 I5.n11 0.00133438
R21133 I5.n8 I5.n7 0.00101192
R21134 I5.n15 I5.n11 0.00100001
R21135 I5.n24 I5.n23 0.000507778
R21136 I5.n28 I5.n27 0.000504658
R21137 OUT2.n122 OUT2.n120 145.809
R21138 OUT2.n65 OUT2.n63 145.809
R21139 OUT2.n25 OUT2.n23 145.809
R21140 OUT2.n102 OUT2.n100 145.808
R21141 OUT2.n65 OUT2.n64 107.409
R21142 OUT2.n67 OUT2.n66 107.409
R21143 OUT2.n69 OUT2.n68 107.409
R21144 OUT2.n71 OUT2.n70 107.409
R21145 OUT2.n73 OUT2.n72 107.409
R21146 OUT2.n75 OUT2.n74 107.409
R21147 OUT2.n25 OUT2.n24 107.409
R21148 OUT2.n27 OUT2.n26 107.409
R21149 OUT2.n29 OUT2.n28 107.409
R21150 OUT2.n31 OUT2.n30 107.409
R21151 OUT2.n33 OUT2.n32 107.409
R21152 OUT2.n35 OUT2.n34 107.409
R21153 OUT2.n122 OUT2.n121 107.407
R21154 OUT2.n124 OUT2.n123 107.407
R21155 OUT2.n126 OUT2.n125 107.407
R21156 OUT2.n128 OUT2.n127 107.407
R21157 OUT2.n130 OUT2.n129 107.407
R21158 OUT2.n132 OUT2.n131 107.407
R21159 OUT2.n102 OUT2.n101 107.407
R21160 OUT2.n104 OUT2.n103 107.407
R21161 OUT2.n106 OUT2.n105 107.407
R21162 OUT2.n108 OUT2.n107 107.407
R21163 OUT2.n110 OUT2.n109 107.407
R21164 OUT2.n112 OUT2.n111 107.407
R21165 OUT2.n138 OUT2.n136 87.1779
R21166 OUT2.n83 OUT2.n81 87.1779
R21167 OUT2.n44 OUT2.n42 87.1779
R21168 OUT2.n4 OUT2.n2 87.1779
R21169 OUT2.n54 OUT2.n53 52.82
R21170 OUT2.n14 OUT2.n13 52.82
R21171 OUT2.n138 OUT2.n137 52.82
R21172 OUT2.n140 OUT2.n139 52.82
R21173 OUT2.n142 OUT2.n141 52.82
R21174 OUT2.n144 OUT2.n143 52.82
R21175 OUT2.n146 OUT2.n145 52.82
R21176 OUT2.n148 OUT2.n147 52.82
R21177 OUT2.n83 OUT2.n82 52.82
R21178 OUT2.n85 OUT2.n84 52.82
R21179 OUT2.n87 OUT2.n86 52.82
R21180 OUT2.n89 OUT2.n88 52.82
R21181 OUT2.n91 OUT2.n90 52.82
R21182 OUT2.n93 OUT2.n92 52.82
R21183 OUT2.n44 OUT2.n43 52.82
R21184 OUT2.n46 OUT2.n45 52.82
R21185 OUT2.n48 OUT2.n47 52.82
R21186 OUT2.n50 OUT2.n49 52.82
R21187 OUT2.n52 OUT2.n51 52.82
R21188 OUT2.n4 OUT2.n3 52.82
R21189 OUT2.n6 OUT2.n5 52.82
R21190 OUT2.n8 OUT2.n7 52.82
R21191 OUT2.n10 OUT2.n9 52.82
R21192 OUT2.n12 OUT2.n11 52.82
R21193 OUT2 OUT2.n149 51.0745
R21194 OUT2 OUT2.n94 51.0745
R21195 OUT2.n124 OUT2.n122 38.4005
R21196 OUT2.n126 OUT2.n124 38.4005
R21197 OUT2.n128 OUT2.n126 38.4005
R21198 OUT2.n130 OUT2.n128 38.4005
R21199 OUT2.n132 OUT2.n130 38.4005
R21200 OUT2.n133 OUT2.n132 38.4005
R21201 OUT2.n104 OUT2.n102 38.4005
R21202 OUT2.n106 OUT2.n104 38.4005
R21203 OUT2.n108 OUT2.n106 38.4005
R21204 OUT2.n110 OUT2.n108 38.4005
R21205 OUT2.n112 OUT2.n110 38.4005
R21206 OUT2.n113 OUT2.n112 38.4005
R21207 OUT2.n67 OUT2.n65 38.4005
R21208 OUT2.n69 OUT2.n67 38.4005
R21209 OUT2.n71 OUT2.n69 38.4005
R21210 OUT2.n73 OUT2.n71 38.4005
R21211 OUT2.n75 OUT2.n73 38.4005
R21212 OUT2.n76 OUT2.n75 38.4005
R21213 OUT2.n27 OUT2.n25 38.4005
R21214 OUT2.n29 OUT2.n27 38.4005
R21215 OUT2.n31 OUT2.n29 38.4005
R21216 OUT2.n33 OUT2.n31 38.4005
R21217 OUT2.n35 OUT2.n33 38.4005
R21218 OUT2.n36 OUT2.n35 38.4005
R21219 OUT2.n140 OUT2.n138 34.3584
R21220 OUT2.n142 OUT2.n140 34.3584
R21221 OUT2.n144 OUT2.n142 34.3584
R21222 OUT2.n146 OUT2.n144 34.3584
R21223 OUT2.n148 OUT2.n146 34.3584
R21224 OUT2.n150 OUT2.n148 34.3584
R21225 OUT2.n85 OUT2.n83 34.3584
R21226 OUT2.n87 OUT2.n85 34.3584
R21227 OUT2.n89 OUT2.n87 34.3584
R21228 OUT2.n91 OUT2.n89 34.3584
R21229 OUT2.n93 OUT2.n91 34.3584
R21230 OUT2.n95 OUT2.n93 34.3584
R21231 OUT2.n46 OUT2.n44 34.3584
R21232 OUT2.n48 OUT2.n46 34.3584
R21233 OUT2.n50 OUT2.n48 34.3584
R21234 OUT2.n52 OUT2.n50 34.3584
R21235 OUT2.n54 OUT2.n52 34.3584
R21236 OUT2.n58 OUT2.n54 34.3584
R21237 OUT2.n6 OUT2.n4 34.3584
R21238 OUT2.n8 OUT2.n6 34.3584
R21239 OUT2.n10 OUT2.n8 34.3584
R21240 OUT2.n12 OUT2.n10 34.3584
R21241 OUT2.n14 OUT2.n12 34.3584
R21242 OUT2.n18 OUT2.n14 34.3584
R21243 OUT2.n118 OUT2.t116 26.5955
R21244 OUT2.n118 OUT2.t65 26.5955
R21245 OUT2.n120 OUT2.t114 26.5955
R21246 OUT2.n120 OUT2.t86 26.5955
R21247 OUT2.n121 OUT2.t72 26.5955
R21248 OUT2.n121 OUT2.t102 26.5955
R21249 OUT2.n123 OUT2.t81 26.5955
R21250 OUT2.n123 OUT2.t122 26.5955
R21251 OUT2.n125 OUT2.t92 26.5955
R21252 OUT2.n125 OUT2.t110 26.5955
R21253 OUT2.n127 OUT2.t108 26.5955
R21254 OUT2.n127 OUT2.t125 26.5955
R21255 OUT2.n129 OUT2.t67 26.5955
R21256 OUT2.n129 OUT2.t97 26.5955
R21257 OUT2.n131 OUT2.t78 26.5955
R21258 OUT2.n131 OUT2.t118 26.5955
R21259 OUT2.n99 OUT2.t77 26.5955
R21260 OUT2.n99 OUT2.t106 26.5955
R21261 OUT2.n100 OUT2.t96 26.5955
R21262 OUT2.n100 OUT2.t105 26.5955
R21263 OUT2.n101 OUT2.t112 26.5955
R21264 OUT2.n101 OUT2.t85 26.5955
R21265 OUT2.n103 OUT2.t127 26.5955
R21266 OUT2.n103 OUT2.t99 26.5955
R21267 OUT2.n105 OUT2.t98 26.5955
R21268 OUT2.n105 OUT2.t111 26.5955
R21269 OUT2.n107 OUT2.t119 26.5955
R21270 OUT2.n107 OUT2.t69 26.5955
R21271 OUT2.n109 OUT2.t68 26.5955
R21272 OUT2.n109 OUT2.t87 26.5955
R21273 OUT2.n111 OUT2.t121 26.5955
R21274 OUT2.n111 OUT2.t89 26.5955
R21275 OUT2.n62 OUT2.t83 26.5955
R21276 OUT2.n62 OUT2.t117 26.5955
R21277 OUT2.n63 OUT2.t103 26.5955
R21278 OUT2.n63 OUT2.t115 26.5955
R21279 OUT2.n64 OUT2.t113 26.5955
R21280 OUT2.n64 OUT2.t73 26.5955
R21281 OUT2.n66 OUT2.t70 26.5955
R21282 OUT2.n66 OUT2.t100 26.5955
R21283 OUT2.n68 OUT2.t126 26.5955
R21284 OUT2.n68 OUT2.t94 26.5955
R21285 OUT2.n70 OUT2.t91 26.5955
R21286 OUT2.n70 OUT2.t109 26.5955
R21287 OUT2.n72 OUT2.t107 26.5955
R21288 OUT2.n72 OUT2.t124 26.5955
R21289 OUT2.n74 OUT2.t66 26.5955
R21290 OUT2.n74 OUT2.t79 26.5955
R21291 OUT2.n22 OUT2.t82 26.5955
R21292 OUT2.n22 OUT2.t95 26.5955
R21293 OUT2.n23 OUT2.t101 26.5955
R21294 OUT2.n23 OUT2.t123 26.5955
R21295 OUT2.n24 OUT2.t120 26.5955
R21296 OUT2.n24 OUT2.t71 26.5955
R21297 OUT2.n26 OUT2.t76 26.5955
R21298 OUT2.n26 OUT2.t88 26.5955
R21299 OUT2.n28 OUT2.t93 26.5955
R21300 OUT2.n28 OUT2.t64 26.5955
R21301 OUT2.n30 OUT2.t104 26.5955
R21302 OUT2.n30 OUT2.t75 26.5955
R21303 OUT2.n32 OUT2.t80 26.5955
R21304 OUT2.n32 OUT2.t90 26.5955
R21305 OUT2.n34 OUT2.t74 26.5955
R21306 OUT2.n34 OUT2.t84 26.5955
R21307 OUT2.n149 OUT2.t6 24.9236
R21308 OUT2.n149 OUT2.t19 24.9236
R21309 OUT2.n136 OUT2.t4 24.9236
R21310 OUT2.n136 OUT2.t40 24.9236
R21311 OUT2.n137 OUT2.t26 24.9236
R21312 OUT2.n137 OUT2.t56 24.9236
R21313 OUT2.n139 OUT2.t35 24.9236
R21314 OUT2.n139 OUT2.t12 24.9236
R21315 OUT2.n141 OUT2.t46 24.9236
R21316 OUT2.n141 OUT2.t0 24.9236
R21317 OUT2.n143 OUT2.t62 24.9236
R21318 OUT2.n143 OUT2.t15 24.9236
R21319 OUT2.n145 OUT2.t21 24.9236
R21320 OUT2.n145 OUT2.t51 24.9236
R21321 OUT2.n147 OUT2.t32 24.9236
R21322 OUT2.n147 OUT2.t8 24.9236
R21323 OUT2.n94 OUT2.t31 24.9236
R21324 OUT2.n94 OUT2.t60 24.9236
R21325 OUT2.n81 OUT2.t50 24.9236
R21326 OUT2.n81 OUT2.t59 24.9236
R21327 OUT2.n82 OUT2.t2 24.9236
R21328 OUT2.n82 OUT2.t39 24.9236
R21329 OUT2.n84 OUT2.t17 24.9236
R21330 OUT2.n84 OUT2.t53 24.9236
R21331 OUT2.n86 OUT2.t52 24.9236
R21332 OUT2.n86 OUT2.t1 24.9236
R21333 OUT2.n88 OUT2.t9 24.9236
R21334 OUT2.n88 OUT2.t23 24.9236
R21335 OUT2.n90 OUT2.t22 24.9236
R21336 OUT2.n90 OUT2.t41 24.9236
R21337 OUT2.n92 OUT2.t11 24.9236
R21338 OUT2.n92 OUT2.t43 24.9236
R21339 OUT2.n55 OUT2.t37 24.9236
R21340 OUT2.n55 OUT2.t7 24.9236
R21341 OUT2.n42 OUT2.t57 24.9236
R21342 OUT2.n42 OUT2.t5 24.9236
R21343 OUT2.n43 OUT2.t3 24.9236
R21344 OUT2.n43 OUT2.t27 24.9236
R21345 OUT2.n45 OUT2.t24 24.9236
R21346 OUT2.n45 OUT2.t54 24.9236
R21347 OUT2.n47 OUT2.t16 24.9236
R21348 OUT2.n47 OUT2.t48 24.9236
R21349 OUT2.n49 OUT2.t44 24.9236
R21350 OUT2.n49 OUT2.t63 24.9236
R21351 OUT2.n51 OUT2.t61 24.9236
R21352 OUT2.n51 OUT2.t14 24.9236
R21353 OUT2.n53 OUT2.t20 24.9236
R21354 OUT2.n53 OUT2.t33 24.9236
R21355 OUT2.n15 OUT2.t36 24.9236
R21356 OUT2.n15 OUT2.t49 24.9236
R21357 OUT2.n2 OUT2.t55 24.9236
R21358 OUT2.n2 OUT2.t13 24.9236
R21359 OUT2.n3 OUT2.t10 24.9236
R21360 OUT2.n3 OUT2.t25 24.9236
R21361 OUT2.n5 OUT2.t30 24.9236
R21362 OUT2.n5 OUT2.t42 24.9236
R21363 OUT2.n7 OUT2.t47 24.9236
R21364 OUT2.n7 OUT2.t18 24.9236
R21365 OUT2.n9 OUT2.t58 24.9236
R21366 OUT2.n9 OUT2.t29 24.9236
R21367 OUT2.n11 OUT2.t34 24.9236
R21368 OUT2.n11 OUT2.t45 24.9236
R21369 OUT2.n13 OUT2.t28 24.9236
R21370 OUT2.n13 OUT2.t38 24.9236
R21371 OUT2 OUT2.n150 11.4429
R21372 OUT2 OUT2.n95 11.4429
R21373 OUT2 OUT2.n58 11.4429
R21374 OUT2 OUT2.n18 11.4429
R21375 OUT2.n77 OUT2.n62 8.55118
R21376 OUT2.n37 OUT2.n22 8.55118
R21377 OUT2.n114 OUT2.n99 8.55117
R21378 OUT2.n119 OUT2.n118 8.47293
R21379 OUT2.n56 OUT2.n55 7.80093
R21380 OUT2.n16 OUT2.n15 7.80093
R21381 OUT2.n78 OUT2.n77 3.20954
R21382 OUT2.n38 OUT2.n37 3.20953
R21383 OUT2.n115 OUT2.n114 3.20289
R21384 OUT2.n151 OUT2 3.10353
R21385 OUT2.n96 OUT2 3.10353
R21386 OUT2.n59 OUT2 3.10353
R21387 OUT2.n19 OUT2 3.10353
R21388 OUT2.n135 OUT2.n134 3.1005
R21389 OUT2.n57 OUT2.n41 3.1005
R21390 OUT2.n17 OUT2.n1 3.1005
R21391 OUT2.n134 OUT2.n133 2.71565
R21392 OUT2.n114 OUT2.n113 2.13383
R21393 OUT2.n77 OUT2.n76 2.13383
R21394 OUT2.n37 OUT2.n36 2.13383
R21395 OUT2.n150 OUT2 1.74595
R21396 OUT2.n95 OUT2 1.74595
R21397 OUT2.n58 OUT2.n57 1.16414
R21398 OUT2.n18 OUT2.n17 1.16414
R21399 OUT2.n157 OUT2.n156 1.07337
R21400 OUT2.n158 OUT2.n157 0.69375
R21401 OUT2.n159 OUT2.n158 0.68905
R21402 OUT2.n56 OUT2 0.488972
R21403 OUT2.n16 OUT2 0.488972
R21404 OUT2.n158 OUT2.n79 0.414635
R21405 OUT2.n157 OUT2.n116 0.382465
R21406 OUT2.n159 OUT2.n39 0.368576
R21407 OUT2 OUT2.n159 0.281623
R21408 OUT2.n134 OUT2.n119 0.196887
R21409 OUT2.n79 OUT2.n78 0.157252
R21410 OUT2.n39 OUT2.n38 0.139891
R21411 OUT2.n156 OUT2.n155 0.139389
R21412 OUT2.n116 OUT2.n115 0.132946
R21413 OUT2.n60 OUT2.n41 0.113
R21414 OUT2.n20 OUT2.n1 0.113
R21415 OUT2.n154 OUT2.n135 0.101889
R21416 OUT2.n57 OUT2.n56 0.0893205
R21417 OUT2.n17 OUT2.n16 0.0893205
R21418 OUT2.n154 OUT2.n152 0.0282778
R21419 OUT2.n135 OUT2.n117 0.0268889
R21420 OUT2.n98 OUT2.n97 0.0213333
R21421 OUT2.n61 OUT2.n60 0.0143889
R21422 OUT2.n21 OUT2.n20 0.0143889
R21423 OUT2.n115 OUT2.n98 0.00100004
R21424 OUT2.n38 OUT2.n21 0.00100004
R21425 OUT2.n78 OUT2.n61 0.00100004
R21426 OUT2.n152 OUT2.n151 0.000513335
R21427 OUT2.n97 OUT2.n96 0.000513335
R21428 OUT2.n60 OUT2.n59 0.000513218
R21429 OUT2.n20 OUT2.n19 0.000513218
R21430 OUT2.n98 OUT2.n80 0.00050517
R21431 OUT2.n154 OUT2.n153 0.000504838
R21432 OUT2.n61 OUT2.n40 0.000504838
R21433 OUT2.n21 OUT2.n0 0.000504838
R21434 OUT2.n155 OUT2.n154 0.000501713
R21435 VFS.n3 VFS 0.239679
R21436 VFS.n4 VFS.t2 0.0274553
R21437 VFS.n0 VFS.t5 0.0274553
R21438 VFS.n1 VFS.n0 0.0274531
R21439 VFS.n2 VFS.n1 0.0274531
R21440 VFS.n6 VFS.n5 0.0274531
R21441 VFS.n5 VFS.n4 0.0274531
R21442 VFS VFS.n6 0.014671
R21443 VFS.n3 VFS.n2 0.011546
R21444 VFS VFS.n3 0.00223611
R21445 VFS.n4 VFS.t7 0.000502142
R21446 VFS.n5 VFS.t4 0.000502142
R21447 VFS.n6 VFS.t6 0.000502142
R21448 VFS.n2 VFS.t3 0.000502142
R21449 VFS.n1 VFS.t1 0.000502142
R21450 VFS.n0 VFS.t0 0.000502142
R21451 VV16.n0 VV16.t17 167.365
R21452 VV16.n0 VV16.t16 92.4496
R21453 VV16.n1 VV16.n0 2.07493
R21454 VV16.n17 VV16 0.8559
R21455 VV16 VV16.n17 0.356917
R21456 VV16.n15 VV16.n14 0.141409
R21457 VV16.n13 VV16.n12 0.141409
R21458 VV16.n11 VV16.n10 0.141409
R21459 VV16.n9 VV16.n8 0.141409
R21460 VV16.n7 VV16.n6 0.141409
R21461 VV16.n5 VV16.n4 0.141409
R21462 VV16.n3 VV16.n2 0.141409
R21463 VV16.n1 VV16 0.12425
R21464 VV16 VV16.n16 0.105614
R21465 VV16 VV16.n1 0.05
R21466 VV16.n17 VV16 0.0193
R21467 VV16.n17 VV16 0.00833333
R21468 VV16.n2 VV16.t13 0.000729415
R21469 VV16.n16 VV16.n15 0.000727273
R21470 VV16.n14 VV16.n13 0.000727273
R21471 VV16.n12 VV16.n11 0.000727273
R21472 VV16.n10 VV16.n9 0.000727273
R21473 VV16.n8 VV16.n7 0.000727273
R21474 VV16.n6 VV16.n5 0.000727273
R21475 VV16.n4 VV16.n3 0.000727273
R21476 VV16.n3 VV16.t14 0.000502142
R21477 VV16.n5 VV16.t15 0.000502142
R21478 VV16.n7 VV16.t5 0.000502142
R21479 VV16.n9 VV16.t7 0.000502142
R21480 VV16.n11 VV16.t0 0.000502142
R21481 VV16.n13 VV16.t2 0.000502142
R21482 VV16.n15 VV16.t1 0.000502142
R21483 VV16.n16 VV16.t10 0.000502142
R21484 VV16.n14 VV16.t3 0.000502142
R21485 VV16.n12 VV16.t4 0.000502142
R21486 VV16.n10 VV16.t8 0.000502142
R21487 VV16.n8 VV16.t11 0.000502142
R21488 VV16.n6 VV16.t9 0.000502142
R21489 VV16.n4 VV16.t12 0.000502142
R21490 VV16.n2 VV16.t6 0.000502142
R21491 a_16599_n13205.n12 a_16599_n13205.t21 182.77
R21492 a_16599_n13205.n13 a_16599_n13205.t14 182.77
R21493 a_16599_n13205.n14 a_16599_n13205.t6 182.77
R21494 a_16599_n13205.n15 a_16599_n13205.t10 182.77
R21495 a_16599_n13205.n16 a_16599_n13205.t18 182.77
R21496 a_16599_n13205.n17 a_16599_n13205.t4 182.77
R21497 a_16599_n13205.n18 a_16599_n13205.t19 182.77
R21498 a_16599_n13205.n19 a_16599_n13205.t9 182.77
R21499 a_16599_n13205.n20 a_16599_n13205.t5 182.77
R21500 a_16599_n13205.n21 a_16599_n13205.t2 182.77
R21501 a_16599_n13205.n2 a_16599_n13205.t8 182.77
R21502 a_16599_n13205.n3 a_16599_n13205.t23 182.77
R21503 a_16599_n13205.n4 a_16599_n13205.t12 182.77
R21504 a_16599_n13205.n5 a_16599_n13205.t20 182.77
R21505 a_16599_n13205.n6 a_16599_n13205.t13 182.77
R21506 a_16599_n13205.n7 a_16599_n13205.t7 182.77
R21507 a_16599_n13205.n8 a_16599_n13205.t22 182.77
R21508 a_16599_n13205.n9 a_16599_n13205.t11 182.77
R21509 a_16599_n13205.n10 a_16599_n13205.t16 182.77
R21510 a_16599_n13205.n11 a_16599_n13205.t17 90.7933
R21511 a_16599_n13205.n1 a_16599_n13205.t15 90.7875
R21512 a_16599_n13205.n43 a_16599_n13205.t0 42.4202
R21513 a_16599_n13205.n0 a_16599_n13205.t3 4.35105
R21514 a_16599_n13205.t1 a_16599_n13205.n43 2.70045
R21515 a_16599_n13205.n2 a_16599_n13205.n1 2.03273
R21516 a_16599_n13205.n12 a_16599_n13205.n11 2.02124
R21517 a_16599_n13205.n41 a_16599_n13205.n40 0.835222
R21518 a_16599_n13205.n40 a_16599_n13205.n39 0.835222
R21519 a_16599_n13205.n39 a_16599_n13205.n38 0.835222
R21520 a_16599_n13205.n38 a_16599_n13205.n37 0.835222
R21521 a_16599_n13205.n37 a_16599_n13205.n36 0.835222
R21522 a_16599_n13205.n36 a_16599_n13205.n35 0.835222
R21523 a_16599_n13205.n35 a_16599_n13205.n34 0.835222
R21524 a_16599_n13205.n34 a_16599_n13205.n33 0.835222
R21525 a_16599_n13205.n33 a_16599_n13205.n32 0.835222
R21526 a_16599_n13205.n13 a_16599_n13205.n12 0.835222
R21527 a_16599_n13205.n14 a_16599_n13205.n13 0.835222
R21528 a_16599_n13205.n15 a_16599_n13205.n14 0.835222
R21529 a_16599_n13205.n16 a_16599_n13205.n15 0.835222
R21530 a_16599_n13205.n17 a_16599_n13205.n16 0.835222
R21531 a_16599_n13205.n18 a_16599_n13205.n17 0.835222
R21532 a_16599_n13205.n19 a_16599_n13205.n18 0.835222
R21533 a_16599_n13205.n20 a_16599_n13205.n19 0.835222
R21534 a_16599_n13205.n21 a_16599_n13205.n20 0.835222
R21535 a_16599_n13205.n10 a_16599_n13205.n9 0.835222
R21536 a_16599_n13205.n9 a_16599_n13205.n8 0.835222
R21537 a_16599_n13205.n8 a_16599_n13205.n7 0.835222
R21538 a_16599_n13205.n7 a_16599_n13205.n6 0.835222
R21539 a_16599_n13205.n6 a_16599_n13205.n5 0.835222
R21540 a_16599_n13205.n5 a_16599_n13205.n4 0.835222
R21541 a_16599_n13205.n4 a_16599_n13205.n3 0.835222
R21542 a_16599_n13205.n3 a_16599_n13205.n2 0.835222
R21543 a_16599_n13205.n24 a_16599_n13205.n23 0.835222
R21544 a_16599_n13205.n25 a_16599_n13205.n24 0.835222
R21545 a_16599_n13205.n26 a_16599_n13205.n25 0.835222
R21546 a_16599_n13205.n27 a_16599_n13205.n26 0.835222
R21547 a_16599_n13205.n28 a_16599_n13205.n27 0.835222
R21548 a_16599_n13205.n29 a_16599_n13205.n28 0.835222
R21549 a_16599_n13205.n30 a_16599_n13205.n29 0.835222
R21550 a_16599_n13205.n31 a_16599_n13205.n30 0.835222
R21551 a_16599_n13205.n0 a_16599_n13205.n42 0.750184
R21552 a_16599_n13205.n0 a_16599_n13205.n22 0.715064
R21553 a_16599_n13205.n22 a_16599_n13205.n10 0.553972
R21554 a_16599_n13205.n42 a_16599_n13205.n31 0.553972
R21555 a_16599_n13205.n43 a_16599_n13205.n0 0.403234
R21556 a_16599_n13205.n42 a_16599_n13205.n41 0.233139
R21557 a_16599_n13205.n22 a_16599_n13205.n21 0.233139
R21558 a_16541_n13117.n0 a_16541_n13117.t16 5.73525
R21559 a_16541_n13117.n18 a_16541_n13117.t14 5.34571
R21560 a_16541_n13117.n0 a_16541_n13117.t4 5.18362
R21561 a_16541_n13117.n1 a_16541_n13117.t8 5.18362
R21562 a_16541_n13117.n2 a_16541_n13117.t19 5.18362
R21563 a_16541_n13117.n3 a_16541_n13117.t11 5.18362
R21564 a_16541_n13117.n4 a_16541_n13117.t18 5.18362
R21565 a_16541_n13117.n5 a_16541_n13117.t5 5.18362
R21566 a_16541_n13117.n6 a_16541_n13117.t9 5.18362
R21567 a_16541_n13117.n7 a_16541_n13117.t20 5.18362
R21568 a_16541_n13117.n8 a_16541_n13117.t15 5.18362
R21569 a_16541_n13117.n9 a_16541_n13117.t7 5.18362
R21570 a_16541_n13117.n10 a_16541_n13117.t3 5.18362
R21571 a_16541_n13117.n11 a_16541_n13117.t12 5.18362
R21572 a_16541_n13117.n12 a_16541_n13117.t21 5.18362
R21573 a_16541_n13117.n13 a_16541_n13117.t13 5.18362
R21574 a_16541_n13117.n14 a_16541_n13117.t2 5.18362
R21575 a_16541_n13117.n15 a_16541_n13117.t6 5.18362
R21576 a_16541_n13117.n16 a_16541_n13117.t17 5.18362
R21577 a_16541_n13117.n17 a_16541_n13117.t10 5.18362
R21578 a_16541_n13117.t0 a_16541_n13117.n19 2.79552
R21579 a_16541_n13117.n19 a_16541_n13117.t1 2.38201
R21580 a_16541_n13117.n9 a_16541_n13117.n8 1.10376
R21581 a_16541_n13117.n1 a_16541_n13117.n0 0.55213
R21582 a_16541_n13117.n2 a_16541_n13117.n1 0.55213
R21583 a_16541_n13117.n3 a_16541_n13117.n2 0.55213
R21584 a_16541_n13117.n4 a_16541_n13117.n3 0.55213
R21585 a_16541_n13117.n5 a_16541_n13117.n4 0.55213
R21586 a_16541_n13117.n6 a_16541_n13117.n5 0.55213
R21587 a_16541_n13117.n7 a_16541_n13117.n6 0.55213
R21588 a_16541_n13117.n8 a_16541_n13117.n7 0.55213
R21589 a_16541_n13117.n10 a_16541_n13117.n9 0.55213
R21590 a_16541_n13117.n11 a_16541_n13117.n10 0.55213
R21591 a_16541_n13117.n12 a_16541_n13117.n11 0.55213
R21592 a_16541_n13117.n13 a_16541_n13117.n12 0.55213
R21593 a_16541_n13117.n14 a_16541_n13117.n13 0.55213
R21594 a_16541_n13117.n15 a_16541_n13117.n14 0.55213
R21595 a_16541_n13117.n16 a_16541_n13117.n15 0.55213
R21596 a_16541_n13117.n17 a_16541_n13117.n16 0.512683
R21597 a_16541_n13117.n19 a_16541_n13117.n18 0.168655
R21598 a_16541_n13117.n18 a_16541_n13117.n17 0.0581389
R21599 a_16719_n13117.n15 a_16719_n13117.t24 473.437
R21600 a_16719_n13117.n19 a_16719_n13117.t25 473.332
R21601 a_16719_n13117.n0 a_16719_n13117.t0 473.329
R21602 a_16719_n13117.n18 a_16719_n13117.t2 140.444
R21603 a_16719_n13117.n18 a_16719_n13117.t3 41.6504
R21604 a_16719_n13117.n2 a_16719_n13117.t12 5.95597
R21605 a_16719_n13117.n26 a_16719_n13117.t10 5.95597
R21606 a_16719_n13117.n8 a_16719_n13117.t5 5.32159
R21607 a_16719_n13117.n7 a_16719_n13117.t20 5.32159
R21608 a_16719_n13117.n6 a_16719_n13117.t14 5.32159
R21609 a_16719_n13117.n5 a_16719_n13117.t7 5.32159
R21610 a_16719_n13117.n4 a_16719_n13117.t15 5.32159
R21611 a_16719_n13117.n3 a_16719_n13117.t4 5.32159
R21612 a_16719_n13117.n2 a_16719_n13117.t19 5.32159
R21613 a_16719_n13117.n1 a_16719_n13117.t11 5.32159
R21614 a_16719_n13117.n11 a_16719_n13117.t16 5.32159
R21615 a_16719_n13117.n26 a_16719_n13117.t6 5.32159
R21616 a_16719_n13117.n27 a_16719_n13117.t13 5.32159
R21617 a_16719_n13117.n28 a_16719_n13117.t21 5.32159
R21618 a_16719_n13117.n29 a_16719_n13117.t17 5.32159
R21619 a_16719_n13117.n30 a_16719_n13117.t9 5.32159
R21620 a_16719_n13117.n25 a_16719_n13117.t8 5.32159
R21621 a_16719_n13117.n24 a_16719_n13117.t18 5.32159
R21622 a_16719_n13117.n23 a_16719_n13117.t22 5.32159
R21623 a_16719_n13117.t23 a_16719_n13117.n31 5.32059
R21624 a_16719_n13117.n14 a_16719_n13117.n13 2.75606
R21625 a_16719_n13117.n17 a_16719_n13117.n14 2.75328
R21626 a_16719_n13117.n14 a_16719_n13117.t1 1.50409
R21627 a_16719_n13117.n19 a_16719_n13117.n18 1.23545
R21628 a_16719_n13117.n23 a_16719_n13117.n22 1.02772
R21629 a_16719_n13117.n3 a_16719_n13117.n2 0.634875
R21630 a_16719_n13117.n4 a_16719_n13117.n3 0.634875
R21631 a_16719_n13117.n5 a_16719_n13117.n4 0.634875
R21632 a_16719_n13117.n6 a_16719_n13117.n5 0.634875
R21633 a_16719_n13117.n7 a_16719_n13117.n6 0.634875
R21634 a_16719_n13117.n8 a_16719_n13117.n7 0.634875
R21635 a_16719_n13117.n24 a_16719_n13117.n23 0.634875
R21636 a_16719_n13117.n25 a_16719_n13117.n24 0.634875
R21637 a_16719_n13117.n31 a_16719_n13117.n25 0.634875
R21638 a_16719_n13117.n31 a_16719_n13117.n30 0.634875
R21639 a_16719_n13117.n30 a_16719_n13117.n29 0.634875
R21640 a_16719_n13117.n29 a_16719_n13117.n28 0.634875
R21641 a_16719_n13117.n28 a_16719_n13117.n27 0.634875
R21642 a_16719_n13117.n27 a_16719_n13117.n26 0.634875
R21643 a_16719_n13117.n0 a_16719_n13117.n21 0.376529
R21644 a_16719_n13117.n16 a_16719_n13117.n15 0.271346
R21645 a_16719_n13117.n21 a_16719_n13117.n20 0.253053
R21646 a_16719_n13117.n9 a_16719_n13117.n8 0.202227
R21647 a_16719_n13117.n20 a_16719_n13117.n19 0.124538
R21648 a_16719_n13117.n17 a_16719_n13117.n16 0.119076
R21649 a_16719_n13117.n13 a_16719_n13117.n12 0.113872
R21650 a_16719_n13117.n0 a_16719_n13117.n17 0.10111
R21651 a_16719_n13117.n1 a_16719_n13117.n0 0.0537895
R21652 a_16719_n13117.n10 a_16719_n13117.n9 0.0386579
R21653 a_16719_n13117.n22 a_16719_n13117.n1 0.0360263
R21654 a_16719_n13117.n0 a_16719_n13117.n11 0.035794
R21655 a_16719_n13117.n11 a_16719_n13117.n10 0.0202368
R21656 CLK.t85 CLK.t89 344.122
R21657 CLK.t72 CLK.t34 344.122
R21658 CLK.t60 CLK.t16 344.122
R21659 CLK.t7 CLK.t57 344.122
R21660 CLK.t87 CLK.t36 344.122
R21661 CLK.t28 CLK.t80 344.122
R21662 CLK.t13 CLK.t70 344.122
R21663 CLK.t51 CLK.t6 344.122
R21664 CLK.t39 CLK.t95 344.122
R21665 CLK.t74 CLK.t71 344.122
R21666 CLK.t64 CLK.t18 344.122
R21667 CLK.t47 CLK.t5 344.122
R21668 CLK.t90 CLK.t38 344.122
R21669 CLK.t73 CLK.t27 344.122
R21670 CLK.t14 CLK.t63 344.122
R21671 CLK.t48 CLK.t46 344.122
R21672 CLK.n3 CLK.t50 232.299
R21673 CLK.n130 CLK.t42 232.299
R21674 CLK.n121 CLK.t84 232.299
R21675 CLK.n112 CLK.t67 232.299
R21676 CLK.n103 CLK.t52 232.299
R21677 CLK.n94 CLK.t1 232.299
R21678 CLK.n85 CLK.t75 232.299
R21679 CLK.n76 CLK.t21 232.299
R21680 CLK.n67 CLK.t3 232.299
R21681 CLK.n58 CLK.t43 232.299
R21682 CLK.n49 CLK.t31 232.299
R21683 CLK.n40 CLK.t68 232.299
R21684 CLK.n31 CLK.t55 232.299
R21685 CLK.n22 CLK.t93 232.299
R21686 CLK.n13 CLK.t77 232.299
R21687 CLK.n152 CLK.t22 232.299
R21688 CLK.n6 CLK.t94 182.915
R21689 CLK.n133 CLK.t81 182.915
R21690 CLK.n124 CLK.t61 182.915
R21691 CLK.n115 CLK.t8 182.915
R21692 CLK.n106 CLK.t88 182.915
R21693 CLK.n97 CLK.t29 182.915
R21694 CLK.n88 CLK.t19 182.915
R21695 CLK.n79 CLK.t53 182.915
R21696 CLK.n70 CLK.t40 182.915
R21697 CLK.n61 CLK.t76 182.915
R21698 CLK.n52 CLK.t65 182.915
R21699 CLK.n43 CLK.t10 182.915
R21700 CLK.n34 CLK.t91 182.915
R21701 CLK.n25 CLK.t32 182.915
R21702 CLK.n16 CLK.t15 182.915
R21703 CLK.n155 CLK.t49 182.915
R21704 CLK.n6 CLK.t85 182.91
R21705 CLK.n133 CLK.t72 182.91
R21706 CLK.n124 CLK.t60 182.91
R21707 CLK.n115 CLK.t7 182.91
R21708 CLK.n106 CLK.t87 182.91
R21709 CLK.n97 CLK.t28 182.91
R21710 CLK.n88 CLK.t13 182.91
R21711 CLK.n79 CLK.t51 182.91
R21712 CLK.n70 CLK.t39 182.91
R21713 CLK.n61 CLK.t74 182.91
R21714 CLK.n52 CLK.t64 182.91
R21715 CLK.n43 CLK.t47 182.91
R21716 CLK.n34 CLK.t90 182.91
R21717 CLK.n25 CLK.t73 182.91
R21718 CLK.n16 CLK.t14 182.91
R21719 CLK.n155 CLK.t48 182.91
R21720 CLK.t94 CLK.n5 182.769
R21721 CLK.t81 CLK.n132 182.769
R21722 CLK.t61 CLK.n123 182.769
R21723 CLK.t8 CLK.n114 182.769
R21724 CLK.t88 CLK.n105 182.769
R21725 CLK.t29 CLK.n96 182.769
R21726 CLK.t19 CLK.n87 182.769
R21727 CLK.t53 CLK.n78 182.769
R21728 CLK.t40 CLK.n69 182.769
R21729 CLK.t76 CLK.n60 182.769
R21730 CLK.t65 CLK.n51 182.769
R21731 CLK.t10 CLK.n42 182.769
R21732 CLK.t91 CLK.n33 182.769
R21733 CLK.t32 CLK.n24 182.769
R21734 CLK.t15 CLK.n15 182.769
R21735 CLK.t49 CLK.n154 182.769
R21736 CLK.n1 CLK.t26 161.262
R21737 CLK.n128 CLK.t59 161.262
R21738 CLK.n119 CLK.t37 161.262
R21739 CLK.n110 CLK.t82 161.262
R21740 CLK.n101 CLK.t62 161.262
R21741 CLK.n92 CLK.t9 161.262
R21742 CLK.n83 CLK.t0 161.262
R21743 CLK.n74 CLK.t30 161.262
R21744 CLK.n65 CLK.t20 161.262
R21745 CLK.n56 CLK.t54 161.262
R21746 CLK.n47 CLK.t41 161.262
R21747 CLK.n38 CLK.t83 161.262
R21748 CLK.n29 CLK.t66 161.262
R21749 CLK.n20 CLK.t11 161.262
R21750 CLK.n11 CLK.t92 161.262
R21751 CLK.n150 CLK.t86 161.262
R21752 CLK.n7 CLK.t23 159.958
R21753 CLK.n134 CLK.t24 159.958
R21754 CLK.n125 CLK.t12 159.958
R21755 CLK.n116 CLK.t44 159.958
R21756 CLK.n107 CLK.t33 159.958
R21757 CLK.n98 CLK.t69 159.958
R21758 CLK.n89 CLK.t56 159.958
R21759 CLK.n80 CLK.t2 159.958
R21760 CLK.n71 CLK.t79 159.958
R21761 CLK.n62 CLK.t25 159.958
R21762 CLK.n53 CLK.t4 159.958
R21763 CLK.n44 CLK.t45 159.958
R21764 CLK.n35 CLK.t35 159.958
R21765 CLK.n26 CLK.t17 159.958
R21766 CLK.n17 CLK.t58 159.958
R21767 CLK.n156 CLK.t78 159.958
R21768 CLK.n136 CLK.n135 1.5536
R21769 CLK.n9 CLK.n8 1.06552
R21770 CLK.n136 CLK.n126 1.06552
R21771 CLK.n137 CLK.n117 1.06552
R21772 CLK.n138 CLK.n108 1.06552
R21773 CLK.n139 CLK.n99 1.06552
R21774 CLK.n140 CLK.n90 1.06552
R21775 CLK.n141 CLK.n81 1.06552
R21776 CLK.n142 CLK.n72 1.06552
R21777 CLK.n143 CLK.n63 1.06552
R21778 CLK.n144 CLK.n54 1.06552
R21779 CLK.n145 CLK.n45 1.06552
R21780 CLK.n146 CLK.n36 1.06552
R21781 CLK.n147 CLK.n27 1.06552
R21782 CLK.n148 CLK.n18 1.06552
R21783 CLK.n157 CLK.n149 1.06552
R21784 CLK.n7 CLK.n6 0.56781
R21785 CLK.n134 CLK.n133 0.56781
R21786 CLK.n125 CLK.n124 0.56781
R21787 CLK.n116 CLK.n115 0.56781
R21788 CLK.n107 CLK.n106 0.56781
R21789 CLK.n98 CLK.n97 0.56781
R21790 CLK.n89 CLK.n88 0.56781
R21791 CLK.n80 CLK.n79 0.56781
R21792 CLK.n71 CLK.n70 0.56781
R21793 CLK.n62 CLK.n61 0.56781
R21794 CLK.n53 CLK.n52 0.56781
R21795 CLK.n44 CLK.n43 0.56781
R21796 CLK.n35 CLK.n34 0.56781
R21797 CLK.n26 CLK.n25 0.56781
R21798 CLK.n17 CLK.n16 0.56781
R21799 CLK.n156 CLK.n155 0.56781
R21800 CLK.n149 CLK.n9 0.488577
R21801 CLK.n149 CLK.n148 0.488577
R21802 CLK.n148 CLK.n147 0.488577
R21803 CLK.n147 CLK.n146 0.488577
R21804 CLK.n146 CLK.n145 0.488577
R21805 CLK.n145 CLK.n144 0.488577
R21806 CLK.n144 CLK.n143 0.488577
R21807 CLK.n143 CLK.n142 0.488577
R21808 CLK.n142 CLK.n141 0.488577
R21809 CLK.n141 CLK.n140 0.488577
R21810 CLK.n140 CLK.n139 0.488577
R21811 CLK.n139 CLK.n138 0.488577
R21812 CLK.n138 CLK.n137 0.488577
R21813 CLK.n137 CLK.n136 0.488577
R21814 CLK.n8 CLK.n7 0.428385
R21815 CLK.n135 CLK.n134 0.428385
R21816 CLK.n126 CLK.n125 0.428385
R21817 CLK.n117 CLK.n116 0.428385
R21818 CLK.n108 CLK.n107 0.428385
R21819 CLK.n99 CLK.n98 0.428385
R21820 CLK.n90 CLK.n89 0.428385
R21821 CLK.n81 CLK.n80 0.428385
R21822 CLK.n72 CLK.n71 0.428385
R21823 CLK.n63 CLK.n62 0.428385
R21824 CLK.n54 CLK.n53 0.428385
R21825 CLK.n45 CLK.n44 0.428385
R21826 CLK.n36 CLK.n35 0.428385
R21827 CLK.n27 CLK.n26 0.428385
R21828 CLK.n18 CLK.n17 0.428385
R21829 CLK.n157 CLK.n156 0.428385
R21830 CLK.n9 CLK 0.316644
R21831 CLK.n0 CLK 0.12425
R21832 CLK.n127 CLK 0.12425
R21833 CLK.n118 CLK 0.12425
R21834 CLK.n109 CLK 0.12425
R21835 CLK.n100 CLK 0.12425
R21836 CLK.n91 CLK 0.12425
R21837 CLK.n82 CLK 0.12425
R21838 CLK.n73 CLK 0.12425
R21839 CLK.n64 CLK 0.12425
R21840 CLK.n55 CLK 0.12425
R21841 CLK.n46 CLK 0.12425
R21842 CLK.n37 CLK 0.12425
R21843 CLK.n28 CLK 0.12425
R21844 CLK.n19 CLK 0.12425
R21845 CLK.n10 CLK 0.12425
R21846 CLK.n158 CLK 0.12425
R21847 CLK.n0 CLK 0.0636313
R21848 CLK.n127 CLK 0.0636313
R21849 CLK.n118 CLK 0.0636313
R21850 CLK.n109 CLK 0.0636313
R21851 CLK.n100 CLK 0.0636313
R21852 CLK.n91 CLK 0.0636313
R21853 CLK.n82 CLK 0.0636313
R21854 CLK.n73 CLK 0.0636313
R21855 CLK.n64 CLK 0.0636313
R21856 CLK.n55 CLK 0.0636313
R21857 CLK.n46 CLK 0.0636313
R21858 CLK.n37 CLK 0.0636313
R21859 CLK.n28 CLK 0.0636313
R21860 CLK.n19 CLK 0.0636313
R21861 CLK.n10 CLK 0.0636313
R21862 CLK CLK.n158 0.0636313
R21863 CLK.n0 CLK 0.0484798
R21864 CLK.n127 CLK 0.0484798
R21865 CLK.n118 CLK 0.0484798
R21866 CLK.n109 CLK 0.0484798
R21867 CLK.n100 CLK 0.0484798
R21868 CLK.n91 CLK 0.0484798
R21869 CLK.n82 CLK 0.0484798
R21870 CLK.n73 CLK 0.0484798
R21871 CLK.n64 CLK 0.0484798
R21872 CLK.n55 CLK 0.0484798
R21873 CLK.n46 CLK 0.0484798
R21874 CLK.n37 CLK 0.0484798
R21875 CLK.n28 CLK 0.0484798
R21876 CLK.n19 CLK 0.0484798
R21877 CLK.n10 CLK 0.0484798
R21878 CLK.n158 CLK 0.0484798
R21879 CLK.n2 CLK.n1 0.0178077
R21880 CLK.n129 CLK.n128 0.0178077
R21881 CLK.n120 CLK.n119 0.0178077
R21882 CLK.n111 CLK.n110 0.0178077
R21883 CLK.n102 CLK.n101 0.0178077
R21884 CLK.n93 CLK.n92 0.0178077
R21885 CLK.n84 CLK.n83 0.0178077
R21886 CLK.n75 CLK.n74 0.0178077
R21887 CLK.n66 CLK.n65 0.0178077
R21888 CLK.n57 CLK.n56 0.0178077
R21889 CLK.n48 CLK.n47 0.0178077
R21890 CLK.n39 CLK.n38 0.0178077
R21891 CLK.n30 CLK.n29 0.0178077
R21892 CLK.n21 CLK.n20 0.0178077
R21893 CLK.n12 CLK.n11 0.0178077
R21894 CLK.n151 CLK.n150 0.0178077
R21895 CLK.n5 CLK.n2 0.00531334
R21896 CLK.n132 CLK.n129 0.00531334
R21897 CLK.n123 CLK.n120 0.00531334
R21898 CLK.n114 CLK.n111 0.00531334
R21899 CLK.n105 CLK.n102 0.00531334
R21900 CLK.n96 CLK.n93 0.00531334
R21901 CLK.n87 CLK.n84 0.00531334
R21902 CLK.n78 CLK.n75 0.00531334
R21903 CLK.n69 CLK.n66 0.00531334
R21904 CLK.n60 CLK.n57 0.00531334
R21905 CLK.n51 CLK.n48 0.00531334
R21906 CLK.n42 CLK.n39 0.00531334
R21907 CLK.n33 CLK.n30 0.00531334
R21908 CLK.n24 CLK.n21 0.00531334
R21909 CLK.n15 CLK.n12 0.00531334
R21910 CLK.n154 CLK.n151 0.00531334
R21911 CLK.n5 CLK.n4 0.00224847
R21912 CLK.n132 CLK.n131 0.00224847
R21913 CLK.n123 CLK.n122 0.00224847
R21914 CLK.n114 CLK.n113 0.00224847
R21915 CLK.n105 CLK.n104 0.00224847
R21916 CLK.n96 CLK.n95 0.00224847
R21917 CLK.n87 CLK.n86 0.00224847
R21918 CLK.n78 CLK.n77 0.00224847
R21919 CLK.n69 CLK.n68 0.00224847
R21920 CLK.n60 CLK.n59 0.00224847
R21921 CLK.n51 CLK.n50 0.00224847
R21922 CLK.n42 CLK.n41 0.00224847
R21923 CLK.n33 CLK.n32 0.00224847
R21924 CLK.n24 CLK.n23 0.00224847
R21925 CLK.n15 CLK.n14 0.00224847
R21926 CLK.n154 CLK.n153 0.00224847
R21927 CLK.n4 CLK.n3 0.00100535
R21928 CLK.n131 CLK.n130 0.00100535
R21929 CLK.n122 CLK.n121 0.00100535
R21930 CLK.n113 CLK.n112 0.00100535
R21931 CLK.n104 CLK.n103 0.00100535
R21932 CLK.n95 CLK.n94 0.00100535
R21933 CLK.n86 CLK.n85 0.00100535
R21934 CLK.n77 CLK.n76 0.00100535
R21935 CLK.n68 CLK.n67 0.00100535
R21936 CLK.n59 CLK.n58 0.00100535
R21937 CLK.n50 CLK.n49 0.00100535
R21938 CLK.n41 CLK.n40 0.00100535
R21939 CLK.n32 CLK.n31 0.00100535
R21940 CLK.n23 CLK.n22 0.00100535
R21941 CLK.n14 CLK.n13 0.00100535
R21942 CLK.n153 CLK.n152 0.00100535
R21943 CLK.n8 CLK.n0 0.000500711
R21944 CLK.n135 CLK.n127 0.000500711
R21945 CLK.n126 CLK.n118 0.000500711
R21946 CLK.n117 CLK.n109 0.000500711
R21947 CLK.n108 CLK.n100 0.000500711
R21948 CLK.n99 CLK.n91 0.000500711
R21949 CLK.n90 CLK.n82 0.000500711
R21950 CLK.n81 CLK.n73 0.000500711
R21951 CLK.n72 CLK.n64 0.000500711
R21952 CLK.n63 CLK.n55 0.000500711
R21953 CLK.n54 CLK.n46 0.000500711
R21954 CLK.n45 CLK.n37 0.000500711
R21955 CLK.n36 CLK.n28 0.000500711
R21956 CLK.n27 CLK.n19 0.000500711
R21957 CLK.n18 CLK.n10 0.000500711
R21958 CLK.n158 CLK.n157 0.000500711
R21959 frontAnalog_v0p0p1_10.x65.A.n1 frontAnalog_v0p0p1_10.x65.A.t4 260.322
R21960 frontAnalog_v0p0p1_10.x65.A.n3 frontAnalog_v0p0p1_10.x65.A.t7 233.929
R21961 frontAnalog_v0p0p1_10.x65.A.n1 frontAnalog_v0p0p1_10.x65.A.t6 175.169
R21962 frontAnalog_v0p0p1_10.x65.A.n2 frontAnalog_v0p0p1_10.x65.A.t5 160.416
R21963 frontAnalog_v0p0p1_10.x65.A.n4 frontAnalog_v0p0p1_10.x65.A.t3 17.4109
R21964 frontAnalog_v0p0p1_10.x65.A.n4 frontAnalog_v0p0p1_10.x65.A.t2 10.2053
R21965 frontAnalog_v0p0p1_10.x65.A.n0 frontAnalog_v0p0p1_10.x65.A 2.78715
R21966 frontAnalog_v0p0p1_10.x65.A.n0 frontAnalog_v0p0p1_10.x65.A.n1 9.09103
R21967 frontAnalog_v0p0p1_10.x65.A.n6 frontAnalog_v0p0p1_10.x65.A.t0 7.94569
R21968 frontAnalog_v0p0p1_10.x65.A.n2 frontAnalog_v0p0p1_10.x65.A.t1 7.55846
R21969 frontAnalog_v0p0p1_10.x65.A.n5 frontAnalog_v0p0p1_10.x65.A.n3 1.4614
R21970 frontAnalog_v0p0p1_10.x65.A.n3 frontAnalog_v0p0p1_10.x65.A.n2 1.19626
R21971 frontAnalog_v0p0p1_10.x65.A.n6 frontAnalog_v0p0p1_10.x65.A.n5 0.836961
R21972 frontAnalog_v0p0p1_10.x65.A frontAnalog_v0p0p1_10.x65.A.n0 0.390342
R21973 frontAnalog_v0p0p1_10.x65.A.n5 frontAnalog_v0p0p1_10.x65.A.n4 0.154668
R21974 frontAnalog_v0p0p1_10.x65.A frontAnalog_v0p0p1_10.x65.A.n6 0.08175
R21975 VV4.n0 VV4.t17 167.365
R21976 VV4.n0 VV4.t16 92.4488
R21977 VV4.n1 VV4.n0 2.07493
R21978 VV4.n10 VV4 0.572333
R21979 VV4 VV4.n10 0.429375
R21980 VV4.n9 VV4.n8 0.141636
R21981 VV4.n8 VV4.n7 0.141636
R21982 VV4.n7 VV4.n6 0.141636
R21983 VV4.n6 VV4.n5 0.141636
R21984 VV4.n5 VV4.n4 0.141636
R21985 VV4.n4 VV4.n3 0.141636
R21986 VV4.n3 VV4.n2 0.141636
R21987 VV4.n1 VV4 0.12425
R21988 VV4 VV4.n9 0.103284
R21989 VV4 VV4.n1 0.0314375
R21990 VV4.n10 VV4 0.00833333
R21991 VV4.n10 VV4 0.006375
R21992 VV4.n3 VV4.t1 0.000502142
R21993 VV4.n4 VV4.t7 0.000502142
R21994 VV4.n5 VV4.t11 0.000502142
R21995 VV4.n6 VV4.t2 0.000502142
R21996 VV4.n7 VV4.t14 0.000502142
R21997 VV4.n8 VV4.t4 0.000502142
R21998 VV4.n9 VV4.t15 0.000502142
R21999 VV4.n2 VV4.t13 0.000502142
R22000 VV4.n3 VV4.t9 0.000502142
R22001 VV4.n4 VV4.t8 0.000502142
R22002 VV4.n5 VV4.t12 0.000502142
R22003 VV4.n6 VV4.t3 0.000502142
R22004 VV4.n7 VV4.t10 0.000502142
R22005 VV4.n8 VV4.t6 0.000502142
R22006 VV4.n9 VV4.t0 0.000502142
R22007 VV4.n2 VV4.t5 0.000502142
R22008 VV3.n0 VV3.t17 167.365
R22009 VV3.n0 VV3.t16 92.4488
R22010 VV3.n1 VV3.n0 2.07493
R22011 VV3.n17 VV3 0.607583
R22012 VV3 VV3.n17 0.455812
R22013 VV3.n15 VV3.n14 0.141409
R22014 VV3.n13 VV3.n12 0.141409
R22015 VV3.n11 VV3.n10 0.141409
R22016 VV3.n9 VV3.n8 0.141409
R22017 VV3.n7 VV3.n6 0.141409
R22018 VV3.n5 VV3.n4 0.141409
R22019 VV3.n3 VV3.n2 0.141409
R22020 VV3.n1 VV3 0.12425
R22021 VV3 VV3.n16 0.100973
R22022 VV3 VV3.n1 0.0314375
R22023 VV3.n17 VV3 0.00833333
R22024 VV3.n17 VV3 0.006375
R22025 VV3.n2 VV3.t14 0.000729415
R22026 VV3.n16 VV3.n15 0.000727273
R22027 VV3.n14 VV3.n13 0.000727273
R22028 VV3.n12 VV3.n11 0.000727273
R22029 VV3.n10 VV3.n9 0.000727273
R22030 VV3.n8 VV3.n7 0.000727273
R22031 VV3.n6 VV3.n5 0.000727273
R22032 VV3.n4 VV3.n3 0.000727273
R22033 VV3.n3 VV3.t9 0.000502142
R22034 VV3.n5 VV3.t7 0.000502142
R22035 VV3.n7 VV3.t12 0.000502142
R22036 VV3.n9 VV3.t3 0.000502142
R22037 VV3.n11 VV3.t10 0.000502142
R22038 VV3.n13 VV3.t6 0.000502142
R22039 VV3.n15 VV3.t1 0.000502142
R22040 VV3.n2 VV3.t4 0.000502142
R22041 VV3.n4 VV3.t11 0.000502142
R22042 VV3.n6 VV3.t2 0.000502142
R22043 VV3.n8 VV3.t8 0.000502142
R22044 VV3.n10 VV3.t0 0.000502142
R22045 VV3.n12 VV3.t15 0.000502142
R22046 VV3.n14 VV3.t13 0.000502142
R22047 VV3.n16 VV3.t5 0.000502142
R22048 R1.n0 R1.t7 260.322
R22049 R1.n5 R1.t4 233.888
R22050 R1.n0 R1.t5 175.169
R22051 R1.n4 R1.t6 159.725
R22052 R1.n6 R1.t2 17.4109
R22053 R1.n1 R1.n0 9.75129
R22054 R1.n6 R1.t3 9.6037
R22055 R1.n2 R1 9.3005
R22056 R1.n8 R1.t1 8.40929
R22057 R1.n4 R1.t0 8.06629
R22058 R1 R1.n1 3.11453
R22059 R1.n5 R1.n4 1.73501
R22060 R1.n7 R1.n5 0.99025
R22061 R1.n8 R1.n7 0.853186
R22062 R1.n3 R1 0.241354
R22063 R1 R1.n9 0.232207
R22064 R1.n3 R1.n2 0.195812
R22065 R1.n8 R1 0.0945934
R22066 R1 R1.n3 0.0691813
R22067 R1.n2 R1.n1 0.0292043
R22068 R1.n9 R1 0.0142195
R22069 R1.n9 R1.n8 0.0108022
R22070 R1.n9 R1 0.00668132
R22071 R1.n7 R1.n6 0.000500726
R22072 S1.n4 S1.t7 260.322
R22073 S1.n1 S1.t5 233.929
R22074 S1.n4 S1.t4 175.169
R22075 S1.n0 S1.t6 160.416
R22076 S1.n2 S1.t2 17.4109
R22077 S1.n2 S1.t3 10.2053
R22078 S1.n6 S1 9.3005
R22079 S1.n5 S1.n4 9.09103
R22080 S1 S1.t1 7.94569
R22081 S1.n0 S1.t0 7.55846
R22082 S1 S1.n5 3.97938
R22083 S1 S1.n9 1.763
R22084 S1.n9 S1 1.763
R22085 S1.n3 S1.n1 1.4614
R22086 S1.n1 S1.n0 1.19626
R22087 S1.n8 S1.n3 0.808836
R22088 S1.n7 S1.n6 0.223714
R22089 S1.n3 S1.n2 0.154668
R22090 S1.n9 S1 0.0789574
R22091 S1.n9 S1 0.0434878
R22092 S1.n9 S1 0.0434878
R22093 S1.n6 S1.n5 0.0421278
R22094 S1.n7 S1 0.0306829
R22095 S1 S1.n8 0.013
R22096 S1.n8 S1.n7 0.0114756
R22097 frontAnalog_v0p0p1_5.RSfetsym_0.QN.n1 frontAnalog_v0p0p1_5.RSfetsym_0.QN.t6 117.511
R22098 frontAnalog_v0p0p1_5.RSfetsym_0.QN.n1 frontAnalog_v0p0p1_5.RSfetsym_0.QN.t5 110.698
R22099 frontAnalog_v0p0p1_5.RSfetsym_0.QN.n2 frontAnalog_v0p0p1_5.RSfetsym_0.QN.t4 19.1963
R22100 frontAnalog_v0p0p1_5.RSfetsym_0.QN.n3 frontAnalog_v0p0p1_5.RSfetsym_0.QN.t0 14.5206
R22101 frontAnalog_v0p0p1_5.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_5.RSfetsym_0.QN.t3 14.283
R22102 frontAnalog_v0p0p1_5.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_5.RSfetsym_0.QN.t2 14.283
R22103 frontAnalog_v0p0p1_5.RSfetsym_0.QN frontAnalog_v0p0p1_5.RSfetsym_0.QN.t1 9.14075
R22104 frontAnalog_v0p0p1_5.RSfetsym_0.QN.n2 frontAnalog_v0p0p1_5.RSfetsym_0.QN.n1 0.826818
R22105 frontAnalog_v0p0p1_5.RSfetsym_0.QN frontAnalog_v0p0p1_5.RSfetsym_0.QN.n0 0.74645
R22106 frontAnalog_v0p0p1_5.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_5.RSfetsym_0.QN.n3 0.249509
R22107 frontAnalog_v0p0p1_5.RSfetsym_0.QN.n3 frontAnalog_v0p0p1_5.RSfetsym_0.QN.n2 0.0968646
R22108 VV11.n0 VV11.t17 167.365
R22109 VV11.n0 VV11.t16 92.4496
R22110 VV11.n1 VV11.n0 2.07493
R22111 VV11.n17 VV11 0.5175
R22112 VV11 VV11.n17 0.38825
R22113 VV11.n15 VV11.n14 0.141409
R22114 VV11.n13 VV11.n12 0.141409
R22115 VV11.n11 VV11.n10 0.141409
R22116 VV11.n9 VV11.n8 0.141409
R22117 VV11.n7 VV11.n6 0.141409
R22118 VV11.n5 VV11.n4 0.141409
R22119 VV11.n3 VV11.n2 0.141409
R22120 VV11.n1 VV11 0.12425
R22121 VV11 VV11.n16 0.104098
R22122 VV11 VV11.n1 0.0314375
R22123 VV11.n17 VV11 0.00833333
R22124 VV11.n17 VV11 0.006375
R22125 VV11.n2 VV11.t15 0.000729415
R22126 VV11.n16 VV11.n15 0.000727273
R22127 VV11.n14 VV11.n13 0.000727273
R22128 VV11.n12 VV11.n11 0.000727273
R22129 VV11.n10 VV11.n9 0.000727273
R22130 VV11.n8 VV11.n7 0.000727273
R22131 VV11.n6 VV11.n5 0.000727273
R22132 VV11.n4 VV11.n3 0.000727273
R22133 VV11.n3 VV11.t4 0.000502142
R22134 VV11.n5 VV11.t12 0.000502142
R22135 VV11.n7 VV11.t6 0.000502142
R22136 VV11.n9 VV11.t1 0.000502142
R22137 VV11.n11 VV11.t10 0.000502142
R22138 VV11.n13 VV11.t3 0.000502142
R22139 VV11.n15 VV11.t9 0.000502142
R22140 VV11.n16 VV11.t11 0.000502142
R22141 VV11.n14 VV11.t5 0.000502142
R22142 VV11.n12 VV11.t0 0.000502142
R22143 VV11.n10 VV11.t14 0.000502142
R22144 VV11.n8 VV11.t8 0.000502142
R22145 VV11.n6 VV11.t13 0.000502142
R22146 VV11.n4 VV11.t2 0.000502142
R22147 VV11.n2 VV11.t7 0.000502142
R22148 VV10.n0 VV10.t16 167.365
R22149 VV10.n0 VV10.t17 92.4496
R22150 VV10.n1 VV10.n0 2.07493
R22151 VV10.n10 VV10 0.474417
R22152 VV10 VV10.n10 0.355937
R22153 VV10.n9 VV10.n8 0.141636
R22154 VV10.n8 VV10.n7 0.141636
R22155 VV10.n7 VV10.n6 0.141636
R22156 VV10.n6 VV10.n5 0.141636
R22157 VV10.n5 VV10.n4 0.141636
R22158 VV10.n4 VV10.n3 0.141636
R22159 VV10.n3 VV10.n2 0.141636
R22160 VV10.n1 VV10 0.12425
R22161 VV10 VV10.n9 0.104326
R22162 VV10 VV10.n1 0.028
R22163 VV10.n10 VV10 0.00833333
R22164 VV10.n10 VV10 0.006375
R22165 VV10.n2 VV10.t15 0.000502142
R22166 VV10.n3 VV10.t7 0.000502142
R22167 VV10.n4 VV10.t0 0.000502142
R22168 VV10.n5 VV10.t2 0.000502142
R22169 VV10.n6 VV10.t5 0.000502142
R22170 VV10.n7 VV10.t13 0.000502142
R22171 VV10.n8 VV10.t11 0.000502142
R22172 VV10.n9 VV10.t14 0.000502142
R22173 VV10.n9 VV10.t8 0.000502142
R22174 VV10.n8 VV10.t3 0.000502142
R22175 VV10.n7 VV10.t9 0.000502142
R22176 VV10.n6 VV10.t1 0.000502142
R22177 VV10.n5 VV10.t6 0.000502142
R22178 VV10.n4 VV10.t10 0.000502142
R22179 VV10.n3 VV10.t4 0.000502142
R22180 VV10.n2 VV10.t12 0.000502142
R22181 VV2.n0 VV2.t16 167.365
R22182 VV2.n0 VV2.t17 92.4488
R22183 VV2.n1 VV2.n0 2.07493
R22184 VV2.n17 VV2 0.64675
R22185 VV2 VV2.n17 0.485188
R22186 VV2.n15 VV2.n14 0.141409
R22187 VV2.n13 VV2.n12 0.141409
R22188 VV2.n11 VV2.n10 0.141409
R22189 VV2.n9 VV2.n8 0.141409
R22190 VV2.n7 VV2.n6 0.141409
R22191 VV2.n5 VV2.n4 0.141409
R22192 VV2.n3 VV2.n2 0.141409
R22193 VV2.n1 VV2 0.12425
R22194 VV2 VV2.n16 0.0968068
R22195 VV2 VV2.n1 0.028
R22196 VV2.n17 VV2 0.00833333
R22197 VV2.n17 VV2 0.006375
R22198 VV2.n2 VV2.t7 0.000729415
R22199 VV2.n16 VV2.n15 0.000727273
R22200 VV2.n14 VV2.n13 0.000727273
R22201 VV2.n12 VV2.n11 0.000727273
R22202 VV2.n10 VV2.n9 0.000727273
R22203 VV2.n8 VV2.n7 0.000727273
R22204 VV2.n6 VV2.n5 0.000727273
R22205 VV2.n4 VV2.n3 0.000727273
R22206 VV2.n4 VV2.t11 0.000502142
R22207 VV2.n6 VV2.t1 0.000502142
R22208 VV2.n8 VV2.t8 0.000502142
R22209 VV2.n10 VV2.t0 0.000502142
R22210 VV2.n12 VV2.t14 0.000502142
R22211 VV2.n14 VV2.t12 0.000502142
R22212 VV2.n16 VV2.t4 0.000502142
R22213 VV2.n3 VV2.t13 0.000502142
R22214 VV2.n5 VV2.t3 0.000502142
R22215 VV2.n7 VV2.t9 0.000502142
R22216 VV2.n9 VV2.t6 0.000502142
R22217 VV2.n11 VV2.t15 0.000502142
R22218 VV2.n13 VV2.t5 0.000502142
R22219 VV2.n15 VV2.t10 0.000502142
R22220 VV2.n2 VV2.t2 0.000502142
R22221 VV1.n0 VV1.t17 167.365
R22222 VV1.n0 VV1.t16 92.4488
R22223 VV1.n1 VV1.n0 2.07493
R22224 VV1.n10 VV1 0.8277
R22225 VV1 VV1.n10 0.591357
R22226 VV1.n9 VV1.n8 0.141636
R22227 VV1.n8 VV1.n7 0.141636
R22228 VV1.n7 VV1.n6 0.141636
R22229 VV1.n6 VV1.n5 0.141636
R22230 VV1.n5 VV1.n4 0.141636
R22231 VV1.n4 VV1.n3 0.141636
R22232 VV1.n3 VV1.n2 0.141636
R22233 VV1.n1 VV1 0.12425
R22234 VV1 VV1.n9 0.0980758
R22235 VV1 VV1.n1 0.0314375
R22236 VV1.n10 VV1 0.0099
R22237 VV1.n10 VV1 0.00721429
R22238 VV1.n3 VV1.t14 0.000502142
R22239 VV1.n4 VV1.t2 0.000502142
R22240 VV1.n5 VV1.t11 0.000502142
R22241 VV1.n6 VV1.t4 0.000502142
R22242 VV1.n7 VV1.t15 0.000502142
R22243 VV1.n8 VV1.t3 0.000502142
R22244 VV1.n9 VV1.t12 0.000502142
R22245 VV1.n2 VV1.t6 0.000502142
R22246 VV1.n3 VV1.t9 0.000502142
R22247 VV1.n4 VV1.t10 0.000502142
R22248 VV1.n5 VV1.t7 0.000502142
R22249 VV1.n6 VV1.t13 0.000502142
R22250 VV1.n7 VV1.t1 0.000502142
R22251 VV1.n8 VV1.t0 0.000502142
R22252 VV1.n9 VV1.t8 0.000502142
R22253 VV1.n2 VV1.t5 0.000502142
R22254 I0.n0 I0.t5 196.549
R22255 I0.n0 I0.t7 148.35
R22256 I0.n4 I0.t8 117.314
R22257 I0.n4 I0.t6 110.853
R22258 I0.n6 I0.t1 17.6181
R22259 I0.n7 I0.t0 14.2865
R22260 I0.n9 I0.t2 14.283
R22261 I0.n9 I0.t3 14.283
R22262 I0 I0.n12 9.77614
R22263 I0.n1 I0.n0 9.49592
R22264 I0.n11 I0.t4 8.77744
R22265 I0.n2 I0.n1 7.58085
R22266 I0.n1 I0 6.44187
R22267 I0.n3 I0.n2 2.50858
R22268 I0.n11 I0.n10 1.20426
R22269 I0.n2 I0 0.88934
R22270 I0.n12 I0.n11 0.32511
R22271 I0.n7 I0.n6 0.314673
R22272 I0.n8 I0.n7 0.299251
R22273 I0.n13 I0 0.204167
R22274 I0.n3 I0 0.2005
R22275 I0 I0.n3 0.1932
R22276 I0.n5 I0.n4 0.159555
R22277 I0 I0.n13 0.15325
R22278 I0.n10 I0.n9 0.106617
R22279 I0.n8 I0.n5 0.0796167
R22280 I0.n10 I0.n8 0.0480595
R22281 I0.n12 I0 0.046937
R22282 I0.n13 I0 0.0161667
R22283 I0.n13 I0 0.01225
R22284 I0.n6 I0.n5 0.000504658
R22285 I2.n6 I2.t5 323.342
R22286 I2.n0 I2.t9 228.927
R22287 I2.n3 I2.t7 196.549
R22288 I2.n6 I2.t8 194.809
R22289 I2.n0 I2.t6 159.391
R22290 I2.n3 I2.t11 148.35
R22291 I2.n10 I2.t12 117.314
R22292 I2.n10 I2.t10 110.853
R22293 I2.n7 I2.n6 76.0005
R22294 I2.n4 I2.n3 76.0005
R22295 I2.n8 I2.n7 29.2624
R22296 I2.n12 I2.t0 17.6181
R22297 I2.n13 I2.t4 14.2865
R22298 I2.n15 I2.t1 14.283
R22299 I2.n15 I2.t2 14.283
R22300 I2.n5 I2 9.11
R22301 I2.n17 I2.t3 8.77744
R22302 I2.n1 I2.n0 8.68501
R22303 I2 I2.n18 7.11948
R22304 I2.n4 I2 5.78114
R22305 I2.n2 I2.n1 4.26764
R22306 I2 I2.n4 3.71663
R22307 I2.n1 I2 1.99697
R22308 I2.n7 I2 1.92927
R22309 I2.n8 I2.n5 1.79514
R22310 I2.n17 I2.n16 1.20426
R22311 I2.n5 I2.n2 0.570143
R22312 I2.n19 I2 0.360833
R22313 I2 I2.n9 0.349867
R22314 I2.n18 I2.n17 0.32511
R22315 I2.n13 I2.n12 0.314673
R22316 I2.n14 I2.n13 0.299251
R22317 I2 I2.n19 0.27075
R22318 I2.n9 I2.n8 0.226885
R22319 I2.n2 I2 0.221483
R22320 I2.n9 I2 0.20675
R22321 I2.n11 I2.n10 0.159555
R22322 I2.n16 I2.n15 0.106617
R22323 I2.n14 I2.n11 0.0796167
R22324 I2.n16 I2.n14 0.0480595
R22325 I2.n18 I2 0.046937
R22326 I2.n19 I2 0.0161667
R22327 I2.n19 I2 0.01225
R22328 I2.n12 I2.n11 0.000504658
R22329 OUT1.n122 OUT1.n120 145.809
R22330 OUT1.n65 OUT1.n63 145.809
R22331 OUT1.n25 OUT1.n23 145.809
R22332 OUT1.n102 OUT1.n100 145.808
R22333 OUT1.n65 OUT1.n64 107.409
R22334 OUT1.n67 OUT1.n66 107.409
R22335 OUT1.n69 OUT1.n68 107.409
R22336 OUT1.n71 OUT1.n70 107.409
R22337 OUT1.n73 OUT1.n72 107.409
R22338 OUT1.n75 OUT1.n74 107.409
R22339 OUT1.n25 OUT1.n24 107.409
R22340 OUT1.n27 OUT1.n26 107.409
R22341 OUT1.n29 OUT1.n28 107.409
R22342 OUT1.n31 OUT1.n30 107.409
R22343 OUT1.n33 OUT1.n32 107.409
R22344 OUT1.n35 OUT1.n34 107.409
R22345 OUT1.n122 OUT1.n121 107.407
R22346 OUT1.n124 OUT1.n123 107.407
R22347 OUT1.n126 OUT1.n125 107.407
R22348 OUT1.n128 OUT1.n127 107.407
R22349 OUT1.n130 OUT1.n129 107.407
R22350 OUT1.n132 OUT1.n131 107.407
R22351 OUT1.n102 OUT1.n101 107.407
R22352 OUT1.n104 OUT1.n103 107.407
R22353 OUT1.n106 OUT1.n105 107.407
R22354 OUT1.n108 OUT1.n107 107.407
R22355 OUT1.n110 OUT1.n109 107.407
R22356 OUT1.n112 OUT1.n111 107.407
R22357 OUT1.n138 OUT1.n136 87.1779
R22358 OUT1.n83 OUT1.n81 87.1779
R22359 OUT1.n44 OUT1.n42 87.1779
R22360 OUT1.n4 OUT1.n2 87.1779
R22361 OUT1.n54 OUT1.n53 52.82
R22362 OUT1.n14 OUT1.n13 52.82
R22363 OUT1.n138 OUT1.n137 52.82
R22364 OUT1.n140 OUT1.n139 52.82
R22365 OUT1.n142 OUT1.n141 52.82
R22366 OUT1.n144 OUT1.n143 52.82
R22367 OUT1.n146 OUT1.n145 52.82
R22368 OUT1.n148 OUT1.n147 52.82
R22369 OUT1.n83 OUT1.n82 52.82
R22370 OUT1.n85 OUT1.n84 52.82
R22371 OUT1.n87 OUT1.n86 52.82
R22372 OUT1.n89 OUT1.n88 52.82
R22373 OUT1.n91 OUT1.n90 52.82
R22374 OUT1.n93 OUT1.n92 52.82
R22375 OUT1.n44 OUT1.n43 52.82
R22376 OUT1.n46 OUT1.n45 52.82
R22377 OUT1.n48 OUT1.n47 52.82
R22378 OUT1.n50 OUT1.n49 52.82
R22379 OUT1.n52 OUT1.n51 52.82
R22380 OUT1.n4 OUT1.n3 52.82
R22381 OUT1.n6 OUT1.n5 52.82
R22382 OUT1.n8 OUT1.n7 52.82
R22383 OUT1.n10 OUT1.n9 52.82
R22384 OUT1.n12 OUT1.n11 52.82
R22385 OUT1 OUT1.n149 51.0745
R22386 OUT1 OUT1.n94 51.0745
R22387 OUT1.n124 OUT1.n122 38.4005
R22388 OUT1.n126 OUT1.n124 38.4005
R22389 OUT1.n128 OUT1.n126 38.4005
R22390 OUT1.n130 OUT1.n128 38.4005
R22391 OUT1.n132 OUT1.n130 38.4005
R22392 OUT1.n133 OUT1.n132 38.4005
R22393 OUT1.n104 OUT1.n102 38.4005
R22394 OUT1.n106 OUT1.n104 38.4005
R22395 OUT1.n108 OUT1.n106 38.4005
R22396 OUT1.n110 OUT1.n108 38.4005
R22397 OUT1.n112 OUT1.n110 38.4005
R22398 OUT1.n113 OUT1.n112 38.4005
R22399 OUT1.n67 OUT1.n65 38.4005
R22400 OUT1.n69 OUT1.n67 38.4005
R22401 OUT1.n71 OUT1.n69 38.4005
R22402 OUT1.n73 OUT1.n71 38.4005
R22403 OUT1.n75 OUT1.n73 38.4005
R22404 OUT1.n76 OUT1.n75 38.4005
R22405 OUT1.n27 OUT1.n25 38.4005
R22406 OUT1.n29 OUT1.n27 38.4005
R22407 OUT1.n31 OUT1.n29 38.4005
R22408 OUT1.n33 OUT1.n31 38.4005
R22409 OUT1.n35 OUT1.n33 38.4005
R22410 OUT1.n36 OUT1.n35 38.4005
R22411 OUT1.n140 OUT1.n138 34.3584
R22412 OUT1.n142 OUT1.n140 34.3584
R22413 OUT1.n144 OUT1.n142 34.3584
R22414 OUT1.n146 OUT1.n144 34.3584
R22415 OUT1.n148 OUT1.n146 34.3584
R22416 OUT1.n150 OUT1.n148 34.3584
R22417 OUT1.n85 OUT1.n83 34.3584
R22418 OUT1.n87 OUT1.n85 34.3584
R22419 OUT1.n89 OUT1.n87 34.3584
R22420 OUT1.n91 OUT1.n89 34.3584
R22421 OUT1.n93 OUT1.n91 34.3584
R22422 OUT1.n95 OUT1.n93 34.3584
R22423 OUT1.n46 OUT1.n44 34.3584
R22424 OUT1.n48 OUT1.n46 34.3584
R22425 OUT1.n50 OUT1.n48 34.3584
R22426 OUT1.n52 OUT1.n50 34.3584
R22427 OUT1.n54 OUT1.n52 34.3584
R22428 OUT1.n58 OUT1.n54 34.3584
R22429 OUT1.n6 OUT1.n4 34.3584
R22430 OUT1.n8 OUT1.n6 34.3584
R22431 OUT1.n10 OUT1.n8 34.3584
R22432 OUT1.n12 OUT1.n10 34.3584
R22433 OUT1.n14 OUT1.n12 34.3584
R22434 OUT1.n18 OUT1.n14 34.3584
R22435 OUT1.n118 OUT1.t99 26.5955
R22436 OUT1.n118 OUT1.t112 26.5955
R22437 OUT1.n120 OUT1.t97 26.5955
R22438 OUT1.n120 OUT1.t69 26.5955
R22439 OUT1.n121 OUT1.t119 26.5955
R22440 OUT1.n121 OUT1.t85 26.5955
R22441 OUT1.n123 OUT1.t64 26.5955
R22442 OUT1.n123 OUT1.t105 26.5955
R22443 OUT1.n125 OUT1.t75 26.5955
R22444 OUT1.n125 OUT1.t93 26.5955
R22445 OUT1.n127 OUT1.t91 26.5955
R22446 OUT1.n127 OUT1.t108 26.5955
R22447 OUT1.n129 OUT1.t114 26.5955
R22448 OUT1.n129 OUT1.t80 26.5955
R22449 OUT1.n131 OUT1.t125 26.5955
R22450 OUT1.n131 OUT1.t101 26.5955
R22451 OUT1.n99 OUT1.t124 26.5955
R22452 OUT1.n99 OUT1.t89 26.5955
R22453 OUT1.n100 OUT1.t79 26.5955
R22454 OUT1.n100 OUT1.t88 26.5955
R22455 OUT1.n101 OUT1.t95 26.5955
R22456 OUT1.n101 OUT1.t68 26.5955
R22457 OUT1.n103 OUT1.t110 26.5955
R22458 OUT1.n103 OUT1.t82 26.5955
R22459 OUT1.n105 OUT1.t81 26.5955
R22460 OUT1.n105 OUT1.t94 26.5955
R22461 OUT1.n107 OUT1.t102 26.5955
R22462 OUT1.n107 OUT1.t116 26.5955
R22463 OUT1.n109 OUT1.t115 26.5955
R22464 OUT1.n109 OUT1.t70 26.5955
R22465 OUT1.n111 OUT1.t104 26.5955
R22466 OUT1.n111 OUT1.t72 26.5955
R22467 OUT1.n62 OUT1.t66 26.5955
R22468 OUT1.n62 OUT1.t100 26.5955
R22469 OUT1.n63 OUT1.t86 26.5955
R22470 OUT1.n63 OUT1.t98 26.5955
R22471 OUT1.n64 OUT1.t96 26.5955
R22472 OUT1.n64 OUT1.t120 26.5955
R22473 OUT1.n66 OUT1.t117 26.5955
R22474 OUT1.n66 OUT1.t83 26.5955
R22475 OUT1.n68 OUT1.t109 26.5955
R22476 OUT1.n68 OUT1.t76 26.5955
R22477 OUT1.n70 OUT1.t74 26.5955
R22478 OUT1.n70 OUT1.t92 26.5955
R22479 OUT1.n72 OUT1.t90 26.5955
R22480 OUT1.n72 OUT1.t107 26.5955
R22481 OUT1.n74 OUT1.t113 26.5955
R22482 OUT1.n74 OUT1.t126 26.5955
R22483 OUT1.n22 OUT1.t65 26.5955
R22484 OUT1.n22 OUT1.t78 26.5955
R22485 OUT1.n23 OUT1.t84 26.5955
R22486 OUT1.n23 OUT1.t106 26.5955
R22487 OUT1.n24 OUT1.t103 26.5955
R22488 OUT1.n24 OUT1.t118 26.5955
R22489 OUT1.n26 OUT1.t123 26.5955
R22490 OUT1.n26 OUT1.t71 26.5955
R22491 OUT1.n28 OUT1.t77 26.5955
R22492 OUT1.n28 OUT1.t111 26.5955
R22493 OUT1.n30 OUT1.t87 26.5955
R22494 OUT1.n30 OUT1.t122 26.5955
R22495 OUT1.n32 OUT1.t127 26.5955
R22496 OUT1.n32 OUT1.t73 26.5955
R22497 OUT1.n34 OUT1.t121 26.5955
R22498 OUT1.n34 OUT1.t67 26.5955
R22499 OUT1.n149 OUT1.t46 24.9236
R22500 OUT1.n149 OUT1.t59 24.9236
R22501 OUT1.n136 OUT1.t44 24.9236
R22502 OUT1.n136 OUT1.t16 24.9236
R22503 OUT1.n137 OUT1.t2 24.9236
R22504 OUT1.n137 OUT1.t32 24.9236
R22505 OUT1.n139 OUT1.t11 24.9236
R22506 OUT1.n139 OUT1.t52 24.9236
R22507 OUT1.n141 OUT1.t22 24.9236
R22508 OUT1.n141 OUT1.t40 24.9236
R22509 OUT1.n143 OUT1.t38 24.9236
R22510 OUT1.n143 OUT1.t55 24.9236
R22511 OUT1.n145 OUT1.t61 24.9236
R22512 OUT1.n145 OUT1.t27 24.9236
R22513 OUT1.n147 OUT1.t8 24.9236
R22514 OUT1.n147 OUT1.t48 24.9236
R22515 OUT1.n94 OUT1.t7 24.9236
R22516 OUT1.n94 OUT1.t36 24.9236
R22517 OUT1.n81 OUT1.t26 24.9236
R22518 OUT1.n81 OUT1.t35 24.9236
R22519 OUT1.n82 OUT1.t42 24.9236
R22520 OUT1.n82 OUT1.t15 24.9236
R22521 OUT1.n84 OUT1.t57 24.9236
R22522 OUT1.n84 OUT1.t29 24.9236
R22523 OUT1.n86 OUT1.t28 24.9236
R22524 OUT1.n86 OUT1.t41 24.9236
R22525 OUT1.n88 OUT1.t49 24.9236
R22526 OUT1.n88 OUT1.t63 24.9236
R22527 OUT1.n90 OUT1.t62 24.9236
R22528 OUT1.n90 OUT1.t17 24.9236
R22529 OUT1.n92 OUT1.t51 24.9236
R22530 OUT1.n92 OUT1.t19 24.9236
R22531 OUT1.n55 OUT1.t13 24.9236
R22532 OUT1.n55 OUT1.t47 24.9236
R22533 OUT1.n42 OUT1.t33 24.9236
R22534 OUT1.n42 OUT1.t45 24.9236
R22535 OUT1.n43 OUT1.t43 24.9236
R22536 OUT1.n43 OUT1.t3 24.9236
R22537 OUT1.n45 OUT1.t0 24.9236
R22538 OUT1.n45 OUT1.t30 24.9236
R22539 OUT1.n47 OUT1.t56 24.9236
R22540 OUT1.n47 OUT1.t24 24.9236
R22541 OUT1.n49 OUT1.t20 24.9236
R22542 OUT1.n49 OUT1.t39 24.9236
R22543 OUT1.n51 OUT1.t37 24.9236
R22544 OUT1.n51 OUT1.t54 24.9236
R22545 OUT1.n53 OUT1.t60 24.9236
R22546 OUT1.n53 OUT1.t9 24.9236
R22547 OUT1.n15 OUT1.t12 24.9236
R22548 OUT1.n15 OUT1.t25 24.9236
R22549 OUT1.n2 OUT1.t31 24.9236
R22550 OUT1.n2 OUT1.t53 24.9236
R22551 OUT1.n3 OUT1.t50 24.9236
R22552 OUT1.n3 OUT1.t1 24.9236
R22553 OUT1.n5 OUT1.t6 24.9236
R22554 OUT1.n5 OUT1.t18 24.9236
R22555 OUT1.n7 OUT1.t23 24.9236
R22556 OUT1.n7 OUT1.t58 24.9236
R22557 OUT1.n9 OUT1.t34 24.9236
R22558 OUT1.n9 OUT1.t5 24.9236
R22559 OUT1.n11 OUT1.t10 24.9236
R22560 OUT1.n11 OUT1.t21 24.9236
R22561 OUT1.n13 OUT1.t4 24.9236
R22562 OUT1.n13 OUT1.t14 24.9236
R22563 OUT1 OUT1.n150 11.4429
R22564 OUT1 OUT1.n95 11.4429
R22565 OUT1 OUT1.n58 11.4429
R22566 OUT1 OUT1.n18 11.4429
R22567 OUT1.n77 OUT1.n62 8.55024
R22568 OUT1.n37 OUT1.n22 8.55024
R22569 OUT1.n114 OUT1.n99 8.55024
R22570 OUT1.n119 OUT1.n118 8.46262
R22571 OUT1.n56 OUT1.n55 7.77479
R22572 OUT1.n16 OUT1.n15 7.77479
R22573 OUT1.n135 OUT1.n134 4.6505
R22574 OUT1.n151 OUT1 3.29747
R22575 OUT1.n96 OUT1 3.29747
R22576 OUT1.n78 OUT1.n77 3.20821
R22577 OUT1.n38 OUT1.n37 3.2082
R22578 OUT1.n115 OUT1.n114 3.20156
R22579 OUT1.n59 OUT1 3.10353
R22580 OUT1.n19 OUT1 3.10353
R22581 OUT1.n57 OUT1.n41 3.1005
R22582 OUT1.n17 OUT1.n1 3.1005
R22583 OUT1.n134 OUT1.n133 2.71565
R22584 OUT1.n114 OUT1.n113 2.32777
R22585 OUT1.n77 OUT1.n76 2.32777
R22586 OUT1.n37 OUT1.n36 2.32777
R22587 OUT1.n150 OUT1 1.74595
R22588 OUT1.n95 OUT1 1.74595
R22589 OUT1.n157 OUT1.n156 1.07337
R22590 OUT1.n58 OUT1.n57 0.970197
R22591 OUT1.n18 OUT1.n17 0.970197
R22592 OUT1.n158 OUT1.n157 0.69375
R22593 OUT1.n159 OUT1.n158 0.68905
R22594 OUT1.n56 OUT1 0.649449
R22595 OUT1.n16 OUT1 0.649449
R22596 OUT1.n158 OUT1.n79 0.414635
R22597 OUT1.n157 OUT1.n116 0.382465
R22598 OUT1.n159 OUT1.n39 0.368576
R22599 OUT1 OUT1.n159 0.279743
R22600 OUT1.n134 OUT1.n119 0.207197
R22601 OUT1.n79 OUT1.n78 0.157252
R22602 OUT1.n39 OUT1.n38 0.139891
R22603 OUT1.n156 OUT1.n155 0.139389
R22604 OUT1.n116 OUT1.n115 0.132946
R22605 OUT1.n57 OUT1.n56 0.118507
R22606 OUT1.n17 OUT1.n16 0.118507
R22607 OUT1.n60 OUT1.n41 0.111611
R22608 OUT1.n20 OUT1.n1 0.111611
R22609 OUT1.n154 OUT1.n135 0.0991111
R22610 OUT1.n154 OUT1.n152 0.0296667
R22611 OUT1.n135 OUT1.n117 0.0282778
R22612 OUT1.n98 OUT1.n97 0.0227222
R22613 OUT1.n61 OUT1.n60 0.0171667
R22614 OUT1.n21 OUT1.n20 0.0171667
R22615 OUT1.n115 OUT1.n98 0.00100004
R22616 OUT1.n38 OUT1.n21 0.00100004
R22617 OUT1.n78 OUT1.n61 0.00100004
R22618 OUT1.n152 OUT1.n151 0.000513563
R22619 OUT1.n97 OUT1.n96 0.000513563
R22620 OUT1.n60 OUT1.n59 0.000513218
R22621 OUT1.n20 OUT1.n19 0.000513218
R22622 OUT1.n98 OUT1.n80 0.00050517
R22623 OUT1.n154 OUT1.n153 0.000504838
R22624 OUT1.n61 OUT1.n40 0.000504838
R22625 OUT1.n21 OUT1.n0 0.000504838
R22626 OUT1.n155 OUT1.n154 0.000501713
R22627 frontAnalog_v0p0p1_8.RSfetsym_0.QN.n1 frontAnalog_v0p0p1_8.RSfetsym_0.QN.t5 117.511
R22628 frontAnalog_v0p0p1_8.RSfetsym_0.QN.n1 frontAnalog_v0p0p1_8.RSfetsym_0.QN.t6 110.698
R22629 frontAnalog_v0p0p1_8.RSfetsym_0.QN.n2 frontAnalog_v0p0p1_8.RSfetsym_0.QN.t2 19.1963
R22630 frontAnalog_v0p0p1_8.RSfetsym_0.QN.n3 frontAnalog_v0p0p1_8.RSfetsym_0.QN.t1 14.5206
R22631 frontAnalog_v0p0p1_8.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_8.RSfetsym_0.QN.t3 14.283
R22632 frontAnalog_v0p0p1_8.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_8.RSfetsym_0.QN.t4 14.283
R22633 frontAnalog_v0p0p1_8.RSfetsym_0.QN frontAnalog_v0p0p1_8.RSfetsym_0.QN.t0 9.14075
R22634 frontAnalog_v0p0p1_8.RSfetsym_0.QN.n2 frontAnalog_v0p0p1_8.RSfetsym_0.QN.n1 0.826818
R22635 frontAnalog_v0p0p1_8.RSfetsym_0.QN frontAnalog_v0p0p1_8.RSfetsym_0.QN.n0 0.74645
R22636 frontAnalog_v0p0p1_8.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_8.RSfetsym_0.QN.n3 0.249509
R22637 frontAnalog_v0p0p1_8.RSfetsym_0.QN.n3 frontAnalog_v0p0p1_8.RSfetsym_0.QN.n2 0.0968646
R22638 VV9.n0 VV9.t17 167.365
R22639 VV9.n0 VV9.t16 92.4496
R22640 VV9.n1 VV9.n0 2.07493
R22641 VV9.n10 VV9 0.431333
R22642 VV9 VV9.n10 0.287722
R22643 VV9.n9 VV9.n8 0.141636
R22644 VV9.n8 VV9.n7 0.141636
R22645 VV9.n7 VV9.n6 0.141636
R22646 VV9.n6 VV9.n5 0.141636
R22647 VV9.n5 VV9.n4 0.141636
R22648 VV9.n4 VV9.n3 0.141636
R22649 VV9.n3 VV9.n2 0.141636
R22650 VV9.n1 VV9 0.12425
R22651 VV9 VV9.n9 0.102242
R22652 VV9 VV9.n1 0.0314375
R22653 VV9.n10 VV9 0.00833333
R22654 VV9.n10 VV9 0.00572222
R22655 VV9.n2 VV9.t12 0.000502142
R22656 VV9.n3 VV9.t4 0.000502142
R22657 VV9.n4 VV9.t6 0.000502142
R22658 VV9.n5 VV9.t2 0.000502142
R22659 VV9.n6 VV9.t8 0.000502142
R22660 VV9.n7 VV9.t10 0.000502142
R22661 VV9.n8 VV9.t15 0.000502142
R22662 VV9.n9 VV9.t3 0.000502142
R22663 VV9.n9 VV9.t13 0.000502142
R22664 VV9.n8 VV9.t9 0.000502142
R22665 VV9.n7 VV9.t11 0.000502142
R22666 VV9.n6 VV9.t5 0.000502142
R22667 VV9.n5 VV9.t1 0.000502142
R22668 VV9.n4 VV9.t0 0.000502142
R22669 VV9.n3 VV9.t7 0.000502142
R22670 VV9.n2 VV9.t14 0.000502142
R22671 VV15.n0 VV15.t16 167.365
R22672 VV15.n0 VV15.t17 92.4496
R22673 VV15.n1 VV15.n0 2.07493
R22674 VV15.n9 VV15.n8 0.141636
R22675 VV15.n8 VV15.n7 0.141636
R22676 VV15.n7 VV15.n6 0.141636
R22677 VV15.n6 VV15.n5 0.141636
R22678 VV15.n5 VV15.n4 0.141636
R22679 VV15.n4 VV15.n3 0.141636
R22680 VV15.n3 VV15.n2 0.141636
R22681 VV15.n1 VV15 0.12425
R22682 VV15 VV15.n9 0.100159
R22683 VV15 VV15.n1 0.0358571
R22684 VV15.n2 VV15.t12 0.000502142
R22685 VV15.n3 VV15.t11 0.000502142
R22686 VV15.n4 VV15.t14 0.000502142
R22687 VV15.n5 VV15.t1 0.000502142
R22688 VV15.n6 VV15.t3 0.000502142
R22689 VV15.n7 VV15.t4 0.000502142
R22690 VV15.n8 VV15.t5 0.000502142
R22691 VV15.n9 VV15.t7 0.000502142
R22692 VV15.n9 VV15.t2 0.000502142
R22693 VV15.n8 VV15.t6 0.000502142
R22694 VV15.n7 VV15.t0 0.000502142
R22695 VV15.n6 VV15.t9 0.000502142
R22696 VV15.n5 VV15.t8 0.000502142
R22697 VV15.n4 VV15.t15 0.000502142
R22698 VV15.n3 VV15.t13 0.000502142
R22699 VV15.n2 VV15.t10 0.000502142
R22700 frontAnalog_v0p0p1_2.x63.A.n2 frontAnalog_v0p0p1_2.x63.A.t5 260.322
R22701 frontAnalog_v0p0p1_2.x63.A.n4 frontAnalog_v0p0p1_2.x63.A.t4 233.888
R22702 frontAnalog_v0p0p1_2.x63.A.n2 frontAnalog_v0p0p1_2.x63.A.t6 175.169
R22703 frontAnalog_v0p0p1_2.x63.A.n3 frontAnalog_v0p0p1_2.x63.A.t7 159.725
R22704 frontAnalog_v0p0p1_2.x63.A.n1 frontAnalog_v0p0p1_2.x63.A.t0 17.4109
R22705 frontAnalog_v0p0p1_2.x63.A.n0 frontAnalog_v0p0p1_2.x63.A.n2 9.75129
R22706 frontAnalog_v0p0p1_2.x63.A.n1 frontAnalog_v0p0p1_2.x63.A.t3 9.6037
R22707 frontAnalog_v0p0p1_2.x63.A.n0 frontAnalog_v0p0p1_2.x63.A 2.33338
R22708 frontAnalog_v0p0p1_2.x63.A.n5 frontAnalog_v0p0p1_2.x63.A.t2 8.40929
R22709 frontAnalog_v0p0p1_2.x63.A.n3 frontAnalog_v0p0p1_2.x63.A.t1 8.06629
R22710 frontAnalog_v0p0p1_2.x63.A.n4 frontAnalog_v0p0p1_2.x63.A.n3 1.73501
R22711 frontAnalog_v0p0p1_2.x63.A.n1 frontAnalog_v0p0p1_2.x63.A.n4 0.99025
R22712 frontAnalog_v0p0p1_2.x63.A.n5 frontAnalog_v0p0p1_2.x63.A.n1 0.853186
R22713 frontAnalog_v0p0p1_2.x63.A frontAnalog_v0p0p1_2.x63.A.n0 0.349517
R22714 frontAnalog_v0p0p1_2.x63.A frontAnalog_v0p0p1_2.x63.A.n5 0.24425
R22715 frontAnalog_v0p0p1_2.x65.A.n1 frontAnalog_v0p0p1_2.x65.A.t4 260.322
R22716 frontAnalog_v0p0p1_2.x65.A.n4 frontAnalog_v0p0p1_2.x65.A.t6 233.929
R22717 frontAnalog_v0p0p1_2.x65.A.n1 frontAnalog_v0p0p1_2.x65.A.t5 175.169
R22718 frontAnalog_v0p0p1_2.x65.A.n3 frontAnalog_v0p0p1_2.x65.A.t7 160.416
R22719 frontAnalog_v0p0p1_2.x65.A.n2 frontAnalog_v0p0p1_2.x65.A.t2 17.4109
R22720 frontAnalog_v0p0p1_2.x65.A.n2 frontAnalog_v0p0p1_2.x65.A.t3 10.2053
R22721 frontAnalog_v0p0p1_2.x65.A.n0 frontAnalog_v0p0p1_2.x65.A 2.78715
R22722 frontAnalog_v0p0p1_2.x65.A.n0 frontAnalog_v0p0p1_2.x65.A.n1 9.09103
R22723 frontAnalog_v0p0p1_2.x65.A.n6 frontAnalog_v0p0p1_2.x65.A.t1 7.94569
R22724 frontAnalog_v0p0p1_2.x65.A.n3 frontAnalog_v0p0p1_2.x65.A.t0 7.55846
R22725 frontAnalog_v0p0p1_2.x65.A.n5 frontAnalog_v0p0p1_2.x65.A.n4 1.4614
R22726 frontAnalog_v0p0p1_2.x65.A.n4 frontAnalog_v0p0p1_2.x65.A.n3 1.19626
R22727 frontAnalog_v0p0p1_2.x65.A.n6 frontAnalog_v0p0p1_2.x65.A.n5 0.836961
R22728 frontAnalog_v0p0p1_2.x65.A frontAnalog_v0p0p1_2.x65.A.n0 0.390342
R22729 frontAnalog_v0p0p1_2.x65.A.n5 frontAnalog_v0p0p1_2.x65.A.n2 0.154668
R22730 frontAnalog_v0p0p1_2.x65.A frontAnalog_v0p0p1_2.x65.A.n6 0.08175
R22731 frontAnalog_v0p0p1_15.RSfetsym_0.QN.n1 frontAnalog_v0p0p1_15.RSfetsym_0.QN.t6 117.511
R22732 frontAnalog_v0p0p1_15.RSfetsym_0.QN.n1 frontAnalog_v0p0p1_15.RSfetsym_0.QN.t5 110.698
R22733 frontAnalog_v0p0p1_15.RSfetsym_0.QN.n2 frontAnalog_v0p0p1_15.RSfetsym_0.QN.t2 19.1963
R22734 frontAnalog_v0p0p1_15.RSfetsym_0.QN.n3 frontAnalog_v0p0p1_15.RSfetsym_0.QN.t4 14.5206
R22735 frontAnalog_v0p0p1_15.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_15.RSfetsym_0.QN.t1 14.283
R22736 frontAnalog_v0p0p1_15.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_15.RSfetsym_0.QN.t0 14.283
R22737 frontAnalog_v0p0p1_15.RSfetsym_0.QN frontAnalog_v0p0p1_15.RSfetsym_0.QN.t3 9.14075
R22738 frontAnalog_v0p0p1_15.RSfetsym_0.QN.n2 frontAnalog_v0p0p1_15.RSfetsym_0.QN.n1 0.826818
R22739 frontAnalog_v0p0p1_15.RSfetsym_0.QN frontAnalog_v0p0p1_15.RSfetsym_0.QN.n0 0.74645
R22740 frontAnalog_v0p0p1_15.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_15.RSfetsym_0.QN.n3 0.249509
R22741 frontAnalog_v0p0p1_15.RSfetsym_0.QN.n3 frontAnalog_v0p0p1_15.RSfetsym_0.QN.n2 0.0968646
R22742 VV6.n0 VV6.t17 167.365
R22743 VV6.n0 VV6.t16 92.4488
R22744 VV6.n1 VV6.n0 2.07493
R22745 VV6.n10 VV6 0.501833
R22746 VV6 VV6.n10 0.3765
R22747 VV6.n9 VV6.n8 0.141636
R22748 VV6.n8 VV6.n7 0.141636
R22749 VV6.n7 VV6.n6 0.141636
R22750 VV6.n6 VV6.n5 0.141636
R22751 VV6.n5 VV6.n4 0.141636
R22752 VV6.n4 VV6.n3 0.141636
R22753 VV6.n3 VV6.n2 0.141636
R22754 VV6.n1 VV6 0.12425
R22755 VV6 VV6.n9 0.0991174
R22756 VV6 VV6.n1 0.0314375
R22757 VV6.n10 VV6 0.00833333
R22758 VV6.n10 VV6 0.006375
R22759 VV6.n3 VV6.t7 0.000502142
R22760 VV6.n4 VV6.t11 0.000502142
R22761 VV6.n5 VV6.t1 0.000502142
R22762 VV6.n6 VV6.t5 0.000502142
R22763 VV6.n7 VV6.t12 0.000502142
R22764 VV6.n8 VV6.t0 0.000502142
R22765 VV6.n9 VV6.t8 0.000502142
R22766 VV6.n2 VV6.t4 0.000502142
R22767 VV6.n3 VV6.t6 0.000502142
R22768 VV6.n4 VV6.t3 0.000502142
R22769 VV6.n5 VV6.t9 0.000502142
R22770 VV6.n6 VV6.t2 0.000502142
R22771 VV6.n7 VV6.t13 0.000502142
R22772 VV6.n8 VV6.t15 0.000502142
R22773 VV6.n9 VV6.t14 0.000502142
R22774 VV6.n2 VV6.t10 0.000502142
R22775 VV5.n0 VV5.t17 167.365
R22776 VV5.n0 VV5.t16 92.4488
R22777 VV5.n1 VV5.n0 2.07493
R22778 VV5.n10 VV5 0.537083
R22779 VV5 VV5.n10 0.402938
R22780 VV5.n9 VV5.n8 0.141636
R22781 VV5.n8 VV5.n7 0.141636
R22782 VV5.n7 VV5.n6 0.141636
R22783 VV5.n6 VV5.n5 0.141636
R22784 VV5.n5 VV5.n4 0.141636
R22785 VV5.n4 VV5.n3 0.141636
R22786 VV5.n3 VV5.n2 0.141636
R22787 VV5.n1 VV5 0.12425
R22788 VV5 VV5.n9 0.103284
R22789 VV5 VV5.n1 0.0314375
R22790 VV5.n10 VV5 0.00833333
R22791 VV5.n10 VV5 0.006375
R22792 VV5.n3 VV5.t7 0.000502142
R22793 VV5.n4 VV5.t3 0.000502142
R22794 VV5.n5 VV5.t9 0.000502142
R22795 VV5.n6 VV5.t2 0.000502142
R22796 VV5.n7 VV5.t11 0.000502142
R22797 VV5.n8 VV5.t13 0.000502142
R22798 VV5.n9 VV5.t12 0.000502142
R22799 VV5.n2 VV5.t6 0.000502142
R22800 VV5.n3 VV5.t0 0.000502142
R22801 VV5.n4 VV5.t8 0.000502142
R22802 VV5.n5 VV5.t10 0.000502142
R22803 VV5.n6 VV5.t1 0.000502142
R22804 VV5.n7 VV5.t14 0.000502142
R22805 VV5.n8 VV5.t5 0.000502142
R22806 VV5.n9 VV5.t15 0.000502142
R22807 VV5.n2 VV5.t4 0.000502142
R22808 I10.n6 I10.t12 323.342
R22809 I10.n0 I10.t11 228.927
R22810 I10.n3 I10.t6 196.549
R22811 I10.n6 I10.t10 194.809
R22812 I10.n0 I10.t8 159.391
R22813 I10.n3 I10.t9 148.35
R22814 I10.n10 I10.t7 117.314
R22815 I10.n10 I10.t5 110.852
R22816 I10.n7 I10.n6 76.0005
R22817 I10.n4 I10.n3 76.0005
R22818 I10.n8 I10.n7 29.3651
R22819 I10.n12 I10.t3 17.6181
R22820 I10.n13 I10.t0 14.2865
R22821 I10.n15 I10.t1 14.283
R22822 I10.n15 I10.t2 14.283
R22823 I10.n5 I10 9.11
R22824 I10.n17 I10.t4 8.77592
R22825 I10.n1 I10.n0 8.6846
R22826 I10.n4 I10 5.78114
R22827 I10.n2 I10.n1 4.26809
R22828 I10 I10.n4 3.71663
R22829 I10 I10.n18 2.22491
R22830 I10.n1 I10 1.99652
R22831 I10.n7 I10 1.92927
R22832 I10.n8 I10.n5 1.69246
R22833 I10.n17 I10.n16 1.20426
R22834 I10.n19 I10 0.760333
R22835 I10 I10.n9 0.7337
R22836 I10.n5 I10.n2 0.570143
R22837 I10 I10.n19 0.4564
R22838 I10.n18 I10.n17 0.336084
R22839 I10.n13 I10.n12 0.314673
R22840 I10.n14 I10.n13 0.300251
R22841 I10.n9 I10.n8 0.224535
R22842 I10.n2 I10 0.221483
R22843 I10.n9 I10 0.2005
R22844 I10.n11 I10.n10 0.159555
R22845 I10.n16 I10.n15 0.106617
R22846 I10.n14 I10.n11 0.0796167
R22847 I10.n16 I10.n14 0.0480595
R22848 I10.n19 I10 0.0161667
R22849 I10.n19 I10 0.0099
R22850 I10.n18 I10 0.00658123
R22851 I10.n12 I10.n11 0.000504658
R22852 frontAnalog_v0p0p1_6.RSfetsym_0.QN.n1 frontAnalog_v0p0p1_6.RSfetsym_0.QN.t6 117.511
R22853 frontAnalog_v0p0p1_6.RSfetsym_0.QN.n1 frontAnalog_v0p0p1_6.RSfetsym_0.QN.t5 110.698
R22854 frontAnalog_v0p0p1_6.RSfetsym_0.QN.n2 frontAnalog_v0p0p1_6.RSfetsym_0.QN.t0 19.1963
R22855 frontAnalog_v0p0p1_6.RSfetsym_0.QN.n3 frontAnalog_v0p0p1_6.RSfetsym_0.QN.t4 14.5206
R22856 frontAnalog_v0p0p1_6.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_6.RSfetsym_0.QN.t1 14.283
R22857 frontAnalog_v0p0p1_6.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_6.RSfetsym_0.QN.t2 14.283
R22858 frontAnalog_v0p0p1_6.RSfetsym_0.QN frontAnalog_v0p0p1_6.RSfetsym_0.QN.t3 9.14075
R22859 frontAnalog_v0p0p1_6.RSfetsym_0.QN.n2 frontAnalog_v0p0p1_6.RSfetsym_0.QN.n1 0.826818
R22860 frontAnalog_v0p0p1_6.RSfetsym_0.QN frontAnalog_v0p0p1_6.RSfetsym_0.QN.n0 0.74645
R22861 frontAnalog_v0p0p1_6.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_6.RSfetsym_0.QN.n3 0.249509
R22862 frontAnalog_v0p0p1_6.RSfetsym_0.QN.n3 frontAnalog_v0p0p1_6.RSfetsym_0.QN.n2 0.0968646
R22863 I13.t9 I13.t13 618.109
R22864 I13.n12 I13.t14 259.74
R22865 I13 I13.t9 253.56
R22866 I13.n0 I13.t11 228.899
R22867 I13.n19 I13.t6 180.286
R22868 I13.n0 I13.t10 159.411
R22869 I13.n12 I13.t8 157.083
R22870 I13.n26 I13.t5 117.314
R22871 I13.n20 I13.t7 111.091
R22872 I13.n26 I13.t12 110.852
R22873 I13.n23 I13 37.7071
R22874 I13.n28 I13.t1 17.6181
R22875 I13.n29 I13.t0 14.2865
R22876 I13.n31 I13.t2 14.283
R22877 I13.n31 I13.t3 14.283
R22878 I13.n21 I13.n20 9.3005
R22879 I13 I13.n11 9.3005
R22880 I13.n33 I13.t4 8.77592
R22881 I13.n22 I13.n21 7.80966
R22882 I13.n13 I13.n12 7.57248
R22883 I13.n1 I13.n0 7.36885
R22884 I13.n20 I13.n19 6.53562
R22885 I13 I13.n34 4.95588
R22886 I13.n13 I13 4.8645
R22887 I13.n3 I13.n2 3.46717
R22888 I13.n4 I13.n3 3.03286
R22889 I13.n18 I13.n17 2.32777
R22890 I13.n22 I13.n16 2.19001
R22891 I13.n17 I13 1.4966
R22892 I13.n33 I13.n32 1.20426
R22893 I13.n24 I13.n9 1.16836
R22894 I13.n23 I13.n22 1.07639
R22895 I13.n3 I13.n1 1.06717
R22896 I13.n2 I13 1.06717
R22897 I13 I13.n25 0.889055
R22898 I13.n9 I13.n8 0.71595
R22899 I13.n21 I13.n18 0.499201
R22900 I13.n25 I13.n24 0.458555
R22901 I13.n34 I13.n33 0.336084
R22902 I13.n29 I13.n28 0.314673
R22903 I13.n30 I13.n29 0.300251
R22904 I13.n9 I13 0.221483
R22905 I13.n25 I13 0.2005
R22906 I13.n24 I13.n23 0.192464
R22907 I13.n27 I13.n26 0.159555
R22908 I13.n32 I13.n31 0.106617
R22909 I13.n30 I13.n27 0.0796167
R22910 I13.n32 I13.n30 0.0480595
R22911 I13.n11 I13.n10 0.0301875
R22912 I13.n16 I13.n15 0.0205312
R22913 I13.n34 I13 0.00658123
R22914 I13.n6 I13.n5 0.00618182
R22915 I13.n5 I13.n4 0.00555107
R22916 I13.n7 I13.n6 0.00430477
R22917 I13.n15 I13.n14 0.00210765
R22918 I13.n14 I13.n13 0.00133438
R22919 I13.n8 I13.n7 0.00101192
R22920 I13.n14 I13.n10 0.00100001
R22921 I13.n28 I13.n27 0.000504658
R22922 frontAnalog_v0p0p1_10.IB.n0 frontAnalog_v0p0p1_10.IB.t1 182.794
R22923 frontAnalog_v0p0p1_10.IB.n1 frontAnalog_v0p0p1_10.IB.t12 91.7714
R22924 frontAnalog_v0p0p1_10.IB.n17 frontAnalog_v0p0p1_10.IB.t17 91.7714
R22925 frontAnalog_v0p0p1_10.IB.n16 frontAnalog_v0p0p1_10.IB.t14 91.7714
R22926 frontAnalog_v0p0p1_10.IB.n15 frontAnalog_v0p0p1_10.IB.t27 91.7714
R22927 frontAnalog_v0p0p1_10.IB.n14 frontAnalog_v0p0p1_10.IB.t21 91.7714
R22928 frontAnalog_v0p0p1_10.IB.n13 frontAnalog_v0p0p1_10.IB.t4 91.7714
R22929 frontAnalog_v0p0p1_10.IB.n12 frontAnalog_v0p0p1_10.IB.t31 91.7714
R22930 frontAnalog_v0p0p1_10.IB.n11 frontAnalog_v0p0p1_10.IB.t10 91.7714
R22931 frontAnalog_v0p0p1_10.IB.n10 frontAnalog_v0p0p1_10.IB.t7 91.7714
R22932 frontAnalog_v0p0p1_10.IB.n9 frontAnalog_v0p0p1_10.IB.t18 91.7714
R22933 frontAnalog_v0p0p1_10.IB.n8 frontAnalog_v0p0p1_10.IB.t15 91.7714
R22934 frontAnalog_v0p0p1_10.IB.n7 frontAnalog_v0p0p1_10.IB.t26 91.7714
R22935 frontAnalog_v0p0p1_10.IB.n6 frontAnalog_v0p0p1_10.IB.t22 91.7714
R22936 frontAnalog_v0p0p1_10.IB.n5 frontAnalog_v0p0p1_10.IB.t5 91.7714
R22937 frontAnalog_v0p0p1_10.IB.n4 frontAnalog_v0p0p1_10.IB.t32 91.7714
R22938 frontAnalog_v0p0p1_10.IB.n2 frontAnalog_v0p0p1_10.IB.t3 91.7714
R22939 frontAnalog_v0p0p1_10.IB.n17 frontAnalog_v0p0p1_10.IB.t28 91.3136
R22940 frontAnalog_v0p0p1_10.IB.n16 frontAnalog_v0p0p1_10.IB.t24 91.3136
R22941 frontAnalog_v0p0p1_10.IB.n15 frontAnalog_v0p0p1_10.IB.t6 91.3136
R22942 frontAnalog_v0p0p1_10.IB.n14 frontAnalog_v0p0p1_10.IB.t33 91.3136
R22943 frontAnalog_v0p0p1_10.IB.n13 frontAnalog_v0p0p1_10.IB.t13 91.3136
R22944 frontAnalog_v0p0p1_10.IB.n12 frontAnalog_v0p0p1_10.IB.t8 91.3136
R22945 frontAnalog_v0p0p1_10.IB.n11 frontAnalog_v0p0p1_10.IB.t20 91.3136
R22946 frontAnalog_v0p0p1_10.IB.n10 frontAnalog_v0p0p1_10.IB.t16 91.3136
R22947 frontAnalog_v0p0p1_10.IB.n9 frontAnalog_v0p0p1_10.IB.t30 91.3136
R22948 frontAnalog_v0p0p1_10.IB.n8 frontAnalog_v0p0p1_10.IB.t25 91.3136
R22949 frontAnalog_v0p0p1_10.IB.n7 frontAnalog_v0p0p1_10.IB.t19 91.3136
R22950 frontAnalog_v0p0p1_10.IB.n6 frontAnalog_v0p0p1_10.IB.t34 91.3136
R22951 frontAnalog_v0p0p1_10.IB.n5 frontAnalog_v0p0p1_10.IB.t29 91.3136
R22952 frontAnalog_v0p0p1_10.IB.n4 frontAnalog_v0p0p1_10.IB.t9 91.3136
R22953 frontAnalog_v0p0p1_10.IB.n2 frontAnalog_v0p0p1_10.IB.t11 91.3136
R22954 frontAnalog_v0p0p1_10.IB.n1 frontAnalog_v0p0p1_10.IB.t23 91.3136
R22955 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_10.IB.n17 45.9747
R22956 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_10.IB.n16 45.9747
R22957 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_10.IB.n15 45.9747
R22958 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_10.IB.n14 45.9747
R22959 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_10.IB.n13 45.9747
R22960 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_10.IB.n12 45.9747
R22961 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_10.IB.n11 45.9747
R22962 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_10.IB.n10 45.9747
R22963 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_10.IB.n9 45.9747
R22964 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_10.IB.n8 45.9747
R22965 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_10.IB.n7 45.9747
R22966 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_10.IB.n6 45.9747
R22967 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_10.IB.n5 45.9747
R22968 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_10.IB.n4 45.9747
R22969 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_10.IB.n2 45.9747
R22970 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_10.IB.n1 45.973
R22971 frontAnalog_v0p0p1_10.IB.n34 frontAnalog_v0p0p1_10.IB.t0 5.91044
R22972 frontAnalog_v0p0p1_10.IB.n32 frontAnalog_v0p0p1_10.IB.t2 4.35136
R22973 frontAnalog_v0p0p1_10.IB.n18 frontAnalog_v0p0p1_10.IB 1.53808
R22974 frontAnalog_v0p0p1_10.IB.n34 frontAnalog_v0p0p1_10.IB.n31 1.41054
R22975 frontAnalog_v0p0p1_10.IB.n3 frontAnalog_v0p0p1_10.IB 1.28321
R22976 frontAnalog_v0p0p1_10.IB.n29 frontAnalog_v0p0p1_10.IB 1.15021
R22977 frontAnalog_v0p0p1_10.IB.n28 frontAnalog_v0p0p1_10.IB 1.14904
R22978 frontAnalog_v0p0p1_10.IB.n26 frontAnalog_v0p0p1_10.IB 1.14883
R22979 frontAnalog_v0p0p1_10.IB.n30 frontAnalog_v0p0p1_10.IB 1.14802
R22980 frontAnalog_v0p0p1_10.IB.n19 frontAnalog_v0p0p1_10.IB 1.14536
R22981 frontAnalog_v0p0p1_10.IB.n25 frontAnalog_v0p0p1_10.IB 1.14495
R22982 frontAnalog_v0p0p1_10.IB.n27 frontAnalog_v0p0p1_10.IB 1.14447
R22983 frontAnalog_v0p0p1_10.IB.n21 frontAnalog_v0p0p1_10.IB 1.14439
R22984 frontAnalog_v0p0p1_10.IB.n22 frontAnalog_v0p0p1_10.IB 1.14419
R22985 frontAnalog_v0p0p1_10.IB.n24 frontAnalog_v0p0p1_10.IB 1.14189
R22986 frontAnalog_v0p0p1_10.IB.n23 frontAnalog_v0p0p1_10.IB 1.14114
R22987 frontAnalog_v0p0p1_10.IB.n18 frontAnalog_v0p0p1_10.IB 1.13988
R22988 frontAnalog_v0p0p1_10.IB.n20 frontAnalog_v0p0p1_10.IB 1.13929
R22989 frontAnalog_v0p0p1_10.IB.n3 frontAnalog_v0p0p1_10.IB 0.957022
R22990 frontAnalog_v0p0p1_10.IB.n33 frontAnalog_v0p0p1_10.IB.n32 0.807781
R22991 frontAnalog_v0p0p1_10.IB.n34 frontAnalog_v0p0p1_10.IB.n0 0.504831
R22992 frontAnalog_v0p0p1_10.IB.n30 frontAnalog_v0p0p1_10.IB.n29 0.399765
R22993 frontAnalog_v0p0p1_10.IB.n28 frontAnalog_v0p0p1_10.IB.n27 0.399029
R22994 frontAnalog_v0p0p1_10.IB.n25 frontAnalog_v0p0p1_10.IB.n24 0.399029
R22995 frontAnalog_v0p0p1_10.IB.n23 frontAnalog_v0p0p1_10.IB.n22 0.398294
R22996 frontAnalog_v0p0p1_10.IB.n21 frontAnalog_v0p0p1_10.IB.n20 0.398294
R22997 frontAnalog_v0p0p1_10.IB.n26 frontAnalog_v0p0p1_10.IB.n25 0.397559
R22998 frontAnalog_v0p0p1_10.IB.n22 frontAnalog_v0p0p1_10.IB.n21 0.396824
R22999 frontAnalog_v0p0p1_10.IB.n20 frontAnalog_v0p0p1_10.IB.n19 0.396824
R23000 frontAnalog_v0p0p1_10.IB.n19 frontAnalog_v0p0p1_10.IB.n18 0.396824
R23001 frontAnalog_v0p0p1_10.IB.n27 frontAnalog_v0p0p1_10.IB.n26 0.396088
R23002 frontAnalog_v0p0p1_10.IB.n24 frontAnalog_v0p0p1_10.IB.n23 0.396088
R23003 frontAnalog_v0p0p1_10.IB.n29 frontAnalog_v0p0p1_10.IB.n28 0.395353
R23004 frontAnalog_v0p0p1_10.IB.n31 frontAnalog_v0p0p1_10.IB.n30 0.249029
R23005 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_10.IB.n34 0.168769
R23006 frontAnalog_v0p0p1_10.IB.n31 frontAnalog_v0p0p1_10.IB.n3 0.151971
R23007 frontAnalog_v0p0p1_10.IB.n0 frontAnalog_v0p0p1_10.IB.n33 0.0762967
R23008 VV14.n0 VV14.t17 167.365
R23009 VV14.n0 VV14.t16 92.4496
R23010 VV14.n1 VV14.n0 2.07493
R23011 VV14.n10 VV14 0.638917
R23012 VV14 VV14.n10 0.479312
R23013 VV14.n9 VV14.n8 0.141636
R23014 VV14.n8 VV14.n7 0.141636
R23015 VV14.n7 VV14.n6 0.141636
R23016 VV14.n6 VV14.n5 0.141636
R23017 VV14.n5 VV14.n4 0.141636
R23018 VV14.n4 VV14.n3 0.141636
R23019 VV14.n3 VV14.n2 0.141636
R23020 VV14.n1 VV14 0.12425
R23021 VV14 VV14.n9 0.102242
R23022 VV14 VV14.n1 0.0358571
R23023 VV14.n10 VV14 0.00833333
R23024 VV14.n10 VV14 0.006375
R23025 VV14.n2 VV14.t9 0.000502142
R23026 VV14.n3 VV14.t10 0.000502142
R23027 VV14.n4 VV14.t6 0.000502142
R23028 VV14.n5 VV14.t11 0.000502142
R23029 VV14.n6 VV14.t1 0.000502142
R23030 VV14.n7 VV14.t5 0.000502142
R23031 VV14.n8 VV14.t12 0.000502142
R23032 VV14.n9 VV14.t8 0.000502142
R23033 VV14.n9 VV14.t7 0.000502142
R23034 VV14.n8 VV14.t4 0.000502142
R23035 VV14.n7 VV14.t3 0.000502142
R23036 VV14.n6 VV14.t2 0.000502142
R23037 VV14.n5 VV14.t0 0.000502142
R23038 VV14.n4 VV14.t15 0.000502142
R23039 VV14.n3 VV14.t13 0.000502142
R23040 VV14.n2 VV14.t14 0.000502142
R23041 VV13.n0 VV13.t16 167.365
R23042 VV13.n0 VV13.t17 92.4496
R23043 VV13.n1 VV13.n0 2.07493
R23044 VV13.n10 VV13 0.59975
R23045 VV13 VV13.n10 0.449937
R23046 VV13.n9 VV13.n8 0.141636
R23047 VV13.n8 VV13.n7 0.141636
R23048 VV13.n7 VV13.n6 0.141636
R23049 VV13.n6 VV13.n5 0.141636
R23050 VV13.n5 VV13.n4 0.141636
R23051 VV13.n4 VV13.n3 0.141636
R23052 VV13.n3 VV13.n2 0.141636
R23053 VV13.n1 VV13 0.12425
R23054 VV13 VV13.n9 0.0991174
R23055 VV13 VV13.n1 0.0314375
R23056 VV13.n10 VV13 0.00833333
R23057 VV13.n10 VV13 0.006375
R23058 VV13.n2 VV13.t6 0.000502142
R23059 VV13.n3 VV13.t4 0.000502142
R23060 VV13.n4 VV13.t1 0.000502142
R23061 VV13.n5 VV13.t15 0.000502142
R23062 VV13.n6 VV13.t8 0.000502142
R23063 VV13.n7 VV13.t13 0.000502142
R23064 VV13.n8 VV13.t9 0.000502142
R23065 VV13.n9 VV13.t2 0.000502142
R23066 VV13.n9 VV13.t7 0.000502142
R23067 VV13.n8 VV13.t14 0.000502142
R23068 VV13.n7 VV13.t3 0.000502142
R23069 VV13.n6 VV13.t0 0.000502142
R23070 VV13.n5 VV13.t12 0.000502142
R23071 VV13.n4 VV13.t5 0.000502142
R23072 VV13.n3 VV13.t11 0.000502142
R23073 VV13.n2 VV13.t10 0.000502142
R23074 VIN.n3 VIN.t19 167.326
R23075 VIN.n18 VIN.t11 167.326
R23076 VIN.n17 VIN.t5 167.326
R23077 VIN.n16 VIN.t20 167.326
R23078 VIN.n15 VIN.t15 167.326
R23079 VIN.n14 VIN.t26 167.326
R23080 VIN.n13 VIN.t23 167.326
R23081 VIN.n12 VIN.t1 167.326
R23082 VIN.n11 VIN.t28 167.326
R23083 VIN.n10 VIN.t13 167.326
R23084 VIN.n9 VIN.t6 167.326
R23085 VIN.n8 VIN.t31 167.326
R23086 VIN.n7 VIN.t16 167.326
R23087 VIN.n6 VIN.t10 167.326
R23088 VIN.n5 VIN.t24 167.326
R23089 VIN.n0 VIN.t4 167.326
R23090 VIN.n3 VIN.t17 92.4649
R23091 VIN.n18 VIN.t7 92.4649
R23092 VIN.n17 VIN.t0 92.4649
R23093 VIN.n16 VIN.t18 92.4649
R23094 VIN.n15 VIN.t12 92.4649
R23095 VIN.n14 VIN.t25 92.4649
R23096 VIN.n13 VIN.t21 92.4649
R23097 VIN.n12 VIN.t30 92.4649
R23098 VIN.n11 VIN.t27 92.4649
R23099 VIN.n10 VIN.t9 92.4649
R23100 VIN.n9 VIN.t2 92.4649
R23101 VIN.n8 VIN.t29 92.4649
R23102 VIN.n7 VIN.t14 92.4649
R23103 VIN.n6 VIN.t8 92.4649
R23104 VIN.n5 VIN.t22 92.4649
R23105 VIN.n0 VIN.t3 92.4649
R23106 VIN.n1 VIN 4.6255
R23107 VIN.n2 VIN.n1 1.6255
R23108 VIN VIN.n18 1.49913
R23109 VIN VIN.n17 1.49913
R23110 VIN VIN.n16 1.49913
R23111 VIN VIN.n15 1.49913
R23112 VIN VIN.n14 1.49913
R23113 VIN VIN.n13 1.49913
R23114 VIN VIN.n12 1.49913
R23115 VIN VIN.n11 1.49913
R23116 VIN VIN.n10 1.49913
R23117 VIN VIN.n9 1.49913
R23118 VIN VIN.n8 1.49913
R23119 VIN VIN.n7 1.49913
R23120 VIN VIN.n5 1.49913
R23121 VIN.n1 VIN.n0 1.49913
R23122 VIN VIN.n3 1.46056
R23123 VIN VIN.n6 1.46056
R23124 VIN.n19 VIN 1.04323
R23125 VIN.n32 VIN.n4 0.573417
R23126 VIN.n32 VIN.n31 0.563
R23127 VIN.n31 VIN.n30 0.563
R23128 VIN.n30 VIN.n29 0.563
R23129 VIN.n29 VIN.n28 0.563
R23130 VIN.n28 VIN.n27 0.563
R23131 VIN.n27 VIN.n26 0.563
R23132 VIN.n26 VIN.n25 0.563
R23133 VIN.n25 VIN.n24 0.563
R23134 VIN.n24 VIN.n23 0.563
R23135 VIN.n23 VIN.n22 0.563
R23136 VIN.n22 VIN.n21 0.563
R23137 VIN.n21 VIN.n20 0.563
R23138 VIN.n20 VIN.n19 0.563
R23139 VIN.n4 VIN 0.517333
R23140 VIN.n25 VIN 0.496386
R23141 VIN.n20 VIN 0.484963
R23142 VIN.n22 VIN 0.484963
R23143 VIN.n23 VIN 0.484963
R23144 VIN.n24 VIN 0.484963
R23145 VIN.n26 VIN 0.484963
R23146 VIN.n27 VIN 0.484963
R23147 VIN.n28 VIN 0.484963
R23148 VIN.n21 VIN 0.480732
R23149 VIN.n29 VIN 0.480732
R23150 VIN.n33 VIN.n32 0.47425
R23151 VIN.n19 VIN 0.473007
R23152 VIN.n31 VIN 0.473007
R23153 VIN.n30 VIN 0.45875
R23154 VIN.n2 VIN 0.316289
R23155 VIN.n4 VIN 0.169571
R23156 VIN VIN.n33 0.01
R23157 VIN.n33 VIN.n2 0.00707895
R23158 frontAnalog_v0p0p1_4.x65.A.n1 frontAnalog_v0p0p1_4.x65.A.t4 260.322
R23159 frontAnalog_v0p0p1_4.x65.A.n3 frontAnalog_v0p0p1_4.x65.A.t7 233.929
R23160 frontAnalog_v0p0p1_4.x65.A.n1 frontAnalog_v0p0p1_4.x65.A.t5 175.169
R23161 frontAnalog_v0p0p1_4.x65.A.n2 frontAnalog_v0p0p1_4.x65.A.t6 160.416
R23162 frontAnalog_v0p0p1_4.x65.A.n4 frontAnalog_v0p0p1_4.x65.A.t2 17.4109
R23163 frontAnalog_v0p0p1_4.x65.A.n4 frontAnalog_v0p0p1_4.x65.A.t3 10.2053
R23164 frontAnalog_v0p0p1_4.x65.A.n0 frontAnalog_v0p0p1_4.x65.A 2.78715
R23165 frontAnalog_v0p0p1_4.x65.A.n0 frontAnalog_v0p0p1_4.x65.A.n1 9.09103
R23166 frontAnalog_v0p0p1_4.x65.A.n6 frontAnalog_v0p0p1_4.x65.A.t0 7.94569
R23167 frontAnalog_v0p0p1_4.x65.A.n2 frontAnalog_v0p0p1_4.x65.A.t1 7.55846
R23168 frontAnalog_v0p0p1_4.x65.A.n5 frontAnalog_v0p0p1_4.x65.A.n3 1.4614
R23169 frontAnalog_v0p0p1_4.x65.A.n3 frontAnalog_v0p0p1_4.x65.A.n2 1.19626
R23170 frontAnalog_v0p0p1_4.x65.A.n6 frontAnalog_v0p0p1_4.x65.A.n5 0.836961
R23171 frontAnalog_v0p0p1_4.x65.A frontAnalog_v0p0p1_4.x65.A.n0 0.390342
R23172 frontAnalog_v0p0p1_4.x65.A.n5 frontAnalog_v0p0p1_4.x65.A.n4 0.154668
R23173 frontAnalog_v0p0p1_4.x65.A frontAnalog_v0p0p1_4.x65.A.n6 0.08175
R23174 VV12.n0 VV12.t17 167.365
R23175 VV12.n0 VV12.t16 92.4496
R23176 VV12.n1 VV12.n0 2.07493
R23177 VV12.n17 VV12 0.560583
R23178 VV12 VV12.n17 0.420563
R23179 VV12.n15 VV12.n14 0.141409
R23180 VV12.n13 VV12.n12 0.141409
R23181 VV12.n11 VV12.n10 0.141409
R23182 VV12.n9 VV12.n8 0.141409
R23183 VV12.n7 VV12.n6 0.141409
R23184 VV12.n5 VV12.n4 0.141409
R23185 VV12.n3 VV12.n2 0.141409
R23186 VV12.n1 VV12 0.12425
R23187 VV12 VV12.n16 0.100973
R23188 VV12 VV12.n1 0.0314375
R23189 VV12.n17 VV12 0.00833333
R23190 VV12.n17 VV12 0.006375
R23191 VV12.n2 VV12.t5 0.000729415
R23192 VV12.n16 VV12.n15 0.000727273
R23193 VV12.n14 VV12.n13 0.000727273
R23194 VV12.n12 VV12.n11 0.000727273
R23195 VV12.n10 VV12.n9 0.000727273
R23196 VV12.n8 VV12.n7 0.000727273
R23197 VV12.n6 VV12.n5 0.000727273
R23198 VV12.n4 VV12.n3 0.000727273
R23199 VV12.n2 VV12.t8 0.000502142
R23200 VV12.n4 VV12.t3 0.000502142
R23201 VV12.n6 VV12.t12 0.000502142
R23202 VV12.n8 VV12.t10 0.000502142
R23203 VV12.n10 VV12.t13 0.000502142
R23204 VV12.n12 VV12.t1 0.000502142
R23205 VV12.n14 VV12.t7 0.000502142
R23206 VV12.n16 VV12.t11 0.000502142
R23207 VV12.n15 VV12.t2 0.000502142
R23208 VV12.n13 VV12.t9 0.000502142
R23209 VV12.n11 VV12.t14 0.000502142
R23210 VV12.n9 VV12.t6 0.000502142
R23211 VV12.n7 VV12.t15 0.000502142
R23212 VV12.n5 VV12.t0 0.000502142
R23213 VV12.n3 VV12.t4 0.000502142
R23214 frontAnalog_v0p0p1_9.x63.A.n2 frontAnalog_v0p0p1_9.x63.A.t5 260.322
R23215 frontAnalog_v0p0p1_9.x63.A.n4 frontAnalog_v0p0p1_9.x63.A.t6 233.888
R23216 frontAnalog_v0p0p1_9.x63.A.n2 frontAnalog_v0p0p1_9.x63.A.t7 175.169
R23217 frontAnalog_v0p0p1_9.x63.A.n3 frontAnalog_v0p0p1_9.x63.A.t4 159.725
R23218 frontAnalog_v0p0p1_9.x63.A.n1 frontAnalog_v0p0p1_9.x63.A.t2 17.4109
R23219 frontAnalog_v0p0p1_9.x63.A.n0 frontAnalog_v0p0p1_9.x63.A.n2 9.75129
R23220 frontAnalog_v0p0p1_9.x63.A.n1 frontAnalog_v0p0p1_9.x63.A.t3 9.6037
R23221 frontAnalog_v0p0p1_9.x63.A.n0 frontAnalog_v0p0p1_9.x63.A 2.33338
R23222 frontAnalog_v0p0p1_9.x63.A.n5 frontAnalog_v0p0p1_9.x63.A.t1 8.40929
R23223 frontAnalog_v0p0p1_9.x63.A.n3 frontAnalog_v0p0p1_9.x63.A.t0 8.06629
R23224 frontAnalog_v0p0p1_9.x63.A.n4 frontAnalog_v0p0p1_9.x63.A.n3 1.73501
R23225 frontAnalog_v0p0p1_9.x63.A.n1 frontAnalog_v0p0p1_9.x63.A.n4 0.99025
R23226 frontAnalog_v0p0p1_9.x63.A.n5 frontAnalog_v0p0p1_9.x63.A.n1 0.853186
R23227 frontAnalog_v0p0p1_9.x63.A frontAnalog_v0p0p1_9.x63.A.n0 0.349517
R23228 frontAnalog_v0p0p1_9.x63.A frontAnalog_v0p0p1_9.x63.A.n5 0.24425
R23229 frontAnalog_v0p0p1_9.x65.A.n1 frontAnalog_v0p0p1_9.x65.A.t6 260.322
R23230 frontAnalog_v0p0p1_9.x65.A.n3 frontAnalog_v0p0p1_9.x65.A.t5 233.929
R23231 frontAnalog_v0p0p1_9.x65.A.n1 frontAnalog_v0p0p1_9.x65.A.t4 175.169
R23232 frontAnalog_v0p0p1_9.x65.A.n2 frontAnalog_v0p0p1_9.x65.A.t7 160.416
R23233 frontAnalog_v0p0p1_9.x65.A.n4 frontAnalog_v0p0p1_9.x65.A.t0 17.4109
R23234 frontAnalog_v0p0p1_9.x65.A.n4 frontAnalog_v0p0p1_9.x65.A.t1 10.2053
R23235 frontAnalog_v0p0p1_9.x65.A.n0 frontAnalog_v0p0p1_9.x65.A 2.78715
R23236 frontAnalog_v0p0p1_9.x65.A.n0 frontAnalog_v0p0p1_9.x65.A.n1 9.09103
R23237 frontAnalog_v0p0p1_9.x65.A.n6 frontAnalog_v0p0p1_9.x65.A.t2 7.94569
R23238 frontAnalog_v0p0p1_9.x65.A.n2 frontAnalog_v0p0p1_9.x65.A.t3 7.55846
R23239 frontAnalog_v0p0p1_9.x65.A.n5 frontAnalog_v0p0p1_9.x65.A.n3 1.4614
R23240 frontAnalog_v0p0p1_9.x65.A.n3 frontAnalog_v0p0p1_9.x65.A.n2 1.19626
R23241 frontAnalog_v0p0p1_9.x65.A.n6 frontAnalog_v0p0p1_9.x65.A.n5 0.836961
R23242 frontAnalog_v0p0p1_9.x65.A frontAnalog_v0p0p1_9.x65.A.n0 0.390342
R23243 frontAnalog_v0p0p1_9.x65.A.n5 frontAnalog_v0p0p1_9.x65.A.n4 0.154668
R23244 frontAnalog_v0p0p1_9.x65.A frontAnalog_v0p0p1_9.x65.A.n6 0.08175
R23245 I1.t8 I1.t9 618.109
R23246 I1.n1 I1.t7 334.723
R23247 I1 I1.t8 253.56
R23248 I1.n1 I1.t6 206.19
R23249 I1.n5 I1.t10 117.314
R23250 I1.n5 I1.t5 110.853
R23251 I1 I1.n1 90.4462
R23252 I1.n0 I1 39.0702
R23253 I1.n7 I1.t0 17.6181
R23254 I1.n8 I1.t4 14.2865
R23255 I1.n10 I1.t1 14.283
R23256 I1.n10 I1.t2 14.283
R23257 I1.n12 I1.t3 8.77744
R23258 I1 I1.n13 8.44781
R23259 I1.n2 I1 7.13193
R23260 I1.n2 I1 5.30336
R23261 I1.n3 I1.n2 5.16688
R23262 I1.n3 I1.n0 2.29514
R23263 I1.n12 I1.n11 1.20426
R23264 I1.n0 I1 0.692911
R23265 I1.n13 I1.n12 0.32511
R23266 I1.n8 I1.n7 0.314673
R23267 I1.n9 I1.n8 0.299251
R23268 I1.n14 I1 0.2825
R23269 I1 I1.n4 0.271533
R23270 I1 I1.n14 0.212
R23271 I1.n4 I1 0.20675
R23272 I1.n6 I1.n5 0.159555
R23273 I1.n4 I1.n3 0.153447
R23274 I1.n11 I1.n10 0.106617
R23275 I1.n9 I1.n6 0.0796167
R23276 I1.n11 I1.n9 0.0480595
R23277 I1.n13 I1 0.046937
R23278 I1.n14 I1 0.0161667
R23279 I1.n14 I1 0.01225
R23280 I1.n7 I1.n6 0.000504658
R23281 frontAnalog_v0p0p1_9.RSfetsym_0.QN.n1 frontAnalog_v0p0p1_9.RSfetsym_0.QN.t6 117.511
R23282 frontAnalog_v0p0p1_9.RSfetsym_0.QN.n1 frontAnalog_v0p0p1_9.RSfetsym_0.QN.t5 110.698
R23283 frontAnalog_v0p0p1_9.RSfetsym_0.QN.n2 frontAnalog_v0p0p1_9.RSfetsym_0.QN.t2 19.1963
R23284 frontAnalog_v0p0p1_9.RSfetsym_0.QN.n3 frontAnalog_v0p0p1_9.RSfetsym_0.QN.t1 14.5206
R23285 frontAnalog_v0p0p1_9.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_9.RSfetsym_0.QN.t3 14.283
R23286 frontAnalog_v0p0p1_9.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_9.RSfetsym_0.QN.t4 14.283
R23287 frontAnalog_v0p0p1_9.RSfetsym_0.QN frontAnalog_v0p0p1_9.RSfetsym_0.QN.t0 9.14075
R23288 frontAnalog_v0p0p1_9.RSfetsym_0.QN.n2 frontAnalog_v0p0p1_9.RSfetsym_0.QN.n1 0.826818
R23289 frontAnalog_v0p0p1_9.RSfetsym_0.QN frontAnalog_v0p0p1_9.RSfetsym_0.QN.n0 0.74645
R23290 frontAnalog_v0p0p1_9.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_9.RSfetsym_0.QN.n3 0.249509
R23291 frontAnalog_v0p0p1_9.RSfetsym_0.QN.n3 frontAnalog_v0p0p1_9.RSfetsym_0.QN.n2 0.0968646
R23292 I6.n17 I6.t6 260.435
R23293 I6.n2 I6.t10 229.433
R23294 I6.n12 I6.t11 196.549
R23295 I6.n2 I6.t7 158.885
R23296 I6.n17 I6.t8 156.403
R23297 I6.n12 I6.t12 148.35
R23298 I6.n25 I6.t9 117.314
R23299 I6.n25 I6.t5 110.853
R23300 I6.n13 I6.n12 76.0005
R23301 I6.n27 I6.t1 17.6181
R23302 I6.n28 I6.t0 14.2865
R23303 I6.n30 I6.t2 14.283
R23304 I6.n30 I6.t3 14.283
R23305 I6.n5 I6.n4 9.3005
R23306 I6.n9 I6.n8 9.3005
R23307 I6.n5 I6.n3 9.3005
R23308 I6 I6.n16 9.3005
R23309 I6.n32 I6.t4 8.77744
R23310 I6.n18 I6.n17 7.60183
R23311 I6.n3 I6.n2 7.39171
R23312 I6.n22 I6.n14 6.24391
R23313 I6.n13 I6 5.78114
R23314 I6.n18 I6 4.8645
R23315 I6.n19 I6.n15 4.54557
R23316 I6.n10 I6.n9 4.51698
R23317 I6.n16 I6.n15 4.51121
R23318 I6.n8 I6.n7 4.5005
R23319 I6.n22 I6.n21 3.53643
R23320 I6.n14 I6.n13 3.51018
R23321 I6.n8 I6.n4 3.46717
R23322 I6 I6.n33 1.82181
R23323 I6.n32 I6.n31 1.20426
R23324 I6.n6 I6.n0 1.13339
R23325 I6.n11 I6.n10 1.11384
R23326 I6.n8 I6.n3 1.06717
R23327 I6.n4 I6 1.06717
R23328 I6.n23 I6.n11 0.874607
R23329 I6.n34 I6 0.6585
R23330 I6 I6.n24 0.647533
R23331 I6.n24 I6.n23 0.520635
R23332 I6 I6.n34 0.494
R23333 I6.n11 I6 0.372375
R23334 I6.n33 I6.n32 0.32511
R23335 I6.n28 I6.n27 0.314673
R23336 I6.n29 I6.n28 0.299251
R23337 I6.n23 I6.n22 0.214786
R23338 I6.n14 I6 0.206952
R23339 I6.n24 I6 0.20675
R23340 I6.n26 I6.n25 0.159555
R23341 I6.n31 I6.n30 0.106617
R23342 I6.n29 I6.n26 0.0796167
R23343 I6.n31 I6.n29 0.0480595
R23344 I6.n33 I6 0.046937
R23345 I6.n20 I6.n16 0.0344286
R23346 I6.n10 I6.n0 0.028
R23347 I6.n34 I6 0.0161667
R23348 I6.n9 I6.n1 0.0142363
R23349 I6.n34 I6 0.01225
R23350 I6.n7 I6.n1 0.00599451
R23351 I6.n6 I6.n5 0.00484776
R23352 I6.n7 I6.n6 0.00226981
R23353 I6.n21 I6.n15 0.00182856
R23354 I6.n21 I6.n20 0.00149885
R23355 I6.n19 I6.n18 0.00133362
R23356 I6.n20 I6.n19 0.00100077
R23357 I6.n1 I6.n0 0.000617139
R23358 I6.n27 I6.n26 0.000504658
R23359 frontAnalog_v0p0p1_13.RSfetsym_0.QN.n1 frontAnalog_v0p0p1_13.RSfetsym_0.QN.t6 117.511
R23360 frontAnalog_v0p0p1_13.RSfetsym_0.QN.n1 frontAnalog_v0p0p1_13.RSfetsym_0.QN.t5 110.698
R23361 frontAnalog_v0p0p1_13.RSfetsym_0.QN.n2 frontAnalog_v0p0p1_13.RSfetsym_0.QN.t1 19.1963
R23362 frontAnalog_v0p0p1_13.RSfetsym_0.QN.n3 frontAnalog_v0p0p1_13.RSfetsym_0.QN.t0 14.5206
R23363 frontAnalog_v0p0p1_13.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_13.RSfetsym_0.QN.t3 14.283
R23364 frontAnalog_v0p0p1_13.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_13.RSfetsym_0.QN.t2 14.283
R23365 frontAnalog_v0p0p1_13.RSfetsym_0.QN frontAnalog_v0p0p1_13.RSfetsym_0.QN.t4 9.14075
R23366 frontAnalog_v0p0p1_13.RSfetsym_0.QN.n2 frontAnalog_v0p0p1_13.RSfetsym_0.QN.n1 0.826818
R23367 frontAnalog_v0p0p1_13.RSfetsym_0.QN frontAnalog_v0p0p1_13.RSfetsym_0.QN.n0 0.74645
R23368 frontAnalog_v0p0p1_13.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_13.RSfetsym_0.QN.n3 0.249509
R23369 frontAnalog_v0p0p1_13.RSfetsym_0.QN.n3 frontAnalog_v0p0p1_13.RSfetsym_0.QN.n2 0.0968646
R23370 frontAnalog_v0p0p1_7.x65.A.n1 frontAnalog_v0p0p1_7.x65.A.t7 260.322
R23371 frontAnalog_v0p0p1_7.x65.A.n3 frontAnalog_v0p0p1_7.x65.A.t6 233.929
R23372 frontAnalog_v0p0p1_7.x65.A.n1 frontAnalog_v0p0p1_7.x65.A.t5 175.169
R23373 frontAnalog_v0p0p1_7.x65.A.n2 frontAnalog_v0p0p1_7.x65.A.t4 160.416
R23374 frontAnalog_v0p0p1_7.x65.A.n4 frontAnalog_v0p0p1_7.x65.A.t1 17.4109
R23375 frontAnalog_v0p0p1_7.x65.A.n4 frontAnalog_v0p0p1_7.x65.A.t0 10.2053
R23376 frontAnalog_v0p0p1_7.x65.A.n0 frontAnalog_v0p0p1_7.x65.A 2.78715
R23377 frontAnalog_v0p0p1_7.x65.A.n0 frontAnalog_v0p0p1_7.x65.A.n1 9.09103
R23378 frontAnalog_v0p0p1_7.x65.A.n6 frontAnalog_v0p0p1_7.x65.A.t3 7.94569
R23379 frontAnalog_v0p0p1_7.x65.A.n2 frontAnalog_v0p0p1_7.x65.A.t2 7.55846
R23380 frontAnalog_v0p0p1_7.x65.A.n5 frontAnalog_v0p0p1_7.x65.A.n3 1.4614
R23381 frontAnalog_v0p0p1_7.x65.A.n3 frontAnalog_v0p0p1_7.x65.A.n2 1.19626
R23382 frontAnalog_v0p0p1_7.x65.A.n6 frontAnalog_v0p0p1_7.x65.A.n5 0.836961
R23383 frontAnalog_v0p0p1_7.x65.A frontAnalog_v0p0p1_7.x65.A.n0 0.390342
R23384 frontAnalog_v0p0p1_7.x65.A.n5 frontAnalog_v0p0p1_7.x65.A.n4 0.154668
R23385 frontAnalog_v0p0p1_7.x65.A frontAnalog_v0p0p1_7.x65.A.n6 0.08175
R23386 frontAnalog_v0p0p1_7.x63.A.n2 frontAnalog_v0p0p1_7.x63.A.t6 260.322
R23387 frontAnalog_v0p0p1_7.x63.A.n4 frontAnalog_v0p0p1_7.x63.A.t7 233.888
R23388 frontAnalog_v0p0p1_7.x63.A.n2 frontAnalog_v0p0p1_7.x63.A.t4 175.169
R23389 frontAnalog_v0p0p1_7.x63.A.n3 frontAnalog_v0p0p1_7.x63.A.t5 159.725
R23390 frontAnalog_v0p0p1_7.x63.A.n1 frontAnalog_v0p0p1_7.x63.A.t2 17.4109
R23391 frontAnalog_v0p0p1_7.x63.A.n0 frontAnalog_v0p0p1_7.x63.A.n2 9.75129
R23392 frontAnalog_v0p0p1_7.x63.A.n1 frontAnalog_v0p0p1_7.x63.A.t3 9.6037
R23393 frontAnalog_v0p0p1_7.x63.A.n0 frontAnalog_v0p0p1_7.x63.A 2.33338
R23394 frontAnalog_v0p0p1_7.x63.A.n5 frontAnalog_v0p0p1_7.x63.A.t1 8.40929
R23395 frontAnalog_v0p0p1_7.x63.A.n3 frontAnalog_v0p0p1_7.x63.A.t0 8.06629
R23396 frontAnalog_v0p0p1_7.x63.A.n4 frontAnalog_v0p0p1_7.x63.A.n3 1.73501
R23397 frontAnalog_v0p0p1_7.x63.A.n1 frontAnalog_v0p0p1_7.x63.A.n4 0.99025
R23398 frontAnalog_v0p0p1_7.x63.A.n5 frontAnalog_v0p0p1_7.x63.A.n1 0.853186
R23399 frontAnalog_v0p0p1_7.x63.A frontAnalog_v0p0p1_7.x63.A.n0 0.349517
R23400 frontAnalog_v0p0p1_7.x63.A frontAnalog_v0p0p1_7.x63.A.n5 0.24425
R23401 I9.t7 I9.t9 618.109
R23402 I9.n1 I9.t8 334.723
R23403 I9 I9.t7 253.56
R23404 I9.n1 I9.t5 206.19
R23405 I9.n5 I9.t10 117.314
R23406 I9.n5 I9.t6 110.852
R23407 I9 I9.n1 90.4462
R23408 I9.n0 I9 39.0702
R23409 I9.n7 I9.t2 17.6181
R23410 I9.n8 I9.t3 14.2865
R23411 I9.n10 I9.t0 14.283
R23412 I9.n10 I9.t1 14.283
R23413 I9.n12 I9.t4 8.77592
R23414 I9.n2 I9 7.13193
R23415 I9.n2 I9 5.30336
R23416 I9.n3 I9.n2 5.27402
R23417 I9.n3 I9.n0 2.188
R23418 I9.n14 I9 1.2225
R23419 I9 I9.n4 1.20605
R23420 I9.n12 I9.n11 1.20426
R23421 I9 I9.n13 1.08107
R23422 I9.n0 I9 0.692911
R23423 I9 I9.n14 0.6115
R23424 I9.n13 I9.n12 0.338241
R23425 I9.n8 I9.n7 0.314673
R23426 I9.n9 I9.n8 0.300251
R23427 I9.n4 I9 0.2005
R23428 I9.n4 I9.n3 0.166764
R23429 I9.n6 I9.n5 0.159555
R23430 I9.n11 I9.n10 0.106617
R23431 I9.n9 I9.n6 0.0796167
R23432 I9.n11 I9.n9 0.0480595
R23433 I9.n14 I9 0.024
R23434 I9.n14 I9 0.01225
R23435 I9.n13 I9 0.00440792
R23436 I9.n7 I9.n6 0.000504658
R23437 VV7.n0 VV7.t16 167.365
R23438 VV7.n0 VV7.t17 92.4488
R23439 VV7.n1 VV7.n0 2.07493
R23440 VV7.n10 VV7 0.462667
R23441 VV7 VV7.n10 0.347125
R23442 VV7.n9 VV7.n8 0.141636
R23443 VV7.n8 VV7.n7 0.141636
R23444 VV7.n7 VV7.n6 0.141636
R23445 VV7.n6 VV7.n5 0.141636
R23446 VV7.n5 VV7.n4 0.141636
R23447 VV7.n4 VV7.n3 0.141636
R23448 VV7.n3 VV7.n2 0.141636
R23449 VV7.n1 VV7 0.12425
R23450 VV7 VV7.n9 0.101201
R23451 VV7 VV7.n1 0.028
R23452 VV7.n10 VV7 0.00833333
R23453 VV7.n10 VV7 0.006375
R23454 VV7.n3 VV7.t11 0.000502142
R23455 VV7.n4 VV7.t9 0.000502142
R23456 VV7.n5 VV7.t14 0.000502142
R23457 VV7.n6 VV7.t5 0.000502142
R23458 VV7.n7 VV7.t13 0.000502142
R23459 VV7.n8 VV7.t3 0.000502142
R23460 VV7.n9 VV7.t15 0.000502142
R23461 VV7.n2 VV7.t8 0.000502142
R23462 VV7.n3 VV7.t6 0.000502142
R23463 VV7.n4 VV7.t10 0.000502142
R23464 VV7.n5 VV7.t1 0.000502142
R23465 VV7.n6 VV7.t2 0.000502142
R23466 VV7.n7 VV7.t12 0.000502142
R23467 VV7.n8 VV7.t0 0.000502142
R23468 VV7.n9 VV7.t7 0.000502142
R23469 VV7.n2 VV7.t4 0.000502142
R23470 frontAnalog_v0p0p1_13.x63.A.n2 frontAnalog_v0p0p1_13.x63.A.t4 260.322
R23471 frontAnalog_v0p0p1_13.x63.A.n4 frontAnalog_v0p0p1_13.x63.A.t5 233.888
R23472 frontAnalog_v0p0p1_13.x63.A.n2 frontAnalog_v0p0p1_13.x63.A.t6 175.169
R23473 frontAnalog_v0p0p1_13.x63.A.n3 frontAnalog_v0p0p1_13.x63.A.t7 159.725
R23474 frontAnalog_v0p0p1_13.x63.A.n1 frontAnalog_v0p0p1_13.x63.A.t3 17.4109
R23475 frontAnalog_v0p0p1_13.x63.A.n0 frontAnalog_v0p0p1_13.x63.A.n2 9.75129
R23476 frontAnalog_v0p0p1_13.x63.A.n1 frontAnalog_v0p0p1_13.x63.A.t2 9.6037
R23477 frontAnalog_v0p0p1_13.x63.A.n0 frontAnalog_v0p0p1_13.x63.A 2.33338
R23478 frontAnalog_v0p0p1_13.x63.A.n5 frontAnalog_v0p0p1_13.x63.A.t0 8.40929
R23479 frontAnalog_v0p0p1_13.x63.A.n3 frontAnalog_v0p0p1_13.x63.A.t1 8.06629
R23480 frontAnalog_v0p0p1_13.x63.A.n4 frontAnalog_v0p0p1_13.x63.A.n3 1.73501
R23481 frontAnalog_v0p0p1_13.x63.A.n1 frontAnalog_v0p0p1_13.x63.A.n4 0.99025
R23482 frontAnalog_v0p0p1_13.x63.A.n5 frontAnalog_v0p0p1_13.x63.A.n1 0.853186
R23483 frontAnalog_v0p0p1_13.x63.A frontAnalog_v0p0p1_13.x63.A.n0 0.349517
R23484 frontAnalog_v0p0p1_13.x63.A frontAnalog_v0p0p1_13.x63.A.n5 0.24425
R23485 frontAnalog_v0p0p1_10.x63.A.n2 frontAnalog_v0p0p1_10.x63.A.t5 260.322
R23486 frontAnalog_v0p0p1_10.x63.A.n4 frontAnalog_v0p0p1_10.x63.A.t6 233.888
R23487 frontAnalog_v0p0p1_10.x63.A.n2 frontAnalog_v0p0p1_10.x63.A.t7 175.169
R23488 frontAnalog_v0p0p1_10.x63.A.n3 frontAnalog_v0p0p1_10.x63.A.t4 159.725
R23489 frontAnalog_v0p0p1_10.x63.A.n1 frontAnalog_v0p0p1_10.x63.A.t0 17.4109
R23490 frontAnalog_v0p0p1_10.x63.A.n0 frontAnalog_v0p0p1_10.x63.A.n2 9.75129
R23491 frontAnalog_v0p0p1_10.x63.A.n1 frontAnalog_v0p0p1_10.x63.A.t1 9.6027
R23492 frontAnalog_v0p0p1_10.x63.A.n0 frontAnalog_v0p0p1_10.x63.A 2.33338
R23493 frontAnalog_v0p0p1_10.x63.A.n5 frontAnalog_v0p0p1_10.x63.A.t2 8.40929
R23494 frontAnalog_v0p0p1_10.x63.A.n3 frontAnalog_v0p0p1_10.x63.A.t3 8.06629
R23495 frontAnalog_v0p0p1_10.x63.A.n4 frontAnalog_v0p0p1_10.x63.A.n3 1.73501
R23496 frontAnalog_v0p0p1_10.x63.A.n1 frontAnalog_v0p0p1_10.x63.A.n4 0.99025
R23497 frontAnalog_v0p0p1_10.x63.A.n5 frontAnalog_v0p0p1_10.x63.A.n1 0.853186
R23498 frontAnalog_v0p0p1_10.x63.A frontAnalog_v0p0p1_10.x63.A.n0 0.349517
R23499 frontAnalog_v0p0p1_10.x63.A frontAnalog_v0p0p1_10.x63.A.n5 0.24425
R23500 frontAnalog_v0p0p1_5.x63.A.n2 frontAnalog_v0p0p1_5.x63.A.t4 260.322
R23501 frontAnalog_v0p0p1_5.x63.A.n4 frontAnalog_v0p0p1_5.x63.A.t5 233.888
R23502 frontAnalog_v0p0p1_5.x63.A.n2 frontAnalog_v0p0p1_5.x63.A.t6 175.169
R23503 frontAnalog_v0p0p1_5.x63.A.n3 frontAnalog_v0p0p1_5.x63.A.t7 159.725
R23504 frontAnalog_v0p0p1_5.x63.A.n1 frontAnalog_v0p0p1_5.x63.A.t1 17.4109
R23505 frontAnalog_v0p0p1_5.x63.A.n0 frontAnalog_v0p0p1_5.x63.A.n2 9.75129
R23506 frontAnalog_v0p0p1_5.x63.A.n1 frontAnalog_v0p0p1_5.x63.A.t0 9.6027
R23507 frontAnalog_v0p0p1_5.x63.A.n0 frontAnalog_v0p0p1_5.x63.A 2.33338
R23508 frontAnalog_v0p0p1_5.x63.A.n5 frontAnalog_v0p0p1_5.x63.A.t3 8.40929
R23509 frontAnalog_v0p0p1_5.x63.A.n3 frontAnalog_v0p0p1_5.x63.A.t2 8.06629
R23510 frontAnalog_v0p0p1_5.x63.A.n4 frontAnalog_v0p0p1_5.x63.A.n3 1.73501
R23511 frontAnalog_v0p0p1_5.x63.A.n1 frontAnalog_v0p0p1_5.x63.A.n4 0.99025
R23512 frontAnalog_v0p0p1_5.x63.A.n5 frontAnalog_v0p0p1_5.x63.A.n1 0.853186
R23513 frontAnalog_v0p0p1_5.x63.A frontAnalog_v0p0p1_5.x63.A.n0 0.349517
R23514 frontAnalog_v0p0p1_5.x63.A frontAnalog_v0p0p1_5.x63.A.n5 0.24425
R23515 frontAnalog_v0p0p1_3.x63.A.n2 frontAnalog_v0p0p1_3.x63.A.t5 260.322
R23516 frontAnalog_v0p0p1_3.x63.A.n4 frontAnalog_v0p0p1_3.x63.A.t6 233.888
R23517 frontAnalog_v0p0p1_3.x63.A.n2 frontAnalog_v0p0p1_3.x63.A.t7 175.169
R23518 frontAnalog_v0p0p1_3.x63.A.n3 frontAnalog_v0p0p1_3.x63.A.t4 159.725
R23519 frontAnalog_v0p0p1_3.x63.A.n1 frontAnalog_v0p0p1_3.x63.A.t3 17.4109
R23520 frontAnalog_v0p0p1_3.x63.A.n0 frontAnalog_v0p0p1_3.x63.A.n2 9.75129
R23521 frontAnalog_v0p0p1_3.x63.A.n1 frontAnalog_v0p0p1_3.x63.A.t2 9.6037
R23522 frontAnalog_v0p0p1_3.x63.A.n0 frontAnalog_v0p0p1_3.x63.A 2.33338
R23523 frontAnalog_v0p0p1_3.x63.A.n5 frontAnalog_v0p0p1_3.x63.A.t0 8.40929
R23524 frontAnalog_v0p0p1_3.x63.A.n3 frontAnalog_v0p0p1_3.x63.A.t1 8.06629
R23525 frontAnalog_v0p0p1_3.x63.A.n4 frontAnalog_v0p0p1_3.x63.A.n3 1.73501
R23526 frontAnalog_v0p0p1_3.x63.A.n1 frontAnalog_v0p0p1_3.x63.A.n4 0.99025
R23527 frontAnalog_v0p0p1_3.x63.A.n5 frontAnalog_v0p0p1_3.x63.A.n1 0.853186
R23528 frontAnalog_v0p0p1_3.x63.A frontAnalog_v0p0p1_3.x63.A.n0 0.349517
R23529 frontAnalog_v0p0p1_3.x63.A frontAnalog_v0p0p1_3.x63.A.n5 0.24425
R23530 frontAnalog_v0p0p1_3.x65.A.n1 frontAnalog_v0p0p1_3.x65.A.t4 260.322
R23531 frontAnalog_v0p0p1_3.x65.A.n4 frontAnalog_v0p0p1_3.x65.A.t7 233.929
R23532 frontAnalog_v0p0p1_3.x65.A.n1 frontAnalog_v0p0p1_3.x65.A.t6 175.169
R23533 frontAnalog_v0p0p1_3.x65.A.n3 frontAnalog_v0p0p1_3.x65.A.t5 160.416
R23534 frontAnalog_v0p0p1_3.x65.A.n2 frontAnalog_v0p0p1_3.x65.A.t2 17.4109
R23535 frontAnalog_v0p0p1_3.x65.A.n2 frontAnalog_v0p0p1_3.x65.A.t3 10.2053
R23536 frontAnalog_v0p0p1_3.x65.A.n0 frontAnalog_v0p0p1_3.x65.A 2.78715
R23537 frontAnalog_v0p0p1_3.x65.A.n0 frontAnalog_v0p0p1_3.x65.A.n1 9.09103
R23538 frontAnalog_v0p0p1_3.x65.A.n6 frontAnalog_v0p0p1_3.x65.A.t1 7.94569
R23539 frontAnalog_v0p0p1_3.x65.A.n3 frontAnalog_v0p0p1_3.x65.A.t0 7.55846
R23540 frontAnalog_v0p0p1_3.x65.A.n5 frontAnalog_v0p0p1_3.x65.A.n4 1.4614
R23541 frontAnalog_v0p0p1_3.x65.A.n4 frontAnalog_v0p0p1_3.x65.A.n3 1.19626
R23542 frontAnalog_v0p0p1_3.x65.A.n6 frontAnalog_v0p0p1_3.x65.A.n5 0.836961
R23543 frontAnalog_v0p0p1_3.x65.A frontAnalog_v0p0p1_3.x65.A.n0 0.390342
R23544 frontAnalog_v0p0p1_3.x65.A.n5 frontAnalog_v0p0p1_3.x65.A.n2 0.154668
R23545 frontAnalog_v0p0p1_3.x65.A frontAnalog_v0p0p1_3.x65.A.n6 0.08175
R23546 S0.n0 S0.t4 260.322
R23547 S0.n7 S0.t7 233.929
R23548 S0.n0 S0.t6 175.169
R23549 S0.n6 S0.t5 160.416
R23550 S0.n8 S0.t0 17.4109
R23551 S0.n8 S0.t1 10.2053
R23552 S0.n2 S0 9.3005
R23553 S0.n1 S0.n0 9.09103
R23554 S0 S0.t2 7.94569
R23555 S0.n6 S0.t3 7.55846
R23556 S0 S0.n1 3.97938
R23557 S0.n3 S0 2.5505
R23558 S0.n9 S0.n7 1.4614
R23559 S0.n7 S0.n6 1.19626
R23560 S0.n10 S0.n9 0.808836
R23561 S0.n11 S0.n2 0.223714
R23562 S0.n9 S0.n8 0.154668
R23563 S0.n4 S0 0.140229
R23564 S0.n5 S0 0.119808
R23565 S0.n5 S0 0.0988607
R23566 S0.n2 S0.n1 0.0421278
R23567 S0.n5 S0.n4 0.0341093
R23568 S0 S0.n5 0.033122
R23569 S0 S0.n11 0.0306829
R23570 S0.n10 S0 0.0233659
R23571 S0.n11 S0.n10 0.0114756
R23572 S0.n3 S0 0.00354878
R23573 S0.n4 S0.n3 0.00306933
R23574 frontAnalog_v0p0p1_4.x63.A.n2 frontAnalog_v0p0p1_4.x63.A.t6 260.322
R23575 frontAnalog_v0p0p1_4.x63.A.n4 frontAnalog_v0p0p1_4.x63.A.t4 233.888
R23576 frontAnalog_v0p0p1_4.x63.A.n2 frontAnalog_v0p0p1_4.x63.A.t5 175.169
R23577 frontAnalog_v0p0p1_4.x63.A.n3 frontAnalog_v0p0p1_4.x63.A.t7 159.725
R23578 frontAnalog_v0p0p1_4.x63.A.n1 frontAnalog_v0p0p1_4.x63.A.t0 17.4109
R23579 frontAnalog_v0p0p1_4.x63.A.n0 frontAnalog_v0p0p1_4.x63.A.n2 9.75129
R23580 frontAnalog_v0p0p1_4.x63.A.n1 frontAnalog_v0p0p1_4.x63.A.t1 9.6027
R23581 frontAnalog_v0p0p1_4.x63.A.n0 frontAnalog_v0p0p1_4.x63.A 2.33338
R23582 frontAnalog_v0p0p1_4.x63.A.n5 frontAnalog_v0p0p1_4.x63.A.t2 8.40929
R23583 frontAnalog_v0p0p1_4.x63.A.n3 frontAnalog_v0p0p1_4.x63.A.t3 8.06629
R23584 frontAnalog_v0p0p1_4.x63.A.n4 frontAnalog_v0p0p1_4.x63.A.n3 1.73501
R23585 frontAnalog_v0p0p1_4.x63.A.n1 frontAnalog_v0p0p1_4.x63.A.n4 0.99025
R23586 frontAnalog_v0p0p1_4.x63.A.n5 frontAnalog_v0p0p1_4.x63.A.n1 0.853186
R23587 frontAnalog_v0p0p1_4.x63.A frontAnalog_v0p0p1_4.x63.A.n0 0.349517
R23588 frontAnalog_v0p0p1_4.x63.A frontAnalog_v0p0p1_4.x63.A.n5 0.24425
R23589 frontAnalog_v0p0p1_1.x65.A.n1 frontAnalog_v0p0p1_1.x65.A.t4 260.322
R23590 frontAnalog_v0p0p1_1.x65.A.n3 frontAnalog_v0p0p1_1.x65.A.t7 233.929
R23591 frontAnalog_v0p0p1_1.x65.A.n1 frontAnalog_v0p0p1_1.x65.A.t6 175.169
R23592 frontAnalog_v0p0p1_1.x65.A.n2 frontAnalog_v0p0p1_1.x65.A.t5 160.416
R23593 frontAnalog_v0p0p1_1.x65.A.n4 frontAnalog_v0p0p1_1.x65.A.t2 17.4109
R23594 frontAnalog_v0p0p1_1.x65.A.n4 frontAnalog_v0p0p1_1.x65.A.t3 10.2053
R23595 frontAnalog_v0p0p1_1.x65.A.n0 frontAnalog_v0p0p1_1.x65.A 2.78715
R23596 frontAnalog_v0p0p1_1.x65.A.n0 frontAnalog_v0p0p1_1.x65.A.n1 9.09103
R23597 frontAnalog_v0p0p1_1.x65.A.n6 frontAnalog_v0p0p1_1.x65.A.t0 7.94569
R23598 frontAnalog_v0p0p1_1.x65.A.n2 frontAnalog_v0p0p1_1.x65.A.t1 7.55846
R23599 frontAnalog_v0p0p1_1.x65.A.n5 frontAnalog_v0p0p1_1.x65.A.n3 1.4614
R23600 frontAnalog_v0p0p1_1.x65.A.n3 frontAnalog_v0p0p1_1.x65.A.n2 1.19626
R23601 frontAnalog_v0p0p1_1.x65.A.n6 frontAnalog_v0p0p1_1.x65.A.n5 0.836961
R23602 frontAnalog_v0p0p1_1.x65.A frontAnalog_v0p0p1_1.x65.A.n0 0.390342
R23603 frontAnalog_v0p0p1_1.x65.A.n5 frontAnalog_v0p0p1_1.x65.A.n4 0.154668
R23604 frontAnalog_v0p0p1_1.x65.A frontAnalog_v0p0p1_1.x65.A.n6 0.08175
R23605 frontAnalog_v0p0p1_10.RSfetsym_0.QN.n1 frontAnalog_v0p0p1_10.RSfetsym_0.QN.t6 117.511
R23606 frontAnalog_v0p0p1_10.RSfetsym_0.QN.n1 frontAnalog_v0p0p1_10.RSfetsym_0.QN.t5 110.698
R23607 frontAnalog_v0p0p1_10.RSfetsym_0.QN.n2 frontAnalog_v0p0p1_10.RSfetsym_0.QN.t1 19.1963
R23608 frontAnalog_v0p0p1_10.RSfetsym_0.QN.n3 frontAnalog_v0p0p1_10.RSfetsym_0.QN.t4 14.5206
R23609 frontAnalog_v0p0p1_10.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_10.RSfetsym_0.QN.t2 14.283
R23610 frontAnalog_v0p0p1_10.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_10.RSfetsym_0.QN.t3 14.283
R23611 frontAnalog_v0p0p1_10.RSfetsym_0.QN frontAnalog_v0p0p1_10.RSfetsym_0.QN.t0 9.14075
R23612 frontAnalog_v0p0p1_10.RSfetsym_0.QN.n2 frontAnalog_v0p0p1_10.RSfetsym_0.QN.n1 0.826818
R23613 frontAnalog_v0p0p1_10.RSfetsym_0.QN frontAnalog_v0p0p1_10.RSfetsym_0.QN.n0 0.74645
R23614 frontAnalog_v0p0p1_10.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_10.RSfetsym_0.QN.n3 0.249509
R23615 frontAnalog_v0p0p1_10.RSfetsym_0.QN.n3 frontAnalog_v0p0p1_10.RSfetsym_0.QN.n2 0.0968646
R23616 I4.n2 I4.t5 260.435
R23617 I4.n7 I4.t11 230.576
R23618 I4.n10 I4.t7 196.549
R23619 I4.n7 I4.t8 158.275
R23620 I4.n2 I4.t10 156.403
R23621 I4.n10 I4.t9 148.35
R23622 I4.n15 I4.t6 117.314
R23623 I4.n15 I4.t12 110.853
R23624 I4.n17 I4.t1 17.6181
R23625 I4.n18 I4.t4 14.2865
R23626 I4.n20 I4.t3 14.283
R23627 I4.n20 I4.t2 14.283
R23628 I4.n11 I4.n10 9.49829
R23629 I4 I4.n1 9.3005
R23630 I4.n22 I4.t0 8.77744
R23631 I4.n8 I4.n7 8.76429
R23632 I4.n12 I4.n11 7.9582
R23633 I4.n9 I4.n8 7.74345
R23634 I4.n3 I4.n2 7.60183
R23635 I4.n8 I4 6.66717
R23636 I4.n11 I4 6.44139
R23637 I4.n3 I4 4.8645
R23638 I4.n4 I4.n0 4.54557
R23639 I4.n1 I4.n0 4.51121
R23640 I4 I4.n23 4.47065
R23641 I4.n13 I4.n6 2.33148
R23642 I4.n22 I4.n21 1.20426
R23643 I4.n12 I4.n9 1.0005
R23644 I4.n24 I4 0.509667
R23645 I4 I4.n14 0.4987
R23646 I4.n13 I4.n12 0.446956
R23647 I4 I4.n24 0.382375
R23648 I4.n9 I4 0.380411
R23649 I4.n14 I4.n13 0.368862
R23650 I4.n23 I4.n22 0.32511
R23651 I4.n18 I4.n17 0.314673
R23652 I4.n19 I4.n18 0.299251
R23653 I4.n14 I4 0.20675
R23654 I4.n16 I4.n15 0.159555
R23655 I4.n21 I4.n20 0.106617
R23656 I4.n19 I4.n16 0.0796167
R23657 I4.n21 I4.n19 0.0480595
R23658 I4.n23 I4 0.046937
R23659 I4.n5 I4.n1 0.0344286
R23660 I4.n24 I4 0.0161667
R23661 I4.n24 I4 0.01225
R23662 I4.n6 I4.n0 0.00182856
R23663 I4.n6 I4.n5 0.00149885
R23664 I4.n4 I4.n3 0.00133362
R23665 I4.n5 I4.n4 0.00100077
R23666 I4.n17 I4.n16 0.000504658
R23667 frontAnalog_v0p0p1_3.RSfetsym_0.QN.n1 frontAnalog_v0p0p1_3.RSfetsym_0.QN.t6 117.511
R23668 frontAnalog_v0p0p1_3.RSfetsym_0.QN.n1 frontAnalog_v0p0p1_3.RSfetsym_0.QN.t5 110.698
R23669 frontAnalog_v0p0p1_3.RSfetsym_0.QN.n2 frontAnalog_v0p0p1_3.RSfetsym_0.QN.t3 19.1963
R23670 frontAnalog_v0p0p1_3.RSfetsym_0.QN.n3 frontAnalog_v0p0p1_3.RSfetsym_0.QN.t0 14.5206
R23671 frontAnalog_v0p0p1_3.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_3.RSfetsym_0.QN.t1 14.283
R23672 frontAnalog_v0p0p1_3.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_3.RSfetsym_0.QN.t2 14.283
R23673 frontAnalog_v0p0p1_3.RSfetsym_0.QN frontAnalog_v0p0p1_3.RSfetsym_0.QN.t4 9.14075
R23674 frontAnalog_v0p0p1_3.RSfetsym_0.QN.n2 frontAnalog_v0p0p1_3.RSfetsym_0.QN.n1 0.826818
R23675 frontAnalog_v0p0p1_3.RSfetsym_0.QN frontAnalog_v0p0p1_3.RSfetsym_0.QN.n0 0.74645
R23676 frontAnalog_v0p0p1_3.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_3.RSfetsym_0.QN.n3 0.249509
R23677 frontAnalog_v0p0p1_3.RSfetsym_0.QN.n3 frontAnalog_v0p0p1_3.RSfetsym_0.QN.n2 0.0968646
R23678 frontAnalog_v0p0p1_6.x63.A.n2 frontAnalog_v0p0p1_6.x63.A.t4 260.322
R23679 frontAnalog_v0p0p1_6.x63.A.n4 frontAnalog_v0p0p1_6.x63.A.t7 233.888
R23680 frontAnalog_v0p0p1_6.x63.A.n2 frontAnalog_v0p0p1_6.x63.A.t6 175.169
R23681 frontAnalog_v0p0p1_6.x63.A.n3 frontAnalog_v0p0p1_6.x63.A.t5 159.725
R23682 frontAnalog_v0p0p1_6.x63.A.n1 frontAnalog_v0p0p1_6.x63.A.t1 17.4109
R23683 frontAnalog_v0p0p1_6.x63.A.n0 frontAnalog_v0p0p1_6.x63.A.n2 9.75129
R23684 frontAnalog_v0p0p1_6.x63.A.n1 frontAnalog_v0p0p1_6.x63.A.t0 9.6027
R23685 frontAnalog_v0p0p1_6.x63.A.n0 frontAnalog_v0p0p1_6.x63.A 2.33338
R23686 frontAnalog_v0p0p1_6.x63.A.n5 frontAnalog_v0p0p1_6.x63.A.t2 8.40929
R23687 frontAnalog_v0p0p1_6.x63.A.n3 frontAnalog_v0p0p1_6.x63.A.t3 8.06629
R23688 frontAnalog_v0p0p1_6.x63.A.n4 frontAnalog_v0p0p1_6.x63.A.n3 1.73501
R23689 frontAnalog_v0p0p1_6.x63.A.n1 frontAnalog_v0p0p1_6.x63.A.n4 0.99025
R23690 frontAnalog_v0p0p1_6.x63.A.n5 frontAnalog_v0p0p1_6.x63.A.n1 0.853186
R23691 frontAnalog_v0p0p1_6.x63.A frontAnalog_v0p0p1_6.x63.A.n0 0.349517
R23692 frontAnalog_v0p0p1_6.x63.A frontAnalog_v0p0p1_6.x63.A.n5 0.24425
R23693 frontAnalog_v0p0p1_12.RSfetsym_0.QN.n1 frontAnalog_v0p0p1_12.RSfetsym_0.QN.t6 117.511
R23694 frontAnalog_v0p0p1_12.RSfetsym_0.QN.n1 frontAnalog_v0p0p1_12.RSfetsym_0.QN.t5 110.698
R23695 frontAnalog_v0p0p1_12.RSfetsym_0.QN.n2 frontAnalog_v0p0p1_12.RSfetsym_0.QN.t0 19.1963
R23696 frontAnalog_v0p0p1_12.RSfetsym_0.QN.n3 frontAnalog_v0p0p1_12.RSfetsym_0.QN.t4 14.5206
R23697 frontAnalog_v0p0p1_12.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_12.RSfetsym_0.QN.t2 14.283
R23698 frontAnalog_v0p0p1_12.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_12.RSfetsym_0.QN.t1 14.283
R23699 frontAnalog_v0p0p1_12.RSfetsym_0.QN frontAnalog_v0p0p1_12.RSfetsym_0.QN.t3 9.14075
R23700 frontAnalog_v0p0p1_12.RSfetsym_0.QN.n2 frontAnalog_v0p0p1_12.RSfetsym_0.QN.n1 0.826818
R23701 frontAnalog_v0p0p1_12.RSfetsym_0.QN frontAnalog_v0p0p1_12.RSfetsym_0.QN.n0 0.74645
R23702 frontAnalog_v0p0p1_12.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_12.RSfetsym_0.QN.n3 0.249509
R23703 frontAnalog_v0p0p1_12.RSfetsym_0.QN.n3 frontAnalog_v0p0p1_12.RSfetsym_0.QN.n2 0.0968646
R23704 VL.n6 VL 0.23241
R23705 VL.n3 VL.t2 0.0203551
R23706 VL.n0 VL.t4 0.0203551
R23707 VL.n1 VL.n0 0.0203529
R23708 VL.n2 VL.n1 0.0203529
R23709 VL.n5 VL.n4 0.0203529
R23710 VL.n4 VL.n3 0.0203529
R23711 VL VL.n2 0.0111618
R23712 VL VL.n6 0.00913171
R23713 VL.n6 VL.n5 0.00105946
R23714 VL.n3 VL.t5 0.000502142
R23715 VL.n4 VL.t6 0.000502142
R23716 VL.n5 VL.t3 0.000502142
R23717 VL.n2 VL.t7 0.000502142
R23718 VL.n1 VL.t1 0.000502142
R23719 VL.n0 VL.t0 0.000502142
R23720 frontAnalog_v0p0p1_11.x65.A.n1 frontAnalog_v0p0p1_11.x65.A.t4 260.322
R23721 frontAnalog_v0p0p1_11.x65.A.n3 frontAnalog_v0p0p1_11.x65.A.t7 233.929
R23722 frontAnalog_v0p0p1_11.x65.A.n1 frontAnalog_v0p0p1_11.x65.A.t6 175.169
R23723 frontAnalog_v0p0p1_11.x65.A.n2 frontAnalog_v0p0p1_11.x65.A.t5 160.416
R23724 frontAnalog_v0p0p1_11.x65.A.n4 frontAnalog_v0p0p1_11.x65.A.t2 17.4109
R23725 frontAnalog_v0p0p1_11.x65.A.n4 frontAnalog_v0p0p1_11.x65.A.t3 10.2053
R23726 frontAnalog_v0p0p1_11.x65.A.n0 frontAnalog_v0p0p1_11.x65.A 2.78715
R23727 frontAnalog_v0p0p1_11.x65.A.n0 frontAnalog_v0p0p1_11.x65.A.n1 9.09103
R23728 frontAnalog_v0p0p1_11.x65.A.n6 frontAnalog_v0p0p1_11.x65.A.t0 7.94569
R23729 frontAnalog_v0p0p1_11.x65.A.n2 frontAnalog_v0p0p1_11.x65.A.t1 7.55846
R23730 frontAnalog_v0p0p1_11.x65.A.n5 frontAnalog_v0p0p1_11.x65.A.n3 1.4614
R23731 frontAnalog_v0p0p1_11.x65.A.n3 frontAnalog_v0p0p1_11.x65.A.n2 1.19626
R23732 frontAnalog_v0p0p1_11.x65.A.n6 frontAnalog_v0p0p1_11.x65.A.n5 0.836961
R23733 frontAnalog_v0p0p1_11.x65.A frontAnalog_v0p0p1_11.x65.A.n0 0.390342
R23734 frontAnalog_v0p0p1_11.x65.A.n5 frontAnalog_v0p0p1_11.x65.A.n4 0.154668
R23735 frontAnalog_v0p0p1_11.x65.A frontAnalog_v0p0p1_11.x65.A.n6 0.08175
R23736 VV8.n0 VV8.t17 167.365
R23737 VV8.n0 VV8.t16 92.4488
R23738 VV8.n1 VV8.n0 2.07493
R23739 VV8.n10 VV8 0.431333
R23740 VV8 VV8.n10 0.323625
R23741 VV8.n9 VV8.n8 0.141636
R23742 VV8.n8 VV8.n7 0.141636
R23743 VV8.n7 VV8.n6 0.141636
R23744 VV8.n6 VV8.n5 0.141636
R23745 VV8.n5 VV8.n4 0.141636
R23746 VV8.n4 VV8.n3 0.141636
R23747 VV8.n3 VV8.n2 0.141636
R23748 VV8.n1 VV8 0.12425
R23749 VV8 VV8.n9 0.100159
R23750 VV8 VV8.n1 0.0314375
R23751 VV8.n10 VV8 0.00833333
R23752 VV8.n10 VV8 0.006375
R23753 VV8.n3 VV8.t5 0.000502142
R23754 VV8.n4 VV8.t7 0.000502142
R23755 VV8.n5 VV8.t1 0.000502142
R23756 VV8.n6 VV8.t8 0.000502142
R23757 VV8.n7 VV8.t10 0.000502142
R23758 VV8.n8 VV8.t15 0.000502142
R23759 VV8.n9 VV8.t4 0.000502142
R23760 VV8.n2 VV8.t2 0.000502142
R23761 VV8.n3 VV8.t9 0.000502142
R23762 VV8.n4 VV8.t6 0.000502142
R23763 VV8.n5 VV8.t12 0.000502142
R23764 VV8.n6 VV8.t3 0.000502142
R23765 VV8.n7 VV8.t11 0.000502142
R23766 VV8.n8 VV8.t0 0.000502142
R23767 VV8.n9 VV8.t14 0.000502142
R23768 VV8.n2 VV8.t13 0.000502142
R23769 I12.n2 I12.t11 260.435
R23770 I12.n7 I12.t12 230.576
R23771 I12.n10 I12.t6 196.549
R23772 I12.n7 I12.t9 158.275
R23773 I12.n2 I12.t8 156.403
R23774 I12.n10 I12.t5 148.35
R23775 I12.n17 I12.t10 117.314
R23776 I12.n17 I12.t7 110.852
R23777 I12.n19 I12.t0 17.6181
R23778 I12.n20 I12.t3 14.2865
R23779 I12.n22 I12.t2 14.283
R23780 I12.n22 I12.t1 14.283
R23781 I12.n11 I12.n10 9.49829
R23782 I12 I12.n1 9.3005
R23783 I12.n24 I12.t4 8.77592
R23784 I12.n8 I12.n7 8.76429
R23785 I12.n12 I12.n11 7.9582
R23786 I12.n9 I12.n8 7.74345
R23787 I12.n3 I12.n2 7.60183
R23788 I12.n8 I12 6.66717
R23789 I12.n11 I12 6.44139
R23790 I12.n3 I12 4.8645
R23791 I12.n4 I12.n0 4.54557
R23792 I12.n1 I12.n0 4.51121
R23793 I12 I12.n25 3.93116
R23794 I12.n13 I12.n6 2.33638
R23795 I12.n24 I12.n23 1.20426
R23796 I12.n12 I12.n9 1.0005
R23797 I12.n26 I12 0.992722
R23798 I12.n14 I12 0.979667
R23799 I12 I12.n16 0.917
R23800 I12.n16 I12 0.82535
R23801 I12 I12.n26 0.447
R23802 I12.n13 I12.n12 0.446956
R23803 I12.n9 I12 0.380411
R23804 I12.n14 I12.n13 0.356917
R23805 I12.n25 I12.n24 0.336084
R23806 I12.n20 I12.n19 0.314673
R23807 I12.n21 I12.n20 0.300251
R23808 I12.n15 I12 0.2005
R23809 I12.n18 I12.n17 0.159555
R23810 I12.n23 I12.n22 0.106617
R23811 I12.n21 I12.n18 0.0796167
R23812 I12.n23 I12.n21 0.0480595
R23813 I12.n5 I12.n1 0.0344286
R23814 I12.n15 I12.n14 0.0287
R23815 I12.n16 I12.n15 0.0287
R23816 I12.n26 I12 0.0266111
R23817 I12.n26 I12 0.01225
R23818 I12.n25 I12 0.00658123
R23819 I12.n6 I12.n0 0.00182856
R23820 I12.n6 I12.n5 0.00149885
R23821 I12.n4 I12.n3 0.00133362
R23822 I12.n5 I12.n4 0.00100077
R23823 I12.n19 I12.n18 0.000504658
R23824 frontAnalog_v0p0p1_1.x63.A.n2 frontAnalog_v0p0p1_1.x63.A.t7 260.322
R23825 frontAnalog_v0p0p1_1.x63.A.n4 frontAnalog_v0p0p1_1.x63.A.t4 233.888
R23826 frontAnalog_v0p0p1_1.x63.A.n2 frontAnalog_v0p0p1_1.x63.A.t6 175.169
R23827 frontAnalog_v0p0p1_1.x63.A.n3 frontAnalog_v0p0p1_1.x63.A.t5 159.725
R23828 frontAnalog_v0p0p1_1.x63.A.n1 frontAnalog_v0p0p1_1.x63.A.t0 17.4109
R23829 frontAnalog_v0p0p1_1.x63.A.n0 frontAnalog_v0p0p1_1.x63.A.n2 9.75129
R23830 frontAnalog_v0p0p1_1.x63.A.n1 frontAnalog_v0p0p1_1.x63.A.t1 9.6027
R23831 frontAnalog_v0p0p1_1.x63.A.n0 frontAnalog_v0p0p1_1.x63.A 2.33338
R23832 frontAnalog_v0p0p1_1.x63.A.n5 frontAnalog_v0p0p1_1.x63.A.t3 8.40929
R23833 frontAnalog_v0p0p1_1.x63.A.n3 frontAnalog_v0p0p1_1.x63.A.t2 8.06629
R23834 frontAnalog_v0p0p1_1.x63.A.n4 frontAnalog_v0p0p1_1.x63.A.n3 1.73501
R23835 frontAnalog_v0p0p1_1.x63.A.n1 frontAnalog_v0p0p1_1.x63.A.n4 0.99025
R23836 frontAnalog_v0p0p1_1.x63.A.n5 frontAnalog_v0p0p1_1.x63.A.n1 0.853186
R23837 frontAnalog_v0p0p1_1.x63.A frontAnalog_v0p0p1_1.x63.A.n0 0.349517
R23838 frontAnalog_v0p0p1_1.x63.A frontAnalog_v0p0p1_1.x63.A.n5 0.24425
R23839 frontAnalog_v0p0p1_5.x65.A.n1 frontAnalog_v0p0p1_5.x65.A.t4 260.322
R23840 frontAnalog_v0p0p1_5.x65.A.n4 frontAnalog_v0p0p1_5.x65.A.t7 233.929
R23841 frontAnalog_v0p0p1_5.x65.A.n1 frontAnalog_v0p0p1_5.x65.A.t6 175.169
R23842 frontAnalog_v0p0p1_5.x65.A.n3 frontAnalog_v0p0p1_5.x65.A.t5 160.416
R23843 frontAnalog_v0p0p1_5.x65.A.n2 frontAnalog_v0p0p1_5.x65.A.t2 17.4109
R23844 frontAnalog_v0p0p1_5.x65.A.n2 frontAnalog_v0p0p1_5.x65.A.t3 10.2053
R23845 frontAnalog_v0p0p1_5.x65.A.n0 frontAnalog_v0p0p1_5.x65.A 2.78715
R23846 frontAnalog_v0p0p1_5.x65.A.n0 frontAnalog_v0p0p1_5.x65.A.n1 9.09103
R23847 frontAnalog_v0p0p1_5.x65.A.n6 frontAnalog_v0p0p1_5.x65.A.t1 7.94569
R23848 frontAnalog_v0p0p1_5.x65.A.n3 frontAnalog_v0p0p1_5.x65.A.t0 7.55846
R23849 frontAnalog_v0p0p1_5.x65.A.n5 frontAnalog_v0p0p1_5.x65.A.n4 1.4614
R23850 frontAnalog_v0p0p1_5.x65.A.n4 frontAnalog_v0p0p1_5.x65.A.n3 1.19626
R23851 frontAnalog_v0p0p1_5.x65.A.n6 frontAnalog_v0p0p1_5.x65.A.n5 0.836961
R23852 frontAnalog_v0p0p1_5.x65.A frontAnalog_v0p0p1_5.x65.A.n0 0.390342
R23853 frontAnalog_v0p0p1_5.x65.A.n5 frontAnalog_v0p0p1_5.x65.A.n2 0.154668
R23854 frontAnalog_v0p0p1_5.x65.A frontAnalog_v0p0p1_5.x65.A.n6 0.08175
R23855 frontAnalog_v0p0p1_14.RSfetsym_0.QN.n1 frontAnalog_v0p0p1_14.RSfetsym_0.QN.t6 117.511
R23856 frontAnalog_v0p0p1_14.RSfetsym_0.QN.n1 frontAnalog_v0p0p1_14.RSfetsym_0.QN.t5 110.698
R23857 frontAnalog_v0p0p1_14.RSfetsym_0.QN.n2 frontAnalog_v0p0p1_14.RSfetsym_0.QN.t2 19.1963
R23858 frontAnalog_v0p0p1_14.RSfetsym_0.QN.n3 frontAnalog_v0p0p1_14.RSfetsym_0.QN.t1 14.5206
R23859 frontAnalog_v0p0p1_14.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_14.RSfetsym_0.QN.t3 14.283
R23860 frontAnalog_v0p0p1_14.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_14.RSfetsym_0.QN.t4 14.283
R23861 frontAnalog_v0p0p1_14.RSfetsym_0.QN frontAnalog_v0p0p1_14.RSfetsym_0.QN.t0 9.14075
R23862 frontAnalog_v0p0p1_14.RSfetsym_0.QN.n2 frontAnalog_v0p0p1_14.RSfetsym_0.QN.n1 0.826818
R23863 frontAnalog_v0p0p1_14.RSfetsym_0.QN frontAnalog_v0p0p1_14.RSfetsym_0.QN.n0 0.74645
R23864 frontAnalog_v0p0p1_14.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_14.RSfetsym_0.QN.n3 0.249509
R23865 frontAnalog_v0p0p1_14.RSfetsym_0.QN.n3 frontAnalog_v0p0p1_14.RSfetsym_0.QN.n2 0.0968646
R23866 frontAnalog_v0p0p1_7.RSfetsym_0.QN.n1 frontAnalog_v0p0p1_7.RSfetsym_0.QN.t6 117.511
R23867 frontAnalog_v0p0p1_7.RSfetsym_0.QN.n1 frontAnalog_v0p0p1_7.RSfetsym_0.QN.t5 110.698
R23868 frontAnalog_v0p0p1_7.RSfetsym_0.QN.n2 frontAnalog_v0p0p1_7.RSfetsym_0.QN.t2 19.1963
R23869 frontAnalog_v0p0p1_7.RSfetsym_0.QN.n3 frontAnalog_v0p0p1_7.RSfetsym_0.QN.t0 14.5206
R23870 frontAnalog_v0p0p1_7.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_7.RSfetsym_0.QN.t3 14.283
R23871 frontAnalog_v0p0p1_7.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_7.RSfetsym_0.QN.t4 14.283
R23872 frontAnalog_v0p0p1_7.RSfetsym_0.QN frontAnalog_v0p0p1_7.RSfetsym_0.QN.t1 9.14075
R23873 frontAnalog_v0p0p1_7.RSfetsym_0.QN.n2 frontAnalog_v0p0p1_7.RSfetsym_0.QN.n1 0.826818
R23874 frontAnalog_v0p0p1_7.RSfetsym_0.QN frontAnalog_v0p0p1_7.RSfetsym_0.QN.n0 0.74645
R23875 frontAnalog_v0p0p1_7.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_7.RSfetsym_0.QN.n3 0.249509
R23876 frontAnalog_v0p0p1_7.RSfetsym_0.QN.n3 frontAnalog_v0p0p1_7.RSfetsym_0.QN.n2 0.0968646
R23877 frontAnalog_v0p0p1_0.RSfetsym_0.QN.n1 frontAnalog_v0p0p1_0.RSfetsym_0.QN.t5 117.511
R23878 frontAnalog_v0p0p1_0.RSfetsym_0.QN.n1 frontAnalog_v0p0p1_0.RSfetsym_0.QN.t6 110.698
R23879 frontAnalog_v0p0p1_0.RSfetsym_0.QN.n2 frontAnalog_v0p0p1_0.RSfetsym_0.QN.t2 19.1963
R23880 frontAnalog_v0p0p1_0.RSfetsym_0.QN.n3 frontAnalog_v0p0p1_0.RSfetsym_0.QN.t3 14.5206
R23881 frontAnalog_v0p0p1_0.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_0.RSfetsym_0.QN.t1 14.283
R23882 frontAnalog_v0p0p1_0.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_0.RSfetsym_0.QN.t0 14.283
R23883 frontAnalog_v0p0p1_0.RSfetsym_0.QN frontAnalog_v0p0p1_0.RSfetsym_0.QN.t4 9.14075
R23884 frontAnalog_v0p0p1_0.RSfetsym_0.QN.n2 frontAnalog_v0p0p1_0.RSfetsym_0.QN.n1 0.826818
R23885 frontAnalog_v0p0p1_0.RSfetsym_0.QN frontAnalog_v0p0p1_0.RSfetsym_0.QN.n0 0.74645
R23886 frontAnalog_v0p0p1_0.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_0.RSfetsym_0.QN.n3 0.249509
R23887 frontAnalog_v0p0p1_0.RSfetsym_0.QN.n3 frontAnalog_v0p0p1_0.RSfetsym_0.QN.n2 0.0968646
R23888 I8.n0 I8.t8 196.549
R23889 I8.n0 I8.t6 148.35
R23890 I8.n4 I8.t7 117.314
R23891 I8.n4 I8.t5 110.853
R23892 I8.n6 I8.t0 17.6181
R23893 I8.n7 I8.t3 14.2865
R23894 I8.n9 I8.t1 14.283
R23895 I8.n9 I8.t2 14.283
R23896 I8.n1 I8.n0 9.49592
R23897 I8.n11 I8.t4 8.77744
R23898 I8.n2 I8.n1 7.58085
R23899 I8.n1 I8 6.44187
R23900 I8.n3 I8.n2 2.34543
R23901 I8.n11 I8.n10 1.20426
R23902 I8.n2 I8 0.88934
R23903 I8 I8.n11 0.357737
R23904 I8 I8.n3 0.336158
R23905 I8.n7 I8.n6 0.314673
R23906 I8.n8 I8.n7 0.299251
R23907 I8.n3 I8 0.200892
R23908 I8.n5 I8.n4 0.159555
R23909 I8.n10 I8.n9 0.106617
R23910 I8.n8 I8.n5 0.0796167
R23911 I8.n10 I8.n8 0.0480595
R23912 I8.n6 I8.n5 0.000504658
R23913 frontAnalog_v0p0p1_13.x65.A.n1 frontAnalog_v0p0p1_13.x65.A.t4 260.322
R23914 frontAnalog_v0p0p1_13.x65.A.n3 frontAnalog_v0p0p1_13.x65.A.t7 233.929
R23915 frontAnalog_v0p0p1_13.x65.A.n1 frontAnalog_v0p0p1_13.x65.A.t6 175.169
R23916 frontAnalog_v0p0p1_13.x65.A.n2 frontAnalog_v0p0p1_13.x65.A.t5 160.416
R23917 frontAnalog_v0p0p1_13.x65.A.n4 frontAnalog_v0p0p1_13.x65.A.t1 17.4109
R23918 frontAnalog_v0p0p1_13.x65.A.n4 frontAnalog_v0p0p1_13.x65.A.t0 10.2053
R23919 frontAnalog_v0p0p1_13.x65.A.n0 frontAnalog_v0p0p1_13.x65.A 2.78715
R23920 frontAnalog_v0p0p1_13.x65.A.n0 frontAnalog_v0p0p1_13.x65.A.n1 9.09103
R23921 frontAnalog_v0p0p1_13.x65.A.n6 frontAnalog_v0p0p1_13.x65.A.t2 7.94569
R23922 frontAnalog_v0p0p1_13.x65.A.n2 frontAnalog_v0p0p1_13.x65.A.t3 7.55846
R23923 frontAnalog_v0p0p1_13.x65.A.n5 frontAnalog_v0p0p1_13.x65.A.n3 1.4614
R23924 frontAnalog_v0p0p1_13.x65.A.n3 frontAnalog_v0p0p1_13.x65.A.n2 1.19626
R23925 frontAnalog_v0p0p1_13.x65.A.n6 frontAnalog_v0p0p1_13.x65.A.n5 0.836961
R23926 frontAnalog_v0p0p1_13.x65.A frontAnalog_v0p0p1_13.x65.A.n0 0.390342
R23927 frontAnalog_v0p0p1_13.x65.A.n5 frontAnalog_v0p0p1_13.x65.A.n4 0.154668
R23928 frontAnalog_v0p0p1_13.x65.A frontAnalog_v0p0p1_13.x65.A.n6 0.08175
R23929 frontAnalog_v0p0p1_11.RSfetsym_0.QN.n1 frontAnalog_v0p0p1_11.RSfetsym_0.QN.t6 117.511
R23930 frontAnalog_v0p0p1_11.RSfetsym_0.QN.n1 frontAnalog_v0p0p1_11.RSfetsym_0.QN.t5 110.698
R23931 frontAnalog_v0p0p1_11.RSfetsym_0.QN.n2 frontAnalog_v0p0p1_11.RSfetsym_0.QN.t4 19.1963
R23932 frontAnalog_v0p0p1_11.RSfetsym_0.QN.n3 frontAnalog_v0p0p1_11.RSfetsym_0.QN.t0 14.5206
R23933 frontAnalog_v0p0p1_11.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_11.RSfetsym_0.QN.t2 14.283
R23934 frontAnalog_v0p0p1_11.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_11.RSfetsym_0.QN.t3 14.283
R23935 frontAnalog_v0p0p1_11.RSfetsym_0.QN frontAnalog_v0p0p1_11.RSfetsym_0.QN.t1 9.14075
R23936 frontAnalog_v0p0p1_11.RSfetsym_0.QN.n2 frontAnalog_v0p0p1_11.RSfetsym_0.QN.n1 0.826818
R23937 frontAnalog_v0p0p1_11.RSfetsym_0.QN frontAnalog_v0p0p1_11.RSfetsym_0.QN.n0 0.74645
R23938 frontAnalog_v0p0p1_11.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_11.RSfetsym_0.QN.n3 0.249509
R23939 frontAnalog_v0p0p1_11.RSfetsym_0.QN.n3 frontAnalog_v0p0p1_11.RSfetsym_0.QN.n2 0.0968646
R23940 frontAnalog_v0p0p1_12.x63.A.n2 frontAnalog_v0p0p1_12.x63.A.t4 260.322
R23941 frontAnalog_v0p0p1_12.x63.A.n4 frontAnalog_v0p0p1_12.x63.A.t5 233.888
R23942 frontAnalog_v0p0p1_12.x63.A.n2 frontAnalog_v0p0p1_12.x63.A.t6 175.169
R23943 frontAnalog_v0p0p1_12.x63.A.n3 frontAnalog_v0p0p1_12.x63.A.t7 159.725
R23944 frontAnalog_v0p0p1_12.x63.A.n1 frontAnalog_v0p0p1_12.x63.A.t3 17.4109
R23945 frontAnalog_v0p0p1_12.x63.A.n0 frontAnalog_v0p0p1_12.x63.A.n2 9.75129
R23946 frontAnalog_v0p0p1_12.x63.A.n1 frontAnalog_v0p0p1_12.x63.A.t2 9.6037
R23947 frontAnalog_v0p0p1_12.x63.A.n0 frontAnalog_v0p0p1_12.x63.A 2.33338
R23948 frontAnalog_v0p0p1_12.x63.A.n5 frontAnalog_v0p0p1_12.x63.A.t0 8.40929
R23949 frontAnalog_v0p0p1_12.x63.A.n3 frontAnalog_v0p0p1_12.x63.A.t1 8.06629
R23950 frontAnalog_v0p0p1_12.x63.A.n4 frontAnalog_v0p0p1_12.x63.A.n3 1.73501
R23951 frontAnalog_v0p0p1_12.x63.A.n1 frontAnalog_v0p0p1_12.x63.A.n4 0.99025
R23952 frontAnalog_v0p0p1_12.x63.A.n5 frontAnalog_v0p0p1_12.x63.A.n1 0.853186
R23953 frontAnalog_v0p0p1_12.x63.A frontAnalog_v0p0p1_12.x63.A.n0 0.349517
R23954 frontAnalog_v0p0p1_12.x63.A frontAnalog_v0p0p1_12.x63.A.n5 0.24425
R23955 frontAnalog_v0p0p1_4.RSfetsym_0.QN.n1 frontAnalog_v0p0p1_4.RSfetsym_0.QN.t6 117.511
R23956 frontAnalog_v0p0p1_4.RSfetsym_0.QN.n1 frontAnalog_v0p0p1_4.RSfetsym_0.QN.t5 110.698
R23957 frontAnalog_v0p0p1_4.RSfetsym_0.QN.n2 frontAnalog_v0p0p1_4.RSfetsym_0.QN.t0 19.1963
R23958 frontAnalog_v0p0p1_4.RSfetsym_0.QN.n3 frontAnalog_v0p0p1_4.RSfetsym_0.QN.t4 14.5206
R23959 frontAnalog_v0p0p1_4.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_4.RSfetsym_0.QN.t1 14.283
R23960 frontAnalog_v0p0p1_4.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_4.RSfetsym_0.QN.t2 14.283
R23961 frontAnalog_v0p0p1_4.RSfetsym_0.QN frontAnalog_v0p0p1_4.RSfetsym_0.QN.t3 9.14075
R23962 frontAnalog_v0p0p1_4.RSfetsym_0.QN.n2 frontAnalog_v0p0p1_4.RSfetsym_0.QN.n1 0.826818
R23963 frontAnalog_v0p0p1_4.RSfetsym_0.QN frontAnalog_v0p0p1_4.RSfetsym_0.QN.n0 0.74645
R23964 frontAnalog_v0p0p1_4.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_4.RSfetsym_0.QN.n3 0.249509
R23965 frontAnalog_v0p0p1_4.RSfetsym_0.QN.n3 frontAnalog_v0p0p1_4.RSfetsym_0.QN.n2 0.0968646
R23966 I7.n4 I7.t5 261.116
R23967 I7.n0 I7.t7 186.03
R23968 I7.n4 I7.t10 155.746
R23969 I7.n0 I7.t8 137.829
R23970 I7.n12 I7.t6 117.314
R23971 I7.n12 I7.t9 110.852
R23972 I7 I7.n0 78.5605
R23973 I7.n9 I7 47.2619
R23974 I7.n14 I7.t1 17.6181
R23975 I7.n15 I7.t0 14.2865
R23976 I7.n17 I7.t3 14.283
R23977 I7.n17 I7.t2 14.283
R23978 I7.n6 I7.n5 9.3005
R23979 I7.n19 I7.t4 8.77592
R23980 I7.n5 I7.n4 7.65549
R23981 I7.n5 I7.n2 4.64342
R23982 I7.n2 I7.n1 4.52687
R23983 I7.n6 I7.n1 4.513
R23984 I7.n9 I7.n8 4.04922
R23985 I7.n3 I7 2.46419
R23986 I7.n19 I7.n18 1.20426
R23987 I7.n10 I7 0.808983
R23988 I7.n5 I7.n3 0.754023
R23989 I7 I7.n11 0.748897
R23990 I7.n21 I7 0.713803
R23991 I7 I7.n21 0.711434
R23992 I7.n11 I7.n10 0.674526
R23993 I7.n10 I7.n9 0.478179
R23994 I7 I7.n20 0.462023
R23995 I7.n20 I7.n19 0.32511
R23996 I7.n15 I7.n14 0.314673
R23997 I7.n16 I7.n15 0.300251
R23998 I7.n11 I7 0.20675
R23999 I7.n13 I7.n12 0.159555
R24000 I7.n18 I7.n17 0.106617
R24001 I7.n16 I7.n13 0.0796167
R24002 I7.n21 I7 0.0626967
R24003 I7.n21 I7 0.06249
R24004 I7.n18 I7.n16 0.0480595
R24005 I7.n20 I7 0.046937
R24006 I7.n7 I7.n6 0.0326429
R24007 I7.n7 I7.n2 0.0197253
R24008 I7.n8 I7.n1 0.00182856
R24009 I7.n8 I7.n7 0.00149885
R24010 I7.n7 I7.n3 0.00125261
R24011 I7.n14 I7.n13 0.000504658
R24012 frontAnalog_v0p0p1_11.x63.A.n2 frontAnalog_v0p0p1_11.x63.A.t5 260.322
R24013 frontAnalog_v0p0p1_11.x63.A.n4 frontAnalog_v0p0p1_11.x63.A.t6 233.888
R24014 frontAnalog_v0p0p1_11.x63.A.n2 frontAnalog_v0p0p1_11.x63.A.t7 175.169
R24015 frontAnalog_v0p0p1_11.x63.A.n3 frontAnalog_v0p0p1_11.x63.A.t4 159.725
R24016 frontAnalog_v0p0p1_11.x63.A.n1 frontAnalog_v0p0p1_11.x63.A.t2 17.4109
R24017 frontAnalog_v0p0p1_11.x63.A.n0 frontAnalog_v0p0p1_11.x63.A.n2 9.75129
R24018 frontAnalog_v0p0p1_11.x63.A.n1 frontAnalog_v0p0p1_11.x63.A.t3 9.6037
R24019 frontAnalog_v0p0p1_11.x63.A.n0 frontAnalog_v0p0p1_11.x63.A 2.33338
R24020 frontAnalog_v0p0p1_11.x63.A.n5 frontAnalog_v0p0p1_11.x63.A.t1 8.40929
R24021 frontAnalog_v0p0p1_11.x63.A.n3 frontAnalog_v0p0p1_11.x63.A.t0 8.06629
R24022 frontAnalog_v0p0p1_11.x63.A.n4 frontAnalog_v0p0p1_11.x63.A.n3 1.73501
R24023 frontAnalog_v0p0p1_11.x63.A.n1 frontAnalog_v0p0p1_11.x63.A.n4 0.99025
R24024 frontAnalog_v0p0p1_11.x63.A.n5 frontAnalog_v0p0p1_11.x63.A.n1 0.853186
R24025 frontAnalog_v0p0p1_11.x63.A frontAnalog_v0p0p1_11.x63.A.n0 0.349517
R24026 frontAnalog_v0p0p1_11.x63.A frontAnalog_v0p0p1_11.x63.A.n5 0.24425
R24027 frontAnalog_v0p0p1_8.x65.A.n1 frontAnalog_v0p0p1_8.x65.A.t4 260.322
R24028 frontAnalog_v0p0p1_8.x65.A.n4 frontAnalog_v0p0p1_8.x65.A.t7 233.929
R24029 frontAnalog_v0p0p1_8.x65.A.n1 frontAnalog_v0p0p1_8.x65.A.t6 175.169
R24030 frontAnalog_v0p0p1_8.x65.A.n3 frontAnalog_v0p0p1_8.x65.A.t5 160.416
R24031 frontAnalog_v0p0p1_8.x65.A.n2 frontAnalog_v0p0p1_8.x65.A.t3 17.4109
R24032 frontAnalog_v0p0p1_8.x65.A.n2 frontAnalog_v0p0p1_8.x65.A.t2 10.2053
R24033 frontAnalog_v0p0p1_8.x65.A.n0 frontAnalog_v0p0p1_8.x65.A 2.78715
R24034 frontAnalog_v0p0p1_8.x65.A.n0 frontAnalog_v0p0p1_8.x65.A.n1 9.09103
R24035 frontAnalog_v0p0p1_8.x65.A.n6 frontAnalog_v0p0p1_8.x65.A.t1 7.94569
R24036 frontAnalog_v0p0p1_8.x65.A.n3 frontAnalog_v0p0p1_8.x65.A.t0 7.55846
R24037 frontAnalog_v0p0p1_8.x65.A.n5 frontAnalog_v0p0p1_8.x65.A.n4 1.4614
R24038 frontAnalog_v0p0p1_8.x65.A.n4 frontAnalog_v0p0p1_8.x65.A.n3 1.19626
R24039 frontAnalog_v0p0p1_8.x65.A.n6 frontAnalog_v0p0p1_8.x65.A.n5 0.836961
R24040 frontAnalog_v0p0p1_8.x65.A frontAnalog_v0p0p1_8.x65.A.n0 0.390342
R24041 frontAnalog_v0p0p1_8.x65.A.n5 frontAnalog_v0p0p1_8.x65.A.n2 0.154668
R24042 frontAnalog_v0p0p1_8.x65.A frontAnalog_v0p0p1_8.x65.A.n6 0.08175
R24043 I14.n17 I14.t11 260.435
R24044 I14.n2 I14.t12 229.433
R24045 I14.n12 I14.t9 196.549
R24046 I14.n2 I14.t6 158.886
R24047 I14.n17 I14.t5 156.403
R24048 I14.n12 I14.t7 148.35
R24049 I14.n27 I14.t10 117.314
R24050 I14.n27 I14.t8 110.852
R24051 I14.n13 I14.n12 76.0005
R24052 I14.n29 I14.t0 17.6181
R24053 I14.n30 I14.t4 14.2865
R24054 I14.n32 I14.t1 14.283
R24055 I14.n32 I14.t2 14.283
R24056 I14 I14.n16 9.3005
R24057 I14.n5 I14.n3 9.3005
R24058 I14.n5 I14.n4 9.3005
R24059 I14.n9 I14.n8 9.3005
R24060 I14.n34 I14.t3 8.77592
R24061 I14.n18 I14.n17 7.60183
R24062 I14.n3 I14.n2 7.39078
R24063 I14.n22 I14.n14 6.24391
R24064 I14.n13 I14 5.78114
R24065 I14.n18 I14 4.8645
R24066 I14.n19 I14.n15 4.54557
R24067 I14.n10 I14.n9 4.51698
R24068 I14.n16 I14.n15 4.51121
R24069 I14.n8 I14.n7 4.5005
R24070 I14.n22 I14.n21 3.53643
R24071 I14.n14 I14.n13 3.51018
R24072 I14.n8 I14.n4 3.46717
R24073 I14.n34 I14.n33 1.20426
R24074 I14.n6 I14.n0 1.13339
R24075 I14.n11 I14.n10 1.11384
R24076 I14.n8 I14.n3 1.06717
R24077 I14.n4 I14 1.06717
R24078 I14.n23 I14.n11 0.767464
R24079 I14.n35 I14 0.731611
R24080 I14.n24 I14 0.718556
R24081 I14 I14.n26 0.655889
R24082 I14.n26 I14 0.59035
R24083 I14.n24 I14.n23 0.503793
R24084 I14.n11 I14 0.372375
R24085 I14 I14.n34 0.370547
R24086 I14.n23 I14.n22 0.321929
R24087 I14.n30 I14.n29 0.314673
R24088 I14.n31 I14.n30 0.300251
R24089 I14 I14.n35 0.299591
R24090 I14.n14 I14 0.206952
R24091 I14.n25 I14 0.2005
R24092 I14.n28 I14.n27 0.159555
R24093 I14.n33 I14.n32 0.106617
R24094 I14.n31 I14.n28 0.0796167
R24095 I14.n33 I14.n31 0.0480595
R24096 I14.n20 I14.n16 0.0344286
R24097 I14.n25 I14.n24 0.0287
R24098 I14.n26 I14.n25 0.0287
R24099 I14.n10 I14.n0 0.028
R24100 I14.n35 I14 0.0266111
R24101 I14.n9 I14.n1 0.0142363
R24102 I14.n35 I14 0.0111818
R24103 I14.n7 I14.n1 0.00599451
R24104 I14.n6 I14.n5 0.00409723
R24105 I14.n7 I14.n6 0.00202085
R24106 I14.n21 I14.n15 0.00182856
R24107 I14.n21 I14.n20 0.00149885
R24108 I14.n19 I14.n18 0.00133362
R24109 I14.n20 I14.n19 0.00100077
R24110 I14.n1 I14.n0 0.000617139
R24111 I14.n29 I14.n28 0.000504658
R24112 I15.n4 I15.t5 261.116
R24113 I15.n0 I15.t7 186.03
R24114 I15.n4 I15.t9 155.746
R24115 I15.n0 I15.t6 137.829
R24116 I15.n14 I15.t10 117.314
R24117 I15.n14 I15.t8 110.852
R24118 I15 I15.n0 78.5605
R24119 I15.n9 I15 47.2619
R24120 I15.n16 I15.t0 17.6181
R24121 I15.n17 I15.t3 14.2865
R24122 I15.n19 I15.t2 14.283
R24123 I15.n19 I15.t1 14.283
R24124 I15.n6 I15.n5 9.3005
R24125 I15.n21 I15.t4 8.77592
R24126 I15.n5 I15.n4 7.65549
R24127 I15.n5 I15.n2 4.64342
R24128 I15.n2 I15.n1 4.52687
R24129 I15.n6 I15.n1 4.513
R24130 I15.n9 I15.n8 4.04922
R24131 I15.n3 I15 2.46419
R24132 I15.n21 I15.n20 1.20426
R24133 I15.n5 I15.n3 0.754023
R24134 I15.n10 I15 0.70184
R24135 I15.n11 I15.n10 0.662978
R24136 I15.n10 I15.n9 0.585321
R24137 I15.n11 I15 0.577556
R24138 I15.n22 I15 0.559278
R24139 I15 I15.n13 0.514889
R24140 I15.n13 I15 0.46345
R24141 I15 I15.n21 0.370547
R24142 I15.n17 I15.n16 0.314673
R24143 I15.n18 I15.n17 0.300251
R24144 I15 I15.n22 0.25195
R24145 I15.n12 I15 0.2005
R24146 I15.n15 I15.n14 0.159555
R24147 I15.n20 I15.n19 0.106617
R24148 I15.n18 I15.n15 0.0796167
R24149 I15.n20 I15.n18 0.0480595
R24150 I15.n7 I15.n6 0.0326429
R24151 I15.n12 I15.n11 0.0287
R24152 I15.n13 I15.n12 0.0287
R24153 I15.n22 I15 0.0266111
R24154 I15.n7 I15.n2 0.0197253
R24155 I15.n22 I15 0.01225
R24156 I15.n8 I15.n1 0.00182856
R24157 I15.n8 I15.n7 0.00149885
R24158 I15.n7 I15.n3 0.00125261
R24159 I15.n16 I15.n15 0.000504658
R24160 I3.n4 I3.t7 334.723
R24161 I3.n3 I3.t10 323.342
R24162 I3.n4 I3.t9 206.19
R24163 I3.n3 I3.t6 194.809
R24164 I3.n0 I3.t5 186.03
R24165 I3.n0 I3.t11 137.829
R24166 I3.n8 I3.t12 117.314
R24167 I3.n8 I3.t8 110.853
R24168 I3 I3.n4 84.2291
R24169 I3 I3.n3 82.1338
R24170 I3.n1 I3.n0 76.0005
R24171 I3.n2 I3 66.7187
R24172 I3.n5 I3 26.4877
R24173 I3.n10 I3.t1 17.6181
R24174 I3.n11 I3.t4 14.2865
R24175 I3.n13 I3.t2 14.283
R24176 I3.n13 I3.t3 14.283
R24177 I3.n15 I3.t0 8.77744
R24178 I3.n1 I3 7.31479
R24179 I3 I3.n16 5.79898
R24180 I3.n5 I3 4.36044
R24181 I3 I3.n1 4.02336
R24182 I3.n6 I3.n5 2.61211
R24183 I3.n6 I3.n2 1.25943
R24184 I3.n15 I3.n14 1.20426
R24185 I3.n2 I3 0.969697
R24186 I3.n17 I3 0.431333
R24187 I3 I3.n7 0.420367
R24188 I3.n16 I3.n15 0.32511
R24189 I3 I3.n17 0.323625
R24190 I3.n11 I3.n10 0.314673
R24191 I3.n7 I3.n6 0.300322
R24192 I3.n12 I3.n11 0.299251
R24193 I3.n7 I3 0.20675
R24194 I3.n9 I3.n8 0.159555
R24195 I3.n14 I3.n13 0.106617
R24196 I3.n12 I3.n9 0.0796167
R24197 I3.n14 I3.n12 0.0480595
R24198 I3.n16 I3 0.046937
R24199 I3.n17 I3 0.0161667
R24200 I3.n17 I3 0.01225
R24201 I3.n10 I3.n9 0.000504658
R24202 frontAnalog_v0p0p1_1.RSfetsym_0.QN.n1 frontAnalog_v0p0p1_1.RSfetsym_0.QN.t6 117.511
R24203 frontAnalog_v0p0p1_1.RSfetsym_0.QN.n1 frontAnalog_v0p0p1_1.RSfetsym_0.QN.t5 110.698
R24204 frontAnalog_v0p0p1_1.RSfetsym_0.QN.n2 frontAnalog_v0p0p1_1.RSfetsym_0.QN.t1 19.1963
R24205 frontAnalog_v0p0p1_1.RSfetsym_0.QN.n3 frontAnalog_v0p0p1_1.RSfetsym_0.QN.t4 14.5206
R24206 frontAnalog_v0p0p1_1.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_1.RSfetsym_0.QN.t3 14.283
R24207 frontAnalog_v0p0p1_1.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_1.RSfetsym_0.QN.t2 14.283
R24208 frontAnalog_v0p0p1_1.RSfetsym_0.QN frontAnalog_v0p0p1_1.RSfetsym_0.QN.t0 9.14075
R24209 frontAnalog_v0p0p1_1.RSfetsym_0.QN.n2 frontAnalog_v0p0p1_1.RSfetsym_0.QN.n1 0.826818
R24210 frontAnalog_v0p0p1_1.RSfetsym_0.QN frontAnalog_v0p0p1_1.RSfetsym_0.QN.n0 0.74645
R24211 frontAnalog_v0p0p1_1.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_1.RSfetsym_0.QN.n3 0.249509
R24212 frontAnalog_v0p0p1_1.RSfetsym_0.QN.n3 frontAnalog_v0p0p1_1.RSfetsym_0.QN.n2 0.0968646
R24213 I11.n4 I11.t7 334.723
R24214 I11.n3 I11.t9 323.342
R24215 I11.n4 I11.t11 206.19
R24216 I11.n3 I11.t6 194.809
R24217 I11.n0 I11.t5 186.03
R24218 I11.n0 I11.t10 137.829
R24219 I11.n10 I11.t12 117.314
R24220 I11.n10 I11.t8 110.852
R24221 I11 I11.n4 84.2291
R24222 I11 I11.n3 82.1338
R24223 I11.n1 I11.n0 76.0005
R24224 I11.n2 I11 66.7187
R24225 I11.n5 I11 26.4877
R24226 I11.n12 I11.t0 17.6181
R24227 I11.n13 I11.t3 14.2865
R24228 I11.n15 I11.t1 14.283
R24229 I11.n15 I11.t2 14.283
R24230 I11.n17 I11.t4 8.77592
R24231 I11.n1 I11 7.31479
R24232 I11.n5 I11 4.36044
R24233 I11 I11.n1 4.02336
R24234 I11 I11.n18 3.30508
R24235 I11.n6 I11.n5 2.71925
R24236 I11.n17 I11.n16 1.20426
R24237 I11.n19 I11 1.17028
R24238 I11.n6 I11.n2 1.15229
R24239 I11.n7 I11 1.14156
R24240 I11 I11.n9 1.07889
R24241 I11.n9 I11 0.97105
R24242 I11.n2 I11 0.969697
R24243 I11 I11.n19 0.957591
R24244 I11.n18 I11.n17 0.33431
R24245 I11.n13 I11.n12 0.314673
R24246 I11.n14 I11.n13 0.300251
R24247 I11.n7 I11.n6 0.28348
R24248 I11.n8 I11 0.2005
R24249 I11.n11 I11.n10 0.159555
R24250 I11.n16 I11.n15 0.106617
R24251 I11.n14 I11.n11 0.0796167
R24252 I11.n16 I11.n14 0.0480595
R24253 I11.n8 I11.n7 0.0287
R24254 I11.n9 I11.n8 0.0287
R24255 I11.n19 I11 0.0109444
R24256 I11.n19 I11 0.00904545
R24257 I11.n18 I11 0.0087668
R24258 I11.n12 I11.n11 0.000504658
R24259 frontAnalog_v0p0p1_8.x63.A.n2 frontAnalog_v0p0p1_8.x63.A.t5 260.322
R24260 frontAnalog_v0p0p1_8.x63.A.n4 frontAnalog_v0p0p1_8.x63.A.t6 233.888
R24261 frontAnalog_v0p0p1_8.x63.A.n2 frontAnalog_v0p0p1_8.x63.A.t7 175.169
R24262 frontAnalog_v0p0p1_8.x63.A.n3 frontAnalog_v0p0p1_8.x63.A.t4 159.725
R24263 frontAnalog_v0p0p1_8.x63.A.n1 frontAnalog_v0p0p1_8.x63.A.t2 17.4109
R24264 frontAnalog_v0p0p1_8.x63.A.n0 frontAnalog_v0p0p1_8.x63.A.n2 9.75129
R24265 frontAnalog_v0p0p1_8.x63.A.n1 frontAnalog_v0p0p1_8.x63.A.t3 9.6037
R24266 frontAnalog_v0p0p1_8.x63.A.n0 frontAnalog_v0p0p1_8.x63.A 2.33338
R24267 frontAnalog_v0p0p1_8.x63.A.n5 frontAnalog_v0p0p1_8.x63.A.t0 8.40929
R24268 frontAnalog_v0p0p1_8.x63.A.n3 frontAnalog_v0p0p1_8.x63.A.t1 8.06629
R24269 frontAnalog_v0p0p1_8.x63.A.n4 frontAnalog_v0p0p1_8.x63.A.n3 1.73501
R24270 frontAnalog_v0p0p1_8.x63.A.n1 frontAnalog_v0p0p1_8.x63.A.n4 0.99025
R24271 frontAnalog_v0p0p1_8.x63.A.n5 frontAnalog_v0p0p1_8.x63.A.n1 0.853186
R24272 frontAnalog_v0p0p1_8.x63.A frontAnalog_v0p0p1_8.x63.A.n0 0.349517
R24273 frontAnalog_v0p0p1_8.x63.A frontAnalog_v0p0p1_8.x63.A.n5 0.24425
R24274 frontAnalog_v0p0p1_2.RSfetsym_0.QN.n1 frontAnalog_v0p0p1_2.RSfetsym_0.QN.t5 117.511
R24275 frontAnalog_v0p0p1_2.RSfetsym_0.QN.n1 frontAnalog_v0p0p1_2.RSfetsym_0.QN.t6 110.698
R24276 frontAnalog_v0p0p1_2.RSfetsym_0.QN.n2 frontAnalog_v0p0p1_2.RSfetsym_0.QN.t2 19.1963
R24277 frontAnalog_v0p0p1_2.RSfetsym_0.QN.n3 frontAnalog_v0p0p1_2.RSfetsym_0.QN.t1 14.5206
R24278 frontAnalog_v0p0p1_2.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_2.RSfetsym_0.QN.t3 14.283
R24279 frontAnalog_v0p0p1_2.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_2.RSfetsym_0.QN.t4 14.283
R24280 frontAnalog_v0p0p1_2.RSfetsym_0.QN frontAnalog_v0p0p1_2.RSfetsym_0.QN.t0 9.14075
R24281 frontAnalog_v0p0p1_2.RSfetsym_0.QN.n2 frontAnalog_v0p0p1_2.RSfetsym_0.QN.n1 0.826818
R24282 frontAnalog_v0p0p1_2.RSfetsym_0.QN frontAnalog_v0p0p1_2.RSfetsym_0.QN.n0 0.74645
R24283 frontAnalog_v0p0p1_2.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_2.RSfetsym_0.QN.n3 0.249509
R24284 frontAnalog_v0p0p1_2.RSfetsym_0.QN.n3 frontAnalog_v0p0p1_2.RSfetsym_0.QN.n2 0.0968646
R24285 frontAnalog_v0p0p1_12.x65.A.n1 frontAnalog_v0p0p1_12.x65.A.t4 260.322
R24286 frontAnalog_v0p0p1_12.x65.A.n3 frontAnalog_v0p0p1_12.x65.A.t7 233.929
R24287 frontAnalog_v0p0p1_12.x65.A.n1 frontAnalog_v0p0p1_12.x65.A.t6 175.169
R24288 frontAnalog_v0p0p1_12.x65.A.n2 frontAnalog_v0p0p1_12.x65.A.t5 160.416
R24289 frontAnalog_v0p0p1_12.x65.A.n4 frontAnalog_v0p0p1_12.x65.A.t0 17.4109
R24290 frontAnalog_v0p0p1_12.x65.A.n4 frontAnalog_v0p0p1_12.x65.A.t1 10.2053
R24291 frontAnalog_v0p0p1_12.x65.A.n0 frontAnalog_v0p0p1_12.x65.A 2.78715
R24292 frontAnalog_v0p0p1_12.x65.A.n0 frontAnalog_v0p0p1_12.x65.A.n1 9.09103
R24293 frontAnalog_v0p0p1_12.x65.A.n6 frontAnalog_v0p0p1_12.x65.A.t2 7.94569
R24294 frontAnalog_v0p0p1_12.x65.A.n2 frontAnalog_v0p0p1_12.x65.A.t3 7.55846
R24295 frontAnalog_v0p0p1_12.x65.A.n5 frontAnalog_v0p0p1_12.x65.A.n3 1.4614
R24296 frontAnalog_v0p0p1_12.x65.A.n3 frontAnalog_v0p0p1_12.x65.A.n2 1.19626
R24297 frontAnalog_v0p0p1_12.x65.A.n6 frontAnalog_v0p0p1_12.x65.A.n5 0.836961
R24298 frontAnalog_v0p0p1_12.x65.A frontAnalog_v0p0p1_12.x65.A.n0 0.390342
R24299 frontAnalog_v0p0p1_12.x65.A.n5 frontAnalog_v0p0p1_12.x65.A.n4 0.154668
R24300 frontAnalog_v0p0p1_12.x65.A frontAnalog_v0p0p1_12.x65.A.n6 0.08175
R24301 frontAnalog_v0p0p1_6.x65.A.n1 frontAnalog_v0p0p1_6.x65.A.t6 260.322
R24302 frontAnalog_v0p0p1_6.x65.A.n4 frontAnalog_v0p0p1_6.x65.A.t5 233.929
R24303 frontAnalog_v0p0p1_6.x65.A.n1 frontAnalog_v0p0p1_6.x65.A.t7 175.169
R24304 frontAnalog_v0p0p1_6.x65.A.n3 frontAnalog_v0p0p1_6.x65.A.t4 160.416
R24305 frontAnalog_v0p0p1_6.x65.A.n2 frontAnalog_v0p0p1_6.x65.A.t2 17.4109
R24306 frontAnalog_v0p0p1_6.x65.A.n2 frontAnalog_v0p0p1_6.x65.A.t3 10.2053
R24307 frontAnalog_v0p0p1_6.x65.A.n0 frontAnalog_v0p0p1_6.x65.A 2.78715
R24308 frontAnalog_v0p0p1_6.x65.A.n0 frontAnalog_v0p0p1_6.x65.A.n1 9.09103
R24309 frontAnalog_v0p0p1_6.x65.A.n6 frontAnalog_v0p0p1_6.x65.A.t1 7.94569
R24310 frontAnalog_v0p0p1_6.x65.A.n3 frontAnalog_v0p0p1_6.x65.A.t0 7.55846
R24311 frontAnalog_v0p0p1_6.x65.A.n5 frontAnalog_v0p0p1_6.x65.A.n4 1.4614
R24312 frontAnalog_v0p0p1_6.x65.A.n4 frontAnalog_v0p0p1_6.x65.A.n3 1.19626
R24313 frontAnalog_v0p0p1_6.x65.A.n6 frontAnalog_v0p0p1_6.x65.A.n5 0.836961
R24314 frontAnalog_v0p0p1_6.x65.A frontAnalog_v0p0p1_6.x65.A.n0 0.390342
R24315 frontAnalog_v0p0p1_6.x65.A.n5 frontAnalog_v0p0p1_6.x65.A.n2 0.154668
R24316 frontAnalog_v0p0p1_6.x65.A frontAnalog_v0p0p1_6.x65.A.n6 0.08175
R24317 frontAnalog_v0p0p1_0.x65.A.n1 frontAnalog_v0p0p1_0.x65.A.t5 260.322
R24318 frontAnalog_v0p0p1_0.x65.A.n4 frontAnalog_v0p0p1_0.x65.A.t7 233.929
R24319 frontAnalog_v0p0p1_0.x65.A.n1 frontAnalog_v0p0p1_0.x65.A.t6 175.169
R24320 frontAnalog_v0p0p1_0.x65.A.n3 frontAnalog_v0p0p1_0.x65.A.t4 160.416
R24321 frontAnalog_v0p0p1_0.x65.A.n2 frontAnalog_v0p0p1_0.x65.A.t3 17.4109
R24322 frontAnalog_v0p0p1_0.x65.A.n2 frontAnalog_v0p0p1_0.x65.A.t2 10.2053
R24323 frontAnalog_v0p0p1_0.x65.A.n0 frontAnalog_v0p0p1_0.x65.A 2.78715
R24324 frontAnalog_v0p0p1_0.x65.A.n0 frontAnalog_v0p0p1_0.x65.A.n1 9.09103
R24325 frontAnalog_v0p0p1_0.x65.A.n6 frontAnalog_v0p0p1_0.x65.A.t1 7.94569
R24326 frontAnalog_v0p0p1_0.x65.A.n3 frontAnalog_v0p0p1_0.x65.A.t0 7.55846
R24327 frontAnalog_v0p0p1_0.x65.A.n5 frontAnalog_v0p0p1_0.x65.A.n4 1.4614
R24328 frontAnalog_v0p0p1_0.x65.A.n4 frontAnalog_v0p0p1_0.x65.A.n3 1.19626
R24329 frontAnalog_v0p0p1_0.x65.A.n6 frontAnalog_v0p0p1_0.x65.A.n5 0.836961
R24330 frontAnalog_v0p0p1_0.x65.A frontAnalog_v0p0p1_0.x65.A.n0 0.390342
R24331 frontAnalog_v0p0p1_0.x65.A.n5 frontAnalog_v0p0p1_0.x65.A.n2 0.154668
R24332 frontAnalog_v0p0p1_0.x65.A frontAnalog_v0p0p1_0.x65.A.n6 0.08175
R24333 frontAnalog_v0p0p1_0.x63.A.n2 frontAnalog_v0p0p1_0.x63.A.t5 260.322
R24334 frontAnalog_v0p0p1_0.x63.A.n4 frontAnalog_v0p0p1_0.x63.A.t4 233.888
R24335 frontAnalog_v0p0p1_0.x63.A.n2 frontAnalog_v0p0p1_0.x63.A.t6 175.169
R24336 frontAnalog_v0p0p1_0.x63.A.n3 frontAnalog_v0p0p1_0.x63.A.t7 159.725
R24337 frontAnalog_v0p0p1_0.x63.A.n1 frontAnalog_v0p0p1_0.x63.A.t2 17.4109
R24338 frontAnalog_v0p0p1_0.x63.A.n0 frontAnalog_v0p0p1_0.x63.A.n2 9.75129
R24339 frontAnalog_v0p0p1_0.x63.A.n1 frontAnalog_v0p0p1_0.x63.A.t3 9.6037
R24340 frontAnalog_v0p0p1_0.x63.A.n0 frontAnalog_v0p0p1_0.x63.A 2.33338
R24341 frontAnalog_v0p0p1_0.x63.A.n5 frontAnalog_v0p0p1_0.x63.A.t0 8.40929
R24342 frontAnalog_v0p0p1_0.x63.A.n3 frontAnalog_v0p0p1_0.x63.A.t1 8.06629
R24343 frontAnalog_v0p0p1_0.x63.A.n4 frontAnalog_v0p0p1_0.x63.A.n3 1.73501
R24344 frontAnalog_v0p0p1_0.x63.A.n1 frontAnalog_v0p0p1_0.x63.A.n4 0.99025
R24345 frontAnalog_v0p0p1_0.x63.A.n5 frontAnalog_v0p0p1_0.x63.A.n1 0.853186
R24346 frontAnalog_v0p0p1_0.x63.A frontAnalog_v0p0p1_0.x63.A.n0 0.349517
R24347 frontAnalog_v0p0p1_0.x63.A frontAnalog_v0p0p1_0.x63.A.n5 0.24425
C0 frontAnalog_v0p0p1_9.x65.A a_57123_n51159# 0.214f
C1 CLK VV15 0.618f
C2 w_55000_n25150# frontAnalog_v0p0p1_10.IB 0.0217f
C3 a_57123_n34959# frontAnalog_v0p0p1_7.x65.X 0.119f
C4 frontAnalog_v0p0p1_5.x63.A VDD 3.67f
C5 frontAnalog_v0p0p1_10.IB VV4 3.88f
C6 CLK VIN 5.84f
C7 a_77605_n40069# I13 0.16f
C8 16to4_PriorityEncoder_v0p0p1_0.x5.x19.C a_77605_n43295# 0.173f
C9 frontAnalog_v0p0p1_6.x63.A frontAnalog_v0p0p1_6.x65.A 3.16f
C10 frontAnalog_v0p0p1_13.x65.A a_57123_n67359# 0.214f
C11 w_55000_n30550# CLK 0.535f
C12 frontAnalog_v0p0p1_2.x65.X VDD 3.46f
C13 16to4_PriorityEncoder_v0p0p1_0.x5.x16.C I12 0.202f
C14 a_55268_n84936# CLK 0.235f
C15 a_57123_n78159# frontAnalog_v0p0p1_14.x65.X 0.119f
C16 16to4_PriorityEncoder_v0p0p1_0.x5.x22.A I15 0.0853f
C17 frontAnalog_v0p0p1_8.RSfetsym_0.QN a_59577_n46683# 0.418f
C18 a_59577_n73683# I2 0.29f
C19 frontAnalog_v0p0p1_2.x65.X frontAnalog_v0p0p1_2.x63.X 0.143f
C20 frontAnalog_v0p0p1_2.x63.A VIN 0.187f
C21 VDD VV3 1.84f
C22 w_55000_n2928# VDD 0.854f
C23 I15 I13 1.14f
C24 16to4_PriorityEncoder_v0p0p1_0.x3.x21.B a_78097_n53777# 0.186f
C25 m3_58396_n58350# CLK 0.189f
C26 a_78065_n49349# VDD 0.156f
C27 a_59578_n78570# I1 0.42f
C28 w_55000_n41350# VV9 0.751f
C29 frontAnalog_v0p0p1_7.x65.X a_59578_n35370# 0.436f
C30 w_55000_n84550# VV1 0.751f
C31 w_55000_n19128# a_53630_n20196# 0.359f
C32 frontAnalog_v0p0p1_2.RSfetsym_0.QN frontAnalog_v0p0p1_2.RSfetsym_0.x1.Y 0.17f
C33 w_55000_n57550# a_55268_n57936# 0.12f
C34 frontAnalog_v0p0p1_12.x63.A a_57123_n74279# 0.212f
C35 a_59577_n84483# VDD 0.0173f
C36 a_77605_n51335# VDD 0.435f
C37 16to4_PriorityEncoder_v0p0p1_0.x3.x4.A VDD 1.55f
C38 a_53630_n57996# a_55268_n57936# 0.015f
C39 16to4_PriorityEncoder_v0p0p1_0.x3.x19.D I0 0.122f
C40 frontAnalog_v0p0p1_2.x63.X VDD 3.13f
C41 frontAnalog_v0p0p1_14.x65.X a_59578_n78570# 0.436f
C42 a_53630_n52596# CLK 0.0136f
C43 frontAnalog_v0p0p1_10.x63.A CLK 1.8f
C44 frontAnalog_v0p0p1_10.x65.A VV6 0.253f
C45 frontAnalog_v0p0p1_4.x63.A frontAnalog_v0p0p1_4.x65.A 3.16f
C46 frontAnalog_v0p0p1_13.x65.A VV4 0.253f
C47 w_55000_n19750# frontAnalog_v0p0p1_4.x65.A 0.0988f
C48 16to4_PriorityEncoder_v0p0p1_0.x5.x16.C 16to4_PriorityEncoder_v0p0p1_0.x5.x15.X 0.0319f
C49 a_53630_n41796# VIN 0.265f
C50 frontAnalog_v0p0p1_13.x63.A frontAnalog_v0p0p1_13.x63.X 0.0301f
C51 w_55000_n13728# VIN 0.866f
C52 I9 I8 3.07f
C53 w_55000_n67728# frontAnalog_v0p0p1_10.IB 0.0216f
C54 a_59577_n35883# I9 0.29f
C55 16to4_PriorityEncoder_v0p0p1_0.x5.x19.D VDD 3.27f
C56 16to4_PriorityEncoder_v0p0p1_0.x5.x16.X a_77605_n43545# 0.102f
C57 16to4_PriorityEncoder_v0p0p1_0.x3.x19.D I4 0.206f
C58 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2 8.68f
C59 frontAnalog_v0p0p1_2.RSfetsym_0.x1.Y frontAnalog_v0p0p1_2.RSfetsym_0.x2.Y 0.0254f
C60 frontAnalog_v0p0p1_1.x63.A a_57123_n41879# 0.212f
C61 a_55268_n63336# VDD 0.565f
C62 a_82906_n51645# 16to4_PriorityEncoder_v0p0p1_0.x2.X 0.12f
C63 16to4_PriorityEncoder_v0p0p1_0.x3.x19.C 16to4_PriorityEncoder_v0p0p1_0.x3.x21.B 0.0127f
C64 frontAnalog_v0p0p1_12.x65.A frontAnalog_v0p0p1_12.x65.X 0.0236f
C65 VV1 VL 1.96f
C66 frontAnalog_v0p0p1_14.x63.X R1 0.0401f
C67 VIN S0 0.655f
C68 w_55000_n73128# CLK 0.57f
C69 frontAnalog_v0p0p1_9.x65.A VDD 3.44f
C70 frontAnalog_v0p0p1_14.RSfetsym_0.x1.Y I1 0.0436f
C71 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_7.x65.A 0.0352f
C72 frontAnalog_v0p0p1_7.x65.X frontAnalog_v0p0p1_7.RSfetsym_0.x1.Y 0.182f
C73 frontAnalog_v0p0p1_11.x63.A a_57123_n63479# 0.212f
C74 frontAnalog_v0p0p1_7.x63.X m3_58396_n36750# 0.134f
C75 w_55000_n41350# VDD 0.829f
C76 frontAnalog_v0p0p1_12.x63.A CLK 1.8f
C77 16to4_PriorityEncoder_v0p0p1_0.x3.x16.X VDD 0.505f
C78 a_55268_n84936# S0 0.461f
C79 a_53630_n47196# a_55268_n47136# 0.015f
C80 frontAnalog_v0p0p1_9.RSfetsym_0.QN VDD 2.55f
C81 a_77605_n51335# 16to4_PriorityEncoder_v0p0p1_0.x3.x16.X 0.0121f
C82 a_57123_n20279# CLK 0.0108f
C83 w_55000_n51528# VV7 0.798f
C84 frontAnalog_v0p0p1_10.IB VV11 3.87f
C85 frontAnalog_v0p0p1_14.x65.X frontAnalog_v0p0p1_14.RSfetsym_0.x1.Y 0.182f
C86 w_55000_n35950# VV10 0.751f
C87 a_53630_n3996# VV16 0.28f
C88 frontAnalog_v0p0p1_9.x63.X m3_58396_n52950# 0.134f
C89 m3_58396_n79950# VDD 1.25f
C90 a_55268_n3936# CLK 0.235f
C91 16to4_PriorityEncoder_v0p0p1_0.x3.x17.A a_78065_n49349# 0.2f
C92 frontAnalog_v0p0p1_4.RSfetsym_0.QN CLK 0.0457f
C93 frontAnalog_v0p0p1_8.x65.A frontAnalog_v0p0p1_8.x65.X 0.0236f
C94 w_55000_n67728# frontAnalog_v0p0p1_13.x65.A 0.658f
C95 16to4_PriorityEncoder_v0p0p1_0.x5.x19.C 16to4_PriorityEncoder_v0p0p1_0.x5.x21.B 0.0127f
C96 16to4_PriorityEncoder_v0p0p1_0.x3.x17.A VDD 1.34f
C97 a_77637_n49127# VDD 0.218f
C98 frontAnalog_v0p0p1_7.RSfetsym_0.x1.Y frontAnalog_v0p0p1_7.x63.X 0.883f
C99 a_53630_n79596# VIN 0.265f
C100 I13 I8 0.331f
C101 frontAnalog_v0p0p1_11.x65.A frontAnalog_v0p0p1_11.x65.X 0.0236f
C102 frontAnalog_v0p0p1_2.RSfetsym_0.QN frontAnalog_v0p0p1_2.RSfetsym_0.x2.Y 0.018f
C103 frontAnalog_v0p0p1_7.x65.A a_55268_n36336# 0.461f
C104 VIN VV8 3.41f
C105 a_77605_n53805# 16to4_PriorityEncoder_v0p0p1_0.x3.x20.X 0.0895f
C106 frontAnalog_v0p0p1_3.x65.A a_55268_n14736# 0.461f
C107 w_55000_n52150# VIN 0.737f
C108 frontAnalog_v0p0p1_2.x63.A a_55268_n3936# 1.24f
C109 a_59577_n3483# VDD 0.0172f
C110 16to4_PriorityEncoder_v0p0p1_0.x3.x16.C I0 0.12f
C111 a_57123_n72759# VDD 0.222f
C112 w_55000_n68350# frontAnalog_v0p0p1_13.x63.A 0.659f
C113 frontAnalog_v0p0p1_14.RSfetsym_0.x1.Y frontAnalog_v0p0p1_14.x63.X 0.883f
C114 frontAnalog_v0p0p1_14.RSfetsym_0.QN I1 2.02f
C115 16to4_PriorityEncoder_v0p0p1_0.x5.x19.C I12 0.405f
C116 a_53630_n25596# VDD 0.134f
C117 frontAnalog_v0p0p1_7.x65.X frontAnalog_v0p0p1_7.RSfetsym_0.QN 2.28f
C118 frontAnalog_v0p0p1_1.x65.A CLK 2.63f
C119 frontAnalog_v0p0p1_2.x63.X a_59577_n3483# 0.28f
C120 16to4_PriorityEncoder_v0p0p1_0.x3.x18.C 16to4_PriorityEncoder_v0p0p1_0.x3.x21.B 0.014f
C121 a_78649_n47567# VDD 0.235f
C122 16to4_PriorityEncoder_v0p0p1_0.x3.x19.D VDD 1.32f
C123 16to4_PriorityEncoder_v0p0p1_0.x3.x19.D 16to4_PriorityEncoder_v0p0p1_0.x3.x4.A 0.0516f
C124 16to4_PriorityEncoder_v0p0p1_0.x5.x16.C VDD 2.83f
C125 frontAnalog_v0p0p1_7.x63.X a_57123_n36479# 0.121f
C126 frontAnalog_v0p0p1_10.IB S1 0.0352f
C127 frontAnalog_v0p0p1_14.x65.X frontAnalog_v0p0p1_14.RSfetsym_0.QN 2.28f
C128 16to4_PriorityEncoder_v0p0p1_0.x3.x16.C I4 0.202f
C129 w_55000_n83928# VDD 0.854f
C130 frontAnalog_v0p0p1_1.x65.X I8 0.445f
C131 frontAnalog_v0p0p1_10.IB VV15 4.52f
C132 frontAnalog_v0p0p1_10.IB VIN 32.9f
C133 frontAnalog_v0p0p1_11.x63.A VV5 0.587f
C134 16to4_PriorityEncoder_v0p0p1_0.x3.x15.X VDD 0.26f
C135 frontAnalog_v0p0p1_3.x65.A VV14 0.253f
C136 a_77605_n51335# 16to4_PriorityEncoder_v0p0p1_0.x3.x15.X 0.0951f
C137 frontAnalog_v0p0p1_11.x65.X I4 0.446f
C138 a_59578_n46170# VDD 0.0209f
C139 VV10 VV9 2.78f
C140 CLK I12 0.0757f
C141 a_59578_n73170# VDD 0.0209f
C142 frontAnalog_v0p0p1_14.x63.X a_57123_n79679# 0.121f
C143 frontAnalog_v0p0p1_14.RSfetsym_0.x2.Y I1 0.198f
C144 16to4_PriorityEncoder_v0p0p1_0.x3.x17.A 16to4_PriorityEncoder_v0p0p1_0.x3.x16.X 0.0198f
C145 frontAnalog_v0p0p1_7.x65.X frontAnalog_v0p0p1_7.RSfetsym_0.x2.Y 0.526f
C146 frontAnalog_v0p0p1_5.x65.A VV12 0.253f
C147 frontAnalog_v0p0p1_7.RSfetsym_0.QN frontAnalog_v0p0p1_7.x63.X 0.378f
C148 w_55000_n30550# frontAnalog_v0p0p1_10.IB 0.0217f
C149 a_82906_n51645# 16to4_PriorityEncoder_v0p0p1_0.x3.A0 0.119f
C150 frontAnalog_v0p0p1_10.IB a_55268_n84936# 0.0848f
C151 frontAnalog_v0p0p1_4.x63.A VV13 0.587f
C152 w_55000_n19750# VV13 0.751f
C153 w_55000_n51528# a_55268_n52536# 0.149f
C154 w_55000_n52150# a_53630_n52596# 0.394f
C155 16to4_PriorityEncoder_v0p0p1_0.x5.x16.C 16to4_PriorityEncoder_v0p0p1_0.x5.x19.D 1.24f
C156 frontAnalog_v0p0p1_8.x65.A VIN 0.654f
C157 w_55000_n35950# CLK 0.535f
C158 frontAnalog_v0p0p1_11.x65.A CLK 2.63f
C159 frontAnalog_v0p0p1_14.RSfetsym_0.QN frontAnalog_v0p0p1_14.x63.X 0.378f
C160 frontAnalog_v0p0p1_14.x65.X frontAnalog_v0p0p1_14.RSfetsym_0.x2.Y 0.526f
C161 16to4_PriorityEncoder_v0p0p1_0.x5.x18.C 16to4_PriorityEncoder_v0p0p1_0.x5.x21.B 0.014f
C162 frontAnalog_v0p0p1_3.x65.A CLK 2.63f
C163 16to4_PriorityEncoder_v0p0p1_0.x1.A 16to4_PriorityEncoder_v0p0p1_0.x2.A 0.304f
C164 frontAnalog_v0p0p1_15.x65.X CLK 0.442f
C165 frontAnalog_v0p0p1_8.RSfetsym_0.x1.Y frontAnalog_v0p0p1_8.RSfetsym_0.x2.Y 0.0254f
C166 16to4_PriorityEncoder_v0p0p1_0.x3.x19.X 16to4_PriorityEncoder_v0p0p1_0.x3.x20.X 0.145f
C167 w_55000_n8328# VDD 0.854f
C168 frontAnalog_v0p0p1_11.x63.X I4 1.85f
C169 a_77605_n52819# 16to4_PriorityEncoder_v0p0p1_0.x3.x19.X 0.0873f
C170 a_55268_n36336# VIN 0.177f
C171 m3_58396_n69150# CLK 0.189f
C172 frontAnalog_v0p0p1_7.x63.X frontAnalog_v0p0p1_7.RSfetsym_0.x2.Y 0.0923f
C173 16to4_PriorityEncoder_v0p0p1_0.x5.x18.C I12 0.432f
C174 w_55000_n62328# w_55000_n62950# 0.327f
C175 a_59578_n40770# VDD 0.0209f
C176 CLK I0 0.0499f
C177 frontAnalog_v0p0p1_4.x63.A a_55268_n20136# 1.24f
C178 a_55268_n68736# VV4 0.215f
C179 w_55000_n35328# a_53630_n36396# 0.359f
C180 frontAnalog_v0p0p1_10.IB a_53630_n52596# 0.473f
C181 w_55000_n19750# a_55268_n20136# 0.12f
C182 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_10.x63.A 0.0926f
C183 m3_58396_n9750# VDD 1.24f
C184 frontAnalog_v0p0p1_13.x65.A VIN 0.655f
C185 16to4_PriorityEncoder_v0p0p1_0.x3.x22.A a_78065_n49349# 0.077f
C186 frontAnalog_v0p0p1_9.RSfetsym_0.x1.Y VDD 0.733f
C187 16to4_PriorityEncoder_v0p0p1_0.x3.x15.X 16to4_PriorityEncoder_v0p0p1_0.x3.x16.X 0.253f
C188 frontAnalog_v0p0p1_1.x63.A a_55268_n41736# 1.24f
C189 frontAnalog_v0p0p1_12.RSfetsym_0.x1.Y VDD 0.733f
C190 frontAnalog_v0p0p1_14.x63.X frontAnalog_v0p0p1_14.RSfetsym_0.x2.Y 0.0923f
C191 a_57123_n7959# frontAnalog_v0p0p1_0.x65.X 0.119f
C192 a_77605_n45765# I13 0.193f
C193 16to4_PriorityEncoder_v0p0p1_0.x3.x22.A VDD 3.23f
C194 a_57123_n51159# CLK 0.0108f
C195 16to4_PriorityEncoder_v0p0p1_0.x3.x22.A a_77605_n51335# 0.0116f
C196 VDD VV10 1.87f
C197 CLK I4 0.0837f
C198 a_53630_n74196# CLK 0.0136f
C199 a_77605_n43545# VDD 0.571f
C200 16to4_PriorityEncoder_v0p0p1_0.x3.x16.C VDD 0.834f
C201 frontAnalog_v0p0p1_12.x63.X m3_58396_n74550# 0.134f
C202 16to4_PriorityEncoder_v0p0p1_0.x3.x16.C a_77605_n51335# 0.0949f
C203 w_55000_n19128# VIN 0.868f
C204 frontAnalog_v0p0p1_6.x63.A VV11 0.587f
C205 w_55000_n73128# frontAnalog_v0p0p1_10.IB 0.0216f
C206 16to4_PriorityEncoder_v0p0p1_0.x5.A2 16to4_PriorityEncoder_v0p0p1_0.x3.A2 0.358f
C207 16to4_PriorityEncoder_v0p0p1_0.x3.x17.A 16to4_PriorityEncoder_v0p0p1_0.x3.x15.X 0.0789f
C208 frontAnalog_v0p0p1_11.x65.X VDD 3.46f
C209 m3_58396_n20550# I12 0.0416f
C210 w_55000_n24528# w_55000_n25150# 0.327f
C211 a_55268_n14736# VDD 0.565f
C212 CLK VV9 0.645f
C213 w_55000_n13728# frontAnalog_v0p0p1_3.x65.A 0.658f
C214 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_12.x63.A 0.0926f
C215 w_55000_n78528# CLK 0.57f
C216 a_57123_n47279# VDD 0.222f
C217 frontAnalog_v0p0p1_5.x65.A a_55268_n25536# 0.461f
C218 a_57123_n74279# VDD 0.222f
C219 16to4_PriorityEncoder_v0p0p1_0.x3.x19.C I0 0.12f
C220 frontAnalog_v0p0p1_0.x65.X a_59578_n8370# 0.436f
C221 frontAnalog_v0p0p1_7.RSfetsym_0.QN a_59577_n35883# 0.418f
C222 a_77639_n42341# I15 0.192f
C223 w_55000_n84550# R0 0.659f
C224 frontAnalog_v0p0p1_7.x63.A a_57123_n36479# 0.212f
C225 w_55000_n46750# VDD 0.829f
C226 frontAnalog_v0p0p1_3.x63.A a_57123_n14879# 0.212f
C227 frontAnalog_v0p0p1_15.x65.X S0 0.0362f
C228 frontAnalog_v0p0p1_10.IB a_55268_n3936# 0.0848f
C229 w_55000_n14350# frontAnalog_v0p0p1_3.x63.A 0.659f
C230 frontAnalog_v0p0p1_5.x63.A CLK 1.8f
C231 frontAnalog_v0p0p1_9.RSfetsym_0.QN frontAnalog_v0p0p1_9.RSfetsym_0.x1.Y 0.17f
C232 frontAnalog_v0p0p1_0.RSfetsym_0.QN I15 0.0512f
C233 frontAnalog_v0p0p1_12.RSfetsym_0.QN VDD 2.55f
C234 w_55000_n67728# a_55268_n68736# 0.149f
C235 w_55000_n68350# a_53630_n68796# 0.394f
C236 frontAnalog_v0p0p1_14.RSfetsym_0.QN a_59577_n79083# 0.418f
C237 16to4_PriorityEncoder_v0p0p1_0.x5.x19.C VDD 2.86f
C238 16to4_PriorityEncoder_v0p0p1_0.x3.x22.A 16to4_PriorityEncoder_v0p0p1_0.x3.x16.X 0.0732f
C239 16to4_PriorityEncoder_v0p0p1_0.x3.x19.C I4 0.405f
C240 frontAnalog_v0p0p1_11.x63.X VDD 3.13f
C241 frontAnalog_v0p0p1_2.x65.X CLK 0.512f
C242 16to4_PriorityEncoder_v0p0p1_0.x3.A2 16to4_PriorityEncoder_v0p0p1_0.x3.EO 0.162f
C243 VDD VV14 1.76f
C244 16to4_PriorityEncoder_v0p0p1_0.x3.x11.X a_78065_n49349# 0.202f
C245 frontAnalog_v0p0p1_2.x65.A a_57123_n2559# 0.214f
C246 frontAnalog_v0p0p1_9.x65.X a_59578_n51570# 0.436f
C247 a_59577_n62883# I4 0.29f
C248 16to4_PriorityEncoder_v0p0p1_0.x3.x16.C 16to4_PriorityEncoder_v0p0p1_0.x3.x16.X 0.07f
C249 16to4_PriorityEncoder_v0p0p1_0.x5.x16.X I11 0.0148f
C250 a_57123_n78159# S1 0.239f
C251 frontAnalog_v0p0p1_0.x65.A VDD 3.44f
C252 a_55268_n30936# VDD 0.565f
C253 w_55000_n29928# frontAnalog_v0p0p1_6.x65.A 0.658f
C254 16to4_PriorityEncoder_v0p0p1_0.x3.x11.X VDD 0.507f
C255 CLK VV3 0.645f
C256 w_55000_n2928# CLK 0.57f
C257 frontAnalog_v0p0p1_1.RSfetsym_0.QN I8 2.02f
C258 a_77605_n44527# I9 0.147f
C259 16to4_PriorityEncoder_v0p0p1_0.x5.x21.B I11 0.0112f
C260 frontAnalog_v0p0p1_6.x63.A VIN 0.187f
C261 frontAnalog_v0p0p1_7.x65.A frontAnalog_v0p0p1_7.x65.X 0.0236f
C262 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_1.x65.A 0.0352f
C263 16to4_PriorityEncoder_v0p0p1_0.x5.x17.A a_78349_n43045# 0.213f
C264 VV2 S1 0.253f
C265 a_78525_n53555# 16to4_PriorityEncoder_v0p0p1_0.x3.x20.X 0.0765f
C266 16to4_PriorityEncoder_v0p0p1_0.x3.x19.X 16to4_PriorityEncoder_v0p0p1_0.x3.x21.X 0.131f
C267 a_77605_n52567# I1 0.147f
C268 a_53630_n63396# VV5 0.28f
C269 16to4_PriorityEncoder_v0p0p1_0.x3.x22.A 16to4_PriorityEncoder_v0p0p1_0.x3.x17.A 1.27f
C270 frontAnalog_v0p0p1_3.x65.A frontAnalog_v0p0p1_3.x65.X 0.0236f
C271 w_55000_n57550# VIN 0.737f
C272 a_77637_n49127# 16to4_PriorityEncoder_v0p0p1_0.x3.x22.A 0.0288f
C273 16to4_PriorityEncoder_v0p0p1_0.x5.x19.C 16to4_PriorityEncoder_v0p0p1_0.x5.x19.D 0.996f
C274 frontAnalog_v0p0p1_8.RSfetsym_0.x2.Y VDD 0.926f
C275 VIN VV2 3.41f
C276 frontAnalog_v0p0p1_12.RSfetsym_0.x2.Y VDD 0.926f
C277 a_55268_n9336# VV15 0.215f
C278 a_53630_n57996# VIN 0.265f
C279 VDD CLK 91.3f
C280 w_55000_n30550# frontAnalog_v0p0p1_6.x63.A 0.659f
C281 frontAnalog_v0p0p1_0.x65.X frontAnalog_v0p0p1_0.RSfetsym_0.x1.Y 0.182f
C282 a_78097_n53777# VDD 0.219f
C283 a_55268_n9336# VIN 0.177f
C284 a_57123_n24159# VDD 0.222f
C285 a_53630_n41796# VV9 0.28f
C286 w_55000_n2928# frontAnalog_v0p0p1_2.x63.A 0.0792f
C287 I12 I11 5.01f
C288 a_53630_n20196# VV13 0.28f
C289 frontAnalog_v0p0p1_2.x63.X CLK 0.46f
C290 R1 S1 3.16f
C291 16to4_PriorityEncoder_v0p0p1_0.x1.A 16to4_PriorityEncoder_v0p0p1_0.x3.A1 0.426f
C292 w_55000_n51528# frontAnalog_v0p0p1_9.x63.A 0.0792f
C293 16to4_PriorityEncoder_v0p0p1_0.x3.x2.X I0 0.0265f
C294 VIN R1 0.19f
C295 16to4_PriorityEncoder_v0p0p1_0.x3.x18.C I0 0.119f
C296 I1 I3 1.73f
C297 I6 I0 0.364f
C298 a_55268_n25536# VV12 0.215f
C299 frontAnalog_v0p0p1_2.x63.A VDD 3.67f
C300 16to4_PriorityEncoder_v0p0p1_0.x3.x19.D 16to4_PriorityEncoder_v0p0p1_0.x3.x22.A 0.0292f
C301 a_53630_n47196# VIN 0.265f
C302 w_55000_n56928# frontAnalog_v0p0p1_10.x65.A 0.658f
C303 frontAnalog_v0p0p1_2.x63.A frontAnalog_v0p0p1_2.x63.X 0.0301f
C304 a_82906_n43855# 16to4_PriorityEncoder_v0p0p1_0.x3.A2 0.119f
C305 a_57123_n67359# frontAnalog_v0p0p1_13.x65.X 0.119f
C306 16to4_PriorityEncoder_v0p0p1_0.x3.x16.C 16to4_PriorityEncoder_v0p0p1_0.x3.x19.D 1.24f
C307 a_55268_n63336# CLK 0.235f
C308 frontAnalog_v0p0p1_0.RSfetsym_0.x1.Y frontAnalog_v0p0p1_0.x63.X 0.883f
C309 16to4_PriorityEncoder_v0p0p1_0.x3.x2.X I4 0.0262f
C310 w_55000_n35950# frontAnalog_v0p0p1_10.IB 0.0217f
C311 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_11.x65.A 0.0352f
C312 a_59578_n24570# VDD 0.0209f
C313 16to4_PriorityEncoder_v0p0p1_0.x5.x18.C VDD 2.22f
C314 16to4_PriorityEncoder_v0p0p1_0.x3.x22.A 16to4_PriorityEncoder_v0p0p1_0.x3.x15.X 0.209f
C315 16to4_PriorityEncoder_v0p0p1_0.x3.x18.C I4 0.432f
C316 a_53630_n20196# a_55268_n20136# 0.015f
C317 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_3.x65.A 0.0352f
C318 I7 I3 1.25f
C319 I4 I6 2.39f
C320 I2 I1 8.04f
C321 16to4_PriorityEncoder_v0p0p1_0.x5.x16.C a_77605_n43545# 0.0677f
C322 frontAnalog_v0p0p1_9.x65.A CLK 2.63f
C323 w_55000_n57550# frontAnalog_v0p0p1_10.x63.A 0.659f
C324 a_59578_n29970# I10 0.42f
C325 a_77605_n47345# 16to4_PriorityEncoder_v0p0p1_0.x3.x2.X 0.0313f
C326 16to4_PriorityEncoder_v0p0p1_0.x3.x19.C VDD 1.19f
C327 16to4_PriorityEncoder_v0p0p1_0.x5.x19.X a_78525_n45515# 0.193f
C328 16to4_PriorityEncoder_v0p0p1_0.x3.x16.C 16to4_PriorityEncoder_v0p0p1_0.x3.x15.X 0.0319f
C329 16to4_PriorityEncoder_v0p0p1_0.x3.x19.C a_77605_n51335# 0.173f
C330 w_55000_n41350# CLK 0.535f
C331 frontAnalog_v0p0p1_1.RSfetsym_0.x1.Y frontAnalog_v0p0p1_1.x63.X 0.883f
C332 frontAnalog_v0p0p1_0.x65.X frontAnalog_v0p0p1_0.RSfetsym_0.QN 2.28f
C333 frontAnalog_v0p0p1_9.RSfetsym_0.QN CLK 0.0457f
C334 frontAnalog_v0p0p1_4.x65.A a_57123_n18759# 0.214f
C335 a_59577_n62883# VDD 0.0172f
C336 I7 I2 0.468f
C337 frontAnalog_v0p0p1_8.RSfetsym_0.QN I7 2.02f
C338 a_53630_n41796# VDD 0.134f
C339 w_55000_n13728# VDD 0.854f
C340 a_55268_n68736# VIN 0.177f
C341 w_55000_n78528# a_53630_n79596# 0.359f
C342 16to4_PriorityEncoder_v0p0p1_0.x3.x11.X 16to4_PriorityEncoder_v0p0p1_0.x3.x17.A 0.125f
C343 16to4_PriorityEncoder_v0p0p1_0.x3.EI I3 1.97f
C344 16to4_PriorityEncoder_v0p0p1_0.x5.x18.C 16to4_PriorityEncoder_v0p0p1_0.x5.x19.D 0.491f
C345 a_77637_n49127# 16to4_PriorityEncoder_v0p0p1_0.x3.x11.X 0.109f
C346 VV9 VV8 3.01f
C347 frontAnalog_v0p0p1_1.x65.A a_57123_n40359# 0.214f
C348 frontAnalog_v0p0p1_13.x65.X a_59578_n67770# 0.436f
C349 m3_58396_n79950# CLK 0.189f
C350 frontAnalog_v0p0p1_0.x63.X a_57123_n9479# 0.121f
C351 16to4_PriorityEncoder_v0p0p1_0.x5.x4.A I11 0.0406f
C352 a_77637_n40777# 16to4_PriorityEncoder_v0p0p1_0.x5.x14.A 0.135f
C353 a_77637_n50057# VDD 0.234f
C354 w_55000_n35950# a_55268_n36336# 0.12f
C355 a_77605_n51585# VDD 0.432f
C356 VDD S0 3.8f
C357 16to4_PriorityEncoder_v0p0p1_0.x3.A1 a_78349_n51085# 0.151f
C358 a_77605_n53805# I5 0.193f
C359 m3_58396_n20550# VDD 1.25f
C360 16to4_PriorityEncoder_v0p0p1_0.x5.x22.A a_78525_n45515# 0.209f
C361 a_57123_n56559# frontAnalog_v0p0p1_10.x65.X 0.119f
C362 frontAnalog_v0p0p1_10.IB a_53630_n74196# 0.473f
C363 frontAnalog_v0p0p1_4.x65.A VIN 0.657f
C364 16to4_PriorityEncoder_v0p0p1_0.x5.x19.C 16to4_PriorityEncoder_v0p0p1_0.x5.x16.C 1.95f
C365 frontAnalog_v0p0p1_5.x63.A a_57123_n25679# 0.212f
C366 16to4_PriorityEncoder_v0p0p1_0.x3.EI I2 1.27f
C367 frontAnalog_v0p0p1_0.RSfetsym_0.QN frontAnalog_v0p0p1_0.x63.X 0.378f
C368 frontAnalog_v0p0p1_0.x65.X frontAnalog_v0p0p1_0.RSfetsym_0.x2.Y 0.526f
C369 frontAnalog_v0p0p1_5.RSfetsym_0.x1.Y VDD 0.733f
C370 a_59577_n41283# VDD 0.0172f
C371 frontAnalog_v0p0p1_12.RSfetsym_0.QN a_59578_n73170# 0.255f
C372 a_78525_n53555# 16to4_PriorityEncoder_v0p0p1_0.x3.x21.X 0.202f
C373 16to4_PriorityEncoder_v0p0p1_0.x5.x22.A a_78349_n43045# 0.17f
C374 a_57123_n72759# CLK 0.0108f
C375 frontAnalog_v0p0p1_6.RSfetsym_0.x1.Y I10 0.0436f
C376 a_53630_n25596# CLK 0.0136f
C377 frontAnalog_v0p0p1_10.IB VV9 3.87f
C378 w_55000_n24528# VIN 0.866f
C379 w_55000_n78528# frontAnalog_v0p0p1_10.IB 0.0216f
C380 frontAnalog_v0p0p1_4.x63.A frontAnalog_v0p0p1_4.x63.X 0.0301f
C381 w_55000_n40728# a_55268_n41736# 0.149f
C382 w_55000_n41350# a_53630_n41796# 0.394f
C383 16to4_PriorityEncoder_v0p0p1_0.x3.x2.X VDD 0.371f
C384 frontAnalog_v0p0p1_3.x65.X VDD 3.46f
C385 frontAnalog_v0p0p1_10.x65.X a_59578_n56970# 0.436f
C386 a_77605_n47345# 16to4_PriorityEncoder_v0p0p1_0.x3.x1.X 0.0991f
C387 16to4_PriorityEncoder_v0p0p1_0.x3.x4.A 16to4_PriorityEncoder_v0p0p1_0.x3.x2.X 0.125f
C388 w_55000_n83928# CLK 0.57f
C389 16to4_PriorityEncoder_v0p0p1_0.x2.A 16to4_PriorityEncoder_v0p0p1_0.x3.A1 1.21f
C390 16to4_PriorityEncoder_v0p0p1_0.x3.x18.C VDD 0.691f
C391 frontAnalog_v0p0p1_8.x65.X I8 0.0353f
C392 frontAnalog_v0p0p1_13.x65.X frontAnalog_v0p0p1_13.RSfetsym_0.x1.Y 0.182f
C393 VDD I6 4.09f
C394 a_53630_n79596# VDD 0.134f
C395 frontAnalog_v0p0p1_5.x65.A frontAnalog_v0p0p1_5.x65.X 0.0236f
C396 frontAnalog_v0p0p1_0.x63.X frontAnalog_v0p0p1_0.RSfetsym_0.x2.Y 0.0923f
C397 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_5.x63.A 0.0926f
C398 a_57123_n25679# VDD 0.222f
C399 VDD VV8 1.84f
C400 a_78159_n39549# 16to4_PriorityEncoder_v0p0p1_0.x5.x2.X 0.121f
C401 w_55000_n52150# VDD 0.829f
C402 frontAnalog_v0p0p1_12.x65.X frontAnalog_v0p0p1_12.x63.X 0.143f
C403 16to4_PriorityEncoder_v0p0p1_0.x3.x16.X a_77605_n51585# 0.102f
C404 16to4_PriorityEncoder_v0p0p1_0.x3.GS VDD 0.608f
C405 frontAnalog_v0p0p1_7.x63.A frontAnalog_v0p0p1_7.x65.A 3.16f
C406 a_57123_n45759# frontAnalog_v0p0p1_8.x65.X 0.119f
C407 frontAnalog_v0p0p1_9.x63.A frontAnalog_v0p0p1_9.x63.X 0.0301f
C408 w_55000_n8328# frontAnalog_v0p0p1_0.x65.A 0.658f
C409 frontAnalog_v0p0p1_5.RSfetsym_0.QN VDD 2.55f
C410 frontAnalog_v0p0p1_11.RSfetsym_0.QN a_59578_n62370# 0.255f
C411 frontAnalog_v0p0p1_10.IB VV3 3.87f
C412 w_55000_n2928# frontAnalog_v0p0p1_10.IB 0.0216f
C413 VDD I11 5.49f
C414 frontAnalog_v0p0p1_12.RSfetsym_0.QN frontAnalog_v0p0p1_12.RSfetsym_0.x1.Y 0.17f
C415 a_59578_n67770# I3 0.42f
C416 frontAnalog_v0p0p1_3.x63.X VDD 3.13f
C417 16to4_PriorityEncoder_v0p0p1_0.x3.x17.A a_77637_n50057# 0.14f
C418 frontAnalog_v0p0p1_6.RSfetsym_0.QN I10 2.02f
C419 frontAnalog_v0p0p1_11.RSfetsym_0.QN I5 0.0512f
C420 frontAnalog_v0p0p1_13.RSfetsym_0.x1.Y frontAnalog_v0p0p1_13.x63.X 0.883f
C421 w_55000_n3550# VV16 0.751f
C422 frontAnalog_v0p0p1_6.x65.X VDD 3.46f
C423 w_55000_n8950# frontAnalog_v0p0p1_0.x63.A 0.659f
C424 16to4_PriorityEncoder_v0p0p1_0.x3.x19.C 16to4_PriorityEncoder_v0p0p1_0.x3.x19.D 0.996f
C425 w_55000_n8328# CLK 0.57f
C426 frontAnalog_v0p0p1_10.IB VDD 19.5f
C427 w_55000_n3550# frontAnalog_v0p0p1_2.x65.A 0.0988f
C428 16to4_PriorityEncoder_v0p0p1_0.x5.x19.C a_77605_n43545# 0.176f
C429 frontAnalog_v0p0p1_9.x65.X frontAnalog_v0p0p1_9.x63.X 0.143f
C430 VDD OUT0 6.72f
C431 frontAnalog_v0p0p1_10.x65.X frontAnalog_v0p0p1_10.RSfetsym_0.x1.Y 0.182f
C432 frontAnalog_v0p0p1_3.RSfetsym_0.QN I14 0.0554f
C433 w_55000_n62950# VIN 0.737f
C434 w_55000_n52150# frontAnalog_v0p0p1_9.x65.A 0.0988f
C435 16to4_PriorityEncoder_v0p0p1_0.x3.x11.X 16to4_PriorityEncoder_v0p0p1_0.x3.x22.A 0.0936f
C436 frontAnalog_v0p0p1_13.x65.X frontAnalog_v0p0p1_13.RSfetsym_0.QN 2.28f
C437 frontAnalog_v0p0p1_0.RSfetsym_0.QN a_59577_n8883# 0.418f
C438 16to4_PriorityEncoder_v0p0p1_0.x5.x19.D I11 1.27f
C439 frontAnalog_v0p0p1_9.RSfetsym_0.QN I6 2.02f
C440 m3_58396_n9750# CLK 0.189f
C441 16to4_PriorityEncoder_v0p0p1_0.x5.A2 VDD 3.08f
C442 frontAnalog_v0p0p1_5.RSfetsym_0.x2.Y VDD 0.926f
C443 I10 I9 7.73f
C444 16to4_PriorityEncoder_v0p0p1_0.x5.x17.A I14 0.0474f
C445 frontAnalog_v0p0p1_11.x65.X frontAnalog_v0p0p1_11.x63.X 0.143f
C446 frontAnalog_v0p0p1_8.x65.A VDD 3.44f
C447 frontAnalog_v0p0p1_12.RSfetsym_0.x1.Y frontAnalog_v0p0p1_12.RSfetsym_0.x2.Y 0.0254f
C448 w_55000_n68350# VV4 0.751f
C449 16to4_PriorityEncoder_v0p0p1_0.x3.x1.X VDD 0.393f
C450 frontAnalog_v0p0p1_6.RSfetsym_0.x2.Y I10 0.196f
C451 a_55268_n14736# VV14 0.215f
C452 frontAnalog_v0p0p1_13.x63.X a_57123_n68879# 0.121f
C453 16to4_PriorityEncoder_v0p0p1_0.x3.x4.A 16to4_PriorityEncoder_v0p0p1_0.x3.x1.X 0.118f
C454 CLK VV10 0.645f
C455 frontAnalog_v0p0p1_1.x63.X a_57123_n41879# 0.121f
C456 frontAnalog_v0p0p1_6.x63.X VDD 3.13f
C457 frontAnalog_v0p0p1_1.RSfetsym_0.x1.Y frontAnalog_v0p0p1_1.RSfetsym_0.x2.Y 0.0254f
C458 frontAnalog_v0p0p1_10.IB a_55268_n63336# 0.0848f
C459 w_55000_n83928# S0 0.658f
C460 frontAnalog_v0p0p1_11.RSfetsym_0.QN frontAnalog_v0p0p1_11.RSfetsym_0.x1.Y 0.17f
C461 a_78159_n39549# 16to4_PriorityEncoder_v0p0p1_0.x5.x1.X 0.192f
C462 w_55000_n62328# frontAnalog_v0p0p1_11.x63.A 0.0792f
C463 16to4_PriorityEncoder_v0p0p1_0.x5.x17.A 16to4_PriorityEncoder_v0p0p1_0.x1.A 0.115f
C464 16to4_PriorityEncoder_v0p0p1_0.x3.x17.A I6 0.0474f
C465 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD 17f
C466 frontAnalog_v0p0p1_13.RSfetsym_0.x1.Y I3 0.0436f
C467 a_55268_n36336# VDD 0.565f
C468 16to4_PriorityEncoder_v0p0p1_0.x5.x4.A a_77605_n39305# 0.0112f
C469 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_9.x65.A 0.0352f
C470 frontAnalog_v0p0p1_10.RSfetsym_0.x1.Y frontAnalog_v0p0p1_10.x63.X 0.883f
C471 frontAnalog_v0p0p1_13.x65.X frontAnalog_v0p0p1_13.RSfetsym_0.x2.Y 0.526f
C472 frontAnalog_v0p0p1_13.RSfetsym_0.QN frontAnalog_v0p0p1_13.x63.X 0.378f
C473 frontAnalog_v0p0p1_10.x65.A a_55268_n57936# 0.461f
C474 VIN VV13 3.41f
C475 frontAnalog_v0p0p1_11.x65.X CLK 0.443f
C476 frontAnalog_v0p0p1_7.x63.A VIN 0.187f
C477 a_55268_n14736# CLK 0.235f
C478 w_55000_n41350# frontAnalog_v0p0p1_10.IB 0.0217f
C479 frontAnalog_v0p0p1_13.x65.A VDD 3.44f
C480 a_57123_n47279# CLK 0.0108f
C481 w_55000_n29928# VV11 0.798f
C482 a_57123_n74279# CLK 0.0108f
C483 16to4_PriorityEncoder_v0p0p1_0.x3.EO VDD 0.761f
C484 frontAnalog_v0p0p1_10.x65.X frontAnalog_v0p0p1_10.RSfetsym_0.QN 2.28f
C485 16to4_PriorityEncoder_v0p0p1_0.x3.x4.A 16to4_PriorityEncoder_v0p0p1_0.x3.EO 0.0491f
C486 16to4_PriorityEncoder_v0p0p1_0.x3.x19.D 16to4_PriorityEncoder_v0p0p1_0.x3.x2.X 0.014f
C487 w_55000_n46750# CLK 0.535f
C488 16to4_PriorityEncoder_v0p0p1_0.x3.x18.C 16to4_PriorityEncoder_v0p0p1_0.x3.x19.D 0.491f
C489 16to4_PriorityEncoder_v0p0p1_0.x3.x19.D I6 0.464f
C490 frontAnalog_v0p0p1_11.RSfetsym_0.x1.Y frontAnalog_v0p0p1_11.RSfetsym_0.x2.Y 0.0254f
C491 a_78159_n39549# 16to4_PriorityEncoder_v0p0p1_0.x5.EO 0.128f
C492 frontAnalog_v0p0p1_12.RSfetsym_0.QN frontAnalog_v0p0p1_12.RSfetsym_0.x2.Y 0.018f
C493 I14 I9 0.258f
C494 I13 I10 0.644f
C495 frontAnalog_v0p0p1_12.RSfetsym_0.QN CLK 0.0457f
C496 a_77605_n40069# I12 0.208f
C497 a_82906_n47995# VDD 0.179f
C498 a_59577_n14283# VDD 0.0172f
C499 frontAnalog_v0p0p1_10.x63.X a_57123_n58079# 0.121f
C500 a_57123_n40359# VDD 0.222f
C501 w_55000_n19128# VDD 0.854f
C502 w_55000_n79150# a_55268_n79536# 0.12f
C503 a_78649_n47567# 16to4_PriorityEncoder_v0p0p1_0.x3.GS 0.136f
C504 frontAnalog_v0p0p1_13.x63.X frontAnalog_v0p0p1_13.RSfetsym_0.x2.Y 0.0923f
C505 a_55268_n20136# VIN 0.177f
C506 frontAnalog_v0p0p1_11.x63.X CLK 0.46f
C507 frontAnalog_v0p0p1_1.x63.X frontAnalog_v0p0p1_1.RSfetsym_0.x2.Y 0.0923f
C508 16to4_PriorityEncoder_v0p0p1_0.x3.x19.C 16to4_PriorityEncoder_v0p0p1_0.x3.x16.C 1.95f
C509 CLK VV14 0.618f
C510 frontAnalog_v0p0p1_8.x63.X a_59577_n46683# 0.28f
C511 w_55000_n67728# w_55000_n68350# 0.327f
C512 VV6 VV5 4.54f
C513 w_55000_n46128# frontAnalog_v0p0p1_8.x63.A 0.0792f
C514 frontAnalog_v0p0p1_12.x63.X a_59577_n73683# 0.28f
C515 w_55000_n78528# VV2 0.798f
C516 frontAnalog_v0p0p1_0.x65.A CLK 2.63f
C517 a_55268_n30936# CLK 0.235f
C518 frontAnalog_v0p0p1_13.RSfetsym_0.QN I3 2.02f
C519 m3_58396_n31350# VDD 1.25f
C520 frontAnalog_v0p0p1_10.RSfetsym_0.QN frontAnalog_v0p0p1_10.x63.X 0.378f
C521 frontAnalog_v0p0p1_10.x65.X frontAnalog_v0p0p1_10.RSfetsym_0.x2.Y 0.526f
C522 I15 I12 0.786f
C523 frontAnalog_v0p0p1_10.IB a_53630_n25596# 0.473f
C524 16to4_PriorityEncoder_v0p0p1_0.x5.x16.C I11 0.132f
C525 w_55000_n78528# R1 0.0792f
C526 16to4_PriorityEncoder_v0p0p1_0.x22.A VDD 1.52f
C527 16to4_PriorityEncoder_v0p0p1_0.x3.x16.C a_77605_n51585# 0.0677f
C528 frontAnalog_v0p0p1_8.x65.X frontAnalog_v0p0p1_8.RSfetsym_0.QN 2.28f
C529 w_55000_n13728# a_55268_n14736# 0.149f
C530 w_55000_n14350# a_53630_n14796# 0.394f
C531 a_57123_n24159# CLK 0.0108f
C532 a_82906_n43855# VDD 0.181f
C533 16to4_PriorityEncoder_v0p0p1_0.x1.A 16to4_PriorityEncoder_v0p0p1_0.x28.A 0.0126f
C534 16to4_PriorityEncoder_v0p0p1_0.x5.EO 16to4_PriorityEncoder_v0p0p1_0.x3.EI 0.644f
C535 a_59577_n30483# VDD 0.0172f
C536 16to4_PriorityEncoder_v0p0p1_0.x5.x18.C 16to4_PriorityEncoder_v0p0p1_0.x5.x19.C 2.6f
C537 w_55000_n29928# VIN 0.866f
C538 w_55000_n83928# frontAnalog_v0p0p1_10.IB 0.0216f
C539 a_77605_n39305# VDD 0.149f
C540 a_53630_n84996# VIN 0.265f
C541 frontAnalog_v0p0p1_11.RSfetsym_0.QN frontAnalog_v0p0p1_11.RSfetsym_0.x2.Y 0.018f
C542 16to4_PriorityEncoder_v0p0p1_0.x5.x22.A I14 0.0536f
C543 a_77605_n44779# 16to4_PriorityEncoder_v0p0p1_0.x5.x19.X 0.0873f
C544 frontAnalog_v0p0p1_13.RSfetsym_0.x2.Y I3 0.198f
C545 w_55000_n29928# w_55000_n30550# 0.327f
C546 frontAnalog_v0p0p1_10.x63.X frontAnalog_v0p0p1_10.RSfetsym_0.x2.Y 0.0923f
C547 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1 8.67f
C548 I14 I13 10.5f
C549 VV3 VV2 4.95f
C550 frontAnalog_v0p0p1_2.x63.A CLK 1.8f
C551 frontAnalog_v0p0p1_13.RSfetsym_0.QN a_59577_n68283# 0.418f
C552 a_57123_n78159# VDD 0.22f
C553 a_53630_n84996# a_55268_n84936# 0.015f
C554 frontAnalog_v0p0p1_9.RSfetsym_0.x1.Y I6 0.0436f
C555 frontAnalog_v0p0p1_15.RSfetsym_0.QN I1 0.0512f
C556 frontAnalog_v0p0p1_6.x63.A VDD 3.67f
C557 frontAnalog_v0p0p1_11.x63.X a_59577_n62883# 0.28f
C558 16to4_PriorityEncoder_v0p0p1_0.x5.x22.A 16to4_PriorityEncoder_v0p0p1_0.x1.A 0.492f
C559 w_55000_n57550# VDD 0.829f
C560 16to4_PriorityEncoder_v0p0p1_0.x3.x22.A I6 0.0536f
C561 VDD VV2 1.93f
C562 a_53630_n57996# VDD 0.134f
C563 w_55000_n13728# VV14 0.798f
C564 a_55268_n9336# VDD 0.565f
C565 a_77605_n48109# I5 0.16f
C566 16to4_PriorityEncoder_v0p0p1_0.x3.EI 16to4_PriorityEncoder_v0p0p1_0.x3.x20.X 0.208f
C567 a_77605_n52567# 16to4_PriorityEncoder_v0p0p1_0.x3.x21.B 0.116f
C568 a_77637_n48817# 16to4_PriorityEncoder_v0p0p1_0.x3.x14.A 0.135f
C569 16to4_PriorityEncoder_v0p0p1_0.x3.x16.C I6 0.491f
C570 16to4_PriorityEncoder_v0p0p1_0.x3.EI a_77605_n52819# 0.175f
C571 w_55000_n8328# frontAnalog_v0p0p1_10.IB 0.0216f
C572 VDD R1 4f
C573 a_78649_n47567# 16to4_PriorityEncoder_v0p0p1_0.x3.EO 0.135f
C574 frontAnalog_v0p0p1_8.x63.A frontAnalog_v0p0p1_8.x63.X 0.0301f
C575 a_59578_n78570# VDD 0.0209f
C576 a_53630_n41796# CLK 0.0136f
C577 w_55000_n13728# CLK 0.57f
C578 a_53630_n47196# VDD 0.134f
C579 w_55000_n62328# a_53630_n63396# 0.359f
C580 16to4_PriorityEncoder_v0p0p1_0.x21.A VDD 0.539f
C581 16to4_PriorityEncoder_v0p0p1_0.x3.x21.B I3 0.0112f
C582 frontAnalog_v0p0p1_10.RSfetsym_0.QN a_59577_n57483# 0.418f
C583 a_77605_n43545# I11 0.162f
C584 w_55000_n68350# VIN 0.737f
C585 16to4_PriorityEncoder_v0p0p1_0.x3.x19.X a_78525_n53555# 0.193f
C586 16to4_PriorityEncoder_v0p0p1_0.x1.A 16to4_PriorityEncoder_v0p0p1_0.x1.X 0.0412f
C587 16to4_PriorityEncoder_v0p0p1_0.x5.x14.A a_78065_n41309# 0.197f
C588 frontAnalog_v0p0p1_10.x63.A a_57123_n58079# 0.212f
C589 CLK S0 2.64f
C590 frontAnalog_v0p0p1_10.IB VV10 3.87f
C591 m3_58396_n20550# CLK 0.189f
C592 w_55000_n46750# VV8 0.751f
C593 a_77637_n42017# I14 0.186f
C594 I12 I8 0.558f
C595 w_55000_n62950# frontAnalog_v0p0p1_11.x65.A 0.0988f
C596 frontAnalog_v0p0p1_2.x65.X I15 0.445f
C597 a_55268_n68736# VDD 0.565f
C598 frontAnalog_v0p0p1_10.IB a_55268_n14736# 0.0848f
C599 w_55000_n24528# frontAnalog_v0p0p1_5.x63.A 0.0792f
C600 a_53630_n3996# VIN 0.265f
C601 frontAnalog_v0p0p1_7.x65.X VDD 3.46f
C602 w_55000_n35328# frontAnalog_v0p0p1_7.x65.A 0.658f
C603 a_77605_n40069# VDD 0.156f
C604 16to4_PriorityEncoder_v0p0p1_0.x5.x19.X 16to4_PriorityEncoder_v0p0p1_0.x2.A 0.0122f
C605 frontAnalog_v0p0p1_10.x65.A frontAnalog_v0p0p1_10.x65.X 0.0236f
C606 frontAnalog_v0p0p1_14.RSfetsym_0.x1.Y VDD 0.733f
C607 16to4_PriorityEncoder_v0p0p1_0.x5.x19.C I11 0.921f
C608 frontAnalog_v0p0p1_3.x65.X CLK 0.443f
C609 w_55000_n46750# frontAnalog_v0p0p1_10.IB 0.0217f
C610 a_55268_n36336# VV10 0.215f
C611 a_57123_n18759# frontAnalog_v0p0p1_4.x65.X 0.119f
C612 CLK I6 0.0837f
C613 a_53630_n79596# CLK 0.0136f
C614 frontAnalog_v0p0p1_4.x65.A VDD 3.44f
C615 w_55000_n35950# frontAnalog_v0p0p1_7.x63.A 0.659f
C616 a_57123_n25679# CLK 0.0108f
C617 CLK VV8 0.645f
C618 16to4_PriorityEncoder_v0p0p1_0.x3.x19.C a_77605_n51585# 0.176f
C619 frontAnalog_v0p0p1_9.x63.A a_57123_n52679# 0.212f
C620 VDD I15 8.2f
C621 w_55000_n52150# CLK 0.535f
C622 frontAnalog_v0p0p1_2.x63.X I15 1.78f
C623 w_55000_n46750# frontAnalog_v0p0p1_8.x65.A 0.0988f
C624 frontAnalog_v0p0p1_10.IB VV14 3.88f
C625 frontAnalog_v0p0p1_7.x63.X VDD 3.13f
C626 VIN VV7 3.42f
C627 16to4_PriorityEncoder_v0p0p1_0.x5.x22.A 16to4_PriorityEncoder_v0p0p1_0.x2.A 0.132f
C628 16to4_PriorityEncoder_v0p0p1_0.x2.X VDD 0.351f
C629 w_55000_n24528# VDD 0.854f
C630 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_0.x65.A 0.0352f
C631 frontAnalog_v0p0p1_10.IB a_55268_n30936# 0.0848f
C632 frontAnalog_v0p0p1_5.RSfetsym_0.QN CLK 0.0457f
C633 a_57123_n79679# VDD 0.221f
C634 CLK I11 0.0837f
C635 w_55000_n56928# VV6 0.798f
C636 frontAnalog_v0p0p1_1.x63.X I9 0.015f
C637 frontAnalog_v0p0p1_3.x63.X CLK 0.46f
C638 frontAnalog_v0p0p1_1.x63.A VIN 0.187f
C639 frontAnalog_v0p0p1_4.x65.X a_59578_n19170# 0.436f
C640 16to4_PriorityEncoder_v0p0p1_0.x5.x19.D I15 0.244f
C641 frontAnalog_v0p0p1_6.x65.X CLK 0.443f
C642 a_77605_n45765# 16to4_PriorityEncoder_v0p0p1_0.x5.x20.X 0.0895f
C643 m3_58396_n42150# VDD 1.25f
C644 frontAnalog_v0p0p1_10.IB CLK 0.873f
C645 16to4_PriorityEncoder_v0p0p1_0.x3.EI 16to4_PriorityEncoder_v0p0p1_0.x1.A 0.534f
C646 16to4_PriorityEncoder_v0p0p1_0.x5.x14.A 16to4_PriorityEncoder_v0p0p1_0.x5.x17.A 0.105f
C647 frontAnalog_v0p0p1_14.RSfetsym_0.QN VDD 2.55f
C648 a_59578_n8370# I14 0.42f
C649 16to4_PriorityEncoder_v0p0p1_0.x3.x18.C 16to4_PriorityEncoder_v0p0p1_0.x3.x19.C 2.6f
C650 16to4_PriorityEncoder_v0p0p1_0.x3.x19.C I6 0.304f
C651 frontAnalog_v0p0p1_2.x65.A VV16 0.252f
C652 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3 7.92f
C653 frontAnalog_v0p0p1_5.RSfetsym_0.QN a_59578_n24570# 0.255f
C654 w_55000_n35328# VIN 0.866f
C655 16to4_PriorityEncoder_v0p0p1_0.x2.A a_82906_n51645# 0.207f
C656 frontAnalog_v0p0p1_8.x65.A CLK 2.63f
C657 VIN VV1 2.01f
C658 frontAnalog_v0p0p1_2.x63.A frontAnalog_v0p0p1_10.IB 0.0784f
C659 I13 I5 0.0641f
C660 a_78649_n39527# VDD 0.414f
C661 a_59578_n24570# I11 0.42f
C662 16to4_PriorityEncoder_v0p0p1_0.x5.x18.C I11 0.251f
C663 frontAnalog_v0p0p1_1.x65.X frontAnalog_v0p0p1_1.RSfetsym_0.x1.Y 0.182f
C664 a_53630_n52596# VV7 0.28f
C665 frontAnalog_v0p0p1_6.x63.X CLK 0.46f
C666 a_77637_n50057# I6 0.186f
C667 a_55268_n84936# VV1 0.214f
C668 frontAnalog_v0p0p1_14.RSfetsym_0.x2.Y VDD 0.926f
C669 frontAnalog_v0p0p1_11.x63.A VIN 0.187f
C670 a_55268_n36336# CLK 0.235f
C671 w_55000_n8328# a_55268_n9336# 0.149f
C672 w_55000_n8950# a_53630_n9396# 0.394f
C673 frontAnalog_v0p0p1_3.x63.A VIN 0.19f
C674 frontAnalog_v0p0p1_13.x63.X m3_58396_n69150# 0.134f
C675 frontAnalog_v0p0p1_10.x65.A VIN 0.655f
C676 16to4_PriorityEncoder_v0p0p1_0.x3.EI 16to4_PriorityEncoder_v0p0p1_0.x3.x14.A 0.0111f
C677 frontAnalog_v0p0p1_4.x65.X frontAnalog_v0p0p1_4.RSfetsym_0.x1.Y 0.182f
C678 w_55000_n62950# VDD 0.829f
C679 frontAnalog_v0p0p1_9.x65.X frontAnalog_v0p0p1_9.RSfetsym_0.x2.Y 0.526f
C680 a_53630_n3996# a_55268_n3936# 0.015f
C681 a_57123_n56559# VDD 0.222f
C682 frontAnalog_v0p0p1_13.x65.A CLK 2.63f
C683 frontAnalog_v0p0p1_0.x65.X VDD 3.46f
C684 frontAnalog_v0p0p1_5.x65.X frontAnalog_v0p0p1_5.x63.X 0.143f
C685 frontAnalog_v0p0p1_0.RSfetsym_0.x1.Y I14 0.0432f
C686 a_59577_n3483# I15 0.29f
C687 a_55268_n52536# VIN 0.177f
C688 VDD I8 5.2f
C689 frontAnalog_v0p0p1_10.IB a_53630_n41796# 0.473f
C690 w_55000_n13728# frontAnalog_v0p0p1_10.IB 0.0216f
C691 a_59577_n35883# VDD 0.0172f
C692 a_77639_n50381# I7 0.192f
C693 frontAnalog_v0p0p1_3.RSfetsym_0.QN a_59578_n13770# 0.255f
C694 frontAnalog_v0p0p1_5.RSfetsym_0.QN frontAnalog_v0p0p1_5.RSfetsym_0.x1.Y 0.17f
C695 16to4_PriorityEncoder_v0p0p1_0.x3.x2.X I6 0.0177f
C696 w_55000_n19128# CLK 0.57f
C697 frontAnalog_v0p0p1_5.RSfetsym_0.x1.Y I11 0.0436f
C698 a_57123_n40359# CLK 0.0108f
C699 frontAnalog_v0p0p1_10.IB S0 0.0352f
C700 a_57123_n45759# VDD 0.222f
C701 frontAnalog_v0p0p1_4.RSfetsym_0.x1.Y frontAnalog_v0p0p1_4.x63.X 0.883f
C702 16to4_PriorityEncoder_v0p0p1_0.x3.x18.C I6 0.3f
C703 frontAnalog_v0p0p1_1.x65.X frontAnalog_v0p0p1_1.x63.X 0.143f
C704 w_55000_n62950# a_55268_n63336# 0.12f
C705 w_55000_n24528# a_53630_n25596# 0.359f
C706 16to4_PriorityEncoder_v0p0p1_0.x5.x16.C I15 0.26f
C707 16to4_PriorityEncoder_v0p0p1_0.x3.A0 VDD 0.829f
C708 frontAnalog_v0p0p1_12.x65.A VIN 0.655f
C709 VDD VV13 1.84f
C710 a_59578_n56970# VDD 0.0209f
C711 frontAnalog_v0p0p1_7.x63.A VDD 3.67f
C712 w_55000_n73750# VIN 0.737f
C713 m3_58396_n69150# I3 0.0416f
C714 frontAnalog_v0p0p1_0.x63.X VDD 3.13f
C715 16to4_PriorityEncoder_v0p0p1_0.x3.EI a_77639_n50381# 0.088f
C716 16to4_PriorityEncoder_v0p0p1_0.x5.x19.D I8 0.122f
C717 frontAnalog_v0p0p1_10.x63.A frontAnalog_v0p0p1_10.x65.A 3.16f
C718 I3 I0 0.677f
C719 m3_58396_n31350# CLK 0.189f
C720 I5 I1 0.378f
C721 frontAnalog_v0p0p1_4.x65.X frontAnalog_v0p0p1_4.RSfetsym_0.QN 2.28f
C722 w_55000_n25150# frontAnalog_v0p0p1_5.x65.A 0.0988f
C723 frontAnalog_v0p0p1_8.RSfetsym_0.QN frontAnalog_v0p0p1_8.RSfetsym_0.x1.Y 0.17f
C724 frontAnalog_v0p0p1_3.x65.X frontAnalog_v0p0p1_3.x63.X 0.143f
C725 16to4_PriorityEncoder_v0p0p1_0.x5.x17.A a_78065_n41309# 0.2f
C726 frontAnalog_v0p0p1_5.RSfetsym_0.x1.Y frontAnalog_v0p0p1_5.RSfetsym_0.x2.Y 0.0254f
C727 16to4_PriorityEncoder_v0p0p1_0.x5.x14.A 16to4_PriorityEncoder_v0p0p1_0.x5.x22.A 0.0179f
C728 16to4_PriorityEncoder_v0p0p1_0.x3.EI 16to4_PriorityEncoder_v0p0p1_0.x2.A 0.645f
C729 frontAnalog_v0p0p1_0.RSfetsym_0.QN I14 2.02f
C730 a_53630_n52596# a_55268_n52536# 0.015f
C731 frontAnalog_v0p0p1_4.x63.X a_57123_n20279# 0.121f
C732 I2 I0 2.46f
C733 I4 I3 5.52f
C734 frontAnalog_v0p0p1_13.x65.X VDD 3.46f
C735 a_55268_n20136# VDD 0.565f
C736 I7 I5 1.12f
C737 frontAnalog_v0p0p1_6.x63.A a_55268_n30936# 1.24f
C738 frontAnalog_v0p0p1_10.IB a_53630_n79596# 0.473f
C739 frontAnalog_v0p0p1_3.RSfetsym_0.QN frontAnalog_v0p0p1_3.RSfetsym_0.x1.Y 0.17f
C740 m3_58396_n15150# I13 0.0416f
C741 frontAnalog_v0p0p1_10.IB VV8 3.87f
C742 a_77605_n47345# I3 0.0597f
C743 frontAnalog_v0p0p1_1.RSfetsym_0.x2.Y I9 0.0165f
C744 w_55000_n46750# a_53630_n47196# 0.394f
C745 w_55000_n46128# a_55268_n47136# 0.149f
C746 w_55000_n52150# frontAnalog_v0p0p1_10.IB 0.0217f
C747 frontAnalog_v0p0p1_5.RSfetsym_0.QN I11 2.02f
C748 frontAnalog_v0p0p1_1.x63.A frontAnalog_v0p0p1_1.x65.A 3.16f
C749 frontAnalog_v0p0p1_5.x63.X m3_58396_n25950# 0.134f
C750 frontAnalog_v0p0p1_4.RSfetsym_0.QN frontAnalog_v0p0p1_4.x63.X 0.378f
C751 frontAnalog_v0p0p1_0.x65.A a_55268_n9336# 0.461f
C752 frontAnalog_v0p0p1_4.x65.X frontAnalog_v0p0p1_4.RSfetsym_0.x2.Y 0.526f
C753 16to4_PriorityEncoder_v0p0p1_0.x29.A 16to4_PriorityEncoder_v0p0p1_0.x29.Y 1.51f
C754 a_57123_n78159# CLK 0.0108f
C755 I2 I4 0.848f
C756 a_77605_n44527# 16to4_PriorityEncoder_v0p0p1_0.x5.x21.B 0.116f
C757 frontAnalog_v0p0p1_6.x63.A CLK 1.8f
C758 frontAnalog_v0p0p1_10.RSfetsym_0.x1.Y VDD 0.733f
C759 16to4_PriorityEncoder_v0p0p1_0.x3.x1.X 16to4_PriorityEncoder_v0p0p1_0.x3.x2.X 0.129f
C760 frontAnalog_v0p0p1_0.RSfetsym_0.x2.Y I14 0.195f
C761 w_55000_n57550# CLK 0.535f
C762 16to4_PriorityEncoder_v0p0p1_0.x3.EI I5 3.69f
C763 frontAnalog_v0p0p1_8.x65.A VV8 0.253f
C764 CLK VV2 0.648f
C765 VDD OUT2 6.68f
C766 a_53630_n57996# CLK 0.0136f
C767 a_77605_n47345# I2 0.216f
C768 frontAnalog_v0p0p1_13.x63.X VDD 3.13f
C769 frontAnalog_v0p0p1_6.RSfetsym_0.QN a_59578_n29970# 0.255f
C770 a_55268_n9336# CLK 0.235f
C771 frontAnalog_v0p0p1_4.x65.X I12 0.446f
C772 frontAnalog_v0p0p1_3.RSfetsym_0.x1.Y frontAnalog_v0p0p1_3.RSfetsym_0.x2.Y 0.0254f
C773 w_55000_n29928# VDD 0.854f
C774 16to4_PriorityEncoder_v0p0p1_0.x3.x21.B 16to4_PriorityEncoder_v0p0p1_0.x3.x20.X 0.0561f
C775 a_53630_n84996# VDD 0.134f
C776 frontAnalog_v0p0p1_5.RSfetsym_0.QN frontAnalog_v0p0p1_5.RSfetsym_0.x2.Y 0.018f
C777 16to4_PriorityEncoder_v0p0p1_0.x5.x2.X I12 0.0262f
C778 w_55000_n73128# frontAnalog_v0p0p1_12.x65.A 0.658f
C779 16to4_PriorityEncoder_v0p0p1_0.x3.x21.B a_77605_n52819# 0.0141f
C780 frontAnalog_v0p0p1_5.RSfetsym_0.x2.Y I11 0.198f
C781 CLK R1 1.82f
C782 a_77605_n45765# VDD 0.552f
C783 w_55000_n73128# w_55000_n73750# 0.327f
C784 16to4_PriorityEncoder_v0p0p1_0.x3.EI a_77605_n53805# 0.343f
C785 frontAnalog_v0p0p1_4.x63.X frontAnalog_v0p0p1_4.RSfetsym_0.x2.Y 0.0923f
C786 a_55268_n57936# VV6 0.215f
C787 frontAnalog_v0p0p1_1.RSfetsym_0.QN frontAnalog_v0p0p1_1.RSfetsym_0.x1.Y 0.17f
C788 a_77605_n52567# VDD 0.432f
C789 frontAnalog_v0p0p1_8.x63.X I7 1.85f
C790 w_55000_n25150# VV12 0.751f
C791 a_78525_n45515# 16to4_PriorityEncoder_v0p0p1_0.x5.x20.X 0.0765f
C792 m3_58396_n52950# VDD 1.25f
C793 a_57123_n58079# VDD 0.222f
C794 16to4_PriorityEncoder_v0p0p1_0.x3.x2.X 16to4_PriorityEncoder_v0p0p1_0.x3.EO 0.0749f
C795 frontAnalog_v0p0p1_12.x63.A frontAnalog_v0p0p1_12.x65.A 3.16f
C796 a_53630_n47196# CLK 0.0136f
C797 frontAnalog_v0p0p1_5.x63.X a_59577_n25083# 0.28f
C798 a_59577_n8883# VDD 0.0172f
C799 a_53630_n63396# VIN 0.265f
C800 16to4_PriorityEncoder_v0p0p1_0.x5.x14.A 16to4_PriorityEncoder_v0p0p1_0.x5.x11.X 0.0721f
C801 16to4_PriorityEncoder_v0p0p1_0.x5.x16.C I8 0.12f
C802 w_55000_n73750# frontAnalog_v0p0p1_12.x63.A 0.659f
C803 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_8.x65.A 0.0352f
C804 frontAnalog_v0p0p1_6.x65.X frontAnalog_v0p0p1_6.x63.X 0.143f
C805 frontAnalog_v0p0p1_4.x63.X I12 1.85f
C806 a_78349_n43045# 16to4_PriorityEncoder_v0p0p1_0.x5.x16.X 0.0673f
C807 16to4_PriorityEncoder_v0p0p1_0.x3.EO 16to4_PriorityEncoder_v0p0p1_0.x3.GS 0.9f
C808 a_59578_n13770# I13 0.42f
C809 frontAnalog_v0p0p1_10.RSfetsym_0.QN VDD 2.55f
C810 16to4_PriorityEncoder_v0p0p1_0.x5.x19.D a_77605_n45765# 0.0838f
C811 VDD I3 3.69f
C812 w_55000_n40728# VIN 0.866f
C813 16to4_PriorityEncoder_v0p0p1_0.x3.x4.A I3 0.0406f
C814 frontAnalog_v0p0p1_10.IB a_55268_n36336# 0.0848f
C815 frontAnalog_v0p0p1_6.RSfetsym_0.QN frontAnalog_v0p0p1_6.RSfetsym_0.x1.Y 0.17f
C816 frontAnalog_v0p0p1_9.x63.A VIN 0.187f
C817 16to4_PriorityEncoder_v0p0p1_0.x5.x19.C I15 0.239f
C818 w_55000_n35328# w_55000_n35950# 0.327f
C819 frontAnalog_v0p0p1_3.RSfetsym_0.QN frontAnalog_v0p0p1_3.RSfetsym_0.x2.Y 0.018f
C820 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0 8.68f
C821 16to4_PriorityEncoder_v0p0p1_0.x5.x22.A a_78065_n41309# 0.077f
C822 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD 11.4f
C823 a_55268_n68736# CLK 0.235f
C824 a_77605_n43295# I10 0.167f
C825 16to4_PriorityEncoder_v0p0p1_0.x36.A 16to4_PriorityEncoder_v0p0p1_0.x36.Y 1.51f
C826 a_57123_n83559# frontAnalog_v0p0p1_15.x65.X 0.119f
C827 frontAnalog_v0p0p1_7.x65.X CLK 0.443f
C828 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_13.x65.A 0.0352f
C829 VDD I2 3.99f
C830 frontAnalog_v0p0p1_8.RSfetsym_0.QN VDD 2.55f
C831 frontAnalog_v0p0p1_4.RSfetsym_0.QN a_59577_n19683# 0.418f
C832 a_77605_n51335# I2 0.167f
C833 frontAnalog_v0p0p1_1.x65.X frontAnalog_v0p0p1_1.RSfetsym_0.x2.Y 0.526f
C834 frontAnalog_v0p0p1_1.RSfetsym_0.QN frontAnalog_v0p0p1_1.x63.X 0.378f
C835 16to4_PriorityEncoder_v0p0p1_0.x3.x4.A I2 0.0109f
C836 w_55000_n68350# VDD 0.829f
C837 frontAnalog_v0p0p1_11.x63.A frontAnalog_v0p0p1_11.x65.A 3.16f
C838 16to4_PriorityEncoder_v0p0p1_0.x5.x4.A 16to4_PriorityEncoder_v0p0p1_0.x5.x2.X 0.125f
C839 frontAnalog_v0p0p1_3.x63.X a_59577_n14283# 0.28f
C840 frontAnalog_v0p0p1_10.RSfetsym_0.x2.Y VDD 0.926f
C841 frontAnalog_v0p0p1_3.x63.A frontAnalog_v0p0p1_3.x65.A 3.16f
C842 frontAnalog_v0p0p1_4.x65.A CLK 2.63f
C843 a_59578_n40770# I8 0.42f
C844 16to4_PriorityEncoder_v0p0p1_0.x3.EI 16to4_PriorityEncoder_v0p0p1_0.x3.x19.X 0.0149f
C845 a_59577_n68283# VDD 0.0172f
C846 frontAnalog_v0p0p1_6.RSfetsym_0.x1.Y frontAnalog_v0p0p1_6.RSfetsym_0.x2.Y 0.0254f
C847 w_55000_n2928# a_53630_n3996# 0.359f
C848 CLK I15 0.0832f
C849 16to4_PriorityEncoder_v0p0p1_0.x3.EI 16to4_PriorityEncoder_v0p0p1_0.x5.x14.A 0.0145f
C850 w_55000_n19128# frontAnalog_v0p0p1_10.IB 0.0216f
C851 a_55268_n74136# VIN 0.177f
C852 frontAnalog_v0p0p1_1.x63.A VV9 0.587f
C853 frontAnalog_v0p0p1_3.RSfetsym_0.x1.Y I13 0.0436f
C854 frontAnalog_v0p0p1_7.x63.X CLK 0.46f
C855 frontAnalog_v0p0p1_15.x65.X a_59578_n83970# 0.436f
C856 VIN R0 0.188f
C857 16to4_PriorityEncoder_v0p0p1_0.x3.x16.X I3 0.0148f
C858 w_55000_n24528# CLK 0.57f
C859 a_53630_n3996# VDD 0.134f
C860 w_55000_n25150# a_55268_n25536# 0.12f
C861 w_55000_n79150# S1 0.0988f
C862 a_57123_n79679# CLK 0.0108f
C863 a_78349_n43045# 16to4_PriorityEncoder_v0p0p1_0.x5.x15.X 0.219f
C864 a_59577_n46683# I7 0.29f
C865 frontAnalog_v0p0p1_5.x65.A VIN 0.655f
C866 w_55000_n79150# VIN 0.737f
C867 16to4_PriorityEncoder_v0p0p1_0.x3.x21.B 16to4_PriorityEncoder_v0p0p1_0.x3.x21.X 0.0197f
C868 a_55268_n84936# R0 1.24f
C869 frontAnalog_v0p0p1_0.x63.X m3_58396_n9750# 0.134f
C870 a_77605_n39305# I11 0.0597f
C871 16to4_PriorityEncoder_v0p0p1_0.x3.x22.A 16to4_PriorityEncoder_v0p0p1_0.x3.A0 0.132f
C872 m3_58396_n63750# I4 0.0416f
C873 a_59578_n83970# I0 0.42f
C874 a_53630_n79596# VV2 0.28f
C875 m3_58396_n42150# CLK 0.189f
C876 frontAnalog_v0p0p1_0.x63.A a_57123_n9479# 0.212f
C877 a_59577_n19683# I12 0.29f
C878 VV12 VV11 3.43f
C879 frontAnalog_v0p0p1_14.RSfetsym_0.QN CLK 0.0457f
C880 frontAnalog_v0p0p1_7.x63.A VV10 0.587f
C881 16to4_PriorityEncoder_v0p0p1_0.x28.A 16to4_PriorityEncoder_v0p0p1_0.x29.A 0.392f
C882 16to4_PriorityEncoder_v0p0p1_0.x5.x18.C I15 0.229f
C883 frontAnalog_v0p0p1_6.x65.A a_57123_n29559# 0.214f
C884 16to4_PriorityEncoder_v0p0p1_0.x3.x19.D a_77605_n52567# 0.14f
C885 a_78525_n45515# 16to4_PriorityEncoder_v0p0p1_0.x5.x21.X 0.202f
C886 w_55000_n83928# a_53630_n84996# 0.359f
C887 w_55000_n62328# VV5 0.798f
C888 16to4_PriorityEncoder_v0p0p1_0.x5.x11.X a_78065_n41309# 0.202f
C889 16to4_PriorityEncoder_v0p0p1_0.x43.A VDD 1.46f
C890 frontAnalog_v0p0p1_6.x63.X m3_58396_n31350# 0.134f
C891 VDD VV7 1.87f
C892 frontAnalog_v0p0p1_6.RSfetsym_0.QN frontAnalog_v0p0p1_6.RSfetsym_0.x2.Y 0.018f
C893 16to4_PriorityEncoder_v0p0p1_0.x5.A2 a_82906_n43855# 0.208f
C894 frontAnalog_v0p0p1_4.x65.X VDD 3.46f
C895 16to4_PriorityEncoder_v0p0p1_0.x5.x4.A 16to4_PriorityEncoder_v0p0p1_0.x5.x1.X 0.118f
C896 a_77605_n44527# VDD 0.439f
C897 frontAnalog_v0p0p1_3.RSfetsym_0.QN I13 2.02f
C898 16to4_PriorityEncoder_v0p0p1_0.x5.x22.A 16to4_PriorityEncoder_v0p0p1_0.x5.x17.A 1.27f
C899 a_77637_n41087# 16to4_PriorityEncoder_v0p0p1_0.x5.x22.A 0.0288f
C900 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_6.x63.A 0.0926f
C901 a_53630_n47196# VV8 0.28f
C902 frontAnalog_v0p0p1_8.x63.X m3_58396_n47550# 0.134f
C903 frontAnalog_v0p0p1_1.x63.A VDD 3.67f
C904 frontAnalog_v0p0p1_15.x65.X frontAnalog_v0p0p1_15.RSfetsym_0.x1.Y 0.182f
C905 16to4_PriorityEncoder_v0p0p1_0.x5.x19.C I8 0.12f
C906 16to4_PriorityEncoder_v0p0p1_0.x5.x2.X VDD 0.367f
C907 16to4_PriorityEncoder_v0p0p1_0.x3.x19.D I3 1.27f
C908 w_55000_n3550# VIN 0.735f
C909 frontAnalog_v0p0p1_10.x65.X I5 0.446f
C910 w_55000_n57550# frontAnalog_v0p0p1_10.IB 0.0217f
C911 frontAnalog_v0p0p1_6.x63.X a_59577_n30483# 0.28f
C912 frontAnalog_v0p0p1_0.x65.A frontAnalog_v0p0p1_0.x65.X 0.0236f
C913 a_77637_n41087# I13 0.194f
C914 frontAnalog_v0p0p1_10.IB VV2 3.87f
C915 frontAnalog_v0p0p1_10.IB a_53630_n57996# 0.473f
C916 16to4_PriorityEncoder_v0p0p1_0.x22.A 16to4_PriorityEncoder_v0p0p1_0.x22.Y 1.51f
C917 frontAnalog_v0p0p1_10.IB a_55268_n9336# 0.0848f
C918 VV16 VFS 4.16f
C919 w_55000_n62950# CLK 0.535f
C920 w_55000_n73750# a_53630_n74196# 0.394f
C921 16to4_PriorityEncoder_v0p0p1_0.x1.A 16to4_PriorityEncoder_v0p0p1_0.x3.A2 1.46f
C922 w_55000_n73128# a_55268_n74136# 0.149f
C923 frontAnalog_v0p0p1_15.RSfetsym_0.x1.Y I0 0.0436f
C924 a_57123_n56559# CLK 0.0108f
C925 16to4_PriorityEncoder_v0p0p1_0.x5.x19.D a_77605_n44527# 0.14f
C926 16to4_PriorityEncoder_v0p0p1_0.x3.x19.D I2 0.196f
C927 frontAnalog_v0p0p1_10.IB R1 0.0926f
C928 frontAnalog_v0p0p1_0.x65.X CLK 0.443f
C929 frontAnalog_v0p0p1_4.x63.X VDD 3.13f
C930 frontAnalog_v0p0p1_6.x63.A frontAnalog_v0p0p1_6.x63.X 0.0301f
C931 16to4_PriorityEncoder_v0p0p1_0.x5.x4.A 16to4_PriorityEncoder_v0p0p1_0.x5.EO 0.0491f
C932 frontAnalog_v0p0p1_9.x65.A VV7 0.252f
C933 16to4_PriorityEncoder_v0p0p1_0.x5.x19.D 16to4_PriorityEncoder_v0p0p1_0.x5.x2.X 0.014f
C934 w_55000_n35328# VDD 0.854f
C935 frontAnalog_v0p0p1_3.RSfetsym_0.x2.Y I13 0.196f
C936 VDD VV1 1.57f
C937 frontAnalog_v0p0p1_12.x63.A a_55268_n74136# 1.24f
C938 VV14 VV13 4.07f
C939 w_55000_n40728# frontAnalog_v0p0p1_1.x65.A 0.658f
C940 a_57123_n83559# VDD 0.218f
C941 CLK I8 0.112f
C942 a_53630_n30996# VV11 0.28f
C943 frontAnalog_v0p0p1_10.IB a_53630_n47196# 0.473f
C944 frontAnalog_v0p0p1_15.RSfetsym_0.x1.Y frontAnalog_v0p0p1_15.x63.X 0.883f
C945 VIN VV12 3.41f
C946 frontAnalog_v0p0p1_10.x63.X I5 1.85f
C947 a_78525_n45515# VDD 0.165f
C948 I12 I10 0.849f
C949 frontAnalog_v0p0p1_8.RSfetsym_0.QN a_59578_n46170# 0.255f
C950 m3_58396_n63750# VDD 1.25f
C951 frontAnalog_v0p0p1_11.x63.A VDD 3.67f
C952 a_59578_n73170# I2 0.42f
C953 a_57123_n45759# CLK 0.0108f
C954 frontAnalog_v0p0p1_3.x63.A VDD 3.67f
C955 w_55000_n41350# frontAnalog_v0p0p1_1.x63.A 0.659f
C956 16to4_PriorityEncoder_v0p0p1_0.x42.A VDD 0.536f
C957 frontAnalog_v0p0p1_10.x65.A VDD 3.44f
C958 16to4_PriorityEncoder_v0p0p1_0.x35.A 16to4_PriorityEncoder_v0p0p1_0.x36.A 0.392f
C959 frontAnalog_v0p0p1_15.x65.X frontAnalog_v0p0p1_15.RSfetsym_0.QN 2.28f
C960 a_78349_n43045# VDD 0.164f
C961 a_53630_n14796# VIN 0.265f
C962 CLK VV13 0.645f
C963 frontAnalog_v0p0p1_7.x63.A CLK 1.8f
C964 frontAnalog_v0p0p1_1.RSfetsym_0.QN frontAnalog_v0p0p1_1.RSfetsym_0.x2.Y 0.018f
C965 16to4_PriorityEncoder_v0p0p1_0.x3.A2 16to4_PriorityEncoder_v0p0p1_0.x3.x14.A 0.074f
C966 frontAnalog_v0p0p1_0.x63.X CLK 0.46f
C967 I13 I9 0.376f
C968 16to4_PriorityEncoder_v0p0p1_0.x5.x17.A a_77637_n42017# 0.14f
C969 a_59578_n83970# VDD 0.0209f
C970 16to4_PriorityEncoder_v0p0p1_0.x5.x11.X 16to4_PriorityEncoder_v0p0p1_0.x5.x17.A 0.125f
C971 a_55268_n52536# VDD 0.565f
C972 frontAnalog_v0p0p1_15.x63.X a_57123_n85079# 0.121f
C973 a_77637_n41087# 16to4_PriorityEncoder_v0p0p1_0.x5.x11.X 0.109f
C974 w_55000_n46128# VIN 0.866f
C975 16to4_PriorityEncoder_v0p0p1_0.x5.x1.X VDD 0.39f
C976 16to4_PriorityEncoder_v0p0p1_0.x5.x18.C I8 0.119f
C977 frontAnalog_v0p0p1_15.RSfetsym_0.QN I0 2.02f
C978 frontAnalog_v0p0p1_10.IB a_55268_n68736# 0.0848f
C979 16to4_PriorityEncoder_v0p0p1_0.x5.x22.A 16to4_PriorityEncoder_v0p0p1_0.x5.x19.X 0.418f
C980 frontAnalog_v0p0p1_8.x63.A a_55268_n47136# 1.24f
C981 a_77605_n48109# I7 0.0614f
C982 frontAnalog_v0p0p1_12.x65.A VV3 0.253f
C983 frontAnalog_v0p0p1_11.x63.A a_55268_n63336# 1.24f
C984 w_55000_n73750# VV3 0.751f
C985 frontAnalog_v0p0p1_8.x65.X frontAnalog_v0p0p1_8.x63.X 0.143f
C986 I15 I11 1.03f
C987 frontAnalog_v0p0p1_13.x65.X CLK 0.443f
C988 frontAnalog_v0p0p1_15.RSfetsym_0.QN frontAnalog_v0p0p1_15.x63.X 0.378f
C989 frontAnalog_v0p0p1_15.x65.X frontAnalog_v0p0p1_15.RSfetsym_0.x2.Y 0.526f
C990 VV5 VV4 5.09f
C991 a_55268_n20136# CLK 0.235f
C992 16to4_PriorityEncoder_v0p0p1_0.x3.x16.C I3 0.132f
C993 frontAnalog_v0p0p1_12.x65.A VDD 3.44f
C994 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_4.x65.A 0.0352f
C995 a_59578_n35370# I9 0.42f
C996 16to4_PriorityEncoder_v0p0p1_0.x5.x16.X 16to4_PriorityEncoder_v0p0p1_0.x1.A 0.0159f
C997 a_53630_n30996# VIN 0.265f
C998 frontAnalog_v0p0p1_1.x65.X I9 0.0396f
C999 w_55000_n73750# VDD 0.829f
C1000 frontAnalog_v0p0p1_12.RSfetsym_0.x1.Y I2 0.0436f
C1001 a_57123_n2559# frontAnalog_v0p0p1_2.x65.X 0.119f
C1002 I14 I12 2.36f
C1003 16to4_PriorityEncoder_v0p0p1_0.x5.EO VDD 1.06f
C1004 frontAnalog_v0p0p1_15.RSfetsym_0.x2.Y I0 0.198f
C1005 w_55000_n30550# a_53630_n30996# 0.394f
C1006 w_55000_n29928# a_55268_n30936# 0.149f
C1007 16to4_PriorityEncoder_v0p0p1_0.x5.x4.A I10 0.0109f
C1008 frontAnalog_v0p0p1_0.x63.A VV15 0.587f
C1009 frontAnalog_v0p0p1_9.x65.A a_55268_n52536# 0.461f
C1010 16to4_PriorityEncoder_v0p0p1_0.x5.x22.A I13 0.066f
C1011 w_55000_n3550# a_55268_n3936# 0.12f
C1012 16to4_PriorityEncoder_v0p0p1_0.x3.x16.C I2 0.925f
C1013 w_55000_n24528# frontAnalog_v0p0p1_10.IB 0.0216f
C1014 m3_58396_n36750# I9 0.0416f
C1015 frontAnalog_v0p0p1_0.x63.A VIN 0.19f
C1016 a_59577_n19683# VDD 0.0172f
C1017 16to4_PriorityEncoder_v0p0p1_0.x5.x21.B a_77605_n44779# 0.0141f
C1018 16to4_PriorityEncoder_v0p0p1_0.x1.X 16to4_PriorityEncoder_v0p0p1_0.x28.A 0.0747f
C1019 a_55268_n25536# VIN 0.177f
C1020 frontAnalog_v0p0p1_13.x63.X CLK 0.46f
C1021 frontAnalog_v0p0p1_15.RSfetsym_0.x1.Y VDD 0.733f
C1022 frontAnalog_v0p0p1_15.x63.X frontAnalog_v0p0p1_15.RSfetsym_0.x2.Y 0.0923f
C1023 m3_58396_n58350# I5 0.0416f
C1024 a_59577_n57483# I5 0.29f
C1025 a_59577_n41283# I8 0.29f
C1026 16to4_PriorityEncoder_v0p0p1_0.x3.A2 16to4_PriorityEncoder_v0p0p1_0.x2.A 0.401f
C1027 frontAnalog_v0p0p1_13.x65.A a_55268_n68736# 0.461f
C1028 w_55000_n29928# CLK 0.57f
C1029 16to4_PriorityEncoder_v0p0p1_0.x3.EI 16to4_PriorityEncoder_v0p0p1_0.x5.x17.A 0.0296f
C1030 a_57123_n2559# VDD 0.222f
C1031 frontAnalog_v0p0p1_9.x63.X a_57123_n52679# 0.121f
C1032 a_53630_n84996# CLK 0.0136f
C1033 frontAnalog_v0p0p1_12.RSfetsym_0.QN I3 0.0512f
C1034 VIN VV6 3.41f
C1035 frontAnalog_v0p0p1_2.x65.X a_59578_n2970# 0.436f
C1036 w_55000_n84550# VIN 0.737f
C1037 16to4_PriorityEncoder_v0p0p1_0.x5.GS VDD 0.771f
C1038 m3_58396_n52950# CLK 0.189f
C1039 16to4_PriorityEncoder_v0p0p1_0.x3.x20.X VDD 0.242f
C1040 a_57123_n58079# CLK 0.0108f
C1041 frontAnalog_v0p0p1_7.RSfetsym_0.x1.Y I9 0.0433f
C1042 w_55000_n40728# VV9 0.798f
C1043 a_77605_n52819# VDD 0.435f
C1044 w_55000_n83928# VV1 0.798f
C1045 16to4_PriorityEncoder_v0p0p1_0.x21.A 16to4_PriorityEncoder_v0p0p1_0.x22.A 0.392f
C1046 w_55000_n84550# a_55268_n84936# 0.12f
C1047 w_55000_n56928# a_55268_n57936# 0.149f
C1048 frontAnalog_v0p0p1_12.RSfetsym_0.QN I2 2.02f
C1049 w_55000_n57550# a_53630_n57996# 0.394f
C1050 a_57123_n85079# VDD 0.221f
C1051 a_57123_n51159# frontAnalog_v0p0p1_9.x65.X 0.119f
C1052 a_59578_n2970# VDD 0.0209f
C1053 frontAnalog_v0p0p1_10.RSfetsym_0.QN CLK 0.0457f
C1054 16to4_PriorityEncoder_v0p0p1_0.x5.x15.X 16to4_PriorityEncoder_v0p0p1_0.x1.A 0.0206f
C1055 CLK I3 0.0837f
C1056 w_55000_n19128# frontAnalog_v0p0p1_4.x65.A 0.658f
C1057 frontAnalog_v0p0p1_15.x63.X R0 0.0402f
C1058 a_53630_n74196# a_55268_n74136# 0.015f
C1059 VV2 R1 0.587f
C1060 frontAnalog_v0p0p1_15.RSfetsym_0.QN VDD 2.56f
C1061 16to4_PriorityEncoder_v0p0p1_0.x5.x11.X 16to4_PriorityEncoder_v0p0p1_0.x5.x22.A 0.0936f
C1062 w_55000_n8950# VV15 0.751f
C1063 frontAnalog_v0p0p1_15.RSfetsym_0.QN a_59577_n84483# 0.418f
C1064 w_55000_n8950# VIN 0.737f
C1065 w_55000_n62950# frontAnalog_v0p0p1_10.IB 0.0217f
C1066 16to4_PriorityEncoder_v0p0p1_0.x5.x11.X I13 0.0201f
C1067 I11 I8 0.672f
C1068 frontAnalog_v0p0p1_9.x63.X frontAnalog_v0p0p1_9.RSfetsym_0.x2.Y 0.0923f
C1069 a_77637_n40777# I12 0.188f
C1070 frontAnalog_v0p0p1_10.x63.A VV6 0.587f
C1071 VDD I10 5.31f
C1072 frontAnalog_v0p0p1_8.RSfetsym_0.QN frontAnalog_v0p0p1_8.RSfetsym_0.x2.Y 0.018f
C1073 frontAnalog_v0p0p1_12.RSfetsym_0.x2.Y I2 0.198f
C1074 frontAnalog_v0p0p1_13.x63.A VV4 0.587f
C1075 a_53630_n63396# VDD 0.134f
C1076 w_55000_n19750# frontAnalog_v0p0p1_4.x63.A 0.659f
C1077 frontAnalog_v0p0p1_2.x65.X frontAnalog_v0p0p1_2.RSfetsym_0.x1.Y 0.182f
C1078 CLK I2 0.0837f
C1079 16to4_PriorityEncoder_v0p0p1_0.x3.x19.C a_77605_n52567# 0.157f
C1080 frontAnalog_v0p0p1_8.RSfetsym_0.QN CLK 0.0457f
C1081 frontAnalog_v0p0p1_12.x65.A a_57123_n72759# 0.214f
C1082 w_55000_n68350# CLK 0.535f
C1083 16to4_PriorityEncoder_v0p0p1_0.x34.A 16to4_PriorityEncoder_v0p0p1_0.x35.A 0.0737f
C1084 frontAnalog_v0p0p1_7.RSfetsym_0.QN I9 2.02f
C1085 16to4_PriorityEncoder_v0p0p1_0.x3.EI a_77637_n48817# 0.0883f
C1086 16to4_PriorityEncoder_v0p0p1_0.x5.x20.X 16to4_PriorityEncoder_v0p0p1_0.x2.A 0.0148f
C1087 w_55000_n40728# VDD 0.854f
C1088 frontAnalog_v0p0p1_15.RSfetsym_0.x2.Y VDD 0.926f
C1089 16to4_PriorityEncoder_v0p0p1_0.x3.x21.B 16to4_PriorityEncoder_v0p0p1_0.x3.x19.X 0.262f
C1090 frontAnalog_v0p0p1_9.x63.A VDD 3.67f
C1091 16to4_PriorityEncoder_v0p0p1_0.x5.x19.D I10 0.196f
C1092 frontAnalog_v0p0p1_2.RSfetsym_0.x1.Y VDD 0.733f
C1093 w_55000_n78528# w_55000_n79150# 0.327f
C1094 16to4_PriorityEncoder_v0p0p1_0.x3.x19.C I3 0.921f
C1095 frontAnalog_v0p0p1_9.x63.X a_59577_n52083# 0.28f
C1096 frontAnalog_v0p0p1_10.IB VV13 3.88f
C1097 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_7.x63.A 0.0926f
C1098 w_55000_n35328# VV10 0.798f
C1099 a_53630_n63396# a_55268_n63336# 0.015f
C1100 frontAnalog_v0p0p1_2.RSfetsym_0.x1.Y frontAnalog_v0p0p1_2.x63.X 0.883f
C1101 m3_58396_n74550# VDD 1.25f
C1102 a_53630_n3996# CLK 0.0136f
C1103 16to4_PriorityEncoder_v0p0p1_0.x3.x14.A I4 0.0493f
C1104 frontAnalog_v0p0p1_8.x65.A a_57123_n45759# 0.214f
C1105 frontAnalog_v0p0p1_5.x63.A frontAnalog_v0p0p1_5.x65.A 3.16f
C1106 16to4_PriorityEncoder_v0p0p1_0.x3.EI 16to4_PriorityEncoder_v0p0p1_0.x5.x22.A 0.208f
C1107 frontAnalog_v0p0p1_7.RSfetsym_0.x2.Y I9 0.192f
C1108 16to4_PriorityEncoder_v0p0p1_0.x5.x19.C a_77605_n44527# 0.157f
C1109 a_55268_n74136# VV3 0.215f
C1110 16to4_PriorityEncoder_v0p0p1_0.x3.x19.C I2 0.447f
C1111 frontAnalog_v0p0p1_11.x65.A a_57123_n61959# 0.214f
C1112 frontAnalog_v0p0p1_2.x65.X frontAnalog_v0p0p1_2.RSfetsym_0.QN 2.28f
C1113 frontAnalog_v0p0p1_12.x63.A frontAnalog_v0p0p1_12.x63.X 0.0301f
C1114 VDD I14 5.92f
C1115 a_77605_n51585# I3 0.162f
C1116 frontAnalog_v0p0p1_9.x65.X VDD 3.46f
C1117 w_55000_n51528# VIN 0.866f
C1118 16to4_PriorityEncoder_v0p0p1_0.x3.x21.X VDD 0.501f
C1119 a_57123_n4079# VDD 0.222f
C1120 VIN VV5 3.41f
C1121 a_55268_n74136# VDD 0.565f
C1122 w_55000_n67728# frontAnalog_v0p0p1_13.x63.A 0.0792f
C1123 frontAnalog_v0p0p1_10.IB a_55268_n20136# 0.0848f
C1124 frontAnalog_v0p0p1_9.x63.A frontAnalog_v0p0p1_9.x65.A 3.16f
C1125 frontAnalog_v0p0p1_2.x63.X a_57123_n4079# 0.121f
C1126 16to4_PriorityEncoder_v0p0p1_0.x3.A2 16to4_PriorityEncoder_v0p0p1_0.x3.A1 0.787f
C1127 w_55000_n40728# w_55000_n41350# 0.327f
C1128 16to4_PriorityEncoder_v0p0p1_0.x3.x19.D a_77605_n52819# 0.148f
C1129 frontAnalog_v0p0p1_7.x63.A a_55268_n36336# 1.24f
C1130 VDD R0 3.89f
C1131 16to4_PriorityEncoder_v0p0p1_0.x3.x18.C a_77605_n52567# 0.117f
C1132 CLK VV7 0.645f
C1133 a_78159_n47589# VDD 0.152f
C1134 frontAnalog_v0p0p1_3.x63.A a_55268_n14736# 1.24f
C1135 16to4_PriorityEncoder_v0p0p1_0.x3.x4.A a_78159_n47589# 0.299f
C1136 m3_58396_n52950# I6 0.0416f
C1137 16to4_PriorityEncoder_v0p0p1_0.x1.A VDD 2.17f
C1138 frontAnalog_v0p0p1_4.x65.X CLK 0.443f
C1139 frontAnalog_v0p0p1_13.x63.A a_57123_n68879# 0.212f
C1140 frontAnalog_v0p0p1_2.RSfetsym_0.QN VDD 2.55f
C1141 16to4_PriorityEncoder_v0p0p1_0.x5.x19.D I14 0.464f
C1142 w_55000_n79150# VDD 0.829f
C1143 frontAnalog_v0p0p1_5.x65.A VDD 3.44f
C1144 frontAnalog_v0p0p1_1.x63.A CLK 1.8f
C1145 frontAnalog_v0p0p1_2.RSfetsym_0.QN frontAnalog_v0p0p1_2.x63.X 0.378f
C1146 frontAnalog_v0p0p1_2.x65.X frontAnalog_v0p0p1_2.RSfetsym_0.x2.Y 0.526f
C1147 a_77605_n44779# VDD 0.614f
C1148 a_57123_n79679# R1 0.222f
C1149 VV16 VV15 4.68f
C1150 frontAnalog_v0p0p1_10.RSfetsym_0.QN I6 0.0512f
C1151 frontAnalog_v0p0p1_9.x65.A frontAnalog_v0p0p1_9.x65.X 0.0236f
C1152 16to4_PriorityEncoder_v0p0p1_0.x3.x18.C I3 0.251f
C1153 VIN VV16 3.02f
C1154 I6 I3 0.602f
C1155 frontAnalog_v0p0p1_14.x65.X I1 0.446f
C1156 frontAnalog_v0p0p1_7.RSfetsym_0.QN a_59578_n35370# 0.255f
C1157 w_55000_n29928# frontAnalog_v0p0p1_10.IB 0.0216f
C1158 frontAnalog_v0p0p1_11.x63.X m3_58396_n63750# 0.134f
C1159 frontAnalog_v0p0p1_11.x63.A frontAnalog_v0p0p1_11.x63.X 0.0301f
C1160 I7 I1 0.244f
C1161 frontAnalog_v0p0p1_10.IB a_53630_n84996# 0.473f
C1162 16to4_PriorityEncoder_v0p0p1_0.x2.X 16to4_PriorityEncoder_v0p0p1_0.x21.A 0.0749f
C1163 w_55000_n19128# VV13 0.798f
C1164 frontAnalog_v0p0p1_2.x65.A VIN 0.653f
C1165 w_55000_n51528# a_53630_n52596# 0.359f
C1166 m3_58396_n85350# I0 0.0416f
C1167 16to4_PriorityEncoder_v0p0p1_0.x3.x14.A a_78065_n49349# 0.197f
C1168 frontAnalog_v0p0p1_3.x63.A VV14 0.587f
C1169 w_55000_n2928# w_55000_n3550# 0.327f
C1170 frontAnalog_v0p0p1_4.x63.X CLK 0.46f
C1171 frontAnalog_v0p0p1_9.x65.X frontAnalog_v0p0p1_9.RSfetsym_0.QN 2.28f
C1172 frontAnalog_v0p0p1_2.RSfetsym_0.x2.Y VDD 0.926f
C1173 frontAnalog_v0p0p1_13.x65.A frontAnalog_v0p0p1_13.x65.X 0.0236f
C1174 16to4_PriorityEncoder_v0p0p1_0.x5.x16.C I10 0.925f
C1175 16to4_PriorityEncoder_v0p0p1_0.x5.x19.D a_77605_n44779# 0.148f
C1176 w_55000_n35328# CLK 0.57f
C1177 CLK VV1 0.618f
C1178 16to4_PriorityEncoder_v0p0p1_0.x5.x18.C a_77605_n44527# 0.117f
C1179 frontAnalog_v0p0p1_14.RSfetsym_0.QN a_59578_n78570# 0.255f
C1180 I5 I0 0.344f
C1181 frontAnalog_v0p0p1_5.x63.A VV12 0.587f
C1182 a_57123_n83559# CLK 0.0108f
C1183 16to4_PriorityEncoder_v0p0p1_0.x3.x14.A VDD 0.462f
C1184 16to4_PriorityEncoder_v0p0p1_0.x3.x18.C I2 0.341f
C1185 I2 I6 0.441f
C1186 frontAnalog_v0p0p1_2.x63.X frontAnalog_v0p0p1_2.RSfetsym_0.x2.Y 0.0923f
C1187 frontAnalog_v0p0p1_15.x63.X m3_58396_n85350# 0.139f
C1188 w_55000_n3550# VDD 0.829f
C1189 a_77605_n39305# I8 0.211f
C1190 a_77605_n40069# I15 0.0614f
C1191 frontAnalog_v0p0p1_8.x63.A VIN 0.186f
C1192 a_59578_n62370# I4 0.42f
C1193 a_53630_n36396# VIN 0.265f
C1194 16to4_PriorityEncoder_v0p0p1_0.x3.EI I1 0.437f
C1195 m3_58396_n63750# CLK 0.189f
C1196 frontAnalog_v0p0p1_11.x63.A CLK 1.8f
C1197 frontAnalog_v0p0p1_14.x63.X I1 1.85f
C1198 frontAnalog_v0p0p1_3.x63.A CLK 1.8f
C1199 frontAnalog_v0p0p1_7.x65.X frontAnalog_v0p0p1_7.x63.X 0.143f
C1200 frontAnalog_v0p0p1_10.x65.A CLK 2.63f
C1201 a_77637_n40777# VDD 0.318f
C1202 I4 I5 6.86f
C1203 a_53630_n68796# VV4 0.28f
C1204 w_55000_n19128# a_55268_n20136# 0.149f
C1205 w_55000_n19750# a_53630_n20196# 0.394f
C1206 frontAnalog_v0p0p1_1.x65.X frontAnalog_v0p0p1_1.RSfetsym_0.QN 2.28f
C1207 m3_58396_n4350# VDD 1.25f
C1208 a_78349_n51085# VDD 0.164f
C1209 frontAnalog_v0p0p1_2.x63.X m3_58396_n4350# 0.134f
C1210 16to4_PriorityEncoder_v0p0p1_0.x3.EI I7 4.79f
C1211 frontAnalog_v0p0p1_14.x65.X frontAnalog_v0p0p1_14.x63.X 0.143f
C1212 a_55268_n52536# CLK 0.235f
C1213 frontAnalog_v0p0p1_7.RSfetsym_0.QN frontAnalog_v0p0p1_7.RSfetsym_0.x1.Y 0.17f
C1214 frontAnalog_v0p0p1_8.RSfetsym_0.x1.Y frontAnalog_v0p0p1_8.x63.X 0.883f
C1215 VDD VV12 1.84f
C1216 16to4_PriorityEncoder_v0p0p1_0.x5.x22.A a_77639_n42341# 0.155f
C1217 frontAnalog_v0p0p1_13.x63.A VIN 0.188f
C1218 a_77639_n50381# VDD 0.23f
C1219 w_55000_n14350# VIN 0.737f
C1220 a_55268_n41736# VIN 0.177f
C1221 w_55000_n68350# frontAnalog_v0p0p1_10.IB 0.0217f
C1222 frontAnalog_v0p0p1_14.RSfetsym_0.QN frontAnalog_v0p0p1_14.RSfetsym_0.x1.Y 0.17f
C1223 16to4_PriorityEncoder_v0p0p1_0.x43.Y 16to4_PriorityEncoder_v0p0p1_0.x5.A2 0.0114f
C1224 16to4_PriorityEncoder_v0p0p1_0.x5.x14.A I12 0.0493f
C1225 16to4_PriorityEncoder_v0p0p1_0.x5.x16.C I14 0.491f
C1226 frontAnalog_v0p0p1_2.RSfetsym_0.QN a_59577_n3483# 0.418f
C1227 a_57123_n61959# VDD 0.222f
C1228 frontAnalog_v0p0p1_12.x65.A CLK 2.63f
C1229 a_53630_n14796# VDD 0.134f
C1230 w_55000_n73750# CLK 0.535f
C1231 frontAnalog_v0p0p1_11.RSfetsym_0.x1.Y I4 0.0436f
C1232 16to4_PriorityEncoder_v0p0p1_0.x2.A VDD 1.89f
C1233 frontAnalog_v0p0p1_7.RSfetsym_0.x1.Y frontAnalog_v0p0p1_7.RSfetsym_0.x2.Y 0.0254f
C1234 w_55000_n83928# R0 0.0792f
C1235 frontAnalog_v0p0p1_1.RSfetsym_0.x1.Y VDD 0.733f
C1236 frontAnalog_v0p0p1_4.x63.X m3_58396_n20550# 0.134f
C1237 w_55000_n46128# VDD 0.854f
C1238 VV1 S0 0.252f
C1239 a_57123_n83559# S0 0.229f
C1240 VV8 VV7 3.46f
C1241 a_78349_n51085# 16to4_PriorityEncoder_v0p0p1_0.x3.x16.X 0.0673f
C1242 w_55000_n13728# frontAnalog_v0p0p1_3.x63.A 0.0792f
C1243 frontAnalog_v0p0p1_10.IB a_53630_n3996# 0.472f
C1244 16to4_PriorityEncoder_v0p0p1_0.x3.x14.A 16to4_PriorityEncoder_v0p0p1_0.x3.x17.A 0.105f
C1245 w_55000_n52150# VV7 0.751f
C1246 frontAnalog_v0p0p1_5.x63.A a_55268_n25536# 1.24f
C1247 w_55000_n67728# a_53630_n68796# 0.359f
C1248 frontAnalog_v0p0p1_14.RSfetsym_0.x1.Y frontAnalog_v0p0p1_14.RSfetsym_0.x2.Y 0.0254f
C1249 a_55268_n3936# VV16 0.214f
C1250 a_59578_n62370# VDD 0.0209f
C1251 m3_58396_n85350# VDD 1.3f
C1252 a_57123_n2559# CLK 0.0108f
C1253 frontAnalog_v0p0p1_2.x65.A a_55268_n3936# 0.461f
C1254 a_55268_n79536# S1 0.461f
C1255 a_53630_n30996# VDD 0.134f
C1256 VDD I5 4.26f
C1257 w_55000_n68350# frontAnalog_v0p0p1_13.x65.A 0.0988f
C1258 a_59577_n79083# I1 0.29f
C1259 16to4_PriorityEncoder_v0p0p1_0.x3.x4.A I5 0.0107f
C1260 16to4_PriorityEncoder_v0p0p1_0.x3.x17.A a_78349_n51085# 0.213f
C1261 a_55268_n79536# VIN 0.177f
C1262 frontAnalog_v0p0p1_7.x65.A a_57123_n34959# 0.214f
C1263 a_78097_n53777# 16to4_PriorityEncoder_v0p0p1_0.x3.x20.X 0.137f
C1264 m3_58396_n9750# I14 0.0416f
C1265 VDD OUT1 6.71f
C1266 w_55000_n56928# VIN 0.866f
C1267 frontAnalog_v0p0p1_3.x65.A a_57123_n13359# 0.214f
C1268 frontAnalog_v0p0p1_10.IB VV7 3.87f
C1269 frontAnalog_v0p0p1_9.x65.X frontAnalog_v0p0p1_9.RSfetsym_0.x1.Y 0.182f
C1270 frontAnalog_v0p0p1_11.RSfetsym_0.QN I4 2.02f
C1271 frontAnalog_v0p0p1_0.x63.A VDD 3.67f
C1272 a_53630_n9396# VV15 0.28f
C1273 16to4_PriorityEncoder_v0p0p1_0.x5.x19.C I10 0.447f
C1274 frontAnalog_v0p0p1_12.x65.X VDD 3.46f
C1275 w_55000_n29928# frontAnalog_v0p0p1_6.x63.A 0.0792f
C1276 a_77605_n53805# VDD 0.201f
C1277 frontAnalog_v0p0p1_7.RSfetsym_0.QN frontAnalog_v0p0p1_7.RSfetsym_0.x2.Y 0.018f
C1278 a_53630_n9396# VIN 0.265f
C1279 a_55268_n25536# VDD 0.565f
C1280 frontAnalog_v0p0p1_1.x63.X VDD 3.13f
C1281 I15 I8 0.342f
C1282 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_1.x63.A 0.0926f
C1283 16to4_PriorityEncoder_v0p0p1_0.x3.x22.A 16to4_PriorityEncoder_v0p0p1_0.x3.x21.X 0.0749f
C1284 frontAnalog_v0p0p1_11.x65.A VV5 0.253f
C1285 m3_58396_n47550# I7 0.0416f
C1286 VDD VV6 1.84f
C1287 frontAnalog_v0p0p1_7.x63.X a_59577_n35883# 0.28f
C1288 frontAnalog_v0p0p1_14.RSfetsym_0.QN frontAnalog_v0p0p1_14.RSfetsym_0.x2.Y 0.018f
C1289 a_53630_n25596# VV12 0.28f
C1290 w_55000_n84550# VDD 0.829f
C1291 frontAnalog_v0p0p1_11.RSfetsym_0.x1.Y VDD 0.733f
C1292 frontAnalog_v0p0p1_4.x65.A VV13 0.253f
C1293 a_78349_n51085# 16to4_PriorityEncoder_v0p0p1_0.x3.x15.X 0.219f
C1294 frontAnalog_v0p0p1_11.RSfetsym_0.x2.Y I4 0.198f
C1295 frontAnalog_v0p0p1_8.x63.X VDD 3.13f
C1296 CLK I10 0.0757f
C1297 a_53630_n63396# CLK 0.0136f
C1298 frontAnalog_v0p0p1_12.x63.X VDD 3.13f
C1299 frontAnalog_v0p0p1_14.x63.X a_59577_n79083# 0.28f
C1300 w_55000_n35328# frontAnalog_v0p0p1_10.IB 0.0216f
C1301 frontAnalog_v0p0p1_10.IB VV1 0.0595f
C1302 m3_58396_n42150# I8 0.0416f
C1303 frontAnalog_v0p0p1_7.x63.A frontAnalog_v0p0p1_7.x63.X 0.0301f
C1304 16to4_PriorityEncoder_v0p0p1_0.x3.x19.C a_77605_n52819# 0.102f
C1305 w_55000_n52150# a_55268_n52536# 0.12f
C1306 frontAnalog_v0p0p1_3.x63.A frontAnalog_v0p0p1_3.x63.X 0.0301f
C1307 w_55000_n56928# frontAnalog_v0p0p1_10.x63.A 0.0792f
C1308 w_55000_n40728# CLK 0.57f
C1309 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_11.x63.A 0.0926f
C1310 16to4_PriorityEncoder_v0p0p1_0.x5.x19.C I14 0.305f
C1311 frontAnalog_v0p0p1_4.x65.A a_55268_n20136# 0.461f
C1312 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_3.x63.A 0.0926f
C1313 a_57123_n63479# VDD 0.222f
C1314 frontAnalog_v0p0p1_9.x63.A CLK 1.8f
C1315 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_10.x65.A 0.0352f
C1316 a_59578_n51570# VDD 0.0209f
C1317 a_77637_n49127# I5 0.194f
C1318 w_55000_n8950# VDD 0.829f
C1319 a_53630_n68796# VIN 0.265f
C1320 16to4_PriorityEncoder_v0p0p1_0.x3.x14.A 16to4_PriorityEncoder_v0p0p1_0.x3.x22.A 0.0179f
C1321 frontAnalog_v0p0p1_1.x65.A a_55268_n41736# 0.461f
C1322 m3_58396_n74550# CLK 0.189f
C1323 16to4_PriorityEncoder_v0p0p1_0.x5.x18.C I10 0.341f
C1324 16to4_PriorityEncoder_v0p0p1_0.x3.x19.X VDD 0.892f
C1325 16to4_PriorityEncoder_v0p0p1_0.x5.x14.A VDD 0.487f
C1326 16to4_PriorityEncoder_v0p0p1_0.x3.A1 VDD 1.93f
C1327 w_55000_n35328# a_55268_n36336# 0.149f
C1328 w_55000_n35950# a_53630_n36396# 0.394f
C1329 frontAnalog_v0p0p1_10.IB a_55268_n52536# 0.0848f
C1330 frontAnalog_v0p0p1_11.RSfetsym_0.QN VDD 2.55f
C1331 m3_58396_n15150# VDD 1.25f
C1332 frontAnalog_v0p0p1_6.x65.A VV11 0.253f
C1333 frontAnalog_v0p0p1_0.RSfetsym_0.QN a_59578_n8370# 0.255f
C1334 16to4_PriorityEncoder_v0p0p1_0.x5.x19.C a_77605_n44779# 0.102f
C1335 16to4_PriorityEncoder_v0p0p1_0.x3.x19.D I5 0.551f
C1336 CLK I14 0.089f
C1337 a_57123_n41879# VDD 0.222f
C1338 frontAnalog_v0p0p1_9.x65.X CLK 0.443f
C1339 16to4_PriorityEncoder_v0p0p1_0.x3.x22.A a_78349_n51085# 0.17f
C1340 a_57123_n4079# CLK 0.0108f
C1341 16to4_PriorityEncoder_v0p0p1_0.x5.x17.A 16to4_PriorityEncoder_v0p0p1_0.x5.x16.X 0.0198f
C1342 a_78097_n53777# 16to4_PriorityEncoder_v0p0p1_0.x3.x21.X 0.109f
C1343 a_57123_n72759# frontAnalog_v0p0p1_12.x65.X 0.119f
C1344 16to4_PriorityEncoder_v0p0p1_0.x5.x22.A a_77605_n43295# 0.0116f
C1345 a_55268_n74136# CLK 0.235f
C1346 frontAnalog_v0p0p1_8.x65.X I7 0.446f
C1347 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_12.x65.A 0.0352f
C1348 frontAnalog_v0p0p1_4.x63.A VIN 0.194f
C1349 w_55000_n19750# VIN 0.737f
C1350 a_53630_n25596# a_55268_n25536# 0.015f
C1351 CLK R0 1.81f
C1352 w_55000_n73750# frontAnalog_v0p0p1_10.IB 0.0217f
C1353 16to4_PriorityEncoder_v0p0p1_0.x3.x19.D a_77605_n53805# 0.0838f
C1354 frontAnalog_v0p0p1_11.RSfetsym_0.x2.Y VDD 0.926f
C1355 16to4_PriorityEncoder_v0p0p1_0.x3.x22.A a_77639_n50381# 0.155f
C1356 frontAnalog_v0p0p1_2.RSfetsym_0.QN CLK 0.0457f
C1357 w_55000_n40728# a_53630_n41796# 0.359f
C1358 a_57123_n13359# VDD 0.222f
C1359 frontAnalog_v0p0p1_2.x63.A a_57123_n4079# 0.212f
C1360 w_55000_n14350# frontAnalog_v0p0p1_3.x65.A 0.0988f
C1361 frontAnalog_v0p0p1_9.RSfetsym_0.QN a_59578_n51570# 0.255f
C1362 frontAnalog_v0p0p1_5.x65.A CLK 2.63f
C1363 w_55000_n79150# CLK 0.535f
C1364 a_59577_n46683# VDD 0.0172f
C1365 frontAnalog_v0p0p1_5.x65.A a_57123_n24159# 0.214f
C1366 a_59577_n73683# VDD 0.0172f
C1367 frontAnalog_v0p0p1_0.x65.X frontAnalog_v0p0p1_0.x63.X 0.143f
C1368 16to4_PriorityEncoder_v0p0p1_0.x5.x18.C I14 0.301f
C1369 a_77605_n39305# 16to4_PriorityEncoder_v0p0p1_0.x5.x2.X 0.0313f
C1370 16to4_PriorityEncoder_v0p0p1_0.x5.EO 16to4_PriorityEncoder_v0p0p1_0.x5.A2 0.136f
C1371 w_55000_n51528# VDD 0.854f
C1372 frontAnalog_v0p0p1_12.x65.X a_59578_n73170# 0.436f
C1373 16to4_PriorityEncoder_v0p0p1_0.x3.A1 16to4_PriorityEncoder_v0p0p1_0.x3.x16.X 0.0159f
C1374 VDD VV5 1.84f
C1375 16to4_PriorityEncoder_v0p0p1_0.x3.x14.A 16to4_PriorityEncoder_v0p0p1_0.x3.x11.X 0.0721f
C1376 w_55000_n83928# w_55000_n84550# 0.327f
C1377 frontAnalog_v0p0p1_0.RSfetsym_0.QN frontAnalog_v0p0p1_0.RSfetsym_0.x1.Y 0.17f
C1378 w_55000_n68350# a_55268_n68736# 0.12f
C1379 frontAnalog_v0p0p1_1.RSfetsym_0.x2.Y VDD 0.926f
C1380 a_57123_n61959# frontAnalog_v0p0p1_11.x65.X 0.119f
C1381 frontAnalog_v0p0p1_6.x65.A VIN 0.655f
C1382 a_59578_n13770# VDD 0.0209f
C1383 a_53630_n14796# a_55268_n14736# 0.015f
C1384 frontAnalog_v0p0p1_2.x65.A frontAnalog_v0p0p1_2.x65.X 0.0236f
C1385 frontAnalog_v0p0p1_14.x65.X S1 0.0378f
C1386 w_55000_n2928# VV16 0.798f
C1387 a_57123_n29559# VDD 0.222f
C1388 16to4_PriorityEncoder_v0p0p1_0.x3.A1 16to4_PriorityEncoder_v0p0p1_0.x3.x17.A 0.115f
C1389 a_77605_n48109# I4 0.208f
C1390 w_55000_n8328# frontAnalog_v0p0p1_0.x63.A 0.0792f
C1391 w_55000_n30550# frontAnalog_v0p0p1_6.x65.A 0.0988f
C1392 w_55000_n3550# CLK 0.535f
C1393 w_55000_n2928# frontAnalog_v0p0p1_2.x65.A 0.658f
C1394 16to4_PriorityEncoder_v0p0p1_0.x5.x17.A 16to4_PriorityEncoder_v0p0p1_0.x5.x15.X 0.0789f
C1395 16to4_PriorityEncoder_v0p0p1_0.x3.x22.A I5 0.066f
C1396 a_55268_n63336# VV5 0.215f
C1397 w_55000_n62328# VIN 0.866f
C1398 VDD VV16 2.41f
C1399 w_55000_n51528# frontAnalog_v0p0p1_9.x65.A 0.658f
C1400 16to4_PriorityEncoder_v0p0p1_0.x5.x19.X 16to4_PriorityEncoder_v0p0p1_0.x5.x20.X 0.145f
C1401 frontAnalog_v0p0p1_5.x63.A frontAnalog_v0p0p1_5.x63.X 0.0301f
C1402 frontAnalog_v0p0p1_0.RSfetsym_0.x1.Y frontAnalog_v0p0p1_0.RSfetsym_0.x2.Y 0.0254f
C1403 a_55268_n57936# VIN 0.177f
C1404 a_78065_n41309# VDD 0.161f
C1405 m3_58396_n4350# CLK 0.189f
C1406 a_78525_n53555# VDD 0.151f
C1407 16to4_PriorityEncoder_v0p0p1_0.x3.x16.C I5 0.415f
C1408 a_55268_n41736# VV9 0.215f
C1409 frontAnalog_v0p0p1_5.x65.X VDD 3.46f
C1410 frontAnalog_v0p0p1_2.x65.A VDD 3.44f
C1411 frontAnalog_v0p0p1_11.x65.X a_59578_n62370# 0.436f
C1412 I11 I10 7.54f
C1413 I12 I9 0.43f
C1414 16to4_PriorityEncoder_v0p0p1_0.x5.x21.B 16to4_PriorityEncoder_v0p0p1_0.x5.x19.X 0.262f
C1415 w_55000_n46128# w_55000_n46750# 0.327f
C1416 w_55000_n3550# frontAnalog_v0p0p1_2.x63.A 0.659f
C1417 16to4_PriorityEncoder_v0p0p1_0.x3.x19.D 16to4_PriorityEncoder_v0p0p1_0.x3.x19.X 0.0195f
C1418 a_55268_n20136# VV13 0.215f
C1419 R0 S0 3.16f
C1420 frontAnalog_v0p0p1_12.x65.X frontAnalog_v0p0p1_12.RSfetsym_0.x1.Y 0.182f
C1421 w_55000_n67728# VV4 0.798f
C1422 VV2 VV1 4.46f
C1423 a_53630_n14796# VV14 0.28f
C1424 frontAnalog_v0p0p1_6.x65.X I10 0.446f
C1425 w_55000_n52150# frontAnalog_v0p0p1_9.x63.A 0.659f
C1426 a_59578_n29970# VDD 0.0209f
C1427 CLK VV12 0.645f
C1428 frontAnalog_v0p0p1_10.IB a_53630_n63396# 0.473f
C1429 frontAnalog_v0p0p1_4.x63.A a_57123_n20279# 0.212f
C1430 frontAnalog_v0p0p1_14.RSfetsym_0.QN I2 0.0512f
C1431 a_77605_n39305# 16to4_PriorityEncoder_v0p0p1_0.x5.x1.X 0.0991f
C1432 frontAnalog_v0p0p1_8.x63.A VDD 3.67f
C1433 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD 16.6f
C1434 a_53630_n36396# VDD 0.134f
C1435 a_55268_n47136# VIN 0.177f
C1436 16to4_PriorityEncoder_v0p0p1_0.x5.x22.A 16to4_PriorityEncoder_v0p0p1_0.x5.x16.X 0.0732f
C1437 16to4_PriorityEncoder_v0p0p1_0.x3.A1 16to4_PriorityEncoder_v0p0p1_0.x3.x15.X 0.0206f
C1438 frontAnalog_v0p0p1_3.RSfetsym_0.x1.Y VDD 0.733f
C1439 w_55000_n57550# frontAnalog_v0p0p1_10.x65.A 0.0988f
C1440 frontAnalog_v0p0p1_13.RSfetsym_0.QN a_59578_n67770# 0.255f
C1441 a_57123_n61959# CLK 0.0108f
C1442 frontAnalog_v0p0p1_9.x65.X I6 0.446f
C1443 16to4_PriorityEncoder_v0p0p1_0.x5.x22.A 16to4_PriorityEncoder_v0p0p1_0.x5.x21.B 0.064f
C1444 a_53630_n14796# CLK 0.0136f
C1445 w_55000_n40728# frontAnalog_v0p0p1_10.IB 0.0216f
C1446 frontAnalog_v0p0p1_5.x63.X VDD 3.13f
C1447 16to4_PriorityEncoder_v0p0p1_0.x3.EI 16to4_PriorityEncoder_v0p0p1_0.x3.x21.B 0.187f
C1448 frontAnalog_v0p0p1_12.RSfetsym_0.x1.Y frontAnalog_v0p0p1_12.x63.X 0.883f
C1449 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_9.x63.A 0.0926f
C1450 frontAnalog_v0p0p1_6.x63.X I10 1.85f
C1451 w_55000_n8328# w_55000_n8950# 0.327f
C1452 a_78159_n47589# 16to4_PriorityEncoder_v0p0p1_0.x3.x2.X 0.121f
C1453 16to4_PriorityEncoder_v0p0p1_0.x5.x2.X a_77605_n40069# 0.134f
C1454 frontAnalog_v0p0p1_10.x63.A a_55268_n57936# 1.24f
C1455 w_55000_n46128# CLK 0.57f
C1456 frontAnalog_v0p0p1_0.RSfetsym_0.QN frontAnalog_v0p0p1_0.RSfetsym_0.x2.Y 0.018f
C1457 frontAnalog_v0p0p1_11.x65.X frontAnalog_v0p0p1_11.RSfetsym_0.x1.Y 0.182f
C1458 frontAnalog_v0p0p1_4.x65.A frontAnalog_v0p0p1_4.x65.X 0.0236f
C1459 frontAnalog_v0p0p1_13.x63.A VDD 3.67f
C1460 a_53630_n30996# a_55268_n30936# 0.015f
C1461 a_57123_n14879# VDD 0.222f
C1462 frontAnalog_v0p0p1_12.x65.X frontAnalog_v0p0p1_12.RSfetsym_0.QN 2.28f
C1463 a_77605_n48109# VDD 0.154f
C1464 16to4_PriorityEncoder_v0p0p1_0.x3.x11.X I5 0.0201f
C1465 I14 I11 0.782f
C1466 a_55268_n41736# VDD 0.565f
C1467 I13 I12 7.14f
C1468 w_55000_n14350# VDD 0.829f
C1469 w_55000_n78528# a_55268_n79536# 0.149f
C1470 w_55000_n79150# a_53630_n79596# 0.394f
C1471 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD 16.6f
C1472 frontAnalog_v0p0p1_1.x65.A frontAnalog_v0p0p1_1.x65.X 0.0236f
C1473 a_53630_n20196# VIN 0.265f
C1474 16to4_PriorityEncoder_v0p0p1_0.x5.x4.A I9 0.0154f
C1475 frontAnalog_v0p0p1_13.x65.X frontAnalog_v0p0p1_13.x63.X 0.143f
C1476 frontAnalog_v0p0p1_6.RSfetsym_0.x1.Y VDD 0.733f
C1477 frontAnalog_v0p0p1_0.x63.X a_59577_n8883# 0.28f
C1478 16to4_PriorityEncoder_v0p0p1_0.x5.x2.X I15 0.0129f
C1479 frontAnalog_v0p0p1_8.x63.X a_57123_n47279# 0.121f
C1480 frontAnalog_v0p0p1_0.x63.A frontAnalog_v0p0p1_0.x65.A 3.16f
C1481 frontAnalog_v0p0p1_12.x63.X a_57123_n74279# 0.121f
C1482 frontAnalog_v0p0p1_9.x63.X VDD 3.13f
C1483 a_53630_n30996# CLK 0.0136f
C1484 CLK I5 0.0837f
C1485 m3_58396_n25950# VDD 1.25f
C1486 frontAnalog_v0p0p1_3.RSfetsym_0.QN VDD 2.55f
C1487 frontAnalog_v0p0p1_10.RSfetsym_0.QN a_59578_n56970# 0.255f
C1488 16to4_PriorityEncoder_v0p0p1_0.x3.x22.A 16to4_PriorityEncoder_v0p0p1_0.x3.x19.X 0.418f
C1489 frontAnalog_v0p0p1_10.IB a_55268_n74136# 0.0848f
C1490 a_77637_n48817# I4 0.188f
C1491 frontAnalog_v0p0p1_8.RSfetsym_0.QN I8 0.0774f
C1492 frontAnalog_v0p0p1_13.RSfetsym_0.QN frontAnalog_v0p0p1_13.RSfetsym_0.x1.Y 0.17f
C1493 16to4_PriorityEncoder_v0p0p1_0.x3.A1 16to4_PriorityEncoder_v0p0p1_0.x3.x22.A 0.519f
C1494 16to4_PriorityEncoder_v0p0p1_0.x5.x17.A VDD 1.36f
C1495 frontAnalog_v0p0p1_10.IB R0 0.0926f
C1496 a_77637_n41087# VDD 0.307f
C1497 frontAnalog_v0p0p1_11.RSfetsym_0.x1.Y frontAnalog_v0p0p1_11.x63.X 0.883f
C1498 a_77605_n44779# I11 0.15f
C1499 frontAnalog_v0p0p1_0.x63.A CLK 1.8f
C1500 frontAnalog_v0p0p1_12.RSfetsym_0.QN frontAnalog_v0p0p1_12.x63.X 0.378f
C1501 frontAnalog_v0p0p1_12.x65.X frontAnalog_v0p0p1_12.RSfetsym_0.x2.Y 0.526f
C1502 16to4_PriorityEncoder_v0p0p1_0.x29.A VDD 1.52f
C1503 frontAnalog_v0p0p1_12.x65.X CLK 0.443f
C1504 16to4_PriorityEncoder_v0p0p1_0.x5.x22.A 16to4_PriorityEncoder_v0p0p1_0.x5.x15.X 0.209f
C1505 w_55000_n13728# a_53630_n14796# 0.359f
C1506 a_55268_n25536# CLK 0.235f
C1507 frontAnalog_v0p0p1_1.x63.X CLK 0.46f
C1508 16to4_PriorityEncoder_v0p0p1_0.x5.x19.X 16to4_PriorityEncoder_v0p0p1_0.x5.x21.X 0.131f
C1509 a_57123_n31079# VDD 0.222f
C1510 w_55000_n25150# VIN 0.737f
C1511 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_5.x65.A 0.0352f
C1512 w_55000_n79150# frontAnalog_v0p0p1_10.IB 0.0217f
C1513 VIN VV4 3.41f
C1514 frontAnalog_v0p0p1_11.x65.X frontAnalog_v0p0p1_11.RSfetsym_0.QN 2.28f
C1515 16to4_PriorityEncoder_v0p0p1_0.x5.A2 16to4_PriorityEncoder_v0p0p1_0.x1.A 0.38f
C1516 m3_58396_n31350# I10 0.0416f
C1517 w_55000_n41350# a_55268_n41736# 0.12f
C1518 frontAnalog_v0p0p1_13.x65.X I3 0.446f
C1519 frontAnalog_v0p0p1_3.RSfetsym_0.x2.Y VDD 0.926f
C1520 CLK VV6 0.645f
C1521 frontAnalog_v0p0p1_10.x65.X frontAnalog_v0p0p1_10.x63.X 0.143f
C1522 a_78159_n47589# 16to4_PriorityEncoder_v0p0p1_0.x3.x1.X 0.192f
C1523 w_55000_n84550# CLK 0.535f
C1524 frontAnalog_v0p0p1_13.RSfetsym_0.x1.Y frontAnalog_v0p0p1_13.RSfetsym_0.x2.Y 0.0254f
C1525 a_55268_n79536# VDD 0.565f
C1526 frontAnalog_v0p0p1_6.RSfetsym_0.QN VDD 2.55f
C1527 a_59577_n25083# VDD 0.0172f
C1528 frontAnalog_v0p0p1_11.x63.X a_57123_n63479# 0.121f
C1529 16to4_PriorityEncoder_v0p0p1_0.x5.x4.A I13 0.0107f
C1530 frontAnalog_v0p0p1_8.x63.X frontAnalog_v0p0p1_8.RSfetsym_0.x2.Y 0.0923f
C1531 16to4_PriorityEncoder_v0p0p1_0.x3.x19.C I5 0.407f
C1532 frontAnalog_v0p0p1_8.x63.X CLK 0.46f
C1533 frontAnalog_v0p0p1_12.x63.X frontAnalog_v0p0p1_12.RSfetsym_0.x2.Y 0.0923f
C1534 w_55000_n56928# VDD 0.854f
C1535 frontAnalog_v0p0p1_12.x63.X CLK 0.46f
C1536 16to4_PriorityEncoder_v0p0p1_0.x5.x22.A 16to4_PriorityEncoder_v0p0p1_0.x5.x21.X 0.0749f
C1537 frontAnalog_v0p0p1_9.RSfetsym_0.QN frontAnalog_v0p0p1_9.x63.X 0.378f
C1538 frontAnalog_v0p0p1_10.RSfetsym_0.QN frontAnalog_v0p0p1_10.RSfetsym_0.x1.Y 0.17f
C1539 a_59577_n30483# I10 0.29f
C1540 16to4_PriorityEncoder_v0p0p1_0.x36.A VDD 1.52f
C1541 a_77605_n39305# I10 0.216f
C1542 a_53630_n9396# VDD 0.134f
C1543 w_55000_n8950# frontAnalog_v0p0p1_0.x65.A 0.0988f
C1544 frontAnalog_v0p0p1_11.x65.X frontAnalog_v0p0p1_11.RSfetsym_0.x2.Y 0.526f
C1545 frontAnalog_v0p0p1_11.RSfetsym_0.QN frontAnalog_v0p0p1_11.x63.X 0.378f
C1546 VDD I9 5.25f
C1547 w_55000_n3550# frontAnalog_v0p0p1_10.IB 0.0217f
C1548 frontAnalog_v0p0p1_13.x63.X I3 1.85f
C1549 a_78159_n47589# 16to4_PriorityEncoder_v0p0p1_0.x3.EO 0.128f
C1550 a_57123_n63479# CLK 0.0108f
C1551 frontAnalog_v0p0p1_6.RSfetsym_0.x2.Y VDD 0.926f
C1552 w_55000_n8950# CLK 0.535f
C1553 a_77637_n48817# VDD 0.23f
C1554 16to4_PriorityEncoder_v0p0p1_0.x5.x19.X VDD 0.938f
C1555 16to4_PriorityEncoder_v0p0p1_0.x28.A VDD 0.538f
C1556 frontAnalog_v0p0p1_10.RSfetsym_0.x1.Y frontAnalog_v0p0p1_10.RSfetsym_0.x2.Y 0.0254f
C1557 16to4_PriorityEncoder_v0p0p1_0.x5.x2.X I8 0.0265f
C1558 w_55000_n67728# VIN 0.866f
C1559 frontAnalog_v0p0p1_13.RSfetsym_0.QN frontAnalog_v0p0p1_13.RSfetsym_0.x2.Y 0.018f
C1560 16to4_PriorityEncoder_v0p0p1_0.x1.A a_82906_n47995# 0.206f
C1561 frontAnalog_v0p0p1_11.RSfetsym_0.QN CLK 0.0457f
C1562 16to4_PriorityEncoder_v0p0p1_0.x5.x19.D I9 0.937f
C1563 16to4_PriorityEncoder_v0p0p1_0.x2.A 16to4_PriorityEncoder_v0p0p1_0.x3.GS 0.0652f
C1564 m3_58396_n15150# CLK 0.189f
C1565 I1 I0 6.2f
C1566 w_55000_n46128# VV8 0.798f
C1567 frontAnalog_v0p0p1_10.IB VV12 3.87f
C1568 frontAnalog_v0p0p1_11.x63.X frontAnalog_v0p0p1_11.RSfetsym_0.x2.Y 0.0923f
C1569 w_55000_n62328# frontAnalog_v0p0p1_11.x65.A 0.658f
C1570 frontAnalog_v0p0p1_12.RSfetsym_0.QN a_59577_n73683# 0.418f
C1571 frontAnalog_v0p0p1_8.RSfetsym_0.x1.Y I7 0.0436f
C1572 a_57123_n41879# CLK 0.0108f
C1573 16to4_PriorityEncoder_v0p0p1_0.x3.x22.A a_78525_n53555# 0.209f
C1574 frontAnalog_v0p0p1_13.x63.X a_59577_n68283# 0.28f
C1575 frontAnalog_v0p0p1_1.x63.X a_59577_n41283# 0.28f
C1576 16to4_PriorityEncoder_v0p0p1_0.x5.x19.D 16to4_PriorityEncoder_v0p0p1_0.x5.x19.X 0.0195f
C1577 frontAnalog_v0p0p1_7.x65.A VIN 0.655f
C1578 16to4_PriorityEncoder_v0p0p1_0.x5.x22.A VDD 3.25f
C1579 16to4_PriorityEncoder_v0p0p1_0.x3.x18.C I5 0.299f
C1580 w_55000_n84550# S0 0.0988f
C1581 a_53630_n68796# VDD 0.134f
C1582 I4 I1 0.432f
C1583 w_55000_n62950# frontAnalog_v0p0p1_11.x63.A 0.659f
C1584 I7 I0 0.403f
C1585 I5 I6 8.44f
C1586 frontAnalog_v0p0p1_10.IB a_53630_n14796# 0.473f
C1587 a_57123_n34959# VDD 0.222f
C1588 16to4_PriorityEncoder_v0p0p1_0.x5.x4.A a_78159_n39549# 0.299f
C1589 VDD I13 8.01f
C1590 16to4_PriorityEncoder_v0p0p1_0.x35.A VDD 0.539f
C1591 VIN VV11 3.41f
C1592 frontAnalog_v0p0p1_10.x65.A a_57123_n56559# 0.214f
C1593 a_77605_n47345# I1 0.159f
C1594 a_57123_n13359# CLK 0.0108f
C1595 w_55000_n46128# frontAnalog_v0p0p1_10.IB 0.0216f
C1596 a_53630_n36396# VV10 0.28f
C1597 I2 I3 7.24f
C1598 w_55000_n30550# VV11 0.751f
C1599 I7 I4 0.77f
C1600 w_55000_n35328# frontAnalog_v0p0p1_7.x63.A 0.0792f
C1601 frontAnalog_v0p0p1_10.RSfetsym_0.QN frontAnalog_v0p0p1_10.RSfetsym_0.x2.Y 0.018f
C1602 16to4_PriorityEncoder_v0p0p1_0.x5.x19.D 16to4_PriorityEncoder_v0p0p1_0.x5.x22.A 0.0292f
C1603 16to4_PriorityEncoder_v0p0p1_0.x3.EI I0 0.365f
C1604 w_55000_n51528# CLK 0.57f
C1605 frontAnalog_v0p0p1_11.RSfetsym_0.QN a_59577_n62883# 0.418f
C1606 16to4_PriorityEncoder_v0p0p1_0.x5.x19.D I13 0.551f
C1607 a_59578_n2970# I15 0.42f
C1608 CLK VV5 0.645f
C1609 a_78649_n39527# 16to4_PriorityEncoder_v0p0p1_0.x5.EO 0.135f
C1610 w_55000_n46128# frontAnalog_v0p0p1_8.x65.A 0.658f
C1611 a_59578_n35370# VDD 0.0209f
C1612 a_59577_n68283# I3 0.29f
C1613 frontAnalog_v0p0p1_10.x63.X m3_58396_n58350# 0.134f
C1614 16to4_PriorityEncoder_v0p0p1_0.x1.X VDD 0.347f
C1615 frontAnalog_v0p0p1_4.x63.A VDD 3.67f
C1616 a_82906_n51645# VDD 0.18f
C1617 frontAnalog_v0p0p1_10.x63.X a_59577_n57483# 0.28f
C1618 frontAnalog_v0p0p1_1.x65.X VDD 3.46f
C1619 w_55000_n19750# VDD 0.829f
C1620 frontAnalog_v0p0p1_10.IB a_53630_n30996# 0.473f
C1621 frontAnalog_v0p0p1_8.x63.A a_57123_n47279# 0.212f
C1622 16to4_PriorityEncoder_v0p0p1_0.x3.EI I4 1.8f
C1623 w_55000_n46750# frontAnalog_v0p0p1_8.x63.A 0.659f
C1624 w_55000_n79150# VV2 0.751f
C1625 a_57123_n29559# CLK 0.0108f
C1626 frontAnalog_v0p0p1_9.RSfetsym_0.x1.Y frontAnalog_v0p0p1_9.x63.X 0.883f
C1627 m3_58396_n36750# VDD 1.25f
C1628 I15 I10 0.444f
C1629 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_0.x63.A 0.0858f
C1630 frontAnalog_v0p0p1_10.x63.A frontAnalog_v0p0p1_10.x63.X 0.0301f
C1631 VIN S1 0.655f
C1632 16to4_PriorityEncoder_v0p0p1_0.x5.x16.C I9 0.0914f
C1633 frontAnalog_v0p0p1_10.IB a_55268_n25536# 0.0848f
C1634 16to4_PriorityEncoder_v0p0p1_0.x2.A 16to4_PriorityEncoder_v0p0p1_0.x3.EO 0.02f
C1635 a_77637_n42017# VDD 0.322f
C1636 VIN VV15 3.42f
C1637 16to4_PriorityEncoder_v0p0p1_0.x5.x11.X VDD 0.514f
C1638 a_78649_n39527# 16to4_PriorityEncoder_v0p0p1_0.x5.GS 0.136f
C1639 CLK VV16 0.618f
C1640 w_55000_n79150# R1 0.659f
C1641 w_55000_n14350# a_55268_n14736# 0.12f
C1642 frontAnalog_v0p0p1_5.x65.X CLK 0.443f
C1643 16to4_PriorityEncoder_v0p0p1_0.x34.A VDD 0.347f
C1644 frontAnalog_v0p0p1_2.x65.A CLK 2.63f
C1645 frontAnalog_v0p0p1_10.IB VV6 3.88f
C1646 VDD I1 4.6f
C1647 w_55000_n30550# VIN 0.737f
C1648 a_57123_n24159# frontAnalog_v0p0p1_5.x65.X 0.119f
C1649 a_59578_n51570# I6 0.42f
C1650 w_55000_n84550# frontAnalog_v0p0p1_10.IB 0.0217f
C1651 a_78159_n39549# VDD 0.155f
C1652 16to4_PriorityEncoder_v0p0p1_0.x3.x4.A I1 0.0154f
C1653 frontAnalog_v0p0p1_6.x65.A VDD 3.44f
C1654 a_55268_n84936# VIN 0.177f
C1655 frontAnalog_v0p0p1_2.RSfetsym_0.x1.Y I15 0.0432f
C1656 frontAnalog_v0p0p1_7.RSfetsym_0.x1.Y VDD 0.733f
C1657 frontAnalog_v0p0p1_2.x63.A VV16 0.587f
C1658 a_77605_n40069# I14 0.214f
C1659 a_53630_n84996# VV1 0.28f
C1660 frontAnalog_v0p0p1_8.x63.A CLK 1.8f
C1661 frontAnalog_v0p0p1_14.x65.X VDD 3.45f
C1662 16to4_PriorityEncoder_v0p0p1_0.x43.A 16to4_PriorityEncoder_v0p0p1_0.x43.Y 1.52f
C1663 w_55000_n8328# a_53630_n9396# 0.359f
C1664 a_53630_n36396# CLK 0.0136f
C1665 frontAnalog_v0p0p1_2.x63.A frontAnalog_v0p0p1_2.x65.A 3.16f
C1666 VDD I7 4.42f
C1667 w_55000_n62328# VDD 0.854f
C1668 frontAnalog_v0p0p1_5.x63.X CLK 0.46f
C1669 a_55268_n57936# VDD 0.565f
C1670 w_55000_n14350# VV14 0.751f
C1671 a_57123_n7959# VDD 0.222f
C1672 I15 I14 5.72f
C1673 frontAnalog_v0p0p1_5.x65.X a_59578_n24570# 0.436f
C1674 a_53630_n52596# VIN 0.265f
C1675 frontAnalog_v0p0p1_10.x63.A VIN 0.187f
C1676 16to4_PriorityEncoder_v0p0p1_0.x5.x16.C I13 0.415f
C1677 w_55000_n8950# frontAnalog_v0p0p1_10.IB 0.0217f
C1678 a_57123_n36479# VDD 0.222f
C1679 16to4_PriorityEncoder_v0p0p1_0.x3.EI VDD 7.86f
C1680 frontAnalog_v0p0p1_3.x63.X m3_58396_n15150# 0.134f
C1681 16to4_PriorityEncoder_v0p0p1_0.x3.EI a_77605_n51335# 0.122f
C1682 16to4_PriorityEncoder_v0p0p1_0.x3.EI 16to4_PriorityEncoder_v0p0p1_0.x3.x4.A 0.547f
C1683 a_57123_n13359# frontAnalog_v0p0p1_3.x65.X 0.119f
C1684 frontAnalog_v0p0p1_13.x63.A CLK 1.8f
C1685 16to4_PriorityEncoder_v0p0p1_0.x3.A0 16to4_PriorityEncoder_v0p0p1_0.x3.x20.X 0.0149f
C1686 frontAnalog_v0p0p1_14.x63.X VDD 3.13f
C1687 a_57123_n14879# CLK 0.0108f
C1688 a_55268_n41736# CLK 0.235f
C1689 w_55000_n14350# CLK 0.535f
C1690 a_55268_n47136# VDD 0.565f
C1691 frontAnalog_v0p0p1_2.RSfetsym_0.QN I15 2.02f
C1692 w_55000_n62950# a_53630_n63396# 0.394f
C1693 w_55000_n62328# a_55268_n63336# 0.149f
C1694 a_57123_n52679# VDD 0.222f
C1695 frontAnalog_v0p0p1_7.RSfetsym_0.QN VDD 2.55f
C1696 w_55000_n73128# VIN 0.866f
C1697 m3_58396_n79950# I1 0.0416f
C1698 16to4_PriorityEncoder_v0p0p1_0.x5.x14.A 16to4_PriorityEncoder_v0p0p1_0.x5.A2 0.074f
C1699 a_59578_n8370# VDD 0.0209f
C1700 frontAnalog_v0p0p1_9.x63.X CLK 0.46f
C1701 m3_58396_n25950# CLK 0.189f
C1702 I10 I8 2.5f
C1703 frontAnalog_v0p0p1_3.RSfetsym_0.QN CLK 0.0457f
C1704 frontAnalog_v0p0p1_9.RSfetsym_0.QN I7 0.0512f
C1705 w_55000_n24528# frontAnalog_v0p0p1_5.x65.A 0.658f
C1706 w_55000_n51528# w_55000_n52150# 0.327f
C1707 frontAnalog_v0p0p1_12.x63.A VIN 0.187f
C1708 frontAnalog_v0p0p1_3.x65.X a_59578_n13770# 0.436f
C1709 frontAnalog_v0p0p1_5.x65.X frontAnalog_v0p0p1_5.RSfetsym_0.x1.Y 0.182f
C1710 frontAnalog_v0p0p1_2.RSfetsym_0.x2.Y I15 0.194f
C1711 a_57123_n67359# VDD 0.222f
C1712 w_55000_n25150# frontAnalog_v0p0p1_5.x63.A 0.659f
C1713 frontAnalog_v0p0p1_7.RSfetsym_0.x2.Y VDD 0.926f
C1714 a_57123_n31079# CLK 0.0108f
C1715 a_55268_n3936# VIN 0.177f
C1716 a_53630_n20196# VDD 0.134f
C1717 w_55000_n35950# frontAnalog_v0p0p1_7.x65.A 0.0988f
C1718 frontAnalog_v0p0p1_1.RSfetsym_0.QN VDD 2.55f
C1719 16to4_PriorityEncoder_v0p0p1_0.x3.EI 16to4_PriorityEncoder_v0p0p1_0.x3.x16.X 0.076f
C1720 16to4_PriorityEncoder_v0p0p1_0.x2.A 16to4_PriorityEncoder_v0p0p1_0.x21.A 0.0121f
C1721 16to4_PriorityEncoder_v0p0p1_0.x5.x19.C I9 0.347f
C1722 w_55000_n46128# a_53630_n47196# 0.359f
C1723 16to4_PriorityEncoder_v0p0p1_0.x3.x19.D I1 0.937f
C1724 w_55000_n51528# frontAnalog_v0p0p1_10.IB 0.0216f
C1725 frontAnalog_v0p0p1_4.RSfetsym_0.QN a_59578_n19170# 0.255f
C1726 frontAnalog_v0p0p1_9.RSfetsym_0.x2.Y VDD 0.926f
C1727 a_55268_n79536# CLK 0.235f
C1728 frontAnalog_v0p0p1_6.RSfetsym_0.QN CLK 0.0457f
C1729 frontAnalog_v0p0p1_10.IB VV5 3.87f
C1730 frontAnalog_v0p0p1_8.x65.X frontAnalog_v0p0p1_8.RSfetsym_0.x1.Y 0.182f
C1731 a_53630_n41796# a_55268_n41736# 0.015f
C1732 w_55000_n13728# w_55000_n14350# 0.327f
C1733 frontAnalog_v0p0p1_14.x63.X m3_58396_n79950# 0.134f
C1734 VV4 VV3 5.64f
C1735 frontAnalog_v0p0p1_0.RSfetsym_0.x1.Y VDD 0.733f
C1736 frontAnalog_v0p0p1_5.RSfetsym_0.x1.Y frontAnalog_v0p0p1_5.x63.X 0.883f
C1737 m3_58396_n4350# I15 0.0416f
C1738 w_55000_n56928# CLK 0.57f
C1739 frontAnalog_v0p0p1_0.x65.X I14 0.445f
C1740 16to4_PriorityEncoder_v0p0p1_0.x3.EI 16to4_PriorityEncoder_v0p0p1_0.x3.x17.A 0.02f
C1741 16to4_PriorityEncoder_v0p0p1_0.x3.EI a_77637_n49127# 0.0829f
C1742 frontAnalog_v0p0p1_1.x65.A VIN 0.655f
C1743 a_59578_n67770# VDD 0.0209f
C1744 frontAnalog_v0p0p1_0.x63.A a_55268_n9336# 1.24f
C1745 16to4_PriorityEncoder_v0p0p1_0.x3.x19.D I7 0.244f
C1746 frontAnalog_v0p0p1_1.x65.X a_59578_n40770# 0.436f
C1747 a_57123_n29559# frontAnalog_v0p0p1_6.x65.X 0.119f
C1748 a_82906_n47995# 16to4_PriorityEncoder_v0p0p1_0.x3.A1 0.121f
C1749 a_53630_n9396# CLK 0.0136f
C1750 I14 I8 0.358f
C1751 w_55000_n25150# VDD 0.829f
C1752 frontAnalog_v0p0p1_3.x65.X frontAnalog_v0p0p1_3.RSfetsym_0.x1.Y 0.182f
C1753 VDD VV4 1.84f
C1754 a_59577_n79083# VDD 0.0172f
C1755 CLK I9 0.069f
C1756 frontAnalog_v0p0p1_5.x65.X frontAnalog_v0p0p1_5.RSfetsym_0.QN 2.28f
C1757 w_55000_n57550# VV6 0.751f
C1758 frontAnalog_v0p0p1_8.x63.A VV8 0.587f
C1759 frontAnalog_v0p0p1_5.x65.X I11 0.446f
C1760 a_53630_n57996# VV6 0.28f
C1761 frontAnalog_v0p0p1_4.x65.X frontAnalog_v0p0p1_4.x63.X 0.143f
C1762 a_59577_n52083# VDD 0.0172f
C1763 a_59578_n46170# I7 0.42f
C1764 frontAnalog_v0p0p1_10.IB VV16 6.18f
C1765 w_55000_n24528# VV12 0.798f
C1766 a_78097_n45737# 16to4_PriorityEncoder_v0p0p1_0.x5.x20.X 0.137f
C1767 m3_58396_n47550# VDD 1.25f
C1768 16to4_PriorityEncoder_v0p0p1_0.x3.EI a_78649_n47567# 0.181f
C1769 frontAnalog_v0p0p1_13.RSfetsym_0.QN I4 0.0512f
C1770 16to4_PriorityEncoder_v0p0p1_0.x3.EI 16to4_PriorityEncoder_v0p0p1_0.x3.x19.D 1.93f
C1771 a_57123_n9479# VDD 0.222f
C1772 frontAnalog_v0p0p1_5.x63.X a_57123_n25679# 0.121f
C1773 frontAnalog_v0p0p1_0.x63.X I14 1.78f
C1774 w_55000_n73128# frontAnalog_v0p0p1_12.x63.A 0.0792f
C1775 frontAnalog_v0p0p1_2.x65.A frontAnalog_v0p0p1_10.IB 0.0352f
C1776 16to4_PriorityEncoder_v0p0p1_0.x42.A 16to4_PriorityEncoder_v0p0p1_0.x43.A 0.392f
C1777 a_77639_n42341# VDD 0.318f
C1778 16to4_PriorityEncoder_v0p0p1_0.x5.x21.B a_78097_n45737# 0.186f
C1779 frontAnalog_v0p0p1_4.RSfetsym_0.QN frontAnalog_v0p0p1_4.RSfetsym_0.x1.Y 0.17f
C1780 frontAnalog_v0p0p1_6.x65.X a_59578_n29970# 0.436f
C1781 16to4_PriorityEncoder_v0p0p1_0.x5.x19.C I13 0.407f
C1782 a_77605_n43295# 16to4_PriorityEncoder_v0p0p1_0.x5.x16.X 0.0121f
C1783 a_59578_n19170# I12 0.42f
C1784 frontAnalog_v0p0p1_9.RSfetsym_0.QN frontAnalog_v0p0p1_9.RSfetsym_0.x2.Y 0.018f
C1785 a_77605_n52819# I3 0.15f
C1786 frontAnalog_v0p0p1_3.RSfetsym_0.x1.Y frontAnalog_v0p0p1_3.x63.X 0.883f
C1787 16to4_PriorityEncoder_v0p0p1_0.x3.x2.X a_77605_n48109# 0.134f
C1788 a_78065_n41309# 16to4_PriorityEncoder_v0p0p1_0.x5.A2 0.144f
C1789 16to4_PriorityEncoder_v0p0p1_0.x3.EI 16to4_PriorityEncoder_v0p0p1_0.x3.x15.X 0.0245f
C1790 frontAnalog_v0p0p1_5.RSfetsym_0.QN frontAnalog_v0p0p1_5.x63.X 0.378f
C1791 frontAnalog_v0p0p1_0.RSfetsym_0.QN VDD 2.55f
C1792 frontAnalog_v0p0p1_5.x65.X frontAnalog_v0p0p1_5.RSfetsym_0.x2.Y 0.526f
C1793 w_55000_n35950# VIN 0.737f
C1794 frontAnalog_v0p0p1_11.x65.A VIN 0.655f
C1795 16to4_PriorityEncoder_v0p0p1_0.x2.A 16to4_PriorityEncoder_v0p0p1_0.x2.X 0.0402f
C1796 a_77605_n48109# I6 0.214f
C1797 16to4_PriorityEncoder_v0p0p1_0.x5.x18.C I9 0.495f
C1798 frontAnalog_v0p0p1_3.x65.A VIN 0.655f
C1799 frontAnalog_v0p0p1_5.x63.X I11 1.93f
C1800 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_8.x63.A 0.0926f
C1801 frontAnalog_v0p0p1_10.IB a_53630_n36396# 0.473f
C1802 frontAnalog_v0p0p1_13.RSfetsym_0.x1.Y VDD 0.733f
C1803 a_55268_n52536# VV7 0.215f
C1804 frontAnalog_v0p0p1_3.x65.X frontAnalog_v0p0p1_3.RSfetsym_0.QN 2.28f
C1805 frontAnalog_v0p0p1_9.x63.X I6 1.85f
C1806 a_53630_n68796# CLK 0.0136f
C1807 a_57123_n34959# CLK 0.0108f
C1808 w_55000_n8950# a_55268_n9336# 0.12f
C1809 16to4_PriorityEncoder_v0p0p1_0.x3.x16.C I1 0.0914f
C1810 CLK I13 0.0757f
C1811 frontAnalog_v0p0p1_4.RSfetsym_0.x1.Y frontAnalog_v0p0p1_4.RSfetsym_0.x2.Y 0.0254f
C1812 frontAnalog_v0p0p1_8.x63.A frontAnalog_v0p0p1_8.x65.A 3.16f
C1813 16to4_PriorityEncoder_v0p0p1_0.x5.x1.X 16to4_PriorityEncoder_v0p0p1_0.x5.x2.X 0.129f
C1814 w_55000_n67728# VDD 0.854f
C1815 frontAnalog_v0p0p1_9.RSfetsym_0.QN a_59577_n52083# 0.418f
C1816 frontAnalog_v0p0p1_3.x63.X a_57123_n14879# 0.121f
C1817 frontAnalog_v0p0p1_10.x65.X VDD 3.46f
C1818 16to4_PriorityEncoder_v0p0p1_0.x3.x22.A I7 0.0853f
C1819 frontAnalog_v0p0p1_0.RSfetsym_0.x2.Y VDD 0.926f
C1820 frontAnalog_v0p0p1_5.x63.X frontAnalog_v0p0p1_5.RSfetsym_0.x2.Y 0.0923f
C1821 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_13.x63.A 0.0926f
C1822 a_57123_n68879# VDD 0.222f
C1823 frontAnalog_v0p0p1_10.IB a_55268_n41736# 0.0848f
C1824 frontAnalog_v0p0p1_6.x65.X frontAnalog_v0p0p1_6.RSfetsym_0.x1.Y 0.182f
C1825 w_55000_n14350# frontAnalog_v0p0p1_10.IB 0.0217f
C1826 16to4_PriorityEncoder_v0p0p1_0.x3.x16.C I7 0.26f
C1827 frontAnalog_v0p0p1_4.RSfetsym_0.x1.Y I12 0.0436f
C1828 a_53630_n36396# a_55268_n36336# 0.015f
C1829 a_53630_n74196# VIN 0.265f
C1830 m3_58396_n25950# I11 0.0416f
C1831 frontAnalog_v0p0p1_3.RSfetsym_0.QN frontAnalog_v0p0p1_3.x63.X 0.378f
C1832 frontAnalog_v0p0p1_3.x65.X frontAnalog_v0p0p1_3.RSfetsym_0.x2.Y 0.526f
C1833 frontAnalog_v0p0p1_7.x65.A VDD 3.44f
C1834 frontAnalog_v0p0p1_4.x63.A CLK 1.8f
C1835 frontAnalog_v0p0p1_1.x65.X CLK 0.443f
C1836 w_55000_n19750# CLK 0.535f
C1837 frontAnalog_v0p0p1_8.x65.X VDD 3.46f
C1838 16to4_PriorityEncoder_v0p0p1_0.x3.EI 16to4_PriorityEncoder_v0p0p1_0.x3.x22.A 0.0483f
C1839 16to4_PriorityEncoder_v0p0p1_0.x5.x2.X 16to4_PriorityEncoder_v0p0p1_0.x5.EO 0.0749f
C1840 frontAnalog_v0p0p1_13.RSfetsym_0.QN VDD 2.55f
C1841 w_55000_n25150# a_53630_n25596# 0.394f
C1842 w_55000_n24528# a_55268_n25536# 0.149f
C1843 16to4_PriorityEncoder_v0p0p1_0.x5.x18.C I13 0.3f
C1844 w_55000_n78528# S1 0.658f
C1845 a_53630_n79596# a_55268_n79536# 0.015f
C1846 a_77605_n43295# 16to4_PriorityEncoder_v0p0p1_0.x5.x15.X 0.0951f
C1847 VDD VV11 1.84f
C1848 VIN VV9 3.41f
C1849 frontAnalog_v0p0p1_10.x63.X VDD 3.13f
C1850 w_55000_n78528# VIN 0.866f
C1851 16to4_PriorityEncoder_v0p0p1_0.x3.EI 16to4_PriorityEncoder_v0p0p1_0.x3.x16.C 2.08f
C1852 a_59577_n8883# I14 0.29f
C1853 16to4_PriorityEncoder_v0p0p1_0.x5.GS 16to4_PriorityEncoder_v0p0p1_0.x43.A 0.0166f
C1854 m3_58396_n36750# CLK 0.189f
C1855 frontAnalog_v0p0p1_4.RSfetsym_0.QN frontAnalog_v0p0p1_4.RSfetsym_0.x2.Y 0.018f
C1856 frontAnalog_v0p0p1_6.RSfetsym_0.x1.Y frontAnalog_v0p0p1_6.x63.X 0.883f
C1857 frontAnalog_v0p0p1_1.x63.X m3_58396_n42150# 0.134f
C1858 frontAnalog_v0p0p1_3.x63.X frontAnalog_v0p0p1_3.RSfetsym_0.x2.Y 0.0923f
C1859 a_78097_n45737# 16to4_PriorityEncoder_v0p0p1_0.x5.x21.X 0.109f
C1860 VV13 VV12 4.41f
C1861 frontAnalog_v0p0p1_6.x65.A a_55268_n30936# 0.461f
C1862 frontAnalog_v0p0p1_5.x63.A VIN 0.188f
C1863 16to4_PriorityEncoder_v0p0p1_0.x5.x17.A 16to4_PriorityEncoder_v0p0p1_0.x5.A2 0.047f
C1864 frontAnalog_v0p0p1_5.RSfetsym_0.QN a_59577_n25083# 0.418f
C1865 frontAnalog_v0p0p1_6.RSfetsym_0.QN I11 0.0512f
C1866 m3_58396_n74550# I2 0.0416f
C1867 a_59577_n25083# I11 0.29f
C1868 frontAnalog_v0p0p1_1.RSfetsym_0.x1.Y I8 0.0439f
C1869 frontAnalog_v0p0p1_13.x63.A frontAnalog_v0p0p1_13.x65.A 3.16f
C1870 frontAnalog_v0p0p1_4.x63.X a_59577_n19683# 0.28f
C1871 frontAnalog_v0p0p1_13.RSfetsym_0.x2.Y VDD 0.926f
C1872 frontAnalog_v0p0p1_1.RSfetsym_0.QN a_59578_n40770# 0.255f
C1873 frontAnalog_v0p0p1_6.x65.X frontAnalog_v0p0p1_6.RSfetsym_0.QN 2.28f
C1874 frontAnalog_v0p0p1_4.RSfetsym_0.QN I12 2.02f
C1875 CLK I1 0.0837f
C1876 a_57123_n18759# VDD 0.222f
C1877 frontAnalog_v0p0p1_6.x65.A CLK 2.63f
C1878 frontAnalog_v0p0p1_10.IB a_55268_n79536# 0.0848f
C1879 16to4_PriorityEncoder_v0p0p1_0.x2.A 16to4_PriorityEncoder_v0p0p1_0.x3.A0 0.398f
C1880 16to4_PriorityEncoder_v0p0p1_0.x5.x16.X 16to4_PriorityEncoder_v0p0p1_0.x5.x21.B 0.0218f
C1881 16to4_PriorityEncoder_v0p0p1_0.x5.x21.B 16to4_PriorityEncoder_v0p0p1_0.x5.x20.X 0.0561f
C1882 VIN VV3 3.42f
C1883 w_55000_n2928# VIN 0.867f
C1884 w_55000_n46750# a_55268_n47136# 0.12f
C1885 w_55000_n56928# frontAnalog_v0p0p1_10.IB 0.0216f
C1886 frontAnalog_v0p0p1_6.x63.X a_57123_n31079# 0.121f
C1887 frontAnalog_v0p0p1_0.x65.A a_57123_n7959# 0.214f
C1888 I11 I9 1.73f
C1889 frontAnalog_v0p0p1_14.x65.X CLK 0.443f
C1890 frontAnalog_v0p0p1_8.RSfetsym_0.x2.Y I7 0.198f
C1891 frontAnalog_v0p0p1_9.RSfetsym_0.x1.Y frontAnalog_v0p0p1_9.RSfetsym_0.x2.Y 0.0254f
C1892 VDD S1 3.89f
C1893 frontAnalog_v0p0p1_10.IB a_53630_n9396# 0.473f
C1894 CLK I7 0.0837f
C1895 VDD VV15 1.75f
C1896 w_55000_n62328# CLK 0.57f
C1897 w_55000_n73128# a_53630_n74196# 0.359f
C1898 VDD VIN 28.5f
C1899 a_55268_n57936# CLK 0.235f
C1900 frontAnalog_v0p0p1_6.x65.X frontAnalog_v0p0p1_6.RSfetsym_0.x2.Y 0.526f
C1901 frontAnalog_v0p0p1_6.RSfetsym_0.QN frontAnalog_v0p0p1_6.x63.X 0.378f
C1902 frontAnalog_v0p0p1_4.RSfetsym_0.x2.Y I12 0.196f
C1903 a_57123_n7959# CLK 0.0108f
C1904 a_59578_n19170# VDD 0.0209f
C1905 frontAnalog_v0p0p1_3.RSfetsym_0.QN a_59577_n14283# 0.418f
C1906 w_55000_n30550# VDD 0.829f
C1907 frontAnalog_v0p0p1_3.x65.X I13 0.446f
C1908 a_55268_n84936# VDD 0.565f
C1909 a_57123_n36479# CLK 0.0108f
C1910 w_55000_n73750# frontAnalog_v0p0p1_12.x65.A 0.0988f
C1911 frontAnalog_v0p0p1_1.x63.X I8 1.86f
C1912 a_59578_n56970# I5 0.42f
C1913 16to4_PriorityEncoder_v0p0p1_0.x5.GS 16to4_PriorityEncoder_v0p0p1_0.x42.A 0.098f
C1914 a_78097_n45737# VDD 0.332f
C1915 16to4_PriorityEncoder_v0p0p1_0.x3.EI a_78097_n53777# 0.106f
C1916 16to4_PriorityEncoder_v0p0p1_0.x3.x19.C I1 0.347f
C1917 16to4_PriorityEncoder_v0p0p1_0.x3.x21.B VDD 0.721f
C1918 frontAnalog_v0p0p1_14.x63.X CLK 0.46f
C1919 a_59577_n57483# VDD 0.0172f
C1920 m3_58396_n58350# VDD 1.25f
C1921 frontAnalog_v0p0p1_9.x63.A VV7 0.587f
C1922 a_55268_n47136# CLK 0.235f
C1923 w_55000_n40728# frontAnalog_v0p0p1_1.x63.A 0.0792f
C1924 a_55268_n63336# VIN 0.177f
C1925 a_57123_n52679# CLK 0.0108f
C1926 frontAnalog_v0p0p1_7.RSfetsym_0.QN CLK 0.0457f
C1927 a_77605_n43295# VDD 0.551f
C1928 frontAnalog_v0p0p1_0.x63.A frontAnalog_v0p0p1_0.x63.X 0.0301f
C1929 frontAnalog_v0p0p1_6.x63.X frontAnalog_v0p0p1_6.RSfetsym_0.x2.Y 0.0923f
C1930 frontAnalog_v0p0p1_9.x65.A VIN 0.655f
C1931 16to4_PriorityEncoder_v0p0p1_0.x5.x15.X 16to4_PriorityEncoder_v0p0p1_0.x5.x16.X 0.253f
C1932 16to4_PriorityEncoder_v0p0p1_0.x3.x19.C I7 0.239f
C1933 I13 I11 1.27f
C1934 frontAnalog_v0p0p1_3.x63.X I13 1.85f
C1935 a_53630_n52596# VDD 0.134f
C1936 frontAnalog_v0p0p1_10.x63.A VDD 3.67f
C1937 w_55000_n41350# VIN 0.737f
C1938 frontAnalog_v0p0p1_10.IB a_53630_n68796# 0.473f
C1939 16to4_PriorityEncoder_v0p0p1_0.x3.A2 a_78065_n49349# 0.144f
C1940 frontAnalog_v0p0p1_4.RSfetsym_0.x1.Y VDD 0.733f
C1941 frontAnalog_v0p0p1_8.x65.X a_59578_n46170# 0.436f
C1942 w_55000_n73128# VV3 0.798f
C1943 16to4_PriorityEncoder_v0p0p1_0.x3.A2 VDD 1.79f
C1944 16to4_PriorityEncoder_v0p0p1_0.x5.x22.A 16to4_PriorityEncoder_v0p0p1_0.x5.A2 0.0408f
C1945 a_57123_n67359# CLK 0.0108f
C1946 16to4_PriorityEncoder_v0p0p1_0.x3.EI 16to4_PriorityEncoder_v0p0p1_0.x3.x19.C 1.71f
C1947 frontAnalog_v0p0p1_15.RSfetsym_0.QN a_59578_n83970# 0.255f
C1948 a_53630_n20196# CLK 0.0136f
C1949 frontAnalog_v0p0p1_1.RSfetsym_0.QN CLK 0.0457f
C1950 16to4_PriorityEncoder_v0p0p1_0.x5.x2.X I14 0.0177f
C1951 frontAnalog_v0p0p1_10.RSfetsym_0.x1.Y I5 0.0436f
C1952 16to4_PriorityEncoder_v0p0p1_0.x5.EO 16to4_PriorityEncoder_v0p0p1_0.x5.GS 0.927f
C1953 frontAnalog_v0p0p1_12.x63.A VV3 0.587f
C1954 16to4_PriorityEncoder_v0p0p1_0.x5.A2 16to4_PriorityEncoder_v0p0p1_0.x35.A 0.0138f
C1955 16to4_PriorityEncoder_v0p0p1_0.x3.x16.X 16to4_PriorityEncoder_v0p0p1_0.x3.x21.B 0.0218f
C1956 w_55000_n73128# VDD 0.854f
C1957 16to4_PriorityEncoder_v0p0p1_0.x5.x20.X 16to4_PriorityEncoder_v0p0p1_0.x5.x21.X 0.122f
C1958 frontAnalog_v0p0p1_1.x65.A VV9 0.253f
C1959 w_55000_n29928# a_53630_n30996# 0.359f
C1960 16to4_PriorityEncoder_v0p0p1_0.x5.x21.B 16to4_PriorityEncoder_v0p0p1_0.x5.x21.X 0.0197f
C1961 frontAnalog_v0p0p1_15.x65.X I0 0.446f
C1962 16to4_PriorityEncoder_v0p0p1_0.x3.EI a_77637_n50057# 0.0878f
C1963 16to4_PriorityEncoder_v0p0p1_0.x3.x18.C I1 0.495f
C1964 frontAnalog_v0p0p1_12.x63.A VDD 3.67f
C1965 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_4.x63.A 0.0926f
C1966 frontAnalog_v0p0p1_6.RSfetsym_0.QN a_59577_n30483# 0.418f
C1967 w_55000_n3550# a_53630_n3996# 0.394f
C1968 w_55000_n2928# a_55268_n3936# 0.149f
C1969 I6 I1 0.26f
C1970 w_55000_n19750# frontAnalog_v0p0p1_10.IB 0.0217f
C1971 a_57123_n20279# VDD 0.222f
C1972 frontAnalog_v0p0p1_6.x63.A a_57123_n31079# 0.212f
C1973 16to4_PriorityEncoder_v0p0p1_0.x3.EI a_77605_n51585# 0.14f
C1974 a_53630_n25596# VIN 0.265f
C1975 frontAnalog_v0p0p1_15.x65.X frontAnalog_v0p0p1_15.x63.X 0.143f
C1976 16to4_PriorityEncoder_v0p0p1_0.x3.A0 16to4_PriorityEncoder_v0p0p1_0.x3.x19.X 0.0123f
C1977 w_55000_n25150# CLK 0.535f
C1978 a_55268_n3936# VDD 0.565f
C1979 16to4_PriorityEncoder_v0p0p1_0.x3.x2.X I7 0.0129f
C1980 frontAnalog_v0p0p1_9.x63.A a_55268_n52536# 1.24f
C1981 CLK VV4 0.645f
C1982 VDD OUT3 7.1f
C1983 16to4_PriorityEncoder_v0p0p1_0.x3.x18.C I7 0.229f
C1984 frontAnalog_v0p0p1_7.x65.A VV10 0.252f
C1985 frontAnalog_v0p0p1_4.RSfetsym_0.QN VDD 2.55f
C1986 I7 I6 5.92f
C1987 VV1 R0 0.587f
C1988 w_55000_n83928# VIN 0.866f
C1989 a_77605_n39305# I9 0.159f
C1990 frontAnalog_v0p0p1_15.RSfetsym_0.QN frontAnalog_v0p0p1_15.RSfetsym_0.x1.Y 0.17f
C1991 frontAnalog_v0p0p1_15.x63.X I0 1.85f
C1992 a_55268_n79536# VV2 0.215f
C1993 frontAnalog_v0p0p1_10.RSfetsym_0.QN I5 2.02f
C1994 m3_58396_n47550# CLK 0.189f
C1995 frontAnalog_v0p0p1_13.x63.A a_55268_n68736# 1.24f
C1996 VV11 VV10 3.38f
C1997 I5 I3 1.27f
C1998 a_57123_n9479# CLK 0.0108f
C1999 I4 I0 0.575f
C2000 w_55000_n56928# w_55000_n57550# 0.327f
C2001 frontAnalog_v0p0p1_6.x65.A frontAnalog_v0p0p1_6.x65.X 0.0236f
C2002 16to4_PriorityEncoder_v0p0p1_0.x3.x19.D 16to4_PriorityEncoder_v0p0p1_0.x3.x21.B 0.151f
C2003 w_55000_n83928# a_55268_n84936# 0.149f
C2004 w_55000_n84550# a_53630_n84996# 0.394f
C2005 a_59577_n14283# I13 0.29f
C2006 w_55000_n56928# a_53630_n57996# 0.359f
C2007 w_55000_n62950# VV5 0.751f
C2008 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_6.x65.A 0.0352f
C2009 16to4_PriorityEncoder_v0p0p1_0.x3.EI 16to4_PriorityEncoder_v0p0p1_0.x3.x18.C 1.56f
C2010 frontAnalog_v0p0p1_1.x65.A VDD 3.44f
C2011 16to4_PriorityEncoder_v0p0p1_0.x3.EI I6 2.13f
C2012 16to4_PriorityEncoder_v0p0p1_0.x5.x16.X VDD 0.556f
C2013 a_55268_n79536# R1 1.24f
C2014 a_77605_n47345# I0 0.211f
C2015 16to4_PriorityEncoder_v0p0p1_0.x5.x20.X VDD 0.473f
C2016 16to4_PriorityEncoder_v0p0p1_0.x3.A2 16to4_PriorityEncoder_v0p0p1_0.x3.x17.A 0.047f
C2017 a_53630_n9396# a_55268_n9336# 0.015f
C2018 16to4_PriorityEncoder_v0p0p1_0.x5.A2 16to4_PriorityEncoder_v0p0p1_0.x34.A 0.0422f
C2019 a_78349_n43045# 16to4_PriorityEncoder_v0p0p1_0.x1.A 0.151f
C2020 frontAnalog_v0p0p1_0.RSfetsym_0.QN CLK 0.0457f
C2021 frontAnalog_v0p0p1_4.RSfetsym_0.x2.Y VDD 0.926f
C2022 I2 I5 0.649f
C2023 16to4_PriorityEncoder_v0p0p1_0.x3.EI 16to4_PriorityEncoder_v0p0p1_0.x3.GS 0.123f
C2024 16to4_PriorityEncoder_v0p0p1_0.x5.x21.B VDD 0.923f
C2025 16to4_PriorityEncoder_v0p0p1_0.x5.x16.C a_77605_n43295# 0.0949f
C2026 a_55268_n47136# VV8 0.215f
C2027 w_55000_n8328# VV15 0.798f
C2028 frontAnalog_v0p0p1_15.RSfetsym_0.x1.Y frontAnalog_v0p0p1_15.RSfetsym_0.x2.Y 0.0254f
C2029 frontAnalog_v0p0p1_10.RSfetsym_0.x2.Y I5 0.198f
C2030 frontAnalog_v0p0p1_1.RSfetsym_0.x2.Y I8 0.199f
C2031 w_55000_n8328# VIN 0.866f
C2032 w_55000_n62328# frontAnalog_v0p0p1_10.IB 0.0216f
C2033 frontAnalog_v0p0p1_1.RSfetsym_0.QN a_59577_n41283# 0.418f
C2034 frontAnalog_v0p0p1_10.IB a_55268_n57936# 0.0848f
C2035 a_82906_n47995# 16to4_PriorityEncoder_v0p0p1_0.x1.X 0.12f
C2036 frontAnalog_v0p0p1_12.x65.X I2 0.446f
C2037 w_55000_n19128# frontAnalog_v0p0p1_4.x63.A 0.0792f
C2038 a_57123_n40359# frontAnalog_v0p0p1_1.x65.X 0.119f
C2039 VDD I12 5.33f
C2040 frontAnalog_v0p0p1_12.x65.A a_55268_n74136# 0.461f
C2041 w_55000_n19128# w_55000_n19750# 0.327f
C2042 w_55000_n67728# CLK 0.57f
C2043 w_55000_n73750# a_55268_n74136# 0.12f
C2044 16to4_PriorityEncoder_v0p0p1_0.x5.x19.D 16to4_PriorityEncoder_v0p0p1_0.x5.x21.B 0.151f
C2045 frontAnalog_v0p0p1_10.x65.X CLK 0.443f
C2046 frontAnalog_v0p0p1_11.x65.A VDD 3.44f
C2047 w_55000_n35950# VDD 0.829f
C2048 a_57123_n68879# CLK 0.0108f
C2049 frontAnalog_v0p0p1_3.x65.A VDD 3.44f
C2050 VIN VV10 3.42f
C2051 w_55000_n41350# frontAnalog_v0p0p1_1.x65.A 0.0988f
C2052 frontAnalog_v0p0p1_15.x65.X VDD 3.45f
C2053 frontAnalog_v0p0p1_10.IB a_55268_n47136# 0.0848f
C2054 a_55268_n30936# VV11 0.215f
C2055 16to4_PriorityEncoder_v0p0p1_0.x3.EI 16to4_PriorityEncoder_v0p0p1_0.x5.A2 0.507f
C2056 frontAnalog_v0p0p1_8.RSfetsym_0.x1.Y VDD 0.733f
C2057 frontAnalog_v0p0p1_7.x65.A CLK 2.63f
C2058 16to4_PriorityEncoder_v0p0p1_0.x5.x19.D I12 0.206f
C2059 frontAnalog_v0p0p1_8.RSfetsym_0.QN frontAnalog_v0p0p1_8.x63.X 0.378f
C2060 frontAnalog_v0p0p1_8.x65.X frontAnalog_v0p0p1_8.RSfetsym_0.x2.Y 0.526f
C2061 frontAnalog_v0p0p1_12.x63.X I2 1.85f
C2062 m3_58396_n69150# VDD 1.25f
C2063 frontAnalog_v0p0p1_8.x65.X CLK 0.443f
C2064 frontAnalog_v0p0p1_9.RSfetsym_0.x2.Y I6 0.198f
C2065 frontAnalog_v0p0p1_13.RSfetsym_0.QN CLK 0.0457f
C2066 frontAnalog_v0p0p1_15.RSfetsym_0.QN frontAnalog_v0p0p1_15.RSfetsym_0.x2.Y 0.018f
C2067 VDD I0 3.92f
C2068 a_59577_n84483# I0 0.29f
C2069 16to4_PriorityEncoder_v0p0p1_0.x3.x22.A 16to4_PriorityEncoder_v0p0p1_0.x3.x21.B 0.064f
C2070 16to4_PriorityEncoder_v0p0p1_0.x3.A0 a_78525_n53555# 0.149f
C2071 CLK VV11 0.645f
C2072 16to4_PriorityEncoder_v0p0p1_0.x5.x15.X VDD 0.272f
C2073 frontAnalog_v0p0p1_8.x65.A a_55268_n47136# 0.461f
C2074 a_55268_n14736# VIN 0.177f
C2075 frontAnalog_v0p0p1_10.x63.X CLK 0.46f
C2076 a_53630_n74196# VV3 0.28f
C2077 frontAnalog_v0p0p1_7.x65.X I9 0.445f
C2078 frontAnalog_v0p0p1_11.x65.A a_55268_n63336# 0.461f
C2079 16to4_PriorityEncoder_v0p0p1_0.x3.x20.X 16to4_PriorityEncoder_v0p0p1_0.x3.x21.X 0.122f
C2080 frontAnalog_v0p0p1_15.x63.X VDD 3.18f
C2081 a_57123_n51159# VDD 0.222f
C2082 frontAnalog_v0p0p1_15.x63.X a_59577_n84483# 0.28f
C2083 w_55000_n46750# VIN 0.737f
C2084 VDD I4 3.6f
C2085 a_53630_n74196# VDD 0.134f
C2086 frontAnalog_v0p0p1_10.IB a_53630_n20196# 0.473f
C2087 16to4_PriorityEncoder_v0p0p1_0.x5.x4.A VDD 1.92f
C2088 a_78525_n45515# 16to4_PriorityEncoder_v0p0p1_0.x2.A 0.148f
C2089 16to4_PriorityEncoder_v0p0p1_0.x3.EI 16to4_PriorityEncoder_v0p0p1_0.x3.EO 0.187f
C2090 I15 I9 0.29f
C2091 a_57123_n85079# R0 0.223f
C2092 a_59577_n52083# I6 0.29f
C2093 a_77605_n47345# VDD 0.152f
C2094 VV15 VV14 5.48f
C2095 16to4_PriorityEncoder_v0p0p1_0.x3.x4.A a_77605_n47345# 0.0112f
C2096 a_57123_n18759# CLK 0.0108f
C2097 a_82906_n43855# 16to4_PriorityEncoder_v0p0p1_0.x34.A 0.12f
C2098 VIN VV14 3.42f
C2099 16to4_PriorityEncoder_v0p0p1_0.x5.x21.X VDD 0.514f
C2100 frontAnalog_v0p0p1_0.x65.A VV15 0.253f
C2101 frontAnalog_v0p0p1_7.x63.X I9 1.73f
C2102 16to4_PriorityEncoder_v0p0p1_0.x3.A2 16to4_PriorityEncoder_v0p0p1_0.x3.x22.A 0.0408f
C2103 VDD VV9 1.84f
C2104 frontAnalog_v0p0p1_0.x65.A VIN 0.655f
C2105 a_55268_n30936# VIN 0.177f
C2106 w_55000_n78528# VDD 0.854f
C2107 frontAnalog_v0p0p1_2.RSfetsym_0.QN a_59578_n2970# 0.255f
C2108 I14 I10 0.443f
C2109 frontAnalog_v0p0p1_1.x63.A frontAnalog_v0p0p1_1.x63.X 0.0301f
C2110 16to4_PriorityEncoder_v0p0p1_0.x5.x16.C 16to4_PriorityEncoder_v0p0p1_0.x5.x16.X 0.07f
C2111 VV7 VV6 4.01f
C2112 16to4_PriorityEncoder_v0p0p1_0.x5.x19.D 16to4_PriorityEncoder_v0p0p1_0.x5.x4.A 0.0516f
C2113 w_55000_n30550# a_55268_n30936# 0.12f
C2114 a_53630_n68796# a_55268_n68736# 0.015f
C2115 CLK S1 2.64f
C2116 S0 GND 3.47f
C2117 R0 GND 2.53f
C2118 S1 GND 3.81f
C2119 R1 GND 2.55f
C2120 VL GND 0.131p
C2121 VV1 GND 82.8f
C2122 VV2 GND 94.7f
C2123 OUT0 GND 30.2f
C2124 VV3 GND 90.4f
C2125 VV4 GND 86.4f
C2126 VV5 GND 85.2f
C2127 OUT1 GND 30.3f
C2128 I0 GND 50.2f
C2129 I3 GND 51.4f
C2130 I1 GND 59.2f
C2131 I6 GND 34.6f
C2132 I5 GND 42.5f
C2133 I4 GND 44.9f
C2134 I2 GND 56.5f
C2135 I7 GND 30.2f
C2136 VV6 GND 83.7f
C2137 VV7 GND 80.6f
C2138 OUT2 GND 30.2f
C2139 VV8 GND 76.6f
C2140 VV9 GND 74.9f
C2141 OUT3 GND 31.9f
C2142 I8 GND 47.1f
C2143 I9 GND 29.9f
C2144 VV10 GND 77.9f
C2145 I10 GND 36.3f
C2146 VV11 GND 82.6f
C2147 VFS GND 0.114p
C2148 I11 GND 41.4f
C2149 VV12 GND 87.1f
C2150 I12 GND 48.4f
C2151 VV13 GND 88.7f
C2152 I13 GND 59.1f
C2153 VV14 GND 87.8f
C2154 I14 GND 76.8f
C2155 VV15 GND 89.4f
C2156 I15 GND 78.8f
C2157 VV16 GND 89.6f
C2158 VIN GND 0.251p
C2159 CLK GND 0.147p
C2160 VDD GND 3.05p
C2161 m3_58396_n85350# GND 0.227f $ **FLOATING
C2162 m3_58396_n79950# GND 0.157f $ **FLOATING
C2163 m3_58396_n74550# GND 0.157f $ **FLOATING
C2164 m3_58396_n69150# GND 0.157f $ **FLOATING
C2165 m3_58396_n63750# GND 0.157f $ **FLOATING
C2166 m3_58396_n58350# GND 0.157f $ **FLOATING
C2167 m3_58396_n52950# GND 0.157f $ **FLOATING
C2168 m3_58396_n47550# GND 0.157f $ **FLOATING
C2169 m3_58396_n42150# GND 0.157f $ **FLOATING
C2170 m3_58396_n36750# GND 0.157f $ **FLOATING
C2171 m3_58396_n31350# GND 0.157f $ **FLOATING
C2172 m3_58396_n25950# GND 0.157f $ **FLOATING
C2173 m3_58396_n20550# GND 0.157f $ **FLOATING
C2174 m3_58396_n15150# GND 0.157f $ **FLOATING
C2175 m3_58396_n9750# GND 0.157f $ **FLOATING
C2176 m3_58396_n4350# GND 0.157f $ **FLOATING
C2177 a_59577_n84483# GND 0.561f
C2178 a_57123_n85079# GND 0.319f
C2179 frontAnalog_v0p0p1_15.RSfetsym_0.x2.Y GND 1.53f
C2180 frontAnalog_v0p0p1_15.x63.X GND 5.21f
C2181 a_59578_n83970# GND 0.555f
C2182 frontAnalog_v0p0p1_15.RSfetsym_0.x1.Y GND 1.93f
C2183 frontAnalog_v0p0p1_15.RSfetsym_0.QN GND 6.32f
C2184 frontAnalog_v0p0p1_15.x65.X GND 5.08f
C2185 a_57123_n83559# GND 0.318f
C2186 a_55268_n84936# GND 1.17f
C2187 a_53630_n84996# GND 2.61f
C2188 a_59577_n79083# GND 0.561f
C2189 a_57123_n79679# GND 0.319f
C2190 frontAnalog_v0p0p1_14.RSfetsym_0.x2.Y GND 1.53f
C2191 frontAnalog_v0p0p1_14.x63.X GND 5.13f
C2192 a_59578_n78570# GND 0.555f
C2193 frontAnalog_v0p0p1_14.RSfetsym_0.x1.Y GND 1.93f
C2194 frontAnalog_v0p0p1_14.RSfetsym_0.QN GND 6.23f
C2195 frontAnalog_v0p0p1_14.x65.X GND 5.08f
C2196 a_57123_n78159# GND 0.318f
C2197 a_55268_n79536# GND 1.17f
C2198 a_53630_n79596# GND 2.61f
C2199 a_59577_n73683# GND 0.561f
C2200 a_57123_n74279# GND 0.319f
C2201 frontAnalog_v0p0p1_12.RSfetsym_0.x2.Y GND 1.53f
C2202 frontAnalog_v0p0p1_12.x63.X GND 5.13f
C2203 a_59578_n73170# GND 0.555f
C2204 frontAnalog_v0p0p1_12.RSfetsym_0.x1.Y GND 1.93f
C2205 frontAnalog_v0p0p1_12.RSfetsym_0.QN GND 6.23f
C2206 frontAnalog_v0p0p1_12.x65.X GND 5.09f
C2207 a_57123_n72759# GND 0.318f
C2208 a_55268_n74136# GND 1.17f
C2209 a_53630_n74196# GND 2.61f
C2210 frontAnalog_v0p0p1_12.x65.A GND 2.64f
C2211 frontAnalog_v0p0p1_12.x63.A GND 2.48f
C2212 a_59577_n68283# GND 0.561f
C2213 a_57123_n68879# GND 0.319f
C2214 frontAnalog_v0p0p1_13.RSfetsym_0.x2.Y GND 1.53f
C2215 frontAnalog_v0p0p1_13.x63.X GND 5.13f
C2216 a_59578_n67770# GND 0.555f
C2217 frontAnalog_v0p0p1_13.RSfetsym_0.x1.Y GND 1.93f
C2218 frontAnalog_v0p0p1_13.RSfetsym_0.QN GND 6.23f
C2219 frontAnalog_v0p0p1_13.x65.X GND 5.09f
C2220 a_57123_n67359# GND 0.318f
C2221 a_55268_n68736# GND 1.17f
C2222 a_53630_n68796# GND 2.61f
C2223 frontAnalog_v0p0p1_13.x65.A GND 2.64f
C2224 frontAnalog_v0p0p1_13.x63.A GND 2.48f
C2225 a_59577_n62883# GND 0.561f
C2226 a_57123_n63479# GND 0.319f
C2227 frontAnalog_v0p0p1_11.RSfetsym_0.x2.Y GND 1.53f
C2228 frontAnalog_v0p0p1_11.x63.X GND 5.13f
C2229 a_59578_n62370# GND 0.555f
C2230 frontAnalog_v0p0p1_11.RSfetsym_0.x1.Y GND 1.93f
C2231 frontAnalog_v0p0p1_11.RSfetsym_0.QN GND 6.23f
C2232 frontAnalog_v0p0p1_11.x65.X GND 5.09f
C2233 a_57123_n61959# GND 0.318f
C2234 a_55268_n63336# GND 1.17f
C2235 a_53630_n63396# GND 2.61f
C2236 frontAnalog_v0p0p1_11.x65.A GND 2.64f
C2237 frontAnalog_v0p0p1_11.x63.A GND 2.48f
C2238 a_59577_n57483# GND 0.561f
C2239 a_57123_n58079# GND 0.319f
C2240 frontAnalog_v0p0p1_10.RSfetsym_0.x2.Y GND 1.53f
C2241 frontAnalog_v0p0p1_10.x63.X GND 5.13f
C2242 a_59578_n56970# GND 0.555f
C2243 frontAnalog_v0p0p1_10.RSfetsym_0.x1.Y GND 1.93f
C2244 frontAnalog_v0p0p1_10.RSfetsym_0.QN GND 6.23f
C2245 frontAnalog_v0p0p1_10.x65.X GND 5.09f
C2246 a_57123_n56559# GND 0.318f
C2247 a_55268_n57936# GND 1.17f
C2248 a_53630_n57996# GND 2.61f
C2249 frontAnalog_v0p0p1_10.x65.A GND 2.64f
C2250 frontAnalog_v0p0p1_10.x63.A GND 2.47f
C2251 16to4_PriorityEncoder_v0p0p1_0.x3.x21.X GND 0.245f
C2252 16to4_PriorityEncoder_v0p0p1_0.x3.x20.X GND 0.69f
C2253 a_78525_n53555# GND 0.366f
C2254 a_78097_n53777# GND 0.22f
C2255 a_77605_n53805# GND 0.296f
C2256 16to4_PriorityEncoder_v0p0p1_0.x3.x19.X GND 0.443f
C2257 a_77605_n52819# GND 0.295f
C2258 16to4_PriorityEncoder_v0p0p1_0.x3.x21.B GND 0.662f
C2259 a_77605_n52567# GND 0.295f
C2260 a_59577_n52083# GND 0.561f
C2261 16to4_PriorityEncoder_v0p0p1_0.x3.A0 GND 7.55f
C2262 a_57123_n52679# GND 0.319f
C2263 frontAnalog_v0p0p1_9.RSfetsym_0.x2.Y GND 1.53f
C2264 frontAnalog_v0p0p1_9.x63.X GND 5.13f
C2265 a_77605_n51585# GND 0.297f
C2266 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND 9.85f
C2267 16to4_PriorityEncoder_v0p0p1_0.x22.A GND 2.13f
C2268 16to4_PriorityEncoder_v0p0p1_0.x21.A GND 0.663f
C2269 16to4_PriorityEncoder_v0p0p1_0.x2.X GND 0.382f
C2270 a_82906_n51645# GND 0.263f
C2271 a_59578_n51570# GND 0.555f
C2272 16to4_PriorityEncoder_v0p0p1_0.x3.x16.X GND 0.871f
C2273 16to4_PriorityEncoder_v0p0p1_0.x3.x15.X GND 0.334f
C2274 frontAnalog_v0p0p1_9.RSfetsym_0.x1.Y GND 1.93f
C2275 a_78349_n51085# GND 0.369f
C2276 a_77605_n51335# GND 0.296f
C2277 frontAnalog_v0p0p1_9.RSfetsym_0.QN GND 6.23f
C2278 frontAnalog_v0p0p1_9.x65.X GND 5.09f
C2279 a_57123_n51159# GND 0.318f
C2280 a_55268_n52536# GND 1.17f
C2281 a_53630_n52596# GND 2.61f
C2282 a_77639_n50381# GND 0.286f
C2283 frontAnalog_v0p0p1_9.x65.A GND 2.64f
C2284 frontAnalog_v0p0p1_9.x63.A GND 2.48f
C2285 a_77637_n50057# GND 0.288f
C2286 a_78065_n49349# GND 0.367f
C2287 16to4_PriorityEncoder_v0p0p1_0.x3.x17.A GND 0.917f
C2288 16to4_PriorityEncoder_v0p0p1_0.x3.x22.A GND 2.02f
C2289 16to4_PriorityEncoder_v0p0p1_0.x3.x11.X GND 0.263f
C2290 a_77637_n49127# GND 0.28f
C2291 16to4_PriorityEncoder_v0p0p1_0.x3.x14.A GND 0.978f
C2292 a_77637_n48817# GND 0.289f
C2293 16to4_PriorityEncoder_v0p0p1_0.x3.A1 GND 5.12f
C2294 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND 9.86f
C2295 16to4_PriorityEncoder_v0p0p1_0.x29.A GND 2.13f
C2296 16to4_PriorityEncoder_v0p0p1_0.x28.A GND 0.665f
C2297 16to4_PriorityEncoder_v0p0p1_0.x1.X GND 0.383f
C2298 a_82906_n47995# GND 0.265f
C2299 a_77605_n48109# GND 0.388f
C2300 16to4_PriorityEncoder_v0p0p1_0.x3.GS GND 2.06f
C2301 16to4_PriorityEncoder_v0p0p1_0.x3.EO GND 2.32f
C2302 16to4_PriorityEncoder_v0p0p1_0.x3.x2.X GND 0.676f
C2303 16to4_PriorityEncoder_v0p0p1_0.x3.x1.X GND 0.162f
C2304 a_78649_n47567# GND 0.258f
C2305 a_78159_n47589# GND 0.343f
C2306 a_77605_n47345# GND 0.379f
C2307 16to4_PriorityEncoder_v0p0p1_0.x3.x4.A GND 1.07f
C2308 16to4_PriorityEncoder_v0p0p1_0.x3.x19.D GND 4.1f
C2309 16to4_PriorityEncoder_v0p0p1_0.x3.x16.C GND 1.84f
C2310 16to4_PriorityEncoder_v0p0p1_0.x3.x19.C GND 4.41f
C2311 16to4_PriorityEncoder_v0p0p1_0.x3.x18.C GND 1.88f
C2312 a_59577_n46683# GND 0.561f
C2313 a_57123_n47279# GND 0.319f
C2314 frontAnalog_v0p0p1_8.RSfetsym_0.x2.Y GND 1.53f
C2315 frontAnalog_v0p0p1_8.x63.X GND 5.13f
C2316 a_59578_n46170# GND 0.555f
C2317 16to4_PriorityEncoder_v0p0p1_0.x2.A GND 6.65f
C2318 16to4_PriorityEncoder_v0p0p1_0.x5.x21.X GND 0.242f
C2319 16to4_PriorityEncoder_v0p0p1_0.x5.x20.X GND 0.684f
C2320 frontAnalog_v0p0p1_8.RSfetsym_0.x1.Y GND 1.93f
C2321 a_78525_n45515# GND 0.364f
C2322 a_78097_n45737# GND 0.217f
C2323 a_77605_n45765# GND 0.291f
C2324 frontAnalog_v0p0p1_8.RSfetsym_0.QN GND 6.21f
C2325 frontAnalog_v0p0p1_8.x65.X GND 5.04f
C2326 a_57123_n45759# GND 0.318f
C2327 a_55268_n47136# GND 1.17f
C2328 a_53630_n47196# GND 2.61f
C2329 16to4_PriorityEncoder_v0p0p1_0.x5.x19.X GND 0.434f
C2330 frontAnalog_v0p0p1_8.x65.A GND 2.64f
C2331 frontAnalog_v0p0p1_8.x63.A GND 2.48f
C2332 a_77605_n44779# GND 0.293f
C2333 16to4_PriorityEncoder_v0p0p1_0.x5.x21.B GND 0.652f
C2334 a_77605_n44527# GND 0.295f
C2335 16to4_PriorityEncoder_v0p0p1_0.x3.A2 GND 7.64f
C2336 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND 9.83f
C2337 16to4_PriorityEncoder_v0p0p1_0.x36.A GND 2.12f
C2338 16to4_PriorityEncoder_v0p0p1_0.x35.A GND 0.662f
C2339 16to4_PriorityEncoder_v0p0p1_0.x34.A GND 0.379f
C2340 a_82906_n43855# GND 0.263f
C2341 a_77605_n43545# GND 0.297f
C2342 16to4_PriorityEncoder_v0p0p1_0.x1.A GND 5.67f
C2343 16to4_PriorityEncoder_v0p0p1_0.x5.x16.X GND 0.871f
C2344 16to4_PriorityEncoder_v0p0p1_0.x5.x15.X GND 0.334f
C2345 a_78349_n43045# GND 0.369f
C2346 a_77605_n43295# GND 0.296f
C2347 a_77639_n42341# GND 0.286f
C2348 a_77637_n42017# GND 0.288f
C2349 16to4_PriorityEncoder_v0p0p1_0.x5.A2 GND 5.29f
C2350 a_78065_n41309# GND 0.367f
C2351 16to4_PriorityEncoder_v0p0p1_0.x5.x17.A GND 0.876f
C2352 16to4_PriorityEncoder_v0p0p1_0.x5.x22.A GND 1.77f
C2353 16to4_PriorityEncoder_v0p0p1_0.x5.x11.X GND 0.263f
C2354 a_77637_n41087# GND 0.28f
C2355 a_59577_n41283# GND 0.561f
C2356 a_57123_n41879# GND 0.319f
C2357 frontAnalog_v0p0p1_1.RSfetsym_0.x2.Y GND 1.51f
C2358 frontAnalog_v0p0p1_1.x63.X GND 5.12f
C2359 16to4_PriorityEncoder_v0p0p1_0.x5.x14.A GND 0.958f
C2360 a_59578_n40770# GND 0.555f
C2361 a_77637_n40777# GND 0.289f
C2362 frontAnalog_v0p0p1_1.RSfetsym_0.x1.Y GND 1.92f
C2363 16to4_PriorityEncoder_v0p0p1_0.x3.EI GND 18.6f
C2364 frontAnalog_v0p0p1_1.RSfetsym_0.QN GND 6.3f
C2365 a_77605_n40069# GND 0.391f
C2366 frontAnalog_v0p0p1_1.x65.X GND 5.01f
C2367 a_57123_n40359# GND 0.318f
C2368 a_55268_n41736# GND 1.17f
C2369 a_53630_n41796# GND 2.61f
C2370 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND 9.88f
C2371 16to4_PriorityEncoder_v0p0p1_0.x43.A GND 2.02f
C2372 16to4_PriorityEncoder_v0p0p1_0.x42.A GND 0.633f
C2373 16to4_PriorityEncoder_v0p0p1_0.x5.GS GND 2.51f
C2374 frontAnalog_v0p0p1_1.x65.A GND 2.64f
C2375 frontAnalog_v0p0p1_1.x63.A GND 2.47f
C2376 16to4_PriorityEncoder_v0p0p1_0.x5.EO GND 2.62f
C2377 16to4_PriorityEncoder_v0p0p1_0.x5.x2.X GND 0.684f
C2378 16to4_PriorityEncoder_v0p0p1_0.x5.x1.X GND 0.167f
C2379 a_78649_n39527# GND 0.262f
C2380 a_78159_n39549# GND 0.347f
C2381 a_77605_n39305# GND 0.384f
C2382 16to4_PriorityEncoder_v0p0p1_0.x5.x4.A GND 1.5f
C2383 16to4_PriorityEncoder_v0p0p1_0.x5.x19.D GND 4.1f
C2384 16to4_PriorityEncoder_v0p0p1_0.x5.x16.C GND 1.85f
C2385 16to4_PriorityEncoder_v0p0p1_0.x5.x19.C GND 4.42f
C2386 16to4_PriorityEncoder_v0p0p1_0.x5.x18.C GND 1.89f
C2387 a_59577_n35883# GND 0.561f
C2388 a_57123_n36479# GND 0.319f
C2389 frontAnalog_v0p0p1_7.RSfetsym_0.x2.Y GND 1.54f
C2390 frontAnalog_v0p0p1_7.x63.X GND 5.21f
C2391 a_59578_n35370# GND 0.555f
C2392 frontAnalog_v0p0p1_7.RSfetsym_0.x1.Y GND 1.93f
C2393 frontAnalog_v0p0p1_7.RSfetsym_0.QN GND 6.3f
C2394 frontAnalog_v0p0p1_7.x65.X GND 5.09f
C2395 a_57123_n34959# GND 0.318f
C2396 a_55268_n36336# GND 1.17f
C2397 a_53630_n36396# GND 2.61f
C2398 frontAnalog_v0p0p1_7.x65.A GND 2.64f
C2399 frontAnalog_v0p0p1_7.x63.A GND 2.48f
C2400 a_59577_n30483# GND 0.561f
C2401 a_57123_n31079# GND 0.319f
C2402 frontAnalog_v0p0p1_6.RSfetsym_0.x2.Y GND 1.53f
C2403 frontAnalog_v0p0p1_6.x63.X GND 5.15f
C2404 a_59578_n29970# GND 0.555f
C2405 frontAnalog_v0p0p1_6.RSfetsym_0.x1.Y GND 1.93f
C2406 frontAnalog_v0p0p1_6.RSfetsym_0.QN GND 6.23f
C2407 frontAnalog_v0p0p1_6.x65.X GND 5.09f
C2408 a_57123_n29559# GND 0.318f
C2409 a_55268_n30936# GND 1.17f
C2410 a_53630_n30996# GND 2.61f
C2411 frontAnalog_v0p0p1_6.x65.A GND 2.64f
C2412 frontAnalog_v0p0p1_6.x63.A GND 2.48f
C2413 a_59577_n25083# GND 0.561f
C2414 a_57123_n25679# GND 0.319f
C2415 frontAnalog_v0p0p1_5.RSfetsym_0.x2.Y GND 1.53f
C2416 frontAnalog_v0p0p1_5.x63.X GND 5.11f
C2417 a_59578_n24570# GND 0.555f
C2418 frontAnalog_v0p0p1_5.RSfetsym_0.x1.Y GND 1.93f
C2419 frontAnalog_v0p0p1_5.RSfetsym_0.QN GND 6.3f
C2420 frontAnalog_v0p0p1_5.x65.X GND 5.09f
C2421 a_57123_n24159# GND 0.318f
C2422 a_55268_n25536# GND 1.17f
C2423 a_53630_n25596# GND 2.61f
C2424 frontAnalog_v0p0p1_5.x65.A GND 2.64f
C2425 frontAnalog_v0p0p1_5.x63.A GND 2.48f
C2426 a_59577_n19683# GND 0.561f
C2427 a_57123_n20279# GND 0.319f
C2428 frontAnalog_v0p0p1_4.RSfetsym_0.x2.Y GND 1.53f
C2429 frontAnalog_v0p0p1_4.x63.X GND 5.15f
C2430 a_59578_n19170# GND 0.555f
C2431 frontAnalog_v0p0p1_4.RSfetsym_0.x1.Y GND 1.93f
C2432 frontAnalog_v0p0p1_4.RSfetsym_0.QN GND 6.3f
C2433 frontAnalog_v0p0p1_4.x65.X GND 5.09f
C2434 a_57123_n18759# GND 0.318f
C2435 a_55268_n20136# GND 1.17f
C2436 a_53630_n20196# GND 2.61f
C2437 frontAnalog_v0p0p1_4.x65.A GND 2.64f
C2438 frontAnalog_v0p0p1_4.x63.A GND 2.47f
C2439 a_59577_n14283# GND 0.561f
C2440 a_57123_n14879# GND 0.319f
C2441 frontAnalog_v0p0p1_3.RSfetsym_0.x2.Y GND 1.53f
C2442 frontAnalog_v0p0p1_3.x63.X GND 5.15f
C2443 a_59578_n13770# GND 0.555f
C2444 frontAnalog_v0p0p1_3.RSfetsym_0.x1.Y GND 1.93f
C2445 frontAnalog_v0p0p1_3.RSfetsym_0.QN GND 6.23f
C2446 frontAnalog_v0p0p1_3.x65.X GND 5.09f
C2447 a_57123_n13359# GND 0.318f
C2448 a_55268_n14736# GND 1.17f
C2449 a_53630_n14796# GND 2.61f
C2450 frontAnalog_v0p0p1_3.x65.A GND 2.64f
C2451 frontAnalog_v0p0p1_3.x63.A GND 2.47f
C2452 a_59577_n8883# GND 0.561f
C2453 a_57123_n9479# GND 0.319f
C2454 frontAnalog_v0p0p1_0.RSfetsym_0.x2.Y GND 1.54f
C2455 frontAnalog_v0p0p1_0.x63.X GND 5.16f
C2456 a_59578_n8370# GND 0.555f
C2457 frontAnalog_v0p0p1_0.RSfetsym_0.x1.Y GND 1.93f
C2458 frontAnalog_v0p0p1_0.RSfetsym_0.QN GND 6.23f
C2459 frontAnalog_v0p0p1_0.x65.X GND 5.09f
C2460 a_57123_n7959# GND 0.318f
C2461 a_55268_n9336# GND 1.17f
C2462 a_53630_n9396# GND 2.61f
C2463 frontAnalog_v0p0p1_0.x65.A GND 2.64f
C2464 frontAnalog_v0p0p1_0.x63.A GND 2.47f
C2465 a_59577_n3483# GND 0.561f
C2466 a_57123_n4079# GND 0.319f
C2467 frontAnalog_v0p0p1_2.RSfetsym_0.x2.Y GND 1.54f
C2468 frontAnalog_v0p0p1_2.x63.X GND 5.16f
C2469 a_59578_n2970# GND 0.555f
C2470 frontAnalog_v0p0p1_2.RSfetsym_0.x1.Y GND 1.93f
C2471 frontAnalog_v0p0p1_2.RSfetsym_0.QN GND 6.3f
C2472 frontAnalog_v0p0p1_2.x65.X GND 5.01f
C2473 a_57123_n2559# GND 0.318f
C2474 a_55268_n3936# GND 1.17f
C2475 a_53630_n3996# GND 2.61f
C2476 frontAnalog_v0p0p1_10.IB GND 0.389p
C2477 frontAnalog_v0p0p1_2.x65.A GND 2.64f
C2478 frontAnalog_v0p0p1_2.x63.A GND 2.46f
C2479 w_55000_n84550# GND 2.69f
C2480 w_55000_n83928# GND 2.69f
C2481 w_55000_n79150# GND 2.69f
C2482 w_55000_n78528# GND 2.69f
C2483 w_55000_n73750# GND 2.69f
C2484 w_55000_n73128# GND 2.69f
C2485 w_55000_n68350# GND 2.69f
C2486 w_55000_n67728# GND 2.69f
C2487 w_55000_n62950# GND 2.69f
C2488 w_55000_n62328# GND 2.69f
C2489 w_55000_n57550# GND 2.69f
C2490 w_55000_n56928# GND 2.69f
C2491 w_55000_n52150# GND 2.69f
C2492 w_55000_n51528# GND 2.69f
C2493 w_55000_n46750# GND 2.69f
C2494 w_55000_n46128# GND 2.69f
C2495 w_55000_n41350# GND 2.69f
C2496 w_55000_n40728# GND 2.69f
C2497 w_55000_n35950# GND 2.69f
C2498 w_55000_n35328# GND 2.69f
C2499 w_55000_n30550# GND 2.69f
C2500 w_55000_n29928# GND 2.69f
C2501 w_55000_n25150# GND 2.69f
C2502 w_55000_n24528# GND 2.69f
C2503 w_55000_n19750# GND 2.69f
C2504 w_55000_n19128# GND 2.68f
C2505 w_55000_n14350# GND 2.69f
C2506 w_55000_n13728# GND 2.69f
C2507 w_55000_n8950# GND 2.69f
C2508 w_55000_n8328# GND 2.69f
C2509 w_55000_n3550# GND 2.69f
C2510 w_55000_n2928# GND 2.68f
C2511 frontAnalog_v0p0p1_0.x63.A.n0 GND 0.12f
C2512 frontAnalog_v0p0p1_0.x63.A.n1 GND 2.22f
C2513 frontAnalog_v0p0p1_0.x63.A.t6 GND 0.014f
C2514 frontAnalog_v0p0p1_0.x63.A.t5 GND 0.0225f
C2515 frontAnalog_v0p0p1_0.x63.A.n2 GND 0.0465f
C2516 frontAnalog_v0p0p1_0.x63.A.t4 GND 0.0256f
C2517 frontAnalog_v0p0p1_0.x63.A.t1 GND 0.173f
C2518 frontAnalog_v0p0p1_0.x63.A.t7 GND 0.175f
C2519 frontAnalog_v0p0p1_0.x63.A.n3 GND 1f
C2520 frontAnalog_v0p0p1_0.x63.A.n4 GND 0.953f
C2521 frontAnalog_v0p0p1_0.x63.A.t2 GND 0.0156f
C2522 frontAnalog_v0p0p1_0.x63.A.t3 GND 0.335f
C2523 frontAnalog_v0p0p1_0.x63.A.t0 GND 0.151f
C2524 frontAnalog_v0p0p1_0.x63.A.n5 GND 1.25f
C2525 frontAnalog_v0p0p1_0.x65.A.n0 GND 0.139f
C2526 frontAnalog_v0p0p1_0.x65.A.t5 GND 0.028f
C2527 frontAnalog_v0p0p1_0.x65.A.t6 GND 0.0175f
C2528 frontAnalog_v0p0p1_0.x65.A.n1 GND 0.0568f
C2529 frontAnalog_v0p0p1_0.x65.A.t1 GND 0.149f
C2530 frontAnalog_v0p0p1_0.x65.A.t2 GND 0.463f
C2531 frontAnalog_v0p0p1_0.x65.A.t3 GND 0.0194f
C2532 frontAnalog_v0p0p1_0.x65.A.n2 GND 1.6f
C2533 frontAnalog_v0p0p1_0.x65.A.t7 GND 0.0318f
C2534 frontAnalog_v0p0p1_0.x65.A.t0 GND 0.141f
C2535 frontAnalog_v0p0p1_0.x65.A.t4 GND 0.219f
C2536 frontAnalog_v0p0p1_0.x65.A.n3 GND 1.37f
C2537 frontAnalog_v0p0p1_0.x65.A.n4 GND 0.898f
C2538 frontAnalog_v0p0p1_0.x65.A.n5 GND 2.01f
C2539 frontAnalog_v0p0p1_0.x65.A.n6 GND 1.72f
C2540 frontAnalog_v0p0p1_6.x65.A.n0 GND 0.139f
C2541 frontAnalog_v0p0p1_6.x65.A.t6 GND 0.028f
C2542 frontAnalog_v0p0p1_6.x65.A.t7 GND 0.0175f
C2543 frontAnalog_v0p0p1_6.x65.A.n1 GND 0.0568f
C2544 frontAnalog_v0p0p1_6.x65.A.t1 GND 0.149f
C2545 frontAnalog_v0p0p1_6.x65.A.t3 GND 0.463f
C2546 frontAnalog_v0p0p1_6.x65.A.t2 GND 0.0194f
C2547 frontAnalog_v0p0p1_6.x65.A.n2 GND 1.6f
C2548 frontAnalog_v0p0p1_6.x65.A.t5 GND 0.0318f
C2549 frontAnalog_v0p0p1_6.x65.A.t0 GND 0.141f
C2550 frontAnalog_v0p0p1_6.x65.A.t4 GND 0.219f
C2551 frontAnalog_v0p0p1_6.x65.A.n3 GND 1.37f
C2552 frontAnalog_v0p0p1_6.x65.A.n4 GND 0.898f
C2553 frontAnalog_v0p0p1_6.x65.A.n5 GND 2.01f
C2554 frontAnalog_v0p0p1_6.x65.A.n6 GND 1.72f
C2555 frontAnalog_v0p0p1_12.x65.A.n0 GND 0.139f
C2556 frontAnalog_v0p0p1_12.x65.A.t4 GND 0.028f
C2557 frontAnalog_v0p0p1_12.x65.A.t6 GND 0.0175f
C2558 frontAnalog_v0p0p1_12.x65.A.n1 GND 0.0568f
C2559 frontAnalog_v0p0p1_12.x65.A.t2 GND 0.149f
C2560 frontAnalog_v0p0p1_12.x65.A.t7 GND 0.0318f
C2561 frontAnalog_v0p0p1_12.x65.A.t3 GND 0.141f
C2562 frontAnalog_v0p0p1_12.x65.A.t5 GND 0.219f
C2563 frontAnalog_v0p0p1_12.x65.A.n2 GND 1.37f
C2564 frontAnalog_v0p0p1_12.x65.A.n3 GND 0.898f
C2565 frontAnalog_v0p0p1_12.x65.A.t1 GND 0.463f
C2566 frontAnalog_v0p0p1_12.x65.A.t0 GND 0.0194f
C2567 frontAnalog_v0p0p1_12.x65.A.n4 GND 1.6f
C2568 frontAnalog_v0p0p1_12.x65.A.n5 GND 2.01f
C2569 frontAnalog_v0p0p1_12.x65.A.n6 GND 1.72f
C2570 frontAnalog_v0p0p1_2.RSfetsym_0.QN.n0 GND 0.993f
C2571 frontAnalog_v0p0p1_2.RSfetsym_0.QN.t5 GND 0.0317f
C2572 frontAnalog_v0p0p1_2.RSfetsym_0.QN.t6 GND 0.0933f
C2573 frontAnalog_v0p0p1_2.RSfetsym_0.QN.n1 GND 1.47f
C2574 frontAnalog_v0p0p1_2.RSfetsym_0.QN.n2 GND 0.587f
C2575 frontAnalog_v0p0p1_2.RSfetsym_0.QN.t1 GND 0.0363f
C2576 frontAnalog_v0p0p1_2.RSfetsym_0.QN.n3 GND 0.622f
C2577 frontAnalog_v0p0p1_2.RSfetsym_0.QN.t3 GND 0.0317f
C2578 frontAnalog_v0p0p1_2.RSfetsym_0.QN.t4 GND 0.0317f
C2579 frontAnalog_v0p0p1_2.RSfetsym_0.QN.t0 GND 0.0558f
C2580 frontAnalog_v0p0p1_8.x63.A.n0 GND 0.12f
C2581 frontAnalog_v0p0p1_8.x63.A.n1 GND 2.22f
C2582 frontAnalog_v0p0p1_8.x63.A.t7 GND 0.014f
C2583 frontAnalog_v0p0p1_8.x63.A.t5 GND 0.0225f
C2584 frontAnalog_v0p0p1_8.x63.A.n2 GND 0.0465f
C2585 frontAnalog_v0p0p1_8.x63.A.t6 GND 0.0256f
C2586 frontAnalog_v0p0p1_8.x63.A.t1 GND 0.173f
C2587 frontAnalog_v0p0p1_8.x63.A.t4 GND 0.175f
C2588 frontAnalog_v0p0p1_8.x63.A.n3 GND 1f
C2589 frontAnalog_v0p0p1_8.x63.A.n4 GND 0.953f
C2590 frontAnalog_v0p0p1_8.x63.A.t2 GND 0.0156f
C2591 frontAnalog_v0p0p1_8.x63.A.t3 GND 0.335f
C2592 frontAnalog_v0p0p1_8.x63.A.t0 GND 0.151f
C2593 frontAnalog_v0p0p1_8.x63.A.n5 GND 1.25f
C2594 I11.n2 GND 0.538f
C2595 I11.n3 GND 0.0114f
C2596 I11.n5 GND 0.965f
C2597 I11.n6 GND 0.443f
C2598 I11.n7 GND 0.551f
C2599 I11.n8 GND 0.145f
C2600 I11.n9 GND 0.9f
C2601 I11.t8 GND 0.0195f
C2602 I11.n10 GND 0.306f
C2603 I11.n11 GND 0.0405f
C2604 I11.n12 GND 0.0919f
C2605 I11.n13 GND 0.061f
C2606 I11.n14 GND 0.0652f
C2607 I11.n15 GND 0.0898f
C2608 I11.n16 GND 0.085f
C2609 I11.n17 GND 0.205f
C2610 I11.n18 GND 8.8f
C2611 I11.n19 GND 1.02f
C2612 frontAnalog_v0p0p1_1.RSfetsym_0.QN.n0 GND 0.993f
C2613 frontAnalog_v0p0p1_1.RSfetsym_0.QN.t6 GND 0.0317f
C2614 frontAnalog_v0p0p1_1.RSfetsym_0.QN.t5 GND 0.0933f
C2615 frontAnalog_v0p0p1_1.RSfetsym_0.QN.n1 GND 1.47f
C2616 frontAnalog_v0p0p1_1.RSfetsym_0.QN.n2 GND 0.587f
C2617 frontAnalog_v0p0p1_1.RSfetsym_0.QN.t4 GND 0.0363f
C2618 frontAnalog_v0p0p1_1.RSfetsym_0.QN.n3 GND 0.622f
C2619 frontAnalog_v0p0p1_1.RSfetsym_0.QN.t3 GND 0.0317f
C2620 frontAnalog_v0p0p1_1.RSfetsym_0.QN.t2 GND 0.0317f
C2621 frontAnalog_v0p0p1_1.RSfetsym_0.QN.t0 GND 0.0558f
C2622 I3.n2 GND 0.411f
C2623 I3.n5 GND 0.717f
C2624 I3.n6 GND 0.337f
C2625 I3.n7 GND 0.528f
C2626 I3.t8 GND 0.0146f
C2627 I3.n8 GND 0.23f
C2628 I3.n9 GND 0.0304f
C2629 I3.n10 GND 0.0689f
C2630 I3.n11 GND 0.0457f
C2631 I3.n12 GND 0.0489f
C2632 I3.n13 GND 0.0674f
C2633 I3.n14 GND 0.0637f
C2634 I3.n15 GND 0.147f
C2635 I3.n16 GND 8.52f
C2636 I3.n17 GND 0.845f
C2637 I15.n8 GND 0.134f
C2638 I15.n9 GND 0.29f
C2639 I15.n10 GND 0.12f
C2640 I15.n11 GND 0.167f
C2641 I15.n12 GND 0.0609f
C2642 I15.n13 GND 0.184f
C2643 I15.n14 GND 0.129f
C2644 I15.n15 GND 0.0171f
C2645 I15.n16 GND 0.0387f
C2646 I15.n17 GND 0.0257f
C2647 I15.n18 GND 0.0275f
C2648 I15.n19 GND 0.0379f
C2649 I15.n20 GND 0.0358f
C2650 I15.n21 GND 0.0936f
C2651 I15.n22 GND 0.309f
C2652 I14.n10 GND 0.0646f
C2653 I14.n11 GND 0.157f
C2654 I14.n14 GND 0.0845f
C2655 I14.n21 GND 0.203f
C2656 I14.n22 GND 0.338f
C2657 I14.n23 GND 0.202f
C2658 I14.n24 GND 0.348f
C2659 I14.n25 GND 0.111f
C2660 I14.n26 GND 0.423f
C2661 I14.t8 GND 0.015f
C2662 I14.n27 GND 0.234f
C2663 I14.n28 GND 0.031f
C2664 I14.n29 GND 0.0704f
C2665 I14.n30 GND 0.0467f
C2666 I14.n31 GND 0.0499f
C2667 I14.n32 GND 0.0688f
C2668 I14.n33 GND 0.0651f
C2669 I14.n34 GND 0.17f
C2670 I14.n35 GND 0.778f
C2671 frontAnalog_v0p0p1_8.x65.A.n0 GND 0.139f
C2672 frontAnalog_v0p0p1_8.x65.A.t4 GND 0.028f
C2673 frontAnalog_v0p0p1_8.x65.A.t6 GND 0.0175f
C2674 frontAnalog_v0p0p1_8.x65.A.n1 GND 0.0568f
C2675 frontAnalog_v0p0p1_8.x65.A.t1 GND 0.149f
C2676 frontAnalog_v0p0p1_8.x65.A.t2 GND 0.463f
C2677 frontAnalog_v0p0p1_8.x65.A.t3 GND 0.0194f
C2678 frontAnalog_v0p0p1_8.x65.A.n2 GND 1.6f
C2679 frontAnalog_v0p0p1_8.x65.A.t7 GND 0.0318f
C2680 frontAnalog_v0p0p1_8.x65.A.t0 GND 0.141f
C2681 frontAnalog_v0p0p1_8.x65.A.t5 GND 0.219f
C2682 frontAnalog_v0p0p1_8.x65.A.n3 GND 1.37f
C2683 frontAnalog_v0p0p1_8.x65.A.n4 GND 0.898f
C2684 frontAnalog_v0p0p1_8.x65.A.n5 GND 2.01f
C2685 frontAnalog_v0p0p1_8.x65.A.n6 GND 1.72f
C2686 frontAnalog_v0p0p1_11.x63.A.n0 GND 0.12f
C2687 frontAnalog_v0p0p1_11.x63.A.n1 GND 2.22f
C2688 frontAnalog_v0p0p1_11.x63.A.t7 GND 0.014f
C2689 frontAnalog_v0p0p1_11.x63.A.t5 GND 0.0225f
C2690 frontAnalog_v0p0p1_11.x63.A.n2 GND 0.0465f
C2691 frontAnalog_v0p0p1_11.x63.A.t1 GND 0.151f
C2692 frontAnalog_v0p0p1_11.x63.A.t2 GND 0.0156f
C2693 frontAnalog_v0p0p1_11.x63.A.t3 GND 0.335f
C2694 frontAnalog_v0p0p1_11.x63.A.t6 GND 0.0256f
C2695 frontAnalog_v0p0p1_11.x63.A.t0 GND 0.173f
C2696 frontAnalog_v0p0p1_11.x63.A.t4 GND 0.175f
C2697 frontAnalog_v0p0p1_11.x63.A.n3 GND 1f
C2698 frontAnalog_v0p0p1_11.x63.A.n4 GND 0.953f
C2699 frontAnalog_v0p0p1_11.x63.A.n5 GND 1.25f
C2700 I7.n0 GND 0.0133f
C2701 I7.n4 GND 0.0124f
C2702 I7.n8 GND 0.484f
C2703 I7.n9 GND 1.04f
C2704 I7.n10 GND 0.441f
C2705 I7.n11 GND 1.73f
C2706 I7.t9 GND 0.0298f
C2707 I7.n12 GND 0.467f
C2708 I7.n13 GND 0.0619f
C2709 I7.t0 GND 0.01f
C2710 I7.n14 GND 0.14f
C2711 I7.n15 GND 0.093f
C2712 I7.n16 GND 0.0995f
C2713 I7.n17 GND 0.137f
C2714 I7.n18 GND 0.13f
C2715 I7.t4 GND 0.011f
C2716 I7.n19 GND 0.299f
C2717 I7.n20 GND 4.39f
C2718 I7.n21 GND 2.56f
C2719 frontAnalog_v0p0p1_4.RSfetsym_0.QN.n0 GND 0.993f
C2720 frontAnalog_v0p0p1_4.RSfetsym_0.QN.t6 GND 0.0317f
C2721 frontAnalog_v0p0p1_4.RSfetsym_0.QN.t5 GND 0.0933f
C2722 frontAnalog_v0p0p1_4.RSfetsym_0.QN.n1 GND 1.47f
C2723 frontAnalog_v0p0p1_4.RSfetsym_0.QN.n2 GND 0.587f
C2724 frontAnalog_v0p0p1_4.RSfetsym_0.QN.t4 GND 0.0363f
C2725 frontAnalog_v0p0p1_4.RSfetsym_0.QN.n3 GND 0.622f
C2726 frontAnalog_v0p0p1_4.RSfetsym_0.QN.t1 GND 0.0317f
C2727 frontAnalog_v0p0p1_4.RSfetsym_0.QN.t2 GND 0.0317f
C2728 frontAnalog_v0p0p1_4.RSfetsym_0.QN.t3 GND 0.0558f
C2729 frontAnalog_v0p0p1_12.x63.A.n0 GND 0.12f
C2730 frontAnalog_v0p0p1_12.x63.A.n1 GND 2.22f
C2731 frontAnalog_v0p0p1_12.x63.A.t6 GND 0.014f
C2732 frontAnalog_v0p0p1_12.x63.A.t4 GND 0.0225f
C2733 frontAnalog_v0p0p1_12.x63.A.n2 GND 0.0465f
C2734 frontAnalog_v0p0p1_12.x63.A.t5 GND 0.0256f
C2735 frontAnalog_v0p0p1_12.x63.A.t1 GND 0.173f
C2736 frontAnalog_v0p0p1_12.x63.A.t7 GND 0.175f
C2737 frontAnalog_v0p0p1_12.x63.A.n3 GND 1f
C2738 frontAnalog_v0p0p1_12.x63.A.n4 GND 0.953f
C2739 frontAnalog_v0p0p1_12.x63.A.t3 GND 0.0156f
C2740 frontAnalog_v0p0p1_12.x63.A.t2 GND 0.335f
C2741 frontAnalog_v0p0p1_12.x63.A.t0 GND 0.151f
C2742 frontAnalog_v0p0p1_12.x63.A.n5 GND 1.25f
C2743 frontAnalog_v0p0p1_11.RSfetsym_0.QN.n0 GND 0.993f
C2744 frontAnalog_v0p0p1_11.RSfetsym_0.QN.t6 GND 0.0317f
C2745 frontAnalog_v0p0p1_11.RSfetsym_0.QN.t5 GND 0.0933f
C2746 frontAnalog_v0p0p1_11.RSfetsym_0.QN.n1 GND 1.47f
C2747 frontAnalog_v0p0p1_11.RSfetsym_0.QN.n2 GND 0.587f
C2748 frontAnalog_v0p0p1_11.RSfetsym_0.QN.t0 GND 0.0363f
C2749 frontAnalog_v0p0p1_11.RSfetsym_0.QN.n3 GND 0.622f
C2750 frontAnalog_v0p0p1_11.RSfetsym_0.QN.t2 GND 0.0317f
C2751 frontAnalog_v0p0p1_11.RSfetsym_0.QN.t3 GND 0.0317f
C2752 frontAnalog_v0p0p1_11.RSfetsym_0.QN.t1 GND 0.0558f
C2753 frontAnalog_v0p0p1_13.x65.A.n0 GND 0.139f
C2754 frontAnalog_v0p0p1_13.x65.A.t4 GND 0.028f
C2755 frontAnalog_v0p0p1_13.x65.A.t6 GND 0.0175f
C2756 frontAnalog_v0p0p1_13.x65.A.n1 GND 0.0568f
C2757 frontAnalog_v0p0p1_13.x65.A.t2 GND 0.149f
C2758 frontAnalog_v0p0p1_13.x65.A.t7 GND 0.0318f
C2759 frontAnalog_v0p0p1_13.x65.A.t3 GND 0.141f
C2760 frontAnalog_v0p0p1_13.x65.A.t5 GND 0.219f
C2761 frontAnalog_v0p0p1_13.x65.A.n2 GND 1.37f
C2762 frontAnalog_v0p0p1_13.x65.A.n3 GND 0.898f
C2763 frontAnalog_v0p0p1_13.x65.A.t0 GND 0.463f
C2764 frontAnalog_v0p0p1_13.x65.A.t1 GND 0.0194f
C2765 frontAnalog_v0p0p1_13.x65.A.n4 GND 1.6f
C2766 frontAnalog_v0p0p1_13.x65.A.n5 GND 2.01f
C2767 frontAnalog_v0p0p1_13.x65.A.n6 GND 1.72f
C2768 I8.n1 GND 0.123f
C2769 I8.n2 GND 0.318f
C2770 I8.n3 GND 2.5f
C2771 I8.t5 GND 0.0121f
C2772 I8.n4 GND 0.189f
C2773 I8.n5 GND 0.0251f
C2774 I8.n6 GND 0.0568f
C2775 I8.n7 GND 0.0377f
C2776 I8.n8 GND 0.0403f
C2777 I8.n9 GND 0.0556f
C2778 I8.n10 GND 0.0526f
C2779 I8.n11 GND 0.137f
C2780 frontAnalog_v0p0p1_0.RSfetsym_0.QN.n0 GND 0.993f
C2781 frontAnalog_v0p0p1_0.RSfetsym_0.QN.t5 GND 0.0317f
C2782 frontAnalog_v0p0p1_0.RSfetsym_0.QN.t6 GND 0.0933f
C2783 frontAnalog_v0p0p1_0.RSfetsym_0.QN.n1 GND 1.47f
C2784 frontAnalog_v0p0p1_0.RSfetsym_0.QN.n2 GND 0.587f
C2785 frontAnalog_v0p0p1_0.RSfetsym_0.QN.t3 GND 0.0363f
C2786 frontAnalog_v0p0p1_0.RSfetsym_0.QN.n3 GND 0.622f
C2787 frontAnalog_v0p0p1_0.RSfetsym_0.QN.t1 GND 0.0317f
C2788 frontAnalog_v0p0p1_0.RSfetsym_0.QN.t0 GND 0.0317f
C2789 frontAnalog_v0p0p1_0.RSfetsym_0.QN.t4 GND 0.0558f
C2790 frontAnalog_v0p0p1_7.RSfetsym_0.QN.n0 GND 0.993f
C2791 frontAnalog_v0p0p1_7.RSfetsym_0.QN.t6 GND 0.0317f
C2792 frontAnalog_v0p0p1_7.RSfetsym_0.QN.t5 GND 0.0933f
C2793 frontAnalog_v0p0p1_7.RSfetsym_0.QN.n1 GND 1.47f
C2794 frontAnalog_v0p0p1_7.RSfetsym_0.QN.n2 GND 0.587f
C2795 frontAnalog_v0p0p1_7.RSfetsym_0.QN.t0 GND 0.0363f
C2796 frontAnalog_v0p0p1_7.RSfetsym_0.QN.n3 GND 0.622f
C2797 frontAnalog_v0p0p1_7.RSfetsym_0.QN.t3 GND 0.0317f
C2798 frontAnalog_v0p0p1_7.RSfetsym_0.QN.t4 GND 0.0317f
C2799 frontAnalog_v0p0p1_7.RSfetsym_0.QN.t1 GND 0.0558f
C2800 frontAnalog_v0p0p1_14.RSfetsym_0.QN.n0 GND 0.993f
C2801 frontAnalog_v0p0p1_14.RSfetsym_0.QN.t6 GND 0.0317f
C2802 frontAnalog_v0p0p1_14.RSfetsym_0.QN.t5 GND 0.0933f
C2803 frontAnalog_v0p0p1_14.RSfetsym_0.QN.n1 GND 1.47f
C2804 frontAnalog_v0p0p1_14.RSfetsym_0.QN.n2 GND 0.587f
C2805 frontAnalog_v0p0p1_14.RSfetsym_0.QN.t1 GND 0.0363f
C2806 frontAnalog_v0p0p1_14.RSfetsym_0.QN.n3 GND 0.622f
C2807 frontAnalog_v0p0p1_14.RSfetsym_0.QN.t3 GND 0.0317f
C2808 frontAnalog_v0p0p1_14.RSfetsym_0.QN.t4 GND 0.0317f
C2809 frontAnalog_v0p0p1_14.RSfetsym_0.QN.t0 GND 0.0558f
C2810 frontAnalog_v0p0p1_5.x65.A.n0 GND 0.139f
C2811 frontAnalog_v0p0p1_5.x65.A.t4 GND 0.028f
C2812 frontAnalog_v0p0p1_5.x65.A.t6 GND 0.0175f
C2813 frontAnalog_v0p0p1_5.x65.A.n1 GND 0.0568f
C2814 frontAnalog_v0p0p1_5.x65.A.t1 GND 0.149f
C2815 frontAnalog_v0p0p1_5.x65.A.t3 GND 0.463f
C2816 frontAnalog_v0p0p1_5.x65.A.t2 GND 0.0194f
C2817 frontAnalog_v0p0p1_5.x65.A.n2 GND 1.6f
C2818 frontAnalog_v0p0p1_5.x65.A.t7 GND 0.0318f
C2819 frontAnalog_v0p0p1_5.x65.A.t0 GND 0.141f
C2820 frontAnalog_v0p0p1_5.x65.A.t5 GND 0.219f
C2821 frontAnalog_v0p0p1_5.x65.A.n3 GND 1.37f
C2822 frontAnalog_v0p0p1_5.x65.A.n4 GND 0.898f
C2823 frontAnalog_v0p0p1_5.x65.A.n5 GND 2.01f
C2824 frontAnalog_v0p0p1_5.x65.A.n6 GND 1.72f
C2825 frontAnalog_v0p0p1_1.x63.A.n0 GND 0.12f
C2826 frontAnalog_v0p0p1_1.x63.A.n1 GND 2.22f
C2827 frontAnalog_v0p0p1_1.x63.A.t6 GND 0.014f
C2828 frontAnalog_v0p0p1_1.x63.A.t7 GND 0.0225f
C2829 frontAnalog_v0p0p1_1.x63.A.n2 GND 0.0465f
C2830 frontAnalog_v0p0p1_1.x63.A.t3 GND 0.151f
C2831 frontAnalog_v0p0p1_1.x63.A.t4 GND 0.0256f
C2832 frontAnalog_v0p0p1_1.x63.A.t2 GND 0.173f
C2833 frontAnalog_v0p0p1_1.x63.A.t5 GND 0.175f
C2834 frontAnalog_v0p0p1_1.x63.A.n3 GND 1f
C2835 frontAnalog_v0p0p1_1.x63.A.n4 GND 0.953f
C2836 frontAnalog_v0p0p1_1.x63.A.t0 GND 0.0156f
C2837 frontAnalog_v0p0p1_1.x63.A.t1 GND 0.334f
C2838 frontAnalog_v0p0p1_1.x63.A.n5 GND 1.25f
C2839 I12.n6 GND 0.144f
C2840 I12.n8 GND 0.0234f
C2841 I12.n9 GND 0.253f
C2842 I12.n11 GND 0.11f
C2843 I12.n12 GND 0.235f
C2844 I12.n13 GND 0.31f
C2845 I12.n14 GND 0.459f
C2846 I12.n15 GND 0.13f
C2847 I12.n16 GND 0.69f
C2848 I12.t7 GND 0.0176f
C2849 I12.n17 GND 0.275f
C2850 I12.n18 GND 0.0365f
C2851 I12.n19 GND 0.0827f
C2852 I12.n20 GND 0.0549f
C2853 I12.n21 GND 0.0587f
C2854 I12.n22 GND 0.0808f
C2855 I12.n23 GND 0.0765f
C2856 I12.n24 GND 0.184f
C2857 I12.n25 GND 9.69f
C2858 I12.n26 GND 1.15f
C2859 VV8.t16 GND 0.0135f
C2860 VV8.n0 GND 0.111f
C2861 VV8.n1 GND 0.0535f
C2862 VV8.t4 GND 0.176f
C2863 VV8.t14 GND 0.176f
C2864 VV8.t15 GND 0.176f
C2865 VV8.t0 GND 0.176f
C2866 VV8.t10 GND 0.176f
C2867 VV8.t11 GND 0.176f
C2868 VV8.t8 GND 0.176f
C2869 VV8.t3 GND 0.176f
C2870 VV8.t1 GND 0.176f
C2871 VV8.t12 GND 0.176f
C2872 VV8.t7 GND 0.176f
C2873 VV8.t6 GND 0.176f
C2874 VV8.t5 GND 0.176f
C2875 VV8.t9 GND 0.176f
C2876 VV8.t2 GND 0.176f
C2877 VV8.t13 GND 0.176f
C2878 VV8.n2 GND 0.422f
C2879 VV8.n3 GND 0.433f
C2880 VV8.n4 GND 0.433f
C2881 VV8.n5 GND 0.433f
C2882 VV8.n6 GND 0.433f
C2883 VV8.n7 GND 0.433f
C2884 VV8.n8 GND 0.433f
C2885 VV8.n9 GND 0.387f
C2886 VV8.n10 GND 0.921f
C2887 frontAnalog_v0p0p1_11.x65.A.n0 GND 0.139f
C2888 frontAnalog_v0p0p1_11.x65.A.t4 GND 0.028f
C2889 frontAnalog_v0p0p1_11.x65.A.t6 GND 0.0175f
C2890 frontAnalog_v0p0p1_11.x65.A.n1 GND 0.0568f
C2891 frontAnalog_v0p0p1_11.x65.A.t7 GND 0.0318f
C2892 frontAnalog_v0p0p1_11.x65.A.t1 GND 0.141f
C2893 frontAnalog_v0p0p1_11.x65.A.t5 GND 0.219f
C2894 frontAnalog_v0p0p1_11.x65.A.n2 GND 1.37f
C2895 frontAnalog_v0p0p1_11.x65.A.n3 GND 0.898f
C2896 frontAnalog_v0p0p1_11.x65.A.t3 GND 0.463f
C2897 frontAnalog_v0p0p1_11.x65.A.t2 GND 0.0194f
C2898 frontAnalog_v0p0p1_11.x65.A.n4 GND 1.6f
C2899 frontAnalog_v0p0p1_11.x65.A.n5 GND 2.01f
C2900 frontAnalog_v0p0p1_11.x65.A.t0 GND 0.149f
C2901 frontAnalog_v0p0p1_11.x65.A.n6 GND 1.72f
C2902 frontAnalog_v0p0p1_12.RSfetsym_0.QN.n0 GND 0.993f
C2903 frontAnalog_v0p0p1_12.RSfetsym_0.QN.t6 GND 0.0317f
C2904 frontAnalog_v0p0p1_12.RSfetsym_0.QN.t5 GND 0.0933f
C2905 frontAnalog_v0p0p1_12.RSfetsym_0.QN.n1 GND 1.47f
C2906 frontAnalog_v0p0p1_12.RSfetsym_0.QN.n2 GND 0.587f
C2907 frontAnalog_v0p0p1_12.RSfetsym_0.QN.t4 GND 0.0363f
C2908 frontAnalog_v0p0p1_12.RSfetsym_0.QN.n3 GND 0.622f
C2909 frontAnalog_v0p0p1_12.RSfetsym_0.QN.t2 GND 0.0317f
C2910 frontAnalog_v0p0p1_12.RSfetsym_0.QN.t1 GND 0.0317f
C2911 frontAnalog_v0p0p1_12.RSfetsym_0.QN.t3 GND 0.0558f
C2912 frontAnalog_v0p0p1_6.x63.A.n0 GND 0.12f
C2913 frontAnalog_v0p0p1_6.x63.A.n1 GND 2.22f
C2914 frontAnalog_v0p0p1_6.x63.A.t6 GND 0.014f
C2915 frontAnalog_v0p0p1_6.x63.A.t4 GND 0.0225f
C2916 frontAnalog_v0p0p1_6.x63.A.n2 GND 0.0465f
C2917 frontAnalog_v0p0p1_6.x63.A.t2 GND 0.151f
C2918 frontAnalog_v0p0p1_6.x63.A.t7 GND 0.0256f
C2919 frontAnalog_v0p0p1_6.x63.A.t3 GND 0.173f
C2920 frontAnalog_v0p0p1_6.x63.A.t5 GND 0.175f
C2921 frontAnalog_v0p0p1_6.x63.A.n3 GND 1f
C2922 frontAnalog_v0p0p1_6.x63.A.n4 GND 0.953f
C2923 frontAnalog_v0p0p1_6.x63.A.t1 GND 0.0156f
C2924 frontAnalog_v0p0p1_6.x63.A.t0 GND 0.334f
C2925 frontAnalog_v0p0p1_6.x63.A.n5 GND 1.25f
C2926 frontAnalog_v0p0p1_3.RSfetsym_0.QN.n0 GND 0.993f
C2927 frontAnalog_v0p0p1_3.RSfetsym_0.QN.t6 GND 0.0317f
C2928 frontAnalog_v0p0p1_3.RSfetsym_0.QN.t5 GND 0.0933f
C2929 frontAnalog_v0p0p1_3.RSfetsym_0.QN.n1 GND 1.47f
C2930 frontAnalog_v0p0p1_3.RSfetsym_0.QN.n2 GND 0.587f
C2931 frontAnalog_v0p0p1_3.RSfetsym_0.QN.t0 GND 0.0363f
C2932 frontAnalog_v0p0p1_3.RSfetsym_0.QN.n3 GND 0.622f
C2933 frontAnalog_v0p0p1_3.RSfetsym_0.QN.t1 GND 0.0317f
C2934 frontAnalog_v0p0p1_3.RSfetsym_0.QN.t2 GND 0.0317f
C2935 frontAnalog_v0p0p1_3.RSfetsym_0.QN.t4 GND 0.0558f
C2936 I4.n6 GND 0.16f
C2937 I4.n8 GND 0.026f
C2938 I4.n9 GND 0.282f
C2939 I4.n11 GND 0.123f
C2940 I4.n12 GND 0.262f
C2941 I4.n13 GND 0.361f
C2942 I4.n14 GND 0.813f
C2943 I4.t12 GND 0.0196f
C2944 I4.n15 GND 0.307f
C2945 I4.n16 GND 0.0406f
C2946 I4.n17 GND 0.0921f
C2947 I4.n18 GND 0.0611f
C2948 I4.n19 GND 0.0654f
C2949 I4.n20 GND 0.09f
C2950 I4.n21 GND 0.0852f
C2951 I4.n22 GND 0.196f
C2952 I4.n23 GND 9.38f
C2953 I4.n24 GND 1.33f
C2954 frontAnalog_v0p0p1_10.RSfetsym_0.QN.n0 GND 0.993f
C2955 frontAnalog_v0p0p1_10.RSfetsym_0.QN.t6 GND 0.0317f
C2956 frontAnalog_v0p0p1_10.RSfetsym_0.QN.t5 GND 0.0933f
C2957 frontAnalog_v0p0p1_10.RSfetsym_0.QN.n1 GND 1.47f
C2958 frontAnalog_v0p0p1_10.RSfetsym_0.QN.n2 GND 0.587f
C2959 frontAnalog_v0p0p1_10.RSfetsym_0.QN.t4 GND 0.0363f
C2960 frontAnalog_v0p0p1_10.RSfetsym_0.QN.n3 GND 0.622f
C2961 frontAnalog_v0p0p1_10.RSfetsym_0.QN.t2 GND 0.0317f
C2962 frontAnalog_v0p0p1_10.RSfetsym_0.QN.t3 GND 0.0317f
C2963 frontAnalog_v0p0p1_10.RSfetsym_0.QN.t0 GND 0.0558f
C2964 frontAnalog_v0p0p1_1.x65.A.n0 GND 0.139f
C2965 frontAnalog_v0p0p1_1.x65.A.t4 GND 0.028f
C2966 frontAnalog_v0p0p1_1.x65.A.t6 GND 0.0175f
C2967 frontAnalog_v0p0p1_1.x65.A.n1 GND 0.0568f
C2968 frontAnalog_v0p0p1_1.x65.A.t7 GND 0.0318f
C2969 frontAnalog_v0p0p1_1.x65.A.t1 GND 0.141f
C2970 frontAnalog_v0p0p1_1.x65.A.t5 GND 0.219f
C2971 frontAnalog_v0p0p1_1.x65.A.n2 GND 1.37f
C2972 frontAnalog_v0p0p1_1.x65.A.n3 GND 0.898f
C2973 frontAnalog_v0p0p1_1.x65.A.t3 GND 0.463f
C2974 frontAnalog_v0p0p1_1.x65.A.t2 GND 0.0194f
C2975 frontAnalog_v0p0p1_1.x65.A.n4 GND 1.6f
C2976 frontAnalog_v0p0p1_1.x65.A.n5 GND 2.01f
C2977 frontAnalog_v0p0p1_1.x65.A.t0 GND 0.149f
C2978 frontAnalog_v0p0p1_1.x65.A.n6 GND 1.72f
C2979 frontAnalog_v0p0p1_4.x63.A.n0 GND 0.12f
C2980 frontAnalog_v0p0p1_4.x63.A.n1 GND 2.22f
C2981 frontAnalog_v0p0p1_4.x63.A.t5 GND 0.014f
C2982 frontAnalog_v0p0p1_4.x63.A.t6 GND 0.0225f
C2983 frontAnalog_v0p0p1_4.x63.A.n2 GND 0.0465f
C2984 frontAnalog_v0p0p1_4.x63.A.t2 GND 0.151f
C2985 frontAnalog_v0p0p1_4.x63.A.t4 GND 0.0256f
C2986 frontAnalog_v0p0p1_4.x63.A.t3 GND 0.173f
C2987 frontAnalog_v0p0p1_4.x63.A.t7 GND 0.175f
C2988 frontAnalog_v0p0p1_4.x63.A.n3 GND 1f
C2989 frontAnalog_v0p0p1_4.x63.A.n4 GND 0.953f
C2990 frontAnalog_v0p0p1_4.x63.A.t0 GND 0.0156f
C2991 frontAnalog_v0p0p1_4.x63.A.t1 GND 0.334f
C2992 frontAnalog_v0p0p1_4.x63.A.n5 GND 1.25f
C2993 S0.t2 GND 0.144f
C2994 S0.t4 GND 0.0271f
C2995 S0.t6 GND 0.0169f
C2996 S0.n0 GND 0.0551f
C2997 S0.n1 GND 0.0448f
C2998 S0.n2 GND 0.0338f
C2999 S0.n3 GND 0.175f
C3000 S0.n5 GND 0.627f
C3001 S0.t7 GND 0.0309f
C3002 S0.t3 GND 0.137f
C3003 S0.t5 GND 0.213f
C3004 S0.n6 GND 1.33f
C3005 S0.n7 GND 0.871f
C3006 S0.t1 GND 0.449f
C3007 S0.t0 GND 0.0188f
C3008 S0.n8 GND 1.55f
C3009 S0.n9 GND 1.93f
C3010 S0.n10 GND 0.661f
C3011 S0.n11 GND 0.207f
C3012 frontAnalog_v0p0p1_3.x65.A.n0 GND 0.139f
C3013 frontAnalog_v0p0p1_3.x65.A.t4 GND 0.028f
C3014 frontAnalog_v0p0p1_3.x65.A.t6 GND 0.0175f
C3015 frontAnalog_v0p0p1_3.x65.A.n1 GND 0.0568f
C3016 frontAnalog_v0p0p1_3.x65.A.t1 GND 0.149f
C3017 frontAnalog_v0p0p1_3.x65.A.t3 GND 0.463f
C3018 frontAnalog_v0p0p1_3.x65.A.t2 GND 0.0194f
C3019 frontAnalog_v0p0p1_3.x65.A.n2 GND 1.6f
C3020 frontAnalog_v0p0p1_3.x65.A.t7 GND 0.0318f
C3021 frontAnalog_v0p0p1_3.x65.A.t0 GND 0.141f
C3022 frontAnalog_v0p0p1_3.x65.A.t5 GND 0.219f
C3023 frontAnalog_v0p0p1_3.x65.A.n3 GND 1.37f
C3024 frontAnalog_v0p0p1_3.x65.A.n4 GND 0.898f
C3025 frontAnalog_v0p0p1_3.x65.A.n5 GND 2.01f
C3026 frontAnalog_v0p0p1_3.x65.A.n6 GND 1.72f
C3027 frontAnalog_v0p0p1_3.x63.A.n0 GND 0.12f
C3028 frontAnalog_v0p0p1_3.x63.A.n1 GND 2.22f
C3029 frontAnalog_v0p0p1_3.x63.A.t7 GND 0.014f
C3030 frontAnalog_v0p0p1_3.x63.A.t5 GND 0.0225f
C3031 frontAnalog_v0p0p1_3.x63.A.n2 GND 0.0465f
C3032 frontAnalog_v0p0p1_3.x63.A.t6 GND 0.0256f
C3033 frontAnalog_v0p0p1_3.x63.A.t1 GND 0.173f
C3034 frontAnalog_v0p0p1_3.x63.A.t4 GND 0.175f
C3035 frontAnalog_v0p0p1_3.x63.A.n3 GND 1f
C3036 frontAnalog_v0p0p1_3.x63.A.n4 GND 0.953f
C3037 frontAnalog_v0p0p1_3.x63.A.t3 GND 0.0156f
C3038 frontAnalog_v0p0p1_3.x63.A.t2 GND 0.335f
C3039 frontAnalog_v0p0p1_3.x63.A.t0 GND 0.151f
C3040 frontAnalog_v0p0p1_3.x63.A.n5 GND 1.25f
C3041 frontAnalog_v0p0p1_5.x63.A.n0 GND 0.12f
C3042 frontAnalog_v0p0p1_5.x63.A.n1 GND 2.22f
C3043 frontAnalog_v0p0p1_5.x63.A.t6 GND 0.014f
C3044 frontAnalog_v0p0p1_5.x63.A.t4 GND 0.0225f
C3045 frontAnalog_v0p0p1_5.x63.A.n2 GND 0.0465f
C3046 frontAnalog_v0p0p1_5.x63.A.t3 GND 0.151f
C3047 frontAnalog_v0p0p1_5.x63.A.t5 GND 0.0256f
C3048 frontAnalog_v0p0p1_5.x63.A.t2 GND 0.173f
C3049 frontAnalog_v0p0p1_5.x63.A.t7 GND 0.175f
C3050 frontAnalog_v0p0p1_5.x63.A.n3 GND 1f
C3051 frontAnalog_v0p0p1_5.x63.A.n4 GND 0.953f
C3052 frontAnalog_v0p0p1_5.x63.A.t1 GND 0.0156f
C3053 frontAnalog_v0p0p1_5.x63.A.t0 GND 0.334f
C3054 frontAnalog_v0p0p1_5.x63.A.n5 GND 1.25f
C3055 frontAnalog_v0p0p1_10.x63.A.n0 GND 0.12f
C3056 frontAnalog_v0p0p1_10.x63.A.n1 GND 2.22f
C3057 frontAnalog_v0p0p1_10.x63.A.t7 GND 0.014f
C3058 frontAnalog_v0p0p1_10.x63.A.t5 GND 0.0225f
C3059 frontAnalog_v0p0p1_10.x63.A.n2 GND 0.0465f
C3060 frontAnalog_v0p0p1_10.x63.A.t2 GND 0.151f
C3061 frontAnalog_v0p0p1_10.x63.A.t6 GND 0.0256f
C3062 frontAnalog_v0p0p1_10.x63.A.t3 GND 0.173f
C3063 frontAnalog_v0p0p1_10.x63.A.t4 GND 0.175f
C3064 frontAnalog_v0p0p1_10.x63.A.n3 GND 1f
C3065 frontAnalog_v0p0p1_10.x63.A.n4 GND 0.953f
C3066 frontAnalog_v0p0p1_10.x63.A.t0 GND 0.0156f
C3067 frontAnalog_v0p0p1_10.x63.A.t1 GND 0.334f
C3068 frontAnalog_v0p0p1_10.x63.A.n5 GND 1.25f
C3069 frontAnalog_v0p0p1_13.x63.A.n0 GND 0.12f
C3070 frontAnalog_v0p0p1_13.x63.A.n1 GND 2.22f
C3071 frontAnalog_v0p0p1_13.x63.A.t6 GND 0.014f
C3072 frontAnalog_v0p0p1_13.x63.A.t4 GND 0.0225f
C3073 frontAnalog_v0p0p1_13.x63.A.n2 GND 0.0465f
C3074 frontAnalog_v0p0p1_13.x63.A.t5 GND 0.0256f
C3075 frontAnalog_v0p0p1_13.x63.A.t1 GND 0.173f
C3076 frontAnalog_v0p0p1_13.x63.A.t7 GND 0.175f
C3077 frontAnalog_v0p0p1_13.x63.A.n3 GND 1f
C3078 frontAnalog_v0p0p1_13.x63.A.n4 GND 0.953f
C3079 frontAnalog_v0p0p1_13.x63.A.t3 GND 0.0156f
C3080 frontAnalog_v0p0p1_13.x63.A.t2 GND 0.335f
C3081 frontAnalog_v0p0p1_13.x63.A.t0 GND 0.151f
C3082 frontAnalog_v0p0p1_13.x63.A.n5 GND 1.25f
C3083 VV7.t17 GND 0.0142f
C3084 VV7.n0 GND 0.116f
C3085 VV7.n1 GND 0.0587f
C3086 VV7.t15 GND 0.186f
C3087 VV7.t7 GND 0.186f
C3088 VV7.t3 GND 0.186f
C3089 VV7.t0 GND 0.186f
C3090 VV7.t13 GND 0.186f
C3091 VV7.t12 GND 0.186f
C3092 VV7.t5 GND 0.186f
C3093 VV7.t2 GND 0.186f
C3094 VV7.t14 GND 0.186f
C3095 VV7.t1 GND 0.186f
C3096 VV7.t9 GND 0.186f
C3097 VV7.t10 GND 0.186f
C3098 VV7.t11 GND 0.186f
C3099 VV7.t6 GND 0.186f
C3100 VV7.t8 GND 0.186f
C3101 VV7.t4 GND 0.186f
C3102 VV7.n2 GND 0.444f
C3103 VV7.n3 GND 0.456f
C3104 VV7.n4 GND 0.456f
C3105 VV7.n5 GND 0.456f
C3106 VV7.n6 GND 0.456f
C3107 VV7.n7 GND 0.456f
C3108 VV7.n8 GND 0.456f
C3109 VV7.n9 GND 0.408f
C3110 VV7.n10 GND 1.04f
C3111 I9.t7 GND 0.0136f
C3112 I9.n0 GND 0.809f
C3113 I9.n1 GND 0.0145f
C3114 I9.n2 GND 0.626f
C3115 I9.n3 GND 1.09f
C3116 I9.n4 GND 1.2f
C3117 I9.t10 GND 0.01f
C3118 I9.t6 GND 0.0307f
C3119 I9.n5 GND 0.481f
C3120 I9.n6 GND 0.0638f
C3121 I9.t3 GND 0.0103f
C3122 I9.n7 GND 0.145f
C3123 I9.n8 GND 0.0959f
C3124 I9.n9 GND 0.103f
C3125 I9.t0 GND 0.0103f
C3126 I9.t1 GND 0.0103f
C3127 I9.n10 GND 0.141f
C3128 I9.n11 GND 0.134f
C3129 I9.t4 GND 0.0113f
C3130 I9.n12 GND 0.32f
C3131 I9.n13 GND 4.81f
C3132 I9.n14 GND 2.83f
C3133 frontAnalog_v0p0p1_7.x63.A.n0 GND 0.12f
C3134 frontAnalog_v0p0p1_7.x63.A.n1 GND 2.22f
C3135 frontAnalog_v0p0p1_7.x63.A.t4 GND 0.014f
C3136 frontAnalog_v0p0p1_7.x63.A.t6 GND 0.0225f
C3137 frontAnalog_v0p0p1_7.x63.A.n2 GND 0.0465f
C3138 frontAnalog_v0p0p1_7.x63.A.t1 GND 0.151f
C3139 frontAnalog_v0p0p1_7.x63.A.t2 GND 0.0156f
C3140 frontAnalog_v0p0p1_7.x63.A.t3 GND 0.335f
C3141 frontAnalog_v0p0p1_7.x63.A.t7 GND 0.0256f
C3142 frontAnalog_v0p0p1_7.x63.A.t0 GND 0.173f
C3143 frontAnalog_v0p0p1_7.x63.A.t5 GND 0.175f
C3144 frontAnalog_v0p0p1_7.x63.A.n3 GND 1f
C3145 frontAnalog_v0p0p1_7.x63.A.n4 GND 0.953f
C3146 frontAnalog_v0p0p1_7.x63.A.n5 GND 1.25f
C3147 frontAnalog_v0p0p1_7.x65.A.n0 GND 0.139f
C3148 frontAnalog_v0p0p1_7.x65.A.t7 GND 0.028f
C3149 frontAnalog_v0p0p1_7.x65.A.t5 GND 0.0175f
C3150 frontAnalog_v0p0p1_7.x65.A.n1 GND 0.0568f
C3151 frontAnalog_v0p0p1_7.x65.A.t3 GND 0.149f
C3152 frontAnalog_v0p0p1_7.x65.A.t6 GND 0.0318f
C3153 frontAnalog_v0p0p1_7.x65.A.t2 GND 0.141f
C3154 frontAnalog_v0p0p1_7.x65.A.t4 GND 0.219f
C3155 frontAnalog_v0p0p1_7.x65.A.n2 GND 1.37f
C3156 frontAnalog_v0p0p1_7.x65.A.n3 GND 0.898f
C3157 frontAnalog_v0p0p1_7.x65.A.t0 GND 0.463f
C3158 frontAnalog_v0p0p1_7.x65.A.t1 GND 0.0194f
C3159 frontAnalog_v0p0p1_7.x65.A.n4 GND 1.6f
C3160 frontAnalog_v0p0p1_7.x65.A.n5 GND 2.01f
C3161 frontAnalog_v0p0p1_7.x65.A.n6 GND 1.72f
C3162 frontAnalog_v0p0p1_13.RSfetsym_0.QN.n0 GND 0.993f
C3163 frontAnalog_v0p0p1_13.RSfetsym_0.QN.t6 GND 0.0317f
C3164 frontAnalog_v0p0p1_13.RSfetsym_0.QN.t5 GND 0.0933f
C3165 frontAnalog_v0p0p1_13.RSfetsym_0.QN.n1 GND 1.47f
C3166 frontAnalog_v0p0p1_13.RSfetsym_0.QN.n2 GND 0.587f
C3167 frontAnalog_v0p0p1_13.RSfetsym_0.QN.t0 GND 0.0363f
C3168 frontAnalog_v0p0p1_13.RSfetsym_0.QN.n3 GND 0.622f
C3169 frontAnalog_v0p0p1_13.RSfetsym_0.QN.t3 GND 0.0317f
C3170 frontAnalog_v0p0p1_13.RSfetsym_0.QN.t2 GND 0.0317f
C3171 frontAnalog_v0p0p1_13.RSfetsym_0.QN.t4 GND 0.0558f
C3172 I6.n0 GND 0.0119f
C3173 I6.n2 GND 0.0166f
C3174 I6.n10 GND 0.147f
C3175 I6.n11 GND 0.372f
C3176 I6.n12 GND 0.0108f
C3177 I6.n13 GND 0.011f
C3178 I6.n14 GND 0.192f
C3179 I6.n17 GND 0.0141f
C3180 I6.n21 GND 0.461f
C3181 I6.n22 GND 0.751f
C3182 I6.n23 GND 0.47f
C3183 I6.n24 GND 1.77f
C3184 I6.t9 GND 0.0111f
C3185 I6.t5 GND 0.034f
C3186 I6.n25 GND 0.533f
C3187 I6.n26 GND 0.0706f
C3188 I6.t0 GND 0.0114f
C3189 I6.n27 GND 0.16f
C3190 I6.n28 GND 0.106f
C3191 I6.n29 GND 0.114f
C3192 I6.t2 GND 0.0114f
C3193 I6.t3 GND 0.0114f
C3194 I6.n30 GND 0.156f
C3195 I6.n31 GND 0.148f
C3196 I6.t4 GND 0.0125f
C3197 I6.n32 GND 0.341f
C3198 I6.n33 GND 9.31f
C3199 I6.n34 GND 2.96f
C3200 frontAnalog_v0p0p1_9.RSfetsym_0.QN.n0 GND 0.993f
C3201 frontAnalog_v0p0p1_9.RSfetsym_0.QN.t6 GND 0.0317f
C3202 frontAnalog_v0p0p1_9.RSfetsym_0.QN.t5 GND 0.0933f
C3203 frontAnalog_v0p0p1_9.RSfetsym_0.QN.n1 GND 1.47f
C3204 frontAnalog_v0p0p1_9.RSfetsym_0.QN.n2 GND 0.587f
C3205 frontAnalog_v0p0p1_9.RSfetsym_0.QN.t1 GND 0.0363f
C3206 frontAnalog_v0p0p1_9.RSfetsym_0.QN.n3 GND 0.622f
C3207 frontAnalog_v0p0p1_9.RSfetsym_0.QN.t3 GND 0.0317f
C3208 frontAnalog_v0p0p1_9.RSfetsym_0.QN.t4 GND 0.0317f
C3209 frontAnalog_v0p0p1_9.RSfetsym_0.QN.t0 GND 0.0558f
C3210 I1.n0 GND 0.361f
C3211 I1.n2 GND 0.268f
C3212 I1.n3 GND 0.476f
C3213 I1.n4 GND 0.342f
C3214 I1.t5 GND 0.0134f
C3215 I1.n5 GND 0.211f
C3216 I1.n6 GND 0.0279f
C3217 I1.n7 GND 0.0633f
C3218 I1.n8 GND 0.042f
C3219 I1.n9 GND 0.0449f
C3220 I1.n10 GND 0.0619f
C3221 I1.n11 GND 0.0585f
C3222 I1.n12 GND 0.135f
C3223 I1.n13 GND 10.5f
C3224 I1.n14 GND 0.517f
C3225 frontAnalog_v0p0p1_9.x65.A.n0 GND 0.139f
C3226 frontAnalog_v0p0p1_9.x65.A.t6 GND 0.028f
C3227 frontAnalog_v0p0p1_9.x65.A.t4 GND 0.0175f
C3228 frontAnalog_v0p0p1_9.x65.A.n1 GND 0.0568f
C3229 frontAnalog_v0p0p1_9.x65.A.t2 GND 0.149f
C3230 frontAnalog_v0p0p1_9.x65.A.t5 GND 0.0318f
C3231 frontAnalog_v0p0p1_9.x65.A.t3 GND 0.141f
C3232 frontAnalog_v0p0p1_9.x65.A.t7 GND 0.219f
C3233 frontAnalog_v0p0p1_9.x65.A.n2 GND 1.37f
C3234 frontAnalog_v0p0p1_9.x65.A.n3 GND 0.898f
C3235 frontAnalog_v0p0p1_9.x65.A.t1 GND 0.463f
C3236 frontAnalog_v0p0p1_9.x65.A.t0 GND 0.0194f
C3237 frontAnalog_v0p0p1_9.x65.A.n4 GND 1.6f
C3238 frontAnalog_v0p0p1_9.x65.A.n5 GND 2.01f
C3239 frontAnalog_v0p0p1_9.x65.A.n6 GND 1.72f
C3240 frontAnalog_v0p0p1_9.x63.A.n0 GND 0.12f
C3241 frontAnalog_v0p0p1_9.x63.A.n1 GND 2.22f
C3242 frontAnalog_v0p0p1_9.x63.A.t7 GND 0.014f
C3243 frontAnalog_v0p0p1_9.x63.A.t5 GND 0.0225f
C3244 frontAnalog_v0p0p1_9.x63.A.n2 GND 0.0465f
C3245 frontAnalog_v0p0p1_9.x63.A.t1 GND 0.151f
C3246 frontAnalog_v0p0p1_9.x63.A.t2 GND 0.0156f
C3247 frontAnalog_v0p0p1_9.x63.A.t3 GND 0.335f
C3248 frontAnalog_v0p0p1_9.x63.A.t6 GND 0.0256f
C3249 frontAnalog_v0p0p1_9.x63.A.t0 GND 0.173f
C3250 frontAnalog_v0p0p1_9.x63.A.t4 GND 0.175f
C3251 frontAnalog_v0p0p1_9.x63.A.n3 GND 1f
C3252 frontAnalog_v0p0p1_9.x63.A.n4 GND 0.953f
C3253 frontAnalog_v0p0p1_9.x63.A.n5 GND 1.25f
C3254 VV12.t16 GND 0.0144f
C3255 VV12.n0 GND 0.118f
C3256 VV12.n1 GND 0.0572f
C3257 VV12.t11 GND 0.189f
C3258 VV12.t2 GND 0.189f
C3259 VV12.t7 GND 0.189f
C3260 VV12.t9 GND 0.189f
C3261 VV12.t1 GND 0.189f
C3262 VV12.t14 GND 0.189f
C3263 VV12.t13 GND 0.189f
C3264 VV12.t6 GND 0.189f
C3265 VV12.t10 GND 0.189f
C3266 VV12.t15 GND 0.189f
C3267 VV12.t12 GND 0.189f
C3268 VV12.t0 GND 0.189f
C3269 VV12.t3 GND 0.189f
C3270 VV12.t4 GND 0.189f
C3271 VV12.t8 GND 0.189f
C3272 VV12.t5 GND 0.407f
C3273 VV12.n2 GND 0.234f
C3274 VV12.n3 GND 0.232f
C3275 VV12.n4 GND 0.232f
C3276 VV12.n5 GND 0.232f
C3277 VV12.n6 GND 0.232f
C3278 VV12.n7 GND 0.232f
C3279 VV12.n8 GND 0.232f
C3280 VV12.n9 GND 0.232f
C3281 VV12.n10 GND 0.232f
C3282 VV12.n11 GND 0.232f
C3283 VV12.n12 GND 0.232f
C3284 VV12.n13 GND 0.232f
C3285 VV12.n14 GND 0.232f
C3286 VV12.n15 GND 0.232f
C3287 VV12.n16 GND 0.183f
C3288 VV12.n17 GND 1.28f
C3289 frontAnalog_v0p0p1_4.x65.A.n0 GND 0.139f
C3290 frontAnalog_v0p0p1_4.x65.A.t4 GND 0.028f
C3291 frontAnalog_v0p0p1_4.x65.A.t5 GND 0.0175f
C3292 frontAnalog_v0p0p1_4.x65.A.n1 GND 0.0568f
C3293 frontAnalog_v0p0p1_4.x65.A.t7 GND 0.0318f
C3294 frontAnalog_v0p0p1_4.x65.A.t1 GND 0.141f
C3295 frontAnalog_v0p0p1_4.x65.A.t6 GND 0.219f
C3296 frontAnalog_v0p0p1_4.x65.A.n2 GND 1.37f
C3297 frontAnalog_v0p0p1_4.x65.A.n3 GND 0.898f
C3298 frontAnalog_v0p0p1_4.x65.A.t3 GND 0.463f
C3299 frontAnalog_v0p0p1_4.x65.A.t2 GND 0.0194f
C3300 frontAnalog_v0p0p1_4.x65.A.n4 GND 1.6f
C3301 frontAnalog_v0p0p1_4.x65.A.n5 GND 2.01f
C3302 frontAnalog_v0p0p1_4.x65.A.t0 GND 0.149f
C3303 frontAnalog_v0p0p1_4.x65.A.n6 GND 1.72f
C3304 VIN.t3 GND 0.0442f
C3305 VIN.n0 GND 0.357f
C3306 VIN.n1 GND 0.0997f
C3307 VIN.t17 GND 0.0442f
C3308 VIN.n3 GND 0.354f
C3309 VIN.n4 GND 4.47f
C3310 VIN.t22 GND 0.0442f
C3311 VIN.n5 GND 0.357f
C3312 VIN.t8 GND 0.0442f
C3313 VIN.n6 GND 0.354f
C3314 VIN.t14 GND 0.0442f
C3315 VIN.n7 GND 0.357f
C3316 VIN.t29 GND 0.0442f
C3317 VIN.n8 GND 0.357f
C3318 VIN.t2 GND 0.0442f
C3319 VIN.n9 GND 0.357f
C3320 VIN.t9 GND 0.0442f
C3321 VIN.n10 GND 0.357f
C3322 VIN.t27 GND 0.0442f
C3323 VIN.n11 GND 0.357f
C3324 VIN.t30 GND 0.0442f
C3325 VIN.n12 GND 0.357f
C3326 VIN.t21 GND 0.0442f
C3327 VIN.n13 GND 0.357f
C3328 VIN.t25 GND 0.0442f
C3329 VIN.n14 GND 0.357f
C3330 VIN.t12 GND 0.0442f
C3331 VIN.n15 GND 0.357f
C3332 VIN.t18 GND 0.0442f
C3333 VIN.n16 GND 0.357f
C3334 VIN.t0 GND 0.0442f
C3335 VIN.n17 GND 0.357f
C3336 VIN.t7 GND 0.0442f
C3337 VIN.n18 GND 0.357f
C3338 VIN.n19 GND 9.36f
C3339 VIN.n20 GND 5.84f
C3340 VIN.n21 GND 5.83f
C3341 VIN.n22 GND 5.84f
C3342 VIN.n23 GND 5.84f
C3343 VIN.n24 GND 5.84f
C3344 VIN.n25 GND 5.85f
C3345 VIN.n26 GND 5.84f
C3346 VIN.n27 GND 5.84f
C3347 VIN.n28 GND 5.84f
C3348 VIN.n29 GND 5.83f
C3349 VIN.n30 GND 5.81f
C3350 VIN.n31 GND 5.84f
C3351 VIN.n32 GND 5.9f
C3352 VIN.n33 GND 0.932f
C3353 VV13.t17 GND 0.0152f
C3354 VV13.n0 GND 0.125f
C3355 VV13.n1 GND 0.0603f
C3356 VV13.t2 GND 0.199f
C3357 VV13.t7 GND 0.199f
C3358 VV13.t9 GND 0.199f
C3359 VV13.t14 GND 0.199f
C3360 VV13.t13 GND 0.199f
C3361 VV13.t3 GND 0.199f
C3362 VV13.t8 GND 0.199f
C3363 VV13.t0 GND 0.199f
C3364 VV13.t15 GND 0.199f
C3365 VV13.t12 GND 0.199f
C3366 VV13.t1 GND 0.199f
C3367 VV13.t5 GND 0.199f
C3368 VV13.t4 GND 0.199f
C3369 VV13.t11 GND 0.199f
C3370 VV13.t6 GND 0.199f
C3371 VV13.t10 GND 0.199f
C3372 VV13.n2 GND 0.476f
C3373 VV13.n3 GND 0.489f
C3374 VV13.n4 GND 0.489f
C3375 VV13.n5 GND 0.489f
C3376 VV13.n6 GND 0.489f
C3377 VV13.n7 GND 0.489f
C3378 VV13.n8 GND 0.489f
C3379 VV13.n9 GND 0.434f
C3380 VV13.n10 GND 1.44f
C3381 VV14.t16 GND 0.0161f
C3382 VV14.n0 GND 0.132f
C3383 VV14.n1 GND 0.061f
C3384 VV14.t8 GND 0.21f
C3385 VV14.t7 GND 0.21f
C3386 VV14.t12 GND 0.21f
C3387 VV14.t4 GND 0.21f
C3388 VV14.t5 GND 0.21f
C3389 VV14.t3 GND 0.21f
C3390 VV14.t1 GND 0.21f
C3391 VV14.t2 GND 0.21f
C3392 VV14.t11 GND 0.21f
C3393 VV14.t0 GND 0.21f
C3394 VV14.t6 GND 0.21f
C3395 VV14.t15 GND 0.21f
C3396 VV14.t10 GND 0.21f
C3397 VV14.t13 GND 0.21f
C3398 VV14.t9 GND 0.21f
C3399 VV14.t14 GND 0.21f
C3400 VV14.n2 GND 0.504f
C3401 VV14.n3 GND 0.517f
C3402 VV14.n4 GND 0.517f
C3403 VV14.n5 GND 0.517f
C3404 VV14.n6 GND 0.517f
C3405 VV14.n7 GND 0.517f
C3406 VV14.n8 GND 0.517f
C3407 VV14.n9 GND 0.464f
C3408 VV14.n10 GND 1.62f
C3409 frontAnalog_v0p0p1_10.IB.n0 GND 0.0481f
C3410 frontAnalog_v0p0p1_10.IB.t12 GND 0.0551f
C3411 frontAnalog_v0p0p1_10.IB.t23 GND 0.0545f
C3412 frontAnalog_v0p0p1_10.IB.t3 GND 0.0551f
C3413 frontAnalog_v0p0p1_10.IB.t11 GND 0.0545f
C3414 frontAnalog_v0p0p1_10.IB.n3 GND 5.42f
C3415 frontAnalog_v0p0p1_10.IB.t32 GND 0.0551f
C3416 frontAnalog_v0p0p1_10.IB.t9 GND 0.0545f
C3417 frontAnalog_v0p0p1_10.IB.t5 GND 0.0551f
C3418 frontAnalog_v0p0p1_10.IB.t29 GND 0.0545f
C3419 frontAnalog_v0p0p1_10.IB.t22 GND 0.0551f
C3420 frontAnalog_v0p0p1_10.IB.t34 GND 0.0545f
C3421 frontAnalog_v0p0p1_10.IB.t26 GND 0.0551f
C3422 frontAnalog_v0p0p1_10.IB.t19 GND 0.0545f
C3423 frontAnalog_v0p0p1_10.IB.t15 GND 0.0551f
C3424 frontAnalog_v0p0p1_10.IB.t25 GND 0.0545f
C3425 frontAnalog_v0p0p1_10.IB.t18 GND 0.0551f
C3426 frontAnalog_v0p0p1_10.IB.t30 GND 0.0545f
C3427 frontAnalog_v0p0p1_10.IB.t7 GND 0.0551f
C3428 frontAnalog_v0p0p1_10.IB.t16 GND 0.0545f
C3429 frontAnalog_v0p0p1_10.IB.t10 GND 0.0551f
C3430 frontAnalog_v0p0p1_10.IB.t20 GND 0.0545f
C3431 frontAnalog_v0p0p1_10.IB.t31 GND 0.0551f
C3432 frontAnalog_v0p0p1_10.IB.t8 GND 0.0545f
C3433 frontAnalog_v0p0p1_10.IB.t4 GND 0.0551f
C3434 frontAnalog_v0p0p1_10.IB.t13 GND 0.0545f
C3435 frontAnalog_v0p0p1_10.IB.t21 GND 0.0551f
C3436 frontAnalog_v0p0p1_10.IB.t33 GND 0.0545f
C3437 frontAnalog_v0p0p1_10.IB.t27 GND 0.0551f
C3438 frontAnalog_v0p0p1_10.IB.t6 GND 0.0545f
C3439 frontAnalog_v0p0p1_10.IB.t14 GND 0.0551f
C3440 frontAnalog_v0p0p1_10.IB.t24 GND 0.0545f
C3441 frontAnalog_v0p0p1_10.IB.t17 GND 0.0551f
C3442 frontAnalog_v0p0p1_10.IB.t28 GND 0.0545f
C3443 frontAnalog_v0p0p1_10.IB.n18 GND 8.11f
C3444 frontAnalog_v0p0p1_10.IB.n19 GND 5.61f
C3445 frontAnalog_v0p0p1_10.IB.n20 GND 5.58f
C3446 frontAnalog_v0p0p1_10.IB.n21 GND 5.65f
C3447 frontAnalog_v0p0p1_10.IB.n22 GND 5.58f
C3448 frontAnalog_v0p0p1_10.IB.n23 GND 5.62f
C3449 frontAnalog_v0p0p1_10.IB.n24 GND 5.59f
C3450 frontAnalog_v0p0p1_10.IB.n25 GND 5.61f
C3451 frontAnalog_v0p0p1_10.IB.n26 GND 5.57f
C3452 frontAnalog_v0p0p1_10.IB.n27 GND 5.58f
C3453 frontAnalog_v0p0p1_10.IB.n28 GND 5.62f
C3454 frontAnalog_v0p0p1_10.IB.n29 GND 5.65f
C3455 frontAnalog_v0p0p1_10.IB.n30 GND 4.67f
C3456 frontAnalog_v0p0p1_10.IB.n31 GND 9.74f
C3457 frontAnalog_v0p0p1_10.IB.t1 GND 0.0307f
C3458 frontAnalog_v0p0p1_10.IB.n32 GND 0.0823f
C3459 frontAnalog_v0p0p1_10.IB.t0 GND 0.42f
C3460 frontAnalog_v0p0p1_10.IB.n34 GND 7.2f
C3461 I13.n8 GND 0.0978f
C3462 I13.n9 GND 0.228f
C3463 I13.n16 GND 0.139f
C3464 I13.n21 GND 0.369f
C3465 I13.n22 GND 0.874f
C3466 I13.n23 GND 0.408f
C3467 I13.n24 GND 0.253f
C3468 I13.n25 GND 0.578f
C3469 I13.t12 GND 0.018f
C3470 I13.n26 GND 0.282f
C3471 I13.n27 GND 0.0373f
C3472 I13.n28 GND 0.0846f
C3473 I13.n29 GND 0.0561f
C3474 I13.n30 GND 0.06f
C3475 I13.n31 GND 0.0827f
C3476 I13.n32 GND 0.0783f
C3477 I13.n33 GND 0.188f
C3478 I13.n34 GND 12.1f
C3479 frontAnalog_v0p0p1_6.RSfetsym_0.QN.n0 GND 0.993f
C3480 frontAnalog_v0p0p1_6.RSfetsym_0.QN.t6 GND 0.0317f
C3481 frontAnalog_v0p0p1_6.RSfetsym_0.QN.t5 GND 0.0933f
C3482 frontAnalog_v0p0p1_6.RSfetsym_0.QN.n1 GND 1.47f
C3483 frontAnalog_v0p0p1_6.RSfetsym_0.QN.n2 GND 0.587f
C3484 frontAnalog_v0p0p1_6.RSfetsym_0.QN.t4 GND 0.0363f
C3485 frontAnalog_v0p0p1_6.RSfetsym_0.QN.n3 GND 0.622f
C3486 frontAnalog_v0p0p1_6.RSfetsym_0.QN.t1 GND 0.0317f
C3487 frontAnalog_v0p0p1_6.RSfetsym_0.QN.t2 GND 0.0317f
C3488 frontAnalog_v0p0p1_6.RSfetsym_0.QN.t3 GND 0.0558f
C3489 I10.n0 GND 0.0143f
C3490 I10.n1 GND 0.103f
C3491 I10.n2 GND 0.21f
C3492 I10.n5 GND 0.523f
C3493 I10.n6 GND 0.0163f
C3494 I10.n7 GND 0.076f
C3495 I10.n8 GND 1.27f
C3496 I10.n9 GND 1.53f
C3497 I10.t5 GND 0.0289f
C3498 I10.n10 GND 0.452f
C3499 I10.n11 GND 0.0599f
C3500 I10.n12 GND 0.136f
C3501 I10.n13 GND 0.0901f
C3502 I10.n14 GND 0.0963f
C3503 I10.n15 GND 0.133f
C3504 I10.n16 GND 0.126f
C3505 I10.t4 GND 0.0106f
C3506 I10.n17 GND 0.302f
C3507 I10.n18 GND 8.36f
C3508 I10.n19 GND 3.31f
C3509 VV5.t16 GND 0.0157f
C3510 VV5.n0 GND 0.129f
C3511 VV5.n1 GND 0.0622f
C3512 VV5.t12 GND 0.205f
C3513 VV5.t15 GND 0.205f
C3514 VV5.t13 GND 0.205f
C3515 VV5.t5 GND 0.205f
C3516 VV5.t11 GND 0.205f
C3517 VV5.t14 GND 0.205f
C3518 VV5.t2 GND 0.205f
C3519 VV5.t1 GND 0.205f
C3520 VV5.t9 GND 0.205f
C3521 VV5.t10 GND 0.205f
C3522 VV5.t3 GND 0.205f
C3523 VV5.t8 GND 0.205f
C3524 VV5.t7 GND 0.205f
C3525 VV5.t0 GND 0.205f
C3526 VV5.t6 GND 0.205f
C3527 VV5.t4 GND 0.205f
C3528 VV5.n2 GND 0.491f
C3529 VV5.n3 GND 0.504f
C3530 VV5.n4 GND 0.504f
C3531 VV5.n5 GND 0.504f
C3532 VV5.n6 GND 0.504f
C3533 VV5.n7 GND 0.504f
C3534 VV5.n8 GND 0.504f
C3535 VV5.n9 GND 0.454f
C3536 VV5.n10 GND 1.33f
C3537 VV6.t16 GND 0.0149f
C3538 VV6.n0 GND 0.122f
C3539 VV6.n1 GND 0.0591f
C3540 VV6.t8 GND 0.195f
C3541 VV6.t14 GND 0.195f
C3542 VV6.t0 GND 0.195f
C3543 VV6.t15 GND 0.195f
C3544 VV6.t12 GND 0.195f
C3545 VV6.t13 GND 0.195f
C3546 VV6.t5 GND 0.195f
C3547 VV6.t2 GND 0.195f
C3548 VV6.t1 GND 0.195f
C3549 VV6.t9 GND 0.195f
C3550 VV6.t11 GND 0.195f
C3551 VV6.t3 GND 0.195f
C3552 VV6.t7 GND 0.195f
C3553 VV6.t6 GND 0.195f
C3554 VV6.t4 GND 0.195f
C3555 VV6.t10 GND 0.195f
C3556 VV6.n2 GND 0.467f
C3557 VV6.n3 GND 0.479f
C3558 VV6.n4 GND 0.479f
C3559 VV6.n5 GND 0.479f
C3560 VV6.n6 GND 0.479f
C3561 VV6.n7 GND 0.479f
C3562 VV6.n8 GND 0.479f
C3563 VV6.n9 GND 0.426f
C3564 VV6.n10 GND 1.18f
C3565 frontAnalog_v0p0p1_15.RSfetsym_0.QN.n0 GND 1.01f
C3566 frontAnalog_v0p0p1_15.RSfetsym_0.QN.t6 GND 0.0321f
C3567 frontAnalog_v0p0p1_15.RSfetsym_0.QN.t5 GND 0.0947f
C3568 frontAnalog_v0p0p1_15.RSfetsym_0.QN.n1 GND 1.49f
C3569 frontAnalog_v0p0p1_15.RSfetsym_0.QN.n2 GND 0.595f
C3570 frontAnalog_v0p0p1_15.RSfetsym_0.QN.t4 GND 0.0368f
C3571 frontAnalog_v0p0p1_15.RSfetsym_0.QN.n3 GND 0.631f
C3572 frontAnalog_v0p0p1_15.RSfetsym_0.QN.t1 GND 0.0322f
C3573 frontAnalog_v0p0p1_15.RSfetsym_0.QN.t0 GND 0.0322f
C3574 frontAnalog_v0p0p1_15.RSfetsym_0.QN.t3 GND 0.0566f
C3575 frontAnalog_v0p0p1_2.x65.A.n0 GND 0.139f
C3576 frontAnalog_v0p0p1_2.x65.A.t4 GND 0.028f
C3577 frontAnalog_v0p0p1_2.x65.A.t5 GND 0.0175f
C3578 frontAnalog_v0p0p1_2.x65.A.n1 GND 0.0568f
C3579 frontAnalog_v0p0p1_2.x65.A.t1 GND 0.149f
C3580 frontAnalog_v0p0p1_2.x65.A.t3 GND 0.463f
C3581 frontAnalog_v0p0p1_2.x65.A.t2 GND 0.0194f
C3582 frontAnalog_v0p0p1_2.x65.A.n2 GND 1.6f
C3583 frontAnalog_v0p0p1_2.x65.A.t6 GND 0.0318f
C3584 frontAnalog_v0p0p1_2.x65.A.t0 GND 0.141f
C3585 frontAnalog_v0p0p1_2.x65.A.t7 GND 0.219f
C3586 frontAnalog_v0p0p1_2.x65.A.n3 GND 1.37f
C3587 frontAnalog_v0p0p1_2.x65.A.n4 GND 0.898f
C3588 frontAnalog_v0p0p1_2.x65.A.n5 GND 2.01f
C3589 frontAnalog_v0p0p1_2.x65.A.n6 GND 1.72f
C3590 frontAnalog_v0p0p1_2.x63.A.n0 GND 0.12f
C3591 frontAnalog_v0p0p1_2.x63.A.n1 GND 2.22f
C3592 frontAnalog_v0p0p1_2.x63.A.t6 GND 0.014f
C3593 frontAnalog_v0p0p1_2.x63.A.t5 GND 0.0225f
C3594 frontAnalog_v0p0p1_2.x63.A.n2 GND 0.0465f
C3595 frontAnalog_v0p0p1_2.x63.A.t2 GND 0.151f
C3596 frontAnalog_v0p0p1_2.x63.A.t0 GND 0.0156f
C3597 frontAnalog_v0p0p1_2.x63.A.t3 GND 0.335f
C3598 frontAnalog_v0p0p1_2.x63.A.t4 GND 0.0256f
C3599 frontAnalog_v0p0p1_2.x63.A.t1 GND 0.173f
C3600 frontAnalog_v0p0p1_2.x63.A.t7 GND 0.175f
C3601 frontAnalog_v0p0p1_2.x63.A.n3 GND 1f
C3602 frontAnalog_v0p0p1_2.x63.A.n4 GND 0.953f
C3603 frontAnalog_v0p0p1_2.x63.A.n5 GND 1.25f
C3604 VV15.t17 GND 0.017f
C3605 VV15.n0 GND 0.139f
C3606 VV15.n1 GND 0.0644f
C3607 VV15.t7 GND 0.222f
C3608 VV15.t2 GND 0.222f
C3609 VV15.t5 GND 0.222f
C3610 VV15.t6 GND 0.222f
C3611 VV15.t4 GND 0.222f
C3612 VV15.t0 GND 0.222f
C3613 VV15.t3 GND 0.222f
C3614 VV15.t9 GND 0.222f
C3615 VV15.t1 GND 0.222f
C3616 VV15.t8 GND 0.222f
C3617 VV15.t14 GND 0.222f
C3618 VV15.t15 GND 0.222f
C3619 VV15.t11 GND 0.222f
C3620 VV15.t13 GND 0.222f
C3621 VV15.t12 GND 0.222f
C3622 VV15.t10 GND 0.222f
C3623 VV15.n2 GND 0.532f
C3624 VV15.n3 GND 0.546f
C3625 VV15.n4 GND 0.546f
C3626 VV15.n5 GND 0.546f
C3627 VV15.n6 GND 0.546f
C3628 VV15.n7 GND 0.546f
C3629 VV15.n8 GND 0.546f
C3630 VV15.n9 GND 0.487f
C3631 VV9.t16 GND 0.013f
C3632 VV9.n0 GND 0.107f
C3633 VV9.n1 GND 0.0517f
C3634 VV9.t3 GND 0.171f
C3635 VV9.t13 GND 0.171f
C3636 VV9.t15 GND 0.171f
C3637 VV9.t9 GND 0.171f
C3638 VV9.t10 GND 0.171f
C3639 VV9.t11 GND 0.171f
C3640 VV9.t8 GND 0.171f
C3641 VV9.t5 GND 0.171f
C3642 VV9.t2 GND 0.171f
C3643 VV9.t1 GND 0.171f
C3644 VV9.t6 GND 0.171f
C3645 VV9.t0 GND 0.171f
C3646 VV9.t4 GND 0.171f
C3647 VV9.t7 GND 0.171f
C3648 VV9.t12 GND 0.171f
C3649 VV9.t14 GND 0.171f
C3650 VV9.n2 GND 0.408f
C3651 VV9.n3 GND 0.419f
C3652 VV9.n4 GND 0.419f
C3653 VV9.n5 GND 0.419f
C3654 VV9.n6 GND 0.419f
C3655 VV9.n7 GND 0.419f
C3656 VV9.n8 GND 0.419f
C3657 VV9.n9 GND 0.376f
C3658 VV9.n10 GND 0.954f
C3659 frontAnalog_v0p0p1_8.RSfetsym_0.QN.n0 GND 0.993f
C3660 frontAnalog_v0p0p1_8.RSfetsym_0.QN.t5 GND 0.0317f
C3661 frontAnalog_v0p0p1_8.RSfetsym_0.QN.t6 GND 0.0933f
C3662 frontAnalog_v0p0p1_8.RSfetsym_0.QN.n1 GND 1.47f
C3663 frontAnalog_v0p0p1_8.RSfetsym_0.QN.n2 GND 0.587f
C3664 frontAnalog_v0p0p1_8.RSfetsym_0.QN.t1 GND 0.0363f
C3665 frontAnalog_v0p0p1_8.RSfetsym_0.QN.n3 GND 0.622f
C3666 frontAnalog_v0p0p1_8.RSfetsym_0.QN.t3 GND 0.0317f
C3667 frontAnalog_v0p0p1_8.RSfetsym_0.QN.t4 GND 0.0317f
C3668 frontAnalog_v0p0p1_8.RSfetsym_0.QN.t0 GND 0.0558f
C3669 OUT1.n2 GND 0.0114f
C3670 OUT1.n4 GND 0.0242f
C3671 OUT1.n6 GND 0.0161f
C3672 OUT1.n8 GND 0.0161f
C3673 OUT1.n10 GND 0.0161f
C3674 OUT1.n12 GND 0.0161f
C3675 OUT1.n14 GND 0.0161f
C3676 OUT1.n23 GND 0.014f
C3677 OUT1.n25 GND 0.0348f
C3678 OUT1.n27 GND 0.021f
C3679 OUT1.n29 GND 0.021f
C3680 OUT1.n31 GND 0.021f
C3681 OUT1.n33 GND 0.021f
C3682 OUT1.n35 GND 0.021f
C3683 OUT1.n37 GND 0.0147f
C3684 OUT1.n38 GND 0.0297f
C3685 OUT1.n39 GND 0.0229f
C3686 OUT1.n42 GND 0.0114f
C3687 OUT1.n44 GND 0.0242f
C3688 OUT1.n46 GND 0.0161f
C3689 OUT1.n48 GND 0.0161f
C3690 OUT1.n50 GND 0.0161f
C3691 OUT1.n52 GND 0.0161f
C3692 OUT1.n54 GND 0.0161f
C3693 OUT1.n63 GND 0.014f
C3694 OUT1.n65 GND 0.0348f
C3695 OUT1.n67 GND 0.021f
C3696 OUT1.n69 GND 0.021f
C3697 OUT1.n71 GND 0.021f
C3698 OUT1.n73 GND 0.021f
C3699 OUT1.n75 GND 0.021f
C3700 OUT1.n77 GND 0.0147f
C3701 OUT1.n78 GND 0.0274f
C3702 OUT1.n79 GND 0.0203f
C3703 OUT1.n81 GND 0.0114f
C3704 OUT1.n83 GND 0.0242f
C3705 OUT1.n85 GND 0.0161f
C3706 OUT1.n87 GND 0.0161f
C3707 OUT1.n89 GND 0.0161f
C3708 OUT1.n91 GND 0.0161f
C3709 OUT1.n93 GND 0.0161f
C3710 OUT1.n97 GND 0.0126f
C3711 OUT1.n100 GND 0.014f
C3712 OUT1.n102 GND 0.0348f
C3713 OUT1.n104 GND 0.021f
C3714 OUT1.n106 GND 0.021f
C3715 OUT1.n108 GND 0.021f
C3716 OUT1.n110 GND 0.021f
C3717 OUT1.n112 GND 0.021f
C3718 OUT1.n114 GND 0.0147f
C3719 OUT1.n115 GND 0.0284f
C3720 OUT1.n116 GND 0.0234f
C3721 OUT1.n120 GND 0.014f
C3722 OUT1.n122 GND 0.0348f
C3723 OUT1.n124 GND 0.021f
C3724 OUT1.n126 GND 0.021f
C3725 OUT1.n128 GND 0.021f
C3726 OUT1.n130 GND 0.021f
C3727 OUT1.n132 GND 0.021f
C3728 OUT1.n136 GND 0.0114f
C3729 OUT1.n138 GND 0.0242f
C3730 OUT1.n140 GND 0.0161f
C3731 OUT1.n142 GND 0.0161f
C3732 OUT1.n144 GND 0.0161f
C3733 OUT1.n146 GND 0.0161f
C3734 OUT1.n148 GND 0.0161f
C3735 OUT1.n152 GND 0.0129f
C3736 OUT1.n155 GND 0.0204f
C3737 OUT1.n156 GND 0.108f
C3738 OUT1.n157 GND 0.275f
C3739 OUT1.n158 GND 0.224f
C3740 OUT1.n159 GND 0.228f
C3741 I2.n1 GND 0.0614f
C3742 I2.n2 GND 0.125f
C3743 I2.n5 GND 0.319f
C3744 I2.n7 GND 0.0432f
C3745 I2.n8 GND 0.756f
C3746 I2.n9 GND 0.531f
C3747 I2.t10 GND 0.0171f
C3748 I2.n10 GND 0.269f
C3749 I2.n11 GND 0.0356f
C3750 I2.n12 GND 0.0807f
C3751 I2.n13 GND 0.0535f
C3752 I2.n14 GND 0.0572f
C3753 I2.n15 GND 0.0789f
C3754 I2.n16 GND 0.0746f
C3755 I2.n17 GND 0.172f
C3756 I2.n18 GND 11.7f
C3757 I2.n19 GND 0.833f
C3758 I0.n1 GND 0.0888f
C3759 I0.n2 GND 0.237f
C3760 I0.n3 GND 0.291f
C3761 I0.n4 GND 0.137f
C3762 I0.n5 GND 0.0181f
C3763 I0.n6 GND 0.0411f
C3764 I0.n7 GND 0.0272f
C3765 I0.n8 GND 0.0292f
C3766 I0.n9 GND 0.0402f
C3767 I0.n10 GND 0.038f
C3768 I0.n11 GND 0.0875f
C3769 I0.n12 GND 7.73f
C3770 I0.n13 GND 0.247f
C3771 VV1.n0 GND 0.0483f
C3772 VV1.n1 GND 0.0234f
C3773 VV1.t12 GND 0.0771f
C3774 VV1.t8 GND 0.0771f
C3775 VV1.t3 GND 0.0771f
C3776 VV1.t0 GND 0.0771f
C3777 VV1.t15 GND 0.0771f
C3778 VV1.t1 GND 0.0771f
C3779 VV1.t4 GND 0.0771f
C3780 VV1.t13 GND 0.0771f
C3781 VV1.t11 GND 0.0771f
C3782 VV1.t7 GND 0.0771f
C3783 VV1.t2 GND 0.0771f
C3784 VV1.t10 GND 0.0771f
C3785 VV1.t14 GND 0.0771f
C3786 VV1.t9 GND 0.0771f
C3787 VV1.t6 GND 0.0771f
C3788 VV1.t5 GND 0.0771f
C3789 VV1.n2 GND 0.185f
C3790 VV1.n3 GND 0.189f
C3791 VV1.n4 GND 0.189f
C3792 VV1.n5 GND 0.189f
C3793 VV1.n6 GND 0.189f
C3794 VV1.n7 GND 0.189f
C3795 VV1.n8 GND 0.189f
C3796 VV1.n9 GND 0.168f
C3797 VV1.n10 GND 0.548f
C3798 VV2.t17 GND 0.0148f
C3799 VV2.n0 GND 0.121f
C3800 VV2.n1 GND 0.0611f
C3801 VV2.t4 GND 0.193f
C3802 VV2.t10 GND 0.193f
C3803 VV2.t12 GND 0.193f
C3804 VV2.t5 GND 0.193f
C3805 VV2.t14 GND 0.193f
C3806 VV2.t15 GND 0.193f
C3807 VV2.t0 GND 0.193f
C3808 VV2.t6 GND 0.193f
C3809 VV2.t8 GND 0.193f
C3810 VV2.t9 GND 0.193f
C3811 VV2.t1 GND 0.193f
C3812 VV2.t3 GND 0.193f
C3813 VV2.t11 GND 0.193f
C3814 VV2.t13 GND 0.193f
C3815 VV2.t7 GND 0.416f
C3816 VV2.t2 GND 0.193f
C3817 VV2.n2 GND 0.239f
C3818 VV2.n3 GND 0.237f
C3819 VV2.n4 GND 0.237f
C3820 VV2.n5 GND 0.237f
C3821 VV2.n6 GND 0.237f
C3822 VV2.n7 GND 0.237f
C3823 VV2.n8 GND 0.237f
C3824 VV2.n9 GND 0.237f
C3825 VV2.n10 GND 0.237f
C3826 VV2.n11 GND 0.237f
C3827 VV2.n12 GND 0.237f
C3828 VV2.n13 GND 0.237f
C3829 VV2.n14 GND 0.237f
C3830 VV2.n15 GND 0.237f
C3831 VV2.n16 GND 0.182f
C3832 VV2.n17 GND 1.5f
C3833 VV10.t17 GND 0.0124f
C3834 VV10.n0 GND 0.102f
C3835 VV10.n1 GND 0.0513f
C3836 VV10.t14 GND 0.162f
C3837 VV10.t8 GND 0.162f
C3838 VV10.t11 GND 0.162f
C3839 VV10.t3 GND 0.162f
C3840 VV10.t13 GND 0.162f
C3841 VV10.t9 GND 0.162f
C3842 VV10.t5 GND 0.162f
C3843 VV10.t1 GND 0.162f
C3844 VV10.t2 GND 0.162f
C3845 VV10.t6 GND 0.162f
C3846 VV10.t0 GND 0.162f
C3847 VV10.t10 GND 0.162f
C3848 VV10.t7 GND 0.162f
C3849 VV10.t4 GND 0.162f
C3850 VV10.t15 GND 0.162f
C3851 VV10.t12 GND 0.162f
C3852 VV10.n2 GND 0.388f
C3853 VV10.n3 GND 0.398f
C3854 VV10.n4 GND 0.398f
C3855 VV10.n5 GND 0.398f
C3856 VV10.n6 GND 0.398f
C3857 VV10.n7 GND 0.398f
C3858 VV10.n8 GND 0.398f
C3859 VV10.n9 GND 0.36f
C3860 VV10.n10 GND 0.93f
C3861 VV11.t16 GND 0.0137f
C3862 VV11.n0 GND 0.112f
C3863 VV11.n1 GND 0.0544f
C3864 VV11.t11 GND 0.179f
C3865 VV11.t9 GND 0.179f
C3866 VV11.t5 GND 0.179f
C3867 VV11.t3 GND 0.179f
C3868 VV11.t0 GND 0.179f
C3869 VV11.t10 GND 0.179f
C3870 VV11.t14 GND 0.179f
C3871 VV11.t1 GND 0.179f
C3872 VV11.t8 GND 0.179f
C3873 VV11.t6 GND 0.179f
C3874 VV11.t13 GND 0.179f
C3875 VV11.t12 GND 0.179f
C3876 VV11.t2 GND 0.179f
C3877 VV11.t4 GND 0.179f
C3878 VV11.t7 GND 0.179f
C3879 VV11.t15 GND 0.387f
C3880 VV11.n2 GND 0.222f
C3881 VV11.n3 GND 0.22f
C3882 VV11.n4 GND 0.22f
C3883 VV11.n5 GND 0.22f
C3884 VV11.n6 GND 0.22f
C3885 VV11.n7 GND 0.22f
C3886 VV11.n8 GND 0.22f
C3887 VV11.n9 GND 0.22f
C3888 VV11.n10 GND 0.22f
C3889 VV11.n11 GND 0.22f
C3890 VV11.n12 GND 0.22f
C3891 VV11.n13 GND 0.22f
C3892 VV11.n14 GND 0.22f
C3893 VV11.n15 GND 0.22f
C3894 VV11.n16 GND 0.178f
C3895 VV11.n17 GND 1.12f
C3896 frontAnalog_v0p0p1_5.RSfetsym_0.QN.n0 GND 0.993f
C3897 frontAnalog_v0p0p1_5.RSfetsym_0.QN.t6 GND 0.0317f
C3898 frontAnalog_v0p0p1_5.RSfetsym_0.QN.t5 GND 0.0933f
C3899 frontAnalog_v0p0p1_5.RSfetsym_0.QN.n1 GND 1.47f
C3900 frontAnalog_v0p0p1_5.RSfetsym_0.QN.n2 GND 0.587f
C3901 frontAnalog_v0p0p1_5.RSfetsym_0.QN.t0 GND 0.0363f
C3902 frontAnalog_v0p0p1_5.RSfetsym_0.QN.n3 GND 0.622f
C3903 frontAnalog_v0p0p1_5.RSfetsym_0.QN.t3 GND 0.0317f
C3904 frontAnalog_v0p0p1_5.RSfetsym_0.QN.t2 GND 0.0317f
C3905 frontAnalog_v0p0p1_5.RSfetsym_0.QN.t1 GND 0.0558f
C3906 S1.t5 GND 0.0307f
C3907 S1.t0 GND 0.136f
C3908 S1.t6 GND 0.212f
C3909 S1.n0 GND 1.33f
C3910 S1.n1 GND 0.867f
C3911 S1.t3 GND 0.447f
C3912 S1.t2 GND 0.0187f
C3913 S1.n2 GND 1.54f
C3914 S1.n3 GND 1.92f
C3915 S1.t7 GND 0.027f
C3916 S1.t4 GND 0.0168f
C3917 S1.n4 GND 0.0548f
C3918 S1.n5 GND 0.0446f
C3919 S1.n6 GND 0.0337f
C3920 S1.t1 GND 0.144f
C3921 S1.n7 GND 0.206f
C3922 S1.n8 GND 0.613f
C3923 S1.n9 GND 0.661f
C3924 R1.t1 GND 0.145f
C3925 R1.t5 GND 0.0135f
C3926 R1.t7 GND 0.0217f
C3927 R1.n0 GND 0.0449f
C3928 R1.n1 GND 0.0354f
C3929 R1.n2 GND 0.0299f
C3930 R1.n3 GND 0.353f
C3931 R1.t4 GND 0.0246f
C3932 R1.t0 GND 0.167f
C3933 R1.t6 GND 0.169f
C3934 R1.n4 GND 0.964f
C3935 R1.n5 GND 0.919f
C3936 R1.t2 GND 0.015f
C3937 R1.t3 GND 0.323f
C3938 R1.n6 GND 1.28f
C3939 R1.n7 GND 0.859f
C3940 R1.n8 GND 1.26f
C3941 R1.n9 GND 0.181f
C3942 VV3.t16 GND 0.016f
C3943 VV3.n0 GND 0.131f
C3944 VV3.n1 GND 0.0634f
C3945 VV3.t5 GND 0.209f
C3946 VV3.t1 GND 0.209f
C3947 VV3.t13 GND 0.209f
C3948 VV3.t6 GND 0.209f
C3949 VV3.t15 GND 0.209f
C3950 VV3.t10 GND 0.209f
C3951 VV3.t0 GND 0.209f
C3952 VV3.t3 GND 0.209f
C3953 VV3.t8 GND 0.209f
C3954 VV3.t12 GND 0.209f
C3955 VV3.t2 GND 0.209f
C3956 VV3.t7 GND 0.209f
C3957 VV3.t11 GND 0.209f
C3958 VV3.t9 GND 0.209f
C3959 VV3.t4 GND 0.209f
C3960 VV3.t14 GND 0.451f
C3961 VV3.n2 GND 0.259f
C3962 VV3.n3 GND 0.257f
C3963 VV3.n4 GND 0.257f
C3964 VV3.n5 GND 0.257f
C3965 VV3.n6 GND 0.257f
C3966 VV3.n7 GND 0.257f
C3967 VV3.n8 GND 0.257f
C3968 VV3.n9 GND 0.257f
C3969 VV3.n10 GND 0.257f
C3970 VV3.n11 GND 0.257f
C3971 VV3.n12 GND 0.257f
C3972 VV3.n13 GND 0.257f
C3973 VV3.n14 GND 0.257f
C3974 VV3.n15 GND 0.257f
C3975 VV3.n16 GND 0.203f
C3976 VV3.n17 GND 1.53f
C3977 VV4.t16 GND 0.0164f
C3978 VV4.n0 GND 0.135f
C3979 VV4.n1 GND 0.0652f
C3980 VV4.t15 GND 0.215f
C3981 VV4.t0 GND 0.215f
C3982 VV4.t4 GND 0.215f
C3983 VV4.t6 GND 0.215f
C3984 VV4.t14 GND 0.215f
C3985 VV4.t10 GND 0.215f
C3986 VV4.t2 GND 0.215f
C3987 VV4.t3 GND 0.215f
C3988 VV4.t11 GND 0.215f
C3989 VV4.t12 GND 0.215f
C3990 VV4.t7 GND 0.215f
C3991 VV4.t8 GND 0.215f
C3992 VV4.t1 GND 0.215f
C3993 VV4.t9 GND 0.215f
C3994 VV4.t13 GND 0.215f
C3995 VV4.t5 GND 0.215f
C3996 VV4.n2 GND 0.515f
C3997 VV4.n3 GND 0.528f
C3998 VV4.n4 GND 0.528f
C3999 VV4.n5 GND 0.528f
C4000 VV4.n6 GND 0.528f
C4001 VV4.n7 GND 0.528f
C4002 VV4.n8 GND 0.528f
C4003 VV4.n9 GND 0.475f
C4004 VV4.n10 GND 1.48f
C4005 frontAnalog_v0p0p1_10.x65.A.n0 GND 0.139f
C4006 frontAnalog_v0p0p1_10.x65.A.t4 GND 0.028f
C4007 frontAnalog_v0p0p1_10.x65.A.t6 GND 0.0175f
C4008 frontAnalog_v0p0p1_10.x65.A.n1 GND 0.0568f
C4009 frontAnalog_v0p0p1_10.x65.A.t7 GND 0.0318f
C4010 frontAnalog_v0p0p1_10.x65.A.t1 GND 0.141f
C4011 frontAnalog_v0p0p1_10.x65.A.t5 GND 0.219f
C4012 frontAnalog_v0p0p1_10.x65.A.n2 GND 1.37f
C4013 frontAnalog_v0p0p1_10.x65.A.n3 GND 0.898f
C4014 frontAnalog_v0p0p1_10.x65.A.t2 GND 0.463f
C4015 frontAnalog_v0p0p1_10.x65.A.t3 GND 0.0194f
C4016 frontAnalog_v0p0p1_10.x65.A.n4 GND 1.6f
C4017 frontAnalog_v0p0p1_10.x65.A.n5 GND 2.01f
C4018 frontAnalog_v0p0p1_10.x65.A.t0 GND 0.149f
C4019 frontAnalog_v0p0p1_10.x65.A.n6 GND 1.72f
C4020 CLK.n0 GND 0.0667f
C4021 CLK.t23 GND 0.0549f
C4022 CLK.t89 GND 0.318f
C4023 CLK.t85 GND 0.321f
C4024 CLK.t26 GND 0.0578f
C4025 CLK.n1 GND 0.453f
C4026 CLK.n3 GND 0.28f
C4027 CLK.n5 GND 0.0661f
C4028 CLK.t94 GND 0.092f
C4029 CLK.n6 GND 0.386f
C4030 CLK.n7 GND 0.352f
C4031 CLK.n8 GND 0.156f
C4032 CLK.n9 GND 5.21f
C4033 CLK.n10 GND 0.0667f
C4034 CLK.t58 GND 0.0549f
C4035 CLK.t63 GND 0.318f
C4036 CLK.t14 GND 0.321f
C4037 CLK.t92 GND 0.0578f
C4038 CLK.n11 GND 0.453f
C4039 CLK.n13 GND 0.28f
C4040 CLK.n15 GND 0.0661f
C4041 CLK.t15 GND 0.092f
C4042 CLK.n16 GND 0.386f
C4043 CLK.n17 GND 0.352f
C4044 CLK.n18 GND 0.156f
C4045 CLK.n19 GND 0.0667f
C4046 CLK.t17 GND 0.0549f
C4047 CLK.t27 GND 0.318f
C4048 CLK.t73 GND 0.321f
C4049 CLK.t11 GND 0.0578f
C4050 CLK.n20 GND 0.453f
C4051 CLK.n22 GND 0.28f
C4052 CLK.n24 GND 0.0661f
C4053 CLK.t32 GND 0.092f
C4054 CLK.n25 GND 0.386f
C4055 CLK.n26 GND 0.352f
C4056 CLK.n27 GND 0.156f
C4057 CLK.n28 GND 0.0667f
C4058 CLK.t35 GND 0.0549f
C4059 CLK.t38 GND 0.318f
C4060 CLK.t90 GND 0.321f
C4061 CLK.t66 GND 0.0578f
C4062 CLK.n29 GND 0.453f
C4063 CLK.n31 GND 0.28f
C4064 CLK.n33 GND 0.0661f
C4065 CLK.t91 GND 0.092f
C4066 CLK.n34 GND 0.386f
C4067 CLK.n35 GND 0.352f
C4068 CLK.n36 GND 0.156f
C4069 CLK.n37 GND 0.0667f
C4070 CLK.t45 GND 0.0549f
C4071 CLK.t5 GND 0.318f
C4072 CLK.t47 GND 0.321f
C4073 CLK.t83 GND 0.0578f
C4074 CLK.n38 GND 0.453f
C4075 CLK.n40 GND 0.28f
C4076 CLK.n42 GND 0.0661f
C4077 CLK.t10 GND 0.092f
C4078 CLK.n43 GND 0.386f
C4079 CLK.n44 GND 0.352f
C4080 CLK.n45 GND 0.156f
C4081 CLK.n46 GND 0.0667f
C4082 CLK.t4 GND 0.0549f
C4083 CLK.t18 GND 0.318f
C4084 CLK.t64 GND 0.321f
C4085 CLK.t41 GND 0.0578f
C4086 CLK.n47 GND 0.453f
C4087 CLK.n49 GND 0.28f
C4088 CLK.n51 GND 0.0661f
C4089 CLK.t65 GND 0.092f
C4090 CLK.n52 GND 0.386f
C4091 CLK.n53 GND 0.352f
C4092 CLK.n54 GND 0.156f
C4093 CLK.n55 GND 0.0667f
C4094 CLK.t25 GND 0.0549f
C4095 CLK.t71 GND 0.318f
C4096 CLK.t74 GND 0.321f
C4097 CLK.t54 GND 0.0578f
C4098 CLK.n56 GND 0.453f
C4099 CLK.n58 GND 0.28f
C4100 CLK.n60 GND 0.0661f
C4101 CLK.t76 GND 0.092f
C4102 CLK.n61 GND 0.386f
C4103 CLK.n62 GND 0.352f
C4104 CLK.n63 GND 0.156f
C4105 CLK.n64 GND 0.0667f
C4106 CLK.t79 GND 0.0549f
C4107 CLK.t95 GND 0.318f
C4108 CLK.t39 GND 0.321f
C4109 CLK.t20 GND 0.0578f
C4110 CLK.n65 GND 0.453f
C4111 CLK.n67 GND 0.28f
C4112 CLK.n69 GND 0.0661f
C4113 CLK.t40 GND 0.092f
C4114 CLK.n70 GND 0.386f
C4115 CLK.n71 GND 0.352f
C4116 CLK.n72 GND 0.156f
C4117 CLK.n73 GND 0.0667f
C4118 CLK.t2 GND 0.0549f
C4119 CLK.t6 GND 0.318f
C4120 CLK.t51 GND 0.321f
C4121 CLK.t30 GND 0.0578f
C4122 CLK.n74 GND 0.453f
C4123 CLK.n76 GND 0.28f
C4124 CLK.n78 GND 0.0661f
C4125 CLK.t53 GND 0.092f
C4126 CLK.n79 GND 0.386f
C4127 CLK.n80 GND 0.352f
C4128 CLK.n81 GND 0.156f
C4129 CLK.n82 GND 0.0667f
C4130 CLK.t56 GND 0.0549f
C4131 CLK.t70 GND 0.318f
C4132 CLK.t13 GND 0.321f
C4133 CLK.t0 GND 0.0578f
C4134 CLK.n83 GND 0.453f
C4135 CLK.n85 GND 0.28f
C4136 CLK.n87 GND 0.0661f
C4137 CLK.t19 GND 0.092f
C4138 CLK.n88 GND 0.386f
C4139 CLK.n89 GND 0.352f
C4140 CLK.n90 GND 0.156f
C4141 CLK.n91 GND 0.0667f
C4142 CLK.t69 GND 0.0549f
C4143 CLK.t80 GND 0.318f
C4144 CLK.t28 GND 0.321f
C4145 CLK.t9 GND 0.0578f
C4146 CLK.n92 GND 0.453f
C4147 CLK.n94 GND 0.28f
C4148 CLK.n96 GND 0.0661f
C4149 CLK.t29 GND 0.092f
C4150 CLK.n97 GND 0.386f
C4151 CLK.n98 GND 0.352f
C4152 CLK.n99 GND 0.156f
C4153 CLK.n100 GND 0.0667f
C4154 CLK.t33 GND 0.0549f
C4155 CLK.t36 GND 0.318f
C4156 CLK.t87 GND 0.321f
C4157 CLK.t62 GND 0.0578f
C4158 CLK.n101 GND 0.453f
C4159 CLK.n103 GND 0.28f
C4160 CLK.n105 GND 0.0661f
C4161 CLK.t88 GND 0.092f
C4162 CLK.n106 GND 0.386f
C4163 CLK.n107 GND 0.352f
C4164 CLK.n108 GND 0.156f
C4165 CLK.n109 GND 0.0667f
C4166 CLK.t44 GND 0.0549f
C4167 CLK.t57 GND 0.318f
C4168 CLK.t7 GND 0.321f
C4169 CLK.t82 GND 0.0578f
C4170 CLK.n110 GND 0.453f
C4171 CLK.n112 GND 0.28f
C4172 CLK.n114 GND 0.0661f
C4173 CLK.t8 GND 0.092f
C4174 CLK.n115 GND 0.386f
C4175 CLK.n116 GND 0.352f
C4176 CLK.n117 GND 0.156f
C4177 CLK.n118 GND 0.0667f
C4178 CLK.t12 GND 0.0549f
C4179 CLK.t16 GND 0.318f
C4180 CLK.t60 GND 0.321f
C4181 CLK.t37 GND 0.0578f
C4182 CLK.n119 GND 0.453f
C4183 CLK.n121 GND 0.28f
C4184 CLK.n123 GND 0.0661f
C4185 CLK.t61 GND 0.092f
C4186 CLK.n124 GND 0.386f
C4187 CLK.n125 GND 0.352f
C4188 CLK.n126 GND 0.156f
C4189 CLK.n127 GND 0.0667f
C4190 CLK.t24 GND 0.0549f
C4191 CLK.t34 GND 0.318f
C4192 CLK.t72 GND 0.321f
C4193 CLK.t59 GND 0.0578f
C4194 CLK.n128 GND 0.453f
C4195 CLK.n130 GND 0.28f
C4196 CLK.n132 GND 0.0661f
C4197 CLK.t81 GND 0.092f
C4198 CLK.n133 GND 0.386f
C4199 CLK.n134 GND 0.352f
C4200 CLK.n135 GND 0.967f
C4201 CLK.n136 GND 6.67f
C4202 CLK.n137 GND 4.9f
C4203 CLK.n138 GND 4.9f
C4204 CLK.n139 GND 4.9f
C4205 CLK.n140 GND 4.9f
C4206 CLK.n141 GND 4.9f
C4207 CLK.n142 GND 4.9f
C4208 CLK.n143 GND 4.9f
C4209 CLK.n144 GND 4.9f
C4210 CLK.n145 GND 4.9f
C4211 CLK.n146 GND 4.9f
C4212 CLK.n147 GND 4.9f
C4213 CLK.n148 GND 4.9f
C4214 CLK.n149 GND 4.9f
C4215 CLK.t78 GND 0.0549f
C4216 CLK.t46 GND 0.318f
C4217 CLK.t48 GND 0.321f
C4218 CLK.t86 GND 0.0578f
C4219 CLK.n150 GND 0.453f
C4220 CLK.n152 GND 0.28f
C4221 CLK.n154 GND 0.0661f
C4222 CLK.t49 GND 0.092f
C4223 CLK.n155 GND 0.386f
C4224 CLK.n156 GND 0.352f
C4225 CLK.n157 GND 0.156f
C4226 CLK.n158 GND 0.0667f
C4227 a_16719_n13117.n0 GND 1.47f
C4228 a_16719_n13117.n1 GND 1.14f
C4229 a_16719_n13117.t8 GND 0.177f
C4230 a_16719_n13117.t18 GND 0.177f
C4231 a_16719_n13117.t22 GND 0.177f
C4232 a_16719_n13117.t11 GND 0.177f
C4233 a_16719_n13117.t16 GND 0.177f
C4234 a_16719_n13117.t5 GND 0.177f
C4235 a_16719_n13117.t20 GND 0.177f
C4236 a_16719_n13117.t14 GND 0.177f
C4237 a_16719_n13117.t7 GND 0.177f
C4238 a_16719_n13117.t15 GND 0.177f
C4239 a_16719_n13117.t4 GND 0.177f
C4240 a_16719_n13117.t19 GND 0.177f
C4241 a_16719_n13117.t12 GND 0.252f
C4242 a_16719_n13117.n2 GND 1.4f
C4243 a_16719_n13117.n3 GND 0.768f
C4244 a_16719_n13117.n4 GND 0.768f
C4245 a_16719_n13117.n5 GND 0.768f
C4246 a_16719_n13117.n6 GND 0.768f
C4247 a_16719_n13117.n7 GND 0.768f
C4248 a_16719_n13117.n8 GND 0.72f
C4249 a_16719_n13117.n9 GND 0.273f
C4250 a_16719_n13117.n10 GND 0.325f
C4251 a_16719_n13117.n11 GND 0.912f
C4252 a_16719_n13117.n12 GND 2.03f
C4253 a_16719_n13117.n13 GND 1.47f
C4254 a_16719_n13117.t1 GND 0.238f
C4255 a_16719_n13117.n14 GND 2.05f
C4256 a_16719_n13117.t24 GND 1.7f
C4257 a_16719_n13117.n15 GND 0.991f
C4258 a_16719_n13117.n16 GND 0.0433f
C4259 a_16719_n13117.n17 GND 0.426f
C4260 a_16719_n13117.t0 GND 1.7f
C4261 a_16719_n13117.t2 GND 0.0103f
C4262 a_16719_n13117.n18 GND 0.213f
C4263 a_16719_n13117.t25 GND 1.7f
C4264 a_16719_n13117.n19 GND 1.05f
C4265 a_16719_n13117.n20 GND 0.0503f
C4266 a_16719_n13117.n21 GND 0.0699f
C4267 a_16719_n13117.n22 GND 0.308f
C4268 a_16719_n13117.n23 GND 0.811f
C4269 a_16719_n13117.n24 GND 0.768f
C4270 a_16719_n13117.n25 GND 0.768f
C4271 a_16719_n13117.t9 GND 0.177f
C4272 a_16719_n13117.t17 GND 0.177f
C4273 a_16719_n13117.t21 GND 0.177f
C4274 a_16719_n13117.t13 GND 0.177f
C4275 a_16719_n13117.t6 GND 0.177f
C4276 a_16719_n13117.t10 GND 0.252f
C4277 a_16719_n13117.n26 GND 1.4f
C4278 a_16719_n13117.n27 GND 0.768f
C4279 a_16719_n13117.n28 GND 0.768f
C4280 a_16719_n13117.n29 GND 0.768f
C4281 a_16719_n13117.n30 GND 0.768f
C4282 a_16719_n13117.n31 GND 0.768f
C4283 a_16719_n13117.t23 GND 0.177f
C4284 a_16541_n13117.t10 GND 0.112f
C4285 a_16541_n13117.t17 GND 0.112f
C4286 a_16541_n13117.t6 GND 0.112f
C4287 a_16541_n13117.t2 GND 0.112f
C4288 a_16541_n13117.t13 GND 0.112f
C4289 a_16541_n13117.t21 GND 0.112f
C4290 a_16541_n13117.t12 GND 0.112f
C4291 a_16541_n13117.t3 GND 0.112f
C4292 a_16541_n13117.t7 GND 0.112f
C4293 a_16541_n13117.t15 GND 0.112f
C4294 a_16541_n13117.t20 GND 0.112f
C4295 a_16541_n13117.t9 GND 0.112f
C4296 a_16541_n13117.t5 GND 0.112f
C4297 a_16541_n13117.t18 GND 0.112f
C4298 a_16541_n13117.t11 GND 0.112f
C4299 a_16541_n13117.t19 GND 0.112f
C4300 a_16541_n13117.t8 GND 0.112f
C4301 a_16541_n13117.t4 GND 0.112f
C4302 a_16541_n13117.t16 GND 0.161f
C4303 a_16541_n13117.n0 GND 1.02f
C4304 a_16541_n13117.n1 GND 0.558f
C4305 a_16541_n13117.n2 GND 0.558f
C4306 a_16541_n13117.n3 GND 0.558f
C4307 a_16541_n13117.n4 GND 0.558f
C4308 a_16541_n13117.n5 GND 0.558f
C4309 a_16541_n13117.n6 GND 0.558f
C4310 a_16541_n13117.n7 GND 0.558f
C4311 a_16541_n13117.n8 GND 0.614f
C4312 a_16541_n13117.n9 GND 0.614f
C4313 a_16541_n13117.n10 GND 0.558f
C4314 a_16541_n13117.n11 GND 0.558f
C4315 a_16541_n13117.n12 GND 0.558f
C4316 a_16541_n13117.n13 GND 0.558f
C4317 a_16541_n13117.n14 GND 0.558f
C4318 a_16541_n13117.n15 GND 0.558f
C4319 a_16541_n13117.n16 GND 0.554f
C4320 a_16541_n13117.n17 GND 0.627f
C4321 a_16541_n13117.t14 GND 0.127f
C4322 a_16541_n13117.n18 GND 1.13f
C4323 a_16541_n13117.t1 GND 0.376f
C4324 a_16541_n13117.n19 GND 10.1f
C4325 a_16541_n13117.t0 GND 1.21f
C4326 a_16599_n13205.n0 GND 0.681f
C4327 a_16599_n13205.t15 GND 0.179f
C4328 a_16599_n13205.n1 GND 0.251f
C4329 a_16599_n13205.t8 GND 0.179f
C4330 a_16599_n13205.n2 GND 0.378f
C4331 a_16599_n13205.t23 GND 0.179f
C4332 a_16599_n13205.n3 GND 0.197f
C4333 a_16599_n13205.t12 GND 0.179f
C4334 a_16599_n13205.n4 GND 0.197f
C4335 a_16599_n13205.t20 GND 0.179f
C4336 a_16599_n13205.n5 GND 0.197f
C4337 a_16599_n13205.t13 GND 0.179f
C4338 a_16599_n13205.n6 GND 0.197f
C4339 a_16599_n13205.t7 GND 0.179f
C4340 a_16599_n13205.n7 GND 0.197f
C4341 a_16599_n13205.t22 GND 0.179f
C4342 a_16599_n13205.n8 GND 0.197f
C4343 a_16599_n13205.t11 GND 0.179f
C4344 a_16599_n13205.n9 GND 0.197f
C4345 a_16599_n13205.t16 GND 0.179f
C4346 a_16599_n13205.n10 GND 0.184f
C4347 a_16599_n13205.t2 GND 0.179f
C4348 a_16599_n13205.t5 GND 0.179f
C4349 a_16599_n13205.t9 GND 0.179f
C4350 a_16599_n13205.t19 GND 0.179f
C4351 a_16599_n13205.t4 GND 0.179f
C4352 a_16599_n13205.t18 GND 0.179f
C4353 a_16599_n13205.t10 GND 0.179f
C4354 a_16599_n13205.t6 GND 0.179f
C4355 a_16599_n13205.t14 GND 0.179f
C4356 a_16599_n13205.t21 GND 0.179f
C4357 a_16599_n13205.t17 GND 0.179f
C4358 a_16599_n13205.n11 GND 0.252f
C4359 a_16599_n13205.n12 GND 0.376f
C4360 a_16599_n13205.n13 GND 0.197f
C4361 a_16599_n13205.n14 GND 0.197f
C4362 a_16599_n13205.n15 GND 0.197f
C4363 a_16599_n13205.n16 GND 0.197f
C4364 a_16599_n13205.n17 GND 0.197f
C4365 a_16599_n13205.n18 GND 0.197f
C4366 a_16599_n13205.n19 GND 0.197f
C4367 a_16599_n13205.n20 GND 0.197f
C4368 a_16599_n13205.n21 GND 0.169f
C4369 a_16599_n13205.n22 GND 0.102f
C4370 a_16599_n13205.n23 GND 0.377f
C4371 a_16599_n13205.n24 GND 0.197f
C4372 a_16599_n13205.n25 GND 0.197f
C4373 a_16599_n13205.n26 GND 0.197f
C4374 a_16599_n13205.n27 GND 0.197f
C4375 a_16599_n13205.n28 GND 0.197f
C4376 a_16599_n13205.n29 GND 0.197f
C4377 a_16599_n13205.n30 GND 0.197f
C4378 a_16599_n13205.n31 GND 0.184f
C4379 a_16599_n13205.n32 GND 0.376f
C4380 a_16599_n13205.n33 GND 0.197f
C4381 a_16599_n13205.n34 GND 0.197f
C4382 a_16599_n13205.n35 GND 0.197f
C4383 a_16599_n13205.n36 GND 0.197f
C4384 a_16599_n13205.n37 GND 0.197f
C4385 a_16599_n13205.n38 GND 0.197f
C4386 a_16599_n13205.n39 GND 0.197f
C4387 a_16599_n13205.n40 GND 0.197f
C4388 a_16599_n13205.n41 GND 0.169f
C4389 a_16599_n13205.n42 GND 0.108f
C4390 a_16599_n13205.t3 GND 0.0381f
C4391 a_16599_n13205.n43 GND 2.83f
C4392 a_16599_n13205.t1 GND 1.94f
C4393 VV16.t16 GND 0.0172f
C4394 VV16.n0 GND 0.141f
C4395 VV16.n1 GND 0.0593f
C4396 VV16.t10 GND 0.225f
C4397 VV16.t1 GND 0.225f
C4398 VV16.t3 GND 0.225f
C4399 VV16.t2 GND 0.225f
C4400 VV16.t4 GND 0.225f
C4401 VV16.t0 GND 0.225f
C4402 VV16.t8 GND 0.225f
C4403 VV16.t7 GND 0.225f
C4404 VV16.t11 GND 0.225f
C4405 VV16.t5 GND 0.225f
C4406 VV16.t9 GND 0.225f
C4407 VV16.t15 GND 0.225f
C4408 VV16.t12 GND 0.225f
C4409 VV16.t14 GND 0.225f
C4410 VV16.t6 GND 0.225f
C4411 VV16.t13 GND 0.485f
C4412 VV16.n2 GND 0.279f
C4413 VV16.n3 GND 0.276f
C4414 VV16.n4 GND 0.276f
C4415 VV16.n5 GND 0.276f
C4416 VV16.n6 GND 0.276f
C4417 VV16.n7 GND 0.276f
C4418 VV16.n8 GND 0.276f
C4419 VV16.n9 GND 0.276f
C4420 VV16.n10 GND 0.276f
C4421 VV16.n11 GND 0.276f
C4422 VV16.n12 GND 0.276f
C4423 VV16.n13 GND 0.276f
C4424 VV16.n14 GND 0.276f
C4425 VV16.n15 GND 0.276f
C4426 VV16.n16 GND 0.224f
C4427 VV16.n17 GND 2.37f
C4428 VFS.t5 GND 0.108f
C4429 VFS.n0 GND 0.0961f
C4430 VFS.n1 GND 0.0961f
C4431 VFS.n2 GND 0.0687f
C4432 VFS.n3 GND 2.49f
C4433 VFS.t2 GND 0.0898f
C4434 VFS.n4 GND 0.0961f
C4435 VFS.n5 GND 0.0961f
C4436 VFS.n6 GND 0.0741f
C4437 OUT2.n2 GND 0.0114f
C4438 OUT2.n4 GND 0.0241f
C4439 OUT2.n6 GND 0.0161f
C4440 OUT2.n8 GND 0.0161f
C4441 OUT2.n10 GND 0.0161f
C4442 OUT2.n12 GND 0.0161f
C4443 OUT2.n14 GND 0.0161f
C4444 OUT2.n23 GND 0.014f
C4445 OUT2.n25 GND 0.0348f
C4446 OUT2.n27 GND 0.021f
C4447 OUT2.n29 GND 0.021f
C4448 OUT2.n31 GND 0.021f
C4449 OUT2.n33 GND 0.021f
C4450 OUT2.n35 GND 0.021f
C4451 OUT2.n37 GND 0.0147f
C4452 OUT2.n38 GND 0.0296f
C4453 OUT2.n39 GND 0.0229f
C4454 OUT2.n42 GND 0.0114f
C4455 OUT2.n44 GND 0.0241f
C4456 OUT2.n46 GND 0.0161f
C4457 OUT2.n48 GND 0.0161f
C4458 OUT2.n50 GND 0.0161f
C4459 OUT2.n52 GND 0.0161f
C4460 OUT2.n54 GND 0.0161f
C4461 OUT2.n63 GND 0.014f
C4462 OUT2.n65 GND 0.0348f
C4463 OUT2.n67 GND 0.021f
C4464 OUT2.n69 GND 0.021f
C4465 OUT2.n71 GND 0.021f
C4466 OUT2.n73 GND 0.021f
C4467 OUT2.n75 GND 0.021f
C4468 OUT2.n77 GND 0.0147f
C4469 OUT2.n78 GND 0.0273f
C4470 OUT2.n79 GND 0.0203f
C4471 OUT2.n81 GND 0.0114f
C4472 OUT2.n83 GND 0.0241f
C4473 OUT2.n85 GND 0.0161f
C4474 OUT2.n87 GND 0.0161f
C4475 OUT2.n89 GND 0.0161f
C4476 OUT2.n91 GND 0.0161f
C4477 OUT2.n93 GND 0.0161f
C4478 OUT2.n97 GND 0.0126f
C4479 OUT2.n100 GND 0.014f
C4480 OUT2.n102 GND 0.0348f
C4481 OUT2.n104 GND 0.021f
C4482 OUT2.n106 GND 0.021f
C4483 OUT2.n108 GND 0.021f
C4484 OUT2.n110 GND 0.021f
C4485 OUT2.n112 GND 0.021f
C4486 OUT2.n114 GND 0.0147f
C4487 OUT2.n115 GND 0.0284f
C4488 OUT2.n116 GND 0.0234f
C4489 OUT2.n120 GND 0.014f
C4490 OUT2.n122 GND 0.0348f
C4491 OUT2.n124 GND 0.021f
C4492 OUT2.n126 GND 0.021f
C4493 OUT2.n128 GND 0.021f
C4494 OUT2.n130 GND 0.021f
C4495 OUT2.n132 GND 0.021f
C4496 OUT2.n136 GND 0.0114f
C4497 OUT2.n138 GND 0.0241f
C4498 OUT2.n140 GND 0.0161f
C4499 OUT2.n142 GND 0.0161f
C4500 OUT2.n144 GND 0.0161f
C4501 OUT2.n146 GND 0.0161f
C4502 OUT2.n148 GND 0.0161f
C4503 OUT2.n152 GND 0.013f
C4504 OUT2.n155 GND 0.0204f
C4505 OUT2.n156 GND 0.108f
C4506 OUT2.n157 GND 0.275f
C4507 OUT2.n158 GND 0.224f
C4508 OUT2.n159 GND 0.228f
C4509 I5.t11 GND 0.0118f
C4510 I5.n3 GND 0.0129f
C4511 I5.n8 GND 0.144f
C4512 I5.n9 GND 0.36f
C4513 I5.n12 GND 0.011f
C4514 I5.n16 GND 0.205f
C4515 I5.n21 GND 0.545f
C4516 I5.n22 GND 1.29f
C4517 I5.n23 GND 0.293f
C4518 I5.n24 GND 0.66f
C4519 I5.n25 GND 1.24f
C4520 I5.t12 GND 0.0265f
C4521 I5.n26 GND 0.416f
C4522 I5.n27 GND 0.0551f
C4523 I5.n28 GND 0.125f
C4524 I5.n29 GND 0.0829f
C4525 I5.n30 GND 0.0886f
C4526 I5.n31 GND 0.122f
C4527 I5.n32 GND 0.116f
C4528 I5.n33 GND 0.266f
C4529 I5.n34 GND 9.98f
C4530 I5.n35 GND 2.07f
C4531 OUT0.n2 GND 0.0114f
C4532 OUT0.n4 GND 0.0241f
C4533 OUT0.n6 GND 0.0161f
C4534 OUT0.n8 GND 0.0161f
C4535 OUT0.n10 GND 0.0161f
C4536 OUT0.n12 GND 0.0161f
C4537 OUT0.n14 GND 0.0161f
C4538 OUT0.n23 GND 0.014f
C4539 OUT0.n25 GND 0.0348f
C4540 OUT0.n27 GND 0.021f
C4541 OUT0.n29 GND 0.021f
C4542 OUT0.n31 GND 0.021f
C4543 OUT0.n33 GND 0.021f
C4544 OUT0.n35 GND 0.021f
C4545 OUT0.n37 GND 0.0147f
C4546 OUT0.n38 GND 0.0296f
C4547 OUT0.n39 GND 0.0229f
C4548 OUT0.n42 GND 0.0114f
C4549 OUT0.n44 GND 0.0241f
C4550 OUT0.n46 GND 0.0161f
C4551 OUT0.n48 GND 0.0161f
C4552 OUT0.n50 GND 0.0161f
C4553 OUT0.n52 GND 0.0161f
C4554 OUT0.n54 GND 0.0161f
C4555 OUT0.n63 GND 0.014f
C4556 OUT0.n65 GND 0.0348f
C4557 OUT0.n67 GND 0.021f
C4558 OUT0.n69 GND 0.021f
C4559 OUT0.n71 GND 0.021f
C4560 OUT0.n73 GND 0.021f
C4561 OUT0.n75 GND 0.021f
C4562 OUT0.n77 GND 0.0147f
C4563 OUT0.n78 GND 0.0273f
C4564 OUT0.n79 GND 0.0203f
C4565 OUT0.n81 GND 0.0114f
C4566 OUT0.n83 GND 0.0241f
C4567 OUT0.n85 GND 0.0161f
C4568 OUT0.n87 GND 0.0161f
C4569 OUT0.n89 GND 0.0161f
C4570 OUT0.n91 GND 0.0161f
C4571 OUT0.n93 GND 0.0161f
C4572 OUT0.n97 GND 0.0126f
C4573 OUT0.n100 GND 0.014f
C4574 OUT0.n102 GND 0.0348f
C4575 OUT0.n104 GND 0.021f
C4576 OUT0.n106 GND 0.021f
C4577 OUT0.n108 GND 0.021f
C4578 OUT0.n110 GND 0.021f
C4579 OUT0.n112 GND 0.021f
C4580 OUT0.n114 GND 0.0147f
C4581 OUT0.n115 GND 0.0284f
C4582 OUT0.n116 GND 0.0234f
C4583 OUT0.n120 GND 0.014f
C4584 OUT0.n122 GND 0.0348f
C4585 OUT0.n124 GND 0.021f
C4586 OUT0.n126 GND 0.021f
C4587 OUT0.n128 GND 0.021f
C4588 OUT0.n130 GND 0.021f
C4589 OUT0.n132 GND 0.021f
C4590 OUT0.n136 GND 0.0114f
C4591 OUT0.n138 GND 0.0241f
C4592 OUT0.n140 GND 0.0161f
C4593 OUT0.n142 GND 0.0161f
C4594 OUT0.n144 GND 0.0161f
C4595 OUT0.n146 GND 0.0161f
C4596 OUT0.n148 GND 0.0161f
C4597 OUT0.n152 GND 0.013f
C4598 OUT0.n155 GND 0.0204f
C4599 OUT0.n156 GND 0.108f
C4600 OUT0.n157 GND 0.275f
C4601 OUT0.n158 GND 0.224f
C4602 OUT0.n159 GND 0.228f
C4603 R0.t2 GND 0.146f
C4604 R0.t6 GND 0.0136f
C4605 R0.t4 GND 0.0218f
C4606 R0.n0 GND 0.0451f
C4607 R0.n1 GND 0.0356f
C4608 R0.n2 GND 0.0301f
C4609 R0.n3 GND 0.3f
C4610 R0.t5 GND 0.0248f
C4611 R0.t3 GND 0.168f
C4612 R0.t7 GND 0.17f
C4613 R0.n4 GND 0.969f
C4614 R0.n5 GND 0.924f
C4615 R0.t1 GND 0.0151f
C4616 R0.t0 GND 0.324f
C4617 R0.n6 GND 1.29f
C4618 R0.n7 GND 0.864f
C4619 R0.n8 GND 1.24f
C4620 R0.n9 GND 0.133f
C4621 OUT3.n5 GND 0.0122f
C4622 OUT3.n7 GND 0.0305f
C4623 OUT3.n9 GND 0.0184f
C4624 OUT3.n11 GND 0.0184f
C4625 OUT3.n13 GND 0.0184f
C4626 OUT3.n15 GND 0.0184f
C4627 OUT3.n17 GND 0.0184f
C4628 OUT3.n26 GND 0.0212f
C4629 OUT3.n28 GND 0.0141f
C4630 OUT3.n30 GND 0.0141f
C4631 OUT3.n32 GND 0.0141f
C4632 OUT3.n34 GND 0.0141f
C4633 OUT3.n36 GND 0.0141f
C4634 OUT3.n44 GND 0.027f
C4635 OUT3.n45 GND 0.0219f
C4636 OUT3.n51 GND 0.0122f
C4637 OUT3.n53 GND 0.0305f
C4638 OUT3.n55 GND 0.0184f
C4639 OUT3.n57 GND 0.0184f
C4640 OUT3.n59 GND 0.0184f
C4641 OUT3.n61 GND 0.0184f
C4642 OUT3.n63 GND 0.0184f
C4643 OUT3.n66 GND 0.0157f
C4644 OUT3.n72 GND 0.0212f
C4645 OUT3.n74 GND 0.0141f
C4646 OUT3.n76 GND 0.0141f
C4647 OUT3.n78 GND 0.0141f
C4648 OUT3.n80 GND 0.0141f
C4649 OUT3.n82 GND 0.0141f
C4650 OUT3.n85 GND 0.015f
C4651 OUT3.n86 GND 0.0477f
C4652 OUT3.n87 GND 0.0111f
C4653 OUT3.n89 GND 0.0122f
C4654 OUT3.n91 GND 0.0305f
C4655 OUT3.n93 GND 0.0184f
C4656 OUT3.n95 GND 0.0184f
C4657 OUT3.n97 GND 0.0184f
C4658 OUT3.n99 GND 0.0184f
C4659 OUT3.n101 GND 0.0184f
C4660 OUT3.n114 GND 0.0212f
C4661 OUT3.n116 GND 0.0141f
C4662 OUT3.n118 GND 0.0141f
C4663 OUT3.n120 GND 0.0141f
C4664 OUT3.n122 GND 0.0141f
C4665 OUT3.n124 GND 0.0141f
C4666 OUT3.n133 GND 0.0282f
C4667 OUT3.n134 GND 0.0213f
C4668 OUT3.n140 GND 0.0122f
C4669 OUT3.n142 GND 0.0305f
C4670 OUT3.n144 GND 0.0184f
C4671 OUT3.n146 GND 0.0184f
C4672 OUT3.n148 GND 0.0184f
C4673 OUT3.n150 GND 0.0184f
C4674 OUT3.n152 GND 0.0184f
C4675 OUT3.n160 GND 0.0212f
C4676 OUT3.n162 GND 0.0141f
C4677 OUT3.n164 GND 0.0141f
C4678 OUT3.n166 GND 0.0141f
C4679 OUT3.n168 GND 0.0141f
C4680 OUT3.n170 GND 0.0141f
C4681 OUT3.n179 GND 0.027f
C4682 OUT3.n180 GND 0.119f
C4683 OUT3.n181 GND 0.304f
C4684 OUT3.n182 GND 0.264f
C4685 OUT3.n183 GND 0.577f
C4686 VDD.t336 GND 0.0102f
C4687 VDD.t1247 GND 0.0213f
C4688 VDD.t696 GND 0.0367f
C4689 VDD.t200 GND 0.0151f
C4690 VDD.t1281 GND 0.0158f
C4691 VDD.t1467 GND 0.0158f
C4692 VDD.t17 GND 0.0183f
C4693 VDD.t1282 GND 0.0297f
C4694 VDD.n0 GND 0.0145f
C4695 VDD.n26 GND 0.0234f
C4696 VDD.n34 GND 0.0903f
C4697 VDD.n35 GND 0.283f
C4698 VDD.n37 GND 0.013f
C4699 VDD.n40 GND 0.0109f
C4700 VDD.n43 GND 0.0109f
C4701 VDD.n50 GND 0.0253f
C4702 VDD.t963 GND 0.0318f
C4703 VDD.t989 GND 0.0138f
C4704 VDD.t947 GND 0.0138f
C4705 VDD.t967 GND 0.0138f
C4706 VDD.t959 GND 0.0138f
C4707 VDD.n53 GND 0.0163f
C4708 VDD.n55 GND 0.102f
C4709 VDD.n59 GND 0.0233f
C4710 VDD.n60 GND 0.0137f
C4711 VDD.n66 GND 0.0257f
C4712 VDD.n70 GND 0.0257f
C4713 VDD.n72 GND 0.0257f
C4714 VDD.n73 GND 0.0193f
C4715 VDD.n74 GND 0.0152f
C4716 VDD.n76 GND 0.0257f
C4717 VDD.n80 GND 0.0257f
C4718 VDD.n82 GND 0.0257f
C4719 VDD.n86 GND 0.0257f
C4720 VDD.n88 GND 0.0257f
C4721 VDD.n92 GND 0.0257f
C4722 VDD.n94 GND 0.0257f
C4723 VDD.n98 GND 0.0214f
C4724 VDD.n99 GND 0.0137f
C4725 VDD.n104 GND 0.0128f
C4726 VDD.n105 GND 0.0109f
C4727 VDD.n106 GND 0.0112f
C4728 VDD.t1007 GND 0.011f
C4729 VDD.t949 GND 0.0138f
C4730 VDD.t985 GND 0.0138f
C4731 VDD.t927 GND 0.0138f
C4732 VDD.t951 GND 0.0138f
C4733 VDD.t975 GND 0.0138f
C4734 VDD.t1039 GND 0.0138f
C4735 VDD.t941 GND 0.0138f
C4736 VDD.t1001 GND 0.0138f
C4737 VDD.t1045 GND 0.0133f
C4738 VDD.t965 GND 0.0179f
C4739 VDD.t1015 GND 0.0138f
C4740 VDD.t931 GND 0.0138f
C4741 VDD.t957 GND 0.0138f
C4742 VDD.t1013 GND 0.0115f
C4743 VDD.t935 GND 0.0138f
C4744 VDD.t977 GND 0.0138f
C4745 VDD.t1041 GND 0.0138f
C4746 VDD.t1011 GND 0.0138f
C4747 VDD.t953 GND 0.0179f
C4748 VDD.t1031 GND 0.0133f
C4749 VDD.t1005 GND 0.0138f
C4750 VDD.t945 GND 0.0138f
C4751 VDD.t1027 GND 0.0138f
C4752 VDD.t999 GND 0.0138f
C4753 VDD.t939 GND 0.0138f
C4754 VDD.t987 GND 0.0138f
C4755 VDD.t1051 GND 0.0138f
C4756 VDD.t1019 GND 0.0138f
C4757 VDD.t981 GND 0.0138f
C4758 VDD.n107 GND 0.0112f
C4759 VDD.n108 GND 0.0109f
C4760 VDD.n111 GND 0.013f
C4761 VDD.n112 GND 0.0137f
C4762 VDD.n116 GND 0.0172f
C4763 VDD.n120 GND 0.0257f
C4764 VDD.n122 GND 0.0257f
C4765 VDD.n126 GND 0.0257f
C4766 VDD.n128 GND 0.0257f
C4767 VDD.n132 GND 0.0257f
C4768 VDD.n134 GND 0.0257f
C4769 VDD.n138 GND 0.0257f
C4770 VDD.n140 GND 0.0257f
C4771 VDD.n141 GND 0.0152f
C4772 VDD.n144 GND 0.0193f
C4773 VDD.n146 GND 0.0257f
C4774 VDD.n150 GND 0.0257f
C4775 VDD.n152 GND 0.0257f
C4776 VDD.n156 GND 0.0214f
C4777 VDD.n157 GND 0.0137f
C4778 VDD.n163 GND 0.0257f
C4779 VDD.n165 GND 0.0257f
C4780 VDD.n169 GND 0.0257f
C4781 VDD.n171 GND 0.0257f
C4782 VDD.n175 GND 0.0257f
C4783 VDD.n177 GND 0.0257f
C4784 VDD.n181 GND 0.0233f
C4785 VDD.n182 GND 0.0137f
C4786 VDD.n187 GND 0.0128f
C4787 VDD.n188 GND 0.0109f
C4788 VDD.n189 GND 0.0112f
C4789 VDD.t1037 GND 0.0122f
C4790 VDD.t937 GND 0.0138f
C4791 VDD.t995 GND 0.0138f
C4792 VDD.t1023 GND 0.0138f
C4793 VDD.t1053 GND 0.0138f
C4794 VDD.t997 GND 0.0138f
C4795 VDD.t1025 GND 0.0138f
C4796 VDD.t969 GND 0.0138f
C4797 VDD.t991 GND 0.0138f
C4798 VDD.t1009 GND 0.0133f
C4799 VDD.t1033 GND 0.0179f
C4800 VDD.t929 GND 0.0138f
C4801 VDD.t955 GND 0.0138f
C4802 VDD.n190 GND 0.0112f
C4803 VDD.t933 GND 0.0133f
C4804 VDD.t993 GND 0.0138f
C4805 VDD.t1017 GND 0.0138f
C4806 VDD.t1049 GND 0.0138f
C4807 VDD.t983 GND 0.0138f
C4808 VDD.t1021 GND 0.0138f
C4809 VDD.t961 GND 0.0138f
C4810 VDD.t1043 GND 0.0138f
C4811 VDD.t943 GND 0.0138f
C4812 VDD.t1003 GND 0.0138f
C4813 VDD.t1029 GND 0.0138f
C4814 VDD.t971 GND 0.0133f
C4815 VDD.t1486 GND 0.0179f
C4816 VDD.t1468 GND 0.0137f
C4817 VDD.n191 GND 0.0112f
C4818 VDD.t1488 GND 0.0138f
C4819 VDD.t1498 GND 0.0138f
C4820 VDD.t1494 GND 0.0138f
C4821 VDD.t1470 GND 0.0138f
C4822 VDD.t1482 GND 0.0138f
C4823 VDD.t1496 GND 0.0138f
C4824 VDD.t1472 GND 0.0138f
C4825 VDD.t1484 GND 0.0138f
C4826 VDD.t1490 GND 0.0138f
C4827 VDD.t1474 GND 0.0138f
C4828 VDD.t1478 GND 0.0138f
C4829 VDD.t1492 GND 0.0138f
C4830 VDD.t1476 GND 0.0133f
C4831 VDD.t64 GND 0.0178f
C4832 VDD.t66 GND 0.0138f
C4833 VDD.t60 GND 0.0138f
C4834 VDD.t62 GND 0.0131f
C4835 VDD.t1255 GND 0.0146f
C4836 VDD.t391 GND 0.0139f
C4837 VDD.t1057 GND 0.0232f
C4838 VDD.t50 GND 0.0171f
C4839 VDD.n192 GND 0.0182f
C4840 VDD.n196 GND 0.0384f
C4841 VDD.n198 GND 0.0299f
C4842 VDD.n199 GND 0.0193f
C4843 VDD.n202 GND 0.0152f
C4844 VDD.n204 GND 0.0169f
C4845 VDD.n205 GND 0.0137f
C4846 VDD.n209 GND 0.0109f
C4847 VDD.n211 GND 0.0149f
C4848 VDD.n213 GND 0.0257f
C4849 VDD.n216 GND 0.0257f
C4850 VDD.n218 GND 0.0257f
C4851 VDD.n219 GND 0.0193f
C4852 VDD.n220 GND 0.0152f
C4853 VDD.n222 GND 0.0257f
C4854 VDD.n226 GND 0.0257f
C4855 VDD.n228 GND 0.0257f
C4856 VDD.n232 GND 0.0257f
C4857 VDD.n234 GND 0.0257f
C4858 VDD.n238 GND 0.0257f
C4859 VDD.n240 GND 0.0257f
C4860 VDD.n244 GND 0.0257f
C4861 VDD.n248 GND 0.0257f
C4862 VDD.n250 GND 0.0257f
C4863 VDD.n254 GND 0.023f
C4864 VDD.n255 GND 0.0137f
C4865 VDD.n258 GND 0.0128f
C4866 VDD.n263 GND 0.0137f
C4867 VDD.n265 GND 0.0216f
C4868 VDD.n266 GND 0.0193f
C4869 VDD.n267 GND 0.0152f
C4870 VDD.n269 GND 0.0257f
C4871 VDD.n273 GND 0.0257f
C4872 VDD.n275 GND 0.0257f
C4873 VDD.n279 GND 0.0257f
C4874 VDD.n281 GND 0.0257f
C4875 VDD.n285 GND 0.0257f
C4876 VDD.n287 GND 0.0257f
C4877 VDD.n291 GND 0.0257f
C4878 VDD.n295 GND 0.0257f
C4879 VDD.n297 GND 0.023f
C4880 VDD.n298 GND 0.0137f
C4881 VDD.n303 GND 0.0128f
C4882 VDD.n306 GND 0.0137f
C4883 VDD.n310 GND 0.0216f
C4884 VDD.n312 GND 0.0257f
C4885 VDD.n313 GND 0.0193f
C4886 VDD.n314 GND 0.0151f
C4887 VDD.n315 GND 10f
C4888 VDD.n316 GND 2.42f
C4889 VDD.t766 GND 0.0102f
C4890 VDD.t1180 GND 0.0213f
C4891 VDD.t135 GND 0.0367f
C4892 VDD.t798 GND 0.0151f
C4893 VDD.t167 GND 0.0158f
C4894 VDD.t409 GND 0.0158f
C4895 VDD.t1324 GND 0.0183f
C4896 VDD.t1326 GND 0.0297f
C4897 VDD.n317 GND 0.0145f
C4898 VDD.n343 GND 0.0234f
C4899 VDD.n351 GND 0.0903f
C4900 VDD.n352 GND 0.449f
C4901 VDD.t796 GND 0.0874f
C4902 VDD.t741 GND 0.0422f
C4903 VDD.t101 GND 0.0884f
C4904 VDD.t659 GND 0.0334f
C4905 VDD.n377 GND 0.0358f
C4906 VDD.n378 GND 0.0516f
C4907 VDD.n379 GND 0.555f
C4908 VDD.t731 GND 0.0144f
C4909 VDD.t1153 GND 0.0101f
C4910 VDD.t661 GND 0.0119f
C4911 VDD.t1169 GND 0.012f
C4912 VDD.t1132 GND 0.0186f
C4913 VDD.t48 GND 0.0268f
C4914 VDD.t728 GND 0.0155f
C4915 VDD.t456 GND 0.0163f
C4916 VDD.t1059 GND 0.0163f
C4917 VDD.t407 GND 0.0188f
C4918 VDD.t729 GND 0.0309f
C4919 VDD.n396 GND 0.0104f
C4920 VDD.n426 GND 0.0652f
C4921 VDD.n427 GND 0.556f
C4922 VDD.n431 GND 0.0253f
C4923 VDD.n434 GND 0.0109f
C4924 VDD.n437 GND 0.0109f
C4925 VDD.n444 GND 0.0247f
C4926 VDD.t1339 GND 0.0324f
C4927 VDD.t1365 GND 0.0138f
C4928 VDD.t1451 GND 0.0138f
C4929 VDD.t1343 GND 0.0138f
C4930 VDD.t1463 GND 0.0138f
C4931 VDD.n447 GND 0.0165f
C4932 VDD.n449 GND 0.103f
C4933 VDD.n453 GND 0.0227f
C4934 VDD.n454 GND 0.0137f
C4935 VDD.n460 GND 0.0257f
C4936 VDD.n464 GND 0.0257f
C4937 VDD.n466 GND 0.0257f
C4938 VDD.n467 GND 0.0193f
C4939 VDD.n468 GND 0.0152f
C4940 VDD.n470 GND 0.0257f
C4941 VDD.n474 GND 0.0257f
C4942 VDD.n476 GND 0.0257f
C4943 VDD.n480 GND 0.0257f
C4944 VDD.n482 GND 0.0257f
C4945 VDD.n486 GND 0.0257f
C4946 VDD.n488 GND 0.0257f
C4947 VDD.n492 GND 0.0219f
C4948 VDD.n493 GND 0.0137f
C4949 VDD.n498 GND 0.0128f
C4950 VDD.n499 GND 0.0109f
C4951 VDD.n500 GND 0.0112f
C4952 VDD.t1383 GND 0.0114f
C4953 VDD.t1453 GND 0.0138f
C4954 VDD.t1363 GND 0.0138f
C4955 VDD.t1431 GND 0.0138f
C4956 VDD.t1455 GND 0.0138f
C4957 VDD.t1351 GND 0.0138f
C4958 VDD.t1415 GND 0.0138f
C4959 VDD.t1445 GND 0.0138f
C4960 VDD.t1377 GND 0.0138f
C4961 VDD.t1421 GND 0.0133f
C4962 VDD.t1341 GND 0.0179f
C4963 VDD.t1409 GND 0.0138f
C4964 VDD.t1435 GND 0.0138f
C4965 VDD.t1461 GND 0.0138f
C4966 VDD.t1389 GND 0.0112f
C4967 VDD.t1439 GND 0.0138f
C4968 VDD.t1353 GND 0.0138f
C4969 VDD.t1417 GND 0.0138f
C4970 VDD.t1387 GND 0.0138f
C4971 VDD.t1457 GND 0.0179f
C4972 VDD.t1405 GND 0.0133f
C4973 VDD.t1381 GND 0.0138f
C4974 VDD.t1449 GND 0.0138f
C4975 VDD.t1401 GND 0.0138f
C4976 VDD.t1375 GND 0.0138f
C4977 VDD.t1443 GND 0.0138f
C4978 VDD.t1361 GND 0.0138f
C4979 VDD.t1427 GND 0.0138f
C4980 VDD.t1393 GND 0.0138f
C4981 VDD.t1357 GND 0.0138f
C4982 VDD.n501 GND 0.0112f
C4983 VDD.n502 GND 0.0109f
C4984 VDD.n503 GND 0.0103f
C4985 VDD.n505 GND 0.0124f
C4986 VDD.n506 GND 0.0137f
C4987 VDD.n510 GND 0.0177f
C4988 VDD.n514 GND 0.0257f
C4989 VDD.n516 GND 0.0257f
C4990 VDD.n520 GND 0.0257f
C4991 VDD.n522 GND 0.0257f
C4992 VDD.n526 GND 0.0257f
C4993 VDD.n528 GND 0.0257f
C4994 VDD.n532 GND 0.0257f
C4995 VDD.n534 GND 0.0257f
C4996 VDD.n535 GND 0.0152f
C4997 VDD.n538 GND 0.0193f
C4998 VDD.n540 GND 0.0257f
C4999 VDD.n544 GND 0.0257f
C5000 VDD.n546 GND 0.0257f
C5001 VDD.n550 GND 0.0208f
C5002 VDD.n551 GND 0.0137f
C5003 VDD.n555 GND 0.0257f
C5004 VDD.n559 GND 0.0257f
C5005 VDD.n561 GND 0.0257f
C5006 VDD.n565 GND 0.0257f
C5007 VDD.n567 GND 0.0257f
C5008 VDD.n571 GND 0.0239f
C5009 VDD.n572 GND 0.0137f
C5010 VDD.n577 GND 0.0128f
C5011 VDD.n578 GND 0.0109f
C5012 VDD.n579 GND 0.0112f
C5013 VDD.t1413 GND 0.0125f
C5014 VDD.t1441 GND 0.0138f
C5015 VDD.t1371 GND 0.0138f
C5016 VDD.t1397 GND 0.0138f
C5017 VDD.t1429 GND 0.0138f
C5018 VDD.t1373 GND 0.0138f
C5019 VDD.t1399 GND 0.0138f
C5020 VDD.t1345 GND 0.0138f
C5021 VDD.t1367 GND 0.0138f
C5022 VDD.t1385 GND 0.0133f
C5023 VDD.t1407 GND 0.0179f
C5024 VDD.t1433 GND 0.0138f
C5025 VDD.t1459 GND 0.0138f
C5026 VDD.n580 GND 0.0112f
C5027 VDD.t1437 GND 0.0137f
C5028 VDD.t1369 GND 0.0138f
C5029 VDD.t1391 GND 0.0138f
C5030 VDD.t1425 GND 0.0138f
C5031 VDD.t1359 GND 0.0138f
C5032 VDD.t1395 GND 0.0138f
C5033 VDD.t1337 GND 0.0138f
C5034 VDD.t1419 GND 0.0138f
C5035 VDD.t1447 GND 0.0138f
C5036 VDD.t1379 GND 0.0138f
C5037 VDD.t1403 GND 0.0138f
C5038 VDD.t1347 GND 0.0133f
C5039 VDD.t518 GND 0.0179f
C5040 VDD.t532 GND 0.0133f
C5041 VDD.n581 GND 0.0112f
C5042 VDD.t520 GND 0.0138f
C5043 VDD.t530 GND 0.0138f
C5044 VDD.t526 GND 0.0138f
C5045 VDD.t534 GND 0.0138f
C5046 VDD.t514 GND 0.0138f
C5047 VDD.t528 GND 0.0138f
C5048 VDD.t536 GND 0.0138f
C5049 VDD.t516 GND 0.0138f
C5050 VDD.t522 GND 0.0138f
C5051 VDD.t506 GND 0.0138f
C5052 VDD.t510 GND 0.0138f
C5053 VDD.t524 GND 0.0138f
C5054 VDD.t508 GND 0.0133f
C5055 VDD.t1073 GND 0.0178f
C5056 VDD.t1075 GND 0.0138f
C5057 VDD.t1077 GND 0.0138f
C5058 VDD.t1079 GND 0.0131f
C5059 VDD.t47 GND 0.0146f
C5060 VDD.t152 GND 0.0139f
C5061 VDD.t1304 GND 0.0232f
C5062 VDD.t663 GND 0.0174f
C5063 VDD.n582 GND 0.0182f
C5064 VDD.n586 GND 0.0384f
C5065 VDD.n588 GND 0.0299f
C5066 VDD.n589 GND 0.0193f
C5067 VDD.n592 GND 0.0152f
C5068 VDD.n594 GND 0.0174f
C5069 VDD.n595 GND 0.0137f
C5070 VDD.n599 GND 0.0109f
C5071 VDD.n601 GND 0.0144f
C5072 VDD.n603 GND 0.0257f
C5073 VDD.n606 GND 0.0257f
C5074 VDD.n608 GND 0.0257f
C5075 VDD.n609 GND 0.0193f
C5076 VDD.n610 GND 0.0152f
C5077 VDD.n612 GND 0.0257f
C5078 VDD.n616 GND 0.0257f
C5079 VDD.n618 GND 0.0257f
C5080 VDD.n622 GND 0.0257f
C5081 VDD.n624 GND 0.0257f
C5082 VDD.n628 GND 0.0257f
C5083 VDD.n630 GND 0.0257f
C5084 VDD.n634 GND 0.0257f
C5085 VDD.n638 GND 0.0257f
C5086 VDD.n640 GND 0.0257f
C5087 VDD.n644 GND 0.0236f
C5088 VDD.n645 GND 0.0137f
C5089 VDD.n648 GND 0.0128f
C5090 VDD.n653 GND 0.0137f
C5091 VDD.n655 GND 0.0211f
C5092 VDD.n656 GND 0.0193f
C5093 VDD.n657 GND 0.0152f
C5094 VDD.n659 GND 0.0257f
C5095 VDD.n663 GND 0.0257f
C5096 VDD.n665 GND 0.0257f
C5097 VDD.n669 GND 0.0257f
C5098 VDD.n671 GND 0.0257f
C5099 VDD.n675 GND 0.0257f
C5100 VDD.n677 GND 0.0257f
C5101 VDD.n681 GND 0.0257f
C5102 VDD.n685 GND 0.0257f
C5103 VDD.n687 GND 0.0236f
C5104 VDD.n688 GND 0.0137f
C5105 VDD.n693 GND 0.0128f
C5106 VDD.n696 GND 0.0137f
C5107 VDD.n700 GND 0.0211f
C5108 VDD.n702 GND 0.0257f
C5109 VDD.n703 GND 0.0193f
C5110 VDD.n704 GND 0.0152f
C5111 VDD.n706 GND 0.0133f
C5112 VDD.n707 GND 8.99f
C5113 VDD.t1060 GND 0.0102f
C5114 VDD.t0 GND 0.0128f
C5115 VDD.t745 GND 0.0352f
C5116 VDD.n723 GND 0.0116f
C5117 VDD.n724 GND 0.195f
C5118 VDD.t16 GND 0.0342f
C5119 VDD.t45 GND 0.0118f
C5120 VDD.t698 GND 0.0262f
C5121 VDD.t1250 GND 0.0489f
C5122 VDD.t459 GND 0.0208f
C5123 VDD.n725 GND 0.0157f
C5124 VDD.n755 GND 0.121f
C5125 VDD.t1209 GND 0.0874f
C5126 VDD.t176 GND 0.0422f
C5127 VDD.t155 GND 0.0884f
C5128 VDD.t139 GND 0.0334f
C5129 VDD.n780 GND 0.0358f
C5130 VDD.n781 GND 0.0516f
C5131 VDD.t700 GND 0.0144f
C5132 VDD.t1232 GND 0.0101f
C5133 VDD.t1206 GND 0.0119f
C5134 VDD.t1238 GND 0.012f
C5135 VDD.t1276 GND 0.0186f
C5136 VDD.t161 GND 0.0268f
C5137 VDD.t359 GND 0.0155f
C5138 VDD.t86 GND 0.0163f
C5139 VDD.t695 GND 0.0163f
C5140 VDD.t1465 GND 0.0188f
C5141 VDD.t1107 GND 0.0309f
C5142 VDD.n798 GND 0.0104f
C5143 VDD.n828 GND 0.0652f
C5144 VDD.n829 GND 0.354f
C5145 VDD.n830 GND 0.446f
C5146 VDD.n832 GND 0.013f
C5147 VDD.n835 GND 0.0109f
C5148 VDD.n838 GND 0.0109f
C5149 VDD.n845 GND 0.0253f
C5150 VDD.t813 GND 0.0318f
C5151 VDD.t839 GND 0.0138f
C5152 VDD.t925 GND 0.0138f
C5153 VDD.t817 GND 0.0138f
C5154 VDD.t809 GND 0.0138f
C5155 VDD.n848 GND 0.0163f
C5156 VDD.n850 GND 0.102f
C5157 VDD.n854 GND 0.0233f
C5158 VDD.n855 GND 0.0137f
C5159 VDD.n861 GND 0.0257f
C5160 VDD.n865 GND 0.0257f
C5161 VDD.n867 GND 0.0257f
C5162 VDD.n868 GND 0.0193f
C5163 VDD.n869 GND 0.0152f
C5164 VDD.n871 GND 0.0257f
C5165 VDD.n875 GND 0.0257f
C5166 VDD.n877 GND 0.0257f
C5167 VDD.n881 GND 0.0257f
C5168 VDD.n883 GND 0.0257f
C5169 VDD.n887 GND 0.0257f
C5170 VDD.n889 GND 0.0257f
C5171 VDD.n893 GND 0.0214f
C5172 VDD.n894 GND 0.0137f
C5173 VDD.n899 GND 0.0128f
C5174 VDD.n900 GND 0.0109f
C5175 VDD.n901 GND 0.0112f
C5176 VDD.t857 GND 0.011f
C5177 VDD.t799 GND 0.0138f
C5178 VDD.t835 GND 0.0138f
C5179 VDD.t905 GND 0.0138f
C5180 VDD.t801 GND 0.0138f
C5181 VDD.t825 GND 0.0138f
C5182 VDD.t889 GND 0.0138f
C5183 VDD.t919 GND 0.0138f
C5184 VDD.t851 GND 0.0138f
C5185 VDD.t895 GND 0.0133f
C5186 VDD.t815 GND 0.0179f
C5187 VDD.t883 GND 0.0138f
C5188 VDD.t909 GND 0.0138f
C5189 VDD.t807 GND 0.0138f
C5190 VDD.t863 GND 0.0115f
C5191 VDD.t913 GND 0.0138f
C5192 VDD.t827 GND 0.0138f
C5193 VDD.t891 GND 0.0138f
C5194 VDD.t861 GND 0.0138f
C5195 VDD.t803 GND 0.0179f
C5196 VDD.t879 GND 0.0133f
C5197 VDD.t855 GND 0.0138f
C5198 VDD.t923 GND 0.0138f
C5199 VDD.t875 GND 0.0138f
C5200 VDD.t849 GND 0.0138f
C5201 VDD.t917 GND 0.0138f
C5202 VDD.t837 GND 0.0138f
C5203 VDD.t901 GND 0.0138f
C5204 VDD.t867 GND 0.0138f
C5205 VDD.t829 GND 0.0138f
C5206 VDD.n902 GND 0.0112f
C5207 VDD.n903 GND 0.0109f
C5208 VDD.n906 GND 0.013f
C5209 VDD.n907 GND 0.0137f
C5210 VDD.n911 GND 0.0172f
C5211 VDD.n915 GND 0.0257f
C5212 VDD.n917 GND 0.0257f
C5213 VDD.n921 GND 0.0257f
C5214 VDD.n923 GND 0.0257f
C5215 VDD.n927 GND 0.0257f
C5216 VDD.n929 GND 0.0257f
C5217 VDD.n933 GND 0.0257f
C5218 VDD.n935 GND 0.0257f
C5219 VDD.n936 GND 0.0152f
C5220 VDD.n939 GND 0.0193f
C5221 VDD.n941 GND 0.0257f
C5222 VDD.n945 GND 0.0257f
C5223 VDD.n947 GND 0.0257f
C5224 VDD.n951 GND 0.0214f
C5225 VDD.n952 GND 0.0137f
C5226 VDD.n958 GND 0.0257f
C5227 VDD.n960 GND 0.0257f
C5228 VDD.n964 GND 0.0257f
C5229 VDD.n966 GND 0.0257f
C5230 VDD.n970 GND 0.0257f
C5231 VDD.n972 GND 0.0257f
C5232 VDD.n976 GND 0.0233f
C5233 VDD.n977 GND 0.0137f
C5234 VDD.n982 GND 0.0128f
C5235 VDD.n983 GND 0.0109f
C5236 VDD.n984 GND 0.0112f
C5237 VDD.t887 GND 0.0122f
C5238 VDD.t915 GND 0.0138f
C5239 VDD.t845 GND 0.0138f
C5240 VDD.t871 GND 0.0138f
C5241 VDD.t903 GND 0.0138f
C5242 VDD.t847 GND 0.0138f
C5243 VDD.t873 GND 0.0138f
C5244 VDD.t819 GND 0.0138f
C5245 VDD.t841 GND 0.0138f
C5246 VDD.t859 GND 0.0133f
C5247 VDD.t881 GND 0.0179f
C5248 VDD.t907 GND 0.0138f
C5249 VDD.t805 GND 0.0138f
C5250 VDD.n985 GND 0.0112f
C5251 VDD.t911 GND 0.0133f
C5252 VDD.t843 GND 0.0138f
C5253 VDD.t865 GND 0.0138f
C5254 VDD.t899 GND 0.0138f
C5255 VDD.t833 GND 0.0138f
C5256 VDD.t869 GND 0.0138f
C5257 VDD.t811 GND 0.0138f
C5258 VDD.t893 GND 0.0138f
C5259 VDD.t921 GND 0.0138f
C5260 VDD.t853 GND 0.0138f
C5261 VDD.t877 GND 0.0138f
C5262 VDD.t821 GND 0.0133f
C5263 VDD.t436 GND 0.0179f
C5264 VDD.t450 GND 0.0137f
C5265 VDD.n986 GND 0.0112f
C5266 VDD.t438 GND 0.0138f
C5267 VDD.t448 GND 0.0138f
C5268 VDD.t444 GND 0.0138f
C5269 VDD.t452 GND 0.0138f
C5270 VDD.t432 GND 0.0138f
C5271 VDD.t446 GND 0.0138f
C5272 VDD.t454 GND 0.0138f
C5273 VDD.t434 GND 0.0138f
C5274 VDD.t440 GND 0.0138f
C5275 VDD.t424 GND 0.0138f
C5276 VDD.t428 GND 0.0138f
C5277 VDD.t442 GND 0.0138f
C5278 VDD.t426 GND 0.0133f
C5279 VDD.t1291 GND 0.0178f
C5280 VDD.t1293 GND 0.0138f
C5281 VDD.t1295 GND 0.0138f
C5282 VDD.t1289 GND 0.0131f
C5283 VDD.t154 GND 0.0146f
C5284 VDD.t546 GND 0.0139f
C5285 VDD.t1134 GND 0.0232f
C5286 VDD.t735 GND 0.0171f
C5287 VDD.n987 GND 0.0182f
C5288 VDD.n991 GND 0.0384f
C5289 VDD.n993 GND 0.0299f
C5290 VDD.n994 GND 0.0193f
C5291 VDD.n997 GND 0.0152f
C5292 VDD.n999 GND 0.0169f
C5293 VDD.n1000 GND 0.0137f
C5294 VDD.n1004 GND 0.0109f
C5295 VDD.n1006 GND 0.0149f
C5296 VDD.n1008 GND 0.0257f
C5297 VDD.n1011 GND 0.0257f
C5298 VDD.n1013 GND 0.0257f
C5299 VDD.n1014 GND 0.0193f
C5300 VDD.n1015 GND 0.0152f
C5301 VDD.n1017 GND 0.0257f
C5302 VDD.n1021 GND 0.0257f
C5303 VDD.n1023 GND 0.0257f
C5304 VDD.n1027 GND 0.0257f
C5305 VDD.n1029 GND 0.0257f
C5306 VDD.n1033 GND 0.0257f
C5307 VDD.n1035 GND 0.0257f
C5308 VDD.n1039 GND 0.0257f
C5309 VDD.n1043 GND 0.0257f
C5310 VDD.n1045 GND 0.0257f
C5311 VDD.n1049 GND 0.023f
C5312 VDD.n1050 GND 0.0137f
C5313 VDD.n1053 GND 0.0128f
C5314 VDD.n1058 GND 0.0137f
C5315 VDD.n1060 GND 0.0216f
C5316 VDD.n1061 GND 0.0193f
C5317 VDD.n1062 GND 0.0152f
C5318 VDD.n1064 GND 0.0257f
C5319 VDD.n1068 GND 0.0257f
C5320 VDD.n1070 GND 0.0257f
C5321 VDD.n1074 GND 0.0257f
C5322 VDD.n1076 GND 0.0257f
C5323 VDD.n1080 GND 0.0257f
C5324 VDD.n1082 GND 0.0257f
C5325 VDD.n1086 GND 0.0257f
C5326 VDD.n1090 GND 0.0257f
C5327 VDD.n1092 GND 0.023f
C5328 VDD.n1093 GND 0.0137f
C5329 VDD.n1098 GND 0.0128f
C5330 VDD.n1101 GND 0.0137f
C5331 VDD.n1105 GND 0.0216f
C5332 VDD.n1107 GND 0.0257f
C5333 VDD.n1108 GND 0.0193f
C5334 VDD.n1109 GND 0.0151f
C5335 VDD.n1110 GND 8.98f
C5336 VDD.n1111 GND 2.82f
C5337 VDD.n1112 GND 0.393f
C5338 VDD.n1113 GND 0.451f
C5339 VDD.n1114 GND 2.13f
C5340 VDD.n1115 GND 0.763f
C5341 VDD.n1124 GND 0.0105f
C5342 VDD.n1125 GND 0.0424f
C5343 VDD.n1137 GND 0.0245f
C5344 VDD.n1170 GND 0.0181f
C5345 VDD.t1243 GND 0.0195f
C5346 VDD.t89 GND 0.0188f
C5347 VDD.t1147 GND 0.0228f
C5348 VDD.t99 GND 0.0197f
C5349 VDD.t682 GND 0.0171f
C5350 VDD.t191 GND 0.0142f
C5351 VDD.t653 GND 0.0225f
C5352 VDD.t1069 GND 0.0197f
C5353 VDD.t141 GND 0.0171f
C5354 VDD.t795 GND 0.0171f
C5355 VDD.t178 GND 0.0162f
C5356 VDD.t791 GND 0.0175f
C5357 VDD.t2 GND 0.0173f
C5358 VDD.t702 GND 0.0175f
C5359 VDD.t1256 GND 0.0175f
C5360 VDD.t1241 GND 0.022f
C5361 VDD.n1174 GND 0.0533f
C5362 VDD.n1178 GND 0.0148f
C5363 VDD.n1179 GND 0.052f
C5364 VDD.n1180 GND 3.66f
C5365 VDD.n1181 GND 3.55f
C5366 VDD.n1190 GND 0.0105f
C5367 VDD.n1191 GND 0.0424f
C5368 VDD.n1203 GND 0.0245f
C5369 VDD.n1236 GND 0.0181f
C5370 VDD.t1174 GND 0.0195f
C5371 VDD.t649 GND 0.0188f
C5372 VDD.t672 GND 0.0228f
C5373 VDD.t137 GND 0.0197f
C5374 VDD.t578 GND 0.0171f
C5375 VDD.t1071 GND 0.0142f
C5376 VDD.t56 GND 0.0225f
C5377 VDD.t501 GND 0.0197f
C5378 VDD.t777 GND 0.0171f
C5379 VDD.t127 GND 0.0171f
C5380 VDD.t1137 GND 0.0162f
C5381 VDD.t1211 GND 0.0175f
C5382 VDD.t1322 GND 0.0173f
C5383 VDD.t68 GND 0.0175f
C5384 VDD.t1314 GND 0.0175f
C5385 VDD.t1166 GND 0.022f
C5386 VDD.n1240 GND 0.0533f
C5387 VDD.n1244 GND 0.0148f
C5388 VDD.n1245 GND 0.453f
C5389 VDD.n1246 GND 0.313f
C5390 VDD.n1249 GND 0.0147f
C5391 VDD.n1251 GND 0.1f
C5392 VDD.n1255 GND 0.0213f
C5393 VDD.n1270 GND 0.0227f
C5394 VDD.n1274 GND 0.0373f
C5395 VDD.n1276 GND 0.0373f
C5396 VDD.n1280 GND 0.0373f
C5397 VDD.n1282 GND 0.0373f
C5398 VDD.n1283 GND 0.111f
C5399 VDD.n1285 GND 0.0127f
C5400 VDD.t317 GND 0.018f
C5401 VDD.t241 GND 0.018f
C5402 VDD.t293 GND 0.018f
C5403 VDD.t219 GND 0.018f
C5404 VDD.t245 GND 0.018f
C5405 VDD.t277 GND 0.018f
C5406 VDD.t213 GND 0.018f
C5407 VDD.t303 GND 0.0157f
C5408 VDD.n1291 GND 0.0332f
C5409 VDD.n1295 GND 0.0373f
C5410 VDD.n1297 GND 0.0373f
C5411 VDD.n1301 GND 0.0373f
C5412 VDD.n1303 GND 0.0268f
C5413 VDD.n1304 GND 0.0689f
C5414 VDD.n1310 GND 0.0127f
C5415 VDD.n1314 GND 0.0117f
C5416 VDD.t255 GND 0.018f
C5417 VDD.t287 GND 0.018f
C5418 VDD.t331 GND 0.018f
C5419 VDD.t259 GND 0.0172f
C5420 VDD.t631 GND 0.018f
C5421 VDD.t621 GND 0.018f
C5422 VDD.t643 GND 0.018f
C5423 VDD.n1331 GND 0.0127f
C5424 VDD.n1333 GND 0.0127f
C5425 VDD.n1337 GND 0.0127f
C5426 VDD.n1339 GND 0.0127f
C5427 VDD.t617 GND 0.018f
C5428 VDD.t627 GND 0.018f
C5429 VDD.t635 GND 0.0165f
C5430 VDD.n1351 GND 0.0127f
C5431 VDD.n1354 GND 0.0127f
C5432 VDD.n1356 GND 0.0127f
C5433 VDD.t393 GND 0.0223f
C5434 VDD.n1371 GND 0.0227f
C5435 VDD.t401 GND 0.017f
C5436 VDD.t397 GND 0.018f
C5437 VDD.t395 GND 0.018f
C5438 VDD.t399 GND 0.0233f
C5439 VDD.n1372 GND 0.0135f
C5440 VDD.n1383 GND 0.0127f
C5441 VDD.n1387 GND 0.0127f
C5442 VDD.n1389 GND 0.0127f
C5443 VDD.n1393 GND 0.01f
C5444 VDD.t641 GND 0.018f
C5445 VDD.t623 GND 0.018f
C5446 VDD.t633 GND 0.018f
C5447 VDD.t613 GND 0.0152f
C5448 VDD.t639 GND 0.018f
C5449 VDD.t625 GND 0.018f
C5450 VDD.t629 GND 0.018f
C5451 VDD.t619 GND 0.0118f
C5452 VDD.n1397 GND 0.0135f
C5453 VDD.n1410 GND 0.0117f
C5454 VDD.n1412 GND 0.0127f
C5455 VDD.n1416 GND 0.0127f
C5456 VDD.n1418 GND 0.0127f
C5457 VDD.n1422 GND 0.0104f
C5458 VDD.n1428 GND 0.0189f
C5459 VDD.t325 GND 0.0174f
C5460 VDD.t247 GND 0.018f
C5461 VDD.t221 GND 0.018f
C5462 VDD.t275 GND 0.018f
C5463 VDD.t243 GND 0.018f
C5464 VDD.t217 GND 0.018f
C5465 VDD.n1429 GND 0.0135f
C5466 VDD.n1433 GND 0.0121f
C5467 VDD.n1437 GND 0.0127f
C5468 VDD.n1441 GND 0.0127f
C5469 VDD.n1443 GND 0.0127f
C5470 VDD.n1447 GND 0.0127f
C5471 VDD.n1449 GND 0.0127f
C5472 VDD.n1453 GND 0.0131f
C5473 VDD.t327 GND 0.018f
C5474 VDD.t231 GND 0.018f
C5475 VDD.t309 GND 0.018f
C5476 VDD.t279 GND 0.0139f
C5477 VDD.n1456 GND 0.0135f
C5478 VDD.t227 GND 0.0184f
C5479 VDD.t301 GND 0.0174f
C5480 VDD.t249 GND 0.018f
C5481 VDD.t223 GND 0.0276f
C5482 VDD.t297 GND 0.0395f
C5483 VDD.t265 GND 0.04f
C5484 VDD.t205 GND 0.04f
C5485 VDD.t239 GND 0.04f
C5486 VDD.t207 GND 0.04f
C5487 VDD.t271 GND 0.04f
C5488 VDD.t235 GND 0.04f
C5489 VDD.t313 GND 0.04f
C5490 VDD.t285 GND 0.04f
C5491 VDD.t253 GND 0.04f
C5492 VDD.t323 GND 0.0402f
C5493 VDD.t281 GND 0.0181f
C5494 VDD.t209 GND 0.0234f
C5495 VDD.n1457 GND 0.0129f
C5496 VDD.n1467 GND 0.0127f
C5497 VDD.n1469 GND 0.0127f
C5498 VDD.n1473 GND 0.0127f
C5499 VDD.n1475 GND 0.0127f
C5500 VDD.n1479 GND 0.0127f
C5501 VDD.n1481 GND 0.0127f
C5502 VDD.n1485 GND 0.0127f
C5503 VDD.n1489 GND 0.0127f
C5504 VDD.n1491 GND 0.0127f
C5505 VDD.n1495 GND 0.0127f
C5506 VDD.n1497 GND 0.0127f
C5507 VDD.n1501 GND 0.0127f
C5508 VDD.n1503 GND 0.0116f
C5509 VDD.t321 GND 0.0414f
C5510 VDD.t211 GND 0.018f
C5511 VDD.t283 GND 0.018f
C5512 VDD.t311 GND 0.018f
C5513 VDD.t233 GND 0.018f
C5514 VDD.t269 GND 0.018f
C5515 VDD.t315 GND 0.018f
C5516 VDD.t237 GND 0.018f
C5517 VDD.t273 GND 0.018f
C5518 VDD.t261 GND 0.018f
C5519 VDD.t295 GND 0.018f
C5520 VDD.t319 GND 0.018f
C5521 VDD.t267 GND 0.018f
C5522 VDD.t299 GND 0.018f
C5523 VDD.t225 GND 0.018f
C5524 VDD.t251 GND 0.0174f
C5525 VDD.t289 GND 0.018f
C5526 VDD.t257 GND 0.018f
C5527 VDD.t329 GND 0.018f
C5528 VDD.t305 GND 0.018f
C5529 VDD.t215 GND 0.018f
C5530 VDD.t263 GND 0.018f
C5531 VDD.t229 GND 0.018f
C5532 VDD.t307 GND 0.0217f
C5533 VDD.n1507 GND 0.0189f
C5534 VDD.n1513 GND 0.0101f
C5535 VDD.n1517 GND 0.0127f
C5536 VDD.n1519 GND 0.0127f
C5537 VDD.n1523 GND 0.0127f
C5538 VDD.n1526 GND 0.0904f
C5539 VDD.n1527 GND 0.0258f
C5540 VDD.n1529 GND 0.0276f
C5541 VDD.n1533 GND 0.0276f
C5542 VDD.n1537 GND 0.0276f
C5543 VDD.n1539 GND 0.0201f
C5544 VDD.n1540 GND 0.308f
C5545 VDD.t651 GND 0.0247f
C5546 VDD.n1541 GND 0.0356f
C5547 VDD.n1548 GND 0.0874f
C5548 VDD.t1093 GND 0.0102f
C5549 VDD.t1222 GND 0.0128f
C5550 VDD.t389 GND 0.0352f
C5551 VDD.n1564 GND 0.0116f
C5552 VDD.n1565 GND 0.195f
C5553 VDD.t410 GND 0.0342f
C5554 VDD.t52 GND 0.0118f
C5555 VDD.t72 GND 0.0262f
C5556 VDD.t345 GND 0.0489f
C5557 VDD.t1163 GND 0.0208f
C5558 VDD.n1566 GND 0.0157f
C5559 VDD.n1596 GND 0.121f
C5560 VDD.n1597 GND 0.454f
C5561 VDD.n1598 GND 0.439f
C5562 VDD.n1599 GND 0.337f
C5563 VDD.n1600 GND 2.47f
C5564 VDD.n1601 GND 1.96f
C5565 VDD.n1602 GND 3.55f
C5566 VDD.n1603 GND 10.2f
C5567 VDD.n1613 GND 0.0185f
C5568 VDD.n1622 GND 0.0562f
C5569 VDD.n1623 GND 0.0449f
C5570 VDD.n1642 GND 0.0348f
C5571 VDD.n1646 GND 0.03f
C5572 VDD.n1652 GND 0.0265f
C5573 VDD.n1653 GND 0.118f
C5574 VDD.n1654 GND 0.0985f
C5575 VDD.n1655 GND 0.0705f
C5576 VDD.n1656 GND 0.0906f
C5577 VDD.n1657 GND 0.112f
C5578 VDD.n1658 GND 0.111f
C5579 VDD.n1659 GND 0.101f
C5580 VDD.n1660 GND 0.115f
C5581 VDD.n1661 GND 0.0861f
C5582 VDD.n1662 GND 0.226f
C5583 VDD.n1663 GND 8.71f
C5584 VDD.n1664 GND 0.208f
C5585 VDD.n1665 GND 0.0179f
C5586 VDD.n1666 GND 0.035f
C5587 VDD.t1227 GND 0.0452f
C5588 VDD.n1678 GND 0.0265f
C5589 VDD.n1686 GND 0.0331f
C5590 VDD.n1687 GND 0.0115f
C5591 VDD.n1695 GND 0.0381f
C5592 VDD.n1711 GND 0.0556f
C5593 VDD.t37 GND 0.0452f
C5594 VDD.n1712 GND 0.0265f
C5595 VDD.n1721 GND 0.0371f
C5596 VDD.n1723 GND 0.0102f
C5597 VDD.n1737 GND 0.0366f
C5598 VDD.n1738 GND 0.044f
C5599 VDD.n1744 GND 0.0442f
C5600 VDD.n1748 GND 0.0101f
C5601 VDD.n1749 GND 0.0356f
C5602 VDD.n1753 GND 0.0219f
C5603 VDD.n1754 GND 0.0102f
C5604 VDD.t753 GND 0.128f
C5605 VDD.n1764 GND 0.0556f
C5606 VDD.n1770 GND 0.0102f
C5607 VDD.n1771 GND 0.0217f
C5608 VDD.n1773 GND 0.0188f
C5609 VDD.n1774 GND 0.0982f
C5610 VDD.n1775 GND 0.323f
C5611 VDD.n1801 GND 0.0336f
C5612 VDD.t39 GND 0.0141f
C5613 VDD.n1802 GND 0.0147f
C5614 VDD.n1803 GND 0.0181f
C5615 VDD.t1224 GND 0.014f
C5616 VDD.n1804 GND 0.121f
C5617 VDD.n1805 GND 0.731f
C5618 VDD.n1806 GND 0.0776f
C5619 VDD.n1807 GND 0.867f
C5620 VDD.n1808 GND 0.697f
C5621 VDD.t1095 GND 0.029f
C5622 VDD.t54 GND 0.0101f
C5623 VDD.n1809 GND 0.0529f
C5624 VDD.n1816 GND 0.0439f
C5625 VDD.n1817 GND 0.0168f
C5626 VDD.n1821 GND 0.0516f
C5627 VDD.n1823 GND 0.059f
C5628 VDD.t382 GND 0.0218f
C5629 VDD.n1836 GND 0.03f
C5630 VDD.n1839 GND 0.0152f
C5631 VDD.n1840 GND 0.0101f
C5632 VDD.n1841 GND 0.0865f
C5633 VDD.n1842 GND 0.0289f
C5634 VDD.n1847 GND 0.0515f
C5635 VDD.n1849 GND 0.068f
C5636 VDD.n1857 GND 0.0655f
C5637 VDD.n1858 GND 0.0292f
C5638 VDD.n1863 GND 0.0317f
C5639 VDD.t355 GND 0.0515f
C5640 VDD.n1872 GND 0.223f
C5641 VDD.n1873 GND 0.125f
C5642 VDD.n1874 GND 0.0503f
C5643 VDD.n1875 GND 0.0163f
C5644 VDD.t417 GND 0.0647f
C5645 VDD.n1886 GND 0.0344f
C5646 VDD.n1887 GND 0.0851f
C5647 VDD.n1892 GND 0.0649f
C5648 VDD.n1893 GND 0.068f
C5649 VDD.n1901 GND 0.0323f
C5650 VDD.n1905 GND 0.0292f
C5651 VDD.t420 GND 0.0515f
C5652 VDD.n1914 GND 0.0515f
C5653 VDD.n1916 GND 0.0662f
C5654 VDD.n1917 GND 0.212f
C5655 VDD.n1918 GND 0.126f
C5656 VDD.n1919 GND 0.148f
C5657 VDD.n1920 GND 0.0593f
C5658 VDD.n1921 GND 1.58f
C5659 VDD.n1922 GND 0.12f
C5660 VDD.n1923 GND 0.105f
C5661 VDD.t1056 GND 0.0162f
C5662 VDD.t1288 GND 0.0162f
C5663 VDD.n1924 GND 0.247f
C5664 VDD.n1925 GND 0.0132f
C5665 VDD.n1927 GND 0.303f
C5666 VDD.n1930 GND 0.0229f
C5667 VDD.n1931 GND 0.24f
C5668 VDD.n1933 GND 0.0959f
C5669 VDD.n1935 GND 0.0102f
C5670 VDD.n1939 GND 0.151f
C5671 VDD.n1940 GND 0.0102f
C5672 VDD.n1942 GND 0.0229f
C5673 VDD.n1943 GND 0.0137f
C5674 VDD.t1286 GND 0.0162f
C5675 VDD.n1945 GND 0.124f
C5676 VDD.n1946 GND 0.0645f
C5677 VDD.n1948 GND 0.0102f
C5678 VDD.n1949 GND 0.24f
C5679 VDD.n1950 GND 0.0128f
C5680 VDD.n1951 GND 0.0128f
C5681 VDD.t1285 GND 0.302f
C5682 VDD.n1952 GND 0.0106f
C5683 VDD.n1953 GND 0.151f
C5684 VDD.n1957 GND 0.0669f
C5685 VDD.n1960 GND 0.0128f
C5686 VDD.n1961 GND 0.0128f
C5687 VDD.t1055 GND 0.293f
C5688 VDD.n1967 GND 0.0128f
C5689 VDD.n1968 GND 0.0128f
C5690 VDD.t1287 GND 0.303f
C5691 VDD.n1970 GND 0.0128f
C5692 VDD.n1971 GND 0.0128f
C5693 VDD.n1974 GND 0.0102f
C5694 VDD.n1979 GND 0.153f
C5695 VDD.n1980 GND 0.0958f
C5696 VDD.n1981 GND 0.0249f
C5697 VDD.n1982 GND 7.24f
C5698 VDD.n1983 GND 0.208f
C5699 VDD.n2009 GND 0.0336f
C5700 VDD.t362 GND 0.0141f
C5701 VDD.n2010 GND 0.0147f
C5702 VDD.n2011 GND 0.0181f
C5703 VDD.t31 GND 0.014f
C5704 VDD.n2012 GND 0.463f
C5705 VDD.n2013 GND 0.349f
C5706 VDD.n2014 GND 0.0179f
C5707 VDD.n2015 GND 0.035f
C5708 VDD.t29 GND 0.0452f
C5709 VDD.n2027 GND 0.0265f
C5710 VDD.n2035 GND 0.0331f
C5711 VDD.n2036 GND 0.0115f
C5712 VDD.n2044 GND 0.0381f
C5713 VDD.n2060 GND 0.0556f
C5714 VDD.t365 GND 0.0452f
C5715 VDD.n2061 GND 0.0265f
C5716 VDD.n2070 GND 0.0371f
C5717 VDD.n2072 GND 0.0102f
C5718 VDD.n2086 GND 0.0366f
C5719 VDD.n2087 GND 0.044f
C5720 VDD.n2093 GND 0.0442f
C5721 VDD.n2097 GND 0.0101f
C5722 VDD.n2098 GND 0.0356f
C5723 VDD.n2102 GND 0.0219f
C5724 VDD.n2103 GND 0.0102f
C5725 VDD.t129 GND 0.128f
C5726 VDD.n2113 GND 0.0556f
C5727 VDD.n2119 GND 0.0102f
C5728 VDD.n2120 GND 0.0217f
C5729 VDD.n2122 GND 0.0188f
C5730 VDD.n2123 GND 0.0982f
C5731 VDD.n2124 GND 0.323f
C5732 VDD.n2125 GND 0.0366f
C5733 VDD.n2126 GND 0.0776f
C5734 VDD.n2127 GND 0.442f
C5735 VDD.n2128 GND 0.836f
C5736 VDD.n2129 GND 0.33f
C5737 VDD.t683 GND 0.029f
C5738 VDD.t647 GND 0.0101f
C5739 VDD.n2130 GND 0.0529f
C5740 VDD.n2137 GND 0.0439f
C5741 VDD.n2138 GND 0.0168f
C5742 VDD.n2142 GND 0.0516f
C5743 VDD.n2144 GND 0.059f
C5744 VDD.t1139 GND 0.0218f
C5745 VDD.n2157 GND 0.03f
C5746 VDD.n2160 GND 0.0152f
C5747 VDD.n2161 GND 0.0101f
C5748 VDD.n2162 GND 0.0865f
C5749 VDD.n2163 GND 0.0289f
C5750 VDD.n2168 GND 0.0515f
C5751 VDD.n2170 GND 0.068f
C5752 VDD.n2178 GND 0.0655f
C5753 VDD.n2179 GND 0.0292f
C5754 VDD.n2184 GND 0.0317f
C5755 VDD.t574 GND 0.0515f
C5756 VDD.n2193 GND 0.223f
C5757 VDD.n2194 GND 0.125f
C5758 VDD.n2195 GND 0.0503f
C5759 VDD.n2196 GND 0.0163f
C5760 VDD.t1085 GND 0.0647f
C5761 VDD.n2207 GND 0.0344f
C5762 VDD.n2208 GND 0.0851f
C5763 VDD.n2213 GND 0.0649f
C5764 VDD.n2214 GND 0.068f
C5765 VDD.n2222 GND 0.0323f
C5766 VDD.n2226 GND 0.0292f
C5767 VDD.t148 GND 0.0515f
C5768 VDD.n2235 GND 0.0515f
C5769 VDD.n2237 GND 0.0662f
C5770 VDD.n2238 GND 0.212f
C5771 VDD.n2239 GND 0.126f
C5772 VDD.n2240 GND 0.148f
C5773 VDD.n2241 GND 0.0593f
C5774 VDD.n2242 GND 1.58f
C5775 VDD.n2243 GND 0.208f
C5776 VDD.n2244 GND 0.0179f
C5777 VDD.n2245 GND 0.035f
C5778 VDD.t541 GND 0.0452f
C5779 VDD.n2257 GND 0.0265f
C5780 VDD.n2265 GND 0.0331f
C5781 VDD.n2266 GND 0.0115f
C5782 VDD.n2274 GND 0.0381f
C5783 VDD.n2290 GND 0.0556f
C5784 VDD.t466 GND 0.0452f
C5785 VDD.n2291 GND 0.0265f
C5786 VDD.n2300 GND 0.0371f
C5787 VDD.n2302 GND 0.0102f
C5788 VDD.n2316 GND 0.0366f
C5789 VDD.n2317 GND 0.044f
C5790 VDD.n2323 GND 0.0442f
C5791 VDD.n2327 GND 0.0101f
C5792 VDD.n2328 GND 0.0356f
C5793 VDD.n2332 GND 0.0219f
C5794 VDD.n2333 GND 0.0102f
C5795 VDD.t70 GND 0.128f
C5796 VDD.n2343 GND 0.0556f
C5797 VDD.n2349 GND 0.0102f
C5798 VDD.n2350 GND 0.0217f
C5799 VDD.n2352 GND 0.0188f
C5800 VDD.n2353 GND 0.0982f
C5801 VDD.n2354 GND 0.323f
C5802 VDD.n2380 GND 0.0336f
C5803 VDD.t464 GND 0.0141f
C5804 VDD.n2381 GND 0.0147f
C5805 VDD.n2382 GND 0.0181f
C5806 VDD.t538 GND 0.014f
C5807 VDD.n2383 GND 0.121f
C5808 VDD.n2384 GND 0.731f
C5809 VDD.n2385 GND 0.0776f
C5810 VDD.n2386 GND 0.867f
C5811 VDD.n2387 GND 0.697f
C5812 VDD.t74 GND 0.029f
C5813 VDD.t105 GND 0.0101f
C5814 VDD.n2388 GND 0.0529f
C5815 VDD.n2395 GND 0.0439f
C5816 VDD.n2396 GND 0.0168f
C5817 VDD.n2400 GND 0.0516f
C5818 VDD.n2402 GND 0.059f
C5819 VDD.t1297 GND 0.0218f
C5820 VDD.n2415 GND 0.03f
C5821 VDD.n2418 GND 0.0152f
C5822 VDD.n2419 GND 0.0101f
C5823 VDD.n2420 GND 0.0865f
C5824 VDD.n2421 GND 0.0289f
C5825 VDD.n2426 GND 0.0515f
C5826 VDD.n2428 GND 0.068f
C5827 VDD.n2436 GND 0.0655f
C5828 VDD.n2437 GND 0.0292f
C5829 VDD.n2442 GND 0.0317f
C5830 VDD.t103 GND 0.0515f
C5831 VDD.n2451 GND 0.223f
C5832 VDD.n2452 GND 0.125f
C5833 VDD.n2453 GND 0.0503f
C5834 VDD.n2454 GND 0.0163f
C5835 VDD.t567 GND 0.0647f
C5836 VDD.n2465 GND 0.0344f
C5837 VDD.n2466 GND 0.0851f
C5838 VDD.n2471 GND 0.0649f
C5839 VDD.n2472 GND 0.068f
C5840 VDD.n2480 GND 0.0323f
C5841 VDD.n2484 GND 0.0292f
C5842 VDD.t676 GND 0.0515f
C5843 VDD.n2493 GND 0.0515f
C5844 VDD.n2495 GND 0.0662f
C5845 VDD.n2496 GND 0.212f
C5846 VDD.n2497 GND 0.126f
C5847 VDD.n2498 GND 0.148f
C5848 VDD.n2499 GND 0.0593f
C5849 VDD.n2500 GND 1.58f
C5850 VDD.n2501 GND 0.208f
C5851 VDD.n2502 GND 0.0179f
C5852 VDD.n2503 GND 0.035f
C5853 VDD.t472 GND 0.0452f
C5854 VDD.n2515 GND 0.0265f
C5855 VDD.n2523 GND 0.0331f
C5856 VDD.n2524 GND 0.0115f
C5857 VDD.n2532 GND 0.0381f
C5858 VDD.n2548 GND 0.0556f
C5859 VDD.t117 GND 0.0452f
C5860 VDD.n2549 GND 0.0265f
C5861 VDD.n2558 GND 0.0371f
C5862 VDD.n2560 GND 0.0102f
C5863 VDD.n2574 GND 0.0366f
C5864 VDD.n2575 GND 0.044f
C5865 VDD.n2581 GND 0.0442f
C5866 VDD.n2585 GND 0.0101f
C5867 VDD.n2586 GND 0.0356f
C5868 VDD.n2590 GND 0.0219f
C5869 VDD.n2591 GND 0.0102f
C5870 VDD.t680 GND 0.128f
C5871 VDD.n2601 GND 0.0556f
C5872 VDD.n2607 GND 0.0102f
C5873 VDD.n2608 GND 0.0217f
C5874 VDD.n2610 GND 0.0188f
C5875 VDD.n2611 GND 0.0982f
C5876 VDD.n2612 GND 0.323f
C5877 VDD.n2638 GND 0.0336f
C5878 VDD.t119 GND 0.0141f
C5879 VDD.n2639 GND 0.0147f
C5880 VDD.n2640 GND 0.0181f
C5881 VDD.t474 GND 0.014f
C5882 VDD.n2641 GND 0.121f
C5883 VDD.n2642 GND 0.731f
C5884 VDD.n2643 GND 0.0776f
C5885 VDD.n2644 GND 0.867f
C5886 VDD.n2645 GND 0.697f
C5887 VDD.t499 GND 0.029f
C5888 VDD.t1118 GND 0.0101f
C5889 VDD.n2646 GND 0.0529f
C5890 VDD.n2653 GND 0.0439f
C5891 VDD.n2654 GND 0.0168f
C5892 VDD.n2658 GND 0.0516f
C5893 VDD.n2660 GND 0.059f
C5894 VDD.t95 GND 0.0218f
C5895 VDD.n2673 GND 0.03f
C5896 VDD.n2676 GND 0.0152f
C5897 VDD.n2677 GND 0.0101f
C5898 VDD.n2678 GND 0.0865f
C5899 VDD.n2679 GND 0.0289f
C5900 VDD.n2684 GND 0.0515f
C5901 VDD.n2686 GND 0.068f
C5902 VDD.n2694 GND 0.0655f
C5903 VDD.n2695 GND 0.0292f
C5904 VDD.n2700 GND 0.0317f
C5905 VDD.t421 GND 0.0515f
C5906 VDD.n2709 GND 0.223f
C5907 VDD.n2710 GND 0.125f
C5908 VDD.n2711 GND 0.0503f
C5909 VDD.n2712 GND 0.0163f
C5910 VDD.t387 GND 0.0647f
C5911 VDD.n2723 GND 0.0344f
C5912 VDD.n2724 GND 0.0851f
C5913 VDD.n2729 GND 0.0649f
C5914 VDD.n2730 GND 0.068f
C5915 VDD.n2738 GND 0.0323f
C5916 VDD.n2742 GND 0.0292f
C5917 VDD.t689 GND 0.0515f
C5918 VDD.n2751 GND 0.0515f
C5919 VDD.n2753 GND 0.0662f
C5920 VDD.n2754 GND 0.212f
C5921 VDD.n2755 GND 0.126f
C5922 VDD.n2756 GND 0.148f
C5923 VDD.n2757 GND 0.0593f
C5924 VDD.n2758 GND 1.58f
C5925 VDD.n2759 GND 0.208f
C5926 VDD.n2760 GND 0.0179f
C5927 VDD.n2761 GND 0.035f
C5928 VDD.t1309 GND 0.0452f
C5929 VDD.n2773 GND 0.0265f
C5930 VDD.n2781 GND 0.0331f
C5931 VDD.n2782 GND 0.0115f
C5932 VDD.n2790 GND 0.0381f
C5933 VDD.n2806 GND 0.0556f
C5934 VDD.t21 GND 0.0452f
C5935 VDD.n2807 GND 0.0265f
C5936 VDD.n2816 GND 0.0371f
C5937 VDD.n2818 GND 0.0102f
C5938 VDD.n2832 GND 0.0366f
C5939 VDD.n2833 GND 0.044f
C5940 VDD.n2839 GND 0.0442f
C5941 VDD.n2843 GND 0.0101f
C5942 VDD.n2844 GND 0.0356f
C5943 VDD.n2848 GND 0.0219f
C5944 VDD.n2849 GND 0.0102f
C5945 VDD.t733 GND 0.128f
C5946 VDD.n2859 GND 0.0556f
C5947 VDD.n2865 GND 0.0102f
C5948 VDD.n2866 GND 0.0217f
C5949 VDD.n2868 GND 0.0188f
C5950 VDD.n2869 GND 0.0982f
C5951 VDD.n2870 GND 0.323f
C5952 VDD.n2896 GND 0.0336f
C5953 VDD.t19 GND 0.0141f
C5954 VDD.n2897 GND 0.0147f
C5955 VDD.n2898 GND 0.0181f
C5956 VDD.t1306 GND 0.014f
C5957 VDD.n2899 GND 0.121f
C5958 VDD.n2900 GND 0.731f
C5959 VDD.n2901 GND 0.0776f
C5960 VDD.n2902 GND 0.867f
C5961 VDD.n2903 GND 0.697f
C5962 VDD.t714 GND 0.029f
C5963 VDD.t403 GND 0.0101f
C5964 VDD.n2904 GND 0.0529f
C5965 VDD.n2911 GND 0.0439f
C5966 VDD.n2912 GND 0.0168f
C5967 VDD.n2916 GND 0.0516f
C5968 VDD.n2918 GND 0.059f
C5969 VDD.t462 GND 0.0218f
C5970 VDD.n2931 GND 0.03f
C5971 VDD.n2934 GND 0.0152f
C5972 VDD.n2935 GND 0.0101f
C5973 VDD.n2936 GND 0.0865f
C5974 VDD.n2937 GND 0.0289f
C5975 VDD.n2942 GND 0.0515f
C5976 VDD.n2944 GND 0.068f
C5977 VDD.n2952 GND 0.0655f
C5978 VDD.n2953 GND 0.0292f
C5979 VDD.n2958 GND 0.0317f
C5980 VDD.t405 GND 0.0515f
C5981 VDD.n2967 GND 0.223f
C5982 VDD.n2968 GND 0.125f
C5983 VDD.n2969 GND 0.0503f
C5984 VDD.n2970 GND 0.0163f
C5985 VDD.t560 GND 0.0647f
C5986 VDD.n2981 GND 0.0344f
C5987 VDD.n2982 GND 0.0851f
C5988 VDD.n2987 GND 0.0649f
C5989 VDD.n2988 GND 0.068f
C5990 VDD.n2996 GND 0.0323f
C5991 VDD.n3000 GND 0.0292f
C5992 VDD.t93 GND 0.0515f
C5993 VDD.n3009 GND 0.0515f
C5994 VDD.n3011 GND 0.0662f
C5995 VDD.n3012 GND 0.212f
C5996 VDD.n3013 GND 0.126f
C5997 VDD.n3014 GND 0.148f
C5998 VDD.n3015 GND 0.0593f
C5999 VDD.n3016 GND 1.58f
C6000 VDD.n3017 GND 0.208f
C6001 VDD.n3018 GND 0.0179f
C6002 VDD.n3019 GND 0.035f
C6003 VDD.t6 GND 0.0452f
C6004 VDD.n3031 GND 0.0265f
C6005 VDD.n3039 GND 0.0331f
C6006 VDD.n3040 GND 0.0115f
C6007 VDD.n3048 GND 0.0381f
C6008 VDD.n3064 GND 0.0556f
C6009 VDD.t590 GND 0.0452f
C6010 VDD.n3065 GND 0.0265f
C6011 VDD.n3074 GND 0.0371f
C6012 VDD.n3076 GND 0.0102f
C6013 VDD.n3090 GND 0.0366f
C6014 VDD.n3091 GND 0.044f
C6015 VDD.n3097 GND 0.0442f
C6016 VDD.n3101 GND 0.0101f
C6017 VDD.n3102 GND 0.0356f
C6018 VDD.n3106 GND 0.0219f
C6019 VDD.n3107 GND 0.0102f
C6020 VDD.t125 GND 0.128f
C6021 VDD.n3117 GND 0.0556f
C6022 VDD.n3123 GND 0.0102f
C6023 VDD.n3124 GND 0.0217f
C6024 VDD.n3126 GND 0.0188f
C6025 VDD.n3127 GND 0.0982f
C6026 VDD.n3128 GND 0.323f
C6027 VDD.n3154 GND 0.0336f
C6028 VDD.t588 GND 0.0141f
C6029 VDD.n3155 GND 0.0147f
C6030 VDD.n3156 GND 0.0181f
C6031 VDD.t8 GND 0.014f
C6032 VDD.n3157 GND 0.121f
C6033 VDD.n3158 GND 0.731f
C6034 VDD.n3159 GND 0.0776f
C6035 VDD.n3160 GND 0.867f
C6036 VDD.n3161 GND 0.697f
C6037 VDD.t685 GND 0.029f
C6038 VDD.t774 GND 0.0101f
C6039 VDD.n3162 GND 0.0529f
C6040 VDD.n3169 GND 0.0439f
C6041 VDD.n3170 GND 0.0168f
C6042 VDD.n3174 GND 0.0516f
C6043 VDD.n3176 GND 0.059f
C6044 VDD.t1105 GND 0.0218f
C6045 VDD.n3189 GND 0.03f
C6046 VDD.n3192 GND 0.0152f
C6047 VDD.n3193 GND 0.0101f
C6048 VDD.n3194 GND 0.0865f
C6049 VDD.n3195 GND 0.0289f
C6050 VDD.n3200 GND 0.0515f
C6051 VDD.n3202 GND 0.068f
C6052 VDD.n3210 GND 0.0655f
C6053 VDD.n3211 GND 0.0292f
C6054 VDD.n3216 GND 0.0317f
C6055 VDD.t144 GND 0.0515f
C6056 VDD.n3225 GND 0.223f
C6057 VDD.n3226 GND 0.125f
C6058 VDD.n3227 GND 0.0503f
C6059 VDD.n3228 GND 0.0163f
C6060 VDD.t573 GND 0.0647f
C6061 VDD.n3239 GND 0.0344f
C6062 VDD.n3240 GND 0.0851f
C6063 VDD.n3245 GND 0.0649f
C6064 VDD.n3246 GND 0.068f
C6065 VDD.n3254 GND 0.0323f
C6066 VDD.n3258 GND 0.0292f
C6067 VDD.t76 GND 0.0515f
C6068 VDD.n3267 GND 0.0515f
C6069 VDD.n3269 GND 0.0662f
C6070 VDD.n3270 GND 0.212f
C6071 VDD.n3271 GND 0.126f
C6072 VDD.n3272 GND 0.148f
C6073 VDD.n3273 GND 0.0593f
C6074 VDD.n3274 GND 1.58f
C6075 VDD.n3275 GND 0.208f
C6076 VDD.n3276 GND 0.0179f
C6077 VDD.n3277 GND 0.035f
C6078 VDD.t1194 GND 0.0452f
C6079 VDD.n3289 GND 0.0265f
C6080 VDD.n3297 GND 0.0331f
C6081 VDD.n3298 GND 0.0115f
C6082 VDD.n3306 GND 0.0381f
C6083 VDD.n3322 GND 0.0556f
C6084 VDD.t550 GND 0.0452f
C6085 VDD.n3323 GND 0.0265f
C6086 VDD.n3332 GND 0.0371f
C6087 VDD.n3334 GND 0.0102f
C6088 VDD.n3348 GND 0.0366f
C6089 VDD.n3349 GND 0.044f
C6090 VDD.n3355 GND 0.0442f
C6091 VDD.n3359 GND 0.0101f
C6092 VDD.n3360 GND 0.0356f
C6093 VDD.n3364 GND 0.0219f
C6094 VDD.n3365 GND 0.0102f
C6095 VDD.t504 GND 0.128f
C6096 VDD.n3375 GND 0.0556f
C6097 VDD.n3381 GND 0.0102f
C6098 VDD.n3382 GND 0.0217f
C6099 VDD.n3384 GND 0.0188f
C6100 VDD.n3385 GND 0.0982f
C6101 VDD.n3386 GND 0.323f
C6102 VDD.n3412 GND 0.0336f
C6103 VDD.t548 GND 0.0141f
C6104 VDD.n3413 GND 0.0147f
C6105 VDD.n3414 GND 0.0181f
C6106 VDD.t1196 GND 0.014f
C6107 VDD.n3415 GND 0.121f
C6108 VDD.n3416 GND 0.731f
C6109 VDD.n3417 GND 0.0776f
C6110 VDD.n3418 GND 0.867f
C6111 VDD.n3419 GND 0.697f
C6112 VDD.t360 GND 0.029f
C6113 VDD.t181 GND 0.0101f
C6114 VDD.n3420 GND 0.0529f
C6115 VDD.n3427 GND 0.0439f
C6116 VDD.n3428 GND 0.0168f
C6117 VDD.n3432 GND 0.0516f
C6118 VDD.n3434 GND 0.059f
C6119 VDD.t1259 GND 0.0218f
C6120 VDD.n3447 GND 0.03f
C6121 VDD.n3450 GND 0.0152f
C6122 VDD.n3451 GND 0.0101f
C6123 VDD.n3452 GND 0.0865f
C6124 VDD.n3453 GND 0.0289f
C6125 VDD.n3458 GND 0.0515f
C6126 VDD.n3460 GND 0.068f
C6127 VDD.n3468 GND 0.0655f
C6128 VDD.n3469 GND 0.0292f
C6129 VDD.n3474 GND 0.0317f
C6130 VDD.t179 GND 0.0515f
C6131 VDD.n3483 GND 0.223f
C6132 VDD.n3484 GND 0.125f
C6133 VDD.n3485 GND 0.0503f
C6134 VDD.n3486 GND 0.0163f
C6135 VDD.t143 GND 0.0647f
C6136 VDD.n3497 GND 0.0344f
C6137 VDD.n3498 GND 0.0851f
C6138 VDD.n3503 GND 0.0649f
C6139 VDD.n3504 GND 0.068f
C6140 VDD.n3512 GND 0.0323f
C6141 VDD.n3516 GND 0.0292f
C6142 VDD.t1186 GND 0.0515f
C6143 VDD.n3525 GND 0.0515f
C6144 VDD.n3527 GND 0.0662f
C6145 VDD.n3528 GND 0.212f
C6146 VDD.n3529 GND 0.126f
C6147 VDD.n3530 GND 0.148f
C6148 VDD.n3531 GND 0.0593f
C6149 VDD.n3532 GND 1.58f
C6150 VDD.n3533 GND 0.208f
C6151 VDD.n3534 GND 0.0179f
C6152 VDD.n3535 GND 0.035f
C6153 VDD.t1268 GND 0.0452f
C6154 VDD.n3547 GND 0.0265f
C6155 VDD.n3555 GND 0.0331f
C6156 VDD.n3556 GND 0.0115f
C6157 VDD.n3564 GND 0.0381f
C6158 VDD.n3580 GND 0.0556f
C6159 VDD.t1100 GND 0.0452f
C6160 VDD.n3581 GND 0.0265f
C6161 VDD.n3590 GND 0.0371f
C6162 VDD.n3592 GND 0.0102f
C6163 VDD.n3606 GND 0.0366f
C6164 VDD.n3607 GND 0.044f
C6165 VDD.n3613 GND 0.0442f
C6166 VDD.n3617 GND 0.0101f
C6167 VDD.n3618 GND 0.0356f
C6168 VDD.n3622 GND 0.0219f
C6169 VDD.n3623 GND 0.0102f
C6170 VDD.t1141 GND 0.128f
C6171 VDD.n3633 GND 0.0556f
C6172 VDD.n3639 GND 0.0102f
C6173 VDD.n3640 GND 0.0217f
C6174 VDD.n3642 GND 0.0188f
C6175 VDD.n3643 GND 0.0982f
C6176 VDD.n3644 GND 0.323f
C6177 VDD.n3670 GND 0.0336f
C6178 VDD.t1097 GND 0.0141f
C6179 VDD.n3671 GND 0.0147f
C6180 VDD.n3672 GND 0.0181f
C6181 VDD.t1270 GND 0.014f
C6182 VDD.n3673 GND 0.121f
C6183 VDD.n3674 GND 0.731f
C6184 VDD.n3675 GND 0.0776f
C6185 VDD.n3676 GND 0.867f
C6186 VDD.n3677 GND 0.697f
C6187 VDD.t1182 GND 0.029f
C6188 VDD.t343 GND 0.0101f
C6189 VDD.n3678 GND 0.0529f
C6190 VDD.n3685 GND 0.0439f
C6191 VDD.n3686 GND 0.0168f
C6192 VDD.n3690 GND 0.0516f
C6193 VDD.n3692 GND 0.059f
C6194 VDD.t1187 GND 0.0218f
C6195 VDD.n3705 GND 0.03f
C6196 VDD.n3708 GND 0.0152f
C6197 VDD.n3709 GND 0.0101f
C6198 VDD.n3710 GND 0.0865f
C6199 VDD.n3711 GND 0.0289f
C6200 VDD.n3716 GND 0.0515f
C6201 VDD.n3718 GND 0.068f
C6202 VDD.n3726 GND 0.0655f
C6203 VDD.n3727 GND 0.0292f
C6204 VDD.n3732 GND 0.0317f
C6205 VDD.t145 GND 0.0515f
C6206 VDD.n3741 GND 0.223f
C6207 VDD.n3742 GND 0.125f
C6208 VDD.n3743 GND 0.0503f
C6209 VDD.n3744 GND 0.0163f
C6210 VDD.t142 GND 0.0647f
C6211 VDD.n3755 GND 0.0344f
C6212 VDD.n3756 GND 0.0851f
C6213 VDD.n3761 GND 0.0649f
C6214 VDD.n3762 GND 0.068f
C6215 VDD.n3770 GND 0.0323f
C6216 VDD.n3774 GND 0.0292f
C6217 VDD.t556 GND 0.0515f
C6218 VDD.n3783 GND 0.0515f
C6219 VDD.n3785 GND 0.0662f
C6220 VDD.n3786 GND 0.212f
C6221 VDD.n3787 GND 0.126f
C6222 VDD.n3788 GND 0.148f
C6223 VDD.n3789 GND 0.0593f
C6224 VDD.n3790 GND 1.58f
C6225 VDD.n3791 GND 0.208f
C6226 VDD.n3792 GND 0.0179f
C6227 VDD.n3793 GND 0.035f
C6228 VDD.t81 GND 0.0452f
C6229 VDD.n3805 GND 0.0265f
C6230 VDD.n3813 GND 0.0331f
C6231 VDD.n3814 GND 0.0115f
C6232 VDD.n3822 GND 0.0381f
C6233 VDD.n3838 GND 0.0556f
C6234 VDD.t785 GND 0.0452f
C6235 VDD.n3839 GND 0.0265f
C6236 VDD.n3848 GND 0.0371f
C6237 VDD.n3850 GND 0.0102f
C6238 VDD.n3864 GND 0.0366f
C6239 VDD.n3865 GND 0.044f
C6240 VDD.n3871 GND 0.0442f
C6241 VDD.n3875 GND 0.0101f
C6242 VDD.n3876 GND 0.0356f
C6243 VDD.n3880 GND 0.0219f
C6244 VDD.n3881 GND 0.0102f
C6245 VDD.t1061 GND 0.128f
C6246 VDD.n3891 GND 0.0556f
C6247 VDD.n3897 GND 0.0102f
C6248 VDD.n3898 GND 0.0217f
C6249 VDD.n3900 GND 0.0188f
C6250 VDD.n3901 GND 0.0982f
C6251 VDD.n3902 GND 0.323f
C6252 VDD.n3928 GND 0.0336f
C6253 VDD.t783 GND 0.0141f
C6254 VDD.n3929 GND 0.0147f
C6255 VDD.n3930 GND 0.0181f
C6256 VDD.t78 GND 0.014f
C6257 VDD.n3931 GND 0.121f
C6258 VDD.n3932 GND 0.731f
C6259 VDD.n3933 GND 0.0776f
C6260 VDD.n3934 GND 0.867f
C6261 VDD.n3935 GND 0.697f
C6262 VDD.t655 GND 0.029f
C6263 VDD.t565 GND 0.0101f
C6264 VDD.n3936 GND 0.0529f
C6265 VDD.n3943 GND 0.0439f
C6266 VDD.n3944 GND 0.0168f
C6267 VDD.n3948 GND 0.0516f
C6268 VDD.n3950 GND 0.059f
C6269 VDD.t58 GND 0.0218f
C6270 VDD.n3963 GND 0.03f
C6271 VDD.n3966 GND 0.0152f
C6272 VDD.n3967 GND 0.0101f
C6273 VDD.n3968 GND 0.0865f
C6274 VDD.n3969 GND 0.0289f
C6275 VDD.n3974 GND 0.0515f
C6276 VDD.n3976 GND 0.068f
C6277 VDD.n3984 GND 0.0655f
C6278 VDD.n3985 GND 0.0292f
C6279 VDD.n3990 GND 0.0317f
C6280 VDD.t563 GND 0.0515f
C6281 VDD.n3999 GND 0.223f
C6282 VDD.n4000 GND 0.125f
C6283 VDD.n4001 GND 0.0503f
C6284 VDD.n4002 GND 0.0163f
C6285 VDD.t782 GND 0.0647f
C6286 VDD.n4013 GND 0.0344f
C6287 VDD.n4014 GND 0.0851f
C6288 VDD.n4019 GND 0.0649f
C6289 VDD.n4020 GND 0.068f
C6290 VDD.n4028 GND 0.0323f
C6291 VDD.n4032 GND 0.0292f
C6292 VDD.t562 GND 0.0515f
C6293 VDD.n4041 GND 0.0515f
C6294 VDD.n4043 GND 0.0662f
C6295 VDD.n4044 GND 0.212f
C6296 VDD.n4045 GND 0.126f
C6297 VDD.n4046 GND 0.148f
C6298 VDD.n4047 GND 0.0593f
C6299 VDD.n4048 GND 1.58f
C6300 VDD.n4049 GND 0.208f
C6301 VDD.n4050 GND 0.0179f
C6302 VDD.n4051 GND 0.035f
C6303 VDD.t723 GND 0.0452f
C6304 VDD.n4063 GND 0.0265f
C6305 VDD.n4071 GND 0.0331f
C6306 VDD.n4072 GND 0.0115f
C6307 VDD.n4080 GND 0.0381f
C6308 VDD.n4096 GND 0.0556f
C6309 VDD.t490 GND 0.0452f
C6310 VDD.n4097 GND 0.0265f
C6311 VDD.n4106 GND 0.0371f
C6312 VDD.n4108 GND 0.0102f
C6313 VDD.n4122 GND 0.0366f
C6314 VDD.n4123 GND 0.044f
C6315 VDD.n4129 GND 0.0442f
C6316 VDD.n4133 GND 0.0101f
C6317 VDD.n4134 GND 0.0356f
C6318 VDD.n4138 GND 0.0219f
C6319 VDD.n4139 GND 0.0102f
C6320 VDD.t414 GND 0.128f
C6321 VDD.n4149 GND 0.0556f
C6322 VDD.n4155 GND 0.0102f
C6323 VDD.n4156 GND 0.0217f
C6324 VDD.n4158 GND 0.0188f
C6325 VDD.n4159 GND 0.0982f
C6326 VDD.n4160 GND 0.323f
C6327 VDD.n4186 GND 0.0336f
C6328 VDD.t492 GND 0.0141f
C6329 VDD.n4187 GND 0.0147f
C6330 VDD.n4188 GND 0.0181f
C6331 VDD.t720 GND 0.014f
C6332 VDD.n4189 GND 0.121f
C6333 VDD.n4190 GND 0.731f
C6334 VDD.n4191 GND 0.0776f
C6335 VDD.n4192 GND 0.867f
C6336 VDD.n4193 GND 0.697f
C6337 VDD.t488 GND 0.029f
C6338 VDD.t1217 GND 0.0101f
C6339 VDD.n4194 GND 0.0529f
C6340 VDD.n4201 GND 0.0439f
C6341 VDD.n4202 GND 0.0168f
C6342 VDD.n4206 GND 0.0516f
C6343 VDD.n4208 GND 0.059f
C6344 VDD.t718 GND 0.0218f
C6345 VDD.n4221 GND 0.03f
C6346 VDD.n4224 GND 0.0152f
C6347 VDD.n4225 GND 0.0101f
C6348 VDD.n4226 GND 0.0865f
C6349 VDD.n4227 GND 0.0289f
C6350 VDD.n4232 GND 0.0515f
C6351 VDD.n4234 GND 0.068f
C6352 VDD.n4242 GND 0.0655f
C6353 VDD.n4243 GND 0.0292f
C6354 VDD.n4248 GND 0.0317f
C6355 VDD.t668 GND 0.0515f
C6356 VDD.n4257 GND 0.223f
C6357 VDD.n4258 GND 0.125f
C6358 VDD.n4259 GND 0.0503f
C6359 VDD.n4260 GND 0.0163f
C6360 VDD.t1087 GND 0.0647f
C6361 VDD.n4271 GND 0.0344f
C6362 VDD.n4272 GND 0.0851f
C6363 VDD.n4277 GND 0.0649f
C6364 VDD.n4278 GND 0.068f
C6365 VDD.n4286 GND 0.0323f
C6366 VDD.n4290 GND 0.0292f
C6367 VDD.t687 GND 0.0515f
C6368 VDD.n4299 GND 0.0515f
C6369 VDD.n4301 GND 0.0662f
C6370 VDD.n4302 GND 0.212f
C6371 VDD.n4303 GND 0.126f
C6372 VDD.n4304 GND 0.148f
C6373 VDD.n4305 GND 0.0593f
C6374 VDD.n4306 GND 1.58f
C6375 VDD.n4307 GND 0.208f
C6376 VDD.n4308 GND 0.0179f
C6377 VDD.n4309 GND 0.035f
C6378 VDD.t1112 GND 0.0452f
C6379 VDD.n4321 GND 0.0265f
C6380 VDD.n4329 GND 0.0331f
C6381 VDD.n4330 GND 0.0115f
C6382 VDD.n4338 GND 0.0381f
C6383 VDD.n4354 GND 0.0556f
C6384 VDD.t374 GND 0.0452f
C6385 VDD.n4355 GND 0.0265f
C6386 VDD.n4364 GND 0.0371f
C6387 VDD.n4366 GND 0.0102f
C6388 VDD.n4380 GND 0.0366f
C6389 VDD.n4381 GND 0.044f
C6390 VDD.n4387 GND 0.0442f
C6391 VDD.n4391 GND 0.0101f
C6392 VDD.n4392 GND 0.0356f
C6393 VDD.n4396 GND 0.0219f
C6394 VDD.n4397 GND 0.0102f
C6395 VDD.t165 GND 0.128f
C6396 VDD.n4407 GND 0.0556f
C6397 VDD.n4413 GND 0.0102f
C6398 VDD.n4414 GND 0.0217f
C6399 VDD.n4416 GND 0.0188f
C6400 VDD.n4417 GND 0.0982f
C6401 VDD.n4418 GND 0.323f
C6402 VDD.n4444 GND 0.0336f
C6403 VDD.t372 GND 0.0141f
C6404 VDD.n4445 GND 0.0147f
C6405 VDD.n4446 GND 0.0181f
C6406 VDD.t1109 GND 0.014f
C6407 VDD.n4447 GND 0.121f
C6408 VDD.n4448 GND 0.731f
C6409 VDD.n4449 GND 0.0776f
C6410 VDD.n4450 GND 0.867f
C6411 VDD.n4451 GND 0.697f
C6412 VDD.t87 GND 0.029f
C6413 VDD.t579 GND 0.0101f
C6414 VDD.n4452 GND 0.0529f
C6415 VDD.n4459 GND 0.0439f
C6416 VDD.n4460 GND 0.0168f
C6417 VDD.n4464 GND 0.0516f
C6418 VDD.n4466 GND 0.059f
C6419 VDD.t1202 GND 0.0218f
C6420 VDD.n4479 GND 0.03f
C6421 VDD.n4482 GND 0.0152f
C6422 VDD.n4483 GND 0.0101f
C6423 VDD.n4484 GND 0.0865f
C6424 VDD.n4485 GND 0.0289f
C6425 VDD.n4490 GND 0.0515f
C6426 VDD.n4492 GND 0.068f
C6427 VDD.n4500 GND 0.0655f
C6428 VDD.n4501 GND 0.0292f
C6429 VDD.n4506 GND 0.0317f
C6430 VDD.t561 GND 0.0515f
C6431 VDD.n4515 GND 0.223f
C6432 VDD.n4516 GND 0.125f
C6433 VDD.n4517 GND 0.0503f
C6434 VDD.n4518 GND 0.0163f
C6435 VDD.t558 GND 0.0647f
C6436 VDD.n4529 GND 0.0344f
C6437 VDD.n4530 GND 0.0851f
C6438 VDD.n4535 GND 0.0649f
C6439 VDD.n4536 GND 0.068f
C6440 VDD.n4544 GND 0.0323f
C6441 VDD.n4548 GND 0.0292f
C6442 VDD.t570 GND 0.0515f
C6443 VDD.n4557 GND 0.0515f
C6444 VDD.n4559 GND 0.0662f
C6445 VDD.n4560 GND 0.212f
C6446 VDD.n4561 GND 0.126f
C6447 VDD.n4562 GND 0.148f
C6448 VDD.n4563 GND 0.0593f
C6449 VDD.n4564 GND 1.58f
C6450 VDD.n4565 GND 0.208f
C6451 VDD.n4566 GND 0.0179f
C6452 VDD.n4567 GND 0.035f
C6453 VDD.t183 GND 0.0452f
C6454 VDD.n4579 GND 0.0265f
C6455 VDD.n4587 GND 0.0331f
C6456 VDD.n4588 GND 0.0115f
C6457 VDD.n4596 GND 0.0381f
C6458 VDD.n4612 GND 0.0556f
C6459 VDD.t111 GND 0.0452f
C6460 VDD.n4613 GND 0.0265f
C6461 VDD.n4622 GND 0.0371f
C6462 VDD.n4624 GND 0.0102f
C6463 VDD.n4638 GND 0.0366f
C6464 VDD.n4639 GND 0.044f
C6465 VDD.n4645 GND 0.0442f
C6466 VDD.n4649 GND 0.0101f
C6467 VDD.n4650 GND 0.0356f
C6468 VDD.n4654 GND 0.0219f
C6469 VDD.n4655 GND 0.0102f
C6470 VDD.t793 GND 0.128f
C6471 VDD.n4665 GND 0.0556f
C6472 VDD.n4671 GND 0.0102f
C6473 VDD.n4672 GND 0.0217f
C6474 VDD.n4674 GND 0.0188f
C6475 VDD.n4675 GND 0.0982f
C6476 VDD.n4676 GND 0.323f
C6477 VDD.n4702 GND 0.0336f
C6478 VDD.t109 GND 0.0141f
C6479 VDD.n4703 GND 0.0147f
C6480 VDD.n4704 GND 0.0181f
C6481 VDD.t185 GND 0.014f
C6482 VDD.n4705 GND 0.121f
C6483 VDD.n4706 GND 0.731f
C6484 VDD.n4707 GND 0.0776f
C6485 VDD.n4708 GND 0.867f
C6486 VDD.n4709 GND 0.697f
C6487 VDD.t1189 GND 0.029f
C6488 VDD.t14 GND 0.0101f
C6489 VDD.n4710 GND 0.0529f
C6490 VDD.n4717 GND 0.0439f
C6491 VDD.n4718 GND 0.0168f
C6492 VDD.n4722 GND 0.0516f
C6493 VDD.n4724 GND 0.059f
C6494 VDD.t602 GND 0.0218f
C6495 VDD.n4737 GND 0.03f
C6496 VDD.n4740 GND 0.0152f
C6497 VDD.n4741 GND 0.0101f
C6498 VDD.n4742 GND 0.0865f
C6499 VDD.n4743 GND 0.0289f
C6500 VDD.n4748 GND 0.0515f
C6501 VDD.n4750 GND 0.068f
C6502 VDD.n4758 GND 0.0655f
C6503 VDD.n4759 GND 0.0292f
C6504 VDD.n4764 GND 0.0317f
C6505 VDD.t750 GND 0.0515f
C6506 VDD.n4773 GND 0.223f
C6507 VDD.n4774 GND 0.125f
C6508 VDD.n4775 GND 0.0503f
C6509 VDD.n4776 GND 0.0163f
C6510 VDD.t572 GND 0.0647f
C6511 VDD.n4787 GND 0.0344f
C6512 VDD.n4788 GND 0.0851f
C6513 VDD.n4793 GND 0.0649f
C6514 VDD.n4794 GND 0.068f
C6515 VDD.n4802 GND 0.0323f
C6516 VDD.n4806 GND 0.0292f
C6517 VDD.t670 GND 0.0515f
C6518 VDD.n4815 GND 0.0515f
C6519 VDD.n4817 GND 0.0662f
C6520 VDD.n4818 GND 0.212f
C6521 VDD.n4819 GND 0.126f
C6522 VDD.n4820 GND 0.148f
C6523 VDD.n4821 GND 0.0593f
C6524 VDD.n4822 GND 1.58f
C6525 VDD.n4823 GND 0.21f
C6526 VDD.n4824 GND 0.0179f
C6527 VDD.n4825 GND 0.035f
C6528 VDD.t1121 GND 0.0452f
C6529 VDD.n4837 GND 0.0265f
C6530 VDD.n4845 GND 0.0331f
C6531 VDD.n4846 GND 0.0115f
C6532 VDD.n4854 GND 0.0381f
C6533 VDD.n4870 GND 0.0556f
C6534 VDD.t349 GND 0.0452f
C6535 VDD.n4871 GND 0.0265f
C6536 VDD.n4880 GND 0.0371f
C6537 VDD.n4882 GND 0.0102f
C6538 VDD.n4896 GND 0.0366f
C6539 VDD.n4897 GND 0.044f
C6540 VDD.n4903 GND 0.0442f
C6541 VDD.n4907 GND 0.0101f
C6542 VDD.n4908 GND 0.0356f
C6543 VDD.n4912 GND 0.0219f
C6544 VDD.n4913 GND 0.0102f
C6545 VDD.t1065 GND 0.128f
C6546 VDD.n4923 GND 0.0556f
C6547 VDD.n4929 GND 0.0102f
C6548 VDD.n4930 GND 0.0217f
C6549 VDD.n4932 GND 0.0188f
C6550 VDD.n4933 GND 0.641f
C6551 VDD.n4935 GND 0.275f
C6552 VDD.n4961 GND 0.0336f
C6553 VDD.t347 GND 0.0141f
C6554 VDD.n4962 GND 0.0147f
C6555 VDD.n4963 GND 0.0181f
C6556 VDD.t1123 GND 0.014f
C6557 VDD.n4964 GND 0.117f
C6558 VDD.n4965 GND 0.597f
C6559 VDD.n4966 GND 0.0801f
C6560 VDD.n4967 GND 0.131f
C6561 VDD.n4968 GND 0.0487f
C6562 VDD.n4969 GND 0.0141f
C6563 VDD.n4970 GND 0.557f
C6564 VDD.t1266 GND 0.029f
C6565 VDD.t769 GND 0.0101f
C6566 VDD.n4971 GND 0.0529f
C6567 VDD.n4978 GND 0.0439f
C6568 VDD.n4979 GND 0.0168f
C6569 VDD.n4983 GND 0.0516f
C6570 VDD.n4985 GND 0.059f
C6571 VDD.t1261 GND 0.0218f
C6572 VDD.n4998 GND 0.03f
C6573 VDD.n5001 GND 0.0152f
C6574 VDD.n5002 GND 0.0101f
C6575 VDD.n5003 GND 0.0865f
C6576 VDD.n5004 GND 0.0289f
C6577 VDD.n5009 GND 0.0515f
C6578 VDD.n5011 GND 0.068f
C6579 VDD.n5019 GND 0.0655f
C6580 VDD.n5020 GND 0.0292f
C6581 VDD.n5025 GND 0.0317f
C6582 VDD.t386 GND 0.0515f
C6583 VDD.n5034 GND 0.223f
C6584 VDD.n5035 GND 0.125f
C6585 VDD.n5036 GND 0.0503f
C6586 VDD.n5037 GND 0.0163f
C6587 VDD.t690 GND 0.0647f
C6588 VDD.n5048 GND 0.0344f
C6589 VDD.n5049 GND 0.0851f
C6590 VDD.n5054 GND 0.0649f
C6591 VDD.n5055 GND 0.068f
C6592 VDD.n5063 GND 0.0323f
C6593 VDD.n5067 GND 0.0292f
C6594 VDD.t581 GND 0.0515f
C6595 VDD.n5076 GND 0.0515f
C6596 VDD.n5078 GND 0.0662f
C6597 VDD.n5079 GND 0.212f
C6598 VDD.n5080 GND 0.126f
C6599 VDD.n5081 GND 0.208f
C6600 VDD.n5082 GND 0.305f
C6601 VDD.n5083 GND 1.62f
C6602 VDD.n5084 GND 0.226f
C6603 VDD.n5085 GND 0.254f
C6604 VDD.n5111 GND 0.0336f
C6605 VDD.t480 GND 0.0141f
C6606 VDD.n5112 GND 0.0147f
C6607 VDD.n5113 GND 0.0181f
C6608 VDD.t192 GND 0.014f
C6609 VDD.n5114 GND 0.117f
C6610 VDD.n5115 GND 0.6f
C6611 VDD.n5116 GND 0.0179f
C6612 VDD.n5117 GND 0.035f
C6613 VDD.t195 GND 0.0452f
C6614 VDD.n5129 GND 0.0265f
C6615 VDD.n5137 GND 0.0331f
C6616 VDD.n5138 GND 0.0115f
C6617 VDD.n5146 GND 0.0381f
C6618 VDD.n5162 GND 0.0556f
C6619 VDD.t482 GND 0.0452f
C6620 VDD.n5163 GND 0.0265f
C6621 VDD.n5172 GND 0.0371f
C6622 VDD.n5174 GND 0.0102f
C6623 VDD.n5188 GND 0.0366f
C6624 VDD.n5189 GND 0.044f
C6625 VDD.n5195 GND 0.0442f
C6626 VDD.n5199 GND 0.0101f
C6627 VDD.n5200 GND 0.0356f
C6628 VDD.n5204 GND 0.0219f
C6629 VDD.n5205 GND 0.0102f
C6630 VDD.t107 GND 0.128f
C6631 VDD.n5215 GND 0.0556f
C6632 VDD.n5221 GND 0.0102f
C6633 VDD.n5222 GND 0.0217f
C6634 VDD.n5224 GND 0.0188f
C6635 VDD.n5225 GND 0.399f
C6636 VDD.n5226 GND 0.453f
C6637 VDD.n5227 GND 0.142f
C6638 VDD.n5228 GND 0.0801f
C6639 VDD.n5229 GND 0.0277f
C6640 VDD.n5230 GND 0.0203f
C6641 VDD.n5231 GND 0.0141f
C6642 VDD.n5232 GND 0.544f
C6643 VDD.t1500 GND 0.029f
C6644 VDD.t131 GND 0.0101f
C6645 VDD.n5233 GND 0.0529f
C6646 VDD.n5240 GND 0.0439f
C6647 VDD.n5241 GND 0.0168f
C6648 VDD.n5245 GND 0.0516f
C6649 VDD.n5247 GND 0.059f
C6650 VDD.t771 GND 0.0218f
C6651 VDD.n5260 GND 0.03f
C6652 VDD.n5263 GND 0.0152f
C6653 VDD.n5264 GND 0.0101f
C6654 VDD.n5265 GND 0.0865f
C6655 VDD.n5266 GND 0.0289f
C6656 VDD.n5271 GND 0.0515f
C6657 VDD.n5273 GND 0.068f
C6658 VDD.n5281 GND 0.0655f
C6659 VDD.n5282 GND 0.0292f
C6660 VDD.n5287 GND 0.0317f
C6661 VDD.t559 GND 0.0515f
C6662 VDD.n5296 GND 0.223f
C6663 VDD.n5297 GND 0.125f
C6664 VDD.n5298 GND 0.0503f
C6665 VDD.n5299 GND 0.0163f
C6666 VDD.t418 GND 0.0647f
C6667 VDD.n5310 GND 0.0344f
C6668 VDD.n5311 GND 0.0851f
C6669 VDD.n5316 GND 0.0649f
C6670 VDD.n5317 GND 0.068f
C6671 VDD.n5325 GND 0.0323f
C6672 VDD.n5329 GND 0.0292f
C6673 VDD.t97 GND 0.0515f
C6674 VDD.n5338 GND 0.0515f
C6675 VDD.n5340 GND 0.0662f
C6676 VDD.n5341 GND 0.212f
C6677 VDD.n5342 GND 0.126f
C6678 VDD.n5343 GND 0.208f
C6679 VDD.n5344 GND 0.373f
C6680 VDD.n5345 GND 6.4f
C6681 VDD.n5346 GND 27.5f
C6682 VDD.n5347 GND 18.2f
C6683 VDD.n5348 GND 18.2f
C6684 VDD.n5349 GND 18.2f
C6685 VDD.n5350 GND 18.2f
C6686 VDD.n5351 GND 18.9f
C6687 VDD.n5352 GND 0.0179f
C6688 VDD.n5353 GND 0.035f
C6689 VDD.t1331 GND 0.0452f
C6690 VDD.n5365 GND 0.0265f
C6691 VDD.n5373 GND 0.0331f
C6692 VDD.n5374 GND 0.0115f
C6693 VDD.n5382 GND 0.0381f
C6694 VDD.n5398 GND 0.0556f
C6695 VDD.t757 GND 0.0452f
C6696 VDD.n5399 GND 0.0265f
C6697 VDD.n5408 GND 0.0371f
C6698 VDD.n5410 GND 0.0102f
C6699 VDD.n5424 GND 0.0366f
C6700 VDD.n5425 GND 0.044f
C6701 VDD.n5431 GND 0.0442f
C6702 VDD.n5435 GND 0.0101f
C6703 VDD.n5436 GND 0.0356f
C6704 VDD.n5440 GND 0.0219f
C6705 VDD.n5441 GND 0.0102f
C6706 VDD.t665 GND 0.128f
C6707 VDD.n5451 GND 0.0556f
C6708 VDD.n5457 GND 0.0102f
C6709 VDD.n5458 GND 0.0217f
C6710 VDD.n5460 GND 0.0188f
C6711 VDD.n5461 GND 0.701f
C6712 VDD.n5462 GND 0.582f
C6713 VDD.n5488 GND 0.0336f
C6714 VDD.t759 GND 0.0141f
C6715 VDD.n5489 GND 0.0147f
C6716 VDD.n5490 GND 0.0181f
C6717 VDD.t1329 GND 0.014f
C6718 VDD.n5491 GND 0.128f
C6719 VDD.n5492 GND 0.95f
C6720 VDD.t1316 GND 0.029f
C6721 VDD.t598 GND 0.0101f
C6722 VDD.n5493 GND 0.0529f
C6723 VDD.n5500 GND 0.0439f
C6724 VDD.n5501 GND 0.0168f
C6725 VDD.n5505 GND 0.0516f
C6726 VDD.n5507 GND 0.059f
C6727 VDD.t1299 GND 0.0218f
C6728 VDD.n5520 GND 0.03f
C6729 VDD.n5523 GND 0.0152f
C6730 VDD.n5524 GND 0.0101f
C6731 VDD.n5525 GND 0.0865f
C6732 VDD.n5526 GND 0.0289f
C6733 VDD.n5531 GND 0.0515f
C6734 VDD.n5533 GND 0.068f
C6735 VDD.n5541 GND 0.0655f
C6736 VDD.n5542 GND 0.0292f
C6737 VDD.n5547 GND 0.0317f
C6738 VDD.t596 GND 0.0515f
C6739 VDD.n5556 GND 0.223f
C6740 VDD.n5557 GND 0.125f
C6741 VDD.n5558 GND 0.0503f
C6742 VDD.n5559 GND 0.0163f
C6743 VDD.t667 GND 0.0647f
C6744 VDD.n5570 GND 0.0344f
C6745 VDD.n5571 GND 0.0851f
C6746 VDD.n5576 GND 0.0649f
C6747 VDD.n5577 GND 0.068f
C6748 VDD.n5585 GND 0.0323f
C6749 VDD.n5589 GND 0.0292f
C6750 VDD.t203 GND 0.0515f
C6751 VDD.n5598 GND 0.0515f
C6752 VDD.n5600 GND 0.0662f
C6753 VDD.n5601 GND 0.212f
C6754 VDD.n5602 GND 0.126f
C6755 VDD.n5603 GND 0.983f
C6756 VDD.n5604 GND 1.81f
C6757 VDD.n5605 GND 17.1f
C6758 VDD.n5606 GND 0.0179f
C6759 VDD.n5607 GND 0.035f
C6760 VDD.t707 GND 0.0452f
C6761 VDD.n5619 GND 0.0265f
C6762 VDD.n5627 GND 0.0331f
C6763 VDD.n5628 GND 0.0115f
C6764 VDD.n5636 GND 0.0381f
C6765 VDD.n5652 GND 0.0556f
C6766 VDD.t170 GND 0.0452f
C6767 VDD.n5653 GND 0.0265f
C6768 VDD.n5662 GND 0.0371f
C6769 VDD.n5664 GND 0.0102f
C6770 VDD.n5678 GND 0.0366f
C6771 VDD.n5679 GND 0.044f
C6772 VDD.n5685 GND 0.0442f
C6773 VDD.n5689 GND 0.0101f
C6774 VDD.n5690 GND 0.0356f
C6775 VDD.n5694 GND 0.0219f
C6776 VDD.n5695 GND 0.0102f
C6777 VDD.t4 GND 0.128f
C6778 VDD.n5705 GND 0.0556f
C6779 VDD.n5711 GND 0.0102f
C6780 VDD.n5712 GND 0.0217f
C6781 VDD.n5714 GND 0.0188f
C6782 VDD.n5715 GND 0.701f
C6783 VDD.n5716 GND 0.582f
C6784 VDD.n5742 GND 0.0336f
C6785 VDD.t168 GND 0.0141f
C6786 VDD.n5743 GND 0.0147f
C6787 VDD.n5744 GND 0.0181f
C6788 VDD.t704 GND 0.014f
C6789 VDD.n5745 GND 0.128f
C6790 VDD.n5746 GND 0.95f
C6791 VDD.t338 GND 0.029f
C6792 VDD.t712 GND 0.0101f
C6793 VDD.n5747 GND 0.0529f
C6794 VDD.n5754 GND 0.0439f
C6795 VDD.n5755 GND 0.0168f
C6796 VDD.n5759 GND 0.0516f
C6797 VDD.n5761 GND 0.059f
C6798 VDD.t1279 GND 0.0218f
C6799 VDD.n5774 GND 0.03f
C6800 VDD.n5777 GND 0.0152f
C6801 VDD.n5778 GND 0.0101f
C6802 VDD.n5779 GND 0.0865f
C6803 VDD.n5780 GND 0.0289f
C6804 VDD.n5785 GND 0.0515f
C6805 VDD.n5787 GND 0.068f
C6806 VDD.n5795 GND 0.0655f
C6807 VDD.n5796 GND 0.0292f
C6808 VDD.n5801 GND 0.0317f
C6809 VDD.t1088 GND 0.0515f
C6810 VDD.n5810 GND 0.223f
C6811 VDD.n5811 GND 0.125f
C6812 VDD.n5812 GND 0.0503f
C6813 VDD.n5813 GND 0.0163f
C6814 VDD.t419 GND 0.0647f
C6815 VDD.n5824 GND 0.0344f
C6816 VDD.n5825 GND 0.0851f
C6817 VDD.n5830 GND 0.0649f
C6818 VDD.n5831 GND 0.068f
C6819 VDD.n5839 GND 0.0323f
C6820 VDD.n5843 GND 0.0292f
C6821 VDD.t159 GND 0.0515f
C6822 VDD.n5852 GND 0.0515f
C6823 VDD.n5854 GND 0.0662f
C6824 VDD.n5855 GND 0.212f
C6825 VDD.n5856 GND 0.126f
C6826 VDD.n5857 GND 0.983f
C6827 VDD.n5858 GND 1.81f
C6828 VDD.n5859 GND 17.2f
C6829 VDD.n5860 GND 19f
C6830 VDD.n5861 GND 18.2f
C6831 VDD.n5862 GND 18.2f
C6832 VDD.n5863 GND 18.2f
C6833 VDD.n5864 GND 18.2f
C6834 VDD.n5865 GND 10.2f
C6835 VDD.n5866 GND 10.8f
C6836 VDD.n5867 GND 21.5f
C6837 VDD.n5868 GND 25.9f
C6838 VDD.n5869 GND 7.19f
C6839 VDD.n5870 GND 10.3f
.ends

