* NGSPICE file created from flashADC_flat.ext - technology: sky130A

.subckt flashADC_flat VFS OUT3 OUT2 OUT1 OUT0 VL VDD CLK VIN GND
X0 GND.t1394 frontAnalog_v0p0p1_7.x65.X frontAnalog_v0p0p1_7.RSfetsym_0.x2.Y GND.t1393 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 OUT3.t63 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD.t1330 VDD.t1329 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 VDD.t1185 frontAnalog_v0p0p1_15.x63.A.t4 a_57123_n85079# VDD.t1184 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X3 GND.t1224 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t127 GND.t1223 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 VDD.t178 frontAnalog_v0p0p1_10.x63.X frontAnalog_v0p0p1_10.Q.t1 VDD.t173 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.25
X5 VDD.t1023 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t63 VDD.t1022 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 VFS.t0 resistorDivider_v0p0p1_0.V16.t2 GND.t506 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X7 a_78315_n41309# 16to4_PriorityEncoder_v0p0p1_0.x5.x14.B a_78243_n41309# VDD.t556 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X8 a_16719_n13117.t19 a_16599_n13205.t4 a_16541_n13117.t18 GND.t213 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X9 w_55000_n56928# CLK.t0 frontAnalog_v0p0p1_10.x65.A.t2 VDD.t409 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X10 resistorDivider_v0p0p1_0.V4.t14 resistorDivider_v0p0p1_0.V3.t9 GND.t84 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X11 frontAnalog_v0p0p1_3.x65.X a_57123_n13359# VDD.t1501 VDD.t1500 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X12 VDD.t198 frontAnalog_v0p0p1_9.x63.X frontAnalog_v0p0p1_9.RSfetsym_0.x1.Y VDD.t191 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13 OUT3.t127 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND.t1385 GND.t1384 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X14 frontAnalog_v0p0p1_14.x65.A.t0 frontAnalog_v0p0p1_14.x63.A.t4 a_55268_n79536# GND.t1089 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X15 OUT2.t127 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND.t1077 GND.t1076 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X16 frontAnalog_v0p0p1_5.RSfetsym_0.QN.t3 frontAnalog_v0p0p1_5.RSfetsym_0.x1.Y GND.t1252 GND.t423 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.25
X17 16to4_PriorityEncoder_v0p0p1_0.x29.A 16to4_PriorityEncoder_v0p0p1_0.x28.A VDD.t71 VDD.t70 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X18 resistorDivider_v0p0p1_0.V11.t3 resistorDivider_v0p0p1_0.V10.t4 GND.t59 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X19 frontAnalog_v0p0p1_6.x63.X a_57123_n31079# GND.t586 GND.t585 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X20 GND.t1383 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t126 GND.t1382 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X21 GND.t567 frontAnalog_v0p0p1_8.x63.X frontAnalog_v0p0p1_8.RSfetsym_0.x1.Y GND.t562 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X22 GND.t1075 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t126 GND.t1074 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X23 OUT3.t62 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD.t1328 VDD.t1327 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X24 resistorDivider_v0p0p1_0.V2.t0 resistorDivider_v0p0p1_0.V1.t0 GND.t26 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X25 a_53630_n84996# resistorDivider_v0p0p1_0.V1.t16 w_55000_n83928# GND.t192 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X26 16to4_PriorityEncoder_v0p0p1_0.x29.Y 16to4_PriorityEncoder_v0p0p1_0.x29.A GND.t481 GND.t480 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X27 GND.t394 frontAnalog_v0p0p1_15.Q.t5 a_77605_n47345# GND.t65 sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X28 VDD.t1174 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t63 VDD.t1173 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X29 VDD.t1326 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t61 VDD.t1325 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X30 a_55268_n63336# CLK.t1 GND.t430 GND.t429 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X31 GND.t1504 16to4_PriorityEncoder_v0p0p1_0.x5.x17.A a_78349_n43045# GND.t252 sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X32 frontAnalog_v0p0p1_14.RSfetsym_0.x1.Y frontAnalog_v0p0p1_14.x63.X VDD.t584 VDD.t577 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X33 a_77605_n51335# frontAnalog_v0p0p1_12.Q.t5 VDD.t217 VDD.t216 sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.109 ps=1.36 w=0.42 l=0.15
X34 frontAnalog_v0p0p1_5.RSfetsym_0.x1.Y frontAnalog_v0p0p1_5.x63.X GND.t650 GND.t646 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X35 VDD.t177 frontAnalog_v0p0p1_10.x63.X frontAnalog_v0p0p1_10.RSfetsym_0.x1.Y VDD.t171 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X36 VDD.t782 VDD.t780 a_77605_n43295# VDD.t781 sky130_fd_pr__pfet_01v8_hvt ad=0.312 pd=1.68 as=0.0588 ps=0.7 w=0.42 l=0.15
X37 VDD.t380 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t63 VDD.t379 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X38 GND.t1381 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t125 GND.t1380 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X39 GND.t788 frontAnalog_v0p0p1_8.RSfetsym_0.QN.t5 a_59577_n46683# GND.t787 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X40 GND.t1073 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t125 GND.t1072 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X41 GND.t32 frontAnalog_v0p0p1_10.Q.t5 a_59578_n56970# GND.t31 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X42 a_53630_n41796# resistorDivider_v0p0p1_0.V9.t16 w_55000_n40728# GND.t70 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X43 VDD.t1021 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t62 VDD.t1020 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X44 resistorDivider_v0p0p1_0.V16.t15 resistorDivider_v0p0p1_0.V15.t15 GND.t102 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X45 OUT1.t127 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND.t393 GND.t392 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X46 GND.t101 frontAnalog_v0p0p1_12.x65.X frontAnalog_v0p0p1_12.RSfetsym_0.x2.Y GND.t100 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X47 OUT2.t61 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD.t1019 VDD.t1018 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X48 GND.t479 16to4_PriorityEncoder_v0p0p1_0.x29.A 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND.t478 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X49 frontAnalog_v0p0p1_7.RSfetsym_0.x1.Y frontAnalog_v0p0p1_7.x63.X VDD.t736 VDD.t729 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X50 OUT0.t126 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND.t1222 GND.t1221 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X51 a_77637_n50057# 16to4_PriorityEncoder_v0p0p1_0.x3.EI VDD.t812 VDD.t37 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X52 frontAnalog_v0p0p1_2.x65.A.t2 frontAnalog_v0p0p1_2.x63.A.t4 a_55268_n3936# GND.t679 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X53 VDD.t1378 frontAnalog_v0p0p1_15.x65.X frontAnalog_v0p0p1_15.RSfetsym_0.QN.t3 VDD.t1374 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.25
X54 GND.t1379 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t124 GND.t1378 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X55 GND.t1220 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t125 GND.t1219 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X56 a_82906_n51645# 16to4_PriorityEncoder_v0p0p1_0.x3.A0 GND.t880 GND.t879 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X57 OUT3.t60 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD.t1324 VDD.t1323 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X58 frontAnalog_v0p0p1_6.RSfetsym_0.QN.t3 frontAnalog_v0p0p1_6.Q.t5 VDD.t648 VDD.t647 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.3
X59 a_77881_n44527# 16to4_PriorityEncoder_v0p0p1_0.x5.x18.C a_77775_n44527# GND.t154 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X60 GND.t438 16to4_PriorityEncoder_v0p0p1_0.I13.t5 a_59578_n13770# GND.t437 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X61 OUT3.t123 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND.t1377 GND.t1376 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X62 16to4_PriorityEncoder_v0p0p1_0.x36.Y 16to4_PriorityEncoder_v0p0p1_0.x36.A GND.t1482 GND.t1481 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X63 a_53630_n9396# frontAnalog_v0p0p1_10.IB.t3 GND.t504 GND.t503 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X64 VDD.t1322 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t59 VDD.t1321 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X65 VDD.t609 frontAnalog_v0p0p1_2.x63.A.t5 a_57123_n4079# VDD.t608 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X66 frontAnalog_v0p0p1_11.x63.X a_57123_n63479# VDD.t895 VDD.t894 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X67 a_77723_n41087# VDD.t1502 a_77637_n41087# GND.t661 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X68 resistorDivider_v0p0p1_0.V14.t8 resistorDivider_v0p0p1_0.V13.t7 GND.t59 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X69 GND.t521 frontAnalog_v0p0p1_6.x65.X frontAnalog_v0p0p1_6.RSfetsym_0.x2.Y GND.t520 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X70 GND.t612 16to4_PriorityEncoder_v0p0p1_0.x21.A 16to4_PriorityEncoder_v0p0p1_0.x22.A GND.t611 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X71 w_55000_n79150# VIN.t0 a_53630_n79596# GND.t613 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X72 GND.t913 frontAnalog_v0p0p1_15.x63.X frontAnalog_v0p0p1_15.RSfetsym_0.x1.Y GND.t908 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X73 VIN.t1 w_55000_n51528# error sky130_fd_pr__cap_var_lvt w=2 l=0.18
X74 GND.t391 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t126 GND.t390 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X75 16to4_PriorityEncoder_v0p0p1_0.x5.x22.C a_77605_n44779# VDD.t748 VDD.t747 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.312 ps=1.68 w=1 l=0.15
X76 OUT2.t60 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD.t1017 VDD.t1016 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X77 resistorDivider_v0p0p1_0.V4.t10 resistorDivider_v0p0p1_0.V3.t6 GND.t399 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X78 16to4_PriorityEncoder_v0p0p1_0.x43.Y 16to4_PriorityEncoder_v0p0p1_0.x43.A VDD.t698 VDD.t697 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X79 VDD.t602 frontAnalog_v0p0p1_4.x65.A.t4 a_57123_n18759# VDD.t601 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X80 resistorDivider_v0p0p1_0.V10.t1 resistorDivider_v0p0p1_0.V9.t2 GND.t26 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X81 OUT0.t62 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD.t1172 VDD.t1171 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X82 a_78065_n41309# 16to4_PriorityEncoder_v0p0p1_0.x5.x22.A GND.t594 GND.t593 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X83 OUT0.t124 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND.t1218 GND.t1217 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X84 GND.t1216 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t123 GND.t1215 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X85 resistorDivider_v0p0p1_0.V3.t4 resistorDivider_v0p0p1_0.V2.t2 GND.t212 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X86 VDD.t811 16to4_PriorityEncoder_v0p0p1_0.x3.EI a_77605_n51335# VDD.t810 sky130_fd_pr__pfet_01v8_hvt ad=0.312 pd=1.68 as=0.0588 ps=0.7 w=0.42 l=0.15
X87 resistorDivider_v0p0p1_0.V13.t14 resistorDivider_v0p0p1_0.V12.t15 GND.t26 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X88 VDD.t1170 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t61 VDD.t1169 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X89 OUT3.t122 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND.t1375 GND.t1374 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X90 frontAnalog_v0p0p1_9.x65.A.t2 CLK.t2 frontAnalog_v0p0p1_9.x63.A.t2 VDD.t410 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X91 OUT2.t124 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND.t1071 GND.t1070 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X92 frontAnalog_v0p0p1_12.RSfetsym_0.x2.Y frontAnalog_v0p0p1_12.x65.X VDD.t79 VDD.t74 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X93 VDD.t1320 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t58 VDD.t1319 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X94 frontAnalog_v0p0p1_4.x63.X a_57123_n20279# VDD.t873 VDD.t872 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X95 GND.t389 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t125 GND.t388 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X96 w_55000_n35950# VIN.t2 a_53630_n36396# GND.t405 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X97 GND.t178 frontAnalog_v0p0p1_1.x63.X frontAnalog_v0p0p1_1.RSfetsym_0.x1.Y GND.t173 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X98 frontAnalog_v0p0p1_10.RSfetsym_0.x2.Y frontAnalog_v0p0p1_10.x65.X GND.t1446 GND.t1445 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X99 GND.t1373 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t121 GND.t1372 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X100 VDD.t547 frontAnalog_v0p0p1_10.Q.t6 a_77637_n49127# VDD.t546 sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X101 GND.t1480 16to4_PriorityEncoder_v0p0p1_0.x36.A 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND.t1479 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X102 VDD.t571 16to4_PriorityEncoder_v0p0p1_0.x21.A 16to4_PriorityEncoder_v0p0p1_0.x22.A VDD.t570 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X103 frontAnalog_v0p0p1_2.RSfetsym_0.x1.Y frontAnalog_v0p0p1_2.x63.X GND.t1412 GND.t1407 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X104 VDD.t1429 16to4_PriorityEncoder_v0p0p1_0.x36.A 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD.t1428 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X105 a_16541_n13117.t21 GND.t1402 GND.t799 sky130_fd_pr__res_xhigh_po_5p73 l=85.8
X106 frontAnalog_v0p0p1_14.Q.t4 frontAnalog_v0p0p1_14.RSfetsym_0.x2.Y GND.t1508 GND.t914 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.25
X107 GND.t483 frontAnalog_v0p0p1_9.x65.A.t4 a_57123_n51159# GND.t482 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X108 resistorDivider_v0p0p1_0.V3.t14 resistorDivider_v0p0p1_0.V2.t14 GND.t693 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X109 VDD.t416 16to4_PriorityEncoder_v0p0p1_0.I13.t6 a_77605_n45765# VDD.t415 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X110 a_77881_n52567# 16to4_PriorityEncoder_v0p0p1_0.x3.x18.C a_77775_n52567# GND.t131 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X111 16to4_PriorityEncoder_v0p0p1_0.x22.Y 16to4_PriorityEncoder_v0p0p1_0.x22.A GND.t1548 GND.t1547 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X112 frontAnalog_v0p0p1_9.x63.A.t0 frontAnalog_v0p0p1_9.x65.A.t5 a_55268_n52536# GND.t484 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X113 OUT2.t59 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD.t1015 VDD.t1014 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X114 OUT0.t60 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD.t1168 VDD.t1167 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X115 VDD.t1166 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t59 VDD.t1165 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X116 frontAnalog_v0p0p1_9.Q.t3 frontAnalog_v0p0p1_9.RSfetsym_0.QN.t5 VDD.t215 VDD.t214 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.3
X117 frontAnalog_v0p0p1_6.RSfetsym_0.x2.Y frontAnalog_v0p0p1_6.x65.X VDD.t480 VDD.t475 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X118 GND.t782 16to4_PriorityEncoder_v0p0p1_0.x43.A 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND.t781 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X119 GND.t387 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t124 GND.t386 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X120 OUT2.t58 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD.t1013 VDD.t1012 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X121 frontAnalog_v0p0p1_3.RSfetsym_0.x2.Y frontAnalog_v0p0p1_3.x65.X GND.t702 GND.t701 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X122 a_77639_n42341# VDD.t777 VDD.t779 VDD.t778 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X123 frontAnalog_v0p0p1_13.RSfetsym_0.x1.Y frontAnalog_v0p0p1_13.x63.X GND.t543 GND.t539 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X124 a_59577_n57483# frontAnalog_v0p0p1_10.x63.X frontAnalog_v0p0p1_10.Q.t2 GND.t185 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X125 a_59578_n67770# frontAnalog_v0p0p1_13.x65.X frontAnalog_v0p0p1_13.RSfetsym_0.QN.t2 GND.t141 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.315 ps=2.72 w=1 l=0.15
X126 a_77687_n45765# 16to4_PriorityEncoder_v0p0p1_0.I13.t7 a_77605_n45765# GND.t658 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X127 16to4_PriorityEncoder_v0p0p1_0.x42.A 16to4_PriorityEncoder_v0p0p1_0.x5.GS VDD.t1499 VDD.t1498 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X128 16to4_PriorityEncoder_v0p0p1_0.x3.x22.C a_77605_n52819# VDD.t712 VDD.t711 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.312 ps=1.68 w=1 l=0.15
X129 resistorDivider_v0p0p1_0.V2.t5 resistorDivider_v0p0p1_0.V1.t8 GND.t60 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X130 VDD.t1011 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t57 VDD.t1010 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X131 OUT1.t123 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND.t385 GND.t384 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X132 frontAnalog_v0p0p1_7.x63.A.t3 frontAnalog_v0p0p1_7.x65.A.t4 VDD.t1446 VDD.t18 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X133 frontAnalog_v0p0p1_7.Q.t4 frontAnalog_v0p0p1_7.RSfetsym_0.x2.Y GND.t1569 GND.t623 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.25
X134 resistorDivider_v0p0p1_0.V7.t16 w_55000_n52150# error sky130_fd_pr__cap_var_lvt w=2 l=0.18
X135 a_16719_n13117.t18 a_16599_n13205.t5 a_16541_n13117.t17 GND.t214 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X136 16to4_PriorityEncoder_v0p0p1_0.x5.x14.B a_77637_n41087# GND.t121 GND.t120 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.112 ps=1.04 w=0.65 l=0.15
X137 OUT0.t122 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND.t1214 GND.t1213 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X138 GND.t1449 16to4_PriorityEncoder_v0p0p1_0.x3.x14.A a_78065_n49349# GND.t1448 sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X139 a_78703_n45515# 16to4_PriorityEncoder_v0p0p1_0.x5.x22.C a_78607_n45515# VDD.t152 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X140 frontAnalog_v0p0p1_2.x65.X a_57123_n2559# GND.t225 GND.t224 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X141 16to4_PriorityEncoder_v0p0p1_0.x22.Y 16to4_PriorityEncoder_v0p0p1_0.x22.A VDD.t1481 VDD.t1480 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X142 a_16719_n13117.t21 a_16719_n13117.t20 a_16599_n13205.t2 GND.t916 sky130_fd_pr__nfet_01v8_lvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X143 resistorDivider_v0p0p1_0.V6.t15 resistorDivider_v0p0p1_0.V5.t15 GND.t506 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X144 VDD.t11 frontAnalog_v0p0p1_8.x65.X frontAnalog_v0p0p1_8.RSfetsym_0.x2.Y VDD.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X145 GND.t1371 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t120 GND.t1370 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X146 GND.t1546 16to4_PriorityEncoder_v0p0p1_0.x22.A 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND.t1545 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X147 VDD.t1009 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t56 VDD.t1008 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X148 VDD.t1187 frontAnalog_v0p0p1_13.x63.A.t4 a_57123_n68879# VDD.t1186 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X149 a_59577_n14283# frontAnalog_v0p0p1_3.x63.X 16to4_PriorityEncoder_v0p0p1_0.I13.t2 GND.t242 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X150 a_59578_n24570# frontAnalog_v0p0p1_5.x65.X frontAnalog_v0p0p1_5.RSfetsym_0.QN.t0 GND.t150 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.315 ps=2.72 w=1 l=0.15
X151 16to4_PriorityEncoder_v0p0p1_0.x29.Y 16to4_PriorityEncoder_v0p0p1_0.x29.A GND.t477 GND.t476 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X152 resistorDivider_v0p0p1_0.V7.t12 resistorDivider_v0p0p1_0.V6.t10 GND.t75 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X153 frontAnalog_v0p0p1_9.Q.t1 frontAnalog_v0p0p1_9.x63.X VDD.t197 VDD.t194 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.25
X154 a_53630_n63396# frontAnalog_v0p0p1_10.IB.t4 GND.t505 GND.t186 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X155 16to4_PriorityEncoder_v0p0p1_0.x5.x22.A a_77639_n42341# VDD.t573 VDD.t572 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.167 ps=1.39 w=1 l=0.15
X156 frontAnalog_v0p0p1_0.RSfetsym_0.x1.Y frontAnalog_v0p0p1_0.x63.X GND.t1559 GND.t1555 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X157 16to4_PriorityEncoder_v0p0p1_0.x43.Y 16to4_PriorityEncoder_v0p0p1_0.x43.A GND.t780 GND.t779 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X158 VDD.t239 frontAnalog_v0p0p1_10.x63.A.t4 frontAnalog_v0p0p1_10.x65.A.t0 VDD.t108 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X159 OUT2.t123 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND.t1069 GND.t1068 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X160 frontAnalog_v0p0p1_0.RSfetsym_0.x2.Y frontAnalog_v0p0p1_0.x65.X GND.t263 GND.t262 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X161 OUT1.t62 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD.t378 VDD.t377 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X162 w_55000_n8950# VIN.t3 a_53630_n9396# GND.t558 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X163 VDD.t549 frontAnalog_v0p0p1_10.Q.t7 a_77605_n53805# VDD.t548 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X164 frontAnalog_v0p0p1_12.x65.X a_57123_n72759# GND.t926 GND.t17 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X165 VDD.t376 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t61 VDD.t375 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X166 OUT0.t58 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD.t1164 VDD.t1163 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X167 frontAnalog_v0p0p1_4.RSfetsym_0.x2.Y frontAnalog_v0p0p1_4.x65.X GND.t903 GND.t902 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X168 GND.t1369 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t119 GND.t1368 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X169 VDD.t407 frontAnalog_v0p0p1_5.x63.A.t4 a_57123_n25679# VDD.t406 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X170 GND.t1212 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t121 GND.t1211 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X171 a_53630_n20196# frontAnalog_v0p0p1_10.IB.t5 GND.t441 GND.t186 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X172 a_77639_n50381# 16to4_PriorityEncoder_v0p0p1_0.x3.EI VDD.t809 VDD.t808 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X173 VDD.t1427 16to4_PriorityEncoder_v0p0p1_0.x36.A 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD.t1426 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X174 VDD.t1479 16to4_PriorityEncoder_v0p0p1_0.x22.A 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD.t1478 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X175 VDD.t817 frontAnalog_v0p0p1_3.x63.A.t4 frontAnalog_v0p0p1_3.x65.A.t2 VDD.t485 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X176 OUT3.t118 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND.t1367 GND.t1366 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X177 VDD.t237 frontAnalog_v0p0p1_15.x65.A.t4 a_57123_n83559# VDD.t236 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X178 GND.t1090 frontAnalog_v0p0p1_14.x63.A.t5 a_57123_n79679# GND.t433 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X179 a_55268_n47136# CLK.t3 GND.t432 GND.t431 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X180 frontAnalog_v0p0p1_1.RSfetsym_0.x2.Y frontAnalog_v0p0p1_1.x65.X GND.t688 GND.t687 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X181 VDD.t78 frontAnalog_v0p0p1_12.x65.X frontAnalog_v0p0p1_12.RSfetsym_0.x2.Y VDD.t74 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X182 GND.t221 16to4_PriorityEncoder_v0p0p1_0.x3.x17.C a_78349_n51085# GND.t165 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X183 frontAnalog_v0p0p1_4.x65.A.t2 frontAnalog_v0p0p1_4.x63.A.t4 a_55268_n20136# GND.t1241 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X184 frontAnalog_v0p0p1_9.RSfetsym_0.QN.t4 frontAnalog_v0p0p1_9.Q.t5 VDD.t1445 VDD.t214 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.3
X185 OUT3.t57 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD.t1318 VDD.t1317 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X186 resistorDivider_v0p0p1_0.V10.t0 resistorDivider_v0p0p1_0.V9.t1 GND.t60 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X187 a_78703_n53555# 16to4_PriorityEncoder_v0p0p1_0.x3.x22.C a_78607_n53555# VDD.t574 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X188 GND.t1210 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t120 GND.t1209 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X189 OUT1.t122 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND.t383 GND.t382 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X190 resistorDivider_v0p0p1_0.V12.t9 resistorDivider_v0p0p1_0.V11.t9 GND.t211 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X191 resistorDivider_v0p0p1_0.V3.t10 resistorDivider_v0p0p1_0.V2.t9 GND.t615 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X192 a_77775_n51335# 16to4_PriorityEncoder_v0p0p1_0.x3.x19.C a_77687_n51335# GND.t157 sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
X193 16to4_PriorityEncoder_v0p0p1_0.x43.A 16to4_PriorityEncoder_v0p0p1_0.x42.A VDD.t662 VDD.t661 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X194 a_53630_n25596# resistorDivider_v0p0p1_0.V12.t16 w_55000_n24528# GND.t63 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X195 resistorDivider_v0p0p1_0.V13.t4 resistorDivider_v0p0p1_0.V12.t3 GND.t60 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X196 OUT3.t117 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND.t1365 GND.t1364 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X197 16to4_PriorityEncoder_v0p0p1_0.x28.A 16to4_PriorityEncoder_v0p0p1_0.x1.X GND.t883 GND.t882 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X198 VDD.t1162 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t57 VDD.t1161 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X199 VDD.t1007 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t55 VDD.t1006 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X200 frontAnalog_v0p0p1_9.RSfetsym_0.x2.Y frontAnalog_v0p0p1_9.x65.X VDD.t638 VDD.t633 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X201 VDD.t1196 frontAnalog_v0p0p1_1.x65.A.t4 a_57123_n40359# VDD.t1195 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X202 GND.t733 frontAnalog_v0p0p1_7.x63.A.t4 a_57123_n36479# GND.t732 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X203 frontAnalog_v0p0p1_10.RSfetsym_0.QN.t3 frontAnalog_v0p0p1_10.x65.X VDD.t1390 VDD.t1386 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.25
X204 frontAnalog_v0p0p1_9.RSfetsym_0.x1.Y frontAnalog_v0p0p1_9.x63.X GND.t205 GND.t200 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X205 VDD.t479 frontAnalog_v0p0p1_6.x65.X frontAnalog_v0p0p1_6.RSfetsym_0.x2.Y VDD.t475 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X206 16to4_PriorityEncoder_v0p0p1_0.x36.Y 16to4_PriorityEncoder_v0p0p1_0.x36.A VDD.t1425 VDD.t1424 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X207 VDD.t1202 frontAnalog_v0p0p1_11.Q.t5 a_77637_n48817# VDD.t1201 sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X208 VDD.t374 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t60 VDD.t373 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X209 VDD.t130 frontAnalog_v0p0p1_13.x65.X frontAnalog_v0p0p1_13.RSfetsym_0.QN.t1 VDD.t126 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.25
X210 GND.t1208 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t119 GND.t1207 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X211 VDD.t1160 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t56 VDD.t1159 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X212 frontAnalog_v0p0p1_11.RSfetsym_0.x1.Y frontAnalog_v0p0p1_11.x63.X VDD.t99 VDD.t94 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X213 OUT0.t118 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND.t1206 GND.t1205 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X214 VFS.t3 resistorDivider_v0p0p1_0.V16.t6 GND.t196 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X215 frontAnalog_v0p0p1_3.RSfetsym_0.QN.t3 frontAnalog_v0p0p1_3.x65.X VDD.t628 VDD.t624 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.25
X216 VDD.t660 16to4_PriorityEncoder_v0p0p1_0.x42.A 16to4_PriorityEncoder_v0p0p1_0.x43.A VDD.t659 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X217 VDD.t372 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t59 VDD.t371 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X218 resistorDivider_v0p0p1_0.V4.t8 resistorDivider_v0p0p1_0.V3.t5 GND.t102 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X219 resistorDivider_v0p0p1_0.V15.t16 w_55000_n8950# error sky130_fd_pr__cap_var_lvt w=2 l=0.18
X220 16to4_PriorityEncoder_v0p0p1_0.x5.x17.A a_77637_n42017# GND.t928 GND.t927 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.112 ps=1.04 w=0.65 l=0.15
X221 VDD.t138 frontAnalog_v0p0p1_5.x65.X frontAnalog_v0p0p1_5.RSfetsym_0.QN.t2 VDD.t134 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.25
X222 resistorDivider_v0p0p1_0.V15.t10 resistorDivider_v0p0p1_0.V14.t12 GND.t84 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X223 GND.t1558 frontAnalog_v0p0p1_0.x63.X frontAnalog_v0p0p1_0.RSfetsym_0.x1.Y GND.t1555 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X224 VDD.t1316 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t56 VDD.t1315 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X225 16to4_PriorityEncoder_v0p0p1_0.x22.Y 16to4_PriorityEncoder_v0p0p1_0.x22.A GND.t1544 GND.t1543 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X226 VDD.t1158 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t55 VDD.t1157 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X227 a_16719_n13117.t17 a_16599_n13205.t6 a_16541_n13117.t16 GND.t215 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X228 frontAnalog_v0p0p1_7.x65.A.t0 CLK.t4 frontAnalog_v0p0p1_7.x63.A.t1 VDD.t411 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X229 resistorDivider_v0p0p1_0.V7.t7 resistorDivider_v0p0p1_0.V6.t4 GND.t119 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X230 VDD.t583 frontAnalog_v0p0p1_14.x63.X frontAnalog_v0p0p1_14.RSfetsym_0.x1.Y VDD.t577 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X231 frontAnalog_v0p0p1_6.x63.A.t3 CLK.t5 w_55000_n30550# VDD.t412 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X232 GND.t649 frontAnalog_v0p0p1_5.x63.X frontAnalog_v0p0p1_5.RSfetsym_0.x1.Y GND.t646 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X233 OUT2.t54 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD.t1005 VDD.t1004 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X234 OUT0.t54 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD.t1156 VDD.t1155 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X235 a_78607_n45515# 16to4_PriorityEncoder_v0p0p1_0.x5.x22.D a_78525_n45515# VDD.t161 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X236 VDD.t27 frontAnalog_v0p0p1_2.x65.A.t4 a_57123_n2559# VDD.t26 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X237 frontAnalog_v0p0p1_11.x65.X a_57123_n61959# VDD.t605 VDD.t604 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X238 GND.t901 frontAnalog_v0p0p1_4.x65.X frontAnalog_v0p0p1_4.RSfetsym_0.x2.Y GND.t900 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X239 frontAnalog_v0p0p1_10.x63.X a_57123_n58079# GND.t486 GND.t485 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X240 OUT1.t58 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD.t370 VDD.t369 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X241 frontAnalog_v0p0p1_9.x63.A.t3 CLK.t6 w_55000_n52150# VDD.t413 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X242 VDD.t1350 CLK.t7 w_55000_n73128# GND.t125 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X243 GND.t1512 frontAnalog_v0p0p1_7.x65.A.t5 a_57123_n34959# GND.t732 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X244 frontAnalog_v0p0p1_12.RSfetsym_0.QN.t4 frontAnalog_v0p0p1_12.RSfetsym_0.x1.Y GND.t1493 GND.t1403 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.25
X245 GND.t1067 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t122 GND.t1066 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X246 16to4_PriorityEncoder_v0p0p1_0.x5.x17.D a_77605_n43545# GND.t164 GND.t163 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.196 ps=1.33 w=0.65 l=0.15
X247 GND.t365 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t121 GND.t364 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X248 GND.t686 frontAnalog_v0p0p1_1.x65.X frontAnalog_v0p0p1_1.RSfetsym_0.x2.Y GND.t685 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X249 frontAnalog_v0p0p1_15.RSfetsym_0.x2.Y frontAnalog_v0p0p1_15.x65.X GND.t1428 GND.t1427 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X250 frontAnalog_v0p0p1_3.RSfetsym_0.x2.Y frontAnalog_v0p0p1_3.x65.X VDD.t627 VDD.t621 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X251 VDD.t735 frontAnalog_v0p0p1_7.x63.X frontAnalog_v0p0p1_7.RSfetsym_0.x1.Y VDD.t729 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X252 VDD.t98 frontAnalog_v0p0p1_11.x63.X frontAnalog_v0p0p1_11.Q.t2 VDD.t92 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.25
X253 VDD.t1351 CLK.t8 w_55000_n73750# GND.t132 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X254 16to4_PriorityEncoder_v0p0p1_0.x22.Y 16to4_PriorityEncoder_v0p0p1_0.x22.A VDD.t1477 VDD.t1476 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X255 resistorDivider_v0p0p1_0.V1.t2 VL.t0 GND.t26 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X256 w_55000_n62328# CLK.t9 frontAnalog_v0p0p1_11.x65.A.t2 VDD.t727 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X257 a_78243_n41309# 16to4_PriorityEncoder_v0p0p1_0.x5.x17.A a_78147_n41309# VDD.t556 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X258 OUT2.t53 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD.t983 VDD.t982 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X259 VDD.t776 VDD.t774 a_78649_n39527# VDD.t775 sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X260 frontAnalog_v0p0p1_3.x63.X a_57123_n14879# GND.t1432 GND.t1431 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X261 OUT3.t116 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND.t1363 GND.t1362 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X262 resistorDivider_v0p0p1_0.V10.t16 w_55000_n35950# error sky130_fd_pr__cap_var_lvt w=2 l=0.18
X263 frontAnalog_v0p0p1_15.x65.A.t0 frontAnalog_v0p0p1_15.x63.A.t5 a_55268_n84936# GND.t500 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X264 a_53630_n68796# resistorDivider_v0p0p1_0.V4.t16 w_55000_n67728# GND.t61 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X265 VDD.t1003 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t52 VDD.t1002 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X266 resistorDivider_v0p0p1_0.V9.t0 resistorDivider_v0p0p1_0.V8.t2 GND.t26 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X267 VDD.t1314 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t55 VDD.t1313 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X268 16to4_PriorityEncoder_v0p0p1_0.x3.x17.A a_77637_n50057# GND.t229 GND.t228 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.112 ps=1.04 w=0.65 l=0.15
X269 OUT0.t117 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND.t1204 GND.t1203 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X270 GND.t1361 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t115 GND.t1360 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X271 GND.t204 frontAnalog_v0p0p1_9.x63.X frontAnalog_v0p0p1_9.RSfetsym_0.x1.Y GND.t200 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X272 OUT3.t54 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD.t1312 VDD.t1311 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X273 16to4_PriorityEncoder_v0p0p1_0.x21.A 16to4_PriorityEncoder_v0p0p1_0.x2.X GND.t560 GND.t559 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X274 VIN.t4 w_55000_n8328# error sky130_fd_pr__cap_var_lvt w=2 l=0.18
X275 GND.t1551 16to4_PriorityEncoder_v0p0p1_0.x5.x21.B a_78183_n45737# GND.t1550 sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X276 VDD.t1352 CLK.t10 w_55000_n30550# GND.t527 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X277 VDD.t62 frontAnalog_v0p0p1_4.x63.X 16to4_PriorityEncoder_v0p0p1_0.I12.t1 VDD.t55 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.25
X278 w_55000_n19128# CLK.t11 frontAnalog_v0p0p1_4.x65.A.t1 VDD.t184 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X279 VDD.t696 16to4_PriorityEncoder_v0p0p1_0.x43.A 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD.t695 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X280 GND.t748 16to4_PriorityEncoder_v0p0p1_0.x42.A 16to4_PriorityEncoder_v0p0p1_0.x43.A GND.t747 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X281 GND.t1065 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t121 GND.t1064 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X282 a_78607_n53555# 16to4_PriorityEncoder_v0p0p1_0.x3.x22.D a_78525_n53555# VDD.t620 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X283 frontAnalog_v0p0p1_1.x65.A.t2 frontAnalog_v0p0p1_1.x63.A.t4 a_55268_n41736# GND.t947 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X284 OUT2.t120 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND.t1063 GND.t1062 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X285 VDD.t97 frontAnalog_v0p0p1_11.x63.X frontAnalog_v0p0p1_11.RSfetsym_0.x1.Y VDD.t94 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X286 GND.t381 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t120 GND.t380 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X287 resistorDivider_v0p0p1_0.V15.t14 resistorDivider_v0p0p1_0.V14.t14 GND.t399 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X288 16to4_PriorityEncoder_v0p0p1_0.x3.x16.C frontAnalog_v0p0p1_10.Q.t8 GND.t588 GND.t587 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X289 OUT0.t53 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD.t1154 VDD.t1153 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X290 OUT3.t53 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD.t1310 VDD.t1309 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X291 GND.t1444 frontAnalog_v0p0p1_10.x65.X frontAnalog_v0p0p1_10.RSfetsym_0.x2.Y GND.t1443 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X292 VIN.t5 w_55000_n78528# error sky130_fd_pr__cap_var_lvt w=2 l=0.18
X293 OUT1.t119 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND.t379 GND.t378 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X294 frontAnalog_v0p0p1_4.RSfetsym_0.x1.Y frontAnalog_v0p0p1_4.x63.X VDD.t61 VDD.t57 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X295 VDD.t399 16to4_PriorityEncoder_v0p0p1_0.x1.A a_82988_n47995# VDD.t398 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X296 GND.t1411 frontAnalog_v0p0p1_2.x63.X frontAnalog_v0p0p1_2.RSfetsym_0.x1.Y GND.t1407 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X297 16to4_PriorityEncoder_v0p0p1_0.x21.A 16to4_PriorityEncoder_v0p0p1_0.x2.X VDD.t513 VDD.t512 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X298 a_77687_n44779# VDD.t1503 a_77605_n44779# GND.t155 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.109 ps=1.36 w=0.42 l=0.15
X299 a_77723_n42017# VDD.t1504 a_77637_n42017# GND.t662 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X300 VDD.t807 16to4_PriorityEncoder_v0p0p1_0.x3.EI a_78649_n47567# VDD.t806 sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X301 GND.t1061 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t119 GND.t1060 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X302 OUT2.t118 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND.t1059 GND.t1058 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X303 frontAnalog_v0p0p1_14.x65.A.t2 CLK.t12 frontAnalog_v0p0p1_14.x63.A.t1 VDD.t1353 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X304 OUT2.t51 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD.t1001 VDD.t1000 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X305 16to4_PriorityEncoder_v0p0p1_0.x43.Y 16to4_PriorityEncoder_v0p0p1_0.x43.A VDD.t694 VDD.t693 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X306 frontAnalog_v0p0p1_8.x63.X a_57123_n47279# VDD.t1487 VDD.t1486 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X307 GND.t700 frontAnalog_v0p0p1_3.x65.X frontAnalog_v0p0p1_3.RSfetsym_0.x2.Y GND.t699 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X308 VIN.t6 w_55000_n35328# error sky130_fd_pr__cap_var_lvt w=2 l=0.18
X309 GND.t542 frontAnalog_v0p0p1_13.x63.X frontAnalog_v0p0p1_13.RSfetsym_0.x1.Y GND.t539 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X310 16to4_PriorityEncoder_v0p0p1_0.x43.Y 16to4_PriorityEncoder_v0p0p1_0.x43.A GND.t778 GND.t777 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X311 OUT1.t118 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND.t377 GND.t376 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X312 VDD.t999 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t50 VDD.t998 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X313 VDD.t1308 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t52 VDD.t1307 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X314 GND.t571 16to4_PriorityEncoder_v0p0p1_0.x3.x21.B a_78183_n53777# GND.t570 sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X315 a_53630_n74196# frontAnalog_v0p0p1_10.IB.t6 GND.t442 GND.t186 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X316 w_55000_n84550# VIN.t7 a_53630_n84996# GND.t192 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X317 GND.t434 frontAnalog_v0p0p1_14.x65.A.t4 a_57123_n78159# GND.t433 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X318 OUT2.t117 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND.t1057 GND.t1056 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X319 VDD.t1025 frontAnalog_v0p0p1_5.x65.A.t4 a_57123_n24159# VDD.t1024 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X320 GND.t1242 frontAnalog_v0p0p1_4.x63.A.t5 a_57123_n20279# GND.t197 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X321 frontAnalog_v0p0p1_14.x63.A.t2 frontAnalog_v0p0p1_14.x65.A.t5 a_55268_n79536# GND.t822 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X322 GND.t1426 frontAnalog_v0p0p1_15.x65.X frontAnalog_v0p0p1_15.RSfetsym_0.x2.Y GND.t1425 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X323 VDD.t368 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t57 VDD.t367 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X324 VDD.t626 frontAnalog_v0p0p1_3.x65.X frontAnalog_v0p0p1_3.RSfetsym_0.x2.Y VDD.t621 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X325 GND.t1359 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t114 GND.t1358 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X326 frontAnalog_v0p0p1_14.Q.t3 frontAnalog_v0p0p1_14.RSfetsym_0.QN.t5 VDD.t1035 VDD.t532 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.3
X327 frontAnalog_v0p0p1_10.RSfetsym_0.x2.Y frontAnalog_v0p0p1_10.x65.X VDD.t1389 VDD.t1383 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X328 GND.t1202 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t116 GND.t1201 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X329 GND.t1478 16to4_PriorityEncoder_v0p0p1_0.x36.A 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND.t1477 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X330 w_55000_n19750# VIN.t8 a_53630_n20196# GND.t69 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X331 VDD.t1423 16to4_PriorityEncoder_v0p0p1_0.x36.A 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD.t1422 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X332 OUT3.t113 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND.t1357 GND.t1356 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X333 a_77881_n43295# 16to4_PriorityEncoder_v0p0p1_0.x5.x16.C a_77775_n43295# GND.t156 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X334 resistorDivider_v0p0p1_0.V6.t9 resistorDivider_v0p0p1_0.V5.t11 GND.t196 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X335 VDD.t997 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t49 VDD.t996 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X336 VDD.t1306 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t51 VDD.t1305 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X337 resistorDivider_v0p0p1_0.V2.t1 resistorDivider_v0p0p1_0.V1.t1 GND.t59 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X338 GND.t475 16to4_PriorityEncoder_v0p0p1_0.x29.A 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND.t474 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X339 resistorDivider_v0p0p1_0.V2.t16 w_55000_n79150# error sky130_fd_pr__cap_var_lvt w=2 l=0.18
X340 w_55000_n41350# VIN.t9 a_53630_n41796# GND.t70 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X341 GND.t261 frontAnalog_v0p0p1_0.x65.X frontAnalog_v0p0p1_0.RSfetsym_0.x2.Y GND.t260 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X342 frontAnalog_v0p0p1_11.RSfetsym_0.x2.Y frontAnalog_v0p0p1_11.x65.X GND.t946 GND.t945 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X343 a_77723_n50057# 16to4_PriorityEncoder_v0p0p1_0.x3.EI a_77637_n50057# GND.t867 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X344 GND.t907 16to4_PriorityEncoder_v0p0p1_0.x5.x20.B a_77881_n44779# GND.t155 sky130_fd_pr__nfet_01v8 ad=0.196 pd=1.33 as=0.0693 ps=0.75 w=0.42 l=0.15
X345 frontAnalog_v0p0p1_7.x63.A.t2 frontAnalog_v0p0p1_7.x65.A.t6 a_55268_n36336# GND.t1513 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X346 resistorDivider_v0p0p1_0.V1.t9 VL.t4 GND.t60 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X347 resistorDivider_v0p0p1_0.V11.t2 resistorDivider_v0p0p1_0.V10.t3 GND.t84 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X348 frontAnalog_v0p0p1_15.Q.t1 frontAnalog_v0p0p1_15.RSfetsym_0.x2.Y GND.t821 GND.t820 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.25
X349 OUT1.t117 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND.t375 GND.t374 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X350 a_77775_n44527# frontAnalog_v0p0p1_7.Q.t5 a_77687_n44527# GND.t154 sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
X351 frontAnalog_v0p0p1_7.Q.t0 frontAnalog_v0p0p1_7.RSfetsym_0.QN.t5 VDD.t190 VDD.t30 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.3
X352 a_59578_n8370# frontAnalog_v0p0p1_0.x65.X frontAnalog_v0p0p1_0.RSfetsym_0.QN.t1 GND.t259 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.315 ps=2.72 w=1 l=0.15
X353 GND.t1055 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t116 GND.t1054 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X354 VDD.t995 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t48 VDD.t994 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X355 a_78147_n41309# 16to4_PriorityEncoder_v0p0p1_0.x5.x22.A a_78065_n41309# VDD.t556 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X356 VDD.t1152 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t52 VDD.t1151 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X357 OUT1.t116 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND.t373 GND.t372 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X358 OUT3.t112 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND.t1355 GND.t1354 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X359 frontAnalog_v0p0p1_14.Q.t2 frontAnalog_v0p0p1_14.x63.X VDD.t582 VDD.t579 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.25
X360 resistorDivider_v0p0p1_0.V9.t6 resistorDivider_v0p0p1_0.V8.t9 GND.t60 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X361 16to4_PriorityEncoder_v0p0p1_0.x36.Y 16to4_PriorityEncoder_v0p0p1_0.x36.A GND.t1476 GND.t1475 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X362 16to4_PriorityEncoder_v0p0p1_0.x36.Y 16to4_PriorityEncoder_v0p0p1_0.x36.A VDD.t1421 VDD.t1420 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X363 GND.t371 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t115 GND.t370 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X364 frontAnalog_v0p0p1_12.RSfetsym_0.x1.Y frontAnalog_v0p0p1_12.x63.X GND.t644 GND.t640 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X365 a_59577_n62883# frontAnalog_v0p0p1_11.x63.X frontAnalog_v0p0p1_11.Q.t0 GND.t118 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X366 frontAnalog_v0p0p1_1.Q.t3 frontAnalog_v0p0p1_1.RSfetsym_0.x2.Y GND.t254 GND.t0 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.25
X367 GND.t1200 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t115 GND.t1199 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X368 16to4_PriorityEncoder_v0p0p1_0.x3.x17.C a_77605_n51335# GND.t152 GND.t151 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.196 ps=1.33 w=0.65 l=0.15
X369 16to4_PriorityEncoder_v0p0p1_0.x43.Y 16to4_PriorityEncoder_v0p0p1_0.x43.A GND.t776 GND.t775 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X370 OUT0.t114 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND.t1198 GND.t1197 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X371 VDD.t1354 CLK.t13 w_55000_n56928# GND.t833 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X372 GND.t369 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t114 GND.t368 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X373 a_53630_n47196# frontAnalog_v0p0p1_10.IB.t7 GND.t443 GND.t186 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X374 frontAnalog_v0p0p1_7.Q.t2 frontAnalog_v0p0p1_7.x63.X VDD.t734 VDD.t731 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.25
X375 OUT1.t56 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD.t366 VDD.t365 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X376 frontAnalog_v0p0p1_15.RSfetsym_0.x1.Y frontAnalog_v0p0p1_15.x63.X VDD.t862 VDD.t855 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X377 VDD.t637 frontAnalog_v0p0p1_9.x65.X frontAnalog_v0p0p1_9.RSfetsym_0.x2.Y VDD.t633 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X378 VDD.t893 frontAnalog_v0p0p1_1.x63.A.t5 frontAnalog_v0p0p1_1.x65.A.t3 VDD.t109 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X379 OUT2.t47 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD.t993 VDD.t992 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X380 frontAnalog_v0p0p1_6.RSfetsym_0.x1.Y frontAnalog_v0p0p1_6.x63.X GND.t44 GND.t40 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X381 frontAnalog_v0p0p1_13.RSfetsym_0.x2.Y frontAnalog_v0p0p1_13.x65.X GND.t140 GND.t139 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X382 16to4_PriorityEncoder_v0p0p1_0.x5.x14.A a_77637_n40777# VDD.t213 VDD.t212 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.167 ps=1.39 w=1 l=0.15
X383 VDD.t364 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t55 VDD.t363 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X384 16to4_PriorityEncoder_v0p0p1_0.x34.A a_82906_n43855# VDD.t1368 VDD.t1367 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.146 ps=1.34 w=1 l=0.15
X385 frontAnalog_v0p0p1_14.RSfetsym_0.QN.t4 frontAnalog_v0p0p1_14.Q.t5 VDD.t533 VDD.t532 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.3
X386 frontAnalog_v0p0p1_10.x65.X a_57123_n56559# GND.t924 GND.t485 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X387 GND.t1256 frontAnalog_v0p0p1_11.Q.t6 a_59578_n62370# GND.t1255 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X388 GND.t232 frontAnalog_v0p0p1_9.RSfetsym_0.QN.t6 a_59577_n52083# GND.t231 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X389 GND.t1351 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t111 GND.t1350 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X390 16to4_PriorityEncoder_v0p0p1_0.x5.x9.Y VDD.t1505 GND.t664 GND.t663 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X391 a_77775_n52567# frontAnalog_v0p0p1_14.Q.t6 a_77687_n52567# GND.t131 sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
X392 resistorDivider_v0p0p1_0.V10.t15 resistorDivider_v0p0p1_0.V9.t15 GND.t59 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X393 a_16719_n13117.t16 a_16599_n13205.t7 a_16541_n13117.t5 GND.t216 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X394 VDD.t1150 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t51 VDD.t1149 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X395 VDD.t69 16to4_PriorityEncoder_v0p0p1_0.x28.A 16to4_PriorityEncoder_v0p0p1_0.x29.A VDD.t68 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X396 VDD.t649 CLK.t14 w_55000_n13728# GND.t736 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X397 OUT3.t110 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND.t1353 GND.t1352 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X398 resistorDivider_v0p0p1_0.V3.t13 resistorDivider_v0p0p1_0.V2.t13 GND.t211 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X399 OUT0.t113 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND.t1196 GND.t1195 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X400 OUT2.t115 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND.t1053 GND.t1052 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X401 resistorDivider_v0p0p1_0.V14.t7 resistorDivider_v0p0p1_0.V13.t6 GND.t84 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X402 resistorDivider_v0p0p1_0.V13.t8 resistorDivider_v0p0p1_0.V12.t8 GND.t59 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X403 16to4_PriorityEncoder_v0p0p1_0.x36.A 16to4_PriorityEncoder_v0p0p1_0.x35.A GND.t55 GND.t54 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X404 VDD.t1304 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t50 VDD.t1303 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X405 OUT0.t50 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD.t1148 VDD.t1147 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X406 GND.t473 16to4_PriorityEncoder_v0p0p1_0.x29.A 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND.t472 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X407 OUT2.t46 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD.t991 VDD.t990 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X408 frontAnalog_v0p0p1_1.RSfetsym_0.x1.Y frontAnalog_v0p0p1_1.x63.X VDD.t169 VDD.t162 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X409 frontAnalog_v0p0p1_14.RSfetsym_0.x2.Y frontAnalog_v0p0p1_14.x65.X VDD.t790 VDD.t785 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X410 GND.t1349 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t109 GND.t1348 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X411 GND.t774 16to4_PriorityEncoder_v0p0p1_0.x43.A 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND.t773 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X412 frontAnalog_v0p0p1_5.RSfetsym_0.x2.Y frontAnalog_v0p0p1_5.x65.X GND.t149 GND.t148 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X413 VDD.t883 frontAnalog_v0p0p1_13.x65.A.t4 a_57123_n67359# VDD.t882 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X414 frontAnalog_v0p0p1_14.RSfetsym_0.x1.Y frontAnalog_v0p0p1_14.x63.X GND.t638 GND.t633 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X415 VDD.t650 CLK.t15 w_55000_n14350# GND.t127 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X416 16to4_PriorityEncoder_v0p0p1_0.x5.x17.D a_77605_n43545# VDD.t156 VDD.t155 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.312 ps=1.68 w=1 l=0.15
X417 VDD.t1388 frontAnalog_v0p0p1_10.x65.X frontAnalog_v0p0p1_10.RSfetsym_0.x2.Y VDD.t1383 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X418 OUT1.t54 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD.t362 VDD.t361 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X419 VDD.t360 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t53 VDD.t359 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X420 frontAnalog_v0p0p1_7.RSfetsym_0.QN.t4 frontAnalog_v0p0p1_7.Q.t6 VDD.t31 VDD.t30 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.3
X421 frontAnalog_v0p0p1_3.x65.X a_57123_n13359# GND.t1567 GND.t1431 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X422 GND.t74 frontAnalog_v0p0p1_15.x63.A.t6 a_57123_n85079# GND.t73 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X423 resistorDivider_v0p0p1_0.V11.t1 resistorDivider_v0p0p1_0.V10.t2 GND.t399 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X424 OUT3.t108 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND.t1347 GND.t1346 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X425 VDD.t534 frontAnalog_v0p0p1_14.Q.t7 a_77605_n52567# VDD.t114 sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X426 resistorDivider_v0p0p1_0.V15.t3 resistorDivider_v0p0p1_0.V14.t4 GND.t102 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X427 GND.t1542 16to4_PriorityEncoder_v0p0p1_0.x22.A 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND.t1541 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X428 OUT2.t45 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD.t989 VDD.t988 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X429 frontAnalog_v0p0p1_7.RSfetsym_0.x2.Y frontAnalog_v0p0p1_7.x65.X VDD.t1338 VDD.t1333 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X430 OUT0.t49 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD.t1146 VDD.t1145 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X431 GND.t367 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t113 GND.t366 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X432 frontAnalog_v0p0p1_7.RSfetsym_0.x1.Y frontAnalog_v0p0p1_7.x63.X GND.t815 GND.t810 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X433 VDD.t987 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t44 VDD.t986 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X434 16to4_PriorityEncoder_v0p0p1_0.x29.Y 16to4_PriorityEncoder_v0p0p1_0.x29.A GND.t471 GND.t470 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X435 OUT0.t112 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND.t1194 GND.t1193 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X436 16to4_PriorityEncoder_v0p0p1_0.x29.Y 16to4_PriorityEncoder_v0p0p1_0.x29.A VDD.t456 VDD.t455 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X437 GND.t112 frontAnalog_v0p0p1_1.x63.A.t6 a_57123_n41879# GND.t111 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X438 frontAnalog_v0p0p1_11.RSfetsym_0.QN.t3 frontAnalog_v0p0p1_11.x65.X VDD.t892 VDD.t888 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.25
X439 VDD.t38 frontAnalog_v0p0p1_9.Q.t6 a_77637_n50057# VDD.t37 sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X440 a_16719_n13117.t15 a_16599_n13205.t8 a_16541_n13117.t4 GND.t217 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X441 frontAnalog_v0p0p1_2.RSfetsym_0.x2.Y frontAnalog_v0p0p1_2.x65.X VDD.t646 VDD.t639 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X442 a_77723_n40777# VDD.t1506 a_77637_n40777# GND.t661 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X443 OUT0.t111 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND.t1192 GND.t1191 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X444 16to4_PriorityEncoder_v0p0p1_0.x3.EI 16to4_PriorityEncoder_v0p0p1_0.x5.EO VDD.t835 VDD.t834 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X445 frontAnalog_v0p0p1_8.RSfetsym_0.x1.Y frontAnalog_v0p0p1_8.x63.X VDD.t524 VDD.t519 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X446 GND.t1345 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t107 GND.t1344 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X447 GND.t1190 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t110 GND.t1189 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X448 GND.t1474 16to4_PriorityEncoder_v0p0p1_0.x36.A 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND.t1473 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X449 VDD.t1475 16to4_PriorityEncoder_v0p0p1_0.x22.A 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD.t1474 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X450 GND.t660 16to4_PriorityEncoder_v0p0p1_0.I13.t8 a_77723_n41087# GND.t659 sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X451 VIN.t10 w_55000_n19128# error sky130_fd_pr__cap_var_lvt w=2 l=0.18
X452 frontAnalog_v0p0p1_15.x63.A.t1 frontAnalog_v0p0p1_15.x65.A.t5 VDD.t238 VDD.t119 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X453 VDD.t250 frontAnalog_v0p0p1_0.x65.X frontAnalog_v0p0p1_0.RSfetsym_0.QN.t3 VDD.t243 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.25
X454 16to4_PriorityEncoder_v0p0p1_0.x3.x17.D a_77605_n51585# VDD.t463 VDD.t462 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.312 ps=1.68 w=1 l=0.15
X455 VDD.t985 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t43 VDD.t984 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X456 VDD.t692 16to4_PriorityEncoder_v0p0p1_0.x43.A 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD.t691 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X457 a_53630_n57996# frontAnalog_v0p0p1_10.IB.t8 GND.t444 GND.t186 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X458 frontAnalog_v0p0p1_14.x63.A.t0 CLK.t16 w_55000_n79150# VDD.t651 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X459 OUT1.t52 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD.t358 VDD.t357 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X460 OUT0.t48 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD.t1144 VDD.t1143 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X461 GND.t1188 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t109 GND.t1187 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X462 VDD.t454 16to4_PriorityEncoder_v0p0p1_0.x29.A 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD.t453 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X463 GND.t138 frontAnalog_v0p0p1_13.x65.X frontAnalog_v0p0p1_13.RSfetsym_0.x2.Y GND.t137 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X464 16to4_PriorityEncoder_v0p0p1_0.x3.x20.B frontAnalog_v0p0p1_9.Q.t7 GND.t34 GND.t33 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X465 frontAnalog_v0p0p1_4.x65.A.t0 CLK.t17 frontAnalog_v0p0p1_4.x63.A.t2 VDD.t652 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X466 a_59578_n73170# frontAnalog_v0p0p1_12.x65.X frontAnalog_v0p0p1_12.RSfetsym_0.QN.t2 GND.t99 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.315 ps=2.72 w=1 l=0.15
X467 OUT0.t47 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD.t1142 VDD.t1141 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X468 resistorDivider_v0p0p1_0.V16.t3 resistorDivider_v0p0p1_0.V15.t6 GND.t75 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X469 a_77605_n52567# 16to4_PriorityEncoder_v0p0p1_0.x3.x19.C VDD.t704 VDD.t114 sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.109 ps=1.36 w=0.42 l=0.15
X470 GND.t1343 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t106 GND.t1342 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X471 resistorDivider_v0p0p1_0.V14.t11 resistorDivider_v0p0p1_0.V13.t10 GND.t399 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X472 frontAnalog_v0p0p1_1.x63.A.t0 frontAnalog_v0p0p1_1.x65.A.t5 VDD.t1197 VDD.t746 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X473 VDD.t1140 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t46 VDD.t1139 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X474 OUT1.t112 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND.t363 GND.t362 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X475 OUT3.t105 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND.t1341 GND.t1340 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X476 frontAnalog_v0p0p1_8.x65.X a_57123_n45759# VDD.t814 VDD.t813 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X477 a_53630_n14796# frontAnalog_v0p0p1_10.IB.t9 GND.t445 GND.t186 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X478 frontAnalog_v0p0p1_7.x63.A.t0 CLK.t18 w_55000_n35950# VDD.t538 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X479 16to4_PriorityEncoder_v0p0p1_0.x36.Y 16to4_PriorityEncoder_v0p0p1_0.x36.A VDD.t1419 VDD.t1418 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X480 GND.t198 frontAnalog_v0p0p1_4.x65.A.t5 a_57123_n18759# GND.t197 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X481 frontAnalog_v0p0p1_10.RSfetsym_0.QN.t4 frontAnalog_v0p0p1_10.RSfetsym_0.x1.Y GND.t1552 GND.t936 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.25
X482 GND.t168 16to4_PriorityEncoder_v0p0p1_0.x3.x17.A a_78065_n49349# GND.t167 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X483 GND.t179 frontAnalog_v0p0p1_2.x63.A.t6 a_57123_n4079# GND.t21 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X484 frontAnalog_v0p0p1_0.RSfetsym_0.x2.Y frontAnalog_v0p0p1_0.x65.X VDD.t249 VDD.t245 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X485 OUT3.t49 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD.t1302 VDD.t1301 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X486 GND.t147 frontAnalog_v0p0p1_5.x65.X frontAnalog_v0p0p1_5.RSfetsym_0.x2.Y GND.t146 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X487 GND.t637 frontAnalog_v0p0p1_14.x63.X frontAnalog_v0p0p1_14.RSfetsym_0.x1.Y GND.t633 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X488 VDD.t356 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t51 VDD.t355 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X489 VDD.t1370 frontAnalog_v0p0p1_12.x63.A.t4 a_57123_n74279# VDD.t1369 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X490 16to4_PriorityEncoder_v0p0p1_0.I12.t4 frontAnalog_v0p0p1_4.RSfetsym_0.QN.t5 VDD.t714 VDD.t713 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.3
X491 GND.t1540 16to4_PriorityEncoder_v0p0p1_0.x22.A 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND.t1539 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X492 VDD.t60 frontAnalog_v0p0p1_4.x63.X frontAnalog_v0p0p1_4.RSfetsym_0.x1.Y VDD.t57 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X493 VDD.t1138 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t45 VDD.t1137 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X494 VDD.t653 CLK.t19 w_55000_n57550# GND.t103 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X495 VDD.t523 frontAnalog_v0p0p1_8.x63.X frontAnalog_v0p0p1_8.Q.t2 VDD.t517 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.25
X496 VDD.t1 frontAnalog_v0p0p1_11.x63.A.t4 frontAnalog_v0p0p1_11.x65.A.t0 VDD.t0 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X497 w_55000_n46128# CLK.t20 frontAnalog_v0p0p1_8.x65.A.t3 VDD.t88 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X498 16to4_PriorityEncoder_v0p0p1_0.x43.Y 16to4_PriorityEncoder_v0p0p1_0.x43.A GND.t772 GND.t771 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X499 16to4_PriorityEncoder_v0p0p1_0.I14.t1 frontAnalog_v0p0p1_0.RSfetsym_0.x2.Y GND.t881 GND.t568 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.25
X500 OUT1.t111 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND.t361 GND.t360 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X501 VDD.t1178 16to4_PriorityEncoder_v0p0p1_0.I15.t5 a_77639_n42341# VDD.t1177 sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X502 resistorDivider_v0p0p1_0.V13.t16 w_55000_n19750# error sky130_fd_pr__cap_var_lvt w=2 l=0.18
X503 a_16719_n13117.t14 a_16599_n13205.t9 a_16541_n13117.t3 GND.t218 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X504 frontAnalog_v0p0p1_13.x65.A.t2 frontAnalog_v0p0p1_13.x63.A.t5 a_55268_n68736# GND.t1239 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X505 OUT2.t42 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD.t981 VDD.t980 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X506 GND.t359 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t110 GND.t358 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X507 OUT3.t48 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD.t1300 VDD.t1299 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X508 frontAnalog_v0p0p1_3.RSfetsym_0.QN.t0 frontAnalog_v0p0p1_3.RSfetsym_0.x1.Y GND.t569 GND.t568 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.25
X509 VDD.t354 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t50 VDD.t353 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X510 GND.t814 frontAnalog_v0p0p1_7.x63.X frontAnalog_v0p0p1_7.RSfetsym_0.x1.Y GND.t810 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X511 VDD.t1366 frontAnalog_v0p0p1_2.x63.X 16to4_PriorityEncoder_v0p0p1_0.I15.t3 VDD.t1359 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.25
X512 VDD.t828 frontAnalog_v0p0p1_6.x63.A.t4 a_57123_n31079# VDD.t827 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X513 VDD.t1417 16to4_PriorityEncoder_v0p0p1_0.x36.A 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD.t1416 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X514 a_53630_n74196# resistorDivider_v0p0p1_0.V3.t16 w_55000_n73128# GND.t1078 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X515 resistorDivider_v0p0p1_0.V5.t1 resistorDivider_v0p0p1_0.V4.t3 GND.t26 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X516 VDD.t690 16to4_PriorityEncoder_v0p0p1_0.x43.A 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD.t689 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X517 resistorDivider_v0p0p1_0.V12.t10 resistorDivider_v0p0p1_0.V11.t10 GND.t506 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X518 GND.t1186 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t108 GND.t1185 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X519 VDD.t1473 16to4_PriorityEncoder_v0p0p1_0.x22.A 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD.t1472 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X520 OUT3.t104 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND.t1339 GND.t1338 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X521 VDD.t494 16to4_PriorityEncoder_v0p0p1_0.x3.x20.B a_77605_n52567# VDD.t114 sky130_fd_pr__pfet_01v8_hvt ad=0.312 pd=1.68 as=0.0588 ps=0.7 w=0.42 l=0.15
X522 a_55268_n52536# CLK.t21 GND.t573 GND.t572 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X523 16to4_PriorityEncoder_v0p0p1_0.x22.Y 16to4_PriorityEncoder_v0p0p1_0.x22.A GND.t1538 GND.t1537 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X524 frontAnalog_v0p0p1_5.x65.A.t0 frontAnalog_v0p0p1_5.x63.A.t5 a_55268_n25536# GND.t427 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X525 GND.t770 16to4_PriorityEncoder_v0p0p1_0.x43.A 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND.t769 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X526 GND.t1051 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t114 GND.t1050 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X527 VDD.t522 frontAnalog_v0p0p1_8.x63.X frontAnalog_v0p0p1_8.RSfetsym_0.x1.Y VDD.t519 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X528 OUT3.t47 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD.t1298 VDD.t1297 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X529 VDD.t352 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t49 VDD.t351 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X530 GND.t824 frontAnalog_v0p0p1_7.RSfetsym_0.QN.t6 a_59577_n35883# GND.t823 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X531 a_53630_n30996# resistorDivider_v0p0p1_0.V11.t16 w_55000_n29928# GND.t490 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X532 16to4_PriorityEncoder_v0p0p1_0.x36.Y 16to4_PriorityEncoder_v0p0p1_0.x36.A GND.t1472 GND.t1471 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X533 VDD.t1296 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t46 VDD.t1295 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X534 OUT1.t48 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD.t350 VDD.t349 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X535 VDD.t1136 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t44 VDD.t1135 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X536 a_55268_n9336# CLK.t22 GND.t575 GND.t574 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X537 GND.t944 frontAnalog_v0p0p1_11.x65.X frontAnalog_v0p0p1_11.RSfetsym_0.x2.Y GND.t943 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X538 VIN.t11 w_55000_n83928# error sky130_fd_pr__cap_var_lvt w=2 l=0.18
X539 frontAnalog_v0p0p1_5.RSfetsym_0.x1.Y frontAnalog_v0p0p1_5.x63.X VDD.t600 VDD.t593 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X540 VDD.t233 frontAnalog_v0p0p1_8.Q.t5 a_77639_n50381# VDD.t232 sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X541 16to4_PriorityEncoder_v0p0p1_0.x22.Y 16to4_PriorityEncoder_v0p0p1_0.x22.A VDD.t1471 VDD.t1470 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X542 VDD.t170 frontAnalog_v0p0p1_2.x63.A.t7 frontAnalog_v0p0p1_2.x65.A.t3 VDD.t106 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X543 VDD.t77 frontAnalog_v0p0p1_12.x65.X frontAnalog_v0p0p1_12.RSfetsym_0.QN.t1 VDD.t72 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.25
X544 16to4_PriorityEncoder_v0p0p1_0.x5.x21.B a_77605_n44527# GND.t170 GND.t169 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.196 ps=1.33 w=0.65 l=0.15
X545 OUT1.t109 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND.t357 GND.t356 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X546 16to4_PriorityEncoder_v0p0p1_0.x29.Y 16to4_PriorityEncoder_v0p0p1_0.x29.A VDD.t452 VDD.t451 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X547 frontAnalog_v0p0p1_2.x65.A.t1 CLK.t23 frontAnalog_v0p0p1_2.x63.A.t2 VDD.t528 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X548 resistorDivider_v0p0p1_0.V11.t15 resistorDivider_v0p0p1_0.V10.t14 GND.t102 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X549 VDD.t1294 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t45 VDD.t1293 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X550 OUT2.t41 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD.t979 VDD.t978 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X551 GND.t355 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t108 GND.t354 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X552 resistorDivider_v0p0p1_0.V16.t11 resistorDivider_v0p0p1_0.V15.t11 GND.t119 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X553 frontAnalog_v0p0p1_15.x65.A.t3 CLK.t24 frontAnalog_v0p0p1_15.x63.A.t3 VDD.t529 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X554 frontAnalog_v0p0p1_9.x63.X a_57123_n52679# VDD.t516 VDD.t515 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X555 OUT0.t107 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND.t1184 GND.t1183 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X556 w_55000_n68350# VIN.t12 a_53630_n68796# GND.t61 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X557 OUT2.t113 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND.t1049 GND.t1048 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X558 GND.t495 frontAnalog_v0p0p1_6.Q.t6 a_77605_n39305# GND.t24 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X559 GND.t643 frontAnalog_v0p0p1_12.x63.X frontAnalog_v0p0p1_12.RSfetsym_0.x1.Y GND.t640 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X560 VIN.t13 w_55000_n40728# error sky130_fd_pr__cap_var_lvt w=2 l=0.18
X561 VDD.t248 frontAnalog_v0p0p1_0.x65.X frontAnalog_v0p0p1_0.RSfetsym_0.x2.Y VDD.t245 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X562 VDD.t466 16to4_PriorityEncoder_v0p0p1_0.x5.x9.Y a_78313_n39305# VDD.t465 sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X563 VDD.t1193 16to4_PriorityEncoder_v0p0p1_0.I12.t5 a_77855_n40069# VDD.t1192 sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X564 resistorDivider_v0p0p1_0.V1.t13 VL.t6 GND.t59 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X565 GND.t247 frontAnalog_v0p0p1_15.x65.A.t6 a_57123_n83559# GND.t73 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X566 16to4_PriorityEncoder_v0p0p1_0.x3.x18.C frontAnalog_v0p0p1_12.Q.t6 GND.t234 GND.t233 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X567 a_77723_n49127# 16to4_PriorityEncoder_v0p0p1_0.x3.EI a_77637_n49127# GND.t865 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X568 VDD.t1292 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t44 VDD.t1291 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X569 GND.t469 16to4_PriorityEncoder_v0p0p1_0.x29.A 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND.t468 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X570 frontAnalog_v0p0p1_15.x63.A.t2 frontAnalog_v0p0p1_15.x65.A.t7 a_55268_n84936# GND.t248 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X571 16to4_PriorityEncoder_v0p0p1_0.x3.A2 a_78065_n49349# VDD.t387 VDD.t386 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.148 ps=1.34 w=1 l=0.15
X572 frontAnalog_v0p0p1_15.Q.t0 frontAnalog_v0p0p1_15.RSfetsym_0.QN.t5 VDD.t514 VDD.t381 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.3
X573 resistorDivider_v0p0p1_0.V9.t8 resistorDivider_v0p0p1_0.V8.t12 GND.t59 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X574 frontAnalog_v0p0p1_1.x65.A.t0 CLK.t25 frontAnalog_v0p0p1_1.x63.A.t2 VDD.t530 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X575 frontAnalog_v0p0p1_11.RSfetsym_0.x2.Y frontAnalog_v0p0p1_11.x65.X VDD.t891 VDD.t885 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X576 VDD.t861 frontAnalog_v0p0p1_15.x63.X frontAnalog_v0p0p1_15.RSfetsym_0.x1.Y VDD.t855 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X577 GND.t353 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t107 GND.t352 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X578 OUT3.t43 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD.t1290 VDD.t1289 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X579 frontAnalog_v0p0p1_2.RSfetsym_0.x1.Y frontAnalog_v0p0p1_2.x63.X VDD.t1365 VDD.t1361 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X580 w_55000_n25150# VIN.t14 a_53630_n25596# GND.t63 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X581 GND.t43 frontAnalog_v0p0p1_6.x63.X frontAnalog_v0p0p1_6.RSfetsym_0.x1.Y GND.t40 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X582 OUT0.t106 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND.t1182 GND.t1181 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X583 frontAnalog_v0p0p1_8.RSfetsym_0.x2.Y frontAnalog_v0p0p1_8.x65.X GND.t10 GND.t9 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X584 OUT0.t43 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD.t1134 VDD.t1133 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X585 a_78065_n49349# 16to4_PriorityEncoder_v0p0p1_0.x3.x22.A GND.t921 GND.t920 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X586 frontAnalog_v0p0p1_11.x63.X a_57123_n63479# GND.t948 GND.t675 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X587 a_53630_n3996# resistorDivider_v0p0p1_0.V16.t16 w_55000_n2928# GND.t1236 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X588 GND.t1180 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t105 GND.t1179 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X589 frontAnalog_v0p0p1_13.Q.t4 frontAnalog_v0p0p1_13.RSfetsym_0.x2.Y GND.t1404 GND.t1403 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.25
X590 resistorDivider_v0p0p1_0.V1.t17 w_55000_n84550# error sky130_fd_pr__cap_var_lvt w=2 l=0.18
X591 a_78065_n41309# 16to4_PriorityEncoder_v0p0p1_0.x5.x14.B GND.t930 GND.t929 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X592 OUT1.t47 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD.t348 VDD.t347 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X593 GND.t1249 frontAnalog_v0p0p1_1.x65.A.t6 a_57123_n40359# GND.t111 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X594 16to4_PriorityEncoder_v0p0p1_0.x3.x21.B a_77605_n52567# GND.t426 GND.t425 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.196 ps=1.33 w=0.65 l=0.15
X595 OUT3.t103 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND.t1337 GND.t1336 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X596 OUT2.t112 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND.t1047 GND.t1046 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X597 a_82988_n43855# 16to4_PriorityEncoder_v0p0p1_0.x3.A2 a_82906_n43855# VDD.t603 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X598 GND.t1045 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t111 GND.t1044 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X599 16to4_PriorityEncoder_v0p0p1_0.x28.A 16to4_PriorityEncoder_v0p0p1_0.x1.X VDD.t831 VDD.t830 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X600 frontAnalog_v0p0p1_1.x63.A.t1 frontAnalog_v0p0p1_1.x65.A.t7 a_55268_n41736# GND.t1243 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X601 GND.t351 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t106 GND.t350 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X602 frontAnalog_v0p0p1_1.Q.t4 frontAnalog_v0p0p1_1.RSfetsym_0.QN.t5 VDD.t1180 VDD.t870 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.3
X603 GND.t1335 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t102 GND.t1334 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X604 VDD.t168 frontAnalog_v0p0p1_1.x63.X frontAnalog_v0p0p1_1.RSfetsym_0.x1.Y VDD.t162 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X605 GND.t1043 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t110 GND.t1042 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X606 VDD.t789 frontAnalog_v0p0p1_14.x65.X frontAnalog_v0p0p1_14.RSfetsym_0.x2.Y VDD.t785 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X607 OUT3.t42 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD.t1288 VDD.t1287 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X608 16to4_PriorityEncoder_v0p0p1_0.x29.Y 16to4_PriorityEncoder_v0p0p1_0.x29.A GND.t467 GND.t466 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X609 frontAnalog_v0p0p1_10.RSfetsym_0.x1.Y frontAnalog_v0p0p1_10.x63.X GND.t184 GND.t180 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X610 a_59577_n46683# frontAnalog_v0p0p1_8.x63.X frontAnalog_v0p0p1_8.Q.t3 GND.t566 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X611 resistorDivider_v0p0p1_0.V14.t5 resistorDivider_v0p0p1_0.V13.t2 GND.t102 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X612 a_59578_n56970# frontAnalog_v0p0p1_10.x65.X frontAnalog_v0p0p1_10.RSfetsym_0.QN.t1 GND.t1442 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.315 ps=2.72 w=1 l=0.15
X613 resistorDivider_v0p0p1_0.V5.t8 resistorDivider_v0p0p1_0.V4.t13 GND.t60 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X614 GND.t1447 frontAnalog_v0p0p1_12.Q.t7 a_77605_n47345# GND.t65 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X615 16to4_PriorityEncoder_v0p0p1_0.x3.x9.Y 16to4_PriorityEncoder_v0p0p1_0.x3.EI VDD.t805 VDD.t804 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X616 OUT0.t42 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD.t1132 VDD.t1131 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X617 VDD.t202 16to4_PriorityEncoder_v0p0p1_0.x3.x9.Y a_78313_n47345# VDD.t201 sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X618 VDD.t1286 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t41 VDD.t1285 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X619 16to4_PriorityEncoder_v0p0p1_0.I11.t4 frontAnalog_v0p0p1_5.RSfetsym_0.x2.Y GND.t1509 GND.t1488 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.25
X620 resistorDivider_v0p0p1_0.V9.t17 w_55000_n41350# error sky130_fd_pr__cap_var_lvt w=2 l=0.18
X621 GND.t1083 frontAnalog_v0p0p1_14.RSfetsym_0.QN.t6 a_59577_n79083# GND.t1082 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X622 GND.t253 16to4_PriorityEncoder_v0p0p1_0.x5.x17.C a_78349_n43045# GND.t252 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X623 VDD.t1130 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t41 VDD.t1129 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X624 16to4_PriorityEncoder_v0p0p1_0.x3.x21.B a_77605_n52567# VDD.t405 VDD.t404 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.312 ps=1.68 w=1 l=0.15
X625 GND.t1333 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t101 GND.t1332 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X626 VDD.t1337 frontAnalog_v0p0p1_7.x65.X frontAnalog_v0p0p1_7.RSfetsym_0.x2.Y VDD.t1333 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X627 frontAnalog_v0p0p1_13.RSfetsym_0.x1.Y frontAnalog_v0p0p1_13.x63.X VDD.t502 VDD.t495 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X628 a_77775_n43295# 16to4_PriorityEncoder_v0p0p1_0.x5.x19.C a_77687_n43295# GND.t156 sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
X629 OUT2.t109 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND.t1041 GND.t1040 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X630 GND.t1039 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t108 GND.t1038 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X631 frontAnalog_v0p0p1_3.RSfetsym_0.x1.Y frontAnalog_v0p0p1_3.x63.X GND.t241 GND.t237 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X632 OUT1.t105 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND.t349 GND.t348 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X633 VDD.t688 16to4_PriorityEncoder_v0p0p1_0.x43.A 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD.t687 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X634 a_59578_n13770# frontAnalog_v0p0p1_3.x65.X frontAnalog_v0p0p1_3.RSfetsym_0.QN.t1 GND.t698 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.315 ps=2.72 w=1 l=0.15
X635 a_53630_n52596# frontAnalog_v0p0p1_10.IB.t10 GND.t652 GND.t186 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X636 frontAnalog_v0p0p1_1.Q.t1 frontAnalog_v0p0p1_1.x63.X VDD.t167 VDD.t164 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.25
X637 16to4_PriorityEncoder_v0p0p1_0.x1.X a_82906_n47995# GND.t784 GND.t783 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1 ps=0.985 w=0.65 l=0.15
X638 16to4_PriorityEncoder_v0p0p1_0.x5.x17.A a_77637_n42017# VDD.t877 VDD.t876 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.167 ps=1.39 w=1 l=0.15
X639 VFS.t5 resistorDivider_v0p0p1_0.V16.t9 GND.t889 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X640 VDD.t187 frontAnalog_v0p0p1_8.x63.A.t4 frontAnalog_v0p0p1_8.x65.A.t1 VDD.t186 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X641 GND.t817 frontAnalog_v0p0p1_8.Q.t6 a_59578_n46170# GND.t816 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X642 16to4_PriorityEncoder_v0p0p1_0.x3.EI 16to4_PriorityEncoder_v0p0p1_0.x5.EO GND.t887 GND.t886 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X643 OUT0.t104 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND.t1178 GND.t1177 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X644 frontAnalog_v0p0p1_2.RSfetsym_0.QN.t0 frontAnalog_v0p0p1_2.RSfetsym_0.x1.Y GND.t626 GND.t625 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.25
X645 resistorDivider_v0p0p1_0.V4.t12 resistorDivider_v0p0p1_0.V3.t8 GND.t75 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X646 VDD.t645 frontAnalog_v0p0p1_2.x65.X frontAnalog_v0p0p1_2.RSfetsym_0.x2.Y VDD.t639 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X647 GND.t22 frontAnalog_v0p0p1_2.x65.A.t5 a_57123_n2559# GND.t21 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X648 frontAnalog_v0p0p1_15.RSfetsym_0.QN.t0 frontAnalog_v0p0p1_15.Q.t6 VDD.t382 VDD.t381 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.3
X649 resistorDivider_v0p0p1_0.V8.t0 resistorDivider_v0p0p1_0.V7.t0 GND.t26 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X650 GND.t1331 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t100 GND.t1330 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X651 frontAnalog_v0p0p1_11.x65.X a_57123_n61959# GND.t676 GND.t675 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X652 GND.t1176 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t103 GND.t1175 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X653 OUT1.t104 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND.t347 GND.t346 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X654 a_77605_n43295# 16to4_PriorityEncoder_v0p0p1_0.x5.x16.C VDD.t505 VDD.t504 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X655 VDD.t819 frontAnalog_v0p0p1_3.x63.A.t5 a_57123_n14879# VDD.t818 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X656 OUT3.t99 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND.t1329 GND.t1328 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X657 VDD.t1284 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t40 VDD.t1283 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X658 GND.t1250 16to4_PriorityEncoder_v0p0p1_0.I12.t6 a_77605_n40069# GND.t243 sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X659 frontAnalog_v0p0p1_4.RSfetsym_0.QN.t4 16to4_PriorityEncoder_v0p0p1_0.I12.t7 VDD.t1198 VDD.t713 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.3
X660 VDD.t1348 frontAnalog_v0p0p1_12.x65.A.t4 a_57123_n72759# VDD.t1347 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X661 GND.t1240 frontAnalog_v0p0p1_13.x63.A.t6 a_57123_n68879# GND.t56 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X662 VDD.t977 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t40 VDD.t976 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X663 16to4_PriorityEncoder_v0p0p1_0.x43.Y 16to4_PriorityEncoder_v0p0p1_0.x43.A VDD.t686 VDD.t685 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X664 VDD.t346 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t46 VDD.t345 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X665 VDD.t890 frontAnalog_v0p0p1_11.x65.X frontAnalog_v0p0p1_11.RSfetsym_0.x2.Y VDD.t885 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X666 VDD.t1364 frontAnalog_v0p0p1_2.x63.X frontAnalog_v0p0p1_2.RSfetsym_0.x1.Y VDD.t1361 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X667 GND.t1536 16to4_PriorityEncoder_v0p0p1_0.x22.A 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND.t1535 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X668 frontAnalog_v0p0p1_1.RSfetsym_0.QN.t4 frontAnalog_v0p0p1_1.Q.t5 VDD.t871 VDD.t870 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.3
X669 OUT0.t40 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD.t1128 VDD.t1127 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X670 a_77605_n39305# 16to4_PriorityEncoder_v0p0p1_0.I11.t5 GND.t1087 GND.t24 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X671 GND.t1174 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t102 GND.t1173 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X672 frontAnalog_v0p0p1_4.RSfetsym_0.x2.Y frontAnalog_v0p0p1_4.x65.X VDD.t849 VDD.t844 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X673 VDD.t1126 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t39 VDD.t1125 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X674 OUT1.t103 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND.t345 GND.t344 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X675 frontAnalog_v0p0p1_4.RSfetsym_0.x1.Y frontAnalog_v0p0p1_4.x63.X GND.t81 GND.t76 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X676 OUT3.t98 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND.t1327 GND.t1326 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X677 a_77855_n40069# 16to4_PriorityEncoder_v0p0p1_0.I13.t9 a_77783_n40069# VDD.t414 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X678 resistorDivider_v0p0p1_0.V2.t8 resistorDivider_v0p0p1_0.V1.t12 GND.t84 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X679 OUT2.t107 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND.t1037 GND.t1036 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X680 VDD.t1282 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t39 VDD.t1281 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X681 a_16719_n13117.t13 a_16599_n13205.t10 a_16541_n13117.t2 GND.t1561 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X682 GND.t343 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t102 GND.t342 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X683 GND.t428 frontAnalog_v0p0p1_5.x63.A.t6 a_57123_n25679# GND.t45 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X684 frontAnalog_v0p0p1_8.RSfetsym_0.QN.t3 frontAnalog_v0p0p1_8.x65.X VDD.t10 VDD.t6 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.25
X685 frontAnalog_v0p0p1_1.RSfetsym_0.x1.Y frontAnalog_v0p0p1_1.x63.X GND.t177 GND.t173 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X686 OUT3.t38 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD.t1280 VDD.t1279 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X687 GND.t1092 16to4_PriorityEncoder_v0p0p1_0.I14.t5 a_77723_n42017# GND.t1091 sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X688 frontAnalog_v0p0p1_2.x63.A.t0 frontAnalog_v0p0p1_2.x65.A.t6 a_55268_n3936# GND.t23 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X689 GND.t1172 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t101 GND.t1171 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X690 VDD.t1469 16to4_PriorityEncoder_v0p0p1_0.x22.A 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD.t1468 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X691 VDD.t401 frontAnalog_v0p0p1_1.Q.t6 a_77855_n39305# VDD.t400 sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X692 OUT3.t97 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND.t1325 GND.t1324 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X693 16to4_PriorityEncoder_v0p0p1_0.x22.Y 16to4_PriorityEncoder_v0p0p1_0.x22.A GND.t1534 GND.t1533 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X694 VDD.t975 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t39 VDD.t974 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X695 VDD.t1124 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t38 VDD.t1123 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X696 a_77605_n51335# 16to4_PriorityEncoder_v0p0p1_0.x3.x16.C VDD.t151 VDD.t150 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X697 frontAnalog_v0p0p1_13.x63.A.t3 frontAnalog_v0p0p1_13.x65.A.t5 VDD.t884 VDD.t122 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X698 a_77881_n52819# 16to4_PriorityEncoder_v0p0p1_0.x3.x19.C a_77775_n52819# GND.t532 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X699 frontAnalog_v0p0p1_2.RSfetsym_0.QN.t3 frontAnalog_v0p0p1_2.x65.X VDD.t644 VDD.t642 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.25
X700 GND.t768 16to4_PriorityEncoder_v0p0p1_0.x43.A 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND.t767 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X701 frontAnalog_v0p0p1_9.RSfetsym_0.x1.Y frontAnalog_v0p0p1_9.x63.X VDD.t196 VDD.t191 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X702 GND.t341 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t101 GND.t340 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X703 GND.t1257 frontAnalog_v0p0p1_11.Q.t7 a_77605_n48109# GND.t818 sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X704 OUT2.t38 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD.t973 VDD.t972 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X705 OUT3.t37 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD.t1278 VDD.t1277 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X706 VDD.t344 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t45 VDD.t343 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X707 OUT1.t44 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD.t342 VDD.t341 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X708 VDD.t625 frontAnalog_v0p0p1_3.x65.X frontAnalog_v0p0p1_3.RSfetsym_0.QN.t2 VDD.t624 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.25
X709 VDD.t1122 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t37 VDD.t1121 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X710 frontAnalog_v0p0p1_15.Q.t4 frontAnalog_v0p0p1_15.x63.X VDD.t860 VDD.t857 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.25
X711 a_77605_n47345# frontAnalog_v0p0p1_13.Q.t5 GND.t1437 GND.t65 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X712 OUT3.t96 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND.t1323 GND.t1322 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X713 frontAnalog_v0p0p1_5.x63.A.t3 frontAnalog_v0p0p1_5.x65.A.t5 VDD.t1026 VDD.t488 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X714 OUT0.t100 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND.t1170 GND.t1169 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X715 a_59577_n3483# frontAnalog_v0p0p1_2.x63.X 16to4_PriorityEncoder_v0p0p1_0.I15.t1 GND.t1410 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X716 resistorDivider_v0p0p1_0.V12.t1 resistorDivider_v0p0p1_0.V11.t0 GND.t196 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X717 16to4_PriorityEncoder_v0p0p1_0.x2.X a_82906_n51645# GND.t236 GND.t235 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1 ps=0.985 w=0.65 l=0.15
X718 16to4_PriorityEncoder_v0p0p1_0.x22.Y 16to4_PriorityEncoder_v0p0p1_0.x22.A VDD.t1467 VDD.t1466 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X719 w_55000_n2928# CLK.t26 frontAnalog_v0p0p1_2.x65.A.t0 VDD.t28 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X720 frontAnalog_v0p0p1_6.x65.X a_57123_n29559# VDD.t841 VDD.t840 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X721 GND.t1321 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t95 GND.t1320 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X722 frontAnalog_v0p0p1_4.x63.A.t3 CLK.t27 w_55000_n19750# VDD.t531 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X723 VDD.t971 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t37 VDD.t970 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X724 OUT2.t36 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD.t969 VDD.t968 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X725 16to4_PriorityEncoder_v0p0p1_0.x29.Y 16to4_PriorityEncoder_v0p0p1_0.x29.A GND.t465 GND.t464 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X726 GND.t36 frontAnalog_v0p0p1_9.Q.t8 a_77723_n50057# GND.t35 sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X727 frontAnalog_v0p0p1_9.x65.X a_57123_n51159# VDD.t391 VDD.t390 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X728 resistorDivider_v0p0p1_0.V4.t4 resistorDivider_v0p0p1_0.V3.t2 GND.t119 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X729 frontAnalog_v0p0p1_8.x63.X a_57123_n47279# GND.t1553 GND.t870 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X730 VDD.t241 frontAnalog_v0p0p1_10.x63.A.t5 a_57123_n58079# VDD.t240 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X731 OUT1.t43 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD.t340 VDD.t339 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X732 resistorDivider_v0p0p1_0.V10.t12 resistorDivider_v0p0p1_0.V9.t12 GND.t84 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X733 VDD.t80 CLK.t28 w_55000_n62328# GND.t103 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X734 OUT0.t99 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND.t1168 GND.t1167 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X735 frontAnalog_v0p0p1_11.RSfetsym_0.QN.t0 frontAnalog_v0p0p1_11.RSfetsym_0.x1.Y GND.t632 GND.t621 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.25
X736 16to4_PriorityEncoder_v0p0p1_0.x5.x16.C 16to4_PriorityEncoder_v0p0p1_0.I13.t10 GND.t436 GND.t435 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X737 a_78349_n51085# 16to4_PriorityEncoder_v0p0p1_0.x3.x17.D GND.t1395 GND.t165 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X738 VDD.t384 frontAnalog_v0p0p1_15.Q.t7 a_77855_n47345# VDD.t383 sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X739 resistorDivider_v0p0p1_0.V3.t12 resistorDivider_v0p0p1_0.V2.t12 GND.t506 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X740 a_77687_n43545# 16to4_PriorityEncoder_v0p0p1_0.I11.t6 a_77605_n43545# GND.t153 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.109 ps=1.36 w=0.42 l=0.15
X741 resistorDivider_v0p0p1_0.V13.t3 resistorDivider_v0p0p1_0.V12.t2 GND.t84 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X742 a_53630_n9396# frontAnalog_v0p0p1_10.IB.t11 GND.t653 GND.t503 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X743 frontAnalog_v0p0p1_12.RSfetsym_0.x2.Y frontAnalog_v0p0p1_12.x65.X GND.t98 GND.t97 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X744 VDD.t207 16to4_PriorityEncoder_v0p0p1_0.I11.t7 a_77605_n44779# VDD.t206 sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X745 resistorDivider_v0p0p1_0.V8.t4 resistorDivider_v0p0p1_0.V7.t5 GND.t60 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X746 OUT2.t35 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD.t967 VDD.t966 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X747 VDD.t599 frontAnalog_v0p0p1_5.x63.X frontAnalog_v0p0p1_5.RSfetsym_0.x1.Y VDD.t593 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X748 resistorDivider_v0p0p1_0.V2.t11 resistorDivider_v0p0p1_0.V1.t14 GND.t399 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X749 OUT0.t36 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD.t1120 VDD.t1119 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X750 VDD.t1438 16to4_PriorityEncoder_v0p0p1_0.x5.x17.A a_78599_n43045# VDD.t1437 sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X751 VDD.t195 frontAnalog_v0p0p1_9.x63.X frontAnalog_v0p0p1_9.Q.t0 VDD.t194 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.25
X752 VDD.t81 CLK.t29 w_55000_n62950# GND.t104 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X753 GND.t1319 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t94 GND.t1318 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X754 16to4_PriorityEncoder_v0p0p1_0.x2.X a_82906_n51645# VDD.t219 VDD.t218 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.146 ps=1.34 w=1 l=0.15
X755 w_55000_n51528# CLK.t30 frontAnalog_v0p0p1_9.x65.A.t3 VDD.t82 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X756 OUT1.t100 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND.t339 GND.t338 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X757 VDD.t1415 16to4_PriorityEncoder_v0p0p1_0.x36.A 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD.t1414 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X758 GND.t80 frontAnalog_v0p0p1_4.x63.X frontAnalog_v0p0p1_4.RSfetsym_0.x1.Y GND.t76 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X759 16to4_PriorityEncoder_v0p0p1_0.x3.x19.C frontAnalog_v0p0p1_11.Q.t8 GND.t447 GND.t446 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X760 frontAnalog_v0p0p1_12.x65.A.t2 frontAnalog_v0p0p1_12.x63.A.t5 a_55268_n74136# GND.t1415 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X761 a_53630_n57996# resistorDivider_v0p0p1_0.V6.t16 w_55000_n56928# GND.t737 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X762 GND.t463 16to4_PriorityEncoder_v0p0p1_0.x29.A 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND.t462 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X763 VDD.t450 16to4_PriorityEncoder_v0p0p1_0.x29.A 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD.t449 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X764 OUT0.t98 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND.t1166 GND.t1165 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X765 frontAnalog_v0p0p1_15.RSfetsym_0.x2.Y frontAnalog_v0p0p1_15.x65.X VDD.t1377 VDD.t1371 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X766 OUT0.t35 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD.t1118 VDD.t1117 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X767 GND.t176 frontAnalog_v0p0p1_1.x63.X frontAnalog_v0p0p1_1.RSfetsym_0.x1.Y GND.t173 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X768 frontAnalog_v0p0p1_0.x63.X a_57123_n9479# VDD.t816 VDD.t815 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X769 frontAnalog_v0p0p1_6.RSfetsym_0.x2.Y frontAnalog_v0p0p1_6.x65.X GND.t519 GND.t518 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X770 a_55268_n36336# CLK.t31 GND.t106 GND.t105 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X771 frontAnalog_v0p0p1_15.RSfetsym_0.x1.Y frontAnalog_v0p0p1_15.x63.X GND.t912 GND.t908 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X772 GND.t766 16to4_PriorityEncoder_v0p0p1_0.x43.A 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND.t765 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X773 GND.t1164 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t97 GND.t1163 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X774 VDD.t83 CLK.t32 w_55000_n19750# GND.t107 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X775 VFS.t6 resistorDivider_v0p0p1_0.V16.t10 GND.t552 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X776 resistorDivider_v0p0p1_0.V6.t8 resistorDivider_v0p0p1_0.V5.t10 GND.t889 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X777 OUT1.t42 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD.t338 VDD.t337 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X778 OUT3.t93 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND.t1317 GND.t1316 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X779 VDD.t961 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t34 VDD.t960 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X780 GND.t1227 frontAnalog_v0p0p1_0.RSfetsym_0.QN.t5 a_59577_n8883# GND.t1226 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X781 OUT1.t41 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD.t336 VDD.t335 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X782 a_53630_n14796# resistorDivider_v0p0p1_0.V14.t16 w_55000_n13728# GND.t546 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X783 GND.t731 frontAnalog_v0p0p1_4.RSfetsym_0.QN.t6 a_59577_n19683# GND.t730 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X784 GND.t497 frontAnalog_v0p0p1_6.Q.t7 a_59578_n29970# GND.t496 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X785 16to4_PriorityEncoder_v0p0p1_0.x36.Y 16to4_PriorityEncoder_v0p0p1_0.x36.A VDD.t1413 VDD.t1412 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X786 OUT3.t36 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD.t1276 VDD.t1275 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X787 VDD.t193 frontAnalog_v0p0p1_9.x63.X frontAnalog_v0p0p1_9.RSfetsym_0.x1.Y VDD.t191 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X788 VDD.t334 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t40 VDD.t333 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X789 frontAnalog_v0p0p1_1.RSfetsym_0.x2.Y frontAnalog_v0p0p1_1.x65.X VDD.t617 VDD.t610 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X790 frontAnalog_v0p0p1_14.x63.X a_57123_n79679# VDD.t708 VDD.t707 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X791 a_77687_n51585# frontAnalog_v0p0p1_13.Q.t6 a_77605_n51585# GND.t158 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.109 ps=1.36 w=0.42 l=0.15
X792 OUT0.t34 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD.t1116 VDD.t1115 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X793 a_78735_n39527# 16to4_PriorityEncoder_v0p0p1_0.x5.EO a_78649_n39527# GND.t885 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X794 GND.t8 frontAnalog_v0p0p1_8.x65.X frontAnalog_v0p0p1_8.RSfetsym_0.x2.Y GND.t7 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X795 16to4_PriorityEncoder_v0p0p1_0.x5.x14.B a_77637_n41087# VDD.t101 VDD.t100 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.167 ps=1.39 w=1 l=0.15
X796 VDD.t1274 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t35 VDD.t1273 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X797 VIN.t15 w_55000_n67728# error sky130_fd_pr__cap_var_lvt w=2 l=0.18
X798 GND.t665 VDD.t1507 a_77881_n43545# GND.t153 sky130_fd_pr__nfet_01v8 ad=0.196 pd=1.33 as=0.0693 ps=0.75 w=0.42 l=0.15
X799 GND.t1162 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t96 GND.t1161 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X800 VDD.t1030 frontAnalog_v0p0p1_13.Q.t7 a_77605_n52819# VDD.t1029 sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X801 a_77605_n44779# VDD.t772 VDD.t773 VDD.t415 sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.109 ps=1.36 w=0.42 l=0.15
X802 VDD.t158 16to4_PriorityEncoder_v0p0p1_0.x3.x17.A a_78599_n51085# VDD.t157 sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X803 GND.t53 16to4_PriorityEncoder_v0p0p1_0.x35.A 16to4_PriorityEncoder_v0p0p1_0.x36.A GND.t52 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X804 VDD.t1114 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t33 VDD.t1113 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X805 VDD.t1387 frontAnalog_v0p0p1_10.x65.X frontAnalog_v0p0p1_10.RSfetsym_0.QN.t2 VDD.t1386 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.25
X806 OUT3.t92 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND.t1315 GND.t1314 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X807 a_77855_n39305# frontAnalog_v0p0p1_7.Q.t7 a_77783_n39305# VDD.t32 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X808 a_78097_n45737# VDD.t769 VDD.t771 VDD.t770 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X809 VDD.t658 16to4_PriorityEncoder_v0p0p1_0.x42.A 16to4_PriorityEncoder_v0p0p1_0.x43.A VDD.t657 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X810 VDD.t332 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t39 VDD.t331 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X811 GND.t1313 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t91 GND.t1312 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X812 resistorDivider_v0p0p1_0.V10.t11 resistorDivider_v0p0p1_0.V9.t10 GND.t399 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X813 OUT2.t106 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND.t1035 GND.t1034 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X814 frontAnalog_v0p0p1_13.x65.A.t1 CLK.t33 frontAnalog_v0p0p1_13.x63.A.t1 VDD.t84 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X815 OUT1.t99 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND.t337 GND.t336 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X816 frontAnalog_v0p0p1_7.x63.X a_57123_n36479# VDD.t619 VDD.t618 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X817 GND.t183 frontAnalog_v0p0p1_10.x63.X frontAnalog_v0p0p1_10.RSfetsym_0.x1.Y GND.t180 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X818 VIN.t16 w_55000_n24528# error sky130_fd_pr__cap_var_lvt w=2 l=0.18
X819 resistorDivider_v0p0p1_0.V13.t12 resistorDivider_v0p0p1_0.V12.t13 GND.t399 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X820 a_53630_n3996# frontAnalog_v0p0p1_10.IB.t12 GND.t654 GND.t503 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X821 16to4_PriorityEncoder_v0p0p1_0.x22.Y 16to4_PriorityEncoder_v0p0p1_0.x22.A GND.t1532 GND.t1531 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X822 a_53630_n63396# frontAnalog_v0p0p1_10.IB.t13 GND.t655 GND.t186 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X823 VDD.t1112 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t32 VDD.t1111 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X824 frontAnalog_v0p0p1_15.x63.A.t0 CLK.t34 w_55000_n84550# VDD.t85 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X825 GND.t57 frontAnalog_v0p0p1_13.x65.A.t6 a_57123_n67359# GND.t56 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X826 OUT2.t33 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD.t965 VDD.t964 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X827 frontAnalog_v0p0p1_13.x63.A.t0 frontAnalog_v0p0p1_13.x65.A.t7 a_55268_n68736# GND.t58 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X828 GND.t96 frontAnalog_v0p0p1_12.x65.X frontAnalog_v0p0p1_12.RSfetsym_0.x2.Y GND.t95 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X829 16to4_PriorityEncoder_v0p0p1_0.x36.A 16to4_PriorityEncoder_v0p0p1_0.x35.A VDD.t54 VDD.t53 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X830 VDD.t448 16to4_PriorityEncoder_v0p0p1_0.x29.A 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD.t447 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X831 frontAnalog_v0p0p1_5.x65.A.t2 CLK.t35 frontAnalog_v0p0p1_5.x63.A.t1 VDD.t12 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X832 frontAnalog_v0p0p1_13.Q.t0 frontAnalog_v0p0p1_13.RSfetsym_0.QN.t5 VDD.t1449 VDD.t1031 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.3
X833 VDD.t501 frontAnalog_v0p0p1_13.x63.X frontAnalog_v0p0p1_13.RSfetsym_0.x1.Y VDD.t495 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X834 frontAnalog_v0p0p1_8.RSfetsym_0.x2.Y frontAnalog_v0p0p1_8.x65.X VDD.t9 VDD.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X835 16to4_PriorityEncoder_v0p0p1_0.x5.x17.C a_77605_n43295# GND.t409 GND.t408 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.196 ps=1.33 w=0.65 l=0.15
X836 GND.t240 frontAnalog_v0p0p1_3.x63.X frontAnalog_v0p0p1_3.RSfetsym_0.x1.Y GND.t237 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X837 GND.t1251 16to4_PriorityEncoder_v0p0p1_0.I12.t8 a_77723_n40777# GND.t659 sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X838 a_78735_n47567# 16to4_PriorityEncoder_v0p0p1_0.x3.EO a_78649_n47567# GND.t1084 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X839 GND.t866 16to4_PriorityEncoder_v0p0p1_0.x3.EI a_77881_n51585# GND.t158 sky130_fd_pr__nfet_01v8 ad=0.196 pd=1.33 as=0.0693 ps=0.75 w=0.42 l=0.15
X840 a_77605_n52819# 16to4_PriorityEncoder_v0p0p1_0.x3.EI VDD.t803 VDD.t548 sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.109 ps=1.36 w=0.42 l=0.15
X841 resistorDivider_v0p0p1_0.V5.t7 resistorDivider_v0p0p1_0.V4.t11 GND.t59 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X842 16to4_PriorityEncoder_v0p0p1_0.x43.Y 16to4_PriorityEncoder_v0p0p1_0.x43.A VDD.t684 VDD.t683 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X843 resistorDivider_v0p0p1_0.V4.t17 w_55000_n68350# error sky130_fd_pr__cap_var_lvt w=2 l=0.18
X844 OUT0.t95 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND.t1160 GND.t1159 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X845 VDD.t854 16to4_PriorityEncoder_v0p0p1_0.x5.x20.B a_77605_n44779# VDD.t853 sky130_fd_pr__pfet_01v8_hvt ad=0.312 pd=1.68 as=0.0588 ps=0.7 w=0.42 l=0.15
X846 GND.t46 frontAnalog_v0p0p1_5.x65.A.t6 a_57123_n24159# GND.t45 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X847 frontAnalog_v0p0p1_9.RSfetsym_0.x2.Y frontAnalog_v0p0p1_9.x65.X GND.t718 GND.t717 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X848 16to4_PriorityEncoder_v0p0p1_0.x22.Y 16to4_PriorityEncoder_v0p0p1_0.x22.A VDD.t1465 VDD.t1464 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X849 frontAnalog_v0p0p1_5.x63.A.t0 frontAnalog_v0p0p1_5.x65.A.t7 a_55268_n25536# GND.t47 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X850 a_78097_n53777# 16to4_PriorityEncoder_v0p0p1_0.x3.EI VDD.t802 VDD.t801 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X851 GND.t1530 16to4_PriorityEncoder_v0p0p1_0.x22.A 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND.t1529 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X852 a_77855_n47345# frontAnalog_v0p0p1_14.Q.t8 a_77783_n47345# VDD.t535 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X853 GND.t517 frontAnalog_v0p0p1_6.x65.X frontAnalog_v0p0p1_6.RSfetsym_0.x2.Y GND.t516 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X854 GND.t911 frontAnalog_v0p0p1_15.x63.X frontAnalog_v0p0p1_15.RSfetsym_0.x1.Y GND.t908 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X855 16to4_PriorityEncoder_v0p0p1_0.I11.t3 frontAnalog_v0p0p1_5.RSfetsym_0.QN.t5 VDD.t543 VDD.t542 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.3
X856 VDD.t330 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t38 VDD.t329 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X857 a_78599_n43045# 16to4_PriorityEncoder_v0p0p1_0.x5.x22.A a_78527_n43045# VDD.t555 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X858 OUT2.t105 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND.t1033 GND.t1032 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X859 VDD.t1272 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t34 VDD.t1271 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X860 16to4_PriorityEncoder_v0p0p1_0.x29.Y 16to4_PriorityEncoder_v0p0p1_0.x29.A VDD.t446 VDD.t445 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X861 16to4_PriorityEncoder_v0p0p1_0.x5.x17.C a_77605_n43295# VDD.t393 VDD.t392 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.312 ps=1.68 w=1 l=0.15
X862 frontAnalog_v0p0p1_13.Q.t3 frontAnalog_v0p0p1_13.x63.X VDD.t500 VDD.t497 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.25
X863 a_53630_n79596# frontAnalog_v0p0p1_10.IB.t14 GND.t656 GND.t186 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X864 resistorDivider_v0p0p1_0.V15.t0 resistorDivider_v0p0p1_0.V14.t1 GND.t75 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X865 OUT3.t33 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD.t1270 VDD.t1269 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X866 resistorDivider_v0p0p1_0.V12.t17 w_55000_n25150# error sky130_fd_pr__cap_var_lvt w=2 l=0.18
X867 frontAnalog_v0p0p1_11.RSfetsym_0.x1.Y frontAnalog_v0p0p1_11.x63.X GND.t117 GND.t113 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X868 OUT0.t31 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD.t1110 VDD.t1109 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X869 frontAnalog_v0p0p1_6.Q.t4 frontAnalog_v0p0p1_6.RSfetsym_0.x2.Y GND.t904 GND.t536 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.25
X870 GND.t735 frontAnalog_v0p0p1_15.RSfetsym_0.QN.t6 a_59577_n84483# GND.t734 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X871 VDD.t1463 16to4_PriorityEncoder_v0p0p1_0.x22.A 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD.t1462 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X872 VDD.t1411 16to4_PriorityEncoder_v0p0p1_0.x36.A 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD.t1410 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X873 VDD.t848 frontAnalog_v0p0p1_4.x65.X frontAnalog_v0p0p1_4.RSfetsym_0.x2.Y VDD.t844 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X874 16to4_PriorityEncoder_v0p0p1_0.x3.x14.A a_77637_n48817# GND.t549 GND.t548 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.112 ps=1.04 w=0.65 l=0.15
X875 OUT2.t104 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND.t1031 GND.t1030 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X876 VDD.t34 frontAnalog_v0p0p1_7.Q.t8 a_77605_n44527# VDD.t33 sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X877 16to4_PriorityEncoder_v0p0p1_0.I11.t2 frontAnalog_v0p0p1_5.x63.X VDD.t598 VDD.t595 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.25
X878 a_53630_n36396# frontAnalog_v0p0p1_10.IB.t15 GND.t931 GND.t186 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X879 16to4_PriorityEncoder_v0p0p1_0.x3.x4.C a_77605_n48109# GND.t704 GND.t703 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.102 ps=0.99 w=0.65 l=0.15
X880 frontAnalog_v0p0p1_12.RSfetsym_0.x1.Y frontAnalog_v0p0p1_12.x63.X VDD.t592 VDD.t585 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X881 VDD.t829 frontAnalog_v0p0p1_6.x63.A.t5 frontAnalog_v0p0p1_6.x65.A.t2 VDD.t412 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X882 OUT3.t32 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD.t1268 VDD.t1267 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X883 a_16541_n13117.t20 GND.t800 GND.t799 sky130_fd_pr__res_xhigh_po_5p73 l=85.8
X884 resistorDivider_v0p0p1_0.V2.t7 resistorDivider_v0p0p1_0.V1.t11 GND.t102 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X885 VDD.t493 16to4_PriorityEncoder_v0p0p1_0.x3.x20.B a_77605_n52819# VDD.t492 sky130_fd_pr__pfet_01v8_hvt ad=0.312 pd=1.68 as=0.0588 ps=0.7 w=0.42 l=0.15
X886 GND.t592 16to4_PriorityEncoder_v0p0p1_0.x5.x22.A a_78525_n45515# GND.t591 sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X887 frontAnalog_v0p0p1_13.RSfetsym_0.QN.t4 frontAnalog_v0p0p1_13.Q.t8 VDD.t1032 VDD.t1031 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.3
X888 GND.t38 frontAnalog_v0p0p1_9.Q.t9 a_59578_n51570# GND.t37 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X889 frontAnalog_v0p0p1_8.x65.X a_57123_n45759# GND.t871 GND.t870 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X890 GND.t1229 frontAnalog_v0p0p1_1.RSfetsym_0.QN.t6 a_59577_n41283# GND.t1228 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X891 OUT0.t94 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND.t1158 GND.t1157 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X892 16to4_PriorityEncoder_v0p0p1_0.x36.Y 16to4_PriorityEncoder_v0p0p1_0.x36.A GND.t1470 GND.t1469 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X893 a_78599_n51085# 16to4_PriorityEncoder_v0p0p1_0.x3.x22.A a_78527_n51085# VDD.t867 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X894 OUT1.t37 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD.t328 VDD.t327 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X895 w_55000_n3550# VIN.t17 a_53630_n3996# GND.t1236 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X896 resistorDivider_v0p0p1_0.V6.t6 resistorDivider_v0p0p1_0.V5.t9 GND.t552 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X897 16to4_PriorityEncoder_v0p0p1_0.x3.x17.C a_77605_n51335# VDD.t140 VDD.t139 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.312 ps=1.68 w=1 l=0.15
X898 16to4_PriorityEncoder_v0p0p1_0.x43.Y 16to4_PriorityEncoder_v0p0p1_0.x43.A VDD.t682 VDD.t681 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X899 frontAnalog_v0p0p1_6.RSfetsym_0.x1.Y frontAnalog_v0p0p1_6.x63.X VDD.t46 VDD.t39 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X900 VDD.t1442 frontAnalog_v0p0p1_10.x65.A.t4 a_57123_n56559# VDD.t1441 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X901 VDD.t1395 16to4_PriorityEncoder_v0p0p1_0.x3.x14.A a_78315_n49349# VDD.t63 sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X902 frontAnalog_v0p0p1_0.RSfetsym_0.x1.Y frontAnalog_v0p0p1_0.x63.X VDD.t1497 VDD.t1490 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X903 frontAnalog_v0p0p1_3.RSfetsym_0.x2.Y frontAnalog_v0p0p1_3.x65.X GND.t697 GND.t696 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X904 frontAnalog_v0p0p1_13.RSfetsym_0.x1.Y frontAnalog_v0p0p1_13.x63.X GND.t541 GND.t539 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X905 resistorDivider_v0p0p1_0.V7.t13 resistorDivider_v0p0p1_0.V6.t11 GND.t26 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X906 GND.t335 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t98 GND.t334 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X907 VDD.t8 frontAnalog_v0p0p1_8.x65.X frontAnalog_v0p0p1_8.RSfetsym_0.x2.Y VDD.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X908 GND.t802 16to4_PriorityEncoder_v0p0p1_0.x5.x4.C a_78159_n39549# GND.t801 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X909 frontAnalog_v0p0p1_5.RSfetsym_0.QN.t4 16to4_PriorityEncoder_v0p0p1_0.I11.t8 VDD.t1488 VDD.t542 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.3
X910 resistorDivider_v0p0p1_0.V1.t4 VL.t1 GND.t84 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X911 GND.t195 frontAnalog_v0p0p1_12.x63.A.t6 a_57123_n74279# GND.t194 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X912 OUT2.t103 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND.t1029 GND.t1028 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X913 VDD.t1266 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t31 VDD.t1265 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X914 16to4_PriorityEncoder_v0p0p1_0.x5.x20.B 16to4_PriorityEncoder_v0p0p1_0.I14.t6 GND.t20 GND.t19 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X915 OUT0.t30 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD.t1108 VDD.t1107 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X916 OUT1.t36 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD.t326 VDD.t325 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X917 w_55000_n73750# VIN.t18 a_53630_n74196# GND.t1078 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X918 resistorDivider_v0p0p1_0.V9.t14 resistorDivider_v0p0p1_0.V8.t14 GND.t84 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X919 a_77605_n44527# 16to4_PriorityEncoder_v0p0p1_0.x5.x19.C VDD.t147 VDD.t33 sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.109 ps=1.36 w=0.42 l=0.15
X920 OUT2.t102 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND.t1027 GND.t1026 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X921 GND.t1025 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t101 GND.t1024 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X922 GND.t1468 16to4_PriorityEncoder_v0p0p1_0.x36.A 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND.t1467 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X923 frontAnalog_v0p0p1_14.RSfetsym_0.x1.Y frontAnalog_v0p0p1_14.x63.X VDD.t581 VDD.t577 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X924 OUT3.t30 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD.t1264 VDD.t1263 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X925 VDD.t723 frontAnalog_v0p0p1_3.x65.A.t4 a_57123_n13359# VDD.t722 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X926 frontAnalog_v0p0p1_5.RSfetsym_0.x2.Y frontAnalog_v0p0p1_5.x65.X VDD.t137 VDD.t131 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X927 VDD.t324 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t35 VDD.t323 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X928 frontAnalog_v0p0p1_5.RSfetsym_0.x1.Y frontAnalog_v0p0p1_5.x63.X GND.t648 GND.t646 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X929 frontAnalog_v0p0p1_6.RSfetsym_0.QN.t2 frontAnalog_v0p0p1_6.x65.X VDD.t478 VDD.t473 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.25
X930 VDD.t1262 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t29 VDD.t1261 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X931 VDD.t680 16to4_PriorityEncoder_v0p0p1_0.x43.A 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD.t679 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X932 GND.t919 16to4_PriorityEncoder_v0p0p1_0.x3.x22.A a_78525_n53555# GND.t918 sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X933 frontAnalog_v0p0p1_0.x65.X a_57123_n7959# VDD.t837 VDD.t836 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X934 GND.t1418 frontAnalog_v0p0p1_6.x63.A.t6 a_57123_n31079# GND.t1417 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X935 frontAnalog_v0p0p1_9.RSfetsym_0.QN.t2 frontAnalog_v0p0p1_9.x65.X VDD.t636 VDD.t631 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.25
X936 VDD.t616 frontAnalog_v0p0p1_1.x65.X frontAnalog_v0p0p1_1.RSfetsym_0.QN.t3 VDD.t613 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.25
X937 16to4_PriorityEncoder_v0p0p1_0.x5.GS a_78649_n39527# GND.t14 GND.t13 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.112 ps=1.04 w=0.65 l=0.15
X938 GND.t333 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t97 GND.t332 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X939 resistorDivider_v0p0p1_0.V10.t7 resistorDivider_v0p0p1_0.V9.t4 GND.t102 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X940 frontAnalog_v0p0p1_7.RSfetsym_0.x1.Y frontAnalog_v0p0p1_7.x63.X VDD.t733 VDD.t729 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X941 resistorDivider_v0p0p1_0.V15.t2 resistorDivider_v0p0p1_0.V14.t3 GND.t119 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X942 resistorDivider_v0p0p1_0.V3.t7 resistorDivider_v0p0p1_0.V2.t6 GND.t196 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X943 OUT3.t28 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD.t1260 VDD.t1259 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X944 OUT1.t96 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND.t331 GND.t330 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X945 VDD.t963 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t32 VDD.t962 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X946 resistorDivider_v0p0p1_0.V13.t11 resistorDivider_v0p0p1_0.V12.t11 GND.t102 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X947 frontAnalog_v0p0p1_12.x63.A.t3 frontAnalog_v0p0p1_12.x65.A.t5 VDD.t1349 VDD.t484 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X948 frontAnalog_v0p0p1_12.Q.t4 frontAnalog_v0p0p1_12.RSfetsym_0.x2.Y GND.t949 GND.t868 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.25
X949 GND.t1023 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t100 GND.t1022 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X950 a_77605_n39305# frontAnalog_v0p0p1_7.Q.t9 GND.t25 GND.t24 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X951 frontAnalog_v0p0p1_14.x65.X a_57123_n78159# VDD.t1436 VDD.t1435 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X952 GND.t1254 16to4_PriorityEncoder_v0p0p1_0.x3.x4.C a_78159_n47589# GND.t1253 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X953 16to4_PriorityEncoder_v0p0p1_0.x3.x16.C frontAnalog_v0p0p1_10.Q.t9 VDD.t551 VDD.t550 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X954 16to4_PriorityEncoder_v0p0p1_0.x36.Y 16to4_PriorityEncoder_v0p0p1_0.x36.A VDD.t1409 VDD.t1408 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X955 a_77723_n48817# 16to4_PriorityEncoder_v0p0p1_0.x3.EI a_77637_n48817# GND.t865 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X956 frontAnalog_v0p0p1_13.x63.A.t2 CLK.t36 w_55000_n68350# VDD.t13 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X957 a_82988_n51645# 16to4_PriorityEncoder_v0p0p1_0.x3.A0 a_82906_n51645# VDD.t826 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X958 VDD.t1376 frontAnalog_v0p0p1_15.x65.X frontAnalog_v0p0p1_15.RSfetsym_0.x2.Y VDD.t1371 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X959 GND.t1021 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t99 GND.t1020 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X960 GND.t589 frontAnalog_v0p0p1_10.Q.t10 a_77723_n49127# GND.t448 sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X961 16to4_PriorityEncoder_v0p0p1_0.x5.GS a_78649_n39527# VDD.t20 VDD.t19 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.167 ps=1.39 w=1 l=0.15
X962 a_59578_n62370# frontAnalog_v0p0p1_11.x65.X frontAnalog_v0p0p1_11.RSfetsym_0.QN.t1 GND.t942 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.315 ps=2.72 w=1 l=0.15
X963 a_59577_n52083# frontAnalog_v0p0p1_9.x63.X frontAnalog_v0p0p1_9.Q.t2 GND.t203 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X964 resistorDivider_v0p0p1_0.V8.t15 resistorDivider_v0p0p1_0.V7.t15 GND.t59 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X965 VDD.t580 frontAnalog_v0p0p1_14.x63.X frontAnalog_v0p0p1_14.Q.t1 VDD.t579 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.25
X966 16to4_PriorityEncoder_v0p0p1_0.x43.Y 16to4_PriorityEncoder_v0p0p1_0.x43.A GND.t764 GND.t763 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X967 frontAnalog_v0p0p1_6.x63.A.t0 frontAnalog_v0p0p1_6.x65.A.t4 VDD.t235 VDD.t234 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X968 GND.t329 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t95 GND.t328 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X969 OUT1.t94 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND.t327 GND.t326 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X970 VDD.t852 16to4_PriorityEncoder_v0p0p1_0.x5.x20.B a_77605_n44527# VDD.t33 sky130_fd_pr__pfet_01v8_hvt ad=0.312 pd=1.68 as=0.0588 ps=0.7 w=0.42 l=0.15
X971 VDD.t1258 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t27 VDD.t1257 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X972 w_55000_n78528# CLK.t37 frontAnalog_v0p0p1_14.x65.A.t3 VDD.t14 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X973 OUT1.t34 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD.t322 VDD.t321 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X974 16to4_PriorityEncoder_v0p0p1_0.x5.A2 a_78065_n41309# GND.t1511 GND.t1510 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.102 ps=0.99 w=0.65 l=0.15
X975 frontAnalog_v0p0p1_7.x65.X a_57123_n34959# VDD.t1356 VDD.t1355 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X976 frontAnalog_v0p0p1_5.x63.A.t2 CLK.t38 w_55000_n25150# VDD.t15 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X977 resistorDivider_v0p0p1_0.V1.t10 VL.t5 GND.t399 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X978 VDD.t16 CLK.t39 w_55000_n46128# GND.t11 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X979 VDD.t320 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t33 VDD.t319 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X980 frontAnalog_v0p0p1_8.RSfetsym_0.QN.t0 frontAnalog_v0p0p1_8.RSfetsym_0.x1.Y GND.t1 GND.t0 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.25
X981 VDD.t615 frontAnalog_v0p0p1_1.x65.X frontAnalog_v0p0p1_1.RSfetsym_0.x2.Y VDD.t610 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X982 16to4_PriorityEncoder_v0p0p1_0.x3.GS a_78649_n47567# GND.t598 GND.t597 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.112 ps=1.04 w=0.65 l=0.15
X983 OUT2.t31 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD.t959 VDD.t958 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X984 GND.t695 frontAnalog_v0p0p1_3.x65.X frontAnalog_v0p0p1_3.RSfetsym_0.x2.Y GND.t694 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X985 GND.t1311 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t90 GND.t1310 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X986 frontAnalog_v0p0p1_10.RSfetsym_0.x2.Y frontAnalog_v0p0p1_10.x65.X GND.t1441 GND.t1440 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X987 GND.t540 frontAnalog_v0p0p1_13.x63.X frontAnalog_v0p0p1_13.RSfetsym_0.x1.Y GND.t539 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X988 VDD.t3 frontAnalog_v0p0p1_11.x63.A.t5 a_57123_n63479# VDD.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X989 resistorDivider_v0p0p1_0.V9.t11 resistorDivider_v0p0p1_0.V8.t13 GND.t399 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X990 resistorDivider_v0p0p1_0.V11.t13 resistorDivider_v0p0p1_0.V10.t10 GND.t75 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X991 OUT1.t93 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND.t325 GND.t324 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X992 VDD.t17 CLK.t40 w_55000_n46750# GND.t12 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X993 frontAnalog_v0p0p1_2.RSfetsym_0.x1.Y frontAnalog_v0p0p1_2.x63.X GND.t1409 GND.t1407 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X994 VDD.t732 frontAnalog_v0p0p1_7.x63.X frontAnalog_v0p0p1_7.Q.t1 VDD.t731 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.25
X995 a_77775_n52819# frontAnalog_v0p0p1_13.Q.t9 a_77687_n52819# GND.t532 sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
X996 OUT3.t89 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND.t1309 GND.t1308 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X997 w_55000_n35328# CLK.t41 frontAnalog_v0p0p1_7.x65.A.t1 VDD.t18 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X998 GND.t1156 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t93 GND.t1155 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X999 VDD.t1344 frontAnalog_v0p0p1_9.x63.A.t4 frontAnalog_v0p0p1_9.x65.A.t1 VDD.t413 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1000 VDD.t1256 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t26 VDD.t1255 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1001 frontAnalog_v0p0p1_2.RSfetsym_0.x2.Y frontAnalog_v0p0p1_2.x65.X GND.t729 GND.t728 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1002 16to4_PriorityEncoder_v0p0p1_0.x36.A 16to4_PriorityEncoder_v0p0p1_0.x35.A GND.t51 GND.t50 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1003 a_55268_n84936# CLK.t42 GND.t804 GND.t803 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1004 GND.t461 16to4_PriorityEncoder_v0p0p1_0.x29.A 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND.t460 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1005 VDD.t444 16to4_PriorityEncoder_v0p0p1_0.x29.A 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD.t443 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1006 a_77605_n47345# frontAnalog_v0p0p1_14.Q.t9 GND.t66 GND.t65 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1007 frontAnalog_v0p0p1_10.x65.A.t1 frontAnalog_v0p0p1_10.x63.A.t6 a_55268_n57936# GND.t249 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1008 OUT3.t25 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD.t1254 VDD.t1253 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1009 VDD.t318 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t32 VDD.t317 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1010 VDD.t578 frontAnalog_v0p0p1_14.x63.X frontAnalog_v0p0p1_14.RSfetsym_0.x1.Y VDD.t577 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1011 resistorDivider_v0p0p1_0.V7.t2 resistorDivider_v0p0p1_0.V6.t0 GND.t60 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1012 frontAnalog_v0p0p1_13.RSfetsym_0.x2.Y frontAnalog_v0p0p1_13.x65.X VDD.t129 VDD.t123 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1013 GND.t647 frontAnalog_v0p0p1_5.x63.X frontAnalog_v0p0p1_5.RSfetsym_0.x1.Y GND.t646 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1014 a_78315_n49349# 16to4_PriorityEncoder_v0p0p1_0.x3.x14.B a_78243_n49349# VDD.t63 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X1015 VDD.t1190 frontAnalog_v0p0p1_4.x63.A.t6 a_57123_n20279# VDD.t1189 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1016 a_53630_n63396# resistorDivider_v0p0p1_0.V5.t16 w_55000_n62328# GND.t792 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1017 16to4_PriorityEncoder_v0p0p1_0.x3.GS a_78649_n47567# VDD.t560 VDD.t559 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.167 ps=1.39 w=1 l=0.15
X1018 OUT3.t88 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND.t1307 GND.t1306 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1019 GND.t1019 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t98 GND.t1018 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1020 a_55268_n41736# CLK.t43 GND.t806 GND.t805 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1021 VIN.t19 w_55000_n2928# error sky130_fd_pr__cap_var_lvt w=2 l=0.18
X1022 OUT2.t30 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD.t957 VDD.t956 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1023 VDD.t1106 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t29 VDD.t1105 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1024 GND.t323 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t92 GND.t322 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1025 VDD.t955 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t29 VDD.t954 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1026 16to4_PriorityEncoder_v0p0p1_0.x43.Y 16to4_PriorityEncoder_v0p0p1_0.x43.A VDD.t678 VDD.t677 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1027 frontAnalog_v0p0p1_3.x65.A.t3 frontAnalog_v0p0p1_3.x63.A.t6 a_55268_n14736# GND.t874 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1028 VDD.t316 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t31 VDD.t315 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1029 VDD.t730 frontAnalog_v0p0p1_7.x63.X frontAnalog_v0p0p1_7.RSfetsym_0.x1.Y VDD.t729 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1030 16to4_PriorityEncoder_v0p0p1_0.x29.Y 16to4_PriorityEncoder_v0p0p1_0.x29.A GND.t459 GND.t458 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1031 VDD.t953 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t28 VDD.t952 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1032 16to4_PriorityEncoder_v0p0p1_0.x5.x18.C frontAnalog_v0p0p1_6.Q.t8 GND.t499 GND.t498 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1033 16to4_PriorityEncoder_v0p0p1_0.x29.Y 16to4_PriorityEncoder_v0p0p1_0.x29.A VDD.t442 VDD.t441 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1034 GND.t1154 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t92 GND.t1153 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1035 OUT3.t87 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND.t1305 GND.t1304 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1036 OUT0.t91 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND.t1152 GND.t1151 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1037 frontAnalog_v0p0p1_0.RSfetsym_0.x2.Y frontAnalog_v0p0p1_0.x65.X GND.t258 GND.t257 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1038 GND.t716 frontAnalog_v0p0p1_9.x65.X frontAnalog_v0p0p1_9.RSfetsym_0.x2.Y GND.t715 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1039 GND.t1303 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t86 GND.t1302 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1040 VIN.t20 w_55000_n73128# error sky130_fd_pr__cap_var_lvt w=2 l=0.18
X1041 resistorDivider_v0p0p1_0.V14.t10 resistorDivider_v0p0p1_0.V13.t9 GND.t75 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1042 OUT3.t24 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD.t1252 VDD.t1251 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1043 VDD.t889 frontAnalog_v0p0p1_11.x65.X frontAnalog_v0p0p1_11.RSfetsym_0.QN.t2 VDD.t888 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.25
X1044 VDD.t951 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t27 VDD.t950 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1045 OUT2.t26 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD.t949 VDD.t948 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1046 VDD.t676 16to4_PriorityEncoder_v0p0p1_0.x43.A 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD.t675 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1047 OUT1.t30 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD.t314 VDD.t313 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1048 16to4_PriorityEncoder_v0p0p1_0.x1.X a_82906_n47995# VDD.t706 VDD.t705 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.146 ps=1.34 w=1 l=0.15
X1049 a_16599_n13205.t1 a_16599_n13205.t0 GND.t828 GND.t827 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1050 VDD.t1104 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t28 VDD.t1103 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1051 frontAnalog_v0p0p1_12.x65.A.t1 CLK.t44 frontAnalog_v0p0p1_12.x63.A.t1 VDD.t717 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1052 GND.t1150 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t90 GND.t1149 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1053 OUT0.t89 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND.t1148 GND.t1147 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1054 frontAnalog_v0p0p1_1.x63.X a_57123_n41879# VDD.t576 VDD.t575 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1055 a_53630_n47196# frontAnalog_v0p0p1_10.IB.t16 GND.t932 GND.t186 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1056 w_55000_n57550# VIN.t21 a_53630_n57996# GND.t545 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1057 GND.t116 frontAnalog_v0p0p1_11.x63.X frontAnalog_v0p0p1_11.RSfetsym_0.x1.Y GND.t113 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1058 OUT0.t27 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD.t1102 VDD.t1101 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1059 16to4_PriorityEncoder_v0p0p1_0.x5.x9.Y VDD.t766 VDD.t768 VDD.t767 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1060 frontAnalog_v0p0p1_14.RSfetsym_0.x2.Y frontAnalog_v0p0p1_14.x65.X GND.t851 GND.t850 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1061 frontAnalog_v0p0p1_0.x63.A.t3 frontAnalog_v0p0p1_0.x65.A.t4 VDD.t1181 VDD.t103 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1062 GND.t1439 frontAnalog_v0p0p1_10.x65.X frontAnalog_v0p0p1_10.RSfetsym_0.x2.Y GND.t1438 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1063 OUT1.t91 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND.t321 GND.t320 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1064 resistorDivider_v0p0p1_0.V16.t17 w_55000_n3550# error sky130_fd_pr__cap_var_lvt w=2 l=0.18
X1065 16to4_PriorityEncoder_v0p0p1_0.x29.A 16to4_PriorityEncoder_v0p0p1_0.x28.A GND.t92 GND.t91 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1066 OUT1.t29 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD.t312 VDD.t311 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1067 GND.t1408 frontAnalog_v0p0p1_2.x63.X frontAnalog_v0p0p1_2.RSfetsym_0.x1.Y GND.t1407 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1068 GND.t825 frontAnalog_v0p0p1_12.x65.A.t6 a_57123_n72759# GND.t194 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X1069 16to4_PriorityEncoder_v0p0p1_0.x5.x21.B a_77605_n44527# VDD.t160 VDD.t159 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.312 ps=1.68 w=1 l=0.15
X1070 OUT0.t88 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND.t1146 GND.t1145 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1071 a_16719_n13117.t12 a_16599_n13205.t11 a_16541_n13117.t1 GND.t1562 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1072 resistorDivider_v0p0p1_0.V11.t4 resistorDivider_v0p0p1_0.V10.t5 GND.t119 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1073 frontAnalog_v0p0p1_6.x65.A.t1 CLK.t45 frontAnalog_v0p0p1_6.x63.A.t2 VDD.t718 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1074 frontAnalog_v0p0p1_12.Q.t0 frontAnalog_v0p0p1_12.RSfetsym_0.QN.t5 VDD.t403 VDD.t402 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.3
X1075 VDD.t591 frontAnalog_v0p0p1_12.x63.X frontAnalog_v0p0p1_12.RSfetsym_0.x1.Y VDD.t585 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1076 frontAnalog_v0p0p1_9.RSfetsym_0.x2.Y frontAnalog_v0p0p1_9.x65.X VDD.t635 VDD.t633 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1077 w_55000_n14350# VIN.t22 a_53630_n14796# GND.t546 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1078 frontAnalog_v0p0p1_7.RSfetsym_0.x2.Y frontAnalog_v0p0p1_7.x65.X GND.t1392 GND.t1391 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1079 GND.t1528 16to4_PriorityEncoder_v0p0p1_0.x22.A 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND.t1527 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1080 VDD.t1100 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t26 VDD.t1099 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1081 OUT0.t25 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD.t1098 VDD.t1097 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1082 VDD.t420 frontAnalog_v0p0p1_11.Q.t9 a_77855_n48109# VDD.t419 sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X1083 VDD.t146 16to4_PriorityEncoder_v0p0p1_0.x5.x19.C a_77605_n43545# VDD.t145 sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X1084 frontAnalog_v0p0p1_9.x63.X a_57123_n52679# GND.t561 GND.t406 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1085 16to4_PriorityEncoder_v0p0p1_0.x43.Y 16to4_PriorityEncoder_v0p0p1_0.x43.A GND.t762 GND.t761 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1086 frontAnalog_v0p0p1_10.Q.t3 frontAnalog_v0p0p1_10.RSfetsym_0.x2.Y GND.t622 GND.t621 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.25
X1087 resistorDivider_v0p0p1_0.V3.t17 w_55000_n73750# error sky130_fd_pr__cap_var_lvt w=2 l=0.18
X1088 OUT1.t28 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD.t310 VDD.t309 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1089 frontAnalog_v0p0p1_6.x63.A.t1 frontAnalog_v0p0p1_6.x65.A.t5 a_55268_n30936# GND.t246 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1090 OUT2.t25 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD.t947 VDD.t946 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1091 a_77687_n51335# frontAnalog_v0p0p1_12.Q.t8 a_77605_n51335# GND.t157 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.109 ps=1.36 w=0.42 l=0.15
X1092 VDD.t308 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t27 VDD.t307 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1093 frontAnalog_v0p0p1_6.Q.t3 frontAnalog_v0p0p1_6.RSfetsym_0.QN.t5 VDD.t654 VDD.t647 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.3
X1094 VDD.t45 frontAnalog_v0p0p1_6.x63.X frontAnalog_v0p0p1_6.RSfetsym_0.x1.Y VDD.t39 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1095 a_59578_n2970# frontAnalog_v0p0p1_2.x65.X frontAnalog_v0p0p1_2.RSfetsym_0.QN.t4 GND.t727 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.315 ps=2.72 w=1 l=0.15
X1096 OUT0.t24 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD.t1096 VDD.t1095 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1097 VDD.t1496 frontAnalog_v0p0p1_0.x63.X frontAnalog_v0p0p1_0.RSfetsym_0.x1.Y VDD.t1490 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1098 frontAnalog_v0p0p1_8.RSfetsym_0.x1.Y frontAnalog_v0p0p1_8.x63.X GND.t565 GND.t562 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1099 GND.t1144 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t87 GND.t1143 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1100 a_78065_n49349# 16to4_PriorityEncoder_v0p0p1_0.x3.x14.B GND.t83 GND.t82 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1101 a_59577_n35883# frontAnalog_v0p0p1_7.x63.X frontAnalog_v0p0p1_7.Q.t3 GND.t813 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1102 a_53630_n84996# frontAnalog_v0p0p1_10.IB.t17 GND.t933 GND.t186 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1103 VDD.t1461 16to4_PriorityEncoder_v0p0p1_0.x22.A 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD.t1460 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1104 a_77637_n42017# VDD.t763 VDD.t765 VDD.t764 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X1105 16to4_PriorityEncoder_v0p0p1_0.I13.t3 frontAnalog_v0p0p1_3.RSfetsym_0.x2.Y GND.t551 GND.t550 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.25
X1106 resistorDivider_v0p0p1_0.V11.t17 w_55000_n30550# error sky130_fd_pr__cap_var_lvt w=2 l=0.18
X1107 frontAnalog_v0p0p1_0.x63.A.t0 CLK.t46 w_55000_n8950# VDD.t719 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1108 GND.t1515 frontAnalog_v0p0p1_13.RSfetsym_0.QN.t6 a_59577_n68283# GND.t1514 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1109 16to4_PriorityEncoder_v0p0p1_0.x22.Y 16to4_PriorityEncoder_v0p0p1_0.x22.A GND.t1526 GND.t1525 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1110 GND.t68 frontAnalog_v0p0p1_14.Q.t10 a_59578_n78570# GND.t67 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1111 GND.t457 16to4_PriorityEncoder_v0p0p1_0.x29.A 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND.t456 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1112 16to4_PriorityEncoder_v0p0p1_0.I14.t3 frontAnalog_v0p0p1_0.x63.X VDD.t1495 VDD.t1493 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.25
X1113 resistorDivider_v0p0p1_0.V1.t15 VL.t7 GND.t102 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1114 GND.t256 frontAnalog_v0p0p1_0.x65.X frontAnalog_v0p0p1_0.RSfetsym_0.x2.Y GND.t255 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1115 VDD.t720 CLK.t47 w_55000_n29928# GND.t509 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1116 a_16719_n13117.t11 a_16599_n13205.t12 a_16541_n13117.t0 GND.t1563 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1117 OUT3.t23 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD.t1250 VDD.t1249 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1118 VDD.t306 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t26 VDD.t305 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1119 VDD.t136 frontAnalog_v0p0p1_5.x65.X frontAnalog_v0p0p1_5.RSfetsym_0.x2.Y VDD.t131 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1120 frontAnalog_v0p0p1_10.RSfetsym_0.x1.Y frontAnalog_v0p0p1_10.x63.X VDD.t176 VDD.t171 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1121 OUT2.t97 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND.t1017 GND.t1016 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1122 VDD.t1248 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t22 VDD.t1247 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1123 resistorDivider_v0p0p1_0.V9.t7 resistorDivider_v0p0p1_0.V8.t11 GND.t102 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1124 a_53630_n41796# frontAnalog_v0p0p1_10.IB.t18 GND.t934 GND.t186 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1125 16to4_PriorityEncoder_v0p0p1_0.x3.x14.B a_77637_n49127# GND.t840 GND.t548 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.112 ps=1.04 w=0.65 l=0.15
X1126 16to4_PriorityEncoder_v0p0p1_0.I14.t0 frontAnalog_v0p0p1_0.RSfetsym_0.QN.t6 VDD.t1179 VDD.t228 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.3
X1127 VDD.t703 16to4_PriorityEncoder_v0p0p1_0.x3.x19.C a_77605_n51585# VDD.t148 sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X1128 a_77605_n43545# 16to4_PriorityEncoder_v0p0p1_0.I11.t9 VDD.t1489 VDD.t145 sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.109 ps=1.36 w=0.42 l=0.15
X1129 resistorDivider_v0p0p1_0.V14.t13 resistorDivider_v0p0p1_0.V13.t13 GND.t119 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1130 VDD.t1094 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t23 VDD.t1093 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1131 GND.t1015 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t96 GND.t1014 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1132 GND.t584 frontAnalog_v0p0p1_5.RSfetsym_0.QN.t6 a_59577_n25083# GND.t583 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1133 frontAnalog_v0p0p1_6.x65.X a_57123_n29559# GND.t894 GND.t585 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1134 16to4_PriorityEncoder_v0p0p1_0.x3.x20.B frontAnalog_v0p0p1_9.Q.t10 VDD.t1341 VDD.t1340 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1135 GND.t740 frontAnalog_v0p0p1_7.Q.t10 a_59578_n35370# GND.t739 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1136 16to4_PriorityEncoder_v0p0p1_0.x5.x4.C a_77605_n40069# VDD.t558 VDD.t557 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.148 ps=1.34 w=1 l=0.15
X1137 a_77605_n52567# 16to4_PriorityEncoder_v0p0p1_0.x3.x18.C VDD.t115 VDD.t114 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X1138 16to4_PriorityEncoder_v0p0p1_0.x22.Y 16to4_PriorityEncoder_v0p0p1_0.x22.A VDD.t1459 VDD.t1458 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1139 frontAnalog_v0p0p1_15.x63.X a_57123_n85079# VDD.t200 VDD.t199 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1140 frontAnalog_v0p0p1_3.RSfetsym_0.x1.Y frontAnalog_v0p0p1_3.x63.X VDD.t227 VDD.t220 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1141 VDD.t1246 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t21 VDD.t1245 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1142 16to4_PriorityEncoder_v0p0p1_0.x29.Y 16to4_PriorityEncoder_v0p0p1_0.x29.A VDD.t440 VDD.t439 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1143 GND.t864 16to4_PriorityEncoder_v0p0p1_0.x3.EI a_77881_n51335# GND.t157 sky130_fd_pr__nfet_01v8 ad=0.196 pd=1.33 as=0.0693 ps=0.75 w=0.42 l=0.15
X1144 16to4_PriorityEncoder_v0p0p1_0.x3.x17.A a_77637_n50057# VDD.t211 VDD.t210 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.167 ps=1.39 w=1 l=0.15
X1145 a_77881_n44779# 16to4_PriorityEncoder_v0p0p1_0.x5.x19.C a_77775_n44779# GND.t155 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X1146 16to4_PriorityEncoder_v0p0p1_0.x3.x22.D a_77605_n53805# GND.t554 GND.t553 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X1147 resistorDivider_v0p0p1_0.V12.t12 resistorDivider_v0p0p1_0.V11.t12 GND.t889 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1148 OUT0.t86 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND.t1142 GND.t1141 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1149 VDD.t726 frontAnalog_v0p0p1_11.x65.A.t4 a_57123_n61959# VDD.t725 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1150 16to4_PriorityEncoder_v0p0p1_0.x22.A 16to4_PriorityEncoder_v0p0p1_0.x21.A GND.t610 GND.t609 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1151 GND.t251 frontAnalog_v0p0p1_10.x63.A.t7 a_57123_n58079# GND.t250 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X1152 frontAnalog_v0p0p1_14.RSfetsym_0.QN.t2 frontAnalog_v0p0p1_14.x65.X VDD.t788 VDD.t783 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.25
X1153 VDD.t634 frontAnalog_v0p0p1_9.x65.X frontAnalog_v0p0p1_9.RSfetsym_0.x2.Y VDD.t633 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1154 a_77783_n40069# 16to4_PriorityEncoder_v0p0p1_0.I14.t7 a_77687_n40069# VDD.t25 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X1155 VDD.t1244 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t20 VDD.t1243 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1156 VDD.t721 CLK.t48 w_55000_n8328# GND.t512 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1157 OUT1.t25 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD.t304 VDD.t303 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1158 resistorDivider_v0p0p1_0.V5.t0 resistorDivider_v0p0p1_0.V4.t2 GND.t84 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1159 GND.t1013 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t95 GND.t1012 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1160 OUT3.t19 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD.t1242 VDD.t1241 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1161 a_77605_n51585# frontAnalog_v0p0p1_13.Q.t10 VDD.t1033 VDD.t148 sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.109 ps=1.36 w=0.42 l=0.15
X1162 VDD.t438 16to4_PriorityEncoder_v0p0p1_0.x29.A 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD.t437 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1163 GND.t875 frontAnalog_v0p0p1_3.x63.A.t7 a_57123_n14879# GND.t807 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X1164 VDD.t743 CLK.t49 w_55000_n8950# GND.t736 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1165 frontAnalog_v0p0p1_7.RSfetsym_0.QN.t2 frontAnalog_v0p0p1_7.x65.X VDD.t1336 VDD.t1331 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.25
X1166 frontAnalog_v0p0p1_12.x63.A.t2 frontAnalog_v0p0p1_12.x65.A.t7 a_55268_n74136# GND.t826 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1167 OUT0.t22 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD.t1092 VDD.t1091 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1168 VDD.t762 VDD.t761 a_77605_n43545# VDD.t145 sky130_fd_pr__pfet_01v8_hvt ad=0.312 pd=1.68 as=0.0588 ps=0.7 w=0.42 l=0.15
X1169 16to4_PriorityEncoder_v0p0p1_0.x22.A 16to4_PriorityEncoder_v0p0p1_0.x21.A VDD.t569 VDD.t568 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1170 VDD.t1485 16to4_PriorityEncoder_v0p0p1_0.x5.x21.B a_78097_n45737# VDD.t1484 sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X1171 frontAnalog_v0p0p1_4.RSfetsym_0.x1.Y frontAnalog_v0p0p1_4.x63.X VDD.t59 VDD.t57 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1172 a_59577_n79083# frontAnalog_v0p0p1_14.x63.X frontAnalog_v0p0p1_14.Q.t0 GND.t636 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1173 a_77855_n48109# frontAnalog_v0p0p1_10.Q.t11 a_77783_n48109# VDD.t552 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X1174 a_78349_n43045# 16to4_PriorityEncoder_v0p0p1_0.x5.x17.D GND.t492 GND.t252 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X1175 GND.t1011 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t94 GND.t1010 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1176 a_77605_n45765# 16to4_PriorityEncoder_v0p0p1_0.x5.x20.B VDD.t851 VDD.t850 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X1177 GND.t319 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t90 GND.t318 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1178 frontAnalog_v0p0p1_0.RSfetsym_0.QN.t0 16to4_PriorityEncoder_v0p0p1_0.I14.t8 VDD.t229 VDD.t228 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.3
X1179 frontAnalog_v0p0p1_10.x63.A.t2 frontAnalog_v0p0p1_10.x65.A.t5 VDD.t1443 VDD.t409 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1180 GND.t726 frontAnalog_v0p0p1_2.x65.X frontAnalog_v0p0p1_2.RSfetsym_0.x2.Y GND.t725 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1181 a_55268_n3936# CLK.t50 GND.t830 GND.t829 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1182 frontAnalog_v0p0p1_1.RSfetsym_0.x1.Y frontAnalog_v0p0p1_1.x63.X VDD.t166 VDD.t162 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1183 OUT3.t18 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD.t1240 VDD.t1239 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1184 a_53630_n30996# frontAnalog_v0p0p1_10.IB.t19 GND.t935 GND.t186 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1185 16to4_PriorityEncoder_v0p0p1_0.x29.Y 16to4_PriorityEncoder_v0p0p1_0.x29.A GND.t455 GND.t454 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1186 GND.t1524 16to4_PriorityEncoder_v0p0p1_0.x22.A 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND.t1523 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1187 OUT3.t85 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND.t1301 GND.t1300 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1188 16to4_PriorityEncoder_v0p0p1_0.x5.x19.C 16to4_PriorityEncoder_v0p0p1_0.I12.t9 GND.t28 GND.t27 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1189 VDD.t128 frontAnalog_v0p0p1_13.x65.X frontAnalog_v0p0p1_13.RSfetsym_0.x2.Y VDD.t123 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1190 a_59578_n46170# frontAnalog_v0p0p1_8.x65.X frontAnalog_v0p0p1_8.RSfetsym_0.QN.t1 GND.t6 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.315 ps=2.72 w=1 l=0.15
X1191 VDD.t52 16to4_PriorityEncoder_v0p0p1_0.x35.A 16to4_PriorityEncoder_v0p0p1_0.x36.A VDD.t51 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1192 frontAnalog_v0p0p1_12.Q.t3 frontAnalog_v0p0p1_12.x63.X VDD.t590 VDD.t587 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.25
X1193 frontAnalog_v0p0p1_3.x63.A.t2 frontAnalog_v0p0p1_3.x65.A.t5 VDD.t724 VDD.t471 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1194 VDD.t1046 frontAnalog_v0p0p1_14.x63.A.t6 frontAnalog_v0p0p1_14.x65.A.t1 VDD.t651 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1195 OUT3.t17 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD.t1238 VDD.t1237 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1196 frontAnalog_v0p0p1_4.x65.X a_57123_n18759# VDD.t666 VDD.t665 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1197 OUT2.t93 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND.t1009 GND.t1008 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1198 OUT2.t24 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD.t945 VDD.t944 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1199 VDD.t674 16to4_PriorityEncoder_v0p0p1_0.x43.A 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD.t673 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1200 OUT1.t24 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD.t302 VDD.t301 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1201 frontAnalog_v0p0p1_6.RSfetsym_0.QN.t4 frontAnalog_v0p0p1_6.RSfetsym_0.x1.Y GND.t1489 GND.t1488 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.25
X1202 VDD.t800 16to4_PriorityEncoder_v0p0p1_0.x3.EI a_77605_n51585# VDD.t148 sky130_fd_pr__pfet_01v8_hvt ad=0.312 pd=1.68 as=0.0588 ps=0.7 w=0.42 l=0.15
X1203 16to4_PriorityEncoder_v0p0p1_0.x3.A1 a_78349_n51085# GND.t876 GND.t151 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.102 ps=0.99 w=0.65 l=0.15
X1204 resistorDivider_v0p0p1_0.V7.t14 resistorDivider_v0p0p1_0.V6.t14 GND.t59 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1205 VDD.t1457 16to4_PriorityEncoder_v0p0p1_0.x22.A 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD.t1456 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1206 OUT1.t89 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND.t317 GND.t316 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1207 VDD.t189 frontAnalog_v0p0p1_8.x63.A.t5 a_57123_n47279# VDD.t188 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1208 VDD.t527 16to4_PriorityEncoder_v0p0p1_0.x3.x21.B a_78097_n53777# VDD.t526 sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X1209 VDD.t744 CLK.t51 w_55000_n51528# GND.t12 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1210 frontAnalog_v0p0p1_6.Q.t2 frontAnalog_v0p0p1_6.x63.X VDD.t44 VDD.t41 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.25
X1211 VDD.t539 frontAnalog_v0p0p1_7.x63.A.t5 frontAnalog_v0p0p1_7.x65.A.t2 VDD.t538 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1212 GND.t1299 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t84 GND.t1298 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1213 a_77605_n53805# 16to4_PriorityEncoder_v0p0p1_0.x3.x20.B VDD.t491 VDD.t490 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X1214 frontAnalog_v0p0p1_11.RSfetsym_0.x2.Y frontAnalog_v0p0p1_11.x65.X GND.t941 GND.t940 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1215 a_55268_n68736# CLK.t52 GND.t832 GND.t831 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1216 OUT3.t16 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD.t1236 VDD.t1235 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1217 resistorDivider_v0p0p1_0.V16.t1 resistorDivider_v0p0p1_0.V15.t5 GND.t26 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1218 VDD.t745 CLK.t53 w_55000_n52150# GND.t833 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1219 resistorDivider_v0p0p1_0.V5.t5 resistorDivider_v0p0p1_0.V4.t7 GND.t399 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1220 16to4_PriorityEncoder_v0p0p1_0.x3.x18.C frontAnalog_v0p0p1_12.Q.t9 VDD.t1392 VDD.t1391 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1221 VDD.t165 frontAnalog_v0p0p1_1.x63.X frontAnalog_v0p0p1_1.Q.t0 VDD.t164 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.25
X1222 OUT3.t83 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND.t1297 GND.t1296 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1223 frontAnalog_v0p0p1_12.RSfetsym_0.QN.t3 frontAnalog_v0p0p1_12.Q.t10 VDD.t1393 VDD.t402 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.3
X1224 a_77759_n53805# 16to4_PriorityEncoder_v0p0p1_0.x3.x20.B a_77687_n53805# GND.t535 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X1225 frontAnalog_v0p0p1_9.x65.X a_57123_n51159# GND.t407 GND.t406 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1226 w_55000_n40728# CLK.t54 frontAnalog_v0p0p1_1.x65.A.t1 VDD.t746 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1227 VDD.t1234 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t15 VDD.t1233 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1228 16to4_PriorityEncoder_v0p0p1_0.I15.t4 frontAnalog_v0p0p1_2.RSfetsym_0.x2.Y GND.t1507 GND.t719 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.25
X1229 GND.t244 16to4_PriorityEncoder_v0p0p1_0.I14.t9 a_77605_n40069# GND.t243 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X1230 GND.t1295 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t82 GND.t1294 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1231 frontAnalog_v0p0p1_11.x65.A.t3 frontAnalog_v0p0p1_11.x63.A.t6 a_55268_n63336# GND.t1230 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1232 a_53630_n47196# resistorDivider_v0p0p1_0.V8.t16 w_55000_n46128# GND.t421 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1233 a_78349_n51085# 16to4_PriorityEncoder_v0p0p1_0.x3.x22.A GND.t917 GND.t165 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1234 GND.t1486 16to4_PriorityEncoder_v0p0p1_0.I14.t10 a_59578_n8370# GND.t1485 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1235 frontAnalog_v0p0p1_12.RSfetsym_0.x2.Y frontAnalog_v0p0p1_12.x65.X VDD.t76 VDD.t74 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1236 a_77637_n41087# VDD.t759 VDD.t760 VDD.t230 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X1237 a_55268_n25536# CLK.t55 GND.t835 GND.t834 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1238 frontAnalog_v0p0p1_12.RSfetsym_0.x1.Y frontAnalog_v0p0p1_12.x63.X GND.t642 GND.t640 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1239 a_78243_n49349# 16to4_PriorityEncoder_v0p0p1_0.x3.x17.A a_78147_n49349# VDD.t63 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X1240 GND.t849 frontAnalog_v0p0p1_14.x65.X frontAnalog_v0p0p1_14.RSfetsym_0.x2.Y GND.t848 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1241 OUT1.t88 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND.t315 GND.t314 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1242 a_82988_n47995# 16to4_PriorityEncoder_v0p0p1_0.x3.A1 a_82906_n47995# VDD.t1343 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X1243 GND.t313 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t87 GND.t312 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1244 a_77687_n40069# 16to4_PriorityEncoder_v0p0p1_0.I15.t6 a_77605_n40069# VDD.t1396 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X1245 VDD.t58 frontAnalog_v0p0p1_4.x63.X frontAnalog_v0p0p1_4.RSfetsym_0.x1.Y VDD.t57 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1246 VDD.t1232 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t14 VDD.t1231 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1247 frontAnalog_v0p0p1_0.x65.A.t3 frontAnalog_v0p0p1_0.x63.A.t4 a_55268_n9336# GND.t1225 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1248 GND.t311 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t86 GND.t310 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1249 OUT2.t23 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD.t943 VDD.t942 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1250 a_77687_n44527# 16to4_PriorityEncoder_v0p0p1_0.x5.x19.C a_77605_n44527# GND.t154 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.109 ps=1.36 w=0.42 l=0.15
X1251 GND.t878 16to4_PriorityEncoder_v0p0p1_0.x5.A2 a_82906_n43855# GND.t877 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X1252 VDD.t163 frontAnalog_v0p0p1_1.x63.X frontAnalog_v0p0p1_1.RSfetsym_0.x1.Y VDD.t162 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1253 frontAnalog_v0p0p1_15.RSfetsym_0.x1.Y frontAnalog_v0p0p1_15.x63.X VDD.t859 VDD.t855 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1254 VDD.t1176 frontAnalog_v0p0p1_0.x63.A.t5 a_57123_n9479# VDD.t1175 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1255 frontAnalog_v0p0p1_6.RSfetsym_0.x2.Y frontAnalog_v0p0p1_6.x65.X VDD.t477 VDD.t475 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1256 GND.t1140 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t85 GND.t1139 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1257 frontAnalog_v0p0p1_13.x63.X a_57123_n68879# VDD.t794 VDD.t793 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1258 frontAnalog_v0p0p1_6.RSfetsym_0.x1.Y frontAnalog_v0p0p1_6.x63.X GND.t42 GND.t40 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1259 GND.t1390 frontAnalog_v0p0p1_7.x65.X frontAnalog_v0p0p1_7.RSfetsym_0.x2.Y GND.t1389 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1260 resistorDivider_v0p0p1_0.V12.t4 resistorDivider_v0p0p1_0.V11.t5 GND.t552 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1261 a_77783_n39305# frontAnalog_v0p0p1_6.Q.t9 a_77687_n39305# VDD.t467 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X1262 VIN.t23 w_55000_n56928# error sky130_fd_pr__cap_var_lvt w=2 l=0.18
X1263 16to4_PriorityEncoder_v0p0p1_0.x22.Y 16to4_PriorityEncoder_v0p0p1_0.x22.A GND.t1522 GND.t1521 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1264 VDD.t672 16to4_PriorityEncoder_v0p0p1_0.x43.A 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD.t671 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1265 frontAnalog_v0p0p1_0.x63.X a_57123_n9479# GND.t873 GND.t872 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1266 VDD.t7 frontAnalog_v0p0p1_8.x65.X frontAnalog_v0p0p1_8.RSfetsym_0.QN.t2 VDD.t6 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.25
X1267 GND.t1396 frontAnalog_v0p0p1_9.Q.t11 a_77605_n48109# GND.t818 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X1268 OUT1.t85 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND.t309 GND.t308 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1269 GND.t307 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t84 GND.t306 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1270 OUT2.t22 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD.t941 VDD.t940 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1271 OUT3.t13 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD.t1230 VDD.t1229 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1272 frontAnalog_v0p0p1_10.x65.A.t3 CLK.t56 frontAnalog_v0p0p1_10.x63.A.t1 VDD.t116 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1273 frontAnalog_v0p0p1_5.x63.X a_57123_n25679# VDD.t395 VDD.t394 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1274 frontAnalog_v0p0p1_14.RSfetsym_0.x2.Y frontAnalog_v0p0p1_14.x65.X VDD.t787 VDD.t785 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1275 GND.t564 frontAnalog_v0p0p1_8.x63.X frontAnalog_v0p0p1_8.RSfetsym_0.x1.Y GND.t562 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1276 resistorDivider_v0p0p1_0.V8.t10 resistorDivider_v0p0p1_0.V7.t10 GND.t84 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1277 VIN.t24 w_55000_n13728# error sky130_fd_pr__cap_var_lvt w=2 l=0.18
X1278 frontAnalog_v0p0p1_14.x63.A.t3 frontAnalog_v0p0p1_14.x65.A.t6 VDD.t738 VDD.t14 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1279 VDD.t1090 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t21 VDD.t1089 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1280 VDD.t643 frontAnalog_v0p0p1_2.x65.X frontAnalog_v0p0p1_2.RSfetsym_0.QN.t2 VDD.t642 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.25
X1281 frontAnalog_v0p0p1_0.RSfetsym_0.x1.Y frontAnalog_v0p0p1_0.x63.X GND.t1557 GND.t1555 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1282 frontAnalog_v0p0p1_15.x65.X a_57123_n83559# VDD.t154 VDD.t153 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1283 GND.t1007 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t92 GND.t1006 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1284 frontAnalog_v0p0p1_14.x63.X a_57123_n79679# GND.t786 GND.t785 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1285 a_53630_n52596# frontAnalog_v0p0p1_10.IB.t20 GND.t705 GND.t186 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1286 16to4_PriorityEncoder_v0p0p1_0.x36.Y 16to4_PriorityEncoder_v0p0p1_0.x36.A VDD.t1407 VDD.t1406 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1287 frontAnalog_v0p0p1_12.x63.A.t0 CLK.t57 w_55000_n73750# VDD.t117 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1288 16to4_PriorityEncoder_v0p0p1_0.x22.Y 16to4_PriorityEncoder_v0p0p1_0.x22.A VDD.t1455 VDD.t1454 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1289 GND.t1293 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t81 GND.t1292 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1290 resistorDivider_v0p0p1_0.V2.t4 resistorDivider_v0p0p1_0.V1.t5 GND.t75 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1291 GND.t1506 frontAnalog_v0p0p1_10.x65.A.t6 a_57123_n56559# GND.t250 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X1292 OUT0.t84 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND.t1138 GND.t1137 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1293 a_77687_n52567# 16to4_PriorityEncoder_v0p0p1_0.x3.x19.C a_77605_n52567# GND.t131 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.109 ps=1.36 w=0.42 l=0.15
X1294 OUT3.t12 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD.t1228 VDD.t1227 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1295 frontAnalog_v0p0p1_10.x63.A.t3 frontAnalog_v0p0p1_10.x65.A.t7 a_55268_n57936# GND.t576 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1296 GND.t939 frontAnalog_v0p0p1_11.x65.X frontAnalog_v0p0p1_11.RSfetsym_0.x2.Y GND.t938 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1297 GND.t906 16to4_PriorityEncoder_v0p0p1_0.x5.x20.B a_77881_n44527# GND.t154 sky130_fd_pr__nfet_01v8 ad=0.196 pd=1.33 as=0.0693 ps=0.75 w=0.42 l=0.15
X1298 frontAnalog_v0p0p1_3.x65.A.t0 CLK.t58 frontAnalog_v0p0p1_3.x63.A.t1 VDD.t118 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1299 frontAnalog_v0p0p1_10.Q.t4 frontAnalog_v0p0p1_10.RSfetsym_0.QN.t5 VDD.t1194 VDD.t1027 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.3
X1300 frontAnalog_v0p0p1_7.RSfetsym_0.x2.Y frontAnalog_v0p0p1_7.x65.X VDD.t1335 VDD.t1333 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1301 VDD.t175 frontAnalog_v0p0p1_10.x63.X frontAnalog_v0p0p1_10.RSfetsym_0.x1.Y VDD.t171 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1302 VDD.t1226 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t11 VDD.t1225 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1303 VDD.t858 frontAnalog_v0p0p1_15.x63.X frontAnalog_v0p0p1_15.Q.t3 VDD.t857 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.25
X1304 VDD.t300 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t23 VDD.t299 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1305 frontAnalog_v0p0p1_4.RSfetsym_0.x2.Y frontAnalog_v0p0p1_4.x65.X GND.t899 GND.t898 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1306 w_55000_n83928# CLK.t59 frontAnalog_v0p0p1_15.x65.A.t2 VDD.t119 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1307 16to4_PriorityEncoder_v0p0p1_0.x5.x4.C a_77605_n40069# GND.t596 GND.t595 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.102 ps=0.99 w=0.65 l=0.15
X1308 a_77783_n47345# frontAnalog_v0p0p1_12.Q.t11 a_77687_n47345# VDD.t1394 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X1309 frontAnalog_v0p0p1_1.x65.X a_57123_n40359# VDD.t418 VDD.t417 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1310 a_16719_n13117.t10 a_16599_n13205.t13 a_16541_n13117.t15 GND.t1564 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1311 frontAnalog_v0p0p1_7.x63.X a_57123_n36479# GND.t690 GND.t689 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1312 resistorDivider_v0p0p1_0.V6.t17 w_55000_n57550# error sky130_fd_pr__cap_var_lvt w=2 l=0.18
X1313 OUT2.t21 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD.t939 VDD.t938 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1314 GND.t808 frontAnalog_v0p0p1_3.x65.A.t6 a_57123_n13359# GND.t807 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X1315 a_78527_n43045# 16to4_PriorityEncoder_v0p0p1_0.x5.x17.C a_78431_n43045# VDD.t242 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X1316 frontAnalog_v0p0p1_9.RSfetsym_0.QN.t0 frontAnalog_v0p0p1_9.RSfetsym_0.x1.Y GND.t227 GND.t226 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.25
X1317 frontAnalog_v0p0p1_2.RSfetsym_0.x2.Y frontAnalog_v0p0p1_2.x65.X VDD.t641 VDD.t639 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1318 resistorDivider_v0p0p1_0.V16.t7 resistorDivider_v0p0p1_0.V15.t9 GND.t60 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1319 frontAnalog_v0p0p1_3.x63.A.t3 frontAnalog_v0p0p1_3.x65.A.t7 a_55268_n14736# GND.t809 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1320 GND.t641 frontAnalog_v0p0p1_12.x63.X frontAnalog_v0p0p1_12.RSfetsym_0.x1.Y GND.t640 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1321 OUT1.t83 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND.t305 GND.t304 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1322 OUT2.t20 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD.t937 VDD.t936 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1323 VDD.t935 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t19 VDD.t934 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1324 VDD.t1405 16to4_PriorityEncoder_v0p0p1_0.x36.A 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD.t1404 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1325 OUT0.t20 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD.t1088 VDD.t1087 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1326 GND.t449 frontAnalog_v0p0p1_11.Q.t10 a_77723_n48817# GND.t448 sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X1327 16to4_PriorityEncoder_v0p0p1_0.I13.t4 frontAnalog_v0p0p1_3.RSfetsym_0.QN.t5 VDD.t1036 VDD.t181 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.3
X1328 frontAnalog_v0p0p1_0.x65.X a_57123_n7959# GND.t888 GND.t872 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1329 VDD.t226 frontAnalog_v0p0p1_3.x63.X frontAnalog_v0p0p1_3.RSfetsym_0.x1.Y VDD.t220 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1330 a_59577_n19683# frontAnalog_v0p0p1_4.x63.X 16to4_PriorityEncoder_v0p0p1_0.I12.t2 GND.t79 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1331 OUT0.t83 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND.t1136 GND.t1135 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1332 a_59578_n29970# frontAnalog_v0p0p1_6.x65.X frontAnalog_v0p0p1_6.RSfetsym_0.QN.t0 GND.t515 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.315 ps=2.72 w=1 l=0.15
X1333 a_53630_n68796# frontAnalog_v0p0p1_10.IB.t21 GND.t706 GND.t186 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1334 GND.t1134 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t82 GND.t1133 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1335 a_77605_n40069# 16to4_PriorityEncoder_v0p0p1_0.I15.t7 GND.t1450 GND.t243 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X1336 resistorDivider_v0p0p1_0.V14.t17 w_55000_n14350# error sky130_fd_pr__cap_var_lvt w=2 l=0.18
X1337 GND.t1132 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t81 GND.t1131 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1338 frontAnalog_v0p0p1_9.RSfetsym_0.x1.Y frontAnalog_v0p0p1_9.x63.X GND.t202 GND.t200 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1339 a_16719_n13117.t9 a_16599_n13205.t14 a_16541_n13117.t14 GND.t1565 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1340 a_77637_n40777# VDD.t756 VDD.t758 VDD.t757 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X1341 VDD.t856 frontAnalog_v0p0p1_15.x63.X frontAnalog_v0p0p1_15.RSfetsym_0.x1.Y VDD.t855 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1342 VDD.t298 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t22 VDD.t297 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1343 GND.t41 frontAnalog_v0p0p1_6.x63.X frontAnalog_v0p0p1_6.RSfetsym_0.x1.Y GND.t40 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1344 16to4_PriorityEncoder_v0p0p1_0.x43.A 16to4_PriorityEncoder_v0p0p1_0.x42.A GND.t746 GND.t745 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1345 GND.t420 frontAnalog_v0p0p1_12.RSfetsym_0.QN.t6 a_59577_n73683# GND.t419 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1346 OUT2.t91 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND.t1005 GND.t1004 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1347 GND.t396 frontAnalog_v0p0p1_15.Q.t8 a_59578_n83970# GND.t395 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1348 a_78147_n49349# 16to4_PriorityEncoder_v0p0p1_0.x3.x22.A a_78065_n49349# VDD.t63 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X1349 GND.t534 16to4_PriorityEncoder_v0p0p1_0.x3.x20.B a_77881_n52567# GND.t131 sky130_fd_pr__nfet_01v8 ad=0.196 pd=1.33 as=0.0693 ps=0.75 w=0.42 l=0.15
X1350 OUT1.t21 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD.t296 VDD.t295 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1351 16to4_PriorityEncoder_v0p0p1_0.x5.x22.C a_77605_n44779# GND.t837 GND.t836 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.196 ps=1.33 w=0.65 l=0.15
X1352 GND.t1003 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t90 GND.t1002 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1353 a_82906_n43855# 16to4_PriorityEncoder_v0p0p1_0.x3.A2 GND.t674 GND.t673 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1354 VDD.t933 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t18 VDD.t932 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1355 a_78313_n39305# 16to4_PriorityEncoder_v0p0p1_0.x5.x4.B a_78241_n39305# VDD.t838 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X1356 resistorDivider_v0p0p1_0.V8.t5 resistorDivider_v0p0p1_0.V7.t6 GND.t399 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1357 resistorDivider_v0p0p1_0.V10.t9 resistorDivider_v0p0p1_0.V9.t9 GND.t75 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1358 16to4_PriorityEncoder_v0p0p1_0.I13.t1 frontAnalog_v0p0p1_3.x63.X VDD.t225 VDD.t222 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.25
X1359 a_53630_n25596# frontAnalog_v0p0p1_10.IB.t22 GND.t707 GND.t186 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1360 a_16719_n13117.t8 a_16599_n13205.t15 a_16541_n13117.t13 GND.t1566 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1361 VDD.t1191 frontAnalog_v0p0p1_4.x63.A.t7 frontAnalog_v0p0p1_4.x65.A.t3 VDD.t531 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1362 frontAnalog_v0p0p1_11.RSfetsym_0.x1.Y frontAnalog_v0p0p1_11.x63.X VDD.t96 VDD.t94 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1363 OUT0.t19 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD.t1086 VDD.t1085 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1364 GND.t30 16to4_PriorityEncoder_v0p0p1_0.I12.t10 a_59578_n19170# GND.t29 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1365 resistorDivider_v0p0p1_0.V3.t11 resistorDivider_v0p0p1_0.V2.t10 GND.t889 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1366 VDD.t1084 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t18 VDD.t1083 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1367 resistorDivider_v0p0p1_0.V13.t1 resistorDivider_v0p0p1_0.V12.t0 GND.t75 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1368 OUT0.t80 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND.t1130 GND.t1129 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1369 GND.t1128 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t79 GND.t1127 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1370 resistorDivider_v0p0p1_0.V5.t6 resistorDivider_v0p0p1_0.V4.t9 GND.t102 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1371 VDD.t786 frontAnalog_v0p0p1_14.x65.X frontAnalog_v0p0p1_14.RSfetsym_0.x2.Y VDD.t785 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1372 a_78527_n51085# 16to4_PriorityEncoder_v0p0p1_0.x3.x17.C a_78431_n51085# VDD.t205 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X1373 GND.t49 16to4_PriorityEncoder_v0p0p1_0.x35.A 16to4_PriorityEncoder_v0p0p1_0.x36.A GND.t48 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1374 VDD.t931 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t17 VDD.t930 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1375 VDD.t1082 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t17 VDD.t1081 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1376 16to4_PriorityEncoder_v0p0p1_0.x3.A0 a_78525_n53555# GND.t1484 GND.t1483 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.102 ps=0.99 w=0.65 l=0.15
X1377 GND.t1234 frontAnalog_v0p0p1_6.RSfetsym_0.QN.t6 a_59577_n30483# GND.t1233 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1378 frontAnalog_v0p0p1_10.RSfetsym_0.QN.t0 frontAnalog_v0p0p1_10.Q.t12 VDD.t1028 VDD.t1027 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.3
X1379 frontAnalog_v0p0p1_7.x65.X a_57123_n34959# GND.t1405 GND.t689 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1380 GND.t417 frontAnalog_v0p0p1_1.Q.t7 a_59578_n40770# GND.t416 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1381 frontAnalog_v0p0p1_10.IB.t2 a_16719_n13117.t24 VDD.t1042 VDD.t1041 sky130_fd_pr__pfet_01v8_lvt ad=5.51 pd=38.6 as=5.51 ps=38.6 w=19 l=1
X1382 a_77687_n39305# 16to4_PriorityEncoder_v0p0p1_0.I11.t10 a_77605_n39305# VDD.t1199 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X1383 VDD.t294 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t20 VDD.t293 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1384 OUT1.t19 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD.t292 VDD.t291 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1385 OUT2.t89 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND.t1001 GND.t1000 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1386 GND.t999 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t88 GND.t998 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1387 16to4_PriorityEncoder_v0p0p1_0.x3.x14.A a_77637_n48817# VDD.t507 VDD.t506 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.167 ps=1.39 w=1 l=0.15
X1388 a_77605_n48109# frontAnalog_v0p0p1_8.Q.t7 GND.t819 GND.t818 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X1389 VDD.t87 frontAnalog_v0p0p1_8.x65.A.t4 a_57123_n45759# VDD.t86 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1390 VDD.t1334 frontAnalog_v0p0p1_7.x65.X frontAnalog_v0p0p1_7.RSfetsym_0.x2.Y VDD.t1333 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1391 16to4_PriorityEncoder_v0p0p1_0.x5.x16.C 16to4_PriorityEncoder_v0p0p1_0.I13.t11 VDD.t180 VDD.t179 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1392 resistorDivider_v0p0p1_0.V2.t3 resistorDivider_v0p0p1_0.V1.t3 GND.t119 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1393 VFS.t7 resistorDivider_v0p0p1_0.V16.t13 GND.t212 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1394 frontAnalog_v0p0p1_3.RSfetsym_0.QN.t4 16to4_PriorityEncoder_v0p0p1_0.I13.t12 VDD.t182 VDD.t181 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.3
X1395 OUT0.t16 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD.t1080 VDD.t1079 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1396 VDD.t1078 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t15 VDD.t1077 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1397 GND.t667 VDD.t1508 a_78735_n39527# GND.t666 sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X1398 VDD.t1044 a_16719_n13117.t25 a_16599_n13205.t3 VDD.t1043 sky130_fd_pr__pfet_01v8_lvt ad=5.51 pd=38.6 as=5.51 ps=38.6 w=19 l=1
X1399 OUT1.t18 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD.t290 VDD.t289 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1400 resistorDivider_v0p0p1_0.V4.t5 resistorDivider_v0p0p1_0.V3.t3 GND.t26 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1401 16to4_PriorityEncoder_v0p0p1_0.x3.x22.C a_77605_n52819# GND.t790 GND.t789 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.196 ps=1.33 w=0.65 l=0.15
X1402 16to4_PriorityEncoder_v0p0p1_0.x36.A 16to4_PriorityEncoder_v0p0p1_0.x35.A VDD.t50 VDD.t49 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1403 VDD.t436 16to4_PriorityEncoder_v0p0p1_0.x29.A 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD.t435 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1404 16to4_PriorityEncoder_v0p0p1_0.x3.x22.B a_78097_n53777# GND.t16 GND.t15 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.112 ps=1.04 w=0.65 l=0.15
X1405 w_55000_n62950# VIN.t25 a_53630_n63396# GND.t792 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1406 frontAnalog_v0p0p1_15.RSfetsym_0.x2.Y frontAnalog_v0p0p1_15.x65.X GND.t1424 GND.t1423 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1407 a_78313_n47345# 16to4_PriorityEncoder_v0p0p1_0.x3.x4.B a_78241_n47345# VDD.t563 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X1408 16to4_PriorityEncoder_v0p0p1_0.x36.Y 16to4_PriorityEncoder_v0p0p1_0.x36.A GND.t1466 GND.t1465 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1409 VDD.t640 frontAnalog_v0p0p1_2.x65.X frontAnalog_v0p0p1_2.RSfetsym_0.x2.Y VDD.t639 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1410 frontAnalog_v0p0p1_13.RSfetsym_0.x1.Y frontAnalog_v0p0p1_13.x63.X VDD.t499 VDD.t495 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1411 16to4_PriorityEncoder_v0p0p1_0.x3.x19.C frontAnalog_v0p0p1_11.Q.t11 VDD.t422 VDD.t421 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1412 frontAnalog_v0p0p1_4.RSfetsym_0.QN.t2 frontAnalog_v0p0p1_4.x65.X VDD.t847 VDD.t842 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.25
X1413 frontAnalog_v0p0p1_3.RSfetsym_0.x1.Y frontAnalog_v0p0p1_3.x63.X GND.t239 GND.t237 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1414 VFS.t4 resistorDivider_v0p0p1_0.V16.t8 GND.t693 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1415 OUT0.t78 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND.t1126 GND.t1125 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1416 a_77687_n47345# frontAnalog_v0p0p1_13.Q.t11 a_77605_n47345# VDD.t1034 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X1417 VDD.t929 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t16 VDD.t928 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1418 VDD.t288 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t17 VDD.t287 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1419 frontAnalog_v0p0p1_1.RSfetsym_0.x2.Y frontAnalog_v0p0p1_1.x65.X GND.t684 GND.t683 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1420 frontAnalog_v0p0p1_5.RSfetsym_0.x1.Y frontAnalog_v0p0p1_5.x63.X VDD.t597 VDD.t593 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1421 a_59577_n84483# frontAnalog_v0p0p1_15.x63.X frontAnalog_v0p0p1_15.Q.t2 GND.t910 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1422 a_77775_n44779# 16to4_PriorityEncoder_v0p0p1_0.I11.t11 a_77687_n44779# GND.t155 sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
X1423 OUT2.t87 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND.t997 GND.t996 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1424 frontAnalog_v0p0p1_11.Q.t4 frontAnalog_v0p0p1_11.RSfetsym_0.x2.Y GND.t1490 GND.t525 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.25
X1425 16to4_PriorityEncoder_v0p0p1_0.x29.Y 16to4_PriorityEncoder_v0p0p1_0.x29.A VDD.t434 VDD.t433 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1426 frontAnalog_v0p0p1_11.x63.A.t3 frontAnalog_v0p0p1_11.x65.A.t5 VDD.t728 VDD.t727 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1427 VDD.t1183 frontAnalog_v0p0p1_0.x65.A.t5 a_57123_n7959# VDD.t1182 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1428 GND.t1464 16to4_PriorityEncoder_v0p0p1_0.x36.A 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND.t1463 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1429 GND.t863 16to4_PriorityEncoder_v0p0p1_0.x3.EI a_78735_n47567# GND.t862 sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X1430 VDD.t120 CLK.t60 w_55000_n78528# GND.t132 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1431 OUT0.t14 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD.t1076 VDD.t1075 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1432 frontAnalog_v0p0p1_10.Q.t0 frontAnalog_v0p0p1_10.x63.X VDD.t174 VDD.t173 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.25
X1433 GND.t90 16to4_PriorityEncoder_v0p0p1_0.x28.A 16to4_PriorityEncoder_v0p0p1_0.x29.A GND.t89 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1434 a_77605_n44779# 16to4_PriorityEncoder_v0p0p1_0.x5.x19.C VDD.t144 VDD.t143 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X1435 VDD.t75 frontAnalog_v0p0p1_12.x65.X frontAnalog_v0p0p1_12.RSfetsym_0.x2.Y VDD.t74 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1436 GND.t861 16to4_PriorityEncoder_v0p0p1_0.x3.EI a_77759_n53805# GND.t860 sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X1437 a_59577_n41283# frontAnalog_v0p0p1_1.x63.X frontAnalog_v0p0p1_1.Q.t2 GND.t175 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1438 resistorDivider_v0p0p1_0.V10.t13 resistorDivider_v0p0p1_0.V9.t13 GND.t119 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1439 a_59578_n51570# frontAnalog_v0p0p1_9.x65.X frontAnalog_v0p0p1_9.RSfetsym_0.QN.t3 GND.t714 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.315 ps=2.72 w=1 l=0.15
X1440 VDD.t498 frontAnalog_v0p0p1_13.x63.X frontAnalog_v0p0p1_13.Q.t2 VDD.t497 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.25
X1441 VDD.t121 CLK.t61 w_55000_n79150# GND.t126 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1442 frontAnalog_v0p0p1_4.x63.A.t1 frontAnalog_v0p0p1_4.x65.A.t6 VDD.t185 VDD.t184 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1443 16to4_PriorityEncoder_v0p0p1_0.I12.t3 frontAnalog_v0p0p1_4.RSfetsym_0.x2.Y GND.t424 GND.t423 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.25
X1444 w_55000_n67728# CLK.t62 frontAnalog_v0p0p1_13.x65.A.t0 VDD.t122 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1445 VDD.t525 frontAnalog_v0p0p1_15.x63.A.t7 frontAnalog_v0p0p1_15.x65.A.t1 VDD.t85 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1446 OUT1.t82 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND.t303 GND.t302 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1447 frontAnalog_v0p0p1_14.x65.X a_57123_n78159# GND.t1492 GND.t785 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1448 resistorDivider_v0p0p1_0.V13.t5 resistorDivider_v0p0p1_0.V12.t5 GND.t119 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1449 frontAnalog_v0p0p1_5.x65.X a_57123_n24159# VDD.t562 VDD.t561 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1450 frontAnalog_v0p0p1_4.x63.X a_57123_n20279# GND.t925 GND.t749 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1451 GND.t995 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t86 GND.t994 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1452 frontAnalog_v0p0p1_3.x63.A.t0 CLK.t63 w_55000_n14350# VDD.t485 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1453 VDD.t486 CLK.t64 w_55000_n35328# GND.t527 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1454 GND.t160 16to4_PriorityEncoder_v0p0p1_0.x5.x22.C a_78525_n45515# GND.t159 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X1455 frontAnalog_v0p0p1_7.RSfetsym_0.QN.t0 frontAnalog_v0p0p1_7.RSfetsym_0.x1.Y GND.t537 GND.t536 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.25
X1456 VDD.t476 frontAnalog_v0p0p1_6.x65.X frontAnalog_v0p0p1_6.RSfetsym_0.x2.Y VDD.t475 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1457 frontAnalog_v0p0p1_8.RSfetsym_0.x2.Y frontAnalog_v0p0p1_8.x65.X GND.t5 GND.t4 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1458 VDD.t1346 frontAnalog_v0p0p1_9.x63.A.t5 a_57123_n52679# VDD.t1345 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1459 VDD.t596 frontAnalog_v0p0p1_5.x63.X 16to4_PriorityEncoder_v0p0p1_0.I11.t1 VDD.t595 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.25
X1460 VDD.t487 CLK.t65 w_55000_n35950# GND.t128 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1461 OUT1.t16 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD.t286 VDD.t285 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1462 16to4_PriorityEncoder_v0p0p1_0.x29.A 16to4_PriorityEncoder_v0p0p1_0.x28.A VDD.t67 VDD.t66 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1463 w_55000_n24528# CLK.t66 frontAnalog_v0p0p1_5.x65.A.t3 VDD.t488 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1464 GND.t1291 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t80 GND.t1290 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1465 a_16719_n13117.t23 a_16719_n13117.t22 VDD.t864 VDD.t863 sky130_fd_pr__pfet_01v8_lvt ad=5.51 pd=38.6 as=5.51 ps=38.6 w=19 l=1
X1466 a_53630_n3996# frontAnalog_v0p0p1_10.IB.t23 GND.t708 GND.t503 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1467 GND.t993 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t85 GND.t992 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1468 a_55268_n74136# CLK.t67 GND.t529 GND.t528 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1469 16to4_PriorityEncoder_v0p0p1_0.x43.Y 16to4_PriorityEncoder_v0p0p1_0.x43.A VDD.t670 VDD.t669 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1470 frontAnalog_v0p0p1_8.x65.A.t0 frontAnalog_v0p0p1_8.x63.A.t6 a_55268_n47136# GND.t108 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1471 VDD.t1432 16to4_PriorityEncoder_v0p0p1_0.I14.t11 a_77637_n42017# VDD.t764 sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X1472 16to4_PriorityEncoder_v0p0p1_0.x5.EO a_78159_n39549# GND.t220 GND.t219 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.102 ps=0.99 w=0.65 l=0.15
X1473 VDD.t496 frontAnalog_v0p0p1_13.x63.X frontAnalog_v0p0p1_13.RSfetsym_0.x1.Y VDD.t495 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1474 a_77605_n52819# 16to4_PriorityEncoder_v0p0p1_0.x3.x19.C VDD.t702 VDD.t701 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X1475 GND.t238 frontAnalog_v0p0p1_3.x63.X frontAnalog_v0p0p1_3.RSfetsym_0.x1.Y GND.t237 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1476 frontAnalog_v0p0p1_10.RSfetsym_0.x2.Y frontAnalog_v0p0p1_10.x65.X VDD.t1385 VDD.t1383 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1477 VFS.t2 resistorDivider_v0p0p1_0.V16.t5 GND.t615 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1478 frontAnalog_v0p0p1_10.RSfetsym_0.x1.Y frontAnalog_v0p0p1_10.x63.X GND.t182 GND.t180 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1479 a_53630_n52596# resistorDivider_v0p0p1_0.V7.t17 w_55000_n51528# GND.t210 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1480 a_16719_n13117.t7 a_16599_n13205.t16 a_16541_n13117.t12 GND.t1496 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1481 resistorDivider_v0p0p1_0.V3.t15 resistorDivider_v0p0p1_0.V2.t15 GND.t552 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1482 VDD.t1224 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t10 VDD.t1223 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1483 resistorDivider_v0p0p1_0.V4.t1 resistorDivider_v0p0p1_0.V3.t1 GND.t60 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1484 GND.t1556 frontAnalog_v0p0p1_0.x63.X frontAnalog_v0p0p1_0.RSfetsym_0.x1.Y GND.t1555 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1485 resistorDivider_v0p0p1_0.V8.t1 resistorDivider_v0p0p1_0.V7.t1 GND.t102 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1486 a_55268_n30936# CLK.t68 GND.t531 GND.t530 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1487 GND.t1231 frontAnalog_v0p0p1_11.x63.A.t7 a_57123_n63479# GND.t1094 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X1488 frontAnalog_v0p0p1_15.RSfetsym_0.QN.t2 frontAnalog_v0p0p1_15.x65.X VDD.t1375 VDD.t1374 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.25
X1489 GND.t991 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t84 GND.t990 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1490 OUT3.t9 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD.t1222 VDD.t1221 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1491 OUT1.t81 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND.t301 GND.t300 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1492 OUT2.t83 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND.t989 GND.t988 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1493 VDD.t594 frontAnalog_v0p0p1_5.x63.X frontAnalog_v0p0p1_5.RSfetsym_0.x1.Y VDD.t593 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1494 GND.t630 16to4_PriorityEncoder_v0p0p1_0.x3.x22.C a_78525_n53555# GND.t629 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X1495 frontAnalog_v0p0p1_3.RSfetsym_0.x2.Y frontAnalog_v0p0p1_3.x65.X VDD.t623 VDD.t621 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1496 16to4_PriorityEncoder_v0p0p1_0.x5.EO a_78159_n39549# VDD.t204 VDD.t203 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.148 ps=1.34 w=1 l=0.15
X1497 GND.t897 frontAnalog_v0p0p1_4.x65.X frontAnalog_v0p0p1_4.RSfetsym_0.x2.Y GND.t896 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1498 a_78159_n39549# 16to4_PriorityEncoder_v0p0p1_0.x5.x4.B GND.t891 GND.t890 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1499 OUT3.t8 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD.t1220 VDD.t1219 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1500 a_53630_n79596# frontAnalog_v0p0p1_10.IB.t24 GND.t709 GND.t186 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1501 frontAnalog_v0p0p1_1.RSfetsym_0.QN.t2 frontAnalog_v0p0p1_1.x65.X VDD.t614 VDD.t613 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.25
X1502 VDD.t474 frontAnalog_v0p0p1_6.x65.X frontAnalog_v0p0p1_6.RSfetsym_0.QN.t1 VDD.t473 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.25
X1503 VDD.t432 16to4_PriorityEncoder_v0p0p1_0.x29.A 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD.t431 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1504 OUT3.t79 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND.t1289 GND.t1288 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1505 resistorDivider_v0p0p1_0.V6.t2 resistorDivider_v0p0p1_0.V5.t3 GND.t212 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1506 16to4_PriorityEncoder_v0p0p1_0.x36.Y 16to4_PriorityEncoder_v0p0p1_0.x36.A GND.t1462 GND.t1461 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1507 16to4_PriorityEncoder_v0p0p1_0.x5.x22.A a_77639_n42341# GND.t628 GND.t627 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.112 ps=1.04 w=0.65 l=0.15
X1508 OUT1.t80 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND.t299 GND.t298 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1509 GND.t608 16to4_PriorityEncoder_v0p0p1_0.x21.A 16to4_PriorityEncoder_v0p0p1_0.x22.A GND.t607 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1510 VDD.t632 frontAnalog_v0p0p1_9.x65.X frontAnalog_v0p0p1_9.RSfetsym_0.QN.t1 VDD.t631 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.25
X1511 16to4_PriorityEncoder_v0p0p1_0.x3.EO a_78159_n47589# GND.t1086 GND.t1085 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.102 ps=0.99 w=0.65 l=0.15
X1512 OUT2.t15 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD.t927 VDD.t926 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1513 resistorDivider_v0p0p1_0.V1.t6 VL.t2 GND.t75 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1514 a_77687_n43295# frontAnalog_v0p0p1_6.Q.t10 a_77605_n43295# GND.t156 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.109 ps=1.36 w=0.42 l=0.15
X1515 VDD.t925 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t14 VDD.t924 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1516 frontAnalog_v0p0p1_11.x65.A.t1 CLK.t69 frontAnalog_v0p0p1_11.x63.A.t1 VDD.t489 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1517 frontAnalog_v0p0p1_13.x65.X a_57123_n67359# VDD.t1434 VDD.t1433 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1518 a_53630_n36396# frontAnalog_v0p0p1_10.IB.t25 GND.t616 GND.t186 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1519 OUT0.t77 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND.t1124 GND.t1123 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1520 OUT3.t7 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD.t1218 VDD.t1217 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1521 frontAnalog_v0p0p1_10.x63.A.t0 CLK.t70 w_55000_n57550# VDD.t108 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1522 GND.t201 frontAnalog_v0p0p1_9.x63.X frontAnalog_v0p0p1_9.RSfetsym_0.x1.Y GND.t200 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1523 16to4_PriorityEncoder_v0p0p1_0.x29.Y 16to4_PriorityEncoder_v0p0p1_0.x29.A GND.t453 GND.t452 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1524 resistorDivider_v0p0p1_0.V9.t3 resistorDivider_v0p0p1_0.V8.t7 GND.t75 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1525 frontAnalog_v0p0p1_14.RSfetsym_0.QN.t3 frontAnalog_v0p0p1_14.RSfetsym_0.x1.Y GND.t869 GND.t868 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.25
X1526 resistorDivider_v0p0p1_0.V6.t12 resistorDivider_v0p0p1_0.V5.t13 GND.t693 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1527 OUT3.t78 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND.t1287 GND.t1286 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1528 VDD.t1216 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t6 VDD.t1215 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1529 resistorDivider_v0p0p1_0.V16.t14 resistorDivider_v0p0p1_0.V15.t13 GND.t59 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1530 frontAnalog_v0p0p1_15.x63.X a_57123_n85079# GND.t206 GND.t161 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1531 GND.t3 frontAnalog_v0p0p1_8.x65.X frontAnalog_v0p0p1_8.RSfetsym_0.x2.Y GND.t2 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1532 resistorDivider_v0p0p1_0.V7.t11 resistorDivider_v0p0p1_0.V6.t7 GND.t84 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1533 GND.t1285 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t77 GND.t1284 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1534 frontAnalog_v0p0p1_4.RSfetsym_0.x2.Y frontAnalog_v0p0p1_4.x65.X VDD.t846 VDD.t844 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1535 GND.t1095 frontAnalog_v0p0p1_11.x65.A.t6 a_57123_n61959# GND.t1094 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X1536 VDD.t567 16to4_PriorityEncoder_v0p0p1_0.x21.A 16to4_PriorityEncoder_v0p0p1_0.x22.A VDD.t566 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1537 a_16719_n13117.t6 a_16599_n13205.t17 a_16541_n13117.t11 GND.t1497 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1538 16to4_PriorityEncoder_v0p0p1_0.x3.EO a_78159_n47589# VDD.t1040 VDD.t1039 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.148 ps=1.34 w=1 l=0.15
X1539 a_78159_n47589# 16to4_PriorityEncoder_v0p0p1_0.x3.x4.B GND.t604 GND.t603 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1540 VDD.t95 frontAnalog_v0p0p1_11.x63.X frontAnalog_v0p0p1_11.RSfetsym_0.x1.Y VDD.t94 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1541 frontAnalog_v0p0p1_1.RSfetsym_0.x2.Y frontAnalog_v0p0p1_1.x65.X VDD.t612 VDD.t610 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1542 OUT2.t82 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND.t987 GND.t986 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1543 frontAnalog_v0p0p1_5.RSfetsym_0.x2.Y frontAnalog_v0p0p1_5.x65.X GND.t145 GND.t144 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1544 frontAnalog_v0p0p1_14.RSfetsym_0.x1.Y frontAnalog_v0p0p1_14.x63.X GND.t635 GND.t633 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1545 OUT1.t79 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND.t297 GND.t296 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1546 a_78525_n45515# 16to4_PriorityEncoder_v0p0p1_0.x5.x22.D GND.t172 GND.t171 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X1547 OUT0.t13 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD.t1074 VDD.t1073 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1548 16to4_PriorityEncoder_v0p0p1_0.x5.x20.B 16to4_PriorityEncoder_v0p0p1_0.I14.t12 VDD.t742 VDD.t741 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1549 16to4_PriorityEncoder_v0p0p1_0.x35.A 16to4_PriorityEncoder_v0p0p1_0.x34.A GND.t413 GND.t412 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1550 16to4_PriorityEncoder_v0p0p1_0.x3.x22.A a_77639_n50381# GND.t1434 GND.t1433 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.112 ps=1.04 w=0.65 l=0.15
X1551 frontAnalog_v0p0p1_1.x63.X a_57123_n41879# GND.t631 GND.t439 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1552 GND.t181 frontAnalog_v0p0p1_10.x63.X frontAnalog_v0p0p1_10.RSfetsym_0.x1.Y GND.t180 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1553 resistorDivider_v0p0p1_0.V5.t17 w_55000_n62950# error sky130_fd_pr__cap_var_lvt w=2 l=0.18
X1554 OUT1.t78 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND.t295 GND.t294 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1555 GND.t293 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t77 GND.t292 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1556 GND.t451 16to4_PriorityEncoder_v0p0p1_0.x29.A 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND.t450 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1557 a_77605_n44527# 16to4_PriorityEncoder_v0p0p1_0.x5.x18.C VDD.t1397 VDD.t33 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X1558 VDD.t923 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t13 VDD.t922 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1559 a_77881_n43545# 16to4_PriorityEncoder_v0p0p1_0.x5.x16.C a_77775_n43545# GND.t153 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X1560 GND.t668 VDD.t1509 a_77881_n43295# GND.t156 sky130_fd_pr__nfet_01v8 ad=0.196 pd=1.33 as=0.0693 ps=0.75 w=0.42 l=0.15
X1561 a_77725_n42341# VDD.t1510 a_77639_n42341# GND.t669 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X1562 OUT3.t76 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND.t1283 GND.t1282 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1563 frontAnalog_v0p0p1_7.RSfetsym_0.x1.Y frontAnalog_v0p0p1_7.x63.X GND.t812 GND.t810 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1564 OUT0.t76 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND.t1122 GND.t1121 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1565 16to4_PriorityEncoder_v0p0p1_0.x5.x22.D a_77605_n45765# GND.t853 GND.t852 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X1566 VDD.t554 16to4_PriorityEncoder_v0p0p1_0.x5.x22.A a_78775_n45515# VDD.t553 sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X1567 GND.t1281 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t75 GND.t1280 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1568 GND.t1248 frontAnalog_v0p0p1_10.RSfetsym_0.QN.t6 a_59577_n57483# GND.t1247 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1569 GND.t1436 frontAnalog_v0p0p1_13.Q.t12 a_59578_n67770# GND.t1435 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1570 VDD.t921 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t12 VDD.t920 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1571 16to4_PriorityEncoder_v0p0p1_0.x43.Y 16to4_PriorityEncoder_v0p0p1_0.x43.A VDD.t668 VDD.t667 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1572 VDD.t284 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t15 VDD.t283 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1573 a_16719_n13117.t5 a_16599_n13205.t18 a_16541_n13117.t10 GND.t1498 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1574 16to4_PriorityEncoder_v0p0p1_0.x43.Y 16to4_PriorityEncoder_v0p0p1_0.x43.A GND.t760 GND.t759 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1575 frontAnalog_v0p0p1_2.x63.X a_57123_n4079# VDD.t1358 VDD.t1357 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1576 GND.t291 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t76 GND.t290 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1577 GND.t1422 frontAnalog_v0p0p1_15.x65.X frontAnalog_v0p0p1_15.RSfetsym_0.x2.Y GND.t1421 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1578 16to4_PriorityEncoder_v0p0p1_0.x29.Y 16to4_PriorityEncoder_v0p0p1_0.x29.A VDD.t430 VDD.t429 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1579 frontAnalog_v0p0p1_8.RSfetsym_0.x1.Y frontAnalog_v0p0p1_8.x63.X VDD.t521 VDD.t519 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1580 resistorDivider_v0p0p1_0.V15.t1 resistorDivider_v0p0p1_0.V14.t2 GND.t26 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1581 a_53630_n30996# frontAnalog_v0p0p1_10.IB.t26 GND.t617 GND.t186 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1582 a_78241_n39305# 16to4_PriorityEncoder_v0p0p1_0.x5.x4.C a_78159_n39549# VDD.t716 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X1583 OUT0.t75 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND.t1120 GND.t1119 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1584 GND.t582 frontAnalog_v0p0p1_2.RSfetsym_0.QN.t5 a_59577_n3483# GND.t581 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1585 a_78525_n53555# 16to4_PriorityEncoder_v0p0p1_0.x3.x22.D GND.t692 GND.t691 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X1586 OUT0.t12 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD.t1072 VDD.t1071 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1587 GND.t289 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t75 GND.t288 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1588 16to4_PriorityEncoder_v0p0p1_0.x5.x22.D a_77605_n45765# VDD.t792 VDD.t791 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X1589 GND.t1246 frontAnalog_v0p0p1_3.RSfetsym_0.QN.t6 a_59577_n14283# GND.t1245 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1590 frontAnalog_v0p0p1_4.x65.X a_57123_n18759# GND.t750 GND.t749 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1591 GND.t223 16to4_PriorityEncoder_v0p0p1_0.I11.t12 a_59578_n24570# GND.t222 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1592 GND.t1279 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t74 GND.t1278 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1593 resistorDivider_v0p0p1_0.V7.t4 resistorDivider_v0p0p1_0.V6.t3 GND.t399 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1594 a_77605_n40069# 16to4_PriorityEncoder_v0p0p1_0.I13.t13 GND.t245 GND.t243 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1595 a_16719_n13117.t4 a_16599_n13205.t19 a_16541_n13117.t9 GND.t1499 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1596 frontAnalog_v0p0p1_12.x63.X a_57123_n74279# VDD.t24 VDD.t23 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1597 resistorDivider_v0p0p1_0.V6.t13 resistorDivider_v0p0p1_0.V5.t14 GND.t615 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1598 resistorDivider_v0p0p1_0.V1.t7 VL.t3 GND.t119 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1599 a_77881_n51585# 16to4_PriorityEncoder_v0p0p1_0.x3.x16.C a_77775_n51585# GND.t158 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X1600 16to4_PriorityEncoder_v0p0p1_0.x5.A2 a_78065_n41309# VDD.t1444 VDD.t100 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.148 ps=1.34 w=1 l=0.15
X1601 GND.t682 frontAnalog_v0p0p1_1.x65.X frontAnalog_v0p0p1_1.RSfetsym_0.x2.Y GND.t681 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1602 VIN.t26 w_55000_n62328# error sky130_fd_pr__cap_var_lvt w=2 l=0.18
X1603 OUT2.t11 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD.t919 VDD.t918 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1604 GND.t166 16to4_PriorityEncoder_v0p0p1_0.x3.x17.A a_78349_n51085# GND.t165 sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X1605 VDD.t1483 frontAnalog_v0p0p1_6.x65.A.t6 a_57123_n29559# VDD.t1482 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1606 16to4_PriorityEncoder_v0p0p1_0.x22.Y 16to4_PriorityEncoder_v0p0p1_0.x22.A GND.t1520 GND.t1519 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1607 16to4_PriorityEncoder_v0p0p1_0.x3.x4.C a_77605_n48109# VDD.t630 VDD.t629 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.148 ps=1.34 w=1 l=0.15
X1608 GND.t985 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t81 GND.t984 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1609 a_77725_n50381# 16to4_PriorityEncoder_v0p0p1_0.x3.EI a_77639_n50381# GND.t859 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X1610 VDD.t231 16to4_PriorityEncoder_v0p0p1_0.I13.t14 a_77637_n41087# VDD.t230 sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X1611 VDD.t845 frontAnalog_v0p0p1_4.x65.X frontAnalog_v0p0p1_4.RSfetsym_0.x2.Y VDD.t844 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1612 OUT1.t14 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD.t282 VDD.t281 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1613 resistorDivider_v0p0p1_0.V9.t5 resistorDivider_v0p0p1_0.V8.t8 GND.t119 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1614 VDD.t866 16to4_PriorityEncoder_v0p0p1_0.x3.x22.A a_78775_n53555# VDD.t865 sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X1615 OUT0.t11 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD.t1070 VDD.t1069 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1616 VDD.t458 frontAnalog_v0p0p1_9.x65.A.t6 a_57123_n51159# VDD.t457 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1617 GND.t110 frontAnalog_v0p0p1_8.x63.A.t7 a_57123_n47279# GND.t109 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X1618 VDD.t611 frontAnalog_v0p0p1_1.x65.X frontAnalog_v0p0p1_1.RSfetsym_0.x2.Y VDD.t610 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1619 frontAnalog_v0p0p1_0.RSfetsym_0.x2.Y frontAnalog_v0p0p1_0.x65.X VDD.t247 VDD.t245 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1620 frontAnalog_v0p0p1_6.x63.X a_57123_n31079# VDD.t545 VDD.t544 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1621 frontAnalog_v0p0p1_15.RSfetsym_0.x2.Y frontAnalog_v0p0p1_15.x65.X VDD.t1373 VDD.t1371 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1622 16to4_PriorityEncoder_v0p0p1_0.x42.A 16to4_PriorityEncoder_v0p0p1_0.x5.GS GND.t1560 GND.t743 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1623 16to4_PriorityEncoder_v0p0p1_0.x29.A 16to4_PriorityEncoder_v0p0p1_0.x28.A GND.t88 GND.t87 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1624 w_55000_n46750# VIN.t27 a_53630_n47196# GND.t421 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1625 frontAnalog_v0p0p1_13.RSfetsym_0.x2.Y frontAnalog_v0p0p1_13.x65.X GND.t136 GND.t135 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1626 OUT0.t74 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND.t1118 GND.t1117 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1627 16to4_PriorityEncoder_v0p0p1_0.x22.Y 16to4_PriorityEncoder_v0p0p1_0.x22.A VDD.t1453 VDD.t1452 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1628 a_78241_n47345# 16to4_PriorityEncoder_v0p0p1_0.x3.x4.C a_78159_n47589# VDD.t1200 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X1629 frontAnalog_v0p0p1_5.RSfetsym_0.QN.t1 frontAnalog_v0p0p1_5.x65.X VDD.t135 VDD.t134 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.25
X1630 frontAnalog_v0p0p1_11.x63.A.t2 frontAnalog_v0p0p1_11.x65.A.t7 a_55268_n63336# GND.t1096 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1631 OUT0.t73 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND.t1116 GND.t1115 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1632 GND.t1114 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t72 GND.t1113 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1633 GND.t1518 16to4_PriorityEncoder_v0p0p1_0.x22.A 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND.t1517 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1634 16to4_PriorityEncoder_v0p0p1_0.x3.x22.D a_77605_n53805# VDD.t509 VDD.t508 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X1635 a_77783_n48109# frontAnalog_v0p0p1_9.Q.t12 a_77687_n48109# VDD.t1342 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X1636 16to4_PriorityEncoder_v0p0p1_0.x1.A a_78349_n43045# GND.t1505 GND.t408 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.102 ps=0.99 w=0.65 l=0.15
X1637 frontAnalog_v0p0p1_11.Q.t3 frontAnalog_v0p0p1_11.RSfetsym_0.QN.t5 VDD.t536 VDD.t423 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.3
X1638 a_77605_n48109# frontAnalog_v0p0p1_10.Q.t13 GND.t1080 GND.t818 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1639 GND.t287 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t74 GND.t286 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1640 GND.t839 16to4_PriorityEncoder_v0p0p1_0.x5.x14.A a_78065_n41309# GND.t838 sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X1641 VDD.t280 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t13 VDD.t279 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1642 OUT1.t12 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD.t278 VDD.t277 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1643 a_59577_n68283# frontAnalog_v0p0p1_13.x63.X frontAnalog_v0p0p1_13.Q.t1 GND.t538 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1644 a_59578_n78570# frontAnalog_v0p0p1_14.x65.X frontAnalog_v0p0p1_14.RSfetsym_0.QN.t0 GND.t847 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.315 ps=2.72 w=1 l=0.15
X1645 GND.t983 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t80 GND.t982 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1646 VDD.t276 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t11 VDD.t275 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1647 frontAnalog_v0p0p1_8.Q.t4 frontAnalog_v0p0p1_8.RSfetsym_0.x2.Y GND.t651 GND.t226 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.25
X1648 frontAnalog_v0p0p1_8.x63.A.t3 frontAnalog_v0p0p1_8.x65.A.t5 VDD.t89 VDD.t88 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1649 16to4_PriorityEncoder_v0p0p1_0.x5.x18.C frontAnalog_v0p0p1_6.Q.t11 VDD.t879 VDD.t878 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1650 OUT0.t10 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD.t1068 VDD.t1067 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1651 OUT2.t79 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND.t981 GND.t980 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1652 frontAnalog_v0p0p1_4.x63.A.t0 frontAnalog_v0p0p1_4.x65.A.t7 a_55268_n20136# GND.t199 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1653 a_77759_n45765# 16to4_PriorityEncoder_v0p0p1_0.x5.x20.B a_77687_n45765# GND.t905 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X1654 VDD.t823 16to4_PriorityEncoder_v0p0p1_0.x5.A2 a_82988_n43855# VDD.t822 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X1655 frontAnalog_v0p0p1_1.x63.A.t3 CLK.t71 w_55000_n41350# VDD.t109 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1656 OUT0.t9 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD.t1066 VDD.t1065 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1657 VDD.t1064 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t8 VDD.t1063 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1658 VDD.t1451 16to4_PriorityEncoder_v0p0p1_0.x22.A 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD.t1450 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1659 VDD.t1384 frontAnalog_v0p0p1_10.x65.X frontAnalog_v0p0p1_10.RSfetsym_0.x2.Y VDD.t1383 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1660 a_78649_n39527# 16to4_PriorityEncoder_v0p0p1_0.x5.EO VDD.t833 VDD.t832 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X1661 GND.t1112 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t71 GND.t1111 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1662 16to4_PriorityEncoder_v0p0p1_0.x1.A a_78349_n43045# VDD.t1440 VDD.t1439 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.148 ps=1.34 w=1 l=0.15
X1663 VDD.t541 frontAnalog_v0p0p1_14.x63.A.t7 a_57123_n79679# VDD.t540 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1664 a_78349_n43045# 16to4_PriorityEncoder_v0p0p1_0.x5.x22.A GND.t590 GND.t252 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1665 a_59577_n25083# frontAnalog_v0p0p1_5.x63.X 16to4_PriorityEncoder_v0p0p1_0.I11.t0 GND.t645 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1666 a_59578_n35370# frontAnalog_v0p0p1_7.x65.X frontAnalog_v0p0p1_7.RSfetsym_0.QN.t3 GND.t1388 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.315 ps=2.72 w=1 l=0.15
X1667 VDD.t110 CLK.t72 w_55000_n83928# GND.t126 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1668 frontAnalog_v0p0p1_11.Q.t1 frontAnalog_v0p0p1_11.x63.X VDD.t93 VDD.t92 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.25
X1669 a_53630_n74196# frontAnalog_v0p0p1_10.IB.t27 GND.t618 GND.t186 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1670 a_78775_n45515# 16to4_PriorityEncoder_v0p0p1_0.x5.x22.B a_78703_n45515# VDD.t839 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X1671 VDD.t1188 frontAnalog_v0p0p1_13.x63.A.t7 frontAnalog_v0p0p1_13.x65.A.t3 VDD.t13 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1672 VDD.t274 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t10 VDD.t273 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1673 OUT1.t9 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD.t272 VDD.t271 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1674 GND.t1110 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t70 GND.t1109 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1675 OUT3.t73 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND.t1277 GND.t1276 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1676 OUT2.t78 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND.t979 GND.t978 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1677 VDD.t111 CLK.t73 w_55000_n19128# GND.t127 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1678 frontAnalog_v0p0p1_15.x65.X a_57123_n83559# GND.t162 GND.t161 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1679 frontAnalog_v0p0p1_4.RSfetsym_0.QN.t3 frontAnalog_v0p0p1_4.RSfetsym_0.x1.Y GND.t1491 GND.t550 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.25
X1680 16to4_PriorityEncoder_v0p0p1_0.x43.A 16to4_PriorityEncoder_v0p0p1_0.x42.A GND.t744 GND.t743 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1681 VDD.t622 frontAnalog_v0p0p1_3.x65.X frontAnalog_v0p0p1_3.RSfetsym_0.x2.Y VDD.t621 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1682 resistorDivider_v0p0p1_0.V15.t7 resistorDivider_v0p0p1_0.V14.t6 GND.t60 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1683 OUT3.t5 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD.t1214 VDD.t1213 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1684 VDD.t1494 frontAnalog_v0p0p1_0.x63.X 16to4_PriorityEncoder_v0p0p1_0.I14.t2 VDD.t1493 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.25
X1685 VDD.t664 frontAnalog_v0p0p1_7.x63.A.t6 a_57123_n36479# VDD.t663 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1686 a_53630_n79596# resistorDivider_v0p0p1_0.V2.t17 w_55000_n78528# GND.t613 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1687 VDD.t112 CLK.t74 w_55000_n40728# GND.t128 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1688 16to4_PriorityEncoder_v0p0p1_0.I12.t0 frontAnalog_v0p0p1_4.x63.X VDD.t56 VDD.t55 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.25
X1689 VFS.t1 resistorDivider_v0p0p1_0.V16.t4 GND.t211 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1690 VDD.t917 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t10 VDD.t916 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1691 VDD.t1062 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t7 VDD.t1061 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1692 a_77687_n53805# frontAnalog_v0p0p1_10.Q.t14 a_77605_n53805# GND.t1081 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X1693 VDD.t408 frontAnalog_v0p0p1_5.x63.A.t7 frontAnalog_v0p0p1_5.x65.A.t1 VDD.t15 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1694 resistorDivider_v0p0p1_0.V4.t0 resistorDivider_v0p0p1_0.V3.t0 GND.t59 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1695 frontAnalog_v0p0p1_9.RSfetsym_0.x2.Y frontAnalog_v0p0p1_9.x65.X GND.t713 GND.t712 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1696 a_55268_n57936# CLK.t75 GND.t130 GND.t129 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1697 VDD.t1372 frontAnalog_v0p0p1_15.x65.X frontAnalog_v0p0p1_15.RSfetsym_0.x2.Y VDD.t1371 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1698 VDD.t113 CLK.t76 w_55000_n41350# GND.t11 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1699 frontAnalog_v0p0p1_6.x65.A.t3 frontAnalog_v0p0p1_6.x63.A.t7 a_55268_n30936# GND.t1419 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1700 frontAnalog_v0p0p1_11.RSfetsym_0.QN.t4 frontAnalog_v0p0p1_11.Q.t12 VDD.t424 VDD.t423 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.3
X1701 VDD.t1060 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t6 VDD.t1059 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1702 GND.t1460 16to4_PriorityEncoder_v0p0p1_0.x36.A 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND.t1459 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1703 frontAnalog_v0p0p1_1.x65.X a_57123_n40359# GND.t440 GND.t439 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1704 VDD.t36 16to4_PriorityEncoder_v0p0p1_0.I12.t11 a_77637_n40777# VDD.t35 sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X1705 16to4_PriorityEncoder_v0p0p1_0.x22.A 16to4_PriorityEncoder_v0p0p1_0.x21.A GND.t606 GND.t605 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1706 a_78649_n47567# 16to4_PriorityEncoder_v0p0p1_0.x3.EO VDD.t1038 VDD.t1037 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X1707 a_53630_n36396# resistorDivider_v0p0p1_0.V10.t17 w_55000_n35328# GND.t405 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1708 16to4_PriorityEncoder_v0p0p1_0.x3.A1 a_78349_n51085# VDD.t821 VDD.t820 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.148 ps=1.34 w=1 l=0.15
X1709 GND.t742 16to4_PriorityEncoder_v0p0p1_0.x42.A 16to4_PriorityEncoder_v0p0p1_0.x43.A GND.t741 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1710 OUT2.t77 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND.t977 GND.t976 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1711 16to4_PriorityEncoder_v0p0p1_0.x3.x22.A a_77639_n50381# VDD.t1382 VDD.t1381 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.167 ps=1.39 w=1 l=0.15
X1712 a_78775_n53555# 16to4_PriorityEncoder_v0p0p1_0.x3.x22.B a_78703_n53555# VDD.t385 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X1713 frontAnalog_v0p0p1_11.RSfetsym_0.x2.Y frontAnalog_v0p0p1_11.x65.X VDD.t887 VDD.t885 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1714 frontAnalog_v0p0p1_2.RSfetsym_0.x1.Y frontAnalog_v0p0p1_2.x63.X VDD.t1363 VDD.t1361 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1715 resistorDivider_v0p0p1_0.V11.t6 resistorDivider_v0p0p1_0.V10.t6 GND.t26 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1716 a_55268_n14736# CLK.t77 GND.t523 GND.t522 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1717 frontAnalog_v0p0p1_11.RSfetsym_0.x1.Y frontAnalog_v0p0p1_11.x63.X GND.t115 GND.t113 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1718 frontAnalog_v0p0p1_13.RSfetsym_0.QN.t0 frontAnalog_v0p0p1_13.x65.X VDD.t127 VDD.t126 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.25
X1719 OUT2.t76 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND.t975 GND.t974 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1720 VDD.t1212 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t4 VDD.t1211 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1721 OUT1.t8 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD.t270 VDD.t269 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1722 GND.t1275 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t72 GND.t1274 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1723 GND.t973 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t75 GND.t972 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1724 VDD.t784 frontAnalog_v0p0p1_14.x65.X frontAnalog_v0p0p1_14.RSfetsym_0.QN.t1 VDD.t783 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.25
X1725 OUT3.t3 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD.t1210 VDD.t1209 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1726 GND.t1108 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t69 GND.t1107 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1727 a_77637_n49127# 16to4_PriorityEncoder_v0p0p1_0.x3.EI VDD.t799 VDD.t546 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X1728 frontAnalog_v0p0p1_0.x65.A.t1 CLK.t78 frontAnalog_v0p0p1_0.x63.A.t1 VDD.t481 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1729 resistorDivider_v0p0p1_0.V7.t9 resistorDivider_v0p0p1_0.V6.t5 GND.t102 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1730 VDD.t1208 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t2 VDD.t1207 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1731 16to4_PriorityEncoder_v0p0p1_0.x22.A 16to4_PriorityEncoder_v0p0p1_0.x21.A VDD.t565 VDD.t564 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1732 frontAnalog_v0p0p1_12.RSfetsym_0.x1.Y frontAnalog_v0p0p1_12.x63.X VDD.t589 VDD.t585 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1733 GND.t143 frontAnalog_v0p0p1_5.x65.X frontAnalog_v0p0p1_5.RSfetsym_0.x2.Y GND.t142 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1734 a_77687_n48109# frontAnalog_v0p0p1_8.Q.t8 a_77605_n48109# VDD.t737 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X1735 GND.t634 frontAnalog_v0p0p1_14.x63.X frontAnalog_v0p0p1_14.RSfetsym_0.x1.Y GND.t633 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1736 VIN.t28 w_55000_n46128# error sky130_fd_pr__cap_var_lvt w=2 l=0.18
X1737 GND.t971 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t74 GND.t970 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1738 OUT2.t9 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD.t915 VDD.t914 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1739 frontAnalog_v0p0p1_2.x65.X a_57123_n2559# VDD.t209 VDD.t208 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1740 a_16719_n13117.t3 a_16599_n13205.t20 a_16541_n13117.t8 GND.t1500 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1741 a_53630_n84996# frontAnalog_v0p0p1_10.IB.t28 GND.t619 GND.t186 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1742 VDD.t1332 frontAnalog_v0p0p1_7.x65.X frontAnalog_v0p0p1_7.RSfetsym_0.QN.t1 VDD.t1331 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.25
X1743 a_16719_n13117.t2 a_16599_n13205.t21 a_16541_n13117.t7 GND.t1501 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1744 OUT1.t73 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND.t285 GND.t284 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1745 VDD.t913 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t8 VDD.t912 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1746 VDD.t1058 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t5 VDD.t1057 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1747 16to4_PriorityEncoder_v0p0p1_0.x3.x14.B a_77637_n49127# VDD.t750 VDD.t386 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.167 ps=1.39 w=1 l=0.15
X1748 frontAnalog_v0p0p1_6.RSfetsym_0.x1.Y frontAnalog_v0p0p1_6.x63.X VDD.t43 VDD.t39 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1749 GND.t283 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t72 GND.t282 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1750 frontAnalog_v0p0p1_8.x65.A.t2 CLK.t79 frontAnalog_v0p0p1_8.x63.A.t0 VDD.t482 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1751 a_77605_n43545# 16to4_PriorityEncoder_v0p0p1_0.x5.x16.C VDD.t503 VDD.t145 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X1752 frontAnalog_v0p0p1_3.x63.X a_57123_n14879# VDD.t1380 VDD.t1379 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1753 frontAnalog_v0p0p1_13.RSfetsym_0.x2.Y frontAnalog_v0p0p1_13.x65.X VDD.t125 VDD.t123 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1754 frontAnalog_v0p0p1_0.RSfetsym_0.x1.Y frontAnalog_v0p0p1_0.x63.X VDD.t1492 VDD.t1490 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1755 a_53630_n20196# frontAnalog_v0p0p1_10.IB.t29 GND.t620 GND.t186 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1756 w_55000_n30550# VIN.t29 a_53630_n30996# GND.t490 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1757 GND.t811 frontAnalog_v0p0p1_7.x63.X frontAnalog_v0p0p1_7.RSfetsym_0.x1.Y GND.t810 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1758 VDD.t48 16to4_PriorityEncoder_v0p0p1_0.x35.A 16to4_PriorityEncoder_v0p0p1_0.x36.A VDD.t47 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1759 GND.t1273 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t71 GND.t1272 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1760 GND.t1088 frontAnalog_v0p0p1_0.x63.A.t6 a_57123_n9479# GND.t794 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X1761 frontAnalog_v0p0p1_12.x65.X a_57123_n72759# VDD.t875 VDD.t874 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1762 frontAnalog_v0p0p1_13.x63.X a_57123_n68879# GND.t855 GND.t854 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1763 GND.t1458 16to4_PriorityEncoder_v0p0p1_0.x36.A 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND.t1457 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1764 a_53630_n9396# resistorDivider_v0p0p1_0.V15.t17 w_55000_n8328# GND.t558 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1765 a_53630_n41796# frontAnalog_v0p0p1_10.IB.t30 GND.t187 GND.t186 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1766 frontAnalog_v0p0p1_11.x63.A.t0 CLK.t80 w_55000_n62950# VDD.t0 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1767 16to4_PriorityEncoder_v0p0p1_0.x5.x4.B a_77605_n39305# GND.t556 GND.t555 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.102 ps=0.99 w=0.65 l=0.15
X1768 resistorDivider_v0p0p1_0.V14.t15 resistorDivider_v0p0p1_0.V13.t15 GND.t26 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1769 GND.t577 frontAnalog_v0p0p1_8.x65.A.t6 a_57123_n45759# GND.t109 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X1770 resistorDivider_v0p0p1_0.V5.t4 resistorDivider_v0p0p1_0.V4.t6 GND.t75 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1771 OUT3.t70 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND.t1271 GND.t1270 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1772 frontAnalog_v0p0p1_15.RSfetsym_0.QN.t1 frontAnalog_v0p0p1_15.RSfetsym_0.x1.Y GND.t915 GND.t914 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.25
X1773 OUT2.t7 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD.t911 VDD.t910 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1774 VDD.t909 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t6 VDD.t908 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1775 GND.t711 frontAnalog_v0p0p1_9.x65.X frontAnalog_v0p0p1_9.RSfetsym_0.x2.Y GND.t710 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1776 GND.t758 16to4_PriorityEncoder_v0p0p1_0.x43.A 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND.t757 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1777 frontAnalog_v0p0p1_8.Q.t0 frontAnalog_v0p0p1_8.RSfetsym_0.QN.t6 VDD.t710 VDD.t709 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.3
X1778 frontAnalog_v0p0p1_5.RSfetsym_0.x2.Y frontAnalog_v0p0p1_5.x65.X VDD.t133 VDD.t131 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1779 VDD.t483 CLK.t81 w_55000_n84550# GND.t524 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1780 VDD.t520 frontAnalog_v0p0p1_8.x63.X frontAnalog_v0p0p1_8.RSfetsym_0.x1.Y VDD.t519 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1781 VDD.t588 frontAnalog_v0p0p1_12.x63.X frontAnalog_v0p0p1_12.Q.t2 VDD.t587 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.25
X1782 w_55000_n73128# CLK.t82 frontAnalog_v0p0p1_12.x65.A.t0 VDD.t484 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1783 frontAnalog_v0p0p1_5.x63.X a_57123_n25679# GND.t411 GND.t410 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1784 GND.t502 frontAnalog_v0p0p1_10.IB.t0 frontAnalog_v0p0p1_10.IB.t1 GND.t501 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1785 resistorDivider_v0p0p1_0.V8.t17 w_55000_n46750# error sky130_fd_pr__cap_var_lvt w=2 l=0.18
X1786 GND.t969 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t73 GND.t968 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1787 frontAnalog_v0p0p1_1.RSfetsym_0.QN.t0 frontAnalog_v0p0p1_1.RSfetsym_0.x1.Y GND.t624 GND.t623 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.25
X1788 16to4_PriorityEncoder_v0p0p1_0.x5.x4.B a_77605_n39305# VDD.t511 VDD.t510 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.148 ps=1.34 w=1 l=0.15
X1789 OUT3.t69 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND.t1269 GND.t1268 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1790 16to4_PriorityEncoder_v0p0p1_0.x2.A a_78525_n45515# GND.t678 GND.t677 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.102 ps=0.99 w=0.65 l=0.15
X1791 16to4_PriorityEncoder_v0p0p1_0.x36.Y 16to4_PriorityEncoder_v0p0p1_0.x36.A GND.t1456 GND.t1455 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1792 VDD.t1206 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t1 VDD.t1205 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1793 GND.t114 frontAnalog_v0p0p1_11.x63.X frontAnalog_v0p0p1_11.RSfetsym_0.x1.Y GND.t113 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1794 GND.t281 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t71 GND.t280 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1795 16to4_PriorityEncoder_v0p0p1_0.x36.Y 16to4_PriorityEncoder_v0p0p1_0.x36.A VDD.t1403 VDD.t1402 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1796 VDD.t42 frontAnalog_v0p0p1_6.x63.X frontAnalog_v0p0p1_6.Q.t1 VDD.t41 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.25
X1797 a_77605_n51585# 16to4_PriorityEncoder_v0p0p1_0.x3.x16.C VDD.t149 VDD.t148 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X1798 w_55000_n29928# CLK.t83 frontAnalog_v0p0p1_6.x65.A.t0 VDD.t234 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1799 frontAnalog_v0p0p1_4.RSfetsym_0.x1.Y frontAnalog_v0p0p1_4.x63.X GND.t78 GND.t76 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1800 a_53630_n57996# frontAnalog_v0p0p1_10.IB.t31 GND.t188 GND.t186 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1801 a_55268_n79536# CLK.t84 GND.t123 GND.t122 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1802 frontAnalog_v0p0p1_9.x65.A.t0 frontAnalog_v0p0p1_9.x63.A.t6 a_55268_n52536# GND.t1399 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1803 16to4_PriorityEncoder_v0p0p1_0.x43.Y 16to4_PriorityEncoder_v0p0p1_0.x43.A GND.t756 GND.t755 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1804 16to4_PriorityEncoder_v0p0p1_0.x3.x4.B a_77605_n47345# GND.t508 GND.t507 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.102 ps=0.99 w=0.65 l=0.15
X1805 resistorDivider_v0p0p1_0.V11.t11 resistorDivider_v0p0p1_0.V10.t8 GND.t60 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1806 VDD.t586 frontAnalog_v0p0p1_12.x63.X frontAnalog_v0p0p1_12.RSfetsym_0.x1.Y VDD.t585 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1807 GND.t279 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t70 GND.t278 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1808 frontAnalog_v0p0p1_0.RSfetsym_0.QN.t4 frontAnalog_v0p0p1_0.RSfetsym_0.x1.Y GND.t720 GND.t719 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.25
X1809 VDD.t246 frontAnalog_v0p0p1_0.x65.X frontAnalog_v0p0p1_0.RSfetsym_0.x2.Y VDD.t245 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1810 16to4_PriorityEncoder_v0p0p1_0.x3.x17.D a_77605_n51585# GND.t488 GND.t487 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.196 ps=1.33 w=0.65 l=0.15
X1811 GND.t1267 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t68 GND.t1266 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1812 GND.t795 frontAnalog_v0p0p1_0.x65.A.t6 a_57123_n7959# GND.t794 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X1813 GND.t580 frontAnalog_v0p0p1_11.RSfetsym_0.QN.t6 a_59577_n62883# GND.t579 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1814 GND.t134 frontAnalog_v0p0p1_13.x65.X frontAnalog_v0p0p1_13.RSfetsym_0.x2.Y GND.t133 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1815 resistorDivider_v0p0p1_0.V6.t1 resistorDivider_v0p0p1_0.V5.t2 GND.t211 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1816 16to4_PriorityEncoder_v0p0p1_0.x2.A a_78525_n45515# VDD.t607 VDD.t606 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.148 ps=1.34 w=1 l=0.15
X1817 OUT2.t5 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD.t907 VDD.t906 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1818 a_78525_n45515# 16to4_PriorityEncoder_v0p0p1_0.x5.x22.B GND.t893 GND.t892 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1819 VDD.t1045 frontAnalog_v0p0p1_0.x63.A.t7 frontAnalog_v0p0p1_0.x65.A.t2 VDD.t719 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1820 16to4_PriorityEncoder_v0p0p1_0.x5.x22.B a_78097_n45737# GND.t842 GND.t841 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.112 ps=1.04 w=0.65 l=0.15
X1821 VDD.t1401 16to4_PriorityEncoder_v0p0p1_0.x36.A 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD.t1400 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1822 a_53630_n14796# frontAnalog_v0p0p1_10.IB.t32 GND.t189 GND.t186 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1823 a_77637_n48817# 16to4_PriorityEncoder_v0p0p1_0.x3.EI VDD.t798 VDD.t797 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X1824 16to4_PriorityEncoder_v0p0p1_0.x5.x19.C 16to4_PriorityEncoder_v0p0p1_0.I12.t12 VDD.t825 VDD.t824 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1825 frontAnalog_v0p0p1_9.RSfetsym_0.x1.Y frontAnalog_v0p0p1_9.x63.X VDD.t192 VDD.t191 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1826 VDD.t740 frontAnalog_v0p0p1_14.x65.A.t7 a_57123_n78159# VDD.t739 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1827 VDD.t65 16to4_PriorityEncoder_v0p0p1_0.x28.A 16to4_PriorityEncoder_v0p0p1_0.x29.A VDD.t64 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1828 VDD.t40 frontAnalog_v0p0p1_6.x63.X frontAnalog_v0p0p1_6.RSfetsym_0.x1.Y VDD.t39 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1829 OUT0.t68 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND.t1106 GND.t1105 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1830 OUT2.t72 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND.t967 GND.t966 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1831 16to4_PriorityEncoder_v0p0p1_0.I15.t0 frontAnalog_v0p0p1_2.RSfetsym_0.QN.t6 VDD.t537 VDD.t388 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.3
X1832 VDD.t124 frontAnalog_v0p0p1_13.x65.X frontAnalog_v0p0p1_13.RSfetsym_0.x2.Y VDD.t123 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1833 VDD.t1491 frontAnalog_v0p0p1_0.x63.X frontAnalog_v0p0p1_0.RSfetsym_0.x1.Y VDD.t1490 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1834 frontAnalog_v0p0p1_10.x63.X a_57123_n58079# VDD.t461 VDD.t460 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1835 16to4_PriorityEncoder_v0p0p1_0.x3.x4.B a_77605_n47345# VDD.t469 VDD.t468 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.148 ps=1.34 w=1 l=0.15
X1836 GND.t1265 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t67 GND.t1264 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1837 GND.t1104 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t67 GND.t1103 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1838 OUT1.t69 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND.t277 GND.t276 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1839 a_77775_n43545# 16to4_PriorityEncoder_v0p0p1_0.x5.x19.C a_77687_n43545# GND.t153 sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
X1840 16to4_PriorityEncoder_v0p0p1_0.x43.A 16to4_PriorityEncoder_v0p0p1_0.x42.A VDD.t656 VDD.t655 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1841 OUT1.t7 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD.t268 VDD.t267 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1842 frontAnalog_v0p0p1_2.RSfetsym_0.x2.Y frontAnalog_v0p0p1_2.x65.X GND.t724 GND.t723 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1843 VDD.t905 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t4 VDD.t904 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1844 VDD.t755 VDD.t753 a_77605_n45765# VDD.t754 sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X1845 16to4_PriorityEncoder_v0p0p1_0.x5.x22.B a_78097_n45737# VDD.t752 VDD.t751 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.167 ps=1.39 w=1 l=0.15
X1846 VDD.t1448 frontAnalog_v0p0p1_7.x65.A.t7 a_57123_n34959# VDD.t1447 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1847 VDD.t132 frontAnalog_v0p0p1_5.x65.X frontAnalog_v0p0p1_5.RSfetsym_0.x2.Y VDD.t131 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1848 resistorDivider_v0p0p1_0.V16.t0 resistorDivider_v0p0p1_0.V15.t4 GND.t84 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1849 resistorDivider_v0p0p1_0.V5.t12 resistorDivider_v0p0p1_0.V4.t15 GND.t119 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1850 OUT2.t71 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND.t965 GND.t964 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1851 OUT0.t4 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD.t1056 VDD.t1055 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1852 16to4_PriorityEncoder_v0p0p1_0.x3.A0 a_78525_n53555# VDD.t1431 VDD.t1430 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.148 ps=1.34 w=1 l=0.15
X1853 GND.t963 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t70 GND.t962 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1854 a_78431_n43045# 16to4_PriorityEncoder_v0p0p1_0.x5.x17.D a_78349_n43045# VDD.t464 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X1855 resistorDivider_v0p0p1_0.V14.t0 resistorDivider_v0p0p1_0.V13.t0 GND.t60 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1856 GND.t671 VDD.t1511 a_77759_n45765# GND.t670 sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X1857 VDD.t903 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t3 VDD.t902 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1858 a_78525_n53555# 16to4_PriorityEncoder_v0p0p1_0.x3.x22.B GND.t398 GND.t397 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1859 VDD.t1054 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t3 VDD.t1053 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1860 a_77687_n52819# 16to4_PriorityEncoder_v0p0p1_0.x3.EI a_77605_n52819# GND.t532 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.109 ps=1.36 w=0.42 l=0.15
X1861 w_55000_n52150# VIN.t30 a_53630_n52596# GND.t210 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1862 frontAnalog_v0p0p1_12.RSfetsym_0.x2.Y frontAnalog_v0p0p1_12.x65.X GND.t94 GND.t93 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1863 frontAnalog_v0p0p1_0.RSfetsym_0.QN.t2 frontAnalog_v0p0p1_0.x65.X VDD.t244 VDD.t243 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.25
X1864 GND.t494 16to4_PriorityEncoder_v0p0p1_0.x5.x9.Y a_78159_n39549# GND.t493 sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X1865 frontAnalog_v0p0p1_2.x63.A.t1 frontAnalog_v0p0p1_2.x65.A.t7 VDD.t29 VDD.t28 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1866 VDD.t102 CLK.t85 w_55000_n2928# GND.t124 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1867 frontAnalog_v0p0p1_8.x63.A.t2 frontAnalog_v0p0p1_8.x65.A.t7 a_55268_n47136# GND.t578 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1868 resistorDivider_v0p0p1_0.V12.t14 resistorDivider_v0p0p1_0.V11.t14 GND.t212 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1869 GND.t1102 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t66 GND.t1101 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1870 a_77775_n51585# 16to4_PriorityEncoder_v0p0p1_0.x3.x19.C a_77687_n51585# GND.t158 sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
X1871 16to4_PriorityEncoder_v0p0p1_0.x5.x14.A a_77637_n40777# GND.t230 GND.t120 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.112 ps=1.04 w=0.65 l=0.15
X1872 VDD.t901 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t2 VDD.t900 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1873 frontAnalog_v0p0p1_6.RSfetsym_0.x2.Y frontAnalog_v0p0p1_6.x65.X GND.t514 GND.t513 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1874 frontAnalog_v0p0p1_15.RSfetsym_0.x1.Y frontAnalog_v0p0p1_15.x63.X GND.t909 GND.t908 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1875 OUT1.t6 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD.t266 VDD.t265 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1876 a_59577_n8883# frontAnalog_v0p0p1_0.x63.X 16to4_PriorityEncoder_v0p0p1_0.I14.t4 GND.t1554 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1877 frontAnalog_v0p0p1_3.RSfetsym_0.x1.Y frontAnalog_v0p0p1_3.x63.X VDD.t224 VDD.t220 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1878 w_55000_n8328# CLK.t86 frontAnalog_v0p0p1_0.x65.A.t0 VDD.t103 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1879 a_59577_n73683# frontAnalog_v0p0p1_12.x63.X frontAnalog_v0p0p1_12.Q.t1 GND.t639 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1880 a_59578_n83970# frontAnalog_v0p0p1_15.x65.X frontAnalog_v0p0p1_15.RSfetsym_0.QN.t4 GND.t1420 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.315 ps=2.72 w=1 l=0.15
X1881 VDD.t796 16to4_PriorityEncoder_v0p0p1_0.x3.EI a_77605_n53805# VDD.t795 sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X1882 16to4_PriorityEncoder_v0p0p1_0.x3.x22.B a_78097_n53777# VDD.t22 VDD.t21 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.167 ps=1.39 w=1 l=0.15
X1883 OUT2.t1 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD.t899 VDD.t898 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1884 frontAnalog_v0p0p1_9.Q.t4 frontAnalog_v0p0p1_9.RSfetsym_0.x2.Y GND.t937 GND.t936 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.25
X1885 GND.t415 16to4_PriorityEncoder_v0p0p1_0.x1.A a_82906_n47995# GND.t414 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X1886 frontAnalog_v0p0p1_2.RSfetsym_0.QN.t1 16to4_PriorityEncoder_v0p0p1_0.I15.t8 VDD.t389 VDD.t388 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.3
X1887 GND.t1100 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t65 GND.t1099 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1888 resistorDivider_v0p0p1_0.V12.t7 resistorDivider_v0p0p1_0.V11.t8 GND.t693 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1889 resistorDivider_v0p0p1_0.V8.t6 resistorDivider_v0p0p1_0.V7.t8 GND.t75 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1890 resistorDivider_v0p0p1_0.V15.t8 resistorDivider_v0p0p1_0.V14.t9 GND.t59 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1891 GND.t1263 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t66 GND.t1262 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1892 a_78183_n45737# VDD.t1512 a_78097_n45737# GND.t672 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X1893 VDD.t104 CLK.t87 w_55000_n67728# GND.t104 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1894 a_59578_n19170# frontAnalog_v0p0p1_4.x65.X frontAnalog_v0p0p1_4.RSfetsym_0.QN.t0 GND.t895 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.315 ps=2.72 w=1 l=0.15
X1895 VDD.t1052 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t2 VDD.t1051 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1896 a_77881_n51335# 16to4_PriorityEncoder_v0p0p1_0.x3.x16.C a_77775_n51335# GND.t157 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X1897 frontAnalog_v0p0p1_8.Q.t1 frontAnalog_v0p0p1_8.x63.X VDD.t518 VDD.t517 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.25
X1898 VDD.t886 frontAnalog_v0p0p1_11.x65.X frontAnalog_v0p0p1_11.RSfetsym_0.x2.Y VDD.t885 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1899 a_78431_n51085# 16to4_PriorityEncoder_v0p0p1_0.x3.x17.D a_78349_n51085# VDD.t1339 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X1900 VDD.t1362 frontAnalog_v0p0p1_2.x63.X frontAnalog_v0p0p1_2.RSfetsym_0.x1.Y VDD.t1361 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1901 OUT2.t69 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND.t961 GND.t960 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1902 frontAnalog_v0p0p1_1.RSfetsym_0.x1.Y frontAnalog_v0p0p1_1.x63.X GND.t174 GND.t173 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1903 frontAnalog_v0p0p1_14.RSfetsym_0.x2.Y frontAnalog_v0p0p1_14.x65.X GND.t846 GND.t845 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1904 OUT1.t5 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD.t264 VDD.t263 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1905 16to4_PriorityEncoder_v0p0p1_0.x36.Y 16to4_PriorityEncoder_v0p0p1_0.x36.A VDD.t1399 VDD.t1398 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1906 a_59577_n30483# frontAnalog_v0p0p1_6.x63.X frontAnalog_v0p0p1_6.Q.t0 GND.t39 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1907 a_59578_n40770# frontAnalog_v0p0p1_1.x65.X frontAnalog_v0p0p1_1.RSfetsym_0.QN.t1 GND.t680 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.315 ps=2.72 w=1 l=0.15
X1908 VDD.t105 CLK.t88 w_55000_n68350# GND.t125 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1909 GND.t533 16to4_PriorityEncoder_v0p0p1_0.x3.x20.B a_77881_n52819# GND.t532 sky130_fd_pr__nfet_01v8 ad=0.196 pd=1.33 as=0.0693 ps=0.75 w=0.42 l=0.15
X1910 VDD.t749 16to4_PriorityEncoder_v0p0p1_0.x5.x14.A a_78315_n41309# VDD.t556 sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X1911 GND.t208 16to4_PriorityEncoder_v0p0p1_0.x3.x9.Y a_78159_n47589# GND.t207 sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X1912 GND.t959 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t68 GND.t958 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1913 VDD.t183 frontAnalog_v0p0p1_12.x63.A.t7 frontAnalog_v0p0p1_12.x65.A.t3 VDD.t117 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1914 frontAnalog_v0p0p1_2.x63.A.t3 CLK.t89 w_55000_n3550# VDD.t106 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1915 frontAnalog_v0p0p1_13.x65.X a_57123_n67359# GND.t1487 GND.t854 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1916 GND.t923 frontAnalog_v0p0p1_12.Q.t12 a_59578_n73170# GND.t922 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1917 resistorDivider_v0p0p1_0.V16.t12 resistorDivider_v0p0p1_0.V15.t12 GND.t399 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1918 VDD.t1050 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t1 VDD.t1049 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1919 16to4_PriorityEncoder_v0p0p1_0.I15.t2 frontAnalog_v0p0p1_2.x63.X VDD.t1360 VDD.t1359 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.25
X1920 GND.t722 frontAnalog_v0p0p1_2.x65.X frontAnalog_v0p0p1_2.RSfetsym_0.x2.Y GND.t721 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1921 VDD.t107 CLK.t90 w_55000_n24528# GND.t107 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1922 OUT0.t64 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND.t1098 GND.t1097 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1923 GND.t275 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t68 GND.t274 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1924 16to4_PriorityEncoder_v0p0p1_0.x29.Y 16to4_PriorityEncoder_v0p0p1_0.x29.A VDD.t428 VDD.t427 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1925 frontAnalog_v0p0p1_7.RSfetsym_0.x2.Y frontAnalog_v0p0p1_7.x65.X GND.t1387 GND.t1386 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1926 VDD.t91 frontAnalog_v0p0p1_1.x63.A.t7 a_57123_n41879# VDD.t90 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1927 GND.t1454 16to4_PriorityEncoder_v0p0p1_0.x36.A 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND.t1453 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1928 VDD.t223 frontAnalog_v0p0p1_3.x63.X 16to4_PriorityEncoder_v0p0p1_0.I13.t0 VDD.t222 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.25
X1929 VDD.t470 CLK.t91 w_55000_n25150# GND.t509 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1930 16to4_PriorityEncoder_v0p0p1_0.x3.A2 a_78065_n49349# GND.t401 GND.t400 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.102 ps=0.99 w=0.65 l=0.15
X1931 w_55000_n13728# CLK.t92 frontAnalog_v0p0p1_3.x65.A.t1 VDD.t471 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1932 frontAnalog_v0p0p1_8.RSfetsym_0.QN.t4 frontAnalog_v0p0p1_8.Q.t9 VDD.t715 VDD.t709 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.3
X1933 GND.t957 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t67 GND.t956 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1934 frontAnalog_v0p0p1_5.x65.X a_57123_n24159# GND.t602 GND.t410 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1935 GND.t403 16to4_PriorityEncoder_v0p0p1_0.I15.t9 a_77725_n42341# GND.t402 sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X1936 frontAnalog_v0p0p1_7.x65.A.t3 frontAnalog_v0p0p1_7.x63.A.t7 a_55268_n36336# GND.t657 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1937 a_53630_n20196# resistorDivider_v0p0p1_0.V13.t17 w_55000_n19128# GND.t69 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1938 a_78183_n53777# 16to4_PriorityEncoder_v0p0p1_0.x3.EI a_78097_n53777# GND.t858 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X1939 OUT2.t0 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD.t897 VDD.t896 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1940 OUT0.t0 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD.t1048 VDD.t1047 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1941 frontAnalog_v0p0p1_8.RSfetsym_0.x2.Y frontAnalog_v0p0p1_8.x65.X VDD.t5 VDD.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1942 OUT1.t4 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD.t262 VDD.t261 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1943 frontAnalog_v0p0p1_8.RSfetsym_0.x1.Y frontAnalog_v0p0p1_8.x63.X GND.t563 GND.t562 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1944 16to4_PriorityEncoder_v0p0p1_0.x35.A 16to4_PriorityEncoder_v0p0p1_0.x34.A VDD.t397 VDD.t396 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1945 GND.t754 16to4_PriorityEncoder_v0p0p1_0.x43.A 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND.t753 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1946 GND.t955 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t66 GND.t954 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1947 VDD.t142 16to4_PriorityEncoder_v0p0p1_0.x5.x19.C a_77605_n43295# VDD.t141 sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X1948 frontAnalog_v0p0p1_0.x63.A.t2 frontAnalog_v0p0p1_0.x65.A.t7 a_55268_n9336# GND.t796 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1949 OUT1.t3 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD.t260 VDD.t259 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1950 VDD.t258 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t2 VDD.t257 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1951 VDD.t426 16to4_PriorityEncoder_v0p0p1_0.x29.A 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD.t425 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1952 GND.t1430 16to4_PriorityEncoder_v0p0p1_0.I15.t10 a_59578_n2970# GND.t1429 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1953 GND.t1400 frontAnalog_v0p0p1_9.x63.A.t7 a_57123_n52679# GND.t482 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X1954 a_55268_n20136# CLK.t93 GND.t511 GND.t510 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1955 frontAnalog_v0p0p1_12.RSfetsym_0.QN.t0 frontAnalog_v0p0p1_12.x65.X VDD.t73 VDD.t72 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.25
X1956 16to4_PriorityEncoder_v0p0p1_0.x36.Y 16to4_PriorityEncoder_v0p0p1_0.x36.A GND.t1452 GND.t1451 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1957 a_16719_n13117.t1 a_16599_n13205.t22 a_16541_n13117.t6 GND.t1494 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1958 VDD.t1204 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t0 VDD.t1203 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1959 16to4_PriorityEncoder_v0p0p1_0.x3.x9.Y 16to4_PriorityEncoder_v0p0p1_0.x3.EI GND.t857 GND.t856 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1960 VDD.t221 frontAnalog_v0p0p1_3.x63.X frontAnalog_v0p0p1_3.RSfetsym_0.x1.Y VDD.t220 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1961 frontAnalog_v0p0p1_10.RSfetsym_0.x1.Y frontAnalog_v0p0p1_10.x63.X VDD.t172 VDD.t171 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1962 resistorDivider_v0p0p1_0.V12.t6 resistorDivider_v0p0p1_0.V11.t7 GND.t615 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1963 VIN.t31 w_55000_n29928# error sky130_fd_pr__cap_var_lvt w=2 l=0.18
X1964 GND.t265 16to4_PriorityEncoder_v0p0p1_0.x2.A a_82906_n51645# GND.t264 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X1965 OUT1.t67 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND.t273 GND.t272 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1966 VDD.t472 CLK.t94 w_55000_n3550# GND.t512 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1967 VDD.t843 frontAnalog_v0p0p1_4.x65.X frontAnalog_v0p0p1_4.RSfetsym_0.QN.t1 VDD.t842 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.25
X1968 a_53630_n68796# frontAnalog_v0p0p1_10.IB.t33 GND.t190 GND.t186 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1969 OUT3.t65 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND.t1261 GND.t1260 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1970 resistorDivider_v0p0p1_0.V8.t3 resistorDivider_v0p0p1_0.V7.t3 GND.t119 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1971 OUT2.t65 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND.t953 GND.t952 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1972 GND.t798 frontAnalog_v0p0p1_8.Q.t10 a_77725_n50381# GND.t797 sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X1973 GND.t271 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t66 GND.t270 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1974 a_82906_n47995# 16to4_PriorityEncoder_v0p0p1_0.x3.A1 GND.t1398 GND.t1397 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1975 VDD.t256 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t1 VDD.t255 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1976 16to4_PriorityEncoder_v0p0p1_0.x34.A a_82906_n43855# GND.t1414 GND.t1413 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1 ps=0.985 w=0.65 l=0.15
X1977 frontAnalog_v0p0p1_2.x63.X a_57123_n4079# GND.t1406 GND.t224 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1978 GND.t844 frontAnalog_v0p0p1_14.x65.X frontAnalog_v0p0p1_14.RSfetsym_0.x2.Y GND.t843 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1979 GND.t1503 16to4_PriorityEncoder_v0p0p1_0.x5.x17.A a_78065_n41309# GND.t1502 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X1980 GND.t418 frontAnalog_v0p0p1_1.Q.t8 a_77605_n39305# GND.t24 sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X1981 GND.t77 frontAnalog_v0p0p1_4.x63.X frontAnalog_v0p0p1_4.RSfetsym_0.x1.Y GND.t76 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1982 frontAnalog_v0p0p1_9.x63.A.t1 frontAnalog_v0p0p1_9.x65.A.t7 VDD.t459 VDD.t82 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1983 GND.t86 16to4_PriorityEncoder_v0p0p1_0.x28.A 16to4_PriorityEncoder_v0p0p1_0.x29.A GND.t85 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1984 VDD.t254 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t0 VDD.t253 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1985 frontAnalog_v0p0p1_10.x65.X a_57123_n56559# VDD.t869 VDD.t868 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1986 OUT3.t64 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND.t1259 GND.t1258 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1987 VDD.t700 16to4_PriorityEncoder_v0p0p1_0.x3.x19.C a_77605_n51335# VDD.t699 sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X1988 a_53630_n25596# frontAnalog_v0p0p1_10.IB.t34 GND.t191 GND.t186 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1989 OUT2.t64 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND.t951 GND.t950 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1990 a_77605_n43295# frontAnalog_v0p0p1_6.Q.t12 VDD.t881 VDD.t880 sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.109 ps=1.36 w=0.42 l=0.15
X1991 frontAnalog_v0p0p1_8.x63.A.t1 CLK.t95 w_55000_n46750# VDD.t186 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1992 GND.t1549 frontAnalog_v0p0p1_6.x65.A.t7 a_57123_n29559# GND.t1417 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X1993 VDD.t252 16to4_PriorityEncoder_v0p0p1_0.x2.A a_82988_n51645# VDD.t251 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X1994 a_16719_n13117.t0 a_16599_n13205.t23 a_16541_n13117.t19 GND.t1495 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1995 frontAnalog_v0p0p1_13.RSfetsym_0.QN.t3 frontAnalog_v0p0p1_13.RSfetsym_0.x1.Y GND.t526 GND.t525 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.25
X1996 GND.t752 16to4_PriorityEncoder_v0p0p1_0.x43.A 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND.t751 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1997 frontAnalog_v0p0p1_12.x63.X a_57123_n74279# GND.t18 GND.t17 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1998 OUT1.t65 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND.t269 GND.t268 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1999 GND.t267 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t64 GND.t266 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
R0 GND.n6411 GND.n515 5.63094e+06
R1 GND.n6461 GND 2.276e+06
R2 GND.n6461 GND 2.00869e+06
R3 GND.n6464 GND 334900
R4 GND.n6409 GND 334900
R5 GND.n5649 GND.n1004 273240
R6 GND.n7752 GND 271091
R7 GND GND.n5649 271091
R8 GND.n6464 GND.n716 215600
R9 GND.n6410 GND.n6409 215600
R10 GND.n3906 GND.n3905 98120
R11 GND.n3227 GND.n3225 20340.7
R12 GND.n2087 GND.n2085 20340.7
R13 GND.n2409 GND.n2407 20340.7
R14 GND.n2567 GND.n2565 20340.7
R15 GND.n2730 GND.n2728 20340.7
R16 GND.n7654 GND.n7653 20340.7
R17 GND.n3004 GND.n3002 20340.7
R18 GND.n3113 GND.n3111 20340.7
R19 GND.n5320 GND.n5318 20340.7
R20 GND.n4995 GND.n4993 20340.7
R21 GND.n3601 GND.n3599 20340.7
R22 GND.n4018 GND.n4016 20340.7
R23 GND.n1214 GND.n1212 20340.7
R24 GND.n7652 GND.n172 20169.3
R25 GND.n1419 GND.n1418 15044.8
R26 GND GND.n172 13209.6
R27 GND.n1212 GND 13209.6
R28 GND.n3225 GND 13209.6
R29 GND.n1418 GND 13209.6
R30 GND.n2085 GND 13209.6
R31 GND.n2407 GND 13209.6
R32 GND.n2565 GND 13209.6
R33 GND.n2728 GND 13209.6
R34 GND GND.n7654 13209.6
R35 GND.n3002 GND 13209.6
R36 GND.n3111 GND 13209.6
R37 GND.n5318 GND 13209.6
R38 GND.n4993 GND 13209.6
R39 GND.n3599 GND 13209.6
R40 GND.n4016 GND 13209.6
R41 GND GND.n3800 13209.6
R42 GND.n3800 GND.n171 12525.6
R43 GND.t1433 GND.n5 10105.3
R44 GND.n6415 GND.t627 10105.3
R45 GND.n2882 GND.n2881 8769.23
R46 GND.t545 GND.n1655 6847.68
R47 GND.t400 GND.n6463 5863.39
R48 GND.n6413 GND.t1510 5863.39
R49 GND GND.n7795 4548.57
R50 GND.n4682 GND.n4680 4526.39
R51 GND.n4725 GND.n4717 4526.39
R52 GND.n4725 GND.n4718 4526.07
R53 GND.n4707 GND.n4706 4525.74
R54 GND.n4682 GND.n4681 4525.74
R55 GND.n4659 GND.n4652 4525.74
R56 GND.n4729 GND.n4726 4525.74
R57 GND.n4679 GND.n4668 4525.09
R58 GND.n4699 GND.n4696 4519.41
R59 GND.n4181 GND.n4177 4519.41
R60 GND.n4176 GND.n4172 4519.41
R61 GND.n4176 GND.n4173 4519.41
R62 GND.n4171 GND.n4169 4519.41
R63 GND.n4168 GND.n4164 4519.41
R64 GND.n4701 GND.n4686 4519.41
R65 GND.n4701 GND.n4687 4519.41
R66 GND.n4163 GND.n4159 4519.41
R67 GND.n4163 GND.n4160 4519.41
R68 GND.n4154 GND.n4151 4519.41
R69 GND.n4154 GND.n4152 4519.41
R70 GND.n4147 GND.n4142 4519.41
R71 GND.n4147 GND.n4143 4519.41
R72 GND.n4695 GND.n4692 4519.41
R73 GND.n4695 GND.n4693 4519.41
R74 GND.n4141 GND.n4136 4519.41
R75 GND.n4141 GND.n4137 4519.41
R76 GND.n4135 GND.n4132 4519.41
R77 GND.n4691 GND.n4688 4519.41
R78 GND.n4691 GND.n4689 4519.41
R79 GND.n4131 GND.n4126 4519.41
R80 GND.n4131 GND.n4127 4519.41
R81 GND.n4643 GND.n4639 4377.09
R82 GND.n7652 GND.n173 4215.55
R83 GND.n4250 GND.n4228 3876.26
R84 GND.n4187 GND.n4113 3876.26
R85 GND.n6411 GND.t13 3455.76
R86 GND.t1278 GND.n5654 3428.59
R87 GND.n6409 GND.n6408 3003.29
R88 GND.n6412 GND.n6228 2817.54
R89 GND.n7795 GND.n4 2744.41
R90 GND.n6416 GND.n1004 2744.41
R91 GND.n6462 GND.t597 2656.51
R92 GND.n6459 GND.n6458 2243.42
R93 GND.n6460 GND.n6417 1899.15
R94 GND.n1940 GND.n1939 1773
R95 GND.n2258 GND.n2257 1773
R96 GND.n7186 GND.n7185 1773
R97 GND.n7020 GND.n7019 1773
R98 GND.n6866 GND.n6865 1773
R99 GND.n6712 GND.n6711 1773
R100 GND.n6564 GND.n6563 1773
R101 GND.n6589 GND.n6588 1773
R102 GND.n5486 GND.n5485 1773
R103 GND.n3346 GND.n3345 1773
R104 GND.n5171 GND.n5170 1773
R105 GND.n4847 GND.n4846 1773
R106 GND.n473 GND.n472 1773
R107 GND.n328 GND.n327 1773
R108 GND.n353 GND.n352 1773
R109 GND.n242 GND.n241 1773
R110 GND.n6461 GND.n6460 1742.45
R111 GND.n6463 GND.n6462 1566.95
R112 GND.n6463 GND.n5 1560.68
R113 GND.n6416 GND.n6415 1548.15
R114 GND.n6417 GND.n6416 1548.15
R115 GND.n7795 GND.n5 1535.61
R116 GND.t1423 GND.n1521 1402.22
R117 GND.n1885 GND.n1882 1390.42
R118 GND.n2210 GND.n2207 1390.42
R119 GND.n7141 GND.n7138 1390.42
R120 GND.n614 GND.n611 1390.42
R121 GND.n624 GND.n621 1390.42
R122 GND.n634 GND.n631 1390.42
R123 GND.n641 GND.n638 1390.42
R124 GND.n5553 GND.n5550 1390.42
R125 GND.n3431 GND.n3428 1390.42
R126 GND.n3337 GND.n3334 1390.42
R127 GND.n5118 GND.n5115 1390.42
R128 GND.n4797 GND.n4794 1390.42
R129 GND.n420 GND.n417 1390.42
R130 GND.n309 GND.n306 1390.42
R131 GND.n208 GND.n205 1390.42
R132 GND.n190 GND.n187 1390.42
R133 GND.n1942 GND.n1940 1384.79
R134 GND.n2260 GND.n2258 1384.79
R135 GND.n7188 GND.n7186 1384.79
R136 GND.n7022 GND.n7020 1384.79
R137 GND.n6868 GND.n6866 1384.79
R138 GND.n6714 GND.n6712 1384.79
R139 GND.n6566 GND.n6564 1384.79
R140 GND.n6591 GND.n6589 1384.79
R141 GND.n5488 GND.n5486 1384.79
R142 GND.n3348 GND.n3346 1384.79
R143 GND.n5173 GND.n5171 1384.79
R144 GND.n4849 GND.n4847 1384.79
R145 GND.n475 GND.n473 1384.79
R146 GND.n330 GND.n328 1384.79
R147 GND.n355 GND.n353 1384.79
R148 GND.n244 GND.n242 1384.79
R149 GND.n6414 GND.n6413 1309.97
R150 GND.n6460 GND.t677 1269.38
R151 GND.t548 GND 1255.01
R152 GND.t120 GND 1255.01
R153 GND.n4412 GND.n4406 1176.21
R154 GND.n4387 GND.n4382 1176.21
R155 GND.n4372 GND.n4367 1176.21
R156 GND.n4357 GND.n4352 1176.21
R157 GND.n4342 GND.n4337 1176.21
R158 GND.n4323 GND.n4318 1176.21
R159 GND.n4308 GND.n4303 1176.21
R160 GND.n4293 GND.n4288 1176.21
R161 GND.n4278 GND.n4273 1176.21
R162 GND.n4597 GND.n4222 1176.21
R163 GND.n4590 GND.n4580 1176.21
R164 GND.n4575 GND.n4574 1176.21
R165 GND.n4560 GND.n4559 1176.21
R166 GND.n4545 GND.n4544 1176.21
R167 GND.n4530 GND.n4529 1176.21
R168 GND.n4513 GND.n4512 1176.21
R169 GND.n4498 GND.n4497 1176.21
R170 GND.n4483 GND.n4482 1176.21
R171 GND.n4468 GND.n4467 1176.21
R172 GND.n4453 GND.n4452 1176.21
R173 GND.n4432 GND.n4431 1176.21
R174 GND.n4414 GND.n4413 1176.21
R175 GND.n4389 GND.n4388 1176.21
R176 GND.n4374 GND.n4373 1176.21
R177 GND.n4359 GND.n4358 1176.21
R178 GND.n4344 GND.n4343 1176.21
R179 GND.n4325 GND.n4324 1176.21
R180 GND.n4310 GND.n4309 1176.21
R181 GND.n4295 GND.n4294 1176.21
R182 GND.n4280 GND.n4279 1176.21
R183 GND.n4598 GND.n4218 1176.21
R184 GND.n4589 GND.n4584 1176.21
R185 GND.n4573 GND.n4568 1176.21
R186 GND.n4558 GND.n4553 1176.21
R187 GND.n4543 GND.n4538 1176.21
R188 GND.n4528 GND.n4523 1176.21
R189 GND.n4511 GND.n4506 1176.21
R190 GND.n4496 GND.n4491 1176.21
R191 GND.n4481 GND.n4476 1176.21
R192 GND.n4466 GND.n4461 1176.21
R193 GND.n4451 GND.n4444 1176.21
R194 GND.n4430 GND.n4424 1176.21
R195 GND.n1425 GND.n1395 1153.03
R196 GND.n2154 GND.n2151 1153.03
R197 GND.n2465 GND.n2462 1153.03
R198 GND.n2628 GND.n2625 1153.03
R199 GND.n2799 GND.n2796 1153.03
R200 GND.n2896 GND.n2893 1153.03
R201 GND.n7722 GND.n7719 1153.03
R202 GND.n3045 GND.n3042 1153.03
R203 GND.n3147 GND.n3144 1153.03
R204 GND.n1252 GND.n1249 1153.03
R205 GND.n3254 GND.n3251 1153.03
R206 GND.n5387 GND.n5384 1153.03
R207 GND.n5058 GND.n5055 1153.03
R208 GND.n3664 GND.n3661 1153.03
R209 GND.n4052 GND.n4049 1153.03
R210 GND.n3865 GND.n3862 1153.03
R211 GND.n7373 GND.t1483 1131.09
R212 GND GND.t886 1129.73
R213 GND.n4080 GND.n4073 1077.71
R214 GND.n1602 GND.n1597 1077.71
R215 GND.n1602 GND.n1598 1077.71
R216 GND.n1606 GND.n1603 1077.71
R217 GND.n1371 GND.n1368 1077.71
R218 GND.n1373 GND.n1366 1077.71
R219 GND.n1616 GND.n1612 1077.71
R220 GND.n2119 GND.n2116 1077.71
R221 GND.n2121 GND.n2114 1077.71
R222 GND.n1611 GND.n1607 1077.71
R223 GND.n1611 GND.n1608 1077.71
R224 GND.n1622 GND.n1617 1077.71
R225 GND.n1622 GND.n1618 1077.71
R226 GND.n1626 GND.n1623 1077.71
R227 GND.n2442 GND.n2439 1077.71
R228 GND.n2444 GND.n2437 1077.71
R229 GND.n1636 GND.n1633 1077.71
R230 GND.n2599 GND.n2596 1077.71
R231 GND.n2601 GND.n2594 1077.71
R232 GND.n1632 GND.n1627 1077.71
R233 GND.n1632 GND.n1628 1077.71
R234 GND.n1641 GND.n1637 1077.71
R235 GND.n1641 GND.n1638 1077.71
R236 GND.n1646 GND.n1642 1077.71
R237 GND.n2763 GND.n2760 1077.71
R238 GND.n2765 GND.n2758 1077.71
R239 GND.n1653 GND.n1647 1077.71
R240 GND.n1653 GND.n1648 1077.71
R241 GND.n1661 GND.n1654 1077.71
R242 GND.n2867 GND.n2866 1077.71
R243 GND.n2872 GND.n2871 1077.71
R244 GND.n1665 GND.n1662 1077.71
R245 GND.n1671 GND.n1666 1077.71
R246 GND.n1671 GND.n1667 1077.71
R247 GND.n7695 GND.n7692 1077.71
R248 GND.n7697 GND.n7690 1077.71
R249 GND.n1681 GND.n1676 1077.71
R250 GND.n1681 GND.n1677 1077.71
R251 GND.n3065 GND.n3062 1077.71
R252 GND.n3067 GND.n3060 1077.71
R253 GND.n1675 GND.n1672 1077.71
R254 GND.n1685 GND.n1682 1077.71
R255 GND.n1691 GND.n1686 1077.71
R256 GND.n1691 GND.n1687 1077.71
R257 GND.n3166 GND.n3163 1077.71
R258 GND.n3168 GND.n3161 1077.71
R259 GND.n1701 GND.n1696 1077.71
R260 GND.n1701 GND.n1697 1077.71
R261 GND.n1272 GND.n1269 1077.71
R262 GND.n1274 GND.n1267 1077.71
R263 GND.n1695 GND.n1692 1077.71
R264 GND.n1705 GND.n1702 1077.71
R265 GND.n1711 GND.n1706 1077.71
R266 GND.n1711 GND.n1707 1077.71
R267 GND.n3273 GND.n3270 1077.71
R268 GND.n3275 GND.n3268 1077.71
R269 GND.n1721 GND.n1717 1077.71
R270 GND.n1721 GND.n1718 1077.71
R271 GND.n5352 GND.n5349 1077.71
R272 GND.n5354 GND.n5347 1077.71
R273 GND.n1716 GND.n1712 1077.71
R274 GND.n1725 GND.n1722 1077.71
R275 GND.n1731 GND.n1726 1077.71
R276 GND.n1731 GND.n1727 1077.71
R277 GND.n5028 GND.n5025 1077.71
R278 GND.n5030 GND.n5023 1077.71
R279 GND.n1736 GND.n1732 1077.71
R280 GND.n1741 GND.n1737 1077.71
R281 GND.n1741 GND.n1738 1077.71
R282 GND.n3633 GND.n3630 1077.71
R283 GND.n3635 GND.n3628 1077.71
R284 GND.n4078 GND.n4075 1077.71
R285 GND.n3916 GND.n3911 1077.71
R286 GND.n3916 GND.n3912 1077.71
R287 GND.n3910 GND.n3907 1077.71
R288 GND.n3922 GND.n3917 1077.71
R289 GND.n3922 GND.n3918 1077.71
R290 GND.n3926 GND.n3923 1077.71
R291 GND.n3896 GND.n3888 1077.71
R292 GND.n3898 GND.n3886 1077.71
R293 GND GND.t908 1058.96
R294 GND GND.t633 1058.96
R295 GND GND.t640 1058.96
R296 GND GND.t539 1058.96
R297 GND GND.t113 1058.96
R298 GND GND.t180 1058.96
R299 GND GND.t200 1058.96
R300 GND GND.t562 1058.96
R301 GND GND.t173 1058.96
R302 GND GND.t810 1058.96
R303 GND GND.t40 1058.96
R304 GND GND.t646 1058.96
R305 GND GND.t76 1058.96
R306 GND GND.t237 1058.96
R307 GND GND.t1555 1058.96
R308 GND GND.t1407 1058.96
R309 GND.n4080 GND.n4072 1054.53
R310 GND.n1373 GND.n1365 1054.53
R311 GND.n2121 GND.n2113 1054.53
R312 GND.n2444 GND.n2436 1054.53
R313 GND.n2601 GND.n2593 1054.53
R314 GND.n2765 GND.n2757 1054.53
R315 GND.n2872 GND.n2870 1054.53
R316 GND.n7697 GND.n7689 1054.53
R317 GND.n3067 GND.n3059 1054.53
R318 GND.n3168 GND.n3160 1054.53
R319 GND.n1274 GND.n1266 1054.53
R320 GND.n3275 GND.n3267 1054.53
R321 GND.n5354 GND.n5346 1054.53
R322 GND.n5030 GND.n5022 1054.53
R323 GND.n3635 GND.n3627 1054.53
R324 GND.n3898 GND.n3885 1054.53
R325 GND.n5649 GND.n5648 940.789
R326 GND GND.t1085 917.571
R327 GND GND.t219 917.571
R328 GND.n1924 GND.n1920 915.471
R329 GND.n1950 GND.n1949 915.471
R330 GND.n1491 GND.n1490 915.471
R331 GND.n2247 GND.n2243 915.471
R332 GND.n2273 GND.n2272 915.471
R333 GND.n1908 GND.n1907 915.471
R334 GND.n7173 GND.n7169 915.471
R335 GND.n7203 GND.n7202 915.471
R336 GND.n2231 GND.n2230 915.471
R337 GND.n7007 GND.n7003 915.471
R338 GND.n7042 GND.n7041 915.471
R339 GND.n7157 GND.n7156 915.471
R340 GND.n6853 GND.n6849 915.471
R341 GND.n6888 GND.n6887 915.471
R342 GND.n6991 GND.n6990 915.471
R343 GND.n6699 GND.n6695 915.471
R344 GND.n6734 GND.n6733 915.471
R345 GND.n6837 GND.n6836 915.471
R346 GND.n6629 GND.n6625 915.471
R347 GND.n6576 GND.n6575 915.471
R348 GND.n6683 GND.n6682 915.471
R349 GND.n5526 GND.n5522 915.471
R350 GND.n5473 GND.n5472 915.471
R351 GND.n6613 GND.n6612 915.471
R352 GND.n1092 GND.n1088 915.471
R353 GND.n1046 GND.n1045 915.471
R354 GND.n5510 GND.n5509 915.471
R355 GND.n3400 GND.n3396 915.471
R356 GND.n3356 GND.n3355 915.471
R357 GND.n1076 GND.n1075 915.471
R358 GND.n5160 GND.n5156 915.471
R359 GND.n5183 GND.n5182 915.471
R360 GND.n3384 GND.n3383 915.471
R361 GND.n4836 GND.n4832 915.471
R362 GND.n4859 GND.n4858 915.471
R363 GND.n5144 GND.n5143 915.471
R364 GND.n462 GND.n458 915.471
R365 GND.n488 GND.n487 915.471
R366 GND.n4820 GND.n4819 915.471
R367 GND.n393 GND.n389 915.471
R368 GND.n340 GND.n339 915.471
R369 GND.n446 GND.n445 915.471
R370 GND.n282 GND.n278 915.471
R371 GND.n229 GND.n228 915.471
R372 GND.n377 GND.n376 915.471
R373 GND.n186 GND.n182 915.471
R374 GND.n7637 GND.n7636 915.471
R375 GND.n266 GND.n265 915.471
R376 GND.n1504 GND.n1501 841.244
R377 GND.n1926 GND.n1918 841.244
R378 GND.n2249 GND.n2241 841.244
R379 GND.n7175 GND.n7167 841.244
R380 GND.n7009 GND.n7001 841.244
R381 GND.n6855 GND.n6847 841.244
R382 GND.n6701 GND.n6693 841.244
R383 GND.n6631 GND.n6623 841.244
R384 GND.n5528 GND.n5520 841.244
R385 GND.n1094 GND.n1086 841.244
R386 GND.n3402 GND.n3394 841.244
R387 GND.n5162 GND.n5154 841.244
R388 GND.n4838 GND.n4830 841.244
R389 GND.n464 GND.n456 841.244
R390 GND.n395 GND.n387 841.244
R391 GND.n284 GND.n276 841.244
R392 GND.t728 GND.n7571 808.275
R393 GND.t262 GND.n7508 808.275
R394 GND.t701 GND.n7446 808.275
R395 GND.t898 GND.n4884 808.275
R396 GND.t144 GND.n5208 808.275
R397 GND.t513 GND.n3473 808.275
R398 GND.n5457 GND.t1391 808.275
R399 GND.t448 GND.t548 806.792
R400 GND.t659 GND.t120 806.792
R401 GND.n4636 GND.n4634 806.47
R402 GND GND.t65 784.713
R403 GND GND.t24 784.713
R404 GND.t597 GND.t862 780.297
R405 GND.t13 GND.t666 780.297
R406 GND.n1584 GND.n1580 778.15
R407 GND.n1584 GND.n1581 778.15
R408 GND.n2053 GND.n2048 778.15
R409 GND.n2053 GND.n2049 778.15
R410 GND.n2360 GND.n2355 778.15
R411 GND.n2360 GND.n2356 778.15
R412 GND.n2047 GND.n2042 778.15
R413 GND.n2047 GND.n2043 778.15
R414 GND.n2354 GND.n2349 778.15
R415 GND.n2354 GND.n2350 778.15
R416 GND.n2533 GND.n2528 778.15
R417 GND.n2533 GND.n2529 778.15
R418 GND.n2681 GND.n2676 778.15
R419 GND.n2681 GND.n2677 778.15
R420 GND.n2527 GND.n2522 778.15
R421 GND.n2527 GND.n2523 778.15
R422 GND.n2675 GND.n2670 778.15
R423 GND.n2675 GND.n2671 778.15
R424 GND.n2951 GND.n2946 778.15
R425 GND.n2951 GND.n2947 778.15
R426 GND.n2945 GND.n2940 778.15
R427 GND.n2945 GND.n2941 778.15
R428 GND.n126 GND.n113 778.15
R429 GND.n126 GND.n114 778.15
R430 GND.n112 GND.n107 778.15
R431 GND.n112 GND.n108 778.15
R432 GND.n1335 GND.n1330 778.15
R433 GND.n1335 GND.n1331 778.15
R434 GND.n5610 GND.n5605 778.15
R435 GND.n5610 GND.n5606 778.15
R436 GND.n1329 GND.n1324 778.15
R437 GND.n1329 GND.n1325 778.15
R438 GND.n5604 GND.n5599 778.15
R439 GND.n5604 GND.n5600 778.15
R440 GND.n1173 GND.n1168 778.15
R441 GND.n1173 GND.n1169 778.15
R442 GND.n3547 GND.n3542 778.15
R443 GND.n3547 GND.n3543 778.15
R444 GND.n1167 GND.n1162 778.15
R445 GND.n1167 GND.n1163 778.15
R446 GND.n3541 GND.n3536 778.15
R447 GND.n3541 GND.n3537 778.15
R448 GND.n5286 GND.n5281 778.15
R449 GND.n5286 GND.n5282 778.15
R450 GND.n4947 GND.n4942 778.15
R451 GND.n4947 GND.n4943 778.15
R452 GND.n5280 GND.n5275 778.15
R453 GND.n5280 GND.n5276 778.15
R454 GND.n4941 GND.n4936 778.15
R455 GND.n4941 GND.n4937 778.15
R456 GND.n3705 GND.n3700 778.15
R457 GND.n3705 GND.n3701 778.15
R458 GND.n3699 GND.n3694 778.15
R459 GND.n3699 GND.n3695 778.15
R460 GND.n3984 GND.n3979 778.15
R461 GND.n3984 GND.n3980 778.15
R462 GND.n3978 GND.n3973 778.15
R463 GND.n3978 GND.n3974 778.15
R464 GND.n3761 GND.n3756 778.15
R465 GND.n3761 GND.n3757 778.15
R466 GND.n3755 GND.n3750 778.15
R467 GND.n3755 GND.n3751 778.15
R468 GND.n3850 GND.n3846 778.15
R469 GND.n3850 GND.n3849 778.15
R470 GND.t797 GND.t228 777.333
R471 GND.t927 GND.t402 777.333
R472 GND GND.t865 754.5
R473 GND GND.t661 754.5
R474 GND.t1448 GND.t400 732.088
R475 GND.t838 GND.t1510 732.088
R476 GND.t1084 GND 729.721
R477 GND.t885 GND 729.721
R478 GND GND.t867 726
R479 GND.t662 GND 726
R480 GND.t920 GND.t167 717.149
R481 GND.t593 GND.t1502 717.149
R482 GND.t1085 GND.t207 708.047
R483 GND.t219 GND.t493 708.047
R484 GND.n6822 GND.t1445 706.715
R485 GND.n6976 GND.t945 706.715
R486 GND.t93 GND.n2298 706.715
R487 GND.t850 GND.n1975 706.715
R488 GND GND.t841 654.159
R489 GND.n6228 GND 654.054
R490 GND.t82 GND.t1448 627.505
R491 GND.t167 GND.t82 627.505
R492 GND.t865 GND.t448 627.505
R493 GND.t929 GND.t838 627.505
R494 GND.t1502 GND.t929 627.505
R495 GND.t661 GND.t659 627.505
R496 GND.t862 GND.t1084 606.898
R497 GND.t207 GND.t603 606.898
R498 GND.t603 GND.t1253 606.898
R499 GND.t666 GND.t885 606.898
R500 GND.t493 GND.t890 606.898
R501 GND.t890 GND.t801 606.898
R502 GND.t859 GND.t35 601.333
R503 GND.t1091 GND.t669 601.333
R504 GND.n7229 GND.t135 591.866
R505 GND.n5647 GND.t683 550.154
R506 GND GND.t818 546.497
R507 GND GND.t243 546.497
R508 GND.n1924 GND.n1921 521.471
R509 GND.n2247 GND.n2244 521.471
R510 GND.n7173 GND.n7170 521.471
R511 GND.n7007 GND.n7004 521.471
R512 GND.n6853 GND.n6850 521.471
R513 GND.n6699 GND.n6696 521.471
R514 GND.n6629 GND.n6626 521.471
R515 GND.n5526 GND.n5523 521.471
R516 GND.n1092 GND.n1089 521.471
R517 GND.n3400 GND.n3397 521.471
R518 GND.n5160 GND.n5157 521.471
R519 GND.n4836 GND.n4833 521.471
R520 GND.n462 GND.n459 521.471
R521 GND.n393 GND.n390 521.471
R522 GND.n282 GND.n279 521.471
R523 GND.n186 GND.n183 521.471
R524 GND.n1975 GND.n1974 515.509
R525 GND.n2298 GND.n2297 515.509
R526 GND.n7228 GND.n7227 515.509
R527 GND.n6978 GND.n6976 515.509
R528 GND.n6824 GND.n6822 515.509
R529 GND.n5646 GND.n5645 515.509
R530 GND.n5458 GND.n5457 515.509
R531 GND.n3473 GND.n3472 515.509
R532 GND.n5208 GND.n5207 515.509
R533 GND.n4884 GND.n4883 515.509
R534 GND.n7446 GND.n514 515.509
R535 GND.n7508 GND.n7507 515.509
R536 GND.n7571 GND.n7570 515.509
R537 GND.t741 GND 513.333
R538 GND.t852 GND.t670 498.408
R539 GND.n1887 GND 484.329
R540 GND.n2212 GND 484.329
R541 GND.n7143 GND 484.329
R542 GND.n616 GND 484.329
R543 GND.n626 GND 484.329
R544 GND.n636 GND 484.329
R545 GND.n643 GND 484.329
R546 GND.n5555 GND 484.329
R547 GND.n3433 GND 484.329
R548 GND.n3339 GND 484.329
R549 GND.n5120 GND 484.329
R550 GND.n4799 GND 484.329
R551 GND.n422 GND 484.329
R552 GND.n311 GND 484.329
R553 GND.n210 GND 484.329
R554 GND.n192 GND 484.329
R555 GND.n1429 GND.n1428 480.913
R556 GND.n2160 GND.n2150 480.913
R557 GND.n2469 GND.n2468 480.913
R558 GND.n2634 GND.n2624 480.913
R559 GND.n2803 GND.n2802 480.913
R560 GND.n2899 GND.n2880 480.913
R561 GND.n7726 GND.n7725 480.913
R562 GND.n3051 GND.n3041 480.913
R563 GND.n3151 GND.n3150 480.913
R564 GND.n1258 GND.n1248 480.913
R565 GND.n3258 GND.n3257 480.913
R566 GND.n5393 GND.n5383 480.913
R567 GND.n5062 GND.n5061 480.913
R568 GND.n3668 GND.n3667 480.913
R569 GND.n4058 GND.n4048 480.913
R570 GND.n3871 GND.n3861 480.913
R571 GND GND.t852 478.938
R572 GND GND.t920 478.099
R573 GND GND.t593 478.099
R574 GND.n1504 GND.n1502 473.865
R575 GND.n1926 GND.n1919 473.865
R576 GND.n2249 GND.n2242 473.865
R577 GND.n7175 GND.n7168 473.865
R578 GND.n7009 GND.n7002 473.865
R579 GND.n6855 GND.n6848 473.865
R580 GND.n6701 GND.n6694 473.865
R581 GND.n6631 GND.n6624 473.865
R582 GND.n5528 GND.n5521 473.865
R583 GND.n1094 GND.n1087 473.865
R584 GND.n3402 GND.n3395 473.865
R585 GND.n5162 GND.n5155 473.865
R586 GND.n4838 GND.n4831 473.865
R587 GND.n464 GND.n457 473.865
R588 GND.n395 GND.n388 473.865
R589 GND.n284 GND.n277 473.865
R590 GND.n6413 GND.n6412 445.014
R591 GND GND.t235 426.178
R592 GND.t841 GND.t1550 420.531
R593 GND.n716 GND 420.382
R594 GND.n6410 GND 420.382
R595 GND.t1253 GND.n716 419.048
R596 GND.t801 GND.n6410 419.048
R597 GND.t161 GND.n1355 405.955
R598 GND.t672 GND 393.274
R599 GND.t677 GND.t591 381.594
R600 GND.t159 GND.t171 373.805
R601 GND.n7444 GND.n515 367.533
R602 GND GND.t157 339.942
R603 GND GND.t156 339.942
R604 GND.n1372 GND.n1367 331.909
R605 GND.n2120 GND.n2115 331.909
R606 GND.n2443 GND.n2438 331.909
R607 GND.n2600 GND.n2595 331.909
R608 GND.n2764 GND.n2759 331.909
R609 GND.n7696 GND.n7691 331.909
R610 GND.n3066 GND.n3061 331.909
R611 GND.n3167 GND.n3162 331.909
R612 GND.n1273 GND.n1268 331.909
R613 GND.n3274 GND.n3269 331.909
R614 GND.n5353 GND.n5348 331.909
R615 GND.n5029 GND.n5024 331.909
R616 GND.n3634 GND.n3629 331.909
R617 GND.n4079 GND.n4074 331.909
R618 GND.n3897 GND.n3887 331.909
R619 GND.n3816 GND.n3815 328.866
R620 GND.n4018 GND.n4017 328.866
R621 GND.n3601 GND.n3600 328.866
R622 GND.n4995 GND.n4994 328.866
R623 GND.n5320 GND.n5319 328.866
R624 GND.n3227 GND.n3226 328.866
R625 GND.n1214 GND.n1213 328.866
R626 GND.n3113 GND.n3112 328.866
R627 GND.n3004 GND.n3003 328.866
R628 GND.n7653 GND.n7652 328.866
R629 GND.n2850 GND.n2849 328.866
R630 GND.n2730 GND.n2729 328.866
R631 GND.n2567 GND.n2566 328.866
R632 GND.n2409 GND.n2408 328.866
R633 GND.n2087 GND.n2086 328.866
R634 GND.t591 GND.t892 327.08
R635 GND.t892 GND.t159 327.08
R636 GND.t1550 GND.t672 327.08
R637 GND.t759 GND.t769 324.212
R638 GND.t781 GND.t771 324.212
R639 GND.t761 GND.t781 324.212
R640 GND.t767 GND.t761 324.212
R641 GND.t777 GND.t767 324.212
R642 GND.t773 GND.t777 324.212
R643 GND.t755 GND.t765 324.212
R644 GND.t763 GND.t751 324.212
R645 GND.t745 GND.t741 324.212
R646 GND.t747 GND.t745 324.212
R647 GND.t743 GND.t747 324.212
R648 GND.t1113 GND 308.692
R649 GND GND.t1101 308.692
R650 GND.t1179 GND 308.692
R651 GND.t1529 GND 308.692
R652 GND GND.t607 306.387
R653 GND.n7796 GND.t559 304.084
R654 GND GND.t763 301.053
R655 GND GND.n6459 299.824
R656 GND.n4130 GND.n4128 293.647
R657 GND.n4130 GND.n4129 293.647
R658 GND.n4134 GND.n4133 293.647
R659 GND.n4140 GND.n4138 293.647
R660 GND.n4140 GND.n4139 293.647
R661 GND.n4146 GND.n4144 293.647
R662 GND.n4146 GND.n4145 293.647
R663 GND.n4149 GND.n4148 293.647
R664 GND.n4157 GND.n4155 293.647
R665 GND.n4157 GND.n4156 293.647
R666 GND.n4162 GND.n4161 293.647
R667 GND.n4167 GND.n4165 293.647
R668 GND.n4167 GND.n4166 293.647
R669 GND.n4175 GND.n4174 293.647
R670 GND.n4180 GND.n4178 293.647
R671 GND.n4180 GND.n4179 293.647
R672 GND.n2887 GND.n2884 290.182
R673 GND.n6226 GND.t775 285.615
R674 GND.n2898 GND.n2882 285.455
R675 GND.t670 GND.t905 280.354
R676 GND.t905 GND.t658 280.354
R677 GND.n1420 GND.n1419 271.185
R678 GND.n6159 GND.t757 270.175
R679 GND.n7794 GND.n7793 267.089
R680 GND GND.t131 266.514
R681 GND GND.t154 266.514
R682 GND.t783 GND 263.26
R683 GND.n5647 GND.n5646 258.123
R684 GND.t658 GND 253.097
R685 GND.n6415 GND.n6414 250.713
R686 GND.t171 GND 249.204
R687 GND.t559 GND 244.189
R688 GND GND.t158 230.905
R689 GND GND.t153 230.905
R690 GND GND.t1413 227.501
R691 GND.t235 GND.t264 223.457
R692 GND.t879 GND 216.544
R693 GND.t290 GND.n737 214.877
R694 GND.n7793 GND.n7792 213.671
R695 GND.n6462 GND.n6461 213.106
R696 GND.n6227 GND 211.114
R697 GND.n1658 GND.n1657 209.695
R698 GND.n1651 GND.n1650 209.695
R699 GND.n1423 GND.n1422 203.294
R700 GND.n6412 GND.t773 196.843
R701 GND.n1381 GND.n1380 195.531
R702 GND.n2129 GND.n2128 195.531
R703 GND.n2452 GND.n2451 195.531
R704 GND.n2609 GND.n2608 195.531
R705 GND.n2773 GND.n2772 195.531
R706 GND.n7705 GND.n7704 195.531
R707 GND.n3075 GND.n3074 195.531
R708 GND.n3176 GND.n3175 195.531
R709 GND.n1282 GND.n1281 195.531
R710 GND.n3283 GND.n3282 195.531
R711 GND.n5362 GND.n5361 195.531
R712 GND.n5038 GND.n5037 195.531
R713 GND.n3643 GND.n3642 195.531
R714 GND.n4082 GND.n4070 195.531
R715 GND.n3900 GND.n3883 195.531
R716 GND.n1 GND.t606 193.933
R717 GND.n1436 GND.t911 193.933
R718 GND.n1524 GND.t1426 193.933
R719 GND.n1020 GND.t176 193.933
R720 GND.n1005 GND.t686 193.933
R721 GND.n6528 GND.t567 193.933
R722 GND.n6500 GND.t3 193.933
R723 GND.n7539 GND.t1558 193.933
R724 GND.n7511 GND.t256 193.933
R725 GND.n5076 GND.t647 193.933
R726 GND.n5211 GND.t147 193.933
R727 GND.n3287 GND.t41 193.933
R728 GND.n3476 GND.t517 193.933
R729 GND.n3442 GND.t814 193.933
R730 GND.n1113 GND.t1394 193.933
R731 GND.n6782 GND.t181 193.933
R732 GND.n6767 GND.t1439 193.933
R733 GND.n7105 GND.t540 193.933
R734 GND.n7077 GND.t138 193.933
R735 GND.n1842 GND.t637 193.933
R736 GND.n1978 GND.t844 193.933
R737 GND.n2177 GND.t641 193.933
R738 GND.n2301 GND.t96 193.933
R739 GND.n6936 GND.t114 193.933
R740 GND.n6921 GND.t939 193.933
R741 GND.n66 GND.t204 193.933
R742 GND.n51 GND.t711 193.933
R743 GND.n4755 GND.t80 193.933
R744 GND.n4887 GND.t901 193.933
R745 GND.n7477 GND.t238 193.933
R746 GND.n7449 GND.t695 193.933
R747 GND.n7602 GND.t1408 193.933
R748 GND.n7574 GND.t722 193.933
R749 GND.n6198 GND.t744 193.933
R750 GND.n979 GND.t88 193.933
R751 GND.n6092 GND.t51 193.933
R752 GND.t882 GND.n1003 193.532
R753 GND.t1137 GND.t1111 193.508
R754 GND.t1223 GND.t1137 193.508
R755 GND.t1115 GND.t1223 193.508
R756 GND.t1107 GND.t1115 193.508
R757 GND.t1129 GND.t1107 193.508
R758 GND.t1097 GND.t1155 193.508
R759 GND.t1133 GND.t1097 193.508
R760 GND.t1203 GND.t1133 193.508
R761 GND.t1099 GND.t1203 193.508
R762 GND.t1123 GND.t1099 193.508
R763 GND.t1187 GND.t1123 193.508
R764 GND.t1217 GND.t1187 193.508
R765 GND.t1149 GND.t1217 193.508
R766 GND.t1193 GND.t1149 193.508
R767 GND.t1181 GND.t1113 193.508
R768 GND.t1207 GND.t1181 193.508
R769 GND.t1105 GND.t1207 193.508
R770 GND.t1161 GND.t1195 193.508
R771 GND.t1195 GND.t1127 193.508
R772 GND.t1127 GND.t1165 193.508
R773 GND.t1165 GND.t1199 193.508
R774 GND.t1199 GND.t1135 193.508
R775 GND.t1135 GND.t1215 193.508
R776 GND.t1215 GND.t1147 193.508
R777 GND.t1147 GND.t1173 193.508
R778 GND.t1173 GND.t1221 193.508
R779 GND.t1221 GND.t1153 193.508
R780 GND.t1153 GND.t1177 193.508
R781 GND.t1101 GND.t1159 193.508
R782 GND.t1159 GND.t1189 193.508
R783 GND.t1189 GND.t1125 193.508
R784 GND.t1125 GND.t1211 193.508
R785 GND.t1185 GND.t1121 193.508
R786 GND.t1213 GND.t1185 193.508
R787 GND.t1143 GND.t1213 193.508
R788 GND.t1169 GND.t1143 193.508
R789 GND.t1145 GND.t1201 193.508
R790 GND.t1171 GND.t1145 193.508
R791 GND.t1117 GND.t1171 193.508
R792 GND.t1139 GND.t1117 193.508
R793 GND.t1157 GND.t1139 193.508
R794 GND.t1205 GND.t1179 193.508
R795 GND.t1103 GND.t1205 193.508
R796 GND.t1183 GND.t1103 193.508
R797 GND.t1141 GND.t1209 193.508
R798 GND.t1163 GND.t1141 193.508
R799 GND.t1197 GND.t1163 193.508
R800 GND.t1131 GND.t1197 193.508
R801 GND.t1167 GND.t1131 193.508
R802 GND.t1109 GND.t1167 193.508
R803 GND.t1191 GND.t1109 193.508
R804 GND.t1219 GND.t1191 193.508
R805 GND.t1151 GND.t1219 193.508
R806 GND.t1175 GND.t1151 193.508
R807 GND.t1119 GND.t1175 193.508
R808 GND.t1543 GND.t1529 193.508
R809 GND.t1523 GND.t1543 193.508
R810 GND.t1531 GND.t1541 193.508
R811 GND.t1541 GND.t1537 193.508
R812 GND.t1537 GND.t1545 193.508
R813 GND.t1545 GND.t1525 193.508
R814 GND.t1525 GND.t1539 193.508
R815 GND.t1539 GND.t1547 193.508
R816 GND.t1547 GND.t1527 193.508
R817 GND.t1527 GND.t1533 193.508
R818 GND.t1533 GND.t1517 193.508
R819 GND.t1517 GND.t1521 193.508
R820 GND.t1521 GND.t1535 193.508
R821 GND.t1535 GND.t1519 193.508
R822 GND.t607 GND.t609 193.508
R823 GND.t609 GND.t611 193.508
R824 GND.t611 GND.t605 193.508
R825 GND.t264 GND.t879 193.508
R826 GND.n560 GND.t608 192.982
R827 GND.n1449 GND.t909 192.982
R828 GND.n1539 GND.t1424 192.982
R829 GND.n1032 GND.t174 192.982
R830 GND.n1011 GND.t684 192.982
R831 GND.n6540 GND.t565 192.982
R832 GND.n6511 GND.t10 192.982
R833 GND.n7551 GND.t1557 192.982
R834 GND.n7522 GND.t263 192.982
R835 GND.n5089 GND.t650 192.982
R836 GND.n5222 GND.t145 192.982
R837 GND.n3300 GND.t44 192.982
R838 GND.n3487 GND.t514 192.982
R839 GND.n3454 GND.t812 192.982
R840 GND.n1119 GND.t1392 192.982
R841 GND.n6794 GND.t184 192.982
R842 GND.n6773 GND.t1446 192.982
R843 GND.n7117 GND.t543 192.982
R844 GND.n7088 GND.t136 192.982
R845 GND.n1854 GND.t635 192.982
R846 GND.n1989 GND.t851 192.982
R847 GND.n2186 GND.t644 192.982
R848 GND.n2312 GND.t94 192.982
R849 GND.n6948 GND.t117 192.982
R850 GND.n6927 GND.t946 192.982
R851 GND.n78 GND.t202 192.982
R852 GND.n56 GND.t718 192.982
R853 GND.n4767 GND.t78 192.982
R854 GND.n4898 GND.t899 192.982
R855 GND.n7489 GND.t241 192.982
R856 GND.n7460 GND.t702 192.982
R857 GND.n7614 GND.t1412 192.982
R858 GND.n7585 GND.t729 192.982
R859 GND.n6197 GND.t742 192.982
R860 GND.n969 GND.t90 192.982
R861 GND.n6082 GND.t53 192.982
R862 GND GND.t292 190.686
R863 GND.t280 GND 190.686
R864 GND GND.t358 190.686
R865 GND.t462 GND 190.686
R866 GND GND.t89 189.263
R867 GND.t1022 GND.n5858 185.69
R868 GND GND.t73 185.418
R869 GND GND.t433 185.418
R870 GND GND.t194 185.418
R871 GND GND.t56 185.418
R872 GND GND.t1094 185.418
R873 GND.t482 GND 185.418
R874 GND GND.t109 185.418
R875 GND GND.t111 185.418
R876 GND GND.t45 185.418
R877 GND GND.t197 185.418
R878 GND GND.t807 185.418
R879 GND GND.t794 185.418
R880 GND.t21 GND 185.418
R881 GND GND.t1417 185.418
R882 GND.t250 GND 185.418
R883 GND GND.t732 185.418
R884 GND.n716 GND 182.167
R885 GND.n6410 GND 182.167
R886 GND GND.t532 181.03
R887 GND GND.t155 181.03
R888 GND GND.t1193 179.686
R889 GND.t1177 GND 179.686
R890 GND GND.t1157 179.686
R891 GND.t1209 GND.n7374 179.686
R892 GND GND.t1119 179.686
R893 GND.t1519 GND 179.686
R894 GND.n4 GND 176.386
R895 GND.n1004 GND 176.386
R896 GND.t605 GND 172.775
R897 GND.n2093 GND.n2092 171.047
R898 GND.n2416 GND.n2414 171.047
R899 GND.n2573 GND.n2572 171.047
R900 GND.n2737 GND.n2735 171.047
R901 GND.n2856 GND.n2855 171.047
R902 GND.n7669 GND.n7667 171.047
R903 GND.n3010 GND.n3009 171.047
R904 GND.n3120 GND.n3118 171.047
R905 GND.n1220 GND.n1219 171.047
R906 GND.n3234 GND.n3232 171.047
R907 GND.n5326 GND.n5325 171.047
R908 GND.n5002 GND.n5000 171.047
R909 GND.n3607 GND.n3606 171.047
R910 GND.n4024 GND.n4023 171.047
R911 GND.n3823 GND.n3821 171.047
R912 GND.n1571 GND.n1568 170.613
R913 GND.t1024 GND 164.786
R914 GND GND.t1012 164.786
R915 GND.t962 GND 164.786
R916 GND GND.t1479 164.786
R917 GND GND.t52 163.555
R918 GND.n6116 GND.t412 162.326
R919 GND.n4412 GND.n4405 162.236
R920 GND.t1121 GND.n7372 161.257
R921 GND.n7787 GND.t717 159.185
R922 GND.n7816 GND.t880 154.006
R923 GND.n982 GND.t1398 154.006
R924 GND.n6095 GND.t674 154.006
R925 GND.n5380 GND.n5371 153.601
R926 GND.n1245 GND.n1236 153.601
R927 GND.n3038 GND.n3029 153.601
R928 GND.n2621 GND.n2618 153.601
R929 GND.n2147 GND.n2138 153.601
R930 GND.n1389 GND.n1387 153.601
R931 GND.n1389 GND.n1388 153.601
R932 GND.n2147 GND.n2146 153.601
R933 GND.n2456 GND.n2454 153.601
R934 GND.n2456 GND.n2455 153.601
R935 GND.n2621 GND.n2620 153.601
R936 GND.n2790 GND.n2781 153.601
R937 GND.n2790 GND.n2789 153.601
R938 GND.n2877 GND.n2876 153.601
R939 GND.n7713 GND.n7707 153.601
R940 GND.n7713 GND.n7712 153.601
R941 GND.n3038 GND.n3037 153.601
R942 GND.n3138 GND.n3136 153.601
R943 GND.n3138 GND.n3137 153.601
R944 GND.n1245 GND.n1244 153.601
R945 GND.n3245 GND.n3243 153.601
R946 GND.n3245 GND.n3244 153.601
R947 GND.n5380 GND.n5379 153.601
R948 GND.n5049 GND.n5040 153.601
R949 GND.n5049 GND.n5048 153.601
R950 GND.n3655 GND.n3645 153.601
R951 GND.n3655 GND.n3654 153.601
R952 GND.n4045 GND.n4044 153.601
R953 GND.n3858 GND.n3853 153.601
R954 GND.n3858 GND.n3857 153.601
R955 GND GND.t882 150.841
R956 GND.n28 GND.t692 150.465
R957 GND.n6352 GND.t172 150.465
R958 GND.n7767 GND.t1395 150.465
R959 GND.n663 GND.t921 150.465
R960 GND.n679 GND.t819 150.465
R961 GND.n712 GND.t1437 150.465
R962 GND.n6307 GND.t492 150.465
R963 GND.n6278 GND.t594 150.465
R964 GND.n6230 GND.t1450 150.465
R965 GND.n6263 GND.t1087 150.465
R966 GND.t1264 GND 149.645
R967 GND.t1294 GND 149.645
R968 GND GND.t1312 149.645
R969 GND GND.t753 149.645
R970 GND.n2092 GND.n2087 148.436
R971 GND.n2414 GND.n2409 148.436
R972 GND.n2572 GND.n2567 148.436
R973 GND.n2735 GND.n2730 148.436
R974 GND.n2855 GND.n2850 148.436
R975 GND.n3009 GND.n3004 148.436
R976 GND.n3118 GND.n3113 148.436
R977 GND.n1219 GND.n1214 148.436
R978 GND.n3232 GND.n3227 148.436
R979 GND.n5325 GND.n5320 148.436
R980 GND.n5000 GND.n4995 148.436
R981 GND.n3606 GND.n3601 148.436
R982 GND.n4023 GND.n4018 148.436
R983 GND.n3821 GND.n3816 148.436
R984 GND.t9 GND.n6497 140.822
R985 GND.n7795 GND 138.286
R986 GND.n6417 GND 138.286
R987 GND.t414 GND.t783 138.035
R988 GND.n3894 GND.n3893 137.827
R989 GND.n7753 GND.n7752 137.55
R990 GND GND.t1397 133.766
R991 GND.n4123 GND.n4114 130.844
R992 GND.t412 GND 130.352
R993 GND.n7375 GND.t1531 129.006
R994 GND.n6412 GND.n6411 128.821
R995 GND.n6414 GND.t759 127.368
R996 GND.n6412 GND.t755 127.368
R997 GND.n7285 GND.t1129 124.398
R998 GND.n7286 GND.t1161 124.398
R999 GND.n1356 GND.t161 123.612
R1000 GND.n2104 GND.t785 123.612
R1001 GND.n2427 GND.t17 123.612
R1002 GND.n2584 GND.t854 123.612
R1003 GND.n2748 GND.t675 123.612
R1004 GND.n7680 GND.t406 123.612
R1005 GND.n3021 GND.t870 123.612
R1006 GND.n3131 GND.t439 123.612
R1007 GND.n5337 GND.t410 123.612
R1008 GND.n5013 GND.t749 123.612
R1009 GND.n3618 GND.t1431 123.612
R1010 GND.n4035 GND.t872 123.612
R1011 GND.n3834 GND.t224 123.612
R1012 GND.n3202 GND.t585 123.612
R1013 GND.n2845 GND.t485 123.612
R1014 GND.n1188 GND.t689 123.612
R1015 GND.n3843 GND.n3842 123.472
R1016 GND.n1444 GND.n1443 121.112
R1017 GND.n1536 GND.n1535 121.112
R1018 GND.n1028 GND.n1027 121.112
R1019 GND.n5627 GND.n5626 121.112
R1020 GND.n6536 GND.n6535 121.112
R1021 GND.n6521 GND.n6520 121.112
R1022 GND.n7547 GND.n7546 121.112
R1023 GND.n7532 GND.n7531 121.112
R1024 GND.n5084 GND.n5083 121.112
R1025 GND.n5232 GND.n5231 121.112
R1026 GND.n3295 GND.n3294 121.112
R1027 GND.n3497 GND.n3496 121.112
R1028 GND.n3450 GND.n3449 121.112
R1029 GND.n5445 GND.n5444 121.112
R1030 GND.n6790 GND.n6789 121.112
R1031 GND.n6810 GND.n6809 121.112
R1032 GND.n7113 GND.n7112 121.112
R1033 GND.n7098 GND.n7097 121.112
R1034 GND.n1850 GND.n1849 121.112
R1035 GND.n1999 GND.n1998 121.112
R1036 GND.n2194 GND.n2193 121.112
R1037 GND.n2322 GND.n2321 121.112
R1038 GND.n6944 GND.n6943 121.112
R1039 GND.n6964 GND.n6963 121.112
R1040 GND.n74 GND.n73 121.112
R1041 GND.n53 GND.n52 121.112
R1042 GND.n4763 GND.n4762 121.112
R1043 GND.n4908 GND.n4907 121.112
R1044 GND.n7485 GND.n7484 121.112
R1045 GND.n7470 GND.n7469 121.112
R1046 GND.n7610 GND.n7609 121.112
R1047 GND.n7595 GND.n7594 121.112
R1048 GND.t73 GND.n1417 120.669
R1049 GND.t433 GND.n2084 120.669
R1050 GND.t194 GND.n2406 120.669
R1051 GND.t56 GND.n2564 120.669
R1052 GND.t1094 GND.n2727 120.669
R1053 GND.n7655 GND.t482 120.669
R1054 GND.t109 GND.n3001 120.669
R1055 GND.t111 GND.n3110 120.669
R1056 GND.t45 GND.n5317 120.669
R1057 GND.t197 GND.n4992 120.669
R1058 GND.t807 GND.n3598 120.669
R1059 GND.t794 GND.n4015 120.669
R1060 GND.n3801 GND.t21 120.669
R1061 GND.t1417 GND.n3224 120.669
R1062 GND.n2834 GND.t250 120.669
R1063 GND.t732 GND.n1211 120.669
R1064 GND.t316 GND.t290 119.534
R1065 GND.t274 GND.t316 119.534
R1066 GND.t294 GND.t274 119.534
R1067 GND.t286 GND.t294 119.534
R1068 GND.t308 GND.t286 119.534
R1069 GND.t334 GND.t276 119.534
R1070 GND.t276 GND.t312 119.534
R1071 GND.t312 GND.t382 119.534
R1072 GND.t382 GND.t278 119.534
R1073 GND.t278 GND.t302 119.534
R1074 GND.t302 GND.t368 119.534
R1075 GND.t368 GND.t268 119.534
R1076 GND.t268 GND.t328 119.534
R1077 GND.t328 GND.t374 119.534
R1078 GND.t292 GND.t360 119.534
R1079 GND.t360 GND.t386 119.534
R1080 GND.t386 GND.t284 119.534
R1081 GND.t376 GND.t340 119.534
R1082 GND.t306 GND.t376 119.534
R1083 GND.t344 GND.t306 119.534
R1084 GND.t380 GND.t344 119.534
R1085 GND.t314 GND.t380 119.534
R1086 GND.t266 GND.t314 119.534
R1087 GND.t326 GND.t266 119.534
R1088 GND.t352 GND.t326 119.534
R1089 GND.t272 GND.t352 119.534
R1090 GND.t332 GND.t272 119.534
R1091 GND.t356 GND.t332 119.534
R1092 GND.t338 GND.t280 119.534
R1093 GND.t370 GND.t338 119.534
R1094 GND.t304 GND.t370 119.534
R1095 GND.t390 GND.t304 119.534
R1096 GND.t300 GND.t366 119.534
R1097 GND.t366 GND.t392 119.534
R1098 GND.t392 GND.t322 119.534
R1099 GND.t322 GND.t348 119.534
R1100 GND.t348 GND.t364 119.534
R1101 GND.t364 GND.t324 119.534
R1102 GND.t324 GND.t350 119.534
R1103 GND.t350 GND.t296 119.534
R1104 GND.t296 GND.t318 119.534
R1105 GND.t318 GND.t336 119.534
R1106 GND.t358 GND.t384 119.534
R1107 GND.t384 GND.t282 119.534
R1108 GND.t282 GND.t362 119.534
R1109 GND.t320 GND.t388 119.534
R1110 GND.t342 GND.t320 119.534
R1111 GND.t378 GND.t342 119.534
R1112 GND.t310 GND.t378 119.534
R1113 GND.t346 GND.t310 119.534
R1114 GND.t288 GND.t346 119.534
R1115 GND.t372 GND.t288 119.534
R1116 GND.t270 GND.t372 119.534
R1117 GND.t330 GND.t270 119.534
R1118 GND.t354 GND.t330 119.534
R1119 GND.t298 GND.t354 119.534
R1120 GND.t476 GND.t462 119.534
R1121 GND.t456 GND.t476 119.534
R1122 GND.t464 GND.t474 119.534
R1123 GND.t474 GND.t470 119.534
R1124 GND.t470 GND.t478 119.534
R1125 GND.t478 GND.t458 119.534
R1126 GND.t458 GND.t472 119.534
R1127 GND.t472 GND.t480 119.534
R1128 GND.t480 GND.t460 119.534
R1129 GND.t460 GND.t466 119.534
R1130 GND.t466 GND.t450 119.534
R1131 GND.t450 GND.t454 119.534
R1132 GND.t454 GND.t468 119.534
R1133 GND.t468 GND.t452 119.534
R1134 GND.t89 GND.t91 119.534
R1135 GND.t91 GND.t85 119.534
R1136 GND.t85 GND.t87 119.534
R1137 GND.t1397 GND.t414 119.534
R1138 GND.t1413 GND.t877 119.285
R1139 GND.t65 GND.t507 119.109
R1140 GND.t818 GND.t703 119.109
R1141 GND.t24 GND.t555 119.109
R1142 GND.t243 GND.t595 119.109
R1143 GND.n7811 GND.n7810 118.1
R1144 GND.n987 GND.n986 118.1
R1145 GND.n6100 GND.n6099 118.1
R1146 GND.n690 GND.n689 117.984
R1147 GND.n6241 GND.n6240 117.984
R1148 GND.n7234 GND.t1112 117.626
R1149 GND.n727 GND.t291 117.626
R1150 GND.n5861 GND.t1023 117.626
R1151 GND.n5657 GND.t1279 117.007
R1152 GND.t388 GND.n926 116.689
R1153 GND.n4402 GND.n4401 116.329
R1154 GND.n48 GND.n47 116.052
R1155 GND.n6372 GND.n6371 116.052
R1156 GND.t673 GND 115.596
R1157 GND.n1935 GND.n1934 115.201
R1158 GND.n2264 GND.n2263 115.201
R1159 GND.n7194 GND.n7193 115.201
R1160 GND.n7033 GND.n7032 115.201
R1161 GND.n6879 GND.n6878 115.201
R1162 GND.n6725 GND.n6724 115.201
R1163 GND.n6668 GND.n6667 115.201
R1164 GND.n6598 GND.n6597 115.201
R1165 GND.n5495 GND.n5494 115.201
R1166 GND.n1061 GND.n1060 115.201
R1167 GND.n3369 GND.n3368 115.201
R1168 GND.n5129 GND.n5128 115.201
R1169 GND.n479 GND.n478 115.201
R1170 GND.n431 GND.n430 115.201
R1171 GND.n362 GND.n361 115.201
R1172 GND.n251 GND.n250 115.201
R1173 GND.n7229 GND.n7228 114.849
R1174 GND.n564 GND.n563 114.713
R1175 GND.n7379 GND.n7378 114.713
R1176 GND.n601 GND.n600 114.713
R1177 GND.n595 GND.n594 114.713
R1178 GND.n591 GND.n590 114.713
R1179 GND.n585 GND.n584 114.713
R1180 GND.n579 GND.n578 114.713
R1181 GND.n573 GND.n572 114.713
R1182 GND.n7426 GND.n7425 114.713
R1183 GND.n7418 GND.n7417 114.713
R1184 GND.n7411 GND.n7410 114.713
R1185 GND.n7407 GND.n7406 114.713
R1186 GND.n7401 GND.n7400 114.713
R1187 GND.n7395 GND.n7394 114.713
R1188 GND.n7389 GND.n7388 114.713
R1189 GND.n7331 GND.n7330 114.713
R1190 GND.n7338 GND.n7337 114.713
R1191 GND.n7364 GND.n7363 114.713
R1192 GND.n7360 GND.n7359 114.713
R1193 GND.n7354 GND.n7353 114.713
R1194 GND.n7348 GND.n7347 114.713
R1195 GND.n7342 GND.n7341 114.713
R1196 GND.n7247 GND.n7246 114.713
R1197 GND.n7290 GND.n7289 114.713
R1198 GND.n7297 GND.n7296 114.713
R1199 GND.n7301 GND.n7300 114.713
R1200 GND.n7307 GND.n7306 114.713
R1201 GND.n7313 GND.n7312 114.713
R1202 GND.n7319 GND.n7318 114.713
R1203 GND.n7233 GND.n7232 114.713
R1204 GND.n7238 GND.n7237 114.713
R1205 GND.n7280 GND.n7279 114.713
R1206 GND.n7275 GND.n7274 114.713
R1207 GND.n7269 GND.n7268 114.713
R1208 GND.n7263 GND.n7262 114.713
R1209 GND.n7257 GND.n7256 114.713
R1210 GND.n6214 GND.n6213 114.713
R1211 GND.n5817 GND.n5816 114.713
R1212 GND.n5811 GND.n5810 114.713
R1213 GND.n5805 GND.n5804 114.713
R1214 GND.n5801 GND.n5800 114.713
R1215 GND.n5795 GND.n5794 114.713
R1216 GND.n5787 GND.n5786 114.713
R1217 GND.n5781 GND.n5780 114.713
R1218 GND.n5771 GND.n5770 114.713
R1219 GND.n5765 GND.n5764 114.713
R1220 GND.n5758 GND.n5757 114.713
R1221 GND.n5689 GND.n5688 114.713
R1222 GND.n5698 GND.n5697 114.713
R1223 GND.n5704 GND.n5703 114.713
R1224 GND.n5710 GND.n5709 114.713
R1225 GND.n5722 GND.n5721 114.713
R1226 GND.n5728 GND.n5727 114.713
R1227 GND.n5748 GND.n5747 114.713
R1228 GND.n5743 GND.n5742 114.713
R1229 GND.n5736 GND.n5735 114.713
R1230 GND.n5651 GND.n5650 114.713
R1231 GND.n6140 GND.n6139 114.713
R1232 GND.n6153 GND.n6152 114.713
R1233 GND.n6163 GND.n6162 114.713
R1234 GND.n6170 GND.n6169 114.713
R1235 GND.n6174 GND.n6173 114.713
R1236 GND.n6180 GND.n6179 114.713
R1237 GND.n6186 GND.n6185 114.713
R1238 GND.n6193 GND.n6192 114.713
R1239 GND.n5660 GND.n5659 114.713
R1240 GND.n5668 GND.n5667 114.713
R1241 GND.n5674 GND.n5673 114.713
R1242 GND.n5678 GND.n5677 114.713
R1243 GND.n5844 GND.n5843 114.713
R1244 GND.n5838 GND.n5837 114.713
R1245 GND.n5832 GND.n5831 114.713
R1246 GND.n974 GND.n973 114.713
R1247 GND.n718 GND.n717 114.713
R1248 GND.n934 GND.n933 114.713
R1249 GND.n940 GND.n939 114.713
R1250 GND.n944 GND.n943 114.713
R1251 GND.n950 GND.n949 114.713
R1252 GND.n956 GND.n955 114.713
R1253 GND.n962 GND.n961 114.713
R1254 GND.n876 GND.n875 114.713
R1255 GND.n921 GND.n920 114.713
R1256 GND.n914 GND.n913 114.713
R1257 GND.n910 GND.n909 114.713
R1258 GND.n904 GND.n903 114.713
R1259 GND.n898 GND.n897 114.713
R1260 GND.n892 GND.n891 114.713
R1261 GND.n789 GND.n788 114.713
R1262 GND.n722 GND.n721 114.713
R1263 GND.n841 GND.n840 114.713
R1264 GND.n845 GND.n844 114.713
R1265 GND.n851 GND.n850 114.713
R1266 GND.n857 GND.n856 114.713
R1267 GND.n863 GND.n862 114.713
R1268 GND.n777 GND.n776 114.713
R1269 GND.n828 GND.n827 114.713
R1270 GND.n821 GND.n820 114.713
R1271 GND.n817 GND.n816 114.713
R1272 GND.n811 GND.n810 114.713
R1273 GND.n805 GND.n804 114.713
R1274 GND.n799 GND.n798 114.713
R1275 GND.n726 GND.n725 114.713
R1276 GND.n731 GND.n730 114.713
R1277 GND.n742 GND.n741 114.713
R1278 GND.n747 GND.n746 114.713
R1279 GND.n753 GND.n752 114.713
R1280 GND.n759 GND.n758 114.713
R1281 GND.n765 GND.n764 114.713
R1282 GND.n6087 GND.n6086 114.713
R1283 GND.n6039 GND.n6038 114.713
R1284 GND.n6047 GND.n6046 114.713
R1285 GND.n6053 GND.n6052 114.713
R1286 GND.n6057 GND.n6056 114.713
R1287 GND.n6063 GND.n6062 114.713
R1288 GND.n6069 GND.n6068 114.713
R1289 GND.n6075 GND.n6074 114.713
R1290 GND.n6125 GND.n6124 114.713
R1291 GND.n5853 GND.n5852 114.713
R1292 GND.n6005 GND.n6004 114.713
R1293 GND.n6009 GND.n6008 114.713
R1294 GND.n6015 GND.n6014 114.713
R1295 GND.n6021 GND.n6020 114.713
R1296 GND.n6027 GND.n6026 114.713
R1297 GND.n5958 GND.n5957 114.713
R1298 GND.n5965 GND.n5964 114.713
R1299 GND.n5991 GND.n5990 114.713
R1300 GND.n5987 GND.n5986 114.713
R1301 GND.n5981 GND.n5980 114.713
R1302 GND.n5975 GND.n5974 114.713
R1303 GND.n5969 GND.n5968 114.713
R1304 GND.n5874 GND.n5873 114.713
R1305 GND.n5917 GND.n5916 114.713
R1306 GND.n5924 GND.n5923 114.713
R1307 GND.n5928 GND.n5927 114.713
R1308 GND.n5934 GND.n5933 114.713
R1309 GND.n5940 GND.n5939 114.713
R1310 GND.n5946 GND.n5945 114.713
R1311 GND.n5860 GND.n5859 114.713
R1312 GND.n5865 GND.n5864 114.713
R1313 GND.n5907 GND.n5906 114.713
R1314 GND.n5902 GND.n5901 114.713
R1315 GND.n5896 GND.n5895 114.713
R1316 GND.n5890 GND.n5889 114.713
R1317 GND.n5884 GND.n5883 114.713
R1318 GND.n558 GND.t1530 113.734
R1319 GND.n555 GND.t1180 113.734
R1320 GND.n7326 GND.t1102 113.734
R1321 GND.n7244 GND.t1114 113.734
R1322 GND.n5823 GND.t1265 113.734
R1323 GND.n5687 GND.t1295 113.734
R1324 GND.n5717 GND.t1313 113.734
R1325 GND.n6148 GND.t754 113.734
R1326 GND.n883 GND.t463 113.734
R1327 GND.n871 GND.t359 113.734
R1328 GND.n784 GND.t281 113.734
R1329 GND.n772 GND.t293 113.734
R1330 GND.n6034 GND.t1480 113.734
R1331 GND.n5851 GND.t963 113.734
R1332 GND.n5953 GND.t1013 113.734
R1333 GND.n5871 GND.t1025 113.734
R1334 GND.n7373 GND.t1169 112.88
R1335 GND.n40 GND.n39 111.957
R1336 GND.n6364 GND.n6363 111.957
R1337 GND.n6479 GND.n6478 111.957
R1338 GND.n6481 GND.n6480 111.957
R1339 GND.n665 GND.n664 111.957
R1340 GND.n670 GND.n655 111.957
R1341 GND.n6389 GND.n6388 111.957
R1342 GND.n6391 GND.n6390 111.957
R1343 GND.n6280 GND.n6279 111.957
R1344 GND.n6285 GND.n6270 111.957
R1345 GND.n0 GND.t560 111.924
R1346 GND.n6203 GND.t1560 111.924
R1347 GND.n6200 GND.t887 111.924
R1348 GND.n981 GND.t883 111.924
R1349 GND.n6420 GND.t857 111.924
R1350 GND.n6421 GND.t34 111.924
R1351 GND.n6422 GND.t588 111.924
R1352 GND.n6423 GND.t447 111.924
R1353 GND.n6424 GND.t234 111.924
R1354 GND.n517 GND.t664 111.924
R1355 GND.n518 GND.t20 111.924
R1356 GND.n519 GND.t436 111.924
R1357 GND.n520 GND.t28 111.924
R1358 GND.n521 GND.t499 111.924
R1359 GND.n6094 GND.t413 111.924
R1360 GND.n559 GND.t1520 111.296
R1361 GND.n557 GND.t1120 111.296
R1362 GND.n554 GND.t1158 111.296
R1363 GND.n7325 GND.t1178 111.296
R1364 GND.n7243 GND.t1194 111.296
R1365 GND.n5824 GND.t1337 111.296
R1366 GND.n5686 GND.t1261 111.296
R1367 GND.n5716 GND.t1259 111.296
R1368 GND.n6147 GND.t1283 111.296
R1369 GND.n6196 GND.t764 111.296
R1370 GND.n968 GND.t453 111.296
R1371 GND.n882 GND.t299 111.296
R1372 GND.n870 GND.t337 111.296
R1373 GND.n783 GND.t357 111.296
R1374 GND.n771 GND.t375 111.296
R1375 GND.n6081 GND.t1470 111.296
R1376 GND.n6033 GND.t1031 111.296
R1377 GND.n5850 GND.t1069 111.296
R1378 GND.n5952 GND.t961 111.296
R1379 GND.n5870 GND.t977 111.296
R1380 GND.t374 GND 110.996
R1381 GND GND.t356 110.996
R1382 GND.t336 GND 110.996
R1383 GND GND.t298 110.996
R1384 GND.t452 GND 110.996
R1385 GND.n6465 GND.n6464 110.841
R1386 GND.n2842 GND.n2841 109.394
R1387 GND.n1352 GND.n1351 109.394
R1388 GND.n2101 GND.n2100 109.394
R1389 GND.n2424 GND.n2423 109.394
R1390 GND.n2581 GND.n2580 109.394
R1391 GND.n2745 GND.n2744 109.394
R1392 GND.n7677 GND.n7676 109.394
R1393 GND.n3018 GND.n3017 109.394
R1394 GND.n3128 GND.n3127 109.394
R1395 GND.n1185 GND.n1184 109.394
R1396 GND.n3199 GND.n3198 109.394
R1397 GND.n5334 GND.n5333 109.394
R1398 GND.n5010 GND.n5009 109.394
R1399 GND.n3615 GND.n3614 109.394
R1400 GND.n4032 GND.n4031 109.394
R1401 GND.n3831 GND.n3830 109.394
R1402 GND.n30 GND.n29 109.359
R1403 GND.n6354 GND.n6353 109.359
R1404 GND.n7764 GND.n7763 109.314
R1405 GND.n660 GND.n659 109.314
R1406 GND.n6304 GND.n6303 109.314
R1407 GND.n6275 GND.n6274 109.314
R1408 GND.n12 GND.t534 108.505
R1409 GND.n9 GND.t533 108.505
R1410 GND.n7760 GND.t866 108.505
R1411 GND.n7757 GND.t864 108.505
R1412 GND.n6334 GND.t906 108.505
R1413 GND.n6331 GND.t907 108.505
R1414 GND.n6300 GND.t665 108.505
R1415 GND.n6297 GND.t668 108.505
R1416 GND.n32 GND.n31 108.016
R1417 GND.n6356 GND.n6355 108.016
R1418 GND.n7765 GND.n7762 108.016
R1419 GND.n658 GND.n657 108.016
R1420 GND.n706 GND.n705 108.016
R1421 GND.n710 GND.n680 108.016
R1422 GND.n686 GND.n685 108.016
R1423 GND.n6305 GND.n6302 108.016
R1424 GND.n6273 GND.n6272 108.016
R1425 GND.n6257 GND.n6256 108.016
R1426 GND.n6261 GND.n6231 108.016
R1427 GND.n6237 GND.n6236 108.016
R1428 GND.n1197 GND.n1196 107.24
R1429 GND.n3210 GND.n3209 107.24
R1430 GND.n4001 GND.n4000 107.24
R1431 GND.n5303 GND.n5302 107.24
R1432 GND.n2987 GND.n2986 107.24
R1433 GND.n2550 GND.n2549 107.24
R1434 GND.n2070 GND.n2069 107.24
R1435 GND.n1401 GND.n1400 107.24
R1436 GND.n2392 GND.n2391 107.24
R1437 GND.n2713 GND.n2712 107.24
R1438 GND.n2826 GND.n2825 107.24
R1439 GND.n157 GND.n156 107.24
R1440 GND.n3096 GND.n3095 107.24
R1441 GND.n4978 GND.n4977 107.24
R1442 GND.n3584 GND.n3583 107.24
R1443 GND.n3792 GND.n3791 107.24
R1444 GND.t87 GND 106.728
R1445 GND.n703 GND.n702 105.975
R1446 GND.n683 GND.n682 105.975
R1447 GND.n693 GND.n688 105.975
R1448 GND.n6254 GND.n6253 105.975
R1449 GND.n6234 GND.n6233 105.975
R1450 GND.n6244 GND.n6239 105.975
R1451 GND.n834 GND.t300 105.305
R1452 GND.n5648 GND.t856 103.51
R1453 GND.t1048 GND.t1022 103.299
R1454 GND.t1006 GND.t1048 103.299
R1455 GND.t1026 GND.t1006 103.299
R1456 GND.t1018 GND.t1026 103.299
R1457 GND.t1040 GND.t1018 103.299
R1458 GND.t1008 GND.t1066 103.299
R1459 GND.t1044 GND.t1008 103.299
R1460 GND.t986 GND.t1044 103.299
R1461 GND.t1010 GND.t986 103.299
R1462 GND.t1034 GND.t1010 103.299
R1463 GND.t970 GND.t1034 103.299
R1464 GND.t1000 GND.t970 103.299
R1465 GND.t1060 GND.t1000 103.299
R1466 GND.t976 GND.t1060 103.299
R1467 GND.t964 GND.t1024 103.299
R1468 GND.t990 GND.t964 103.299
R1469 GND.t1016 GND.t990 103.299
R1470 GND.t1072 GND.t978 103.299
R1471 GND.t978 GND.t1038 103.299
R1472 GND.t1038 GND.t1076 103.299
R1473 GND.t1076 GND.t982 103.299
R1474 GND.t982 GND.t1046 103.299
R1475 GND.t1046 GND.t998 103.299
R1476 GND.t998 GND.t1058 103.299
R1477 GND.t1058 GND.t956 103.299
R1478 GND.t956 GND.t1004 103.299
R1479 GND.t1004 GND.t1064 103.299
R1480 GND.t1064 GND.t960 103.299
R1481 GND.t1012 GND.t1070 103.299
R1482 GND.t1070 GND.t972 103.299
R1483 GND.t972 GND.t1036 103.299
R1484 GND.t1036 GND.t994 103.299
R1485 GND.t968 GND.t1032 103.299
R1486 GND.t996 GND.t968 103.299
R1487 GND.t1054 GND.t996 103.299
R1488 GND.t952 GND.t1054 103.299
R1489 GND.t984 GND.t952 103.299
R1490 GND.t1056 GND.t984 103.299
R1491 GND.t954 GND.t1056 103.299
R1492 GND.t1028 GND.t954 103.299
R1493 GND.t1050 GND.t1028 103.299
R1494 GND.t1068 GND.t1050 103.299
R1495 GND.t988 GND.t962 103.299
R1496 GND.t1014 GND.t988 103.299
R1497 GND.t966 GND.t1014 103.299
R1498 GND.t992 GND.t1052 103.299
R1499 GND.t1052 GND.t1074 103.299
R1500 GND.t1074 GND.t980 103.299
R1501 GND.t980 GND.t1042 103.299
R1502 GND.t1042 GND.t950 103.299
R1503 GND.t950 GND.t1020 103.299
R1504 GND.t1020 GND.t974 103.299
R1505 GND.t974 GND.t1002 103.299
R1506 GND.t1002 GND.t1062 103.299
R1507 GND.t1062 GND.t958 103.299
R1508 GND.t958 GND.t1030 103.299
R1509 GND.t1479 GND.t1461 103.299
R1510 GND.t1461 GND.t1473 103.299
R1511 GND.t1481 GND.t1459 103.299
R1512 GND.t1459 GND.t1455 103.299
R1513 GND.t1455 GND.t1463 103.299
R1514 GND.t1463 GND.t1475 103.299
R1515 GND.t1475 GND.t1457 103.299
R1516 GND.t1457 GND.t1465 103.299
R1517 GND.t1465 GND.t1477 103.299
R1518 GND.t1477 GND.t1451 103.299
R1519 GND.t1451 GND.t1467 103.299
R1520 GND.t1467 GND.t1471 103.299
R1521 GND.t1471 GND.t1453 103.299
R1522 GND.t1453 GND.t1469 103.299
R1523 GND.t52 GND.t54 103.299
R1524 GND.t54 GND.t48 103.299
R1525 GND.t48 GND.t50 103.299
R1526 GND.t877 GND.t673 103.299
R1527 GND.n3810 GND.n3809 101.948
R1528 GND.n47 GND.t861 101.43
R1529 GND.n6371 GND.t671 101.43
R1530 GND.n3953 GND.n3944 100.894
R1531 GND.n5255 GND.n5246 100.894
R1532 GND.n3516 GND.n3507 100.894
R1533 GND.n1140 GND.n1131 100.894
R1534 GND.n5579 GND.n5570 100.894
R1535 GND.n1304 GND.n1295 100.894
R1536 GND.n2918 GND.n2909 100.894
R1537 GND.n2502 GND.n2493 100.894
R1538 GND.n2022 GND.n2013 100.894
R1539 GND.n1562 GND.n1555 100.894
R1540 GND.n2341 GND.n2332 100.894
R1541 GND.n2662 GND.n2653 100.894
R1542 GND.n99 GND.n90 100.894
R1543 GND.n4928 GND.n4919 100.894
R1544 GND.n3686 GND.n3677 100.894
R1545 GND.n3742 GND.n3733 100.894
R1546 GND.n7652 GND.n175 100.692
R1547 GND GND.t33 98.3051
R1548 GND GND.t587 98.3051
R1549 GND GND.t233 98.3051
R1550 GND GND.t446 97.1486
R1551 GND GND.t976 95.92
R1552 GND.t960 GND 95.92
R1553 GND GND.t1068 95.92
R1554 GND.n6118 GND.t992 95.92
R1555 GND.t1030 GND 95.92
R1556 GND.t1469 GND 95.92
R1557 GND.t1296 GND.t1278 93.8076
R1558 GND.t1368 GND.t1268 93.8076
R1559 GND.t1268 GND.t1318 93.8076
R1560 GND.t1318 GND.t1354 93.8076
R1561 GND.t1354 GND.t1272 93.8076
R1562 GND.t1272 GND.t1322 93.8076
R1563 GND.t1322 GND.t1358 93.8076
R1564 GND.t1380 GND.t1346 93.8076
R1565 GND.t1276 GND.t1380 93.8076
R1566 GND.t1350 GND.t1276 93.8076
R1567 GND.t1384 GND.t1350 93.8076
R1568 GND.t1310 GND.t1384 93.8076
R1569 GND.t1314 GND.t1264 93.8076
R1570 GND.t1348 GND.t1314 93.8076
R1571 GND.t1300 GND.t1348 93.8076
R1572 GND.t1262 GND.t1300 93.8076
R1573 GND.t1286 GND.t1262 93.8076
R1574 GND.t1342 GND.t1286 93.8076
R1575 GND.t1374 GND.t1342 93.8076
R1576 GND.t1274 GND.t1374 93.8076
R1577 GND.t1326 GND.t1274 93.8076
R1578 GND.t1378 GND.t1326 93.8076
R1579 GND.t1330 GND.t1304 93.8076
R1580 GND.t1362 GND.t1330 93.8076
R1581 GND.t1298 GND.t1362 93.8076
R1582 GND.t1260 GND.t1298 93.8076
R1583 GND.t1366 GND.t1294 93.8076
R1584 GND.t1280 GND.t1366 93.8076
R1585 GND.t1338 GND.t1280 93.8076
R1586 GND.t1370 GND.t1338 93.8076
R1587 GND.t1270 GND.t1370 93.8076
R1588 GND.t1320 GND.t1270 93.8076
R1589 GND.t1356 GND.t1292 93.8076
R1590 GND.t1292 GND.t1324 93.8076
R1591 GND.t1324 GND.t1290 93.8076
R1592 GND.t1290 GND.t1352 93.8076
R1593 GND.t1352 GND.t1382 93.8076
R1594 GND.t1382 GND.t1308 93.8076
R1595 GND.t1308 GND.t1334 93.8076
R1596 GND.t1334 GND.t1258 93.8076
R1597 GND.t1312 GND.t1364 93.8076
R1598 GND.t1364 GND.t1266 93.8076
R1599 GND.t1266 GND.t1316 93.8076
R1600 GND.t1316 GND.t1284 93.8076
R1601 GND.t1284 GND.t1340 93.8076
R1602 GND.t1372 GND.t1288 93.8076
R1603 GND.t1288 GND.t1344 93.8076
R1604 GND.t1344 GND.t1376 93.8076
R1605 GND.t1376 GND.t1302 93.8076
R1606 GND.t1302 GND.t1328 93.8076
R1607 GND.t1328 GND.t1360 93.8076
R1608 GND.t1360 GND.t1306 93.8076
R1609 GND.t1306 GND.t1332 93.8076
R1610 GND.t1332 GND.t1282 93.8076
R1611 GND.t50 GND 92.2308
R1612 GND.n3970 GND.n3967 91.8593
R1613 GND.n5272 GND.n5269 91.8593
R1614 GND.n3533 GND.n3530 91.8593
R1615 GND.n1159 GND.n1156 91.8593
R1616 GND.n5596 GND.n5593 91.8593
R1617 GND.n1321 GND.n1318 91.8593
R1618 GND.n2937 GND.n2934 91.8593
R1619 GND.n2519 GND.n2516 91.8593
R1620 GND.n2039 GND.n2036 91.8593
R1621 GND.n1577 GND.n1574 91.8593
R1622 GND.n2376 GND.n2373 91.8593
R1623 GND.n2697 GND.n2694 91.8593
R1624 GND.n142 GND.n139 91.8593
R1625 GND.n4963 GND.n4960 91.8593
R1626 GND.n3721 GND.n3718 91.8593
R1627 GND.n3777 GND.n3774 91.8593
R1628 GND.n1500 GND.n1499 90.3534
R1629 GND.n1917 GND.n1916 90.3534
R1630 GND.n2240 GND.n2239 90.3534
R1631 GND.n7166 GND.n7165 90.3534
R1632 GND.n7000 GND.n6999 90.3534
R1633 GND.n6846 GND.n6845 90.3534
R1634 GND.n6692 GND.n6691 90.3534
R1635 GND.n6622 GND.n6621 90.3534
R1636 GND.n5519 GND.n5518 90.3534
R1637 GND.n1085 GND.n1084 90.3534
R1638 GND.n3393 GND.n3392 90.3534
R1639 GND.n5153 GND.n5152 90.3534
R1640 GND.n4829 GND.n4828 90.3534
R1641 GND.n455 GND.n454 90.3534
R1642 GND.n386 GND.n385 90.3534
R1643 GND.n275 GND.n274 90.3534
R1644 GND.n1884 GND.n1883 90.3427
R1645 GND.n3430 GND.n3429 90.3427
R1646 GND.n5552 GND.n5551 90.3427
R1647 GND.n207 GND.n206 90.3427
R1648 GND.n4796 GND.n4795 90.3427
R1649 GND.n5117 GND.n5116 90.3427
R1650 GND.n3336 GND.n3335 90.3427
R1651 GND.n633 GND.n632 90.3427
R1652 GND.n613 GND.n612 90.3427
R1653 GND.n2209 GND.n2208 90.3427
R1654 GND.n7140 GND.n7139 90.3427
R1655 GND.n623 GND.n622 90.3427
R1656 GND.n640 GND.n639 90.3427
R1657 GND.n419 GND.n418 90.3427
R1658 GND.n308 GND.n307 90.3427
R1659 GND.n189 GND.n188 90.3427
R1660 GND.n7796 GND 87.5398
R1661 GND.n5692 GND.t1310 87.1071
R1662 GND GND.t1336 87.1071
R1663 GND GND.t1260 87.1071
R1664 GND.t1258 GND 87.1071
R1665 GND.t1282 GND 87.1071
R1666 GND.n1467 GND.n1466 86.1558
R1667 GND.n5461 GND.n5460 86.1558
R1668 GND.n5642 GND.n5641 86.1558
R1669 GND.n7567 GND.n7566 86.1558
R1670 GND.n5106 GND.n5105 86.1558
R1671 GND.n3315 GND.n3314 86.1558
R1672 GND.n3470 GND.n3469 86.1558
R1673 GND.n629 GND.n628 86.1558
R1674 GND.n609 GND.n608 86.1558
R1675 GND.n1872 GND.n1871 86.1558
R1676 GND.n7130 GND.n7129 86.1558
R1677 GND.n619 GND.n618 86.1558
R1678 GND.n6653 GND.n6652 86.1558
R1679 GND.n4785 GND.n4784 86.1558
R1680 GND.n7505 GND.n7504 86.1558
R1681 GND.n199 GND.n198 86.1558
R1682 GND.n1519 GND.n1518 86.1558
R1683 GND.n1972 GND.n1971 86.1558
R1684 GND.n2295 GND.n2294 86.1558
R1685 GND.n7225 GND.n7224 86.1558
R1686 GND.n6981 GND.n6980 86.1558
R1687 GND.n6827 GND.n6826 86.1558
R1688 GND.n6663 GND.n6662 86.1558
R1689 GND.n647 GND.n646 86.1558
R1690 GND.n5466 GND.n5465 86.1558
R1691 GND.n3423 GND.n3422 86.1558
R1692 GND.n3321 GND.n3320 86.1558
R1693 GND.n5205 GND.n5204 86.1558
R1694 GND.n4881 GND.n4880 86.1558
R1695 GND.n512 GND.n511 86.1558
R1696 GND.n315 GND.n314 86.1558
R1697 GND.n213 GND.n212 86.1558
R1698 GND.t1032 GND.n5999 86.0821
R1699 GND.n927 GND.t464 85.3821
R1700 GND.t803 GND.t248 84.4087
R1701 GND.n2031 GND.n2030 83.5572
R1702 GND.n2368 GND.n2365 83.5572
R1703 GND.n2511 GND.n2510 83.5572
R1704 GND.n2689 GND.n2686 83.5572
R1705 GND.n2929 GND.n2926 83.5572
R1706 GND.n134 GND.n131 83.5572
R1707 GND.n1313 GND.n1310 83.5572
R1708 GND.n5588 GND.n5585 83.5572
R1709 GND.n1151 GND.n1148 83.5572
R1710 GND.n3525 GND.n3522 83.5572
R1711 GND.n5264 GND.n5263 83.5572
R1712 GND.n4955 GND.n4952 83.5572
R1713 GND.n3713 GND.n3710 83.5572
R1714 GND.n3962 GND.n3959 83.5572
R1715 GND.n3769 GND.n3766 83.5572
R1716 GND.t340 GND.n833 82.5361
R1717 GND.n2093 GND.n2064 81.2313
R1718 GND.n2573 GND.n2544 81.2313
R1719 GND.n2856 GND.n2848 81.2313
R1720 GND.n3010 GND.n2981 81.2313
R1721 GND.n1220 GND.n1191 81.2313
R1722 GND.n5326 GND.n5297 81.2313
R1723 GND.n3607 GND.n3578 81.2313
R1724 GND.n4024 GND.n3995 81.2313
R1725 GND.t1201 GND.n7373 80.6288
R1726 GND.t1304 GND.n5693 80.4066
R1727 GND.n7652 GND.n179 79.3342
R1728 GND.n1557 GND.n1556 78.6829
R1729 GND.n3893 GND.n3892 78.6829
R1730 GND.n4051 GND.n4050 74.9181
R1731 GND.n1424 GND.n1423 74.9181
R1732 GND.n2153 GND.n2152 74.9181
R1733 GND.n2464 GND.n2463 74.9181
R1734 GND.n2627 GND.n2626 74.9181
R1735 GND.n2798 GND.n2797 74.9181
R1736 GND.n2895 GND.n2894 74.9181
R1737 GND.n7721 GND.n7720 74.9181
R1738 GND.n3044 GND.n3043 74.9181
R1739 GND.n3146 GND.n3145 74.9181
R1740 GND.n1251 GND.n1250 74.9181
R1741 GND.n3253 GND.n3252 74.9181
R1742 GND.n5386 GND.n5385 74.9181
R1743 GND.n5057 GND.n5056 74.9181
R1744 GND.n3663 GND.n3662 74.9181
R1745 GND.n3864 GND.n3863 74.9181
R1746 GND.t158 GND.t487 73.7614
R1747 GND.t153 GND.t163 73.7614
R1748 GND.n39 GND.t571 72.8576
R1749 GND.n6363 GND.t1551 72.8576
R1750 GND.n6478 GND.t798 72.8576
R1751 GND.n6480 GND.t36 72.8576
R1752 GND.n664 GND.t589 72.8576
R1753 GND.n655 GND.t449 72.8576
R1754 GND.n689 GND.t863 72.8576
R1755 GND.n6388 GND.t403 72.8576
R1756 GND.n6390 GND.t1092 72.8576
R1757 GND.n6279 GND.t660 72.8576
R1758 GND.n6270 GND.t1251 72.8576
R1759 GND.n6240 GND.t667 72.8576
R1760 GND.t399 GND.t211 72.6261
R1761 GND.t59 GND.t196 72.6261
R1762 GND.t506 GND.t75 72.6261
R1763 GND.t693 GND.t84 72.6261
R1764 GND.t615 GND.t119 72.6261
R1765 GND.n716 GND 72.2501
R1766 GND.n6410 GND 72.2501
R1767 GND.t914 GND.n1888 71.7802
R1768 GND.t868 GND.n2213 71.7802
R1769 GND.t1403 GND.n7144 71.7802
R1770 GND.t525 GND.n617 71.7802
R1771 GND.t621 GND.n627 71.7802
R1772 GND.t936 GND.n637 71.7802
R1773 GND.t226 GND.n644 71.7802
R1774 GND.t0 GND.n5556 71.7802
R1775 GND.t623 GND.n3434 71.7802
R1776 GND.t536 GND.n3340 71.7802
R1777 GND.t1488 GND.n5121 71.7802
R1778 GND.t423 GND.n4800 71.7802
R1779 GND.t550 GND.n423 71.7802
R1780 GND.t568 GND.n312 71.7802
R1781 GND.t719 GND.n211 71.7802
R1782 GND.n738 GND.t308 71.1519
R1783 GND.n3909 GND.n3908 70.024
R1784 GND.n4077 GND.n4076 70.024
R1785 GND.n1275 GND.n1265 70.024
R1786 GND.n3068 GND.n3058 70.024
R1787 GND.n1374 GND.n1364 70.024
R1788 GND.n1370 GND.n1369 70.024
R1789 GND.n1605 GND.n1604 70.024
R1790 GND.n1601 GND.n1599 70.024
R1791 GND.n1601 GND.n1600 70.024
R1792 GND.n2122 GND.n2112 70.024
R1793 GND.n2118 GND.n2117 70.024
R1794 GND.n1615 GND.n1613 70.024
R1795 GND.n1615 GND.n1614 70.024
R1796 GND.n1610 GND.n1609 70.024
R1797 GND.n2445 GND.n2435 70.024
R1798 GND.n2441 GND.n2440 70.024
R1799 GND.n1625 GND.n1624 70.024
R1800 GND.n1621 GND.n1619 70.024
R1801 GND.n1621 GND.n1620 70.024
R1802 GND.n2602 GND.n2592 70.024
R1803 GND.n2598 GND.n2597 70.024
R1804 GND.n1635 GND.n1634 70.024
R1805 GND.n1631 GND.n1629 70.024
R1806 GND.n1631 GND.n1630 70.024
R1807 GND.n2766 GND.n2756 70.024
R1808 GND.n2762 GND.n2761 70.024
R1809 GND.n1645 GND.n1643 70.024
R1810 GND.n1645 GND.n1644 70.024
R1811 GND.n1640 GND.n1639 70.024
R1812 GND.n1660 GND.n1658 70.024
R1813 GND.n1660 GND.n1659 70.024
R1814 GND.n2868 GND.n2865 70.024
R1815 GND.n2873 GND.n2869 70.024
R1816 GND.n1652 GND.n1651 70.024
R1817 GND.n7698 GND.n7688 70.024
R1818 GND.n7694 GND.n7693 70.024
R1819 GND.n1670 GND.n1668 70.024
R1820 GND.n1670 GND.n1669 70.024
R1821 GND.n1664 GND.n1663 70.024
R1822 GND.n3064 GND.n3063 70.024
R1823 GND.n1680 GND.n1678 70.024
R1824 GND.n1680 GND.n1679 70.024
R1825 GND.n1674 GND.n1673 70.024
R1826 GND.n3169 GND.n3159 70.024
R1827 GND.n3165 GND.n3164 70.024
R1828 GND.n1690 GND.n1688 70.024
R1829 GND.n1690 GND.n1689 70.024
R1830 GND.n1684 GND.n1683 70.024
R1831 GND.n1271 GND.n1270 70.024
R1832 GND.n1700 GND.n1698 70.024
R1833 GND.n1700 GND.n1699 70.024
R1834 GND.n1694 GND.n1693 70.024
R1835 GND.n3276 GND.n3266 70.024
R1836 GND.n3272 GND.n3271 70.024
R1837 GND.n1710 GND.n1708 70.024
R1838 GND.n1710 GND.n1709 70.024
R1839 GND.n1704 GND.n1703 70.024
R1840 GND.n5355 GND.n5345 70.024
R1841 GND.n5351 GND.n5350 70.024
R1842 GND.n1720 GND.n1719 70.024
R1843 GND.n1715 GND.n1713 70.024
R1844 GND.n1715 GND.n1714 70.024
R1845 GND.n5031 GND.n5021 70.024
R1846 GND.n5027 GND.n5026 70.024
R1847 GND.n1730 GND.n1728 70.024
R1848 GND.n1730 GND.n1729 70.024
R1849 GND.n1724 GND.n1723 70.024
R1850 GND.n1735 GND.n1733 70.024
R1851 GND.n1735 GND.n1734 70.024
R1852 GND.n1740 GND.n1739 70.024
R1853 GND.n3632 GND.n3631 70.024
R1854 GND.n3636 GND.n3626 70.024
R1855 GND.n3915 GND.n3913 70.024
R1856 GND.n3915 GND.n3914 70.024
R1857 GND.n4081 GND.n4071 70.024
R1858 GND.n3895 GND.n3894 70.024
R1859 GND.n3921 GND.n3919 70.024
R1860 GND.n3921 GND.n3920 70.024
R1861 GND.n3925 GND.n3924 70.024
R1862 GND.n3899 GND.n3884 70.024
R1863 GND.t1155 GND.n7285 69.1104
R1864 GND.n7286 GND.t1105 69.1104
R1865 GND.n6117 GND.t1481 68.8658
R1866 GND.n6497 GND.n6496 68.1084
R1867 GND.n13 GND.n12 67.973
R1868 GND.n10 GND.n9 67.973
R1869 GND.n7771 GND.n7760 67.973
R1870 GND.n7758 GND.n7757 67.973
R1871 GND.n6335 GND.n6334 67.973
R1872 GND.n6332 GND.n6331 67.973
R1873 GND.n6311 GND.n6300 67.973
R1874 GND.n6298 GND.n6297 67.973
R1875 GND.n123 GND.n122 67.5205
R1876 GND.n3853 GND.n3852 67.5205
R1877 GND.n5655 GND.t1296 67.0056
R1878 GND.n5912 GND.t1040 66.4063
R1879 GND.n5913 GND.t1072 66.4063
R1880 GND.t1340 GND.n5753 64.7721
R1881 GND.n7375 GND.t1523 64.5031
R1882 GND.n7652 GND.n171 64.3169
R1883 GND.t856 GND 61.2963
R1884 GND.t33 GND 61.2963
R1885 GND.t587 GND 61.2963
R1886 GND.t446 GND 61.2963
R1887 GND.t233 GND 61.2963
R1888 GND.n1923 GND.n1922 59.4829
R1889 GND.n1091 GND.n1090 59.4829
R1890 GND.n5525 GND.n5524 59.4829
R1891 GND.n281 GND.n280 59.4829
R1892 GND.n4835 GND.n4834 59.4829
R1893 GND.n5159 GND.n5158 59.4829
R1894 GND.n3399 GND.n3398 59.4829
R1895 GND.n6698 GND.n6697 59.4829
R1896 GND.n7006 GND.n7005 59.4829
R1897 GND.n2246 GND.n2245 59.4829
R1898 GND.n7172 GND.n7171 59.4829
R1899 GND.n6852 GND.n6851 59.4829
R1900 GND.n6628 GND.n6627 59.4829
R1901 GND.n461 GND.n460 59.4829
R1902 GND.n392 GND.n391 59.4829
R1903 GND.n185 GND.n184 59.4829
R1904 GND.n2874 GND.n2868 57.977
R1905 GND.t131 GND.t425 57.8291
R1906 GND.t532 GND.t789 57.8291
R1907 GND.t154 GND.t169 57.8291
R1908 GND.t155 GND.t836 57.8291
R1909 GND.n1282 GND.n1275 57.224
R1910 GND.n3075 GND.n3068 57.224
R1911 GND.n1381 GND.n1374 57.224
R1912 GND.n2129 GND.n2122 57.224
R1913 GND.n2452 GND.n2445 57.224
R1914 GND.n2609 GND.n2602 57.224
R1915 GND.n2773 GND.n2766 57.224
R1916 GND.n2874 GND.n2873 57.224
R1917 GND.n7705 GND.n7698 57.224
R1918 GND.n3176 GND.n3169 57.224
R1919 GND.n3283 GND.n3276 57.224
R1920 GND.n5362 GND.n5355 57.224
R1921 GND.n5038 GND.n5031 57.224
R1922 GND.n3643 GND.n3636 57.224
R1923 GND.n4082 GND.n4081 57.224
R1924 GND.n3900 GND.n3899 57.224
R1925 GND.n6414 GND.t753 56.9548
R1926 GND.n7810 GND.t265 55.7148
R1927 GND.n986 GND.t415 55.7148
R1928 GND.n6099 GND.t878 55.7148
R1929 GND.n3890 GND.n3889 54.813
R1930 GND.n1505 GND.n1500 54.66
R1931 GND.n1927 GND.n1917 54.66
R1932 GND.n2250 GND.n2240 54.66
R1933 GND.n7176 GND.n7166 54.66
R1934 GND.n7010 GND.n7000 54.66
R1935 GND.n6856 GND.n6846 54.66
R1936 GND.n6702 GND.n6692 54.66
R1937 GND.n6632 GND.n6622 54.66
R1938 GND.n5529 GND.n5519 54.66
R1939 GND.n1095 GND.n1085 54.66
R1940 GND.n3403 GND.n3393 54.66
R1941 GND.n5163 GND.n5153 54.66
R1942 GND.n4839 GND.n4829 54.66
R1943 GND.n465 GND.n455 54.66
R1944 GND.n396 GND.n386 54.66
R1945 GND.n285 GND.n275 54.66
R1946 GND.t165 GND.t151 54.5194
R1947 GND.n4 GND 54.5194
R1948 GND.t252 GND.t408 54.5194
R1949 GND.n1004 GND 54.5194
R1950 GND.n6159 GND.t779 54.0356
R1951 GND.n5754 GND.t1356 53.6046
R1952 GND.t503 GND.n3927 52.9309
R1953 GND.n4099 GND.t503 52.9309
R1954 GND.n29 GND.t919 52.8576
R1955 GND.n6353 GND.t592 52.8576
R1956 GND.n7763 GND.t166 52.8576
R1957 GND.n659 GND.t1449 52.8576
R1958 GND.n702 GND.t1257 52.8576
R1959 GND.n682 GND.t394 52.8576
R1960 GND.n688 GND.t208 52.8576
R1961 GND.n6303 GND.t1504 52.8576
R1962 GND.n6274 GND.t839 52.8576
R1963 GND.n6253 GND.t1250 52.8576
R1964 GND.n6233 GND.t418 52.8576
R1965 GND.n6239 GND.t494 52.8576
R1966 GND.n7652 GND.n174 51.4154
R1967 GND.n7652 GND.n176 51.4154
R1968 GND.n7652 GND.n177 51.4154
R1969 GND.n7652 GND.n178 51.4154
R1970 GND.n7652 GND.n180 51.4154
R1971 GND.n7652 GND.n181 51.4154
R1972 GND.n7652 GND.n168 51.4154
R1973 GND.n7652 GND.n167 51.4154
R1974 GND.n7652 GND.n166 51.4154
R1975 GND.n7652 GND.n165 51.4154
R1976 GND.n7652 GND.n169 51.4154
R1977 GND.n7652 GND.n170 51.4154
R1978 GND.n1583 GND.n1582 50.5605
R1979 GND.n2052 GND.n2050 50.5605
R1980 GND.n2052 GND.n2051 50.5605
R1981 GND.n2046 GND.n2044 50.5605
R1982 GND.n2046 GND.n2045 50.5605
R1983 GND.n2359 GND.n2357 50.5605
R1984 GND.n2359 GND.n2358 50.5605
R1985 GND.n2353 GND.n2351 50.5605
R1986 GND.n2353 GND.n2352 50.5605
R1987 GND.n2532 GND.n2530 50.5605
R1988 GND.n2532 GND.n2531 50.5605
R1989 GND.n2526 GND.n2524 50.5605
R1990 GND.n2526 GND.n2525 50.5605
R1991 GND.n2680 GND.n2678 50.5605
R1992 GND.n2680 GND.n2679 50.5605
R1993 GND.n2674 GND.n2672 50.5605
R1994 GND.n2674 GND.n2673 50.5605
R1995 GND.n2950 GND.n2948 50.5605
R1996 GND.n2950 GND.n2949 50.5605
R1997 GND.n2944 GND.n2942 50.5605
R1998 GND.n2944 GND.n2943 50.5605
R1999 GND.n125 GND.n123 50.5605
R2000 GND.n125 GND.n124 50.5605
R2001 GND.n111 GND.n109 50.5605
R2002 GND.n111 GND.n110 50.5605
R2003 GND.n1334 GND.n1332 50.5605
R2004 GND.n1334 GND.n1333 50.5605
R2005 GND.n1328 GND.n1326 50.5605
R2006 GND.n1328 GND.n1327 50.5605
R2007 GND.n5609 GND.n5607 50.5605
R2008 GND.n5609 GND.n5608 50.5605
R2009 GND.n5603 GND.n5601 50.5605
R2010 GND.n5603 GND.n5602 50.5605
R2011 GND.n1172 GND.n1170 50.5605
R2012 GND.n1172 GND.n1171 50.5605
R2013 GND.n1166 GND.n1164 50.5605
R2014 GND.n1166 GND.n1165 50.5605
R2015 GND.n3546 GND.n3544 50.5605
R2016 GND.n3546 GND.n3545 50.5605
R2017 GND.n3540 GND.n3538 50.5605
R2018 GND.n3540 GND.n3539 50.5605
R2019 GND.n5285 GND.n5283 50.5605
R2020 GND.n5285 GND.n5284 50.5605
R2021 GND.n5279 GND.n5277 50.5605
R2022 GND.n5279 GND.n5278 50.5605
R2023 GND.n4946 GND.n4944 50.5605
R2024 GND.n4946 GND.n4945 50.5605
R2025 GND.n4940 GND.n4938 50.5605
R2026 GND.n4940 GND.n4939 50.5605
R2027 GND.n3704 GND.n3702 50.5605
R2028 GND.n3704 GND.n3703 50.5605
R2029 GND.n3698 GND.n3696 50.5605
R2030 GND.n3698 GND.n3697 50.5605
R2031 GND.n3983 GND.n3981 50.5605
R2032 GND.n3983 GND.n3982 50.5605
R2033 GND.n3977 GND.n3975 50.5605
R2034 GND.n3977 GND.n3976 50.5605
R2035 GND.n3760 GND.n3758 50.5605
R2036 GND.n3760 GND.n3759 50.5605
R2037 GND.n3754 GND.n3752 50.5605
R2038 GND.n3754 GND.n3753 50.5605
R2039 GND.n3852 GND.n3851 50.5605
R2040 GND.n7651 GND.t1429 50.1906
R2041 GND.n738 GND.t334 48.3834
R2042 GND.n1003 GND 48.3834
R2043 GND.n7795 GND 47.7719
R2044 GND.n6417 GND 47.7719
R2045 GND.n4186 GND.t552 47.2072
R2046 GND.n4249 GND.n4248 47.1486
R2047 GND GND.n6116 46.7305
R2048 GND.n1359 GND.n1350 46.2978
R2049 GND.n2430 GND.n2422 46.2978
R2050 GND.n2751 GND.n2743 46.2978
R2051 GND.n7683 GND.n7675 46.2978
R2052 GND.n3024 GND.n3016 46.2978
R2053 GND.n3134 GND.n3126 46.2978
R2054 GND.n5016 GND.n5008 46.2978
R2055 GND.n4038 GND.n4030 46.2978
R2056 GND.n2107 GND.n2099 46.2978
R2057 GND.n2587 GND.n2579 46.2978
R2058 GND.n5340 GND.n5332 46.2978
R2059 GND.n3837 GND.n3829 46.2978
R2060 GND.n2863 GND.n2862 46.2978
R2061 GND.n1227 GND.n1226 46.2978
R2062 GND.n3241 GND.n3240 46.2978
R2063 GND.n3621 GND.n3613 46.2978
R2064 GND.n7572 GND 46.1266
R2065 GND.n7509 GND 46.1266
R2066 GND.n7447 GND 46.1266
R2067 GND.n4885 GND 46.1266
R2068 GND.n5209 GND 46.1266
R2069 GND.n3474 GND 46.1266
R2070 GND GND.n5456 46.1266
R2071 GND GND.n5638 46.1266
R2072 GND.n6498 GND 46.1266
R2073 GND.t625 GND.n192 43.4986
R2074 GND GND.n5647 43.3696
R2075 GND.n2840 GND.n2819 42.8187
R2076 GND.n3577 GND.n3576 42.8187
R2077 GND.n3814 GND.n3813 42.8187
R2078 GND.n3994 GND.n3993 42.8174
R2079 GND.n1407 GND.n1406 42.8174
R2080 GND.n2063 GND.n2062 42.8174
R2081 GND.n2386 GND.n2385 42.8174
R2082 GND.n2543 GND.n2542 42.8174
R2083 GND.n2707 GND.n2706 42.8174
R2084 GND.n7662 GND.n7661 42.8174
R2085 GND.n2980 GND.n2979 42.8174
R2086 GND.n3090 GND.n3089 42.8174
R2087 GND.n1183 GND.n1182 42.8174
R2088 GND.n3197 GND.n3196 42.8174
R2089 GND.n5296 GND.n5295 42.8174
R2090 GND.n4972 GND.n4971 42.8174
R2091 GND.t663 GND.n7444 42.5398
R2092 GND.t524 GND.n1347 40.7031
R2093 GND GND.n6821 40.3307
R2094 GND GND.n6975 40.3307
R2095 GND.n7075 GND 40.3307
R2096 GND.n2299 GND 40.3307
R2097 GND.n1976 GND 40.3307
R2098 GND.n1522 GND 40.3307
R2099 GND.n5754 GND.t1320 40.2035
R2100 GND.t212 GND.n4182 40.0617
R2101 GND.n4700 GND.t60 40.0617
R2102 GND.n1382 GND.n1363 39.6805
R2103 GND.n2130 GND.n2111 39.6805
R2104 GND.n2453 GND.n2434 39.6805
R2105 GND.n2610 GND.n2591 39.6805
R2106 GND.n2774 GND.n2755 39.6805
R2107 GND.n7706 GND.n7687 39.6805
R2108 GND.n3076 GND.n3057 39.6805
R2109 GND.n3177 GND.n3158 39.6805
R2110 GND.n1283 GND.n1264 39.6805
R2111 GND.n3284 GND.n3265 39.6805
R2112 GND.n5363 GND.n5344 39.6805
R2113 GND.n5039 GND.n5020 39.6805
R2114 GND.n3644 GND.n3625 39.6805
R2115 GND.n4083 GND.n4064 39.6805
R2116 GND.n3901 GND.n3877 39.6805
R2117 GND.n6209 GND.n6199 39.2858
R2118 GND.n23 GND.n22 39.2858
R2119 GND.n7781 GND.n7780 39.2858
R2120 GND.n6485 GND.n6475 39.2858
R2121 GND.n6489 GND.n6488 39.2858
R2122 GND.n675 GND.n674 39.2858
R2123 GND.n6345 GND.n6344 39.2858
R2124 GND.n6321 GND.n6320 39.2858
R2125 GND.n6395 GND.n6385 39.2858
R2126 GND.n6399 GND.n6398 39.2858
R2127 GND.n6290 GND.n6289 39.2858
R2128 GND.n19 GND.n6 38.7881
R2129 GND.n7777 GND.n7754 38.7881
R2130 GND.n671 GND.n652 38.7881
R2131 GND.n6341 GND.n6328 38.7881
R2132 GND.n6317 GND.n6294 38.7881
R2133 GND.n6286 GND.n6267 38.7881
R2134 GND.n12 GND.t426 38.7697
R2135 GND.n9 GND.t790 38.7697
R2136 GND.n7760 GND.t488 38.7697
R2137 GND.n7757 GND.t152 38.7697
R2138 GND.n6334 GND.t170 38.7697
R2139 GND.n6331 GND.t837 38.7697
R2140 GND.n6300 GND.t164 38.7697
R2141 GND.n6297 GND.t409 38.7697
R2142 GND.n692 GND.n690 38.7523
R2143 GND.n6243 GND.n6241 38.7523
R2144 GND.t751 GND.n6226 38.597
R2145 GND.n31 GND.t398 38.5719
R2146 GND.n31 GND.t630 38.5719
R2147 GND.n6355 GND.t893 38.5719
R2148 GND.n6355 GND.t160 38.5719
R2149 GND.n7762 GND.t917 38.5719
R2150 GND.n7762 GND.t221 38.5719
R2151 GND.n657 GND.t83 38.5719
R2152 GND.n657 GND.t168 38.5719
R2153 GND.n705 GND.t1080 38.5719
R2154 GND.n705 GND.t1396 38.5719
R2155 GND.n680 GND.t66 38.5719
R2156 GND.n680 GND.t1447 38.5719
R2157 GND.n685 GND.t604 38.5719
R2158 GND.n685 GND.t1254 38.5719
R2159 GND.n6302 GND.t590 38.5719
R2160 GND.n6302 GND.t253 38.5719
R2161 GND.n6272 GND.t930 38.5719
R2162 GND.n6272 GND.t1503 38.5719
R2163 GND.n6256 GND.t245 38.5719
R2164 GND.n6256 GND.t244 38.5719
R2165 GND.n6231 GND.t25 38.5719
R2166 GND.n6231 GND.t495 38.5719
R2167 GND.n6236 GND.t891 38.5719
R2168 GND.n6236 GND.t802 38.5719
R2169 GND.n833 GND.t284 36.9992
R2170 GND.t1066 GND.n5912 36.8926
R2171 GND.n5913 GND.t1016 36.8926
R2172 GND.t122 GND.t500 36.3723
R2173 GND.t528 GND.t1089 36.3723
R2174 GND.t831 GND.t1415 36.3723
R2175 GND.t429 GND.t1239 36.3723
R2176 GND.t129 GND.t1230 36.3723
R2177 GND.t572 GND.t249 36.3723
R2178 GND.t431 GND.t1399 36.3723
R2179 GND.t805 GND.t108 36.3723
R2180 GND.t105 GND.t947 36.3723
R2181 GND.t530 GND.t657 36.3723
R2182 GND.t834 GND.t1419 36.3723
R2183 GND.t510 GND.t427 36.3723
R2184 GND.t522 GND.t1241 36.3723
R2185 GND.t574 GND.t874 36.3723
R2186 GND.t829 GND.t1225 36.3723
R2187 GND.t102 GND.n4185 36.3719
R2188 GND.n2416 GND.n2415 35.6515
R2189 GND.n2737 GND.n2736 35.6515
R2190 GND.n7669 GND.n7668 35.6515
R2191 GND.n3120 GND.n3119 35.6515
R2192 GND.n3234 GND.n3233 35.6515
R2193 GND.n5002 GND.n5001 35.6515
R2194 GND.n3823 GND.n3822 35.6515
R2195 GND.n7806 GND.n7805 34.6358
R2196 GND.n38 GND.n37 34.6358
R2197 GND.n41 GND.n26 34.6358
R2198 GND.n45 GND.n26 34.6358
R2199 GND.n46 GND.n45 34.6358
R2200 GND.n6362 GND.n6361 34.6358
R2201 GND.n6365 GND.n6350 34.6358
R2202 GND.n6369 GND.n6350 34.6358
R2203 GND.n6370 GND.n6369 34.6358
R2204 GND.n994 GND.n993 34.6358
R2205 GND.n15 GND.n14 34.6358
R2206 GND.n14 GND.n7 34.6358
R2207 GND.n22 GND.n7 34.6358
R2208 GND.n18 GND.n17 34.6358
R2209 GND.n19 GND.n18 34.6358
R2210 GND.n7773 GND.n7772 34.6358
R2211 GND.n7772 GND.n7755 34.6358
R2212 GND.n7780 GND.n7755 34.6358
R2213 GND.n7776 GND.n7775 34.6358
R2214 GND.n7777 GND.n7776 34.6358
R2215 GND.n6485 GND.n6484 34.6358
R2216 GND.n6488 GND.n6476 34.6358
R2217 GND.n674 GND.n653 34.6358
R2218 GND.n667 GND.n666 34.6358
R2219 GND.n699 GND.n698 34.6358
R2220 GND.n6448 GND.n6447 34.6358
R2221 GND.n6442 GND.n6441 34.6358
R2222 GND.n6430 GND.n6429 34.6358
R2223 GND.n6337 GND.n6336 34.6358
R2224 GND.n6336 GND.n6329 34.6358
R2225 GND.n6344 GND.n6329 34.6358
R2226 GND.n6340 GND.n6339 34.6358
R2227 GND.n6341 GND.n6340 34.6358
R2228 GND.n6313 GND.n6312 34.6358
R2229 GND.n6312 GND.n6295 34.6358
R2230 GND.n6320 GND.n6295 34.6358
R2231 GND.n6316 GND.n6315 34.6358
R2232 GND.n6317 GND.n6316 34.6358
R2233 GND.n6395 GND.n6394 34.6358
R2234 GND.n6398 GND.n6386 34.6358
R2235 GND.n6289 GND.n6268 34.6358
R2236 GND.n6282 GND.n6281 34.6358
R2237 GND.n6250 GND.n6249 34.6358
R2238 GND.n545 GND.n544 34.6358
R2239 GND.n539 GND.n538 34.6358
R2240 GND.n527 GND.n526 34.6358
R2241 GND.n6107 GND.n6106 34.6358
R2242 GND.t1473 GND.n6117 34.4331
R2243 GND.n927 GND.t456 34.1532
R2244 GND.n1560 GND.n1559 34.1229
R2245 GND.n6436 GND.n6435 33.8829
R2246 GND.n533 GND.n532 33.8829
R2247 GND.n1196 GND.t1405 33.462
R2248 GND.n1196 GND.t1512 33.462
R2249 GND.n3209 GND.t894 33.462
R2250 GND.n3209 GND.t1549 33.462
R2251 GND.n4000 GND.t888 33.462
R2252 GND.n4000 GND.t795 33.462
R2253 GND.n5302 GND.t602 33.462
R2254 GND.n5302 GND.t46 33.462
R2255 GND.n2986 GND.t871 33.462
R2256 GND.n2986 GND.t577 33.462
R2257 GND.n2841 GND.t486 33.462
R2258 GND.n2841 GND.t251 33.462
R2259 GND.n2549 GND.t1487 33.462
R2260 GND.n2549 GND.t57 33.462
R2261 GND.n2069 GND.t1492 33.462
R2262 GND.n2069 GND.t434 33.462
R2263 GND.n1400 GND.t162 33.462
R2264 GND.n1400 GND.t247 33.462
R2265 GND.n1351 GND.t206 33.462
R2266 GND.n1351 GND.t74 33.462
R2267 GND.n2100 GND.t786 33.462
R2268 GND.n2100 GND.t1090 33.462
R2269 GND.n2391 GND.t926 33.462
R2270 GND.n2391 GND.t825 33.462
R2271 GND.n2423 GND.t18 33.462
R2272 GND.n2423 GND.t195 33.462
R2273 GND.n2580 GND.t855 33.462
R2274 GND.n2580 GND.t1240 33.462
R2275 GND.n2712 GND.t676 33.462
R2276 GND.n2712 GND.t1095 33.462
R2277 GND.n2744 GND.t948 33.462
R2278 GND.n2744 GND.t1231 33.462
R2279 GND.n2825 GND.t924 33.462
R2280 GND.n2825 GND.t1506 33.462
R2281 GND.n156 GND.t407 33.462
R2282 GND.n156 GND.t483 33.462
R2283 GND.n7676 GND.t561 33.462
R2284 GND.n7676 GND.t1400 33.462
R2285 GND.n3017 GND.t1553 33.462
R2286 GND.n3017 GND.t110 33.462
R2287 GND.n3095 GND.t440 33.462
R2288 GND.n3095 GND.t1249 33.462
R2289 GND.n3127 GND.t631 33.462
R2290 GND.n3127 GND.t112 33.462
R2291 GND.n1184 GND.t690 33.462
R2292 GND.n1184 GND.t733 33.462
R2293 GND.n3198 GND.t586 33.462
R2294 GND.n3198 GND.t1418 33.462
R2295 GND.n5333 GND.t411 33.462
R2296 GND.n5333 GND.t428 33.462
R2297 GND.n4977 GND.t750 33.462
R2298 GND.n4977 GND.t198 33.462
R2299 GND.n5009 GND.t925 33.462
R2300 GND.n5009 GND.t1242 33.462
R2301 GND.n3583 GND.t1567 33.462
R2302 GND.n3583 GND.t808 33.462
R2303 GND.n3614 GND.t1432 33.462
R2304 GND.n3614 GND.t875 33.462
R2305 GND.n4031 GND.t873 33.462
R2306 GND.n4031 GND.t1088 33.462
R2307 GND.n3791 GND.t225 33.462
R2308 GND.n3791 GND.t22 33.462
R2309 GND.n3830 GND.t1406 33.462
R2310 GND.n3830 GND.t179 33.462
R2311 GND.n7372 GND.t1211 32.2518
R2312 GND.n7771 GND.n7770 32.1329
R2313 GND.n6311 GND.n6310 32.1329
R2314 GND.n7652 GND.n7651 31.7876
R2315 GND.n1506 GND.n1505 30.7897
R2316 GND.n1928 GND.n1927 30.7897
R2317 GND.n2251 GND.n2250 30.7897
R2318 GND.n7177 GND.n7176 30.7897
R2319 GND.n7011 GND.n7010 30.7897
R2320 GND.n6857 GND.n6856 30.7897
R2321 GND.n6703 GND.n6702 30.7897
R2322 GND.n6633 GND.n6632 30.7897
R2323 GND.n5530 GND.n5529 30.7897
R2324 GND.n1096 GND.n1095 30.7897
R2325 GND.n3404 GND.n3403 30.7897
R2326 GND.n5164 GND.n5163 30.7897
R2327 GND.n4840 GND.n4839 30.7897
R2328 GND.n466 GND.n465 30.7897
R2329 GND.n397 GND.n396 30.7897
R2330 GND.n286 GND.n285 30.7897
R2331 GND.n1887 GND.n1881 30.5561
R2332 GND.n5753 GND.t1372 29.036
R2333 GND.n7446 GND.n7445 29.0202
R2334 GND.n3958 GND.n3953 28.9511
R2335 GND.n5260 GND.n5255 28.9511
R2336 GND.n3521 GND.n3516 28.9511
R2337 GND.n1145 GND.n1140 28.9511
R2338 GND.n5584 GND.n5579 28.9511
R2339 GND.n1309 GND.n1304 28.9511
R2340 GND.n2923 GND.n2918 28.9511
R2341 GND.n2507 GND.n2502 28.9511
R2342 GND.n2027 GND.n2022 28.9511
R2343 GND.n1567 GND.n1562 28.9511
R2344 GND.n2346 GND.n2341 28.9511
R2345 GND.n2667 GND.n2662 28.9511
R2346 GND.n104 GND.n99 28.9511
R2347 GND.n4933 GND.n4928 28.9511
R2348 GND.n3691 GND.n3686 28.9511
R2349 GND.n3747 GND.n3742 28.9511
R2350 GND.n1887 GND.n1886 28.8988
R2351 GND.n2212 GND.n2211 28.8988
R2352 GND.n7143 GND.n7142 28.8988
R2353 GND.n616 GND.n615 28.8988
R2354 GND.n626 GND.n625 28.8988
R2355 GND.n636 GND.n635 28.8988
R2356 GND.n643 GND.n642 28.8988
R2357 GND.n5555 GND.n5554 28.8988
R2358 GND.n3433 GND.n3432 28.8988
R2359 GND.n3339 GND.n3338 28.8988
R2360 GND.n5120 GND.n5119 28.8988
R2361 GND.n4799 GND.n4798 28.8988
R2362 GND.n422 GND.n421 28.8988
R2363 GND.n311 GND.n310 28.8988
R2364 GND.n210 GND.n209 28.8988
R2365 GND.n1495 GND.n1494 28.8193
R2366 GND.n1912 GND.n1911 28.8193
R2367 GND.n2235 GND.n2234 28.8193
R2368 GND.n7161 GND.n7160 28.8193
R2369 GND.n6995 GND.n6994 28.8193
R2370 GND.n6841 GND.n6840 28.8193
R2371 GND.n6687 GND.n6686 28.8193
R2372 GND.n6617 GND.n6616 28.8193
R2373 GND.n5514 GND.n5513 28.8193
R2374 GND.n1080 GND.n1079 28.8193
R2375 GND.n3388 GND.n3387 28.8193
R2376 GND.n5148 GND.n5147 28.8193
R2377 GND.n4824 GND.n4823 28.8193
R2378 GND.n450 GND.n449 28.8193
R2379 GND.n381 GND.n380 28.8193
R2380 GND.n270 GND.n269 28.8193
R2381 GND.n558 GND.n557 27.8593
R2382 GND.n555 GND.n554 27.8593
R2383 GND.n7326 GND.n7325 27.8593
R2384 GND.n7244 GND.n7243 27.8593
R2385 GND.n5824 GND.n5823 27.8593
R2386 GND.n5717 GND.n5716 27.8593
R2387 GND.n6148 GND.n6147 27.8593
R2388 GND.n883 GND.n882 27.8593
R2389 GND.n871 GND.n870 27.8593
R2390 GND.n784 GND.n783 27.8593
R2391 GND.n772 GND.n771 27.8593
R2392 GND.n6034 GND.n6033 27.8593
R2393 GND.n5851 GND.n5850 27.8593
R2394 GND.n5953 GND.n5952 27.8593
R2395 GND.n5871 GND.n5870 27.8593
R2396 GND.n29 GND.t1484 27.5691
R2397 GND.n6353 GND.t678 27.5691
R2398 GND.n7763 GND.t876 27.5691
R2399 GND.n659 GND.t401 27.5691
R2400 GND.n702 GND.t704 27.5691
R2401 GND.n682 GND.t508 27.5691
R2402 GND.n688 GND.t1086 27.5691
R2403 GND.n6303 GND.t1505 27.5691
R2404 GND.n6274 GND.t1511 27.5691
R2405 GND.n6253 GND.t596 27.5691
R2406 GND.n6233 GND.t556 27.5691
R2407 GND.n6239 GND.t220 27.5691
R2408 GND.n6207 GND.n6198 27.1064
R2409 GND GND.n7786 26.9763
R2410 GND.n4612 GND.t502 26.8697
R2411 GND.n7810 GND.t236 26.8576
R2412 GND.n986 GND.t784 26.8576
R2413 GND.n6099 GND.t1414 26.8576
R2414 GND.n5655 GND.t1368 26.8025
R2415 GND.n1956 GND.n1955 26.7111
R2416 GND.n1052 GND.n1051 26.7111
R2417 GND.n5479 GND.n5478 26.7111
R2418 GND.n235 GND.n234 26.7111
R2419 GND.n4865 GND.n4864 26.7111
R2420 GND.n5189 GND.n5188 26.7111
R2421 GND.n3362 GND.n3361 26.7111
R2422 GND.n6740 GND.n6739 26.7111
R2423 GND.n7048 GND.n7047 26.7111
R2424 GND.n2279 GND.n2278 26.7111
R2425 GND.n7209 GND.n7208 26.7111
R2426 GND.n6894 GND.n6893 26.7111
R2427 GND.n6582 GND.n6581 26.7111
R2428 GND.n494 GND.n493 26.7111
R2429 GND.n346 GND.n345 26.7111
R2430 GND.n7643 GND.n7642 26.7111
R2431 GND.n6227 GND.t743 26.1036
R2432 GND.n47 GND.t554 25.9346
R2433 GND.n6371 GND.t853 25.9346
R2434 GND.t721 GND.t723 25.66
R2435 GND.t723 GND.t725 25.66
R2436 GND.t725 GND.t728 25.66
R2437 GND.t255 GND.t257 25.66
R2438 GND.t257 GND.t260 25.66
R2439 GND.t260 GND.t262 25.66
R2440 GND.t694 GND.t696 25.66
R2441 GND.t696 GND.t699 25.66
R2442 GND.t699 GND.t701 25.66
R2443 GND.t900 GND.t902 25.66
R2444 GND.t902 GND.t896 25.66
R2445 GND.t896 GND.t898 25.66
R2446 GND.t146 GND.t148 25.66
R2447 GND.t148 GND.t142 25.66
R2448 GND.t142 GND.t144 25.66
R2449 GND.t516 GND.t518 25.66
R2450 GND.t518 GND.t520 25.66
R2451 GND.t520 GND.t513 25.66
R2452 GND.t1386 GND.t1393 25.66
R2453 GND.t1389 GND.t1386 25.66
R2454 GND.t1391 GND.t1389 25.66
R2455 GND.t687 GND.t685 25.66
R2456 GND.t681 GND.t687 25.66
R2457 GND.t683 GND.t681 25.66
R2458 GND.t2 GND.t4 25.66
R2459 GND.t4 GND.t7 25.66
R2460 GND.t7 GND.t9 25.66
R2461 GND.n4186 GND.t26 25.4195
R2462 GND.n3989 GND.n3970 25.0358
R2463 GND.n5291 GND.n5272 25.0358
R2464 GND.n3552 GND.n3533 25.0358
R2465 GND.n1178 GND.n1159 25.0358
R2466 GND.n5615 GND.n5596 25.0358
R2467 GND.n1340 GND.n1321 25.0358
R2468 GND.n2956 GND.n2937 25.0358
R2469 GND.n2538 GND.n2519 25.0358
R2470 GND.n2058 GND.n2039 25.0358
R2471 GND.n1587 GND.n1577 25.0358
R2472 GND.n2377 GND.n2376 25.0358
R2473 GND.n2698 GND.n2697 25.0358
R2474 GND.n143 GND.n142 25.0358
R2475 GND.n4964 GND.n4963 25.0358
R2476 GND.n3722 GND.n3721 25.0358
R2477 GND.n3778 GND.n3777 25.0358
R2478 GND.n563 GND.t610 24.9236
R2479 GND.n563 GND.t612 24.9236
R2480 GND.n7378 GND.t1544 24.9236
R2481 GND.n7378 GND.t1524 24.9236
R2482 GND.n600 GND.t1532 24.9236
R2483 GND.n600 GND.t1542 24.9236
R2484 GND.n594 GND.t1538 24.9236
R2485 GND.n594 GND.t1546 24.9236
R2486 GND.n590 GND.t1526 24.9236
R2487 GND.n590 GND.t1540 24.9236
R2488 GND.n584 GND.t1548 24.9236
R2489 GND.n584 GND.t1528 24.9236
R2490 GND.n578 GND.t1534 24.9236
R2491 GND.n578 GND.t1518 24.9236
R2492 GND.n572 GND.t1522 24.9236
R2493 GND.n572 GND.t1536 24.9236
R2494 GND.n7425 GND.t1206 24.9236
R2495 GND.n7425 GND.t1104 24.9236
R2496 GND.n7417 GND.t1184 24.9236
R2497 GND.n7417 GND.t1210 24.9236
R2498 GND.n7410 GND.t1142 24.9236
R2499 GND.n7410 GND.t1164 24.9236
R2500 GND.n7406 GND.t1198 24.9236
R2501 GND.n7406 GND.t1132 24.9236
R2502 GND.n7400 GND.t1168 24.9236
R2503 GND.n7400 GND.t1110 24.9236
R2504 GND.n7394 GND.t1192 24.9236
R2505 GND.n7394 GND.t1220 24.9236
R2506 GND.n7388 GND.t1152 24.9236
R2507 GND.n7388 GND.t1176 24.9236
R2508 GND.n7330 GND.t1160 24.9236
R2509 GND.n7330 GND.t1190 24.9236
R2510 GND.n7337 GND.t1126 24.9236
R2511 GND.n7337 GND.t1212 24.9236
R2512 GND.n7363 GND.t1122 24.9236
R2513 GND.n7363 GND.t1186 24.9236
R2514 GND.n7359 GND.t1214 24.9236
R2515 GND.n7359 GND.t1144 24.9236
R2516 GND.n7353 GND.t1170 24.9236
R2517 GND.n7353 GND.t1202 24.9236
R2518 GND.n7347 GND.t1146 24.9236
R2519 GND.n7347 GND.t1172 24.9236
R2520 GND.n7341 GND.t1118 24.9236
R2521 GND.n7341 GND.t1140 24.9236
R2522 GND.n7246 GND.t1182 24.9236
R2523 GND.n7246 GND.t1208 24.9236
R2524 GND.n7289 GND.t1106 24.9236
R2525 GND.n7289 GND.t1162 24.9236
R2526 GND.n7296 GND.t1196 24.9236
R2527 GND.n7296 GND.t1128 24.9236
R2528 GND.n7300 GND.t1166 24.9236
R2529 GND.n7300 GND.t1200 24.9236
R2530 GND.n7306 GND.t1136 24.9236
R2531 GND.n7306 GND.t1216 24.9236
R2532 GND.n7312 GND.t1148 24.9236
R2533 GND.n7312 GND.t1174 24.9236
R2534 GND.n7318 GND.t1222 24.9236
R2535 GND.n7318 GND.t1154 24.9236
R2536 GND.n7232 GND.t1138 24.9236
R2537 GND.n7232 GND.t1224 24.9236
R2538 GND.n7237 GND.t1116 24.9236
R2539 GND.n7237 GND.t1108 24.9236
R2540 GND.n7279 GND.t1130 24.9236
R2541 GND.n7279 GND.t1156 24.9236
R2542 GND.n7274 GND.t1098 24.9236
R2543 GND.n7274 GND.t1134 24.9236
R2544 GND.n7268 GND.t1204 24.9236
R2545 GND.n7268 GND.t1100 24.9236
R2546 GND.n7262 GND.t1124 24.9236
R2547 GND.n7262 GND.t1188 24.9236
R2548 GND.n7256 GND.t1218 24.9236
R2549 GND.n7256 GND.t1150 24.9236
R2550 GND.n1443 GND.t912 24.9236
R2551 GND.n1443 GND.t913 24.9236
R2552 GND.n1535 GND.t1428 24.9236
R2553 GND.n1535 GND.t1422 24.9236
R2554 GND.n1027 GND.t177 24.9236
R2555 GND.n1027 GND.t178 24.9236
R2556 GND.n5626 GND.t688 24.9236
R2557 GND.n5626 GND.t682 24.9236
R2558 GND.n6535 GND.t563 24.9236
R2559 GND.n6535 GND.t564 24.9236
R2560 GND.n6520 GND.t5 24.9236
R2561 GND.n6520 GND.t8 24.9236
R2562 GND.n7546 GND.t1559 24.9236
R2563 GND.n7546 GND.t1556 24.9236
R2564 GND.n7531 GND.t258 24.9236
R2565 GND.n7531 GND.t261 24.9236
R2566 GND.n5083 GND.t648 24.9236
R2567 GND.n5083 GND.t649 24.9236
R2568 GND.n5231 GND.t149 24.9236
R2569 GND.n5231 GND.t143 24.9236
R2570 GND.n3294 GND.t42 24.9236
R2571 GND.n3294 GND.t43 24.9236
R2572 GND.n3496 GND.t519 24.9236
R2573 GND.n3496 GND.t521 24.9236
R2574 GND.n3449 GND.t815 24.9236
R2575 GND.n3449 GND.t811 24.9236
R2576 GND.n5444 GND.t1387 24.9236
R2577 GND.n5444 GND.t1390 24.9236
R2578 GND.n6789 GND.t182 24.9236
R2579 GND.n6789 GND.t183 24.9236
R2580 GND.n6809 GND.t1441 24.9236
R2581 GND.n6809 GND.t1444 24.9236
R2582 GND.n7112 GND.t541 24.9236
R2583 GND.n7112 GND.t542 24.9236
R2584 GND.n7097 GND.t140 24.9236
R2585 GND.n7097 GND.t134 24.9236
R2586 GND.n1849 GND.t638 24.9236
R2587 GND.n1849 GND.t634 24.9236
R2588 GND.n1998 GND.t846 24.9236
R2589 GND.n1998 GND.t849 24.9236
R2590 GND.n2193 GND.t642 24.9236
R2591 GND.n2193 GND.t643 24.9236
R2592 GND.n2321 GND.t98 24.9236
R2593 GND.n2321 GND.t101 24.9236
R2594 GND.n6943 GND.t115 24.9236
R2595 GND.n6943 GND.t116 24.9236
R2596 GND.n6963 GND.t941 24.9236
R2597 GND.n6963 GND.t944 24.9236
R2598 GND.n73 GND.t205 24.9236
R2599 GND.n73 GND.t201 24.9236
R2600 GND.n52 GND.t713 24.9236
R2601 GND.n52 GND.t716 24.9236
R2602 GND.n4762 GND.t81 24.9236
R2603 GND.n4762 GND.t77 24.9236
R2604 GND.n4907 GND.t903 24.9236
R2605 GND.n4907 GND.t897 24.9236
R2606 GND.n7484 GND.t239 24.9236
R2607 GND.n7484 GND.t240 24.9236
R2608 GND.n7469 GND.t697 24.9236
R2609 GND.n7469 GND.t700 24.9236
R2610 GND.n7609 GND.t1409 24.9236
R2611 GND.n7609 GND.t1411 24.9236
R2612 GND.n7594 GND.t724 24.9236
R2613 GND.n7594 GND.t726 24.9236
R2614 GND.n6213 GND.t746 24.9236
R2615 GND.n6213 GND.t748 24.9236
R2616 GND.n5816 GND.t1315 24.9236
R2617 GND.n5816 GND.t1349 24.9236
R2618 GND.n5810 GND.t1301 24.9236
R2619 GND.n5810 GND.t1263 24.9236
R2620 GND.n5804 GND.t1287 24.9236
R2621 GND.n5804 GND.t1343 24.9236
R2622 GND.n5800 GND.t1375 24.9236
R2623 GND.n5800 GND.t1275 24.9236
R2624 GND.n5794 GND.t1327 24.9236
R2625 GND.n5794 GND.t1379 24.9236
R2626 GND.n5786 GND.t1305 24.9236
R2627 GND.n5786 GND.t1331 24.9236
R2628 GND.n5780 GND.t1363 24.9236
R2629 GND.n5780 GND.t1299 24.9236
R2630 GND.n5770 GND.t1367 24.9236
R2631 GND.n5770 GND.t1281 24.9236
R2632 GND.n5764 GND.t1339 24.9236
R2633 GND.n5764 GND.t1371 24.9236
R2634 GND.n5757 GND.t1271 24.9236
R2635 GND.n5757 GND.t1321 24.9236
R2636 GND.n5688 GND.t1357 24.9236
R2637 GND.n5688 GND.t1293 24.9236
R2638 GND.n5697 GND.t1325 24.9236
R2639 GND.n5697 GND.t1291 24.9236
R2640 GND.n5703 GND.t1353 24.9236
R2641 GND.n5703 GND.t1383 24.9236
R2642 GND.n5709 GND.t1309 24.9236
R2643 GND.n5709 GND.t1335 24.9236
R2644 GND.n5721 GND.t1365 24.9236
R2645 GND.n5721 GND.t1267 24.9236
R2646 GND.n5727 GND.t1317 24.9236
R2647 GND.n5727 GND.t1285 24.9236
R2648 GND.n5747 GND.t1341 24.9236
R2649 GND.n5747 GND.t1373 24.9236
R2650 GND.n5742 GND.t1289 24.9236
R2651 GND.n5742 GND.t1345 24.9236
R2652 GND.n5735 GND.t1377 24.9236
R2653 GND.n5735 GND.t1303 24.9236
R2654 GND.n5650 GND.t1329 24.9236
R2655 GND.n5650 GND.t1361 24.9236
R2656 GND.n6139 GND.t1307 24.9236
R2657 GND.n6139 GND.t1333 24.9236
R2658 GND.n6152 GND.t760 24.9236
R2659 GND.n6152 GND.t770 24.9236
R2660 GND.n6162 GND.t780 24.9236
R2661 GND.n6162 GND.t758 24.9236
R2662 GND.n6169 GND.t772 24.9236
R2663 GND.n6169 GND.t782 24.9236
R2664 GND.n6173 GND.t762 24.9236
R2665 GND.n6173 GND.t768 24.9236
R2666 GND.n6179 GND.t778 24.9236
R2667 GND.n6179 GND.t774 24.9236
R2668 GND.n6185 GND.t756 24.9236
R2669 GND.n6185 GND.t766 24.9236
R2670 GND.n6192 GND.t776 24.9236
R2671 GND.n6192 GND.t752 24.9236
R2672 GND.n5659 GND.t1297 24.9236
R2673 GND.n5659 GND.t1369 24.9236
R2674 GND.n5667 GND.t1269 24.9236
R2675 GND.n5667 GND.t1319 24.9236
R2676 GND.n5673 GND.t1355 24.9236
R2677 GND.n5673 GND.t1273 24.9236
R2678 GND.n5677 GND.t1323 24.9236
R2679 GND.n5677 GND.t1359 24.9236
R2680 GND.n5843 GND.t1347 24.9236
R2681 GND.n5843 GND.t1381 24.9236
R2682 GND.n5837 GND.t1277 24.9236
R2683 GND.n5837 GND.t1351 24.9236
R2684 GND.n5831 GND.t1385 24.9236
R2685 GND.n5831 GND.t1311 24.9236
R2686 GND.n973 GND.t92 24.9236
R2687 GND.n973 GND.t86 24.9236
R2688 GND.n717 GND.t477 24.9236
R2689 GND.n717 GND.t457 24.9236
R2690 GND.n933 GND.t465 24.9236
R2691 GND.n933 GND.t475 24.9236
R2692 GND.n939 GND.t471 24.9236
R2693 GND.n939 GND.t479 24.9236
R2694 GND.n943 GND.t459 24.9236
R2695 GND.n943 GND.t473 24.9236
R2696 GND.n949 GND.t481 24.9236
R2697 GND.n949 GND.t461 24.9236
R2698 GND.n955 GND.t467 24.9236
R2699 GND.n955 GND.t451 24.9236
R2700 GND.n961 GND.t455 24.9236
R2701 GND.n961 GND.t469 24.9236
R2702 GND.n875 GND.t385 24.9236
R2703 GND.n875 GND.t283 24.9236
R2704 GND.n920 GND.t363 24.9236
R2705 GND.n920 GND.t389 24.9236
R2706 GND.n913 GND.t321 24.9236
R2707 GND.n913 GND.t343 24.9236
R2708 GND.n909 GND.t379 24.9236
R2709 GND.n909 GND.t311 24.9236
R2710 GND.n903 GND.t347 24.9236
R2711 GND.n903 GND.t289 24.9236
R2712 GND.n897 GND.t373 24.9236
R2713 GND.n897 GND.t271 24.9236
R2714 GND.n891 GND.t331 24.9236
R2715 GND.n891 GND.t355 24.9236
R2716 GND.n788 GND.t339 24.9236
R2717 GND.n788 GND.t371 24.9236
R2718 GND.n721 GND.t305 24.9236
R2719 GND.n721 GND.t391 24.9236
R2720 GND.n840 GND.t301 24.9236
R2721 GND.n840 GND.t367 24.9236
R2722 GND.n844 GND.t393 24.9236
R2723 GND.n844 GND.t323 24.9236
R2724 GND.n850 GND.t349 24.9236
R2725 GND.n850 GND.t365 24.9236
R2726 GND.n856 GND.t325 24.9236
R2727 GND.n856 GND.t351 24.9236
R2728 GND.n862 GND.t297 24.9236
R2729 GND.n862 GND.t319 24.9236
R2730 GND.n776 GND.t361 24.9236
R2731 GND.n776 GND.t387 24.9236
R2732 GND.n827 GND.t285 24.9236
R2733 GND.n827 GND.t341 24.9236
R2734 GND.n820 GND.t377 24.9236
R2735 GND.n820 GND.t307 24.9236
R2736 GND.n816 GND.t345 24.9236
R2737 GND.n816 GND.t381 24.9236
R2738 GND.n810 GND.t315 24.9236
R2739 GND.n810 GND.t267 24.9236
R2740 GND.n804 GND.t327 24.9236
R2741 GND.n804 GND.t353 24.9236
R2742 GND.n798 GND.t273 24.9236
R2743 GND.n798 GND.t333 24.9236
R2744 GND.n725 GND.t317 24.9236
R2745 GND.n725 GND.t275 24.9236
R2746 GND.n730 GND.t295 24.9236
R2747 GND.n730 GND.t287 24.9236
R2748 GND.n741 GND.t309 24.9236
R2749 GND.n741 GND.t335 24.9236
R2750 GND.n746 GND.t277 24.9236
R2751 GND.n746 GND.t313 24.9236
R2752 GND.n752 GND.t383 24.9236
R2753 GND.n752 GND.t279 24.9236
R2754 GND.n758 GND.t303 24.9236
R2755 GND.n758 GND.t369 24.9236
R2756 GND.n764 GND.t269 24.9236
R2757 GND.n764 GND.t329 24.9236
R2758 GND.n6086 GND.t55 24.9236
R2759 GND.n6086 GND.t49 24.9236
R2760 GND.n6038 GND.t1462 24.9236
R2761 GND.n6038 GND.t1474 24.9236
R2762 GND.n6046 GND.t1482 24.9236
R2763 GND.n6046 GND.t1460 24.9236
R2764 GND.n6052 GND.t1456 24.9236
R2765 GND.n6052 GND.t1464 24.9236
R2766 GND.n6056 GND.t1476 24.9236
R2767 GND.n6056 GND.t1458 24.9236
R2768 GND.n6062 GND.t1466 24.9236
R2769 GND.n6062 GND.t1478 24.9236
R2770 GND.n6068 GND.t1452 24.9236
R2771 GND.n6068 GND.t1468 24.9236
R2772 GND.n6074 GND.t1472 24.9236
R2773 GND.n6074 GND.t1454 24.9236
R2774 GND.n6124 GND.t989 24.9236
R2775 GND.n6124 GND.t1015 24.9236
R2776 GND.n5852 GND.t967 24.9236
R2777 GND.n5852 GND.t993 24.9236
R2778 GND.n6004 GND.t1053 24.9236
R2779 GND.n6004 GND.t1075 24.9236
R2780 GND.n6008 GND.t981 24.9236
R2781 GND.n6008 GND.t1043 24.9236
R2782 GND.n6014 GND.t951 24.9236
R2783 GND.n6014 GND.t1021 24.9236
R2784 GND.n6020 GND.t975 24.9236
R2785 GND.n6020 GND.t1003 24.9236
R2786 GND.n6026 GND.t1063 24.9236
R2787 GND.n6026 GND.t959 24.9236
R2788 GND.n5957 GND.t1071 24.9236
R2789 GND.n5957 GND.t973 24.9236
R2790 GND.n5964 GND.t1037 24.9236
R2791 GND.n5964 GND.t995 24.9236
R2792 GND.n5990 GND.t1033 24.9236
R2793 GND.n5990 GND.t969 24.9236
R2794 GND.n5986 GND.t997 24.9236
R2795 GND.n5986 GND.t1055 24.9236
R2796 GND.n5980 GND.t953 24.9236
R2797 GND.n5980 GND.t985 24.9236
R2798 GND.n5974 GND.t1057 24.9236
R2799 GND.n5974 GND.t955 24.9236
R2800 GND.n5968 GND.t1029 24.9236
R2801 GND.n5968 GND.t1051 24.9236
R2802 GND.n5873 GND.t965 24.9236
R2803 GND.n5873 GND.t991 24.9236
R2804 GND.n5916 GND.t1017 24.9236
R2805 GND.n5916 GND.t1073 24.9236
R2806 GND.n5923 GND.t979 24.9236
R2807 GND.n5923 GND.t1039 24.9236
R2808 GND.n5927 GND.t1077 24.9236
R2809 GND.n5927 GND.t983 24.9236
R2810 GND.n5933 GND.t1047 24.9236
R2811 GND.n5933 GND.t999 24.9236
R2812 GND.n5939 GND.t1059 24.9236
R2813 GND.n5939 GND.t957 24.9236
R2814 GND.n5945 GND.t1005 24.9236
R2815 GND.n5945 GND.t1065 24.9236
R2816 GND.n5859 GND.t1049 24.9236
R2817 GND.n5859 GND.t1007 24.9236
R2818 GND.n5864 GND.t1027 24.9236
R2819 GND.n5864 GND.t1019 24.9236
R2820 GND.n5906 GND.t1041 24.9236
R2821 GND.n5906 GND.t1067 24.9236
R2822 GND.n5901 GND.t1009 24.9236
R2823 GND.n5901 GND.t1045 24.9236
R2824 GND.n5895 GND.t987 24.9236
R2825 GND.n5895 GND.t1011 24.9236
R2826 GND.n5889 GND.t1035 24.9236
R2827 GND.n5889 GND.t971 24.9236
R2828 GND.n5883 GND.t1001 24.9236
R2829 GND.n5883 GND.t1061 24.9236
R2830 GND.n560 GND.n559 24.4711
R2831 GND.n37 GND.n28 24.4711
R2832 GND.n6361 GND.n6352 24.4711
R2833 GND.n6197 GND.n6196 24.4711
R2834 GND.n969 GND.n968 24.4711
R2835 GND.n667 GND.n663 24.4711
R2836 GND.n693 GND.n692 24.4711
R2837 GND.n6282 GND.n6278 24.4711
R2838 GND.n6244 GND.n6243 24.4711
R2839 GND.n6082 GND.n6081 24.4711
R2840 GND.t132 GND.n2417 23.9028
R2841 GND.t104 GND.n2738 23.9028
R2842 GND.t833 GND.n7670 23.9028
R2843 GND.t11 GND.n3121 23.9028
R2844 GND.t527 GND.n3235 23.9028
R2845 GND.t107 GND.n5003 23.9028
R2846 GND.t512 GND.n3824 23.9028
R2847 GND.n699 GND.n683 23.7181
R2848 GND.n6250 GND.n6234 23.7181
R2849 GND.n1382 GND.n1381 23.4245
R2850 GND.n2130 GND.n2129 23.4245
R2851 GND.n2453 GND.n2452 23.4245
R2852 GND.n2610 GND.n2609 23.4245
R2853 GND.n2774 GND.n2773 23.4245
R2854 GND.n2875 GND.n2874 23.4245
R2855 GND.n7706 GND.n7705 23.4245
R2856 GND.n3076 GND.n3075 23.4245
R2857 GND.n3177 GND.n3176 23.4245
R2858 GND.n1283 GND.n1282 23.4245
R2859 GND.n3284 GND.n3283 23.4245
R2860 GND.n5363 GND.n5362 23.4245
R2861 GND.n5039 GND.n5038 23.4245
R2862 GND.n3644 GND.n3643 23.4245
R2863 GND.n4083 GND.n4082 23.4245
R2864 GND.n3901 GND.n3900 23.4245
R2865 GND.n33 GND.n32 22.9652
R2866 GND.n6357 GND.n6356 22.9652
R2867 GND.n7766 GND.n7765 22.9652
R2868 GND.n662 GND.n658 22.9652
R2869 GND.n706 GND.n704 22.9652
R2870 GND.n711 GND.n710 22.9652
R2871 GND.n6306 GND.n6305 22.9652
R2872 GND.n6277 GND.n6273 22.9652
R2873 GND.n6257 GND.n6255 22.9652
R2874 GND.n6262 GND.n6261 22.9652
R2875 GND.n1507 GND.n1506 22.9087
R2876 GND.n1929 GND.n1928 22.9087
R2877 GND.n2252 GND.n2251 22.9087
R2878 GND.n7178 GND.n7177 22.9087
R2879 GND.n7012 GND.n7011 22.9087
R2880 GND.n6858 GND.n6857 22.9087
R2881 GND.n6704 GND.n6703 22.9087
R2882 GND.n6634 GND.n6633 22.9087
R2883 GND.n5531 GND.n5530 22.9087
R2884 GND.n1097 GND.n1096 22.9087
R2885 GND.n3405 GND.n3404 22.9087
R2886 GND.n5165 GND.n5164 22.9087
R2887 GND.n4841 GND.n4840 22.9087
R2888 GND.n467 GND.n466 22.9087
R2889 GND.n398 GND.n397 22.9087
R2890 GND.n287 GND.n286 22.9087
R2891 GND.t126 GND.n2094 22.765
R2892 GND.t125 GND.n2574 22.765
R2893 GND.t103 GND.n2857 22.765
R2894 GND.t12 GND.n3011 22.765
R2895 GND.t128 GND.n1221 22.765
R2896 GND.t509 GND.n5327 22.765
R2897 GND.t127 GND.n3608 22.765
R2898 GND.t736 GND.n4025 22.765
R2899 GND.n1936 GND.n1935 22.5323
R2900 GND.n6726 GND.n6725 22.5323
R2901 GND.n7034 GND.n7033 22.5323
R2902 GND.n2265 GND.n2264 22.5323
R2903 GND.n7195 GND.n7194 22.5323
R2904 GND.n6880 GND.n6879 22.5323
R2905 GND.n480 GND.n479 22.5323
R2906 GND.t712 GND.t710 22.4359
R2907 GND.t715 GND.t712 22.4359
R2908 GND.t717 GND.t715 22.4359
R2909 GND.t1440 GND.t1438 22.4359
R2910 GND.t1443 GND.t1440 22.4359
R2911 GND.t1445 GND.t1443 22.4359
R2912 GND.t940 GND.t938 22.4359
R2913 GND.t943 GND.t940 22.4359
R2914 GND.t945 GND.t943 22.4359
R2915 GND.t137 GND.t139 22.4359
R2916 GND.t139 GND.t133 22.4359
R2917 GND.t133 GND.t135 22.4359
R2918 GND.t95 GND.t97 22.4359
R2919 GND.t97 GND.t100 22.4359
R2920 GND.t100 GND.t93 22.4359
R2921 GND.t843 GND.t845 22.4359
R2922 GND.t845 GND.t848 22.4359
R2923 GND.t848 GND.t850 22.4359
R2924 GND.t1425 GND.t1427 22.4359
R2925 GND.t1427 GND.t1421 22.4359
R2926 GND.t1421 GND.t1423 22.4359
R2927 GND.n252 GND.n251 22.4086
R2928 GND.n363 GND.n362 22.4086
R2929 GND.n432 GND.n431 22.4086
R2930 GND.n5130 GND.n5129 22.4086
R2931 GND.n3370 GND.n3369 22.4086
R2932 GND.n1062 GND.n1061 22.4086
R2933 GND.n5496 GND.n5495 22.4086
R2934 GND.n6599 GND.n6598 22.4086
R2935 GND.n6669 GND.n6668 22.4086
R2936 GND.n39 GND.t16 22.3257
R2937 GND.n6363 GND.t842 22.3257
R2938 GND.n6478 GND.t1434 22.3257
R2939 GND.n6480 GND.t229 22.3257
R2940 GND.n664 GND.t840 22.3257
R2941 GND.n655 GND.t549 22.3257
R2942 GND.n689 GND.t598 22.3257
R2943 GND.n6388 GND.t628 22.3257
R2944 GND.n6390 GND.t928 22.3257
R2945 GND.n6279 GND.t121 22.3257
R2946 GND.n6270 GND.t230 22.3257
R2947 GND.n6240 GND.t14 22.3257
R2948 GND.n698 GND.n686 22.2123
R2949 GND.n694 GND.n686 22.2123
R2950 GND.n6249 GND.n6237 22.2123
R2951 GND.n6245 GND.n6237 22.2123
R2952 GND GND.t15 22.1322
R2953 GND.n1959 GND.n1958 22.0429
R2954 GND.n1055 GND.n1054 22.0429
R2955 GND.n5482 GND.n5481 22.0429
R2956 GND.n238 GND.n237 22.0429
R2957 GND.n4868 GND.n4867 22.0429
R2958 GND.n5192 GND.n5191 22.0429
R2959 GND.n3365 GND.n3364 22.0429
R2960 GND.n6743 GND.n6742 22.0429
R2961 GND.n7051 GND.n7050 22.0429
R2962 GND.n2282 GND.n2281 22.0429
R2963 GND.n7212 GND.n7211 22.0429
R2964 GND.n6897 GND.n6896 22.0429
R2965 GND.n6585 GND.n6584 22.0429
R2966 GND.n497 GND.n496 22.0429
R2967 GND.n349 GND.n348 22.0429
R2968 GND.n7646 GND.n7645 22.0429
R2969 GND.n1437 GND.n1436 21.8358
R2970 GND.n1021 GND.n1020 21.8358
R2971 GND.n6529 GND.n6528 21.8358
R2972 GND.n7540 GND.n7539 21.8358
R2973 GND.n5077 GND.n5076 21.8358
R2974 GND.n3288 GND.n3287 21.8358
R2975 GND.n3443 GND.n3442 21.8358
R2976 GND.n6783 GND.n6782 21.8358
R2977 GND.n7106 GND.n7105 21.8358
R2978 GND.n1843 GND.n1842 21.8358
R2979 GND.n2178 GND.n2177 21.8358
R2980 GND.n6937 GND.n6936 21.8358
R2981 GND.n67 GND.n66 21.8358
R2982 GND.n4756 GND.n4755 21.8358
R2983 GND.n7478 GND.n7477 21.8358
R2984 GND.n7603 GND.n7602 21.8358
R2985 GND.n48 GND.n46 21.4593
R2986 GND.n6372 GND.n6370 21.4593
R2987 GND.n15 GND.n13 21.4593
R2988 GND.n17 GND.n10 21.4593
R2989 GND.n7773 GND.n7771 21.4593
R2990 GND.n7775 GND.n7758 21.4593
R2991 GND.n707 GND.n706 21.4593
R2992 GND.n710 GND.n709 21.4593
R2993 GND.n6337 GND.n6335 21.4593
R2994 GND.n6339 GND.n6332 21.4593
R2995 GND.n6313 GND.n6311 21.4593
R2996 GND.n6315 GND.n6298 21.4593
R2997 GND.n6258 GND.n6257 21.4593
R2998 GND.n6261 GND.n6260 21.4593
R2999 GND.n7795 GND.n7794 21.3675
R3000 GND.n1426 GND.n1394 20.6255
R3001 GND.n2159 GND.n2158 20.6255
R3002 GND.n2466 GND.n2461 20.6255
R3003 GND.n2633 GND.n2632 20.6255
R3004 GND.n2800 GND.n2795 20.6255
R3005 GND.n7723 GND.n7718 20.6255
R3006 GND.n3050 GND.n3049 20.6255
R3007 GND.n3148 GND.n3143 20.6255
R3008 GND.n1257 GND.n1256 20.6255
R3009 GND.n3255 GND.n3250 20.6255
R3010 GND.n5392 GND.n5391 20.6255
R3011 GND.n5059 GND.n5054 20.6255
R3012 GND.n3665 GND.n3660 20.6255
R3013 GND.n4057 GND.n4056 20.6255
R3014 GND.n3870 GND.n3869 20.6255
R3015 GND.n3927 GND.n3906 20.0775
R3016 GND.n33 GND.n28 19.9534
R3017 GND.n6357 GND.n6352 19.9534
R3018 GND.n7767 GND.n7766 19.9534
R3019 GND.n663 GND.n662 19.9534
R3020 GND.n704 GND.n679 19.9534
R3021 GND.n712 GND.n711 19.9534
R3022 GND.n6307 GND.n6306 19.9534
R3023 GND.n6278 GND.n6277 19.9534
R3024 GND.n6255 GND.n6230 19.9534
R3025 GND.n6263 GND.n6262 19.9534
R3026 GND.t157 GND.t165 19.2425
R3027 GND.t156 GND.t252 19.2425
R3028 GND.n3813 GND.n3812 19.2005
R3029 GND.n1572 GND.n1571 17.9597
R3030 GND.n5565 GND.t417 17.475
R3031 GND.n6550 GND.t817 17.475
R3032 GND.n7561 GND.t1486 17.475
R3033 GND.n5110 GND.t223 17.475
R3034 GND.n3331 GND.t497 17.475
R3035 GND.n3464 GND.t740 17.475
R3036 GND.n6803 GND.t32 17.475
R3037 GND.n7127 GND.t1436 17.475
R3038 GND.n1876 GND.t68 17.475
R3039 GND.n2202 GND.t923 17.475
R3040 GND.n6957 GND.t1256 17.475
R3041 GND.n6657 GND.t38 17.475
R3042 GND.n4789 GND.t30 17.475
R3043 GND.n7499 GND.t438 17.475
R3044 GND.n7624 GND.t1430 17.475
R3045 GND.n1459 GND.t396 17.475
R3046 GND.n3938 GND.t575 17.4601
R3047 GND.n5240 GND.t835 17.4601
R3048 GND.n3553 GND.t531 17.4601
R3049 GND.n1146 GND.t106 17.4601
R3050 GND.n5616 GND.t806 17.4601
R3051 GND.n1289 GND.t432 17.4601
R3052 GND.n2924 GND.t130 17.4601
R3053 GND.n2487 GND.t832 17.4601
R3054 GND.n2007 GND.t123 17.4601
R3055 GND.n1588 GND.t804 17.4601
R3056 GND.n2378 GND.t529 17.4601
R3057 GND.n2699 GND.t430 17.4601
R3058 GND.n144 GND.t573 17.4601
R3059 GND.n4965 GND.t511 17.4601
R3060 GND.n3723 GND.t523 17.4601
R3061 GND.n3779 GND.t830 17.4601
R3062 GND.n5565 GND.t1229 17.4528
R3063 GND.n6550 GND.t788 17.4528
R3064 GND.n7561 GND.t1227 17.4528
R3065 GND.n5110 GND.t584 17.4528
R3066 GND.n3331 GND.t1234 17.4528
R3067 GND.n3464 GND.t824 17.4528
R3068 GND.n6803 GND.t1248 17.4528
R3069 GND.n7127 GND.t1515 17.4528
R3070 GND.n1876 GND.t1083 17.4528
R3071 GND.n2202 GND.t420 17.4528
R3072 GND.n6957 GND.t580 17.4528
R3073 GND.n6657 GND.t232 17.4528
R3074 GND.n4789 GND.t731 17.4528
R3075 GND.n7499 GND.t1246 17.4528
R3076 GND.n7624 GND.t582 17.4528
R3077 GND.n1459 GND.t735 17.4528
R3078 GND.n192 GND.n191 17.2882
R3079 GND.n5999 GND.t994 17.2168
R3080 GND.t19 GND 17.1372
R3081 GND.t435 GND 17.1372
R3082 GND.t498 GND 17.1372
R3083 GND.n592 GND.n591 16.9417
R3084 GND.n7408 GND.n7407 16.9417
R3085 GND.n7361 GND.n7360 16.9417
R3086 GND.n7302 GND.n7301 16.9417
R3087 GND.n7276 GND.n7275 16.9417
R3088 GND.n5802 GND.n5801 16.9417
R3089 GND.n5690 GND.n5689 16.9417
R3090 GND.n5744 GND.n5743 16.9417
R3091 GND.n6175 GND.n6174 16.9417
R3092 GND.n5679 GND.n5678 16.9417
R3093 GND.n945 GND.n944 16.9417
R3094 GND.n911 GND.n910 16.9417
R3095 GND.n846 GND.n845 16.9417
R3096 GND.n818 GND.n817 16.9417
R3097 GND.n748 GND.n747 16.9417
R3098 GND.n707 GND.n703 16.9417
R3099 GND.n709 GND.n683 16.9417
R3100 GND.n6258 GND.n6254 16.9417
R3101 GND.n6260 GND.n6234 16.9417
R3102 GND.n6058 GND.n6057 16.9417
R3103 GND.n6010 GND.n6009 16.9417
R3104 GND.n5988 GND.n5987 16.9417
R3105 GND.n5929 GND.n5928 16.9417
R3106 GND.n5903 GND.n5902 16.9417
R3107 GND.t27 GND 16.9356
R3108 GND.t553 GND.t860 16.8628
R3109 GND GND.t553 16.2041
R3110 GND.n1525 GND.n1524 16.1887
R3111 GND.n5635 GND.n1005 16.1887
R3112 GND.n6501 GND.n6500 16.1887
R3113 GND.n7512 GND.n7511 16.1887
R3114 GND.n5212 GND.n5211 16.1887
R3115 GND.n3477 GND.n3476 16.1887
R3116 GND.n5453 GND.n1113 16.1887
R3117 GND.n6818 GND.n6767 16.1887
R3118 GND.n7078 GND.n7077 16.1887
R3119 GND.n1979 GND.n1978 16.1887
R3120 GND.n2302 GND.n2301 16.1887
R3121 GND.n6972 GND.n6921 16.1887
R3122 GND.n7748 GND.n51 16.1887
R3123 GND.n4888 GND.n4887 16.1887
R3124 GND.n7450 GND.n7449 16.1887
R3125 GND.n7575 GND.n7574 16.1887
R3126 GND.n694 GND.n693 16.1887
R3127 GND.n6245 GND.n6244 16.1887
R3128 GND.n1385 GND.n1383 14.7755
R3129 GND.n2134 GND.n2132 14.7755
R3130 GND.n2144 GND.n2139 14.7755
R3131 GND.n2136 GND.n2131 14.7755
R3132 GND.n2142 GND.n2140 14.7755
R3133 GND.n2614 GND.n2612 14.7755
R3134 GND.n2777 GND.n2776 14.7755
R3135 GND.n2616 GND.n2611 14.7755
R3136 GND.n2779 GND.n2775 14.7755
R3137 GND.n2787 GND.n2782 14.7755
R3138 GND.n2785 GND.n2783 14.7755
R3139 GND.n120 GND.n119 14.7755
R3140 GND.n117 GND.n115 14.7755
R3141 GND.n7710 GND.n7708 14.7755
R3142 GND.n3035 GND.n3030 14.7755
R3143 GND.n3027 GND.n3026 14.7755
R3144 GND.n3033 GND.n3031 14.7755
R3145 GND.n1232 GND.n1230 14.7755
R3146 GND.n1242 GND.n1237 14.7755
R3147 GND.n1234 GND.n1229 14.7755
R3148 GND.n1240 GND.n1238 14.7755
R3149 GND.n5367 GND.n5365 14.7755
R3150 GND.n5377 GND.n5372 14.7755
R3151 GND.n5369 GND.n5364 14.7755
R3152 GND.n5375 GND.n5373 14.7755
R3153 GND.n5046 GND.n5041 14.7755
R3154 GND.n5044 GND.n5042 14.7755
R3155 GND.n3652 GND.n3651 14.7755
R3156 GND.n3649 GND.n3648 14.7755
R3157 GND.n4042 GND.n4040 14.7755
R3158 GND.n3855 GND.n3854 14.7755
R3159 GND.n3844 GND.n3839 14.7755
R3160 GND.t228 GND.t1433 14.6672
R3161 GND.t35 GND.t797 14.6672
R3162 GND.t867 GND.t859 14.6672
R3163 GND.t627 GND.t927 14.6672
R3164 GND.t402 GND.t1091 14.6672
R3165 GND.t669 GND.t662 14.6672
R3166 GND.n7797 GND.n3 14.5711
R3167 GND.n1002 GND.n978 14.5711
R3168 GND.n6115 GND.n6091 14.5711
R3169 GND.t124 GND.n3810 14.4569
R3170 GND.n834 GND.t390 14.2308
R3171 GND.t15 GND.t570 14.228
R3172 GND.n7374 GND.t1183 13.8225
R3173 GND.n6482 GND.n6479 13.5727
R3174 GND.n6392 GND.n6389 13.5727
R3175 GND.n6482 GND.n6481 13.5705
R3176 GND.n6392 GND.n6391 13.5705
R3177 GND.n670 GND.n669 13.5646
R3178 GND.n6285 GND.n6284 13.5646
R3179 GND.n4408 GND.n4407 13.4405
R3180 GND.n5693 GND.t1378 13.4015
R3181 GND.n7786 GND.n7751 13.3549
R3182 GND.t858 GND 13.3059
R3183 GND.t1483 GND.t918 12.9107
R3184 GND.t629 GND.t691 12.6472
R3185 GND.n1585 GND.t803 12.5719
R3186 GND GND.t721 12.5248
R3187 GND GND.t255 12.5248
R3188 GND GND.t694 12.5248
R3189 GND GND.t900 12.5248
R3190 GND GND.t146 12.5248
R3191 GND GND.t516 12.5248
R3192 GND.t1393 GND 12.5248
R3193 GND.t685 GND 12.5248
R3194 GND GND.t2 12.5248
R3195 GND.t186 GND.n1742 11.89
R3196 GND.n5419 GND.t186 11.89
R3197 GND.t501 GND.n4221 11.89
R3198 GND.t1566 GND.n4583 11.89
R3199 GND.t217 GND.n4567 11.89
R3200 GND.t1495 GND.n4552 11.89
R3201 GND.t1563 GND.n4537 11.89
R3202 GND.t1500 GND.n4522 11.89
R3203 GND.t1564 GND.n4505 11.89
R3204 GND.t216 GND.n4490 11.89
R3205 GND.t1494 GND.n4475 11.89
R3206 GND.t1562 GND.n4460 11.89
R3207 GND.t1496 GND.n4443 11.89
R3208 GND.t827 GND.n4423 11.89
R3209 GND.t218 GND.n4381 11.89
R3210 GND.t1499 GND.n4366 11.89
R3211 GND.t213 GND.n4351 11.89
R3212 GND.t1498 GND.n4336 11.89
R3213 GND.t1561 GND.n4317 11.89
R3214 GND.t215 GND.n4302 11.89
R3215 GND.t1565 GND.n4287 11.89
R3216 GND.t1501 GND.n4272 11.89
R3217 GND.n596 GND.n595 11.6711
R3218 GND.n7412 GND.n7411 11.6711
R3219 GND.n7365 GND.n7364 11.6711
R3220 GND.n7298 GND.n7297 11.6711
R3221 GND.n7281 GND.n7280 11.6711
R3222 GND.n5806 GND.n5805 11.6711
R3223 GND.n5759 GND.n5758 11.6711
R3224 GND.n5749 GND.n5748 11.6711
R3225 GND.n6171 GND.n6170 11.6711
R3226 GND.n5675 GND.n5674 11.6711
R3227 GND.n941 GND.n940 11.6711
R3228 GND.n915 GND.n914 11.6711
R3229 GND.n842 GND.n841 11.6711
R3230 GND.n822 GND.n821 11.6711
R3231 GND.n743 GND.n742 11.6711
R3232 GND.n6054 GND.n6053 11.6711
R3233 GND.n6006 GND.n6005 11.6711
R3234 GND.n5992 GND.n5991 11.6711
R3235 GND.n5925 GND.n5924 11.6711
R3236 GND.n5908 GND.n5907 11.6711
R3237 GND.t214 GND.n4396 11.48
R3238 GND.n6203 GND.n6202 11.427
R3239 GND.n6201 GND.n6200 11.427
R3240 GND.n6425 GND.n6424 11.427
R3241 GND.n522 GND.n521 11.427
R3242 GND.t918 GND.t397 11.0664
R3243 GND.t397 GND.t629 11.0664
R3244 GND.t570 GND.t858 11.0664
R3245 GND.t710 GND 10.9511
R3246 GND.t1438 GND 10.9511
R3247 GND.t938 GND 10.9511
R3248 GND GND.t137 10.9511
R3249 GND GND.t95 10.9511
R3250 GND GND.t843 10.9511
R3251 GND GND.t1425 10.9511
R3252 GND.n586 GND.n585 10.9181
R3253 GND.n7402 GND.n7401 10.9181
R3254 GND.n7355 GND.n7354 10.9181
R3255 GND.n7308 GND.n7307 10.9181
R3256 GND.n7270 GND.n7269 10.9181
R3257 GND.n5796 GND.n5795 10.9181
R3258 GND.n5699 GND.n5698 10.9181
R3259 GND.n5737 GND.n5736 10.9181
R3260 GND.n6181 GND.n6180 10.9181
R3261 GND.n5845 GND.n5844 10.9181
R3262 GND.n951 GND.n950 10.9181
R3263 GND.n905 GND.n904 10.9181
R3264 GND.n852 GND.n851 10.9181
R3265 GND.n812 GND.n811 10.9181
R3266 GND.n754 GND.n753 10.9181
R3267 GND.n6064 GND.n6063 10.9181
R3268 GND.n6016 GND.n6015 10.9181
R3269 GND.n5982 GND.n5981 10.9181
R3270 GND.n5935 GND.n5934 10.9181
R3271 GND.n5897 GND.n5896 10.9181
R3272 GND GND.t663 10.6857
R3273 GND GND.t19 10.6857
R3274 GND GND.t435 10.6857
R3275 GND GND.t27 10.6857
R3276 GND GND.t498 10.6857
R3277 GND.n6204 GND.n6203 10.5417
R3278 GND.t799 GND.n4737 10.3672
R3279 GND GND.n7229 10.1442
R3280 GND.n2019 GND.n2016 9.8307
R3281 GND.t500 GND.t822 9.8307
R3282 GND.n2034 GND.n2031 9.8307
R3283 GND.n2338 GND.n2335 9.8307
R3284 GND.t1089 GND.t826 9.8307
R3285 GND.n2371 GND.n2368 9.8307
R3286 GND.n2499 GND.n2496 9.8307
R3287 GND.t1415 GND.t58 9.8307
R3288 GND.n2514 GND.n2511 9.8307
R3289 GND.n2659 GND.n2656 9.8307
R3290 GND.t1239 GND.t1096 9.8307
R3291 GND.n2692 GND.n2689 9.8307
R3292 GND.n2915 GND.n2912 9.8307
R3293 GND.t1230 GND.t576 9.8307
R3294 GND.n2932 GND.n2929 9.8307
R3295 GND.n96 GND.n93 9.8307
R3296 GND.t249 GND.t484 9.8307
R3297 GND.n137 GND.n134 9.8307
R3298 GND.n1301 GND.n1298 9.8307
R3299 GND.t1399 GND.t578 9.8307
R3300 GND.n1316 GND.n1313 9.8307
R3301 GND.n5576 GND.n5573 9.8307
R3302 GND.t108 GND.t1243 9.8307
R3303 GND.n5591 GND.n5588 9.8307
R3304 GND.n1137 GND.n1134 9.8307
R3305 GND.t947 GND.t1513 9.8307
R3306 GND.n1154 GND.n1151 9.8307
R3307 GND.n3513 GND.n3510 9.8307
R3308 GND.t657 GND.t246 9.8307
R3309 GND.n3528 GND.n3525 9.8307
R3310 GND.n5252 GND.n5249 9.8307
R3311 GND.t1419 GND.t47 9.8307
R3312 GND.n5267 GND.n5264 9.8307
R3313 GND.n4925 GND.n4922 9.8307
R3314 GND.t427 GND.t199 9.8307
R3315 GND.n4958 GND.n4955 9.8307
R3316 GND.n3683 GND.n3680 9.8307
R3317 GND.t1241 GND.t809 9.8307
R3318 GND.n3716 GND.n3713 9.8307
R3319 GND.n3950 GND.n3947 9.8307
R3320 GND.t874 GND.t796 9.8307
R3321 GND.n3965 GND.n3962 9.8307
R3322 GND.n3739 GND.n3736 9.8307
R3323 GND.t1225 GND.t23 9.8307
R3324 GND.n3772 GND.n3769 9.8307
R3325 GND.t860 GND.t535 9.48553
R3326 GND.t535 GND.t1081 9.48553
R3327 GND.n40 GND.n38 9.41227
R3328 GND.n6364 GND.n6362 9.41227
R3329 GND.n666 GND.n665 9.41227
R3330 GND.n6281 GND.n6280 9.41227
R3331 GND.n1452 GND.n1451 9.3005
R3332 GND.n1438 GND.n1437 9.3005
R3333 GND.n1440 GND.n1439 9.3005
R3334 GND.n1542 GND.n1541 9.3005
R3335 GND.n1526 GND.n1525 9.3005
R3336 GND.n1035 GND.n1034 9.3005
R3337 GND.n1022 GND.n1021 9.3005
R3338 GND.n1024 GND.n1023 9.3005
R3339 GND.n1037 GND.n1036 9.3005
R3340 GND.n1014 GND.n1013 9.3005
R3341 GND.n5636 GND.n5635 9.3005
R3342 GND.n1042 GND.n1041 9.3005
R3343 GND.n5492 GND.n5491 9.3005
R3344 GND.n1053 GND.n1052 9.3005
R3345 GND.n1044 GND.n1043 9.3005
R3346 GND.n1056 GND.n1055 9.3005
R3347 GND.n1109 GND.n1108 9.3005
R3348 GND.n5462 GND.n5461 9.3005
R3349 GND.n1111 GND.n1110 9.3005
R3350 GND.n6543 GND.n6542 9.3005
R3351 GND.n6530 GND.n6529 9.3005
R3352 GND.n6532 GND.n6531 9.3005
R3353 GND.n6545 GND.n6544 9.3005
R3354 GND.n6514 GND.n6513 9.3005
R3355 GND.n6502 GND.n6501 9.3005
R3356 GND.n5469 GND.n5468 9.3005
R3357 GND.n6595 GND.n6594 9.3005
R3358 GND.n5480 GND.n5479 9.3005
R3359 GND.n5471 GND.n5470 9.3005
R3360 GND.n5483 GND.n5482 9.3005
R3361 GND.n5543 GND.n5542 9.3005
R3362 GND.n5641 GND.n5640 9.3005
R3363 GND.n5545 GND.n5544 9.3005
R3364 GND.n7554 GND.n7553 9.3005
R3365 GND.n7541 GND.n7540 9.3005
R3366 GND.n7543 GND.n7542 9.3005
R3367 GND.n7556 GND.n7555 9.3005
R3368 GND.n7525 GND.n7524 9.3005
R3369 GND.n7513 GND.n7512 9.3005
R3370 GND.n225 GND.n224 9.3005
R3371 GND.n359 GND.n358 9.3005
R3372 GND.n236 GND.n235 9.3005
R3373 GND.n227 GND.n226 9.3005
R3374 GND.n239 GND.n238 9.3005
R3375 GND.n299 GND.n298 9.3005
R3376 GND.n7566 GND.n7565 9.3005
R3377 GND.n301 GND.n300 9.3005
R3378 GND.n5092 GND.n5091 9.3005
R3379 GND.n5078 GND.n5077 9.3005
R3380 GND.n5080 GND.n5079 9.3005
R3381 GND.n5225 GND.n5224 9.3005
R3382 GND.n5213 GND.n5212 9.3005
R3383 GND.n4855 GND.n4854 9.3005
R3384 GND.n4852 GND.n4851 9.3005
R3385 GND.n4866 GND.n4865 9.3005
R3386 GND.n4857 GND.n4856 9.3005
R3387 GND.n4869 GND.n4868 9.3005
R3388 GND.n5100 GND.n5099 9.3005
R3389 GND.n5107 GND.n5106 9.3005
R3390 GND.n5102 GND.n5101 9.3005
R3391 GND.n3303 GND.n3302 9.3005
R3392 GND.n3289 GND.n3288 9.3005
R3393 GND.n3291 GND.n3290 9.3005
R3394 GND.n3490 GND.n3489 9.3005
R3395 GND.n3478 GND.n3477 9.3005
R3396 GND.n5179 GND.n5178 9.3005
R3397 GND.n5176 GND.n5175 9.3005
R3398 GND.n5190 GND.n5189 9.3005
R3399 GND.n5181 GND.n5180 9.3005
R3400 GND.n5193 GND.n5192 9.3005
R3401 GND.n3309 GND.n3308 9.3005
R3402 GND.n3316 GND.n3315 9.3005
R3403 GND.n3311 GND.n3310 9.3005
R3404 GND.n3457 GND.n3456 9.3005
R3405 GND.n3444 GND.n3443 9.3005
R3406 GND.n3446 GND.n3445 9.3005
R3407 GND.n3459 GND.n3458 9.3005
R3408 GND.n1122 GND.n1121 9.3005
R3409 GND.n5454 GND.n5453 9.3005
R3410 GND.n3352 GND.n3351 9.3005
R3411 GND.n1058 GND.n1057 9.3005
R3412 GND.n3363 GND.n3362 9.3005
R3413 GND.n3354 GND.n3353 9.3005
R3414 GND.n3366 GND.n3365 9.3005
R3415 GND.n3417 GND.n3416 9.3005
R3416 GND.n3469 GND.n3468 9.3005
R3417 GND.n3419 GND.n3418 9.3005
R3418 GND.n6797 GND.n6796 9.3005
R3419 GND.n6784 GND.n6783 9.3005
R3420 GND.n6786 GND.n6785 9.3005
R3421 GND.n6799 GND.n6798 9.3005
R3422 GND.n6776 GND.n6775 9.3005
R3423 GND.n6819 GND.n6818 9.3005
R3424 GND.n6730 GND.n6729 9.3005
R3425 GND.n6727 GND.n6726 9.3005
R3426 GND.n6741 GND.n6740 9.3005
R3427 GND.n6732 GND.n6731 9.3005
R3428 GND.n6744 GND.n6743 9.3005
R3429 GND.n6709 GND.n6708 9.3005
R3430 GND.n630 GND.n629 9.3005
R3431 GND.n6762 GND.n6761 9.3005
R3432 GND.n7120 GND.n7119 9.3005
R3433 GND.n7107 GND.n7106 9.3005
R3434 GND.n7109 GND.n7108 9.3005
R3435 GND.n7122 GND.n7121 9.3005
R3436 GND.n7091 GND.n7090 9.3005
R3437 GND.n7079 GND.n7078 9.3005
R3438 GND.n7038 GND.n7037 9.3005
R3439 GND.n7035 GND.n7034 9.3005
R3440 GND.n7049 GND.n7048 9.3005
R3441 GND.n7040 GND.n7039 9.3005
R3442 GND.n7052 GND.n7051 9.3005
R3443 GND.n7017 GND.n7016 9.3005
R3444 GND.n610 GND.n609 9.3005
R3445 GND.n7070 GND.n7069 9.3005
R3446 GND.n1857 GND.n1856 9.3005
R3447 GND.n1844 GND.n1843 9.3005
R3448 GND.n1846 GND.n1845 9.3005
R3449 GND.n1859 GND.n1858 9.3005
R3450 GND.n1992 GND.n1991 9.3005
R3451 GND.n1980 GND.n1979 9.3005
R3452 GND.n2269 GND.n2268 9.3005
R3453 GND.n2266 GND.n2265 9.3005
R3454 GND.n2280 GND.n2279 9.3005
R3455 GND.n2271 GND.n2270 9.3005
R3456 GND.n2283 GND.n2282 9.3005
R3457 GND.n1866 GND.n1865 9.3005
R3458 GND.n1873 GND.n1872 9.3005
R3459 GND.n1868 GND.n1867 9.3005
R3460 GND.n1430 GND.n1429 9.3005
R3461 GND.n2161 GND.n2160 9.3005
R3462 GND.n2160 GND.n2159 9.3005
R3463 GND.n2189 GND.n2188 9.3005
R3464 GND.n2179 GND.n2178 9.3005
R3465 GND.n2181 GND.n2180 9.3005
R3466 GND.n2191 GND.n2190 9.3005
R3467 GND.n2315 GND.n2314 9.3005
R3468 GND.n2303 GND.n2302 9.3005
R3469 GND.n7199 GND.n7198 9.3005
R3470 GND.n7196 GND.n7195 9.3005
R3471 GND.n7210 GND.n7209 9.3005
R3472 GND.n7201 GND.n7200 9.3005
R3473 GND.n7213 GND.n7212 9.3005
R3474 GND.n7183 GND.n7182 9.3005
R3475 GND.n7131 GND.n7130 9.3005
R3476 GND.n7133 GND.n7132 9.3005
R3477 GND.n2470 GND.n2469 9.3005
R3478 GND.n2635 GND.n2634 9.3005
R3479 GND.n2634 GND.n2633 9.3005
R3480 GND.n6951 GND.n6950 9.3005
R3481 GND.n6938 GND.n6937 9.3005
R3482 GND.n6940 GND.n6939 9.3005
R3483 GND.n6953 GND.n6952 9.3005
R3484 GND.n6930 GND.n6929 9.3005
R3485 GND.n6973 GND.n6972 9.3005
R3486 GND.n6884 GND.n6883 9.3005
R3487 GND.n6881 GND.n6880 9.3005
R3488 GND.n6895 GND.n6894 9.3005
R3489 GND.n6886 GND.n6885 9.3005
R3490 GND.n6898 GND.n6897 9.3005
R3491 GND.n6863 GND.n6862 9.3005
R3492 GND.n620 GND.n619 9.3005
R3493 GND.n6916 GND.n6915 9.3005
R3494 GND.n2804 GND.n2803 9.3005
R3495 GND.n2900 GND.n2899 9.3005
R3496 GND.n2899 GND.n2898 9.3005
R3497 GND.n81 GND.n80 9.3005
R3498 GND.n68 GND.n67 9.3005
R3499 GND.n70 GND.n69 9.3005
R3500 GND.n83 GND.n82 9.3005
R3501 GND.n59 GND.n58 9.3005
R3502 GND.n7749 GND.n7748 9.3005
R3503 GND.n6572 GND.n6571 9.3005
R3504 GND.n6569 GND.n6568 9.3005
R3505 GND.n6583 GND.n6582 9.3005
R3506 GND.n6574 GND.n6573 9.3005
R3507 GND.n6586 GND.n6585 9.3005
R3508 GND.n6646 GND.n6645 9.3005
R3509 GND.n6654 GND.n6653 9.3005
R3510 GND.n6648 GND.n6647 9.3005
R3511 GND.n7727 GND.n7726 9.3005
R3512 GND.n3052 GND.n3051 9.3005
R3513 GND.n3051 GND.n3050 9.3005
R3514 GND.n3152 GND.n3151 9.3005
R3515 GND.n1259 GND.n1258 9.3005
R3516 GND.n1258 GND.n1257 9.3005
R3517 GND.n3259 GND.n3258 9.3005
R3518 GND.n5394 GND.n5393 9.3005
R3519 GND.n5393 GND.n5392 9.3005
R3520 GND.n4770 GND.n4769 9.3005
R3521 GND.n4757 GND.n4756 9.3005
R3522 GND.n4759 GND.n4758 9.3005
R3523 GND.n4772 GND.n4771 9.3005
R3524 GND.n4901 GND.n4900 9.3005
R3525 GND.n4889 GND.n4888 9.3005
R3526 GND.n484 GND.n483 9.3005
R3527 GND.n481 GND.n480 9.3005
R3528 GND.n495 GND.n494 9.3005
R3529 GND.n486 GND.n485 9.3005
R3530 GND.n498 GND.n497 9.3005
R3531 GND.n4779 GND.n4778 9.3005
R3532 GND.n4786 GND.n4785 9.3005
R3533 GND.n4781 GND.n4780 9.3005
R3534 GND.n5063 GND.n5062 9.3005
R3535 GND.n7492 GND.n7491 9.3005
R3536 GND.n7479 GND.n7478 9.3005
R3537 GND.n7481 GND.n7480 9.3005
R3538 GND.n7494 GND.n7493 9.3005
R3539 GND.n7463 GND.n7462 9.3005
R3540 GND.n7451 GND.n7450 9.3005
R3541 GND.n336 GND.n335 9.3005
R3542 GND.n333 GND.n332 9.3005
R3543 GND.n347 GND.n346 9.3005
R3544 GND.n338 GND.n337 9.3005
R3545 GND.n350 GND.n349 9.3005
R3546 GND.n410 GND.n409 9.3005
R3547 GND.n7504 GND.n7503 9.3005
R3548 GND.n412 GND.n411 9.3005
R3549 GND.n3669 GND.n3668 9.3005
R3550 GND.n4059 GND.n4058 9.3005
R3551 GND.n4058 GND.n4057 9.3005
R3552 GND.n7617 GND.n7616 9.3005
R3553 GND.n7604 GND.n7603 9.3005
R3554 GND.n7606 GND.n7605 9.3005
R3555 GND.n7619 GND.n7618 9.3005
R3556 GND.n7588 GND.n7587 9.3005
R3557 GND.n7576 GND.n7575 9.3005
R3558 GND.n7633 GND.n7632 9.3005
R3559 GND.n248 GND.n247 9.3005
R3560 GND.n7644 GND.n7643 9.3005
R3561 GND.n7635 GND.n7634 9.3005
R3562 GND.n7647 GND.n7646 9.3005
R3563 GND.n7631 GND.n7630 9.3005
R3564 GND.n200 GND.n199 9.3005
R3565 GND.n7629 GND.n7628 9.3005
R3566 GND.n4332 GND.n4331 9.3005
R3567 GND.n4244 GND.n4243 9.3005
R3568 GND.n4752 GND.n4751 9.3005
R3569 GND.n4519 GND.n4518 9.3005
R3570 GND.n3872 GND.n3871 9.3005
R3571 GND.n3871 GND.n3870 9.3005
R3572 GND.n1468 GND.n1467 9.3005
R3573 GND.n1463 GND.n1462 9.3005
R3574 GND.n1960 GND.n1959 9.3005
R3575 GND.n1461 GND.n1460 9.3005
R3576 GND.n1957 GND.n1956 9.3005
R3577 GND.n1948 GND.n1947 9.3005
R3578 GND.n1946 GND.n1945 9.3005
R3579 GND.n1937 GND.n1936 9.3005
R3580 GND.n1476 GND.n1475 9.3005
R3581 GND.n1518 GND.n1517 9.3005
R3582 GND.n1508 GND.n1507 9.3005
R3583 GND.n1487 GND.n1486 9.3005
R3584 GND.n1496 GND.n1495 9.3005
R3585 GND.n1478 GND.n1477 9.3005
R3586 GND.n1485 GND.n1484 9.3005
R3587 GND.n1893 GND.n1892 9.3005
R3588 GND.n1971 GND.n1970 9.3005
R3589 GND.n1930 GND.n1929 9.3005
R3590 GND.n1904 GND.n1903 9.3005
R3591 GND.n1913 GND.n1912 9.3005
R3592 GND.n1895 GND.n1894 9.3005
R3593 GND.n1902 GND.n1901 9.3005
R3594 GND.n2218 GND.n2217 9.3005
R3595 GND.n2294 GND.n2293 9.3005
R3596 GND.n2253 GND.n2252 9.3005
R3597 GND.n2227 GND.n2226 9.3005
R3598 GND.n2236 GND.n2235 9.3005
R3599 GND.n7191 GND.n7190 9.3005
R3600 GND.n2225 GND.n2224 9.3005
R3601 GND.n7149 GND.n7148 9.3005
R3602 GND.n7224 GND.n7223 9.3005
R3603 GND.n7179 GND.n7178 9.3005
R3604 GND.n7153 GND.n7152 9.3005
R3605 GND.n7162 GND.n7161 9.3005
R3606 GND.n7030 GND.n7029 9.3005
R3607 GND.n7151 GND.n7150 9.3005
R3608 GND.n7062 GND.n7061 9.3005
R3609 GND.n6982 GND.n6981 9.3005
R3610 GND.n7013 GND.n7012 9.3005
R3611 GND.n6987 GND.n6986 9.3005
R3612 GND.n6996 GND.n6995 9.3005
R3613 GND.n6876 GND.n6875 9.3005
R3614 GND.n6985 GND.n6984 9.3005
R3615 GND.n6908 GND.n6907 9.3005
R3616 GND.n6828 GND.n6827 9.3005
R3617 GND.n6859 GND.n6858 9.3005
R3618 GND.n6833 GND.n6832 9.3005
R3619 GND.n6842 GND.n6841 9.3005
R3620 GND.n6722 GND.n6721 9.3005
R3621 GND.n6831 GND.n6830 9.3005
R3622 GND.n6754 GND.n6753 9.3005
R3623 GND.n6664 GND.n6663 9.3005
R3624 GND.n6705 GND.n6704 9.3005
R3625 GND.n6679 GND.n6678 9.3005
R3626 GND.n6688 GND.n6687 9.3005
R3627 GND.n6670 GND.n6669 9.3005
R3628 GND.n6677 GND.n6676 9.3005
R3629 GND.n6555 GND.n6554 9.3005
R3630 GND.n648 GND.n647 9.3005
R3631 GND.n6635 GND.n6634 9.3005
R3632 GND.n6609 GND.n6608 9.3005
R3633 GND.n6618 GND.n6617 9.3005
R3634 GND.n6600 GND.n6599 9.3005
R3635 GND.n6607 GND.n6606 9.3005
R3636 GND.n5561 GND.n5560 9.3005
R3637 GND.n5467 GND.n5466 9.3005
R3638 GND.n5532 GND.n5531 9.3005
R3639 GND.n5506 GND.n5505 9.3005
R3640 GND.n5515 GND.n5514 9.3005
R3641 GND.n5497 GND.n5496 9.3005
R3642 GND.n5504 GND.n5503 9.3005
R3643 GND.n3439 GND.n3438 9.3005
R3644 GND.n3424 GND.n3423 9.3005
R3645 GND.n1098 GND.n1097 9.3005
R3646 GND.n1072 GND.n1071 9.3005
R3647 GND.n1081 GND.n1080 9.3005
R3648 GND.n1063 GND.n1062 9.3005
R3649 GND.n1070 GND.n1069 9.3005
R3650 GND.n3327 GND.n3326 9.3005
R3651 GND.n3322 GND.n3321 9.3005
R3652 GND.n3406 GND.n3405 9.3005
R3653 GND.n3380 GND.n3379 9.3005
R3654 GND.n3389 GND.n3388 9.3005
R3655 GND.n3371 GND.n3370 9.3005
R3656 GND.n3378 GND.n3377 9.3005
R3657 GND.n5126 GND.n5125 9.3005
R3658 GND.n5204 GND.n5203 9.3005
R3659 GND.n5166 GND.n5165 9.3005
R3660 GND.n5140 GND.n5139 9.3005
R3661 GND.n5149 GND.n5148 9.3005
R3662 GND.n5131 GND.n5130 9.3005
R3663 GND.n5138 GND.n5137 9.3005
R3664 GND.n4805 GND.n4804 9.3005
R3665 GND.n4880 GND.n4879 9.3005
R3666 GND.n4842 GND.n4841 9.3005
R3667 GND.n4816 GND.n4815 9.3005
R3668 GND.n4825 GND.n4824 9.3005
R3669 GND.n4807 GND.n4806 9.3005
R3670 GND.n4814 GND.n4813 9.3005
R3671 GND.n428 GND.n427 9.3005
R3672 GND.n511 GND.n510 9.3005
R3673 GND.n468 GND.n467 9.3005
R3674 GND.n442 GND.n441 9.3005
R3675 GND.n451 GND.n450 9.3005
R3676 GND.n433 GND.n432 9.3005
R3677 GND.n440 GND.n439 9.3005
R3678 GND.n319 GND.n318 9.3005
R3679 GND.n316 GND.n315 9.3005
R3680 GND.n399 GND.n398 9.3005
R3681 GND.n373 GND.n372 9.3005
R3682 GND.n382 GND.n381 9.3005
R3683 GND.n364 GND.n363 9.3005
R3684 GND.n371 GND.n370 9.3005
R3685 GND.n217 GND.n216 9.3005
R3686 GND.n214 GND.n213 9.3005
R3687 GND.n288 GND.n287 9.3005
R3688 GND.n262 GND.n261 9.3005
R3689 GND.n271 GND.n270 9.3005
R3690 GND.n253 GND.n252 9.3005
R3691 GND.n260 GND.n259 9.3005
R3692 GND.n4607 GND.n4606 9.2805
R3693 GND.n1429 GND.n1427 9.1766
R3694 GND.n2469 GND.n2467 9.1766
R3695 GND.n2803 GND.n2801 9.1766
R3696 GND.n7726 GND.n7724 9.1766
R3697 GND.n3151 GND.n3149 9.1766
R3698 GND.n3258 GND.n3256 9.1766
R3699 GND.n5062 GND.n5060 9.1766
R3700 GND.n3668 GND.n3666 9.1766
R3701 GND.n2020 GND.n2019 8.84768
R3702 GND.n2339 GND.n2338 8.84768
R3703 GND.n2500 GND.n2499 8.84768
R3704 GND.n2660 GND.n2659 8.84768
R3705 GND.n2916 GND.n2915 8.84768
R3706 GND.n97 GND.n96 8.84768
R3707 GND.n1302 GND.n1301 8.84768
R3708 GND.n5577 GND.n5576 8.84768
R3709 GND.n1138 GND.n1137 8.84768
R3710 GND.n3514 GND.n3513 8.84768
R3711 GND.n5253 GND.n5252 8.84768
R3712 GND.n4926 GND.n4925 8.84768
R3713 GND.n3684 GND.n3683 8.84768
R3714 GND.n3951 GND.n3950 8.84768
R3715 GND.n3740 GND.n3739 8.84768
R3716 GND.n1469 GND.t915 8.70904
R3717 GND.n5463 GND.t624 8.70904
R3718 GND.n5639 GND.t1 8.70904
R3719 GND.n7564 GND.t720 8.70904
R3720 GND.n5108 GND.t1252 8.70904
R3721 GND.n3317 GND.t1489 8.70904
R3722 GND.n3467 GND.t537 8.70904
R3723 GND.n6764 GND.t1552 8.70904
R3724 GND.n7072 GND.t526 8.70904
R3725 GND.n1874 GND.t869 8.70904
R3726 GND.n2200 GND.t1493 8.70904
R3727 GND.n6918 GND.t632 8.70904
R3728 GND.n6655 GND.t227 8.70904
R3729 GND.n4787 GND.t1491 8.70904
R3730 GND.n7502 GND.t569 8.70904
R3731 GND.n201 GND.t626 8.70904
R3732 GND.n1474 GND.t821 8.70236
R3733 GND.n5559 GND.t254 8.70236
R3734 GND.n6556 GND.t651 8.70236
R3735 GND.n320 GND.t881 8.70236
R3736 GND.n5124 GND.t1509 8.70236
R3737 GND.n3325 GND.t904 8.70236
R3738 GND.n3437 GND.t1569 8.70236
R3739 GND.n6909 GND.t622 8.70236
R3740 GND.n7147 GND.t1404 8.70236
R3741 GND.n1891 GND.t1508 8.70236
R3742 GND.n2216 GND.t949 8.70236
R3743 GND.n7063 GND.t1490 8.70236
R3744 GND.n6755 GND.t937 8.70236
R3745 GND.n4803 GND.t424 8.70236
R3746 GND.n426 GND.t551 8.70236
R3747 GND.n218 GND.t1507 8.70236
R3748 GND.t1081 GND 8.56337
R3749 GND.t691 GND 8.43164
R3750 GND.t395 GND.t734 8.20945
R3751 GND.t67 GND.t1082 8.20945
R3752 GND.t922 GND.t419 8.20945
R3753 GND.t1435 GND.t1514 8.20945
R3754 GND.t1255 GND.t579 8.20945
R3755 GND.t31 GND.t1247 8.20945
R3756 GND.t37 GND.t231 8.20945
R3757 GND.t816 GND.t787 8.20945
R3758 GND.t416 GND.t1228 8.20945
R3759 GND.t739 GND.t823 8.20945
R3760 GND.t496 GND.t1233 8.20945
R3761 GND.t222 GND.t583 8.20945
R3762 GND.t29 GND.t730 8.20945
R3763 GND.t437 GND.t1245 8.20945
R3764 GND.t1485 GND.t1226 8.20945
R3765 GND.t1429 GND.t581 8.20945
R3766 GND.n2842 GND 8.05791
R3767 GND.n1352 GND 8.05791
R3768 GND.n2101 GND 8.05791
R3769 GND.n2424 GND 8.05791
R3770 GND.n2581 GND 8.05791
R3771 GND.n2745 GND 8.05791
R3772 GND.n7677 GND 8.05791
R3773 GND.n3018 GND 8.05791
R3774 GND.n3128 GND 8.05791
R3775 GND.n1185 GND 8.05791
R3776 GND.n3199 GND 8.05791
R3777 GND.n5334 GND 8.05791
R3778 GND.n5010 GND 8.05791
R3779 GND.n3615 GND 8.05791
R3780 GND.n4032 GND 8.05791
R3781 GND.n3831 GND 8.05791
R3782 GND.t916 GND.n4404 8.02446
R3783 GND.n4030 GND.n4029 7.90638
R3784 GND.n2862 GND.n2861 7.90638
R3785 GND.n1350 GND.n1349 7.90638
R3786 GND.n2099 GND.n2098 7.90638
R3787 GND.n2422 GND.n2421 7.90638
R3788 GND.n2579 GND.n2578 7.90638
R3789 GND.n2743 GND.n2742 7.90638
R3790 GND.n7675 GND.n7674 7.90638
R3791 GND.n3016 GND.n3015 7.90638
R3792 GND.n3126 GND.n3125 7.90638
R3793 GND.n1226 GND.n1225 7.90638
R3794 GND.n3240 GND.n3239 7.90638
R3795 GND.n5332 GND.n5331 7.90638
R3796 GND.n5008 GND.n5007 7.90638
R3797 GND.n3613 GND.n3612 7.90638
R3798 GND.n3829 GND.n3828 7.90638
R3799 GND.n7445 GND 7.56079
R3800 GND.n6118 GND.t966 7.37892
R3801 GND.n2056 GND.t122 6.88164
R3802 GND.n2363 GND.t528 6.88164
R3803 GND.n2536 GND.t831 6.88164
R3804 GND.n2684 GND.t429 6.88164
R3805 GND.n2954 GND.t129 6.88164
R3806 GND.n129 GND.t572 6.88164
R3807 GND.n1338 GND.t431 6.88164
R3808 GND.n5613 GND.t805 6.88164
R3809 GND.n1176 GND.t105 6.88164
R3810 GND.n3550 GND.t530 6.88164
R3811 GND.n5289 GND.t834 6.88164
R3812 GND.n4950 GND.t510 6.88164
R3813 GND.n3708 GND.t522 6.88164
R3814 GND.n3987 GND.t574 6.88164
R3815 GND.n3764 GND.t829 6.88164
R3816 GND.n7805 GND.n0 6.77697
R3817 GND.n994 GND.n981 6.77697
R3818 GND.n6448 GND.n6420 6.77697
R3819 GND.n6442 GND.n6421 6.77697
R3820 GND.n6436 GND.n6422 6.77697
R3821 GND.n6430 GND.n6423 6.77697
R3822 GND.n545 GND.n517 6.77697
R3823 GND.n539 GND.n518 6.77697
R3824 GND.n533 GND.n519 6.77697
R3825 GND.n527 GND.n520 6.77697
R3826 GND.n6107 GND.n6094 6.77697
R3827 GND.t1336 GND.n5692 6.70101
R3828 GND.n3039 GND.n3038 6.52989
R3829 GND.n1246 GND.n1245 6.52989
R3830 GND.n4046 GND.n4045 6.52989
R3831 GND.n1390 GND.n1389 6.5285
R3832 GND.n2148 GND.n2147 6.5285
R3833 GND.n2457 GND.n2456 6.5285
R3834 GND.n2622 GND.n2621 6.5285
R3835 GND.n2791 GND.n2790 6.5285
R3836 GND.n2878 GND.n2877 6.5285
R3837 GND.n7714 GND.n7713 6.5285
R3838 GND.n3139 GND.n3138 6.5285
R3839 GND.n3246 GND.n3245 6.5285
R3840 GND.n5381 GND.n5380 6.5285
R3841 GND.n5050 GND.n5049 6.5285
R3842 GND.n3656 GND.n3655 6.5285
R3843 GND.n3859 GND.n3858 6.5285
R3844 GND.n41 GND.n40 6.4005
R3845 GND.n6365 GND.n6364 6.4005
R3846 GND.n6484 GND.n6479 6.4005
R3847 GND.n6481 GND.n6476 6.4005
R3848 GND.n665 GND.n653 6.4005
R3849 GND.n671 GND.n670 6.4005
R3850 GND.n6394 GND.n6389 6.4005
R3851 GND.n6391 GND.n6386 6.4005
R3852 GND.n6280 GND.n6268 6.4005
R3853 GND.n6286 GND.n6285 6.4005
R3854 GND.n7817 GND.n7816 6.15638
R3855 GND.n983 GND.n982 6.15638
R3856 GND.n6096 GND.n6095 6.15638
R3857 GND.n7748 GND.n7747 6.02403
R3858 GND.n602 GND.n601 5.64756
R3859 GND.n7419 GND.n7418 5.64756
R3860 GND.n7339 GND.n7338 5.64756
R3861 GND.n7291 GND.n7290 5.64756
R3862 GND.n7239 GND.n7238 5.64756
R3863 GND.n1206 GND 5.64756
R3864 GND.n3219 GND 5.64756
R3865 GND.n4010 GND 5.64756
R3866 GND.n5312 GND 5.64756
R3867 GND.n2996 GND 5.64756
R3868 GND.n2559 GND 5.64756
R3869 GND.n2079 GND 5.64756
R3870 GND.n1412 GND 5.64756
R3871 GND.n2401 GND 5.64756
R3872 GND.n2722 GND 5.64756
R3873 GND.n2830 GND 5.64756
R3874 GND.n161 GND 5.64756
R3875 GND.n3105 GND 5.64756
R3876 GND.n4987 GND 5.64756
R3877 GND.n3593 GND 5.64756
R3878 GND.n3796 GND 5.64756
R3879 GND.n5812 GND.n5811 5.64756
R3880 GND.n5766 GND.n5765 5.64756
R3881 GND.n5729 GND.n5728 5.64756
R3882 GND.n6164 GND.n6163 5.64756
R3883 GND.n5669 GND.n5668 5.64756
R3884 GND.n935 GND.n934 5.64756
R3885 GND.n922 GND.n921 5.64756
R3886 GND.n723 GND.n722 5.64756
R3887 GND.n829 GND.n828 5.64756
R3888 GND.n732 GND.n731 5.64756
R3889 GND.n6048 GND.n6047 5.64756
R3890 GND.n5854 GND.n5853 5.64756
R3891 GND.n5966 GND.n5965 5.64756
R3892 GND.n5918 GND.n5917 5.64756
R3893 GND.n5866 GND.n5865 5.64756
R3894 GND.n1939 GND.n1938 5.62907
R3895 GND.n2257 GND.n2256 5.62907
R3896 GND.n7185 GND.n7184 5.62907
R3897 GND.n7019 GND.n7018 5.62907
R3898 GND.n6865 GND.n6864 5.62907
R3899 GND.n6711 GND.n6710 5.62907
R3900 GND.n6563 GND.n6562 5.62907
R3901 GND.n6588 GND.n6587 5.62907
R3902 GND.n5485 GND.n5484 5.62907
R3903 GND.n3345 GND.n3344 5.62907
R3904 GND.n5170 GND.n5169 5.62907
R3905 GND.n4846 GND.n4845 5.62907
R3906 GND.n472 GND.n471 5.62907
R3907 GND.n327 GND.n326 5.62907
R3908 GND.n352 GND.n351 5.62907
R3909 GND.n241 GND.n240 5.62907
R3910 GND.n3989 GND.n3958 5.1205
R3911 GND.n5291 GND.n5260 5.1205
R3912 GND.n3552 GND.n3521 5.1205
R3913 GND.n1178 GND.n1145 5.1205
R3914 GND.n5615 GND.n5584 5.1205
R3915 GND.n1340 GND.n1309 5.1205
R3916 GND.n2956 GND.n2923 5.1205
R3917 GND.n2538 GND.n2507 5.1205
R3918 GND.n2058 GND.n2027 5.1205
R3919 GND.n1587 GND.n1567 5.1205
R3920 GND.n2377 GND.n2346 5.1205
R3921 GND.n2698 GND.n2667 5.1205
R3922 GND.n143 GND.n104 5.1205
R3923 GND.n4964 GND.n4933 5.1205
R3924 GND.n3722 GND.n3691 5.1205
R3925 GND.n3778 GND.n3747 5.1205
R3926 GND.n4329 GND.n4328 4.90717
R3927 GND.n580 GND.n579 4.89462
R3928 GND.n7396 GND.n7395 4.89462
R3929 GND.n7349 GND.n7348 4.89462
R3930 GND.n7314 GND.n7313 4.89462
R3931 GND.n7264 GND.n7263 4.89462
R3932 GND.n1448 GND.n1447 4.89462
R3933 GND.n5088 GND.n5087 4.89462
R3934 GND.n3299 GND.n3298 4.89462
R3935 GND.n5788 GND.n5787 4.89462
R3936 GND.n5705 GND.n5704 4.89462
R3937 GND.n5652 GND.n5651 4.89462
R3938 GND.n6187 GND.n6186 4.89462
R3939 GND.n5839 GND.n5838 4.89462
R3940 GND.n957 GND.n956 4.89462
R3941 GND.n899 GND.n898 4.89462
R3942 GND.n858 GND.n857 4.89462
R3943 GND.n806 GND.n805 4.89462
R3944 GND.n760 GND.n759 4.89462
R3945 GND.n6070 GND.n6069 4.89462
R3946 GND.n6022 GND.n6021 4.89462
R3947 GND.n5976 GND.n5975 4.89462
R3948 GND.n5941 GND.n5940 4.89462
R3949 GND.n5891 GND.n5890 4.89462
R3950 GND.n4420 GND.t828 4.78444
R3951 GND.n1436 GND 4.66821
R3952 GND.n1020 GND 4.66821
R3953 GND.n6528 GND 4.66821
R3954 GND.n7539 GND 4.66821
R3955 GND.n5076 GND 4.66821
R3956 GND.n3287 GND 4.66821
R3957 GND.n3442 GND 4.66821
R3958 GND.n6782 GND 4.66821
R3959 GND.n7105 GND 4.66821
R3960 GND.n1842 GND 4.66821
R3961 GND.n2177 GND 4.66821
R3962 GND.n6936 GND 4.66821
R3963 GND.n66 GND 4.66821
R3964 GND.n4755 GND 4.66821
R3965 GND.n7477 GND 4.66821
R3966 GND.n7602 GND 4.66821
R3967 GND.n35 GND.n28 4.6505
R3968 GND.n46 GND.n25 4.6505
R3969 GND.n45 GND.n44 4.6505
R3970 GND.n43 GND.n26 4.6505
R3971 GND.n42 GND.n41 4.6505
R3972 GND.n38 GND.n27 4.6505
R3973 GND.n37 GND.n36 4.6505
R3974 GND.n34 GND.n33 4.6505
R3975 GND.n1450 GND.n1449 4.6505
R3976 GND.n1524 GND.n1523 4.6505
R3977 GND.n1540 GND.n1539 4.6505
R3978 GND.n1033 GND.n1032 4.6505
R3979 GND.n5637 GND.n1005 4.6505
R3980 GND.n1012 GND.n1011 4.6505
R3981 GND.n6541 GND.n6540 4.6505
R3982 GND.n6500 GND.n6499 4.6505
R3983 GND.n6512 GND.n6511 4.6505
R3984 GND.n7552 GND.n7551 4.6505
R3985 GND.n7511 GND.n7510 4.6505
R3986 GND.n7523 GND.n7522 4.6505
R3987 GND.n5090 GND.n5089 4.6505
R3988 GND.n5211 GND.n5210 4.6505
R3989 GND.n5223 GND.n5222 4.6505
R3990 GND.n3301 GND.n3300 4.6505
R3991 GND.n3476 GND.n3475 4.6505
R3992 GND.n3488 GND.n3487 4.6505
R3993 GND.n3455 GND.n3454 4.6505
R3994 GND.n5455 GND.n1113 4.6505
R3995 GND.n1120 GND.n1119 4.6505
R3996 GND.n6795 GND.n6794 4.6505
R3997 GND.n6820 GND.n6767 4.6505
R3998 GND.n6774 GND.n6773 4.6505
R3999 GND.n7118 GND.n7117 4.6505
R4000 GND.n7077 GND.n7076 4.6505
R4001 GND.n7089 GND.n7088 4.6505
R4002 GND.n1855 GND.n1854 4.6505
R4003 GND.n1978 GND.n1977 4.6505
R4004 GND.n1990 GND.n1989 4.6505
R4005 GND.n2187 GND.n2186 4.6505
R4006 GND.n2301 GND.n2300 4.6505
R4007 GND.n2313 GND.n2312 4.6505
R4008 GND.n6949 GND.n6948 4.6505
R4009 GND.n6974 GND.n6921 4.6505
R4010 GND.n6928 GND.n6927 4.6505
R4011 GND.n79 GND.n78 4.6505
R4012 GND.n7750 GND.n51 4.6505
R4013 GND.n57 GND.n56 4.6505
R4014 GND.n4768 GND.n4767 4.6505
R4015 GND.n4887 GND.n4886 4.6505
R4016 GND.n4899 GND.n4898 4.6505
R4017 GND.n7490 GND.n7489 4.6505
R4018 GND.n7449 GND.n7448 4.6505
R4019 GND.n7461 GND.n7460 4.6505
R4020 GND.n7615 GND.n7614 4.6505
R4021 GND.n7574 GND.n7573 4.6505
R4022 GND.n7586 GND.n7585 4.6505
R4023 GND.n6359 GND.n6352 4.6505
R4024 GND.n6370 GND.n6349 4.6505
R4025 GND.n6369 GND.n6368 4.6505
R4026 GND.n6367 GND.n6350 4.6505
R4027 GND.n6366 GND.n6365 4.6505
R4028 GND.n6362 GND.n6351 4.6505
R4029 GND.n6361 GND.n6360 4.6505
R4030 GND.n6358 GND.n6357 4.6505
R4031 GND.n6206 GND.n6199 4.6505
R4032 GND.n6218 GND.n6197 4.6505
R4033 GND.n6210 GND.n6198 4.6505
R4034 GND.n6217 GND.n6216 4.6505
R4035 GND.n6215 GND.n6214 4.6505
R4036 GND.n6212 GND.n6211 4.6505
R4037 GND.n6208 GND.n6207 4.6505
R4038 GND.n6205 GND.n6204 4.6505
R4039 GND.n6147 GND.n6146 4.6505
R4040 GND.n6149 GND.n6148 4.6505
R4041 GND.n6220 GND.n6196 4.6505
R4042 GND.n6151 GND.n6150 4.6505
R4043 GND.n6155 GND.n6154 4.6505
R4044 GND.n6158 GND.n6157 4.6505
R4045 GND.n6165 GND.n6164 4.6505
R4046 GND.n6168 GND.n6167 4.6505
R4047 GND.n6172 GND.n6171 4.6505
R4048 GND.n6176 GND.n6175 4.6505
R4049 GND.n6178 GND.n6177 4.6505
R4050 GND.n6182 GND.n6181 4.6505
R4051 GND.n6184 GND.n6183 4.6505
R4052 GND.n6188 GND.n6187 4.6505
R4053 GND.n6190 GND.n6189 4.6505
R4054 GND.n6195 GND.n6194 4.6505
R4055 GND.n6223 GND.n6222 4.6505
R4056 GND.n5740 GND.n5739 4.6505
R4057 GND.n5738 GND.n5737 4.6505
R4058 GND.n5734 GND.n5733 4.6505
R4059 GND.n5653 GND.n5652 4.6505
R4060 GND.n6138 GND.n6137 4.6505
R4061 GND.n6142 GND.n6141 4.6505
R4062 GND.n6144 GND.n6143 4.6505
R4063 GND.n5823 GND.n5822 4.6505
R4064 GND.n5777 GND.n5686 4.6505
R4065 GND.n5776 GND.n5687 4.6505
R4066 GND.n5716 GND.n5715 4.6505
R4067 GND.n5718 GND.n5717 4.6505
R4068 GND.n5821 GND.n5820 4.6505
R4069 GND.n5819 GND.n5818 4.6505
R4070 GND.n5815 GND.n5814 4.6505
R4071 GND.n5813 GND.n5812 4.6505
R4072 GND.n5809 GND.n5808 4.6505
R4073 GND.n5807 GND.n5806 4.6505
R4074 GND.n5803 GND.n5802 4.6505
R4075 GND.n5799 GND.n5798 4.6505
R4076 GND.n5797 GND.n5796 4.6505
R4077 GND.n5792 GND.n5791 4.6505
R4078 GND.n5789 GND.n5788 4.6505
R4079 GND.n5785 GND.n5784 4.6505
R4080 GND.n5783 GND.n5782 4.6505
R4081 GND.n5779 GND.n5778 4.6505
R4082 GND.n5775 GND.n5774 4.6505
R4083 GND.n5773 GND.n5772 4.6505
R4084 GND.n5769 GND.n5768 4.6505
R4085 GND.n5767 GND.n5766 4.6505
R4086 GND.n5763 GND.n5762 4.6505
R4087 GND.n5760 GND.n5759 4.6505
R4088 GND.n5691 GND.n5690 4.6505
R4089 GND.n5696 GND.n5695 4.6505
R4090 GND.n5700 GND.n5699 4.6505
R4091 GND.n5702 GND.n5701 4.6505
R4092 GND.n5706 GND.n5705 4.6505
R4093 GND.n5708 GND.n5707 4.6505
R4094 GND.n5712 GND.n5711 4.6505
R4095 GND.n5714 GND.n5713 4.6505
R4096 GND.n5720 GND.n5719 4.6505
R4097 GND.n5724 GND.n5723 4.6505
R4098 GND.n5726 GND.n5725 4.6505
R4099 GND.n5730 GND.n5729 4.6505
R4100 GND.n5732 GND.n5731 4.6505
R4101 GND.n5750 GND.n5749 4.6505
R4102 GND.n5745 GND.n5744 4.6505
R4103 GND.n5825 GND.n5824 4.6505
R4104 GND.n5828 GND.n5827 4.6505
R4105 GND.n5662 GND.n5661 4.6505
R4106 GND.n5665 GND.n5664 4.6505
R4107 GND.n5670 GND.n5669 4.6505
R4108 GND.n5672 GND.n5671 4.6505
R4109 GND.n5676 GND.n5675 4.6505
R4110 GND.n5680 GND.n5679 4.6505
R4111 GND.n5682 GND.n5681 4.6505
R4112 GND.n5846 GND.n5845 4.6505
R4113 GND.n5842 GND.n5841 4.6505
R4114 GND.n5840 GND.n5839 4.6505
R4115 GND.n5836 GND.n5835 4.6505
R4116 GND.n5834 GND.n5833 4.6505
R4117 GND.n771 GND.n770 4.6505
R4118 GND.n773 GND.n772 4.6505
R4119 GND.n795 GND.n783 4.6505
R4120 GND.n794 GND.n784 4.6505
R4121 GND.n870 GND.n869 4.6505
R4122 GND.n872 GND.n871 4.6505
R4123 GND.n888 GND.n882 4.6505
R4124 GND.n887 GND.n883 4.6505
R4125 GND.n968 GND.n967 4.6505
R4126 GND.n970 GND.n969 4.6505
R4127 GND.n980 GND.n979 4.6505
R4128 GND.n729 GND.n728 4.6505
R4129 GND.n733 GND.n732 4.6505
R4130 GND.n736 GND.n735 4.6505
R4131 GND.n744 GND.n743 4.6505
R4132 GND.n749 GND.n748 4.6505
R4133 GND.n751 GND.n750 4.6505
R4134 GND.n755 GND.n754 4.6505
R4135 GND.n757 GND.n756 4.6505
R4136 GND.n761 GND.n760 4.6505
R4137 GND.n763 GND.n762 4.6505
R4138 GND.n767 GND.n766 4.6505
R4139 GND.n769 GND.n768 4.6505
R4140 GND.n775 GND.n774 4.6505
R4141 GND.n779 GND.n778 4.6505
R4142 GND.n782 GND.n781 4.6505
R4143 GND.n830 GND.n829 4.6505
R4144 GND.n825 GND.n824 4.6505
R4145 GND.n823 GND.n822 4.6505
R4146 GND.n819 GND.n818 4.6505
R4147 GND.n815 GND.n814 4.6505
R4148 GND.n813 GND.n812 4.6505
R4149 GND.n809 GND.n808 4.6505
R4150 GND.n807 GND.n806 4.6505
R4151 GND.n803 GND.n802 4.6505
R4152 GND.n801 GND.n800 4.6505
R4153 GND.n797 GND.n796 4.6505
R4154 GND.n793 GND.n792 4.6505
R4155 GND.n791 GND.n790 4.6505
R4156 GND.n787 GND.n786 4.6505
R4157 GND.n724 GND.n723 4.6505
R4158 GND.n838 GND.n837 4.6505
R4159 GND.n843 GND.n842 4.6505
R4160 GND.n847 GND.n846 4.6505
R4161 GND.n849 GND.n848 4.6505
R4162 GND.n853 GND.n852 4.6505
R4163 GND.n855 GND.n854 4.6505
R4164 GND.n859 GND.n858 4.6505
R4165 GND.n861 GND.n860 4.6505
R4166 GND.n865 GND.n864 4.6505
R4167 GND.n868 GND.n867 4.6505
R4168 GND.n874 GND.n873 4.6505
R4169 GND.n878 GND.n877 4.6505
R4170 GND.n881 GND.n880 4.6505
R4171 GND.n923 GND.n922 4.6505
R4172 GND.n918 GND.n917 4.6505
R4173 GND.n916 GND.n915 4.6505
R4174 GND.n912 GND.n911 4.6505
R4175 GND.n908 GND.n907 4.6505
R4176 GND.n906 GND.n905 4.6505
R4177 GND.n902 GND.n901 4.6505
R4178 GND.n900 GND.n899 4.6505
R4179 GND.n896 GND.n895 4.6505
R4180 GND.n894 GND.n893 4.6505
R4181 GND.n890 GND.n889 4.6505
R4182 GND.n886 GND.n885 4.6505
R4183 GND.n720 GND.n719 4.6505
R4184 GND.n931 GND.n930 4.6505
R4185 GND.n936 GND.n935 4.6505
R4186 GND.n938 GND.n937 4.6505
R4187 GND.n942 GND.n941 4.6505
R4188 GND.n946 GND.n945 4.6505
R4189 GND.n948 GND.n947 4.6505
R4190 GND.n952 GND.n951 4.6505
R4191 GND.n954 GND.n953 4.6505
R4192 GND.n958 GND.n957 4.6505
R4193 GND.n960 GND.n959 4.6505
R4194 GND.n964 GND.n963 4.6505
R4195 GND.n966 GND.n965 4.6505
R4196 GND.n972 GND.n971 4.6505
R4197 GND.n975 GND.n974 4.6505
R4198 GND.n977 GND.n976 4.6505
R4199 GND.n1000 GND.n999 4.6505
R4200 GND.n997 GND.n996 4.6505
R4201 GND.n995 GND.n994 4.6505
R4202 GND.n993 GND.n992 4.6505
R4203 GND.n991 GND.n990 4.6505
R4204 GND.n989 GND.n988 4.6505
R4205 GND.n985 GND.n984 4.6505
R4206 GND.n20 GND.n19 4.6505
R4207 GND.n18 GND.n8 4.6505
R4208 GND.n17 GND.n16 4.6505
R4209 GND.n16 GND.n15 4.6505
R4210 GND.n14 GND.n8 4.6505
R4211 GND.n20 GND.n7 4.6505
R4212 GND.n22 GND.n21 4.6505
R4213 GND.n7766 GND.n7761 4.6505
R4214 GND.n7768 GND.n7767 4.6505
R4215 GND.n7775 GND.n7774 4.6505
R4216 GND.n7776 GND.n7756 4.6505
R4217 GND.n7778 GND.n7777 4.6505
R4218 GND.n7771 GND.n7759 4.6505
R4219 GND.n7774 GND.n7773 4.6505
R4220 GND.n7772 GND.n7756 4.6505
R4221 GND.n7778 GND.n7755 4.6505
R4222 GND.n7780 GND.n7779 4.6505
R4223 GND.n6477 GND.n6476 4.6505
R4224 GND.n6488 GND.n6487 4.6505
R4225 GND.n6484 GND.n6483 4.6505
R4226 GND.n6486 GND.n6485 4.6505
R4227 GND.n672 GND.n671 4.6505
R4228 GND.n663 GND.n656 4.6505
R4229 GND.n662 GND.n661 4.6505
R4230 GND.n668 GND.n667 4.6505
R4231 GND.n666 GND.n654 4.6505
R4232 GND.n672 GND.n653 4.6505
R4233 GND.n674 GND.n673 4.6505
R4234 GND.n693 GND.n687 4.6505
R4235 GND.n696 GND.n686 4.6505
R4236 GND.n684 GND.n683 4.6505
R4237 GND.n710 GND.n681 4.6505
R4238 GND.n692 GND.n691 4.6505
R4239 GND.n695 GND.n694 4.6505
R4240 GND.n698 GND.n697 4.6505
R4241 GND.n700 GND.n699 4.6505
R4242 GND.n709 GND.n708 4.6505
R4243 GND.n711 GND.n678 4.6505
R4244 GND.n713 GND.n712 4.6505
R4245 GND.n706 GND.n681 4.6505
R4246 GND.n708 GND.n707 4.6505
R4247 GND.n704 GND.n678 4.6505
R4248 GND.n713 GND.n679 4.6505
R4249 GND.n6427 GND.n6426 4.6505
R4250 GND.n6429 GND.n6428 4.6505
R4251 GND.n6431 GND.n6430 4.6505
R4252 GND.n6433 GND.n6432 4.6505
R4253 GND.n6435 GND.n6434 4.6505
R4254 GND.n6437 GND.n6436 4.6505
R4255 GND.n6439 GND.n6438 4.6505
R4256 GND.n6441 GND.n6440 4.6505
R4257 GND.n6443 GND.n6442 4.6505
R4258 GND.n6445 GND.n6444 4.6505
R4259 GND.n6447 GND.n6446 4.6505
R4260 GND.n6449 GND.n6448 4.6505
R4261 GND.n6342 GND.n6341 4.6505
R4262 GND.n6340 GND.n6330 4.6505
R4263 GND.n6339 GND.n6338 4.6505
R4264 GND.n6338 GND.n6337 4.6505
R4265 GND.n6336 GND.n6330 4.6505
R4266 GND.n6342 GND.n6329 4.6505
R4267 GND.n6344 GND.n6343 4.6505
R4268 GND.n6306 GND.n6301 4.6505
R4269 GND.n6308 GND.n6307 4.6505
R4270 GND.n6315 GND.n6314 4.6505
R4271 GND.n6316 GND.n6296 4.6505
R4272 GND.n6318 GND.n6317 4.6505
R4273 GND.n6311 GND.n6299 4.6505
R4274 GND.n6314 GND.n6313 4.6505
R4275 GND.n6312 GND.n6296 4.6505
R4276 GND.n6318 GND.n6295 4.6505
R4277 GND.n6320 GND.n6319 4.6505
R4278 GND.n6387 GND.n6386 4.6505
R4279 GND.n6398 GND.n6397 4.6505
R4280 GND.n6394 GND.n6393 4.6505
R4281 GND.n6396 GND.n6395 4.6505
R4282 GND.n6287 GND.n6286 4.6505
R4283 GND.n6278 GND.n6271 4.6505
R4284 GND.n6277 GND.n6276 4.6505
R4285 GND.n6283 GND.n6282 4.6505
R4286 GND.n6281 GND.n6269 4.6505
R4287 GND.n6287 GND.n6268 4.6505
R4288 GND.n6289 GND.n6288 4.6505
R4289 GND.n6244 GND.n6238 4.6505
R4290 GND.n6247 GND.n6237 4.6505
R4291 GND.n6235 GND.n6234 4.6505
R4292 GND.n6261 GND.n6232 4.6505
R4293 GND.n6243 GND.n6242 4.6505
R4294 GND.n6246 GND.n6245 4.6505
R4295 GND.n6249 GND.n6248 4.6505
R4296 GND.n6251 GND.n6250 4.6505
R4297 GND.n6260 GND.n6259 4.6505
R4298 GND.n6262 GND.n6229 4.6505
R4299 GND.n6264 GND.n6263 4.6505
R4300 GND.n6257 GND.n6232 4.6505
R4301 GND.n6259 GND.n6258 4.6505
R4302 GND.n6255 GND.n6229 4.6505
R4303 GND.n6264 GND.n6230 4.6505
R4304 GND.n524 GND.n523 4.6505
R4305 GND.n526 GND.n525 4.6505
R4306 GND.n528 GND.n527 4.6505
R4307 GND.n530 GND.n529 4.6505
R4308 GND.n532 GND.n531 4.6505
R4309 GND.n534 GND.n533 4.6505
R4310 GND.n536 GND.n535 4.6505
R4311 GND.n538 GND.n537 4.6505
R4312 GND.n540 GND.n539 4.6505
R4313 GND.n542 GND.n541 4.6505
R4314 GND.n544 GND.n543 4.6505
R4315 GND.n546 GND.n545 4.6505
R4316 GND.n5880 GND.n5870 4.6505
R4317 GND.n5879 GND.n5871 4.6505
R4318 GND.n5952 GND.n5951 4.6505
R4319 GND.n5954 GND.n5953 4.6505
R4320 GND.n6131 GND.n5850 4.6505
R4321 GND.n6130 GND.n5851 4.6505
R4322 GND.n6033 GND.n6032 4.6505
R4323 GND.n6035 GND.n6034 4.6505
R4324 GND.n6081 GND.n6080 4.6505
R4325 GND.n6083 GND.n6082 4.6505
R4326 GND.n6093 GND.n6092 4.6505
R4327 GND.n5863 GND.n5862 4.6505
R4328 GND.n5867 GND.n5866 4.6505
R4329 GND.n5869 GND.n5868 4.6505
R4330 GND.n5909 GND.n5908 4.6505
R4331 GND.n5904 GND.n5903 4.6505
R4332 GND.n5900 GND.n5899 4.6505
R4333 GND.n5898 GND.n5897 4.6505
R4334 GND.n5894 GND.n5893 4.6505
R4335 GND.n5892 GND.n5891 4.6505
R4336 GND.n5888 GND.n5887 4.6505
R4337 GND.n5886 GND.n5885 4.6505
R4338 GND.n5882 GND.n5881 4.6505
R4339 GND.n5878 GND.n5877 4.6505
R4340 GND.n5876 GND.n5875 4.6505
R4341 GND.n5857 GND.n5856 4.6505
R4342 GND.n5919 GND.n5918 4.6505
R4343 GND.n5922 GND.n5921 4.6505
R4344 GND.n5926 GND.n5925 4.6505
R4345 GND.n5930 GND.n5929 4.6505
R4346 GND.n5932 GND.n5931 4.6505
R4347 GND.n5936 GND.n5935 4.6505
R4348 GND.n5938 GND.n5937 4.6505
R4349 GND.n5942 GND.n5941 4.6505
R4350 GND.n5944 GND.n5943 4.6505
R4351 GND.n5948 GND.n5947 4.6505
R4352 GND.n5950 GND.n5949 4.6505
R4353 GND.n5956 GND.n5955 4.6505
R4354 GND.n5960 GND.n5959 4.6505
R4355 GND.n5962 GND.n5961 4.6505
R4356 GND.n5967 GND.n5966 4.6505
R4357 GND.n5996 GND.n5995 4.6505
R4358 GND.n5993 GND.n5992 4.6505
R4359 GND.n5989 GND.n5988 4.6505
R4360 GND.n5985 GND.n5984 4.6505
R4361 GND.n5983 GND.n5982 4.6505
R4362 GND.n5979 GND.n5978 4.6505
R4363 GND.n5977 GND.n5976 4.6505
R4364 GND.n5973 GND.n5972 4.6505
R4365 GND.n5971 GND.n5970 4.6505
R4366 GND.n5849 GND.n5848 4.6505
R4367 GND.n6129 GND.n6128 4.6505
R4368 GND.n6127 GND.n6126 4.6505
R4369 GND.n6122 GND.n6121 4.6505
R4370 GND.n5855 GND.n5854 4.6505
R4371 GND.n6003 GND.n6002 4.6505
R4372 GND.n6007 GND.n6006 4.6505
R4373 GND.n6011 GND.n6010 4.6505
R4374 GND.n6013 GND.n6012 4.6505
R4375 GND.n6017 GND.n6016 4.6505
R4376 GND.n6019 GND.n6018 4.6505
R4377 GND.n6023 GND.n6022 4.6505
R4378 GND.n6025 GND.n6024 4.6505
R4379 GND.n6029 GND.n6028 4.6505
R4380 GND.n6031 GND.n6030 4.6505
R4381 GND.n6037 GND.n6036 4.6505
R4382 GND.n6041 GND.n6040 4.6505
R4383 GND.n6044 GND.n6043 4.6505
R4384 GND.n6049 GND.n6048 4.6505
R4385 GND.n6051 GND.n6050 4.6505
R4386 GND.n6055 GND.n6054 4.6505
R4387 GND.n6059 GND.n6058 4.6505
R4388 GND.n6061 GND.n6060 4.6505
R4389 GND.n6065 GND.n6064 4.6505
R4390 GND.n6067 GND.n6066 4.6505
R4391 GND.n6071 GND.n6070 4.6505
R4392 GND.n6073 GND.n6072 4.6505
R4393 GND.n6077 GND.n6076 4.6505
R4394 GND.n6079 GND.n6078 4.6505
R4395 GND.n6085 GND.n6084 4.6505
R4396 GND.n6088 GND.n6087 4.6505
R4397 GND.n6090 GND.n6089 4.6505
R4398 GND.n6113 GND.n6112 4.6505
R4399 GND.n6110 GND.n6109 4.6505
R4400 GND.n6108 GND.n6107 4.6505
R4401 GND.n6106 GND.n6105 4.6505
R4402 GND.n6104 GND.n6103 4.6505
R4403 GND.n6102 GND.n6101 4.6505
R4404 GND.n6098 GND.n6097 4.6505
R4405 GND.n7253 GND.n7243 4.6505
R4406 GND.n7252 GND.n7244 4.6505
R4407 GND.n7325 GND.n7324 4.6505
R4408 GND.n7327 GND.n7326 4.6505
R4409 GND.n7432 GND.n554 4.6505
R4410 GND.n7431 GND.n555 4.6505
R4411 GND.n7385 GND.n557 4.6505
R4412 GND.n7384 GND.n558 4.6505
R4413 GND.n569 GND.n559 4.6505
R4414 GND.n568 GND.n560 4.6505
R4415 GND.n2 GND.n1 4.6505
R4416 GND.n7236 GND.n7235 4.6505
R4417 GND.n7240 GND.n7239 4.6505
R4418 GND.n7242 GND.n7241 4.6505
R4419 GND.n7282 GND.n7281 4.6505
R4420 GND.n7277 GND.n7276 4.6505
R4421 GND.n7273 GND.n7272 4.6505
R4422 GND.n7271 GND.n7270 4.6505
R4423 GND.n7267 GND.n7266 4.6505
R4424 GND.n7265 GND.n7264 4.6505
R4425 GND.n7261 GND.n7260 4.6505
R4426 GND.n7259 GND.n7258 4.6505
R4427 GND.n7255 GND.n7254 4.6505
R4428 GND.n7251 GND.n7250 4.6505
R4429 GND.n7249 GND.n7248 4.6505
R4430 GND.n7231 GND.n7230 4.6505
R4431 GND.n7292 GND.n7291 4.6505
R4432 GND.n7295 GND.n7294 4.6505
R4433 GND.n7299 GND.n7298 4.6505
R4434 GND.n7303 GND.n7302 4.6505
R4435 GND.n7305 GND.n7304 4.6505
R4436 GND.n7309 GND.n7308 4.6505
R4437 GND.n7311 GND.n7310 4.6505
R4438 GND.n7315 GND.n7314 4.6505
R4439 GND.n7317 GND.n7316 4.6505
R4440 GND.n7321 GND.n7320 4.6505
R4441 GND.n7323 GND.n7322 4.6505
R4442 GND.n7329 GND.n7328 4.6505
R4443 GND.n7333 GND.n7332 4.6505
R4444 GND.n7335 GND.n7334 4.6505
R4445 GND.n7340 GND.n7339 4.6505
R4446 GND.n7369 GND.n7368 4.6505
R4447 GND.n7366 GND.n7365 4.6505
R4448 GND.n7362 GND.n7361 4.6505
R4449 GND.n7358 GND.n7357 4.6505
R4450 GND.n7356 GND.n7355 4.6505
R4451 GND.n7352 GND.n7351 4.6505
R4452 GND.n7350 GND.n7349 4.6505
R4453 GND.n7346 GND.n7345 4.6505
R4454 GND.n7344 GND.n7343 4.6505
R4455 GND.n553 GND.n552 4.6505
R4456 GND.n7430 GND.n7429 4.6505
R4457 GND.n7428 GND.n7427 4.6505
R4458 GND.n7423 GND.n7422 4.6505
R4459 GND.n7420 GND.n7419 4.6505
R4460 GND.n7415 GND.n7414 4.6505
R4461 GND.n7413 GND.n7412 4.6505
R4462 GND.n7409 GND.n7408 4.6505
R4463 GND.n7405 GND.n7404 4.6505
R4464 GND.n7403 GND.n7402 4.6505
R4465 GND.n7399 GND.n7398 4.6505
R4466 GND.n7397 GND.n7396 4.6505
R4467 GND.n7393 GND.n7392 4.6505
R4468 GND.n7391 GND.n7390 4.6505
R4469 GND.n7387 GND.n7386 4.6505
R4470 GND.n7383 GND.n7382 4.6505
R4471 GND.n7381 GND.n7380 4.6505
R4472 GND.n606 GND.n605 4.6505
R4473 GND.n603 GND.n602 4.6505
R4474 GND.n599 GND.n598 4.6505
R4475 GND.n597 GND.n596 4.6505
R4476 GND.n593 GND.n592 4.6505
R4477 GND.n589 GND.n588 4.6505
R4478 GND.n587 GND.n586 4.6505
R4479 GND.n583 GND.n582 4.6505
R4480 GND.n581 GND.n580 4.6505
R4481 GND.n577 GND.n576 4.6505
R4482 GND.n575 GND.n574 4.6505
R4483 GND.n571 GND.n570 4.6505
R4484 GND.n567 GND.n566 4.6505
R4485 GND.n565 GND.n564 4.6505
R4486 GND.n562 GND.n561 4.6505
R4487 GND.n7800 GND.n7799 4.6505
R4488 GND.n7803 GND.n7802 4.6505
R4489 GND.n7805 GND.n7804 4.6505
R4490 GND.n7807 GND.n7806 4.6505
R4491 GND.n7809 GND.n7808 4.6505
R4492 GND.n7813 GND.n7812 4.6505
R4493 GND.n7815 GND.n7814 4.6505
R4494 GND.n4639 GND.n4638 4.52281
R4495 GND.n1742 GND.n1596 4.51032
R4496 GND.n1442 GND.n1441 4.5005
R4497 GND.n1454 GND.n1448 4.5005
R4498 GND.n1530 GND.n1529 4.5005
R4499 GND.n1544 GND.n1538 4.5005
R4500 GND.n1026 GND.n1025 4.5005
R4501 GND.n1038 GND.n1031 4.5005
R4502 GND.n5633 GND.n1007 4.5005
R4503 GND.n1016 GND.n1010 4.5005
R4504 GND.n6534 GND.n6533 4.5005
R4505 GND.n6546 GND.n6539 4.5005
R4506 GND.n6506 GND.n6505 4.5005
R4507 GND.n6516 GND.n6510 4.5005
R4508 GND.n7545 GND.n7544 4.5005
R4509 GND.n7557 GND.n7550 4.5005
R4510 GND.n7517 GND.n7516 4.5005
R4511 GND.n7527 GND.n7521 4.5005
R4512 GND.n5082 GND.n5081 4.5005
R4513 GND.n5094 GND.n5088 4.5005
R4514 GND.n5217 GND.n5216 4.5005
R4515 GND.n5227 GND.n5221 4.5005
R4516 GND.n3293 GND.n3292 4.5005
R4517 GND.n3305 GND.n3299 4.5005
R4518 GND.n3482 GND.n3481 4.5005
R4519 GND.n3492 GND.n3486 4.5005
R4520 GND.n3448 GND.n3447 4.5005
R4521 GND.n3460 GND.n3453 4.5005
R4522 GND.n5451 GND.n1115 4.5005
R4523 GND.n1124 GND.n1118 4.5005
R4524 GND.n6788 GND.n6787 4.5005
R4525 GND.n6800 GND.n6793 4.5005
R4526 GND.n6816 GND.n6769 4.5005
R4527 GND.n6778 GND.n6772 4.5005
R4528 GND.n7111 GND.n7110 4.5005
R4529 GND.n7123 GND.n7116 4.5005
R4530 GND.n7083 GND.n7082 4.5005
R4531 GND.n7093 GND.n7087 4.5005
R4532 GND.n1848 GND.n1847 4.5005
R4533 GND.n1860 GND.n1853 4.5005
R4534 GND.n1984 GND.n1983 4.5005
R4535 GND.n1994 GND.n1988 4.5005
R4536 GND.n2183 GND.n2182 4.5005
R4537 GND.n2192 GND.n2185 4.5005
R4538 GND.n2307 GND.n2306 4.5005
R4539 GND.n2317 GND.n2311 4.5005
R4540 GND.n6942 GND.n6941 4.5005
R4541 GND.n6954 GND.n6947 4.5005
R4542 GND.n6970 GND.n6923 4.5005
R4543 GND.n6932 GND.n6926 4.5005
R4544 GND.n72 GND.n71 4.5005
R4545 GND.n84 GND.n77 4.5005
R4546 GND.n61 GND.n55 4.5005
R4547 GND.n4761 GND.n4760 4.5005
R4548 GND.n4773 GND.n4766 4.5005
R4549 GND.n4893 GND.n4892 4.5005
R4550 GND.n4903 GND.n4897 4.5005
R4551 GND.n7483 GND.n7482 4.5005
R4552 GND.n7495 GND.n7488 4.5005
R4553 GND.n7455 GND.n7454 4.5005
R4554 GND.n7465 GND.n7459 4.5005
R4555 GND.n7608 GND.n7607 4.5005
R4556 GND.n7620 GND.n7613 4.5005
R4557 GND.n7580 GND.n7579 4.5005
R4558 GND.n7590 GND.n7584 4.5005
R4559 GND.n4420 GND.n4223 4.5005
R4560 GND.n4420 GND.n4419 4.5005
R4561 GND.n4614 GND.n4613 4.4805
R4562 GND.n4602 GND.n4601 4.4805
R4563 GND.n7234 GND.n7233 4.45136
R4564 GND.n727 GND.n726 4.45136
R4565 GND.n5861 GND.n5860 4.45136
R4566 GND.n4089 GND.t653 4.41708
R4567 GND.n5403 GND.t191 4.41708
R4568 GND.n3190 GND.t616 4.41708
R4569 GND.n3083 GND.t932 4.41708
R4570 GND.n2965 GND.t444 4.41708
R4571 GND.n2644 GND.t190 4.41708
R4572 GND.n2170 GND.t709 4.41708
R4573 GND.n5425 GND.t619 4.41708
R4574 GND.n2479 GND.t442 4.41708
R4575 GND.n2813 GND.t655 4.41708
R4576 GND.n2973 GND.t705 4.41708
R4577 GND.n3184 GND.t187 4.41708
R4578 GND.n3564 GND.t935 4.41708
R4579 GND.n5072 GND.t620 4.41708
R4580 GND.n5413 GND.t445 4.41708
R4581 GND.n4105 GND.t708 4.41708
R4582 GND.n1286 GND.t931 4.35136
R4583 GND.n3081 GND.t443 4.35136
R4584 GND.n5426 GND.t933 4.35136
R4585 GND.n1841 GND.t656 4.35136
R4586 GND.n2176 GND.t618 4.35136
R4587 GND.n2485 GND.t706 4.35136
R4588 GND.n2650 GND.t505 4.35136
R4589 GND.n2963 GND.t188 4.35136
R4590 GND.n2971 GND.t652 4.35136
R4591 GND.n3182 GND.t934 4.35136
R4592 GND.n3562 GND.t617 4.35136
R4593 GND.n5404 GND.t707 4.35136
R4594 GND.n5073 GND.t441 4.35136
R4595 GND.n5411 GND.t189 4.35136
R4596 GND.n3937 GND.t504 4.35136
R4597 GND.n4106 GND.t654 4.35136
R4598 GND.n6228 GND.n6227 4.25025
R4599 GND.n49 GND.n48 4.06709
R4600 GND.n6373 GND.n6372 4.06709
R4601 GND.n11 GND.n10 4.06409
R4602 GND.n6333 GND.n6332 4.06409
R4603 GND.n13 GND.n11 4.0631
R4604 GND.n6335 GND.n6333 4.0631
R4605 GND.n7769 GND.n7758 4.05611
R4606 GND.n6309 GND.n6298 4.05611
R4607 GND.n703 GND.n701 3.98881
R4608 GND.n6254 GND.n6252 3.98881
R4609 GND.n3053 GND.n3052 3.9685
R4610 GND.n1260 GND.n1259 3.9685
R4611 GND.n4060 GND.n4059 3.9685
R4612 GND.n3873 GND.n3872 3.9685
R4613 GND.n4611 GND.n4610 3.84205
R4614 GND.n7765 GND.n7764 3.80559
R4615 GND.n660 GND.n658 3.80559
R4616 GND.n6305 GND.n6304 3.80559
R4617 GND.n6275 GND.n6273 3.80559
R4618 GND.n32 GND.n30 3.80083
R4619 GND.n6356 GND.n6354 3.80083
R4620 GND.n4404 GND.n4399 3.69035
R4621 GND.n2898 GND.n2890 3.63686
R4622 GND.n4257 GND.n4224 3.38533
R4623 GND.n4242 GND.n4240 3.20453
R4624 GND.n1445 GND.n1444 3.03311
R4625 GND.n1546 GND.n1536 3.03311
R4626 GND.n1029 GND.n1028 3.03311
R4627 GND.n5628 GND.n5627 3.03311
R4628 GND.n6537 GND.n6536 3.03311
R4629 GND.n6522 GND.n6521 3.03311
R4630 GND.n4002 GND.n4001 3.03311
R4631 GND.n4011 GND.n4010 3.03311
R4632 GND.n7548 GND.n7547 3.03311
R4633 GND.n7533 GND.n7532 3.03311
R4634 GND.n5085 GND.n5084 3.03311
R4635 GND.n5233 GND.n5232 3.03311
R4636 GND.n3296 GND.n3295 3.03311
R4637 GND.n3498 GND.n3497 3.03311
R4638 GND.n3451 GND.n3450 3.03311
R4639 GND.n5446 GND.n5445 3.03311
R4640 GND.n6791 GND.n6790 3.03311
R4641 GND.n6811 GND.n6810 3.03311
R4642 GND.n7114 GND.n7113 3.03311
R4643 GND.n7099 GND.n7098 3.03311
R4644 GND.n1851 GND.n1850 3.03311
R4645 GND.n2000 GND.n1999 3.03311
R4646 GND.n1402 GND.n1401 3.03311
R4647 GND.n1413 GND.n1412 3.03311
R4648 GND.n2071 GND.n2070 3.03311
R4649 GND.n2080 GND.n2079 3.03311
R4650 GND.n2195 GND.n2194 3.03311
R4651 GND.n2323 GND.n2322 3.03311
R4652 GND.n2393 GND.n2392 3.03311
R4653 GND.n2402 GND.n2401 3.03311
R4654 GND.n2551 GND.n2550 3.03311
R4655 GND.n2560 GND.n2559 3.03311
R4656 GND.n6945 GND.n6944 3.03311
R4657 GND.n6965 GND.n6964 3.03311
R4658 GND.n2714 GND.n2713 3.03311
R4659 GND.n2723 GND.n2722 3.03311
R4660 GND.n2827 GND.n2826 3.03311
R4661 GND.n2831 GND.n2830 3.03311
R4662 GND.n75 GND.n74 3.03311
R4663 GND.n64 GND.n53 3.03311
R4664 GND.n158 GND.n157 3.03311
R4665 GND.n162 GND.n161 3.03311
R4666 GND.n2988 GND.n2987 3.03311
R4667 GND.n2997 GND.n2996 3.03311
R4668 GND.n3097 GND.n3096 3.03311
R4669 GND.n3106 GND.n3105 3.03311
R4670 GND.n5304 GND.n5303 3.03311
R4671 GND.n5313 GND.n5312 3.03311
R4672 GND.n4764 GND.n4763 3.03311
R4673 GND.n4909 GND.n4908 3.03311
R4674 GND.n4979 GND.n4978 3.03311
R4675 GND.n4988 GND.n4987 3.03311
R4676 GND.n7486 GND.n7485 3.03311
R4677 GND.n7471 GND.n7470 3.03311
R4678 GND.n3585 GND.n3584 3.03311
R4679 GND.n3594 GND.n3593 3.03311
R4680 GND.n7611 GND.n7610 3.03311
R4681 GND.n7596 GND.n7595 3.03311
R4682 GND.n3793 GND.n3792 3.03311
R4683 GND.n3797 GND.n3796 3.03311
R4684 GND.n3211 GND.n3210 3.03311
R4685 GND.n3220 GND.n3219 3.03311
R4686 GND.n1198 GND.n1197 3.03311
R4687 GND.n1207 GND.n1206 3.03311
R4688 GND.n2844 GND 3.0005
R4689 GND.n1354 GND 3.0005
R4690 GND.n2103 GND 3.0005
R4691 GND.n2426 GND 3.0005
R4692 GND.n2583 GND 3.0005
R4693 GND.n2747 GND 3.0005
R4694 GND.n7679 GND 3.0005
R4695 GND.n3020 GND 3.0005
R4696 GND.n3130 GND 3.0005
R4697 GND.n1187 GND 3.0005
R4698 GND.n3201 GND 3.0005
R4699 GND.n5336 GND 3.0005
R4700 GND.n5012 GND 3.0005
R4701 GND.n3617 GND 3.0005
R4702 GND.n4034 GND 3.0005
R4703 GND.n3833 GND 3.0005
R4704 GND.n926 GND.t362 2.84655
R4705 GND.n2094 GND.n2093 2.5872
R4706 GND.n2574 GND.n2573 2.5872
R4707 GND.n2857 GND.n2856 2.5872
R4708 GND.n3011 GND.n3010 2.5872
R4709 GND.n1221 GND.n1220 2.5872
R4710 GND.n5327 GND.n5326 2.5872
R4711 GND.n3608 GND.n3607 2.5872
R4712 GND.n4025 GND.n4024 2.5872
R4713 GND.n2417 GND.n2416 2.56838
R4714 GND.n2738 GND.n2737 2.56838
R4715 GND.n7670 GND.n7669 2.56838
R4716 GND.n3121 GND.n3120 2.56838
R4717 GND.n3235 GND.n3234 2.56838
R4718 GND.n5003 GND.n5002 2.56838
R4719 GND.n3824 GND.n3823 2.56838
R4720 GND.n4210 GND.t1402 2.36824
R4721 GND.n4207 GND.t800 2.36824
R4722 GND.n7812 GND.n7811 2.25932
R4723 GND.n988 GND.n987 2.25932
R4724 GND.n6101 GND.n6100 2.25932
R4725 GND.n1344 GND.n1343 2.1579
R4726 GND.n1577 GND.n1576 1.93119
R4727 GND.n1576 GND.n1575 1.93119
R4728 GND.n2039 GND.n2038 1.93119
R4729 GND.n2038 GND.n2037 1.93119
R4730 GND.n2376 GND.n2375 1.93119
R4731 GND.n2375 GND.n2374 1.93119
R4732 GND.n2519 GND.n2518 1.93119
R4733 GND.n2518 GND.n2517 1.93119
R4734 GND.n2697 GND.n2696 1.93119
R4735 GND.n2696 GND.n2695 1.93119
R4736 GND.n2937 GND.n2936 1.93119
R4737 GND.n2936 GND.n2935 1.93119
R4738 GND.n142 GND.n141 1.93119
R4739 GND.n141 GND.n140 1.93119
R4740 GND.n1321 GND.n1320 1.93119
R4741 GND.n1320 GND.n1319 1.93119
R4742 GND.n5596 GND.n5595 1.93119
R4743 GND.n5595 GND.n5594 1.93119
R4744 GND.n1159 GND.n1158 1.93119
R4745 GND.n1158 GND.n1157 1.93119
R4746 GND.n3533 GND.n3532 1.93119
R4747 GND.n3532 GND.n3531 1.93119
R4748 GND.n5272 GND.n5271 1.93119
R4749 GND.n5271 GND.n5270 1.93119
R4750 GND.n4963 GND.n4962 1.93119
R4751 GND.n4962 GND.n4961 1.93119
R4752 GND.n3721 GND.n3720 1.93119
R4753 GND.n3720 GND.n3719 1.93119
R4754 GND.n3970 GND.n3969 1.93119
R4755 GND.n3969 GND.n3968 1.93119
R4756 GND.n3777 GND.n3776 1.93119
R4757 GND.n3776 GND.n3775 1.93119
R4758 GND.n4242 GND.n4241 1.85757
R4759 GND.n2890 GND.n2887 1.81868
R4760 GND.n5622 GND.n5621 1.74523
R4761 GND.n1343 GND.n650 1.74523
R4762 GND.n3992 GND.n304 1.71871
R4763 GND.n5294 GND.n5239 1.71871
R4764 GND.n3559 GND.n3504 1.71871
R4765 GND.n5440 GND.n5439 1.71871
R4766 GND.n2541 GND.n2486 1.71871
R4767 GND.n2061 GND.n2006 1.71871
R4768 GND.n2384 GND.n2329 1.71871
R4769 GND.n7735 GND.n7734 1.71871
R4770 GND.n4970 GND.n4915 1.71871
R4771 GND.n3729 GND.n508 1.71871
R4772 GND.n1594 GND.n1552 1.71871
R4773 GND.n4204 GND.n4203 1.70717
R4774 GND GND.n3180 1.65137
R4775 GND GND.n3079 1.65137
R4776 GND.n1432 GND.n1431 1.64041
R4777 GND.n2163 GND.n2162 1.64041
R4778 GND.n2472 GND.n2471 1.64041
R4779 GND.n2637 GND.n2636 1.64041
R4780 GND.n2806 GND.n2805 1.64041
R4781 GND.n2902 GND.n2901 1.64041
R4782 GND.n7729 GND.n7728 1.64041
R4783 GND.n3154 GND.n3153 1.64041
R4784 GND.n3261 GND.n3260 1.64041
R4785 GND.n5396 GND.n5395 1.64041
R4786 GND.n5065 GND.n5064 1.64041
R4787 GND.n3671 GND.n3670 1.64041
R4788 GND.n1431 GND.n1430 1.63319
R4789 GND.n2162 GND.n2161 1.63319
R4790 GND.n2471 GND.n2470 1.63319
R4791 GND.n2636 GND.n2635 1.63319
R4792 GND.n2805 GND.n2804 1.63319
R4793 GND.n2901 GND.n2900 1.63319
R4794 GND.n7728 GND.n7727 1.63319
R4795 GND.n3153 GND.n3152 1.63319
R4796 GND.n3260 GND.n3259 1.63319
R4797 GND.n5395 GND.n5394 1.63319
R4798 GND.n5064 GND.n5063 1.63319
R4799 GND.n3670 GND.n3669 1.63319
R4800 GND.n4426 GND.n4425 1.49383
R4801 GND.n7435 GND 1.48176
R4802 GND.n4256 GND.n4254 1.40675
R4803 GND.n4252 GND.n4227 1.40675
R4804 GND.n4239 GND.n4237 1.3822
R4805 GND.n4245 GND.n4244 1.3822
R4806 GND.n4749 GND.n4628 1.2805
R4807 GND.n4621 GND.n4620 1.2805
R4808 GND.n574 GND.n573 1.12991
R4809 GND.n7390 GND.n7389 1.12991
R4810 GND.n7343 GND.n7342 1.12991
R4811 GND.n7320 GND.n7319 1.12991
R4812 GND.n7258 GND.n7257 1.12991
R4813 GND.n1538 GND.n1537 1.12991
R4814 GND.n1010 GND.n1009 1.12991
R4815 GND.n6510 GND.n6509 1.12991
R4816 GND.n7521 GND.n7520 1.12991
R4817 GND.n5221 GND.n5220 1.12991
R4818 GND.n3486 GND.n3485 1.12991
R4819 GND.n1118 GND.n1117 1.12991
R4820 GND.n6772 GND.n6771 1.12991
R4821 GND.n7087 GND.n7086 1.12991
R4822 GND.n1988 GND.n1987 1.12991
R4823 GND.n2311 GND.n2310 1.12991
R4824 GND.n6926 GND.n6925 1.12991
R4825 GND.n55 GND.n54 1.12991
R4826 GND.n4897 GND.n4896 1.12991
R4827 GND.n7459 GND.n7458 1.12991
R4828 GND.n7584 GND.n7583 1.12991
R4829 GND.n5782 GND.n5781 1.12991
R4830 GND.n5711 GND.n5710 1.12991
R4831 GND.n6141 GND.n6140 1.12991
R4832 GND.n6194 GND.n6193 1.12991
R4833 GND.n5833 GND.n5832 1.12991
R4834 GND.n963 GND.n962 1.12991
R4835 GND.n893 GND.n892 1.12991
R4836 GND.n864 GND.n863 1.12991
R4837 GND.n800 GND.n799 1.12991
R4838 GND.n766 GND.n765 1.12991
R4839 GND.n6076 GND.n6075 1.12991
R4840 GND.n6028 GND.n6027 1.12991
R4841 GND.n5970 GND.n5969 1.12991
R4842 GND.n5947 GND.n5946 1.12991
R4843 GND.n5885 GND.n5884 1.12991
R4844 GND.n3178 GND.n3155 1.10214
R4845 GND.n3285 GND.n3262 1.10214
R4846 GND.n3902 GND.n3874 1.10164
R4847 GND.n5398 GND.n5397 1.10116
R4848 GND.n2904 GND.n2903 1.10116
R4849 GND.n2639 GND.n2638 1.10116
R4850 GND.n2165 GND.n2164 1.10116
R4851 GND.n1434 GND.n1433 1.10116
R4852 GND.n2474 GND.n2473 1.10116
R4853 GND.n2808 GND.n2807 1.10116
R4854 GND.n7731 GND.n7730 1.10116
R4855 GND.n5067 GND.n5066 1.10116
R4856 GND.n3673 GND.n3672 1.10116
R4857 GND.n4084 GND.n4061 1.10114
R4858 GND.n1284 GND.n1261 1.10114
R4859 GND.n3077 GND.n3054 1.10114
R4860 GND.n1387 GND.n1386 0.9605
R4861 GND.n2138 GND.n2137 0.9605
R4862 GND.n2146 GND.n2145 0.9605
R4863 GND.n2618 GND.n2617 0.9605
R4864 GND.n2620 GND.n2619 0.9605
R4865 GND.n2781 GND.n2780 0.9605
R4866 GND.n2789 GND.n2788 0.9605
R4867 GND.n122 GND.n121 0.9605
R4868 GND.n7712 GND.n7711 0.9605
R4869 GND.n3029 GND.n3028 0.9605
R4870 GND.n3037 GND.n3036 0.9605
R4871 GND.n1236 GND.n1235 0.9605
R4872 GND.n1244 GND.n1243 0.9605
R4873 GND.n5371 GND.n5370 0.9605
R4874 GND.n5379 GND.n5378 0.9605
R4875 GND.n5048 GND.n5047 0.9605
R4876 GND.n3654 GND.n3653 0.9605
R4877 GND.n3647 GND.n3646 0.9605
R4878 GND.n4044 GND.n4043 0.9605
R4879 GND.n3857 GND.n3856 0.9605
R4880 GND.n3853 GND.n3845 0.9605
R4881 GND.n1888 GND.n1887 0.932703
R4882 GND.n1925 GND.t395 0.932703
R4883 GND.n2213 GND.n2212 0.932703
R4884 GND.n2248 GND.t67 0.932703
R4885 GND.n7144 GND.n7143 0.932703
R4886 GND.n7174 GND.t922 0.932703
R4887 GND.n617 GND.n616 0.932703
R4888 GND.n7008 GND.t1435 0.932703
R4889 GND.n627 GND.n626 0.932703
R4890 GND.n6854 GND.t1255 0.932703
R4891 GND.n637 GND.n636 0.932703
R4892 GND.n6700 GND.t31 0.932703
R4893 GND.n644 GND.n643 0.932703
R4894 GND.n6630 GND.t37 0.932703
R4895 GND.n5556 GND.n5555 0.932703
R4896 GND.n5527 GND.t816 0.932703
R4897 GND.n3434 GND.n3433 0.932703
R4898 GND.n1093 GND.t416 0.932703
R4899 GND.n3340 GND.n3339 0.932703
R4900 GND.n3401 GND.t739 0.932703
R4901 GND.n5121 GND.n5120 0.932703
R4902 GND.n5161 GND.t496 0.932703
R4903 GND.n4800 GND.n4799 0.932703
R4904 GND.n4837 GND.t222 0.932703
R4905 GND.n423 GND.n422 0.932703
R4906 GND.n463 GND.t29 0.932703
R4907 GND.n312 GND.n311 0.932703
R4908 GND.n394 GND.t437 0.932703
R4909 GND.n211 GND.n210 0.932703
R4910 GND.n283 GND.t1485 0.932703
R4911 GND.n5422 GND.n5421 0.795683
R4912 GND.n2175 GND.n2174 0.795683
R4913 GND.n2484 GND.n2483 0.795683
R4914 GND.n2649 GND.n2648 0.795683
R4915 GND.n2818 GND.n2817 0.795683
R4916 GND.n2970 GND.n2969 0.795683
R4917 GND.n2978 GND.n2977 0.795683
R4918 GND.n3088 GND.n3087 0.795683
R4919 GND.n3189 GND.n3188 0.795683
R4920 GND.n3195 GND.n3194 0.795683
R4921 GND.n3569 GND.n3568 0.795683
R4922 GND.n3572 GND.n3571 0.795683
R4923 GND.n3575 GND.n3574 0.795683
R4924 GND.n5418 GND.n5417 0.795683
R4925 GND.n4102 GND.n4101 0.795683
R4926 GND.n5421 GND.n5420 0.795337
R4927 GND.n2174 GND.n2173 0.795337
R4928 GND.n2483 GND.n2482 0.795337
R4929 GND.n2648 GND.n2647 0.795337
R4930 GND.n2817 GND.n2816 0.795337
R4931 GND.n2969 GND.n2968 0.795337
R4932 GND.n2977 GND.n2976 0.795337
R4933 GND.n3087 GND.n3086 0.795337
R4934 GND.n3188 GND.n3187 0.795337
R4935 GND.n3194 GND.n3193 0.795337
R4936 GND.n3568 GND.n3567 0.795337
R4937 GND.n3571 GND.n3570 0.795337
R4938 GND.n3574 GND.n3573 0.795337
R4939 GND.n5417 GND.n5416 0.795337
R4940 GND.n4101 GND.n4100 0.795337
R4941 GND.n4098 GND.n4097 0.795337
R4942 GND.n4099 GND.n4098 0.795337
R4943 GND.n5658 GND.n5657 0.705542
R4944 GND.n7435 GND.n7434 0.701583
R4945 GND.n4191 GND.n4189 0.6255
R4946 GND.n4198 GND.n4196 0.614587
R4947 GND.n3181 GND.n3179 0.5645
R4948 GND.n3080 GND.n3078 0.5645
R4949 GND.n4234 GND.n4233 0.549071
R4950 GND.n4215 GND.n4214 0.54612
R4951 GND.n5203 GND.n5202 0.533636
R4952 GND.n3329 GND.n3322 0.533636
R4953 GND.n6829 GND.n6828 0.533636
R4954 GND.n7223 GND.n7222 0.533636
R4955 GND.n1970 GND.n1969 0.533636
R4956 GND.n2293 GND.n2292 0.533636
R4957 GND.n6983 GND.n6982 0.533636
R4958 GND.n6665 GND.n6664 0.533636
R4959 GND.n4879 GND.n4878 0.533636
R4960 GND.n510 GND.n507 0.533636
R4961 GND.n1517 GND.n1516 0.533636
R4962 GND.n6135 GND.n5847 0.53211
R4963 GND.n1595 GND.n1435 0.520438
R4964 GND.n2167 GND.n2166 0.520438
R4965 GND.n2476 GND.n2475 0.520438
R4966 GND.n2641 GND.n2640 0.520438
R4967 GND.n2810 GND.n2809 0.520438
R4968 GND.n2961 GND.n2905 0.520438
R4969 GND.n7733 GND.n7732 0.520438
R4970 GND.n5400 GND.n5399 0.520438
R4971 GND.n5069 GND.n5068 0.520438
R4972 GND.n3730 GND.n3674 0.520438
R4973 GND.n4086 GND.n4085 0.520438
R4974 GND.n3904 GND.n3903 0.520438
R4975 GND.n3560 GND.n3286 0.520438
R4976 GND.n5438 GND.n1285 0.520438
R4977 GND.n6760 GND.n630 0.498714
R4978 GND.n7068 GND.n610 0.498714
R4979 GND.n7135 GND.n7131 0.498714
R4980 GND.n6914 GND.n620 0.498714
R4981 GND.n6133 GND.n6132 0.48654
R4982 GND.n866 GND.n551 0.479239
R4983 GND.n1562 GND.n1561 0.436742
R4984 GND.n1561 GND.n1560 0.436742
R4985 GND.n2022 GND.n2021 0.436742
R4986 GND.n2021 GND.n2020 0.436742
R4987 GND.n2341 GND.n2340 0.436742
R4988 GND.n2340 GND.n2339 0.436742
R4989 GND.n2502 GND.n2501 0.436742
R4990 GND.n2501 GND.n2500 0.436742
R4991 GND.n2662 GND.n2661 0.436742
R4992 GND.n2661 GND.n2660 0.436742
R4993 GND.n2918 GND.n2917 0.436742
R4994 GND.n2917 GND.n2916 0.436742
R4995 GND.n99 GND.n98 0.436742
R4996 GND.n98 GND.n97 0.436742
R4997 GND.n1304 GND.n1303 0.436742
R4998 GND.n1303 GND.n1302 0.436742
R4999 GND.n5579 GND.n5578 0.436742
R5000 GND.n5578 GND.n5577 0.436742
R5001 GND.n1140 GND.n1139 0.436742
R5002 GND.n1139 GND.n1138 0.436742
R5003 GND.n3516 GND.n3515 0.436742
R5004 GND.n3515 GND.n3514 0.436742
R5005 GND.n5255 GND.n5254 0.436742
R5006 GND.n5254 GND.n5253 0.436742
R5007 GND.n4928 GND.n4927 0.436742
R5008 GND.n4927 GND.n4926 0.436742
R5009 GND.n3686 GND.n3685 0.436742
R5010 GND.n3685 GND.n3684 0.436742
R5011 GND.n3953 GND.n3952 0.436742
R5012 GND.n3952 GND.n3951 0.436742
R5013 GND.n3742 GND.n3741 0.436742
R5014 GND.n3741 GND.n3740 0.436742
R5015 GND.n4200 GND.n4199 0.427167
R5016 GND.n4436 GND.n4435 0.427167
R5017 GND.n1469 GND.n1468 0.425574
R5018 GND.n5463 GND.n5462 0.425574
R5019 GND.n5640 GND.n5639 0.425574
R5020 GND.n7565 GND.n7564 0.425574
R5021 GND.n5108 GND.n5107 0.425574
R5022 GND.n3317 GND.n3316 0.425574
R5023 GND.n3468 GND.n3467 0.425574
R5024 GND.n1874 GND.n1873 0.425574
R5025 GND.n6655 GND.n6654 0.425574
R5026 GND.n4787 GND.n4786 0.425574
R5027 GND.n7503 GND.n7502 0.425574
R5028 GND.n201 GND.n200 0.425574
R5029 GND.n7791 GND.n7790 0.414845
R5030 GND.n6376 GND.n6375 0.414845
R5031 GND.n5532 GND.n5515 0.38056
R5032 GND.n6635 GND.n6618 0.38056
R5033 GND.n399 GND.n382 0.38056
R5034 GND.n5166 GND.n5149 0.38056
R5035 GND.n3406 GND.n3389 0.38056
R5036 GND.n1098 GND.n1081 0.38056
R5037 GND.n6859 GND.n6842 0.38056
R5038 GND.n7179 GND.n7162 0.38056
R5039 GND.n1930 GND.n1913 0.38056
R5040 GND.n2253 GND.n2236 0.38056
R5041 GND.n7013 GND.n6996 0.38056
R5042 GND.n6705 GND.n6688 0.38056
R5043 GND.n4842 GND.n4825 0.38056
R5044 GND.n468 GND.n451 0.38056
R5045 GND.n288 GND.n271 0.38056
R5046 GND.n1508 GND.n1496 0.38056
R5047 GND.n4086 GND.n3992 0.378813
R5048 GND.n5400 GND.n5294 0.378813
R5049 GND.n3560 GND.n3559 0.378813
R5050 GND.n5439 GND.n5438 0.378813
R5051 GND.n2961 GND.n2960 0.378813
R5052 GND.n2641 GND.n2541 0.378813
R5053 GND.n2167 GND.n2061 0.378813
R5054 GND.n2476 GND.n2384 0.378813
R5055 GND.n2810 GND.n2705 0.378813
R5056 GND.n7734 GND.n7733 0.378813
R5057 GND.n5069 GND.n4970 0.378813
R5058 GND.n3730 GND.n3729 0.378813
R5059 GND.n3904 GND.n3785 0.378813
R5060 GND.n1595 GND.n1594 0.378813
R5061 GND.n5504 GND.n5502 0.377583
R5062 GND.n6607 GND.n6605 0.377583
R5063 GND.n371 GND.n369 0.377583
R5064 GND.n5138 GND.n5136 0.377583
R5065 GND.n3378 GND.n3376 0.377583
R5066 GND.n1070 GND.n1068 0.377583
R5067 GND.n1902 GND.n1900 0.377583
R5068 GND.n2225 GND.n2223 0.377583
R5069 GND.n6677 GND.n6675 0.377583
R5070 GND.n4814 GND.n4812 0.377583
R5071 GND.n440 GND.n438 0.377583
R5072 GND.n260 GND.n258 0.377583
R5073 GND.n1485 GND.n1483 0.377583
R5074 GND.n7380 GND.n7379 0.376971
R5075 GND.n7427 GND.n7426 0.376971
R5076 GND.n7332 GND.n7331 0.376971
R5077 GND.n7248 GND.n7247 0.376971
R5078 GND.n1529 GND.n1528 0.376971
R5079 GND.n1007 GND.n1006 0.376971
R5080 GND.n6505 GND.n6504 0.376971
R5081 GND.n7516 GND.n7515 0.376971
R5082 GND.n5216 GND.n5215 0.376971
R5083 GND.n3481 GND.n3480 0.376971
R5084 GND.n1115 GND.n1114 0.376971
R5085 GND.n6769 GND.n6768 0.376971
R5086 GND.n7082 GND.n7081 0.376971
R5087 GND.n1983 GND.n1982 0.376971
R5088 GND.n2306 GND.n2305 0.376971
R5089 GND.n6923 GND.n6922 0.376971
R5090 GND.n7747 GND.n7746 0.376971
R5091 GND.n4892 GND.n4891 0.376971
R5092 GND.n7454 GND.n7453 0.376971
R5093 GND.n7579 GND.n7578 0.376971
R5094 GND.n5818 GND.n5817 0.376971
R5095 GND.n5772 GND.n5771 0.376971
R5096 GND.n5723 GND.n5722 0.376971
R5097 GND.n6154 GND.n6153 0.376971
R5098 GND.n5661 GND.n5660 0.376971
R5099 GND.n719 GND.n718 0.376971
R5100 GND.n877 GND.n876 0.376971
R5101 GND.n790 GND.n789 0.376971
R5102 GND.n778 GND.n777 0.376971
R5103 GND.n6040 GND.n6039 0.376971
R5104 GND.n6126 GND.n6125 0.376971
R5105 GND.n5959 GND.n5958 0.376971
R5106 GND.n5875 GND.n5874 0.376971
R5107 GND.n7789 GND.n7788 0.375505
R5108 GND.n6377 GND.n6348 0.375505
R5109 GND.n5500 GND.n5497 0.3755
R5110 GND.n6603 GND.n6600 0.3755
R5111 GND.n367 GND.n364 0.3755
R5112 GND.n5134 GND.n5131 0.3755
R5113 GND.n3374 GND.n3371 0.3755
R5114 GND.n1066 GND.n1063 0.3755
R5115 GND.n6722 GND.n6720 0.3755
R5116 GND.n7030 GND.n7028 0.3755
R5117 GND.n1898 GND.n1895 0.3755
R5118 GND.n6876 GND.n6874 0.3755
R5119 GND.n6673 GND.n6670 0.3755
R5120 GND.n4810 GND.n4807 0.3755
R5121 GND.n436 GND.n433 0.3755
R5122 GND.n256 GND.n253 0.3755
R5123 GND.n1481 GND.n1478 0.3755
R5124 GND.n5492 GND.n5490 0.373417
R5125 GND.n6595 GND.n6593 0.373417
R5126 GND.n359 GND.n357 0.373417
R5127 GND.n4855 GND.n4853 0.373417
R5128 GND.n4853 GND.n4852 0.373417
R5129 GND.n5179 GND.n5177 0.373417
R5130 GND.n5177 GND.n5176 0.373417
R5131 GND.n3352 GND.n3350 0.373417
R5132 GND.n6730 GND.n6728 0.373417
R5133 GND.n6728 GND.n6727 0.373417
R5134 GND.n7038 GND.n7036 0.373417
R5135 GND.n7036 GND.n7035 0.373417
R5136 GND.n2269 GND.n2267 0.373417
R5137 GND.n2267 GND.n2266 0.373417
R5138 GND.n7199 GND.n7197 0.373417
R5139 GND.n7197 GND.n7196 0.373417
R5140 GND.n6884 GND.n6882 0.373417
R5141 GND.n6882 GND.n6881 0.373417
R5142 GND.n6572 GND.n6570 0.373417
R5143 GND.n6570 GND.n6569 0.373417
R5144 GND.n484 GND.n482 0.373417
R5145 GND.n482 GND.n481 0.373417
R5146 GND.n336 GND.n334 0.373417
R5147 GND.n334 GND.n333 0.373417
R5148 GND.n248 GND.n246 0.373417
R5149 GND.n1946 GND.n1944 0.373417
R5150 GND.n1944 GND.n1937 0.373417
R5151 GND.n1934 GND.n1933 0.366214
R5152 GND.n2263 GND.n2262 0.366214
R5153 GND.n7193 GND.n7192 0.366214
R5154 GND.n7032 GND.n7031 0.366214
R5155 GND.n6878 GND.n6877 0.366214
R5156 GND.n6724 GND.n6723 0.366214
R5157 GND.n6667 GND.n6666 0.366214
R5158 GND.n6597 GND.n6596 0.366214
R5159 GND.n5494 GND.n5493 0.366214
R5160 GND.n1060 GND.n1059 0.366214
R5161 GND.n3368 GND.n3367 0.366214
R5162 GND.n5128 GND.n5127 0.366214
R5163 GND.n478 GND.n477 0.366214
R5164 GND.n430 GND.n429 0.366214
R5165 GND.n361 GND.n360 0.366214
R5166 GND.n250 GND.n249 0.366214
R5167 GND.n5201 GND.n5200 0.355857
R5168 GND.n6906 GND.n6905 0.355857
R5169 GND.n7221 GND.n7220 0.355857
R5170 GND.n1968 GND.n1967 0.355857
R5171 GND.n2291 GND.n2290 0.355857
R5172 GND.n7060 GND.n7059 0.355857
R5173 GND.n6752 GND.n6751 0.355857
R5174 GND.n4877 GND.n4876 0.355857
R5175 GND.n506 GND.n505 0.355857
R5176 GND.n1515 GND.n1514 0.355857
R5177 GND.n2844 GND 0.354667
R5178 GND.n1354 GND 0.354667
R5179 GND.n2103 GND 0.354667
R5180 GND.n2426 GND 0.354667
R5181 GND.n2583 GND 0.354667
R5182 GND.n2747 GND 0.354667
R5183 GND.n7679 GND 0.354667
R5184 GND.n3020 GND 0.354667
R5185 GND.n3130 GND 0.354667
R5186 GND.n1187 GND 0.354667
R5187 GND.n3201 GND 0.354667
R5188 GND.n5336 GND 0.354667
R5189 GND.n5012 GND 0.354667
R5190 GND.n3617 GND 0.354667
R5191 GND.n4034 GND 0.354667
R5192 GND.n3833 GND 0.354667
R5193 GND.n4600 GND.n4217 0.352931
R5194 GND.n4587 GND.n4586 0.352931
R5195 GND.n4571 GND.n4570 0.352931
R5196 GND.n4556 GND.n4555 0.352931
R5197 GND.n4541 GND.n4540 0.352931
R5198 GND.n4526 GND.n4525 0.352931
R5199 GND.n4509 GND.n4508 0.352931
R5200 GND.n4494 GND.n4493 0.352931
R5201 GND.n4479 GND.n4478 0.352931
R5202 GND.n4464 GND.n4463 0.352931
R5203 GND.n4428 GND.n4427 0.352931
R5204 GND.n4410 GND.n4409 0.352931
R5205 GND.n4385 GND.n4384 0.352931
R5206 GND.n4370 GND.n4369 0.352931
R5207 GND.n4355 GND.n4354 0.352931
R5208 GND.n4340 GND.n4339 0.352931
R5209 GND.n4321 GND.n4320 0.352931
R5210 GND.n4306 GND.n4305 0.352931
R5211 GND.n4291 GND.n4290 0.352931
R5212 GND.n4276 GND.n4275 0.352931
R5213 GND.n4449 GND.n4448 0.347722
R5214 GND.n3425 GND.n1112 0.345738
R5215 GND.n5547 GND.n5546 0.345738
R5216 GND.n302 GND.n223 0.345738
R5217 GND.n3420 GND.n3343 0.345738
R5218 GND.n6763 GND.n6760 0.345738
R5219 GND.n7071 GND.n7068 0.345738
R5220 GND.n7135 GND.n7134 0.345738
R5221 GND.n6917 GND.n6914 0.345738
R5222 GND.n6649 GND.n6561 0.345738
R5223 GND.n413 GND.n325 0.345738
R5224 GND.n7627 GND.n195 0.345738
R5225 GND.n7784 GND.n50 0.33677
R5226 GND.n6378 GND.n6326 0.33677
R5227 GND.n6134 GND.n6133 0.336652
R5228 GND.n6451 GND 0.327423
R5229 GND.n548 GND 0.327423
R5230 GND.n6495 GND.n6494 0.326891
R5231 GND.n6404 GND.n6292 0.326891
R5232 GND.n6468 GND.n6467 0.325812
R5233 GND.n6406 GND.n6405 0.325812
R5234 GND.n4006 GND.n3994 0.321569
R5235 GND.n2863 GND.n2847 0.321569
R5236 GND.n1359 GND.n1358 0.321569
R5237 GND.n1408 GND.n1407 0.321569
R5238 GND.n2107 GND.n2106 0.321569
R5239 GND.n2075 GND.n2063 0.321569
R5240 GND.n2430 GND.n2429 0.321569
R5241 GND.n2397 GND.n2386 0.321569
R5242 GND.n2587 GND.n2586 0.321569
R5243 GND.n2555 GND.n2543 0.321569
R5244 GND.n2751 GND.n2750 0.321569
R5245 GND.n2718 GND.n2707 0.321569
R5246 GND.n2840 GND.n2839 0.321569
R5247 GND.n7683 GND.n7682 0.321569
R5248 GND.n7662 GND.n7660 0.321569
R5249 GND.n3024 GND.n3023 0.321569
R5250 GND.n2992 GND.n2980 0.321569
R5251 GND.n3134 GND.n3133 0.321569
R5252 GND.n3101 GND.n3090 0.321569
R5253 GND.n1227 GND.n1190 0.321569
R5254 GND.n3241 GND.n3204 0.321569
R5255 GND.n5340 GND.n5339 0.321569
R5256 GND.n5308 GND.n5296 0.321569
R5257 GND.n5016 GND.n5015 0.321569
R5258 GND.n4983 GND.n4972 0.321569
R5259 GND.n3621 GND.n3620 0.321569
R5260 GND.n3589 GND.n3577 0.321569
R5261 GND.n4038 GND.n4037 0.321569
R5262 GND.n3814 GND.n3806 0.321569
R5263 GND.n3837 GND.n3836 0.321569
R5264 GND.n3215 GND.n3197 0.321569
R5265 GND.n1202 GND.n1183 0.321569
R5266 GND.n5497 GND.n5492 0.321333
R5267 GND.n6600 GND.n6595 0.321333
R5268 GND.n364 GND.n359 0.321333
R5269 GND.n1063 GND.n1058 0.321333
R5270 GND.n6727 GND.n6722 0.321333
R5271 GND.n7035 GND.n7030 0.321333
R5272 GND.n7196 GND.n7191 0.321333
R5273 GND.n6881 GND.n6876 0.321333
R5274 GND.n253 GND.n248 0.321333
R5275 GND.n4624 GND.n4621 0.3205
R5276 GND.n6135 GND.n6134 0.31982
R5277 GND.n1435 GND.n1360 0.314812
R5278 GND.n2166 GND.n2108 0.314812
R5279 GND.n2475 GND.n2431 0.314812
R5280 GND.n2640 GND.n2588 0.314812
R5281 GND.n2809 GND.n2752 0.314812
R5282 GND.n2905 GND.n2864 0.314812
R5283 GND.n7732 GND.n7684 0.314812
R5284 GND.n5399 GND.n5341 0.314812
R5285 GND.n5068 GND.n5017 0.314812
R5286 GND.n3674 GND.n3622 0.314812
R5287 GND.n4085 GND.n4039 0.314812
R5288 GND.n3903 GND.n3838 0.314812
R5289 GND.n3286 GND.n3242 0.314812
R5290 GND.n1285 GND.n1228 0.314812
R5291 GND.n3179 GND.n3135 0.314812
R5292 GND.n3078 GND.n3025 0.314812
R5293 GND.n1056 GND.n1053 0.313
R5294 GND.n5483 GND.n5480 0.313
R5295 GND.n239 GND.n236 0.313
R5296 GND.n4869 GND.n4866 0.313
R5297 GND.n5193 GND.n5190 0.313
R5298 GND.n3366 GND.n3363 0.313
R5299 GND.n6744 GND.n6741 0.313
R5300 GND.n7052 GND.n7049 0.313
R5301 GND.n2283 GND.n2280 0.313
R5302 GND.n7213 GND.n7210 0.313
R5303 GND.n6898 GND.n6895 0.313
R5304 GND.n6586 GND.n6583 0.313
R5305 GND.n498 GND.n495 0.313
R5306 GND.n350 GND.n347 0.313
R5307 GND.n7647 GND.n7644 0.313
R5308 GND.n1960 GND.n1957 0.313
R5309 GND.n7434 GND.n551 0.309146
R5310 GND.n4603 GND.n4600 0.302583
R5311 GND.n5559 GND.n5467 0.300798
R5312 GND.n6556 GND.n648 0.300798
R5313 GND.n320 GND.n316 0.300798
R5314 GND.n3437 GND.n3424 0.300798
R5315 GND.n218 GND.n214 0.300798
R5316 GND GND.n49 0.295209
R5317 GND GND.n6373 0.295209
R5318 GND.n2844 GND.n2842 0.295052
R5319 GND.n1354 GND.n1352 0.295052
R5320 GND.n2103 GND.n2101 0.295052
R5321 GND.n2426 GND.n2424 0.295052
R5322 GND.n2583 GND.n2581 0.295052
R5323 GND.n2747 GND.n2745 0.295052
R5324 GND.n7679 GND.n7677 0.295052
R5325 GND.n3020 GND.n3018 0.295052
R5326 GND.n3130 GND.n3128 0.295052
R5327 GND.n1187 GND.n1185 0.295052
R5328 GND.n3201 GND.n3199 0.295052
R5329 GND.n5336 GND.n5334 0.295052
R5330 GND.n5012 GND.n5010 0.295052
R5331 GND.n3617 GND.n3615 0.295052
R5332 GND.n4034 GND.n4032 0.295052
R5333 GND.n3833 GND.n3831 0.295052
R5334 GND.n1476 GND.n1474 0.290381
R5335 GND.n5561 GND.n5559 0.290381
R5336 GND.n6556 GND.n6555 0.290381
R5337 GND.n320 GND.n319 0.290381
R5338 GND.n5126 GND.n5124 0.290381
R5339 GND.n3327 GND.n3325 0.290381
R5340 GND.n3439 GND.n3437 0.290381
R5341 GND.n6909 GND.n6908 0.290381
R5342 GND.n7149 GND.n7147 0.290381
R5343 GND.n1893 GND.n1891 0.290381
R5344 GND.n2218 GND.n2216 0.290381
R5345 GND.n7063 GND.n7062 0.290381
R5346 GND.n6755 GND.n6754 0.290381
R5347 GND.n4805 GND.n4803 0.290381
R5348 GND.n428 GND.n426 0.290381
R5349 GND.n218 GND.n217 0.290381
R5350 GND.n7436 GND.n7435 0.283189
R5351 GND.n6133 GND.n551 0.282159
R5352 GND.n6493 GND.n6492 0.280127
R5353 GND.n6403 GND.n6402 0.280127
R5354 GND.n4206 GND.n4205 0.270108
R5355 GND.n3079 GND 0.262544
R5356 GND.n3180 GND 0.262544
R5357 GND.n4637 GND.n4636 0.260982
R5358 GND.n4636 GND.n4635 0.2605
R5359 GND.n5429 GND 0.246986
R5360 GND.n5506 GND.n5504 0.24425
R5361 GND.n6609 GND.n6607 0.24425
R5362 GND.n373 GND.n371 0.24425
R5363 GND.n5140 GND.n5138 0.24425
R5364 GND.n3380 GND.n3378 0.24425
R5365 GND.n1072 GND.n1070 0.24425
R5366 GND.n6833 GND.n6831 0.24425
R5367 GND.n7153 GND.n7151 0.24425
R5368 GND.n1904 GND.n1902 0.24425
R5369 GND.n2227 GND.n2225 0.24425
R5370 GND.n6987 GND.n6985 0.24425
R5371 GND.n6679 GND.n6677 0.24425
R5372 GND.n4816 GND.n4814 0.24425
R5373 GND.n442 GND.n440 0.24425
R5374 GND.n262 GND.n260 0.24425
R5375 GND.n1487 GND.n1485 0.24425
R5376 GND.n5564 GND.n5464 0.243155
R5377 GND.n6551 GND.n649 0.243155
R5378 GND.n7563 GND.n7562 0.243155
R5379 GND.n5111 GND.n5109 0.243155
R5380 GND.n3330 GND.n3318 0.243155
R5381 GND.n3466 GND.n3465 0.243155
R5382 GND.n6766 GND.n6765 0.243155
R5383 GND.n7128 GND.n7073 0.243155
R5384 GND.n1877 GND.n1875 0.243155
R5385 GND.n2203 GND.n2201 0.243155
R5386 GND.n6920 GND.n6919 0.243155
R5387 GND.n6658 GND.n6656 0.243155
R5388 GND.n4790 GND.n4788 0.243155
R5389 GND.n7501 GND.n7500 0.243155
R5390 GND.n7626 GND.n7625 0.243155
R5391 GND.n1471 GND.n1470 0.243155
R5392 GND.n1044 GND.n1042 0.238893
R5393 GND.n5471 GND.n5469 0.238893
R5394 GND.n227 GND.n225 0.238893
R5395 GND.n4857 GND.n4855 0.238893
R5396 GND.n5181 GND.n5179 0.238893
R5397 GND.n3354 GND.n3352 0.238893
R5398 GND.n6732 GND.n6730 0.238893
R5399 GND.n7040 GND.n7038 0.238893
R5400 GND.n2271 GND.n2269 0.238893
R5401 GND.n7201 GND.n7199 0.238893
R5402 GND.n6886 GND.n6884 0.238893
R5403 GND.n6574 GND.n6572 0.238893
R5404 GND.n486 GND.n484 0.238893
R5405 GND.n338 GND.n336 0.238893
R5406 GND.n7635 GND.n7633 0.238893
R5407 GND.n1948 GND.n1946 0.238893
R5408 GND.n5741 GND 0.228789
R5409 GND.n34 GND.n30 0.226583
R5410 GND.n6358 GND.n6354 0.226583
R5411 GND.n5623 GND.n5566 0.224247
R5412 GND.n6549 GND.n6527 0.224247
R5413 GND.n7560 GND.n7538 0.224247
R5414 GND.n5238 GND.n5097 0.224247
R5415 GND.n3503 GND.n3332 0.224247
R5416 GND.n6806 GND.n6804 0.224247
R5417 GND.n7126 GND.n7104 0.224247
R5418 GND.n2005 GND.n1863 0.224247
R5419 GND.n2328 GND.n2198 0.224247
R5420 GND.n6960 GND.n6958 0.224247
R5421 GND.n7736 GND.n87 0.224247
R5422 GND.n4914 GND.n4776 0.224247
R5423 GND.n7498 GND.n7476 0.224247
R5424 GND.n7623 GND.n7601 0.224247
R5425 GND.n1551 GND.n1457 0.224247
R5426 GND.n5666 GND 0.209082
R5427 GND.n5564 GND.n5563 0.202208
R5428 GND.n6552 GND.n6551 0.202208
R5429 GND.n1111 GND.n1109 0.200996
R5430 GND.n5545 GND.n5543 0.200996
R5431 GND.n301 GND.n299 0.200996
R5432 GND.n5102 GND.n5100 0.200996
R5433 GND.n3311 GND.n3309 0.200996
R5434 GND.n3419 GND.n3417 0.200996
R5435 GND.n1868 GND.n1866 0.200996
R5436 GND.n6648 GND.n6646 0.200996
R5437 GND.n4781 GND.n4779 0.200996
R5438 GND.n412 GND.n410 0.200996
R5439 GND.n7631 GND.n7629 0.200996
R5440 GND.n1463 GND.n1461 0.200996
R5441 GND.n4014 GND.n3996 0.197423
R5442 GND.n1416 GND.n1396 0.197423
R5443 GND.n2083 GND.n2065 0.197423
R5444 GND.n2405 GND.n2387 0.197423
R5445 GND.n2563 GND.n2545 0.197423
R5446 GND.n2726 GND.n2708 0.197423
R5447 GND.n2835 GND.n2833 0.197423
R5448 GND.n7656 GND.n164 0.197423
R5449 GND.n3000 GND.n2982 0.197423
R5450 GND.n3109 GND.n3091 0.197423
R5451 GND.n5316 GND.n5298 0.197423
R5452 GND.n4991 GND.n4973 0.197423
R5453 GND.n3597 GND.n3579 0.197423
R5454 GND.n3802 GND.n3799 0.197423
R5455 GND.n3223 GND.n3205 0.197423
R5456 GND.n1210 GND.n1192 0.197423
R5457 GND.n4208 GND.n4207 0.196239
R5458 GND.n4210 GND.n4209 0.190273
R5459 GND.n7764 GND.n7761 0.189094
R5460 GND.n661 GND.n660 0.189094
R5461 GND.n6304 GND.n6301 0.189094
R5462 GND.n6276 GND.n6275 0.189094
R5463 GND.n4215 GND.n4210 0.188284
R5464 GND.n4752 GND.n4750 0.181849
R5465 GND.n1516 GND.n1515 0.181736
R5466 GND.n317 GND.n303 0.181736
R5467 GND.n5202 GND.n5201 0.181736
R5468 GND.n3329 GND.n3328 0.181736
R5469 GND.n3441 GND.n3440 0.181736
R5470 GND.n6906 GND.n6829 0.181736
R5471 GND.n7222 GND.n7221 0.181736
R5472 GND.n1969 GND.n1968 0.181736
R5473 GND.n2292 GND.n2291 0.181736
R5474 GND.n7060 GND.n6983 0.181736
R5475 GND.n6752 GND.n6665 0.181736
R5476 GND.n4878 GND.n4877 0.181736
R5477 GND.n507 GND.n506 0.181736
R5478 GND.n215 GND.n202 0.181736
R5479 GND.n5429 GND 0.180197
R5480 GND.n5430 GND 0.180197
R5481 GND.n5431 GND 0.180197
R5482 GND.n5432 GND 0.180197
R5483 GND.n5433 GND 0.180197
R5484 GND.n5434 GND 0.180197
R5485 GND.n5407 GND 0.180197
R5486 GND.n5408 GND 0.180197
R5487 GND GND.n5409 0.180197
R5488 GND.n4110 GND 0.180197
R5489 GND.n4109 GND 0.180197
R5490 GND GND.n1288 0.180197
R5491 GND GND.n5436 0.180197
R5492 GND.n4207 GND.n4206 0.178057
R5493 GND.n1516 GND.n1471 0.17675
R5494 GND.n7562 GND.n303 0.17675
R5495 GND.n5202 GND.n5111 0.17675
R5496 GND.n3330 GND.n3329 0.17675
R5497 GND.n3465 GND.n3441 0.17675
R5498 GND.n6829 GND.n6766 0.17675
R5499 GND.n7222 GND.n7128 0.17675
R5500 GND.n1969 GND.n1877 0.17675
R5501 GND.n2292 GND.n2203 0.17675
R5502 GND.n6983 GND.n6920 0.17675
R5503 GND.n6665 GND.n6658 0.17675
R5504 GND.n4878 GND.n4790 0.17675
R5505 GND.n7500 GND.n507 0.17675
R5506 GND.n7625 GND.n202 0.17675
R5507 GND.t214 GND.t916 0.176207
R5508 GND.n4249 GND.n4231 0.176207
R5509 GND.n3079 GND 0.175427
R5510 GND.n3180 GND 0.175427
R5511 GND.n5508 GND.n5506 0.171333
R5512 GND.n6611 GND.n6609 0.171333
R5513 GND.n375 GND.n373 0.171333
R5514 GND.n5142 GND.n5140 0.171333
R5515 GND.n3382 GND.n3380 0.171333
R5516 GND.n1074 GND.n1072 0.171333
R5517 GND.n6835 GND.n6833 0.171333
R5518 GND.n7155 GND.n7153 0.171333
R5519 GND.n1906 GND.n1904 0.171333
R5520 GND.n2229 GND.n2227 0.171333
R5521 GND.n6989 GND.n6987 0.171333
R5522 GND.n6681 GND.n6679 0.171333
R5523 GND.n4818 GND.n4816 0.171333
R5524 GND.n444 GND.n442 0.171333
R5525 GND.n264 GND.n262 0.171333
R5526 GND.n1489 GND.n1487 0.171333
R5527 GND.n5515 GND.n5512 0.16925
R5528 GND.n6618 GND.n6615 0.16925
R5529 GND.n382 GND.n379 0.16925
R5530 GND.n5149 GND.n5146 0.16925
R5531 GND.n3389 GND.n3386 0.16925
R5532 GND.n1081 GND.n1078 0.16925
R5533 GND.n6842 GND.n6839 0.16925
R5534 GND.n7162 GND.n7159 0.16925
R5535 GND.n1913 GND.n1910 0.16925
R5536 GND.n2236 GND.n2233 0.16925
R5537 GND.n6996 GND.n6993 0.16925
R5538 GND.n6688 GND.n6685 0.16925
R5539 GND.n4825 GND.n4822 0.16925
R5540 GND.n451 GND.n448 0.16925
R5541 GND.n271 GND.n268 0.16925
R5542 GND.n1496 GND.n1493 0.16925
R5543 GND.n550 GND 0.165163
R5544 GND.n1109 GND.n1107 0.164786
R5545 GND.n1107 GND.n1056 0.164786
R5546 GND.n5543 GND.n5541 0.164786
R5547 GND.n5541 GND.n5483 0.164786
R5548 GND.n299 GND.n297 0.164786
R5549 GND.n297 GND.n239 0.164786
R5550 GND.n4870 GND.n4869 0.164786
R5551 GND.n5194 GND.n5193 0.164786
R5552 GND.n3417 GND.n3415 0.164786
R5553 GND.n3415 GND.n3366 0.164786
R5554 GND.n6745 GND.n6709 0.164786
R5555 GND.n6745 GND.n6744 0.164786
R5556 GND.n7053 GND.n7017 0.164786
R5557 GND.n7053 GND.n7052 0.164786
R5558 GND.n2284 GND.n2283 0.164786
R5559 GND.n7214 GND.n7183 0.164786
R5560 GND.n7214 GND.n7213 0.164786
R5561 GND.n6899 GND.n6863 0.164786
R5562 GND.n6899 GND.n6898 0.164786
R5563 GND.n6646 GND.n6644 0.164786
R5564 GND.n6644 GND.n6586 0.164786
R5565 GND.n499 GND.n498 0.164786
R5566 GND.n410 GND.n408 0.164786
R5567 GND.n408 GND.n350 0.164786
R5568 GND.n7648 GND.n7631 0.164786
R5569 GND.n7648 GND.n7647 0.164786
R5570 GND.n1961 GND.n1960 0.164786
R5571 GND.n5563 GND.n5562 0.160043
R5572 GND.n6553 GND.n6552 0.160043
R5573 GND.n5534 GND.n5532 0.159429
R5574 GND.n6637 GND.n6635 0.159429
R5575 GND.n401 GND.n399 0.159429
R5576 GND.n5168 GND.n5166 0.159429
R5577 GND.n3408 GND.n3406 0.159429
R5578 GND.n1100 GND.n1098 0.159429
R5579 GND.n6861 GND.n6859 0.159429
R5580 GND.n7181 GND.n7179 0.159429
R5581 GND.n1932 GND.n1930 0.159429
R5582 GND.n2255 GND.n2253 0.159429
R5583 GND.n7015 GND.n7013 0.159429
R5584 GND.n6707 GND.n6705 0.159429
R5585 GND.n4844 GND.n4842 0.159429
R5586 GND.n470 GND.n468 0.159429
R5587 GND.n290 GND.n288 0.159429
R5588 GND.n1510 GND.n1508 0.159429
R5589 GND.n6451 GND.n6450 0.15606
R5590 GND.n548 GND.n547 0.15606
R5591 GND.n1053 GND.n1050 0.148714
R5592 GND.n1048 GND.n1044 0.148714
R5593 GND.n5480 GND.n5477 0.148714
R5594 GND.n5475 GND.n5471 0.148714
R5595 GND.n236 GND.n233 0.148714
R5596 GND.n231 GND.n227 0.148714
R5597 GND.n4866 GND.n4863 0.148714
R5598 GND.n4861 GND.n4857 0.148714
R5599 GND.n5190 GND.n5187 0.148714
R5600 GND.n5185 GND.n5181 0.148714
R5601 GND.n3363 GND.n3360 0.148714
R5602 GND.n3358 GND.n3354 0.148714
R5603 GND.n6741 GND.n6738 0.148714
R5604 GND.n6736 GND.n6732 0.148714
R5605 GND.n7049 GND.n7046 0.148714
R5606 GND.n7044 GND.n7040 0.148714
R5607 GND.n2280 GND.n2277 0.148714
R5608 GND.n2275 GND.n2271 0.148714
R5609 GND.n7210 GND.n7207 0.148714
R5610 GND.n7205 GND.n7201 0.148714
R5611 GND.n6895 GND.n6892 0.148714
R5612 GND.n6890 GND.n6886 0.148714
R5613 GND.n6583 GND.n6580 0.148714
R5614 GND.n6578 GND.n6574 0.148714
R5615 GND.n495 GND.n492 0.148714
R5616 GND.n490 GND.n486 0.148714
R5617 GND.n347 GND.n344 0.148714
R5618 GND.n342 GND.n338 0.148714
R5619 GND.n7644 GND.n7641 0.148714
R5620 GND.n7639 GND.n7635 0.148714
R5621 GND.n1957 GND.n1954 0.148714
R5622 GND.n1952 GND.n1948 0.148714
R5623 GND.n4753 GND.n4215 0.148287
R5624 GND.n1287 GND.n1286 0.142154
R5625 GND.n3082 GND.n3081 0.142154
R5626 GND.n5427 GND.n5426 0.142154
R5627 GND.n2169 GND.n1841 0.142154
R5628 GND.n2478 GND.n2176 0.142154
R5629 GND.n2643 GND.n2485 0.142154
R5630 GND.n2812 GND.n2650 0.142154
R5631 GND.n2964 GND.n2963 0.142154
R5632 GND.n2972 GND.n2971 0.142154
R5633 GND.n3183 GND.n3182 0.142154
R5634 GND.n3563 GND.n3562 0.142154
R5635 GND.n5405 GND.n5404 0.142154
R5636 GND.n5074 GND.n5073 0.142154
R5637 GND.n5412 GND.n5411 0.142154
R5638 GND.n4088 GND.n3937 0.142154
R5639 GND.n4107 GND.n4106 0.142154
R5640 GND.n4595 GND.n4594 0.141472
R5641 GND.n4594 GND.n4592 0.141472
R5642 GND.n4592 GND.n4579 0.141472
R5643 GND.n4579 GND.n4577 0.141472
R5644 GND.n4577 GND.n4564 0.141472
R5645 GND.n4564 GND.n4562 0.141472
R5646 GND.n4562 GND.n4549 0.141472
R5647 GND.n4549 GND.n4547 0.141472
R5648 GND.n4547 GND.n4534 0.141472
R5649 GND.n4534 GND.n4532 0.141472
R5650 GND.n4517 GND.n4515 0.141472
R5651 GND.n4515 GND.n4502 0.141472
R5652 GND.n4502 GND.n4500 0.141472
R5653 GND.n4500 GND.n4487 0.141472
R5654 GND.n4487 GND.n4485 0.141472
R5655 GND.n4485 GND.n4472 0.141472
R5656 GND.n4472 GND.n4470 0.141472
R5657 GND.n4470 GND.n4457 0.141472
R5658 GND.n4457 GND.n4455 0.141472
R5659 GND.n4437 GND.n4434 0.141472
R5660 GND.n4418 GND.n4416 0.141472
R5661 GND.n4416 GND.n4393 0.141472
R5662 GND.n4393 GND.n4391 0.141472
R5663 GND.n4391 GND.n4378 0.141472
R5664 GND.n4378 GND.n4376 0.141472
R5665 GND.n4376 GND.n4363 0.141472
R5666 GND.n4363 GND.n4361 0.141472
R5667 GND.n4361 GND.n4348 0.141472
R5668 GND.n4348 GND.n4346 0.141472
R5669 GND.n4330 GND.n4327 0.141472
R5670 GND.n4327 GND.n4314 0.141472
R5671 GND.n4314 GND.n4312 0.141472
R5672 GND.n4312 GND.n4299 0.141472
R5673 GND.n4299 GND.n4297 0.141472
R5674 GND.n4297 GND.n4284 0.141472
R5675 GND.n4284 GND.n4282 0.141472
R5676 GND.n4282 GND.n4269 0.141472
R5677 GND.n4269 GND.n4267 0.141472
R5678 GND.n2884 GND.n2883 0.140883
R5679 GND.n6452 GND 0.140869
R5680 GND.n549 GND 0.140869
R5681 GND.n4455 GND.n4440 0.136611
R5682 GND.n7791 GND 0.134348
R5683 GND.n6375 GND 0.134348
R5684 GND.n4230 GND.n4229 0.134262
R5685 GND.n1425 GND.n1424 0.131784
R5686 GND.n1426 GND.n1425 0.131784
R5687 GND.n2154 GND.n2153 0.131784
R5688 GND.n2465 GND.n2464 0.131784
R5689 GND.n2466 GND.n2465 0.131784
R5690 GND.n2628 GND.n2627 0.131784
R5691 GND.n2799 GND.n2798 0.131784
R5692 GND.n2800 GND.n2799 0.131784
R5693 GND.n2896 GND.n2895 0.131784
R5694 GND.n7722 GND.n7721 0.131784
R5695 GND.n7723 GND.n7722 0.131784
R5696 GND.n3045 GND.n3044 0.131784
R5697 GND.n3147 GND.n3146 0.131784
R5698 GND.n3148 GND.n3147 0.131784
R5699 GND.n1252 GND.n1251 0.131784
R5700 GND.n3254 GND.n3253 0.131784
R5701 GND.n3255 GND.n3254 0.131784
R5702 GND.n5387 GND.n5386 0.131784
R5703 GND.n5058 GND.n5057 0.131784
R5704 GND.n5059 GND.n5058 0.131784
R5705 GND.n3664 GND.n3663 0.131784
R5706 GND.n3665 GND.n3664 0.131784
R5707 GND.n4052 GND.n4051 0.131784
R5708 GND.n3865 GND.n3864 0.131784
R5709 GND.n2157 GND.n2154 0.13084
R5710 GND.n2631 GND.n2628 0.13084
R5711 GND.n2897 GND.n2896 0.13084
R5712 GND.n3048 GND.n3045 0.13084
R5713 GND.n1255 GND.n1252 0.13084
R5714 GND.n5390 GND.n5387 0.13084
R5715 GND.n4055 GND.n4052 0.13084
R5716 GND.n3868 GND.n3865 0.13084
R5717 GND.n6450 GND.n6449 0.12814
R5718 GND.n547 GND.n546 0.12814
R5719 GND.n4244 GND.n4242 0.127732
R5720 GND.n1393 GND.n1392 0.126877
R5721 GND.n2156 GND.n2155 0.126877
R5722 GND.n2460 GND.n2459 0.126877
R5723 GND.n2630 GND.n2629 0.126877
R5724 GND.n2794 GND.n2793 0.126877
R5725 GND.n2892 GND.n2891 0.126877
R5726 GND.n7717 GND.n7716 0.126877
R5727 GND.n3047 GND.n3046 0.126877
R5728 GND.n3142 GND.n3141 0.126877
R5729 GND.n1254 GND.n1253 0.126877
R5730 GND.n3249 GND.n3248 0.126877
R5731 GND.n5389 GND.n5388 0.126877
R5732 GND.n5053 GND.n5052 0.126877
R5733 GND.n3659 GND.n3658 0.126877
R5734 GND.n4054 GND.n4053 0.126877
R5735 GND.n3867 GND.n3866 0.126877
R5736 GND.n2157 GND.n2156 0.125988
R5737 GND.n2631 GND.n2630 0.125988
R5738 GND.n2897 GND.n2892 0.125988
R5739 GND.n3048 GND.n3047 0.125988
R5740 GND.n1255 GND.n1254 0.125988
R5741 GND.n5390 GND.n5389 0.125988
R5742 GND.n4055 GND.n4054 0.125988
R5743 GND.n3868 GND.n3867 0.125988
R5744 GND.n1427 GND.n1393 0.125687
R5745 GND.n2467 GND.n2460 0.125687
R5746 GND.n2801 GND.n2794 0.125687
R5747 GND.n7724 GND.n7717 0.125687
R5748 GND.n3149 GND.n3142 0.125687
R5749 GND.n3256 GND.n3249 0.125687
R5750 GND.n5060 GND.n5053 0.125687
R5751 GND.n3666 GND.n3659 0.125687
R5752 GND.n4346 GND.n4333 0.1255
R5753 GND.n7573 GND.n7572 0.122064
R5754 GND.n7510 GND.n7509 0.122064
R5755 GND.n7448 GND.n7447 0.122064
R5756 GND.n4886 GND.n4885 0.122064
R5757 GND.n5210 GND.n5209 0.122064
R5758 GND.n3475 GND.n3474 0.122064
R5759 GND.n5456 GND.n5455 0.122064
R5760 GND.n5638 GND.n5637 0.122064
R5761 GND.n6499 GND.n6498 0.122064
R5762 GND.n7751 GND.n7750 0.122064
R5763 GND.n6821 GND.n6820 0.122064
R5764 GND.n6975 GND.n6974 0.122064
R5765 GND.n7076 GND.n7075 0.122064
R5766 GND.n2300 GND.n2299 0.122064
R5767 GND.n1977 GND.n1976 0.122064
R5768 GND.n1523 GND.n1522 0.122064
R5769 GND.n4237 GND.n4235 0.118804
R5770 GND.n4754 GND.n4753 0.118
R5771 GND.n4182 GND.n4123 0.117638
R5772 GND.t26 GND.t212 0.117638
R5773 GND.t552 GND.t399 0.117638
R5774 GND.t211 GND.t59 0.117638
R5775 GND.t196 GND.t102 0.117638
R5776 GND.t75 GND.t889 0.117638
R5777 GND.t84 GND.t506 0.117638
R5778 GND.t119 GND.t693 0.117638
R5779 GND.t60 GND.t615 0.117638
R5780 GND.n4267 GND.n4261 0.117167
R5781 GND.n6446 GND.n6445 0.1155
R5782 GND.n6445 GND.n6443 0.1155
R5783 GND.n6440 GND.n6439 0.1155
R5784 GND.n6439 GND.n6437 0.1155
R5785 GND.n6434 GND.n6433 0.1155
R5786 GND.n6433 GND.n6431 0.1155
R5787 GND.n6428 GND.n6427 0.1155
R5788 GND.n6427 GND.n6425 0.1155
R5789 GND.n543 GND.n542 0.1155
R5790 GND.n542 GND.n540 0.1155
R5791 GND.n537 GND.n536 0.1155
R5792 GND.n536 GND.n534 0.1155
R5793 GND.n531 GND.n530 0.1155
R5794 GND.n530 GND.n528 0.1155
R5795 GND.n525 GND.n524 0.1155
R5796 GND.n524 GND.n522 0.1155
R5797 GND.n7563 GND.n302 0.112135
R5798 GND.n5109 GND.n5103 0.112135
R5799 GND.n3318 GND.n3312 0.112135
R5800 GND.n3466 GND.n3420 0.112135
R5801 GND.n6765 GND.n6763 0.112135
R5802 GND.n7073 GND.n7071 0.112135
R5803 GND.n1875 GND.n1869 0.112135
R5804 GND.n6919 GND.n6917 0.112135
R5805 GND.n6656 GND.n6649 0.112135
R5806 GND.n4788 GND.n4782 0.112135
R5807 GND.n7501 GND.n413 0.112135
R5808 GND.n7627 GND.n7626 0.112135
R5809 GND.n1470 GND.n1464 0.112135
R5810 GND.n49 GND.n25 0.110055
R5811 GND.n6373 GND.n6349 0.110055
R5812 GND.n1574 GND.n1573 0.10956
R5813 GND.n1573 GND.n1572 0.10956
R5814 GND.n1555 GND.n1554 0.10956
R5815 GND.n1554 GND.n1553 0.10956
R5816 GND.n1579 GND.n1578 0.10956
R5817 GND.t248 GND.n1579 0.10956
R5818 GND.n1584 GND.n1583 0.10956
R5819 GND.t248 GND.n1584 0.10956
R5820 GND.n2036 GND.n2035 0.10956
R5821 GND.n2035 GND.n2034 0.10956
R5822 GND.n2013 GND.n2012 0.10956
R5823 GND.n2012 GND.n2011 0.10956
R5824 GND.n2055 GND.n2054 0.10956
R5825 GND.t500 GND.n2055 0.10956
R5826 GND.t500 GND.n2053 0.10956
R5827 GND.n2053 GND.n2052 0.10956
R5828 GND.n2041 GND.n2040 0.10956
R5829 GND.t822 GND.n2041 0.10956
R5830 GND.n2047 GND.n2046 0.10956
R5831 GND.t822 GND.n2047 0.10956
R5832 GND.n2373 GND.n2372 0.10956
R5833 GND.n2372 GND.n2371 0.10956
R5834 GND.n2332 GND.n2331 0.10956
R5835 GND.n2331 GND.n2330 0.10956
R5836 GND.n2362 GND.n2361 0.10956
R5837 GND.t1089 GND.n2362 0.10956
R5838 GND.t1089 GND.n2360 0.10956
R5839 GND.n2360 GND.n2359 0.10956
R5840 GND.n2348 GND.n2347 0.10956
R5841 GND.t826 GND.n2348 0.10956
R5842 GND.n2354 GND.n2353 0.10956
R5843 GND.t826 GND.n2354 0.10956
R5844 GND.n2516 GND.n2515 0.10956
R5845 GND.n2515 GND.n2514 0.10956
R5846 GND.n2493 GND.n2492 0.10956
R5847 GND.n2492 GND.n2491 0.10956
R5848 GND.n2535 GND.n2534 0.10956
R5849 GND.t1415 GND.n2535 0.10956
R5850 GND.t1415 GND.n2533 0.10956
R5851 GND.n2533 GND.n2532 0.10956
R5852 GND.n2521 GND.n2520 0.10956
R5853 GND.t58 GND.n2521 0.10956
R5854 GND.n2527 GND.n2526 0.10956
R5855 GND.t58 GND.n2527 0.10956
R5856 GND.n2694 GND.n2693 0.10956
R5857 GND.n2693 GND.n2692 0.10956
R5858 GND.n2653 GND.n2652 0.10956
R5859 GND.n2652 GND.n2651 0.10956
R5860 GND.n2683 GND.n2682 0.10956
R5861 GND.t1239 GND.n2683 0.10956
R5862 GND.t1239 GND.n2681 0.10956
R5863 GND.n2681 GND.n2680 0.10956
R5864 GND.n2669 GND.n2668 0.10956
R5865 GND.t1096 GND.n2669 0.10956
R5866 GND.n2675 GND.n2674 0.10956
R5867 GND.t1096 GND.n2675 0.10956
R5868 GND.n2934 GND.n2933 0.10956
R5869 GND.n2933 GND.n2932 0.10956
R5870 GND.n2909 GND.n2908 0.10956
R5871 GND.n2908 GND.n2907 0.10956
R5872 GND.n2953 GND.n2952 0.10956
R5873 GND.t1230 GND.n2953 0.10956
R5874 GND.t1230 GND.n2951 0.10956
R5875 GND.n2951 GND.n2950 0.10956
R5876 GND.n2939 GND.n2938 0.10956
R5877 GND.t576 GND.n2939 0.10956
R5878 GND.n2945 GND.n2944 0.10956
R5879 GND.t576 GND.n2945 0.10956
R5880 GND.n139 GND.n138 0.10956
R5881 GND.n138 GND.n137 0.10956
R5882 GND.n90 GND.n89 0.10956
R5883 GND.n89 GND.n88 0.10956
R5884 GND.n128 GND.n127 0.10956
R5885 GND.t249 GND.n128 0.10956
R5886 GND.t249 GND.n126 0.10956
R5887 GND.n126 GND.n125 0.10956
R5888 GND.n106 GND.n105 0.10956
R5889 GND.t484 GND.n106 0.10956
R5890 GND.n112 GND.n111 0.10956
R5891 GND.t484 GND.n112 0.10956
R5892 GND.n1318 GND.n1317 0.10956
R5893 GND.n1317 GND.n1316 0.10956
R5894 GND.n1295 GND.n1294 0.10956
R5895 GND.n1294 GND.n1293 0.10956
R5896 GND.n1337 GND.n1336 0.10956
R5897 GND.t1399 GND.n1337 0.10956
R5898 GND.t1399 GND.n1335 0.10956
R5899 GND.n1335 GND.n1334 0.10956
R5900 GND.n1323 GND.n1322 0.10956
R5901 GND.t578 GND.n1323 0.10956
R5902 GND.n1329 GND.n1328 0.10956
R5903 GND.t578 GND.n1329 0.10956
R5904 GND.n5593 GND.n5592 0.10956
R5905 GND.n5592 GND.n5591 0.10956
R5906 GND.n5570 GND.n5569 0.10956
R5907 GND.n5569 GND.n5568 0.10956
R5908 GND.n5612 GND.n5611 0.10956
R5909 GND.t108 GND.n5612 0.10956
R5910 GND.t108 GND.n5610 0.10956
R5911 GND.n5610 GND.n5609 0.10956
R5912 GND.n5598 GND.n5597 0.10956
R5913 GND.t1243 GND.n5598 0.10956
R5914 GND.n5604 GND.n5603 0.10956
R5915 GND.t1243 GND.n5604 0.10956
R5916 GND.n1156 GND.n1155 0.10956
R5917 GND.n1155 GND.n1154 0.10956
R5918 GND.n1131 GND.n1130 0.10956
R5919 GND.n1130 GND.n1129 0.10956
R5920 GND.n1175 GND.n1174 0.10956
R5921 GND.t947 GND.n1175 0.10956
R5922 GND.t947 GND.n1173 0.10956
R5923 GND.n1173 GND.n1172 0.10956
R5924 GND.n1161 GND.n1160 0.10956
R5925 GND.t1513 GND.n1161 0.10956
R5926 GND.n1167 GND.n1166 0.10956
R5927 GND.t1513 GND.n1167 0.10956
R5928 GND.n3530 GND.n3529 0.10956
R5929 GND.n3529 GND.n3528 0.10956
R5930 GND.n3507 GND.n3506 0.10956
R5931 GND.n3506 GND.n3505 0.10956
R5932 GND.n3549 GND.n3548 0.10956
R5933 GND.t657 GND.n3549 0.10956
R5934 GND.t657 GND.n3547 0.10956
R5935 GND.n3547 GND.n3546 0.10956
R5936 GND.n3535 GND.n3534 0.10956
R5937 GND.t246 GND.n3535 0.10956
R5938 GND.n3541 GND.n3540 0.10956
R5939 GND.t246 GND.n3541 0.10956
R5940 GND.n5269 GND.n5268 0.10956
R5941 GND.n5268 GND.n5267 0.10956
R5942 GND.n5246 GND.n5245 0.10956
R5943 GND.n5245 GND.n5244 0.10956
R5944 GND.n5288 GND.n5287 0.10956
R5945 GND.t1419 GND.n5288 0.10956
R5946 GND.t1419 GND.n5286 0.10956
R5947 GND.n5286 GND.n5285 0.10956
R5948 GND.n5274 GND.n5273 0.10956
R5949 GND.t47 GND.n5274 0.10956
R5950 GND.n5280 GND.n5279 0.10956
R5951 GND.t47 GND.n5280 0.10956
R5952 GND.n4960 GND.n4959 0.10956
R5953 GND.n4959 GND.n4958 0.10956
R5954 GND.n4919 GND.n4918 0.10956
R5955 GND.n4918 GND.n4917 0.10956
R5956 GND.n4949 GND.n4948 0.10956
R5957 GND.t427 GND.n4949 0.10956
R5958 GND.t427 GND.n4947 0.10956
R5959 GND.n4947 GND.n4946 0.10956
R5960 GND.n4935 GND.n4934 0.10956
R5961 GND.t199 GND.n4935 0.10956
R5962 GND.n4941 GND.n4940 0.10956
R5963 GND.t199 GND.n4941 0.10956
R5964 GND.n3718 GND.n3717 0.10956
R5965 GND.n3717 GND.n3716 0.10956
R5966 GND.n3677 GND.n3676 0.10956
R5967 GND.n3676 GND.n3675 0.10956
R5968 GND.n3707 GND.n3706 0.10956
R5969 GND.t1241 GND.n3707 0.10956
R5970 GND.t1241 GND.n3705 0.10956
R5971 GND.n3705 GND.n3704 0.10956
R5972 GND.n3693 GND.n3692 0.10956
R5973 GND.t809 GND.n3693 0.10956
R5974 GND.n3699 GND.n3698 0.10956
R5975 GND.t809 GND.n3699 0.10956
R5976 GND.n3967 GND.n3966 0.10956
R5977 GND.n3966 GND.n3965 0.10956
R5978 GND.n3944 GND.n3943 0.10956
R5979 GND.n3943 GND.n3942 0.10956
R5980 GND.n3986 GND.n3985 0.10956
R5981 GND.t874 GND.n3986 0.10956
R5982 GND.t874 GND.n3984 0.10956
R5983 GND.n3984 GND.n3983 0.10956
R5984 GND.n3972 GND.n3971 0.10956
R5985 GND.t796 GND.n3972 0.10956
R5986 GND.n3978 GND.n3977 0.10956
R5987 GND.t796 GND.n3978 0.10956
R5988 GND.n4395 GND.n4394 0.10956
R5989 GND.n4396 GND.n4395 0.10956
R5990 GND.n4403 GND.n4402 0.10956
R5991 GND.n4404 GND.n4403 0.10956
R5992 GND.n3749 GND.n3748 0.10956
R5993 GND.t23 GND.n3749 0.10956
R5994 GND.n3755 GND.n3754 0.10956
R5995 GND.t23 GND.n3755 0.10956
R5996 GND.n3774 GND.n3773 0.10956
R5997 GND.n3773 GND.n3772 0.10956
R5998 GND.n3733 GND.n3732 0.10956
R5999 GND.n3732 GND.n3731 0.10956
R6000 GND.n3763 GND.n3762 0.10956
R6001 GND.t1225 GND.n3763 0.10956
R6002 GND.t1225 GND.n3761 0.10956
R6003 GND.n3761 GND.n3760 0.10956
R6004 GND.n3850 GND.t679 0.10956
R6005 GND.n3848 GND.n3847 0.10956
R6006 GND.t679 GND.n3848 0.10956
R6007 GND.n3851 GND.n3850 0.10956
R6008 GND.n1505 GND.n1504 0.10956
R6009 GND.n1504 GND.n1503 0.10956
R6010 GND.n1924 GND.n1923 0.10956
R6011 GND.t395 GND.n1924 0.10956
R6012 GND.n1927 GND.n1926 0.10956
R6013 GND.n1926 GND.n1925 0.10956
R6014 GND.n2247 GND.n2246 0.10956
R6015 GND.t67 GND.n2247 0.10956
R6016 GND.n2250 GND.n2249 0.10956
R6017 GND.n2249 GND.n2248 0.10956
R6018 GND.n7173 GND.n7172 0.10956
R6019 GND.t922 GND.n7173 0.10956
R6020 GND.n7176 GND.n7175 0.10956
R6021 GND.n7175 GND.n7174 0.10956
R6022 GND.n7007 GND.n7006 0.10956
R6023 GND.t1435 GND.n7007 0.10956
R6024 GND.n7010 GND.n7009 0.10956
R6025 GND.n7009 GND.n7008 0.10956
R6026 GND.n6853 GND.n6852 0.10956
R6027 GND.t1255 GND.n6853 0.10956
R6028 GND.n6856 GND.n6855 0.10956
R6029 GND.n6855 GND.n6854 0.10956
R6030 GND.n6699 GND.n6698 0.10956
R6031 GND.t31 GND.n6699 0.10956
R6032 GND.n6702 GND.n6701 0.10956
R6033 GND.n6701 GND.n6700 0.10956
R6034 GND.n6629 GND.n6628 0.10956
R6035 GND.t37 GND.n6629 0.10956
R6036 GND.n6632 GND.n6631 0.10956
R6037 GND.n6631 GND.n6630 0.10956
R6038 GND.n5526 GND.n5525 0.10956
R6039 GND.t816 GND.n5526 0.10956
R6040 GND.n5529 GND.n5528 0.10956
R6041 GND.n5528 GND.n5527 0.10956
R6042 GND.n1092 GND.n1091 0.10956
R6043 GND.t416 GND.n1092 0.10956
R6044 GND.n1095 GND.n1094 0.10956
R6045 GND.n1094 GND.n1093 0.10956
R6046 GND.n3400 GND.n3399 0.10956
R6047 GND.t739 GND.n3400 0.10956
R6048 GND.n3403 GND.n3402 0.10956
R6049 GND.n3402 GND.n3401 0.10956
R6050 GND.n5160 GND.n5159 0.10956
R6051 GND.t496 GND.n5160 0.10956
R6052 GND.n5163 GND.n5162 0.10956
R6053 GND.n5162 GND.n5161 0.10956
R6054 GND.n4836 GND.n4835 0.10956
R6055 GND.t222 GND.n4836 0.10956
R6056 GND.n4839 GND.n4838 0.10956
R6057 GND.n4838 GND.n4837 0.10956
R6058 GND.n462 GND.n461 0.10956
R6059 GND.t29 GND.n462 0.10956
R6060 GND.n465 GND.n464 0.10956
R6061 GND.n464 GND.n463 0.10956
R6062 GND.n393 GND.n392 0.10956
R6063 GND.t437 GND.n393 0.10956
R6064 GND.n396 GND.n395 0.10956
R6065 GND.n395 GND.n394 0.10956
R6066 GND.n282 GND.n281 0.10956
R6067 GND.t1485 GND.n282 0.10956
R6068 GND.n285 GND.n284 0.10956
R6069 GND.n284 GND.n283 0.10956
R6070 GND.n186 GND.n185 0.10956
R6071 GND.t1429 GND.n186 0.10956
R6072 GND.n5464 GND.n1112 0.107827
R6073 GND.n5546 GND.n649 0.107827
R6074 GND.n4109 GND 0.104579
R6075 GND.n1567 GND.n1566 0.104537
R6076 GND.n1566 GND.n1565 0.104537
R6077 GND.n2027 GND.n2026 0.104537
R6078 GND.n2026 GND.n2025 0.104537
R6079 GND.n2346 GND.n2345 0.104537
R6080 GND.n2345 GND.n2344 0.104537
R6081 GND.n2507 GND.n2506 0.104537
R6082 GND.n2506 GND.n2505 0.104537
R6083 GND.n2667 GND.n2666 0.104537
R6084 GND.n2666 GND.n2665 0.104537
R6085 GND.n2923 GND.n2922 0.104537
R6086 GND.n2922 GND.n2921 0.104537
R6087 GND.n104 GND.n103 0.104537
R6088 GND.n103 GND.n102 0.104537
R6089 GND.n1309 GND.n1308 0.104537
R6090 GND.n1308 GND.n1307 0.104537
R6091 GND.n5584 GND.n5583 0.104537
R6092 GND.n5583 GND.n5582 0.104537
R6093 GND.n1145 GND.n1144 0.104537
R6094 GND.n1144 GND.n1143 0.104537
R6095 GND.n3521 GND.n3520 0.104537
R6096 GND.n3520 GND.n3519 0.104537
R6097 GND.n5260 GND.n5259 0.104537
R6098 GND.n5259 GND.n5258 0.104537
R6099 GND.n4933 GND.n4932 0.104537
R6100 GND.n4932 GND.n4931 0.104537
R6101 GND.n3691 GND.n3690 0.104537
R6102 GND.n3690 GND.n3689 0.104537
R6103 GND.n3958 GND.n3957 0.104537
R6104 GND.n3957 GND.n3956 0.104537
R6105 GND.n3747 GND.n3746 0.104537
R6106 GND.n3746 GND.n3745 0.104537
R6107 GND.n6348 GND.n6327 0.102336
R6108 GND.n7788 GND.n7787 0.102336
R6109 GND.n5464 GND.n5463 0.102333
R6110 GND.n5639 GND.n649 0.102333
R6111 GND.n7564 GND.n7563 0.102333
R6112 GND.n5109 GND.n5108 0.102333
R6113 GND.n3318 GND.n3317 0.102333
R6114 GND.n3467 GND.n3466 0.102333
R6115 GND.n6765 GND.n6764 0.102333
R6116 GND.n7073 GND.n7072 0.102333
R6117 GND.n1875 GND.n1874 0.102333
R6118 GND.n2201 GND.n2200 0.102333
R6119 GND.n6919 GND.n6918 0.102333
R6120 GND.n6656 GND.n6655 0.102333
R6121 GND.n4788 GND.n4787 0.102333
R6122 GND.n7502 GND.n7501 0.102333
R6123 GND.n7626 GND.n201 0.102333
R6124 GND.n1470 GND.n1469 0.102333
R6125 GND.n7770 GND 0.101889
R6126 GND.n6310 GND 0.101889
R6127 GND.n4753 GND 0.0991625
R6128 GND.n35 GND.n34 0.0963333
R6129 GND.n36 GND.n27 0.0963333
R6130 GND.n42 GND.n27 0.0963333
R6131 GND.n43 GND.n42 0.0963333
R6132 GND.n44 GND.n43 0.0963333
R6133 GND.n6359 GND.n6358 0.0963333
R6134 GND.n6360 GND.n6351 0.0963333
R6135 GND.n6366 GND.n6351 0.0963333
R6136 GND.n6367 GND.n6366 0.0963333
R6137 GND.n6368 GND.n6367 0.0963333
R6138 GND.n4401 GND.n4400 0.0944005
R6139 GND.n1520 GND.n1519 0.0944005
R6140 GND.n1521 GND.n1520 0.0944005
R6141 GND.n1466 GND.n1465 0.0944005
R6142 GND.n1973 GND.n1972 0.0944005
R6143 GND.n1974 GND.n1973 0.0944005
R6144 GND.n1871 GND.n1870 0.0944005
R6145 GND.n2296 GND.n2295 0.0944005
R6146 GND.n2297 GND.n2296 0.0944005
R6147 GND.n7227 GND.n607 0.0944005
R6148 GND.n7226 GND.n7225 0.0944005
R6149 GND.n7227 GND.n7226 0.0944005
R6150 GND.n6978 GND.n6977 0.0944005
R6151 GND.n6980 GND.n6979 0.0944005
R6152 GND.n6979 GND.n6978 0.0944005
R6153 GND.n6824 GND.n6823 0.0944005
R6154 GND.n6826 GND.n6825 0.0944005
R6155 GND.n6825 GND.n6824 0.0944005
R6156 GND.n6660 GND.n6659 0.0944005
R6157 GND.n6662 GND.n6661 0.0944005
R6158 GND.n6661 GND.n6660 0.0944005
R6159 GND.n6652 GND.n6651 0.0944005
R6160 GND.n6651 GND.n6650 0.0944005
R6161 GND.n646 GND.n645 0.0944005
R6162 GND.n5643 GND.n5642 0.0944005
R6163 GND.n5645 GND.n5643 0.0944005
R6164 GND.n5645 GND.n5644 0.0944005
R6165 GND.n5460 GND.n5459 0.0944005
R6166 GND.n5459 GND.n5458 0.0944005
R6167 GND.n3422 GND.n3421 0.0944005
R6168 GND.n3471 GND.n3470 0.0944005
R6169 GND.n3472 GND.n3471 0.0944005
R6170 GND.n3320 GND.n3319 0.0944005
R6171 GND.n3314 GND.n3313 0.0944005
R6172 GND.n5206 GND.n5205 0.0944005
R6173 GND.n5207 GND.n5206 0.0944005
R6174 GND.n5105 GND.n5104 0.0944005
R6175 GND.n4882 GND.n4881 0.0944005
R6176 GND.n4883 GND.n4882 0.0944005
R6177 GND.n4784 GND.n4783 0.0944005
R6178 GND.n513 GND.n512 0.0944005
R6179 GND.n514 GND.n513 0.0944005
R6180 GND.n7506 GND.n7505 0.0944005
R6181 GND.n7507 GND.n7506 0.0944005
R6182 GND.n314 GND.n313 0.0944005
R6183 GND.n7568 GND.n7567 0.0944005
R6184 GND.n7570 GND.n7568 0.0944005
R6185 GND.n7570 GND.n7569 0.0944005
R6186 GND.n198 GND.n197 0.0944005
R6187 GND.n197 GND.n196 0.0944005
R6188 GND.n1452 GND.n1450 0.0921667
R6189 GND.n1035 GND.n1033 0.0921667
R6190 GND.n6543 GND.n6541 0.0921667
R6191 GND.n7554 GND.n7552 0.0921667
R6192 GND.n5092 GND.n5090 0.0921667
R6193 GND.n3303 GND.n3301 0.0921667
R6194 GND.n3457 GND.n3455 0.0921667
R6195 GND.n6797 GND.n6795 0.0921667
R6196 GND.n7120 GND.n7118 0.0921667
R6197 GND.n1857 GND.n1855 0.0921667
R6198 GND.n2189 GND.n2187 0.0921667
R6199 GND.n6951 GND.n6949 0.0921667
R6200 GND.n81 GND.n79 0.0921667
R6201 GND.n4770 GND.n4768 0.0921667
R6202 GND.n7492 GND.n7490 0.0921667
R6203 GND.n7617 GND.n7615 0.0921667
R6204 GND.n4605 GND.n4603 0.0920099
R6205 GND.n729 GND.n727 0.0894537
R6206 GND.n5863 GND.n5861 0.0894537
R6207 GND.n7236 GND.n7234 0.0894537
R6208 GND.n1542 GND.n1540 0.0891364
R6209 GND.n1014 GND.n1012 0.0891364
R6210 GND.n6514 GND.n6512 0.0891364
R6211 GND.n7525 GND.n7523 0.0891364
R6212 GND.n5225 GND.n5223 0.0891364
R6213 GND.n3490 GND.n3488 0.0891364
R6214 GND.n1122 GND.n1120 0.0891364
R6215 GND.n6776 GND.n6774 0.0891364
R6216 GND.n7091 GND.n7089 0.0891364
R6217 GND.n1992 GND.n1990 0.0891364
R6218 GND.n2315 GND.n2313 0.0891364
R6219 GND.n6930 GND.n6928 0.0891364
R6220 GND.n59 GND.n57 0.0891364
R6221 GND.n4901 GND.n4899 0.0891364
R6222 GND.n7463 GND.n7461 0.0891364
R6223 GND.n7588 GND.n7586 0.0891364
R6224 GND.n1360 GND.n1359 0.08745
R6225 GND.n2108 GND.n2107 0.08745
R6226 GND.n2431 GND.n2430 0.08745
R6227 GND.n2588 GND.n2587 0.08745
R6228 GND.n2752 GND.n2751 0.08745
R6229 GND.n2864 GND.n2863 0.08745
R6230 GND.n7684 GND.n7683 0.08745
R6231 GND.n3025 GND.n3024 0.08745
R6232 GND.n3135 GND.n3134 0.08745
R6233 GND.n5341 GND.n5340 0.08745
R6234 GND.n5017 GND.n5016 0.08745
R6235 GND.n3622 GND.n3621 0.08745
R6236 GND.n4039 GND.n4038 0.08745
R6237 GND.n3838 GND.n3837 0.08745
R6238 GND.n3242 GND.n3241 0.08745
R6239 GND.n1228 GND.n1227 0.08745
R6240 GND.n4039 GND.n3994 0.0868625
R6241 GND.n5341 GND.n5296 0.0868625
R6242 GND.n3025 GND.n2980 0.0868625
R6243 GND.n2588 GND.n2543 0.0868625
R6244 GND.n2108 GND.n2063 0.0868625
R6245 GND.n1407 GND.n1360 0.0868625
R6246 GND.n2431 GND.n2386 0.0868625
R6247 GND.n2752 GND.n2707 0.0868625
R6248 GND.n2864 GND.n2840 0.0868625
R6249 GND.n7684 GND.n7662 0.0868625
R6250 GND.n3135 GND.n3090 0.0868625
R6251 GND.n5017 GND.n4972 0.0868625
R6252 GND.n3622 GND.n3577 0.0868625
R6253 GND.n3838 GND.n3814 0.0868625
R6254 GND.n3242 GND.n3197 0.0868625
R6255 GND.n1228 GND.n1183 0.0868625
R6256 GND.n4227 GND.n4225 0.0853214
R6257 GND.n5623 GND.n5622 0.0845572
R6258 GND.n6527 GND.n650 0.0845572
R6259 GND.n7538 GND.n304 0.0845572
R6260 GND.n5239 GND.n5238 0.0845572
R6261 GND.n3504 GND.n3503 0.0845572
R6262 GND.n5441 GND.n5440 0.0845572
R6263 GND.n6806 GND.n6805 0.0845572
R6264 GND.n2006 GND.n2005 0.0845572
R6265 GND.n2329 GND.n2328 0.0845572
R6266 GND.n6960 GND.n6959 0.0845572
R6267 GND.n7736 GND.n7735 0.0845572
R6268 GND.n4915 GND.n4914 0.0845572
R6269 GND.n7476 GND.n508 0.0845572
R6270 GND.n7601 GND.n203 0.0845572
R6271 GND.n1552 GND.n1551 0.0845572
R6272 GND.n4532 GND.n4519 0.0838333
R6273 GND.n6495 GND 0.0824444
R6274 GND.n6292 GND 0.0824444
R6275 GND.n3079 GND.n1344 0.0813539
R6276 GND.n3180 GND.n1345 0.0813539
R6277 GND.n1438 GND 0.0775833
R6278 GND.n1022 GND 0.0775833
R6279 GND.n6530 GND 0.0775833
R6280 GND.n7541 GND 0.0775833
R6281 GND.n5078 GND 0.0775833
R6282 GND.n3289 GND 0.0775833
R6283 GND.n3444 GND 0.0775833
R6284 GND.n6784 GND 0.0775833
R6285 GND.n7107 GND 0.0775833
R6286 GND.n1844 GND 0.0775833
R6287 GND.n2179 GND 0.0775833
R6288 GND.n6938 GND 0.0775833
R6289 GND.n68 GND 0.0775833
R6290 GND.n4757 GND 0.0775833
R6291 GND.n7479 GND 0.0775833
R6292 GND.n7604 GND 0.0775833
R6293 GND.n6403 GND.n6378 0.0740087
R6294 GND.n6493 GND.n50 0.0740087
R6295 GND.n5435 GND.n1346 0.0735308
R6296 GND.n6404 GND.n6403 0.0732412
R6297 GND.n6494 GND.n6493 0.0732412
R6298 GND.n6405 GND.n6404 0.0727407
R6299 GND.n6494 GND.n6468 0.0727407
R6300 GND.n4420 GND.n4418 0.0727222
R6301 GND.n6468 GND.n676 0.0714246
R6302 GND.n7434 GND.n7433 0.0711855
R6303 GND.n6454 GND.n6453 0.0696598
R6304 GND.n7438 GND.n7437 0.0696598
R6305 GND.n6378 GND.n6377 0.0692593
R6306 GND.n7789 GND.n50 0.0692593
R6307 GND.n4434 GND.n4420 0.06925
R6308 GND.n1526 GND 0.0675455
R6309 GND GND.n5636 0.0675455
R6310 GND.n6502 GND 0.0675455
R6311 GND.n7513 GND 0.0675455
R6312 GND.n5213 GND 0.0675455
R6313 GND.n3478 GND 0.0675455
R6314 GND GND.n5454 0.0675455
R6315 GND GND.n6819 0.0675455
R6316 GND.n7079 GND 0.0675455
R6317 GND.n1980 GND 0.0675455
R6318 GND.n2303 GND 0.0675455
R6319 GND GND.n6973 0.0675455
R6320 GND GND.n7749 0.0675455
R6321 GND.n4889 GND 0.0675455
R6322 GND.n7451 GND 0.0675455
R6323 GND.n7576 GND 0.0675455
R6324 GND.n4110 GND.n4109 0.0672895
R6325 GND.n5409 GND.n5408 0.0672895
R6326 GND.n5408 GND.n5407 0.0672895
R6327 GND.n5407 GND.n1288 0.0672895
R6328 GND.n5434 GND.n5433 0.0672895
R6329 GND.n5433 GND.n5432 0.0672895
R6330 GND.n5432 GND.n5431 0.0672895
R6331 GND.n5431 GND.n5430 0.0672895
R6332 GND.n5430 GND.n5429 0.0672895
R6333 GND.n16 GND.n11 0.0659695
R6334 GND.n6338 GND.n6333 0.0659695
R6335 GND.n4642 GND.n4641 0.0653227
R6336 GND.n5436 GND.n1288 0.0648158
R6337 GND.n6218 GND.n6217 0.0643889
R6338 GND.n6217 GND.n6215 0.0643889
R6339 GND.n6215 GND.n6212 0.0643889
R6340 GND.n6212 GND.n6210 0.0643889
R6341 GND.n16 GND.n8 0.0643889
R6342 GND.n20 GND.n8 0.0643889
R6343 GND.n21 GND.n20 0.0643889
R6344 GND.n7768 GND.n7761 0.0643889
R6345 GND.n7774 GND.n7759 0.0643889
R6346 GND.n7774 GND.n7756 0.0643889
R6347 GND.n7778 GND.n7756 0.0643889
R6348 GND.n7779 GND.n7778 0.0643889
R6349 GND.n661 GND.n656 0.0643889
R6350 GND.n672 GND.n654 0.0643889
R6351 GND.n673 GND.n672 0.0643889
R6352 GND.n6338 GND.n6330 0.0643889
R6353 GND.n6342 GND.n6330 0.0643889
R6354 GND.n6343 GND.n6342 0.0643889
R6355 GND.n6308 GND.n6301 0.0643889
R6356 GND.n6314 GND.n6299 0.0643889
R6357 GND.n6314 GND.n6296 0.0643889
R6358 GND.n6318 GND.n6296 0.0643889
R6359 GND.n6319 GND.n6318 0.0643889
R6360 GND.n6276 GND.n6271 0.0643889
R6361 GND.n6287 GND.n6269 0.0643889
R6362 GND.n6288 GND.n6287 0.0643889
R6363 GND.n1371 GND.n1370 0.0636886
R6364 GND.n1372 GND.n1371 0.0636886
R6365 GND.n1374 GND.n1373 0.0636886
R6366 GND.n1373 GND.n1372 0.0636886
R6367 GND.n1349 GND.n1348 0.0636886
R6368 GND.n1348 GND.t524 0.0636886
R6369 GND.n2096 GND.n2095 0.0636886
R6370 GND.t126 GND.n2096 0.0636886
R6371 GND.n2098 GND.n2097 0.0636886
R6372 GND.n2097 GND.t126 0.0636886
R6373 GND.n2119 GND.n2118 0.0636886
R6374 GND.n2120 GND.n2119 0.0636886
R6375 GND.n2122 GND.n2121 0.0636886
R6376 GND.n2121 GND.n2120 0.0636886
R6377 GND.n2442 GND.n2441 0.0636886
R6378 GND.n2443 GND.n2442 0.0636886
R6379 GND.n2445 GND.n2444 0.0636886
R6380 GND.n2444 GND.n2443 0.0636886
R6381 GND.t132 GND.n2419 0.0636886
R6382 GND.n2419 GND.n2418 0.0636886
R6383 GND.n2420 GND.t132 0.0636886
R6384 GND.n2421 GND.n2420 0.0636886
R6385 GND.n2576 GND.n2575 0.0636886
R6386 GND.t125 GND.n2576 0.0636886
R6387 GND.n2578 GND.n2577 0.0636886
R6388 GND.n2577 GND.t125 0.0636886
R6389 GND.n2599 GND.n2598 0.0636886
R6390 GND.n2600 GND.n2599 0.0636886
R6391 GND.n2602 GND.n2601 0.0636886
R6392 GND.n2601 GND.n2600 0.0636886
R6393 GND.n2763 GND.n2762 0.0636886
R6394 GND.n2764 GND.n2763 0.0636886
R6395 GND.n2766 GND.n2765 0.0636886
R6396 GND.n2765 GND.n2764 0.0636886
R6397 GND.t104 GND.n2740 0.0636886
R6398 GND.n2740 GND.n2739 0.0636886
R6399 GND.n2741 GND.t104 0.0636886
R6400 GND.n2742 GND.n2741 0.0636886
R6401 GND.n2859 GND.n2858 0.0636886
R6402 GND.t103 GND.n2859 0.0636886
R6403 GND.n2861 GND.n2860 0.0636886
R6404 GND.n2860 GND.t103 0.0636886
R6405 GND.n2868 GND.n2867 0.0636886
R6406 GND.n2873 GND.n2872 0.0636886
R6407 GND.n7695 GND.n7694 0.0636886
R6408 GND.n7696 GND.n7695 0.0636886
R6409 GND.n7698 GND.n7697 0.0636886
R6410 GND.n7697 GND.n7696 0.0636886
R6411 GND.t833 GND.n7672 0.0636886
R6412 GND.n7672 GND.n7671 0.0636886
R6413 GND.n7673 GND.t833 0.0636886
R6414 GND.n7674 GND.n7673 0.0636886
R6415 GND.n3013 GND.n3012 0.0636886
R6416 GND.t12 GND.n3013 0.0636886
R6417 GND.n3014 GND.t12 0.0636886
R6418 GND.n3015 GND.n3014 0.0636886
R6419 GND.n3065 GND.n3064 0.0636886
R6420 GND.n3066 GND.n3065 0.0636886
R6421 GND.n3068 GND.n3067 0.0636886
R6422 GND.n3067 GND.n3066 0.0636886
R6423 GND.n3166 GND.n3165 0.0636886
R6424 GND.n3167 GND.n3166 0.0636886
R6425 GND.n3169 GND.n3168 0.0636886
R6426 GND.n3168 GND.n3167 0.0636886
R6427 GND.t11 GND.n3123 0.0636886
R6428 GND.n3123 GND.n3122 0.0636886
R6429 GND.n3124 GND.t11 0.0636886
R6430 GND.n3125 GND.n3124 0.0636886
R6431 GND.n1223 GND.n1222 0.0636886
R6432 GND.t128 GND.n1223 0.0636886
R6433 GND.n1224 GND.t128 0.0636886
R6434 GND.n1225 GND.n1224 0.0636886
R6435 GND.n1272 GND.n1271 0.0636886
R6436 GND.n1273 GND.n1272 0.0636886
R6437 GND.n1275 GND.n1274 0.0636886
R6438 GND.n1274 GND.n1273 0.0636886
R6439 GND.n3273 GND.n3272 0.0636886
R6440 GND.n3274 GND.n3273 0.0636886
R6441 GND.n3276 GND.n3275 0.0636886
R6442 GND.n3275 GND.n3274 0.0636886
R6443 GND.t527 GND.n3237 0.0636886
R6444 GND.n3237 GND.n3236 0.0636886
R6445 GND.n3238 GND.t527 0.0636886
R6446 GND.n3239 GND.n3238 0.0636886
R6447 GND.n5329 GND.n5328 0.0636886
R6448 GND.t509 GND.n5329 0.0636886
R6449 GND.n5331 GND.n5330 0.0636886
R6450 GND.n5330 GND.t509 0.0636886
R6451 GND.n5352 GND.n5351 0.0636886
R6452 GND.n5353 GND.n5352 0.0636886
R6453 GND.n5355 GND.n5354 0.0636886
R6454 GND.n5354 GND.n5353 0.0636886
R6455 GND.n5028 GND.n5027 0.0636886
R6456 GND.n5029 GND.n5028 0.0636886
R6457 GND.n5031 GND.n5030 0.0636886
R6458 GND.n5030 GND.n5029 0.0636886
R6459 GND.t107 GND.n5005 0.0636886
R6460 GND.n5005 GND.n5004 0.0636886
R6461 GND.n5006 GND.t107 0.0636886
R6462 GND.n5007 GND.n5006 0.0636886
R6463 GND.n3610 GND.n3609 0.0636886
R6464 GND.t127 GND.n3610 0.0636886
R6465 GND.n3611 GND.t127 0.0636886
R6466 GND.n3612 GND.n3611 0.0636886
R6467 GND.n3633 GND.n3632 0.0636886
R6468 GND.n3634 GND.n3633 0.0636886
R6469 GND.n3636 GND.n3635 0.0636886
R6470 GND.n3635 GND.n3634 0.0636886
R6471 GND.n4027 GND.n4026 0.0636886
R6472 GND.t736 GND.n4027 0.0636886
R6473 GND.n4028 GND.t736 0.0636886
R6474 GND.n4029 GND.n4028 0.0636886
R6475 GND.n4078 GND.n4077 0.0636886
R6476 GND.n4079 GND.n4078 0.0636886
R6477 GND.n4081 GND.n4080 0.0636886
R6478 GND.n4080 GND.n4079 0.0636886
R6479 GND.n1606 GND.n1605 0.0636886
R6480 GND.n1742 GND.n1606 0.0636886
R6481 GND.n1602 GND.n1601 0.0636886
R6482 GND.n1742 GND.n1602 0.0636886
R6483 GND.n1744 GND.n1743 0.0636886
R6484 GND.t186 GND.n1744 0.0636886
R6485 GND.n1616 GND.n1615 0.0636886
R6486 GND.n1742 GND.n1616 0.0636886
R6487 GND.n1611 GND.n1610 0.0636886
R6488 GND.n1742 GND.n1611 0.0636886
R6489 GND.n1746 GND.n1745 0.0636886
R6490 GND.t186 GND.n1746 0.0636886
R6491 GND.n1626 GND.n1625 0.0636886
R6492 GND.n1742 GND.n1626 0.0636886
R6493 GND.n1622 GND.n1621 0.0636886
R6494 GND.n1742 GND.n1622 0.0636886
R6495 GND.n1748 GND.n1747 0.0636886
R6496 GND.t186 GND.n1748 0.0636886
R6497 GND.n1636 GND.n1635 0.0636886
R6498 GND.n1742 GND.n1636 0.0636886
R6499 GND.n1632 GND.n1631 0.0636886
R6500 GND.n1742 GND.n1632 0.0636886
R6501 GND.n1750 GND.n1749 0.0636886
R6502 GND.t186 GND.n1750 0.0636886
R6503 GND.n1646 GND.n1645 0.0636886
R6504 GND.n1742 GND.n1646 0.0636886
R6505 GND.n1641 GND.n1640 0.0636886
R6506 GND.n1742 GND.n1641 0.0636886
R6507 GND.n1752 GND.n1751 0.0636886
R6508 GND.t186 GND.n1752 0.0636886
R6509 GND.n1661 GND.n1660 0.0636886
R6510 GND.n1742 GND.n1661 0.0636886
R6511 GND.n1653 GND.n1652 0.0636886
R6512 GND.n1742 GND.n1653 0.0636886
R6513 GND.n1754 GND.n1753 0.0636886
R6514 GND.t186 GND.n1754 0.0636886
R6515 GND.n1671 GND.n1670 0.0636886
R6516 GND.n1742 GND.n1671 0.0636886
R6517 GND.n1665 GND.n1664 0.0636886
R6518 GND.n1742 GND.n1665 0.0636886
R6519 GND.n1756 GND.n1755 0.0636886
R6520 GND.t186 GND.n1756 0.0636886
R6521 GND.n1681 GND.n1680 0.0636886
R6522 GND.n1742 GND.n1681 0.0636886
R6523 GND.n1675 GND.n1674 0.0636886
R6524 GND.n1742 GND.n1675 0.0636886
R6525 GND.n1758 GND.n1757 0.0636886
R6526 GND.t186 GND.n1758 0.0636886
R6527 GND.n1691 GND.n1690 0.0636886
R6528 GND.n1742 GND.n1691 0.0636886
R6529 GND.n1685 GND.n1684 0.0636886
R6530 GND.n1742 GND.n1685 0.0636886
R6531 GND.n1760 GND.n1759 0.0636886
R6532 GND.t186 GND.n1760 0.0636886
R6533 GND.n1701 GND.n1700 0.0636886
R6534 GND.n1742 GND.n1701 0.0636886
R6535 GND.n1695 GND.n1694 0.0636886
R6536 GND.n1742 GND.n1695 0.0636886
R6537 GND.n1762 GND.n1761 0.0636886
R6538 GND.t186 GND.n1762 0.0636886
R6539 GND.n1711 GND.n1710 0.0636886
R6540 GND.n1742 GND.n1711 0.0636886
R6541 GND.n1705 GND.n1704 0.0636886
R6542 GND.n1742 GND.n1705 0.0636886
R6543 GND.n1764 GND.n1763 0.0636886
R6544 GND.t186 GND.n1764 0.0636886
R6545 GND.n1721 GND.n1720 0.0636886
R6546 GND.n1742 GND.n1721 0.0636886
R6547 GND.n1716 GND.n1715 0.0636886
R6548 GND.n1742 GND.n1716 0.0636886
R6549 GND.n1766 GND.n1765 0.0636886
R6550 GND.t186 GND.n1766 0.0636886
R6551 GND.n1731 GND.n1730 0.0636886
R6552 GND.n1742 GND.n1731 0.0636886
R6553 GND.n1725 GND.n1724 0.0636886
R6554 GND.n1742 GND.n1725 0.0636886
R6555 GND.n1768 GND.n1767 0.0636886
R6556 GND.t186 GND.n1768 0.0636886
R6557 GND.n1741 GND.n1740 0.0636886
R6558 GND.n1742 GND.n1741 0.0636886
R6559 GND.n1736 GND.n1735 0.0636886
R6560 GND.n1742 GND.n1736 0.0636886
R6561 GND.n1770 GND.n1769 0.0636886
R6562 GND.t186 GND.n1770 0.0636886
R6563 GND.n3926 GND.n3925 0.0636886
R6564 GND.n3927 GND.n3926 0.0636886
R6565 GND.n3922 GND.n3921 0.0636886
R6566 GND.n3927 GND.n3922 0.0636886
R6567 GND.n3931 GND.n3930 0.0636886
R6568 GND.t503 GND.n3931 0.0636886
R6569 GND.n3916 GND.n3915 0.0636886
R6570 GND.n3927 GND.n3916 0.0636886
R6571 GND.n3910 GND.n3909 0.0636886
R6572 GND.n3927 GND.n3910 0.0636886
R6573 GND.n3929 GND.n3928 0.0636886
R6574 GND.t503 GND.n3929 0.0636886
R6575 GND.n3896 GND.n3895 0.0636886
R6576 GND.n3897 GND.n3896 0.0636886
R6577 GND.n3899 GND.n3898 0.0636886
R6578 GND.n3898 GND.n3897 0.0636886
R6579 GND.n3827 GND.t512 0.0636886
R6580 GND.n3828 GND.n3827 0.0636886
R6581 GND.t512 GND.n3826 0.0636886
R6582 GND.n3826 GND.n3825 0.0636886
R6583 GND.n3812 GND.n3811 0.0636886
R6584 GND.n3811 GND.t124 0.0636886
R6585 GND.n6347 GND.n6346 0.0636834
R6586 GND.n7794 GND.n24 0.0636834
R6587 GND.n6377 GND 0.0628765
R6588 GND GND.n7789 0.0628765
R6589 GND.n691 GND.n687 0.0610263
R6590 GND.n695 GND.n687 0.0610263
R6591 GND.n696 GND.n695 0.0610263
R6592 GND.n697 GND.n696 0.0610263
R6593 GND.n708 GND.n684 0.0610263
R6594 GND.n708 GND.n681 0.0610263
R6595 GND.n681 GND.n678 0.0610263
R6596 GND.n713 GND.n678 0.0610263
R6597 GND.n6242 GND.n6238 0.0610263
R6598 GND.n6246 GND.n6238 0.0610263
R6599 GND.n6247 GND.n6246 0.0610263
R6600 GND.n6248 GND.n6247 0.0610263
R6601 GND.n6259 GND.n6235 0.0610263
R6602 GND.n6259 GND.n6232 0.0610263
R6603 GND.n6232 GND.n6229 0.0610263
R6604 GND.n6264 GND.n6229 0.0610263
R6605 GND.n1552 GND 0.060284
R6606 GND.n5622 GND 0.060284
R6607 GND.n650 GND 0.060284
R6608 GND.n304 GND 0.060284
R6609 GND.n5239 GND 0.060284
R6610 GND.n3504 GND 0.060284
R6611 GND.n5440 GND 0.060284
R6612 GND.n6805 GND 0.060284
R6613 GND.n2486 GND 0.060284
R6614 GND.n2006 GND 0.060284
R6615 GND.n2329 GND 0.060284
R6616 GND.n6959 GND 0.060284
R6617 GND.n7735 GND 0.060284
R6618 GND.n4915 GND 0.060284
R6619 GND.n508 GND 0.060284
R6620 GND.n203 GND 0.060284
R6621 GND.n6405 GND.n550 0.0593951
R6622 GND.n4609 GND.n4608 0.0589677
R6623 GND.n3203 GND.n3202 0.0588369
R6624 GND.n2846 GND.n2845 0.0588369
R6625 GND.n1189 GND.n1188 0.0588369
R6626 GND.n1357 GND.n1356 0.0588344
R6627 GND.n2105 GND.n2104 0.0588344
R6628 GND.n2428 GND.n2427 0.0588344
R6629 GND.n2585 GND.n2584 0.0588344
R6630 GND.n2749 GND.n2748 0.0588344
R6631 GND.n7681 GND.n7680 0.0588344
R6632 GND.n3022 GND.n3021 0.0588344
R6633 GND.n3132 GND.n3131 0.0588344
R6634 GND.n5338 GND.n5337 0.0588344
R6635 GND.n5014 GND.n5013 0.0588344
R6636 GND.n3619 GND.n3618 0.0588344
R6637 GND.n4036 GND.n4035 0.0588344
R6638 GND.n3835 GND.n3834 0.0588344
R6639 GND.n1455 GND.n1454 0.0582982
R6640 GND.n1039 GND.n1038 0.0582982
R6641 GND.n6547 GND.n6546 0.0582982
R6642 GND.n7558 GND.n7557 0.0582982
R6643 GND.n5095 GND.n5094 0.0582982
R6644 GND.n3306 GND.n3305 0.0582982
R6645 GND.n3461 GND.n3460 0.0582982
R6646 GND.n6801 GND.n6800 0.0582982
R6647 GND.n7124 GND.n7123 0.0582982
R6648 GND.n1861 GND.n1860 0.0582982
R6649 GND.n2196 GND.n2192 0.0582982
R6650 GND.n6955 GND.n6954 0.0582982
R6651 GND.n85 GND.n84 0.0582982
R6652 GND.n4774 GND.n4773 0.0582982
R6653 GND.n7496 GND.n7495 0.0582982
R6654 GND.n7621 GND.n7620 0.0582982
R6655 GND.n4519 GND.n4517 0.0581389
R6656 GND.n6483 GND.n6482 0.0580634
R6657 GND.n6393 GND.n6392 0.0580634
R6658 GND.n23 GND.n6 0.0580441
R6659 GND.n7781 GND.n7754 0.0580441
R6660 GND.n669 GND.n668 0.0580441
R6661 GND.n675 GND.n652 0.0580441
R6662 GND.n6345 GND.n6328 0.0580441
R6663 GND.n6321 GND.n6294 0.0580441
R6664 GND.n6284 GND.n6283 0.0580441
R6665 GND.n6290 GND.n6267 0.0580441
R6666 GND.n6446 GND 0.058
R6667 GND.n6440 GND 0.058
R6668 GND.n6428 GND 0.058
R6669 GND.n543 GND 0.058
R6670 GND.n537 GND 0.058
R6671 GND.n525 GND 0.058
R6672 GND.n4205 GND.n4202 0.0570476
R6673 GND.n1532 GND.n1458 0.05675
R6674 GND.n5631 GND.n1008 0.05675
R6675 GND.n6508 GND.n651 0.05675
R6676 GND.n7519 GND.n305 0.05675
R6677 GND.n5219 GND.n5098 0.05675
R6678 GND.n3484 GND.n3333 0.05675
R6679 GND.n5449 GND.n1116 0.05675
R6680 GND.n6814 GND.n6770 0.05675
R6681 GND.n7085 GND.n7074 0.05675
R6682 GND.n1986 GND.n1864 0.05675
R6683 GND.n2309 GND.n2199 0.05675
R6684 GND.n6968 GND.n6924 0.05675
R6685 GND.n7742 GND.n7741 0.05675
R6686 GND.n4895 GND.n4777 0.05675
R6687 GND.n7457 GND.n509 0.05675
R6688 GND.n7582 GND.n204 0.05675
R6689 GND.n6486 GND.n6477 0.05675
R6690 GND.n6487 GND.n6475 0.05675
R6691 GND.n6396 GND.n6387 0.05675
R6692 GND.n6397 GND.n6385 0.05675
R6693 GND.n7770 GND.n7769 0.0567153
R6694 GND.n6310 GND.n6309 0.0567153
R6695 GND.n1018 GND.n1017 0.0560434
R6696 GND.n6518 GND.n6517 0.0560434
R6697 GND.n7529 GND.n7528 0.0560434
R6698 GND.n5229 GND.n5228 0.0560434
R6699 GND.n3494 GND.n3493 0.0560434
R6700 GND.n1126 GND.n1125 0.0560434
R6701 GND.n6780 GND.n6779 0.0560434
R6702 GND.n7095 GND.n7094 0.0560434
R6703 GND.n1996 GND.n1995 0.0560434
R6704 GND.n2319 GND.n2318 0.0560434
R6705 GND.n6934 GND.n6933 0.0560434
R6706 GND.n63 GND.n62 0.0560434
R6707 GND.n4905 GND.n4904 0.0560434
R6708 GND.n7467 GND.n7466 0.0560434
R6709 GND.n7592 GND.n7591 0.0560434
R6710 GND.n6453 GND.n6452 0.0558279
R6711 GND.n7437 GND.n549 0.0558279
R6712 GND.n6434 GND 0.0555
R6713 GND.n531 GND 0.0555
R6714 GND.n1548 GND.n1532 0.05425
R6715 GND.n5631 GND.n5630 0.05425
R6716 GND.n6524 GND.n6508 0.05425
R6717 GND.n7535 GND.n7519 0.05425
R6718 GND.n5235 GND.n5219 0.05425
R6719 GND.n3500 GND.n3484 0.05425
R6720 GND.n5449 GND.n5448 0.05425
R6721 GND.n6814 GND.n6813 0.05425
R6722 GND.n7101 GND.n7085 0.05425
R6723 GND.n2002 GND.n1986 0.05425
R6724 GND.n2325 GND.n2309 0.05425
R6725 GND.n6968 GND.n6967 0.05425
R6726 GND.n4911 GND.n4895 0.05425
R6727 GND.n7473 GND.n7457 0.05425
R6728 GND.n7598 GND.n7582 0.05425
R6729 GND.n4257 GND.n4256 0.0540714
R6730 GND.n1546 GND.n1545 0.0532741
R6731 GND.n64 GND.n63 0.0532741
R6732 GND.n4201 GND.n4198 0.0530794
R6733 GND.n701 GND.n700 0.052907
R6734 GND.n6252 GND.n6251 0.052907
R6735 GND.n1840 GND.n1839 0.0528195
R6736 GND.n1835 GND.n1834 0.0528195
R6737 GND.n1830 GND.n1829 0.0528195
R6738 GND.n1825 GND.n1824 0.0528195
R6739 GND.n1820 GND.n1819 0.0528195
R6740 GND.n1815 GND.n1814 0.0528195
R6741 GND.n1810 GND.n1809 0.0528195
R6742 GND.n1805 GND.n1804 0.0528195
R6743 GND.n1800 GND.n1799 0.0528195
R6744 GND.n1795 GND.n1794 0.0528195
R6745 GND.n1790 GND.n1789 0.0528195
R6746 GND.n1785 GND.n1784 0.0528195
R6747 GND.n1780 GND.n1779 0.0528195
R6748 GND.n1775 GND.n1772 0.0528195
R6749 GND.n3936 GND.n3933 0.0528195
R6750 GND.n1540 GND 0.0527727
R6751 GND.n1012 GND 0.0527727
R6752 GND.n6512 GND 0.0527727
R6753 GND.n7523 GND 0.0527727
R6754 GND.n5223 GND 0.0527727
R6755 GND.n3488 GND 0.0527727
R6756 GND.n1120 GND 0.0527727
R6757 GND.n6774 GND 0.0527727
R6758 GND.n7089 GND 0.0527727
R6759 GND.n1990 GND 0.0527727
R6760 GND.n2313 GND 0.0527727
R6761 GND.n6928 GND 0.0527727
R6762 GND.n57 GND 0.0527727
R6763 GND.n4899 GND 0.0527727
R6764 GND.n7461 GND 0.0527727
R6765 GND.n7586 GND 0.0527727
R6766 GND.n1564 GND.n1563 0.0525185
R6767 GND.n1565 GND.n1564 0.0525185
R6768 GND.n1558 GND.n1557 0.0525185
R6769 GND.n1559 GND.n1558 0.0525185
R6770 GND.n1570 GND.n1569 0.0525185
R6771 GND.n1571 GND.n1570 0.0525185
R6772 GND.n2024 GND.n2023 0.0525185
R6773 GND.n2025 GND.n2024 0.0525185
R6774 GND.n2018 GND.n2017 0.0525185
R6775 GND.n2019 GND.n2018 0.0525185
R6776 GND.n2033 GND.n2032 0.0525185
R6777 GND.n2034 GND.n2033 0.0525185
R6778 GND.n2029 GND.n2028 0.0525185
R6779 GND.n2031 GND.n2029 0.0525185
R6780 GND.n2015 GND.n2014 0.0525185
R6781 GND.n2016 GND.n2015 0.0525185
R6782 GND.n2343 GND.n2342 0.0525185
R6783 GND.n2344 GND.n2343 0.0525185
R6784 GND.n2337 GND.n2336 0.0525185
R6785 GND.n2338 GND.n2337 0.0525185
R6786 GND.n2370 GND.n2369 0.0525185
R6787 GND.n2371 GND.n2370 0.0525185
R6788 GND.n2334 GND.n2333 0.0525185
R6789 GND.n2335 GND.n2334 0.0525185
R6790 GND.n2367 GND.n2366 0.0525185
R6791 GND.n2368 GND.n2367 0.0525185
R6792 GND.n2504 GND.n2503 0.0525185
R6793 GND.n2505 GND.n2504 0.0525185
R6794 GND.n2498 GND.n2497 0.0525185
R6795 GND.n2499 GND.n2498 0.0525185
R6796 GND.n2513 GND.n2512 0.0525185
R6797 GND.n2514 GND.n2513 0.0525185
R6798 GND.n2509 GND.n2508 0.0525185
R6799 GND.n2511 GND.n2509 0.0525185
R6800 GND.n2495 GND.n2494 0.0525185
R6801 GND.n2496 GND.n2495 0.0525185
R6802 GND.n2664 GND.n2663 0.0525185
R6803 GND.n2665 GND.n2664 0.0525185
R6804 GND.n2658 GND.n2657 0.0525185
R6805 GND.n2659 GND.n2658 0.0525185
R6806 GND.n2691 GND.n2690 0.0525185
R6807 GND.n2692 GND.n2691 0.0525185
R6808 GND.n2655 GND.n2654 0.0525185
R6809 GND.n2656 GND.n2655 0.0525185
R6810 GND.n2688 GND.n2687 0.0525185
R6811 GND.n2689 GND.n2688 0.0525185
R6812 GND.n2920 GND.n2919 0.0525185
R6813 GND.n2921 GND.n2920 0.0525185
R6814 GND.n2914 GND.n2913 0.0525185
R6815 GND.n2915 GND.n2914 0.0525185
R6816 GND.n2931 GND.n2930 0.0525185
R6817 GND.n2932 GND.n2931 0.0525185
R6818 GND.n2928 GND.n2927 0.0525185
R6819 GND.n2929 GND.n2928 0.0525185
R6820 GND.n2911 GND.n2910 0.0525185
R6821 GND.n2912 GND.n2911 0.0525185
R6822 GND.n101 GND.n100 0.0525185
R6823 GND.n102 GND.n101 0.0525185
R6824 GND.n95 GND.n94 0.0525185
R6825 GND.n96 GND.n95 0.0525185
R6826 GND.n136 GND.n135 0.0525185
R6827 GND.n137 GND.n136 0.0525185
R6828 GND.n92 GND.n91 0.0525185
R6829 GND.n93 GND.n92 0.0525185
R6830 GND.n133 GND.n132 0.0525185
R6831 GND.n134 GND.n133 0.0525185
R6832 GND.n1306 GND.n1305 0.0525185
R6833 GND.n1307 GND.n1306 0.0525185
R6834 GND.n1300 GND.n1299 0.0525185
R6835 GND.n1301 GND.n1300 0.0525185
R6836 GND.n1315 GND.n1314 0.0525185
R6837 GND.n1316 GND.n1315 0.0525185
R6838 GND.n1312 GND.n1311 0.0525185
R6839 GND.n1313 GND.n1312 0.0525185
R6840 GND.n1297 GND.n1296 0.0525185
R6841 GND.n1298 GND.n1297 0.0525185
R6842 GND.n5581 GND.n5580 0.0525185
R6843 GND.n5582 GND.n5581 0.0525185
R6844 GND.n5575 GND.n5574 0.0525185
R6845 GND.n5576 GND.n5575 0.0525185
R6846 GND.n5590 GND.n5589 0.0525185
R6847 GND.n5591 GND.n5590 0.0525185
R6848 GND.n5572 GND.n5571 0.0525185
R6849 GND.n5573 GND.n5572 0.0525185
R6850 GND.n5587 GND.n5586 0.0525185
R6851 GND.n5588 GND.n5587 0.0525185
R6852 GND.n1142 GND.n1141 0.0525185
R6853 GND.n1143 GND.n1142 0.0525185
R6854 GND.n1136 GND.n1135 0.0525185
R6855 GND.n1137 GND.n1136 0.0525185
R6856 GND.n1153 GND.n1152 0.0525185
R6857 GND.n1154 GND.n1153 0.0525185
R6858 GND.n1150 GND.n1149 0.0525185
R6859 GND.n1151 GND.n1150 0.0525185
R6860 GND.n1133 GND.n1132 0.0525185
R6861 GND.n1134 GND.n1133 0.0525185
R6862 GND.n3518 GND.n3517 0.0525185
R6863 GND.n3519 GND.n3518 0.0525185
R6864 GND.n3512 GND.n3511 0.0525185
R6865 GND.n3513 GND.n3512 0.0525185
R6866 GND.n3527 GND.n3526 0.0525185
R6867 GND.n3528 GND.n3527 0.0525185
R6868 GND.n3509 GND.n3508 0.0525185
R6869 GND.n3510 GND.n3509 0.0525185
R6870 GND.n3524 GND.n3523 0.0525185
R6871 GND.n3525 GND.n3524 0.0525185
R6872 GND.n5257 GND.n5256 0.0525185
R6873 GND.n5258 GND.n5257 0.0525185
R6874 GND.n5251 GND.n5250 0.0525185
R6875 GND.n5252 GND.n5251 0.0525185
R6876 GND.n5266 GND.n5265 0.0525185
R6877 GND.n5267 GND.n5266 0.0525185
R6878 GND.n5262 GND.n5261 0.0525185
R6879 GND.n5264 GND.n5262 0.0525185
R6880 GND.n5248 GND.n5247 0.0525185
R6881 GND.n5249 GND.n5248 0.0525185
R6882 GND.n4930 GND.n4929 0.0525185
R6883 GND.n4931 GND.n4930 0.0525185
R6884 GND.n4924 GND.n4923 0.0525185
R6885 GND.n4925 GND.n4924 0.0525185
R6886 GND.n4957 GND.n4956 0.0525185
R6887 GND.n4958 GND.n4957 0.0525185
R6888 GND.n4921 GND.n4920 0.0525185
R6889 GND.n4922 GND.n4921 0.0525185
R6890 GND.n4954 GND.n4953 0.0525185
R6891 GND.n4955 GND.n4954 0.0525185
R6892 GND.n3688 GND.n3687 0.0525185
R6893 GND.n3689 GND.n3688 0.0525185
R6894 GND.n3682 GND.n3681 0.0525185
R6895 GND.n3683 GND.n3682 0.0525185
R6896 GND.n3715 GND.n3714 0.0525185
R6897 GND.n3716 GND.n3715 0.0525185
R6898 GND.n3679 GND.n3678 0.0525185
R6899 GND.n3680 GND.n3679 0.0525185
R6900 GND.n3712 GND.n3711 0.0525185
R6901 GND.n3713 GND.n3712 0.0525185
R6902 GND.n3955 GND.n3954 0.0525185
R6903 GND.n3956 GND.n3955 0.0525185
R6904 GND.n3949 GND.n3948 0.0525185
R6905 GND.n3950 GND.n3949 0.0525185
R6906 GND.n3964 GND.n3963 0.0525185
R6907 GND.n3965 GND.n3964 0.0525185
R6908 GND.n3961 GND.n3960 0.0525185
R6909 GND.n3962 GND.n3961 0.0525185
R6910 GND.n3946 GND.n3945 0.0525185
R6911 GND.n3947 GND.n3946 0.0525185
R6912 GND.n3735 GND.n3734 0.0525185
R6913 GND.n3736 GND.n3735 0.0525185
R6914 GND.n3768 GND.n3767 0.0525185
R6915 GND.n3769 GND.n3768 0.0525185
R6916 GND.n3744 GND.n3743 0.0525185
R6917 GND.n3745 GND.n3744 0.0525185
R6918 GND.n3738 GND.n3737 0.0525185
R6919 GND.n3739 GND.n3738 0.0525185
R6920 GND.n3771 GND.n3770 0.0525185
R6921 GND.n3772 GND.n3771 0.0525185
R6922 GND.n3841 GND.n3840 0.0525185
R6923 GND.n3842 GND.n3841 0.0525185
R6924 GND.n3892 GND.n3891 0.0525185
R6925 GND.n3891 GND.n3890 0.0525185
R6926 GND.n1839 GND.n1838 0.0523204
R6927 GND.n1834 GND.n1833 0.0523204
R6928 GND.n1829 GND.n1828 0.0523204
R6929 GND.n1824 GND.n1823 0.0523204
R6930 GND.n1819 GND.n1818 0.0523204
R6931 GND.n1814 GND.n1813 0.0523204
R6932 GND.n1809 GND.n1808 0.0523204
R6933 GND.n1804 GND.n1803 0.0523204
R6934 GND.n1799 GND.n1798 0.0523204
R6935 GND.n1794 GND.n1793 0.0523204
R6936 GND.n1789 GND.n1788 0.0523204
R6937 GND.n1784 GND.n1783 0.0523204
R6938 GND.n1779 GND.n1778 0.0523204
R6939 GND.n1772 GND.n1771 0.0523204
R6940 GND.n3933 GND.n3932 0.0523204
R6941 GND.n4096 GND.n4095 0.0523204
R6942 GND.n4099 GND.n4096 0.0523204
R6943 GND.n1531 GND.n1530 0.0516364
R6944 GND.n5633 GND.n5632 0.0516364
R6945 GND.n6507 GND.n6506 0.0516364
R6946 GND.n7518 GND.n7517 0.0516364
R6947 GND.n5218 GND.n5217 0.0516364
R6948 GND.n3483 GND.n3482 0.0516364
R6949 GND.n5451 GND.n5450 0.0516364
R6950 GND.n6816 GND.n6815 0.0516364
R6951 GND.n7084 GND.n7083 0.0516364
R6952 GND.n1985 GND.n1984 0.0516364
R6953 GND.n2308 GND.n2307 0.0516364
R6954 GND.n6970 GND.n6969 0.0516364
R6955 GND.n7744 GND.n7743 0.0516364
R6956 GND.n4894 GND.n4893 0.0516364
R6957 GND.n7456 GND.n7455 0.0516364
R6958 GND.n7581 GND.n7580 0.0516364
R6959 GND.n6376 GND.n676 0.0500734
R6960 GND.n5565 GND.n5564 0.0494583
R6961 GND.n6551 GND.n6550 0.0494583
R6962 GND.n7562 GND.n7561 0.0494583
R6963 GND.n5111 GND.n5110 0.0494583
R6964 GND.n3331 GND.n3330 0.0494583
R6965 GND.n3465 GND.n3464 0.0494583
R6966 GND.n6803 GND.n6766 0.0494583
R6967 GND.n7128 GND.n7127 0.0494583
R6968 GND.n1877 GND.n1876 0.0494583
R6969 GND.n2203 GND.n2202 0.0494583
R6970 GND.n6957 GND.n6920 0.0494583
R6971 GND.n6658 GND.n6657 0.0494583
R6972 GND.n4790 GND.n4789 0.0494583
R6973 GND.n7500 GND.n7499 0.0494583
R6974 GND.n7625 GND.n7624 0.0494583
R6975 GND.n1471 GND.n1459 0.0494583
R6976 GND.n7743 GND.n7740 0.0493636
R6977 GND GND.n690 0.0490201
R6978 GND GND.n6241 0.0490201
R6979 GND.n1456 GND.n1446 0.0486039
R6980 GND.n1040 GND.n1030 0.0486039
R6981 GND.n6548 GND.n6538 0.0486039
R6982 GND.n7559 GND.n7549 0.0486039
R6983 GND.n5096 GND.n5086 0.0486039
R6984 GND.n3307 GND.n3297 0.0486039
R6985 GND.n3462 GND.n3452 0.0486039
R6986 GND.n6802 GND.n6792 0.0486039
R6987 GND.n7125 GND.n7115 0.0486039
R6988 GND.n1862 GND.n1852 0.0486039
R6989 GND.n2197 GND.n2184 0.0486039
R6990 GND.n6956 GND.n6946 0.0486039
R6991 GND.n86 GND.n76 0.0486039
R6992 GND.n4775 GND.n4765 0.0486039
R6993 GND.n7497 GND.n7487 0.0486039
R6994 GND.n7622 GND.n7612 0.0486039
R6995 GND.n36 GND 0.0484167
R6996 GND GND.n25 0.0484167
R6997 GND.n1450 GND 0.0484167
R6998 GND.n1033 GND 0.0484167
R6999 GND.n6541 GND 0.0484167
R7000 GND.n7552 GND 0.0484167
R7001 GND.n5090 GND 0.0484167
R7002 GND.n3301 GND 0.0484167
R7003 GND.n3455 GND 0.0484167
R7004 GND.n6795 GND 0.0484167
R7005 GND.n7118 GND 0.0484167
R7006 GND.n1855 GND 0.0484167
R7007 GND.n2187 GND 0.0484167
R7008 GND.n6949 GND 0.0484167
R7009 GND.n79 GND 0.0484167
R7010 GND.n4768 GND 0.0484167
R7011 GND.n7490 GND 0.0484167
R7012 GND.n7615 GND 0.0484167
R7013 GND.n6360 GND 0.0484167
R7014 GND GND.n6349 0.0484167
R7015 GND.n1545 GND.n1544 0.0483725
R7016 GND.n1017 GND.n1016 0.0483725
R7017 GND.n6517 GND.n6516 0.0483725
R7018 GND.n7528 GND.n7527 0.0483725
R7019 GND.n5228 GND.n5227 0.0483725
R7020 GND.n3493 GND.n3492 0.0483725
R7021 GND.n1125 GND.n1124 0.0483725
R7022 GND.n6779 GND.n6778 0.0483725
R7023 GND.n7094 GND.n7093 0.0483725
R7024 GND.n1995 GND.n1994 0.0483725
R7025 GND.n2318 GND.n2317 0.0483725
R7026 GND.n6933 GND.n6932 0.0483725
R7027 GND.n63 GND.n61 0.0483725
R7028 GND.n4904 GND.n4903 0.0483725
R7029 GND.n7466 GND.n7465 0.0483725
R7030 GND.n7591 GND.n7590 0.0483725
R7031 GND.n4214 GND.n4212 0.048348
R7032 GND.n3190 GND.n1287 0.0483051
R7033 GND.n3083 GND.n3082 0.0483051
R7034 GND.n5427 GND.n5425 0.0483051
R7035 GND.n2170 GND.n2169 0.0483051
R7036 GND.n2479 GND.n2478 0.0483051
R7037 GND.n2644 GND.n2643 0.0483051
R7038 GND.n2813 GND.n2812 0.0483051
R7039 GND.n2965 GND.n2964 0.0483051
R7040 GND.n2973 GND.n2972 0.0483051
R7041 GND.n3184 GND.n3183 0.0483051
R7042 GND.n3564 GND.n3563 0.0483051
R7043 GND.n5405 GND.n5403 0.0483051
R7044 GND.n5074 GND.n5072 0.0483051
R7045 GND.n5413 GND.n5412 0.0483051
R7046 GND.n4089 GND.n4088 0.0483051
R7047 GND.n4107 GND.n4105 0.0483051
R7048 GND.n1446 GND.n1445 0.0464802
R7049 GND.n1030 GND.n1029 0.0464802
R7050 GND.n6538 GND.n6537 0.0464802
R7051 GND.n7549 GND.n7548 0.0464802
R7052 GND.n5086 GND.n5085 0.0464802
R7053 GND.n3297 GND.n3296 0.0464802
R7054 GND.n3452 GND.n3451 0.0464802
R7055 GND.n6792 GND.n6791 0.0464802
R7056 GND.n7115 GND.n7114 0.0464802
R7057 GND.n1852 GND.n1851 0.0464802
R7058 GND.n6946 GND.n6945 0.0464802
R7059 GND.n76 GND.n75 0.0464802
R7060 GND.n4765 GND.n4764 0.0464802
R7061 GND.n7487 GND.n7486 0.0464802
R7062 GND.n7612 GND.n7611 0.0464802
R7063 GND.n7782 GND 0.04425
R7064 GND.n6322 GND 0.04425
R7065 GND.n1499 GND.n1498 0.0425017
R7066 GND.n1498 GND.n1497 0.0425017
R7067 GND.n1885 GND.n1884 0.0425017
R7068 GND.n1886 GND.n1885 0.0425017
R7069 GND.n1916 GND.n1915 0.0425017
R7070 GND.n1915 GND.n1914 0.0425017
R7071 GND.n2210 GND.n2209 0.0425017
R7072 GND.n2211 GND.n2210 0.0425017
R7073 GND.n2239 GND.n2238 0.0425017
R7074 GND.n2238 GND.n2237 0.0425017
R7075 GND.n7141 GND.n7140 0.0425017
R7076 GND.n7142 GND.n7141 0.0425017
R7077 GND.n7165 GND.n7164 0.0425017
R7078 GND.n7164 GND.n7163 0.0425017
R7079 GND.n614 GND.n613 0.0425017
R7080 GND.n615 GND.n614 0.0425017
R7081 GND.n6999 GND.n6998 0.0425017
R7082 GND.n6998 GND.n6997 0.0425017
R7083 GND.n624 GND.n623 0.0425017
R7084 GND.n625 GND.n624 0.0425017
R7085 GND.n6845 GND.n6844 0.0425017
R7086 GND.n6844 GND.n6843 0.0425017
R7087 GND.n634 GND.n633 0.0425017
R7088 GND.n635 GND.n634 0.0425017
R7089 GND.n6691 GND.n6690 0.0425017
R7090 GND.n6690 GND.n6689 0.0425017
R7091 GND.n641 GND.n640 0.0425017
R7092 GND.n642 GND.n641 0.0425017
R7093 GND.n6621 GND.n6620 0.0425017
R7094 GND.n6620 GND.n6619 0.0425017
R7095 GND.n5553 GND.n5552 0.0425017
R7096 GND.n5554 GND.n5553 0.0425017
R7097 GND.n5518 GND.n5517 0.0425017
R7098 GND.n5517 GND.n5516 0.0425017
R7099 GND.n3431 GND.n3430 0.0425017
R7100 GND.n3432 GND.n3431 0.0425017
R7101 GND.n1084 GND.n1083 0.0425017
R7102 GND.n1083 GND.n1082 0.0425017
R7103 GND.n3337 GND.n3336 0.0425017
R7104 GND.n3338 GND.n3337 0.0425017
R7105 GND.n3392 GND.n3391 0.0425017
R7106 GND.n3391 GND.n3390 0.0425017
R7107 GND.n5118 GND.n5117 0.0425017
R7108 GND.n5119 GND.n5118 0.0425017
R7109 GND.n5152 GND.n5151 0.0425017
R7110 GND.n5151 GND.n5150 0.0425017
R7111 GND.n4797 GND.n4796 0.0425017
R7112 GND.n4798 GND.n4797 0.0425017
R7113 GND.n4828 GND.n4827 0.0425017
R7114 GND.n4827 GND.n4826 0.0425017
R7115 GND.n420 GND.n419 0.0425017
R7116 GND.n421 GND.n420 0.0425017
R7117 GND.n454 GND.n453 0.0425017
R7118 GND.n453 GND.n452 0.0425017
R7119 GND.n309 GND.n308 0.0425017
R7120 GND.n310 GND.n309 0.0425017
R7121 GND.n385 GND.n384 0.0425017
R7122 GND.n384 GND.n383 0.0425017
R7123 GND.n208 GND.n207 0.0425017
R7124 GND.n209 GND.n208 0.0425017
R7125 GND.n274 GND.n273 0.0425017
R7126 GND.n273 GND.n272 0.0425017
R7127 GND.n190 GND.n189 0.0425017
R7128 GND.n191 GND.n190 0.0425017
R7129 GND.n4004 GND.n4003 0.0415714
R7130 GND.n1404 GND.n1403 0.0415714
R7131 GND.n2073 GND.n2072 0.0415714
R7132 GND.n2395 GND.n2394 0.0415714
R7133 GND.n2553 GND.n2552 0.0415714
R7134 GND.n2716 GND.n2715 0.0415714
R7135 GND.n2821 GND.n2820 0.0415714
R7136 GND.n152 GND.n151 0.0415714
R7137 GND.n2990 GND.n2989 0.0415714
R7138 GND.n3099 GND.n3098 0.0415714
R7139 GND.n5306 GND.n5305 0.0415714
R7140 GND.n4981 GND.n4980 0.0415714
R7141 GND.n3587 GND.n3586 0.0415714
R7142 GND.n3787 GND.n3786 0.0415714
R7143 GND.n3213 GND.n3212 0.0415714
R7144 GND.n1200 GND.n1199 0.0415714
R7145 GND.n4006 GND.n4005 0.0406786
R7146 GND.n1408 GND.n1405 0.0406786
R7147 GND.n2075 GND.n2074 0.0406786
R7148 GND.n2397 GND.n2396 0.0406786
R7149 GND.n2555 GND.n2554 0.0406786
R7150 GND.n2718 GND.n2717 0.0406786
R7151 GND.n2839 GND.n2838 0.0406786
R7152 GND.n7660 GND.n7659 0.0406786
R7153 GND.n2992 GND.n2991 0.0406786
R7154 GND.n3101 GND.n3100 0.0406786
R7155 GND.n5308 GND.n5307 0.0406786
R7156 GND.n4983 GND.n4982 0.0406786
R7157 GND.n3589 GND.n3588 0.0406786
R7158 GND.n3806 GND.n3805 0.0406786
R7159 GND.n3215 GND.n3214 0.0406786
R7160 GND.n1202 GND.n1201 0.0406786
R7161 GND.n4734 GND.n4731 0.0390862
R7162 GND.n1286 GND 0.0386944
R7163 GND.n3081 GND 0.0386944
R7164 GND.n5426 GND 0.0386944
R7165 GND.n1841 GND 0.0386944
R7166 GND.n2176 GND 0.0386944
R7167 GND.n2485 GND 0.0386944
R7168 GND.n2650 GND 0.0386944
R7169 GND.n2963 GND 0.0386944
R7170 GND.n2971 GND 0.0386944
R7171 GND.n3182 GND 0.0386944
R7172 GND.n3562 GND 0.0386944
R7173 GND.n5404 GND 0.0386944
R7174 GND.n5073 GND 0.0386944
R7175 GND.n5411 GND 0.0386944
R7176 GND.n3937 GND 0.0386944
R7177 GND.n4106 GND 0.0386944
R7178 GND.n4209 GND.n4191 0.0381984
R7179 GND.n4608 GND.n4605 0.0367903
R7180 GND.n4754 GND.n4110 0.0363684
R7181 GND.n7788 GND.n24 0.0356562
R7182 GND.n6348 GND.n6347 0.0356562
R7183 GND.n714 GND 0.0353684
R7184 GND.n6265 GND 0.0353684
R7185 GND.n6206 GND.n6205 0.0352222
R7186 GND.n1112 GND.n1111 0.0345278
R7187 GND.n5546 GND.n5545 0.0345278
R7188 GND.n302 GND.n301 0.0345278
R7189 GND.n5103 GND.n5102 0.0345278
R7190 GND.n3312 GND.n3311 0.0345278
R7191 GND.n3420 GND.n3419 0.0345278
R7192 GND.n6763 GND.n6762 0.0345278
R7193 GND.n7071 GND.n7070 0.0345278
R7194 GND.n1869 GND.n1868 0.0345278
R7195 GND.n7134 GND.n7133 0.0345278
R7196 GND.n6917 GND.n6916 0.0345278
R7197 GND.n6649 GND.n6648 0.0345278
R7198 GND.n4782 GND.n4781 0.0345278
R7199 GND.n413 GND.n412 0.0345278
R7200 GND.n7629 GND.n7627 0.0345278
R7201 GND.n1464 GND.n1463 0.0345278
R7202 GND.n5566 GND.n5565 0.0337917
R7203 GND.n6550 GND.n6549 0.0337917
R7204 GND.n7561 GND.n7560 0.0337917
R7205 GND.n5110 GND.n5097 0.0337917
R7206 GND.n3332 GND.n3331 0.0337917
R7207 GND.n3464 GND.n3463 0.0337917
R7208 GND.n6804 GND.n6803 0.0337917
R7209 GND.n7127 GND.n7126 0.0337917
R7210 GND.n1876 GND.n1863 0.0337917
R7211 GND.n2202 GND.n2198 0.0337917
R7212 GND.n6958 GND.n6957 0.0337917
R7213 GND.n6657 GND.n87 0.0337917
R7214 GND.n4789 GND.n4776 0.0337917
R7215 GND.n7499 GND.n7498 0.0337917
R7216 GND.n7624 GND.n7623 0.0337917
R7217 GND.n1459 GND.n1457 0.0337917
R7218 GND.n6490 GND 0.033625
R7219 GND.n6400 GND 0.033625
R7220 GND.n1446 GND.n1442 0.0335935
R7221 GND.n1030 GND.n1026 0.0335935
R7222 GND.n6538 GND.n6534 0.0335935
R7223 GND.n7549 GND.n7545 0.0335935
R7224 GND.n5086 GND.n5082 0.0335935
R7225 GND.n3297 GND.n3293 0.0335935
R7226 GND.n3452 GND.n3448 0.0335935
R7227 GND.n6792 GND.n6788 0.0335935
R7228 GND.n7115 GND.n7111 0.0335935
R7229 GND.n1852 GND.n1848 0.0335935
R7230 GND.n2184 GND.n2183 0.0335935
R7231 GND.n6946 GND.n6942 0.0335935
R7232 GND.n76 GND.n72 0.0335935
R7233 GND.n4765 GND.n4761 0.0335935
R7234 GND.n7487 GND.n7483 0.0335935
R7235 GND.n7612 GND.n7608 0.0335935
R7236 GND GND.n6218 0.0324444
R7237 GND GND.n6208 0.0324444
R7238 GND.n668 GND 0.0324444
R7239 GND.n6283 GND 0.0324444
R7240 GND.n4245 GND.n4239 0.03175
R7241 GND.n7783 GND.n7782 0.03175
R7242 GND.n6323 GND.n6322 0.03175
R7243 GND.n5409 GND.n4754 0.0314211
R7244 GND.n6151 GND.n6149 0.0307632
R7245 GND.n6155 GND.n6151 0.0307632
R7246 GND.n6172 GND.n6168 0.0307632
R7247 GND.n6176 GND.n6172 0.0307632
R7248 GND.n6178 GND.n6176 0.0307632
R7249 GND.n6182 GND.n6178 0.0307632
R7250 GND.n6184 GND.n6182 0.0307632
R7251 GND.n6188 GND.n6184 0.0307632
R7252 GND.n6190 GND.n6188 0.0307632
R7253 GND.n5822 GND.n5821 0.0307632
R7254 GND.n5821 GND.n5819 0.0307632
R7255 GND.n5819 GND.n5815 0.0307632
R7256 GND.n5815 GND.n5813 0.0307632
R7257 GND.n5813 GND.n5809 0.0307632
R7258 GND.n5809 GND.n5807 0.0307632
R7259 GND.n5807 GND.n5803 0.0307632
R7260 GND.n5803 GND.n5799 0.0307632
R7261 GND.n5799 GND.n5797 0.0307632
R7262 GND.n5789 GND.n5785 0.0307632
R7263 GND.n5785 GND.n5783 0.0307632
R7264 GND.n5783 GND.n5779 0.0307632
R7265 GND.n5779 GND.n5777 0.0307632
R7266 GND.n5776 GND.n5775 0.0307632
R7267 GND.n5775 GND.n5773 0.0307632
R7268 GND.n5773 GND.n5769 0.0307632
R7269 GND.n5769 GND.n5767 0.0307632
R7270 GND.n5767 GND.n5763 0.0307632
R7271 GND.n5700 GND.n5696 0.0307632
R7272 GND.n5702 GND.n5700 0.0307632
R7273 GND.n5706 GND.n5702 0.0307632
R7274 GND.n5708 GND.n5706 0.0307632
R7275 GND.n5712 GND.n5708 0.0307632
R7276 GND.n5714 GND.n5712 0.0307632
R7277 GND.n5715 GND.n5714 0.0307632
R7278 GND.n5720 GND.n5718 0.0307632
R7279 GND.n5724 GND.n5720 0.0307632
R7280 GND.n5726 GND.n5724 0.0307632
R7281 GND.n5730 GND.n5726 0.0307632
R7282 GND.n5732 GND.n5730 0.0307632
R7283 GND.n691 GND 0.0307632
R7284 GND.n700 GND 0.0307632
R7285 GND.n6242 GND 0.0307632
R7286 GND.n6251 GND 0.0307632
R7287 GND.n2379 GND.n2378 0.0307537
R7288 GND.n2700 GND.n2699 0.0307537
R7289 GND.n145 GND.n144 0.0307537
R7290 GND.n4966 GND.n4965 0.0307537
R7291 GND.n3724 GND.n3723 0.0307537
R7292 GND.n3780 GND.n3779 0.0307537
R7293 GND.n715 GND.n714 0.0301053
R7294 GND.n6266 GND.n6265 0.0301053
R7295 GND GND.n4752 0.0300162
R7296 GND.n6208 GND.n6206 0.0296667
R7297 GND.n6205 GND.n6201 0.0296667
R7298 GND.n3939 GND.n3938 0.0296391
R7299 GND.n5241 GND.n5240 0.0296391
R7300 GND.n3554 GND.n3553 0.0296391
R7301 GND.n1147 GND.n1146 0.0296391
R7302 GND.n5617 GND.n5616 0.0296391
R7303 GND.n1290 GND.n1289 0.0296391
R7304 GND.n2925 GND.n2924 0.0296391
R7305 GND.n2488 GND.n2487 0.0296391
R7306 GND.n2008 GND.n2007 0.0296391
R7307 GND.n1589 GND.n1588 0.0296391
R7308 GND.n5745 GND.n5741 0.0294474
R7309 GND.n6491 GND.n6490 0.028625
R7310 GND.n6492 GND.n6491 0.028625
R7311 GND.n6401 GND.n6400 0.028625
R7312 GND.n6402 GND.n6401 0.028625
R7313 GND.n6221 GND.n6220 0.0284605
R7314 GND.n5797 GND.n5793 0.0282663
R7315 GND.n24 GND 0.0268889
R7316 GND.n6347 GND 0.0268889
R7317 GND.n5435 GND.n5434 0.0264737
R7318 GND.n5751 GND.n5732 0.0262926
R7319 GND.n3181 GND 0.024
R7320 GND.n3080 GND 0.024
R7321 GND.n6156 GND.n6155 0.0238553
R7322 GND.n5763 GND.n5761 0.0231974
R7323 GND.n5826 GND.n5825 0.0225395
R7324 GND.n5696 GND.n5694 0.0225395
R7325 GND.n5436 GND.n1344 0.0220137
R7326 GND.n5436 GND.n1345 0.0220137
R7327 GND.n6168 GND.n6166 0.0218816
R7328 GND.n6449 GND 0.02175
R7329 GND.n6443 GND 0.02175
R7330 GND.n6437 GND 0.02175
R7331 GND.n6431 GND 0.02175
R7332 GND.n6425 GND 0.02175
R7333 GND.n546 GND 0.02175
R7334 GND.n540 GND 0.02175
R7335 GND.n534 GND 0.02175
R7336 GND.n528 GND 0.02175
R7337 GND.n522 GND 0.02175
R7338 GND.n6224 GND.n6223 0.0212237
R7339 GND.n6455 GND.n6454 0.0209918
R7340 GND.n7439 GND.n7438 0.0209918
R7341 GND.n3999 GND.n3998 0.0208901
R7342 GND.n4002 GND.n3999 0.0208901
R7343 GND.n4012 GND.n4011 0.0208901
R7344 GND.n1399 GND.n1398 0.0208901
R7345 GND.n1402 GND.n1399 0.0208901
R7346 GND.n1414 GND.n1413 0.0208901
R7347 GND.n2068 GND.n2067 0.0208901
R7348 GND.n2071 GND.n2068 0.0208901
R7349 GND.n2081 GND.n2080 0.0208901
R7350 GND.n2390 GND.n2389 0.0208901
R7351 GND.n2393 GND.n2390 0.0208901
R7352 GND.n2403 GND.n2402 0.0208901
R7353 GND.n2548 GND.n2547 0.0208901
R7354 GND.n2551 GND.n2548 0.0208901
R7355 GND.n2561 GND.n2560 0.0208901
R7356 GND.n2711 GND.n2710 0.0208901
R7357 GND.n2714 GND.n2711 0.0208901
R7358 GND.n2724 GND.n2723 0.0208901
R7359 GND.n2824 GND.n2823 0.0208901
R7360 GND.n2827 GND.n2824 0.0208901
R7361 GND.n2832 GND.n2831 0.0208901
R7362 GND.n155 GND.n154 0.0208901
R7363 GND.n158 GND.n155 0.0208901
R7364 GND.n163 GND.n162 0.0208901
R7365 GND.n2985 GND.n2984 0.0208901
R7366 GND.n2988 GND.n2985 0.0208901
R7367 GND.n2998 GND.n2997 0.0208901
R7368 GND.n3094 GND.n3093 0.0208901
R7369 GND.n3097 GND.n3094 0.0208901
R7370 GND.n3107 GND.n3106 0.0208901
R7371 GND.n5301 GND.n5300 0.0208901
R7372 GND.n5304 GND.n5301 0.0208901
R7373 GND.n5314 GND.n5313 0.0208901
R7374 GND.n4976 GND.n4975 0.0208901
R7375 GND.n4979 GND.n4976 0.0208901
R7376 GND.n4989 GND.n4988 0.0208901
R7377 GND.n3582 GND.n3581 0.0208901
R7378 GND.n3585 GND.n3582 0.0208901
R7379 GND.n3595 GND.n3594 0.0208901
R7380 GND.n3790 GND.n3789 0.0208901
R7381 GND.n3793 GND.n3790 0.0208901
R7382 GND.n3798 GND.n3797 0.0208901
R7383 GND.n3208 GND.n3207 0.0208901
R7384 GND.n3211 GND.n3208 0.0208901
R7385 GND.n3221 GND.n3220 0.0208901
R7386 GND.n1195 GND.n1194 0.0208901
R7387 GND.n1198 GND.n1195 0.0208901
R7388 GND.n1208 GND.n1207 0.0208901
R7389 GND.n5792 GND.n5790 0.0205658
R7390 GND.n4637 GND.n4633 0.0202922
R7391 GND.n2846 GND.n2844 0.0200011
R7392 GND.n1357 GND.n1354 0.0200011
R7393 GND.n2105 GND.n2103 0.0200011
R7394 GND.n2428 GND.n2426 0.0200011
R7395 GND.n2585 GND.n2583 0.0200011
R7396 GND.n2749 GND.n2747 0.0200011
R7397 GND.n7681 GND.n7679 0.0200011
R7398 GND.n3022 GND.n3020 0.0200011
R7399 GND.n3132 GND.n3130 0.0200011
R7400 GND.n1189 GND.n1187 0.0200011
R7401 GND.n3203 GND.n3201 0.0200011
R7402 GND.n5338 GND.n5336 0.0200011
R7403 GND.n5014 GND.n5012 0.0200011
R7404 GND.n3619 GND.n3617 0.0200011
R7405 GND.n4036 GND.n4034 0.0200011
R7406 GND.n3835 GND.n3833 0.0200011
R7407 GND.n1523 GND 0.0198182
R7408 GND.n5637 GND 0.0198182
R7409 GND.n6499 GND 0.0198182
R7410 GND.n7510 GND 0.0198182
R7411 GND.n5210 GND 0.0198182
R7412 GND.n3475 GND 0.0198182
R7413 GND.n5455 GND 0.0198182
R7414 GND.n6820 GND 0.0198182
R7415 GND.n7076 GND 0.0198182
R7416 GND.n1977 GND 0.0198182
R7417 GND.n2300 GND 0.0198182
R7418 GND.n6974 GND 0.0198182
R7419 GND.n7750 GND 0.0198182
R7420 GND.n4886 GND 0.0198182
R7421 GND.n7448 GND 0.0198182
R7422 GND.n7573 GND 0.0198182
R7423 GND.n4633 GND.n4632 0.0197936
R7424 GND.n4013 GND.n4012 0.0195603
R7425 GND.n1415 GND.n1414 0.0195603
R7426 GND.n2082 GND.n2081 0.0195603
R7427 GND.n2404 GND.n2403 0.0195603
R7428 GND.n2562 GND.n2561 0.0195603
R7429 GND.n2725 GND.n2724 0.0195603
R7430 GND.n2836 GND.n2832 0.0195603
R7431 GND.n7657 GND.n163 0.0195603
R7432 GND.n2999 GND.n2998 0.0195603
R7433 GND.n3108 GND.n3107 0.0195603
R7434 GND.n5315 GND.n5314 0.0195603
R7435 GND.n4990 GND.n4989 0.0195603
R7436 GND.n3596 GND.n3595 0.0195603
R7437 GND.n3803 GND.n3798 0.0195603
R7438 GND.n3222 GND.n3221 0.0195603
R7439 GND.n1209 GND.n1208 0.0195603
R7440 GND.n1527 GND.n1526 0.0186818
R7441 GND.n5636 GND.n5634 0.0186818
R7442 GND.n6503 GND.n6502 0.0186818
R7443 GND.n7514 GND.n7513 0.0186818
R7444 GND.n5214 GND.n5213 0.0186818
R7445 GND.n3479 GND.n3478 0.0186818
R7446 GND.n5454 GND.n5452 0.0186818
R7447 GND.n6819 GND.n6817 0.0186818
R7448 GND.n7080 GND.n7079 0.0186818
R7449 GND.n1981 GND.n1980 0.0186818
R7450 GND.n2304 GND.n2303 0.0186818
R7451 GND.n6973 GND.n6971 0.0186818
R7452 GND.n7749 GND.n7745 0.0186818
R7453 GND.n4890 GND.n4889 0.0186818
R7454 GND.n7452 GND.n7451 0.0186818
R7455 GND.n7577 GND.n7576 0.0186818
R7456 GND.n5750 GND.n5746 0.0185921
R7457 GND.n4209 GND.n4201 0.0183571
R7458 GND.n44 GND 0.0182083
R7459 GND.n6368 GND 0.0182083
R7460 GND.n4627 GND.n4626 0.0179743
R7461 GND GND.n6209 0.0178611
R7462 GND.n1391 GND.n1390 0.0176904
R7463 GND.n2149 GND.n2148 0.0176904
R7464 GND.n2458 GND.n2457 0.0176904
R7465 GND.n2623 GND.n2622 0.0176904
R7466 GND.n2792 GND.n2791 0.0176904
R7467 GND.n2879 GND.n2878 0.0176904
R7468 GND.n7715 GND.n7714 0.0176904
R7469 GND.n3140 GND.n3139 0.0176904
R7470 GND.n3247 GND.n3246 0.0176904
R7471 GND.n5382 GND.n5381 0.0176904
R7472 GND.n5051 GND.n5050 0.0176904
R7473 GND.n3657 GND.n3656 0.0176904
R7474 GND.n3860 GND.n3859 0.0176904
R7475 GND.n6191 GND.n6190 0.0172763
R7476 GND.n4047 GND.n4046 0.0172687
R7477 GND.n1247 GND.n1246 0.0172687
R7478 GND.n3040 GND.n3039 0.0172687
R7479 GND GND.n35 0.0171667
R7480 GND.n1442 GND.n1440 0.0171667
R7481 GND.n1026 GND.n1024 0.0171667
R7482 GND.n6534 GND.n6532 0.0171667
R7483 GND.n7545 GND.n7543 0.0171667
R7484 GND.n5082 GND.n5080 0.0171667
R7485 GND.n3293 GND.n3291 0.0171667
R7486 GND.n3448 GND.n3446 0.0171667
R7487 GND.n6788 GND.n6786 0.0171667
R7488 GND.n7111 GND.n7109 0.0171667
R7489 GND.n1848 GND.n1846 0.0171667
R7490 GND.n2183 GND.n2181 0.0171667
R7491 GND.n6942 GND.n6940 0.0171667
R7492 GND.n72 GND.n70 0.0171667
R7493 GND.n4761 GND.n4759 0.0171667
R7494 GND.n7483 GND.n7481 0.0171667
R7495 GND.n7608 GND.n7606 0.0171667
R7496 GND GND.n6359 0.0171667
R7497 GND.n5740 GND.n5738 0.0171667
R7498 GND.n5738 GND.n5734 0.0171667
R7499 GND.n5734 GND.n5653 0.0171667
R7500 GND.n6142 GND.n6138 0.0171667
R7501 GND.n6144 GND.n6142 0.0171667
R7502 GND.n4205 GND.n4204 0.0167601
R7503 GND.n3991 GND.n3990 0.0166817
R7504 GND.n5293 GND.n5292 0.0166817
R7505 GND.n1181 GND.n1180 0.0166817
R7506 GND.n5620 GND.n5619 0.0166817
R7507 GND.n1342 GND.n1341 0.0166817
R7508 GND.n2959 GND.n2958 0.0166817
R7509 GND.n2540 GND.n2539 0.0166817
R7510 GND.n2060 GND.n2059 0.0166817
R7511 GND.n1593 GND.n1592 0.0166817
R7512 GND.n6161 GND.n6158 0.0166184
R7513 GND.n1543 GND.n1542 0.0164091
R7514 GND.n1015 GND.n1014 0.0164091
R7515 GND.n6515 GND.n6514 0.0164091
R7516 GND.n7526 GND.n7525 0.0164091
R7517 GND.n5226 GND.n5225 0.0164091
R7518 GND.n3491 GND.n3490 0.0164091
R7519 GND.n1123 GND.n1122 0.0164091
R7520 GND.n6777 GND.n6776 0.0164091
R7521 GND.n7092 GND.n7091 0.0164091
R7522 GND.n1993 GND.n1992 0.0164091
R7523 GND.n2316 GND.n2315 0.0164091
R7524 GND.n6931 GND.n6930 0.0164091
R7525 GND.n60 GND.n59 0.0164091
R7526 GND.n4902 GND.n4901 0.0164091
R7527 GND.n7464 GND.n7463 0.0164091
R7528 GND.n7589 GND.n7588 0.0164091
R7529 GND.n4254 GND.n4252 0.016125
R7530 GND.n5760 GND.n5756 0.0159605
R7531 GND.n5829 GND 0.0158101
R7532 GND.n6145 GND.n6144 0.0157174
R7533 GND.n4968 GND.n4967 0.0157059
R7534 GND.n6149 GND 0.0156316
R7535 GND.n5822 GND 0.0156316
R7536 GND GND.n5776 0.0156316
R7537 GND.n5718 GND 0.0156316
R7538 GND.n5756 GND.n5691 0.0153026
R7539 GND.n3991 GND.n3941 0.0152059
R7540 GND.n5293 GND.n5243 0.0152059
R7541 GND.n3558 GND.n3557 0.0152059
R7542 GND.n1181 GND.n1128 0.0152059
R7543 GND.n5620 GND.n5567 0.0152059
R7544 GND.n1342 GND.n1292 0.0152059
R7545 GND.n2959 GND.n2906 0.0152059
R7546 GND.n2540 GND.n2490 0.0152059
R7547 GND.n2060 GND.n2010 0.0152059
R7548 GND.n2383 GND.n2381 0.0152059
R7549 GND.n2704 GND.n2702 0.0152059
R7550 GND.n149 GND.n147 0.0152059
R7551 GND.n4969 GND.n4916 0.0152059
R7552 GND.n3728 GND.n3726 0.0152059
R7553 GND.n3784 GND.n3782 0.0152059
R7554 GND.n1380 GND.n1379 0.015169
R7555 GND.n1379 GND.t192 0.015169
R7556 GND.n1378 GND.n1377 0.015169
R7557 GND.t192 GND.n1378 0.015169
R7558 GND.n1376 GND.n1375 0.015169
R7559 GND.t192 GND.n1376 0.015169
R7560 GND.n1422 GND.n1421 0.015169
R7561 GND.n1421 GND.n1420 0.015169
R7562 GND.n1386 GND.n1385 0.015169
R7563 GND.n1385 GND.n1384 0.015169
R7564 GND.n2134 GND.n2133 0.015169
R7565 GND.n2135 GND.n2134 0.015169
R7566 GND.n2089 GND.n2088 0.015169
R7567 GND.n2092 GND.n2089 0.015169
R7568 GND.n2137 GND.n2136 0.015169
R7569 GND.n2136 GND.n2135 0.015169
R7570 GND.n2091 GND.n2090 0.015169
R7571 GND.n2092 GND.n2091 0.015169
R7572 GND.n2128 GND.n2127 0.015169
R7573 GND.n2127 GND.t613 0.015169
R7574 GND.n2126 GND.n2125 0.015169
R7575 GND.t613 GND.n2126 0.015169
R7576 GND.n2124 GND.n2123 0.015169
R7577 GND.t613 GND.n2124 0.015169
R7578 GND.n2451 GND.n2450 0.015169
R7579 GND.n2450 GND.t1078 0.015169
R7580 GND.n2449 GND.n2448 0.015169
R7581 GND.t1078 GND.n2449 0.015169
R7582 GND.n2447 GND.n2446 0.015169
R7583 GND.t1078 GND.n2447 0.015169
R7584 GND.n2145 GND.n2144 0.015169
R7585 GND.n2144 GND.n2143 0.015169
R7586 GND.n2411 GND.n2410 0.015169
R7587 GND.n2414 GND.n2411 0.015169
R7588 GND.n2413 GND.n2412 0.015169
R7589 GND.n2414 GND.n2413 0.015169
R7590 GND.n2142 GND.n2141 0.015169
R7591 GND.n2143 GND.n2142 0.015169
R7592 GND.n2614 GND.n2613 0.015169
R7593 GND.n2615 GND.n2614 0.015169
R7594 GND.n2569 GND.n2568 0.015169
R7595 GND.n2572 GND.n2569 0.015169
R7596 GND.n2617 GND.n2616 0.015169
R7597 GND.n2616 GND.n2615 0.015169
R7598 GND.n2571 GND.n2570 0.015169
R7599 GND.n2572 GND.n2571 0.015169
R7600 GND.n2608 GND.n2607 0.015169
R7601 GND.n2607 GND.t61 0.015169
R7602 GND.n2606 GND.n2605 0.015169
R7603 GND.t61 GND.n2606 0.015169
R7604 GND.n2604 GND.n2603 0.015169
R7605 GND.t61 GND.n2604 0.015169
R7606 GND.n2772 GND.n2771 0.015169
R7607 GND.n2771 GND.t792 0.015169
R7608 GND.n2770 GND.n2769 0.015169
R7609 GND.t792 GND.n2770 0.015169
R7610 GND.n2768 GND.n2767 0.015169
R7611 GND.t792 GND.n2768 0.015169
R7612 GND.n2778 GND.n2777 0.015169
R7613 GND.n2732 GND.n2731 0.015169
R7614 GND.n2735 GND.n2732 0.015169
R7615 GND.n2734 GND.n2733 0.015169
R7616 GND.n2735 GND.n2734 0.015169
R7617 GND.n2780 GND.n2779 0.015169
R7618 GND.n2779 GND.n2778 0.015169
R7619 GND.n2788 GND.n2787 0.015169
R7620 GND.n2787 GND.n2786 0.015169
R7621 GND.n2852 GND.n2851 0.015169
R7622 GND.n2855 GND.n2852 0.015169
R7623 GND.n2785 GND.n2784 0.015169
R7624 GND.n2786 GND.n2785 0.015169
R7625 GND.n2854 GND.n2853 0.015169
R7626 GND.n2855 GND.n2854 0.015169
R7627 GND.n1657 GND.n1656 0.015169
R7628 GND.n1656 GND.t545 0.015169
R7629 GND.n2889 GND.n2888 0.015169
R7630 GND.n2890 GND.n2889 0.015169
R7631 GND.n1650 GND.n1649 0.015169
R7632 GND.n1649 GND.t737 0.015169
R7633 GND.n7704 GND.n7703 0.015169
R7634 GND.n7703 GND.t210 0.015169
R7635 GND.n7702 GND.n7701 0.015169
R7636 GND.t210 GND.n7702 0.015169
R7637 GND.n7700 GND.n7699 0.015169
R7638 GND.t210 GND.n7700 0.015169
R7639 GND.n121 GND.n120 0.015169
R7640 GND.n120 GND.n118 0.015169
R7641 GND.n7664 GND.n7663 0.015169
R7642 GND.n7667 GND.n7664 0.015169
R7643 GND.n7666 GND.n7665 0.015169
R7644 GND.n7667 GND.n7666 0.015169
R7645 GND.n117 GND.n116 0.015169
R7646 GND.n118 GND.n117 0.015169
R7647 GND.n7711 GND.n7710 0.015169
R7648 GND.n7710 GND.n7709 0.015169
R7649 GND.n3006 GND.n3005 0.015169
R7650 GND.n3009 GND.n3006 0.015169
R7651 GND.n3028 GND.n3027 0.015169
R7652 GND.n3008 GND.n3007 0.015169
R7653 GND.n3009 GND.n3008 0.015169
R7654 GND.n3074 GND.n3073 0.015169
R7655 GND.n3073 GND.t421 0.015169
R7656 GND.n3072 GND.n3071 0.015169
R7657 GND.t421 GND.n3072 0.015169
R7658 GND.n3070 GND.n3069 0.015169
R7659 GND.t421 GND.n3070 0.015169
R7660 GND.n3175 GND.n3174 0.015169
R7661 GND.n3174 GND.t70 0.015169
R7662 GND.n3173 GND.n3172 0.015169
R7663 GND.t70 GND.n3173 0.015169
R7664 GND.n3171 GND.n3170 0.015169
R7665 GND.t70 GND.n3171 0.015169
R7666 GND.n3036 GND.n3035 0.015169
R7667 GND.n3035 GND.n3034 0.015169
R7668 GND.n3115 GND.n3114 0.015169
R7669 GND.n3118 GND.n3115 0.015169
R7670 GND.n3117 GND.n3116 0.015169
R7671 GND.n3118 GND.n3117 0.015169
R7672 GND.n3033 GND.n3032 0.015169
R7673 GND.n3034 GND.n3033 0.015169
R7674 GND.n1232 GND.n1231 0.015169
R7675 GND.n1233 GND.n1232 0.015169
R7676 GND.n1216 GND.n1215 0.015169
R7677 GND.n1219 GND.n1216 0.015169
R7678 GND.n1235 GND.n1234 0.015169
R7679 GND.n1234 GND.n1233 0.015169
R7680 GND.n1218 GND.n1217 0.015169
R7681 GND.n1219 GND.n1218 0.015169
R7682 GND.n1281 GND.n1280 0.015169
R7683 GND.n1280 GND.t405 0.015169
R7684 GND.n1279 GND.n1278 0.015169
R7685 GND.t405 GND.n1279 0.015169
R7686 GND.n1277 GND.n1276 0.015169
R7687 GND.t405 GND.n1277 0.015169
R7688 GND.n3282 GND.n3281 0.015169
R7689 GND.n3281 GND.t490 0.015169
R7690 GND.n3280 GND.n3279 0.015169
R7691 GND.t490 GND.n3280 0.015169
R7692 GND.n3278 GND.n3277 0.015169
R7693 GND.t490 GND.n3278 0.015169
R7694 GND.n1243 GND.n1242 0.015169
R7695 GND.n1242 GND.n1241 0.015169
R7696 GND.n3229 GND.n3228 0.015169
R7697 GND.n3232 GND.n3229 0.015169
R7698 GND.n3231 GND.n3230 0.015169
R7699 GND.n3232 GND.n3231 0.015169
R7700 GND.n1240 GND.n1239 0.015169
R7701 GND.n1241 GND.n1240 0.015169
R7702 GND.n5367 GND.n5366 0.015169
R7703 GND.n5368 GND.n5367 0.015169
R7704 GND.n5322 GND.n5321 0.015169
R7705 GND.n5325 GND.n5322 0.015169
R7706 GND.n5370 GND.n5369 0.015169
R7707 GND.n5369 GND.n5368 0.015169
R7708 GND.n5324 GND.n5323 0.015169
R7709 GND.n5325 GND.n5324 0.015169
R7710 GND.n5361 GND.n5360 0.015169
R7711 GND.n5360 GND.t63 0.015169
R7712 GND.n5359 GND.n5358 0.015169
R7713 GND.t63 GND.n5359 0.015169
R7714 GND.n5357 GND.n5356 0.015169
R7715 GND.t63 GND.n5357 0.015169
R7716 GND.n5037 GND.n5036 0.015169
R7717 GND.n5036 GND.t69 0.015169
R7718 GND.n5035 GND.n5034 0.015169
R7719 GND.t69 GND.n5035 0.015169
R7720 GND.n5033 GND.n5032 0.015169
R7721 GND.t69 GND.n5033 0.015169
R7722 GND.n5378 GND.n5377 0.015169
R7723 GND.n5377 GND.n5376 0.015169
R7724 GND.n4997 GND.n4996 0.015169
R7725 GND.n5000 GND.n4997 0.015169
R7726 GND.n4999 GND.n4998 0.015169
R7727 GND.n5000 GND.n4999 0.015169
R7728 GND.n5375 GND.n5374 0.015169
R7729 GND.n5376 GND.n5375 0.015169
R7730 GND.n5047 GND.n5046 0.015169
R7731 GND.n5046 GND.n5045 0.015169
R7732 GND.n3603 GND.n3602 0.015169
R7733 GND.n3606 GND.n3603 0.015169
R7734 GND.n3605 GND.n3604 0.015169
R7735 GND.n3606 GND.n3605 0.015169
R7736 GND.n5044 GND.n5043 0.015169
R7737 GND.n5045 GND.n5044 0.015169
R7738 GND.n3642 GND.n3641 0.015169
R7739 GND.n3641 GND.t546 0.015169
R7740 GND.n3640 GND.n3639 0.015169
R7741 GND.t546 GND.n3640 0.015169
R7742 GND.n3638 GND.n3637 0.015169
R7743 GND.t546 GND.n3638 0.015169
R7744 GND.n3653 GND.n3652 0.015169
R7745 GND.n3652 GND.n3650 0.015169
R7746 GND.n4020 GND.n4019 0.015169
R7747 GND.n4023 GND.n4020 0.015169
R7748 GND.n3649 GND.n3647 0.015169
R7749 GND.n3650 GND.n3649 0.015169
R7750 GND.n4022 GND.n4021 0.015169
R7751 GND.n4023 GND.n4022 0.015169
R7752 GND.n4070 GND.n4069 0.015169
R7753 GND.n4069 GND.t558 0.015169
R7754 GND.n4068 GND.n4067 0.015169
R7755 GND.t558 GND.n4068 0.015169
R7756 GND.n4066 GND.n4065 0.015169
R7757 GND.t558 GND.n4066 0.015169
R7758 GND.n4271 GND.n4270 0.015169
R7759 GND.n4272 GND.n4271 0.015169
R7760 GND.n4286 GND.n4285 0.015169
R7761 GND.n4287 GND.n4286 0.015169
R7762 GND.n4301 GND.n4300 0.015169
R7763 GND.n4302 GND.n4301 0.015169
R7764 GND.n4316 GND.n4315 0.015169
R7765 GND.n4317 GND.n4316 0.015169
R7766 GND.n4335 GND.n4334 0.015169
R7767 GND.n4336 GND.n4335 0.015169
R7768 GND.n4350 GND.n4349 0.015169
R7769 GND.n4351 GND.n4350 0.015169
R7770 GND.n4365 GND.n4364 0.015169
R7771 GND.n4366 GND.n4365 0.015169
R7772 GND.n4380 GND.n4379 0.015169
R7773 GND.n4381 GND.n4380 0.015169
R7774 GND.n4398 GND.n4397 0.015169
R7775 GND.n4399 GND.n4398 0.015169
R7776 GND.n4422 GND.n4421 0.015169
R7777 GND.n4423 GND.n4422 0.015169
R7778 GND.n4442 GND.n4441 0.015169
R7779 GND.n4443 GND.n4442 0.015169
R7780 GND.n4459 GND.n4458 0.015169
R7781 GND.n4460 GND.n4459 0.015169
R7782 GND.n4474 GND.n4473 0.015169
R7783 GND.n4475 GND.n4474 0.015169
R7784 GND.n4489 GND.n4488 0.015169
R7785 GND.n4490 GND.n4489 0.015169
R7786 GND.n4504 GND.n4503 0.015169
R7787 GND.n4505 GND.n4504 0.015169
R7788 GND.n4521 GND.n4520 0.015169
R7789 GND.n4522 GND.n4521 0.015169
R7790 GND.n4536 GND.n4535 0.015169
R7791 GND.n4537 GND.n4536 0.015169
R7792 GND.n4551 GND.n4550 0.015169
R7793 GND.n4552 GND.n4551 0.015169
R7794 GND.n4566 GND.n4565 0.015169
R7795 GND.n4567 GND.n4566 0.015169
R7796 GND.n4231 GND.n4230 0.015169
R7797 GND.n4582 GND.n4581 0.015169
R7798 GND.n4583 GND.n4582 0.015169
R7799 GND.n4220 GND.n4219 0.015169
R7800 GND.n4221 GND.n4220 0.015169
R7801 GND.n3881 GND.n3880 0.015169
R7802 GND.t1236 GND.n3881 0.015169
R7803 GND.n3882 GND.t1236 0.015169
R7804 GND.n3883 GND.n3882 0.015169
R7805 GND.n3879 GND.n3878 0.015169
R7806 GND.t1236 GND.n3879 0.015169
R7807 GND.n3856 GND.n3855 0.015169
R7808 GND.n4043 GND.n4042 0.015169
R7809 GND.n4042 GND.n4041 0.015169
R7810 GND.n3818 GND.n3817 0.015169
R7811 GND.n3821 GND.n3818 0.015169
R7812 GND.n3820 GND.n3819 0.015169
R7813 GND.n3821 GND.n3820 0.015169
R7814 GND.n3845 GND.n3844 0.015169
R7815 GND.n3844 GND.n3843 0.015169
R7816 GND.n3808 GND.n3807 0.015169
R7817 GND.n3809 GND.n3808 0.015169
R7818 GND.n4094 GND.n4093 0.014943
R7819 GND.n1840 GND.n1837 0.014943
R7820 GND.n1835 GND.n1832 0.014943
R7821 GND.n1830 GND.n1827 0.014943
R7822 GND.n1825 GND.n1822 0.014943
R7823 GND.n1820 GND.n1817 0.014943
R7824 GND.n1815 GND.n1812 0.014943
R7825 GND.n1810 GND.n1807 0.014943
R7826 GND.n1805 GND.n1802 0.014943
R7827 GND.n1800 GND.n1797 0.014943
R7828 GND.n1795 GND.n1792 0.014943
R7829 GND.n1790 GND.n1787 0.014943
R7830 GND.n1785 GND.n1782 0.014943
R7831 GND.n1780 GND.n1777 0.014943
R7832 GND.n1775 GND.n1774 0.014943
R7833 GND.n3936 GND.n3935 0.014943
R7834 GND.n6165 GND.n6161 0.0146447
R7835 GND.n5665 GND.n5663 0.0146077
R7836 GND.n1837 GND.n1836 0.0144432
R7837 GND.n1832 GND.n1831 0.0144432
R7838 GND.n1827 GND.n1826 0.0144432
R7839 GND.n1822 GND.n1821 0.0144432
R7840 GND.n1817 GND.n1816 0.0144432
R7841 GND.n1812 GND.n1811 0.0144432
R7842 GND.n1807 GND.n1806 0.0144432
R7843 GND.n1802 GND.n1801 0.0144432
R7844 GND.n1797 GND.n1796 0.0144432
R7845 GND.n1792 GND.n1791 0.0144432
R7846 GND.n1787 GND.n1786 0.0144432
R7847 GND.n1782 GND.n1781 0.0144432
R7848 GND.n1777 GND.n1776 0.0144432
R7849 GND.n1774 GND.n1773 0.0144432
R7850 GND.n3935 GND.n3934 0.0144432
R7851 GND.n4093 GND.n4092 0.0144432
R7852 GND.n4196 GND.n4194 0.0143889
R7853 GND.n1454 GND.n1453 0.0140417
R7854 GND.n1038 GND.n1037 0.0140417
R7855 GND.n6546 GND.n6545 0.0140417
R7856 GND.n7557 GND.n7556 0.0140417
R7857 GND.n5094 GND.n5093 0.0140417
R7858 GND.n3305 GND.n3304 0.0140417
R7859 GND.n3460 GND.n3459 0.0140417
R7860 GND.n6800 GND.n6799 0.0140417
R7861 GND.n7123 GND.n7122 0.0140417
R7862 GND.n1860 GND.n1859 0.0140417
R7863 GND.n2192 GND.n2191 0.0140417
R7864 GND.n6954 GND.n6953 0.0140417
R7865 GND.n84 GND.n83 0.0140417
R7866 GND.n4773 GND.n4772 0.0140417
R7867 GND.n7495 GND.n7494 0.0140417
R7868 GND.n7620 GND.n7619 0.0140417
R7869 GND.n6195 GND.n6191 0.0139868
R7870 GND.n4009 GND.n4008 0.0138596
R7871 GND.n1411 GND.n1410 0.0138596
R7872 GND.n2078 GND.n2077 0.0138596
R7873 GND.n2400 GND.n2399 0.0138596
R7874 GND.n2558 GND.n2557 0.0138596
R7875 GND.n2721 GND.n2720 0.0138596
R7876 GND.n2829 GND.n2828 0.0138596
R7877 GND.n160 GND.n159 0.0138596
R7878 GND.n2995 GND.n2994 0.0138596
R7879 GND.n3104 GND.n3103 0.0138596
R7880 GND.n5311 GND.n5310 0.0138596
R7881 GND.n4986 GND.n4985 0.0138596
R7882 GND.n3592 GND.n3591 0.0138596
R7883 GND.n3795 GND.n3794 0.0138596
R7884 GND.n3218 GND.n3217 0.0138596
R7885 GND.n1205 GND.n1204 0.0138596
R7886 GND.n733 GND.n729 0.012734
R7887 GND.n751 GND.n749 0.012734
R7888 GND.n755 GND.n751 0.012734
R7889 GND.n757 GND.n755 0.012734
R7890 GND.n761 GND.n757 0.012734
R7891 GND.n763 GND.n761 0.012734
R7892 GND.n767 GND.n763 0.012734
R7893 GND.n769 GND.n767 0.012734
R7894 GND.n770 GND.n769 0.012734
R7895 GND.n775 GND.n773 0.012734
R7896 GND.n779 GND.n775 0.012734
R7897 GND.n825 GND.n823 0.012734
R7898 GND.n823 GND.n819 0.012734
R7899 GND.n819 GND.n815 0.012734
R7900 GND.n815 GND.n813 0.012734
R7901 GND.n813 GND.n809 0.012734
R7902 GND.n809 GND.n807 0.012734
R7903 GND.n807 GND.n803 0.012734
R7904 GND.n803 GND.n801 0.012734
R7905 GND.n801 GND.n797 0.012734
R7906 GND.n797 GND.n795 0.012734
R7907 GND.n794 GND.n793 0.012734
R7908 GND.n793 GND.n791 0.012734
R7909 GND.n791 GND.n787 0.012734
R7910 GND.n847 GND.n843 0.012734
R7911 GND.n849 GND.n847 0.012734
R7912 GND.n853 GND.n849 0.012734
R7913 GND.n855 GND.n853 0.012734
R7914 GND.n859 GND.n855 0.012734
R7915 GND.n861 GND.n859 0.012734
R7916 GND.n865 GND.n861 0.012734
R7917 GND.n869 GND.n868 0.012734
R7918 GND.n874 GND.n872 0.012734
R7919 GND.n878 GND.n874 0.012734
R7920 GND.n918 GND.n916 0.012734
R7921 GND.n916 GND.n912 0.012734
R7922 GND.n912 GND.n908 0.012734
R7923 GND.n908 GND.n906 0.012734
R7924 GND.n906 GND.n902 0.012734
R7925 GND.n902 GND.n900 0.012734
R7926 GND.n900 GND.n896 0.012734
R7927 GND.n896 GND.n894 0.012734
R7928 GND.n894 GND.n890 0.012734
R7929 GND.n890 GND.n888 0.012734
R7930 GND.n887 GND.n886 0.012734
R7931 GND.n938 GND.n936 0.012734
R7932 GND.n942 GND.n938 0.012734
R7933 GND.n946 GND.n942 0.012734
R7934 GND.n948 GND.n946 0.012734
R7935 GND.n952 GND.n948 0.012734
R7936 GND.n954 GND.n952 0.012734
R7937 GND.n958 GND.n954 0.012734
R7938 GND.n960 GND.n958 0.012734
R7939 GND.n964 GND.n960 0.012734
R7940 GND.n966 GND.n964 0.012734
R7941 GND.n967 GND.n966 0.012734
R7942 GND.n972 GND.n970 0.012734
R7943 GND.n975 GND.n972 0.012734
R7944 GND.n977 GND.n975 0.012734
R7945 GND.n997 GND.n995 0.012734
R7946 GND.n992 GND.n991 0.012734
R7947 GND.n991 GND.n989 0.012734
R7948 GND.n989 GND.n985 0.012734
R7949 GND.n985 GND.n983 0.012734
R7950 GND.n5867 GND.n5863 0.012734
R7951 GND.n5869 GND.n5867 0.012734
R7952 GND.n5904 GND.n5900 0.012734
R7953 GND.n5900 GND.n5898 0.012734
R7954 GND.n5898 GND.n5894 0.012734
R7955 GND.n5894 GND.n5892 0.012734
R7956 GND.n5892 GND.n5888 0.012734
R7957 GND.n5888 GND.n5886 0.012734
R7958 GND.n5886 GND.n5882 0.012734
R7959 GND.n5882 GND.n5880 0.012734
R7960 GND.n5879 GND.n5878 0.012734
R7961 GND.n5878 GND.n5876 0.012734
R7962 GND.n5926 GND.n5922 0.012734
R7963 GND.n5930 GND.n5926 0.012734
R7964 GND.n5932 GND.n5930 0.012734
R7965 GND.n5936 GND.n5932 0.012734
R7966 GND.n5938 GND.n5936 0.012734
R7967 GND.n5942 GND.n5938 0.012734
R7968 GND.n5944 GND.n5942 0.012734
R7969 GND.n5948 GND.n5944 0.012734
R7970 GND.n5950 GND.n5948 0.012734
R7971 GND.n5951 GND.n5950 0.012734
R7972 GND.n5956 GND.n5954 0.012734
R7973 GND.n5960 GND.n5956 0.012734
R7974 GND.n5962 GND.n5960 0.012734
R7975 GND.n5993 GND.n5989 0.012734
R7976 GND.n5989 GND.n5985 0.012734
R7977 GND.n5985 GND.n5983 0.012734
R7978 GND.n5983 GND.n5979 0.012734
R7979 GND.n5979 GND.n5977 0.012734
R7980 GND.n5977 GND.n5973 0.012734
R7981 GND.n5973 GND.n5971 0.012734
R7982 GND.n5971 GND.n5849 0.012734
R7983 GND.n6130 GND.n6129 0.012734
R7984 GND.n6129 GND.n6127 0.012734
R7985 GND.n6007 GND.n6003 0.012734
R7986 GND.n6011 GND.n6007 0.012734
R7987 GND.n6013 GND.n6011 0.012734
R7988 GND.n6017 GND.n6013 0.012734
R7989 GND.n6019 GND.n6017 0.012734
R7990 GND.n6023 GND.n6019 0.012734
R7991 GND.n6025 GND.n6023 0.012734
R7992 GND.n6029 GND.n6025 0.012734
R7993 GND.n6031 GND.n6029 0.012734
R7994 GND.n6032 GND.n6031 0.012734
R7995 GND.n6037 GND.n6035 0.012734
R7996 GND.n6041 GND.n6037 0.012734
R7997 GND.n6051 GND.n6049 0.012734
R7998 GND.n6055 GND.n6051 0.012734
R7999 GND.n6059 GND.n6055 0.012734
R8000 GND.n6061 GND.n6059 0.012734
R8001 GND.n6065 GND.n6061 0.012734
R8002 GND.n6067 GND.n6065 0.012734
R8003 GND.n6071 GND.n6067 0.012734
R8004 GND.n6073 GND.n6071 0.012734
R8005 GND.n6077 GND.n6073 0.012734
R8006 GND.n6079 GND.n6077 0.012734
R8007 GND.n6080 GND.n6079 0.012734
R8008 GND.n6085 GND.n6083 0.012734
R8009 GND.n6088 GND.n6085 0.012734
R8010 GND.n6090 GND.n6088 0.012734
R8011 GND.n6110 GND.n6108 0.012734
R8012 GND.n6105 GND.n6104 0.012734
R8013 GND.n6104 GND.n6102 0.012734
R8014 GND.n6102 GND.n6098 0.012734
R8015 GND.n6098 GND.n6096 0.012734
R8016 GND.n7240 GND.n7236 0.012734
R8017 GND.n7242 GND.n7240 0.012734
R8018 GND.n7277 GND.n7273 0.012734
R8019 GND.n7273 GND.n7271 0.012734
R8020 GND.n7271 GND.n7267 0.012734
R8021 GND.n7267 GND.n7265 0.012734
R8022 GND.n7265 GND.n7261 0.012734
R8023 GND.n7261 GND.n7259 0.012734
R8024 GND.n7259 GND.n7255 0.012734
R8025 GND.n7255 GND.n7253 0.012734
R8026 GND.n7252 GND.n7251 0.012734
R8027 GND.n7251 GND.n7249 0.012734
R8028 GND.n7299 GND.n7295 0.012734
R8029 GND.n7303 GND.n7299 0.012734
R8030 GND.n7305 GND.n7303 0.012734
R8031 GND.n7309 GND.n7305 0.012734
R8032 GND.n7311 GND.n7309 0.012734
R8033 GND.n7315 GND.n7311 0.012734
R8034 GND.n7317 GND.n7315 0.012734
R8035 GND.n7321 GND.n7317 0.012734
R8036 GND.n7323 GND.n7321 0.012734
R8037 GND.n7324 GND.n7323 0.012734
R8038 GND.n7329 GND.n7327 0.012734
R8039 GND.n7333 GND.n7329 0.012734
R8040 GND.n7335 GND.n7333 0.012734
R8041 GND.n7366 GND.n7362 0.012734
R8042 GND.n7362 GND.n7358 0.012734
R8043 GND.n7358 GND.n7356 0.012734
R8044 GND.n7356 GND.n7352 0.012734
R8045 GND.n7352 GND.n7350 0.012734
R8046 GND.n7350 GND.n7346 0.012734
R8047 GND.n7346 GND.n7344 0.012734
R8048 GND.n7344 GND.n553 0.012734
R8049 GND.n7431 GND.n7430 0.012734
R8050 GND.n7430 GND.n7428 0.012734
R8051 GND.n7415 GND.n7413 0.012734
R8052 GND.n7413 GND.n7409 0.012734
R8053 GND.n7409 GND.n7405 0.012734
R8054 GND.n7405 GND.n7403 0.012734
R8055 GND.n7403 GND.n7399 0.012734
R8056 GND.n7399 GND.n7397 0.012734
R8057 GND.n7397 GND.n7393 0.012734
R8058 GND.n7393 GND.n7391 0.012734
R8059 GND.n7391 GND.n7387 0.012734
R8060 GND.n7387 GND.n7385 0.012734
R8061 GND.n7384 GND.n7383 0.012734
R8062 GND.n7383 GND.n7381 0.012734
R8063 GND.n603 GND.n599 0.012734
R8064 GND.n599 GND.n597 0.012734
R8065 GND.n597 GND.n593 0.012734
R8066 GND.n593 GND.n589 0.012734
R8067 GND.n589 GND.n587 0.012734
R8068 GND.n587 GND.n583 0.012734
R8069 GND.n583 GND.n581 0.012734
R8070 GND.n581 GND.n577 0.012734
R8071 GND.n577 GND.n575 0.012734
R8072 GND.n575 GND.n571 0.012734
R8073 GND.n571 GND.n569 0.012734
R8074 GND.n568 GND.n567 0.012734
R8075 GND.n567 GND.n565 0.012734
R8076 GND.n565 GND.n562 0.012734
R8077 GND.n7804 GND.n7803 0.012734
R8078 GND.n7809 GND.n7807 0.012734
R8079 GND.n7813 GND.n7809 0.012734
R8080 GND.n7815 GND.n7813 0.012734
R8081 GND.n7817 GND.n7815 0.012734
R8082 GND.n5746 GND.n5745 0.0126711
R8083 GND.n734 GND.n733 0.0126011
R8084 GND.n6132 GND.n6131 0.0126011
R8085 GND.n7433 GND.n7432 0.0126011
R8086 GND.n697 GND 0.0123421
R8087 GND.n6248 GND 0.0123421
R8088 GND.n866 GND.n865 0.0123351
R8089 GND.n886 GND.n884 0.0123351
R8090 GND.n6210 GND 0.0123056
R8091 GND GND.n6201 0.0123056
R8092 GND.n6202 GND 0.0123056
R8093 GND GND.n23 0.0123056
R8094 GND GND.n7781 0.0123056
R8095 GND GND.n675 0.0123056
R8096 GND GND.n6345 0.0123056
R8097 GND GND.n6321 0.0123056
R8098 GND GND.n6290 0.0123056
R8099 GND.n2844 GND.n2843 0.0120741
R8100 GND.n1354 GND.n1353 0.0120741
R8101 GND.n2103 GND.n2102 0.0120741
R8102 GND.n2426 GND.n2425 0.0120741
R8103 GND.n2583 GND.n2582 0.0120741
R8104 GND.n2747 GND.n2746 0.0120741
R8105 GND.n7679 GND.n7678 0.0120741
R8106 GND.n3020 GND.n3019 0.0120741
R8107 GND.n3130 GND.n3129 0.0120741
R8108 GND.n1187 GND.n1186 0.0120741
R8109 GND.n3201 GND.n3200 0.0120741
R8110 GND.n5336 GND.n5335 0.0120741
R8111 GND.n5012 GND.n5011 0.0120741
R8112 GND.n3617 GND.n3616 0.0120741
R8113 GND.n4034 GND.n4033 0.0120741
R8114 GND.n3833 GND.n3832 0.0120741
R8115 GND.n5876 GND.n5872 0.0120691
R8116 GND.n7249 GND.n7245 0.0120691
R8117 GND.n6138 GND.n6136 0.0117319
R8118 GND GND.n7768 0.0116111
R8119 GND.n656 GND 0.0116111
R8120 GND GND.n6308 0.0116111
R8121 GND.n6271 GND 0.0116111
R8122 GND.n780 GND.n779 0.0115372
R8123 GND.n5562 GND.n5561 0.0112143
R8124 GND.n6555 GND.n6553 0.0112143
R8125 GND.n319 GND.n317 0.0112143
R8126 GND.n5201 GND.n5126 0.0112143
R8127 GND.n3328 GND.n3327 0.0112143
R8128 GND.n3440 GND.n3439 0.0112143
R8129 GND.n6908 GND.n6906 0.0112143
R8130 GND.n7221 GND.n7149 0.0112143
R8131 GND.n1968 GND.n1893 0.0112143
R8132 GND.n2291 GND.n2218 0.0112143
R8133 GND.n7062 GND.n7060 0.0112143
R8134 GND.n6754 GND.n6752 0.0112143
R8135 GND.n4877 GND.n4805 0.0112143
R8136 GND.n506 GND.n428 0.0112143
R8137 GND.n217 GND.n215 0.0112143
R8138 GND.n1515 GND.n1476 0.0112143
R8139 GND.n2843 GND 0.0111481
R8140 GND.n1353 GND 0.0111481
R8141 GND.n2102 GND 0.0111481
R8142 GND.n2425 GND 0.0111481
R8143 GND.n2582 GND 0.0111481
R8144 GND.n2746 GND 0.0111481
R8145 GND.n7678 GND 0.0111481
R8146 GND.n3019 GND 0.0111481
R8147 GND.n3129 GND 0.0111481
R8148 GND.n1186 GND 0.0111481
R8149 GND.n3200 GND 0.0111481
R8150 GND.n5335 GND 0.0111481
R8151 GND.n5011 GND 0.0111481
R8152 GND.n3616 GND 0.0111481
R8153 GND.n4033 GND 0.0111481
R8154 GND.n3832 GND 0.0111481
R8155 GND GND.n713 0.0110263
R8156 GND GND.n6264 0.0110263
R8157 GND.n4261 GND.n4259 0.0109167
R8158 GND.n843 GND.n839 0.0107394
R8159 GND.n919 GND.n918 0.0107394
R8160 GND.n6091 GND.n6090 0.0107394
R8161 GND.n562 GND.n3 0.0107394
R8162 GND.n5910 GND.n5869 0.0107015
R8163 GND.n7283 GND.n7242 0.0107015
R8164 GND.n5790 GND.n5789 0.0106974
R8165 GND.n6042 GND.n6041 0.0104355
R8166 GND.n7381 GND.n7377 0.0104355
R8167 GND.n4333 GND.n4332 0.0102222
R8168 GND.n978 GND.n977 0.0102074
R8169 GND.n5994 GND.n5993 0.0102074
R8170 GND.n6003 GND.n6001 0.0102074
R8171 GND.n7367 GND.n7366 0.0102074
R8172 GND.n7416 GND.n7415 0.0102074
R8173 GND.n4122 GND.n4121 0.0101468
R8174 GND.n4123 GND.n4122 0.0101468
R8175 GND.n4181 GND.n4180 0.0101468
R8176 GND.n4182 GND.n4181 0.0101468
R8177 GND.n4176 GND.n4175 0.0101468
R8178 GND.n4182 GND.n4176 0.0101468
R8179 GND.n4171 GND.n4170 0.0101468
R8180 GND.n4182 GND.n4171 0.0101468
R8181 GND.n4168 GND.n4167 0.0101468
R8182 GND.n4182 GND.n4168 0.0101468
R8183 GND.n4120 GND.n4119 0.0101468
R8184 GND.n4123 GND.n4120 0.0101468
R8185 GND.n4163 GND.n4162 0.0101468
R8186 GND.n4182 GND.n4163 0.0101468
R8187 GND.n4158 GND.n4157 0.0101468
R8188 GND.n4182 GND.n4158 0.0101468
R8189 GND.n4154 GND.n4153 0.0101468
R8190 GND.n4182 GND.n4154 0.0101468
R8191 GND.n4150 GND.n4149 0.0101468
R8192 GND.n4182 GND.n4150 0.0101468
R8193 GND.n4147 GND.n4146 0.0101468
R8194 GND.n4182 GND.n4147 0.0101468
R8195 GND.n4118 GND.n4117 0.0101468
R8196 GND.n4123 GND.n4118 0.0101468
R8197 GND.n4141 GND.n4140 0.0101468
R8198 GND.n4182 GND.n4141 0.0101468
R8199 GND.n4135 GND.n4134 0.0101468
R8200 GND.n4182 GND.n4135 0.0101468
R8201 GND.n4116 GND.n4115 0.0101468
R8202 GND.n4123 GND.n4116 0.0101468
R8203 GND.n4131 GND.n4130 0.0101468
R8204 GND.n4182 GND.n4131 0.0101468
R8205 GND.n4125 GND.n4124 0.0101468
R8206 GND.n4182 GND.n4125 0.0101468
R8207 GND.n6224 GND.n6195 0.0100395
R8208 GND.n5662 GND.n5658 0.0100149
R8209 GND GND.n6489 0.009875
R8210 GND GND.n6399 0.009875
R8211 GND.n740 GND.n736 0.00967553
R8212 GND.n4261 GND.n4260 0.00959091
R8213 GND.n701 GND.n684 0.00950855
R8214 GND.n6252 GND.n6235 0.00950855
R8215 GND.n5672 GND.n5670 0.00941473
R8216 GND.n5676 GND.n5672 0.00941473
R8217 GND.n5680 GND.n5676 0.00941473
R8218 GND.n5682 GND.n5680 0.00941473
R8219 GND.n5846 GND.n5842 0.00941473
R8220 GND.n5842 GND.n5840 0.00941473
R8221 GND.n5840 GND.n5836 0.00941473
R8222 GND.n5836 GND.n5834 0.00941473
R8223 GND.n929 GND.n720 0.00940957
R8224 GND.n6166 GND.n6165 0.00938158
R8225 GND.n5915 GND.n5857 0.00914362
R8226 GND.n7288 GND.n7231 0.00914362
R8227 GND.n7769 GND.n7759 0.00906279
R8228 GND.n6309 GND.n6299 0.00906279
R8229 GND.n4646 GND.n4645 0.00904142
R8230 GND.n4723 GND.n4720 0.00898517
R8231 GND.n4685 GND.n4683 0.00898517
R8232 GND.n4703 GND.n4685 0.00898517
R8233 GND.n4665 GND.n4664 0.00898517
R8234 GND.n4664 GND.n4662 0.00898517
R8235 GND.n4649 GND.n4648 0.00898517
R8236 GND.n4648 GND.n4646 0.00898517
R8237 GND.n4723 GND.n4722 0.00897458
R8238 GND.n4734 GND.n4733 0.00896398
R8239 GND.n4705 GND.n4703 0.00896398
R8240 GND.n4709 GND.n4705 0.00896398
R8241 GND.n4711 GND.n4709 0.00896398
R8242 GND.n4712 GND.n4711 0.00896398
R8243 GND.n4677 GND.n4676 0.00896398
R8244 GND.n4657 GND.n4654 0.00896398
R8245 GND.n4657 GND.n4656 0.00896398
R8246 GND.n4665 GND.n4661 0.0089428
R8247 GND.n998 GND.n997 0.00887766
R8248 GND.n5963 GND.n5962 0.00887766
R8249 GND.n6127 GND.n6123 0.00887766
R8250 GND.n7336 GND.n7335 0.00887766
R8251 GND.n7428 GND.n7424 0.00887766
R8252 GND.n5828 GND.n5826 0.00872368
R8253 GND.n5694 GND.n5691 0.00872368
R8254 GND.n831 GND.n782 0.0086117
R8255 GND.n4617 GND.n4609 0.00856452
R8256 GND.n787 GND.n785 0.00834574
R8257 GND.n879 GND.n878 0.00834574
R8258 GND.n6111 GND.n6110 0.00834574
R8259 GND.n7803 GND.n7801 0.00834574
R8260 GND.n4676 GND 0.00822246
R8261 GND GND.n6219 0.00806579
R8262 GND.n5761 GND.n5760 0.00806579
R8263 GND.n4011 GND.n4009 0.00783909
R8264 GND.n1413 GND.n1411 0.00783909
R8265 GND.n2080 GND.n2078 0.00783909
R8266 GND.n2402 GND.n2400 0.00783909
R8267 GND.n2560 GND.n2558 0.00783909
R8268 GND.n2723 GND.n2721 0.00783909
R8269 GND.n2831 GND.n2829 0.00783909
R8270 GND.n162 GND.n160 0.00783909
R8271 GND.n2997 GND.n2995 0.00783909
R8272 GND.n3106 GND.n3104 0.00783909
R8273 GND.n5313 GND.n5311 0.00783909
R8274 GND.n4988 GND.n4986 0.00783909
R8275 GND.n3594 GND.n3592 0.00783909
R8276 GND.n3797 GND.n3795 0.00783909
R8277 GND.n3220 GND.n3218 0.00783909
R8278 GND.n1207 GND.n1205 0.00783909
R8279 GND.n4672 GND.n4670 0.00781992
R8280 GND.n838 GND.n836 0.00781383
R8281 GND.n924 GND.n923 0.00781383
R8282 GND.n4214 GND.n4213 0.00779984
R8283 GND.n21 GND.n6 0.00775202
R8284 GND.n7779 GND.n7754 0.00775202
R8285 GND.n669 GND.n654 0.00775202
R8286 GND.n673 GND.n652 0.00775202
R8287 GND.n6343 GND.n6328 0.00775202
R8288 GND.n6319 GND.n6294 0.00775202
R8289 GND.n6284 GND.n6269 0.00775202
R8290 GND.n6288 GND.n6267 0.00775202
R8291 GND.n4615 GND.n4614 0.00769258
R8292 GND.n4603 GND.n4602 0.00769258
R8293 GND.n826 GND.n825 0.00754787
R8294 GND.n4745 GND.n4744 0.00744444
R8295 GND.n4189 GND.n4112 0.00744444
R8296 GND.n6158 GND.n6156 0.00740789
R8297 GND.n3998 GND.n3997 0.00739975
R8298 GND.n1398 GND.n1397 0.00739975
R8299 GND.n2067 GND.n2066 0.00739975
R8300 GND.n2389 GND.n2388 0.00739975
R8301 GND.n2547 GND.n2546 0.00739975
R8302 GND.n2710 GND.n2709 0.00739975
R8303 GND.n2823 GND.n2822 0.00739975
R8304 GND.n154 GND.n153 0.00739975
R8305 GND.n2984 GND.n2983 0.00739975
R8306 GND.n3093 GND.n3092 0.00739975
R8307 GND.n5300 GND.n5299 0.00739975
R8308 GND.n4975 GND.n4974 0.00739975
R8309 GND.n3581 GND.n3580 0.00739975
R8310 GND.n3789 GND.n3788 0.00739975
R8311 GND.n3207 GND.n3206 0.00739975
R8312 GND.n1194 GND.n1193 0.00739975
R8313 GND.n4201 GND.n4200 0.00738379
R8314 GND.n5909 GND.n5905 0.00728191
R8315 GND.n5997 GND.n5996 0.00728191
R8316 GND.n6120 GND.n5855 0.00728191
R8317 GND.n7282 GND.n7278 0.00728191
R8318 GND.n7370 GND.n7369 0.00728191
R8319 GND.n7421 GND.n7420 0.00728191
R8320 GND.n4235 GND.n4232 0.00719643
R8321 GND.n5829 GND.n5828 0.00707895
R8322 GND.n5922 GND.n5920 0.00701596
R8323 GND.n6045 GND.n6044 0.00701596
R8324 GND.n7295 GND.n7293 0.00701596
R8325 GND.n606 GND.n604 0.00701596
R8326 GND.n4332 GND.n4330 0.00675
R8327 GND.n745 GND.n744 0.00675
R8328 GND.n936 GND.n932 0.00675
R8329 GND.n4259 GND.n4258 0.0066794
R8330 GND.n4235 GND.n4234 0.0066794
R8331 GND.n773 GND 0.00661702
R8332 GND GND.n794 0.00661702
R8333 GND.n872 GND 0.00661702
R8334 GND GND.n887 0.00661702
R8335 GND.n970 GND 0.00661702
R8336 GND.n992 GND 0.00661702
R8337 GND GND.n5879 0.00661702
R8338 GND.n5954 GND 0.00661702
R8339 GND GND.n6130 0.00661702
R8340 GND.n6035 GND 0.00661702
R8341 GND.n6083 GND 0.00661702
R8342 GND.n6105 GND 0.00661702
R8343 GND GND.n7252 0.00661702
R8344 GND.n7327 GND 0.00661702
R8345 GND GND.n7431 0.00661702
R8346 GND GND.n7384 0.00661702
R8347 GND GND.n568 0.00661702
R8348 GND.n7807 GND 0.00661702
R8349 GND.n749 GND.n745 0.00648404
R8350 GND.n932 GND.n931 0.00648404
R8351 GND.n5666 GND.n5665 0.00647015
R8352 GND.n5670 GND.n5666 0.00631395
R8353 GND.n5920 GND.n5919 0.00621809
R8354 GND.n6049 GND.n6045 0.00621809
R8355 GND.n7293 GND.n7292 0.00621809
R8356 GND.n604 GND.n603 0.00621809
R8357 GND.n6146 GND 0.00609211
R8358 GND.n6220 GND 0.00609211
R8359 GND.n5777 GND 0.00609211
R8360 GND.n5715 GND 0.00609211
R8361 GND.n4259 GND.n4257 0.00605556
R8362 GND.n1001 GND.n1000 0.00595213
R8363 GND.n5905 GND.n5904 0.00595213
R8364 GND.n5997 GND.n5967 0.00595213
R8365 GND.n6122 GND.n6120 0.00595213
R8366 GND.n7278 GND.n7277 0.00595213
R8367 GND.n7370 GND.n7340 0.00595213
R8368 GND.n7423 GND.n7421 0.00595213
R8369 GND.n6136 GND.n5653 0.00593478
R8370 GND.n5751 GND.n5750 0.00593421
R8371 GND.n1050 GND.n1048 0.00585714
R8372 GND.n5477 GND.n5475 0.00585714
R8373 GND.n233 GND.n231 0.00585714
R8374 GND.n4863 GND.n4861 0.00585714
R8375 GND.n5187 GND.n5185 0.00585714
R8376 GND.n3360 GND.n3358 0.00585714
R8377 GND.n6738 GND.n6736 0.00585714
R8378 GND.n7046 GND.n7044 0.00585714
R8379 GND.n2277 GND.n2275 0.00585714
R8380 GND.n7207 GND.n7205 0.00585714
R8381 GND.n6892 GND.n6890 0.00585714
R8382 GND.n6580 GND.n6578 0.00585714
R8383 GND.n492 GND.n490 0.00585714
R8384 GND.n344 GND.n342 0.00585714
R8385 GND.n7641 GND.n7639 0.00585714
R8386 GND.n1954 GND.n1952 0.00585714
R8387 GND.n4712 GND.n1346 0.00571186
R8388 GND.n4448 GND.n4446 0.00570833
R8389 GND.n830 GND.n826 0.00568617
R8390 GND.n3874 GND.n3860 0.00557093
R8391 GND.n836 GND.n724 0.00542021
R8392 GND.n924 GND.n881 0.00542021
R8393 GND.n6114 GND.n6113 0.00542021
R8394 GND.n7800 GND.n7798 0.00542021
R8395 GND.n5847 GND.n5846 0.00534496
R8396 GND.n5436 GND.n5435 0.00531302
R8397 GND GND.n5684 0.00510526
R8398 GND.n4061 GND.n4047 0.00507317
R8399 GND.n5397 GND.n5382 0.00507317
R8400 GND.n1261 GND.n1247 0.00507317
R8401 GND.n3054 GND.n3040 0.00507317
R8402 GND.n2903 GND.n2879 0.00507317
R8403 GND.n2638 GND.n2623 0.00507317
R8404 GND.n2164 GND.n2149 0.00507317
R8405 GND.n1433 GND.n1391 0.00507317
R8406 GND.n2473 GND.n2458 0.00507317
R8407 GND.n2807 GND.n2792 0.00507317
R8408 GND.n7730 GND.n7715 0.00507317
R8409 GND.n3155 GND.n3140 0.00507317
R8410 GND.n3262 GND.n3247 0.00507317
R8411 GND.n5066 GND.n5051 0.00507317
R8412 GND.n3672 GND.n3657 0.00507317
R8413 GND.n5834 GND.n5830 0.00505426
R8414 GND.n6145 GND 0.00502899
R8415 GND.n7436 GND.n550 0.00498679
R8416 GND.n785 GND.n724 0.0048883
R8417 GND.n881 GND.n879 0.0048883
R8418 GND.n6113 GND.n6111 0.0048883
R8419 GND.n7801 GND.n7800 0.0048883
R8420 GND.n4209 GND.n4208 0.00476136
R8421 GND.n3554 GND.n3552 0.00469846
R8422 GND.n1178 GND.n1147 0.00469846
R8423 GND.n2956 GND.n2925 0.00469846
R8424 GND.n1453 GND.n1452 0.00466667
R8425 GND.n1037 GND.n1035 0.00466667
R8426 GND.n5502 GND.n5500 0.00466667
R8427 GND.n6545 GND.n6543 0.00466667
R8428 GND.n6605 GND.n6603 0.00466667
R8429 GND.n7556 GND.n7554 0.00466667
R8430 GND.n369 GND.n367 0.00466667
R8431 GND.n5093 GND.n5092 0.00466667
R8432 GND.n5136 GND.n5134 0.00466667
R8433 GND.n3304 GND.n3303 0.00466667
R8434 GND.n3376 GND.n3374 0.00466667
R8435 GND.n3459 GND.n3457 0.00466667
R8436 GND.n1068 GND.n1066 0.00466667
R8437 GND.n6799 GND.n6797 0.00466667
R8438 GND.n6720 GND.n6717 0.00466667
R8439 GND.n7122 GND.n7120 0.00466667
R8440 GND.n7028 GND.n7025 0.00466667
R8441 GND.n1859 GND.n1857 0.00466667
R8442 GND.n1900 GND.n1898 0.00466667
R8443 GND.n2191 GND.n2189 0.00466667
R8444 GND.n2223 GND.n2221 0.00466667
R8445 GND.n6953 GND.n6951 0.00466667
R8446 GND.n6874 GND.n6871 0.00466667
R8447 GND.n83 GND.n81 0.00466667
R8448 GND.n6675 GND.n6673 0.00466667
R8449 GND.n4772 GND.n4770 0.00466667
R8450 GND.n4812 GND.n4810 0.00466667
R8451 GND.n7494 GND.n7492 0.00466667
R8452 GND.n438 GND.n436 0.00466667
R8453 GND.n7619 GND.n7617 0.00466667
R8454 GND.n258 GND.n256 0.00466667
R8455 GND.n1483 GND.n1481 0.00466667
R8456 GND.n6219 GND 0.00466667
R8457 GND.n831 GND.n830 0.00462234
R8458 GND.n5847 GND.n5682 0.00456977
R8459 GND.n7790 GND 0.00456173
R8460 GND.n5663 GND.n5662 0.00454478
R8461 GND.n4269 GND.n4268 0.00438796
R8462 GND.n4284 GND.n4283 0.00438796
R8463 GND.n4299 GND.n4298 0.00438796
R8464 GND.n4314 GND.n4313 0.00438796
R8465 GND.n4330 GND.n4329 0.00438796
R8466 GND.n4348 GND.n4347 0.00438796
R8467 GND.n4363 GND.n4362 0.00438796
R8468 GND.n4378 GND.n4377 0.00438796
R8469 GND.n4393 GND.n4392 0.00438796
R8470 GND.n4418 GND.n4417 0.00438796
R8471 GND.n4437 GND.n4436 0.00438796
R8472 GND.n4457 GND.n4456 0.00438796
R8473 GND.n4472 GND.n4471 0.00438796
R8474 GND.n4487 GND.n4486 0.00438796
R8475 GND.n4502 GND.n4501 0.00438796
R8476 GND.n4517 GND.n4516 0.00438796
R8477 GND.n4534 GND.n4533 0.00438796
R8478 GND.n4549 GND.n4548 0.00438796
R8479 GND.n4564 GND.n4563 0.00438796
R8480 GND.n4579 GND.n4578 0.00438796
R8481 GND.n4594 GND.n4593 0.00438796
R8482 GND.n4217 GND.n4216 0.00438796
R8483 GND.n4586 GND.n4585 0.00438796
R8484 GND.n4570 GND.n4569 0.00438796
R8485 GND.n4555 GND.n4554 0.00438796
R8486 GND.n4540 GND.n4539 0.00438796
R8487 GND.n4525 GND.n4524 0.00438796
R8488 GND.n4508 GND.n4507 0.00438796
R8489 GND.n4493 GND.n4492 0.00438796
R8490 GND.n4478 GND.n4477 0.00438796
R8491 GND.n4463 GND.n4462 0.00438796
R8492 GND.n4446 GND.n4445 0.00438796
R8493 GND.n4427 GND.n4426 0.00438796
R8494 GND.n4409 GND.n4408 0.00438796
R8495 GND.n4384 GND.n4383 0.00438796
R8496 GND.n4369 GND.n4368 0.00438796
R8497 GND.n4354 GND.n4353 0.00438796
R8498 GND.n4339 GND.n4338 0.00438796
R8499 GND.n4320 GND.n4319 0.00438796
R8500 GND.n4305 GND.n4304 0.00438796
R8501 GND.n4290 GND.n4289 0.00438796
R8502 GND.n4275 GND.n4274 0.00438796
R8503 GND.n1000 GND.n998 0.00435638
R8504 GND.n5967 GND.n5963 0.00435638
R8505 GND.n6123 GND.n6122 0.00435638
R8506 GND.n7340 GND.n7336 0.00435638
R8507 GND.n7424 GND.n7423 0.00435638
R8508 GND.n1548 GND.n1534 0.00425
R8509 GND.n5630 GND.n1019 0.00425
R8510 GND.n6524 GND.n6519 0.00425
R8511 GND.n7535 GND.n7530 0.00425
R8512 GND.n5235 GND.n5230 0.00425
R8513 GND.n3500 GND.n3495 0.00425
R8514 GND.n5448 GND.n1127 0.00425
R8515 GND.n6813 GND.n6781 0.00425
R8516 GND.n7101 GND.n7096 0.00425
R8517 GND.n2002 GND.n1997 0.00425
R8518 GND.n2325 GND.n2320 0.00425
R8519 GND.n6967 GND.n6935 0.00425
R8520 GND.n7739 GND.n65 0.00425
R8521 GND.n4911 GND.n4906 0.00425
R8522 GND.n7473 GND.n7468 0.00425
R8523 GND.n7598 GND.n7593 0.00425
R8524 GND.n1587 GND.n1586 0.00420666
R8525 GND.n1586 GND.n1585 0.00420666
R8526 GND.n2058 GND.n2057 0.00420666
R8527 GND.n2057 GND.n2056 0.00420666
R8528 GND.n2377 GND.n2364 0.00420666
R8529 GND.n2364 GND.n2363 0.00420666
R8530 GND.n2538 GND.n2537 0.00420666
R8531 GND.n2537 GND.n2536 0.00420666
R8532 GND.n2698 GND.n2685 0.00420666
R8533 GND.n2685 GND.n2684 0.00420666
R8534 GND.n2956 GND.n2955 0.00420666
R8535 GND.n2955 GND.n2954 0.00420666
R8536 GND.n143 GND.n130 0.00420666
R8537 GND.n130 GND.n129 0.00420666
R8538 GND.n1340 GND.n1339 0.00420666
R8539 GND.n1339 GND.n1338 0.00420666
R8540 GND.n5615 GND.n5614 0.00420666
R8541 GND.n5614 GND.n5613 0.00420666
R8542 GND.n1178 GND.n1177 0.00420666
R8543 GND.n1177 GND.n1176 0.00420666
R8544 GND.n3552 GND.n3551 0.00420666
R8545 GND.n3551 GND.n3550 0.00420666
R8546 GND.n5291 GND.n5290 0.00420666
R8547 GND.n5290 GND.n5289 0.00420666
R8548 GND.n4964 GND.n4951 0.00420666
R8549 GND.n4951 GND.n4950 0.00420666
R8550 GND.n3722 GND.n3709 0.00420666
R8551 GND.n3709 GND.n3708 0.00420666
R8552 GND.n3989 GND.n3988 0.00420666
R8553 GND.n3988 GND.n3987 0.00420666
R8554 GND.n3778 GND.n3765 0.00420666
R8555 GND.n3765 GND.n3764 0.00420666
R8556 GND.n5919 GND.n5915 0.00409043
R8557 GND.n7292 GND.n7288 0.00409043
R8558 GND.n4440 GND.n4438 0.00397222
R8559 GND.n1952 GND.n1951 0.00396756
R8560 GND.n1493 GND.n1492 0.00396756
R8561 GND.n2275 GND.n2274 0.00396756
R8562 GND.n1910 GND.n1909 0.00396756
R8563 GND.n7205 GND.n7204 0.00396756
R8564 GND.n2233 GND.n2232 0.00396756
R8565 GND.n7044 GND.n7043 0.00396756
R8566 GND.n7159 GND.n7158 0.00396756
R8567 GND.n6890 GND.n6889 0.00396756
R8568 GND.n6993 GND.n6992 0.00396756
R8569 GND.n6736 GND.n6735 0.00396756
R8570 GND.n6839 GND.n6838 0.00396756
R8571 GND.n6578 GND.n6577 0.00396756
R8572 GND.n6685 GND.n6684 0.00396756
R8573 GND.n5475 GND.n5474 0.00396756
R8574 GND.n6615 GND.n6614 0.00396756
R8575 GND.n1048 GND.n1047 0.00396756
R8576 GND.n5512 GND.n5511 0.00396756
R8577 GND.n3358 GND.n3357 0.00396756
R8578 GND.n1078 GND.n1077 0.00396756
R8579 GND.n5185 GND.n5184 0.00396756
R8580 GND.n3386 GND.n3385 0.00396756
R8581 GND.n4861 GND.n4860 0.00396756
R8582 GND.n5146 GND.n5145 0.00396756
R8583 GND.n490 GND.n489 0.00396756
R8584 GND.n4822 GND.n4821 0.00396756
R8585 GND.n342 GND.n341 0.00396756
R8586 GND.n448 GND.n447 0.00396756
R8587 GND.n231 GND.n230 0.00396756
R8588 GND.n379 GND.n378 0.00396756
R8589 GND.n7639 GND.n7638 0.00396756
R8590 GND.n268 GND.n267 0.00396756
R8591 GND.n5793 GND.n5792 0.00396053
R8592 GND.n5624 GND.n5623 0.00395031
R8593 GND.n6527 GND.n6526 0.00395031
R8594 GND.n7538 GND.n7537 0.00395031
R8595 GND.n5238 GND.n5237 0.00395031
R8596 GND.n3503 GND.n3502 0.00395031
R8597 GND.n5442 GND.n5441 0.00395031
R8598 GND.n6807 GND.n6806 0.00395031
R8599 GND.n7104 GND.n7103 0.00395031
R8600 GND.n2005 GND.n2004 0.00395031
R8601 GND.n2328 GND.n2327 0.00395031
R8602 GND.n6961 GND.n6960 0.00395031
R8603 GND.n7737 GND.n7736 0.00395031
R8604 GND.n4914 GND.n4913 0.00395031
R8605 GND.n7476 GND.n7475 0.00395031
R8606 GND.n7601 GND.n7600 0.00395031
R8607 GND.n1551 GND.n1550 0.00395031
R8608 GND.n1951 GND.n1950 0.0039133
R8609 GND.n1950 GND.t1420 0.0039133
R8610 GND.n1492 GND.n1491 0.0039133
R8611 GND.n1491 GND.t910 0.0039133
R8612 GND.n2274 GND.n2273 0.0039133
R8613 GND.n2273 GND.t847 0.0039133
R8614 GND.n1909 GND.n1908 0.0039133
R8615 GND.n1908 GND.t636 0.0039133
R8616 GND.n7204 GND.n7203 0.0039133
R8617 GND.n7203 GND.t99 0.0039133
R8618 GND.n2232 GND.n2231 0.0039133
R8619 GND.n2231 GND.t639 0.0039133
R8620 GND.n7043 GND.n7042 0.0039133
R8621 GND.n7042 GND.t141 0.0039133
R8622 GND.n7158 GND.n7157 0.0039133
R8623 GND.n7157 GND.t538 0.0039133
R8624 GND.n6889 GND.n6888 0.0039133
R8625 GND.n6888 GND.t942 0.0039133
R8626 GND.n6992 GND.n6991 0.0039133
R8627 GND.n6991 GND.t118 0.0039133
R8628 GND.n6735 GND.n6734 0.0039133
R8629 GND.n6734 GND.t1442 0.0039133
R8630 GND.n6838 GND.n6837 0.0039133
R8631 GND.n6837 GND.t185 0.0039133
R8632 GND.n6577 GND.n6576 0.0039133
R8633 GND.n6576 GND.t714 0.0039133
R8634 GND.n6684 GND.n6683 0.0039133
R8635 GND.n6683 GND.t203 0.0039133
R8636 GND.n5474 GND.n5473 0.0039133
R8637 GND.n5473 GND.t6 0.0039133
R8638 GND.n6614 GND.n6613 0.0039133
R8639 GND.n6613 GND.t566 0.0039133
R8640 GND.n1047 GND.n1046 0.0039133
R8641 GND.n1046 GND.t680 0.0039133
R8642 GND.n5511 GND.n5510 0.0039133
R8643 GND.n5510 GND.t175 0.0039133
R8644 GND.n3357 GND.n3356 0.0039133
R8645 GND.n3356 GND.t1388 0.0039133
R8646 GND.n1077 GND.n1076 0.0039133
R8647 GND.n1076 GND.t813 0.0039133
R8648 GND.n5184 GND.n5183 0.0039133
R8649 GND.n5183 GND.t515 0.0039133
R8650 GND.n3385 GND.n3384 0.0039133
R8651 GND.n3384 GND.t39 0.0039133
R8652 GND.n4860 GND.n4859 0.0039133
R8653 GND.n4859 GND.t150 0.0039133
R8654 GND.n5145 GND.n5144 0.0039133
R8655 GND.n5144 GND.t645 0.0039133
R8656 GND.n489 GND.n488 0.0039133
R8657 GND.n488 GND.t895 0.0039133
R8658 GND.n4821 GND.n4820 0.0039133
R8659 GND.n4820 GND.t79 0.0039133
R8660 GND.n341 GND.n340 0.0039133
R8661 GND.n340 GND.t698 0.0039133
R8662 GND.n447 GND.n446 0.0039133
R8663 GND.n446 GND.t242 0.0039133
R8664 GND.n230 GND.n229 0.0039133
R8665 GND.n229 GND.t259 0.0039133
R8666 GND.n378 GND.n377 0.0039133
R8667 GND.n377 GND.t1554 0.0039133
R8668 GND.n7638 GND.n7637 0.0039133
R8669 GND.n7637 GND.t727 0.0039133
R8670 GND.n267 GND.n266 0.0039133
R8671 GND.n266 GND.t1410 0.0039133
R8672 GND.n1547 GND.n1546 0.00390909
R8673 GND.n1544 GND.n1543 0.00390909
R8674 GND.n5629 GND.n5628 0.00390909
R8675 GND.n1016 GND.n1015 0.00390909
R8676 GND.n6523 GND.n6522 0.00390909
R8677 GND.n6516 GND.n6515 0.00390909
R8678 GND.n7534 GND.n7533 0.00390909
R8679 GND.n7527 GND.n7526 0.00390909
R8680 GND.n5234 GND.n5233 0.00390909
R8681 GND.n5227 GND.n5226 0.00390909
R8682 GND.n3499 GND.n3498 0.00390909
R8683 GND.n3492 GND.n3491 0.00390909
R8684 GND.n5447 GND.n5446 0.00390909
R8685 GND.n1124 GND.n1123 0.00390909
R8686 GND.n6812 GND.n6811 0.00390909
R8687 GND.n6778 GND.n6777 0.00390909
R8688 GND.n7100 GND.n7099 0.00390909
R8689 GND.n7093 GND.n7092 0.00390909
R8690 GND.n2001 GND.n2000 0.00390909
R8691 GND.n1994 GND.n1993 0.00390909
R8692 GND.n2324 GND.n2323 0.00390909
R8693 GND.n2317 GND.n2316 0.00390909
R8694 GND.n6966 GND.n6965 0.00390909
R8695 GND.n6932 GND.n6931 0.00390909
R8696 GND.n7740 GND.n64 0.00390909
R8697 GND.n61 GND.n60 0.00390909
R8698 GND.n4910 GND.n4909 0.00390909
R8699 GND.n4903 GND.n4902 0.00390909
R8700 GND.n7472 GND.n7471 0.00390909
R8701 GND.n7465 GND.n7464 0.00390909
R8702 GND.n7597 GND.n7596 0.00390909
R8703 GND.n7590 GND.n7589 0.00390909
R8704 GND.n931 GND.n929 0.00382447
R8705 GND.n6044 GND.n6042 0.00379255
R8706 GND.n7377 GND.n606 0.00379255
R8707 GND.n4670 GND.n1346 0.00377331
R8708 GND.n744 GND.n740 0.00355851
R8709 GND.n5910 GND.n5909 0.0035266
R8710 GND.n7283 GND.n7282 0.0035266
R8711 GND.n1514 GND.n1513 0.0034846
R8712 GND.n1967 GND.n1966 0.0034846
R8713 GND.n2290 GND.n2289 0.0034846
R8714 GND.n7220 GND.n7219 0.0034846
R8715 GND.n7059 GND.n7058 0.0034846
R8716 GND.n6905 GND.n6904 0.0034846
R8717 GND.n6751 GND.n6750 0.0034846
R8718 GND.n6639 GND.n6638 0.0034846
R8719 GND.n5536 GND.n5535 0.0034846
R8720 GND.n1102 GND.n1101 0.0034846
R8721 GND.n3410 GND.n3409 0.0034846
R8722 GND.n5200 GND.n5199 0.0034846
R8723 GND.n4876 GND.n4875 0.0034846
R8724 GND.n505 GND.n504 0.0034846
R8725 GND.n403 GND.n402 0.0034846
R8726 GND.n292 GND.n291 0.0034846
R8727 GND.n1513 GND.n1512 0.00343883
R8728 GND.n1512 GND.n1511 0.00343883
R8729 GND.n1963 GND.n1962 0.00343883
R8730 GND.n1964 GND.n1963 0.00343883
R8731 GND.n1966 GND.n1965 0.00343883
R8732 GND.n1965 GND.n1964 0.00343883
R8733 GND.n2286 GND.n2285 0.00343883
R8734 GND.n2287 GND.n2286 0.00343883
R8735 GND.n2289 GND.n2288 0.00343883
R8736 GND.n2288 GND.n2287 0.00343883
R8737 GND.n7216 GND.n7215 0.00343883
R8738 GND.n7217 GND.n7216 0.00343883
R8739 GND.n7219 GND.n7218 0.00343883
R8740 GND.n7218 GND.n7217 0.00343883
R8741 GND.n7055 GND.n7054 0.00343883
R8742 GND.n7056 GND.n7055 0.00343883
R8743 GND.n7058 GND.n7057 0.00343883
R8744 GND.n7057 GND.n7056 0.00343883
R8745 GND.n6901 GND.n6900 0.00343883
R8746 GND.n6902 GND.n6901 0.00343883
R8747 GND.n6904 GND.n6903 0.00343883
R8748 GND.n6903 GND.n6902 0.00343883
R8749 GND.n6747 GND.n6746 0.00343883
R8750 GND.n6748 GND.n6747 0.00343883
R8751 GND.n6750 GND.n6749 0.00343883
R8752 GND.n6749 GND.n6748 0.00343883
R8753 GND.n6643 GND.n6642 0.00343883
R8754 GND.n6642 GND.n6641 0.00343883
R8755 GND.n6640 GND.n6639 0.00343883
R8756 GND.n6641 GND.n6640 0.00343883
R8757 GND.n5540 GND.n5539 0.00343883
R8758 GND.n5539 GND.n5538 0.00343883
R8759 GND.n5537 GND.n5536 0.00343883
R8760 GND.n5538 GND.n5537 0.00343883
R8761 GND.n1106 GND.n1105 0.00343883
R8762 GND.n1105 GND.n1104 0.00343883
R8763 GND.n1103 GND.n1102 0.00343883
R8764 GND.n1104 GND.n1103 0.00343883
R8765 GND.n3414 GND.n3413 0.00343883
R8766 GND.n3413 GND.n3412 0.00343883
R8767 GND.n3411 GND.n3410 0.00343883
R8768 GND.n3412 GND.n3411 0.00343883
R8769 GND.n5196 GND.n5195 0.00343883
R8770 GND.n5197 GND.n5196 0.00343883
R8771 GND.n5199 GND.n5198 0.00343883
R8772 GND.n5198 GND.n5197 0.00343883
R8773 GND.n4872 GND.n4871 0.00343883
R8774 GND.n4873 GND.n4872 0.00343883
R8775 GND.n4875 GND.n4874 0.00343883
R8776 GND.n4874 GND.n4873 0.00343883
R8777 GND.n501 GND.n500 0.00343883
R8778 GND.n502 GND.n501 0.00343883
R8779 GND.n504 GND.n503 0.00343883
R8780 GND.n503 GND.n502 0.00343883
R8781 GND.n407 GND.n406 0.00343883
R8782 GND.n406 GND.n405 0.00343883
R8783 GND.n404 GND.n403 0.00343883
R8784 GND.n405 GND.n404 0.00343883
R8785 GND.n296 GND.n295 0.00343883
R8786 GND.n295 GND.n294 0.00343883
R8787 GND.n293 GND.n292 0.00343883
R8788 GND.n294 GND.n293 0.00343883
R8789 GND.n7650 GND.n7649 0.00343883
R8790 GND.n7651 GND.n7650 0.00343883
R8791 GND GND.n6376 0.00340123
R8792 GND.n7790 GND 0.00340123
R8793 GND.n6209 GND 0.00327778
R8794 GND.n6202 GND 0.00327778
R8795 GND.n6146 GND.n6145 0.00313158
R8796 GND.n2196 GND.n2195 0.00308428
R8797 GND.n6419 GND.n6418 0.00307458
R8798 GND.n980 GND.n978 0.0030266
R8799 GND.n5996 GND.n5994 0.0030266
R8800 GND.n6001 GND.n5855 0.0030266
R8801 GND.n7369 GND.n7367 0.0030266
R8802 GND.n7420 GND.n7416 0.0030266
R8803 GND.n1534 GND.n1533 0.003
R8804 GND.n1019 GND.n1018 0.003
R8805 GND.n6519 GND.n6518 0.003
R8806 GND.n7530 GND.n7529 0.003
R8807 GND.n5230 GND.n5229 0.003
R8808 GND.n3495 GND.n3494 0.003
R8809 GND.n1127 GND.n1126 0.003
R8810 GND.n6781 GND.n6780 0.003
R8811 GND.n7096 GND.n7095 0.003
R8812 GND.n1997 GND.n1996 0.003
R8813 GND.n2320 GND.n2319 0.003
R8814 GND.n6935 GND.n6934 0.003
R8815 GND.n4906 GND.n4905 0.003
R8816 GND.n7468 GND.n7467 0.003
R8817 GND.n7593 GND.n7592 0.003
R8818 GND.n4263 GND.n4262 0.00299232
R8819 GND.n5830 GND.n5829 0.00292248
R8820 GND.n6452 GND.n6451 0.00290385
R8821 GND.n549 GND.n548 0.00290385
R8822 GND.n2168 GND.n2167 0.00285
R8823 GND.n2477 GND.n2476 0.00285
R8824 GND.n2642 GND.n2641 0.00285
R8825 GND.n2811 GND.n2810 0.00285
R8826 GND.n2962 GND.n2961 0.00285
R8827 GND.n7733 GND.n150 0.00285
R8828 GND.n5406 GND.n5400 0.00285
R8829 GND.n5075 GND.n5069 0.00285
R8830 GND.n5410 GND.n3730 0.00285
R8831 GND.n4087 GND.n4086 0.00285
R8832 GND.n4108 GND.n3904 0.00285
R8833 GND.n3561 GND.n3560 0.00285
R8834 GND.n5438 GND.n5437 0.00285
R8835 GND.n5428 GND.n1595 0.00285
R8836 GND.n6223 GND.n6221 0.00280263
R8837 GND.n6474 GND.n6471 0.00277946
R8838 GND.n6384 GND.n6381 0.00277946
R8839 GND.n770 GND 0.00276064
R8840 GND.n795 GND 0.00276064
R8841 GND.n869 GND 0.00276064
R8842 GND.n888 GND 0.00276064
R8843 GND.n967 GND 0.00276064
R8844 GND GND.n980 0.00276064
R8845 GND.n995 GND 0.00276064
R8846 GND.n983 GND 0.00276064
R8847 GND.n5880 GND 0.00276064
R8848 GND.n5951 GND 0.00276064
R8849 GND.n6131 GND 0.00276064
R8850 GND.n6032 GND 0.00276064
R8851 GND.n6080 GND 0.00276064
R8852 GND GND.n6093 0.00276064
R8853 GND.n6108 GND 0.00276064
R8854 GND.n6096 GND 0.00276064
R8855 GND.n7253 GND 0.00276064
R8856 GND.n7324 GND 0.00276064
R8857 GND.n7432 GND 0.00276064
R8858 GND.n7385 GND 0.00276064
R8859 GND.n569 GND 0.00276064
R8860 GND.n2 GND 0.00276064
R8861 GND.n7804 GND 0.00276064
R8862 GND GND.n7817 0.00276064
R8863 GND.n1427 GND.n1426 0.00266776
R8864 GND.n2467 GND.n2466 0.00266776
R8865 GND.n2801 GND.n2800 0.00266776
R8866 GND.n7724 GND.n7723 0.00266776
R8867 GND.n3149 GND.n3148 0.00266776
R8868 GND.n3256 GND.n3255 0.00266776
R8869 GND.n5060 GND.n5059 0.00266776
R8870 GND.n3666 GND.n3665 0.00266776
R8871 GND.n5512 GND.n5508 0.00258333
R8872 GND.n6615 GND.n6611 0.00258333
R8873 GND.n379 GND.n375 0.00258333
R8874 GND.n5146 GND.n5142 0.00258333
R8875 GND.n3386 GND.n3382 0.00258333
R8876 GND.n1078 GND.n1074 0.00258333
R8877 GND.n6839 GND.n6835 0.00258333
R8878 GND.n7159 GND.n7155 0.00258333
R8879 GND.n1910 GND.n1906 0.00258333
R8880 GND.n2233 GND.n2229 0.00258333
R8881 GND.n6993 GND.n6989 0.00258333
R8882 GND.n6685 GND.n6681 0.00258333
R8883 GND.n4822 GND.n4818 0.00258333
R8884 GND.n448 GND.n444 0.00258333
R8885 GND.n268 GND.n264 0.00258333
R8886 GND.n1493 GND.n1489 0.00258333
R8887 GND.n4626 GND.n4625 0.00253688
R8888 GND.n4617 GND.n4616 0.00253688
R8889 GND.n4600 GND.n4599 0.00250907
R8890 GND.n4588 GND.n4587 0.00250907
R8891 GND.n4572 GND.n4571 0.00250907
R8892 GND.n4557 GND.n4556 0.00250907
R8893 GND.n4542 GND.n4541 0.00250907
R8894 GND.n4527 GND.n4526 0.00250907
R8895 GND.n4510 GND.n4509 0.00250907
R8896 GND.n4495 GND.n4494 0.00250907
R8897 GND.n4480 GND.n4479 0.00250907
R8898 GND.n4465 GND.n4464 0.00250907
R8899 GND.n4450 GND.n4449 0.00250907
R8900 GND.n4429 GND.n4428 0.00250907
R8901 GND.n4411 GND.n4410 0.00250907
R8902 GND.n4386 GND.n4385 0.00250907
R8903 GND.n4371 GND.n4370 0.00250907
R8904 GND.n4356 GND.n4355 0.00250907
R8905 GND.n4341 GND.n4340 0.00250907
R8906 GND.n4322 GND.n4321 0.00250907
R8907 GND.n4307 GND.n4306 0.00250907
R8908 GND.n4292 GND.n4291 0.00250907
R8909 GND.n4277 GND.n4276 0.00250907
R8910 GND.n4267 GND.n4266 0.00250907
R8911 GND.n4282 GND.n4281 0.00250907
R8912 GND.n4297 GND.n4296 0.00250907
R8913 GND.n4312 GND.n4311 0.00250907
R8914 GND.n4327 GND.n4326 0.00250907
R8915 GND.n4346 GND.n4345 0.00250907
R8916 GND.n4361 GND.n4360 0.00250907
R8917 GND.n4376 GND.n4375 0.00250907
R8918 GND.n4391 GND.n4390 0.00250907
R8919 GND.n4416 GND.n4415 0.00250907
R8920 GND.n4434 GND.n4433 0.00250907
R8921 GND.n4455 GND.n4454 0.00250907
R8922 GND.n4470 GND.n4469 0.00250907
R8923 GND.n4485 GND.n4484 0.00250907
R8924 GND.n4500 GND.n4499 0.00250907
R8925 GND.n4515 GND.n4514 0.00250907
R8926 GND.n4532 GND.n4531 0.00250907
R8927 GND.n4547 GND.n4546 0.00250907
R8928 GND.n4562 GND.n4561 0.00250907
R8929 GND.n4577 GND.n4576 0.00250907
R8930 GND.n4592 GND.n4591 0.00250907
R8931 GND.n4596 GND.n4595 0.00250907
R8932 GND.n839 GND.n838 0.00249468
R8933 GND.n923 GND.n919 0.00249468
R8934 GND.n6093 GND.n6091 0.00249468
R8935 GND.n3 GND.n2 0.00249468
R8936 GND.n4265 GND.t1497 0.00247763
R8937 GND.n4280 GND.t1501 0.00247763
R8938 GND.n4295 GND.t1565 0.00247763
R8939 GND.n4310 GND.t215 0.00247763
R8940 GND.n4325 GND.t1561 0.00247763
R8941 GND.n4344 GND.t1498 0.00247763
R8942 GND.n4359 GND.t213 0.00247763
R8943 GND.n4374 GND.t1499 0.00247763
R8944 GND.n4389 GND.t218 0.00247763
R8945 GND.n4414 GND.t214 0.00247763
R8946 GND.n4432 GND.t827 0.00247763
R8947 GND.n4453 GND.t1496 0.00247763
R8948 GND.n4468 GND.t1562 0.00247763
R8949 GND.n4483 GND.t1494 0.00247763
R8950 GND.n4498 GND.t216 0.00247763
R8951 GND.n4513 GND.t1564 0.00247763
R8952 GND.n4530 GND.t1500 0.00247763
R8953 GND.n4545 GND.t1563 0.00247763
R8954 GND.n4560 GND.t1495 0.00247763
R8955 GND.n4575 GND.t217 0.00247763
R8956 GND.n4573 GND.n4572 0.00247763
R8957 GND.t217 GND.n4573 0.00247763
R8958 GND.n4558 GND.n4557 0.00247763
R8959 GND.t1495 GND.n4558 0.00247763
R8960 GND.n4543 GND.n4542 0.00247763
R8961 GND.t1563 GND.n4543 0.00247763
R8962 GND.n4528 GND.n4527 0.00247763
R8963 GND.t1500 GND.n4528 0.00247763
R8964 GND.n4511 GND.n4510 0.00247763
R8965 GND.t1564 GND.n4511 0.00247763
R8966 GND.n4496 GND.n4495 0.00247763
R8967 GND.t216 GND.n4496 0.00247763
R8968 GND.n4481 GND.n4480 0.00247763
R8969 GND.t1494 GND.n4481 0.00247763
R8970 GND.n4466 GND.n4465 0.00247763
R8971 GND.t1562 GND.n4466 0.00247763
R8972 GND.n4451 GND.n4450 0.00247763
R8973 GND.t1496 GND.n4451 0.00247763
R8974 GND.n4430 GND.n4429 0.00247763
R8975 GND.t827 GND.n4430 0.00247763
R8976 GND.n4412 GND.n4411 0.00247763
R8977 GND.t214 GND.n4412 0.00247763
R8978 GND.n4387 GND.n4386 0.00247763
R8979 GND.t218 GND.n4387 0.00247763
R8980 GND.n4372 GND.n4371 0.00247763
R8981 GND.t1499 GND.n4372 0.00247763
R8982 GND.n4357 GND.n4356 0.00247763
R8983 GND.t213 GND.n4357 0.00247763
R8984 GND.n4342 GND.n4341 0.00247763
R8985 GND.t1498 GND.n4342 0.00247763
R8986 GND.n4323 GND.n4322 0.00247763
R8987 GND.t1561 GND.n4323 0.00247763
R8988 GND.n4308 GND.n4307 0.00247763
R8989 GND.t215 GND.n4308 0.00247763
R8990 GND.n4293 GND.n4292 0.00247763
R8991 GND.t1565 GND.n4293 0.00247763
R8992 GND.n4278 GND.n4277 0.00247763
R8993 GND.t1501 GND.n4278 0.00247763
R8994 GND.n4264 GND.n4263 0.00247763
R8995 GND.t1497 GND.n4264 0.00247763
R8996 GND.n4266 GND.n4265 0.00247763
R8997 GND.n4281 GND.n4280 0.00247763
R8998 GND.n4296 GND.n4295 0.00247763
R8999 GND.n4311 GND.n4310 0.00247763
R9000 GND.n4326 GND.n4325 0.00247763
R9001 GND.n4345 GND.n4344 0.00247763
R9002 GND.n4360 GND.n4359 0.00247763
R9003 GND.n4375 GND.n4374 0.00247763
R9004 GND.n4390 GND.n4389 0.00247763
R9005 GND.n4415 GND.n4414 0.00247763
R9006 GND.n4433 GND.n4432 0.00247763
R9007 GND.n4454 GND.n4453 0.00247763
R9008 GND.n4469 GND.n4468 0.00247763
R9009 GND.n4484 GND.n4483 0.00247763
R9010 GND.n4499 GND.n4498 0.00247763
R9011 GND.n4514 GND.n4513 0.00247763
R9012 GND.n4531 GND.n4530 0.00247763
R9013 GND.n4546 GND.n4545 0.00247763
R9014 GND.n4561 GND.n4560 0.00247763
R9015 GND.n4576 GND.n4575 0.00247763
R9016 GND.n4591 GND.n4590 0.00247763
R9017 GND.n4590 GND.t1566 0.00247763
R9018 GND.n4589 GND.n4588 0.00247763
R9019 GND.t1566 GND.n4589 0.00247763
R9020 GND.n4599 GND.n4598 0.00247763
R9021 GND.n4598 GND.t501 0.00247763
R9022 GND.t501 GND.n4597 0.00247763
R9023 GND.n4597 GND.n4596 0.00247763
R9024 GND.n6219 GND 0.00247368
R9025 GND.n1550 GND.n1549 0.00245833
R9026 GND.n5625 GND.n5624 0.00245833
R9027 GND.n6526 GND.n6525 0.00245833
R9028 GND.n7537 GND.n7536 0.00245833
R9029 GND.n5237 GND.n5236 0.00245833
R9030 GND.n3502 GND.n3501 0.00245833
R9031 GND.n5443 GND.n5442 0.00245833
R9032 GND.n6808 GND.n6807 0.00245833
R9033 GND.n7103 GND.n7102 0.00245833
R9034 GND.n2004 GND.n2003 0.00245833
R9035 GND.n2327 GND.n2326 0.00245833
R9036 GND.n6962 GND.n6961 0.00245833
R9037 GND.n7738 GND.n7737 0.00245833
R9038 GND.n4913 GND.n4912 0.00245833
R9039 GND.n7475 GND.n7474 0.00245833
R9040 GND.n7600 GND.n7599 0.00245833
R9041 GND.n5535 GND.n5534 0.00228571
R9042 GND.n6638 GND.n6637 0.00228571
R9043 GND.n402 GND.n401 0.00228571
R9044 GND.n5200 GND.n5168 0.00228571
R9045 GND.n3409 GND.n3408 0.00228571
R9046 GND.n1101 GND.n1100 0.00228571
R9047 GND.n6905 GND.n6861 0.00228571
R9048 GND.n7220 GND.n7181 0.00228571
R9049 GND.n1967 GND.n1932 0.00228571
R9050 GND.n2290 GND.n2255 0.00228571
R9051 GND.n7059 GND.n7015 0.00228571
R9052 GND.n6751 GND.n6707 0.00228571
R9053 GND.n4876 GND.n4844 0.00228571
R9054 GND.n505 GND.n470 0.00228571
R9055 GND.n291 GND.n290 0.00228571
R9056 GND.n1514 GND.n1510 0.00228571
R9057 GND.n4008 GND 0.00217027
R9058 GND.n1410 GND 0.00217027
R9059 GND.n2077 GND 0.00217027
R9060 GND.n2399 GND 0.00217027
R9061 GND.n2557 GND 0.00217027
R9062 GND.n2720 GND 0.00217027
R9063 GND.n2828 GND 0.00217027
R9064 GND.n159 GND 0.00217027
R9065 GND.n2994 GND 0.00217027
R9066 GND.n3103 GND 0.00217027
R9067 GND.n5310 GND 0.00217027
R9068 GND.n4985 GND 0.00217027
R9069 GND.n3591 GND 0.00217027
R9070 GND.n3794 GND 0.00217027
R9071 GND.n3217 GND 0.00217027
R9072 GND.n1204 GND 0.00217027
R9073 GND.n4085 GND.n4084 0.00199276
R9074 GND.n1285 GND.n1284 0.00199276
R9075 GND.n3078 GND.n3077 0.00199276
R9076 GND.n3903 GND.n3902 0.00199276
R9077 GND.n6384 GND.n6383 0.00193331
R9078 GND.n6474 GND.n6473 0.00193331
R9079 GND.n4438 GND.n4437 0.00188889
R9080 GND.n4184 GND.n4183 0.00186977
R9081 GND.n4185 GND.n4184 0.00186977
R9082 GND.n1481 GND.n1480 0.00183506
R9083 GND.n1898 GND.n1897 0.00183506
R9084 GND.n2221 GND.n2220 0.00183506
R9085 GND.n7028 GND.n7027 0.00183506
R9086 GND.n6874 GND.n6873 0.00183506
R9087 GND.n6720 GND.n6719 0.00183506
R9088 GND.n6673 GND.n6672 0.00183506
R9089 GND.n6603 GND.n6602 0.00183506
R9090 GND.n5500 GND.n5499 0.00183506
R9091 GND.n1066 GND.n1065 0.00183506
R9092 GND.n3374 GND.n3373 0.00183506
R9093 GND.n5134 GND.n5133 0.00183506
R9094 GND.n4810 GND.n4809 0.00183506
R9095 GND.n436 GND.n435 0.00183506
R9096 GND.n367 GND.n366 0.00183506
R9097 GND.n256 GND.n255 0.00183506
R9098 GND.n1480 GND.n1479 0.00181454
R9099 GND.n1943 GND.n1942 0.00181454
R9100 GND.n1942 GND.n1941 0.00181454
R9101 GND.n1897 GND.n1896 0.00181454
R9102 GND.n2261 GND.n2260 0.00181454
R9103 GND.n2260 GND.n2259 0.00181454
R9104 GND.n2220 GND.n2219 0.00181454
R9105 GND.n7189 GND.n7188 0.00181454
R9106 GND.n7188 GND.n7187 0.00181454
R9107 GND.n7027 GND.n7026 0.00181454
R9108 GND.n7023 GND.n7022 0.00181454
R9109 GND.n7022 GND.n7021 0.00181454
R9110 GND.n6873 GND.n6872 0.00181454
R9111 GND.n6869 GND.n6868 0.00181454
R9112 GND.n6868 GND.n6867 0.00181454
R9113 GND.n6719 GND.n6718 0.00181454
R9114 GND.n6715 GND.n6714 0.00181454
R9115 GND.n6714 GND.n6713 0.00181454
R9116 GND.n6672 GND.n6671 0.00181454
R9117 GND.n6567 GND.n6566 0.00181454
R9118 GND.n6566 GND.n6565 0.00181454
R9119 GND.n6602 GND.n6601 0.00181454
R9120 GND.n6592 GND.n6591 0.00181454
R9121 GND.n6591 GND.n6590 0.00181454
R9122 GND.n5499 GND.n5498 0.00181454
R9123 GND.n5489 GND.n5488 0.00181454
R9124 GND.n5488 GND.n5487 0.00181454
R9125 GND.n1065 GND.n1064 0.00181454
R9126 GND.n3349 GND.n3348 0.00181454
R9127 GND.n3348 GND.n3347 0.00181454
R9128 GND.n3373 GND.n3372 0.00181454
R9129 GND.n5174 GND.n5173 0.00181454
R9130 GND.n5173 GND.n5172 0.00181454
R9131 GND.n5133 GND.n5132 0.00181454
R9132 GND.n4850 GND.n4849 0.00181454
R9133 GND.n4849 GND.n4848 0.00181454
R9134 GND.n4809 GND.n4808 0.00181454
R9135 GND.n476 GND.n475 0.00181454
R9136 GND.n475 GND.n474 0.00181454
R9137 GND.n435 GND.n434 0.00181454
R9138 GND.n331 GND.n330 0.00181454
R9139 GND.n330 GND.n329 0.00181454
R9140 GND.n366 GND.n365 0.00181454
R9141 GND.n356 GND.n355 0.00181454
R9142 GND.n355 GND.n354 0.00181454
R9143 GND.n255 GND.n254 0.00181454
R9144 GND.n245 GND.n244 0.00181454
R9145 GND.n244 GND.n243 0.00181454
R9146 GND.n2168 GND 0.00175333
R9147 GND.n2477 GND 0.00175333
R9148 GND.n2642 GND 0.00175333
R9149 GND.n2811 GND 0.00175333
R9150 GND.n2962 GND 0.00175333
R9151 GND GND.n150 0.00175333
R9152 GND GND.n5406 0.00175333
R9153 GND GND.n5075 0.00175333
R9154 GND.n5410 GND 0.00175333
R9155 GND.n4087 GND 0.00175333
R9156 GND GND.n4108 0.00175333
R9157 GND.n3561 GND 0.00175333
R9158 GND.n5437 GND 0.00175333
R9159 GND GND.n5428 0.00175333
R9160 GND.n6483 GND.n6477 0.00175
R9161 GND.n6487 GND.n6486 0.00175
R9162 GND.n6489 GND.n6475 0.00175
R9163 GND.n6393 GND.n6387 0.00175
R9164 GND.n6397 GND.n6396 0.00175
R9165 GND.n6399 GND.n6385 0.00175
R9166 GND.n3940 GND.n3939 0.00174202
R9167 GND.n5242 GND.n5241 0.00174202
R9168 GND.n3556 GND.n3554 0.00174202
R9169 GND.n5618 GND.n5617 0.00174202
R9170 GND.n1291 GND.n1290 0.00174202
R9171 GND.n2489 GND.n2488 0.00174202
R9172 GND.n2009 GND.n2008 0.00174202
R9173 GND.n1591 GND.n1589 0.00174202
R9174 GND.n4740 GND.n4739 0.00172549
R9175 GND.n2159 GND.n2157 0.001708
R9176 GND.n2633 GND.n2631 0.001708
R9177 GND.n2898 GND.n2897 0.001708
R9178 GND.n3050 GND.n3048 0.001708
R9179 GND.n1257 GND.n1255 0.001708
R9180 GND.n5392 GND.n5390 0.001708
R9181 GND.n4057 GND.n4055 0.001708
R9182 GND.n3870 GND.n3868 0.001708
R9183 GND.n782 GND.n780 0.00169681
R9184 GND.n6114 GND 0.00169681
R9185 GND.n7798 GND 0.00169681
R9186 GND.n4674 GND.n4672 0.00166525
R9187 GND.n1530 GND.n1527 0.00163636
R9188 GND.n5634 GND.n5633 0.00163636
R9189 GND.n6506 GND.n6503 0.00163636
R9190 GND.n7517 GND.n7514 0.00163636
R9191 GND.n5217 GND.n5214 0.00163636
R9192 GND.n3482 GND.n3479 0.00163636
R9193 GND.n5452 GND.n5451 0.00163636
R9194 GND.n6817 GND.n6816 0.00163636
R9195 GND.n7083 GND.n7080 0.00163636
R9196 GND.n1984 GND.n1981 0.00163636
R9197 GND.n2307 GND.n2304 0.00163636
R9198 GND.n6971 GND.n6970 0.00163636
R9199 GND.n7745 GND.n7744 0.00163636
R9200 GND.n4893 GND.n4890 0.00163636
R9201 GND.n7455 GND.n7452 0.00163636
R9202 GND.n7580 GND.n7577 0.00163636
R9203 GND.n1440 GND.n1438 0.00154167
R9204 GND.n1024 GND.n1022 0.00154167
R9205 GND.n6532 GND.n6530 0.00154167
R9206 GND.n7543 GND.n7541 0.00154167
R9207 GND.n5080 GND.n5078 0.00154167
R9208 GND.n3291 GND.n3289 0.00154167
R9209 GND.n3446 GND.n3444 0.00154167
R9210 GND.n6786 GND.n6784 0.00154167
R9211 GND.n7109 GND.n7107 0.00154167
R9212 GND.n1846 GND.n1844 0.00154167
R9213 GND.n2181 GND.n2179 0.00154167
R9214 GND.n6940 GND.n6938 0.00154167
R9215 GND.n70 GND.n68 0.00154167
R9216 GND.n4759 GND.n4757 0.00154167
R9217 GND.n7481 GND.n7479 0.00154167
R9218 GND.n7606 GND.n7604 0.00154167
R9219 GND.n1433 GND.n1432 0.00150729
R9220 GND.n2164 GND.n2163 0.00150729
R9221 GND.n2473 GND.n2472 0.00150729
R9222 GND.n2638 GND.n2637 0.00150729
R9223 GND.n2807 GND.n2806 0.00150729
R9224 GND.n2903 GND.n2902 0.00150729
R9225 GND.n7730 GND.n7729 0.00150729
R9226 GND.n3155 GND.n3154 0.00150729
R9227 GND.n3262 GND.n3261 0.00150729
R9228 GND.n5397 GND.n5396 0.00150729
R9229 GND.n5066 GND.n5065 0.00150729
R9230 GND.n2379 GND.n2377 0.00150234
R9231 GND.n2700 GND.n2698 0.00150234
R9232 GND.n145 GND.n143 0.00150234
R9233 GND.n4966 GND.n4964 0.00150234
R9234 GND.n3724 GND.n3722 0.00150234
R9235 GND.n3780 GND.n3778 0.00150234
R9236 GND.n7437 GND.n7436 0.00150166
R9237 GND.n2380 GND.n2379 0.00150164
R9238 GND.n2701 GND.n2700 0.00150164
R9239 GND.n146 GND.n145 0.00150164
R9240 GND.n4967 GND.n4966 0.00150164
R9241 GND.n3725 GND.n3724 0.00150164
R9242 GND.n3781 GND.n3780 0.00150164
R9243 GND.n6453 GND.n676 0.00150121
R9244 GND.n5825 GND.n5684 0.00148684
R9245 GND.n4006 GND.n4004 0.00139286
R9246 GND.n1408 GND.n1404 0.00139286
R9247 GND.n2075 GND.n2073 0.00139286
R9248 GND.n2397 GND.n2395 0.00139286
R9249 GND.n2555 GND.n2553 0.00139286
R9250 GND.n2718 GND.n2716 0.00139286
R9251 GND.n2839 GND.n2821 0.00139286
R9252 GND.n7660 GND.n152 0.00139286
R9253 GND.n2992 GND.n2990 0.00139286
R9254 GND.n3101 GND.n3099 0.00139286
R9255 GND.n5308 GND.n5306 0.00139286
R9256 GND.n4983 GND.n4981 0.00139286
R9257 GND.n3589 GND.n3587 0.00139286
R9258 GND.n3806 GND.n3787 0.00139286
R9259 GND.n3215 GND.n3213 0.00139286
R9260 GND.n1202 GND.n1200 0.00139286
R9261 GND.n4013 GND.n4007 0.00138653
R9262 GND.n1415 GND.n1409 0.00138653
R9263 GND.n2082 GND.n2076 0.00138653
R9264 GND.n2404 GND.n2398 0.00138653
R9265 GND.n2562 GND.n2556 0.00138653
R9266 GND.n2725 GND.n2719 0.00138653
R9267 GND.n2837 GND.n2836 0.00138653
R9268 GND.n7658 GND.n7657 0.00138653
R9269 GND.n2999 GND.n2993 0.00138653
R9270 GND.n3108 GND.n3102 0.00138653
R9271 GND.n5315 GND.n5309 0.00138653
R9272 GND.n4990 GND.n4984 0.00138653
R9273 GND.n3596 GND.n3590 0.00138653
R9274 GND.n3804 GND.n3803 0.00138653
R9275 GND.n3222 GND.n3216 0.00138653
R9276 GND.n1209 GND.n1203 0.00138653
R9277 GND.n4094 GND.n4091 0.00132676
R9278 GND.n5423 GND.n5422 0.0013267
R9279 GND.n2175 GND.n2172 0.0013267
R9280 GND.n2484 GND.n2481 0.0013267
R9281 GND.n2649 GND.n2646 0.0013267
R9282 GND.n2818 GND.n2815 0.0013267
R9283 GND.n2970 GND.n2967 0.0013267
R9284 GND.n2978 GND.n2975 0.0013267
R9285 GND.n3088 GND.n3085 0.0013267
R9286 GND.n3189 GND.n3186 0.0013267
R9287 GND.n3195 GND.n3192 0.0013267
R9288 GND.n3569 GND.n3566 0.0013267
R9289 GND.n5401 GND.n3572 0.0013267
R9290 GND.n5070 GND.n3575 0.0013267
R9291 GND.n5418 GND.n5415 0.0013267
R9292 GND.n4103 GND.n4102 0.0013267
R9293 GND.n1472 GND.t820 0.00131092
R9294 GND.n1473 GND.n1472 0.00131092
R9295 GND.n1880 GND.n1879 0.00131092
R9296 GND.t914 GND.n1880 0.00131092
R9297 GND.n1889 GND.t914 0.00131092
R9298 GND.n1890 GND.n1889 0.00131092
R9299 GND.n2206 GND.n2205 0.00131092
R9300 GND.t868 GND.n2206 0.00131092
R9301 GND.n2214 GND.t868 0.00131092
R9302 GND.n2215 GND.n2214 0.00131092
R9303 GND.n7137 GND.n7136 0.00131092
R9304 GND.t1403 GND.n7137 0.00131092
R9305 GND.n7145 GND.t1403 0.00131092
R9306 GND.n7146 GND.n7145 0.00131092
R9307 GND.n7067 GND.n7066 0.00131092
R9308 GND.n7066 GND.t525 0.00131092
R9309 GND.t525 GND.n7065 0.00131092
R9310 GND.n7065 GND.n7064 0.00131092
R9311 GND.n6913 GND.n6912 0.00131092
R9312 GND.n6912 GND.t621 0.00131092
R9313 GND.t621 GND.n6911 0.00131092
R9314 GND.n6911 GND.n6910 0.00131092
R9315 GND.n6759 GND.n6758 0.00131092
R9316 GND.n6758 GND.t936 0.00131092
R9317 GND.t936 GND.n6757 0.00131092
R9318 GND.n6757 GND.n6756 0.00131092
R9319 GND.n6560 GND.n6559 0.00131092
R9320 GND.n6559 GND.t226 0.00131092
R9321 GND.t226 GND.n6558 0.00131092
R9322 GND.n6558 GND.n6557 0.00131092
R9323 GND.n5549 GND.n5548 0.00131092
R9324 GND.t0 GND.n5549 0.00131092
R9325 GND.n5557 GND.t0 0.00131092
R9326 GND.n5558 GND.n5557 0.00131092
R9327 GND.n3427 GND.n3426 0.00131092
R9328 GND.t623 GND.n3427 0.00131092
R9329 GND.n3435 GND.t623 0.00131092
R9330 GND.n3436 GND.n3435 0.00131092
R9331 GND.n3342 GND.n3341 0.00131092
R9332 GND.n3341 GND.t536 0.00131092
R9333 GND.n3324 GND.n3323 0.00131092
R9334 GND.n5114 GND.n5113 0.00131092
R9335 GND.t1488 GND.n5114 0.00131092
R9336 GND.n5122 GND.t1488 0.00131092
R9337 GND.n5123 GND.n5122 0.00131092
R9338 GND.n4793 GND.n4792 0.00131092
R9339 GND.t423 GND.n4793 0.00131092
R9340 GND.n4801 GND.t423 0.00131092
R9341 GND.n4802 GND.n4801 0.00131092
R9342 GND.n416 GND.n415 0.00131092
R9343 GND.t550 GND.n416 0.00131092
R9344 GND.n424 GND.t550 0.00131092
R9345 GND.n425 GND.n424 0.00131092
R9346 GND.n324 GND.n323 0.00131092
R9347 GND.n323 GND.t568 0.00131092
R9348 GND.t568 GND.n322 0.00131092
R9349 GND.n322 GND.n321 0.00131092
R9350 GND.n222 GND.n221 0.00131092
R9351 GND.n221 GND.t719 0.00131092
R9352 GND.t719 GND.n220 0.00131092
R9353 GND.n220 GND.n219 0.00131092
R9354 GND.n194 GND.n193 0.00131092
R9355 GND.n193 GND.t625 0.00131092
R9356 GND.n4616 GND.n4615 0.00125043
R9357 GND GND.n4674 0.00124153
R9358 GND.n5741 GND.n5740 0.00122464
R9359 GND.n1001 GND 0.00116489
R9360 GND.n5872 GND.n5857 0.00116489
R9361 GND.n7245 GND.n7231 0.00116489
R9362 GND.n7443 GND.n7441 0.00115206
R9363 GND.n7443 GND.n7442 0.00115206
R9364 GND.n4750 GND.n4627 0.00114322
R9365 GND.n6458 GND.n6457 0.00109111
R9366 GND.n6491 GND.n6474 0.00108327
R9367 GND.n6401 GND.n6384 0.00108327
R9368 GND.n6457 GND.n6456 0.00107707
R9369 GND.n7441 GND.n7440 0.00107707
R9370 GND.n6375 GND.n6374 0.00107231
R9371 GND.n7793 GND.n7791 0.00107231
R9372 GND.n2847 GND.n2846 0.00103916
R9373 GND.n1358 GND.n1357 0.00103916
R9374 GND.n2106 GND.n2105 0.00103916
R9375 GND.n2429 GND.n2428 0.00103916
R9376 GND.n2586 GND.n2585 0.00103916
R9377 GND.n2750 GND.n2749 0.00103916
R9378 GND.n7682 GND.n7681 0.00103916
R9379 GND.n3023 GND.n3022 0.00103916
R9380 GND.n3133 GND.n3132 0.00103916
R9381 GND.n1190 GND.n1189 0.00103916
R9382 GND.n3204 GND.n3203 0.00103916
R9383 GND.n5339 GND.n5338 0.00103916
R9384 GND.n5015 GND.n5014 0.00103916
R9385 GND.n3620 GND.n3619 0.00103916
R9386 GND.n4037 GND.n4036 0.00103916
R9387 GND.n3836 GND.n3835 0.00103916
R9388 GND.n4615 GND.n4612 0.00103602
R9389 GND.n4084 GND.n4083 0.00102722
R9390 GND.n1284 GND.n1283 0.00102722
R9391 GND.n3077 GND.n3076 0.00102722
R9392 GND.n3902 GND.n3901 0.00102722
R9393 GND.n5399 GND.n5398 0.00101312
R9394 GND.n2905 GND.n2904 0.00101312
R9395 GND.n2640 GND.n2639 0.00101312
R9396 GND.n2166 GND.n2165 0.00101312
R9397 GND.n1435 GND.n1434 0.00101312
R9398 GND.n2475 GND.n2474 0.00101312
R9399 GND.n2809 GND.n2808 0.00101312
R9400 GND.n7732 GND.n7731 0.00101312
R9401 GND.n5068 GND.n5067 0.00101312
R9402 GND.n3674 GND.n3673 0.00101312
R9403 GND.n3179 GND.n3178 0.00101312
R9404 GND.n3286 GND.n3285 0.00101312
R9405 GND.n3874 GND.n3873 0.00100729
R9406 GND.n3178 GND.n3177 0.00100714
R9407 GND.n3285 GND.n3284 0.00100714
R9408 GND.n5398 GND.n5363 0.00100714
R9409 GND.n2904 GND.n2875 0.00100714
R9410 GND.n2639 GND.n2610 0.00100714
R9411 GND.n2165 GND.n2130 0.00100714
R9412 GND.n1434 GND.n1382 0.00100714
R9413 GND.n2474 GND.n2453 0.00100714
R9414 GND.n2808 GND.n2774 0.00100714
R9415 GND.n7731 GND.n7706 0.00100714
R9416 GND.n5067 GND.n5039 0.00100714
R9417 GND.n3673 GND.n3644 0.00100714
R9418 GND.n4641 GND.n4640 0.00100417
R9419 GND.n3990 GND.n3989 0.001004
R9420 GND.n5292 GND.n5291 0.001004
R9421 GND.n1180 GND.n1178 0.001004
R9422 GND.n5619 GND.n5615 0.001004
R9423 GND.n1341 GND.n1340 0.001004
R9424 GND.n2958 GND.n2956 0.001004
R9425 GND.n2539 GND.n2538 0.001004
R9426 GND.n2059 GND.n2058 0.001004
R9427 GND.n1592 GND.n1587 0.001004
R9428 GND.n4698 GND.n4697 0.00100271
R9429 GND.n7785 GND.n7784 0.00100171
R9430 GND.n6467 GND.n6466 0.00100171
R9431 GND.n6326 GND.n6325 0.00100171
R9432 GND.n6407 GND.n6406 0.00100171
R9433 GND.n7784 GND.n7783 0.00100166
R9434 GND.n6467 GND.n715 0.00100166
R9435 GND.n6326 GND.n6323 0.00100166
R9436 GND.n6406 GND.n6266 0.00100166
R9437 GND.n4737 GND.n4637 0.00100126
R9438 GND.n7377 GND.n7376 0.00100097
R9439 GND.n5911 GND.n5910 0.00100097
R9440 GND.n6042 GND.n6000 0.00100097
R9441 GND.n7284 GND.n7283 0.00100097
R9442 GND.n5663 GND.n5656 0.00100097
R9443 GND.n5793 GND.n5685 0.00100097
R9444 GND.n5752 GND.n5751 0.00100097
R9445 GND.n1456 GND.n1455 0.00100095
R9446 GND.n1040 GND.n1039 0.00100095
R9447 GND.n6548 GND.n6547 0.00100095
R9448 GND.n7559 GND.n7558 0.00100095
R9449 GND.n5096 GND.n5095 0.00100095
R9450 GND.n3307 GND.n3306 0.00100095
R9451 GND.n3462 GND.n3461 0.00100095
R9452 GND.n6802 GND.n6801 0.00100095
R9453 GND.n7125 GND.n7124 0.00100095
R9454 GND.n1862 GND.n1861 0.00100095
R9455 GND.n2197 GND.n2196 0.00100095
R9456 GND.n6956 GND.n6955 0.00100095
R9457 GND.n86 GND.n85 0.00100095
R9458 GND.n4775 GND.n4774 0.00100095
R9459 GND.n7497 GND.n7496 0.00100095
R9460 GND.n7622 GND.n7621 0.00100095
R9461 GND.n6455 GND.n6419 0.00100086
R9462 GND.n7439 GND.n516 0.00100086
R9463 GND.n2383 GND.n2382 0.00100064
R9464 GND.n2704 GND.n2703 0.00100064
R9465 GND.n149 GND.n148 0.00100064
R9466 GND.n4969 GND.n4968 0.00100064
R9467 GND.n3728 GND.n3727 0.00100064
R9468 GND.n3784 GND.n3783 0.00100064
R9469 GND.n5419 GND.n1840 0.00100018
R9470 GND.n5419 GND.n1835 0.00100018
R9471 GND.n5419 GND.n1830 0.00100018
R9472 GND.n5419 GND.n1825 0.00100018
R9473 GND.n5419 GND.n1820 0.00100018
R9474 GND.n5419 GND.n1815 0.00100018
R9475 GND.n5419 GND.n1810 0.00100018
R9476 GND.n5419 GND.n1805 0.00100018
R9477 GND.n5419 GND.n1800 0.00100018
R9478 GND.n5419 GND.n1795 0.00100018
R9479 GND.n5419 GND.n1790 0.00100018
R9480 GND.n5419 GND.n1785 0.00100018
R9481 GND.n5419 GND.n1780 0.00100018
R9482 GND.n5419 GND.n1775 0.00100018
R9483 GND.n4099 GND.n3936 0.00100018
R9484 GND.n7440 GND.n7439 0.00100017
R9485 GND.n6456 GND.n6455 0.00100017
R9486 GND.n5422 GND.n5419 0.00100006
R9487 GND.n5419 GND.n2175 0.00100006
R9488 GND.n5419 GND.n2484 0.00100006
R9489 GND.n5419 GND.n2649 0.00100006
R9490 GND.n5419 GND.n2818 0.00100006
R9491 GND.n5419 GND.n2970 0.00100006
R9492 GND.n5419 GND.n2978 0.00100006
R9493 GND.n5419 GND.n3088 0.00100006
R9494 GND.n5419 GND.n3189 0.00100006
R9495 GND.n5419 GND.n3195 0.00100006
R9496 GND.n5419 GND.n3569 0.00100006
R9497 GND.n5419 GND.n3572 0.00100006
R9498 GND.n5419 GND.n3575 0.00100006
R9499 GND.n5419 GND.n5418 0.00100006
R9500 GND.n4102 GND.n4099 0.00100006
R9501 GND.n4617 GND.n4611 0.00100003
R9502 GND.n3556 GND.n3555 0.00100001
R9503 GND.n1180 GND.n1179 0.00100001
R9504 GND.n5619 GND.n5618 0.00100001
R9505 GND.n2958 GND.n2957 0.00100001
R9506 GND.n1592 GND.n1591 0.00100001
R9507 GND.n4099 GND.n4094 0.001
R9508 GND.n6496 GND.n6495 0.001
R9509 GND.n7444 GND.n7443 0.001
R9510 GND.n6292 GND.n6291 0.001
R9511 GND.n4625 GND.n4624 0.000966399
R9512 GND.n4624 GND.n4623 0.000959101
R9513 GND.n4623 GND.n4622 0.000959101
R9514 GND.n4007 GND.n4002 0.000943262
R9515 GND.n1409 GND.n1402 0.000943262
R9516 GND.n2076 GND.n2071 0.000943262
R9517 GND.n2398 GND.n2393 0.000943262
R9518 GND.n2556 GND.n2551 0.000943262
R9519 GND.n2719 GND.n2714 0.000943262
R9520 GND.n2837 GND.n2827 0.000943262
R9521 GND.n7658 GND.n158 0.000943262
R9522 GND.n2993 GND.n2988 0.000943262
R9523 GND.n3102 GND.n3097 0.000943262
R9524 GND.n5309 GND.n5304 0.000943262
R9525 GND.n4984 GND.n4979 0.000943262
R9526 GND.n3590 GND.n3585 0.000943262
R9527 GND.n3804 GND.n3793 0.000943262
R9528 GND.n3216 GND.n3211 0.000943262
R9529 GND.n1203 GND.n1198 0.000943262
R9530 GND.n868 GND.n866 0.000898936
R9531 GND.n884 GND.n720 0.000898936
R9532 GND.n4246 GND.n4245 0.000864406
R9533 GND.n4252 GND.n4251 0.000864406
R9534 GND.n4247 GND.n4246 0.000858717
R9535 GND.n4249 GND.n4247 0.000858717
R9536 GND.n4251 GND.n4250 0.000858717
R9537 GND.n4250 GND.n4249 0.000858717
R9538 GND.n4188 GND.n4187 0.000858717
R9539 GND.n4187 GND.n4186 0.000858717
R9540 GND.n4193 GND.n4192 0.000858717
R9541 GND.n4643 GND.n4642 0.000840211
R9542 GND.n4737 GND.n4643 0.000840211
R9543 GND.n5424 GND.n5423 0.000826763
R9544 GND.n2172 GND.n2171 0.000826763
R9545 GND.n2481 GND.n2480 0.000826763
R9546 GND.n2646 GND.n2645 0.000826763
R9547 GND.n2815 GND.n2814 0.000826763
R9548 GND.n2967 GND.n2966 0.000826763
R9549 GND.n2975 GND.n2974 0.000826763
R9550 GND.n3085 GND.n3084 0.000826763
R9551 GND.n3186 GND.n3185 0.000826763
R9552 GND.n3192 GND.n3191 0.000826763
R9553 GND.n3566 GND.n3565 0.000826763
R9554 GND.n5402 GND.n5401 0.000826763
R9555 GND.n5071 GND.n5070 0.000826763
R9556 GND.n5415 GND.n5414 0.000826763
R9557 GND.n4104 GND.n4103 0.000826763
R9558 GND.n4091 GND.n4090 0.000826763
R9559 GND.n4699 GND.n4698 0.000801918
R9560 GND.n4700 GND.n4699 0.000801918
R9561 GND.n4736 GND.n4735 0.000801918
R9562 GND.n4737 GND.n4736 0.000801918
R9563 GND.n4729 GND.n4728 0.000801918
R9564 GND.n4737 GND.n4729 0.000801918
R9565 GND.n4725 GND.n4724 0.000801918
R9566 GND.n4737 GND.n4725 0.000801918
R9567 GND.n4716 GND.n4715 0.000801918
R9568 GND.n4737 GND.n4716 0.000801918
R9569 GND.n4702 GND.n4701 0.000801918
R9570 GND.n4701 GND.n4700 0.000801918
R9571 GND.n4708 GND.n4707 0.000801918
R9572 GND.n4714 GND.n4713 0.000801918
R9573 GND.n4737 GND.n4714 0.000801918
R9574 GND.n4737 GND.n4682 0.000801918
R9575 GND.n4679 GND.n4678 0.000801918
R9576 GND.n4737 GND.n4679 0.000801918
R9577 GND.n4667 GND.n4666 0.000801918
R9578 GND.n4737 GND.n4667 0.000801918
R9579 GND.n4695 GND.n4694 0.000801918
R9580 GND.n4700 GND.n4695 0.000801918
R9581 GND.n4659 GND.n4658 0.000801918
R9582 GND.n4737 GND.n4659 0.000801918
R9583 GND.n4651 GND.n4650 0.000801918
R9584 GND.n4737 GND.n4651 0.000801918
R9585 GND.n4691 GND.n4690 0.000801918
R9586 GND.n4700 GND.n4691 0.000801918
R9587 GND.n4631 GND.n4630 0.000801918
R9588 GND.n4737 GND.n4631 0.000801918
R9589 GND.n1363 GND.n1362 0.000756235
R9590 GND.n1362 GND.n1361 0.000756235
R9591 GND.n2111 GND.n2110 0.000756235
R9592 GND.n2110 GND.n2109 0.000756235
R9593 GND.n2434 GND.n2433 0.000756235
R9594 GND.n2433 GND.n2432 0.000756235
R9595 GND.n2591 GND.n2590 0.000756235
R9596 GND.n2590 GND.n2589 0.000756235
R9597 GND.n2755 GND.n2754 0.000756235
R9598 GND.n2754 GND.n2753 0.000756235
R9599 GND.n2886 GND.n2885 0.000756235
R9600 GND.n2887 GND.n2886 0.000756235
R9601 GND.n7687 GND.n7686 0.000756235
R9602 GND.n7686 GND.n7685 0.000756235
R9603 GND.n3057 GND.n3056 0.000756235
R9604 GND.n3056 GND.n3055 0.000756235
R9605 GND.n3158 GND.n3157 0.000756235
R9606 GND.n3157 GND.n3156 0.000756235
R9607 GND.n1264 GND.n1263 0.000756235
R9608 GND.n1263 GND.n1262 0.000756235
R9609 GND.n3265 GND.n3264 0.000756235
R9610 GND.n3264 GND.n3263 0.000756235
R9611 GND.n5344 GND.n5343 0.000756235
R9612 GND.n5343 GND.n5342 0.000756235
R9613 GND.n5020 GND.n5019 0.000756235
R9614 GND.n5019 GND.n5018 0.000756235
R9615 GND.n3625 GND.n3624 0.000756235
R9616 GND.n3624 GND.n3623 0.000756235
R9617 GND.n4064 GND.n4063 0.000756235
R9618 GND.n4063 GND.n4062 0.000756235
R9619 GND.n3877 GND.n3876 0.000756235
R9620 GND.n3876 GND.n3875 0.000756235
R9621 GND.n4625 GND.n4619 0.000714408
R9622 GND.n736 GND.n734 0.000632979
R9623 GND.n6132 GND.n5849 0.000632979
R9624 GND.n7433 GND.n553 0.000632979
R9625 GND.n4619 GND.n4617 0.000607204
R9626 GND.n4605 GND.n4604 0.000567786
R9627 GND.n6323 GND.n6293 0.000560793
R9628 GND.n715 GND.n677 0.000560793
R9629 GND.n7783 GND.n7753 0.000560793
R9630 GND.n6408 GND.n6407 0.000557763
R9631 GND.n6325 GND.n6324 0.000557763
R9632 GND.n6466 GND.n6465 0.000557763
R9633 GND.n7786 GND.n7785 0.000557763
R9634 GND.n4227 GND.n4226 0.000557678
R9635 GND.n1532 GND.n1531 0.000544755
R9636 GND.n5632 GND.n5631 0.000544755
R9637 GND.n6508 GND.n6507 0.000544755
R9638 GND.n7519 GND.n7518 0.000544755
R9639 GND.n5219 GND.n5218 0.000544755
R9640 GND.n3484 GND.n3483 0.000544755
R9641 GND.n5450 GND.n5449 0.000544755
R9642 GND.n6815 GND.n6814 0.000544755
R9643 GND.n7085 GND.n7084 0.000544755
R9644 GND.n1986 GND.n1985 0.000544755
R9645 GND.n2309 GND.n2308 0.000544755
R9646 GND.n6969 GND.n6968 0.000544755
R9647 GND.n7743 GND.n7742 0.000544755
R9648 GND.n4895 GND.n4894 0.000544755
R9649 GND.n7457 GND.n7456 0.000544755
R9650 GND.n7582 GND.n7581 0.000544755
R9651 GND.n4237 GND.n4236 0.000538452
R9652 GND.n4191 GND.n4190 0.000537082
R9653 GND.n1489 GND.n1488 0.000530553
R9654 GND.n1906 GND.n1905 0.000530553
R9655 GND.n2229 GND.n2228 0.000530553
R9656 GND.n7155 GND.n7154 0.000530553
R9657 GND.n6989 GND.n6988 0.000530553
R9658 GND.n6835 GND.n6834 0.000530553
R9659 GND.n6681 GND.n6680 0.000530553
R9660 GND.n6611 GND.n6610 0.000530553
R9661 GND.n5508 GND.n5507 0.000530553
R9662 GND.n1074 GND.n1073 0.000530553
R9663 GND.n3382 GND.n3381 0.000530553
R9664 GND.n5142 GND.n5141 0.000530553
R9665 GND.n4818 GND.n4817 0.000530553
R9666 GND.n444 GND.n443 0.000530553
R9667 GND.n375 GND.n374 0.000530553
R9668 GND.n264 GND.n263 0.000530553
R9669 GND.n6381 GND.n6380 0.000528881
R9670 GND.n6380 GND.n6379 0.000528881
R9671 GND.n6383 GND.n6382 0.000528881
R9672 GND.n6471 GND.n6470 0.000528881
R9673 GND.n6470 GND.n6469 0.000528881
R9674 GND.n6473 GND.n6472 0.000528881
R9675 GND.n1510 GND.n1509 0.00052846
R9676 GND.n1932 GND.n1931 0.00052846
R9677 GND.n2255 GND.n2254 0.00052846
R9678 GND.n7181 GND.n7180 0.00052846
R9679 GND.n7015 GND.n7014 0.00052846
R9680 GND.n6861 GND.n6860 0.00052846
R9681 GND.n6707 GND.n6706 0.00052846
R9682 GND.n6637 GND.n6636 0.00052846
R9683 GND.n5534 GND.n5533 0.00052846
R9684 GND.n1100 GND.n1099 0.00052846
R9685 GND.n3408 GND.n3407 0.00052846
R9686 GND.n5168 GND.n5167 0.00052846
R9687 GND.n4844 GND.n4843 0.00052846
R9688 GND.n470 GND.n469 0.00052846
R9689 GND.n401 GND.n400 0.00052846
R9690 GND.n290 GND.n289 0.00052846
R9691 GND.n1050 GND.n1049 0.00052846
R9692 GND.n5477 GND.n5476 0.00052846
R9693 GND.n233 GND.n232 0.00052846
R9694 GND.n4863 GND.n4862 0.00052846
R9695 GND.n5187 GND.n5186 0.00052846
R9696 GND.n3360 GND.n3359 0.00052846
R9697 GND.n6738 GND.n6737 0.00052846
R9698 GND.n7046 GND.n7045 0.00052846
R9699 GND.n2277 GND.n2276 0.00052846
R9700 GND.n7207 GND.n7206 0.00052846
R9701 GND.n6892 GND.n6891 0.00052846
R9702 GND.n6580 GND.n6579 0.00052846
R9703 GND.n492 GND.n491 0.00052846
R9704 GND.n344 GND.n343 0.00052846
R9705 GND.n7641 GND.n7640 0.00052846
R9706 GND.n1954 GND.n1953 0.00052846
R9707 GND.n4256 GND.n4255 0.000526656
R9708 GND.n1962 GND.n1961 0.0005264
R9709 GND.n1107 GND.n1106 0.0005264
R9710 GND.n5541 GND.n5540 0.0005264
R9711 GND.n297 GND.n296 0.0005264
R9712 GND.n4871 GND.n4870 0.0005264
R9713 GND.n5195 GND.n5194 0.0005264
R9714 GND.n3415 GND.n3414 0.0005264
R9715 GND.n6746 GND.n6745 0.0005264
R9716 GND.n7054 GND.n7053 0.0005264
R9717 GND.n2285 GND.n2284 0.0005264
R9718 GND.n7215 GND.n7214 0.0005264
R9719 GND.n6900 GND.n6899 0.0005264
R9720 GND.n6644 GND.n6643 0.0005264
R9721 GND.n500 GND.n499 0.0005264
R9722 GND.n408 GND.n407 0.0005264
R9723 GND.n7649 GND.n7648 0.0005264
R9724 GND.n4608 GND.n4607 0.000525991
R9725 GND.n4198 GND.n4197 0.000524722
R9726 GND.n4746 GND.n4745 0.000523819
R9727 GND.n4750 GND.n4749 0.000523819
R9728 GND.n4741 GND.n4740 0.000523819
R9729 GND.t799 GND.n4747 0.000523446
R9730 GND.n4749 GND.n4748 0.000523446
R9731 GND.n4748 GND.t799 0.000523446
R9732 GND.n4747 GND.n4746 0.000523446
R9733 GND.n4742 GND.n4741 0.000523446
R9734 GND.t799 GND.n4742 0.000523446
R9735 GND.n4212 GND.n4211 0.000517138
R9736 GND.n5490 GND.n5489 0.000512627
R9737 GND.n6593 GND.n6592 0.000512627
R9738 GND.n357 GND.n356 0.000512627
R9739 GND.n4853 GND.n4850 0.000512627
R9740 GND.n5177 GND.n5174 0.000512627
R9741 GND.n3350 GND.n3349 0.000512627
R9742 GND.n6728 GND.n6715 0.000512627
R9743 GND.n7036 GND.n7023 0.000512627
R9744 GND.n2267 GND.n2261 0.000512627
R9745 GND.n7197 GND.n7189 0.000512627
R9746 GND.n6882 GND.n6869 0.000512627
R9747 GND.n6570 GND.n6567 0.000512627
R9748 GND.n482 GND.n476 0.000512627
R9749 GND.n334 GND.n331 0.000512627
R9750 GND.n246 GND.n245 0.000512627
R9751 GND.n1944 GND.n1943 0.000512627
R9752 GND.n1483 GND.n1482 0.000512369
R9753 GND.n1900 GND.n1899 0.000512369
R9754 GND.n2223 GND.n2222 0.000512369
R9755 GND.n7025 GND.n7024 0.000512369
R9756 GND.n6871 GND.n6870 0.000512369
R9757 GND.n6717 GND.n6716 0.000512369
R9758 GND.n6675 GND.n6674 0.000512369
R9759 GND.n6605 GND.n6604 0.000512369
R9760 GND.n5502 GND.n5501 0.000512369
R9761 GND.n1068 GND.n1067 0.000512369
R9762 GND.n3376 GND.n3375 0.000512369
R9763 GND.n5136 GND.n5135 0.000512369
R9764 GND.n4812 GND.n4811 0.000512369
R9765 GND.n438 GND.n437 0.000512369
R9766 GND.n369 GND.n368 0.000512369
R9767 GND.n258 GND.n257 0.000512369
R9768 GND.n4650 GND.n4649 0.000508571
R9769 GND.n4658 GND.n4657 0.000508571
R9770 GND.n4666 GND.n4665 0.000508571
R9771 GND.n4678 GND.n4677 0.000508571
R9772 GND.n4674 GND.n4673 0.000508571
R9773 GND.n4713 GND.n4712 0.000508571
R9774 GND.n4709 GND.n4708 0.000508571
R9775 GND.n4724 GND.n4723 0.000508571
R9776 GND.n4728 GND.n4727 0.000508571
R9777 GND.n4735 GND.n4734 0.000508571
R9778 GND.n4630 GND.n4629 0.000508571
R9779 GND.n1879 GND.n1878 0.000507826
R9780 GND.n2205 GND.n2204 0.000507826
R9781 GND.n7136 GND.n7135 0.000507826
R9782 GND.n7068 GND.n7067 0.000507826
R9783 GND.n6914 GND.n6913 0.000507826
R9784 GND.n6760 GND.n6759 0.000507826
R9785 GND.n6561 GND.n6560 0.000507826
R9786 GND.n5548 GND.n5547 0.000507826
R9787 GND.n3426 GND.n3425 0.000507826
R9788 GND.n3343 GND.n3342 0.000507826
R9789 GND.n5113 GND.n5112 0.000507826
R9790 GND.n4792 GND.n4791 0.000507826
R9791 GND.n415 GND.n414 0.000507826
R9792 GND.n325 GND.n324 0.000507826
R9793 GND.n223 GND.n222 0.000507826
R9794 GND.n195 GND.n194 0.000507826
R9795 GND.n1474 GND.n1473 0.000507826
R9796 GND.n1891 GND.n1890 0.000507826
R9797 GND.n2216 GND.n2215 0.000507826
R9798 GND.n7147 GND.n7146 0.000507826
R9799 GND.n7064 GND.n7063 0.000507826
R9800 GND.n6910 GND.n6909 0.000507826
R9801 GND.n6756 GND.n6755 0.000507826
R9802 GND.n6557 GND.n6556 0.000507826
R9803 GND.n5559 GND.n5558 0.000507826
R9804 GND.n3437 GND.n3436 0.000507826
R9805 GND.n3325 GND.n3324 0.000507826
R9806 GND.n5124 GND.n5123 0.000507826
R9807 GND.n4803 GND.n4802 0.000507826
R9808 GND.n426 GND.n425 0.000507826
R9809 GND.n321 GND.n320 0.000507826
R9810 GND.n219 GND.n218 0.000507826
R9811 GND.n3054 GND.n3053 0.000507291
R9812 GND.n1261 GND.n1260 0.000507291
R9813 GND.n3672 GND.n3671 0.000507291
R9814 GND.n4061 GND.n4060 0.000507291
R9815 GND.n5912 GND.n5911 0.000506774
R9816 GND.n5914 GND.n5913 0.000506774
R9817 GND.n6117 GND.n6000 0.000506774
R9818 GND.n6116 GND.n6115 0.000506774
R9819 GND.n6119 GND.n6118 0.000506774
R9820 GND.n5999 GND.n5998 0.000506774
R9821 GND.n739 GND.n738 0.000506774
R9822 GND.n833 GND.n832 0.000506774
R9823 GND.n928 GND.n927 0.000506774
R9824 GND.n1003 GND.n1002 0.000506774
R9825 GND.n926 GND.n925 0.000506774
R9826 GND.n835 GND.n834 0.000506774
R9827 GND.n5693 GND.n5685 0.000506774
R9828 GND.n5753 GND.n5752 0.000506774
R9829 GND.n5656 GND.n5655 0.000506774
R9830 GND.n5692 GND.n5683 0.000506774
R9831 GND.n5755 GND.n5754 0.000506774
R9832 GND.n6226 GND.n6225 0.000506774
R9833 GND.n6160 GND.n6159 0.000506774
R9834 GND.n7287 GND.n7286 0.000506774
R9835 GND.n7376 GND.n7375 0.000506774
R9836 GND.n7797 GND.n7796 0.000506774
R9837 GND.n7374 GND.n556 0.000506774
R9838 GND.n7372 GND.n7371 0.000506774
R9839 GND.n7285 GND.n7284 0.000506774
R9840 GND.n1417 GND.n1416 0.000505544
R9841 GND.n2084 GND.n2083 0.000505544
R9842 GND.n2406 GND.n2405 0.000505544
R9843 GND.n2564 GND.n2563 0.000505544
R9844 GND.n2727 GND.n2726 0.000505544
R9845 GND.n7656 GND.n7655 0.000505544
R9846 GND.n3001 GND.n3000 0.000505544
R9847 GND.n3110 GND.n3109 0.000505544
R9848 GND.n5317 GND.n5316 0.000505544
R9849 GND.n4992 GND.n4991 0.000505544
R9850 GND.n3598 GND.n3597 0.000505544
R9851 GND.n4015 GND.n4014 0.000505544
R9852 GND.n3802 GND.n3801 0.000505544
R9853 GND.n3224 GND.n3223 0.000505544
R9854 GND.n2835 GND.n2834 0.000505544
R9855 GND.n1211 GND.n1210 0.000505544
R9856 GND.n1457 GND.n1456 0.000504863
R9857 GND.n5566 GND.n1040 0.000504863
R9858 GND.n6549 GND.n6548 0.000504863
R9859 GND.n7560 GND.n7559 0.000504863
R9860 GND.n5097 GND.n5096 0.000504863
R9861 GND.n3332 GND.n3307 0.000504863
R9862 GND.n3463 GND.n3462 0.000504863
R9863 GND.n6804 GND.n6802 0.000504863
R9864 GND.n7126 GND.n7125 0.000504863
R9865 GND.n1863 GND.n1862 0.000504863
R9866 GND.n2198 GND.n2197 0.000504863
R9867 GND.n6958 GND.n6956 0.000504863
R9868 GND.n87 GND.n86 0.000504863
R9869 GND.n4776 GND.n4775 0.000504863
R9870 GND.n7498 GND.n7497 0.000504863
R9871 GND.n7623 GND.n7622 0.000504863
R9872 GND.n4661 GND.n4660 0.000504378
R9873 GND.n4703 GND.n4702 0.000504346
R9874 GND.n4731 GND.n4730 0.00050424
R9875 GND.n4733 GND.n4732 0.00050424
R9876 GND.n4705 GND.n4704 0.00050424
R9877 GND.n4711 GND.n4710 0.00050424
R9878 GND.n4676 GND.n4675 0.00050424
R9879 GND.n4654 GND.n4653 0.00050424
R9880 GND.n4656 GND.n4655 0.00050424
R9881 GND.n4645 GND.n4644 0.00050424
R9882 GND.n4722 GND.n4721 0.000504176
R9883 GND.n4720 GND.n4719 0.000504112
R9884 GND.n4685 GND.n4684 0.000504112
R9885 GND.n4670 GND.n4669 0.000504112
R9886 GND.n4664 GND.n4663 0.000504112
R9887 GND.n4648 GND.n4647 0.000504112
R9888 GND.n3941 GND.n3940 0.000504005
R9889 GND.n5243 GND.n5242 0.000504005
R9890 GND.n3557 GND.n3556 0.000504005
R9891 GND.n1292 GND.n1291 0.000504005
R9892 GND.n2490 GND.n2489 0.000504005
R9893 GND.n2010 GND.n2009 0.000504005
R9894 GND.n1591 GND.n1590 0.000504005
R9895 GND.n2381 GND.n2380 0.000504005
R9896 GND.n2702 GND.n2701 0.000504005
R9897 GND.n147 GND.n146 0.000504005
R9898 GND.n3726 GND.n3725 0.000504005
R9899 GND.n3782 GND.n3781 0.000504005
R9900 GND.n4619 GND.n4618 0.00050212
R9901 GND.n3992 GND.n3991 0.000501449
R9902 GND.n5294 GND.n5293 0.000501449
R9903 GND.n3559 GND.n3558 0.000501449
R9904 GND.n5439 GND.n1181 0.000501449
R9905 GND.n2960 GND.n2959 0.000501449
R9906 GND.n2541 GND.n2540 0.000501449
R9907 GND.n2061 GND.n2060 0.000501449
R9908 GND.n2384 GND.n2383 0.000501449
R9909 GND.n2705 GND.n2704 0.000501449
R9910 GND.n7734 GND.n149 0.000501449
R9911 GND.n4970 GND.n4969 0.000501449
R9912 GND.n3729 GND.n3728 0.000501449
R9913 GND.n3785 GND.n3784 0.000501449
R9914 GND.n1343 GND.n1342 0.000501449
R9915 GND.n5621 GND.n5620 0.000501449
R9916 GND.n1594 GND.n1593 0.000501449
R9917 GND.n1549 GND.n1548 0.000501292
R9918 GND.n1548 GND.n1547 0.000501292
R9919 GND.n5630 GND.n5625 0.000501292
R9920 GND.n5630 GND.n5629 0.000501292
R9921 GND.n6525 GND.n6524 0.000501292
R9922 GND.n6524 GND.n6523 0.000501292
R9923 GND.n7536 GND.n7535 0.000501292
R9924 GND.n7535 GND.n7534 0.000501292
R9925 GND.n5236 GND.n5235 0.000501292
R9926 GND.n5235 GND.n5234 0.000501292
R9927 GND.n3501 GND.n3500 0.000501292
R9928 GND.n3500 GND.n3499 0.000501292
R9929 GND.n5448 GND.n5443 0.000501292
R9930 GND.n5448 GND.n5447 0.000501292
R9931 GND.n6813 GND.n6808 0.000501292
R9932 GND.n6813 GND.n6812 0.000501292
R9933 GND.n7102 GND.n7101 0.000501292
R9934 GND.n7101 GND.n7100 0.000501292
R9935 GND.n2003 GND.n2002 0.000501292
R9936 GND.n2002 GND.n2001 0.000501292
R9937 GND.n2326 GND.n2325 0.000501292
R9938 GND.n2325 GND.n2324 0.000501292
R9939 GND.n6967 GND.n6962 0.000501292
R9940 GND.n6967 GND.n6966 0.000501292
R9941 GND.n7739 GND.n7738 0.000501292
R9942 GND.n7740 GND.n7739 0.000501292
R9943 GND.n4912 GND.n4911 0.000501292
R9944 GND.n4911 GND.n4910 0.000501292
R9945 GND.n7474 GND.n7473 0.000501292
R9946 GND.n7473 GND.n7472 0.000501292
R9947 GND.n7599 GND.n7598 0.000501292
R9948 GND.n7598 GND.n7597 0.000501292
R9949 GND.n4189 GND.n4188 0.00050117
R9950 GND.n4194 GND.n4193 0.00050117
R9951 GND.n5915 GND.n5914 0.00050097
R9952 GND.n6115 GND.n6114 0.00050097
R9953 GND.n6120 GND.n6119 0.00050097
R9954 GND.n5998 GND.n5997 0.00050097
R9955 GND.n740 GND.n739 0.00050097
R9956 GND.n832 GND.n831 0.00050097
R9957 GND.n929 GND.n928 0.00050097
R9958 GND.n1002 GND.n1001 0.00050097
R9959 GND.n925 GND.n924 0.00050097
R9960 GND.n836 GND.n835 0.00050097
R9961 GND.n5756 GND.n5755 0.00050097
R9962 GND.n6225 GND.n6224 0.00050097
R9963 GND.n6161 GND.n6160 0.00050097
R9964 GND.n7288 GND.n7287 0.00050097
R9965 GND.n7798 GND.n7797 0.00050097
R9966 GND.n7421 GND.n556 0.00050097
R9967 GND.n7371 GND.n7370 0.00050097
R9968 GND.n5826 GND.n5683 0.00050097
R9969 GND.n1416 GND.n1415 0.000500915
R9970 GND.n2083 GND.n2082 0.000500915
R9971 GND.n2405 GND.n2404 0.000500915
R9972 GND.n2563 GND.n2562 0.000500915
R9973 GND.n2726 GND.n2725 0.000500915
R9974 GND.n7657 GND.n7656 0.000500915
R9975 GND.n3000 GND.n2999 0.000500915
R9976 GND.n3109 GND.n3108 0.000500915
R9977 GND.n5316 GND.n5315 0.000500915
R9978 GND.n4991 GND.n4990 0.000500915
R9979 GND.n3597 GND.n3596 0.000500915
R9980 GND.n4014 GND.n4013 0.000500915
R9981 GND.n3803 GND.n3802 0.000500915
R9982 GND.n3223 GND.n3222 0.000500915
R9983 GND.n2836 GND.n2835 0.000500915
R9984 GND.n1210 GND.n1209 0.000500915
R9985 GND.n4239 GND.n4238 0.000500552
R9986 GND.n4254 GND.n4253 0.000500539
R9987 GND.n3191 GND.n3190 0.000500526
R9988 GND.n3084 GND.n3083 0.000500526
R9989 GND.n5425 GND.n5424 0.000500526
R9990 GND.n2171 GND.n2170 0.000500526
R9991 GND.n2480 GND.n2479 0.000500526
R9992 GND.n2645 GND.n2644 0.000500526
R9993 GND.n2814 GND.n2813 0.000500526
R9994 GND.n2966 GND.n2965 0.000500526
R9995 GND.n2974 GND.n2973 0.000500526
R9996 GND.n3185 GND.n3184 0.000500526
R9997 GND.n3565 GND.n3564 0.000500526
R9998 GND.n5403 GND.n5402 0.000500526
R9999 GND.n5072 GND.n5071 0.000500526
R10000 GND.n5414 GND.n5413 0.000500526
R10001 GND.n4090 GND.n4089 0.000500526
R10002 GND.n4105 GND.n4104 0.000500526
R10003 GND.n4196 GND.n4195 0.000500355
R10004 GND.n4112 GND.n4111 0.000500347
R10005 GND.n4007 GND.n4006 0.000500286
R10006 GND.n1409 GND.n1408 0.000500286
R10007 GND.n2076 GND.n2075 0.000500286
R10008 GND.n2398 GND.n2397 0.000500286
R10009 GND.n2556 GND.n2555 0.000500286
R10010 GND.n2719 GND.n2718 0.000500286
R10011 GND.n2839 GND.n2837 0.000500286
R10012 GND.n7660 GND.n7658 0.000500286
R10013 GND.n2993 GND.n2992 0.000500286
R10014 GND.n3102 GND.n3101 0.000500286
R10015 GND.n5309 GND.n5308 0.000500286
R10016 GND.n4984 GND.n4983 0.000500286
R10017 GND.n3590 GND.n3589 0.000500286
R10018 GND.n3806 GND.n3804 0.000500286
R10019 GND.n3216 GND.n3215 0.000500286
R10020 GND.n1203 GND.n1202 0.000500286
R10021 GND.n4440 GND.n4439 0.000500199
R10022 GND.n6136 GND.n6135 0.00050016
R10023 GND.n4448 GND.n4447 0.000500107
R10024 GND.n2169 GND.n2168 0.000500059
R10025 GND.n2478 GND.n2477 0.000500059
R10026 GND.n2643 GND.n2642 0.000500059
R10027 GND.n2812 GND.n2811 0.000500059
R10028 GND.n2964 GND.n2962 0.000500059
R10029 GND.n2972 GND.n150 0.000500059
R10030 GND.n5406 GND.n5405 0.000500059
R10031 GND.n5075 GND.n5074 0.000500059
R10032 GND.n5412 GND.n5410 0.000500059
R10033 GND.n4088 GND.n4087 0.000500059
R10034 GND.n4108 GND.n4107 0.000500059
R10035 GND.n3563 GND.n3561 0.000500059
R10036 GND.n5437 GND.n1287 0.000500059
R10037 GND.n3183 GND.n3181 0.000500059
R10038 GND.n3082 GND.n3080 0.000500059
R10039 GND.n5428 GND.n5427 0.000500059
R10040 GND.n4744 GND.n4743 0.000500053
R10041 GND.n4739 GND.n4738 0.000500023
R10042 GND.n4672 GND.n4671 0.00050002
R10043 VDD.n1970 VDD.n1931 8089.41
R10044 VDD.n1951 VDD.n1949 8089.41
R10045 VDD.n1954 VDD.n1948 6801.18
R10046 VDD.n1913 VDD.n1895 2565.88
R10047 VDD.n1913 VDD.n1896 2565.88
R10048 VDD.n1878 VDD.n1823 2565.88
R10049 VDD.n1859 VDD.n1848 2565.88
R10050 VDD.n1864 VDD.n1848 2565.88
R10051 VDD.n2180 VDD.n2169 2565.88
R10052 VDD.n2185 VDD.n2169 2565.88
R10053 VDD.n2199 VDD.n2144 2565.88
R10054 VDD.n2234 VDD.n2216 2565.88
R10055 VDD.n2234 VDD.n2217 2565.88
R10056 VDD.n2438 VDD.n2427 2565.88
R10057 VDD.n2443 VDD.n2427 2565.88
R10058 VDD.n2457 VDD.n2402 2565.88
R10059 VDD.n2492 VDD.n2474 2565.88
R10060 VDD.n2492 VDD.n2475 2565.88
R10061 VDD.n2696 VDD.n2685 2565.88
R10062 VDD.n2701 VDD.n2685 2565.88
R10063 VDD.n2715 VDD.n2660 2565.88
R10064 VDD.n2750 VDD.n2732 2565.88
R10065 VDD.n2750 VDD.n2733 2565.88
R10066 VDD.n2954 VDD.n2943 2565.88
R10067 VDD.n2959 VDD.n2943 2565.88
R10068 VDD.n2973 VDD.n2918 2565.88
R10069 VDD.n3008 VDD.n2990 2565.88
R10070 VDD.n3008 VDD.n2991 2565.88
R10071 VDD.n3212 VDD.n3201 2565.88
R10072 VDD.n3217 VDD.n3201 2565.88
R10073 VDD.n3231 VDD.n3176 2565.88
R10074 VDD.n3266 VDD.n3248 2565.88
R10075 VDD.n3266 VDD.n3249 2565.88
R10076 VDD.n3470 VDD.n3459 2565.88
R10077 VDD.n3475 VDD.n3459 2565.88
R10078 VDD.n3489 VDD.n3434 2565.88
R10079 VDD.n3524 VDD.n3506 2565.88
R10080 VDD.n3524 VDD.n3507 2565.88
R10081 VDD.n5790 VDD.n5779 2565.88
R10082 VDD.n5795 VDD.n5779 2565.88
R10083 VDD.n5809 VDD.n5754 2565.88
R10084 VDD.n5844 VDD.n5826 2565.88
R10085 VDD.n5844 VDD.n5827 2565.88
R10086 VDD.n5536 VDD.n5525 2565.88
R10087 VDD.n5541 VDD.n5525 2565.88
R10088 VDD.n5555 VDD.n5500 2565.88
R10089 VDD.n5590 VDD.n5572 2565.88
R10090 VDD.n5590 VDD.n5573 2565.88
R10091 VDD.n3728 VDD.n3717 2565.88
R10092 VDD.n3733 VDD.n3717 2565.88
R10093 VDD.n3747 VDD.n3692 2565.88
R10094 VDD.n3782 VDD.n3764 2565.88
R10095 VDD.n3782 VDD.n3765 2565.88
R10096 VDD.n3986 VDD.n3975 2565.88
R10097 VDD.n3991 VDD.n3975 2565.88
R10098 VDD.n4005 VDD.n3950 2565.88
R10099 VDD.n4040 VDD.n4022 2565.88
R10100 VDD.n4040 VDD.n4023 2565.88
R10101 VDD.n4244 VDD.n4233 2565.88
R10102 VDD.n4249 VDD.n4233 2565.88
R10103 VDD.n4263 VDD.n4208 2565.88
R10104 VDD.n4298 VDD.n4280 2565.88
R10105 VDD.n4298 VDD.n4281 2565.88
R10106 VDD.n4502 VDD.n4491 2565.88
R10107 VDD.n4507 VDD.n4491 2565.88
R10108 VDD.n4521 VDD.n4466 2565.88
R10109 VDD.n4556 VDD.n4538 2565.88
R10110 VDD.n4556 VDD.n4539 2565.88
R10111 VDD.n4760 VDD.n4749 2565.88
R10112 VDD.n4765 VDD.n4749 2565.88
R10113 VDD.n4779 VDD.n4724 2565.88
R10114 VDD.n4814 VDD.n4796 2565.88
R10115 VDD.n4814 VDD.n4797 2565.88
R10116 VDD.n5018 VDD.n5007 2565.88
R10117 VDD.n5023 VDD.n5007 2565.88
R10118 VDD.n5037 VDD.n4982 2565.88
R10119 VDD.n5072 VDD.n5054 2565.88
R10120 VDD.n5072 VDD.n5055 2565.88
R10121 VDD.n5276 VDD.n5265 2565.88
R10122 VDD.n5281 VDD.n5265 2565.88
R10123 VDD.n5295 VDD.n5240 2565.88
R10124 VDD.n5330 VDD.n5312 2565.88
R10125 VDD.n5330 VDD.n5313 2565.88
R10126 VDD.n1744 VDD.n1713 2082.55
R10127 VDD.n2093 VDD.n2062 2082.55
R10128 VDD.n2323 VDD.n2292 2082.55
R10129 VDD.n2581 VDD.n2550 2082.55
R10130 VDD.n2839 VDD.n2808 2082.55
R10131 VDD.n3097 VDD.n3066 2082.55
R10132 VDD.n3355 VDD.n3324 2082.55
R10133 VDD.n5678 VDD.n5647 2082.55
R10134 VDD.n5424 VDD.n5393 2082.55
R10135 VDD.n3613 VDD.n3582 2082.55
R10136 VDD.n3871 VDD.n3840 2082.55
R10137 VDD.n4129 VDD.n4098 2082.55
R10138 VDD.n4387 VDD.n4356 2082.55
R10139 VDD.n4645 VDD.n4614 2082.55
R10140 VDD.n4903 VDD.n4872 2082.55
R10141 VDD.n5161 VDD.n5130 2082.55
R10142 VDD.n1694 VDD.n1674 2080.64
R10143 VDD.n2043 VDD.n2023 2080.64
R10144 VDD.n2273 VDD.n2253 2080.64
R10145 VDD.n2531 VDD.n2511 2080.64
R10146 VDD.n2789 VDD.n2769 2080.64
R10147 VDD.n3047 VDD.n3027 2080.64
R10148 VDD.n3305 VDD.n3285 2080.64
R10149 VDD.n5628 VDD.n5608 2080.64
R10150 VDD.n5374 VDD.n5354 2080.64
R10151 VDD.n3563 VDD.n3543 2080.64
R10152 VDD.n3821 VDD.n3801 2080.64
R10153 VDD.n4079 VDD.n4059 2080.64
R10154 VDD.n4337 VDD.n4317 2080.64
R10155 VDD.n4595 VDD.n4575 2080.64
R10156 VDD.n4853 VDD.n4833 2080.64
R10157 VDD.n5111 VDD.n5091 2080.64
R10158 VDD.n1742 VDD.n1712 2015.29
R10159 VDD.n1698 VDD.n1678 2015.29
R10160 VDD.n2091 VDD.n2061 2015.29
R10161 VDD.n2047 VDD.n2027 2015.29
R10162 VDD.n2321 VDD.n2291 2015.29
R10163 VDD.n2277 VDD.n2257 2015.29
R10164 VDD.n2579 VDD.n2549 2015.29
R10165 VDD.n2535 VDD.n2515 2015.29
R10166 VDD.n2837 VDD.n2807 2015.29
R10167 VDD.n2793 VDD.n2773 2015.29
R10168 VDD.n3095 VDD.n3065 2015.29
R10169 VDD.n3051 VDD.n3031 2015.29
R10170 VDD.n3353 VDD.n3323 2015.29
R10171 VDD.n3309 VDD.n3289 2015.29
R10172 VDD.n5676 VDD.n5646 2015.29
R10173 VDD.n5632 VDD.n5612 2015.29
R10174 VDD.n5422 VDD.n5392 2015.29
R10175 VDD.n5378 VDD.n5358 2015.29
R10176 VDD.n3611 VDD.n3581 2015.29
R10177 VDD.n3567 VDD.n3547 2015.29
R10178 VDD.n3869 VDD.n3839 2015.29
R10179 VDD.n3825 VDD.n3805 2015.29
R10180 VDD.n4127 VDD.n4097 2015.29
R10181 VDD.n4083 VDD.n4063 2015.29
R10182 VDD.n4385 VDD.n4355 2015.29
R10183 VDD.n4341 VDD.n4321 2015.29
R10184 VDD.n4643 VDD.n4613 2015.29
R10185 VDD.n4599 VDD.n4579 2015.29
R10186 VDD.n4901 VDD.n4871 2015.29
R10187 VDD.n4857 VDD.n4837 2015.29
R10188 VDD.n5159 VDD.n5129 2015.29
R10189 VDD.n5115 VDD.n5095 2015.29
R10190 VDD.n1904 VDD.n1894 1997.65
R10191 VDD.n1899 VDD.n1894 1997.65
R10192 VDD.n1868 VDD.n1850 1997.65
R10193 VDD.n1868 VDD.n1851 1997.65
R10194 VDD.n2189 VDD.n2171 1997.65
R10195 VDD.n2189 VDD.n2172 1997.65
R10196 VDD.n2225 VDD.n2215 1997.65
R10197 VDD.n2220 VDD.n2215 1997.65
R10198 VDD.n2447 VDD.n2429 1997.65
R10199 VDD.n2447 VDD.n2430 1997.65
R10200 VDD.n2483 VDD.n2473 1997.65
R10201 VDD.n2478 VDD.n2473 1997.65
R10202 VDD.n2705 VDD.n2687 1997.65
R10203 VDD.n2705 VDD.n2688 1997.65
R10204 VDD.n2741 VDD.n2731 1997.65
R10205 VDD.n2736 VDD.n2731 1997.65
R10206 VDD.n2963 VDD.n2945 1997.65
R10207 VDD.n2963 VDD.n2946 1997.65
R10208 VDD.n2999 VDD.n2989 1997.65
R10209 VDD.n2994 VDD.n2989 1997.65
R10210 VDD.n3221 VDD.n3203 1997.65
R10211 VDD.n3221 VDD.n3204 1997.65
R10212 VDD.n3257 VDD.n3247 1997.65
R10213 VDD.n3252 VDD.n3247 1997.65
R10214 VDD.n3479 VDD.n3461 1997.65
R10215 VDD.n3479 VDD.n3462 1997.65
R10216 VDD.n3515 VDD.n3505 1997.65
R10217 VDD.n3510 VDD.n3505 1997.65
R10218 VDD.n5799 VDD.n5781 1997.65
R10219 VDD.n5799 VDD.n5782 1997.65
R10220 VDD.n5835 VDD.n5825 1997.65
R10221 VDD.n5830 VDD.n5825 1997.65
R10222 VDD.n5545 VDD.n5527 1997.65
R10223 VDD.n5545 VDD.n5528 1997.65
R10224 VDD.n5581 VDD.n5571 1997.65
R10225 VDD.n5576 VDD.n5571 1997.65
R10226 VDD.n3737 VDD.n3719 1997.65
R10227 VDD.n3737 VDD.n3720 1997.65
R10228 VDD.n3773 VDD.n3763 1997.65
R10229 VDD.n3768 VDD.n3763 1997.65
R10230 VDD.n3995 VDD.n3977 1997.65
R10231 VDD.n3995 VDD.n3978 1997.65
R10232 VDD.n4031 VDD.n4021 1997.65
R10233 VDD.n4026 VDD.n4021 1997.65
R10234 VDD.n4253 VDD.n4235 1997.65
R10235 VDD.n4253 VDD.n4236 1997.65
R10236 VDD.n4289 VDD.n4279 1997.65
R10237 VDD.n4284 VDD.n4279 1997.65
R10238 VDD.n4511 VDD.n4493 1997.65
R10239 VDD.n4511 VDD.n4494 1997.65
R10240 VDD.n4547 VDD.n4537 1997.65
R10241 VDD.n4542 VDD.n4537 1997.65
R10242 VDD.n4769 VDD.n4751 1997.65
R10243 VDD.n4769 VDD.n4752 1997.65
R10244 VDD.n4805 VDD.n4795 1997.65
R10245 VDD.n4800 VDD.n4795 1997.65
R10246 VDD.n5027 VDD.n5009 1997.65
R10247 VDD.n5027 VDD.n5010 1997.65
R10248 VDD.n5063 VDD.n5053 1997.65
R10249 VDD.n5058 VDD.n5053 1997.65
R10250 VDD.n5285 VDD.n5267 1997.65
R10251 VDD.n5285 VDD.n5268 1997.65
R10252 VDD.n5321 VDD.n5311 1997.65
R10253 VDD.n5316 VDD.n5311 1997.65
R10254 VDD.n1878 VDD.n1819 1814.12
R10255 VDD.n2199 VDD.n2140 1814.12
R10256 VDD.n2457 VDD.n2398 1814.12
R10257 VDD.n2715 VDD.n2656 1814.12
R10258 VDD.n2973 VDD.n2914 1814.12
R10259 VDD.n3231 VDD.n3172 1814.12
R10260 VDD.n3489 VDD.n3430 1814.12
R10261 VDD.n5809 VDD.n5750 1814.12
R10262 VDD.n5555 VDD.n5496 1814.12
R10263 VDD.n3747 VDD.n3688 1814.12
R10264 VDD.n4005 VDD.n3946 1814.12
R10265 VDD.n4263 VDD.n4204 1814.12
R10266 VDD.n4521 VDD.n4462 1814.12
R10267 VDD.n4779 VDD.n4720 1814.12
R10268 VDD.n5037 VDD.n4978 1814.12
R10269 VDD.n5295 VDD.n5236 1814.12
R10270 VDD.n1881 VDD.n1880 1598.82
R10271 VDD.n2202 VDD.n2201 1598.82
R10272 VDD.n2460 VDD.n2459 1598.82
R10273 VDD.n2718 VDD.n2717 1598.82
R10274 VDD.n2976 VDD.n2975 1598.82
R10275 VDD.n3234 VDD.n3233 1598.82
R10276 VDD.n3492 VDD.n3491 1598.82
R10277 VDD.n5812 VDD.n5811 1598.82
R10278 VDD.n5558 VDD.n5557 1598.82
R10279 VDD.n3750 VDD.n3749 1598.82
R10280 VDD.n4008 VDD.n4007 1598.82
R10281 VDD.n4266 VDD.n4265 1598.82
R10282 VDD.n4524 VDD.n4523 1598.82
R10283 VDD.n4782 VDD.n4781 1598.82
R10284 VDD.n5040 VDD.n5039 1598.82
R10285 VDD.n5298 VDD.n5297 1598.82
R10286 VDD.n1698 VDD.n1697 1514.12
R10287 VDD.n2047 VDD.n2046 1514.12
R10288 VDD.n2277 VDD.n2276 1514.12
R10289 VDD.n2535 VDD.n2534 1514.12
R10290 VDD.n2793 VDD.n2792 1514.12
R10291 VDD.n3051 VDD.n3050 1514.12
R10292 VDD.n3309 VDD.n3308 1514.12
R10293 VDD.n5632 VDD.n5631 1514.12
R10294 VDD.n5378 VDD.n5377 1514.12
R10295 VDD.n3567 VDD.n3566 1514.12
R10296 VDD.n3825 VDD.n3824 1514.12
R10297 VDD.n4083 VDD.n4082 1514.12
R10298 VDD.n4341 VDD.n4340 1514.12
R10299 VDD.n4599 VDD.n4598 1514.12
R10300 VDD.n4857 VDD.n4856 1514.12
R10301 VDD.n5115 VDD.n5114 1514.12
R10302 VDD.n1856 VDD.n1844 1440
R10303 VDD.n1869 VDD.n1846 1440
R10304 VDD.n2177 VDD.n2165 1440
R10305 VDD.n2190 VDD.n2167 1440
R10306 VDD.n2435 VDD.n2423 1440
R10307 VDD.n2448 VDD.n2425 1440
R10308 VDD.n2693 VDD.n2681 1440
R10309 VDD.n2706 VDD.n2683 1440
R10310 VDD.n2951 VDD.n2939 1440
R10311 VDD.n2964 VDD.n2941 1440
R10312 VDD.n3209 VDD.n3197 1440
R10313 VDD.n3222 VDD.n3199 1440
R10314 VDD.n3467 VDD.n3455 1440
R10315 VDD.n3480 VDD.n3457 1440
R10316 VDD.n5787 VDD.n5775 1440
R10317 VDD.n5800 VDD.n5777 1440
R10318 VDD.n5533 VDD.n5521 1440
R10319 VDD.n5546 VDD.n5523 1440
R10320 VDD.n3725 VDD.n3713 1440
R10321 VDD.n3738 VDD.n3715 1440
R10322 VDD.n3983 VDD.n3971 1440
R10323 VDD.n3996 VDD.n3973 1440
R10324 VDD.n4241 VDD.n4229 1440
R10325 VDD.n4254 VDD.n4231 1440
R10326 VDD.n4499 VDD.n4487 1440
R10327 VDD.n4512 VDD.n4489 1440
R10328 VDD.n4757 VDD.n4745 1440
R10329 VDD.n4770 VDD.n4747 1440
R10330 VDD.n5015 VDD.n5003 1440
R10331 VDD.n5028 VDD.n5005 1440
R10332 VDD.n5273 VDD.n5261 1440
R10333 VDD.n5286 VDD.n5263 1440
R10334 VDD.n1915 VDD.n1890 1422.35
R10335 VDD.n1900 VDD.n1891 1422.35
R10336 VDD.n2236 VDD.n2211 1422.35
R10337 VDD.n2221 VDD.n2212 1422.35
R10338 VDD.n2494 VDD.n2469 1422.35
R10339 VDD.n2479 VDD.n2470 1422.35
R10340 VDD.n2752 VDD.n2727 1422.35
R10341 VDD.n2737 VDD.n2728 1422.35
R10342 VDD.n3010 VDD.n2985 1422.35
R10343 VDD.n2995 VDD.n2986 1422.35
R10344 VDD.n3268 VDD.n3243 1422.35
R10345 VDD.n3253 VDD.n3244 1422.35
R10346 VDD.n3526 VDD.n3501 1422.35
R10347 VDD.n3511 VDD.n3502 1422.35
R10348 VDD.n5846 VDD.n5821 1422.35
R10349 VDD.n5831 VDD.n5822 1422.35
R10350 VDD.n5592 VDD.n5567 1422.35
R10351 VDD.n5577 VDD.n5568 1422.35
R10352 VDD.n3784 VDD.n3759 1422.35
R10353 VDD.n3769 VDD.n3760 1422.35
R10354 VDD.n4042 VDD.n4017 1422.35
R10355 VDD.n4027 VDD.n4018 1422.35
R10356 VDD.n4300 VDD.n4275 1422.35
R10357 VDD.n4285 VDD.n4276 1422.35
R10358 VDD.n4558 VDD.n4533 1422.35
R10359 VDD.n4543 VDD.n4534 1422.35
R10360 VDD.n4816 VDD.n4791 1422.35
R10361 VDD.n4801 VDD.n4792 1422.35
R10362 VDD.n5074 VDD.n5049 1422.35
R10363 VDD.n5059 VDD.n5050 1422.35
R10364 VDD.n5332 VDD.n5307 1422.35
R10365 VDD.n5317 VDD.n5308 1422.35
R10366 VDD.n857 VDD 1319.65
R10367 VDD.n1240 VDD 1319.65
R10368 VDD.n1713 VDD.n1676 1231.76
R10369 VDD.n2062 VDD.n2025 1231.76
R10370 VDD.n2292 VDD.n2255 1231.76
R10371 VDD.n2550 VDD.n2513 1231.76
R10372 VDD.n2808 VDD.n2771 1231.76
R10373 VDD.n3066 VDD.n3029 1231.76
R10374 VDD.n3324 VDD.n3287 1231.76
R10375 VDD.n5647 VDD.n5610 1231.76
R10376 VDD.n5393 VDD.n5356 1231.76
R10377 VDD.n3582 VDD.n3545 1231.76
R10378 VDD.n3840 VDD.n3803 1231.76
R10379 VDD.n4098 VDD.n4061 1231.76
R10380 VDD.n4356 VDD.n4319 1231.76
R10381 VDD.n4614 VDD.n4577 1231.76
R10382 VDD.n4872 VDD.n4835 1231.76
R10383 VDD.n5130 VDD.n5093 1231.76
R10384 VDD.n1765 VDD.n1674 1228.24
R10385 VDD.n2114 VDD.n2023 1228.24
R10386 VDD.n2344 VDD.n2253 1228.24
R10387 VDD.n2602 VDD.n2511 1228.24
R10388 VDD.n2860 VDD.n2769 1228.24
R10389 VDD.n3118 VDD.n3027 1228.24
R10390 VDD.n3376 VDD.n3285 1228.24
R10391 VDD.n5699 VDD.n5608 1228.24
R10392 VDD.n5445 VDD.n5354 1228.24
R10393 VDD.n3634 VDD.n3543 1228.24
R10394 VDD.n3892 VDD.n3801 1228.24
R10395 VDD.n4150 VDD.n4059 1228.24
R10396 VDD.n4408 VDD.n4317 1228.24
R10397 VDD.n4666 VDD.n4575 1228.24
R10398 VDD.n4924 VDD.n4833 1228.24
R10399 VDD.n5182 VDD.n5091 1228.24
R10400 VDD.n1765 VDD.n1675 1224.71
R10401 VDD.n1676 VDD.n1675 1224.71
R10402 VDD.n2114 VDD.n2024 1224.71
R10403 VDD.n2025 VDD.n2024 1224.71
R10404 VDD.n2344 VDD.n2254 1224.71
R10405 VDD.n2255 VDD.n2254 1224.71
R10406 VDD.n2602 VDD.n2512 1224.71
R10407 VDD.n2513 VDD.n2512 1224.71
R10408 VDD.n2860 VDD.n2770 1224.71
R10409 VDD.n2771 VDD.n2770 1224.71
R10410 VDD.n3118 VDD.n3028 1224.71
R10411 VDD.n3029 VDD.n3028 1224.71
R10412 VDD.n3376 VDD.n3286 1224.71
R10413 VDD.n3287 VDD.n3286 1224.71
R10414 VDD.n5699 VDD.n5609 1224.71
R10415 VDD.n5610 VDD.n5609 1224.71
R10416 VDD.n5445 VDD.n5355 1224.71
R10417 VDD.n5356 VDD.n5355 1224.71
R10418 VDD.n3634 VDD.n3544 1224.71
R10419 VDD.n3545 VDD.n3544 1224.71
R10420 VDD.n3892 VDD.n3802 1224.71
R10421 VDD.n3803 VDD.n3802 1224.71
R10422 VDD.n4150 VDD.n4060 1224.71
R10423 VDD.n4061 VDD.n4060 1224.71
R10424 VDD.n4408 VDD.n4318 1224.71
R10425 VDD.n4319 VDD.n4318 1224.71
R10426 VDD.n4666 VDD.n4576 1224.71
R10427 VDD.n4577 VDD.n4576 1224.71
R10428 VDD.n4924 VDD.n4834 1224.71
R10429 VDD.n4835 VDD.n4834 1224.71
R10430 VDD.n5182 VDD.n5092 1224.71
R10431 VDD.n5093 VDD.n5092 1224.71
R10432 VDD.n1718 VDD.n1675 1153.33
R10433 VDD.n2067 VDD.n2024 1153.33
R10434 VDD.n2297 VDD.n2254 1153.33
R10435 VDD.n2555 VDD.n2512 1153.33
R10436 VDD.n2813 VDD.n2770 1153.33
R10437 VDD.n3071 VDD.n3028 1153.33
R10438 VDD.n3329 VDD.n3286 1153.33
R10439 VDD.n5652 VDD.n5609 1153.33
R10440 VDD.n5398 VDD.n5355 1153.33
R10441 VDD.n3587 VDD.n3544 1153.33
R10442 VDD.n3845 VDD.n3802 1153.33
R10443 VDD.n4103 VDD.n4060 1153.33
R10444 VDD.n4361 VDD.n4318 1153.33
R10445 VDD.n4619 VDD.n4576 1153.33
R10446 VDD.n4877 VDD.n4834 1153.33
R10447 VDD.n5135 VDD.n5092 1153.33
R10448 VDD.n1902 VDD.n1900 1143.53
R10449 VDD.n2223 VDD.n2221 1143.53
R10450 VDD.n2481 VDD.n2479 1143.53
R10451 VDD.n2739 VDD.n2737 1143.53
R10452 VDD.n2997 VDD.n2995 1143.53
R10453 VDD.n3255 VDD.n3253 1143.53
R10454 VDD.n3513 VDD.n3511 1143.53
R10455 VDD.n5833 VDD.n5831 1143.53
R10456 VDD.n5579 VDD.n5577 1143.53
R10457 VDD.n3771 VDD.n3769 1143.53
R10458 VDD.n4029 VDD.n4027 1143.53
R10459 VDD.n4287 VDD.n4285 1143.53
R10460 VDD.n4545 VDD.n4543 1143.53
R10461 VDD.n4803 VDD.n4801 1143.53
R10462 VDD.n5061 VDD.n5059 1143.53
R10463 VDD.n5319 VDD.n5317 1143.53
R10464 VDD.n1862 VDD.n1846 1125.88
R10465 VDD.n2183 VDD.n2167 1125.88
R10466 VDD.n2441 VDD.n2425 1125.88
R10467 VDD.n2699 VDD.n2683 1125.88
R10468 VDD.n2957 VDD.n2941 1125.88
R10469 VDD.n3215 VDD.n3199 1125.88
R10470 VDD.n3473 VDD.n3457 1125.88
R10471 VDD.n5793 VDD.n5777 1125.88
R10472 VDD.n5539 VDD.n5523 1125.88
R10473 VDD.n3731 VDD.n3715 1125.88
R10474 VDD.n3989 VDD.n3973 1125.88
R10475 VDD.n4247 VDD.n4231 1125.88
R10476 VDD.n4505 VDD.n4489 1125.88
R10477 VDD.n4763 VDD.n4747 1125.88
R10478 VDD.n5021 VDD.n5005 1125.88
R10479 VDD.n5279 VDD.n5263 1125.88
R10480 VDD.n1756 VDD.n1718 1072.94
R10481 VDD.n2105 VDD.n2067 1072.94
R10482 VDD.n2335 VDD.n2297 1072.94
R10483 VDD.n2593 VDD.n2555 1072.94
R10484 VDD.n2851 VDD.n2813 1072.94
R10485 VDD.n3109 VDD.n3071 1072.94
R10486 VDD.n3367 VDD.n3329 1072.94
R10487 VDD.n5690 VDD.n5652 1072.94
R10488 VDD.n5436 VDD.n5398 1072.94
R10489 VDD.n3625 VDD.n3587 1072.94
R10490 VDD.n3883 VDD.n3845 1072.94
R10491 VDD.n4141 VDD.n4103 1072.94
R10492 VDD.n4399 VDD.n4361 1072.94
R10493 VDD.n4657 VDD.n4619 1072.94
R10494 VDD.n4915 VDD.n4877 1072.94
R10495 VDD.n5173 VDD.n5135 1072.94
R10496 VDD.n1718 VDD.n1670 1069.41
R10497 VDD.n2067 VDD.n2019 1069.41
R10498 VDD.n2297 VDD.n2249 1069.41
R10499 VDD.n2555 VDD.n2507 1069.41
R10500 VDD.n2813 VDD.n2765 1069.41
R10501 VDD.n3071 VDD.n3023 1069.41
R10502 VDD.n3329 VDD.n3281 1069.41
R10503 VDD.n5652 VDD.n5604 1069.41
R10504 VDD.n5398 VDD.n5350 1069.41
R10505 VDD.n3587 VDD.n3539 1069.41
R10506 VDD.n3845 VDD.n3797 1069.41
R10507 VDD.n4103 VDD.n4055 1069.41
R10508 VDD.n4361 VDD.n4313 1069.41
R10509 VDD.n4619 VDD.n4571 1069.41
R10510 VDD.n4877 VDD.n4829 1069.41
R10511 VDD.n5135 VDD.n5087 1069.41
R10512 VDD.n1906 VDD.n1890 1051.76
R10513 VDD.n1856 VDD.n1855 1051.76
R10514 VDD.n2177 VDD.n2176 1051.76
R10515 VDD.n2227 VDD.n2211 1051.76
R10516 VDD.n2435 VDD.n2434 1051.76
R10517 VDD.n2485 VDD.n2469 1051.76
R10518 VDD.n2693 VDD.n2692 1051.76
R10519 VDD.n2743 VDD.n2727 1051.76
R10520 VDD.n2951 VDD.n2950 1051.76
R10521 VDD.n3001 VDD.n2985 1051.76
R10522 VDD.n3209 VDD.n3208 1051.76
R10523 VDD.n3259 VDD.n3243 1051.76
R10524 VDD.n3467 VDD.n3466 1051.76
R10525 VDD.n3517 VDD.n3501 1051.76
R10526 VDD.n5787 VDD.n5786 1051.76
R10527 VDD.n5837 VDD.n5821 1051.76
R10528 VDD.n5533 VDD.n5532 1051.76
R10529 VDD.n5583 VDD.n5567 1051.76
R10530 VDD.n3725 VDD.n3724 1051.76
R10531 VDD.n3775 VDD.n3759 1051.76
R10532 VDD.n3983 VDD.n3982 1051.76
R10533 VDD.n4033 VDD.n4017 1051.76
R10534 VDD.n4241 VDD.n4240 1051.76
R10535 VDD.n4291 VDD.n4275 1051.76
R10536 VDD.n4499 VDD.n4498 1051.76
R10537 VDD.n4549 VDD.n4533 1051.76
R10538 VDD.n4757 VDD.n4756 1051.76
R10539 VDD.n4807 VDD.n4791 1051.76
R10540 VDD.n5015 VDD.n5014 1051.76
R10541 VDD.n5065 VDD.n5049 1051.76
R10542 VDD.n5273 VDD.n5272 1051.76
R10543 VDD.n5323 VDD.n5307 1051.76
R10544 VDD.n1960 VDD.n1942 862.871
R10545 VDD.n1950 VDD.n1942 862.871
R10546 VDD.n1971 VDD.n1930 862.871
R10547 VDD.n1967 VDD.n1930 862.871
R10548 VDD.n1759 VDD.n1758 861.178
R10549 VDD.n2108 VDD.n2107 861.178
R10550 VDD.n2338 VDD.n2337 861.178
R10551 VDD.n2596 VDD.n2595 861.178
R10552 VDD.n2854 VDD.n2853 861.178
R10553 VDD.n3112 VDD.n3111 861.178
R10554 VDD.n3370 VDD.n3369 861.178
R10555 VDD.n5693 VDD.n5692 861.178
R10556 VDD.n5439 VDD.n5438 861.178
R10557 VDD.n3628 VDD.n3627 861.178
R10558 VDD.n3886 VDD.n3885 861.178
R10559 VDD.n4144 VDD.n4143 861.178
R10560 VDD.n4402 VDD.n4401 861.178
R10561 VDD.n4660 VDD.n4659 861.178
R10562 VDD.n4918 VDD.n4917 861.178
R10563 VDD.n5176 VDD.n5175 861.178
R10564 VDD.n1962 VDD.n1961 857.648
R10565 VDD.n1963 VDD.n1962 857.648
R10566 VDD.n1963 VDD.n1928 857.648
R10567 VDD.n1970 VDD.n1928 857.648
R10568 VDD.n1951 VDD.n1938 857.648
R10569 VDD.n1964 VDD.n1938 857.648
R10570 VDD.n1964 VDD.n1932 857.648
R10571 VDD.n1968 VDD.n1932 857.648
R10572 VDD.n1883 VDD.n1819 751.765
R10573 VDD.n2204 VDD.n2140 751.765
R10574 VDD.n2462 VDD.n2398 751.765
R10575 VDD.n2720 VDD.n2656 751.765
R10576 VDD.n2978 VDD.n2914 751.765
R10577 VDD.n3236 VDD.n3172 751.765
R10578 VDD.n3494 VDD.n3430 751.765
R10579 VDD.n5814 VDD.n5750 751.765
R10580 VDD.n5560 VDD.n5496 751.765
R10581 VDD.n3752 VDD.n3688 751.765
R10582 VDD.n4010 VDD.n3946 751.765
R10583 VDD.n4268 VDD.n4204 751.765
R10584 VDD.n4526 VDD.n4462 751.765
R10585 VDD.n4784 VDD.n4720 751.765
R10586 VDD.n5042 VDD.n4978 751.765
R10587 VDD.n5300 VDD.n5236 751.765
R10588 VDD.n1714 VDD.n1712 723.529
R10589 VDD.n2063 VDD.n2061 723.529
R10590 VDD.n2293 VDD.n2291 723.529
R10591 VDD.n2551 VDD.n2549 723.529
R10592 VDD.n2809 VDD.n2807 723.529
R10593 VDD.n3067 VDD.n3065 723.529
R10594 VDD.n3325 VDD.n3323 723.529
R10595 VDD.n5648 VDD.n5646 723.529
R10596 VDD.n5394 VDD.n5392 723.529
R10597 VDD.n3583 VDD.n3581 723.529
R10598 VDD.n3841 VDD.n3839 723.529
R10599 VDD.n4099 VDD.n4097 723.529
R10600 VDD.n4357 VDD.n4355 723.529
R10601 VDD.n4615 VDD.n4613 723.529
R10602 VDD.n4873 VDD.n4871 723.529
R10603 VDD.n5131 VDD.n5129 723.529
R10604 VDD.n1680 VDD.n1678 720
R10605 VDD.n2029 VDD.n2027 720
R10606 VDD.n2259 VDD.n2257 720
R10607 VDD.n2517 VDD.n2515 720
R10608 VDD.n2775 VDD.n2773 720
R10609 VDD.n3033 VDD.n3031 720
R10610 VDD.n3291 VDD.n3289 720
R10611 VDD.n5614 VDD.n5612 720
R10612 VDD.n5360 VDD.n5358 720
R10613 VDD.n3549 VDD.n3547 720
R10614 VDD.n3807 VDD.n3805 720
R10615 VDD.n4065 VDD.n4063 720
R10616 VDD.n4323 VDD.n4321 720
R10617 VDD.n4581 VDD.n4579 720
R10618 VDD.n4839 VDD.n4837 720
R10619 VDD.n5097 VDD.n5095 720
R10620 VDD.n1695 VDD.t642 632.183
R10621 VDD.n2044 VDD.t243 632.183
R10622 VDD.n2274 VDD.t624 632.183
R10623 VDD.n2532 VDD.t842 632.183
R10624 VDD.n2790 VDD.t134 632.183
R10625 VDD.n3048 VDD.t473 632.183
R10626 VDD.n3306 VDD.t1331 632.183
R10627 VDD.n5629 VDD.t613 632.183
R10628 VDD.n5375 VDD.t6 632.183
R10629 VDD.n3564 VDD.t631 632.183
R10630 VDD.n3822 VDD.t1386 632.183
R10631 VDD.n4080 VDD.t888 632.183
R10632 VDD.n4338 VDD.t126 632.183
R10633 VDD.n4596 VDD.t72 632.183
R10634 VDD.n4854 VDD.t783 632.183
R10635 VDD.n5112 VDD.t1374 632.183
R10636 VDD.n1677 VDD.n1674 593.144
R10637 VDD.n1680 VDD.n1677 593.144
R10638 VDD.n2026 VDD.n2023 593.144
R10639 VDD.n2029 VDD.n2026 593.144
R10640 VDD.n2256 VDD.n2253 593.144
R10641 VDD.n2259 VDD.n2256 593.144
R10642 VDD.n2514 VDD.n2511 593.144
R10643 VDD.n2517 VDD.n2514 593.144
R10644 VDD.n2772 VDD.n2769 593.144
R10645 VDD.n2775 VDD.n2772 593.144
R10646 VDD.n3030 VDD.n3027 593.144
R10647 VDD.n3033 VDD.n3030 593.144
R10648 VDD.n3288 VDD.n3285 593.144
R10649 VDD.n3291 VDD.n3288 593.144
R10650 VDD.n5611 VDD.n5608 593.144
R10651 VDD.n5614 VDD.n5611 593.144
R10652 VDD.n5357 VDD.n5354 593.144
R10653 VDD.n5360 VDD.n5357 593.144
R10654 VDD.n3546 VDD.n3543 593.144
R10655 VDD.n3549 VDD.n3546 593.144
R10656 VDD.n3804 VDD.n3801 593.144
R10657 VDD.n3807 VDD.n3804 593.144
R10658 VDD.n4062 VDD.n4059 593.144
R10659 VDD.n4065 VDD.n4062 593.144
R10660 VDD.n4320 VDD.n4317 593.144
R10661 VDD.n4323 VDD.n4320 593.144
R10662 VDD.n4578 VDD.n4575 593.144
R10663 VDD.n4581 VDD.n4578 593.144
R10664 VDD.n4836 VDD.n4833 593.144
R10665 VDD.n4839 VDD.n4836 593.144
R10666 VDD.n5094 VDD.n5091 593.144
R10667 VDD.n5097 VDD.n5094 593.144
R10668 VDD.n1795 VDD.t1363 584.644
R10669 VDD.n1781 VDD.t646 584.644
R10670 VDD.n2003 VDD.t1497 584.644
R10671 VDD.n1989 VDD.t247 584.644
R10672 VDD.n2374 VDD.t227 584.644
R10673 VDD.n2360 VDD.t623 584.644
R10674 VDD.n2632 VDD.t61 584.644
R10675 VDD.n2618 VDD.t849 584.644
R10676 VDD.n2890 VDD.t600 584.644
R10677 VDD.n2876 VDD.t137 584.644
R10678 VDD.n3148 VDD.t46 584.644
R10679 VDD.n3134 VDD.t477 584.644
R10680 VDD.n3406 VDD.t736 584.644
R10681 VDD.n3392 VDD.t1338 584.644
R10682 VDD.n5729 VDD.t169 584.644
R10683 VDD.n5715 VDD.t617 584.644
R10684 VDD.n5475 VDD.t521 584.644
R10685 VDD.n5461 VDD.t5 584.644
R10686 VDD.n3664 VDD.t192 584.644
R10687 VDD.n3650 VDD.t638 584.644
R10688 VDD.n3922 VDD.t176 584.644
R10689 VDD.n3908 VDD.t1385 584.644
R10690 VDD.n4180 VDD.t96 584.644
R10691 VDD.n4166 VDD.t887 584.644
R10692 VDD.n4438 VDD.t502 584.644
R10693 VDD.n4424 VDD.t129 584.644
R10694 VDD.n4696 VDD.t592 584.644
R10695 VDD.n4682 VDD.t76 584.644
R10696 VDD.n4954 VDD.t584 584.644
R10697 VDD.n4940 VDD.t790 584.644
R10698 VDD.n5212 VDD.t862 584.644
R10699 VDD.n5198 VDD.t1377 584.644
R10700 VDD.n523 VDD.t567 584.644
R10701 VDD.n873 VDD.t52 584.644
R10702 VDD.n122 VDD.t65 584.644
R10703 VDD.n1348 VDD.t660 584.644
R10704 VDD.n1763 VDD.n1713 576.668
R10705 VDD.n1763 VDD.n1714 576.668
R10706 VDD.n2112 VDD.n2062 576.668
R10707 VDD.n2112 VDD.n2063 576.668
R10708 VDD.n2342 VDD.n2292 576.668
R10709 VDD.n2342 VDD.n2293 576.668
R10710 VDD.n2600 VDD.n2550 576.668
R10711 VDD.n2600 VDD.n2551 576.668
R10712 VDD.n2858 VDD.n2808 576.668
R10713 VDD.n2858 VDD.n2809 576.668
R10714 VDD.n3116 VDD.n3066 576.668
R10715 VDD.n3116 VDD.n3067 576.668
R10716 VDD.n3374 VDD.n3324 576.668
R10717 VDD.n3374 VDD.n3325 576.668
R10718 VDD.n5697 VDD.n5647 576.668
R10719 VDD.n5697 VDD.n5648 576.668
R10720 VDD.n5443 VDD.n5393 576.668
R10721 VDD.n5443 VDD.n5394 576.668
R10722 VDD.n3632 VDD.n3582 576.668
R10723 VDD.n3632 VDD.n3583 576.668
R10724 VDD.n3890 VDD.n3840 576.668
R10725 VDD.n3890 VDD.n3841 576.668
R10726 VDD.n4148 VDD.n4098 576.668
R10727 VDD.n4148 VDD.n4099 576.668
R10728 VDD.n4406 VDD.n4356 576.668
R10729 VDD.n4406 VDD.n4357 576.668
R10730 VDD.n4664 VDD.n4614 576.668
R10731 VDD.n4664 VDD.n4615 576.668
R10732 VDD.n4922 VDD.n4872 576.668
R10733 VDD.n4922 VDD.n4873 576.668
R10734 VDD.n5180 VDD.n5130 576.668
R10735 VDD.n5180 VDD.n5131 576.668
R10736 VDD.n1906 VDD.n1904 568.236
R10737 VDD.n1899 VDD.n1896 568.236
R10738 VDD.n1902 VDD.n1899 568.236
R10739 VDD.n1904 VDD.n1895 568.236
R10740 VDD.n1859 VDD.n1850 568.236
R10741 VDD.n1862 VDD.n1851 568.236
R10742 VDD.n1864 VDD.n1851 568.236
R10743 VDD.n1855 VDD.n1850 568.236
R10744 VDD.n2180 VDD.n2171 568.236
R10745 VDD.n2183 VDD.n2172 568.236
R10746 VDD.n2185 VDD.n2172 568.236
R10747 VDD.n2176 VDD.n2171 568.236
R10748 VDD.n2227 VDD.n2225 568.236
R10749 VDD.n2220 VDD.n2217 568.236
R10750 VDD.n2223 VDD.n2220 568.236
R10751 VDD.n2225 VDD.n2216 568.236
R10752 VDD.n2438 VDD.n2429 568.236
R10753 VDD.n2441 VDD.n2430 568.236
R10754 VDD.n2443 VDD.n2430 568.236
R10755 VDD.n2434 VDD.n2429 568.236
R10756 VDD.n2485 VDD.n2483 568.236
R10757 VDD.n2478 VDD.n2475 568.236
R10758 VDD.n2481 VDD.n2478 568.236
R10759 VDD.n2483 VDD.n2474 568.236
R10760 VDD.n2696 VDD.n2687 568.236
R10761 VDD.n2699 VDD.n2688 568.236
R10762 VDD.n2701 VDD.n2688 568.236
R10763 VDD.n2692 VDD.n2687 568.236
R10764 VDD.n2743 VDD.n2741 568.236
R10765 VDD.n2736 VDD.n2733 568.236
R10766 VDD.n2739 VDD.n2736 568.236
R10767 VDD.n2741 VDD.n2732 568.236
R10768 VDD.n2954 VDD.n2945 568.236
R10769 VDD.n2957 VDD.n2946 568.236
R10770 VDD.n2959 VDD.n2946 568.236
R10771 VDD.n2950 VDD.n2945 568.236
R10772 VDD.n3001 VDD.n2999 568.236
R10773 VDD.n2994 VDD.n2991 568.236
R10774 VDD.n2997 VDD.n2994 568.236
R10775 VDD.n2999 VDD.n2990 568.236
R10776 VDD.n3212 VDD.n3203 568.236
R10777 VDD.n3215 VDD.n3204 568.236
R10778 VDD.n3217 VDD.n3204 568.236
R10779 VDD.n3208 VDD.n3203 568.236
R10780 VDD.n3259 VDD.n3257 568.236
R10781 VDD.n3252 VDD.n3249 568.236
R10782 VDD.n3255 VDD.n3252 568.236
R10783 VDD.n3257 VDD.n3248 568.236
R10784 VDD.n3470 VDD.n3461 568.236
R10785 VDD.n3473 VDD.n3462 568.236
R10786 VDD.n3475 VDD.n3462 568.236
R10787 VDD.n3466 VDD.n3461 568.236
R10788 VDD.n3517 VDD.n3515 568.236
R10789 VDD.n3510 VDD.n3507 568.236
R10790 VDD.n3513 VDD.n3510 568.236
R10791 VDD.n3515 VDD.n3506 568.236
R10792 VDD.n5790 VDD.n5781 568.236
R10793 VDD.n5793 VDD.n5782 568.236
R10794 VDD.n5795 VDD.n5782 568.236
R10795 VDD.n5786 VDD.n5781 568.236
R10796 VDD.n5837 VDD.n5835 568.236
R10797 VDD.n5830 VDD.n5827 568.236
R10798 VDD.n5833 VDD.n5830 568.236
R10799 VDD.n5835 VDD.n5826 568.236
R10800 VDD.n5536 VDD.n5527 568.236
R10801 VDD.n5539 VDD.n5528 568.236
R10802 VDD.n5541 VDD.n5528 568.236
R10803 VDD.n5532 VDD.n5527 568.236
R10804 VDD.n5583 VDD.n5581 568.236
R10805 VDD.n5576 VDD.n5573 568.236
R10806 VDD.n5579 VDD.n5576 568.236
R10807 VDD.n5581 VDD.n5572 568.236
R10808 VDD.n3728 VDD.n3719 568.236
R10809 VDD.n3731 VDD.n3720 568.236
R10810 VDD.n3733 VDD.n3720 568.236
R10811 VDD.n3724 VDD.n3719 568.236
R10812 VDD.n3775 VDD.n3773 568.236
R10813 VDD.n3768 VDD.n3765 568.236
R10814 VDD.n3771 VDD.n3768 568.236
R10815 VDD.n3773 VDD.n3764 568.236
R10816 VDD.n3986 VDD.n3977 568.236
R10817 VDD.n3989 VDD.n3978 568.236
R10818 VDD.n3991 VDD.n3978 568.236
R10819 VDD.n3982 VDD.n3977 568.236
R10820 VDD.n4033 VDD.n4031 568.236
R10821 VDD.n4026 VDD.n4023 568.236
R10822 VDD.n4029 VDD.n4026 568.236
R10823 VDD.n4031 VDD.n4022 568.236
R10824 VDD.n4244 VDD.n4235 568.236
R10825 VDD.n4247 VDD.n4236 568.236
R10826 VDD.n4249 VDD.n4236 568.236
R10827 VDD.n4240 VDD.n4235 568.236
R10828 VDD.n4291 VDD.n4289 568.236
R10829 VDD.n4284 VDD.n4281 568.236
R10830 VDD.n4287 VDD.n4284 568.236
R10831 VDD.n4289 VDD.n4280 568.236
R10832 VDD.n4502 VDD.n4493 568.236
R10833 VDD.n4505 VDD.n4494 568.236
R10834 VDD.n4507 VDD.n4494 568.236
R10835 VDD.n4498 VDD.n4493 568.236
R10836 VDD.n4549 VDD.n4547 568.236
R10837 VDD.n4542 VDD.n4539 568.236
R10838 VDD.n4545 VDD.n4542 568.236
R10839 VDD.n4547 VDD.n4538 568.236
R10840 VDD.n4760 VDD.n4751 568.236
R10841 VDD.n4763 VDD.n4752 568.236
R10842 VDD.n4765 VDD.n4752 568.236
R10843 VDD.n4756 VDD.n4751 568.236
R10844 VDD.n4807 VDD.n4805 568.236
R10845 VDD.n4800 VDD.n4797 568.236
R10846 VDD.n4803 VDD.n4800 568.236
R10847 VDD.n4805 VDD.n4796 568.236
R10848 VDD.n5018 VDD.n5009 568.236
R10849 VDD.n5021 VDD.n5010 568.236
R10850 VDD.n5023 VDD.n5010 568.236
R10851 VDD.n5014 VDD.n5009 568.236
R10852 VDD.n5065 VDD.n5063 568.236
R10853 VDD.n5058 VDD.n5055 568.236
R10854 VDD.n5061 VDD.n5058 568.236
R10855 VDD.n5063 VDD.n5054 568.236
R10856 VDD.n5276 VDD.n5267 568.236
R10857 VDD.n5279 VDD.n5268 568.236
R10858 VDD.n5281 VDD.n5268 568.236
R10859 VDD.n5272 VDD.n5267 568.236
R10860 VDD.n5323 VDD.n5321 568.236
R10861 VDD.n5316 VDD.n5313 568.236
R10862 VDD.n5319 VDD.n5316 568.236
R10863 VDD.n5321 VDD.n5312 568.236
R10864 VDD.n857 VDD.t804 533.735
R10865 VDD.n1240 VDD.t767 533.735
R10866 VDD.n1744 VDD.n1743 481.226
R10867 VDD.n2093 VDD.n2092 481.226
R10868 VDD.n2323 VDD.n2322 481.226
R10869 VDD.n2581 VDD.n2580 481.226
R10870 VDD.n2839 VDD.n2838 481.226
R10871 VDD.n3097 VDD.n3096 481.226
R10872 VDD.n3355 VDD.n3354 481.226
R10873 VDD.n5678 VDD.n5677 481.226
R10874 VDD.n5424 VDD.n5423 481.226
R10875 VDD.n3613 VDD.n3612 481.226
R10876 VDD.n3871 VDD.n3870 481.226
R10877 VDD.n4129 VDD.n4128 481.226
R10878 VDD.n4387 VDD.n4386 481.226
R10879 VDD.n4645 VDD.n4644 481.226
R10880 VDD.n4903 VDD.n4902 481.226
R10881 VDD.n5161 VDD.n5160 481.226
R10882 VDD.n1857 VDD.n1847 473.839
R10883 VDD.t106 VDD.n1849 473.839
R10884 VDD.n2178 VDD.n2168 473.839
R10885 VDD.t719 VDD.n2170 473.839
R10886 VDD.n2436 VDD.n2426 473.839
R10887 VDD.t485 VDD.n2428 473.839
R10888 VDD.n2694 VDD.n2684 473.839
R10889 VDD.t531 VDD.n2686 473.839
R10890 VDD.n2952 VDD.n2942 473.839
R10891 VDD.t15 VDD.n2944 473.839
R10892 VDD.n3210 VDD.n3200 473.839
R10893 VDD.t412 VDD.n3202 473.839
R10894 VDD.n3468 VDD.n3458 473.839
R10895 VDD.t538 VDD.n3460 473.839
R10896 VDD.n5788 VDD.n5778 473.839
R10897 VDD.t109 VDD.n5780 473.839
R10898 VDD.n5534 VDD.n5524 473.839
R10899 VDD.t186 VDD.n5526 473.839
R10900 VDD.n3726 VDD.n3716 473.839
R10901 VDD.t413 VDD.n3718 473.839
R10902 VDD.n3984 VDD.n3974 473.839
R10903 VDD.t108 VDD.n3976 473.839
R10904 VDD.n4242 VDD.n4232 473.839
R10905 VDD.t0 VDD.n4234 473.839
R10906 VDD.n4500 VDD.n4490 473.839
R10907 VDD.t13 VDD.n4492 473.839
R10908 VDD.n4758 VDD.n4748 473.839
R10909 VDD.t117 VDD.n4750 473.839
R10910 VDD.n5016 VDD.n5006 473.839
R10911 VDD.t651 VDD.n5008 473.839
R10912 VDD.n5274 VDD.n5264 473.839
R10913 VDD.t85 VDD.n5266 473.839
R10914 VDD.n1914 VDD.n1892 468.033
R10915 VDD.t28 VDD.n1893 468.033
R10916 VDD.n2235 VDD.n2213 468.033
R10917 VDD.t103 VDD.n2214 468.033
R10918 VDD.n2493 VDD.n2471 468.033
R10919 VDD.t471 VDD.n2472 468.033
R10920 VDD.n2751 VDD.n2729 468.033
R10921 VDD.t184 VDD.n2730 468.033
R10922 VDD.n3009 VDD.n2987 468.033
R10923 VDD.t488 VDD.n2988 468.033
R10924 VDD.n3267 VDD.n3245 468.033
R10925 VDD.t234 VDD.n3246 468.033
R10926 VDD.n3525 VDD.n3503 468.033
R10927 VDD.t18 VDD.n3504 468.033
R10928 VDD.n5845 VDD.n5823 468.033
R10929 VDD.t746 VDD.n5824 468.033
R10930 VDD.n5591 VDD.n5569 468.033
R10931 VDD.t88 VDD.n5570 468.033
R10932 VDD.n3783 VDD.n3761 468.033
R10933 VDD.t82 VDD.n3762 468.033
R10934 VDD.n4041 VDD.n4019 468.033
R10935 VDD.t409 VDD.n4020 468.033
R10936 VDD.n4299 VDD.n4277 468.033
R10937 VDD.t727 VDD.n4278 468.033
R10938 VDD.n4557 VDD.n4535 468.033
R10939 VDD.t122 VDD.n4536 468.033
R10940 VDD.n4815 VDD.n4793 468.033
R10941 VDD.t484 VDD.n4794 468.033
R10942 VDD.n5073 VDD.n5051 468.033
R10943 VDD.t14 VDD.n5052 468.033
R10944 VDD.n5331 VDD.n5309 468.033
R10945 VDD.t119 VDD.n5310 468.033
R10946 VDD.n1933 VDD.n1925 459.009
R10947 VDD.n1935 VDD.n1932 437.647
R10948 VDD.n1974 VDD.n1928 430.589
R10949 VDD.n1962 VDD.n1940 430.589
R10950 VDD.n483 VDD.n482 425.228
R10951 VDD.n81 VDD.n80 425.228
R10952 VDD VDD.t834 421.082
R10953 VDD.n1948 VDD.n1938 420
R10954 VDD.n407 VDD.t629 396.079
R10955 VDD.n1565 VDD.t557 396.079
R10956 VDD.n9 VDD.t809 382.793
R10957 VDD.n465 VDD.t802 382.793
R10958 VDD.n412 VDD.t812 382.793
R10959 VDD.n411 VDD.t799 382.793
R10960 VDD.n393 VDD.t798 382.793
R10961 VDD.n63 VDD.t771 382.793
R10962 VDD.n1153 VDD.t779 382.793
R10963 VDD.n1570 VDD.t765 382.793
R10964 VDD.n1569 VDD.t760 382.793
R10965 VDD.n1551 VDD.t758 382.793
R10966 VDD.n805 VDD.t1038 382.793
R10967 VDD.n1188 VDD.t833 382.793
R10968 VDD VDD.t1340 374.711
R10969 VDD VDD.t550 374.711
R10970 VDD VDD.t1391 374.711
R10971 VDD VDD.t741 374.711
R10972 VDD VDD.t179 374.711
R10973 VDD VDD.t878 374.711
R10974 VDD.n1709 VDD.n1680 370.589
R10975 VDD.n1759 VDD.n1714 370.589
R10976 VDD.n2058 VDD.n2029 370.589
R10977 VDD.n2108 VDD.n2063 370.589
R10978 VDD.n2288 VDD.n2259 370.589
R10979 VDD.n2338 VDD.n2293 370.589
R10980 VDD.n2546 VDD.n2517 370.589
R10981 VDD.n2596 VDD.n2551 370.589
R10982 VDD.n2804 VDD.n2775 370.589
R10983 VDD.n2854 VDD.n2809 370.589
R10984 VDD.n3062 VDD.n3033 370.589
R10985 VDD.n3112 VDD.n3067 370.589
R10986 VDD.n3320 VDD.n3291 370.589
R10987 VDD.n3370 VDD.n3325 370.589
R10988 VDD.n5643 VDD.n5614 370.589
R10989 VDD.n5693 VDD.n5648 370.589
R10990 VDD.n5389 VDD.n5360 370.589
R10991 VDD.n5439 VDD.n5394 370.589
R10992 VDD.n3578 VDD.n3549 370.589
R10993 VDD.n3628 VDD.n3583 370.589
R10994 VDD.n3836 VDD.n3807 370.589
R10995 VDD.n3886 VDD.n3841 370.589
R10996 VDD.n4094 VDD.n4065 370.589
R10997 VDD.n4144 VDD.n4099 370.589
R10998 VDD.n4352 VDD.n4323 370.589
R10999 VDD.n4402 VDD.n4357 370.589
R11000 VDD.n4610 VDD.n4581 370.589
R11001 VDD.n4660 VDD.n4615 370.589
R11002 VDD.n4868 VDD.n4839 370.589
R11003 VDD.n4918 VDD.n4873 370.589
R11004 VDD.n5126 VDD.n5097 370.589
R11005 VDD.n5176 VDD.n5131 370.589
R11006 VDD.n12 VDD.t217 370.341
R11007 VDD.n473 VDD.t803 370.341
R11008 VDD.n445 VDD.t1033 370.341
R11009 VDD.n446 VDD.t704 370.341
R11010 VDD.n71 VDD.t773 370.341
R11011 VDD.n42 VDD.t1489 370.341
R11012 VDD.n43 VDD.t147 370.341
R11013 VDD.n1156 VDD.t881 370.341
R11014 VDD VDD.t421 370.303
R11015 VDD VDD.t824 370.303
R11016 VDD.t388 VDD.t642 333.365
R11017 VDD.t388 VDD.t1359 333.365
R11018 VDD.t228 VDD.t243 333.365
R11019 VDD.t228 VDD.t1493 333.365
R11020 VDD.t181 VDD.t624 333.365
R11021 VDD.t181 VDD.t222 333.365
R11022 VDD.t713 VDD.t842 333.365
R11023 VDD.t713 VDD.t55 333.365
R11024 VDD.t542 VDD.t134 333.365
R11025 VDD.t542 VDD.t595 333.365
R11026 VDD.t647 VDD.t473 333.365
R11027 VDD.t647 VDD.t41 333.365
R11028 VDD.t30 VDD.t1331 333.365
R11029 VDD.t30 VDD.t731 333.365
R11030 VDD.t870 VDD.t613 333.365
R11031 VDD.t870 VDD.t164 333.365
R11032 VDD.t709 VDD.t6 333.365
R11033 VDD.t709 VDD.t517 333.365
R11034 VDD.t214 VDD.t631 333.365
R11035 VDD.t214 VDD.t194 333.365
R11036 VDD.t1027 VDD.t1386 333.365
R11037 VDD.t1027 VDD.t173 333.365
R11038 VDD.t423 VDD.t888 333.365
R11039 VDD.t423 VDD.t92 333.365
R11040 VDD.t1031 VDD.t126 333.365
R11041 VDD.t1031 VDD.t497 333.365
R11042 VDD.t402 VDD.t72 333.365
R11043 VDD.t402 VDD.t587 333.365
R11044 VDD.t532 VDD.t783 333.365
R11045 VDD.t532 VDD.t579 333.365
R11046 VDD.t381 VDD.t1374 333.365
R11047 VDD.t381 VDD.t857 333.365
R11048 VDD VDD.t139 331.981
R11049 VDD VDD.t392 331.981
R11050 VDD.n1634 VDD.t780 330.12
R11051 VDD.n1635 VDD.t761 330.002
R11052 VDD.n1541 VDD 323.514
R11053 VDD.n1643 VDD.t772 323.342
R11054 VDD.n34 VDD.t820 321.801
R11055 VDD.n1178 VDD.t1439 321.801
R11056 VDD.n476 VDD.n475 318.678
R11057 VDD.n74 VDD.n73 318.678
R11058 VDD.n511 VDD.t1430 318.108
R11059 VDD.n109 VDD.t606 318.108
R11060 VDD VDD.t218 313.839
R11061 VDD VDD.t1367 313.839
R11062 VDD VDD.t705 313.839
R11063 VDD.n8 VDD.n7 307.24
R11064 VDD.n472 VDD.n471 307.24
R11065 VDD.n442 VDD.n441 307.24
R11066 VDD.n444 VDD.n443 307.24
R11067 VDD.n70 VDD.n69 307.24
R11068 VDD.n39 VDD.n38 307.24
R11069 VDD.n41 VDD.n40 307.24
R11070 VDD.n1152 VDD.n1151 307.24
R11071 VDD.t388 VDD.n1678 298.82
R11072 VDD.t388 VDD.n1712 298.82
R11073 VDD.t228 VDD.n2027 298.82
R11074 VDD.t228 VDD.n2061 298.82
R11075 VDD.t181 VDD.n2257 298.82
R11076 VDD.t181 VDD.n2291 298.82
R11077 VDD.t713 VDD.n2515 298.82
R11078 VDD.t713 VDD.n2549 298.82
R11079 VDD.t542 VDD.n2773 298.82
R11080 VDD.t542 VDD.n2807 298.82
R11081 VDD.t647 VDD.n3031 298.82
R11082 VDD.t647 VDD.n3065 298.82
R11083 VDD.t30 VDD.n3289 298.82
R11084 VDD.t30 VDD.n3323 298.82
R11085 VDD.t870 VDD.n5612 298.82
R11086 VDD.t870 VDD.n5646 298.82
R11087 VDD.t709 VDD.n5358 298.82
R11088 VDD.t709 VDD.n5392 298.82
R11089 VDD.t214 VDD.n3547 298.82
R11090 VDD.t214 VDD.n3581 298.82
R11091 VDD.t1027 VDD.n3805 298.82
R11092 VDD.t1027 VDD.n3839 298.82
R11093 VDD.t423 VDD.n4063 298.82
R11094 VDD.t423 VDD.n4097 298.82
R11095 VDD.t1031 VDD.n4321 298.82
R11096 VDD.t1031 VDD.n4355 298.82
R11097 VDD.t402 VDD.n4579 298.82
R11098 VDD.t402 VDD.n4613 298.82
R11099 VDD.t532 VDD.n4837 298.82
R11100 VDD.t532 VDD.n4871 298.82
R11101 VDD.t381 VDD.n5095 298.82
R11102 VDD.t381 VDD.n5129 298.82
R11103 VDD.n1912 VDD.n1897 273.695
R11104 VDD.n1912 VDD.n1911 273.695
R11105 VDD.n1877 VDD.n1824 273.695
R11106 VDD.n1824 VDD.n1822 273.695
R11107 VDD.n1861 VDD.n1860 273.695
R11108 VDD.n1865 VDD.n1861 273.695
R11109 VDD.n2182 VDD.n2181 273.695
R11110 VDD.n2186 VDD.n2182 273.695
R11111 VDD.n2198 VDD.n2145 273.695
R11112 VDD.n2145 VDD.n2143 273.695
R11113 VDD.n2233 VDD.n2218 273.695
R11114 VDD.n2233 VDD.n2232 273.695
R11115 VDD.n2440 VDD.n2439 273.695
R11116 VDD.n2444 VDD.n2440 273.695
R11117 VDD.n2456 VDD.n2403 273.695
R11118 VDD.n2403 VDD.n2401 273.695
R11119 VDD.n2491 VDD.n2476 273.695
R11120 VDD.n2491 VDD.n2490 273.695
R11121 VDD.n2698 VDD.n2697 273.695
R11122 VDD.n2702 VDD.n2698 273.695
R11123 VDD.n2714 VDD.n2661 273.695
R11124 VDD.n2661 VDD.n2659 273.695
R11125 VDD.n2749 VDD.n2734 273.695
R11126 VDD.n2749 VDD.n2748 273.695
R11127 VDD.n2956 VDD.n2955 273.695
R11128 VDD.n2960 VDD.n2956 273.695
R11129 VDD.n2972 VDD.n2919 273.695
R11130 VDD.n2919 VDD.n2917 273.695
R11131 VDD.n3007 VDD.n2992 273.695
R11132 VDD.n3007 VDD.n3006 273.695
R11133 VDD.n3214 VDD.n3213 273.695
R11134 VDD.n3218 VDD.n3214 273.695
R11135 VDD.n3230 VDD.n3177 273.695
R11136 VDD.n3177 VDD.n3175 273.695
R11137 VDD.n3265 VDD.n3250 273.695
R11138 VDD.n3265 VDD.n3264 273.695
R11139 VDD.n3472 VDD.n3471 273.695
R11140 VDD.n3476 VDD.n3472 273.695
R11141 VDD.n3488 VDD.n3435 273.695
R11142 VDD.n3435 VDD.n3433 273.695
R11143 VDD.n3523 VDD.n3508 273.695
R11144 VDD.n3523 VDD.n3522 273.695
R11145 VDD.n5792 VDD.n5791 273.695
R11146 VDD.n5796 VDD.n5792 273.695
R11147 VDD.n5808 VDD.n5755 273.695
R11148 VDD.n5755 VDD.n5753 273.695
R11149 VDD.n5843 VDD.n5828 273.695
R11150 VDD.n5843 VDD.n5842 273.695
R11151 VDD.n5538 VDD.n5537 273.695
R11152 VDD.n5542 VDD.n5538 273.695
R11153 VDD.n5554 VDD.n5501 273.695
R11154 VDD.n5501 VDD.n5499 273.695
R11155 VDD.n5589 VDD.n5574 273.695
R11156 VDD.n5589 VDD.n5588 273.695
R11157 VDD.n3730 VDD.n3729 273.695
R11158 VDD.n3734 VDD.n3730 273.695
R11159 VDD.n3746 VDD.n3693 273.695
R11160 VDD.n3693 VDD.n3691 273.695
R11161 VDD.n3781 VDD.n3766 273.695
R11162 VDD.n3781 VDD.n3780 273.695
R11163 VDD.n3988 VDD.n3987 273.695
R11164 VDD.n3992 VDD.n3988 273.695
R11165 VDD.n4004 VDD.n3951 273.695
R11166 VDD.n3951 VDD.n3949 273.695
R11167 VDD.n4039 VDD.n4024 273.695
R11168 VDD.n4039 VDD.n4038 273.695
R11169 VDD.n4246 VDD.n4245 273.695
R11170 VDD.n4250 VDD.n4246 273.695
R11171 VDD.n4262 VDD.n4209 273.695
R11172 VDD.n4209 VDD.n4207 273.695
R11173 VDD.n4297 VDD.n4282 273.695
R11174 VDD.n4297 VDD.n4296 273.695
R11175 VDD.n4504 VDD.n4503 273.695
R11176 VDD.n4508 VDD.n4504 273.695
R11177 VDD.n4520 VDD.n4467 273.695
R11178 VDD.n4467 VDD.n4465 273.695
R11179 VDD.n4555 VDD.n4540 273.695
R11180 VDD.n4555 VDD.n4554 273.695
R11181 VDD.n4762 VDD.n4761 273.695
R11182 VDD.n4766 VDD.n4762 273.695
R11183 VDD.n4778 VDD.n4725 273.695
R11184 VDD.n4725 VDD.n4723 273.695
R11185 VDD.n4813 VDD.n4798 273.695
R11186 VDD.n4813 VDD.n4812 273.695
R11187 VDD.n5020 VDD.n5019 273.695
R11188 VDD.n5024 VDD.n5020 273.695
R11189 VDD.n5036 VDD.n4983 273.695
R11190 VDD.n4983 VDD.n4981 273.695
R11191 VDD.n5071 VDD.n5056 273.695
R11192 VDD.n5071 VDD.n5070 273.695
R11193 VDD.n5278 VDD.n5277 273.695
R11194 VDD.n5282 VDD.n5278 273.695
R11195 VDD.n5294 VDD.n5241 273.695
R11196 VDD.n5241 VDD.n5239 273.695
R11197 VDD.n5329 VDD.n5314 273.695
R11198 VDD.n5329 VDD.n5328 273.695
R11199 VDD.n1616 VDD.t774 260.435
R11200 VDD.n1624 VDD.t756 256.07
R11201 VDD.n1627 VDD.t759 256.07
R11202 VDD.n1629 VDD.t763 256.07
R11203 VDD.n1632 VDD.t777 256.07
R11204 VDD.n1649 VDD.t769 251.637
R11205 VDD.t139 VDD.t810 246.023
R11206 VDD.t392 VDD.t781 246.023
R11207 VDD VDD.t21 241.819
R11208 VDD VDD.t751 241.819
R11209 VDD.t804 VDD 233.643
R11210 VDD.t1340 VDD 233.643
R11211 VDD.t550 VDD 233.643
R11212 VDD.t421 VDD 233.643
R11213 VDD.t1391 VDD 233.643
R11214 VDD.t767 VDD 233.643
R11215 VDD.t741 VDD 233.643
R11216 VDD.t179 VDD 233.643
R11217 VDD.t824 VDD 233.643
R11218 VDD.t878 VDD 233.643
R11219 VDD.n1605 VDD.t766 229.433
R11220 VDD.t1063 VDD 227.321
R11221 VDD VDD.t1051 227.321
R11222 VDD.t1129 VDD 227.321
R11223 VDD.t1462 VDD 227.321
R11224 VDD.t934 VDD 227.321
R11225 VDD VDD.t922 227.321
R11226 VDD.t1002 VDD 227.321
R11227 VDD.t1416 VDD 227.321
R11228 VDD.t257 VDD 227.321
R11229 VDD VDD.t373 227.321
R11230 VDD.t323 VDD 227.321
R11231 VDD.t437 VDD 227.321
R11232 VDD.t566 VDD 225.625
R11233 VDD.t51 VDD 225.625
R11234 VDD.t64 VDD 225.625
R11235 VDD.n1909 VDD.n1908 213.083
R11236 VDD.n1910 VDD.n1909 213.083
R11237 VDD.n1867 VDD.n1852 213.083
R11238 VDD.n1867 VDD.n1866 213.083
R11239 VDD.n2188 VDD.n2173 213.083
R11240 VDD.n2188 VDD.n2187 213.083
R11241 VDD.n2230 VDD.n2229 213.083
R11242 VDD.n2231 VDD.n2230 213.083
R11243 VDD.n2446 VDD.n2431 213.083
R11244 VDD.n2446 VDD.n2445 213.083
R11245 VDD.n2488 VDD.n2487 213.083
R11246 VDD.n2489 VDD.n2488 213.083
R11247 VDD.n2704 VDD.n2689 213.083
R11248 VDD.n2704 VDD.n2703 213.083
R11249 VDD.n2746 VDD.n2745 213.083
R11250 VDD.n2747 VDD.n2746 213.083
R11251 VDD.n2962 VDD.n2947 213.083
R11252 VDD.n2962 VDD.n2961 213.083
R11253 VDD.n3004 VDD.n3003 213.083
R11254 VDD.n3005 VDD.n3004 213.083
R11255 VDD.n3220 VDD.n3205 213.083
R11256 VDD.n3220 VDD.n3219 213.083
R11257 VDD.n3262 VDD.n3261 213.083
R11258 VDD.n3263 VDD.n3262 213.083
R11259 VDD.n3478 VDD.n3463 213.083
R11260 VDD.n3478 VDD.n3477 213.083
R11261 VDD.n3520 VDD.n3519 213.083
R11262 VDD.n3521 VDD.n3520 213.083
R11263 VDD.n5798 VDD.n5783 213.083
R11264 VDD.n5798 VDD.n5797 213.083
R11265 VDD.n5840 VDD.n5839 213.083
R11266 VDD.n5841 VDD.n5840 213.083
R11267 VDD.n5544 VDD.n5529 213.083
R11268 VDD.n5544 VDD.n5543 213.083
R11269 VDD.n5586 VDD.n5585 213.083
R11270 VDD.n5587 VDD.n5586 213.083
R11271 VDD.n3736 VDD.n3721 213.083
R11272 VDD.n3736 VDD.n3735 213.083
R11273 VDD.n3778 VDD.n3777 213.083
R11274 VDD.n3779 VDD.n3778 213.083
R11275 VDD.n3994 VDD.n3979 213.083
R11276 VDD.n3994 VDD.n3993 213.083
R11277 VDD.n4036 VDD.n4035 213.083
R11278 VDD.n4037 VDD.n4036 213.083
R11279 VDD.n4252 VDD.n4237 213.083
R11280 VDD.n4252 VDD.n4251 213.083
R11281 VDD.n4294 VDD.n4293 213.083
R11282 VDD.n4295 VDD.n4294 213.083
R11283 VDD.n4510 VDD.n4495 213.083
R11284 VDD.n4510 VDD.n4509 213.083
R11285 VDD.n4552 VDD.n4551 213.083
R11286 VDD.n4553 VDD.n4552 213.083
R11287 VDD.n4768 VDD.n4753 213.083
R11288 VDD.n4768 VDD.n4767 213.083
R11289 VDD.n4810 VDD.n4809 213.083
R11290 VDD.n4811 VDD.n4810 213.083
R11291 VDD.n5026 VDD.n5011 213.083
R11292 VDD.n5026 VDD.n5025 213.083
R11293 VDD.n5068 VDD.n5067 213.083
R11294 VDD.n5069 VDD.n5068 213.083
R11295 VDD.n5284 VDD.n5269 213.083
R11296 VDD.n5284 VDD.n5283 213.083
R11297 VDD.n5326 VDD.n5325 213.083
R11298 VDD.n5327 VDD.n5326 213.083
R11299 VDD.n531 VDD.t1062 204.903
R11300 VDD.n881 VDD.t933 204.903
R11301 VDD.n130 VDD.t256 204.903
R11302 VDD.n1249 VDD.t1320 204.9
R11303 VDD.n1634 VDD.t1509 201.587
R11304 VDD.n542 VDD.t1064 201.012
R11305 VDD.n621 VDD.t1052 201.012
R11306 VDD.n517 VDD.t1130 201.012
R11307 VDD.n520 VDD.t1463 201.012
R11308 VDD.n892 VDD.t935 201.012
R11309 VDD.n971 VDD.t923 201.012
R11310 VDD.n867 VDD.t1003 201.012
R11311 VDD.n870 VDD.t1417 201.012
R11312 VDD.n141 VDD.t258 201.012
R11313 VDD.n220 VDD.t374 201.012
R11314 VDD.n116 VDD.t324 201.012
R11315 VDD.n119 VDD.t438 201.012
R11316 VDD.n1313 VDD.t1226 201.012
R11317 VDD.n1342 VDD.t692 201.012
R11318 VDD.n1263 VDD.t1208 201.012
R11319 VDD.n1260 VDD.t1306 201.012
R11320 VDD.n1635 VDD.t1507 200.782
R11321 VDD.n1643 VDD.t1503 194.809
R11322 VDD.n1901 VDD.n1893 189.304
R11323 VDD.n2222 VDD.n2214 189.304
R11324 VDD.n2480 VDD.n2472 189.304
R11325 VDD.n2738 VDD.n2730 189.304
R11326 VDD.n2996 VDD.n2988 189.304
R11327 VDD.n3254 VDD.n3246 189.304
R11328 VDD.n3512 VDD.n3504 189.304
R11329 VDD.n5832 VDD.n5824 189.304
R11330 VDD.n5578 VDD.n5570 189.304
R11331 VDD.n3770 VDD.n3762 189.304
R11332 VDD.n4028 VDD.n4020 189.304
R11333 VDD.n4286 VDD.n4278 189.304
R11334 VDD.n4544 VDD.n4536 189.304
R11335 VDD.n4802 VDD.n4794 189.304
R11336 VDD.n5060 VDD.n5052 189.304
R11337 VDD.n5318 VDD.n5310 189.304
R11338 VDD.n1954 VDD.n1939 185
R11339 VDD.n1900 VDD.n1898 185
R11340 VDD.n1900 VDD.n1893 185
R11341 VDD.n1890 VDD.n1888 185
R11342 VDD.n1892 VDD.n1890 185
R11343 VDD.n1697 VDD.n1682 185
R11344 VDD.n2046 VDD.n2031 185
R11345 VDD.n2221 VDD.n2219 185
R11346 VDD.n2221 VDD.n2214 185
R11347 VDD.n2211 VDD.n2209 185
R11348 VDD.n2213 VDD.n2211 185
R11349 VDD.n2276 VDD.n2261 185
R11350 VDD.n2479 VDD.n2477 185
R11351 VDD.n2479 VDD.n2472 185
R11352 VDD.n2469 VDD.n2467 185
R11353 VDD.n2471 VDD.n2469 185
R11354 VDD.n2534 VDD.n2519 185
R11355 VDD.n2737 VDD.n2735 185
R11356 VDD.n2737 VDD.n2730 185
R11357 VDD.n2727 VDD.n2725 185
R11358 VDD.n2729 VDD.n2727 185
R11359 VDD.n2792 VDD.n2777 185
R11360 VDD.n2995 VDD.n2993 185
R11361 VDD.n2995 VDD.n2988 185
R11362 VDD.n2985 VDD.n2983 185
R11363 VDD.n2987 VDD.n2985 185
R11364 VDD.n3050 VDD.n3035 185
R11365 VDD.n3253 VDD.n3251 185
R11366 VDD.n3253 VDD.n3246 185
R11367 VDD.n3243 VDD.n3241 185
R11368 VDD.n3245 VDD.n3243 185
R11369 VDD.n3308 VDD.n3293 185
R11370 VDD.n3511 VDD.n3509 185
R11371 VDD.n3511 VDD.n3504 185
R11372 VDD.n3501 VDD.n3499 185
R11373 VDD.n3503 VDD.n3501 185
R11374 VDD.n5631 VDD.n5616 185
R11375 VDD.n5831 VDD.n5829 185
R11376 VDD.n5831 VDD.n5824 185
R11377 VDD.n5821 VDD.n5819 185
R11378 VDD.n5823 VDD.n5821 185
R11379 VDD.n5377 VDD.n5362 185
R11380 VDD.n5577 VDD.n5575 185
R11381 VDD.n5577 VDD.n5570 185
R11382 VDD.n5567 VDD.n5565 185
R11383 VDD.n5569 VDD.n5567 185
R11384 VDD.n3566 VDD.n3551 185
R11385 VDD.n3769 VDD.n3767 185
R11386 VDD.n3769 VDD.n3762 185
R11387 VDD.n3759 VDD.n3757 185
R11388 VDD.n3761 VDD.n3759 185
R11389 VDD.n3824 VDD.n3809 185
R11390 VDD.n4027 VDD.n4025 185
R11391 VDD.n4027 VDD.n4020 185
R11392 VDD.n4017 VDD.n4015 185
R11393 VDD.n4019 VDD.n4017 185
R11394 VDD.n4082 VDD.n4067 185
R11395 VDD.n4285 VDD.n4283 185
R11396 VDD.n4285 VDD.n4278 185
R11397 VDD.n4275 VDD.n4273 185
R11398 VDD.n4277 VDD.n4275 185
R11399 VDD.n4340 VDD.n4325 185
R11400 VDD.n4543 VDD.n4541 185
R11401 VDD.n4543 VDD.n4536 185
R11402 VDD.n4533 VDD.n4531 185
R11403 VDD.n4535 VDD.n4533 185
R11404 VDD.n4598 VDD.n4583 185
R11405 VDD.n4801 VDD.n4799 185
R11406 VDD.n4801 VDD.n4794 185
R11407 VDD.n4791 VDD.n4789 185
R11408 VDD.n4793 VDD.n4791 185
R11409 VDD.n4856 VDD.n4841 185
R11410 VDD.n5059 VDD.n5057 185
R11411 VDD.n5059 VDD.n5052 185
R11412 VDD.n5049 VDD.n5047 185
R11413 VDD.n5051 VDD.n5049 185
R11414 VDD.n5114 VDD.n5099 185
R11415 VDD.n5317 VDD.n5315 185
R11416 VDD.n5317 VDD.n5310 185
R11417 VDD.n5307 VDD.n5305 185
R11418 VDD.n5309 VDD.n5307 185
R11419 VDD.n1863 VDD.n1849 183.496
R11420 VDD.n2184 VDD.n2170 183.496
R11421 VDD.n2442 VDD.n2428 183.496
R11422 VDD.n2700 VDD.n2686 183.496
R11423 VDD.n2958 VDD.n2944 183.496
R11424 VDD.n3216 VDD.n3202 183.496
R11425 VDD.n3474 VDD.n3460 183.496
R11426 VDD.n5794 VDD.n5780 183.496
R11427 VDD.n5540 VDD.n5526 183.496
R11428 VDD.n3732 VDD.n3718 183.496
R11429 VDD.n3990 VDD.n3976 183.496
R11430 VDD.n4248 VDD.n4234 183.496
R11431 VDD.n4506 VDD.n4492 183.496
R11432 VDD.n4764 VDD.n4750 183.496
R11433 VDD.n5022 VDD.n5008 183.496
R11434 VDD.n5280 VDD.n5266 183.496
R11435 VDD.n807 VDD.n806 183.363
R11436 VDD.n1190 VDD.n1189 183.363
R11437 VDD.n1793 VDD.n1792 180.994
R11438 VDD.n1790 VDD.n1788 180.994
R11439 VDD.n2001 VDD.n2000 180.994
R11440 VDD.n1998 VDD.n1996 180.994
R11441 VDD.n2372 VDD.n2371 180.994
R11442 VDD.n2369 VDD.n2367 180.994
R11443 VDD.n2630 VDD.n2629 180.994
R11444 VDD.n2627 VDD.n2625 180.994
R11445 VDD.n2888 VDD.n2887 180.994
R11446 VDD.n2885 VDD.n2883 180.994
R11447 VDD.n3146 VDD.n3145 180.994
R11448 VDD.n3143 VDD.n3141 180.994
R11449 VDD.n3404 VDD.n3403 180.994
R11450 VDD.n3401 VDD.n3399 180.994
R11451 VDD.n5727 VDD.n5726 180.994
R11452 VDD.n5724 VDD.n5722 180.994
R11453 VDD.n5473 VDD.n5472 180.994
R11454 VDD.n5470 VDD.n5468 180.994
R11455 VDD.n3662 VDD.n3661 180.994
R11456 VDD.n3659 VDD.n3657 180.994
R11457 VDD.n3920 VDD.n3919 180.994
R11458 VDD.n3917 VDD.n3915 180.994
R11459 VDD.n4178 VDD.n4177 180.994
R11460 VDD.n4175 VDD.n4173 180.994
R11461 VDD.n4436 VDD.n4435 180.994
R11462 VDD.n4433 VDD.n4431 180.994
R11463 VDD.n4694 VDD.n4693 180.994
R11464 VDD.n4691 VDD.n4689 180.994
R11465 VDD.n4952 VDD.n4951 180.994
R11466 VDD.n4949 VDD.n4947 180.994
R11467 VDD.n5210 VDD.n5209 180.994
R11468 VDD.n5207 VDD.n5205 180.994
R11469 VDD.t512 VDD 179.821
R11470 VDD.t826 VDD 179.821
R11471 VDD.t396 VDD 179.821
R11472 VDD.t603 VDD 179.821
R11473 VDD.n265 VDD.t830 179.821
R11474 VDD.t830 VDD 179.821
R11475 VDD.t1343 VDD 179.821
R11476 VDD.n19 VDD.n5 179.131
R11477 VDD.n495 VDD.n494 179.131
R11478 VDD.n423 VDD.n422 179.131
R11479 VDD.n419 VDD.n418 179.131
R11480 VDD.n402 VDD.n401 179.131
R11481 VDD.n93 VDD.n92 179.131
R11482 VDD.n1163 VDD.n1149 179.131
R11483 VDD.n1581 VDD.n1580 179.131
R11484 VDD.n1577 VDD.n1576 179.131
R11485 VDD.n1560 VDD.n1559 179.131
R11486 VDD.t639 VDD.n1803 174.632
R11487 VDD.t245 VDD.n2011 174.632
R11488 VDD.t621 VDD.n2382 174.632
R11489 VDD.t844 VDD.n2640 174.632
R11490 VDD.t131 VDD.n2898 174.632
R11491 VDD.t475 VDD.n3156 174.632
R11492 VDD.t1333 VDD.n3414 174.632
R11493 VDD.t610 VDD.n5737 174.632
R11494 VDD.t4 VDD.n5483 174.632
R11495 VDD.t633 VDD.n3672 174.632
R11496 VDD.t1383 VDD.n3930 174.632
R11497 VDD.t885 VDD.n4188 174.632
R11498 VDD.t123 VDD.n4446 174.632
R11499 VDD.t74 VDD.n4704 174.632
R11500 VDD.t785 VDD.n4962 174.632
R11501 VDD.t1371 VDD.n5220 174.632
R11502 VDD.t1039 VDD 174.602
R11503 VDD.t203 VDD 174.602
R11504 VDD.n693 VDD.n692 174.595
R11505 VDD.n556 VDD.n555 174.595
R11506 VDD.n562 VDD.n561 174.595
R11507 VDD.n568 VDD.n567 174.595
R11508 VDD.n574 VDD.n573 174.595
R11509 VDD.n579 VDD.n578 174.595
R11510 VDD.n535 VDD.n534 174.595
R11511 VDD.n530 VDD.n529 174.595
R11512 VDD.n614 VDD.n613 174.595
R11513 VDD.n608 VDD.n607 174.595
R11514 VDD.n602 VDD.n601 174.595
R11515 VDD.n596 VDD.n595 174.595
R11516 VDD.n592 VDD.n591 174.595
R11517 VDD.n526 VDD.n525 174.595
R11518 VDD.n546 VDD.n545 174.595
R11519 VDD.n639 VDD.n638 174.595
R11520 VDD.n645 VDD.n644 174.595
R11521 VDD.n651 VDD.n650 174.595
R11522 VDD.n657 VDD.n656 174.595
R11523 VDD.n662 VDD.n661 174.595
R11524 VDD.n632 VDD.n631 174.595
R11525 VDD.n626 VDD.n625 174.595
R11526 VDD.n749 VDD.n748 174.595
R11527 VDD.n755 VDD.n754 174.595
R11528 VDD.n761 VDD.n760 174.595
R11529 VDD.n767 VDD.n766 174.595
R11530 VDD.n771 VDD.n770 174.595
R11531 VDD.n778 VDD.n777 174.595
R11532 VDD.n786 VDD.n785 174.595
R11533 VDD.n702 VDD.n701 174.595
R11534 VDD.n708 VDD.n707 174.595
R11535 VDD.n714 VDD.n713 174.595
R11536 VDD.n720 VDD.n719 174.595
R11537 VDD.n724 VDD.n723 174.595
R11538 VDD.n730 VDD.n729 174.595
R11539 VDD.n738 VDD.n737 174.595
R11540 VDD.n1043 VDD.n1042 174.595
R11541 VDD.n906 VDD.n905 174.595
R11542 VDD.n912 VDD.n911 174.595
R11543 VDD.n918 VDD.n917 174.595
R11544 VDD.n924 VDD.n923 174.595
R11545 VDD.n929 VDD.n928 174.595
R11546 VDD.n885 VDD.n884 174.595
R11547 VDD.n880 VDD.n879 174.595
R11548 VDD.n964 VDD.n963 174.595
R11549 VDD.n958 VDD.n957 174.595
R11550 VDD.n952 VDD.n951 174.595
R11551 VDD.n946 VDD.n945 174.595
R11552 VDD.n942 VDD.n941 174.595
R11553 VDD.n876 VDD.n875 174.595
R11554 VDD.n896 VDD.n895 174.595
R11555 VDD.n989 VDD.n988 174.595
R11556 VDD.n995 VDD.n994 174.595
R11557 VDD.n1001 VDD.n1000 174.595
R11558 VDD.n1007 VDD.n1006 174.595
R11559 VDD.n1012 VDD.n1011 174.595
R11560 VDD.n982 VDD.n981 174.595
R11561 VDD.n976 VDD.n975 174.595
R11562 VDD.n1099 VDD.n1098 174.595
R11563 VDD.n1105 VDD.n1104 174.595
R11564 VDD.n1111 VDD.n1110 174.595
R11565 VDD.n1117 VDD.n1116 174.595
R11566 VDD.n1121 VDD.n1120 174.595
R11567 VDD.n1128 VDD.n1127 174.595
R11568 VDD.n1136 VDD.n1135 174.595
R11569 VDD.n1052 VDD.n1051 174.595
R11570 VDD.n1058 VDD.n1057 174.595
R11571 VDD.n1064 VDD.n1063 174.595
R11572 VDD.n1070 VDD.n1069 174.595
R11573 VDD.n1074 VDD.n1073 174.595
R11574 VDD.n1080 VDD.n1079 174.595
R11575 VDD.n1088 VDD.n1087 174.595
R11576 VDD.n288 VDD.n287 174.595
R11577 VDD.n155 VDD.n154 174.595
R11578 VDD.n161 VDD.n160 174.595
R11579 VDD.n167 VDD.n166 174.595
R11580 VDD.n173 VDD.n172 174.595
R11581 VDD.n178 VDD.n177 174.595
R11582 VDD.n134 VDD.n133 174.595
R11583 VDD.n129 VDD.n128 174.595
R11584 VDD.n213 VDD.n212 174.595
R11585 VDD.n207 VDD.n206 174.595
R11586 VDD.n201 VDD.n200 174.595
R11587 VDD.n195 VDD.n194 174.595
R11588 VDD.n191 VDD.n190 174.595
R11589 VDD.n125 VDD.n124 174.595
R11590 VDD.n145 VDD.n144 174.595
R11591 VDD.n112 VDD.n111 174.595
R11592 VDD.n240 VDD.n239 174.595
R11593 VDD.n246 VDD.n245 174.595
R11594 VDD.n252 VDD.n251 174.595
R11595 VDD.n257 VDD.n256 174.595
R11596 VDD.n231 VDD.n230 174.595
R11597 VDD.n225 VDD.n224 174.595
R11598 VDD.n344 VDD.n343 174.595
R11599 VDD.n350 VDD.n349 174.595
R11600 VDD.n356 VDD.n355 174.595
R11601 VDD.n362 VDD.n361 174.595
R11602 VDD.n366 VDD.n365 174.595
R11603 VDD.n373 VDD.n372 174.595
R11604 VDD.n381 VDD.n380 174.595
R11605 VDD.n297 VDD.n296 174.595
R11606 VDD.n303 VDD.n302 174.595
R11607 VDD.n309 VDD.n308 174.595
R11608 VDD.n315 VDD.n314 174.595
R11609 VDD.n319 VDD.n318 174.595
R11610 VDD.n325 VDD.n324 174.595
R11611 VDD.n333 VDD.n332 174.595
R11612 VDD.n1353 VDD.n1352 174.595
R11613 VDD.n1335 VDD.n1334 174.595
R11614 VDD.n1329 VDD.n1328 174.595
R11615 VDD.n1322 VDD.n1321 174.595
R11616 VDD.n1435 VDD.n1434 174.595
R11617 VDD.n1439 VDD.n1438 174.595
R11618 VDD.n1445 VDD.n1444 174.595
R11619 VDD.n1451 VDD.n1450 174.595
R11620 VDD.n1379 VDD.n1378 174.595
R11621 VDD.n1385 VDD.n1384 174.595
R11622 VDD.n1391 VDD.n1390 174.595
R11623 VDD.n1403 VDD.n1402 174.595
R11624 VDD.n1408 VDD.n1407 174.595
R11625 VDD.n1414 VDD.n1413 174.595
R11626 VDD.n1420 VDD.n1419 174.595
R11627 VDD.n1306 VDD.n1305 174.595
R11628 VDD.n1299 VDD.n1298 174.595
R11629 VDD.n1293 VDD.n1292 174.595
R11630 VDD.n1268 VDD.n1267 174.595
R11631 VDD.n1272 VDD.n1271 174.595
R11632 VDD.n1278 VDD.n1277 174.595
R11633 VDD.n1265 VDD.n1264 174.595
R11634 VDD.n1465 VDD.n1464 174.595
R11635 VDD.n1471 VDD.n1470 174.595
R11636 VDD.n1477 VDD.n1476 174.595
R11637 VDD.n1483 VDD.n1482 174.595
R11638 VDD.n1487 VDD.n1486 174.595
R11639 VDD.n1493 VDD.n1492 174.595
R11640 VDD.n1499 VDD.n1498 174.595
R11641 VDD.n1515 VDD.n1514 174.595
R11642 VDD.n1521 VDD.n1520 174.595
R11643 VDD.n1257 VDD.n1256 174.595
R11644 VDD.n1531 VDD.n1530 174.595
R11645 VDD.n1535 VDD.n1534 174.595
R11646 VDD.n1253 VDD.n1252 174.595
R11647 VDD.n1248 VDD.n1247 174.595
R11648 VDD VDD.t1207 174.385
R11649 VDD VDD.t1225 174.385
R11650 VDD VDD.t659 173.083
R11651 VDD.n670 VDD.t512 173.036
R11652 VDD.n1020 VDD.t396 173.036
R11653 VDD.n1822 VDD.n1820 170.542
R11654 VDD.n2143 VDD.n2141 170.542
R11655 VDD.n2401 VDD.n2399 170.542
R11656 VDD.n2659 VDD.n2657 170.542
R11657 VDD.n2917 VDD.n2915 170.542
R11658 VDD.n3175 VDD.n3173 170.542
R11659 VDD.n3433 VDD.n3431 170.542
R11660 VDD.n5753 VDD.n5751 170.542
R11661 VDD.n5499 VDD.n5497 170.542
R11662 VDD.n3691 VDD.n3689 170.542
R11663 VDD.n3949 VDD.n3947 170.542
R11664 VDD.n4207 VDD.n4205 170.542
R11665 VDD.n4465 VDD.n4463 170.542
R11666 VDD.n4723 VDD.n4721 170.542
R11667 VDD.n4981 VDD.n4979 170.542
R11668 VDD.n5239 VDD.n5237 170.542
R11669 VDD.t468 VDD 170.478
R11670 VDD.t510 VDD 170.478
R11671 VDD VDD.n1428 169.179
R11672 VDD.n32 VDD.n31 169.107
R11673 VDD.n509 VDD.n508 169.107
R11674 VDD.n436 VDD.n435 169.107
R11675 VDD.n405 VDD.n404 169.107
R11676 VDD.n107 VDD.n106 169.107
R11677 VDD.n1176 VDD.n1175 169.107
R11678 VDD.n1594 VDD.n1593 169.107
R11679 VDD.n1563 VDD.n1562 169.107
R11680 VDD.n819 VDD.n800 169.107
R11681 VDD.n812 VDD.n803 169.107
R11682 VDD.n1202 VDD.n1183 169.107
R11683 VDD.n1195 VDD.n1186 169.107
R11684 VDD.n673 VDD.n672 169.017
R11685 VDD.n1023 VDD.n1022 169.017
R11686 VDD.n268 VDD.n267 169.017
R11687 VDD.n1645 VDD.t753 168.561
R11688 VDD.n1689 VDD.n1673 167.234
R11689 VDD.n2038 VDD.n2022 167.234
R11690 VDD.n2268 VDD.n2252 167.234
R11691 VDD.n2526 VDD.n2510 167.234
R11692 VDD.n2784 VDD.n2768 167.234
R11693 VDD.n3042 VDD.n3026 167.234
R11694 VDD.n3300 VDD.n3284 167.234
R11695 VDD.n5623 VDD.n5607 167.234
R11696 VDD.n5369 VDD.n5353 167.234
R11697 VDD.n3558 VDD.n3542 167.234
R11698 VDD.n3816 VDD.n3800 167.234
R11699 VDD.n4074 VDD.n4058 167.234
R11700 VDD.n4332 VDD.n4316 167.234
R11701 VDD.n4590 VDD.n4574 167.234
R11702 VDD.n4848 VDD.n4832 167.234
R11703 VDD.n5106 VDD.n5090 167.234
R11704 VDD.n1746 VDD.n1715 166.812
R11705 VDD.n2095 VDD.n2064 166.812
R11706 VDD.n2325 VDD.n2294 166.812
R11707 VDD.n2583 VDD.n2552 166.812
R11708 VDD.n2841 VDD.n2810 166.812
R11709 VDD.n3099 VDD.n3068 166.812
R11710 VDD.n3357 VDD.n3326 166.812
R11711 VDD.n5680 VDD.n5649 166.812
R11712 VDD.n5426 VDD.n5395 166.812
R11713 VDD.n3615 VDD.n3584 166.812
R11714 VDD.n3873 VDD.n3842 166.812
R11715 VDD.n4131 VDD.n4100 166.812
R11716 VDD.n4389 VDD.n4358 166.812
R11717 VDD.n4647 VDD.n4616 166.812
R11718 VDD.n4905 VDD.n4874 166.812
R11719 VDD.n5163 VDD.n5132 166.812
R11720 VDD.n1645 VDD.t1511 166.328
R11721 VDD.n1834 VDD.n1830 165.767
R11722 VDD.n1814 VDD.n1813 165.767
R11723 VDD.n2135 VDD.n2134 165.767
R11724 VDD.n2155 VDD.n2151 165.767
R11725 VDD.n2393 VDD.n2392 165.767
R11726 VDD.n2413 VDD.n2409 165.767
R11727 VDD.n2651 VDD.n2650 165.767
R11728 VDD.n2671 VDD.n2667 165.767
R11729 VDD.n2909 VDD.n2908 165.767
R11730 VDD.n2929 VDD.n2925 165.767
R11731 VDD.n3167 VDD.n3166 165.767
R11732 VDD.n3187 VDD.n3183 165.767
R11733 VDD.n3425 VDD.n3424 165.767
R11734 VDD.n3445 VDD.n3441 165.767
R11735 VDD.n5745 VDD.n5744 165.767
R11736 VDD.n5765 VDD.n5761 165.767
R11737 VDD.n5491 VDD.n5490 165.767
R11738 VDD.n5511 VDD.n5507 165.767
R11739 VDD.n3683 VDD.n3682 165.767
R11740 VDD.n3703 VDD.n3699 165.767
R11741 VDD.n3941 VDD.n3940 165.767
R11742 VDD.n3961 VDD.n3957 165.767
R11743 VDD.n4199 VDD.n4198 165.767
R11744 VDD.n4219 VDD.n4215 165.767
R11745 VDD.n4457 VDD.n4456 165.767
R11746 VDD.n4477 VDD.n4473 165.767
R11747 VDD.n4715 VDD.n4714 165.767
R11748 VDD.n4735 VDD.n4731 165.767
R11749 VDD.n4973 VDD.n4972 165.767
R11750 VDD.n4993 VDD.n4989 165.767
R11751 VDD.n5231 VDD.n5230 165.767
R11752 VDD.n5251 VDD.n5247 165.767
R11753 VDD.t218 VDD.t251 164.554
R11754 VDD.t1367 VDD.t822 164.554
R11755 VDD.t705 VDD.t398 164.554
R11756 VDD.n24 VDD.n1 164.215
R11757 VDD.n488 VDD.n468 164.215
R11758 VDD.n440 VDD.n439 164.215
R11759 VDD.n460 VDD.n459 164.215
R11760 VDD.n86 VDD.n66 164.215
R11761 VDD.n37 VDD.n36 164.215
R11762 VDD.n57 VDD.n56 164.215
R11763 VDD.n1168 VDD.n1145 164.215
R11764 VDD.n1699 VDD.n1682 161.506
R11765 VDD.n2048 VDD.n2031 161.506
R11766 VDD.n2278 VDD.n2261 161.506
R11767 VDD.n2536 VDD.n2519 161.506
R11768 VDD.n2794 VDD.n2777 161.506
R11769 VDD.n3052 VDD.n3035 161.506
R11770 VDD.n3310 VDD.n3293 161.506
R11771 VDD.n5633 VDD.n5616 161.506
R11772 VDD.n5379 VDD.n5362 161.506
R11773 VDD.n3568 VDD.n3551 161.506
R11774 VDD.n3826 VDD.n3809 161.506
R11775 VDD.n4084 VDD.n4067 161.506
R11776 VDD.n4342 VDD.n4325 161.506
R11777 VDD.n4600 VDD.n4583 161.506
R11778 VDD.n4858 VDD.n4841 161.506
R11779 VDD.n5116 VDD.n5099 161.506
R11780 VDD.n1741 VDD.n1728 159.143
R11781 VDD.n2090 VDD.n2077 159.143
R11782 VDD.n2320 VDD.n2307 159.143
R11783 VDD.n2578 VDD.n2565 159.143
R11784 VDD.n2836 VDD.n2823 159.143
R11785 VDD.n3094 VDD.n3081 159.143
R11786 VDD.n3352 VDD.n3339 159.143
R11787 VDD.n5675 VDD.n5662 159.143
R11788 VDD.n5421 VDD.n5408 159.143
R11789 VDD.n3610 VDD.n3597 159.143
R11790 VDD.n3868 VDD.n3855 159.143
R11791 VDD.n4126 VDD.n4113 159.143
R11792 VDD.n4384 VDD.n4371 159.143
R11793 VDD.n4642 VDD.n4629 159.143
R11794 VDD.n4900 VDD.n4887 159.143
R11795 VDD.n5158 VDD.n5145 159.143
R11796 VDD.n1905 VDD.n1892 159.108
R11797 VDD.n1858 VDD.n1857 159.108
R11798 VDD.n2179 VDD.n2178 159.108
R11799 VDD.n2226 VDD.n2213 159.108
R11800 VDD.n2437 VDD.n2436 159.108
R11801 VDD.n2484 VDD.n2471 159.108
R11802 VDD.n2695 VDD.n2694 159.108
R11803 VDD.n2742 VDD.n2729 159.108
R11804 VDD.n2953 VDD.n2952 159.108
R11805 VDD.n3000 VDD.n2987 159.108
R11806 VDD.n3211 VDD.n3210 159.108
R11807 VDD.n3258 VDD.n3245 159.108
R11808 VDD.n3469 VDD.n3468 159.108
R11809 VDD.n3516 VDD.n3503 159.108
R11810 VDD.n5789 VDD.n5788 159.108
R11811 VDD.n5836 VDD.n5823 159.108
R11812 VDD.n5535 VDD.n5534 159.108
R11813 VDD.n5582 VDD.n5569 159.108
R11814 VDD.n3727 VDD.n3726 159.108
R11815 VDD.n3774 VDD.n3761 159.108
R11816 VDD.n3985 VDD.n3984 159.108
R11817 VDD.n4032 VDD.n4019 159.108
R11818 VDD.n4243 VDD.n4242 159.108
R11819 VDD.n4290 VDD.n4277 159.108
R11820 VDD.n4501 VDD.n4500 159.108
R11821 VDD.n4548 VDD.n4535 159.108
R11822 VDD.n4759 VDD.n4758 159.108
R11823 VDD.n4806 VDD.n4793 159.108
R11824 VDD.n5017 VDD.n5016 159.108
R11825 VDD.n5064 VDD.n5051 159.108
R11826 VDD.n5275 VDD.n5274 159.108
R11827 VDD.n5322 VDD.n5309 159.108
R11828 VDD.n1605 VDD.t1505 158.886
R11829 VDD.n1700 VDD.n1699 158.776
R11830 VDD.n2049 VDD.n2048 158.776
R11831 VDD.n2279 VDD.n2278 158.776
R11832 VDD.n2537 VDD.n2536 158.776
R11833 VDD.n2795 VDD.n2794 158.776
R11834 VDD.n3053 VDD.n3052 158.776
R11835 VDD.n3311 VDD.n3310 158.776
R11836 VDD.n5634 VDD.n5633 158.776
R11837 VDD.n5380 VDD.n5379 158.776
R11838 VDD.n3569 VDD.n3568 158.776
R11839 VDD.n3827 VDD.n3826 158.776
R11840 VDD.n4085 VDD.n4084 158.776
R11841 VDD.n4343 VDD.n4342 158.776
R11842 VDD.n4601 VDD.n4600 158.776
R11843 VDD.n4859 VDD.n4858 158.776
R11844 VDD.n5117 VDD.n5116 158.776
R11845 VDD.n541 VDD.t1144 158.117
R11846 VDD.n620 VDD.t1128 158.117
R11847 VDD.n516 VDD.t1108 158.117
R11848 VDD.n519 VDD.t1070 158.117
R11849 VDD.n522 VDD.t1453 158.117
R11850 VDD.n891 VDD.t1015 158.117
R11851 VDD.n970 VDD.t1001 158.117
R11852 VDD.n866 VDD.t979 158.117
R11853 VDD.n869 VDD.t941 158.117
R11854 VDD.n872 VDD.t1407 158.117
R11855 VDD.n140 VDD.t338 158.117
R11856 VDD.n219 VDD.t322 158.117
R11857 VDD.n115 VDD.t302 158.117
R11858 VDD.n118 VDD.t264 158.117
R11859 VDD.n121 VDD.t428 158.117
R11860 VDD.n1341 VDD.t1324 158.117
R11861 VDD.n1347 VDD.t670 158.117
R11862 VDD.n1312 VDD.t1300 158.117
R11863 VDD.n1262 VDD.t1302 158.117
R11864 VDD.n1259 VDD.t1250 158.117
R11865 VDD.n671 VDD.t513 158.06
R11866 VDD.n1021 VDD.t397 158.06
R11867 VDD.n266 VDD.t831 158.06
R11868 VDD.n1362 VDD.t1499 158.06
R11869 VDD.n826 VDD.t1392 158.06
R11870 VDD.n825 VDD.t422 158.06
R11871 VDD.n824 VDD.t551 158.06
R11872 VDD.n823 VDD.t1341 158.06
R11873 VDD.n822 VDD.t805 158.06
R11874 VDD.n1542 VDD.t835 158.06
R11875 VDD.n1209 VDD.t879 158.06
R11876 VDD.n1208 VDD.t825 158.06
R11877 VDD.n1207 VDD.t180 158.06
R11878 VDD.n1206 VDD.t742 158.06
R11879 VDD.n1205 VDD.t768 158.06
R11880 VDD.n1616 VDD.t1508 156.403
R11881 VDD.t21 VDD.t526 155.456
R11882 VDD.t751 VDD.t1484 155.456
R11883 VDD.n1679 VDD.n1670 155.294
R11884 VDD.n2028 VDD.n2019 155.294
R11885 VDD.n2258 VDD.n2249 155.294
R11886 VDD.n2516 VDD.n2507 155.294
R11887 VDD.n2774 VDD.n2765 155.294
R11888 VDD.n3032 VDD.n3023 155.294
R11889 VDD.n3290 VDD.n3281 155.294
R11890 VDD.n5613 VDD.n5604 155.294
R11891 VDD.n5359 VDD.n5350 155.294
R11892 VDD.n3548 VDD.n3539 155.294
R11893 VDD.n3806 VDD.n3797 155.294
R11894 VDD.n4064 VDD.n4055 155.294
R11895 VDD.n4322 VDD.n4313 155.294
R11896 VDD.n4580 VDD.n4571 155.294
R11897 VDD.n4838 VDD.n4829 155.294
R11898 VDD.n5096 VDD.n5087 155.294
R11899 VDD.n1507 VDD.t1305 153.562
R11900 VDD VDD.t492 151.137
R11901 VDD VDD.t853 151.137
R11902 VDD.n1784 VDD.t1364 151.123
R11903 VDD.n1786 VDD.t640 151.123
R11904 VDD.n1992 VDD.t1491 151.123
R11905 VDD.n1994 VDD.t248 151.123
R11906 VDD.n2363 VDD.t221 151.123
R11907 VDD.n2365 VDD.t626 151.123
R11908 VDD.n2621 VDD.t58 151.123
R11909 VDD.n2623 VDD.t845 151.123
R11910 VDD.n2879 VDD.t594 151.123
R11911 VDD.n2881 VDD.t132 151.123
R11912 VDD.n3137 VDD.t40 151.123
R11913 VDD.n3139 VDD.t479 151.123
R11914 VDD.n3395 VDD.t730 151.123
R11915 VDD.n3397 VDD.t1334 151.123
R11916 VDD.n5718 VDD.t163 151.123
R11917 VDD.n5720 VDD.t611 151.123
R11918 VDD.n5464 VDD.t522 151.123
R11919 VDD.n5466 VDD.t8 151.123
R11920 VDD.n3653 VDD.t193 151.123
R11921 VDD.n3655 VDD.t634 151.123
R11922 VDD.n3911 VDD.t177 151.123
R11923 VDD.n3913 VDD.t1388 151.123
R11924 VDD.n4169 VDD.t97 151.123
R11925 VDD.n4171 VDD.t890 151.123
R11926 VDD.n4427 VDD.t496 151.123
R11927 VDD.n4429 VDD.t124 151.123
R11928 VDD.n4685 VDD.t586 151.123
R11929 VDD.n4687 VDD.t78 151.123
R11930 VDD.n4943 VDD.t578 151.123
R11931 VDD.n4945 VDD.t786 151.123
R11932 VDD.n5201 VDD.t856 151.123
R11933 VDD.n5203 VDD.t1372 151.123
R11934 VDD.n524 VDD.t565 151.123
R11935 VDD.n874 VDD.t50 151.123
R11936 VDD.n123 VDD.t71 151.123
R11937 VDD.n1357 VDD.t662 151.123
R11938 VDD.n1624 VDD.t1506 150.03
R11939 VDD.n1627 VDD.t1502 150.03
R11940 VDD.n1629 VDD.t1504 150.03
R11941 VDD.n1632 VDD.t1510 150.03
R11942 VDD.t806 VDD.t559 148.481
R11943 VDD.t775 VDD.t19 148.481
R11944 VDD.n1802 VDD.t1361 146.691
R11945 VDD.n2010 VDD.t1490 146.691
R11946 VDD.n2381 VDD.t220 146.691
R11947 VDD.n2639 VDD.t57 146.691
R11948 VDD.n2897 VDD.t593 146.691
R11949 VDD.n3155 VDD.t39 146.691
R11950 VDD.n3413 VDD.t729 146.691
R11951 VDD.n5736 VDD.t162 146.691
R11952 VDD.n5482 VDD.t519 146.691
R11953 VDD.n3671 VDD.t191 146.691
R11954 VDD.n3929 VDD.t171 146.691
R11955 VDD.n4187 VDD.t94 146.691
R11956 VDD.n4445 VDD.t495 146.691
R11957 VDD.n4703 VDD.t585 146.691
R11958 VDD.n4961 VDD.t577 146.691
R11959 VDD.n5219 VDD.t855 146.691
R11960 VDD.t820 VDD.t157 145.243
R11961 VDD.t1439 VDD.t1437 145.243
R11962 VDD.n1647 VDD.t1512 145.043
R11963 VDD.n1741 VDD.n1740 143.435
R11964 VDD.n2090 VDD.n2089 143.435
R11965 VDD.n2320 VDD.n2319 143.435
R11966 VDD.n2578 VDD.n2577 143.435
R11967 VDD.n2836 VDD.n2835 143.435
R11968 VDD.n3094 VDD.n3093 143.435
R11969 VDD.n3352 VDD.n3351 143.435
R11970 VDD.n5675 VDD.n5674 143.435
R11971 VDD.n5421 VDD.n5420 143.435
R11972 VDD.n3610 VDD.n3609 143.435
R11973 VDD.n3868 VDD.n3867 143.435
R11974 VDD.n4126 VDD.n4125 143.435
R11975 VDD.n4384 VDD.n4383 143.435
R11976 VDD.n4642 VDD.n4641 143.435
R11977 VDD.n4900 VDD.n4899 143.435
R11978 VDD.n5158 VDD.n5157 143.435
R11979 VDD.t629 VDD.t419 143.232
R11980 VDD.t557 VDD.t1192 143.232
R11981 VDD.t1087 VDD.t1061 142.5
R11982 VDD.t1173 VDD.t1087 142.5
R11983 VDD.t1065 VDD.t1173 142.5
R11984 VDD.t1057 VDD.t1065 142.5
R11985 VDD.t1079 VDD.t1057 142.5
R11986 VDD.t1047 VDD.t1105 142.5
R11987 VDD.t1083 VDD.t1047 142.5
R11988 VDD.t1153 VDD.t1083 142.5
R11989 VDD.t1049 VDD.t1153 142.5
R11990 VDD.t1073 VDD.t1049 142.5
R11991 VDD.t1137 VDD.t1073 142.5
R11992 VDD.t1167 VDD.t1137 142.5
R11993 VDD.t1099 VDD.t1167 142.5
R11994 VDD.t1143 VDD.t1099 142.5
R11995 VDD.t1131 VDD.t1063 142.5
R11996 VDD.t1157 VDD.t1131 142.5
R11997 VDD.t1055 VDD.t1157 142.5
R11998 VDD.t1111 VDD.t1055 142.5
R11999 VDD.t1145 VDD.t1077 142.5
R12000 VDD.t1077 VDD.t1115 142.5
R12001 VDD.t1115 VDD.t1149 142.5
R12002 VDD.t1149 VDD.t1085 142.5
R12003 VDD.t1085 VDD.t1165 142.5
R12004 VDD.t1165 VDD.t1097 142.5
R12005 VDD.t1097 VDD.t1123 142.5
R12006 VDD.t1123 VDD.t1171 142.5
R12007 VDD.t1171 VDD.t1103 142.5
R12008 VDD.t1103 VDD.t1127 142.5
R12009 VDD.t1051 VDD.t1109 142.5
R12010 VDD.t1109 VDD.t1139 142.5
R12011 VDD.t1139 VDD.t1075 142.5
R12012 VDD.t1075 VDD.t1161 142.5
R12013 VDD.t1161 VDD.t1071 142.5
R12014 VDD.t1163 VDD.t1135 142.5
R12015 VDD.t1093 VDD.t1163 142.5
R12016 VDD.t1119 VDD.t1093 142.5
R12017 VDD.t1151 VDD.t1119 142.5
R12018 VDD.t1095 VDD.t1151 142.5
R12019 VDD.t1121 VDD.t1095 142.5
R12020 VDD.t1067 VDD.t1121 142.5
R12021 VDD.t1089 VDD.t1067 142.5
R12022 VDD.t1107 VDD.t1089 142.5
R12023 VDD.t1155 VDD.t1129 142.5
R12024 VDD.t1053 VDD.t1155 142.5
R12025 VDD.t1133 VDD.t1053 142.5
R12026 VDD.t1091 VDD.t1159 142.5
R12027 VDD.t1113 VDD.t1091 142.5
R12028 VDD.t1147 VDD.t1113 142.5
R12029 VDD.t1081 VDD.t1147 142.5
R12030 VDD.t1117 VDD.t1081 142.5
R12031 VDD.t1059 VDD.t1117 142.5
R12032 VDD.t1141 VDD.t1059 142.5
R12033 VDD.t1169 VDD.t1141 142.5
R12034 VDD.t1101 VDD.t1169 142.5
R12035 VDD.t1125 VDD.t1101 142.5
R12036 VDD.t1069 VDD.t1125 142.5
R12037 VDD.t1476 VDD.t1462 142.5
R12038 VDD.t1464 VDD.t1456 142.5
R12039 VDD.t1474 VDD.t1464 142.5
R12040 VDD.t1470 VDD.t1474 142.5
R12041 VDD.t1478 VDD.t1470 142.5
R12042 VDD.t1458 VDD.t1478 142.5
R12043 VDD.t1472 VDD.t1458 142.5
R12044 VDD.t1480 VDD.t1472 142.5
R12045 VDD.t1460 VDD.t1480 142.5
R12046 VDD.t1466 VDD.t1460 142.5
R12047 VDD.t1450 VDD.t1466 142.5
R12048 VDD.t1454 VDD.t1450 142.5
R12049 VDD.t1468 VDD.t1454 142.5
R12050 VDD.t1452 VDD.t1468 142.5
R12051 VDD.t568 VDD.t566 142.5
R12052 VDD.t570 VDD.t568 142.5
R12053 VDD.t564 VDD.t570 142.5
R12054 VDD.t958 VDD.t932 142.5
R12055 VDD.t916 VDD.t958 142.5
R12056 VDD.t936 VDD.t916 142.5
R12057 VDD.t928 VDD.t936 142.5
R12058 VDD.t948 VDD.t928 142.5
R12059 VDD.t918 VDD.t976 142.5
R12060 VDD.t954 VDD.t918 142.5
R12061 VDD.t896 VDD.t954 142.5
R12062 VDD.t920 VDD.t896 142.5
R12063 VDD.t944 VDD.t920 142.5
R12064 VDD.t1008 VDD.t944 142.5
R12065 VDD.t910 VDD.t1008 142.5
R12066 VDD.t970 VDD.t910 142.5
R12067 VDD.t1014 VDD.t970 142.5
R12068 VDD.t982 VDD.t934 142.5
R12069 VDD.t900 VDD.t982 142.5
R12070 VDD.t926 VDD.t900 142.5
R12071 VDD.t984 VDD.t926 142.5
R12072 VDD.t1016 VDD.t950 142.5
R12073 VDD.t950 VDD.t988 142.5
R12074 VDD.t988 VDD.t1020 142.5
R12075 VDD.t1020 VDD.t956 142.5
R12076 VDD.t956 VDD.t908 142.5
R12077 VDD.t908 VDD.t968 142.5
R12078 VDD.t968 VDD.t996 142.5
R12079 VDD.t996 VDD.t914 142.5
R12080 VDD.t914 VDD.t974 142.5
R12081 VDD.t974 VDD.t1000 142.5
R12082 VDD.t922 VDD.t980 142.5
R12083 VDD.t980 VDD.t1010 142.5
R12084 VDD.t1010 VDD.t946 142.5
R12085 VDD.t946 VDD.t904 142.5
R12086 VDD.t904 VDD.t942 142.5
R12087 VDD.t906 VDD.t1006 142.5
R12088 VDD.t960 VDD.t906 142.5
R12089 VDD.t992 VDD.t960 142.5
R12090 VDD.t1022 VDD.t992 142.5
R12091 VDD.t966 VDD.t1022 142.5
R12092 VDD.t994 VDD.t966 142.5
R12093 VDD.t938 VDD.t994 142.5
R12094 VDD.t962 VDD.t938 142.5
R12095 VDD.t978 VDD.t962 142.5
R12096 VDD.t898 VDD.t1002 142.5
R12097 VDD.t924 VDD.t898 142.5
R12098 VDD.t1004 VDD.t924 142.5
R12099 VDD.t964 VDD.t902 142.5
R12100 VDD.t986 VDD.t964 142.5
R12101 VDD.t1018 VDD.t986 142.5
R12102 VDD.t952 VDD.t1018 142.5
R12103 VDD.t990 VDD.t952 142.5
R12104 VDD.t930 VDD.t990 142.5
R12105 VDD.t1012 VDD.t930 142.5
R12106 VDD.t912 VDD.t1012 142.5
R12107 VDD.t972 VDD.t912 142.5
R12108 VDD.t998 VDD.t972 142.5
R12109 VDD.t940 VDD.t998 142.5
R12110 VDD.t1398 VDD.t1416 142.5
R12111 VDD.t1418 VDD.t1410 142.5
R12112 VDD.t1428 VDD.t1418 142.5
R12113 VDD.t1424 VDD.t1428 142.5
R12114 VDD.t1400 VDD.t1424 142.5
R12115 VDD.t1412 VDD.t1400 142.5
R12116 VDD.t1426 VDD.t1412 142.5
R12117 VDD.t1402 VDD.t1426 142.5
R12118 VDD.t1414 VDD.t1402 142.5
R12119 VDD.t1420 VDD.t1414 142.5
R12120 VDD.t1404 VDD.t1420 142.5
R12121 VDD.t1408 VDD.t1404 142.5
R12122 VDD.t1422 VDD.t1408 142.5
R12123 VDD.t1406 VDD.t1422 142.5
R12124 VDD.t53 VDD.t51 142.5
R12125 VDD.t47 VDD.t53 142.5
R12126 VDD.t49 VDD.t47 142.5
R12127 VDD.t281 VDD.t255 142.5
R12128 VDD.t367 VDD.t281 142.5
R12129 VDD.t259 VDD.t367 142.5
R12130 VDD.t379 VDD.t259 142.5
R12131 VDD.t271 VDD.t379 142.5
R12132 VDD.t369 VDD.t299 142.5
R12133 VDD.t279 VDD.t369 142.5
R12134 VDD.t347 VDD.t279 142.5
R12135 VDD.t371 VDD.t347 142.5
R12136 VDD.t267 VDD.t371 142.5
R12137 VDD.t331 VDD.t267 142.5
R12138 VDD.t361 VDD.t331 142.5
R12139 VDD.t293 VDD.t361 142.5
R12140 VDD.t337 VDD.t293 142.5
R12141 VDD.t325 VDD.t257 142.5
R12142 VDD.t351 VDD.t325 142.5
R12143 VDD.t377 VDD.t351 142.5
R12144 VDD.t305 VDD.t377 142.5
R12145 VDD.t339 VDD.t273 142.5
R12146 VDD.t273 VDD.t309 142.5
R12147 VDD.t309 VDD.t343 142.5
R12148 VDD.t343 VDD.t277 142.5
R12149 VDD.t277 VDD.t359 142.5
R12150 VDD.t359 VDD.t291 142.5
R12151 VDD.t291 VDD.t317 142.5
R12152 VDD.t317 VDD.t365 142.5
R12153 VDD.t365 VDD.t297 142.5
R12154 VDD.t297 VDD.t321 142.5
R12155 VDD.t373 VDD.t303 142.5
R12156 VDD.t303 VDD.t333 142.5
R12157 VDD.t333 VDD.t269 142.5
R12158 VDD.t269 VDD.t355 142.5
R12159 VDD.t355 VDD.t265 142.5
R12160 VDD.t357 VDD.t329 142.5
R12161 VDD.t287 VDD.t357 142.5
R12162 VDD.t313 VDD.t287 142.5
R12163 VDD.t345 VDD.t313 142.5
R12164 VDD.t289 VDD.t345 142.5
R12165 VDD.t315 VDD.t289 142.5
R12166 VDD.t261 VDD.t315 142.5
R12167 VDD.t283 VDD.t261 142.5
R12168 VDD.t301 VDD.t283 142.5
R12169 VDD.t349 VDD.t323 142.5
R12170 VDD.t375 VDD.t349 142.5
R12171 VDD.t327 VDD.t375 142.5
R12172 VDD.t285 VDD.t353 142.5
R12173 VDD.t307 VDD.t285 142.5
R12174 VDD.t341 VDD.t307 142.5
R12175 VDD.t275 VDD.t341 142.5
R12176 VDD.t311 VDD.t275 142.5
R12177 VDD.t253 VDD.t311 142.5
R12178 VDD.t335 VDD.t253 142.5
R12179 VDD.t363 VDD.t335 142.5
R12180 VDD.t295 VDD.t363 142.5
R12181 VDD.t319 VDD.t295 142.5
R12182 VDD.t263 VDD.t319 142.5
R12183 VDD.t451 VDD.t437 142.5
R12184 VDD.t439 VDD.t431 142.5
R12185 VDD.t449 VDD.t439 142.5
R12186 VDD.t445 VDD.t449 142.5
R12187 VDD.t453 VDD.t445 142.5
R12188 VDD.t433 VDD.t453 142.5
R12189 VDD.t447 VDD.t433 142.5
R12190 VDD.t455 VDD.t447 142.5
R12191 VDD.t435 VDD.t455 142.5
R12192 VDD.t441 VDD.t435 142.5
R12193 VDD.t425 VDD.t441 142.5
R12194 VDD.t429 VDD.t425 142.5
R12195 VDD.t443 VDD.t429 142.5
R12196 VDD.t427 VDD.t443 142.5
R12197 VDD.t66 VDD.t64 142.5
R12198 VDD.t68 VDD.t66 142.5
R12199 VDD.t70 VDD.t68 142.5
R12200 VDD.t157 VDD.t867 142.279
R12201 VDD.t205 VDD.t1339 142.279
R12202 VDD.t1437 VDD.t555 142.279
R12203 VDD.t242 VDD.t464 142.279
R12204 VDD.t1430 VDD.t865 141.061
R12205 VDD.t606 VDD.t553 141.061
R12206 VDD.n669 VDD.t1476 139.107
R12207 VDD.n1019 VDD.t1398 139.107
R12208 VDD.t353 VDD.n263 139.107
R12209 VDD VDD.t1037 138.857
R12210 VDD VDD.t832 138.857
R12211 VDD.t865 VDD.t385 138.183
R12212 VDD.t574 VDD.t620 138.183
R12213 VDD.t553 VDD.t839 138.183
R12214 VDD.t152 VDD.t161 138.183
R12215 VDD.t1498 VDD 137.946
R12216 VDD.t528 VDD.n1821 136.591
R12217 VDD.t481 VDD.n2142 136.591
R12218 VDD.t118 VDD.n2400 136.591
R12219 VDD.t652 VDD.n2658 136.591
R12220 VDD.t12 VDD.n2916 136.591
R12221 VDD.t718 VDD.n3174 136.591
R12222 VDD.t411 VDD.n3432 136.591
R12223 VDD.t530 VDD.n5752 136.591
R12224 VDD.t482 VDD.n5498 136.591
R12225 VDD.t410 VDD.n3690 136.591
R12226 VDD.t116 VDD.n3948 136.591
R12227 VDD.t489 VDD.n4206 136.591
R12228 VDD.t84 VDD.n4464 136.591
R12229 VDD.t717 VDD.n4722 136.591
R12230 VDD.t1353 VDD.n4980 136.591
R12231 VDD.t529 VDD.n5238 136.591
R12232 VDD.n1697 VDD.n1696 135.117
R12233 VDD.n2046 VDD.n2045 135.117
R12234 VDD.n2276 VDD.n2275 135.117
R12235 VDD.n2534 VDD.n2533 135.117
R12236 VDD.n2792 VDD.n2791 135.117
R12237 VDD.n3050 VDD.n3049 135.117
R12238 VDD.n3308 VDD.n3307 135.117
R12239 VDD.n5631 VDD.n5630 135.117
R12240 VDD.n5377 VDD.n5376 135.117
R12241 VDD.n3566 VDD.n3565 135.117
R12242 VDD.n3824 VDD.n3823 135.117
R12243 VDD.n4082 VDD.n4081 135.117
R12244 VDD.n4340 VDD.n4339 135.117
R12245 VDD.n4598 VDD.n4597 135.117
R12246 VDD.n4856 VDD.n4855 135.117
R12247 VDD.n5114 VDD.n5113 135.117
R12248 VDD.t201 VDD.t1039 134.732
R12249 VDD.t383 VDD.t468 134.732
R12250 VDD.t465 VDD.t203 134.732
R12251 VDD.t400 VDD.t510 134.732
R12252 VDD.n1371 VDD.t1498 132.74
R12253 VDD VDD.t1143 132.321
R12254 VDD.t1127 VDD 132.321
R12255 VDD VDD.t1107 132.321
R12256 VDD.t1159 VDD.n668 132.321
R12257 VDD VDD.t1069 132.321
R12258 VDD VDD.t1452 132.321
R12259 VDD VDD.t1014 132.321
R12260 VDD.t1000 VDD 132.321
R12261 VDD VDD.t978 132.321
R12262 VDD.t902 VDD.n1018 132.321
R12263 VDD VDD.t940 132.321
R12264 VDD VDD.t1406 132.321
R12265 VDD VDD.t337 132.321
R12266 VDD.t321 VDD 132.321
R12267 VDD VDD.t301 132.321
R12268 VDD VDD.t263 132.321
R12269 VDD.n264 VDD.t451 132.321
R12270 VDD VDD.t427 132.321
R12271 VDD.t563 VDD.t201 131.983
R12272 VDD.t535 VDD.t383 131.983
R12273 VDD.t1034 VDD.t1394 131.983
R12274 VDD.t838 VDD.t465 131.983
R12275 VDD.t32 VDD.t400 131.983
R12276 VDD.t1199 VDD.t467 131.983
R12277 VDD.n1715 VDD.n1672 131.388
R12278 VDD.n2064 VDD.n2021 131.388
R12279 VDD.n2294 VDD.n2251 131.388
R12280 VDD.n2552 VDD.n2509 131.388
R12281 VDD.n2810 VDD.n2767 131.388
R12282 VDD.n3068 VDD.n3025 131.388
R12283 VDD.n3326 VDD.n3283 131.388
R12284 VDD.n5649 VDD.n5606 131.388
R12285 VDD.n5395 VDD.n5352 131.388
R12286 VDD.n3584 VDD.n3541 131.388
R12287 VDD.n3842 VDD.n3799 131.388
R12288 VDD.n4100 VDD.n4057 131.388
R12289 VDD.n4358 VDD.n4315 131.388
R12290 VDD.n4616 VDD.n4573 131.388
R12291 VDD.n4874 VDD.n4831 131.388
R12292 VDD.n5132 VDD.n5089 131.388
R12293 VDD.n1766 VDD.n1673 131.012
R12294 VDD.n2115 VDD.n2022 131.012
R12295 VDD.n2345 VDD.n2252 131.012
R12296 VDD.n2603 VDD.n2510 131.012
R12297 VDD.n2861 VDD.n2768 131.012
R12298 VDD.n3119 VDD.n3026 131.012
R12299 VDD.n3377 VDD.n3284 131.012
R12300 VDD.n5700 VDD.n5607 131.012
R12301 VDD.n5446 VDD.n5353 131.012
R12302 VDD.n3635 VDD.n3542 131.012
R12303 VDD.n3893 VDD.n3800 131.012
R12304 VDD.n4151 VDD.n4058 131.012
R12305 VDD.n4409 VDD.n4316 131.012
R12306 VDD.n4667 VDD.n4574 131.012
R12307 VDD.n4925 VDD.n4832 131.012
R12308 VDD.n5183 VDD.n5090 131.012
R12309 VDD.n1767 VDD.n1672 130.636
R12310 VDD.n1767 VDD.n1766 130.636
R12311 VDD.n2116 VDD.n2021 130.636
R12312 VDD.n2116 VDD.n2115 130.636
R12313 VDD.n2346 VDD.n2251 130.636
R12314 VDD.n2346 VDD.n2345 130.636
R12315 VDD.n2604 VDD.n2509 130.636
R12316 VDD.n2604 VDD.n2603 130.636
R12317 VDD.n2862 VDD.n2767 130.636
R12318 VDD.n2862 VDD.n2861 130.636
R12319 VDD.n3120 VDD.n3025 130.636
R12320 VDD.n3120 VDD.n3119 130.636
R12321 VDD.n3378 VDD.n3283 130.636
R12322 VDD.n3378 VDD.n3377 130.636
R12323 VDD.n5701 VDD.n5606 130.636
R12324 VDD.n5701 VDD.n5700 130.636
R12325 VDD.n5447 VDD.n5352 130.636
R12326 VDD.n5447 VDD.n5446 130.636
R12327 VDD.n3636 VDD.n3541 130.636
R12328 VDD.n3636 VDD.n3635 130.636
R12329 VDD.n3894 VDD.n3799 130.636
R12330 VDD.n3894 VDD.n3893 130.636
R12331 VDD.n4152 VDD.n4057 130.636
R12332 VDD.n4152 VDD.n4151 130.636
R12333 VDD.n4410 VDD.n4315 130.636
R12334 VDD.n4410 VDD.n4409 130.636
R12335 VDD.n4668 VDD.n4573 130.636
R12336 VDD.n4668 VDD.n4667 130.636
R12337 VDD.n4926 VDD.n4831 130.636
R12338 VDD.n4926 VDD.n4925 130.636
R12339 VDD.n5184 VDD.n5089 130.636
R12340 VDD.n5184 VDD.n5183 130.636
R12341 VDD.n1879 VDD.n1823 129.691
R12342 VDD.n2200 VDD.n2144 129.691
R12343 VDD.n2458 VDD.n2402 129.691
R12344 VDD.n2716 VDD.n2660 129.691
R12345 VDD.n2974 VDD.n2918 129.691
R12346 VDD.n3232 VDD.n3176 129.691
R12347 VDD.n3490 VDD.n3434 129.691
R12348 VDD.n5810 VDD.n5754 129.691
R12349 VDD.n5556 VDD.n5500 129.691
R12350 VDD.n3748 VDD.n3692 129.691
R12351 VDD.n4006 VDD.n3950 129.691
R12352 VDD.n4264 VDD.n4208 129.691
R12353 VDD.n4522 VDD.n4466 129.691
R12354 VDD.n4780 VDD.n4724 129.691
R12355 VDD.n5038 VDD.n4982 129.691
R12356 VDD.n5296 VDD.n5240 129.691
R12357 VDD VDD.t546 129.228
R12358 VDD VDD.t230 129.228
R12359 VDD VDD.t564 127.233
R12360 VDD VDD.t49 127.233
R12361 VDD VDD.t70 127.233
R12362 VDD.t26 VDD 126.02
R12363 VDD.t1182 VDD 126.02
R12364 VDD.t722 VDD 126.02
R12365 VDD.t601 VDD 126.02
R12366 VDD.t1024 VDD 126.02
R12367 VDD.t1482 VDD 126.02
R12368 VDD.t1447 VDD 126.02
R12369 VDD.t1195 VDD 126.02
R12370 VDD.t86 VDD 126.02
R12371 VDD.t457 VDD 126.02
R12372 VDD.t1441 VDD 126.02
R12373 VDD.t725 VDD 126.02
R12374 VDD.t882 VDD 126.02
R12375 VDD.t1347 VDD 126.02
R12376 VDD.t739 VDD 126.02
R12377 VDD.t236 VDD 126.02
R12378 VDD.t251 VDD.t826 122.144
R12379 VDD.t822 VDD.t603 122.144
R12380 VDD.t398 VDD.t1343 122.144
R12381 VDD.n1903 VDD.n1898 121.977
R12382 VDD.n2224 VDD.n2219 121.977
R12383 VDD.n2482 VDD.n2477 121.977
R12384 VDD.n2740 VDD.n2735 121.977
R12385 VDD.n2998 VDD.n2993 121.977
R12386 VDD.n3256 VDD.n3251 121.977
R12387 VDD.n3514 VDD.n3509 121.977
R12388 VDD.n5834 VDD.n5829 121.977
R12389 VDD.n5580 VDD.n5575 121.977
R12390 VDD.n3772 VDD.n3767 121.977
R12391 VDD.n4030 VDD.n4025 121.977
R12392 VDD.n4288 VDD.n4283 121.977
R12393 VDD.n4546 VDD.n4541 121.977
R12394 VDD.n4804 VDD.n4799 121.977
R12395 VDD.n5062 VDD.n5057 121.977
R12396 VDD.n5320 VDD.n5315 121.977
R12397 VDD.t150 VDD.t232 121.529
R12398 VDD.t504 VDD.t1177 121.529
R12399 VDD.n1764 VDD.t388 121.114
R12400 VDD.t388 VDD.n1711 121.114
R12401 VDD.n2113 VDD.t228 121.114
R12402 VDD.t228 VDD.n2060 121.114
R12403 VDD.n2343 VDD.t181 121.114
R12404 VDD.t181 VDD.n2290 121.114
R12405 VDD.n2601 VDD.t713 121.114
R12406 VDD.t713 VDD.n2548 121.114
R12407 VDD.n2859 VDD.t542 121.114
R12408 VDD.t542 VDD.n2806 121.114
R12409 VDD.n3117 VDD.t647 121.114
R12410 VDD.t647 VDD.n3064 121.114
R12411 VDD.n3375 VDD.t30 121.114
R12412 VDD.t30 VDD.n3322 121.114
R12413 VDD.n5698 VDD.t870 121.114
R12414 VDD.t870 VDD.n5645 121.114
R12415 VDD.n5444 VDD.t709 121.114
R12416 VDD.t709 VDD.n5391 121.114
R12417 VDD.n3633 VDD.t214 121.114
R12418 VDD.t214 VDD.n3580 121.114
R12419 VDD.n3891 VDD.t1027 121.114
R12420 VDD.t1027 VDD.n3838 121.114
R12421 VDD.n4149 VDD.t423 121.114
R12422 VDD.t423 VDD.n4096 121.114
R12423 VDD.n4407 VDD.t1031 121.114
R12424 VDD.t1031 VDD.n4354 121.114
R12425 VDD.n4665 VDD.t402 121.114
R12426 VDD.t402 VDD.n4612 121.114
R12427 VDD.n4923 VDD.t532 121.114
R12428 VDD.t532 VDD.n4870 121.114
R12429 VDD.n5181 VDD.t381 121.114
R12430 VDD.t381 VDD.n5128 121.114
R12431 VDD.t526 VDD.t801 120.909
R12432 VDD.t490 VDD.t548 120.909
R12433 VDD.t1484 VDD.t770 120.909
R12434 VDD.t850 VDD.t415 120.909
R12435 VDD.n1853 VDD.n1845 120.094
R12436 VDD.n2174 VDD.n2166 120.094
R12437 VDD.n2432 VDD.n2424 120.094
R12438 VDD.n2690 VDD.n2682 120.094
R12439 VDD.n2948 VDD.n2940 120.094
R12440 VDD.n3206 VDD.n3198 120.094
R12441 VDD.n3464 VDD.n3456 120.094
R12442 VDD.n5784 VDD.n5776 120.094
R12443 VDD.n5530 VDD.n5522 120.094
R12444 VDD.n3722 VDD.n3714 120.094
R12445 VDD.n3980 VDD.n3972 120.094
R12446 VDD.n4238 VDD.n4230 120.094
R12447 VDD.n4496 VDD.n4488 120.094
R12448 VDD.n4754 VDD.n4746 120.094
R12449 VDD.n5012 VDD.n5004 120.094
R12450 VDD.n5270 VDD.n5262 120.094
R12451 VDD.n1 VDD.t811 117.451
R12452 VDD.n468 VDD.t493 117.451
R12453 VDD.n439 VDD.t800 117.451
R12454 VDD.n459 VDD.t494 117.451
R12455 VDD.n66 VDD.t854 117.451
R12456 VDD.n36 VDD.t762 117.451
R12457 VDD.n56 VDD.t852 117.451
R12458 VDD.n1145 VDD.t782 117.451
R12459 VDD.n5 VDD.t233 116.322
R12460 VDD.n494 VDD.t527 116.322
R12461 VDD.n422 VDD.t38 116.322
R12462 VDD.n418 VDD.t547 116.322
R12463 VDD.n401 VDD.t1202 116.322
R12464 VDD.n92 VDD.t1485 116.322
R12465 VDD.n1149 VDD.t1178 116.322
R12466 VDD.n1580 VDD.t1432 116.322
R12467 VDD.n1576 VDD.t231 116.322
R12468 VDD.n1559 VDD.t36 116.322
R12469 VDD.n806 VDD.t807 116.322
R12470 VDD.n1189 VDD.t776 116.322
R12471 VDD.n1768 VDD.n1767 116.267
R12472 VDD.n2117 VDD.n2116 116.267
R12473 VDD.n2347 VDD.n2346 116.267
R12474 VDD.n2605 VDD.n2604 116.267
R12475 VDD.n2863 VDD.n2862 116.267
R12476 VDD.n3121 VDD.n3120 116.267
R12477 VDD.n3379 VDD.n3378 116.267
R12478 VDD.n5702 VDD.n5701 116.267
R12479 VDD.n5448 VDD.n5447 116.267
R12480 VDD.n3637 VDD.n3636 116.267
R12481 VDD.n3895 VDD.n3894 116.267
R12482 VDD.n4153 VDD.n4152 116.267
R12483 VDD.n4411 VDD.n4410 116.267
R12484 VDD.n4669 VDD.n4668 116.267
R12485 VDD.n4927 VDD.n4926 116.267
R12486 VDD.n5185 VDD.n5184 116.267
R12487 VDD.t1037 VDD.t806 115.486
R12488 VDD.t832 VDD.t775 115.486
R12489 VDD.n670 VDD 115.358
R12490 VDD.n1020 VDD 115.358
R12491 VDD.t329 VDD.n262 115.358
R12492 VDD.n1907 VDD.n1888 112.189
R12493 VDD.n1854 VDD.n1843 112.189
R12494 VDD.n2175 VDD.n2164 112.189
R12495 VDD.n2228 VDD.n2209 112.189
R12496 VDD.n2433 VDD.n2422 112.189
R12497 VDD.n2486 VDD.n2467 112.189
R12498 VDD.n2691 VDD.n2680 112.189
R12499 VDD.n2744 VDD.n2725 112.189
R12500 VDD.n2949 VDD.n2938 112.189
R12501 VDD.n3002 VDD.n2983 112.189
R12502 VDD.n3207 VDD.n3196 112.189
R12503 VDD.n3260 VDD.n3241 112.189
R12504 VDD.n3465 VDD.n3454 112.189
R12505 VDD.n3518 VDD.n3499 112.189
R12506 VDD.n5785 VDD.n5774 112.189
R12507 VDD.n5838 VDD.n5819 112.189
R12508 VDD.n5531 VDD.n5520 112.189
R12509 VDD.n5584 VDD.n5565 112.189
R12510 VDD.n3723 VDD.n3712 112.189
R12511 VDD.n3776 VDD.n3757 112.189
R12512 VDD.n3981 VDD.n3970 112.189
R12513 VDD.n4034 VDD.n4015 112.189
R12514 VDD.n4239 VDD.n4228 112.189
R12515 VDD.n4292 VDD.n4273 112.189
R12516 VDD.n4497 VDD.n4486 112.189
R12517 VDD.n4550 VDD.n4531 112.189
R12518 VDD.n4755 VDD.n4744 112.189
R12519 VDD.n4808 VDD.n4789 112.189
R12520 VDD.n5013 VDD.n5002 112.189
R12521 VDD.n5066 VDD.n5047 112.189
R12522 VDD.n5271 VDD.n5260 112.189
R12523 VDD.n5324 VDD.n5305 112.189
R12524 VDD.t795 VDD.t1029 110.834
R12525 VDD.t754 VDD.t206 110.834
R12526 VDD.t1209 VDD.t1319 109.316
R12527 VDD.t1281 VDD.t1209 109.316
R12528 VDD.t1309 VDD.t1281 109.316
R12529 VDD.t1231 VDD.t1309 109.316
R12530 VDD.t1267 VDD.t1231 109.316
R12531 VDD.t1313 VDD.t1267 109.316
R12532 VDD.t1235 VDD.t1313 109.316
R12533 VDD.t1271 VDD.t1235 109.316
R12534 VDD.t1259 VDD.t1271 109.316
R12535 VDD.t1293 VDD.t1259 109.316
R12536 VDD.t1317 VDD.t1293 109.316
R12537 VDD.t1265 VDD.t1317 109.316
R12538 VDD.t1297 VDD.t1265 109.316
R12539 VDD.t1223 VDD.t1297 109.316
R12540 VDD.t1249 VDD.t1223 109.316
R12541 VDD.t1305 VDD.t1227 109.316
R12542 VDD.t1227 VDD.t1261 109.316
R12543 VDD.t1261 VDD.t1213 109.316
R12544 VDD.t1213 VDD.t1303 109.316
R12545 VDD.t1303 VDD.t1327 109.316
R12546 VDD.t1327 VDD.t1255 109.316
R12547 VDD.t1255 VDD.t1287 109.316
R12548 VDD.t1239 VDD.t1315 109.316
R12549 VDD.t1291 VDD.t1239 109.316
R12550 VDD.t1217 VDD.t1291 109.316
R12551 VDD.t1243 VDD.t1217 109.316
R12552 VDD.t1275 VDD.t1243 109.316
R12553 VDD.t1211 VDD.t1275 109.316
R12554 VDD.t1301 VDD.t1211 109.316
R12555 VDD.t1207 VDD.t1279 109.316
R12556 VDD.t1221 VDD.t1247 109.316
R12557 VDD.t1247 VDD.t1299 109.316
R12558 VDD.t1277 VDD.t1307 109.316
R12559 VDD.t1307 VDD.t1229 109.316
R12560 VDD.t1229 VDD.t1325 109.316
R12561 VDD.t1285 VDD.t1253 109.316
R12562 VDD.t1329 VDD.t1285 109.316
R12563 VDD.t1257 VDD.t1329 109.316
R12564 VDD.t1289 VDD.t1215 109.316
R12565 VDD.t1215 VDD.t1241 109.316
R12566 VDD.t1241 VDD.t1273 109.316
R12567 VDD.t1273 VDD.t1219 109.316
R12568 VDD.t1219 VDD.t1245 109.316
R12569 VDD.t1245 VDD.t1323 109.316
R12570 VDD.t691 VDD.t697 109.316
R12571 VDD.t697 VDD.t675 109.316
R12572 VDD.t675 VDD.t685 109.316
R12573 VDD.t677 VDD.t695 109.316
R12574 VDD.t687 VDD.t677 109.316
R12575 VDD.t667 VDD.t687 109.316
R12576 VDD.t673 VDD.t683 109.316
R12577 VDD.t683 VDD.t679 109.316
R12578 VDD.t679 VDD.t693 109.316
R12579 VDD.t681 VDD.t671 109.316
R12580 VDD.t689 VDD.t681 109.316
R12581 VDD.t659 VDD.t655 109.316
R12582 VDD.t655 VDD.t657 109.316
R12583 VDD.t657 VDD.t661 109.316
R12584 VDD.t1135 VDD.n667 108.572
R12585 VDD.t1006 VDD.n1017 108.572
R12586 VDD.n265 VDD 108.572
R12587 VDD.t867 VDD.t205 106.709
R12588 VDD.t555 VDD.t242 106.709
R12589 VDD.t385 VDD.t574 103.636
R12590 VDD.t839 VDD.t152 103.636
R12591 VDD.n1769 VDD.n1768 102.721
R12592 VDD.n1755 VDD.n1671 102.721
R12593 VDD.n2118 VDD.n2117 102.721
R12594 VDD.n2104 VDD.n2020 102.721
R12595 VDD.n2348 VDD.n2347 102.721
R12596 VDD.n2334 VDD.n2250 102.721
R12597 VDD.n2606 VDD.n2605 102.721
R12598 VDD.n2592 VDD.n2508 102.721
R12599 VDD.n2864 VDD.n2863 102.721
R12600 VDD.n2850 VDD.n2766 102.721
R12601 VDD.n3122 VDD.n3121 102.721
R12602 VDD.n3108 VDD.n3024 102.721
R12603 VDD.n3380 VDD.n3379 102.721
R12604 VDD.n3366 VDD.n3282 102.721
R12605 VDD.n5703 VDD.n5702 102.721
R12606 VDD.n5689 VDD.n5605 102.721
R12607 VDD.n5449 VDD.n5448 102.721
R12608 VDD.n5435 VDD.n5351 102.721
R12609 VDD.n3638 VDD.n3637 102.721
R12610 VDD.n3624 VDD.n3540 102.721
R12611 VDD.n3896 VDD.n3895 102.721
R12612 VDD.n3882 VDD.n3798 102.721
R12613 VDD.n4154 VDD.n4153 102.721
R12614 VDD.n4140 VDD.n4056 102.721
R12615 VDD.n4412 VDD.n4411 102.721
R12616 VDD.n4398 VDD.n4314 102.721
R12617 VDD.n4670 VDD.n4669 102.721
R12618 VDD.n4656 VDD.n4572 102.721
R12619 VDD.n4928 VDD.n4927 102.721
R12620 VDD.n4914 VDD.n4830 102.721
R12621 VDD.n5186 VDD.n5185 102.721
R12622 VDD.n5172 VDD.n5088 102.721
R12623 VDD VDD.t1249 101.507
R12624 VDD.t1299 VDD 101.507
R12625 VDD.t1323 VDD 101.507
R12626 VDD.t669 VDD 101.507
R12627 VDD.t608 VDD 99.5973
R12628 VDD.t1175 VDD 99.5973
R12629 VDD.t818 VDD 99.5973
R12630 VDD.t1189 VDD 99.5973
R12631 VDD.t406 VDD 99.5973
R12632 VDD.t827 VDD 99.5973
R12633 VDD.t663 VDD 99.5973
R12634 VDD.t90 VDD 99.5973
R12635 VDD.t188 VDD 99.5973
R12636 VDD.t1345 VDD 99.5973
R12637 VDD.t240 VDD 99.5973
R12638 VDD.t2 VDD 99.5973
R12639 VDD.t1186 VDD 99.5973
R12640 VDD.t1369 VDD 99.5973
R12641 VDD.t540 VDD 99.5973
R12642 VDD.t1184 VDD 99.5973
R12643 VDD VDD.t37 99.5409
R12644 VDD VDD.t764 99.5409
R12645 VDD.t1200 VDD.t563 98.9875
R12646 VDD.t1394 VDD.t535 98.9875
R12647 VDD.t716 VDD.t838 98.9875
R12648 VDD.t467 VDD.t32 98.9875
R12649 VDD.n1429 VDD.t1257 98.9046
R12650 VDD.t508 VDD.t701 97.8793
R12651 VDD.t791 VDD.t143 97.8793
R12652 VDD.t661 VDD 97.6032
R12653 VDD.n31 VDD.t158 96.1553
R12654 VDD.n672 VDD.t252 96.1553
R12655 VDD.n508 VDD.t866 96.1553
R12656 VDD.n435 VDD.t1395 96.1553
R12657 VDD.n404 VDD.t420 96.1553
R12658 VDD.n106 VDD.t554 96.1553
R12659 VDD.n1175 VDD.t1438 96.1553
R12660 VDD.n1593 VDD.t749 96.1553
R12661 VDD.n1562 VDD.t1193 96.1553
R12662 VDD.n800 VDD.t384 96.1553
R12663 VDD.n803 VDD.t202 96.1553
R12664 VDD.n1022 VDD.t823 96.1553
R12665 VDD.n267 VDD.t399 96.1553
R12666 VDD.n1183 VDD.t401 96.1553
R12667 VDD.n1186 VDD.t466 96.1553
R12668 VDD.n585 VDD.t1111 95.0005
R12669 VDD.n935 VDD.t984 95.0005
R12670 VDD.t1339 VDD 94.8523
R12671 VDD.t464 VDD 94.8523
R12672 VDD.n482 VDD.t796 93.81
R12673 VDD.n80 VDD.t755 93.81
R12674 VDD.t548 VDD 93.5611
R12675 VDD.t415 VDD 93.5611
R12676 VDD.t737 VDD 93.539
R12677 VDD.t1396 VDD 93.539
R12678 VDD VDD.t1200 93.4882
R12679 VDD VDD.t716 93.4882
R12680 VDD.t216 VDD 93.3702
R12681 VDD.t880 VDD 93.3702
R12682 VDD.n1733 VDD.n1730 92.5005
R12683 VDD.n2082 VDD.n2079 92.5005
R12684 VDD.n2312 VDD.n2309 92.5005
R12685 VDD.n2570 VDD.n2567 92.5005
R12686 VDD.n2828 VDD.n2825 92.5005
R12687 VDD.n3086 VDD.n3083 92.5005
R12688 VDD.n3344 VDD.n3341 92.5005
R12689 VDD.n5667 VDD.n5664 92.5005
R12690 VDD.n5413 VDD.n5410 92.5005
R12691 VDD.n3602 VDD.n3599 92.5005
R12692 VDD.n3860 VDD.n3857 92.5005
R12693 VDD.n4118 VDD.n4115 92.5005
R12694 VDD.n4376 VDD.n4373 92.5005
R12695 VDD.n4634 VDD.n4631 92.5005
R12696 VDD.n4892 VDD.n4889 92.5005
R12697 VDD.n5150 VDD.n5147 92.5005
R12698 VDD.t620 VDD 92.1217
R12699 VDD.t161 VDD 92.1217
R12700 VDD.t699 VDD.t808 91.8882
R12701 VDD.t141 VDD.t778 91.8882
R12702 VDD.n1915 VDD.n1891 91.7652
R12703 VDD.n2236 VDD.n2212 91.7652
R12704 VDD.n2494 VDD.n2470 91.7652
R12705 VDD.n2752 VDD.n2728 91.7652
R12706 VDD.n3010 VDD.n2986 91.7652
R12707 VDD.n3268 VDD.n3244 91.7652
R12708 VDD.n3526 VDD.n3502 91.7652
R12709 VDD.n5846 VDD.n5822 91.7652
R12710 VDD.n5592 VDD.n5568 91.7652
R12711 VDD.n3784 VDD.n3760 91.7652
R12712 VDD.n4042 VDD.n4018 91.7652
R12713 VDD.n4300 VDD.n4276 91.7652
R12714 VDD.n4558 VDD.n4534 91.7652
R12715 VDD.n4816 VDD.n4792 91.7652
R12716 VDD.n5074 VDD.n5050 91.7652
R12717 VDD.n5332 VDD.n5308 91.7652
R12718 VDD.t299 VDD.n183 91.6076
R12719 VDD.n1960 VDD.n1959 91.4829
R12720 VDD.n1959 VDD.n1929 91.4829
R12721 VDD.n1972 VDD.n1929 91.4829
R12722 VDD.n1972 VDD.n1971 91.4829
R12723 VDD.n1950 VDD.n1937 91.4829
R12724 VDD.n1965 VDD.n1937 91.4829
R12725 VDD.n1966 VDD.n1965 91.4829
R12726 VDD.n1967 VDD.n1966 91.4829
R12727 VDD.n1884 VDD.n1820 91.343
R12728 VDD.n2205 VDD.n2141 91.343
R12729 VDD.n2463 VDD.n2399 91.343
R12730 VDD.n2721 VDD.n2657 91.343
R12731 VDD.n2979 VDD.n2915 91.343
R12732 VDD.n3237 VDD.n3173 91.343
R12733 VDD.n3495 VDD.n3431 91.343
R12734 VDD.n5815 VDD.n5751 91.343
R12735 VDD.n5561 VDD.n5497 91.343
R12736 VDD.n3753 VDD.n3689 91.343
R12737 VDD.n4011 VDD.n3947 91.343
R12738 VDD.n4269 VDD.n4205 91.343
R12739 VDD.n4527 VDD.n4463 91.343
R12740 VDD.n4785 VDD.n4721 91.343
R12741 VDD.n5043 VDD.n4979 91.343
R12742 VDD.n5301 VDD.n5237 91.343
R12743 VDD.n1372 VDD.t689 91.0964
R12744 VDD.n1827 VDD.t26 89.1694
R12745 VDD.n2148 VDD.t1182 89.1694
R12746 VDD.n2406 VDD.t722 89.1694
R12747 VDD.n2664 VDD.t601 89.1694
R12748 VDD.n2922 VDD.t1024 89.1694
R12749 VDD.n3180 VDD.t1482 89.1694
R12750 VDD.n3438 VDD.t1447 89.1694
R12751 VDD.n5758 VDD.t1195 89.1694
R12752 VDD.n5504 VDD.t86 89.1694
R12753 VDD.n3696 VDD.t457 89.1694
R12754 VDD.n3954 VDD.t1441 89.1694
R12755 VDD.n4212 VDD.t725 89.1694
R12756 VDD.n4470 VDD.t882 89.1694
R12757 VDD.n4728 VDD.t1347 89.1694
R12758 VDD.n4986 VDD.t739 89.1694
R12759 VDD.n5244 VDD.t236 89.1694
R12760 VDD.t810 VDD.t1381 88.9241
R12761 VDD.t781 VDD.t572 88.9241
R12762 VDD VDD.n1371 88.4936
R12763 VDD.n184 VDD.t305 88.2148
R12764 VDD VDD.t1034 87.9889
R12765 VDD VDD.t1199 87.9889
R12766 VDD.t711 VDD 87.8035
R12767 VDD.t747 VDD 87.8035
R12768 VDD.t506 VDD.t552 87.6928
R12769 VDD.t1342 VDD.t797 87.6928
R12770 VDD.t212 VDD.t414 87.6928
R12771 VDD.t25 VDD.t757 87.6928
R12772 VDD.n7 VDD.t151 86.7743
R12773 VDD.n7 VDD.t700 86.7743
R12774 VDD.n471 VDD.t702 86.7743
R12775 VDD.n471 VDD.t1030 86.7743
R12776 VDD.n441 VDD.t149 86.7743
R12777 VDD.n441 VDD.t703 86.7743
R12778 VDD.n443 VDD.t115 86.7743
R12779 VDD.n443 VDD.t534 86.7743
R12780 VDD.n69 VDD.t144 86.7743
R12781 VDD.n69 VDD.t207 86.7743
R12782 VDD.n38 VDD.t503 86.7743
R12783 VDD.n38 VDD.t146 86.7743
R12784 VDD.n40 VDD.t1397 86.7743
R12785 VDD.n40 VDD.t34 86.7743
R12786 VDD.n1151 VDD.t505 86.7743
R12787 VDD.n1151 VDD.t142 86.7743
R12788 VDD.t1105 VDD.n584 84.8219
R12789 VDD.t976 VDD.n934 84.8219
R12790 VDD.n438 VDD.n408 83.3098
R12791 VDD.n1596 VDD.n1566 83.3098
R12792 VDD.n1827 VDD.t208 81.2688
R12793 VDD.n2148 VDD.t836 81.2688
R12794 VDD.n2406 VDD.t1500 81.2688
R12795 VDD.n2664 VDD.t665 81.2688
R12796 VDD.n2922 VDD.t561 81.2688
R12797 VDD.n3180 VDD.t840 81.2688
R12798 VDD.n3438 VDD.t1355 81.2688
R12799 VDD.n5758 VDD.t417 81.2688
R12800 VDD.n5504 VDD.t813 81.2688
R12801 VDD.n3696 VDD.t390 81.2688
R12802 VDD.n3954 VDD.t868 81.2688
R12803 VDD.n4212 VDD.t604 81.2688
R12804 VDD.n4470 VDD.t1433 81.2688
R12805 VDD.n4728 VDD.t874 81.2688
R12806 VDD.n4986 VDD.t1435 81.2688
R12807 VDD.n5244 VDD.t153 81.2688
R12808 VDD.n1457 VDD.t1301 80.6854
R12809 VDD.n1760 VDD.n1717 80.5087
R12810 VDD.n2109 VDD.n2066 80.5087
R12811 VDD.n2339 VDD.n2296 80.5087
R12812 VDD.n2597 VDD.n2554 80.5087
R12813 VDD.n2855 VDD.n2812 80.5087
R12814 VDD.n3113 VDD.n3070 80.5087
R12815 VDD.n3371 VDD.n3328 80.5087
R12816 VDD.n5694 VDD.n5651 80.5087
R12817 VDD.n5440 VDD.n5397 80.5087
R12818 VDD.n3629 VDD.n3586 80.5087
R12819 VDD.n3887 VDD.n3844 80.5087
R12820 VDD.n4145 VDD.n4102 80.5087
R12821 VDD.n4403 VDD.n4360 80.5087
R12822 VDD.n4661 VDD.n4618 80.5087
R12823 VDD.n4919 VDD.n4876 80.5087
R12824 VDD.n5177 VDD.n5134 80.5087
R12825 VDD.n1708 VDD.n1669 80.2452
R12826 VDD.n2057 VDD.n2018 80.2452
R12827 VDD.n2287 VDD.n2248 80.2452
R12828 VDD.n2545 VDD.n2506 80.2452
R12829 VDD.n2803 VDD.n2764 80.2452
R12830 VDD.n3061 VDD.n3022 80.2452
R12831 VDD.n3319 VDD.n3280 80.2452
R12832 VDD.n5642 VDD.n5603 80.2452
R12833 VDD.n5388 VDD.n5349 80.2452
R12834 VDD.n3577 VDD.n3538 80.2452
R12835 VDD.n3835 VDD.n3796 80.2452
R12836 VDD.n4093 VDD.n4054 80.2452
R12837 VDD.n4351 VDD.n4312 80.2452
R12838 VDD.n4609 VDD.n4570 80.2452
R12839 VDD.n4867 VDD.n4828 80.2452
R12840 VDD.n5125 VDD.n5086 80.2452
R12841 VDD VDD.n1643 79.5475
R12842 VDD.t1279 VDD.t1321 78.5727
R12843 VDD VDD.n1634 78.5148
R12844 VDD.n1633 VDD.n1632 77.1383
R12845 VDD.n1870 VDD.n1845 76.5328
R12846 VDD.n2191 VDD.n2166 76.5328
R12847 VDD.n2449 VDD.n2424 76.5328
R12848 VDD.n2707 VDD.n2682 76.5328
R12849 VDD.n2965 VDD.n2940 76.5328
R12850 VDD.n3223 VDD.n3198 76.5328
R12851 VDD.n3481 VDD.n3456 76.5328
R12852 VDD.n5801 VDD.n5776 76.5328
R12853 VDD.n5547 VDD.n5522 76.5328
R12854 VDD.n3739 VDD.n3714 76.5328
R12855 VDD.n3997 VDD.n3972 76.5328
R12856 VDD.n4255 VDD.n4230 76.5328
R12857 VDD.n4513 VDD.n4488 76.5328
R12858 VDD.n4771 VDD.n4746 76.5328
R12859 VDD.n5029 VDD.n5004 76.5328
R12860 VDD.n5287 VDD.n5262 76.5328
R12861 VDD.n1625 VDD.n1624 76.0005
R12862 VDD.n1628 VDD.n1627 76.0005
R12863 VDD.n1630 VDD.n1629 76.0005
R12864 VDD.n1397 VDD.t667 75.48
R12865 VDD.n1869 VDD.n1844 74.1181
R12866 VDD.n2190 VDD.n2165 74.1181
R12867 VDD.n2448 VDD.n2423 74.1181
R12868 VDD.n2706 VDD.n2681 74.1181
R12869 VDD.n2964 VDD.n2939 74.1181
R12870 VDD.n3222 VDD.n3197 74.1181
R12871 VDD.n3480 VDD.n3455 74.1181
R12872 VDD.n5800 VDD.n5775 74.1181
R12873 VDD.n5546 VDD.n5521 74.1181
R12874 VDD.n3738 VDD.n3713 74.1181
R12875 VDD.n3996 VDD.n3971 74.1181
R12876 VDD.n4254 VDD.n4229 74.1181
R12877 VDD.n4512 VDD.n4487 74.1181
R12878 VDD.n4770 VDD.n4745 74.1181
R12879 VDD.n5028 VDD.n5003 74.1181
R12880 VDD.n5286 VDD.n5261 74.1181
R12881 VDD.n1871 VDD.n1843 71.6136
R12882 VDD.n2192 VDD.n2164 71.6136
R12883 VDD.n2450 VDD.n2422 71.6136
R12884 VDD.n2708 VDD.n2680 71.6136
R12885 VDD.n2966 VDD.n2938 71.6136
R12886 VDD.n3224 VDD.n3196 71.6136
R12887 VDD.n3482 VDD.n3454 71.6136
R12888 VDD.n5802 VDD.n5774 71.6136
R12889 VDD.n5548 VDD.n5520 71.6136
R12890 VDD.n3740 VDD.n3712 71.6136
R12891 VDD.n3998 VDD.n3970 71.6136
R12892 VDD.n4256 VDD.n4228 71.6136
R12893 VDD.n4514 VDD.n4486 71.6136
R12894 VDD.n4772 VDD.n4744 71.6136
R12895 VDD.n5030 VDD.n5002 71.6136
R12896 VDD.n5288 VDD.n5260 71.6136
R12897 VDD.n1809 VDD.t608 70.4844
R12898 VDD.n2130 VDD.t1175 70.4844
R12899 VDD.n2388 VDD.t818 70.4844
R12900 VDD.n2646 VDD.t1189 70.4844
R12901 VDD.n2904 VDD.t406 70.4844
R12902 VDD.n3162 VDD.t827 70.4844
R12903 VDD.n3420 VDD.t663 70.4844
R12904 VDD.n5740 VDD.t90 70.4844
R12905 VDD.n5486 VDD.t188 70.4844
R12906 VDD.n3678 VDD.t1345 70.4844
R12907 VDD.n3936 VDD.t240 70.4844
R12908 VDD.n4194 VDD.t2 70.4844
R12909 VDD.n4452 VDD.t1186 70.4844
R12910 VDD.n4710 VDD.t1369 70.4844
R12911 VDD.n4968 VDD.t540 70.4844
R12912 VDD.n5226 VDD.t1184 70.4844
R12913 VDD.t552 VDD.t1201 70.1543
R12914 VDD.t414 VDD.t35 70.1543
R12915 VDD.n1877 VDD.n1876 66.2808
R12916 VDD.n2198 VDD.n2197 66.2808
R12917 VDD.n2456 VDD.n2455 66.2808
R12918 VDD.n2714 VDD.n2713 66.2808
R12919 VDD.n2972 VDD.n2971 66.2808
R12920 VDD.n3230 VDD.n3229 66.2808
R12921 VDD.n3488 VDD.n3487 66.2808
R12922 VDD.n5808 VDD.n5807 66.2808
R12923 VDD.n5554 VDD.n5553 66.2808
R12924 VDD.n3746 VDD.n3745 66.2808
R12925 VDD.n4004 VDD.n4003 66.2808
R12926 VDD.n4262 VDD.n4261 66.2808
R12927 VDD.n4520 VDD.n4519 66.2808
R12928 VDD.n4778 VDD.n4777 66.2808
R12929 VDD.n5036 VDD.n5035 66.2808
R12930 VDD.n5294 VDD.n5293 66.2808
R12931 VDD.n1898 VDD.n1889 65.0929
R12932 VDD.n2219 VDD.n2210 65.0929
R12933 VDD.n2477 VDD.n2468 65.0929
R12934 VDD.n2735 VDD.n2726 65.0929
R12935 VDD.n2993 VDD.n2984 65.0929
R12936 VDD.n3251 VDD.n3242 65.0929
R12937 VDD.n3509 VDD.n3500 65.0929
R12938 VDD.n5829 VDD.n5820 65.0929
R12939 VDD.n5575 VDD.n5566 65.0929
R12940 VDD.n3767 VDD.n3758 65.0929
R12941 VDD.n4025 VDD.n4016 65.0929
R12942 VDD.n4283 VDD.n4274 65.0929
R12943 VDD.n4541 VDD.n4532 65.0929
R12944 VDD.n4799 VDD.n4790 65.0929
R12945 VDD.n5057 VDD.n5048 65.0929
R12946 VDD.n5315 VDD.n5306 65.0929
R12947 VDD.n1809 VDD.t1357 64.3553
R12948 VDD.n2130 VDD.t815 64.3553
R12949 VDD.n2388 VDD.t1379 64.3553
R12950 VDD.n2646 VDD.t872 64.3553
R12951 VDD.n2904 VDD.t394 64.3553
R12952 VDD.n3162 VDD.t544 64.3553
R12953 VDD.n3420 VDD.t618 64.3553
R12954 VDD.n5740 VDD.t575 64.3553
R12955 VDD.n5486 VDD.t1486 64.3553
R12956 VDD.n3678 VDD.t515 64.3553
R12957 VDD.n3936 VDD.t460 64.3553
R12958 VDD.n4194 VDD.t894 64.3553
R12959 VDD.n4452 VDD.t793 64.3553
R12960 VDD.n4710 VDD.t23 64.3553
R12961 VDD.n4968 VDD.t707 64.3553
R12962 VDD.n5226 VDD.t199 64.3553
R12963 VDD.n475 VDD.t491 63.3219
R12964 VDD.n475 VDD.t549 63.3219
R12965 VDD.n73 VDD.t851 63.3219
R12966 VDD.n73 VDD.t416 63.3219
R12967 VDD.n1706 VDD.n1673 63.2691
R12968 VDD.n1707 VDD.n1706 63.2691
R12969 VDD.n2055 VDD.n2022 63.2691
R12970 VDD.n2056 VDD.n2055 63.2691
R12971 VDD.n2285 VDD.n2252 63.2691
R12972 VDD.n2286 VDD.n2285 63.2691
R12973 VDD.n2543 VDD.n2510 63.2691
R12974 VDD.n2544 VDD.n2543 63.2691
R12975 VDD.n2801 VDD.n2768 63.2691
R12976 VDD.n2802 VDD.n2801 63.2691
R12977 VDD.n3059 VDD.n3026 63.2691
R12978 VDD.n3060 VDD.n3059 63.2691
R12979 VDD.n3317 VDD.n3284 63.2691
R12980 VDD.n3318 VDD.n3317 63.2691
R12981 VDD.n5640 VDD.n5607 63.2691
R12982 VDD.n5641 VDD.n5640 63.2691
R12983 VDD.n5386 VDD.n5353 63.2691
R12984 VDD.n5387 VDD.n5386 63.2691
R12985 VDD.n3575 VDD.n3542 63.2691
R12986 VDD.n3576 VDD.n3575 63.2691
R12987 VDD.n3833 VDD.n3800 63.2691
R12988 VDD.n3834 VDD.n3833 63.2691
R12989 VDD.n4091 VDD.n4058 63.2691
R12990 VDD.n4092 VDD.n4091 63.2691
R12991 VDD.n4349 VDD.n4316 63.2691
R12992 VDD.n4350 VDD.n4349 63.2691
R12993 VDD.n4607 VDD.n4574 63.2691
R12994 VDD.n4608 VDD.n4607 63.2691
R12995 VDD.n4865 VDD.n4832 63.2691
R12996 VDD.n4866 VDD.n4865 63.2691
R12997 VDD.n5123 VDD.n5090 63.2691
R12998 VDD.n5124 VDD.n5123 63.2691
R12999 VDD.n1762 VDD.n1715 61.5116
R13000 VDD.n1762 VDD.n1761 61.5116
R13001 VDD.n2111 VDD.n2064 61.5116
R13002 VDD.n2111 VDD.n2110 61.5116
R13003 VDD.n2341 VDD.n2294 61.5116
R13004 VDD.n2341 VDD.n2340 61.5116
R13005 VDD.n2599 VDD.n2552 61.5116
R13006 VDD.n2599 VDD.n2598 61.5116
R13007 VDD.n2857 VDD.n2810 61.5116
R13008 VDD.n2857 VDD.n2856 61.5116
R13009 VDD.n3115 VDD.n3068 61.5116
R13010 VDD.n3115 VDD.n3114 61.5116
R13011 VDD.n3373 VDD.n3326 61.5116
R13012 VDD.n3373 VDD.n3372 61.5116
R13013 VDD.n5696 VDD.n5649 61.5116
R13014 VDD.n5696 VDD.n5695 61.5116
R13015 VDD.n5442 VDD.n5395 61.5116
R13016 VDD.n5442 VDD.n5441 61.5116
R13017 VDD.n3631 VDD.n3584 61.5116
R13018 VDD.n3631 VDD.n3630 61.5116
R13019 VDD.n3889 VDD.n3842 61.5116
R13020 VDD.n3889 VDD.n3888 61.5116
R13021 VDD.n4147 VDD.n4100 61.5116
R13022 VDD.n4147 VDD.n4146 61.5116
R13023 VDD.n4405 VDD.n4358 61.5116
R13024 VDD.n4405 VDD.n4404 61.5116
R13025 VDD.n4663 VDD.n4616 61.5116
R13026 VDD.n4663 VDD.n4662 61.5116
R13027 VDD.n4921 VDD.n4874 61.5116
R13028 VDD.n4921 VDD.n4920 61.5116
R13029 VDD.n5179 VDD.n5132 61.5116
R13030 VDD.n5179 VDD.n5178 61.5116
R13031 VDD.n1908 VDD.n1897 60.6123
R13032 VDD.n1911 VDD.n1910 60.6123
R13033 VDD.n1910 VDD.n1903 60.6123
R13034 VDD.n1908 VDD.n1907 60.6123
R13035 VDD.n1860 VDD.n1852 60.6123
R13036 VDD.n1866 VDD.n1853 60.6123
R13037 VDD.n1866 VDD.n1865 60.6123
R13038 VDD.n1854 VDD.n1852 60.6123
R13039 VDD.n2181 VDD.n2173 60.6123
R13040 VDD.n2187 VDD.n2174 60.6123
R13041 VDD.n2187 VDD.n2186 60.6123
R13042 VDD.n2175 VDD.n2173 60.6123
R13043 VDD.n2229 VDD.n2218 60.6123
R13044 VDD.n2232 VDD.n2231 60.6123
R13045 VDD.n2231 VDD.n2224 60.6123
R13046 VDD.n2229 VDD.n2228 60.6123
R13047 VDD.n2439 VDD.n2431 60.6123
R13048 VDD.n2445 VDD.n2432 60.6123
R13049 VDD.n2445 VDD.n2444 60.6123
R13050 VDD.n2433 VDD.n2431 60.6123
R13051 VDD.n2487 VDD.n2476 60.6123
R13052 VDD.n2490 VDD.n2489 60.6123
R13053 VDD.n2489 VDD.n2482 60.6123
R13054 VDD.n2487 VDD.n2486 60.6123
R13055 VDD.n2697 VDD.n2689 60.6123
R13056 VDD.n2703 VDD.n2690 60.6123
R13057 VDD.n2703 VDD.n2702 60.6123
R13058 VDD.n2691 VDD.n2689 60.6123
R13059 VDD.n2745 VDD.n2734 60.6123
R13060 VDD.n2748 VDD.n2747 60.6123
R13061 VDD.n2747 VDD.n2740 60.6123
R13062 VDD.n2745 VDD.n2744 60.6123
R13063 VDD.n2955 VDD.n2947 60.6123
R13064 VDD.n2961 VDD.n2948 60.6123
R13065 VDD.n2961 VDD.n2960 60.6123
R13066 VDD.n2949 VDD.n2947 60.6123
R13067 VDD.n3003 VDD.n2992 60.6123
R13068 VDD.n3006 VDD.n3005 60.6123
R13069 VDD.n3005 VDD.n2998 60.6123
R13070 VDD.n3003 VDD.n3002 60.6123
R13071 VDD.n3213 VDD.n3205 60.6123
R13072 VDD.n3219 VDD.n3206 60.6123
R13073 VDD.n3219 VDD.n3218 60.6123
R13074 VDD.n3207 VDD.n3205 60.6123
R13075 VDD.n3261 VDD.n3250 60.6123
R13076 VDD.n3264 VDD.n3263 60.6123
R13077 VDD.n3263 VDD.n3256 60.6123
R13078 VDD.n3261 VDD.n3260 60.6123
R13079 VDD.n3471 VDD.n3463 60.6123
R13080 VDD.n3477 VDD.n3464 60.6123
R13081 VDD.n3477 VDD.n3476 60.6123
R13082 VDD.n3465 VDD.n3463 60.6123
R13083 VDD.n3519 VDD.n3508 60.6123
R13084 VDD.n3522 VDD.n3521 60.6123
R13085 VDD.n3521 VDD.n3514 60.6123
R13086 VDD.n3519 VDD.n3518 60.6123
R13087 VDD.n5791 VDD.n5783 60.6123
R13088 VDD.n5797 VDD.n5784 60.6123
R13089 VDD.n5797 VDD.n5796 60.6123
R13090 VDD.n5785 VDD.n5783 60.6123
R13091 VDD.n5839 VDD.n5828 60.6123
R13092 VDD.n5842 VDD.n5841 60.6123
R13093 VDD.n5841 VDD.n5834 60.6123
R13094 VDD.n5839 VDD.n5838 60.6123
R13095 VDD.n5537 VDD.n5529 60.6123
R13096 VDD.n5543 VDD.n5530 60.6123
R13097 VDD.n5543 VDD.n5542 60.6123
R13098 VDD.n5531 VDD.n5529 60.6123
R13099 VDD.n5585 VDD.n5574 60.6123
R13100 VDD.n5588 VDD.n5587 60.6123
R13101 VDD.n5587 VDD.n5580 60.6123
R13102 VDD.n5585 VDD.n5584 60.6123
R13103 VDD.n3729 VDD.n3721 60.6123
R13104 VDD.n3735 VDD.n3722 60.6123
R13105 VDD.n3735 VDD.n3734 60.6123
R13106 VDD.n3723 VDD.n3721 60.6123
R13107 VDD.n3777 VDD.n3766 60.6123
R13108 VDD.n3780 VDD.n3779 60.6123
R13109 VDD.n3779 VDD.n3772 60.6123
R13110 VDD.n3777 VDD.n3776 60.6123
R13111 VDD.n3987 VDD.n3979 60.6123
R13112 VDD.n3993 VDD.n3980 60.6123
R13113 VDD.n3993 VDD.n3992 60.6123
R13114 VDD.n3981 VDD.n3979 60.6123
R13115 VDD.n4035 VDD.n4024 60.6123
R13116 VDD.n4038 VDD.n4037 60.6123
R13117 VDD.n4037 VDD.n4030 60.6123
R13118 VDD.n4035 VDD.n4034 60.6123
R13119 VDD.n4245 VDD.n4237 60.6123
R13120 VDD.n4251 VDD.n4238 60.6123
R13121 VDD.n4251 VDD.n4250 60.6123
R13122 VDD.n4239 VDD.n4237 60.6123
R13123 VDD.n4293 VDD.n4282 60.6123
R13124 VDD.n4296 VDD.n4295 60.6123
R13125 VDD.n4295 VDD.n4288 60.6123
R13126 VDD.n4293 VDD.n4292 60.6123
R13127 VDD.n4503 VDD.n4495 60.6123
R13128 VDD.n4509 VDD.n4496 60.6123
R13129 VDD.n4509 VDD.n4508 60.6123
R13130 VDD.n4497 VDD.n4495 60.6123
R13131 VDD.n4551 VDD.n4540 60.6123
R13132 VDD.n4554 VDD.n4553 60.6123
R13133 VDD.n4553 VDD.n4546 60.6123
R13134 VDD.n4551 VDD.n4550 60.6123
R13135 VDD.n4761 VDD.n4753 60.6123
R13136 VDD.n4767 VDD.n4754 60.6123
R13137 VDD.n4767 VDD.n4766 60.6123
R13138 VDD.n4755 VDD.n4753 60.6123
R13139 VDD.n4809 VDD.n4798 60.6123
R13140 VDD.n4812 VDD.n4811 60.6123
R13141 VDD.n4811 VDD.n4804 60.6123
R13142 VDD.n4809 VDD.n4808 60.6123
R13143 VDD.n5019 VDD.n5011 60.6123
R13144 VDD.n5025 VDD.n5012 60.6123
R13145 VDD.n5025 VDD.n5024 60.6123
R13146 VDD.n5013 VDD.n5011 60.6123
R13147 VDD.n5067 VDD.n5056 60.6123
R13148 VDD.n5070 VDD.n5069 60.6123
R13149 VDD.n5069 VDD.n5062 60.6123
R13150 VDD.n5067 VDD.n5066 60.6123
R13151 VDD.n5277 VDD.n5269 60.6123
R13152 VDD.n5283 VDD.n5270 60.6123
R13153 VDD.n5283 VDD.n5282 60.6123
R13154 VDD.n5271 VDD.n5269 60.6123
R13155 VDD.n5325 VDD.n5314 60.6123
R13156 VDD.n5328 VDD.n5327 60.6123
R13157 VDD.n5327 VDD.n5320 60.6123
R13158 VDD.n5325 VDD.n5324 60.6123
R13159 VDD.n1456 VDD.t1277 59.8635
R13160 VDD.n1916 VDD.n1888 58.0325
R13161 VDD.n2237 VDD.n2209 58.0325
R13162 VDD.n2495 VDD.n2467 58.0325
R13163 VDD.n2753 VDD.n2725 58.0325
R13164 VDD.n3011 VDD.n2983 58.0325
R13165 VDD.n3269 VDD.n3241 58.0325
R13166 VDD.n3527 VDD.n3499 58.0325
R13167 VDD.n5847 VDD.n5819 58.0325
R13168 VDD.n5593 VDD.n5565 58.0325
R13169 VDD.n3785 VDD.n3757 58.0325
R13170 VDD.n4043 VDD.n4015 58.0325
R13171 VDD.n4301 VDD.n4273 58.0325
R13172 VDD.n4559 VDD.n4531 58.0325
R13173 VDD.n4817 VDD.n4789 58.0325
R13174 VDD.n5075 VDD.n5047 58.0325
R13175 VDD.n5333 VDD.n5305 58.0325
R13176 VDD.n584 VDD.t1079 57.6791
R13177 VDD.n934 VDD.t948 57.6791
R13178 VDD.t801 VDD.t711 57.5763
R13179 VDD.t770 VDD.t747 57.5763
R13180 VDD VDD.t148 57.5434
R13181 VDD VDD.t145 57.5434
R13182 VDD.t808 VDD.t216 56.3188
R13183 VDD.t778 VDD.t880 56.3188
R13184 VDD.n1732 VDD.n1731 55.4672
R13185 VDD.n1733 VDD.n1729 55.4672
R13186 VDD.n2081 VDD.n2080 55.4672
R13187 VDD.n2082 VDD.n2078 55.4672
R13188 VDD.n2311 VDD.n2310 55.4672
R13189 VDD.n2312 VDD.n2308 55.4672
R13190 VDD.n2569 VDD.n2568 55.4672
R13191 VDD.n2570 VDD.n2566 55.4672
R13192 VDD.n2827 VDD.n2826 55.4672
R13193 VDD.n2828 VDD.n2824 55.4672
R13194 VDD.n3085 VDD.n3084 55.4672
R13195 VDD.n3086 VDD.n3082 55.4672
R13196 VDD.n3343 VDD.n3342 55.4672
R13197 VDD.n3344 VDD.n3340 55.4672
R13198 VDD.n5666 VDD.n5665 55.4672
R13199 VDD.n5667 VDD.n5663 55.4672
R13200 VDD.n5412 VDD.n5411 55.4672
R13201 VDD.n5413 VDD.n5409 55.4672
R13202 VDD.n3601 VDD.n3600 55.4672
R13203 VDD.n3602 VDD.n3598 55.4672
R13204 VDD.n3859 VDD.n3858 55.4672
R13205 VDD.n3860 VDD.n3856 55.4672
R13206 VDD.n4117 VDD.n4116 55.4672
R13207 VDD.n4118 VDD.n4114 55.4672
R13208 VDD.n4375 VDD.n4374 55.4672
R13209 VDD.n4376 VDD.n4372 55.4672
R13210 VDD.n4633 VDD.n4632 55.4672
R13211 VDD.n4634 VDD.n4630 55.4672
R13212 VDD.n4891 VDD.n4890 55.4672
R13213 VDD.n4892 VDD.n4888 55.4672
R13214 VDD.n5149 VDD.n5148 55.4672
R13215 VDD.n5150 VDD.n5146 55.4672
R13216 VDD.n1803 VDD 54.4858
R13217 VDD.n2011 VDD 54.4858
R13218 VDD.n2382 VDD 54.4858
R13219 VDD.n2640 VDD 54.4858
R13220 VDD.n2898 VDD 54.4858
R13221 VDD.n3156 VDD 54.4858
R13222 VDD.n3414 VDD 54.4858
R13223 VDD.n5737 VDD 54.4858
R13224 VDD.n5483 VDD 54.4858
R13225 VDD.n3672 VDD 54.4858
R13226 VDD.n3930 VDD 54.4858
R13227 VDD.n4188 VDD 54.4858
R13228 VDD.n4446 VDD 54.4858
R13229 VDD.n4704 VDD 54.4858
R13230 VDD.n4962 VDD 54.4858
R13231 VDD.n5220 VDD 54.4858
R13232 VDD.t863 VDD.n1927 54.472
R13233 VDD.t1043 VDD.n1927 54.472
R13234 VDD.n184 VDD.t339 54.2862
R13235 VDD.n1953 VDD.t1041 54.2478
R13236 VDD.n1949 VDD.n1941 54.1098
R13237 VDD.n1969 VDD.n1931 54.1091
R13238 VDD.t419 VDD.t506 52.6159
R13239 VDD.t797 VDD.t737 52.6159
R13240 VDD.t1192 VDD.t212 52.6159
R13241 VDD.t757 VDD.t1396 52.6159
R13242 VDD.n183 VDD.t271 50.8934
R13243 VDD.t863 VDD.n1939 50.8854
R13244 VDD.t386 VDD.t63 50.6439
R13245 VDD.t100 VDD.t556 50.6439
R13246 VDD.n1876 VDD.n1818 50.1034
R13247 VDD.n2197 VDD.n2139 50.1034
R13248 VDD.n2455 VDD.n2397 50.1034
R13249 VDD.n2713 VDD.n2655 50.1034
R13250 VDD.n2971 VDD.n2913 50.1034
R13251 VDD.n3229 VDD.n3171 50.1034
R13252 VDD.n3487 VDD.n3429 50.1034
R13253 VDD.n5807 VDD.n5749 50.1034
R13254 VDD.n5553 VDD.n5495 50.1034
R13255 VDD.n3745 VDD.n3687 50.1034
R13256 VDD.n4003 VDD.n3945 50.1034
R13257 VDD.n4261 VDD.n4203 50.1034
R13258 VDD.n4519 VDD.n4461 50.1034
R13259 VDD.n4777 VDD.n4719 50.1034
R13260 VDD.n5035 VDD.n4977 50.1034
R13261 VDD.n5293 VDD.n5235 50.1034
R13262 VDD.t1225 VDD.n1456 49.4526
R13263 VDD.t1321 VDD.t1251 49.2598
R13264 VDD.t1251 VDD.t1283 49.2598
R13265 VDD.t1283 VDD.t1311 49.2598
R13266 VDD.t1311 VDD.t1233 49.2598
R13267 VDD.t1233 VDD.t1269 49.2598
R13268 VDD.t1269 VDD.t1205 49.2598
R13269 VDD.t1205 VDD.t1237 49.2598
R13270 VDD.t1237 VDD.t1203 49.2598
R13271 VDD.t1203 VDD.t1263 49.2598
R13272 VDD.t1263 VDD.t1295 49.2598
R13273 VDD.t1361 VDD.n1801 49.1183
R13274 VDD.t1490 VDD.n2009 49.1183
R13275 VDD.t220 VDD.n2380 49.1183
R13276 VDD.t57 VDD.n2638 49.1183
R13277 VDD.t593 VDD.n2896 49.1183
R13278 VDD.t39 VDD.n3154 49.1183
R13279 VDD.t729 VDD.n3412 49.1183
R13280 VDD.t162 VDD.n5735 49.1183
R13281 VDD.t519 VDD.n5481 49.1183
R13282 VDD.t191 VDD.n3670 49.1183
R13283 VDD.t171 VDD.n3928 49.1183
R13284 VDD.t94 VDD.n4186 49.1183
R13285 VDD.t495 VDD.n4444 49.1183
R13286 VDD.t585 VDD.n4702 49.1183
R13287 VDD.t577 VDD.n4960 49.1183
R13288 VDD.t855 VDD.n5218 49.1183
R13289 VDD.t1295 VDD.t1221 47.9846
R13290 VDD.n585 VDD.t1145 47.5005
R13291 VDD.n935 VDD.t1016 47.5005
R13292 VDD.n1700 VDD.n1681 47.0405
R13293 VDD.n2049 VDD.n2030 47.0405
R13294 VDD.n2279 VDD.n2260 47.0405
R13295 VDD.n2537 VDD.n2518 47.0405
R13296 VDD.n2795 VDD.n2776 47.0405
R13297 VDD.n3053 VDD.n3034 47.0405
R13298 VDD.n3311 VDD.n3292 47.0405
R13299 VDD.n5634 VDD.n5615 47.0405
R13300 VDD.n5380 VDD.n5361 47.0405
R13301 VDD.n3569 VDD.n3550 47.0405
R13302 VDD.n3827 VDD.n3808 47.0405
R13303 VDD.n4085 VDD.n4066 47.0405
R13304 VDD.n4343 VDD.n4324 47.0405
R13305 VDD.n4601 VDD.n4582 47.0405
R13306 VDD.n4859 VDD.n4840 47.0405
R13307 VDD.n5117 VDD.n5098 47.0405
R13308 VDD.n1966 VDD.n1936 46.6829
R13309 VDD.n1973 VDD.n1972 45.9299
R13310 VDD.n1959 VDD.n1958 45.9299
R13311 VDD.n1705 VDD.n1704 45.7605
R13312 VDD.n1689 VDD.n1685 45.7605
R13313 VDD.n2054 VDD.n2053 45.7605
R13314 VDD.n2038 VDD.n2034 45.7605
R13315 VDD.n2284 VDD.n2283 45.7605
R13316 VDD.n2268 VDD.n2264 45.7605
R13317 VDD.n2542 VDD.n2541 45.7605
R13318 VDD.n2526 VDD.n2522 45.7605
R13319 VDD.n2800 VDD.n2799 45.7605
R13320 VDD.n2784 VDD.n2780 45.7605
R13321 VDD.n3058 VDD.n3057 45.7605
R13322 VDD.n3042 VDD.n3038 45.7605
R13323 VDD.n3316 VDD.n3315 45.7605
R13324 VDD.n3300 VDD.n3296 45.7605
R13325 VDD.n5639 VDD.n5638 45.7605
R13326 VDD.n5623 VDD.n5619 45.7605
R13327 VDD.n5385 VDD.n5384 45.7605
R13328 VDD.n5369 VDD.n5365 45.7605
R13329 VDD.n3574 VDD.n3573 45.7605
R13330 VDD.n3558 VDD.n3554 45.7605
R13331 VDD.n3832 VDD.n3831 45.7605
R13332 VDD.n3816 VDD.n3812 45.7605
R13333 VDD.n4090 VDD.n4089 45.7605
R13334 VDD.n4074 VDD.n4070 45.7605
R13335 VDD.n4348 VDD.n4347 45.7605
R13336 VDD.n4332 VDD.n4328 45.7605
R13337 VDD.n4606 VDD.n4605 45.7605
R13338 VDD.n4590 VDD.n4586 45.7605
R13339 VDD.n4864 VDD.n4863 45.7605
R13340 VDD.n4848 VDD.n4844 45.7605
R13341 VDD.n5122 VDD.n5121 45.7605
R13342 VDD.n5106 VDD.n5102 45.7605
R13343 VDD.n1684 VDD.n1682 45.4405
R13344 VDD.n2033 VDD.n2031 45.4405
R13345 VDD.n2263 VDD.n2261 45.4405
R13346 VDD.n2521 VDD.n2519 45.4405
R13347 VDD.n2779 VDD.n2777 45.4405
R13348 VDD.n3037 VDD.n3035 45.4405
R13349 VDD.n3295 VDD.n3293 45.4405
R13350 VDD.n5618 VDD.n5616 45.4405
R13351 VDD.n5364 VDD.n5362 45.4405
R13352 VDD.n3553 VDD.n3551 45.4405
R13353 VDD.n3811 VDD.n3809 45.4405
R13354 VDD.n4069 VDD.n4067 45.4405
R13355 VDD.n4327 VDD.n4325 45.4405
R13356 VDD.n4585 VDD.n4583 45.4405
R13357 VDD.n4843 VDD.n4841 45.4405
R13358 VDD.n5101 VDD.n5099 45.4405
R13359 VDD.n1947 VDD.n1937 44.8005
R13360 VDD.n408 VDD 43.6586
R13361 VDD.n1566 VDD 43.6586
R13362 VDD.n1 VDD.t140 42.3555
R13363 VDD.n468 VDD.t712 42.3555
R13364 VDD.n439 VDD.t463 42.3555
R13365 VDD.n459 VDD.t405 42.3555
R13366 VDD.n66 VDD.t748 42.3555
R13367 VDD.n36 VDD.t156 42.3555
R13368 VDD.n56 VDD.t160 42.3555
R13369 VDD.n1145 VDD.t393 42.3555
R13370 VDD.n1947 VDD.n1946 41.323
R13371 VDD.n1936 VDD.n1933 41.2617
R13372 VDD.n1708 VDD.n1707 39.5299
R13373 VDD.n1761 VDD.n1760 39.5299
R13374 VDD.n2057 VDD.n2056 39.5299
R13375 VDD.n2110 VDD.n2109 39.5299
R13376 VDD.n2287 VDD.n2286 39.5299
R13377 VDD.n2340 VDD.n2339 39.5299
R13378 VDD.n2545 VDD.n2544 39.5299
R13379 VDD.n2598 VDD.n2597 39.5299
R13380 VDD.n2803 VDD.n2802 39.5299
R13381 VDD.n2856 VDD.n2855 39.5299
R13382 VDD.n3061 VDD.n3060 39.5299
R13383 VDD.n3114 VDD.n3113 39.5299
R13384 VDD.n3319 VDD.n3318 39.5299
R13385 VDD.n3372 VDD.n3371 39.5299
R13386 VDD.n5642 VDD.n5641 39.5299
R13387 VDD.n5695 VDD.n5694 39.5299
R13388 VDD.n5388 VDD.n5387 39.5299
R13389 VDD.n5441 VDD.n5440 39.5299
R13390 VDD.n3577 VDD.n3576 39.5299
R13391 VDD.n3630 VDD.n3629 39.5299
R13392 VDD.n3835 VDD.n3834 39.5299
R13393 VDD.n3888 VDD.n3887 39.5299
R13394 VDD.n4093 VDD.n4092 39.5299
R13395 VDD.n4146 VDD.n4145 39.5299
R13396 VDD.n4351 VDD.n4350 39.5299
R13397 VDD.n4404 VDD.n4403 39.5299
R13398 VDD.n4609 VDD.n4608 39.5299
R13399 VDD.n4662 VDD.n4661 39.5299
R13400 VDD.n4867 VDD.n4866 39.5299
R13401 VDD.n4920 VDD.n4919 39.5299
R13402 VDD.n5125 VDD.n5124 39.5299
R13403 VDD.n5178 VDD.n5177 39.5299
R13404 VDD.n20 VDD.n3 39.2858
R13405 VDD.n1164 VDD.n1147 39.2858
R13406 VDD VDD.t114 39.0862
R13407 VDD VDD.t33 39.0862
R13408 VDD.n1885 VDD.n1884 38.9491
R13409 VDD.n2206 VDD.n2205 38.9491
R13410 VDD.n2464 VDD.n2463 38.9491
R13411 VDD.n2722 VDD.n2721 38.9491
R13412 VDD.n2980 VDD.n2979 38.9491
R13413 VDD.n3238 VDD.n3237 38.9491
R13414 VDD.n3496 VDD.n3495 38.9491
R13415 VDD.n5816 VDD.n5815 38.9491
R13416 VDD.n5562 VDD.n5561 38.9491
R13417 VDD.n3754 VDD.n3753 38.9491
R13418 VDD.n4012 VDD.n4011 38.9491
R13419 VDD.n4270 VDD.n4269 38.9491
R13420 VDD.n4528 VDD.n4527 38.9491
R13421 VDD.n4786 VDD.n4785 38.9491
R13422 VDD.n5044 VDD.n5043 38.9491
R13423 VDD.n5302 VDD.n5301 38.9491
R13424 VDD.t701 VDD.t795 38.8641
R13425 VDD.t143 VDD.t754 38.8641
R13426 VDD.t1381 VDD.t150 38.534
R13427 VDD.t572 VDD.t504 38.534
R13428 VDD.n1746 VDD.n1745 37.3765
R13429 VDD.n1728 VDD.n1725 37.3765
R13430 VDD.n2095 VDD.n2094 37.3765
R13431 VDD.n2077 VDD.n2074 37.3765
R13432 VDD.n2325 VDD.n2324 37.3765
R13433 VDD.n2307 VDD.n2304 37.3765
R13434 VDD.n2583 VDD.n2582 37.3765
R13435 VDD.n2565 VDD.n2562 37.3765
R13436 VDD.n2841 VDD.n2840 37.3765
R13437 VDD.n2823 VDD.n2820 37.3765
R13438 VDD.n3099 VDD.n3098 37.3765
R13439 VDD.n3081 VDD.n3078 37.3765
R13440 VDD.n3357 VDD.n3356 37.3765
R13441 VDD.n3339 VDD.n3336 37.3765
R13442 VDD.n5680 VDD.n5679 37.3765
R13443 VDD.n5662 VDD.n5659 37.3765
R13444 VDD.n5426 VDD.n5425 37.3765
R13445 VDD.n5408 VDD.n5405 37.3765
R13446 VDD.n3615 VDD.n3614 37.3765
R13447 VDD.n3597 VDD.n3594 37.3765
R13448 VDD.n3873 VDD.n3872 37.3765
R13449 VDD.n3855 VDD.n3852 37.3765
R13450 VDD.n4131 VDD.n4130 37.3765
R13451 VDD.n4113 VDD.n4110 37.3765
R13452 VDD.n4389 VDD.n4388 37.3765
R13453 VDD.n4371 VDD.n4368 37.3765
R13454 VDD.n4647 VDD.n4646 37.3765
R13455 VDD.n4629 VDD.n4626 37.3765
R13456 VDD.n4905 VDD.n4904 37.3765
R13457 VDD.n4887 VDD.n4884 37.3765
R13458 VDD.n5163 VDD.n5162 37.3765
R13459 VDD.n5145 VDD.n5142 37.3765
R13460 VDD.n1830 VDD.t209 36.1587
R13461 VDD.n1830 VDD.t27 36.1587
R13462 VDD.n1813 VDD.t1358 36.1587
R13463 VDD.n1813 VDD.t609 36.1587
R13464 VDD.n2134 VDD.t816 36.1587
R13465 VDD.n2134 VDD.t1176 36.1587
R13466 VDD.n2151 VDD.t837 36.1587
R13467 VDD.n2151 VDD.t1183 36.1587
R13468 VDD.n2392 VDD.t1380 36.1587
R13469 VDD.n2392 VDD.t819 36.1587
R13470 VDD.n2409 VDD.t1501 36.1587
R13471 VDD.n2409 VDD.t723 36.1587
R13472 VDD.n2650 VDD.t873 36.1587
R13473 VDD.n2650 VDD.t1190 36.1587
R13474 VDD.n2667 VDD.t666 36.1587
R13475 VDD.n2667 VDD.t602 36.1587
R13476 VDD.n2908 VDD.t395 36.1587
R13477 VDD.n2908 VDD.t407 36.1587
R13478 VDD.n2925 VDD.t562 36.1587
R13479 VDD.n2925 VDD.t1025 36.1587
R13480 VDD.n3166 VDD.t545 36.1587
R13481 VDD.n3166 VDD.t828 36.1587
R13482 VDD.n3183 VDD.t841 36.1587
R13483 VDD.n3183 VDD.t1483 36.1587
R13484 VDD.n3424 VDD.t619 36.1587
R13485 VDD.n3424 VDD.t664 36.1587
R13486 VDD.n3441 VDD.t1356 36.1587
R13487 VDD.n3441 VDD.t1448 36.1587
R13488 VDD.n5744 VDD.t576 36.1587
R13489 VDD.n5744 VDD.t91 36.1587
R13490 VDD.n5761 VDD.t418 36.1587
R13491 VDD.n5761 VDD.t1196 36.1587
R13492 VDD.n5490 VDD.t1487 36.1587
R13493 VDD.n5490 VDD.t189 36.1587
R13494 VDD.n5507 VDD.t814 36.1587
R13495 VDD.n5507 VDD.t87 36.1587
R13496 VDD.n3682 VDD.t516 36.1587
R13497 VDD.n3682 VDD.t1346 36.1587
R13498 VDD.n3699 VDD.t391 36.1587
R13499 VDD.n3699 VDD.t458 36.1587
R13500 VDD.n3940 VDD.t461 36.1587
R13501 VDD.n3940 VDD.t241 36.1587
R13502 VDD.n3957 VDD.t869 36.1587
R13503 VDD.n3957 VDD.t1442 36.1587
R13504 VDD.n4198 VDD.t895 36.1587
R13505 VDD.n4198 VDD.t3 36.1587
R13506 VDD.n4215 VDD.t605 36.1587
R13507 VDD.n4215 VDD.t726 36.1587
R13508 VDD.n4456 VDD.t794 36.1587
R13509 VDD.n4456 VDD.t1187 36.1587
R13510 VDD.n4473 VDD.t1434 36.1587
R13511 VDD.n4473 VDD.t883 36.1587
R13512 VDD.n4714 VDD.t24 36.1587
R13513 VDD.n4714 VDD.t1370 36.1587
R13514 VDD.n4731 VDD.t875 36.1587
R13515 VDD.n4731 VDD.t1348 36.1587
R13516 VDD.n4972 VDD.t708 36.1587
R13517 VDD.n4972 VDD.t541 36.1587
R13518 VDD.n4989 VDD.t1436 36.1587
R13519 VDD.n4989 VDD.t740 36.1587
R13520 VDD.n5230 VDD.t200 36.1587
R13521 VDD.n5230 VDD.t1185 36.1587
R13522 VDD.n5247 VDD.t154 36.1587
R13523 VDD.n5247 VDD.t237 36.1587
R13524 VDD.t1201 VDD.t1342 35.0774
R13525 VDD.t35 VDD.t25 35.0774
R13526 VDD VDD.n1802 34.927
R13527 VDD VDD.n2010 34.927
R13528 VDD VDD.n2381 34.927
R13529 VDD VDD.n2639 34.927
R13530 VDD VDD.n2897 34.927
R13531 VDD VDD.n3155 34.927
R13532 VDD VDD.n3413 34.927
R13533 VDD VDD.n5736 34.927
R13534 VDD VDD.n5482 34.927
R13535 VDD VDD.n3671 34.927
R13536 VDD VDD.n3929 34.927
R13537 VDD VDD.n4187 34.927
R13538 VDD VDD.n4445 34.927
R13539 VDD VDD.n4703 34.927
R13540 VDD VDD.n4961 34.927
R13541 VDD VDD.n5219 34.927
R13542 VDD.n23 VDD.n2 34.6358
R13543 VDD.n18 VDD.n6 34.6358
R13544 VDD.n679 VDD.n678 34.6358
R13545 VDD.n500 VDD.n499 34.6358
R13546 VDD.n427 VDD.n426 34.6358
R13547 VDD.n98 VDD.n97 34.6358
R13548 VDD.n1167 VDD.n1146 34.6358
R13549 VDD.n1162 VDD.n1150 34.6358
R13550 VDD.n1585 VDD.n1584 34.6358
R13551 VDD.n832 VDD.n831 34.6358
R13552 VDD.n844 VDD.n843 34.6358
R13553 VDD.n850 VDD.n849 34.6358
R13554 VDD.n813 VDD.n801 34.6358
R13555 VDD.n817 VDD.n801 34.6358
R13556 VDD.n818 VDD.n817 34.6358
R13557 VDD.n811 VDD.n804 34.6358
R13558 VDD.n1029 VDD.n1028 34.6358
R13559 VDD.n274 VDD.n273 34.6358
R13560 VDD.n1215 VDD.n1214 34.6358
R13561 VDD.n1227 VDD.n1226 34.6358
R13562 VDD.n1233 VDD.n1232 34.6358
R13563 VDD.n1196 VDD.n1184 34.6358
R13564 VDD.n1200 VDD.n1184 34.6358
R13565 VDD.n1201 VDD.n1200 34.6358
R13566 VDD.n1194 VDD.n1187 34.6358
R13567 VDD.n667 VDD.t1071 33.9291
R13568 VDD.n1017 VDD.t942 33.9291
R13569 VDD.n838 VDD.n837 33.8829
R13570 VDD.n1221 VDD.n1220 33.8829
R13571 VDD.n1958 VDD.n1957 33.8422
R13572 VDD.n1397 VDD.t673 33.8361
R13573 VDD.n1973 VDD.n1923 33.6292
R13574 VDD.t232 VDD.t699 32.6058
R13575 VDD.t1177 VDD.t141 32.6058
R13576 VDD.t148 VDD.t462 31.4862
R13577 VDD.t114 VDD.t404 31.4862
R13578 VDD.t145 VDD.t155 31.4862
R13579 VDD.t33 VDD.t159 31.4862
R13580 VDD.n1914 VDD.t28 30.1961
R13581 VDD.n2235 VDD.t103 30.1961
R13582 VDD.n2493 VDD.t471 30.1961
R13583 VDD.n2751 VDD.t184 30.1961
R13584 VDD.n3009 VDD.t488 30.1961
R13585 VDD.n3267 VDD.t234 30.1961
R13586 VDD.n3525 VDD.t18 30.1961
R13587 VDD.n5845 VDD.t746 30.1961
R13588 VDD.n5591 VDD.t88 30.1961
R13589 VDD.n3783 VDD.t82 30.1961
R13590 VDD.n4041 VDD.t409 30.1961
R13591 VDD.n4299 VDD.t727 30.1961
R13592 VDD.n4557 VDD.t122 30.1961
R13593 VDD.n4815 VDD.t484 30.1961
R13594 VDD.n5073 VDD.t14 30.1961
R13595 VDD.n5331 VDD.t119 30.1961
R13596 VDD.n542 VDD.n541 29.3652
R13597 VDD.n621 VDD.n620 29.3652
R13598 VDD.n517 VDD.n516 29.3652
R13599 VDD.n520 VDD.n519 29.3652
R13600 VDD.n892 VDD.n891 29.3652
R13601 VDD.n971 VDD.n970 29.3652
R13602 VDD.n867 VDD.n866 29.3652
R13603 VDD.n870 VDD.n869 29.3652
R13604 VDD.n141 VDD.n140 29.3652
R13605 VDD.n220 VDD.n219 29.3652
R13606 VDD.n116 VDD.n115 29.3652
R13607 VDD.n119 VDD.n118 29.3652
R13608 VDD.n1313 VDD.n1312 29.3652
R13609 VDD.n1342 VDD.n1341 29.3652
R13610 VDD.n523 VDD.n522 28.9887
R13611 VDD.n873 VDD.n872 28.9887
R13612 VDD.n122 VDD.n121 28.9887
R13613 VDD.n1348 VDD.n1347 28.9887
R13614 VDD.n5 VDD.t1382 28.4628
R13615 VDD.n494 VDD.t22 28.4628
R13616 VDD.n422 VDD.t211 28.4628
R13617 VDD.n418 VDD.t750 28.4628
R13618 VDD.n401 VDD.t507 28.4628
R13619 VDD.n92 VDD.t752 28.4628
R13620 VDD.n1149 VDD.t573 28.4628
R13621 VDD.n1580 VDD.t877 28.4628
R13622 VDD.n1576 VDD.t101 28.4628
R13623 VDD.n1559 VDD.t213 28.4628
R13624 VDD.n806 VDD.t560 28.4628
R13625 VDD.n1189 VDD.t20 28.4628
R13626 VDD.n1793 VDD.n1782 28.2358
R13627 VDD.n1794 VDD.n1793 28.2358
R13628 VDD.n1790 VDD.n1787 28.2358
R13629 VDD.n1790 VDD.n1789 28.2358
R13630 VDD.n2001 VDD.n1990 28.2358
R13631 VDD.n2002 VDD.n2001 28.2358
R13632 VDD.n1998 VDD.n1995 28.2358
R13633 VDD.n1998 VDD.n1997 28.2358
R13634 VDD.n2372 VDD.n2361 28.2358
R13635 VDD.n2373 VDD.n2372 28.2358
R13636 VDD.n2369 VDD.n2366 28.2358
R13637 VDD.n2369 VDD.n2368 28.2358
R13638 VDD.n2630 VDD.n2619 28.2358
R13639 VDD.n2631 VDD.n2630 28.2358
R13640 VDD.n2627 VDD.n2624 28.2358
R13641 VDD.n2627 VDD.n2626 28.2358
R13642 VDD.n2888 VDD.n2877 28.2358
R13643 VDD.n2889 VDD.n2888 28.2358
R13644 VDD.n2885 VDD.n2882 28.2358
R13645 VDD.n2885 VDD.n2884 28.2358
R13646 VDD.n3146 VDD.n3135 28.2358
R13647 VDD.n3147 VDD.n3146 28.2358
R13648 VDD.n3143 VDD.n3140 28.2358
R13649 VDD.n3143 VDD.n3142 28.2358
R13650 VDD.n3404 VDD.n3393 28.2358
R13651 VDD.n3405 VDD.n3404 28.2358
R13652 VDD.n3401 VDD.n3398 28.2358
R13653 VDD.n3401 VDD.n3400 28.2358
R13654 VDD.n5727 VDD.n5716 28.2358
R13655 VDD.n5728 VDD.n5727 28.2358
R13656 VDD.n5724 VDD.n5721 28.2358
R13657 VDD.n5724 VDD.n5723 28.2358
R13658 VDD.n5473 VDD.n5462 28.2358
R13659 VDD.n5474 VDD.n5473 28.2358
R13660 VDD.n5470 VDD.n5467 28.2358
R13661 VDD.n5470 VDD.n5469 28.2358
R13662 VDD.n3662 VDD.n3651 28.2358
R13663 VDD.n3663 VDD.n3662 28.2358
R13664 VDD.n3659 VDD.n3656 28.2358
R13665 VDD.n3659 VDD.n3658 28.2358
R13666 VDD.n3920 VDD.n3909 28.2358
R13667 VDD.n3921 VDD.n3920 28.2358
R13668 VDD.n3917 VDD.n3914 28.2358
R13669 VDD.n3917 VDD.n3916 28.2358
R13670 VDD.n4178 VDD.n4167 28.2358
R13671 VDD.n4179 VDD.n4178 28.2358
R13672 VDD.n4175 VDD.n4172 28.2358
R13673 VDD.n4175 VDD.n4174 28.2358
R13674 VDD.n4436 VDD.n4425 28.2358
R13675 VDD.n4437 VDD.n4436 28.2358
R13676 VDD.n4433 VDD.n4430 28.2358
R13677 VDD.n4433 VDD.n4432 28.2358
R13678 VDD.n4694 VDD.n4683 28.2358
R13679 VDD.n4695 VDD.n4694 28.2358
R13680 VDD.n4691 VDD.n4688 28.2358
R13681 VDD.n4691 VDD.n4690 28.2358
R13682 VDD.n4952 VDD.n4941 28.2358
R13683 VDD.n4953 VDD.n4952 28.2358
R13684 VDD.n4949 VDD.n4946 28.2358
R13685 VDD.n4949 VDD.n4948 28.2358
R13686 VDD.n5210 VDD.n5199 28.2358
R13687 VDD.n5211 VDD.n5210 28.2358
R13688 VDD.n5207 VDD.n5204 28.2358
R13689 VDD.n5207 VDD.n5206 28.2358
R13690 VDD.n13 VDD.n8 28.2358
R13691 VDD.n1157 VDD.n1152 28.2358
R13692 VDD.n463 VDD 28.2291
R13693 VDD.n60 VDD 28.2291
R13694 VDD.n262 VDD.t265 27.1434
R13695 VDD.n482 VDD.t509 26.9729
R13696 VDD.n80 VDD.t792 26.9729
R13697 VDD.n1835 VDD.n1834 26.8623
R13698 VDD.n2156 VDD.n2155 26.8623
R13699 VDD.n2414 VDD.n2413 26.8623
R13700 VDD.n2672 VDD.n2671 26.8623
R13701 VDD.n2930 VDD.n2929 26.8623
R13702 VDD.n3188 VDD.n3187 26.8623
R13703 VDD.n3446 VDD.n3445 26.8623
R13704 VDD.n5766 VDD.n5765 26.8623
R13705 VDD.n5512 VDD.n5511 26.8623
R13706 VDD.n3704 VDD.n3703 26.8623
R13707 VDD.n3962 VDD.n3961 26.8623
R13708 VDD.n4220 VDD.n4219 26.8623
R13709 VDD.n4478 VDD.n4477 26.8623
R13710 VDD.n4736 VDD.n4735 26.8623
R13711 VDD.n4994 VDD.n4993 26.8623
R13712 VDD.n5252 VDD.n5251 26.8623
R13713 VDD.n1656 VDD 26.615
R13714 VDD.n31 VDD.t821 26.5955
R13715 VDD.n508 VDD.t1431 26.5955
R13716 VDD.n435 VDD.t387 26.5955
R13717 VDD.n404 VDD.t630 26.5955
R13718 VDD.n106 VDD.t607 26.5955
R13719 VDD.n1175 VDD.t1440 26.5955
R13720 VDD.n1593 VDD.t1444 26.5955
R13721 VDD.n1562 VDD.t558 26.5955
R13722 VDD.n800 VDD.t469 26.5955
R13723 VDD.n803 VDD.t1040 26.5955
R13724 VDD.n1183 VDD.t511 26.5955
R13725 VDD.n1186 VDD.t204 26.5955
R13726 VDD.n1792 VDD.t1365 26.5955
R13727 VDD.n1792 VDD.t1362 26.5955
R13728 VDD.n1788 VDD.t641 26.5955
R13729 VDD.n1788 VDD.t645 26.5955
R13730 VDD.n2000 VDD.t1492 26.5955
R13731 VDD.n2000 VDD.t1496 26.5955
R13732 VDD.n1996 VDD.t249 26.5955
R13733 VDD.n1996 VDD.t246 26.5955
R13734 VDD.n2371 VDD.t224 26.5955
R13735 VDD.n2371 VDD.t226 26.5955
R13736 VDD.n2367 VDD.t627 26.5955
R13737 VDD.n2367 VDD.t622 26.5955
R13738 VDD.n2629 VDD.t59 26.5955
R13739 VDD.n2629 VDD.t60 26.5955
R13740 VDD.n2625 VDD.t846 26.5955
R13741 VDD.n2625 VDD.t848 26.5955
R13742 VDD.n2887 VDD.t597 26.5955
R13743 VDD.n2887 VDD.t599 26.5955
R13744 VDD.n2883 VDD.t133 26.5955
R13745 VDD.n2883 VDD.t136 26.5955
R13746 VDD.n3145 VDD.t43 26.5955
R13747 VDD.n3145 VDD.t45 26.5955
R13748 VDD.n3141 VDD.t480 26.5955
R13749 VDD.n3141 VDD.t476 26.5955
R13750 VDD.n3403 VDD.t733 26.5955
R13751 VDD.n3403 VDD.t735 26.5955
R13752 VDD.n3399 VDD.t1335 26.5955
R13753 VDD.n3399 VDD.t1337 26.5955
R13754 VDD.n5726 VDD.t166 26.5955
R13755 VDD.n5726 VDD.t168 26.5955
R13756 VDD.n5722 VDD.t612 26.5955
R13757 VDD.n5722 VDD.t615 26.5955
R13758 VDD.n5472 VDD.t524 26.5955
R13759 VDD.n5472 VDD.t520 26.5955
R13760 VDD.n5468 VDD.t9 26.5955
R13761 VDD.n5468 VDD.t11 26.5955
R13762 VDD.n3661 VDD.t196 26.5955
R13763 VDD.n3661 VDD.t198 26.5955
R13764 VDD.n3657 VDD.t635 26.5955
R13765 VDD.n3657 VDD.t637 26.5955
R13766 VDD.n3919 VDD.t172 26.5955
R13767 VDD.n3919 VDD.t175 26.5955
R13768 VDD.n3915 VDD.t1389 26.5955
R13769 VDD.n3915 VDD.t1384 26.5955
R13770 VDD.n4177 VDD.t99 26.5955
R13771 VDD.n4177 VDD.t95 26.5955
R13772 VDD.n4173 VDD.t891 26.5955
R13773 VDD.n4173 VDD.t886 26.5955
R13774 VDD.n4435 VDD.t499 26.5955
R13775 VDD.n4435 VDD.t501 26.5955
R13776 VDD.n4431 VDD.t125 26.5955
R13777 VDD.n4431 VDD.t128 26.5955
R13778 VDD.n4693 VDD.t589 26.5955
R13779 VDD.n4693 VDD.t591 26.5955
R13780 VDD.n4689 VDD.t79 26.5955
R13781 VDD.n4689 VDD.t75 26.5955
R13782 VDD.n4951 VDD.t581 26.5955
R13783 VDD.n4951 VDD.t583 26.5955
R13784 VDD.n4947 VDD.t787 26.5955
R13785 VDD.n4947 VDD.t789 26.5955
R13786 VDD.n5209 VDD.t859 26.5955
R13787 VDD.n5209 VDD.t861 26.5955
R13788 VDD.n5205 VDD.t1373 26.5955
R13789 VDD.n5205 VDD.t1376 26.5955
R13790 VDD.n692 VDD.t569 26.5955
R13791 VDD.n692 VDD.t571 26.5955
R13792 VDD.n555 VDD.t1168 26.5955
R13793 VDD.n555 VDD.t1100 26.5955
R13794 VDD.n561 VDD.t1074 26.5955
R13795 VDD.n561 VDD.t1138 26.5955
R13796 VDD.n567 VDD.t1154 26.5955
R13797 VDD.n567 VDD.t1050 26.5955
R13798 VDD.n573 VDD.t1048 26.5955
R13799 VDD.n573 VDD.t1084 26.5955
R13800 VDD.n578 VDD.t1080 26.5955
R13801 VDD.n578 VDD.t1106 26.5955
R13802 VDD.n534 VDD.t1066 26.5955
R13803 VDD.n534 VDD.t1058 26.5955
R13804 VDD.n529 VDD.t1088 26.5955
R13805 VDD.n529 VDD.t1174 26.5955
R13806 VDD.n613 VDD.t1172 26.5955
R13807 VDD.n613 VDD.t1104 26.5955
R13808 VDD.n607 VDD.t1098 26.5955
R13809 VDD.n607 VDD.t1124 26.5955
R13810 VDD.n601 VDD.t1086 26.5955
R13811 VDD.n601 VDD.t1166 26.5955
R13812 VDD.n595 VDD.t1116 26.5955
R13813 VDD.n595 VDD.t1150 26.5955
R13814 VDD.n591 VDD.t1146 26.5955
R13815 VDD.n591 VDD.t1078 26.5955
R13816 VDD.n525 VDD.t1056 26.5955
R13817 VDD.n525 VDD.t1112 26.5955
R13818 VDD.n545 VDD.t1132 26.5955
R13819 VDD.n545 VDD.t1158 26.5955
R13820 VDD.n638 VDD.t1068 26.5955
R13821 VDD.n638 VDD.t1090 26.5955
R13822 VDD.n644 VDD.t1096 26.5955
R13823 VDD.n644 VDD.t1122 26.5955
R13824 VDD.n650 VDD.t1120 26.5955
R13825 VDD.n650 VDD.t1152 26.5955
R13826 VDD.n656 VDD.t1164 26.5955
R13827 VDD.n656 VDD.t1094 26.5955
R13828 VDD.n661 VDD.t1072 26.5955
R13829 VDD.n661 VDD.t1136 26.5955
R13830 VDD.n631 VDD.t1076 26.5955
R13831 VDD.n631 VDD.t1162 26.5955
R13832 VDD.n625 VDD.t1110 26.5955
R13833 VDD.n625 VDD.t1140 26.5955
R13834 VDD.n748 VDD.t1102 26.5955
R13835 VDD.n748 VDD.t1126 26.5955
R13836 VDD.n754 VDD.t1142 26.5955
R13837 VDD.n754 VDD.t1170 26.5955
R13838 VDD.n760 VDD.t1118 26.5955
R13839 VDD.n760 VDD.t1060 26.5955
R13840 VDD.n766 VDD.t1148 26.5955
R13841 VDD.n766 VDD.t1082 26.5955
R13842 VDD.n770 VDD.t1092 26.5955
R13843 VDD.n770 VDD.t1114 26.5955
R13844 VDD.n777 VDD.t1134 26.5955
R13845 VDD.n777 VDD.t1160 26.5955
R13846 VDD.n785 VDD.t1156 26.5955
R13847 VDD.n785 VDD.t1054 26.5955
R13848 VDD.n701 VDD.t1455 26.5955
R13849 VDD.n701 VDD.t1469 26.5955
R13850 VDD.n707 VDD.t1467 26.5955
R13851 VDD.n707 VDD.t1451 26.5955
R13852 VDD.n713 VDD.t1481 26.5955
R13853 VDD.n713 VDD.t1461 26.5955
R13854 VDD.n719 VDD.t1459 26.5955
R13855 VDD.n719 VDD.t1473 26.5955
R13856 VDD.n723 VDD.t1471 26.5955
R13857 VDD.n723 VDD.t1479 26.5955
R13858 VDD.n729 VDD.t1465 26.5955
R13859 VDD.n729 VDD.t1475 26.5955
R13860 VDD.n737 VDD.t1477 26.5955
R13861 VDD.n737 VDD.t1457 26.5955
R13862 VDD.n1042 VDD.t54 26.5955
R13863 VDD.n1042 VDD.t48 26.5955
R13864 VDD.n905 VDD.t911 26.5955
R13865 VDD.n905 VDD.t971 26.5955
R13866 VDD.n911 VDD.t945 26.5955
R13867 VDD.n911 VDD.t1009 26.5955
R13868 VDD.n917 VDD.t897 26.5955
R13869 VDD.n917 VDD.t921 26.5955
R13870 VDD.n923 VDD.t919 26.5955
R13871 VDD.n923 VDD.t955 26.5955
R13872 VDD.n928 VDD.t949 26.5955
R13873 VDD.n928 VDD.t977 26.5955
R13874 VDD.n884 VDD.t937 26.5955
R13875 VDD.n884 VDD.t929 26.5955
R13876 VDD.n879 VDD.t959 26.5955
R13877 VDD.n879 VDD.t917 26.5955
R13878 VDD.n963 VDD.t915 26.5955
R13879 VDD.n963 VDD.t975 26.5955
R13880 VDD.n957 VDD.t969 26.5955
R13881 VDD.n957 VDD.t997 26.5955
R13882 VDD.n951 VDD.t957 26.5955
R13883 VDD.n951 VDD.t909 26.5955
R13884 VDD.n945 VDD.t989 26.5955
R13885 VDD.n945 VDD.t1021 26.5955
R13886 VDD.n941 VDD.t1017 26.5955
R13887 VDD.n941 VDD.t951 26.5955
R13888 VDD.n875 VDD.t927 26.5955
R13889 VDD.n875 VDD.t985 26.5955
R13890 VDD.n895 VDD.t983 26.5955
R13891 VDD.n895 VDD.t901 26.5955
R13892 VDD.n988 VDD.t939 26.5955
R13893 VDD.n988 VDD.t963 26.5955
R13894 VDD.n994 VDD.t967 26.5955
R13895 VDD.n994 VDD.t995 26.5955
R13896 VDD.n1000 VDD.t993 26.5955
R13897 VDD.n1000 VDD.t1023 26.5955
R13898 VDD.n1006 VDD.t907 26.5955
R13899 VDD.n1006 VDD.t961 26.5955
R13900 VDD.n1011 VDD.t943 26.5955
R13901 VDD.n1011 VDD.t1007 26.5955
R13902 VDD.n981 VDD.t947 26.5955
R13903 VDD.n981 VDD.t905 26.5955
R13904 VDD.n975 VDD.t981 26.5955
R13905 VDD.n975 VDD.t1011 26.5955
R13906 VDD.n1098 VDD.t973 26.5955
R13907 VDD.n1098 VDD.t999 26.5955
R13908 VDD.n1104 VDD.t1013 26.5955
R13909 VDD.n1104 VDD.t913 26.5955
R13910 VDD.n1110 VDD.t991 26.5955
R13911 VDD.n1110 VDD.t931 26.5955
R13912 VDD.n1116 VDD.t1019 26.5955
R13913 VDD.n1116 VDD.t953 26.5955
R13914 VDD.n1120 VDD.t965 26.5955
R13915 VDD.n1120 VDD.t987 26.5955
R13916 VDD.n1127 VDD.t1005 26.5955
R13917 VDD.n1127 VDD.t903 26.5955
R13918 VDD.n1135 VDD.t899 26.5955
R13919 VDD.n1135 VDD.t925 26.5955
R13920 VDD.n1051 VDD.t1409 26.5955
R13921 VDD.n1051 VDD.t1423 26.5955
R13922 VDD.n1057 VDD.t1421 26.5955
R13923 VDD.n1057 VDD.t1405 26.5955
R13924 VDD.n1063 VDD.t1403 26.5955
R13925 VDD.n1063 VDD.t1415 26.5955
R13926 VDD.n1069 VDD.t1413 26.5955
R13927 VDD.n1069 VDD.t1427 26.5955
R13928 VDD.n1073 VDD.t1425 26.5955
R13929 VDD.n1073 VDD.t1401 26.5955
R13930 VDD.n1079 VDD.t1419 26.5955
R13931 VDD.n1079 VDD.t1429 26.5955
R13932 VDD.n1087 VDD.t1399 26.5955
R13933 VDD.n1087 VDD.t1411 26.5955
R13934 VDD.n287 VDD.t67 26.5955
R13935 VDD.n287 VDD.t69 26.5955
R13936 VDD.n154 VDD.t362 26.5955
R13937 VDD.n154 VDD.t294 26.5955
R13938 VDD.n160 VDD.t268 26.5955
R13939 VDD.n160 VDD.t332 26.5955
R13940 VDD.n166 VDD.t348 26.5955
R13941 VDD.n166 VDD.t372 26.5955
R13942 VDD.n172 VDD.t370 26.5955
R13943 VDD.n172 VDD.t280 26.5955
R13944 VDD.n177 VDD.t272 26.5955
R13945 VDD.n177 VDD.t300 26.5955
R13946 VDD.n133 VDD.t260 26.5955
R13947 VDD.n133 VDD.t380 26.5955
R13948 VDD.n128 VDD.t282 26.5955
R13949 VDD.n128 VDD.t368 26.5955
R13950 VDD.n212 VDD.t366 26.5955
R13951 VDD.n212 VDD.t298 26.5955
R13952 VDD.n206 VDD.t292 26.5955
R13953 VDD.n206 VDD.t318 26.5955
R13954 VDD.n200 VDD.t278 26.5955
R13955 VDD.n200 VDD.t360 26.5955
R13956 VDD.n194 VDD.t310 26.5955
R13957 VDD.n194 VDD.t344 26.5955
R13958 VDD.n190 VDD.t340 26.5955
R13959 VDD.n190 VDD.t274 26.5955
R13960 VDD.n124 VDD.t378 26.5955
R13961 VDD.n124 VDD.t306 26.5955
R13962 VDD.n144 VDD.t326 26.5955
R13963 VDD.n144 VDD.t352 26.5955
R13964 VDD.n111 VDD.t262 26.5955
R13965 VDD.n111 VDD.t284 26.5955
R13966 VDD.n239 VDD.t290 26.5955
R13967 VDD.n239 VDD.t316 26.5955
R13968 VDD.n245 VDD.t314 26.5955
R13969 VDD.n245 VDD.t346 26.5955
R13970 VDD.n251 VDD.t358 26.5955
R13971 VDD.n251 VDD.t288 26.5955
R13972 VDD.n256 VDD.t266 26.5955
R13973 VDD.n256 VDD.t330 26.5955
R13974 VDD.n230 VDD.t270 26.5955
R13975 VDD.n230 VDD.t356 26.5955
R13976 VDD.n224 VDD.t304 26.5955
R13977 VDD.n224 VDD.t334 26.5955
R13978 VDD.n343 VDD.t296 26.5955
R13979 VDD.n343 VDD.t320 26.5955
R13980 VDD.n349 VDD.t336 26.5955
R13981 VDD.n349 VDD.t364 26.5955
R13982 VDD.n355 VDD.t312 26.5955
R13983 VDD.n355 VDD.t254 26.5955
R13984 VDD.n361 VDD.t342 26.5955
R13985 VDD.n361 VDD.t276 26.5955
R13986 VDD.n365 VDD.t286 26.5955
R13987 VDD.n365 VDD.t308 26.5955
R13988 VDD.n372 VDD.t328 26.5955
R13989 VDD.n372 VDD.t354 26.5955
R13990 VDD.n380 VDD.t350 26.5955
R13991 VDD.n380 VDD.t376 26.5955
R13992 VDD.n296 VDD.t430 26.5955
R13993 VDD.n296 VDD.t444 26.5955
R13994 VDD.n302 VDD.t442 26.5955
R13995 VDD.n302 VDD.t426 26.5955
R13996 VDD.n308 VDD.t456 26.5955
R13997 VDD.n308 VDD.t436 26.5955
R13998 VDD.n314 VDD.t434 26.5955
R13999 VDD.n314 VDD.t448 26.5955
R14000 VDD.n318 VDD.t446 26.5955
R14001 VDD.n318 VDD.t454 26.5955
R14002 VDD.n324 VDD.t440 26.5955
R14003 VDD.n324 VDD.t450 26.5955
R14004 VDD.n332 VDD.t452 26.5955
R14005 VDD.n332 VDD.t432 26.5955
R14006 VDD.n1352 VDD.t656 26.5955
R14007 VDD.n1352 VDD.t658 26.5955
R14008 VDD.n1334 VDD.t1220 26.5955
R14009 VDD.n1334 VDD.t1246 26.5955
R14010 VDD.n1328 VDD.t1242 26.5955
R14011 VDD.n1328 VDD.t1274 26.5955
R14012 VDD.n1321 VDD.t1290 26.5955
R14013 VDD.n1321 VDD.t1216 26.5955
R14014 VDD.n1434 VDD.t1330 26.5955
R14015 VDD.n1434 VDD.t1258 26.5955
R14016 VDD.n1438 VDD.t1254 26.5955
R14017 VDD.n1438 VDD.t1286 26.5955
R14018 VDD.n1444 VDD.t1230 26.5955
R14019 VDD.n1444 VDD.t1326 26.5955
R14020 VDD.n1450 VDD.t1278 26.5955
R14021 VDD.n1450 VDD.t1308 26.5955
R14022 VDD.n1378 VDD.t682 26.5955
R14023 VDD.n1378 VDD.t690 26.5955
R14024 VDD.n1384 VDD.t694 26.5955
R14025 VDD.n1384 VDD.t672 26.5955
R14026 VDD.n1390 VDD.t684 26.5955
R14027 VDD.n1390 VDD.t680 26.5955
R14028 VDD.n1402 VDD.t668 26.5955
R14029 VDD.n1402 VDD.t674 26.5955
R14030 VDD.n1407 VDD.t678 26.5955
R14031 VDD.n1407 VDD.t688 26.5955
R14032 VDD.n1413 VDD.t686 26.5955
R14033 VDD.n1413 VDD.t696 26.5955
R14034 VDD.n1419 VDD.t698 26.5955
R14035 VDD.n1419 VDD.t676 26.5955
R14036 VDD.n1305 VDD.t1222 26.5955
R14037 VDD.n1305 VDD.t1248 26.5955
R14038 VDD.n1298 VDD.t1264 26.5955
R14039 VDD.n1298 VDD.t1296 26.5955
R14040 VDD.n1292 VDD.t1238 26.5955
R14041 VDD.n1292 VDD.t1204 26.5955
R14042 VDD.n1267 VDD.t1270 26.5955
R14043 VDD.n1267 VDD.t1206 26.5955
R14044 VDD.n1271 VDD.t1312 26.5955
R14045 VDD.n1271 VDD.t1234 26.5955
R14046 VDD.n1277 VDD.t1252 26.5955
R14047 VDD.n1277 VDD.t1284 26.5955
R14048 VDD.n1264 VDD.t1280 26.5955
R14049 VDD.n1264 VDD.t1322 26.5955
R14050 VDD.n1464 VDD.t1276 26.5955
R14051 VDD.n1464 VDD.t1212 26.5955
R14052 VDD.n1470 VDD.t1218 26.5955
R14053 VDD.n1470 VDD.t1244 26.5955
R14054 VDD.n1476 VDD.t1240 26.5955
R14055 VDD.n1476 VDD.t1292 26.5955
R14056 VDD.n1482 VDD.t1288 26.5955
R14057 VDD.n1482 VDD.t1316 26.5955
R14058 VDD.n1486 VDD.t1328 26.5955
R14059 VDD.n1486 VDD.t1256 26.5955
R14060 VDD.n1492 VDD.t1214 26.5955
R14061 VDD.n1492 VDD.t1304 26.5955
R14062 VDD.n1498 VDD.t1228 26.5955
R14063 VDD.n1498 VDD.t1262 26.5955
R14064 VDD.n1514 VDD.t1298 26.5955
R14065 VDD.n1514 VDD.t1224 26.5955
R14066 VDD.n1520 VDD.t1318 26.5955
R14067 VDD.n1520 VDD.t1266 26.5955
R14068 VDD.n1256 VDD.t1260 26.5955
R14069 VDD.n1256 VDD.t1294 26.5955
R14070 VDD.n1530 VDD.t1236 26.5955
R14071 VDD.n1530 VDD.t1272 26.5955
R14072 VDD.n1534 VDD.t1268 26.5955
R14073 VDD.n1534 VDD.t1314 26.5955
R14074 VDD.n1252 VDD.t1310 26.5955
R14075 VDD.n1252 VDD.t1232 26.5955
R14076 VDD.n1247 VDD.t1210 26.5955
R14077 VDD.n1247 VDD.t1282 26.5955
R14078 VDD.n812 VDD.n811 25.977
R14079 VDD.n1195 VDD.n1194 25.977
R14080 VDD.t492 VDD.t508 25.9096
R14081 VDD.t853 VDD.t791 25.9096
R14082 VDD.n672 VDD.t219 25.6105
R14083 VDD.n1022 VDD.t1368 25.6105
R14084 VDD.n267 VDD.t706 25.6105
R14085 VDD.n819 VDD.n818 25.224
R14086 VDD.n1202 VDD.n1201 25.224
R14087 VDD.t106 VDD.n1847 24.3893
R14088 VDD.t719 VDD.n2168 24.3893
R14089 VDD.t485 VDD.n2426 24.3893
R14090 VDD.t531 VDD.n2684 24.3893
R14091 VDD.t15 VDD.n2942 24.3893
R14092 VDD.t412 VDD.n3200 24.3893
R14093 VDD.t538 VDD.n3458 24.3893
R14094 VDD.t109 VDD.n5778 24.3893
R14095 VDD.t186 VDD.n5524 24.3893
R14096 VDD.t413 VDD.n3716 24.3893
R14097 VDD.t108 VDD.n3974 24.3893
R14098 VDD.t0 VDD.n4232 24.3893
R14099 VDD.t13 VDD.n4490 24.3893
R14100 VDD.t117 VDD.n4748 24.3893
R14101 VDD.t651 VDD.n5006 24.3893
R14102 VDD.t85 VDD.n5264 24.3893
R14103 VDD.t1029 VDD.t490 23.0308
R14104 VDD.t206 VDD.t850 23.0308
R14105 VDD.n408 VDD 22.7027
R14106 VDD.n1566 VDD 22.7027
R14107 VDD.n1660 VDD.n1626 22.5125
R14108 VDD.n1834 VDD.n1833 22.2123
R14109 VDD.n1814 VDD.n1812 22.2123
R14110 VDD.n1784 VDD.n1782 22.2123
R14111 VDD.n1795 VDD.n1794 22.2123
R14112 VDD.n1787 VDD.n1786 22.2123
R14113 VDD.n1789 VDD.n1781 22.2123
R14114 VDD.n2135 VDD.n2133 22.2123
R14115 VDD.n2155 VDD.n2154 22.2123
R14116 VDD.n1992 VDD.n1990 22.2123
R14117 VDD.n2003 VDD.n2002 22.2123
R14118 VDD.n1995 VDD.n1994 22.2123
R14119 VDD.n1997 VDD.n1989 22.2123
R14120 VDD.n2393 VDD.n2391 22.2123
R14121 VDD.n2413 VDD.n2412 22.2123
R14122 VDD.n2363 VDD.n2361 22.2123
R14123 VDD.n2374 VDD.n2373 22.2123
R14124 VDD.n2366 VDD.n2365 22.2123
R14125 VDD.n2368 VDD.n2360 22.2123
R14126 VDD.n2651 VDD.n2649 22.2123
R14127 VDD.n2671 VDD.n2670 22.2123
R14128 VDD.n2621 VDD.n2619 22.2123
R14129 VDD.n2632 VDD.n2631 22.2123
R14130 VDD.n2624 VDD.n2623 22.2123
R14131 VDD.n2626 VDD.n2618 22.2123
R14132 VDD.n2909 VDD.n2907 22.2123
R14133 VDD.n2929 VDD.n2928 22.2123
R14134 VDD.n2879 VDD.n2877 22.2123
R14135 VDD.n2890 VDD.n2889 22.2123
R14136 VDD.n2882 VDD.n2881 22.2123
R14137 VDD.n2884 VDD.n2876 22.2123
R14138 VDD.n3167 VDD.n3165 22.2123
R14139 VDD.n3187 VDD.n3186 22.2123
R14140 VDD.n3137 VDD.n3135 22.2123
R14141 VDD.n3148 VDD.n3147 22.2123
R14142 VDD.n3140 VDD.n3139 22.2123
R14143 VDD.n3142 VDD.n3134 22.2123
R14144 VDD.n3425 VDD.n3423 22.2123
R14145 VDD.n3445 VDD.n3444 22.2123
R14146 VDD.n3395 VDD.n3393 22.2123
R14147 VDD.n3406 VDD.n3405 22.2123
R14148 VDD.n3398 VDD.n3397 22.2123
R14149 VDD.n3400 VDD.n3392 22.2123
R14150 VDD.n5745 VDD.n5743 22.2123
R14151 VDD.n5765 VDD.n5764 22.2123
R14152 VDD.n5718 VDD.n5716 22.2123
R14153 VDD.n5729 VDD.n5728 22.2123
R14154 VDD.n5721 VDD.n5720 22.2123
R14155 VDD.n5723 VDD.n5715 22.2123
R14156 VDD.n5491 VDD.n5489 22.2123
R14157 VDD.n5511 VDD.n5510 22.2123
R14158 VDD.n5464 VDD.n5462 22.2123
R14159 VDD.n5475 VDD.n5474 22.2123
R14160 VDD.n5467 VDD.n5466 22.2123
R14161 VDD.n5469 VDD.n5461 22.2123
R14162 VDD.n3683 VDD.n3681 22.2123
R14163 VDD.n3703 VDD.n3702 22.2123
R14164 VDD.n3653 VDD.n3651 22.2123
R14165 VDD.n3664 VDD.n3663 22.2123
R14166 VDD.n3656 VDD.n3655 22.2123
R14167 VDD.n3658 VDD.n3650 22.2123
R14168 VDD.n3941 VDD.n3939 22.2123
R14169 VDD.n3961 VDD.n3960 22.2123
R14170 VDD.n3911 VDD.n3909 22.2123
R14171 VDD.n3922 VDD.n3921 22.2123
R14172 VDD.n3914 VDD.n3913 22.2123
R14173 VDD.n3916 VDD.n3908 22.2123
R14174 VDD.n4199 VDD.n4197 22.2123
R14175 VDD.n4219 VDD.n4218 22.2123
R14176 VDD.n4169 VDD.n4167 22.2123
R14177 VDD.n4180 VDD.n4179 22.2123
R14178 VDD.n4172 VDD.n4171 22.2123
R14179 VDD.n4174 VDD.n4166 22.2123
R14180 VDD.n4457 VDD.n4455 22.2123
R14181 VDD.n4477 VDD.n4476 22.2123
R14182 VDD.n4427 VDD.n4425 22.2123
R14183 VDD.n4438 VDD.n4437 22.2123
R14184 VDD.n4430 VDD.n4429 22.2123
R14185 VDD.n4432 VDD.n4424 22.2123
R14186 VDD.n4715 VDD.n4713 22.2123
R14187 VDD.n4735 VDD.n4734 22.2123
R14188 VDD.n4685 VDD.n4683 22.2123
R14189 VDD.n4696 VDD.n4695 22.2123
R14190 VDD.n4688 VDD.n4687 22.2123
R14191 VDD.n4690 VDD.n4682 22.2123
R14192 VDD.n4973 VDD.n4971 22.2123
R14193 VDD.n4993 VDD.n4992 22.2123
R14194 VDD.n4943 VDD.n4941 22.2123
R14195 VDD.n4954 VDD.n4953 22.2123
R14196 VDD.n4946 VDD.n4945 22.2123
R14197 VDD.n4948 VDD.n4940 22.2123
R14198 VDD.n5231 VDD.n5229 22.2123
R14199 VDD.n5251 VDD.n5250 22.2123
R14200 VDD.n5201 VDD.n5199 22.2123
R14201 VDD.n5212 VDD.n5211 22.2123
R14202 VDD.n5204 VDD.n5203 22.2123
R14203 VDD.n5206 VDD.n5198 22.2123
R14204 VDD.n813 VDD.n812 22.2123
R14205 VDD.n1196 VDD.n1195 22.2123
R14206 VDD.n1804 VDD.t639 20.9587
R14207 VDD.n2012 VDD.t245 20.9587
R14208 VDD.n2383 VDD.t621 20.9587
R14209 VDD.n2641 VDD.t844 20.9587
R14210 VDD.n2899 VDD.t131 20.9587
R14211 VDD.n3157 VDD.t475 20.9587
R14212 VDD.n3415 VDD.t1333 20.9587
R14213 VDD.n5738 VDD.t610 20.9587
R14214 VDD.n5484 VDD.t4 20.9587
R14215 VDD.n3673 VDD.t633 20.9587
R14216 VDD.n3931 VDD.t1383 20.9587
R14217 VDD.n4189 VDD.t885 20.9587
R14218 VDD.n4447 VDD.t123 20.9587
R14219 VDD.n4705 VDD.t74 20.9587
R14220 VDD.n4963 VDD.t785 20.9587
R14221 VDD.n5221 VDD.t1371 20.9587
R14222 VDD.n1507 VDD 20.8224
R14223 VDD.n1457 VDD 20.8224
R14224 VDD.n1707 VDD.n1705 20.5934
R14225 VDD.n2056 VDD.n2054 20.5934
R14226 VDD.n2286 VDD.n2284 20.5934
R14227 VDD.n2544 VDD.n2542 20.5934
R14228 VDD.n2802 VDD.n2800 20.5934
R14229 VDD.n3060 VDD.n3058 20.5934
R14230 VDD.n3318 VDD.n3316 20.5934
R14231 VDD.n5641 VDD.n5639 20.5934
R14232 VDD.n5387 VDD.n5385 20.5934
R14233 VDD.n3576 VDD.n3574 20.5934
R14234 VDD.n3834 VDD.n3832 20.5934
R14235 VDD.n4092 VDD.n4090 20.5934
R14236 VDD.n4350 VDD.n4348 20.5934
R14237 VDD.n4608 VDD.n4606 20.5934
R14238 VDD.n4866 VDD.n4864 20.5934
R14239 VDD.n5124 VDD.n5122 20.5934
R14240 VDD.n13 VDD.n12 19.9534
R14241 VDD.n1157 VDD.n1156 19.9534
R14242 VDD.n1840 VDD.n1839 18.6543
R14243 VDD.n2161 VDD.n2160 18.6543
R14244 VDD.n2419 VDD.n2418 18.6543
R14245 VDD.n2677 VDD.n2676 18.6543
R14246 VDD.n2935 VDD.n2934 18.6543
R14247 VDD.n3193 VDD.n3192 18.6543
R14248 VDD.n3451 VDD.n3450 18.6543
R14249 VDD.n5771 VDD.n5770 18.6543
R14250 VDD.n5517 VDD.n5516 18.6543
R14251 VDD.n3709 VDD.n3708 18.6543
R14252 VDD.n3967 VDD.n3966 18.6543
R14253 VDD.n4225 VDD.n4224 18.6543
R14254 VDD.n4483 VDD.n4482 18.6543
R14255 VDD.n4741 VDD.n4740 18.6543
R14256 VDD.n4999 VDD.n4998 18.6543
R14257 VDD.n5257 VDD.n5256 18.6543
R14258 VDD.n1372 VDD.t669 18.2197
R14259 VDD.n1654 VDD 17.4176
R14260 VDD.n1761 VDD.n1716 17.109
R14261 VDD.n2110 VDD.n2065 17.109
R14262 VDD.n2340 VDD.n2295 17.109
R14263 VDD.n2598 VDD.n2553 17.109
R14264 VDD.n2856 VDD.n2811 17.109
R14265 VDD.n3114 VDD.n3069 17.109
R14266 VDD.n3372 VDD.n3327 17.109
R14267 VDD.n5695 VDD.n5650 17.109
R14268 VDD.n5441 VDD.n5396 17.109
R14269 VDD.n3630 VDD.n3585 17.109
R14270 VDD.n3888 VDD.n3843 17.109
R14271 VDD.n4146 VDD.n4101 17.109
R14272 VDD.n4404 VDD.n4359 17.109
R14273 VDD.n4662 VDD.n4617 17.109
R14274 VDD.n4920 VDD.n4875 17.109
R14275 VDD.n5178 VDD.n5133 17.109
R14276 VDD.n24 VDD.n23 16.9417
R14277 VDD.n575 VDD.n574 16.9417
R14278 VDD.n597 VDD.n596 16.9417
R14279 VDD.n658 VDD.n657 16.9417
R14280 VDD.n768 VDD.n767 16.9417
R14281 VDD.n721 VDD.n720 16.9417
R14282 VDD.n488 VDD.n487 16.9417
R14283 VDD.n86 VDD.n85 16.9417
R14284 VDD.n1168 VDD.n1167 16.9417
R14285 VDD.n925 VDD.n924 16.9417
R14286 VDD.n947 VDD.n946 16.9417
R14287 VDD.n1008 VDD.n1007 16.9417
R14288 VDD.n1118 VDD.n1117 16.9417
R14289 VDD.n1071 VDD.n1070 16.9417
R14290 VDD.n174 VDD.n173 16.9417
R14291 VDD.n196 VDD.n195 16.9417
R14292 VDD.n253 VDD.n252 16.9417
R14293 VDD.n363 VDD.n362 16.9417
R14294 VDD.n316 VDD.n315 16.9417
R14295 VDD.n1436 VDD.n1435 16.9417
R14296 VDD.n1404 VDD.n1403 16.9417
R14297 VDD.n1269 VDD.n1268 16.9417
R14298 VDD.n1484 VDD.n1483 16.9417
R14299 VDD.n1532 VDD.n1531 16.9417
R14300 VDD.n8 VDD.n2 16.1887
R14301 VDD.n1152 VDD.n1146 16.1887
R14302 VDD.n688 VDD.n687 14.5711
R14303 VDD.n1038 VDD.n1037 14.5711
R14304 VDD.n283 VDD.n282 14.5711
R14305 VDD.n1659 VDD 14.551
R14306 VDD.n1686 VDD.t643 14.2962
R14307 VDD.n2035 VDD.t250 14.2962
R14308 VDD.n2265 VDD.t625 14.2962
R14309 VDD.n2523 VDD.t843 14.2962
R14310 VDD.n2781 VDD.t138 14.2962
R14311 VDD.n3039 VDD.t474 14.2962
R14312 VDD.n3297 VDD.t1332 14.2962
R14313 VDD.n5620 VDD.t616 14.2962
R14314 VDD.n5366 VDD.t7 14.2962
R14315 VDD.n3555 VDD.t632 14.2962
R14316 VDD.n3813 VDD.t1387 14.2962
R14317 VDD.n4071 VDD.t889 14.2962
R14318 VDD.n4329 VDD.t130 14.2962
R14319 VDD.n4587 VDD.t77 14.2962
R14320 VDD.n4845 VDD.t784 14.2962
R14321 VDD.n5103 VDD.t1378 14.2962
R14322 VDD.n1666 VDD.t644 14.2955
R14323 VDD.n2015 VDD.t244 14.2955
R14324 VDD.n2245 VDD.t628 14.2955
R14325 VDD.n2503 VDD.t847 14.2955
R14326 VDD.n2761 VDD.t135 14.2955
R14327 VDD.n3019 VDD.t478 14.2955
R14328 VDD.n3277 VDD.t1336 14.2955
R14329 VDD.n5600 VDD.t614 14.2955
R14330 VDD.n5346 VDD.t10 14.2955
R14331 VDD.n3535 VDD.t636 14.2955
R14332 VDD.n3793 VDD.t1390 14.2955
R14333 VDD.n4051 VDD.t892 14.2955
R14334 VDD.n4309 VDD.t127 14.2955
R14335 VDD.n4567 VDD.t73 14.2955
R14336 VDD.n4825 VDD.t788 14.2955
R14337 VDD.n5083 VDD.t1375 14.2955
R14338 VDD.n1749 VDD.t1366 14.2865
R14339 VDD.n2098 VDD.t1494 14.2865
R14340 VDD.n2328 VDD.t223 14.2865
R14341 VDD.n2586 VDD.t62 14.2865
R14342 VDD.n2844 VDD.t596 14.2865
R14343 VDD.n3102 VDD.t42 14.2865
R14344 VDD.n3360 VDD.t732 14.2865
R14345 VDD.n5683 VDD.t165 14.2865
R14346 VDD.n5429 VDD.t523 14.2865
R14347 VDD.n3618 VDD.t195 14.2865
R14348 VDD.n3876 VDD.t178 14.2865
R14349 VDD.n4134 VDD.t98 14.2865
R14350 VDD.n4392 VDD.t498 14.2865
R14351 VDD.n4650 VDD.t588 14.2865
R14352 VDD.n4908 VDD.t580 14.2865
R14353 VDD.n5166 VDD.t858 14.2865
R14354 VDD.n1737 VDD.t1360 14.2864
R14355 VDD.n2086 VDD.t1495 14.2864
R14356 VDD.n2316 VDD.t225 14.2864
R14357 VDD.n2574 VDD.t56 14.2864
R14358 VDD.n2832 VDD.t598 14.2864
R14359 VDD.n3090 VDD.t44 14.2864
R14360 VDD.n3348 VDD.t734 14.2864
R14361 VDD.n5671 VDD.t167 14.2864
R14362 VDD.n5417 VDD.t518 14.2864
R14363 VDD.n3606 VDD.t197 14.2864
R14364 VDD.n3864 VDD.t174 14.2864
R14365 VDD.n4122 VDD.t93 14.2864
R14366 VDD.n4380 VDD.t500 14.2864
R14367 VDD.n4638 VDD.t590 14.2864
R14368 VDD.n4896 VDD.t582 14.2864
R14369 VDD.n5154 VDD.t860 14.2864
R14370 VDD.n1771 VDD.t389 14.2849
R14371 VDD.n1753 VDD.t537 14.2849
R14372 VDD.n2120 VDD.t229 14.2849
R14373 VDD.n2102 VDD.t1179 14.2849
R14374 VDD.n2350 VDD.t182 14.2849
R14375 VDD.n2332 VDD.t1036 14.2849
R14376 VDD.n2608 VDD.t1198 14.2849
R14377 VDD.n2590 VDD.t714 14.2849
R14378 VDD.n2866 VDD.t1488 14.2849
R14379 VDD.n2848 VDD.t543 14.2849
R14380 VDD.n3124 VDD.t648 14.2849
R14381 VDD.n3106 VDD.t654 14.2849
R14382 VDD.n3382 VDD.t31 14.2849
R14383 VDD.n3364 VDD.t190 14.2849
R14384 VDD.n5705 VDD.t871 14.2849
R14385 VDD.n5687 VDD.t1180 14.2849
R14386 VDD.n5451 VDD.t715 14.2849
R14387 VDD.n5433 VDD.t710 14.2849
R14388 VDD.n3640 VDD.t1445 14.2849
R14389 VDD.n3622 VDD.t215 14.2849
R14390 VDD.n3898 VDD.t1028 14.2849
R14391 VDD.n3880 VDD.t1194 14.2849
R14392 VDD.n4156 VDD.t424 14.2849
R14393 VDD.n4138 VDD.t536 14.2849
R14394 VDD.n4414 VDD.t1032 14.2849
R14395 VDD.n4396 VDD.t1449 14.2849
R14396 VDD.n4672 VDD.t1393 14.2849
R14397 VDD.n4654 VDD.t403 14.2849
R14398 VDD.n4930 VDD.t533 14.2849
R14399 VDD.n4912 VDD.t1035 14.2849
R14400 VDD.n5188 VDD.t382 14.2849
R14401 VDD.n5170 VDD.t514 14.2849
R14402 VDD.n1620 VDD.n1619 14.1868
R14403 VDD.n1769 VDD.n1669 14.0805
R14404 VDD.n2118 VDD.n2018 14.0805
R14405 VDD.n2348 VDD.n2248 14.0805
R14406 VDD.n2606 VDD.n2506 14.0805
R14407 VDD.n2864 VDD.n2764 14.0805
R14408 VDD.n3122 VDD.n3022 14.0805
R14409 VDD.n3380 VDD.n3280 14.0805
R14410 VDD.n5703 VDD.n5603 14.0805
R14411 VDD.n5449 VDD.n5349 14.0805
R14412 VDD.n3638 VDD.n3538 14.0805
R14413 VDD.n3896 VDD.n3796 14.0805
R14414 VDD.n4154 VDD.n4054 14.0805
R14415 VDD.n4412 VDD.n4312 14.0805
R14416 VDD.n4670 VDD.n4570 14.0805
R14417 VDD.n4928 VDD.n4828 14.0805
R14418 VDD.n5186 VDD.n5086 14.0805
R14419 VDD.t546 VDD.t386 13.9711
R14420 VDD.t37 VDD.t210 13.9711
R14421 VDD.t230 VDD.t100 13.9711
R14422 VDD.t764 VDD.t876 13.9711
R14423 VDD.n1755 VDD.n1717 13.7605
R14424 VDD.n2104 VDD.n2066 13.7605
R14425 VDD.n2334 VDD.n2296 13.7605
R14426 VDD.n2592 VDD.n2554 13.7605
R14427 VDD.n2850 VDD.n2812 13.7605
R14428 VDD.n3108 VDD.n3070 13.7605
R14429 VDD.n3366 VDD.n3328 13.7605
R14430 VDD.n5689 VDD.n5651 13.7605
R14431 VDD.n5435 VDD.n5397 13.7605
R14432 VDD.n3624 VDD.n3586 13.7605
R14433 VDD.n3882 VDD.n3844 13.7605
R14434 VDD.n4140 VDD.n4102 13.7605
R14435 VDD.n4398 VDD.n4360 13.7605
R14436 VDD.n4656 VDD.n4618 13.7605
R14437 VDD.n4914 VDD.n4876 13.7605
R14438 VDD.n5172 VDD.n5134 13.7605
R14439 VDD.n1658 VDD.n1631 13.4428
R14440 VDD.n1657 VDD 13.4235
R14441 VDD.n807 VDD.n805 13.3488
R14442 VDD.n1190 VDD.n1188 13.3488
R14443 VDD.n827 VDD.n826 12.9329
R14444 VDD.n1543 VDD.n1542 12.9329
R14445 VDD.n1363 VDD.n1362 12.9329
R14446 VDD.n1210 VDD.n1209 12.9329
R14447 VDD.n580 VDD.n579 11.6711
R14448 VDD.n593 VDD.n592 11.6711
R14449 VDD.n663 VDD.n662 11.6711
R14450 VDD.n772 VDD.n771 11.6711
R14451 VDD.n725 VDD.n724 11.6711
R14452 VDD.n930 VDD.n929 11.6711
R14453 VDD.n943 VDD.n942 11.6711
R14454 VDD.n1013 VDD.n1012 11.6711
R14455 VDD.n1122 VDD.n1121 11.6711
R14456 VDD.n1075 VDD.n1074 11.6711
R14457 VDD.n179 VDD.n178 11.6711
R14458 VDD.n192 VDD.n191 11.6711
R14459 VDD.n258 VDD.n257 11.6711
R14460 VDD.n367 VDD.n366 11.6711
R14461 VDD.n320 VDD.n319 11.6711
R14462 VDD.n1440 VDD.n1439 11.6711
R14463 VDD.n1409 VDD.n1408 11.6711
R14464 VDD.n1273 VDD.n1272 11.6711
R14465 VDD.n1488 VDD.n1487 11.6711
R14466 VDD.n1536 VDD.n1535 11.6711
R14467 VDD.n569 VDD.n568 10.9181
R14468 VDD.n603 VDD.n602 10.9181
R14469 VDD.n652 VDD.n651 10.9181
R14470 VDD.n762 VDD.n761 10.9181
R14471 VDD.n715 VDD.n714 10.9181
R14472 VDD.n919 VDD.n918 10.9181
R14473 VDD.n953 VDD.n952 10.9181
R14474 VDD.n1002 VDD.n1001 10.9181
R14475 VDD.n1112 VDD.n1111 10.9181
R14476 VDD.n1065 VDD.n1064 10.9181
R14477 VDD.n168 VDD.n167 10.9181
R14478 VDD.n202 VDD.n201 10.9181
R14479 VDD.n247 VDD.n246 10.9181
R14480 VDD.n357 VDD.n356 10.9181
R14481 VDD.n310 VDD.n309 10.9181
R14482 VDD.n1323 VDD.n1322 10.9181
R14483 VDD.n1392 VDD.n1391 10.9181
R14484 VDD.n1294 VDD.n1293 10.9181
R14485 VDD.n1478 VDD.n1477 10.9181
R14486 VDD.n1258 VDD.n1257 10.9181
R14487 VDD.n1957 VDD.n1956 10.8802
R14488 VDD.n463 VDD 10.8576
R14489 VDD.n60 VDD 10.8576
R14490 VDD.n1955 VDD.n1954 10.5887
R14491 VDD.n1429 VDD.t1289 10.4115
R14492 VDD.n668 VDD.t1133 10.1791
R14493 VDD.n1018 VDD.t1004 10.1791
R14494 VDD.t431 VDD.n264 10.1791
R14495 VDD.n1617 VDD 9.58775
R14496 VDD.n9 VDD.n6 9.41227
R14497 VDD.n1153 VDD.n1150 9.41227
R14498 VDD.n1954 VDD.n1953 9.3005
R14499 VDD.n1916 VDD.n1915 9.3005
R14500 VDD.n1915 VDD.n1914 9.3005
R14501 VDD.n1828 VDD.n1826 9.3005
R14502 VDD.n1747 VDD.n1746 9.3005
R14503 VDD.n1728 VDD.n1727 9.3005
R14504 VDD.n1731 VDD.n1722 9.3005
R14505 VDD.n1705 VDD.n1667 9.3005
R14506 VDD.n1690 VDD.n1689 9.3005
R14507 VDD.n2096 VDD.n2095 9.3005
R14508 VDD.n2077 VDD.n2076 9.3005
R14509 VDD.n2080 VDD.n2071 9.3005
R14510 VDD.n2054 VDD.n2016 9.3005
R14511 VDD.n2039 VDD.n2038 9.3005
R14512 VDD.n2237 VDD.n2236 9.3005
R14513 VDD.n2236 VDD.n2235 9.3005
R14514 VDD.n2149 VDD.n2147 9.3005
R14515 VDD.n2326 VDD.n2325 9.3005
R14516 VDD.n2307 VDD.n2306 9.3005
R14517 VDD.n2310 VDD.n2301 9.3005
R14518 VDD.n2284 VDD.n2246 9.3005
R14519 VDD.n2269 VDD.n2268 9.3005
R14520 VDD.n2495 VDD.n2494 9.3005
R14521 VDD.n2494 VDD.n2493 9.3005
R14522 VDD.n2407 VDD.n2405 9.3005
R14523 VDD.n2584 VDD.n2583 9.3005
R14524 VDD.n2565 VDD.n2564 9.3005
R14525 VDD.n2568 VDD.n2559 9.3005
R14526 VDD.n2542 VDD.n2504 9.3005
R14527 VDD.n2527 VDD.n2526 9.3005
R14528 VDD.n2753 VDD.n2752 9.3005
R14529 VDD.n2752 VDD.n2751 9.3005
R14530 VDD.n2665 VDD.n2663 9.3005
R14531 VDD.n2842 VDD.n2841 9.3005
R14532 VDD.n2823 VDD.n2822 9.3005
R14533 VDD.n2826 VDD.n2817 9.3005
R14534 VDD.n2800 VDD.n2762 9.3005
R14535 VDD.n2785 VDD.n2784 9.3005
R14536 VDD.n3011 VDD.n3010 9.3005
R14537 VDD.n3010 VDD.n3009 9.3005
R14538 VDD.n2923 VDD.n2921 9.3005
R14539 VDD.n3100 VDD.n3099 9.3005
R14540 VDD.n3081 VDD.n3080 9.3005
R14541 VDD.n3084 VDD.n3075 9.3005
R14542 VDD.n3058 VDD.n3020 9.3005
R14543 VDD.n3043 VDD.n3042 9.3005
R14544 VDD.n3269 VDD.n3268 9.3005
R14545 VDD.n3268 VDD.n3267 9.3005
R14546 VDD.n3181 VDD.n3179 9.3005
R14547 VDD.n3358 VDD.n3357 9.3005
R14548 VDD.n3339 VDD.n3338 9.3005
R14549 VDD.n3342 VDD.n3333 9.3005
R14550 VDD.n3316 VDD.n3278 9.3005
R14551 VDD.n3301 VDD.n3300 9.3005
R14552 VDD.n3527 VDD.n3526 9.3005
R14553 VDD.n3526 VDD.n3525 9.3005
R14554 VDD.n3439 VDD.n3437 9.3005
R14555 VDD.n5681 VDD.n5680 9.3005
R14556 VDD.n5662 VDD.n5661 9.3005
R14557 VDD.n5665 VDD.n5656 9.3005
R14558 VDD.n5639 VDD.n5601 9.3005
R14559 VDD.n5624 VDD.n5623 9.3005
R14560 VDD.n5847 VDD.n5846 9.3005
R14561 VDD.n5846 VDD.n5845 9.3005
R14562 VDD.n5759 VDD.n5757 9.3005
R14563 VDD.n5427 VDD.n5426 9.3005
R14564 VDD.n5408 VDD.n5407 9.3005
R14565 VDD.n5411 VDD.n5402 9.3005
R14566 VDD.n5385 VDD.n5347 9.3005
R14567 VDD.n5370 VDD.n5369 9.3005
R14568 VDD.n5593 VDD.n5592 9.3005
R14569 VDD.n5592 VDD.n5591 9.3005
R14570 VDD.n5505 VDD.n5503 9.3005
R14571 VDD.n3616 VDD.n3615 9.3005
R14572 VDD.n3597 VDD.n3596 9.3005
R14573 VDD.n3600 VDD.n3591 9.3005
R14574 VDD.n3574 VDD.n3536 9.3005
R14575 VDD.n3559 VDD.n3558 9.3005
R14576 VDD.n3785 VDD.n3784 9.3005
R14577 VDD.n3784 VDD.n3783 9.3005
R14578 VDD.n3697 VDD.n3695 9.3005
R14579 VDD.n3874 VDD.n3873 9.3005
R14580 VDD.n3855 VDD.n3854 9.3005
R14581 VDD.n3858 VDD.n3849 9.3005
R14582 VDD.n3832 VDD.n3794 9.3005
R14583 VDD.n3817 VDD.n3816 9.3005
R14584 VDD.n4043 VDD.n4042 9.3005
R14585 VDD.n4042 VDD.n4041 9.3005
R14586 VDD.n3955 VDD.n3953 9.3005
R14587 VDD.n4132 VDD.n4131 9.3005
R14588 VDD.n4113 VDD.n4112 9.3005
R14589 VDD.n4116 VDD.n4107 9.3005
R14590 VDD.n4090 VDD.n4052 9.3005
R14591 VDD.n4075 VDD.n4074 9.3005
R14592 VDD.n4301 VDD.n4300 9.3005
R14593 VDD.n4300 VDD.n4299 9.3005
R14594 VDD.n4213 VDD.n4211 9.3005
R14595 VDD.n4390 VDD.n4389 9.3005
R14596 VDD.n4371 VDD.n4370 9.3005
R14597 VDD.n4374 VDD.n4365 9.3005
R14598 VDD.n4348 VDD.n4310 9.3005
R14599 VDD.n4333 VDD.n4332 9.3005
R14600 VDD.n4559 VDD.n4558 9.3005
R14601 VDD.n4558 VDD.n4557 9.3005
R14602 VDD.n4471 VDD.n4469 9.3005
R14603 VDD.n4648 VDD.n4647 9.3005
R14604 VDD.n4629 VDD.n4628 9.3005
R14605 VDD.n4632 VDD.n4623 9.3005
R14606 VDD.n4606 VDD.n4568 9.3005
R14607 VDD.n4591 VDD.n4590 9.3005
R14608 VDD.n4817 VDD.n4816 9.3005
R14609 VDD.n4816 VDD.n4815 9.3005
R14610 VDD.n4729 VDD.n4727 9.3005
R14611 VDD.n4906 VDD.n4905 9.3005
R14612 VDD.n4887 VDD.n4886 9.3005
R14613 VDD.n4890 VDD.n4881 9.3005
R14614 VDD.n4864 VDD.n4826 9.3005
R14615 VDD.n4849 VDD.n4848 9.3005
R14616 VDD.n5075 VDD.n5074 9.3005
R14617 VDD.n5074 VDD.n5073 9.3005
R14618 VDD.n4987 VDD.n4985 9.3005
R14619 VDD.n5164 VDD.n5163 9.3005
R14620 VDD.n5145 VDD.n5144 9.3005
R14621 VDD.n5148 VDD.n5139 9.3005
R14622 VDD.n5122 VDD.n5084 9.3005
R14623 VDD.n5107 VDD.n5106 9.3005
R14624 VDD.n5333 VDD.n5332 9.3005
R14625 VDD.n5332 VDD.n5331 9.3005
R14626 VDD.n5245 VDD.n5243 9.3005
R14627 VDD.n1618 VDD.n1617 9.3005
R14628 VDD VDD.n1628 9.22489
R14629 VDD.n1646 VDD.n1645 9.0245
R14630 VDD.n1734 VDD.n1733 8.88939
R14631 VDD.n2083 VDD.n2082 8.88939
R14632 VDD.n2313 VDD.n2312 8.88939
R14633 VDD.n2571 VDD.n2570 8.88939
R14634 VDD.n2829 VDD.n2828 8.88939
R14635 VDD.n3087 VDD.n3086 8.88939
R14636 VDD.n3345 VDD.n3344 8.88939
R14637 VDD.n5668 VDD.n5667 8.88939
R14638 VDD.n5414 VDD.n5413 8.88939
R14639 VDD.n3603 VDD.n3602 8.88939
R14640 VDD.n3861 VDD.n3860 8.88939
R14641 VDD.n4119 VDD.n4118 8.88939
R14642 VDD.n4377 VDD.n4376 8.88939
R14643 VDD.n4635 VDD.n4634 8.88939
R14644 VDD.n4893 VDD.n4892 8.88939
R14645 VDD.n5151 VDD.n5150 8.88939
R14646 VDD.n1954 VDD.n1943 8.85536
R14647 VDD.n10 VDD.n9 8.79168
R14648 VDD.n413 VDD.n412 8.79168
R14649 VDD.n413 VDD.n411 8.79168
R14650 VDD.n394 VDD.n393 8.79168
R14651 VDD.n1154 VDD.n1153 8.79168
R14652 VDD.n1571 VDD.n1570 8.79168
R14653 VDD.n1571 VDD.n1569 8.79168
R14654 VDD.n1552 VDD.n1551 8.79168
R14655 VDD.n1652 VDD.n1649 8.76429
R14656 VDD.n679 VDD.n671 8.28285
R14657 VDD.n832 VDD.n825 8.28285
R14658 VDD.n838 VDD.n824 8.28285
R14659 VDD.n844 VDD.n823 8.28285
R14660 VDD.n850 VDD.n822 8.28285
R14661 VDD.n1029 VDD.n1021 8.28285
R14662 VDD.n274 VDD.n266 8.28285
R14663 VDD.n1215 VDD.n1208 8.28285
R14664 VDD.n1221 VDD.n1207 8.28285
R14665 VDD.n1227 VDD.n1206 8.28285
R14666 VDD.n1233 VDD.n1205 8.28285
R14667 VDD.n1977 VDD.n1923 7.681
R14668 VDD.n1628 VDD 7.6805
R14669 VDD.n1618 VDD.n1616 7.60183
R14670 VDD.n424 VDD.n423 7.54105
R14671 VDD.n403 VDD.n402 7.54105
R14672 VDD.n1582 VDD.n1581 7.54105
R14673 VDD.n1561 VDD.n1560 7.54105
R14674 VDD.n1885 VDD.n1818 7.49764
R14675 VDD.n2206 VDD.n2139 7.49764
R14676 VDD.n2464 VDD.n2397 7.49764
R14677 VDD.n2722 VDD.n2655 7.49764
R14678 VDD.n2980 VDD.n2913 7.49764
R14679 VDD.n3238 VDD.n3171 7.49764
R14680 VDD.n3496 VDD.n3429 7.49764
R14681 VDD.n5816 VDD.n5749 7.49764
R14682 VDD.n5562 VDD.n5495 7.49764
R14683 VDD.n3754 VDD.n3687 7.49764
R14684 VDD.n4012 VDD.n3945 7.49764
R14685 VDD.n4270 VDD.n4203 7.49764
R14686 VDD.n4528 VDD.n4461 7.49764
R14687 VDD.n4786 VDD.n4719 7.49764
R14688 VDD.n5044 VDD.n4977 7.49764
R14689 VDD.n5302 VDD.n5235 7.49764
R14690 VDD.n1606 VDD.n1605 7.39078
R14691 VDD.n1636 VDD.n1635 7.27155
R14692 VDD.n1917 VDD.t29 7.15136
R14693 VDD.n2238 VDD.t1181 7.15136
R14694 VDD.n2496 VDD.t724 7.15136
R14695 VDD.n2754 VDD.t185 7.15136
R14696 VDD.n3012 VDD.t1026 7.15136
R14697 VDD.n3270 VDD.t235 7.15136
R14698 VDD.n3528 VDD.t1446 7.15136
R14699 VDD.n5848 VDD.t1197 7.15136
R14700 VDD.n5594 VDD.t89 7.15136
R14701 VDD.n3786 VDD.t459 7.15136
R14702 VDD.n4044 VDD.t1443 7.15136
R14703 VDD.n4302 VDD.t728 7.15136
R14704 VDD.n4560 VDD.t884 7.15136
R14705 VDD.n4818 VDD.t1349 7.15136
R14706 VDD.n5076 VDD.t738 7.15136
R14707 VDD.n5334 VDD.t238 7.15136
R14708 VDD.n1872 VDD.t170 7.14897
R14709 VDD.n2193 VDD.t1045 7.14897
R14710 VDD.n2451 VDD.t817 7.14897
R14711 VDD.n2709 VDD.t1191 7.14897
R14712 VDD.n2967 VDD.t408 7.14897
R14713 VDD.n3225 VDD.t829 7.14897
R14714 VDD.n3483 VDD.t539 7.14897
R14715 VDD.n5803 VDD.t893 7.14897
R14716 VDD.n5549 VDD.t187 7.14897
R14717 VDD.n3741 VDD.t1344 7.14897
R14718 VDD.n3999 VDD.t239 7.14897
R14719 VDD.n4257 VDD.t1 7.14897
R14720 VDD.n4515 VDD.t1188 7.14897
R14721 VDD.n4773 VDD.t183 7.14897
R14722 VDD.n5031 VDD.t1046 7.14897
R14723 VDD.n5289 VDD.t525 7.14897
R14724 VDD.n1976 VDD.n1926 7.05932
R14725 VDD.n1625 VDD 6.73734
R14726 VDD.n1833 VDD 6.4005
R14727 VDD.n1812 VDD 6.4005
R14728 VDD.n2133 VDD 6.4005
R14729 VDD.n2154 VDD 6.4005
R14730 VDD.n2391 VDD 6.4005
R14731 VDD.n2412 VDD 6.4005
R14732 VDD.n2649 VDD 6.4005
R14733 VDD.n2670 VDD 6.4005
R14734 VDD.n2907 VDD 6.4005
R14735 VDD.n2928 VDD 6.4005
R14736 VDD.n3165 VDD 6.4005
R14737 VDD.n3186 VDD 6.4005
R14738 VDD.n3423 VDD 6.4005
R14739 VDD.n3444 VDD 6.4005
R14740 VDD.n5743 VDD 6.4005
R14741 VDD.n5764 VDD 6.4005
R14742 VDD.n5489 VDD 6.4005
R14743 VDD.n5510 VDD 6.4005
R14744 VDD.n3681 VDD 6.4005
R14745 VDD.n3702 VDD 6.4005
R14746 VDD.n3939 VDD 6.4005
R14747 VDD.n3960 VDD 6.4005
R14748 VDD.n4197 VDD 6.4005
R14749 VDD.n4218 VDD 6.4005
R14750 VDD.n4455 VDD 6.4005
R14751 VDD.n4476 VDD 6.4005
R14752 VDD.n4713 VDD 6.4005
R14753 VDD.n4734 VDD 6.4005
R14754 VDD.n4971 VDD 6.4005
R14755 VDD.n4992 VDD 6.4005
R14756 VDD.n5229 VDD 6.4005
R14757 VDD.n5250 VDD 6.4005
R14758 VDD.n19 VDD.n18 6.4005
R14759 VDD.n1163 VDD.n1162 6.4005
R14760 VDD.n1646 VDD.n1644 6.23487
R14761 VDD.n1652 VDD 5.65631
R14762 VDD.n1631 VDD 5.65631
R14763 VDD.n536 VDD.n535 5.64756
R14764 VDD.n527 VDD.n526 5.64756
R14765 VDD.n633 VDD.n632 5.64756
R14766 VDD.n779 VDD.n778 5.64756
R14767 VDD.n731 VDD.n730 5.64756
R14768 VDD.n886 VDD.n885 5.64756
R14769 VDD.n877 VDD.n876 5.64756
R14770 VDD.n983 VDD.n982 5.64756
R14771 VDD.n1129 VDD.n1128 5.64756
R14772 VDD.n1081 VDD.n1080 5.64756
R14773 VDD.n135 VDD.n134 5.64756
R14774 VDD.n126 VDD.n125 5.64756
R14775 VDD.n232 VDD.n231 5.64756
R14776 VDD.n374 VDD.n373 5.64756
R14777 VDD.n326 VDD.n325 5.64756
R14778 VDD.n1446 VDD.n1445 5.64756
R14779 VDD.n1415 VDD.n1414 5.64756
R14780 VDD.n1279 VDD.n1278 5.64756
R14781 VDD.n1494 VDD.n1493 5.64756
R14782 VDD.n1254 VDD.n1253 5.64756
R14783 VDD.n2128 VDD.n2013 5.34133
R14784 VDD.n1626 VDD 5.31371
R14785 VDD.n1360 VDD.n1359 5.27114
R14786 VDD.n1505 VDD.n1504 5.27114
R14787 VDD.n1288 VDD.n1287 5.27114
R14788 VDD.n1428 VDD.t691 5.20598
R14789 VDD.n1653 VDD.n1652 4.99699
R14790 VDD.n1648 VDD.n1647 4.98671
R14791 VDD.n563 VDD.n562 4.89462
R14792 VDD.n609 VDD.n608 4.89462
R14793 VDD.n646 VDD.n645 4.89462
R14794 VDD.n756 VDD.n755 4.89462
R14795 VDD.n709 VDD.n708 4.89462
R14796 VDD.n913 VDD.n912 4.89462
R14797 VDD.n959 VDD.n958 4.89462
R14798 VDD.n996 VDD.n995 4.89462
R14799 VDD.n1106 VDD.n1105 4.89462
R14800 VDD.n1059 VDD.n1058 4.89462
R14801 VDD.n162 VDD.n161 4.89462
R14802 VDD.n208 VDD.n207 4.89462
R14803 VDD.n241 VDD.n240 4.89462
R14804 VDD.n351 VDD.n350 4.89462
R14805 VDD.n304 VDD.n303 4.89462
R14806 VDD.n1330 VDD.n1329 4.89462
R14807 VDD.n1386 VDD.n1385 4.89462
R14808 VDD.n1300 VDD.n1299 4.89462
R14809 VDD.n1472 VDD.n1471 4.89462
R14810 VDD.n1522 VDD.n1521 4.89462
R14811 VDD.n1618 VDD 4.8645
R14812 VDD.n1833 VDD.n1832 4.6505
R14813 VDD.n1834 VDD.n1829 4.6505
R14814 VDD.n1812 VDD.n1811 4.6505
R14815 VDD.n1796 VDD.n1781 4.6505
R14816 VDD.n1796 VDD.n1795 4.6505
R14817 VDD.n1791 VDD.n1790 4.6505
R14818 VDD.n1793 VDD.n1791 4.6505
R14819 VDD.n1789 VDD.n1780 4.6505
R14820 VDD.n1787 VDD.n1783 4.6505
R14821 VDD.n1786 VDD.n1785 4.6505
R14822 VDD.n1794 VDD.n1780 4.6505
R14823 VDD.n1783 VDD.n1782 4.6505
R14824 VDD.n1785 VDD.n1784 4.6505
R14825 VDD.n2133 VDD.n2132 4.6505
R14826 VDD.n2154 VDD.n2153 4.6505
R14827 VDD.n2155 VDD.n2150 4.6505
R14828 VDD.n2004 VDD.n1989 4.6505
R14829 VDD.n2004 VDD.n2003 4.6505
R14830 VDD.n1999 VDD.n1998 4.6505
R14831 VDD.n2001 VDD.n1999 4.6505
R14832 VDD.n1997 VDD.n1988 4.6505
R14833 VDD.n1995 VDD.n1991 4.6505
R14834 VDD.n1994 VDD.n1993 4.6505
R14835 VDD.n2002 VDD.n1988 4.6505
R14836 VDD.n1991 VDD.n1990 4.6505
R14837 VDD.n1993 VDD.n1992 4.6505
R14838 VDD.n2391 VDD.n2390 4.6505
R14839 VDD.n2412 VDD.n2411 4.6505
R14840 VDD.n2413 VDD.n2408 4.6505
R14841 VDD.n2375 VDD.n2360 4.6505
R14842 VDD.n2375 VDD.n2374 4.6505
R14843 VDD.n2370 VDD.n2369 4.6505
R14844 VDD.n2372 VDD.n2370 4.6505
R14845 VDD.n2368 VDD.n2359 4.6505
R14846 VDD.n2366 VDD.n2362 4.6505
R14847 VDD.n2365 VDD.n2364 4.6505
R14848 VDD.n2373 VDD.n2359 4.6505
R14849 VDD.n2362 VDD.n2361 4.6505
R14850 VDD.n2364 VDD.n2363 4.6505
R14851 VDD.n2649 VDD.n2648 4.6505
R14852 VDD.n2670 VDD.n2669 4.6505
R14853 VDD.n2671 VDD.n2666 4.6505
R14854 VDD.n2633 VDD.n2618 4.6505
R14855 VDD.n2633 VDD.n2632 4.6505
R14856 VDD.n2628 VDD.n2627 4.6505
R14857 VDD.n2630 VDD.n2628 4.6505
R14858 VDD.n2626 VDD.n2617 4.6505
R14859 VDD.n2624 VDD.n2620 4.6505
R14860 VDD.n2623 VDD.n2622 4.6505
R14861 VDD.n2631 VDD.n2617 4.6505
R14862 VDD.n2620 VDD.n2619 4.6505
R14863 VDD.n2622 VDD.n2621 4.6505
R14864 VDD.n2907 VDD.n2906 4.6505
R14865 VDD.n2928 VDD.n2927 4.6505
R14866 VDD.n2929 VDD.n2924 4.6505
R14867 VDD.n2891 VDD.n2876 4.6505
R14868 VDD.n2891 VDD.n2890 4.6505
R14869 VDD.n2886 VDD.n2885 4.6505
R14870 VDD.n2888 VDD.n2886 4.6505
R14871 VDD.n2884 VDD.n2875 4.6505
R14872 VDD.n2882 VDD.n2878 4.6505
R14873 VDD.n2881 VDD.n2880 4.6505
R14874 VDD.n2889 VDD.n2875 4.6505
R14875 VDD.n2878 VDD.n2877 4.6505
R14876 VDD.n2880 VDD.n2879 4.6505
R14877 VDD.n3165 VDD.n3164 4.6505
R14878 VDD.n3186 VDD.n3185 4.6505
R14879 VDD.n3187 VDD.n3182 4.6505
R14880 VDD.n3149 VDD.n3134 4.6505
R14881 VDD.n3149 VDD.n3148 4.6505
R14882 VDD.n3144 VDD.n3143 4.6505
R14883 VDD.n3146 VDD.n3144 4.6505
R14884 VDD.n3142 VDD.n3133 4.6505
R14885 VDD.n3140 VDD.n3136 4.6505
R14886 VDD.n3139 VDD.n3138 4.6505
R14887 VDD.n3147 VDD.n3133 4.6505
R14888 VDD.n3136 VDD.n3135 4.6505
R14889 VDD.n3138 VDD.n3137 4.6505
R14890 VDD.n3423 VDD.n3422 4.6505
R14891 VDD.n3444 VDD.n3443 4.6505
R14892 VDD.n3445 VDD.n3440 4.6505
R14893 VDD.n3407 VDD.n3392 4.6505
R14894 VDD.n3407 VDD.n3406 4.6505
R14895 VDD.n3402 VDD.n3401 4.6505
R14896 VDD.n3404 VDD.n3402 4.6505
R14897 VDD.n3400 VDD.n3391 4.6505
R14898 VDD.n3398 VDD.n3394 4.6505
R14899 VDD.n3397 VDD.n3396 4.6505
R14900 VDD.n3405 VDD.n3391 4.6505
R14901 VDD.n3394 VDD.n3393 4.6505
R14902 VDD.n3396 VDD.n3395 4.6505
R14903 VDD.n5743 VDD.n5742 4.6505
R14904 VDD.n5764 VDD.n5763 4.6505
R14905 VDD.n5765 VDD.n5760 4.6505
R14906 VDD.n5730 VDD.n5715 4.6505
R14907 VDD.n5730 VDD.n5729 4.6505
R14908 VDD.n5725 VDD.n5724 4.6505
R14909 VDD.n5727 VDD.n5725 4.6505
R14910 VDD.n5723 VDD.n5714 4.6505
R14911 VDD.n5721 VDD.n5717 4.6505
R14912 VDD.n5720 VDD.n5719 4.6505
R14913 VDD.n5728 VDD.n5714 4.6505
R14914 VDD.n5717 VDD.n5716 4.6505
R14915 VDD.n5719 VDD.n5718 4.6505
R14916 VDD.n5489 VDD.n5488 4.6505
R14917 VDD.n5510 VDD.n5509 4.6505
R14918 VDD.n5511 VDD.n5506 4.6505
R14919 VDD.n5476 VDD.n5461 4.6505
R14920 VDD.n5476 VDD.n5475 4.6505
R14921 VDD.n5471 VDD.n5470 4.6505
R14922 VDD.n5473 VDD.n5471 4.6505
R14923 VDD.n5469 VDD.n5460 4.6505
R14924 VDD.n5467 VDD.n5463 4.6505
R14925 VDD.n5466 VDD.n5465 4.6505
R14926 VDD.n5474 VDD.n5460 4.6505
R14927 VDD.n5463 VDD.n5462 4.6505
R14928 VDD.n5465 VDD.n5464 4.6505
R14929 VDD.n3681 VDD.n3680 4.6505
R14930 VDD.n3702 VDD.n3701 4.6505
R14931 VDD.n3703 VDD.n3698 4.6505
R14932 VDD.n3665 VDD.n3650 4.6505
R14933 VDD.n3665 VDD.n3664 4.6505
R14934 VDD.n3660 VDD.n3659 4.6505
R14935 VDD.n3662 VDD.n3660 4.6505
R14936 VDD.n3658 VDD.n3649 4.6505
R14937 VDD.n3656 VDD.n3652 4.6505
R14938 VDD.n3655 VDD.n3654 4.6505
R14939 VDD.n3663 VDD.n3649 4.6505
R14940 VDD.n3652 VDD.n3651 4.6505
R14941 VDD.n3654 VDD.n3653 4.6505
R14942 VDD.n3939 VDD.n3938 4.6505
R14943 VDD.n3960 VDD.n3959 4.6505
R14944 VDD.n3961 VDD.n3956 4.6505
R14945 VDD.n3923 VDD.n3908 4.6505
R14946 VDD.n3923 VDD.n3922 4.6505
R14947 VDD.n3918 VDD.n3917 4.6505
R14948 VDD.n3920 VDD.n3918 4.6505
R14949 VDD.n3916 VDD.n3907 4.6505
R14950 VDD.n3914 VDD.n3910 4.6505
R14951 VDD.n3913 VDD.n3912 4.6505
R14952 VDD.n3921 VDD.n3907 4.6505
R14953 VDD.n3910 VDD.n3909 4.6505
R14954 VDD.n3912 VDD.n3911 4.6505
R14955 VDD.n4197 VDD.n4196 4.6505
R14956 VDD.n4218 VDD.n4217 4.6505
R14957 VDD.n4219 VDD.n4214 4.6505
R14958 VDD.n4181 VDD.n4166 4.6505
R14959 VDD.n4181 VDD.n4180 4.6505
R14960 VDD.n4176 VDD.n4175 4.6505
R14961 VDD.n4178 VDD.n4176 4.6505
R14962 VDD.n4174 VDD.n4165 4.6505
R14963 VDD.n4172 VDD.n4168 4.6505
R14964 VDD.n4171 VDD.n4170 4.6505
R14965 VDD.n4179 VDD.n4165 4.6505
R14966 VDD.n4168 VDD.n4167 4.6505
R14967 VDD.n4170 VDD.n4169 4.6505
R14968 VDD.n4455 VDD.n4454 4.6505
R14969 VDD.n4476 VDD.n4475 4.6505
R14970 VDD.n4477 VDD.n4472 4.6505
R14971 VDD.n4439 VDD.n4424 4.6505
R14972 VDD.n4439 VDD.n4438 4.6505
R14973 VDD.n4434 VDD.n4433 4.6505
R14974 VDD.n4436 VDD.n4434 4.6505
R14975 VDD.n4432 VDD.n4423 4.6505
R14976 VDD.n4430 VDD.n4426 4.6505
R14977 VDD.n4429 VDD.n4428 4.6505
R14978 VDD.n4437 VDD.n4423 4.6505
R14979 VDD.n4426 VDD.n4425 4.6505
R14980 VDD.n4428 VDD.n4427 4.6505
R14981 VDD.n4713 VDD.n4712 4.6505
R14982 VDD.n4734 VDD.n4733 4.6505
R14983 VDD.n4735 VDD.n4730 4.6505
R14984 VDD.n4697 VDD.n4682 4.6505
R14985 VDD.n4697 VDD.n4696 4.6505
R14986 VDD.n4692 VDD.n4691 4.6505
R14987 VDD.n4694 VDD.n4692 4.6505
R14988 VDD.n4690 VDD.n4681 4.6505
R14989 VDD.n4688 VDD.n4684 4.6505
R14990 VDD.n4687 VDD.n4686 4.6505
R14991 VDD.n4695 VDD.n4681 4.6505
R14992 VDD.n4684 VDD.n4683 4.6505
R14993 VDD.n4686 VDD.n4685 4.6505
R14994 VDD.n4971 VDD.n4970 4.6505
R14995 VDD.n4992 VDD.n4991 4.6505
R14996 VDD.n4993 VDD.n4988 4.6505
R14997 VDD.n4955 VDD.n4940 4.6505
R14998 VDD.n4955 VDD.n4954 4.6505
R14999 VDD.n4950 VDD.n4949 4.6505
R15000 VDD.n4952 VDD.n4950 4.6505
R15001 VDD.n4948 VDD.n4939 4.6505
R15002 VDD.n4946 VDD.n4942 4.6505
R15003 VDD.n4945 VDD.n4944 4.6505
R15004 VDD.n4953 VDD.n4939 4.6505
R15005 VDD.n4942 VDD.n4941 4.6505
R15006 VDD.n4944 VDD.n4943 4.6505
R15007 VDD.n5229 VDD.n5228 4.6505
R15008 VDD.n5250 VDD.n5249 4.6505
R15009 VDD.n5251 VDD.n5246 4.6505
R15010 VDD.n5213 VDD.n5198 4.6505
R15011 VDD.n5213 VDD.n5212 4.6505
R15012 VDD.n5208 VDD.n5207 4.6505
R15013 VDD.n5210 VDD.n5208 4.6505
R15014 VDD.n5206 VDD.n5197 4.6505
R15015 VDD.n5204 VDD.n5200 4.6505
R15016 VDD.n5203 VDD.n5202 4.6505
R15017 VDD.n5211 VDD.n5197 4.6505
R15018 VDD.n5200 VDD.n5199 4.6505
R15019 VDD.n5202 VDD.n5201 4.6505
R15020 VDD.n12 VDD.n11 4.6505
R15021 VDD.n14 VDD.n13 4.6505
R15022 VDD.n16 VDD.n8 4.6505
R15023 VDD.n4 VDD.n2 4.6505
R15024 VDD.n23 VDD.n22 4.6505
R15025 VDD.n15 VDD.n6 4.6505
R15026 VDD.n18 VDD.n17 4.6505
R15027 VDD.n21 VDD.n20 4.6505
R15028 VDD.n30 VDD.n29 4.6505
R15029 VDD.n689 VDD.n524 4.6505
R15030 VDD.n697 VDD.n523 4.6505
R15031 VDD.n698 VDD.n522 4.6505
R15032 VDD.n744 VDD.n520 4.6505
R15033 VDD.n745 VDD.n519 4.6505
R15034 VDD.n791 VDD.n517 4.6505
R15035 VDD.n792 VDD.n516 4.6505
R15036 VDD.n622 VDD.n621 4.6505
R15037 VDD.n620 VDD.n619 4.6505
R15038 VDD.n551 VDD.n542 4.6505
R15039 VDD.n552 VDD.n541 4.6505
R15040 VDD.n676 VDD.n675 4.6505
R15041 VDD.n678 VDD.n677 4.6505
R15042 VDD.n680 VDD.n679 4.6505
R15043 VDD.n682 VDD.n681 4.6505
R15044 VDD.n685 VDD.n684 4.6505
R15045 VDD.n691 VDD.n690 4.6505
R15046 VDD.n694 VDD.n693 4.6505
R15047 VDD.n696 VDD.n695 4.6505
R15048 VDD.n700 VDD.n699 4.6505
R15049 VDD.n704 VDD.n703 4.6505
R15050 VDD.n706 VDD.n705 4.6505
R15051 VDD.n710 VDD.n709 4.6505
R15052 VDD.n712 VDD.n711 4.6505
R15053 VDD.n716 VDD.n715 4.6505
R15054 VDD.n718 VDD.n717 4.6505
R15055 VDD.n722 VDD.n721 4.6505
R15056 VDD.n726 VDD.n725 4.6505
R15057 VDD.n728 VDD.n727 4.6505
R15058 VDD.n732 VDD.n731 4.6505
R15059 VDD.n735 VDD.n734 4.6505
R15060 VDD.n740 VDD.n739 4.6505
R15061 VDD.n743 VDD.n742 4.6505
R15062 VDD.n747 VDD.n746 4.6505
R15063 VDD.n751 VDD.n750 4.6505
R15064 VDD.n753 VDD.n752 4.6505
R15065 VDD.n757 VDD.n756 4.6505
R15066 VDD.n759 VDD.n758 4.6505
R15067 VDD.n763 VDD.n762 4.6505
R15068 VDD.n765 VDD.n764 4.6505
R15069 VDD.n769 VDD.n768 4.6505
R15070 VDD.n773 VDD.n772 4.6505
R15071 VDD.n775 VDD.n774 4.6505
R15072 VDD.n780 VDD.n779 4.6505
R15073 VDD.n783 VDD.n782 4.6505
R15074 VDD.n788 VDD.n787 4.6505
R15075 VDD.n790 VDD.n789 4.6505
R15076 VDD.n515 VDD.n514 4.6505
R15077 VDD.n641 VDD.n640 4.6505
R15078 VDD.n643 VDD.n642 4.6505
R15079 VDD.n647 VDD.n646 4.6505
R15080 VDD.n649 VDD.n648 4.6505
R15081 VDD.n653 VDD.n652 4.6505
R15082 VDD.n655 VDD.n654 4.6505
R15083 VDD.n659 VDD.n658 4.6505
R15084 VDD.n664 VDD.n663 4.6505
R15085 VDD.n637 VDD.n636 4.6505
R15086 VDD.n634 VDD.n633 4.6505
R15087 VDD.n630 VDD.n629 4.6505
R15088 VDD.n628 VDD.n627 4.6505
R15089 VDD.n624 VDD.n623 4.6505
R15090 VDD.n618 VDD.n617 4.6505
R15091 VDD.n616 VDD.n615 4.6505
R15092 VDD.n612 VDD.n611 4.6505
R15093 VDD.n610 VDD.n609 4.6505
R15094 VDD.n606 VDD.n605 4.6505
R15095 VDD.n604 VDD.n603 4.6505
R15096 VDD.n600 VDD.n599 4.6505
R15097 VDD.n598 VDD.n597 4.6505
R15098 VDD.n594 VDD.n593 4.6505
R15099 VDD.n589 VDD.n588 4.6505
R15100 VDD.n528 VDD.n527 4.6505
R15101 VDD.n544 VDD.n543 4.6505
R15102 VDD.n548 VDD.n547 4.6505
R15103 VDD.n550 VDD.n549 4.6505
R15104 VDD.n554 VDD.n553 4.6505
R15105 VDD.n558 VDD.n557 4.6505
R15106 VDD.n560 VDD.n559 4.6505
R15107 VDD.n564 VDD.n563 4.6505
R15108 VDD.n566 VDD.n565 4.6505
R15109 VDD.n570 VDD.n569 4.6505
R15110 VDD.n572 VDD.n571 4.6505
R15111 VDD.n576 VDD.n575 4.6505
R15112 VDD.n581 VDD.n580 4.6505
R15113 VDD.n540 VDD.n539 4.6505
R15114 VDD.n537 VDD.n536 4.6505
R15115 VDD.n533 VDD.n532 4.6505
R15116 VDD.n474 VDD.n473 4.6505
R15117 VDD.n480 VDD.n472 4.6505
R15118 VDD.n480 VDD.n470 4.6505
R15119 VDD.n479 VDD.n478 4.6505
R15120 VDD.n485 VDD.n483 4.6505
R15121 VDD.n486 VDD.n469 4.6505
R15122 VDD.n467 VDD.n466 4.6505
R15123 VDD.n491 VDD.n490 4.6505
R15124 VDD.n493 VDD.n492 4.6505
R15125 VDD.n497 VDD.n496 4.6505
R15126 VDD.n499 VDD.n498 4.6505
R15127 VDD.n501 VDD.n500 4.6505
R15128 VDD.n503 VDD.n502 4.6505
R15129 VDD.n505 VDD.n504 4.6505
R15130 VDD.n507 VDD.n506 4.6505
R15131 VDD.n485 VDD.n484 4.6505
R15132 VDD.n487 VDD.n486 4.6505
R15133 VDD.n447 VDD.n446 4.6505
R15134 VDD.n451 VDD.n444 4.6505
R15135 VDD.n450 VDD.n448 4.6505
R15136 VDD.n454 VDD.n452 4.6505
R15137 VDD.n457 VDD.n455 4.6505
R15138 VDD.n447 VDD.n445 4.6505
R15139 VDD.n450 VDD.n449 4.6505
R15140 VDD.n451 VDD.n442 4.6505
R15141 VDD.n454 VDD.n453 4.6505
R15142 VDD.n457 VDD.n456 4.6505
R15143 VDD.n458 VDD.n440 4.6505
R15144 VDD.n415 VDD.n410 4.6505
R15145 VDD.n417 VDD.n409 4.6505
R15146 VDD.n415 VDD.n414 4.6505
R15147 VDD.n417 VDD.n416 4.6505
R15148 VDD.n421 VDD.n420 4.6505
R15149 VDD.n426 VDD.n425 4.6505
R15150 VDD.n428 VDD.n427 4.6505
R15151 VDD.n430 VDD.n429 4.6505
R15152 VDD.n432 VDD.n431 4.6505
R15153 VDD.n434 VDD.n433 4.6505
R15154 VDD.n396 VDD.n392 4.6505
R15155 VDD.n398 VDD.n391 4.6505
R15156 VDD.n398 VDD.n397 4.6505
R15157 VDD.n400 VDD.n399 4.6505
R15158 VDD.n72 VDD.n71 4.6505
R15159 VDD.n78 VDD.n70 4.6505
R15160 VDD.n78 VDD.n68 4.6505
R15161 VDD.n77 VDD.n76 4.6505
R15162 VDD.n83 VDD.n81 4.6505
R15163 VDD.n84 VDD.n67 4.6505
R15164 VDD.n65 VDD.n64 4.6505
R15165 VDD.n89 VDD.n88 4.6505
R15166 VDD.n91 VDD.n90 4.6505
R15167 VDD.n95 VDD.n94 4.6505
R15168 VDD.n97 VDD.n96 4.6505
R15169 VDD.n99 VDD.n98 4.6505
R15170 VDD.n101 VDD.n100 4.6505
R15171 VDD.n103 VDD.n102 4.6505
R15172 VDD.n105 VDD.n104 4.6505
R15173 VDD.n83 VDD.n82 4.6505
R15174 VDD.n85 VDD.n84 4.6505
R15175 VDD.n44 VDD.n43 4.6505
R15176 VDD.n48 VDD.n41 4.6505
R15177 VDD.n47 VDD.n45 4.6505
R15178 VDD.n51 VDD.n49 4.6505
R15179 VDD.n54 VDD.n52 4.6505
R15180 VDD.n44 VDD.n42 4.6505
R15181 VDD.n47 VDD.n46 4.6505
R15182 VDD.n48 VDD.n39 4.6505
R15183 VDD.n51 VDD.n50 4.6505
R15184 VDD.n54 VDD.n53 4.6505
R15185 VDD.n55 VDD.n37 4.6505
R15186 VDD.n1156 VDD.n1155 4.6505
R15187 VDD.n1158 VDD.n1157 4.6505
R15188 VDD.n1160 VDD.n1152 4.6505
R15189 VDD.n1148 VDD.n1146 4.6505
R15190 VDD.n1167 VDD.n1166 4.6505
R15191 VDD.n1159 VDD.n1150 4.6505
R15192 VDD.n1162 VDD.n1161 4.6505
R15193 VDD.n1165 VDD.n1164 4.6505
R15194 VDD.n1174 VDD.n1173 4.6505
R15195 VDD.n1573 VDD.n1568 4.6505
R15196 VDD.n1575 VDD.n1567 4.6505
R15197 VDD.n1573 VDD.n1572 4.6505
R15198 VDD.n1575 VDD.n1574 4.6505
R15199 VDD.n1579 VDD.n1578 4.6505
R15200 VDD.n1584 VDD.n1583 4.6505
R15201 VDD.n1586 VDD.n1585 4.6505
R15202 VDD.n1588 VDD.n1587 4.6505
R15203 VDD.n1590 VDD.n1589 4.6505
R15204 VDD.n1592 VDD.n1591 4.6505
R15205 VDD.n1554 VDD.n1550 4.6505
R15206 VDD.n1556 VDD.n1549 4.6505
R15207 VDD.n1556 VDD.n1555 4.6505
R15208 VDD.n1558 VDD.n1557 4.6505
R15209 VDD.n851 VDD.n850 4.6505
R15210 VDD.n849 VDD.n848 4.6505
R15211 VDD.n847 VDD.n846 4.6505
R15212 VDD.n845 VDD.n844 4.6505
R15213 VDD.n843 VDD.n842 4.6505
R15214 VDD.n841 VDD.n840 4.6505
R15215 VDD.n839 VDD.n838 4.6505
R15216 VDD.n837 VDD.n836 4.6505
R15217 VDD.n835 VDD.n834 4.6505
R15218 VDD.n833 VDD.n832 4.6505
R15219 VDD.n831 VDD.n830 4.6505
R15220 VDD.n829 VDD.n828 4.6505
R15221 VDD.n808 VDD.n804 4.6505
R15222 VDD.n812 VDD.n802 4.6505
R15223 VDD.n818 VDD.n799 4.6505
R15224 VDD.n817 VDD.n816 4.6505
R15225 VDD.n815 VDD.n801 4.6505
R15226 VDD.n814 VDD.n813 4.6505
R15227 VDD.n811 VDD.n810 4.6505
R15228 VDD.n1546 VDD.n1545 4.6505
R15229 VDD.n1039 VDD.n874 4.6505
R15230 VDD.n1047 VDD.n873 4.6505
R15231 VDD.n1048 VDD.n872 4.6505
R15232 VDD.n1094 VDD.n870 4.6505
R15233 VDD.n1095 VDD.n869 4.6505
R15234 VDD.n1141 VDD.n867 4.6505
R15235 VDD.n1142 VDD.n866 4.6505
R15236 VDD.n972 VDD.n971 4.6505
R15237 VDD.n970 VDD.n969 4.6505
R15238 VDD.n901 VDD.n892 4.6505
R15239 VDD.n902 VDD.n891 4.6505
R15240 VDD.n1026 VDD.n1025 4.6505
R15241 VDD.n1028 VDD.n1027 4.6505
R15242 VDD.n1030 VDD.n1029 4.6505
R15243 VDD.n1032 VDD.n1031 4.6505
R15244 VDD.n1035 VDD.n1034 4.6505
R15245 VDD.n1041 VDD.n1040 4.6505
R15246 VDD.n1044 VDD.n1043 4.6505
R15247 VDD.n1046 VDD.n1045 4.6505
R15248 VDD.n1050 VDD.n1049 4.6505
R15249 VDD.n1054 VDD.n1053 4.6505
R15250 VDD.n1056 VDD.n1055 4.6505
R15251 VDD.n1060 VDD.n1059 4.6505
R15252 VDD.n1062 VDD.n1061 4.6505
R15253 VDD.n1066 VDD.n1065 4.6505
R15254 VDD.n1068 VDD.n1067 4.6505
R15255 VDD.n1072 VDD.n1071 4.6505
R15256 VDD.n1076 VDD.n1075 4.6505
R15257 VDD.n1078 VDD.n1077 4.6505
R15258 VDD.n1082 VDD.n1081 4.6505
R15259 VDD.n1085 VDD.n1084 4.6505
R15260 VDD.n1090 VDD.n1089 4.6505
R15261 VDD.n1093 VDD.n1092 4.6505
R15262 VDD.n1097 VDD.n1096 4.6505
R15263 VDD.n1101 VDD.n1100 4.6505
R15264 VDD.n1103 VDD.n1102 4.6505
R15265 VDD.n1107 VDD.n1106 4.6505
R15266 VDD.n1109 VDD.n1108 4.6505
R15267 VDD.n1113 VDD.n1112 4.6505
R15268 VDD.n1115 VDD.n1114 4.6505
R15269 VDD.n1119 VDD.n1118 4.6505
R15270 VDD.n1123 VDD.n1122 4.6505
R15271 VDD.n1125 VDD.n1124 4.6505
R15272 VDD.n1130 VDD.n1129 4.6505
R15273 VDD.n1133 VDD.n1132 4.6505
R15274 VDD.n1138 VDD.n1137 4.6505
R15275 VDD.n1140 VDD.n1139 4.6505
R15276 VDD.n865 VDD.n864 4.6505
R15277 VDD.n991 VDD.n990 4.6505
R15278 VDD.n993 VDD.n992 4.6505
R15279 VDD.n997 VDD.n996 4.6505
R15280 VDD.n999 VDD.n998 4.6505
R15281 VDD.n1003 VDD.n1002 4.6505
R15282 VDD.n1005 VDD.n1004 4.6505
R15283 VDD.n1009 VDD.n1008 4.6505
R15284 VDD.n1014 VDD.n1013 4.6505
R15285 VDD.n987 VDD.n986 4.6505
R15286 VDD.n984 VDD.n983 4.6505
R15287 VDD.n980 VDD.n979 4.6505
R15288 VDD.n978 VDD.n977 4.6505
R15289 VDD.n974 VDD.n973 4.6505
R15290 VDD.n968 VDD.n967 4.6505
R15291 VDD.n966 VDD.n965 4.6505
R15292 VDD.n962 VDD.n961 4.6505
R15293 VDD.n960 VDD.n959 4.6505
R15294 VDD.n956 VDD.n955 4.6505
R15295 VDD.n954 VDD.n953 4.6505
R15296 VDD.n950 VDD.n949 4.6505
R15297 VDD.n948 VDD.n947 4.6505
R15298 VDD.n944 VDD.n943 4.6505
R15299 VDD.n939 VDD.n938 4.6505
R15300 VDD.n878 VDD.n877 4.6505
R15301 VDD.n894 VDD.n893 4.6505
R15302 VDD.n898 VDD.n897 4.6505
R15303 VDD.n900 VDD.n899 4.6505
R15304 VDD.n904 VDD.n903 4.6505
R15305 VDD.n908 VDD.n907 4.6505
R15306 VDD.n910 VDD.n909 4.6505
R15307 VDD.n914 VDD.n913 4.6505
R15308 VDD.n916 VDD.n915 4.6505
R15309 VDD.n920 VDD.n919 4.6505
R15310 VDD.n922 VDD.n921 4.6505
R15311 VDD.n926 VDD.n925 4.6505
R15312 VDD.n931 VDD.n930 4.6505
R15313 VDD.n890 VDD.n889 4.6505
R15314 VDD.n887 VDD.n886 4.6505
R15315 VDD.n883 VDD.n882 4.6505
R15316 VDD.n284 VDD.n123 4.6505
R15317 VDD.n292 VDD.n122 4.6505
R15318 VDD.n293 VDD.n121 4.6505
R15319 VDD.n339 VDD.n119 4.6505
R15320 VDD.n340 VDD.n118 4.6505
R15321 VDD.n386 VDD.n116 4.6505
R15322 VDD.n387 VDD.n115 4.6505
R15323 VDD.n221 VDD.n220 4.6505
R15324 VDD.n219 VDD.n218 4.6505
R15325 VDD.n150 VDD.n141 4.6505
R15326 VDD.n151 VDD.n140 4.6505
R15327 VDD.n271 VDD.n270 4.6505
R15328 VDD.n273 VDD.n272 4.6505
R15329 VDD.n275 VDD.n274 4.6505
R15330 VDD.n277 VDD.n276 4.6505
R15331 VDD.n280 VDD.n279 4.6505
R15332 VDD.n286 VDD.n285 4.6505
R15333 VDD.n289 VDD.n288 4.6505
R15334 VDD.n291 VDD.n290 4.6505
R15335 VDD.n295 VDD.n294 4.6505
R15336 VDD.n299 VDD.n298 4.6505
R15337 VDD.n301 VDD.n300 4.6505
R15338 VDD.n305 VDD.n304 4.6505
R15339 VDD.n307 VDD.n306 4.6505
R15340 VDD.n311 VDD.n310 4.6505
R15341 VDD.n313 VDD.n312 4.6505
R15342 VDD.n317 VDD.n316 4.6505
R15343 VDD.n321 VDD.n320 4.6505
R15344 VDD.n323 VDD.n322 4.6505
R15345 VDD.n327 VDD.n326 4.6505
R15346 VDD.n330 VDD.n329 4.6505
R15347 VDD.n335 VDD.n334 4.6505
R15348 VDD.n338 VDD.n337 4.6505
R15349 VDD.n342 VDD.n341 4.6505
R15350 VDD.n346 VDD.n345 4.6505
R15351 VDD.n348 VDD.n347 4.6505
R15352 VDD.n352 VDD.n351 4.6505
R15353 VDD.n354 VDD.n353 4.6505
R15354 VDD.n358 VDD.n357 4.6505
R15355 VDD.n360 VDD.n359 4.6505
R15356 VDD.n364 VDD.n363 4.6505
R15357 VDD.n368 VDD.n367 4.6505
R15358 VDD.n370 VDD.n369 4.6505
R15359 VDD.n375 VDD.n374 4.6505
R15360 VDD.n378 VDD.n377 4.6505
R15361 VDD.n383 VDD.n382 4.6505
R15362 VDD.n385 VDD.n384 4.6505
R15363 VDD.n389 VDD.n388 4.6505
R15364 VDD.n114 VDD.n113 4.6505
R15365 VDD.n238 VDD.n237 4.6505
R15366 VDD.n242 VDD.n241 4.6505
R15367 VDD.n244 VDD.n243 4.6505
R15368 VDD.n248 VDD.n247 4.6505
R15369 VDD.n250 VDD.n249 4.6505
R15370 VDD.n254 VDD.n253 4.6505
R15371 VDD.n259 VDD.n258 4.6505
R15372 VDD.n236 VDD.n235 4.6505
R15373 VDD.n233 VDD.n232 4.6505
R15374 VDD.n229 VDD.n228 4.6505
R15375 VDD.n227 VDD.n226 4.6505
R15376 VDD.n223 VDD.n222 4.6505
R15377 VDD.n217 VDD.n216 4.6505
R15378 VDD.n215 VDD.n214 4.6505
R15379 VDD.n211 VDD.n210 4.6505
R15380 VDD.n209 VDD.n208 4.6505
R15381 VDD.n205 VDD.n204 4.6505
R15382 VDD.n203 VDD.n202 4.6505
R15383 VDD.n199 VDD.n198 4.6505
R15384 VDD.n197 VDD.n196 4.6505
R15385 VDD.n193 VDD.n192 4.6505
R15386 VDD.n188 VDD.n187 4.6505
R15387 VDD.n127 VDD.n126 4.6505
R15388 VDD.n143 VDD.n142 4.6505
R15389 VDD.n147 VDD.n146 4.6505
R15390 VDD.n149 VDD.n148 4.6505
R15391 VDD.n153 VDD.n152 4.6505
R15392 VDD.n157 VDD.n156 4.6505
R15393 VDD.n159 VDD.n158 4.6505
R15394 VDD.n163 VDD.n162 4.6505
R15395 VDD.n165 VDD.n164 4.6505
R15396 VDD.n169 VDD.n168 4.6505
R15397 VDD.n171 VDD.n170 4.6505
R15398 VDD.n175 VDD.n174 4.6505
R15399 VDD.n180 VDD.n179 4.6505
R15400 VDD.n139 VDD.n138 4.6505
R15401 VDD.n136 VDD.n135 4.6505
R15402 VDD.n132 VDD.n131 4.6505
R15403 VDD.n1358 VDD.n1357 4.6505
R15404 VDD.n1349 VDD.n1348 4.6505
R15405 VDD.n1347 VDD.n1346 4.6505
R15406 VDD.n1343 VDD.n1342 4.6505
R15407 VDD.n1341 VDD.n1340 4.6505
R15408 VDD.n1314 VDD.n1313 4.6505
R15409 VDD.n1365 VDD.n1364 4.6505
R15410 VDD.n1368 VDD.n1367 4.6505
R15411 VDD.n1356 VDD.n1355 4.6505
R15412 VDD.n1354 VDD.n1353 4.6505
R15413 VDD.n1351 VDD.n1350 4.6505
R15414 VDD.n1376 VDD.n1375 4.6505
R15415 VDD.n1381 VDD.n1380 4.6505
R15416 VDD.n1383 VDD.n1382 4.6505
R15417 VDD.n1387 VDD.n1386 4.6505
R15418 VDD.n1389 VDD.n1388 4.6505
R15419 VDD.n1393 VDD.n1392 4.6505
R15420 VDD.n1396 VDD.n1395 4.6505
R15421 VDD.n1405 VDD.n1404 4.6505
R15422 VDD.n1410 VDD.n1409 4.6505
R15423 VDD.n1412 VDD.n1411 4.6505
R15424 VDD.n1416 VDD.n1415 4.6505
R15425 VDD.n1418 VDD.n1417 4.6505
R15426 VDD.n1422 VDD.n1421 4.6505
R15427 VDD.n1425 VDD.n1424 4.6505
R15428 VDD.n1339 VDD.n1338 4.6505
R15429 VDD.n1337 VDD.n1336 4.6505
R15430 VDD.n1333 VDD.n1332 4.6505
R15431 VDD.n1331 VDD.n1330 4.6505
R15432 VDD.n1327 VDD.n1326 4.6505
R15433 VDD.n1324 VDD.n1323 4.6505
R15434 VDD.n1433 VDD.n1432 4.6505
R15435 VDD.n1437 VDD.n1436 4.6505
R15436 VDD.n1441 VDD.n1440 4.6505
R15437 VDD.n1443 VDD.n1442 4.6505
R15438 VDD.n1447 VDD.n1446 4.6505
R15439 VDD.n1449 VDD.n1448 4.6505
R15440 VDD.n1453 VDD.n1452 4.6505
R15441 VDD.n1317 VDD.n1316 4.6505
R15442 VDD.n1312 VDD.n1311 4.6505
R15443 VDD.n1310 VDD.n1309 4.6505
R15444 VDD.n1308 VDD.n1307 4.6505
R15445 VDD.n1527 VDD.n1258 4.6505
R15446 VDD.n1529 VDD.n1528 4.6505
R15447 VDD.n1533 VDD.n1532 4.6505
R15448 VDD.n1537 VDD.n1536 4.6505
R15449 VDD.n1539 VDD.n1538 4.6505
R15450 VDD.n1255 VDD.n1254 4.6505
R15451 VDD.n1251 VDD.n1250 4.6505
R15452 VDD.n1286 VDD.n1263 4.6505
R15453 VDD.n1460 VDD.n1262 4.6505
R15454 VDD.n1261 VDD.n1260 4.6505
R15455 VDD.n1510 VDD.n1259 4.6505
R15456 VDD.n1283 VDD.n1266 4.6505
R15457 VDD.n1285 VDD.n1284 4.6505
R15458 VDD.n1463 VDD.n1462 4.6505
R15459 VDD.n1467 VDD.n1466 4.6505
R15460 VDD.n1469 VDD.n1468 4.6505
R15461 VDD.n1473 VDD.n1472 4.6505
R15462 VDD.n1475 VDD.n1474 4.6505
R15463 VDD.n1479 VDD.n1478 4.6505
R15464 VDD.n1481 VDD.n1480 4.6505
R15465 VDD.n1485 VDD.n1484 4.6505
R15466 VDD.n1489 VDD.n1488 4.6505
R15467 VDD.n1491 VDD.n1490 4.6505
R15468 VDD.n1495 VDD.n1494 4.6505
R15469 VDD.n1497 VDD.n1496 4.6505
R15470 VDD.n1501 VDD.n1500 4.6505
R15471 VDD.n1503 VDD.n1502 4.6505
R15472 VDD.n1513 VDD.n1512 4.6505
R15473 VDD.n1517 VDD.n1516 4.6505
R15474 VDD.n1519 VDD.n1518 4.6505
R15475 VDD.n1523 VDD.n1522 4.6505
R15476 VDD.n1525 VDD.n1524 4.6505
R15477 VDD.n1303 VDD.n1302 4.6505
R15478 VDD.n1301 VDD.n1300 4.6505
R15479 VDD.n1297 VDD.n1296 4.6505
R15480 VDD.n1295 VDD.n1294 4.6505
R15481 VDD.n1291 VDD.n1290 4.6505
R15482 VDD.n1270 VDD.n1269 4.6505
R15483 VDD.n1274 VDD.n1273 4.6505
R15484 VDD.n1276 VDD.n1275 4.6505
R15485 VDD.n1280 VDD.n1279 4.6505
R15486 VDD.n1282 VDD.n1281 4.6505
R15487 VDD.n1234 VDD.n1233 4.6505
R15488 VDD.n1232 VDD.n1231 4.6505
R15489 VDD.n1230 VDD.n1229 4.6505
R15490 VDD.n1228 VDD.n1227 4.6505
R15491 VDD.n1226 VDD.n1225 4.6505
R15492 VDD.n1224 VDD.n1223 4.6505
R15493 VDD.n1222 VDD.n1221 4.6505
R15494 VDD.n1220 VDD.n1219 4.6505
R15495 VDD.n1218 VDD.n1217 4.6505
R15496 VDD.n1216 VDD.n1215 4.6505
R15497 VDD.n1214 VDD.n1213 4.6505
R15498 VDD.n1212 VDD.n1211 4.6505
R15499 VDD.n1191 VDD.n1187 4.6505
R15500 VDD.n1195 VDD.n1185 4.6505
R15501 VDD.n1201 VDD.n1182 4.6505
R15502 VDD.n1200 VDD.n1199 4.6505
R15503 VDD.n1198 VDD.n1184 4.6505
R15504 VDD.n1197 VDD.n1196 4.6505
R15505 VDD.n1194 VDD.n1193 4.6505
R15506 VDD.n1653 VDD.n1646 4.61128
R15507 VDD.n1946 VDD.n1943 4.58799
R15508 VDD.n1751 VDD.n1721 4.5005
R15509 VDD.n1751 VDD.n1716 4.5005
R15510 VDD.n1751 VDD.n1750 4.5005
R15511 VDD.n1777 VDD.n1776 4.5005
R15512 VDD.n1800 VDD.n1779 4.5005
R15513 VDD.n1800 VDD.n1799 4.5005
R15514 VDD.n1797 VDD.n1779 4.5005
R15515 VDD.n2100 VDD.n2070 4.5005
R15516 VDD.n2100 VDD.n2065 4.5005
R15517 VDD.n2100 VDD.n2099 4.5005
R15518 VDD.n1985 VDD.n1984 4.5005
R15519 VDD.n2008 VDD.n1987 4.5005
R15520 VDD.n2008 VDD.n2007 4.5005
R15521 VDD.n2005 VDD.n1987 4.5005
R15522 VDD.n2330 VDD.n2300 4.5005
R15523 VDD.n2330 VDD.n2295 4.5005
R15524 VDD.n2330 VDD.n2329 4.5005
R15525 VDD.n2356 VDD.n2355 4.5005
R15526 VDD.n2379 VDD.n2358 4.5005
R15527 VDD.n2379 VDD.n2378 4.5005
R15528 VDD.n2376 VDD.n2358 4.5005
R15529 VDD.n2588 VDD.n2558 4.5005
R15530 VDD.n2588 VDD.n2553 4.5005
R15531 VDD.n2588 VDD.n2587 4.5005
R15532 VDD.n2614 VDD.n2613 4.5005
R15533 VDD.n2637 VDD.n2616 4.5005
R15534 VDD.n2637 VDD.n2636 4.5005
R15535 VDD.n2634 VDD.n2616 4.5005
R15536 VDD.n2846 VDD.n2816 4.5005
R15537 VDD.n2846 VDD.n2811 4.5005
R15538 VDD.n2846 VDD.n2845 4.5005
R15539 VDD.n2872 VDD.n2871 4.5005
R15540 VDD.n2895 VDD.n2874 4.5005
R15541 VDD.n2895 VDD.n2894 4.5005
R15542 VDD.n2892 VDD.n2874 4.5005
R15543 VDD.n3104 VDD.n3074 4.5005
R15544 VDD.n3104 VDD.n3069 4.5005
R15545 VDD.n3104 VDD.n3103 4.5005
R15546 VDD.n3130 VDD.n3129 4.5005
R15547 VDD.n3153 VDD.n3132 4.5005
R15548 VDD.n3153 VDD.n3152 4.5005
R15549 VDD.n3150 VDD.n3132 4.5005
R15550 VDD.n3362 VDD.n3332 4.5005
R15551 VDD.n3362 VDD.n3327 4.5005
R15552 VDD.n3362 VDD.n3361 4.5005
R15553 VDD.n3388 VDD.n3387 4.5005
R15554 VDD.n3411 VDD.n3390 4.5005
R15555 VDD.n3411 VDD.n3410 4.5005
R15556 VDD.n3408 VDD.n3390 4.5005
R15557 VDD.n5685 VDD.n5655 4.5005
R15558 VDD.n5685 VDD.n5650 4.5005
R15559 VDD.n5685 VDD.n5684 4.5005
R15560 VDD.n5711 VDD.n5710 4.5005
R15561 VDD.n5734 VDD.n5713 4.5005
R15562 VDD.n5734 VDD.n5733 4.5005
R15563 VDD.n5731 VDD.n5713 4.5005
R15564 VDD.n5431 VDD.n5401 4.5005
R15565 VDD.n5431 VDD.n5396 4.5005
R15566 VDD.n5431 VDD.n5430 4.5005
R15567 VDD.n5457 VDD.n5456 4.5005
R15568 VDD.n5480 VDD.n5459 4.5005
R15569 VDD.n5480 VDD.n5479 4.5005
R15570 VDD.n5477 VDD.n5459 4.5005
R15571 VDD.n3620 VDD.n3590 4.5005
R15572 VDD.n3620 VDD.n3585 4.5005
R15573 VDD.n3620 VDD.n3619 4.5005
R15574 VDD.n3646 VDD.n3645 4.5005
R15575 VDD.n3669 VDD.n3648 4.5005
R15576 VDD.n3669 VDD.n3668 4.5005
R15577 VDD.n3666 VDD.n3648 4.5005
R15578 VDD.n3878 VDD.n3848 4.5005
R15579 VDD.n3878 VDD.n3843 4.5005
R15580 VDD.n3878 VDD.n3877 4.5005
R15581 VDD.n3904 VDD.n3903 4.5005
R15582 VDD.n3927 VDD.n3906 4.5005
R15583 VDD.n3927 VDD.n3926 4.5005
R15584 VDD.n3924 VDD.n3906 4.5005
R15585 VDD.n4136 VDD.n4106 4.5005
R15586 VDD.n4136 VDD.n4101 4.5005
R15587 VDD.n4136 VDD.n4135 4.5005
R15588 VDD.n4162 VDD.n4161 4.5005
R15589 VDD.n4185 VDD.n4164 4.5005
R15590 VDD.n4185 VDD.n4184 4.5005
R15591 VDD.n4182 VDD.n4164 4.5005
R15592 VDD.n4394 VDD.n4364 4.5005
R15593 VDD.n4394 VDD.n4359 4.5005
R15594 VDD.n4394 VDD.n4393 4.5005
R15595 VDD.n4420 VDD.n4419 4.5005
R15596 VDD.n4443 VDD.n4422 4.5005
R15597 VDD.n4443 VDD.n4442 4.5005
R15598 VDD.n4440 VDD.n4422 4.5005
R15599 VDD.n4652 VDD.n4622 4.5005
R15600 VDD.n4652 VDD.n4617 4.5005
R15601 VDD.n4652 VDD.n4651 4.5005
R15602 VDD.n4678 VDD.n4677 4.5005
R15603 VDD.n4701 VDD.n4680 4.5005
R15604 VDD.n4701 VDD.n4700 4.5005
R15605 VDD.n4698 VDD.n4680 4.5005
R15606 VDD.n4910 VDD.n4880 4.5005
R15607 VDD.n4910 VDD.n4875 4.5005
R15608 VDD.n4910 VDD.n4909 4.5005
R15609 VDD.n4936 VDD.n4935 4.5005
R15610 VDD.n4959 VDD.n4938 4.5005
R15611 VDD.n4959 VDD.n4958 4.5005
R15612 VDD.n4956 VDD.n4938 4.5005
R15613 VDD.n5168 VDD.n5138 4.5005
R15614 VDD.n5168 VDD.n5133 4.5005
R15615 VDD.n5168 VDD.n5167 4.5005
R15616 VDD.n5194 VDD.n5193 4.5005
R15617 VDD.n5217 VDD.n5196 4.5005
R15618 VDD.n5217 VDD.n5216 4.5005
R15619 VDD.n5214 VDD.n5196 4.5005
R15620 VDD.n1249 VDD.n1248 4.45149
R15621 VDD.n531 VDD.n530 4.4514
R15622 VDD.n881 VDD.n880 4.4514
R15623 VDD.n130 VDD.n129 4.4514
R15624 VDD.n1649 VDD.n1648 4.43268
R15625 VDD.n1887 VDD.t472 4.35136
R15626 VDD.n1874 VDD.t102 4.35136
R15627 VDD.n2195 VDD.t721 4.35136
R15628 VDD.n2208 VDD.t743 4.35136
R15629 VDD.n2453 VDD.t649 4.35136
R15630 VDD.n2466 VDD.t650 4.35136
R15631 VDD.n2711 VDD.t111 4.35136
R15632 VDD.n2724 VDD.t83 4.35136
R15633 VDD.n2969 VDD.t107 4.35136
R15634 VDD.n2982 VDD.t470 4.35136
R15635 VDD.n3227 VDD.t720 4.35136
R15636 VDD.n3240 VDD.t1352 4.35136
R15637 VDD.n3485 VDD.t486 4.35136
R15638 VDD.n3498 VDD.t487 4.35136
R15639 VDD.n5805 VDD.t112 4.35136
R15640 VDD.n5818 VDD.t113 4.35136
R15641 VDD.n5551 VDD.t16 4.35136
R15642 VDD.n5564 VDD.t17 4.35136
R15643 VDD.n3743 VDD.t744 4.35136
R15644 VDD.n3756 VDD.t745 4.35136
R15645 VDD.n4001 VDD.t1354 4.35136
R15646 VDD.n4014 VDD.t653 4.35136
R15647 VDD.n4259 VDD.t80 4.35136
R15648 VDD.n4272 VDD.t81 4.35136
R15649 VDD.n4517 VDD.t104 4.35136
R15650 VDD.n4530 VDD.t105 4.35136
R15651 VDD.n4775 VDD.t1350 4.35136
R15652 VDD.n4788 VDD.t1351 4.35136
R15653 VDD.n5033 VDD.t120 4.35136
R15654 VDD.n5046 VDD.t121 4.35136
R15655 VDD.n5291 VDD.t110 4.35136
R15656 VDD.n5304 VDD.t483 4.35136
R15657 VDD.n1633 VDD 4.26717
R15658 VDD.n674 VDD.n673 4.14756
R15659 VDD.n1024 VDD.n1023 4.14756
R15660 VDD.n269 VDD.n268 4.14756
R15661 VDD.n466 VDD.n465 4.14168
R15662 VDD.n64 VDD.n63 4.14168
R15663 VDD.n805 VDD.n804 4.14168
R15664 VDD.n1188 VDD.n1187 4.14168
R15665 VDD.n489 VDD.n488 4.05611
R15666 VDD.n87 VDD.n86 4.05611
R15667 VDD.n25 VDD.n24 4.05569
R15668 VDD.n461 VDD.n460 4.05569
R15669 VDD.n58 VDD.n57 4.05569
R15670 VDD.n1169 VDD.n1168 4.05569
R15671 VDD.n1626 VDD.n1625 4.04261
R15672 VDD.n510 VDD.n509 4.01726
R15673 VDD.n437 VDD.n436 4.01726
R15674 VDD.n406 VDD.n405 4.01726
R15675 VDD.n108 VDD.n107 4.01726
R15676 VDD.n1595 VDD.n1594 4.01726
R15677 VDD.n1564 VDD.n1563 4.01726
R15678 VDD.n33 VDD.n32 4.01682
R15679 VDD.n1177 VDD.n1176 4.01682
R15680 VDD.n1815 VDD.n1814 3.96837
R15681 VDD.n2136 VDD.n2135 3.96837
R15682 VDD.n2394 VDD.n2393 3.96837
R15683 VDD.n2652 VDD.n2651 3.96837
R15684 VDD.n2910 VDD.n2909 3.96837
R15685 VDD.n3168 VDD.n3167 3.96837
R15686 VDD.n3426 VDD.n3425 3.96837
R15687 VDD.n5746 VDD.n5745 3.96837
R15688 VDD.n5492 VDD.n5491 3.96837
R15689 VDD.n3684 VDD.n3683 3.96837
R15690 VDD.n3942 VDD.n3941 3.96837
R15691 VDD.n4200 VDD.n4199 3.96837
R15692 VDD.n4458 VDD.n4457 3.96837
R15693 VDD.n4716 VDD.n4715 3.96837
R15694 VDD.n4974 VDD.n4973 3.96837
R15695 VDD.n5232 VDD.n5231 3.96837
R15696 VDD.n820 VDD.n819 3.96556
R15697 VDD.n1203 VDD.n1202 3.96556
R15698 VDD.n1638 VDD.n1637 3.88621
R15699 VDD.n1952 VDD.n1939 3.5871
R15700 VDD.n1694 VDD.n1683 3.52991
R15701 VDD.n2043 VDD.n2032 3.52991
R15702 VDD.n2273 VDD.n2262 3.52991
R15703 VDD.n2531 VDD.n2520 3.52991
R15704 VDD.n2789 VDD.n2778 3.52991
R15705 VDD.n3047 VDD.n3036 3.52991
R15706 VDD.n3305 VDD.n3294 3.52991
R15707 VDD.n5628 VDD.n5617 3.52991
R15708 VDD.n5374 VDD.n5363 3.52991
R15709 VDD.n3563 VDD.n3552 3.52991
R15710 VDD.n3821 VDD.n3810 3.52991
R15711 VDD.n4079 VDD.n4068 3.52991
R15712 VDD.n4337 VDD.n4326 3.52991
R15713 VDD.n4595 VDD.n4584 3.52991
R15714 VDD.n4853 VDD.n4842 3.52991
R15715 VDD.n5111 VDD.n5100 3.52991
R15716 VDD.n1608 VDD.n1607 3.46717
R15717 VDD.t1456 VDD.n669 3.39336
R15718 VDD.t1410 VDD.n1019 3.39336
R15719 VDD.n263 VDD.t327 3.39336
R15720 VDD.n20 VDD.n19 3.38874
R15721 VDD.n496 VDD.n495 3.38874
R15722 VDD.n420 VDD.n419 3.38874
R15723 VDD.n94 VDD.n93 3.38874
R15724 VDD.n1164 VDD.n1163 3.38874
R15725 VDD.n1578 VDD.n1577 3.38874
R15726 VDD.n1980 VDD.n1922 3.1102
R15727 VDD.n1980 VDD.n1979 3.08146
R15728 VDD.n1701 VDD.n1700 3.03311
R15729 VDD.n2050 VDD.n2049 3.03311
R15730 VDD.n2280 VDD.n2279 3.03311
R15731 VDD.n2538 VDD.n2537 3.03311
R15732 VDD.n2796 VDD.n2795 3.03311
R15733 VDD.n3054 VDD.n3053 3.03311
R15734 VDD.n3312 VDD.n3311 3.03311
R15735 VDD.n5635 VDD.n5634 3.03311
R15736 VDD.n5381 VDD.n5380 3.03311
R15737 VDD.n3570 VDD.n3569 3.03311
R15738 VDD.n3828 VDD.n3827 3.03311
R15739 VDD.n4086 VDD.n4085 3.03311
R15740 VDD.n4344 VDD.n4343 3.03311
R15741 VDD.n4602 VDD.n4601 3.03311
R15742 VDD.n4860 VDD.n4859 3.03311
R15743 VDD.n5118 VDD.n5117 3.03311
R15744 VDD.n1609 VDD.n1608 3.03311
R15745 VDD VDD.n1622 3.02091
R15746 VDD.n1831 VDD 3.0005
R15747 VDD.n2152 VDD 3.0005
R15748 VDD.n2410 VDD 3.0005
R15749 VDD.n2668 VDD 3.0005
R15750 VDD.n2926 VDD 3.0005
R15751 VDD.n3184 VDD 3.0005
R15752 VDD.n3442 VDD 3.0005
R15753 VDD.n5762 VDD 3.0005
R15754 VDD.n5508 VDD 3.0005
R15755 VDD.n3700 VDD 3.0005
R15756 VDD.n3958 VDD 3.0005
R15757 VDD.n4216 VDD 3.0005
R15758 VDD.n4474 VDD 3.0005
R15759 VDD.n4732 VDD 3.0005
R15760 VDD.n4990 VDD 3.0005
R15761 VDD.n5248 VDD 3.0005
R15762 VDD.n1871 VDD.n1870 2.98717
R15763 VDD.n2192 VDD.n2191 2.98717
R15764 VDD.n2450 VDD.n2449 2.98717
R15765 VDD.n2708 VDD.n2707 2.98717
R15766 VDD.n2966 VDD.n2965 2.98717
R15767 VDD.n3224 VDD.n3223 2.98717
R15768 VDD.n3482 VDD.n3481 2.98717
R15769 VDD.n5802 VDD.n5801 2.98717
R15770 VDD.n5548 VDD.n5547 2.98717
R15771 VDD.n3740 VDD.n3739 2.98717
R15772 VDD.n3998 VDD.n3997 2.98717
R15773 VDD.n4256 VDD.n4255 2.98717
R15774 VDD.n4514 VDD.n4513 2.98717
R15775 VDD.n4772 VDD.n4771 2.98717
R15776 VDD.n5030 VDD.n5029 2.98717
R15777 VDD.n5288 VDD.n5287 2.98717
R15778 VDD.n1916 VDD.n1889 2.72837
R15779 VDD.n2237 VDD.n2210 2.72837
R15780 VDD.n2495 VDD.n2468 2.72837
R15781 VDD.n2753 VDD.n2726 2.72837
R15782 VDD.n3011 VDD.n2984 2.72837
R15783 VDD.n3269 VDD.n3242 2.72837
R15784 VDD.n3527 VDD.n3500 2.72837
R15785 VDD.n5847 VDD.n5820 2.72837
R15786 VDD.n5593 VDD.n5566 2.72837
R15787 VDD.n3785 VDD.n3758 2.72837
R15788 VDD.n4043 VDD.n4016 2.72837
R15789 VDD.n4301 VDD.n4274 2.72837
R15790 VDD.n4559 VDD.n4532 2.72837
R15791 VDD.n4817 VDD.n4790 2.72837
R15792 VDD.n5075 VDD.n5048 2.72837
R15793 VDD.n5333 VDD.n5306 2.72837
R15794 VDD.n477 VDD.n476 2.30978
R15795 VDD.n75 VDD.n74 2.30978
R15796 VDD.n1622 VDD.n1614 2.251
R15797 VDD.n1778 VDD.n1777 2.2278
R15798 VDD.n1986 VDD.n1985 2.2278
R15799 VDD.n2357 VDD.n2356 2.2278
R15800 VDD.n2615 VDD.n2614 2.2278
R15801 VDD.n2873 VDD.n2872 2.2278
R15802 VDD.n3131 VDD.n3130 2.2278
R15803 VDD.n3389 VDD.n3388 2.2278
R15804 VDD.n5712 VDD.n5711 2.2278
R15805 VDD.n5458 VDD.n5457 2.2278
R15806 VDD.n3647 VDD.n3646 2.2278
R15807 VDD.n3905 VDD.n3904 2.2278
R15808 VDD.n4163 VDD.n4162 2.2278
R15809 VDD.n4421 VDD.n4420 2.2278
R15810 VDD.n4679 VDD.n4678 2.2278
R15811 VDD.n4937 VDD.n4936 2.2278
R15812 VDD.n5195 VDD.n5194 2.2278
R15813 VDD VDD.n1633 2.13383
R15814 VDD.n1644 VDD 2.11184
R15815 VDD.n1655 VDD.n1642 1.59861
R15816 VDD.n1630 VDD 1.53093
R15817 VDD.n1981 VDD 1.52828
R15818 VDD.n1772 VDD.n1771 1.51475
R15819 VDD.n2121 VDD.n2120 1.51475
R15820 VDD.n2351 VDD.n2350 1.51475
R15821 VDD.n2609 VDD.n2608 1.51475
R15822 VDD.n2867 VDD.n2866 1.51475
R15823 VDD.n3125 VDD.n3124 1.51475
R15824 VDD.n3383 VDD.n3382 1.51475
R15825 VDD.n5706 VDD.n5705 1.51475
R15826 VDD.n5452 VDD.n5451 1.51475
R15827 VDD.n3641 VDD.n3640 1.51475
R15828 VDD.n3899 VDD.n3898 1.51475
R15829 VDD.n4157 VDD.n4156 1.51475
R15830 VDD.n4415 VDD.n4414 1.51475
R15831 VDD.n4673 VDD.n4672 1.51475
R15832 VDD.n4931 VDD.n4930 1.51475
R15833 VDD.n5189 VDD.n5188 1.51475
R15834 VDD.n1945 VDD.t1042 1.50409
R15835 VDD.n1924 VDD.t864 1.50409
R15836 VDD.n1924 VDD.t1044 1.50409
R15837 VDD.n1918 VDD.n1917 1.49778
R15838 VDD.n2239 VDD.n2238 1.49778
R15839 VDD.n2497 VDD.n2496 1.49778
R15840 VDD.n2755 VDD.n2754 1.49778
R15841 VDD.n3013 VDD.n3012 1.49778
R15842 VDD.n3271 VDD.n3270 1.49778
R15843 VDD.n3529 VDD.n3528 1.49778
R15844 VDD.n5849 VDD.n5848 1.49778
R15845 VDD.n5595 VDD.n5594 1.49778
R15846 VDD.n3787 VDD.n3786 1.49778
R15847 VDD.n4045 VDD.n4044 1.49778
R15848 VDD.n4303 VDD.n4302 1.49778
R15849 VDD.n4561 VDD.n4560 1.49778
R15850 VDD.n4819 VDD.n4818 1.49778
R15851 VDD.n5077 VDD.n5076 1.49778
R15852 VDD.n5335 VDD.n5334 1.49778
R15853 VDD.n2013 VDD.n2012 1.47642
R15854 VDD.n1661 VDD.n1660 1.43354
R15855 VDD.n1740 VDD.n1729 1.42272
R15856 VDD.n2089 VDD.n2078 1.42272
R15857 VDD.n2319 VDD.n2308 1.42272
R15858 VDD.n2577 VDD.n2566 1.42272
R15859 VDD.n2835 VDD.n2824 1.42272
R15860 VDD.n3093 VDD.n3082 1.42272
R15861 VDD.n3351 VDD.n3340 1.42272
R15862 VDD.n5674 VDD.n5663 1.42272
R15863 VDD.n5420 VDD.n5409 1.42272
R15864 VDD.n3609 VDD.n3598 1.42272
R15865 VDD.n3867 VDD.n3856 1.42272
R15866 VDD.n4125 VDD.n4114 1.42272
R15867 VDD.n4383 VDD.n4372 1.42272
R15868 VDD.n4641 VDD.n4630 1.42272
R15869 VDD.n4899 VDD.n4888 1.42272
R15870 VDD.n5157 VDD.n5146 1.42272
R15871 VDD.n1663 VDD.n1662 1.39179
R15872 VDD.n1887 VDD.n1886 1.25748
R15873 VDD.n2208 VDD.n2207 1.25748
R15874 VDD.n2466 VDD.n2465 1.25748
R15875 VDD.n2724 VDD.n2723 1.25748
R15876 VDD.n2982 VDD.n2981 1.25748
R15877 VDD.n3240 VDD.n3239 1.25748
R15878 VDD.n3498 VDD.n3497 1.25748
R15879 VDD.n5818 VDD.n5817 1.25748
R15880 VDD.n5564 VDD.n5563 1.25748
R15881 VDD.n3756 VDD.n3755 1.25748
R15882 VDD.n4014 VDD.n4013 1.25748
R15883 VDD.n4272 VDD.n4271 1.25748
R15884 VDD.n4530 VDD.n4529 1.25748
R15885 VDD.n4788 VDD.n4787 1.25748
R15886 VDD.n5046 VDD.n5045 1.25748
R15887 VDD.n5304 VDD.n5303 1.25748
R15888 VDD.n1651 VDD.n1650 1.25267
R15889 VDD.n1655 VDD.n1654 1.21925
R15890 VDD.n557 VDD.n556 1.12991
R15891 VDD.n615 VDD.n614 1.12991
R15892 VDD.n640 VDD.n639 1.12991
R15893 VDD.n750 VDD.n749 1.12991
R15894 VDD.n703 VDD.n702 1.12991
R15895 VDD.n907 VDD.n906 1.12991
R15896 VDD.n965 VDD.n964 1.12991
R15897 VDD.n990 VDD.n989 1.12991
R15898 VDD.n1100 VDD.n1099 1.12991
R15899 VDD.n1053 VDD.n1052 1.12991
R15900 VDD.n156 VDD.n155 1.12991
R15901 VDD.n214 VDD.n213 1.12991
R15902 VDD.n113 VDD.n112 1.12991
R15903 VDD.n345 VDD.n344 1.12991
R15904 VDD.n298 VDD.n297 1.12991
R15905 VDD.n1336 VDD.n1335 1.12991
R15906 VDD.n1380 VDD.n1379 1.12991
R15907 VDD.n1307 VDD.n1306 1.12991
R15908 VDD.n1466 VDD.n1465 1.12991
R15909 VDD.n1516 VDD.n1515 1.12991
R15910 VDD.n1652 VDD.n1651 1.11354
R15911 VDD.n1631 VDD.n1630 1.11354
R15912 VDD.n1623 VDD.n1613 1.10388
R15913 VDD.n1731 VDD.n1716 1.06717
R15914 VDD.n2080 VDD.n2065 1.06717
R15915 VDD.n2310 VDD.n2295 1.06717
R15916 VDD.n2568 VDD.n2553 1.06717
R15917 VDD.n2826 VDD.n2811 1.06717
R15918 VDD.n3084 VDD.n3069 1.06717
R15919 VDD.n3342 VDD.n3327 1.06717
R15920 VDD.n5665 VDD.n5650 1.06717
R15921 VDD.n5411 VDD.n5396 1.06717
R15922 VDD.n3600 VDD.n3585 1.06717
R15923 VDD.n3858 VDD.n3843 1.06717
R15924 VDD.n4116 VDD.n4101 1.06717
R15925 VDD.n4374 VDD.n4359 1.06717
R15926 VDD.n4632 VDD.n4617 1.06717
R15927 VDD.n4890 VDD.n4875 1.06717
R15928 VDD.n5148 VDD.n5133 1.06717
R15929 VDD.n1608 VDD.n1606 1.06717
R15930 VDD.n1607 VDD 1.06717
R15931 VDD.n1873 VDD.n1872 1.00783
R15932 VDD.n2194 VDD.n2193 1.00687
R15933 VDD.n2452 VDD.n2451 1.00687
R15934 VDD.n2710 VDD.n2709 1.00687
R15935 VDD.n2968 VDD.n2967 1.00687
R15936 VDD.n3226 VDD.n3225 1.00687
R15937 VDD.n3484 VDD.n3483 1.00687
R15938 VDD.n5804 VDD.n5803 1.00687
R15939 VDD.n5550 VDD.n5549 1.00687
R15940 VDD.n3742 VDD.n3741 1.00687
R15941 VDD.n4000 VDD.n3999 1.00687
R15942 VDD.n4258 VDD.n4257 1.00687
R15943 VDD.n4516 VDD.n4515 1.00687
R15944 VDD.n4774 VDD.n4773 1.00687
R15945 VDD.n5032 VDD.n5031 1.00687
R15946 VDD.n5290 VDD.n5289 1.00687
R15947 VDD.n1644 VDD 0.970197
R15948 VDD.n1704 VDD.n1681 0.9605
R15949 VDD.n2053 VDD.n2030 0.9605
R15950 VDD.n2283 VDD.n2260 0.9605
R15951 VDD.n2541 VDD.n2518 0.9605
R15952 VDD.n2799 VDD.n2776 0.9605
R15953 VDD.n3057 VDD.n3034 0.9605
R15954 VDD.n3315 VDD.n3292 0.9605
R15955 VDD.n5638 VDD.n5615 0.9605
R15956 VDD.n5384 VDD.n5361 0.9605
R15957 VDD.n3573 VDD.n3550 0.9605
R15958 VDD.n3831 VDD.n3808 0.9605
R15959 VDD.n4089 VDD.n4066 0.9605
R15960 VDD.n4347 VDD.n4324 0.9605
R15961 VDD.n4605 VDD.n4582 0.9605
R15962 VDD.n4863 VDD.n4840 0.9605
R15963 VDD.n5121 VDD.n5098 0.9605
R15964 VDD.n1603 VDD.n1245 0.939577
R15965 VDD.n5859 VDD.n1982 0.885753
R15966 VDD.n1662 VDD.n1661 0.87764
R15967 VDD.n796 VDD.n407 0.826983
R15968 VDD.n1598 VDD.n1565 0.826983
R15969 VDD.n1933 VDD.n1924 0.800961
R15970 VDD.n5861 VDD 0.78236
R15971 VDD.n1619 VDD.n1618 0.7685
R15972 VDD.n1956 VDD.n1943 0.738962
R15973 VDD.n1638 VDD.n1636 0.686214
R15974 VDD.n1657 VDD.n1656 0.683536
R15975 VDD.n1663 VDD.n1603 0.673542
R15976 VDD.n1693 VDD.n1685 0.6405
R15977 VDD.n2042 VDD.n2034 0.6405
R15978 VDD.n2272 VDD.n2264 0.6405
R15979 VDD.n2530 VDD.n2522 0.6405
R15980 VDD.n2788 VDD.n2780 0.6405
R15981 VDD.n3046 VDD.n3038 0.6405
R15982 VDD.n3304 VDD.n3296 0.6405
R15983 VDD.n5627 VDD.n5619 0.6405
R15984 VDD.n5373 VDD.n5365 0.6405
R15985 VDD.n3562 VDD.n3554 0.6405
R15986 VDD.n3820 VDD.n3812 0.6405
R15987 VDD.n4078 VDD.n4070 0.6405
R15988 VDD.n4336 VDD.n4328 0.6405
R15989 VDD.n4594 VDD.n4586 0.6405
R15990 VDD.n4852 VDD.n4844 0.6405
R15991 VDD.n5110 VDD.n5102 0.6405
R15992 VDD.n1688 VDD.n1687 0.590778
R15993 VDD.n2037 VDD.n2036 0.590778
R15994 VDD.n2267 VDD.n2266 0.590778
R15995 VDD.n2525 VDD.n2524 0.590778
R15996 VDD.n2783 VDD.n2782 0.590778
R15997 VDD.n3041 VDD.n3040 0.590778
R15998 VDD.n3299 VDD.n3298 0.590778
R15999 VDD.n5622 VDD.n5621 0.590778
R16000 VDD.n5368 VDD.n5367 0.590778
R16001 VDD.n3557 VDD.n3556 0.590778
R16002 VDD.n3815 VDD.n3814 0.590778
R16003 VDD.n4073 VDD.n4072 0.590778
R16004 VDD.n4331 VDD.n4330 0.590778
R16005 VDD.n4589 VDD.n4588 0.590778
R16006 VDD.n4847 VDD.n4846 0.590778
R16007 VDD.n5105 VDD.n5104 0.590778
R16008 VDD.n5739 VDD.n5738 0.588569
R16009 VDD.n5485 VDD.n5484 0.588569
R16010 VDD.n1805 VDD.n1804 0.580785
R16011 VDD.n2384 VDD.n2383 0.580785
R16012 VDD.n2642 VDD.n2641 0.580785
R16013 VDD.n2900 VDD.n2899 0.580785
R16014 VDD.n3158 VDD.n3157 0.580785
R16015 VDD.n3416 VDD.n3415 0.580785
R16016 VDD.n3674 VDD.n3673 0.580785
R16017 VDD.n3932 VDD.n3931 0.580785
R16018 VDD.n4190 VDD.n4189 0.580785
R16019 VDD.n4448 VDD.n4447 0.580785
R16020 VDD.n4706 VDD.n4705 0.580785
R16021 VDD.n4964 VDD.n4963 0.580785
R16022 VDD.n5222 VDD.n5221 0.580785
R16023 VDD.n1658 VDD.n1657 0.571929
R16024 VDD.n1660 VDD.n1659 0.558536
R16025 VDD.n795 VDD.n438 0.557954
R16026 VDD.n1597 VDD.n1596 0.557954
R16027 VDD.n1659 VDD.n1658 0.549607
R16028 VDD.n1748 VDD.n1723 0.514389
R16029 VDD.n2097 VDD.n2072 0.514389
R16030 VDD.n2327 VDD.n2302 0.514389
R16031 VDD.n2585 VDD.n2560 0.514389
R16032 VDD.n2843 VDD.n2818 0.514389
R16033 VDD.n3101 VDD.n3076 0.514389
R16034 VDD.n3359 VDD.n3334 0.514389
R16035 VDD.n5682 VDD.n5657 0.514389
R16036 VDD.n5428 VDD.n5403 0.514389
R16037 VDD.n3617 VDD.n3592 0.514389
R16038 VDD.n3875 VDD.n3850 0.514389
R16039 VDD.n4133 VDD.n4108 0.514389
R16040 VDD.n4391 VDD.n4366 0.514389
R16041 VDD.n4649 VDD.n4624 0.514389
R16042 VDD.n4907 VDD.n4882 0.514389
R16043 VDD.n5165 VDD.n5140 0.514389
R16044 VDD.n1977 VDD.n1925 0.5125
R16045 VDD.n1839 VDD.n1826 0.492808
R16046 VDD.n2160 VDD.n2147 0.492808
R16047 VDD.n2418 VDD.n2405 0.492808
R16048 VDD.n2676 VDD.n2663 0.492808
R16049 VDD.n2934 VDD.n2921 0.492808
R16050 VDD.n3192 VDD.n3179 0.492808
R16051 VDD.n3450 VDD.n3437 0.492808
R16052 VDD.n5770 VDD.n5757 0.492808
R16053 VDD.n5516 VDD.n5503 0.492808
R16054 VDD.n3708 VDD.n3695 0.492808
R16055 VDD.n3966 VDD.n3953 0.492808
R16056 VDD.n4224 VDD.n4211 0.492808
R16057 VDD.n4482 VDD.n4469 0.492808
R16058 VDD.n4740 VDD.n4727 0.492808
R16059 VDD.n4998 VDD.n4985 0.492808
R16060 VDD.n5256 VDD.n5243 0.492808
R16061 VDD.n26 VDD 0.476404
R16062 VDD.n1170 VDD 0.476404
R16063 VDD.n1686 VDD.n1665 0.471224
R16064 VDD.n2035 VDD.n2014 0.471224
R16065 VDD.n2265 VDD.n2244 0.471224
R16066 VDD.n2523 VDD.n2502 0.471224
R16067 VDD.n2781 VDD.n2760 0.471224
R16068 VDD.n3039 VDD.n3018 0.471224
R16069 VDD.n3297 VDD.n3276 0.471224
R16070 VDD.n5620 VDD.n5599 0.471224
R16071 VDD.n5366 VDD.n5345 0.471224
R16072 VDD.n3555 VDD.n3534 0.471224
R16073 VDD.n3813 VDD.n3792 0.471224
R16074 VDD.n4071 VDD.n4050 0.471224
R16075 VDD.n4329 VDD.n4308 0.471224
R16076 VDD.n4587 VDD.n4566 0.471224
R16077 VDD.n4845 VDD.n4824 0.471224
R16078 VDD.n5103 VDD.n5082 0.471224
R16079 VDD.n1773 VDD.n1666 0.467504
R16080 VDD.n2122 VDD.n2015 0.467504
R16081 VDD.n2352 VDD.n2245 0.467504
R16082 VDD.n2610 VDD.n2503 0.467504
R16083 VDD.n2868 VDD.n2761 0.467504
R16084 VDD.n3126 VDD.n3019 0.467504
R16085 VDD.n3384 VDD.n3277 0.467504
R16086 VDD.n5707 VDD.n5600 0.467504
R16087 VDD.n5453 VDD.n5346 0.467504
R16088 VDD.n3642 VDD.n3535 0.467504
R16089 VDD.n3900 VDD.n3793 0.467504
R16090 VDD.n4158 VDD.n4051 0.467504
R16091 VDD.n4416 VDD.n4309 0.467504
R16092 VDD.n4674 VDD.n4567 0.467504
R16093 VDD.n4932 VDD.n4825 0.467504
R16094 VDD.n5190 VDD.n5083 0.467504
R16095 VDD.n1654 VDD.n1653 0.464786
R16096 VDD.n1637 VDD 0.457643
R16097 VDD.n1661 VDD.n1623 0.424377
R16098 VDD.n1810 VDD 0.411214
R16099 VDD.n2131 VDD 0.411214
R16100 VDD.n2389 VDD 0.411214
R16101 VDD.n2647 VDD 0.411214
R16102 VDD.n2905 VDD 0.411214
R16103 VDD.n3163 VDD 0.411214
R16104 VDD.n3421 VDD 0.411214
R16105 VDD.n5741 VDD 0.411214
R16106 VDD.n5487 VDD 0.411214
R16107 VDD.n3679 VDD 0.411214
R16108 VDD.n3937 VDD 0.411214
R16109 VDD.n4195 VDD 0.411214
R16110 VDD.n4453 VDD 0.411214
R16111 VDD.n4711 VDD 0.411214
R16112 VDD.n4969 VDD 0.411214
R16113 VDD.n5227 VDD 0.411214
R16114 VDD.n1753 VDD.n1752 0.410606
R16115 VDD.n2102 VDD.n2101 0.410606
R16116 VDD.n2332 VDD.n2331 0.410606
R16117 VDD.n2590 VDD.n2589 0.410606
R16118 VDD.n2848 VDD.n2847 0.410606
R16119 VDD.n3106 VDD.n3105 0.410606
R16120 VDD.n3364 VDD.n3363 0.410606
R16121 VDD.n5687 VDD.n5686 0.410606
R16122 VDD.n5433 VDD.n5432 0.410606
R16123 VDD.n3622 VDD.n3621 0.410606
R16124 VDD.n3880 VDD.n3879 0.410606
R16125 VDD.n4138 VDD.n4137 0.410606
R16126 VDD.n4396 VDD.n4395 0.410606
R16127 VDD.n4654 VDD.n4653 0.410606
R16128 VDD.n4912 VDD.n4911 0.410606
R16129 VDD.n5170 VDD.n5169 0.410606
R16130 VDD.n1921 VDD.n1920 0.409102
R16131 VDD.n2242 VDD.n2241 0.409102
R16132 VDD.n2500 VDD.n2499 0.409102
R16133 VDD.n2758 VDD.n2757 0.409102
R16134 VDD.n3016 VDD.n3015 0.409102
R16135 VDD.n3274 VDD.n3273 0.409102
R16136 VDD.n3532 VDD.n3531 0.409102
R16137 VDD.n3790 VDD.n3789 0.409102
R16138 VDD.n4048 VDD.n4047 0.409102
R16139 VDD.n4306 VDD.n4305 0.409102
R16140 VDD.n4564 VDD.n4563 0.409102
R16141 VDD.n4822 VDD.n4821 0.409102
R16142 VDD.n5080 VDD.n5079 0.409102
R16143 VDD.n5338 VDD.n5337 0.409102
R16144 VDD VDD.n26 0.403703
R16145 VDD VDD.n1170 0.403703
R16146 VDD.n1738 VDD.n1737 0.399706
R16147 VDD.n2087 VDD.n2086 0.399706
R16148 VDD.n2317 VDD.n2316 0.399706
R16149 VDD.n2575 VDD.n2574 0.399706
R16150 VDD.n2833 VDD.n2832 0.399706
R16151 VDD.n3091 VDD.n3090 0.399706
R16152 VDD.n3349 VDD.n3348 0.399706
R16153 VDD.n5672 VDD.n5671 0.399706
R16154 VDD.n5418 VDD.n5417 0.399706
R16155 VDD.n3607 VDD.n3606 0.399706
R16156 VDD.n3865 VDD.n3864 0.399706
R16157 VDD.n4123 VDD.n4122 0.399706
R16158 VDD.n4381 VDD.n4380 0.399706
R16159 VDD.n4639 VDD.n4638 0.399706
R16160 VDD.n4897 VDD.n4896 0.399706
R16161 VDD.n5155 VDD.n5154 0.399706
R16162 VDD.n513 VDD.n464 0.399037
R16163 VDD.n62 VDD.n61 0.399037
R16164 VDD.n1749 VDD.n1748 0.398914
R16165 VDD.n2098 VDD.n2097 0.398914
R16166 VDD.n2328 VDD.n2327 0.398914
R16167 VDD.n2586 VDD.n2585 0.398914
R16168 VDD.n2844 VDD.n2843 0.398914
R16169 VDD.n3102 VDD.n3101 0.398914
R16170 VDD.n3360 VDD.n3359 0.398914
R16171 VDD.n5683 VDD.n5682 0.398914
R16172 VDD.n5429 VDD.n5428 0.398914
R16173 VDD.n3618 VDD.n3617 0.398914
R16174 VDD.n3876 VDD.n3875 0.398914
R16175 VDD.n4134 VDD.n4133 0.398914
R16176 VDD.n4392 VDD.n4391 0.398914
R16177 VDD.n4650 VDD.n4649 0.398914
R16178 VDD.n4908 VDD.n4907 0.398914
R16179 VDD.n5166 VDD.n5165 0.398914
R16180 VDD.n1737 VDD.n1723 0.398403
R16181 VDD.n2086 VDD.n2072 0.398403
R16182 VDD.n2316 VDD.n2302 0.398403
R16183 VDD.n2574 VDD.n2560 0.398403
R16184 VDD.n2832 VDD.n2818 0.398403
R16185 VDD.n3090 VDD.n3076 0.398403
R16186 VDD.n3348 VDD.n3334 0.398403
R16187 VDD.n5671 VDD.n5657 0.398403
R16188 VDD.n5417 VDD.n5403 0.398403
R16189 VDD.n3606 VDD.n3592 0.398403
R16190 VDD.n3864 VDD.n3850 0.398403
R16191 VDD.n4122 VDD.n4108 0.398403
R16192 VDD.n4380 VDD.n4366 0.398403
R16193 VDD.n4638 VDD.n4624 0.398403
R16194 VDD.n4896 VDD.n4882 0.398403
R16195 VDD.n5154 VDD.n5140 0.398403
R16196 VDD.n1656 VDD.n1655 0.384429
R16197 VDD.n1807 VDD.n1806 0.3805
R16198 VDD.n2127 VDD.n2126 0.3805
R16199 VDD.n2386 VDD.n2385 0.3805
R16200 VDD.n2644 VDD.n2643 0.3805
R16201 VDD.n2902 VDD.n2901 0.3805
R16202 VDD.n3160 VDD.n3159 0.3805
R16203 VDD.n3418 VDD.n3417 0.3805
R16204 VDD.n3676 VDD.n3675 0.3805
R16205 VDD.n3934 VDD.n3933 0.3805
R16206 VDD.n4192 VDD.n4191 0.3805
R16207 VDD.n4450 VDD.n4449 0.3805
R16208 VDD.n4708 VDD.n4707 0.3805
R16209 VDD.n4966 VDD.n4965 0.3805
R16210 VDD.n5224 VDD.n5223 0.3805
R16211 VDD.n547 VDD.n546 0.376971
R16212 VDD.n627 VDD.n626 0.376971
R16213 VDD.n787 VDD.n786 0.376971
R16214 VDD.n739 VDD.n738 0.376971
R16215 VDD.n897 VDD.n896 0.376971
R16216 VDD.n977 VDD.n976 0.376971
R16217 VDD.n1137 VDD.n1136 0.376971
R16218 VDD.n1089 VDD.n1088 0.376971
R16219 VDD.n146 VDD.n145 0.376971
R16220 VDD.n226 VDD.n225 0.376971
R16221 VDD.n382 VDD.n381 0.376971
R16222 VDD.n334 VDD.n333 0.376971
R16223 VDD.n1452 VDD.n1451 0.376971
R16224 VDD.n1421 VDD.n1420 0.376971
R16225 VDD.n1266 VDD.n1265 0.376971
R16226 VDD.n1500 VDD.n1499 0.376971
R16227 VDD.n1687 VDD.n1686 0.368458
R16228 VDD.n2036 VDD.n2035 0.368458
R16229 VDD.n2266 VDD.n2265 0.368458
R16230 VDD.n2524 VDD.n2523 0.368458
R16231 VDD.n2782 VDD.n2781 0.368458
R16232 VDD.n3040 VDD.n3039 0.368458
R16233 VDD.n3298 VDD.n3297 0.368458
R16234 VDD.n5621 VDD.n5620 0.368458
R16235 VDD.n5367 VDD.n5366 0.368458
R16236 VDD.n3556 VDD.n3555 0.368458
R16237 VDD.n3814 VDD.n3813 0.368458
R16238 VDD.n4072 VDD.n4071 0.368458
R16239 VDD.n4330 VDD.n4329 0.368458
R16240 VDD.n4588 VDD.n4587 0.368458
R16241 VDD.n4846 VDD.n4845 0.368458
R16242 VDD.n5104 VDD.n5103 0.368458
R16243 VDD.n1688 VDD.n1666 0.361663
R16244 VDD.n2037 VDD.n2015 0.361663
R16245 VDD.n2267 VDD.n2245 0.361663
R16246 VDD.n2525 VDD.n2503 0.361663
R16247 VDD.n2783 VDD.n2761 0.361663
R16248 VDD.n3041 VDD.n3019 0.361663
R16249 VDD.n3299 VDD.n3277 0.361663
R16250 VDD.n5622 VDD.n5600 0.361663
R16251 VDD.n5368 VDD.n5346 0.361663
R16252 VDD.n3557 VDD.n3535 0.361663
R16253 VDD.n3815 VDD.n3793 0.361663
R16254 VDD.n4073 VDD.n4051 0.361663
R16255 VDD.n4331 VDD.n4309 0.361663
R16256 VDD.n4589 VDD.n4567 0.361663
R16257 VDD.n4847 VDD.n4825 0.361663
R16258 VDD.n5105 VDD.n5083 0.361663
R16259 VDD.n1750 VDD.n1749 0.357683
R16260 VDD.n2099 VDD.n2098 0.357683
R16261 VDD.n2329 VDD.n2328 0.357683
R16262 VDD.n2587 VDD.n2586 0.357683
R16263 VDD.n2845 VDD.n2844 0.357683
R16264 VDD.n3103 VDD.n3102 0.357683
R16265 VDD.n3361 VDD.n3360 0.357683
R16266 VDD.n5684 VDD.n5683 0.357683
R16267 VDD.n5430 VDD.n5429 0.357683
R16268 VDD.n3619 VDD.n3618 0.357683
R16269 VDD.n3877 VDD.n3876 0.357683
R16270 VDD.n4135 VDD.n4134 0.357683
R16271 VDD.n4393 VDD.n4392 0.357683
R16272 VDD.n4651 VDD.n4650 0.357683
R16273 VDD.n4909 VDD.n4908 0.357683
R16274 VDD.n5167 VDD.n5166 0.357683
R16275 VDD.n1734 VDD.n1732 0.356056
R16276 VDD.n2083 VDD.n2081 0.356056
R16277 VDD.n2313 VDD.n2311 0.356056
R16278 VDD.n2571 VDD.n2569 0.356056
R16279 VDD.n2829 VDD.n2827 0.356056
R16280 VDD.n3087 VDD.n3085 0.356056
R16281 VDD.n3345 VDD.n3343 0.356056
R16282 VDD.n5668 VDD.n5666 0.356056
R16283 VDD.n5414 VDD.n5412 0.356056
R16284 VDD.n3603 VDD.n3601 0.356056
R16285 VDD.n3861 VDD.n3859 0.356056
R16286 VDD.n4119 VDD.n4117 0.356056
R16287 VDD.n4377 VDD.n4375 0.356056
R16288 VDD.n4635 VDD.n4633 0.356056
R16289 VDD.n4893 VDD.n4891 0.356056
R16290 VDD.n5151 VDD.n5149 0.356056
R16291 VDD.n35 VDD.n34 0.35558
R16292 VDD.n1179 VDD.n1178 0.35558
R16293 VDD.n1836 VDD 0.355332
R16294 VDD.n2157 VDD 0.355332
R16295 VDD.n2415 VDD 0.355332
R16296 VDD.n2673 VDD 0.355332
R16297 VDD.n2931 VDD 0.355332
R16298 VDD.n3189 VDD 0.355332
R16299 VDD.n3447 VDD 0.355332
R16300 VDD.n5767 VDD 0.355332
R16301 VDD.n5513 VDD 0.355332
R16302 VDD.n3705 VDD 0.355332
R16303 VDD.n3963 VDD 0.355332
R16304 VDD.n4221 VDD 0.355332
R16305 VDD.n4479 VDD 0.355332
R16306 VDD.n4737 VDD 0.355332
R16307 VDD.n4995 VDD 0.355332
R16308 VDD.n5253 VDD 0.355332
R16309 VDD.n1918 VDD.n1887 0.349136
R16310 VDD.n2239 VDD.n2208 0.349136
R16311 VDD.n2497 VDD.n2466 0.349136
R16312 VDD.n2755 VDD.n2724 0.349136
R16313 VDD.n3013 VDD.n2982 0.349136
R16314 VDD.n3271 VDD.n3240 0.349136
R16315 VDD.n3529 VDD.n3498 0.349136
R16316 VDD.n5849 VDD.n5818 0.349136
R16317 VDD.n5595 VDD.n5564 0.349136
R16318 VDD.n3787 VDD.n3756 0.349136
R16319 VDD.n4045 VDD.n4014 0.349136
R16320 VDD.n4303 VDD.n4272 0.349136
R16321 VDD.n4561 VDD.n4530 0.349136
R16322 VDD.n4819 VDD.n4788 0.349136
R16323 VDD.n5077 VDD.n5046 0.349136
R16324 VDD.n5335 VDD.n5304 0.349136
R16325 VDD.n0 VDD 0.340206
R16326 VDD.n1144 VDD 0.340206
R16327 VDD.n1692 VDD.n1687 0.340142
R16328 VDD.n2041 VDD.n2036 0.340142
R16329 VDD.n2271 VDD.n2266 0.340142
R16330 VDD.n2529 VDD.n2524 0.340142
R16331 VDD.n2787 VDD.n2782 0.340142
R16332 VDD.n3045 VDD.n3040 0.340142
R16333 VDD.n3303 VDD.n3298 0.340142
R16334 VDD.n5626 VDD.n5621 0.340142
R16335 VDD.n5372 VDD.n5367 0.340142
R16336 VDD.n3561 VDD.n3556 0.340142
R16337 VDD.n3819 VDD.n3814 0.340142
R16338 VDD.n4077 VDD.n4072 0.340142
R16339 VDD.n4335 VDD.n4330 0.340142
R16340 VDD.n4593 VDD.n4588 0.340142
R16341 VDD.n4851 VDD.n4846 0.340142
R16342 VDD.n5109 VDD.n5104 0.340142
R16343 VDD.n1283 VDD 0.330819
R16344 VDD.n1768 VDD.n1671 0.3205
R16345 VDD.n1693 VDD.n1684 0.3205
R16346 VDD.n2117 VDD.n2020 0.3205
R16347 VDD.n2042 VDD.n2033 0.3205
R16348 VDD.n2347 VDD.n2250 0.3205
R16349 VDD.n2272 VDD.n2263 0.3205
R16350 VDD.n2605 VDD.n2508 0.3205
R16351 VDD.n2530 VDD.n2521 0.3205
R16352 VDD.n2863 VDD.n2766 0.3205
R16353 VDD.n2788 VDD.n2779 0.3205
R16354 VDD.n3121 VDD.n3024 0.3205
R16355 VDD.n3046 VDD.n3037 0.3205
R16356 VDD.n3379 VDD.n3282 0.3205
R16357 VDD.n3304 VDD.n3295 0.3205
R16358 VDD.n5702 VDD.n5605 0.3205
R16359 VDD.n5627 VDD.n5618 0.3205
R16360 VDD.n5448 VDD.n5351 0.3205
R16361 VDD.n5373 VDD.n5364 0.3205
R16362 VDD.n3637 VDD.n3540 0.3205
R16363 VDD.n3562 VDD.n3553 0.3205
R16364 VDD.n3895 VDD.n3798 0.3205
R16365 VDD.n3820 VDD.n3811 0.3205
R16366 VDD.n4153 VDD.n4056 0.3205
R16367 VDD.n4078 VDD.n4069 0.3205
R16368 VDD.n4411 VDD.n4314 0.3205
R16369 VDD.n4336 VDD.n4327 0.3205
R16370 VDD.n4669 VDD.n4572 0.3205
R16371 VDD.n4594 VDD.n4585 0.3205
R16372 VDD.n4927 VDD.n4830 0.3205
R16373 VDD.n4852 VDD.n4843 0.3205
R16374 VDD.n5185 VDD.n5088 0.3205
R16375 VDD.n5110 VDD.n5101 0.3205
R16376 VDD.n1919 VDD.n1918 0.314572
R16377 VDD.n2240 VDD.n2239 0.314572
R16378 VDD.n2498 VDD.n2497 0.314572
R16379 VDD.n2756 VDD.n2755 0.314572
R16380 VDD.n3014 VDD.n3013 0.314572
R16381 VDD.n3272 VDD.n3271 0.314572
R16382 VDD.n3530 VDD.n3529 0.314572
R16383 VDD.n5850 VDD.n5849 0.314572
R16384 VDD.n5596 VDD.n5595 0.314572
R16385 VDD.n3788 VDD.n3787 0.314572
R16386 VDD.n4046 VDD.n4045 0.314572
R16387 VDD.n4304 VDD.n4303 0.314572
R16388 VDD.n4562 VDD.n4561 0.314572
R16389 VDD.n4820 VDD.n4819 0.314572
R16390 VDD.n5078 VDD.n5077 0.314572
R16391 VDD.n5336 VDD.n5335 0.314572
R16392 VDD.n1874 VDD.n1873 0.311403
R16393 VDD.n2195 VDD.n2194 0.311403
R16394 VDD.n2453 VDD.n2452 0.311403
R16395 VDD.n2711 VDD.n2710 0.311403
R16396 VDD.n2969 VDD.n2968 0.311403
R16397 VDD.n3227 VDD.n3226 0.311403
R16398 VDD.n3485 VDD.n3484 0.311403
R16399 VDD.n5805 VDD.n5804 0.311403
R16400 VDD.n5551 VDD.n5550 0.311403
R16401 VDD.n3743 VDD.n3742 0.311403
R16402 VDD.n4001 VDD.n4000 0.311403
R16403 VDD.n4259 VDD.n4258 0.311403
R16404 VDD.n4517 VDD.n4516 0.311403
R16405 VDD.n4775 VDD.n4774 0.311403
R16406 VDD.n5033 VDD.n5032 0.311403
R16407 VDD.n5291 VDD.n5290 0.311403
R16408 VDD.n1691 VDD.n1690 0.296036
R16409 VDD.n2040 VDD.n2039 0.296036
R16410 VDD.n2270 VDD.n2269 0.296036
R16411 VDD.n2528 VDD.n2527 0.296036
R16412 VDD.n2786 VDD.n2785 0.296036
R16413 VDD.n3044 VDD.n3043 0.296036
R16414 VDD.n3302 VDD.n3301 0.296036
R16415 VDD.n5625 VDD.n5624 0.296036
R16416 VDD.n5371 VDD.n5370 0.296036
R16417 VDD.n3560 VDD.n3559 0.296036
R16418 VDD.n3818 VDD.n3817 0.296036
R16419 VDD.n4076 VDD.n4075 0.296036
R16420 VDD.n4334 VDD.n4333 0.296036
R16421 VDD.n4592 VDD.n4591 0.296036
R16422 VDD.n4850 VDD.n4849 0.296036
R16423 VDD.n5108 VDD.n5107 0.296036
R16424 VDD.n1650 VDD 0.278761
R16425 VDD VDD.n5863 0.269394
R16426 VDD.n1747 VDD.n1724 0.261214
R16427 VDD.n1727 VDD.n1726 0.261214
R16428 VDD.n2096 VDD.n2073 0.261214
R16429 VDD.n2076 VDD.n2075 0.261214
R16430 VDD.n2326 VDD.n2303 0.261214
R16431 VDD.n2306 VDD.n2305 0.261214
R16432 VDD.n2584 VDD.n2561 0.261214
R16433 VDD.n2564 VDD.n2563 0.261214
R16434 VDD.n2842 VDD.n2819 0.261214
R16435 VDD.n2822 VDD.n2821 0.261214
R16436 VDD.n3100 VDD.n3077 0.261214
R16437 VDD.n3080 VDD.n3079 0.261214
R16438 VDD.n3358 VDD.n3335 0.261214
R16439 VDD.n3338 VDD.n3337 0.261214
R16440 VDD.n5681 VDD.n5658 0.261214
R16441 VDD.n5661 VDD.n5660 0.261214
R16442 VDD.n5427 VDD.n5404 0.261214
R16443 VDD.n5407 VDD.n5406 0.261214
R16444 VDD.n3616 VDD.n3593 0.261214
R16445 VDD.n3596 VDD.n3595 0.261214
R16446 VDD.n3874 VDD.n3851 0.261214
R16447 VDD.n3854 VDD.n3853 0.261214
R16448 VDD.n4132 VDD.n4109 0.261214
R16449 VDD.n4112 VDD.n4111 0.261214
R16450 VDD.n4390 VDD.n4367 0.261214
R16451 VDD.n4370 VDD.n4369 0.261214
R16452 VDD.n4648 VDD.n4625 0.261214
R16453 VDD.n4628 VDD.n4627 0.261214
R16454 VDD.n4906 VDD.n4883 0.261214
R16455 VDD.n4886 VDD.n4885 0.261214
R16456 VDD.n5164 VDD.n5141 0.261214
R16457 VDD.n5144 VDD.n5143 0.261214
R16458 VDD.n1745 VDD.n1725 0.2565
R16459 VDD.n2094 VDD.n2074 0.2565
R16460 VDD.n2324 VDD.n2304 0.2565
R16461 VDD.n2582 VDD.n2562 0.2565
R16462 VDD.n2840 VDD.n2820 0.2565
R16463 VDD.n3098 VDD.n3078 0.2565
R16464 VDD.n3356 VDD.n3336 0.2565
R16465 VDD.n5679 VDD.n5659 0.2565
R16466 VDD.n5425 VDD.n5405 0.2565
R16467 VDD.n3614 VDD.n3594 0.2565
R16468 VDD.n3872 VDD.n3852 0.2565
R16469 VDD.n4130 VDD.n4110 0.2565
R16470 VDD.n4388 VDD.n4368 0.2565
R16471 VDD.n4646 VDD.n4626 0.2565
R16472 VDD.n4904 VDD.n4884 0.2565
R16473 VDD.n5162 VDD.n5142 0.2565
R16474 VDD.n1736 VDD.n1735 0.251889
R16475 VDD.n2085 VDD.n2084 0.251889
R16476 VDD.n2315 VDD.n2314 0.251889
R16477 VDD.n2573 VDD.n2572 0.251889
R16478 VDD.n2831 VDD.n2830 0.251889
R16479 VDD.n3089 VDD.n3088 0.251889
R16480 VDD.n3347 VDD.n3346 0.251889
R16481 VDD.n5670 VDD.n5669 0.251889
R16482 VDD.n5416 VDD.n5415 0.251889
R16483 VDD.n3605 VDD.n3604 0.251889
R16484 VDD.n3863 VDD.n3862 0.251889
R16485 VDD.n4121 VDD.n4120 0.251889
R16486 VDD.n4379 VDD.n4378 0.251889
R16487 VDD.n4637 VDD.n4636 0.251889
R16488 VDD.n4895 VDD.n4894 0.251889
R16489 VDD.n5153 VDD.n5152 0.251889
R16490 VDD.n5851 VDD.n5739 0.25042
R16491 VDD.n5597 VDD.n5485 0.25042
R16492 VDD.n1754 VDD.n1719 0.248103
R16493 VDD.n2103 VDD.n2068 0.248103
R16494 VDD.n2333 VDD.n2298 0.248103
R16495 VDD.n2591 VDD.n2556 0.248103
R16496 VDD.n2849 VDD.n2814 0.248103
R16497 VDD.n3107 VDD.n3072 0.248103
R16498 VDD.n3365 VDD.n3330 0.248103
R16499 VDD.n5688 VDD.n5653 0.248103
R16500 VDD.n5434 VDD.n5399 0.248103
R16501 VDD.n3623 VDD.n3588 0.248103
R16502 VDD.n3881 VDD.n3846 0.248103
R16503 VDD.n4139 VDD.n4104 0.248103
R16504 VDD.n4397 VDD.n4362 0.248103
R16505 VDD.n4655 VDD.n4620 0.248103
R16506 VDD.n4913 VDD.n4878 0.248103
R16507 VDD.n5171 VDD.n5136 0.248103
R16508 VDD.n1770 VDD.n1668 0.247868
R16509 VDD.n2119 VDD.n2017 0.247868
R16510 VDD.n2349 VDD.n2247 0.247868
R16511 VDD.n2607 VDD.n2505 0.247868
R16512 VDD.n2865 VDD.n2763 0.247868
R16513 VDD.n3123 VDD.n3021 0.247868
R16514 VDD.n3381 VDD.n3279 0.247868
R16515 VDD.n5704 VDD.n5602 0.247868
R16516 VDD.n5450 VDD.n5348 0.247868
R16517 VDD.n3639 VDD.n3537 0.247868
R16518 VDD.n3897 VDD.n3795 0.247868
R16519 VDD.n4155 VDD.n4053 0.247868
R16520 VDD.n4413 VDD.n4311 0.247868
R16521 VDD.n4671 VDD.n4569 0.247868
R16522 VDD.n4929 VDD.n4827 0.247868
R16523 VDD.n5187 VDD.n5085 0.247868
R16524 VDD.n808 VDD.n807 0.240091
R16525 VDD.n1191 VDD.n1190 0.240091
R16526 VDD.n1738 VDD.n1721 0.232755
R16527 VDD.n2087 VDD.n2070 0.232755
R16528 VDD.n2317 VDD.n2300 0.232755
R16529 VDD.n2575 VDD.n2558 0.232755
R16530 VDD.n2833 VDD.n2816 0.232755
R16531 VDD.n3091 VDD.n3074 0.232755
R16532 VDD.n3349 VDD.n3332 0.232755
R16533 VDD.n5672 VDD.n5655 0.232755
R16534 VDD.n5418 VDD.n5401 0.232755
R16535 VDD.n3607 VDD.n3590 0.232755
R16536 VDD.n3865 VDD.n3848 0.232755
R16537 VDD.n4123 VDD.n4106 0.232755
R16538 VDD.n4381 VDD.n4364 0.232755
R16539 VDD.n4639 VDD.n4622 0.232755
R16540 VDD.n4897 VDD.n4880 0.232755
R16541 VDD.n5155 VDD.n5138 0.232755
R16542 VDD.n1953 VDD.n1952 0.224662
R16543 VDD.n5862 VDD.n1181 0.221061
R16544 VDD.n1730 VDD.n1722 0.217167
R16545 VDD.n2079 VDD.n2071 0.217167
R16546 VDD.n2309 VDD.n2301 0.217167
R16547 VDD.n2567 VDD.n2559 0.217167
R16548 VDD.n2825 VDD.n2817 0.217167
R16549 VDD.n3083 VDD.n3075 0.217167
R16550 VDD.n3341 VDD.n3333 0.217167
R16551 VDD.n5664 VDD.n5656 0.217167
R16552 VDD.n5410 VDD.n5402 0.217167
R16553 VDD.n3599 VDD.n3591 0.217167
R16554 VDD.n3857 VDD.n3849 0.217167
R16555 VDD.n4115 VDD.n4107 0.217167
R16556 VDD.n4373 VDD.n4365 0.217167
R16557 VDD.n4631 VDD.n4623 0.217167
R16558 VDD.n4889 VDD.n4881 0.217167
R16559 VDD.n5147 VDD.n5139 0.217167
R16560 VDD.n512 VDD.n511 0.212557
R16561 VDD.n110 VDD.n109 0.212557
R16562 VDD.n407 VDD.n406 0.211096
R16563 VDD.n1565 VDD.n1564 0.211096
R16564 VDD.n481 VDD 0.210222
R16565 VDD.n79 VDD 0.210222
R16566 VDD.n1702 VDD.n1701 0.204667
R16567 VDD.n2051 VDD.n2050 0.204667
R16568 VDD.n2281 VDD.n2280 0.204667
R16569 VDD.n2539 VDD.n2538 0.204667
R16570 VDD.n2797 VDD.n2796 0.204667
R16571 VDD.n3055 VDD.n3054 0.204667
R16572 VDD.n3313 VDD.n3312 0.204667
R16573 VDD.n5636 VDD.n5635 0.204667
R16574 VDD.n5382 VDD.n5381 0.204667
R16575 VDD.n3571 VDD.n3570 0.204667
R16576 VDD.n3829 VDD.n3828 0.204667
R16577 VDD.n4087 VDD.n4086 0.204667
R16578 VDD.n4345 VDD.n4344 0.204667
R16579 VDD.n4603 VDD.n4602 0.204667
R16580 VDD.n4861 VDD.n4860 0.204667
R16581 VDD.n5119 VDD.n5118 0.204667
R16582 VDD.n1662 VDD 0.2005
R16583 VDD.n1703 VDD.n1667 0.199111
R16584 VDD.n2052 VDD.n2016 0.199111
R16585 VDD.n2282 VDD.n2246 0.199111
R16586 VDD.n2540 VDD.n2504 0.199111
R16587 VDD.n2798 VDD.n2762 0.199111
R16588 VDD.n3056 VDD.n3020 0.199111
R16589 VDD.n3314 VDD.n3278 0.199111
R16590 VDD.n5637 VDD.n5601 0.199111
R16591 VDD.n5383 VDD.n5347 0.199111
R16592 VDD.n3572 VDD.n3536 0.199111
R16593 VDD.n3830 VDD.n3794 0.199111
R16594 VDD.n4088 VDD.n4052 0.199111
R16595 VDD.n4346 VDD.n4310 0.199111
R16596 VDD.n4604 VDD.n4568 0.199111
R16597 VDD.n4862 VDD.n4826 0.199111
R16598 VDD.n5120 VDD.n5084 0.199111
R16599 VDD.n28 VDD 0.196824
R16600 VDD.n1172 VDD 0.196824
R16601 VDD.n1816 VDD.n1815 0.192557
R16602 VDD.n2137 VDD.n2136 0.192557
R16603 VDD.n2395 VDD.n2394 0.192557
R16604 VDD.n2653 VDD.n2652 0.192557
R16605 VDD.n2911 VDD.n2910 0.192557
R16606 VDD.n3169 VDD.n3168 0.192557
R16607 VDD.n3427 VDD.n3426 0.192557
R16608 VDD.n5747 VDD.n5746 0.192557
R16609 VDD.n5493 VDD.n5492 0.192557
R16610 VDD.n3685 VDD.n3684 0.192557
R16611 VDD.n3943 VDD.n3942 0.192557
R16612 VDD.n4201 VDD.n4200 0.192557
R16613 VDD.n4459 VDD.n4458 0.192557
R16614 VDD.n4717 VDD.n4716 0.192557
R16615 VDD.n4975 VDD.n4974 0.192557
R16616 VDD.n5233 VDD.n5232 0.192557
R16617 VDD.n1811 VDD.n1810 0.192167
R16618 VDD.n2132 VDD.n2131 0.192167
R16619 VDD.n2390 VDD.n2389 0.192167
R16620 VDD.n2648 VDD.n2647 0.192167
R16621 VDD.n2906 VDD.n2905 0.192167
R16622 VDD.n3164 VDD.n3163 0.192167
R16623 VDD.n3422 VDD.n3421 0.192167
R16624 VDD.n5742 VDD.n5741 0.192167
R16625 VDD.n5488 VDD.n5487 0.192167
R16626 VDD.n3680 VDD.n3679 0.192167
R16627 VDD.n3938 VDD.n3937 0.192167
R16628 VDD.n4196 VDD.n4195 0.192167
R16629 VDD.n4454 VDD.n4453 0.192167
R16630 VDD.n4712 VDD.n4711 0.192167
R16631 VDD.n4970 VDD.n4969 0.192167
R16632 VDD.n5228 VDD.n5227 0.192167
R16633 VDD.n5863 VDD.n863 0.189
R16634 VDD.n34 VDD.n33 0.183651
R16635 VDD.n1178 VDD.n1177 0.183651
R16636 VDD.n1804 VDD.n1776 0.180841
R16637 VDD.n2012 VDD.n1984 0.180841
R16638 VDD.n2383 VDD.n2355 0.180841
R16639 VDD.n2641 VDD.n2613 0.180841
R16640 VDD.n2899 VDD.n2871 0.180841
R16641 VDD.n3157 VDD.n3129 0.180841
R16642 VDD.n3415 VDD.n3387 0.180841
R16643 VDD.n5738 VDD.n5710 0.180841
R16644 VDD.n5484 VDD.n5456 0.180841
R16645 VDD.n3673 VDD.n3645 0.180841
R16646 VDD.n3931 VDD.n3903 0.180841
R16647 VDD.n4189 VDD.n4161 0.180841
R16648 VDD.n4447 VDD.n4419 0.180841
R16649 VDD.n4705 VDD.n4677 0.180841
R16650 VDD.n4963 VDD.n4935 0.180841
R16651 VDD.n5221 VDD.n5193 0.180841
R16652 VDD.n511 VDD.n510 0.175873
R16653 VDD.n109 VDD.n108 0.175873
R16654 VDD.n1599 VDD.n1548 0.168948
R16655 VDD.n1760 VDD.n1759 0.164944
R16656 VDD.n1759 VDD.n1711 0.164944
R16657 VDD.n2109 VDD.n2108 0.164944
R16658 VDD.n2108 VDD.n2060 0.164944
R16659 VDD.n2339 VDD.n2338 0.164944
R16660 VDD.n2338 VDD.n2290 0.164944
R16661 VDD.n2597 VDD.n2596 0.164944
R16662 VDD.n2596 VDD.n2548 0.164944
R16663 VDD.n2855 VDD.n2854 0.164944
R16664 VDD.n2854 VDD.n2806 0.164944
R16665 VDD.n3113 VDD.n3112 0.164944
R16666 VDD.n3112 VDD.n3064 0.164944
R16667 VDD.n3371 VDD.n3370 0.164944
R16668 VDD.n3370 VDD.n3322 0.164944
R16669 VDD.n5694 VDD.n5693 0.164944
R16670 VDD.n5693 VDD.n5645 0.164944
R16671 VDD.n5440 VDD.n5439 0.164944
R16672 VDD.n5439 VDD.n5391 0.164944
R16673 VDD.n3629 VDD.n3628 0.164944
R16674 VDD.n3628 VDD.n3580 0.164944
R16675 VDD.n3887 VDD.n3886 0.164944
R16676 VDD.n3886 VDD.n3838 0.164944
R16677 VDD.n4145 VDD.n4144 0.164944
R16678 VDD.n4144 VDD.n4096 0.164944
R16679 VDD.n4403 VDD.n4402 0.164944
R16680 VDD.n4402 VDD.n4354 0.164944
R16681 VDD.n4661 VDD.n4660 0.164944
R16682 VDD.n4660 VDD.n4612 0.164944
R16683 VDD.n4919 VDD.n4918 0.164944
R16684 VDD.n4918 VDD.n4870 0.164944
R16685 VDD.n5177 VDD.n5176 0.164944
R16686 VDD.n5176 VDD.n5128 0.164944
R16687 VDD.n1710 VDD.n1709 0.159358
R16688 VDD.n2059 VDD.n2058 0.159358
R16689 VDD.n2289 VDD.n2288 0.159358
R16690 VDD.n2547 VDD.n2546 0.159358
R16691 VDD.n2805 VDD.n2804 0.159358
R16692 VDD.n3063 VDD.n3062 0.159358
R16693 VDD.n3321 VDD.n3320 0.159358
R16694 VDD.n5644 VDD.n5643 0.159358
R16695 VDD.n5390 VDD.n5389 0.159358
R16696 VDD.n3579 VDD.n3578 0.159358
R16697 VDD.n3837 VDD.n3836 0.159358
R16698 VDD.n4095 VDD.n4094 0.159358
R16699 VDD.n4353 VDD.n4352 0.159358
R16700 VDD.n4611 VDD.n4610 0.159358
R16701 VDD.n4869 VDD.n4868 0.159358
R16702 VDD.n5127 VDD.n5126 0.159358
R16703 VDD.n1709 VDD.n1708 0.15889
R16704 VDD.n2058 VDD.n2057 0.15889
R16705 VDD.n2288 VDD.n2287 0.15889
R16706 VDD.n2546 VDD.n2545 0.15889
R16707 VDD.n2804 VDD.n2803 0.15889
R16708 VDD.n3062 VDD.n3061 0.15889
R16709 VDD.n3320 VDD.n3319 0.15889
R16710 VDD.n5643 VDD.n5642 0.15889
R16711 VDD.n5389 VDD.n5388 0.15889
R16712 VDD.n3578 VDD.n3577 0.15889
R16713 VDD.n3836 VDD.n3835 0.15889
R16714 VDD.n4094 VDD.n4093 0.15889
R16715 VDD.n4352 VDD.n4351 0.15889
R16716 VDD.n4610 VDD.n4609 0.15889
R16717 VDD.n4868 VDD.n4867 0.15889
R16718 VDD.n5126 VDD.n5125 0.15889
R16719 VDD.n438 VDD.n437 0.155541
R16720 VDD.n1596 VDD.n1595 0.155541
R16721 VDD.n27 VDD 0.145087
R16722 VDD.n1171 VDD 0.145087
R16723 VDD VDD.n820 0.137071
R16724 VDD VDD.n1203 0.137071
R16725 VDD.n5339 VDD.n5338 0.135642
R16726 VDD.n5861 VDD.n1663 0.134625
R16727 VDD.n852 VDD.n851 0.128415
R16728 VDD.n1235 VDD.n1234 0.128415
R16729 VDD.n464 VDD.n462 0.120987
R16730 VDD.n61 VDD.n59 0.120987
R16731 VDD.n853 VDD.n852 0.119283
R16732 VDD.n1236 VDD.n1235 0.119283
R16733 VDD.n5851 VDD.n5850 0.118114
R16734 VDD.n5597 VDD.n5596 0.118114
R16735 VDD.n1774 VDD.n1773 0.117306
R16736 VDD.n2123 VDD.n2122 0.117306
R16737 VDD.n2353 VDD.n2352 0.117306
R16738 VDD.n2611 VDD.n2610 0.117306
R16739 VDD.n2869 VDD.n2868 0.117306
R16740 VDD.n3127 VDD.n3126 0.117306
R16741 VDD.n3385 VDD.n3384 0.117306
R16742 VDD.n5708 VDD.n5707 0.117306
R16743 VDD.n5454 VDD.n5453 0.117306
R16744 VDD.n3643 VDD.n3642 0.117306
R16745 VDD.n3901 VDD.n3900 0.117306
R16746 VDD.n4159 VDD.n4158 0.117306
R16747 VDD.n4417 VDD.n4416 0.117306
R16748 VDD.n4675 VDD.n4674 0.117306
R16749 VDD.n4933 VDD.n4932 0.117306
R16750 VDD.n5191 VDD.n5190 0.117306
R16751 VDD.n794 VDD.n793 0.116581
R16752 VDD.n848 VDD.n847 0.1155
R16753 VDD.n847 VDD.n845 0.1155
R16754 VDD.n842 VDD.n841 0.1155
R16755 VDD.n841 VDD.n839 0.1155
R16756 VDD.n836 VDD.n835 0.1155
R16757 VDD.n835 VDD.n833 0.1155
R16758 VDD.n830 VDD.n829 0.1155
R16759 VDD.n829 VDD.n827 0.1155
R16760 VDD.n1231 VDD.n1230 0.1155
R16761 VDD.n1230 VDD.n1228 0.1155
R16762 VDD.n1225 VDD.n1224 0.1155
R16763 VDD.n1224 VDD.n1222 0.1155
R16764 VDD.n1219 VDD.n1218 0.1155
R16765 VDD.n1218 VDD.n1216 0.1155
R16766 VDD.n1213 VDD.n1212 0.1155
R16767 VDD.n1212 VDD.n1210 0.1155
R16768 VDD.n862 VDD 0.109094
R16769 VDD.n1245 VDD 0.109094
R16770 VDD.n862 VDD.n861 0.107922
R16771 VDD.n1245 VDD.n1244 0.107922
R16772 VDD.n1948 VDD.n1947 0.107375
R16773 VDD.n1952 VDD.n1948 0.107375
R16774 VDD.n1856 VDD.n1843 0.104784
R16775 VDD.n1857 VDD.n1856 0.104784
R16776 VDD.n2177 VDD.n2164 0.104784
R16777 VDD.n2178 VDD.n2177 0.104784
R16778 VDD.n2435 VDD.n2422 0.104784
R16779 VDD.n2436 VDD.n2435 0.104784
R16780 VDD.n2693 VDD.n2680 0.104784
R16781 VDD.n2694 VDD.n2693 0.104784
R16782 VDD.n2951 VDD.n2938 0.104784
R16783 VDD.n2952 VDD.n2951 0.104784
R16784 VDD.n3209 VDD.n3196 0.104784
R16785 VDD.n3210 VDD.n3209 0.104784
R16786 VDD.n3467 VDD.n3454 0.104784
R16787 VDD.n3468 VDD.n3467 0.104784
R16788 VDD.n5787 VDD.n5774 0.104784
R16789 VDD.n5788 VDD.n5787 0.104784
R16790 VDD.n5533 VDD.n5520 0.104784
R16791 VDD.n5534 VDD.n5533 0.104784
R16792 VDD.n3725 VDD.n3712 0.104784
R16793 VDD.n3726 VDD.n3725 0.104784
R16794 VDD.n3983 VDD.n3970 0.104784
R16795 VDD.n3984 VDD.n3983 0.104784
R16796 VDD.n4241 VDD.n4228 0.104784
R16797 VDD.n4242 VDD.n4241 0.104784
R16798 VDD.n4499 VDD.n4486 0.104784
R16799 VDD.n4500 VDD.n4499 0.104784
R16800 VDD.n4757 VDD.n4744 0.104784
R16801 VDD.n4758 VDD.n4757 0.104784
R16802 VDD.n5015 VDD.n5002 0.104784
R16803 VDD.n5016 VDD.n5015 0.104784
R16804 VDD.n5273 VDD.n5260 0.104784
R16805 VDD.n5274 VDD.n5273 0.104784
R16806 VDD.n797 VDD.n390 0.102139
R16807 VDD.n1975 VDD.n1974 0.100461
R16808 VDD.n1944 VDD.n1940 0.100461
R16809 VDD.n1974 VDD.n1973 0.0999624
R16810 VDD.n1958 VDD.n1940 0.0999624
R16811 VDD.n1873 VDD.n1842 0.0972991
R16812 VDD.n2194 VDD.n2163 0.0972991
R16813 VDD.n2452 VDD.n2421 0.0972991
R16814 VDD.n2710 VDD.n2679 0.0972991
R16815 VDD.n2968 VDD.n2937 0.0972991
R16816 VDD.n3226 VDD.n3195 0.0972991
R16817 VDD.n3484 VDD.n3453 0.0972991
R16818 VDD.n5804 VDD.n5773 0.0972991
R16819 VDD.n5550 VDD.n5519 0.0972991
R16820 VDD.n3742 VDD.n3711 0.0972991
R16821 VDD.n4000 VDD.n3969 0.0972991
R16822 VDD.n4258 VDD.n4227 0.0972991
R16823 VDD.n4516 VDD.n4485 0.0972991
R16824 VDD.n4774 VDD.n4743 0.0972991
R16825 VDD.n5032 VDD.n5001 0.0972991
R16826 VDD.n5290 VDD.n5259 0.0972991
R16827 VDD.n1811 VDD 0.0963333
R16828 VDD.n2132 VDD 0.0963333
R16829 VDD.n2390 VDD 0.0963333
R16830 VDD.n2648 VDD 0.0963333
R16831 VDD.n2906 VDD 0.0963333
R16832 VDD.n3164 VDD 0.0963333
R16833 VDD.n3422 VDD 0.0963333
R16834 VDD.n5742 VDD 0.0963333
R16835 VDD.n5488 VDD 0.0963333
R16836 VDD.n3680 VDD 0.0963333
R16837 VDD.n3938 VDD 0.0963333
R16838 VDD.n4196 VDD 0.0963333
R16839 VDD.n4454 VDD 0.0963333
R16840 VDD.n4712 VDD 0.0963333
R16841 VDD.n4970 VDD 0.0963333
R16842 VDD.n5228 VDD 0.0963333
R16843 VDD.n1935 VDD.n1934 0.0960166
R16844 VDD.n1936 VDD.n1935 0.095518
R16845 VDD.n853 VDD 0.0950313
R16846 VDD.n1236 VDD 0.0950313
R16847 VDD.n1841 VDD 0.0948131
R16848 VDD.n2162 VDD 0.0948131
R16849 VDD.n2420 VDD 0.0948131
R16850 VDD.n2678 VDD 0.0948131
R16851 VDD.n2936 VDD 0.0948131
R16852 VDD.n3194 VDD 0.0948131
R16853 VDD.n3452 VDD 0.0948131
R16854 VDD.n5772 VDD 0.0948131
R16855 VDD.n5518 VDD 0.0948131
R16856 VDD.n3710 VDD 0.0948131
R16857 VDD.n3968 VDD 0.0948131
R16858 VDD.n4226 VDD 0.0948131
R16859 VDD.n4484 VDD 0.0948131
R16860 VDD.n4742 VDD 0.0948131
R16861 VDD.n5000 VDD 0.0948131
R16862 VDD.n5258 VDD 0.0948131
R16863 VDD.n1875 VDD.n1817 0.0945934
R16864 VDD.n2196 VDD.n2138 0.0945934
R16865 VDD.n2454 VDD.n2396 0.0945934
R16866 VDD.n2712 VDD.n2654 0.0945934
R16867 VDD.n2970 VDD.n2912 0.0945934
R16868 VDD.n3228 VDD.n3170 0.0945934
R16869 VDD.n3486 VDD.n3428 0.0945934
R16870 VDD.n5806 VDD.n5748 0.0945934
R16871 VDD.n5552 VDD.n5494 0.0945934
R16872 VDD.n3744 VDD.n3686 0.0945934
R16873 VDD.n4002 VDD.n3944 0.0945934
R16874 VDD.n4260 VDD.n4202 0.0945934
R16875 VDD.n4518 VDD.n4460 0.0945934
R16876 VDD.n4776 VDD.n4718 0.0945934
R16877 VDD.n5034 VDD.n4976 0.0945934
R16878 VDD.n5292 VDD.n5234 0.0945934
R16879 VDD.n5860 VDD.n1921 0.0944319
R16880 VDD.n5858 VDD.n2242 0.0944319
R16881 VDD.n5857 VDD.n2500 0.0944319
R16882 VDD.n5856 VDD.n2758 0.0944319
R16883 VDD.n5855 VDD.n3016 0.0944319
R16884 VDD.n5854 VDD.n3274 0.0944319
R16885 VDD.n5853 VDD.n3532 0.0944319
R16886 VDD.n5344 VDD.n3790 0.0944319
R16887 VDD.n5343 VDD.n4048 0.0944319
R16888 VDD.n5342 VDD.n4306 0.0944319
R16889 VDD.n5341 VDD.n4564 0.0944319
R16890 VDD.n5340 VDD.n4822 0.0944319
R16891 VDD.n5339 VDD.n5080 0.0944319
R16892 VDD.n1836 VDD 0.0902606
R16893 VDD.n2157 VDD 0.0902606
R16894 VDD.n2415 VDD 0.0902606
R16895 VDD.n2673 VDD 0.0902606
R16896 VDD.n2931 VDD 0.0902606
R16897 VDD.n3189 VDD 0.0902606
R16898 VDD.n3447 VDD 0.0902606
R16899 VDD.n5767 VDD 0.0902606
R16900 VDD.n5513 VDD 0.0902606
R16901 VDD.n3705 VDD 0.0902606
R16902 VDD.n3963 VDD 0.0902606
R16903 VDD.n4221 VDD 0.0902606
R16904 VDD.n4479 VDD 0.0902606
R16905 VDD.n4737 VDD 0.0902606
R16906 VDD.n4995 VDD 0.0902606
R16907 VDD.n5253 VDD 0.0902606
R16908 VDD.n794 VDD 0.0900726
R16909 VDD.n533 VDD.n531 0.0892839
R16910 VDD.n883 VDD.n881 0.0892839
R16911 VDD.n132 VDD.n130 0.0892839
R16912 VDD.n1251 VDD.n1249 0.088354
R16913 VDD.n1797 VDD.n1778 0.0864543
R16914 VDD.n1800 VDD.n1778 0.0864543
R16915 VDD.n2005 VDD.n1986 0.0864543
R16916 VDD.n2008 VDD.n1986 0.0864543
R16917 VDD.n2376 VDD.n2357 0.0864543
R16918 VDD.n2379 VDD.n2357 0.0864543
R16919 VDD.n2634 VDD.n2615 0.0864543
R16920 VDD.n2637 VDD.n2615 0.0864543
R16921 VDD.n2892 VDD.n2873 0.0864543
R16922 VDD.n2895 VDD.n2873 0.0864543
R16923 VDD.n3150 VDD.n3131 0.0864543
R16924 VDD.n3153 VDD.n3131 0.0864543
R16925 VDD.n3408 VDD.n3389 0.0864543
R16926 VDD.n3411 VDD.n3389 0.0864543
R16927 VDD.n5731 VDD.n5712 0.0864543
R16928 VDD.n5734 VDD.n5712 0.0864543
R16929 VDD.n5477 VDD.n5458 0.0864543
R16930 VDD.n5480 VDD.n5458 0.0864543
R16931 VDD.n3666 VDD.n3647 0.0864543
R16932 VDD.n3669 VDD.n3647 0.0864543
R16933 VDD.n3924 VDD.n3905 0.0864543
R16934 VDD.n3927 VDD.n3905 0.0864543
R16935 VDD.n4182 VDD.n4163 0.0864543
R16936 VDD.n4185 VDD.n4163 0.0864543
R16937 VDD.n4440 VDD.n4421 0.0864543
R16938 VDD.n4443 VDD.n4421 0.0864543
R16939 VDD.n4698 VDD.n4679 0.0864543
R16940 VDD.n4701 VDD.n4679 0.0864543
R16941 VDD.n4956 VDD.n4937 0.0864543
R16942 VDD.n4959 VDD.n4937 0.0864543
R16943 VDD.n5214 VDD.n5195 0.0864543
R16944 VDD.n5217 VDD.n5195 0.0864543
R16945 VDD.n5862 VDD.n5861 0.0862917
R16946 VDD.n1774 VDD.n1665 0.0855148
R16947 VDD.n2123 VDD.n2014 0.0855148
R16948 VDD.n2353 VDD.n2244 0.0855148
R16949 VDD.n2611 VDD.n2502 0.0855148
R16950 VDD.n2869 VDD.n2760 0.0855148
R16951 VDD.n3127 VDD.n3018 0.0855148
R16952 VDD.n3385 VDD.n3276 0.0855148
R16953 VDD.n5708 VDD.n5599 0.0855148
R16954 VDD.n5454 VDD.n5345 0.0855148
R16955 VDD.n3643 VDD.n3534 0.0855148
R16956 VDD.n3901 VDD.n3792 0.0855148
R16957 VDD.n4159 VDD.n4050 0.0855148
R16958 VDD.n4417 VDD.n4308 0.0855148
R16959 VDD.n4675 VDD.n4566 0.0855148
R16960 VDD.n4933 VDD.n4824 0.0855148
R16961 VDD.n5191 VDD.n5082 0.0855148
R16962 VDD.n26 VDD.n25 0.0849867
R16963 VDD.n1170 VDD.n1169 0.0849867
R16964 VDD.n5851 VDD.n5709 0.0841827
R16965 VDD.n5597 VDD.n5455 0.0841827
R16966 VDD.n1832 VDD.n1825 0.0832206
R16967 VDD.n2153 VDD.n2146 0.0832206
R16968 VDD.n2411 VDD.n2404 0.0832206
R16969 VDD.n2669 VDD.n2662 0.0832206
R16970 VDD.n2927 VDD.n2920 0.0832206
R16971 VDD.n3185 VDD.n3178 0.0832206
R16972 VDD.n3443 VDD.n3436 0.0832206
R16973 VDD.n5763 VDD.n5756 0.0832206
R16974 VDD.n5509 VDD.n5502 0.0832206
R16975 VDD.n3701 VDD.n3694 0.0832206
R16976 VDD.n3959 VDD.n3952 0.0832206
R16977 VDD.n4217 VDD.n4210 0.0832206
R16978 VDD.n4475 VDD.n4468 0.0832206
R16979 VDD.n4733 VDD.n4726 0.0832206
R16980 VDD.n4991 VDD.n4984 0.0832206
R16981 VDD.n5249 VDD.n5242 0.0832206
R16982 VDD.n1180 VDD.n1143 0.082109
R16983 VDD.n1727 VDD.n1723 0.07913
R16984 VDD.n2076 VDD.n2072 0.07913
R16985 VDD.n2306 VDD.n2302 0.07913
R16986 VDD.n2564 VDD.n2560 0.07913
R16987 VDD.n2822 VDD.n2818 0.07913
R16988 VDD.n3080 VDD.n3076 0.07913
R16989 VDD.n3338 VDD.n3334 0.07913
R16990 VDD.n5661 VDD.n5657 0.07913
R16991 VDD.n5407 VDD.n5403 0.07913
R16992 VDD.n3596 VDD.n3592 0.07913
R16993 VDD.n3854 VDD.n3850 0.07913
R16994 VDD.n4112 VDD.n4108 0.07913
R16995 VDD.n4370 VDD.n4366 0.07913
R16996 VDD.n4628 VDD.n4624 0.07913
R16997 VDD.n4886 VDD.n4882 0.07913
R16998 VDD.n5144 VDD.n5140 0.07913
R16999 VDD.n1835 VDD.n1828 0.078625
R17000 VDD.n2156 VDD.n2149 0.078625
R17001 VDD.n2414 VDD.n2407 0.078625
R17002 VDD.n2672 VDD.n2665 0.078625
R17003 VDD.n2930 VDD.n2923 0.078625
R17004 VDD.n3188 VDD.n3181 0.078625
R17005 VDD.n3446 VDD.n3439 0.078625
R17006 VDD.n5766 VDD.n5759 0.078625
R17007 VDD.n5512 VDD.n5505 0.078625
R17008 VDD.n3704 VDD.n3697 0.078625
R17009 VDD.n3962 VDD.n3955 0.078625
R17010 VDD.n4220 VDD.n4213 0.078625
R17011 VDD.n4478 VDD.n4471 0.078625
R17012 VDD.n4736 VDD.n4729 0.078625
R17013 VDD.n4994 VDD.n4987 0.078625
R17014 VDD.n5252 VDD.n5245 0.078625
R17015 VDD.n33 VDD.n30 0.0777407
R17016 VDD.n1177 VDD.n1174 0.0777407
R17017 VDD.n1748 VDD.n1747 0.0773443
R17018 VDD.n2097 VDD.n2096 0.0773443
R17019 VDD.n2327 VDD.n2326 0.0773443
R17020 VDD.n2585 VDD.n2584 0.0773443
R17021 VDD.n2843 VDD.n2842 0.0773443
R17022 VDD.n3101 VDD.n3100 0.0773443
R17023 VDD.n3359 VDD.n3358 0.0773443
R17024 VDD.n5682 VDD.n5681 0.0773443
R17025 VDD.n5428 VDD.n5427 0.0773443
R17026 VDD.n3617 VDD.n3616 0.0773443
R17027 VDD.n3875 VDD.n3874 0.0773443
R17028 VDD.n4133 VDD.n4132 0.0773443
R17029 VDD.n4391 VDD.n4390 0.0773443
R17030 VDD.n4649 VDD.n4648 0.0773443
R17031 VDD.n4907 VDD.n4906 0.0773443
R17032 VDD.n5165 VDD.n5164 0.0773443
R17033 VDD.n1690 VDD.n1688 0.0755586
R17034 VDD.n2039 VDD.n2037 0.0755586
R17035 VDD.n2269 VDD.n2267 0.0755586
R17036 VDD.n2527 VDD.n2525 0.0755586
R17037 VDD.n2785 VDD.n2783 0.0755586
R17038 VDD.n3043 VDD.n3041 0.0755586
R17039 VDD.n3301 VDD.n3299 0.0755586
R17040 VDD.n5624 VDD.n5622 0.0755586
R17041 VDD.n5370 VDD.n5368 0.0755586
R17042 VDD.n3559 VDD.n3557 0.0755586
R17043 VDD.n3817 VDD.n3815 0.0755586
R17044 VDD.n4075 VDD.n4073 0.0755586
R17045 VDD.n4333 VDD.n4331 0.0755586
R17046 VDD.n4591 VDD.n4589 0.0755586
R17047 VDD.n4849 VDD.n4847 0.0755586
R17048 VDD.n5107 VDD.n5105 0.0755586
R17049 VDD.n510 VDD.n507 0.0734782
R17050 VDD.n437 VDD.n434 0.0734782
R17051 VDD.n108 VDD.n105 0.0734782
R17052 VDD.n1595 VDD.n1592 0.0734782
R17053 VDD.n1842 VDD.n1841 0.0710611
R17054 VDD.n2163 VDD.n2162 0.0710611
R17055 VDD.n2421 VDD.n2420 0.0710611
R17056 VDD.n2679 VDD.n2678 0.0710611
R17057 VDD.n2937 VDD.n2936 0.0710611
R17058 VDD.n3195 VDD.n3194 0.0710611
R17059 VDD.n3453 VDD.n3452 0.0710611
R17060 VDD.n5773 VDD.n5772 0.0710611
R17061 VDD.n5519 VDD.n5518 0.0710611
R17062 VDD.n3711 VDD.n3710 0.0710611
R17063 VDD.n3969 VDD.n3968 0.0710611
R17064 VDD.n4227 VDD.n4226 0.0710611
R17065 VDD.n4485 VDD.n4484 0.0710611
R17066 VDD.n4743 VDD.n4742 0.0710611
R17067 VDD.n5001 VDD.n5000 0.0710611
R17068 VDD.n5259 VDD.n5258 0.0710611
R17069 VDD.n1919 VDD.n1816 0.0705353
R17070 VDD.n2240 VDD.n2137 0.0705353
R17071 VDD.n2498 VDD.n2395 0.0705353
R17072 VDD.n2756 VDD.n2653 0.0705353
R17073 VDD.n3014 VDD.n2911 0.0705353
R17074 VDD.n3272 VDD.n3169 0.0705353
R17075 VDD.n3530 VDD.n3427 0.0705353
R17076 VDD.n5850 VDD.n5747 0.0705353
R17077 VDD.n5596 VDD.n5493 0.0705353
R17078 VDD.n3788 VDD.n3685 0.0705353
R17079 VDD.n4046 VDD.n3943 0.0705353
R17080 VDD.n4304 VDD.n4201 0.0705353
R17081 VDD.n4562 VDD.n4459 0.0705353
R17082 VDD.n4820 VDD.n4717 0.0705353
R17083 VDD.n5078 VDD.n4975 0.0705353
R17084 VDD.n5336 VDD.n5233 0.0705353
R17085 VDD.n1846 VDD.n1845 0.0694784
R17086 VDD.n1849 VDD.n1846 0.0694784
R17087 VDD.n2167 VDD.n2166 0.0694784
R17088 VDD.n2170 VDD.n2167 0.0694784
R17089 VDD.n2425 VDD.n2424 0.0694784
R17090 VDD.n2428 VDD.n2425 0.0694784
R17091 VDD.n2683 VDD.n2682 0.0694784
R17092 VDD.n2686 VDD.n2683 0.0694784
R17093 VDD.n2941 VDD.n2940 0.0694784
R17094 VDD.n2944 VDD.n2941 0.0694784
R17095 VDD.n3199 VDD.n3198 0.0694784
R17096 VDD.n3202 VDD.n3199 0.0694784
R17097 VDD.n3457 VDD.n3456 0.0694784
R17098 VDD.n3460 VDD.n3457 0.0694784
R17099 VDD.n5777 VDD.n5776 0.0694784
R17100 VDD.n5780 VDD.n5777 0.0694784
R17101 VDD.n5523 VDD.n5522 0.0694784
R17102 VDD.n5526 VDD.n5523 0.0694784
R17103 VDD.n3715 VDD.n3714 0.0694784
R17104 VDD.n3718 VDD.n3715 0.0694784
R17105 VDD.n3973 VDD.n3972 0.0694784
R17106 VDD.n3976 VDD.n3973 0.0694784
R17107 VDD.n4231 VDD.n4230 0.0694784
R17108 VDD.n4234 VDD.n4231 0.0694784
R17109 VDD.n4489 VDD.n4488 0.0694784
R17110 VDD.n4492 VDD.n4489 0.0694784
R17111 VDD.n4747 VDD.n4746 0.0694784
R17112 VDD.n4750 VDD.n4747 0.0694784
R17113 VDD.n5005 VDD.n5004 0.0694784
R17114 VDD.n5008 VDD.n5005 0.0694784
R17115 VDD.n5263 VDD.n5262 0.0694784
R17116 VDD.n5266 VDD.n5263 0.0694784
R17117 VDD.n458 VDD.n457 0.0681471
R17118 VDD.n457 VDD.n454 0.0681471
R17119 VDD.n454 VDD.n451 0.0681471
R17120 VDD.n451 VDD.n450 0.0681471
R17121 VDD.n450 VDD.n447 0.0681471
R17122 VDD.n55 VDD.n54 0.0681471
R17123 VDD.n54 VDD.n51 0.0681471
R17124 VDD.n51 VDD.n48 0.0681471
R17125 VDD.n48 VDD.n47 0.0681471
R17126 VDD.n47 VDD.n44 0.0681471
R17127 VDD.n406 VDD.n403 0.0671334
R17128 VDD.n1564 VDD.n1561 0.0671334
R17129 VDD.n22 VDD.n21 0.065907
R17130 VDD.n17 VDD.n4 0.065907
R17131 VDD.n16 VDD.n15 0.065907
R17132 VDD.n14 VDD.n10 0.065907
R17133 VDD.n1166 VDD.n1165 0.065907
R17134 VDD.n1161 VDD.n1148 0.065907
R17135 VDD.n1160 VDD.n1159 0.065907
R17136 VDD.n1158 VDD.n1154 0.065907
R17137 VDD.n480 VDD.n479 0.0658409
R17138 VDD.n78 VDD.n77 0.0658409
R17139 VDD.n5739 VDD 0.0644514
R17140 VDD.n5485 VDD 0.0644514
R17141 VDD.n1791 VDD.n1783 0.0643889
R17142 VDD.n1791 VDD.n1780 0.0643889
R17143 VDD.n1796 VDD.n1780 0.0643889
R17144 VDD.n1999 VDD.n1991 0.0643889
R17145 VDD.n1999 VDD.n1988 0.0643889
R17146 VDD.n2004 VDD.n1988 0.0643889
R17147 VDD.n2370 VDD.n2362 0.0643889
R17148 VDD.n2370 VDD.n2359 0.0643889
R17149 VDD.n2375 VDD.n2359 0.0643889
R17150 VDD.n2628 VDD.n2620 0.0643889
R17151 VDD.n2628 VDD.n2617 0.0643889
R17152 VDD.n2633 VDD.n2617 0.0643889
R17153 VDD.n2886 VDD.n2878 0.0643889
R17154 VDD.n2886 VDD.n2875 0.0643889
R17155 VDD.n2891 VDD.n2875 0.0643889
R17156 VDD.n3144 VDD.n3136 0.0643889
R17157 VDD.n3144 VDD.n3133 0.0643889
R17158 VDD.n3149 VDD.n3133 0.0643889
R17159 VDD.n3402 VDD.n3394 0.0643889
R17160 VDD.n3402 VDD.n3391 0.0643889
R17161 VDD.n3407 VDD.n3391 0.0643889
R17162 VDD.n5725 VDD.n5717 0.0643889
R17163 VDD.n5725 VDD.n5714 0.0643889
R17164 VDD.n5730 VDD.n5714 0.0643889
R17165 VDD.n5471 VDD.n5463 0.0643889
R17166 VDD.n5471 VDD.n5460 0.0643889
R17167 VDD.n5476 VDD.n5460 0.0643889
R17168 VDD.n3660 VDD.n3652 0.0643889
R17169 VDD.n3660 VDD.n3649 0.0643889
R17170 VDD.n3665 VDD.n3649 0.0643889
R17171 VDD.n3918 VDD.n3910 0.0643889
R17172 VDD.n3918 VDD.n3907 0.0643889
R17173 VDD.n3923 VDD.n3907 0.0643889
R17174 VDD.n4176 VDD.n4168 0.0643889
R17175 VDD.n4176 VDD.n4165 0.0643889
R17176 VDD.n4181 VDD.n4165 0.0643889
R17177 VDD.n4434 VDD.n4426 0.0643889
R17178 VDD.n4434 VDD.n4423 0.0643889
R17179 VDD.n4439 VDD.n4423 0.0643889
R17180 VDD.n4692 VDD.n4684 0.0643889
R17181 VDD.n4692 VDD.n4681 0.0643889
R17182 VDD.n4697 VDD.n4681 0.0643889
R17183 VDD.n4950 VDD.n4942 0.0643889
R17184 VDD.n4950 VDD.n4939 0.0643889
R17185 VDD.n4955 VDD.n4939 0.0643889
R17186 VDD.n5208 VDD.n5200 0.0643889
R17187 VDD.n5208 VDD.n5197 0.0643889
R17188 VDD.n5213 VDD.n5197 0.0643889
R17189 VDD.n507 VDD.n505 0.0643889
R17190 VDD.n505 VDD.n503 0.0643889
R17191 VDD.n503 VDD.n501 0.0643889
R17192 VDD.n498 VDD.n497 0.0643889
R17193 VDD.n497 VDD.n493 0.0643889
R17194 VDD.n493 VDD.n491 0.0643889
R17195 VDD.n486 VDD.n485 0.0643889
R17196 VDD.n434 VDD.n432 0.0643889
R17197 VDD.n432 VDD.n430 0.0643889
R17198 VDD.n430 VDD.n428 0.0643889
R17199 VDD.n421 VDD.n417 0.0643889
R17200 VDD.n417 VDD.n415 0.0643889
R17201 VDD.n415 VDD.n413 0.0643889
R17202 VDD.n400 VDD.n398 0.0643889
R17203 VDD.n398 VDD.n396 0.0643889
R17204 VDD.n105 VDD.n103 0.0643889
R17205 VDD.n103 VDD.n101 0.0643889
R17206 VDD.n101 VDD.n99 0.0643889
R17207 VDD.n96 VDD.n95 0.0643889
R17208 VDD.n95 VDD.n91 0.0643889
R17209 VDD.n91 VDD.n89 0.0643889
R17210 VDD.n84 VDD.n83 0.0643889
R17211 VDD.n1592 VDD.n1590 0.0643889
R17212 VDD.n1590 VDD.n1588 0.0643889
R17213 VDD.n1588 VDD.n1586 0.0643889
R17214 VDD.n1579 VDD.n1575 0.0643889
R17215 VDD.n1575 VDD.n1573 0.0643889
R17216 VDD.n1573 VDD.n1571 0.0643889
R17217 VDD.n1558 VDD.n1556 0.0643889
R17218 VDD.n1556 VDD.n1554 0.0643889
R17219 VDD.n1526 VDD 0.0639804
R17220 VDD.n1806 VDD 0.0630006
R17221 VDD.n2126 VDD 0.0630006
R17222 VDD.n2385 VDD 0.0630006
R17223 VDD.n2643 VDD 0.0630006
R17224 VDD.n2901 VDD 0.0630006
R17225 VDD.n3159 VDD 0.0630006
R17226 VDD.n3417 VDD 0.0630006
R17227 VDD.n3675 VDD 0.0630006
R17228 VDD.n3933 VDD 0.0630006
R17229 VDD.n4191 VDD 0.0630006
R17230 VDD.n4449 VDD 0.0630006
R17231 VDD.n4707 VDD 0.0630006
R17232 VDD.n4965 VDD 0.0630006
R17233 VDD.n5223 VDD 0.0630006
R17234 VDD.n1623 VDD 0.0604792
R17235 VDD.n462 VDD.n461 0.0599867
R17236 VDD.n59 VDD.n58 0.0599867
R17237 VDD.n1772 VDD.n1667 0.0588333
R17238 VDD.n2121 VDD.n2016 0.0588333
R17239 VDD.n2351 VDD.n2246 0.0588333
R17240 VDD.n2609 VDD.n2504 0.0588333
R17241 VDD.n2867 VDD.n2762 0.0588333
R17242 VDD.n3125 VDD.n3020 0.0588333
R17243 VDD.n3383 VDD.n3278 0.0588333
R17244 VDD.n5706 VDD.n5601 0.0588333
R17245 VDD.n5452 VDD.n5347 0.0588333
R17246 VDD.n3641 VDD.n3536 0.0588333
R17247 VDD.n3899 VDD.n3794 0.0588333
R17248 VDD.n4157 VDD.n4052 0.0588333
R17249 VDD.n4415 VDD.n4310 0.0588333
R17250 VDD.n4673 VDD.n4568 0.0588333
R17251 VDD.n4931 VDD.n4826 0.0588333
R17252 VDD.n5189 VDD.n5084 0.0588333
R17253 VDD.n395 VDD.n394 0.0587674
R17254 VDD.n1553 VDD.n1552 0.0587674
R17255 VDD.n425 VDD.n424 0.0580441
R17256 VDD.n1583 VDD.n1582 0.0580441
R17257 VDD.n848 VDD 0.058
R17258 VDD.n842 VDD 0.058
R17259 VDD.n830 VDD 0.058
R17260 VDD.n1231 VDD 0.058
R17261 VDD.n1225 VDD 0.058
R17262 VDD.n1213 VDD 0.058
R17263 VDD.n491 VDD.n489 0.0567153
R17264 VDD.n89 VDD.n87 0.0567153
R17265 VDD.n5863 VDD.n5862 0.0560833
R17266 VDD.n836 VDD 0.0555
R17267 VDD.n1219 VDD 0.0555
R17268 VDD.n5852 VDD.n5851 0.0554144
R17269 VDD.n5598 VDD.n5597 0.0554144
R17270 VDD VDD.n5860 0.0546184
R17271 VDD VDD.n1783 0.0525833
R17272 VDD VDD.n1991 0.0525833
R17273 VDD VDD.n2362 0.0525833
R17274 VDD VDD.n2620 0.0525833
R17275 VDD VDD.n2878 0.0525833
R17276 VDD VDD.n3136 0.0525833
R17277 VDD VDD.n3394 0.0525833
R17278 VDD VDD.n5717 0.0525833
R17279 VDD VDD.n5463 0.0525833
R17280 VDD VDD.n3652 0.0525833
R17281 VDD VDD.n3910 0.0525833
R17282 VDD VDD.n4168 0.0525833
R17283 VDD VDD.n4426 0.0525833
R17284 VDD VDD.n4684 0.0525833
R17285 VDD VDD.n4942 0.0525833
R17286 VDD VDD.n5200 0.0525833
R17287 VDD.n481 VDD.n480 0.0516364
R17288 VDD.n79 VDD.n78 0.0516364
R17289 VDD.n1799 VDD 0.0470278
R17290 VDD.n2007 VDD 0.0470278
R17291 VDD.n2378 VDD 0.0470278
R17292 VDD.n2636 VDD 0.0470278
R17293 VDD.n2894 VDD 0.0470278
R17294 VDD.n3152 VDD 0.0470278
R17295 VDD.n3410 VDD 0.0470278
R17296 VDD.n5733 VDD 0.0470278
R17297 VDD.n5479 VDD 0.0470278
R17298 VDD.n3668 VDD 0.0470278
R17299 VDD.n3926 VDD 0.0470278
R17300 VDD.n4184 VDD 0.0470278
R17301 VDD.n4442 VDD 0.0470278
R17302 VDD.n4700 VDD 0.0470278
R17303 VDD.n4958 VDD 0.0470278
R17304 VDD.n5216 VDD 0.0470278
R17305 VDD.n5852 VDD.n5598 0.0430009
R17306 VDD.n5853 VDD.n5852 0.0425691
R17307 VDD.n5598 VDD.n5344 0.0421424
R17308 VDD.n25 VDD.n0 0.0418891
R17309 VDD.n1169 VDD.n1144 0.0418891
R17310 VDD.n5858 VDD.n5857 0.0417105
R17311 VDD.n5857 VDD.n5856 0.0417105
R17312 VDD.n5856 VDD.n5855 0.0417105
R17313 VDD.n5855 VDD.n5854 0.0417105
R17314 VDD.n5854 VDD.n5853 0.0417105
R17315 VDD.n5344 VDD.n5343 0.0417105
R17316 VDD.n5343 VDD.n5342 0.0417105
R17317 VDD.n5342 VDD.n5341 0.0417105
R17318 VDD.n5341 VDD.n5340 0.0417105
R17319 VDD.n5340 VDD.n5339 0.0417105
R17320 VDD.n1832 VDD.n1831 0.0409412
R17321 VDD.n2153 VDD.n2152 0.0409412
R17322 VDD.n2411 VDD.n2410 0.0409412
R17323 VDD.n2669 VDD.n2668 0.0409412
R17324 VDD.n2927 VDD.n2926 0.0409412
R17325 VDD.n3185 VDD.n3184 0.0409412
R17326 VDD.n3443 VDD.n3442 0.0409412
R17327 VDD.n5763 VDD.n5762 0.0409412
R17328 VDD.n5509 VDD.n5508 0.0409412
R17329 VDD.n3701 VDD.n3700 0.0409412
R17330 VDD.n3959 VDD.n3958 0.0409412
R17331 VDD.n4217 VDD.n4216 0.0409412
R17332 VDD.n4475 VDD.n4474 0.0409412
R17333 VDD.n4733 VDD.n4732 0.0409412
R17334 VDD.n4991 VDD.n4990 0.0409412
R17335 VDD.n5249 VDD.n5248 0.0409412
R17336 VDD.n30 VDD.n28 0.0409412
R17337 VDD.n1174 VDD.n1172 0.0409412
R17338 VDD.n5709 VDD.n5708 0.0399318
R17339 VDD.n5455 VDD.n5454 0.0399318
R17340 VDD.n5860 VDD.n5859 0.0398026
R17341 VDD.n820 VDD.n799 0.03976
R17342 VDD.n1203 VDD.n1182 0.03976
R17343 VDD.n1797 VDD.n1776 0.0395625
R17344 VDD.n2005 VDD.n1984 0.0395625
R17345 VDD.n2376 VDD.n2355 0.0395625
R17346 VDD.n2634 VDD.n2613 0.0395625
R17347 VDD.n2892 VDD.n2871 0.0395625
R17348 VDD.n3150 VDD.n3129 0.0395625
R17349 VDD.n3408 VDD.n3387 0.0395625
R17350 VDD.n5731 VDD.n5710 0.0395625
R17351 VDD.n5477 VDD.n5456 0.0395625
R17352 VDD.n3666 VDD.n3645 0.0395625
R17353 VDD.n3924 VDD.n3903 0.0395625
R17354 VDD.n4182 VDD.n4161 0.0395625
R17355 VDD.n4440 VDD.n4419 0.0395625
R17356 VDD.n4698 VDD.n4677 0.0395625
R17357 VDD.n4956 VDD.n4935 0.0395625
R17358 VDD.n5214 VDD.n5193 0.0395625
R17359 VDD.n797 VDD 0.0390887
R17360 VDD.n854 VDD.n853 0.0376094
R17361 VDD.n1237 VDD.n1236 0.0376094
R17362 VDD.n1836 VDD.n1835 0.0372647
R17363 VDD.n2157 VDD.n2156 0.0372647
R17364 VDD.n2415 VDD.n2414 0.0372647
R17365 VDD.n2673 VDD.n2672 0.0372647
R17366 VDD.n2931 VDD.n2930 0.0372647
R17367 VDD.n3189 VDD.n3188 0.0372647
R17368 VDD.n3447 VDD.n3446 0.0372647
R17369 VDD.n5767 VDD.n5766 0.0372647
R17370 VDD.n5513 VDD.n5512 0.0372647
R17371 VDD.n3705 VDD.n3704 0.0372647
R17372 VDD.n3963 VDD.n3962 0.0372647
R17373 VDD.n4221 VDD.n4220 0.0372647
R17374 VDD.n4479 VDD.n4478 0.0372647
R17375 VDD.n4737 VDD.n4736 0.0372647
R17376 VDD.n4995 VDD.n4994 0.0372647
R17377 VDD.n5253 VDD.n5252 0.0372647
R17378 VDD.n28 VDD.n27 0.0371297
R17379 VDD.n1172 VDD.n1171 0.0371297
R17380 VDD.n1701 VDD.n1665 0.0364409
R17381 VDD.n2050 VDD.n2014 0.0364409
R17382 VDD.n2280 VDD.n2244 0.0364409
R17383 VDD.n2538 VDD.n2502 0.0364409
R17384 VDD.n2796 VDD.n2760 0.0364409
R17385 VDD.n3054 VDD.n3018 0.0364409
R17386 VDD.n3312 VDD.n3276 0.0364409
R17387 VDD.n5635 VDD.n5599 0.0364409
R17388 VDD.n5381 VDD.n5345 0.0364409
R17389 VDD.n3570 VDD.n3534 0.0364409
R17390 VDD.n3828 VDD.n3792 0.0364409
R17391 VDD.n4086 VDD.n4050 0.0364409
R17392 VDD.n4344 VDD.n4308 0.0364409
R17393 VDD.n4602 VDD.n4566 0.0364409
R17394 VDD.n4860 VDD.n4824 0.0364409
R17395 VDD.n5118 VDD.n5082 0.0364409
R17396 VDD.n1837 VDD.n1836 0.0361152
R17397 VDD.n2158 VDD.n2157 0.0361152
R17398 VDD.n2416 VDD.n2415 0.0361152
R17399 VDD.n2674 VDD.n2673 0.0361152
R17400 VDD.n2932 VDD.n2931 0.0361152
R17401 VDD.n3190 VDD.n3189 0.0361152
R17402 VDD.n3448 VDD.n3447 0.0361152
R17403 VDD.n5768 VDD.n5767 0.0361152
R17404 VDD.n5514 VDD.n5513 0.0361152
R17405 VDD.n3706 VDD.n3705 0.0361152
R17406 VDD.n3964 VDD.n3963 0.0361152
R17407 VDD.n4222 VDD.n4221 0.0361152
R17408 VDD.n4480 VDD.n4479 0.0361152
R17409 VDD.n4738 VDD.n4737 0.0361152
R17410 VDD.n4996 VDD.n4995 0.0361152
R17411 VDD.n5254 VDD.n5253 0.0361152
R17412 VDD.n1752 VDD.n1751 0.0357224
R17413 VDD.n2101 VDD.n2100 0.0357224
R17414 VDD.n2331 VDD.n2330 0.0357224
R17415 VDD.n2589 VDD.n2588 0.0357224
R17416 VDD.n2847 VDD.n2846 0.0357224
R17417 VDD.n3105 VDD.n3104 0.0357224
R17418 VDD.n3363 VDD.n3362 0.0357224
R17419 VDD.n5686 VDD.n5685 0.0357224
R17420 VDD.n5432 VDD.n5431 0.0357224
R17421 VDD.n3621 VDD.n3620 0.0357224
R17422 VDD.n3879 VDD.n3878 0.0357224
R17423 VDD.n4137 VDD.n4136 0.0357224
R17424 VDD.n4395 VDD.n4394 0.0357224
R17425 VDD.n4653 VDD.n4652 0.0357224
R17426 VDD.n4911 VDD.n4910 0.0357224
R17427 VDD.n5169 VDD.n5168 0.0357224
R17428 VDD.n1684 VDD.n1683 0.034445
R17429 VDD.n2033 VDD.n2032 0.034445
R17430 VDD.n2263 VDD.n2262 0.034445
R17431 VDD.n2521 VDD.n2520 0.034445
R17432 VDD.n2779 VDD.n2778 0.034445
R17433 VDD.n3037 VDD.n3036 0.034445
R17434 VDD.n3295 VDD.n3294 0.034445
R17435 VDD.n5618 VDD.n5617 0.034445
R17436 VDD.n5364 VDD.n5363 0.034445
R17437 VDD.n3553 VDD.n3552 0.034445
R17438 VDD.n3811 VDD.n3810 0.034445
R17439 VDD.n4069 VDD.n4068 0.034445
R17440 VDD.n4327 VDD.n4326 0.034445
R17441 VDD.n4585 VDD.n4584 0.034445
R17442 VDD.n4843 VDD.n4842 0.034445
R17443 VDD.n5101 VDD.n5100 0.034445
R17444 VDD.n3 VDD.n0 0.0339302
R17445 VDD.n1147 VDD.n1144 0.0339302
R17446 VDD.n810 VDD.n802 0.033737
R17447 VDD.n814 VDD.n802 0.033737
R17448 VDD.n815 VDD.n814 0.033737
R17449 VDD.n816 VDD.n815 0.033737
R17450 VDD.n1193 VDD.n1185 0.033737
R17451 VDD.n1197 VDD.n1185 0.033737
R17452 VDD.n1198 VDD.n1197 0.033737
R17453 VDD.n1199 VDD.n1198 0.033737
R17454 VDD.n479 VDD.n477 0.0334425
R17455 VDD.n477 VDD.n474 0.0334425
R17456 VDD.n77 VDD.n75 0.0334425
R17457 VDD.n75 VDD.n72 0.0334425
R17458 VDD.n1548 VDD.n1547 0.0333707
R17459 VDD.n863 VDD.n798 0.0325611
R17460 VDD VDD.n1796 0.0324444
R17461 VDD VDD.n2004 0.0324444
R17462 VDD VDD.n2375 0.0324444
R17463 VDD VDD.n2633 0.0324444
R17464 VDD VDD.n2891 0.0324444
R17465 VDD VDD.n3149 0.0324444
R17466 VDD VDD.n3407 0.0324444
R17467 VDD VDD.n5730 0.0324444
R17468 VDD VDD.n5476 0.0324444
R17469 VDD VDD.n3665 0.0324444
R17470 VDD VDD.n3923 0.0324444
R17471 VDD VDD.n4181 0.0324444
R17472 VDD VDD.n4439 0.0324444
R17473 VDD VDD.n4697 0.0324444
R17474 VDD VDD.n4955 0.0324444
R17475 VDD VDD.n5213 0.0324444
R17476 VDD.n498 VDD 0.0324444
R17477 VDD.n486 VDD 0.0324444
R17478 VDD.n425 VDD 0.0324444
R17479 VDD.n96 VDD 0.0324444
R17480 VDD.n84 VDD 0.0324444
R17481 VDD.n1583 VDD 0.0324444
R17482 VDD.n1640 VDD.n1639 0.0308571
R17483 VDD.n110 VDD.n62 0.0299677
R17484 VDD.n798 VDD.n110 0.0299677
R17485 VDD.n513 VDD.n512 0.0299677
R17486 VDD.n1771 VDD.n1770 0.0294474
R17487 VDD.n2120 VDD.n2119 0.0294474
R17488 VDD.n2350 VDD.n2349 0.0294474
R17489 VDD.n2608 VDD.n2607 0.0294474
R17490 VDD.n2866 VDD.n2865 0.0294474
R17491 VDD.n3124 VDD.n3123 0.0294474
R17492 VDD.n3382 VDD.n3381 0.0294474
R17493 VDD.n5705 VDD.n5704 0.0294474
R17494 VDD.n5451 VDD.n5450 0.0294474
R17495 VDD.n3640 VDD.n3639 0.0294474
R17496 VDD.n3898 VDD.n3897 0.0294474
R17497 VDD.n4156 VDD.n4155 0.0294474
R17498 VDD.n4414 VDD.n4413 0.0294474
R17499 VDD.n4672 VDD.n4671 0.0294474
R17500 VDD.n4930 VDD.n4929 0.0294474
R17501 VDD.n5188 VDD.n5187 0.0294474
R17502 VDD.n1598 VDD.n1597 0.0292661
R17503 VDD.n796 VDD.n795 0.0292661
R17504 VDD.n1754 VDD.n1753 0.0287895
R17505 VDD.n2103 VDD.n2102 0.0287895
R17506 VDD.n2333 VDD.n2332 0.0287895
R17507 VDD.n2591 VDD.n2590 0.0287895
R17508 VDD.n2849 VDD.n2848 0.0287895
R17509 VDD.n3107 VDD.n3106 0.0287895
R17510 VDD.n3365 VDD.n3364 0.0287895
R17511 VDD.n5688 VDD.n5687 0.0287895
R17512 VDD.n5434 VDD.n5433 0.0287895
R17513 VDD.n3623 VDD.n3622 0.0287895
R17514 VDD.n3881 VDD.n3880 0.0287895
R17515 VDD.n4139 VDD.n4138 0.0287895
R17516 VDD.n4397 VDD.n4396 0.0287895
R17517 VDD.n4655 VDD.n4654 0.0287895
R17518 VDD.n4913 VDD.n4912 0.0287895
R17519 VDD.n5171 VDD.n5170 0.0287895
R17520 VDD.n1750 VDD.n1720 0.0282778
R17521 VDD.n2099 VDD.n2069 0.0282778
R17522 VDD.n2329 VDD.n2299 0.0282778
R17523 VDD.n2587 VDD.n2557 0.0282778
R17524 VDD.n2845 VDD.n2815 0.0282778
R17525 VDD.n3103 VDD.n3073 0.0282778
R17526 VDD.n3361 VDD.n3331 0.0282778
R17527 VDD.n5684 VDD.n5654 0.0282778
R17528 VDD.n5430 VDD.n5400 0.0282778
R17529 VDD.n3619 VDD.n3589 0.0282778
R17530 VDD.n3877 VDD.n3847 0.0282778
R17531 VDD.n4135 VDD.n4105 0.0282778
R17532 VDD.n4393 VDD.n4363 0.0282778
R17533 VDD.n4651 VDD.n4621 0.0282778
R17534 VDD.n4909 VDD.n4879 0.0282778
R17535 VDD.n5167 VDD.n5137 0.0282778
R17536 VDD.t388 VDD.n1763 0.0282694
R17537 VDD.n1763 VDD.n1762 0.0282694
R17538 VDD.t388 VDD.n1677 0.0282694
R17539 VDD.n1706 VDD.n1677 0.0282694
R17540 VDD.t228 VDD.n2112 0.0282694
R17541 VDD.n2112 VDD.n2111 0.0282694
R17542 VDD.t228 VDD.n2026 0.0282694
R17543 VDD.n2055 VDD.n2026 0.0282694
R17544 VDD.t181 VDD.n2342 0.0282694
R17545 VDD.n2342 VDD.n2341 0.0282694
R17546 VDD.t181 VDD.n2256 0.0282694
R17547 VDD.n2285 VDD.n2256 0.0282694
R17548 VDD.t713 VDD.n2600 0.0282694
R17549 VDD.n2600 VDD.n2599 0.0282694
R17550 VDD.t713 VDD.n2514 0.0282694
R17551 VDD.n2543 VDD.n2514 0.0282694
R17552 VDD.t542 VDD.n2858 0.0282694
R17553 VDD.n2858 VDD.n2857 0.0282694
R17554 VDD.t542 VDD.n2772 0.0282694
R17555 VDD.n2801 VDD.n2772 0.0282694
R17556 VDD.t647 VDD.n3116 0.0282694
R17557 VDD.n3116 VDD.n3115 0.0282694
R17558 VDD.t647 VDD.n3030 0.0282694
R17559 VDD.n3059 VDD.n3030 0.0282694
R17560 VDD.t30 VDD.n3374 0.0282694
R17561 VDD.n3374 VDD.n3373 0.0282694
R17562 VDD.t30 VDD.n3288 0.0282694
R17563 VDD.n3317 VDD.n3288 0.0282694
R17564 VDD.t870 VDD.n5697 0.0282694
R17565 VDD.n5697 VDD.n5696 0.0282694
R17566 VDD.t870 VDD.n5611 0.0282694
R17567 VDD.n5640 VDD.n5611 0.0282694
R17568 VDD.t709 VDD.n5443 0.0282694
R17569 VDD.n5443 VDD.n5442 0.0282694
R17570 VDD.t709 VDD.n5357 0.0282694
R17571 VDD.n5386 VDD.n5357 0.0282694
R17572 VDD.t214 VDD.n3632 0.0282694
R17573 VDD.n3632 VDD.n3631 0.0282694
R17574 VDD.t214 VDD.n3546 0.0282694
R17575 VDD.n3575 VDD.n3546 0.0282694
R17576 VDD.t1027 VDD.n3890 0.0282694
R17577 VDD.n3890 VDD.n3889 0.0282694
R17578 VDD.t1027 VDD.n3804 0.0282694
R17579 VDD.n3833 VDD.n3804 0.0282694
R17580 VDD.t423 VDD.n4148 0.0282694
R17581 VDD.n4148 VDD.n4147 0.0282694
R17582 VDD.t423 VDD.n4062 0.0282694
R17583 VDD.n4091 VDD.n4062 0.0282694
R17584 VDD.t1031 VDD.n4406 0.0282694
R17585 VDD.n4406 VDD.n4405 0.0282694
R17586 VDD.t1031 VDD.n4320 0.0282694
R17587 VDD.n4349 VDD.n4320 0.0282694
R17588 VDD.t402 VDD.n4664 0.0282694
R17589 VDD.n4664 VDD.n4663 0.0282694
R17590 VDD.t402 VDD.n4578 0.0282694
R17591 VDD.n4607 VDD.n4578 0.0282694
R17592 VDD.t532 VDD.n4922 0.0282694
R17593 VDD.n4922 VDD.n4921 0.0282694
R17594 VDD.t532 VDD.n4836 0.0282694
R17595 VDD.n4865 VDD.n4836 0.0282694
R17596 VDD.t381 VDD.n5180 0.0282694
R17597 VDD.n5180 VDD.n5179 0.0282694
R17598 VDD.t381 VDD.n5094 0.0282694
R17599 VDD.n5123 VDD.n5094 0.0282694
R17600 VDD.n674 VDD 0.0279106
R17601 VDD.n1024 VDD 0.0279106
R17602 VDD.n269 VDD 0.0279106
R17603 VDD.n1897 VDD.n1895 0.0265784
R17604 VDD.n1905 VDD.n1895 0.0265784
R17605 VDD.n1911 VDD.n1896 0.0265784
R17606 VDD.n1901 VDD.n1896 0.0265784
R17607 VDD.n1903 VDD.n1902 0.0265784
R17608 VDD.n1902 VDD.n1901 0.0265784
R17609 VDD.n1907 VDD.n1906 0.0265784
R17610 VDD.n1906 VDD.n1905 0.0265784
R17611 VDD.n1878 VDD.n1877 0.0265784
R17612 VDD.t528 VDD.n1878 0.0265784
R17613 VDD.n1880 VDD.n1822 0.0265784
R17614 VDD.n1860 VDD.n1859 0.0265784
R17615 VDD.n1859 VDD.n1858 0.0265784
R17616 VDD.n1862 VDD.n1853 0.0265784
R17617 VDD.n1863 VDD.n1862 0.0265784
R17618 VDD.n1865 VDD.n1864 0.0265784
R17619 VDD.n1864 VDD.n1863 0.0265784
R17620 VDD.n1858 VDD.n1855 0.0265784
R17621 VDD.n1855 VDD.n1854 0.0265784
R17622 VDD.n2181 VDD.n2180 0.0265784
R17623 VDD.n2180 VDD.n2179 0.0265784
R17624 VDD.n2183 VDD.n2174 0.0265784
R17625 VDD.n2184 VDD.n2183 0.0265784
R17626 VDD.n2186 VDD.n2185 0.0265784
R17627 VDD.n2185 VDD.n2184 0.0265784
R17628 VDD.n2179 VDD.n2176 0.0265784
R17629 VDD.n2176 VDD.n2175 0.0265784
R17630 VDD.n2199 VDD.n2198 0.0265784
R17631 VDD.t481 VDD.n2199 0.0265784
R17632 VDD.n2201 VDD.n2143 0.0265784
R17633 VDD.n2218 VDD.n2216 0.0265784
R17634 VDD.n2226 VDD.n2216 0.0265784
R17635 VDD.n2232 VDD.n2217 0.0265784
R17636 VDD.n2222 VDD.n2217 0.0265784
R17637 VDD.n2224 VDD.n2223 0.0265784
R17638 VDD.n2223 VDD.n2222 0.0265784
R17639 VDD.n2228 VDD.n2227 0.0265784
R17640 VDD.n2227 VDD.n2226 0.0265784
R17641 VDD.n2439 VDD.n2438 0.0265784
R17642 VDD.n2438 VDD.n2437 0.0265784
R17643 VDD.n2441 VDD.n2432 0.0265784
R17644 VDD.n2442 VDD.n2441 0.0265784
R17645 VDD.n2444 VDD.n2443 0.0265784
R17646 VDD.n2443 VDD.n2442 0.0265784
R17647 VDD.n2437 VDD.n2434 0.0265784
R17648 VDD.n2434 VDD.n2433 0.0265784
R17649 VDD.n2457 VDD.n2456 0.0265784
R17650 VDD.t118 VDD.n2457 0.0265784
R17651 VDD.n2459 VDD.n2401 0.0265784
R17652 VDD.n2476 VDD.n2474 0.0265784
R17653 VDD.n2484 VDD.n2474 0.0265784
R17654 VDD.n2490 VDD.n2475 0.0265784
R17655 VDD.n2480 VDD.n2475 0.0265784
R17656 VDD.n2482 VDD.n2481 0.0265784
R17657 VDD.n2481 VDD.n2480 0.0265784
R17658 VDD.n2486 VDD.n2485 0.0265784
R17659 VDD.n2485 VDD.n2484 0.0265784
R17660 VDD.n2697 VDD.n2696 0.0265784
R17661 VDD.n2696 VDD.n2695 0.0265784
R17662 VDD.n2699 VDD.n2690 0.0265784
R17663 VDD.n2700 VDD.n2699 0.0265784
R17664 VDD.n2702 VDD.n2701 0.0265784
R17665 VDD.n2701 VDD.n2700 0.0265784
R17666 VDD.n2695 VDD.n2692 0.0265784
R17667 VDD.n2692 VDD.n2691 0.0265784
R17668 VDD.n2715 VDD.n2714 0.0265784
R17669 VDD.t652 VDD.n2715 0.0265784
R17670 VDD.n2717 VDD.n2659 0.0265784
R17671 VDD.n2734 VDD.n2732 0.0265784
R17672 VDD.n2742 VDD.n2732 0.0265784
R17673 VDD.n2748 VDD.n2733 0.0265784
R17674 VDD.n2738 VDD.n2733 0.0265784
R17675 VDD.n2740 VDD.n2739 0.0265784
R17676 VDD.n2739 VDD.n2738 0.0265784
R17677 VDD.n2744 VDD.n2743 0.0265784
R17678 VDD.n2743 VDD.n2742 0.0265784
R17679 VDD.n2955 VDD.n2954 0.0265784
R17680 VDD.n2954 VDD.n2953 0.0265784
R17681 VDD.n2957 VDD.n2948 0.0265784
R17682 VDD.n2958 VDD.n2957 0.0265784
R17683 VDD.n2960 VDD.n2959 0.0265784
R17684 VDD.n2959 VDD.n2958 0.0265784
R17685 VDD.n2953 VDD.n2950 0.0265784
R17686 VDD.n2950 VDD.n2949 0.0265784
R17687 VDD.n2973 VDD.n2972 0.0265784
R17688 VDD.t12 VDD.n2973 0.0265784
R17689 VDD.n2975 VDD.n2917 0.0265784
R17690 VDD.n2992 VDD.n2990 0.0265784
R17691 VDD.n3000 VDD.n2990 0.0265784
R17692 VDD.n3006 VDD.n2991 0.0265784
R17693 VDD.n2996 VDD.n2991 0.0265784
R17694 VDD.n2998 VDD.n2997 0.0265784
R17695 VDD.n2997 VDD.n2996 0.0265784
R17696 VDD.n3002 VDD.n3001 0.0265784
R17697 VDD.n3001 VDD.n3000 0.0265784
R17698 VDD.n3213 VDD.n3212 0.0265784
R17699 VDD.n3212 VDD.n3211 0.0265784
R17700 VDD.n3215 VDD.n3206 0.0265784
R17701 VDD.n3216 VDD.n3215 0.0265784
R17702 VDD.n3218 VDD.n3217 0.0265784
R17703 VDD.n3217 VDD.n3216 0.0265784
R17704 VDD.n3211 VDD.n3208 0.0265784
R17705 VDD.n3208 VDD.n3207 0.0265784
R17706 VDD.n3231 VDD.n3230 0.0265784
R17707 VDD.t718 VDD.n3231 0.0265784
R17708 VDD.n3233 VDD.n3175 0.0265784
R17709 VDD.n3250 VDD.n3248 0.0265784
R17710 VDD.n3258 VDD.n3248 0.0265784
R17711 VDD.n3264 VDD.n3249 0.0265784
R17712 VDD.n3254 VDD.n3249 0.0265784
R17713 VDD.n3256 VDD.n3255 0.0265784
R17714 VDD.n3255 VDD.n3254 0.0265784
R17715 VDD.n3260 VDD.n3259 0.0265784
R17716 VDD.n3259 VDD.n3258 0.0265784
R17717 VDD.n3471 VDD.n3470 0.0265784
R17718 VDD.n3470 VDD.n3469 0.0265784
R17719 VDD.n3473 VDD.n3464 0.0265784
R17720 VDD.n3474 VDD.n3473 0.0265784
R17721 VDD.n3476 VDD.n3475 0.0265784
R17722 VDD.n3475 VDD.n3474 0.0265784
R17723 VDD.n3469 VDD.n3466 0.0265784
R17724 VDD.n3466 VDD.n3465 0.0265784
R17725 VDD.n3489 VDD.n3488 0.0265784
R17726 VDD.t411 VDD.n3489 0.0265784
R17727 VDD.n3491 VDD.n3433 0.0265784
R17728 VDD.n3508 VDD.n3506 0.0265784
R17729 VDD.n3516 VDD.n3506 0.0265784
R17730 VDD.n3522 VDD.n3507 0.0265784
R17731 VDD.n3512 VDD.n3507 0.0265784
R17732 VDD.n3514 VDD.n3513 0.0265784
R17733 VDD.n3513 VDD.n3512 0.0265784
R17734 VDD.n3518 VDD.n3517 0.0265784
R17735 VDD.n3517 VDD.n3516 0.0265784
R17736 VDD.n5791 VDD.n5790 0.0265784
R17737 VDD.n5790 VDD.n5789 0.0265784
R17738 VDD.n5793 VDD.n5784 0.0265784
R17739 VDD.n5794 VDD.n5793 0.0265784
R17740 VDD.n5796 VDD.n5795 0.0265784
R17741 VDD.n5795 VDD.n5794 0.0265784
R17742 VDD.n5789 VDD.n5786 0.0265784
R17743 VDD.n5786 VDD.n5785 0.0265784
R17744 VDD.n5809 VDD.n5808 0.0265784
R17745 VDD.t530 VDD.n5809 0.0265784
R17746 VDD.n5811 VDD.n5753 0.0265784
R17747 VDD.n5828 VDD.n5826 0.0265784
R17748 VDD.n5836 VDD.n5826 0.0265784
R17749 VDD.n5842 VDD.n5827 0.0265784
R17750 VDD.n5832 VDD.n5827 0.0265784
R17751 VDD.n5834 VDD.n5833 0.0265784
R17752 VDD.n5833 VDD.n5832 0.0265784
R17753 VDD.n5838 VDD.n5837 0.0265784
R17754 VDD.n5837 VDD.n5836 0.0265784
R17755 VDD.n5537 VDD.n5536 0.0265784
R17756 VDD.n5536 VDD.n5535 0.0265784
R17757 VDD.n5539 VDD.n5530 0.0265784
R17758 VDD.n5540 VDD.n5539 0.0265784
R17759 VDD.n5542 VDD.n5541 0.0265784
R17760 VDD.n5541 VDD.n5540 0.0265784
R17761 VDD.n5535 VDD.n5532 0.0265784
R17762 VDD.n5532 VDD.n5531 0.0265784
R17763 VDD.n5555 VDD.n5554 0.0265784
R17764 VDD.t482 VDD.n5555 0.0265784
R17765 VDD.n5557 VDD.n5499 0.0265784
R17766 VDD.n5574 VDD.n5572 0.0265784
R17767 VDD.n5582 VDD.n5572 0.0265784
R17768 VDD.n5588 VDD.n5573 0.0265784
R17769 VDD.n5578 VDD.n5573 0.0265784
R17770 VDD.n5580 VDD.n5579 0.0265784
R17771 VDD.n5579 VDD.n5578 0.0265784
R17772 VDD.n5584 VDD.n5583 0.0265784
R17773 VDD.n5583 VDD.n5582 0.0265784
R17774 VDD.n3729 VDD.n3728 0.0265784
R17775 VDD.n3728 VDD.n3727 0.0265784
R17776 VDD.n3731 VDD.n3722 0.0265784
R17777 VDD.n3732 VDD.n3731 0.0265784
R17778 VDD.n3734 VDD.n3733 0.0265784
R17779 VDD.n3733 VDD.n3732 0.0265784
R17780 VDD.n3727 VDD.n3724 0.0265784
R17781 VDD.n3724 VDD.n3723 0.0265784
R17782 VDD.n3747 VDD.n3746 0.0265784
R17783 VDD.t410 VDD.n3747 0.0265784
R17784 VDD.n3749 VDD.n3691 0.0265784
R17785 VDD.n3766 VDD.n3764 0.0265784
R17786 VDD.n3774 VDD.n3764 0.0265784
R17787 VDD.n3780 VDD.n3765 0.0265784
R17788 VDD.n3770 VDD.n3765 0.0265784
R17789 VDD.n3772 VDD.n3771 0.0265784
R17790 VDD.n3771 VDD.n3770 0.0265784
R17791 VDD.n3776 VDD.n3775 0.0265784
R17792 VDD.n3775 VDD.n3774 0.0265784
R17793 VDD.n3987 VDD.n3986 0.0265784
R17794 VDD.n3986 VDD.n3985 0.0265784
R17795 VDD.n3989 VDD.n3980 0.0265784
R17796 VDD.n3990 VDD.n3989 0.0265784
R17797 VDD.n3992 VDD.n3991 0.0265784
R17798 VDD.n3991 VDD.n3990 0.0265784
R17799 VDD.n3985 VDD.n3982 0.0265784
R17800 VDD.n3982 VDD.n3981 0.0265784
R17801 VDD.n4005 VDD.n4004 0.0265784
R17802 VDD.t116 VDD.n4005 0.0265784
R17803 VDD.n4007 VDD.n3949 0.0265784
R17804 VDD.n4024 VDD.n4022 0.0265784
R17805 VDD.n4032 VDD.n4022 0.0265784
R17806 VDD.n4038 VDD.n4023 0.0265784
R17807 VDD.n4028 VDD.n4023 0.0265784
R17808 VDD.n4030 VDD.n4029 0.0265784
R17809 VDD.n4029 VDD.n4028 0.0265784
R17810 VDD.n4034 VDD.n4033 0.0265784
R17811 VDD.n4033 VDD.n4032 0.0265784
R17812 VDD.n4245 VDD.n4244 0.0265784
R17813 VDD.n4244 VDD.n4243 0.0265784
R17814 VDD.n4247 VDD.n4238 0.0265784
R17815 VDD.n4248 VDD.n4247 0.0265784
R17816 VDD.n4250 VDD.n4249 0.0265784
R17817 VDD.n4249 VDD.n4248 0.0265784
R17818 VDD.n4243 VDD.n4240 0.0265784
R17819 VDD.n4240 VDD.n4239 0.0265784
R17820 VDD.n4263 VDD.n4262 0.0265784
R17821 VDD.t489 VDD.n4263 0.0265784
R17822 VDD.n4265 VDD.n4207 0.0265784
R17823 VDD.n4282 VDD.n4280 0.0265784
R17824 VDD.n4290 VDD.n4280 0.0265784
R17825 VDD.n4296 VDD.n4281 0.0265784
R17826 VDD.n4286 VDD.n4281 0.0265784
R17827 VDD.n4288 VDD.n4287 0.0265784
R17828 VDD.n4287 VDD.n4286 0.0265784
R17829 VDD.n4292 VDD.n4291 0.0265784
R17830 VDD.n4291 VDD.n4290 0.0265784
R17831 VDD.n4503 VDD.n4502 0.0265784
R17832 VDD.n4502 VDD.n4501 0.0265784
R17833 VDD.n4505 VDD.n4496 0.0265784
R17834 VDD.n4506 VDD.n4505 0.0265784
R17835 VDD.n4508 VDD.n4507 0.0265784
R17836 VDD.n4507 VDD.n4506 0.0265784
R17837 VDD.n4501 VDD.n4498 0.0265784
R17838 VDD.n4498 VDD.n4497 0.0265784
R17839 VDD.n4521 VDD.n4520 0.0265784
R17840 VDD.t84 VDD.n4521 0.0265784
R17841 VDD.n4523 VDD.n4465 0.0265784
R17842 VDD.n4540 VDD.n4538 0.0265784
R17843 VDD.n4548 VDD.n4538 0.0265784
R17844 VDD.n4554 VDD.n4539 0.0265784
R17845 VDD.n4544 VDD.n4539 0.0265784
R17846 VDD.n4546 VDD.n4545 0.0265784
R17847 VDD.n4545 VDD.n4544 0.0265784
R17848 VDD.n4550 VDD.n4549 0.0265784
R17849 VDD.n4549 VDD.n4548 0.0265784
R17850 VDD.n4761 VDD.n4760 0.0265784
R17851 VDD.n4760 VDD.n4759 0.0265784
R17852 VDD.n4763 VDD.n4754 0.0265784
R17853 VDD.n4764 VDD.n4763 0.0265784
R17854 VDD.n4766 VDD.n4765 0.0265784
R17855 VDD.n4765 VDD.n4764 0.0265784
R17856 VDD.n4759 VDD.n4756 0.0265784
R17857 VDD.n4756 VDD.n4755 0.0265784
R17858 VDD.n4779 VDD.n4778 0.0265784
R17859 VDD.t717 VDD.n4779 0.0265784
R17860 VDD.n4781 VDD.n4723 0.0265784
R17861 VDD.n4798 VDD.n4796 0.0265784
R17862 VDD.n4806 VDD.n4796 0.0265784
R17863 VDD.n4812 VDD.n4797 0.0265784
R17864 VDD.n4802 VDD.n4797 0.0265784
R17865 VDD.n4804 VDD.n4803 0.0265784
R17866 VDD.n4803 VDD.n4802 0.0265784
R17867 VDD.n4808 VDD.n4807 0.0265784
R17868 VDD.n4807 VDD.n4806 0.0265784
R17869 VDD.n5019 VDD.n5018 0.0265784
R17870 VDD.n5018 VDD.n5017 0.0265784
R17871 VDD.n5021 VDD.n5012 0.0265784
R17872 VDD.n5022 VDD.n5021 0.0265784
R17873 VDD.n5024 VDD.n5023 0.0265784
R17874 VDD.n5023 VDD.n5022 0.0265784
R17875 VDD.n5017 VDD.n5014 0.0265784
R17876 VDD.n5014 VDD.n5013 0.0265784
R17877 VDD.n5037 VDD.n5036 0.0265784
R17878 VDD.t1353 VDD.n5037 0.0265784
R17879 VDD.n5039 VDD.n4981 0.0265784
R17880 VDD.n5056 VDD.n5054 0.0265784
R17881 VDD.n5064 VDD.n5054 0.0265784
R17882 VDD.n5070 VDD.n5055 0.0265784
R17883 VDD.n5060 VDD.n5055 0.0265784
R17884 VDD.n5062 VDD.n5061 0.0265784
R17885 VDD.n5061 VDD.n5060 0.0265784
R17886 VDD.n5066 VDD.n5065 0.0265784
R17887 VDD.n5065 VDD.n5064 0.0265784
R17888 VDD.n5277 VDD.n5276 0.0265784
R17889 VDD.n5276 VDD.n5275 0.0265784
R17890 VDD.n5279 VDD.n5270 0.0265784
R17891 VDD.n5280 VDD.n5279 0.0265784
R17892 VDD.n5282 VDD.n5281 0.0265784
R17893 VDD.n5281 VDD.n5280 0.0265784
R17894 VDD.n5275 VDD.n5272 0.0265784
R17895 VDD.n5272 VDD.n5271 0.0265784
R17896 VDD.n5295 VDD.n5294 0.0265784
R17897 VDD.t529 VDD.n5295 0.0265784
R17898 VDD.n5297 VDD.n5239 0.0265784
R17899 VDD.n5314 VDD.n5312 0.0265784
R17900 VDD.n5322 VDD.n5312 0.0265784
R17901 VDD.n5328 VDD.n5313 0.0265784
R17902 VDD.n5318 VDD.n5313 0.0265784
R17903 VDD.n5320 VDD.n5319 0.0265784
R17904 VDD.n5319 VDD.n5318 0.0265784
R17905 VDD.n5324 VDD.n5323 0.0265784
R17906 VDD.n5323 VDD.n5322 0.0265784
R17907 VDD.n1840 VDD.n1825 0.0261194
R17908 VDD.n2161 VDD.n2146 0.0261194
R17909 VDD.n2419 VDD.n2404 0.0261194
R17910 VDD.n2677 VDD.n2662 0.0261194
R17911 VDD.n2935 VDD.n2920 0.0261194
R17912 VDD.n3193 VDD.n3178 0.0261194
R17913 VDD.n3451 VDD.n3436 0.0261194
R17914 VDD.n5771 VDD.n5756 0.0261194
R17915 VDD.n5517 VDD.n5502 0.0261194
R17916 VDD.n3709 VDD.n3694 0.0261194
R17917 VDD.n3967 VDD.n3952 0.0261194
R17918 VDD.n4225 VDD.n4210 0.0261194
R17919 VDD.n4483 VDD.n4468 0.0261194
R17920 VDD.n4741 VDD.n4726 0.0261194
R17921 VDD.n4999 VDD.n4984 0.0261194
R17922 VDD.n5257 VDD.n5242 0.0261194
R17923 VDD.n1304 VDD 0.0260435
R17924 VDD.n1945 VDD.n1922 0.0258165
R17925 VDD.n1696 VDD.n1683 0.0257918
R17926 VDD.n2045 VDD.n2032 0.0257918
R17927 VDD.n2275 VDD.n2262 0.0257918
R17928 VDD.n2533 VDD.n2520 0.0257918
R17929 VDD.n2791 VDD.n2778 0.0257918
R17930 VDD.n3049 VDD.n3036 0.0257918
R17931 VDD.n3307 VDD.n3294 0.0257918
R17932 VDD.n5630 VDD.n5617 0.0257918
R17933 VDD.n5376 VDD.n5363 0.0257918
R17934 VDD.n3565 VDD.n3552 0.0257918
R17935 VDD.n3823 VDD.n3810 0.0257918
R17936 VDD.n4081 VDD.n4068 0.0257918
R17937 VDD.n4339 VDD.n4326 0.0257918
R17938 VDD.n4597 VDD.n4584 0.0257918
R17939 VDD.n4855 VDD.n4842 0.0257918
R17940 VDD.n5113 VDD.n5100 0.0257918
R17941 VDD.n1880 VDD.n1879 0.02576
R17942 VDD.n2201 VDD.n2200 0.02576
R17943 VDD.n2459 VDD.n2458 0.02576
R17944 VDD.n2717 VDD.n2716 0.02576
R17945 VDD.n2975 VDD.n2974 0.02576
R17946 VDD.n3233 VDD.n3232 0.02576
R17947 VDD.n3491 VDD.n3490 0.02576
R17948 VDD.n5811 VDD.n5810 0.02576
R17949 VDD.n5557 VDD.n5556 0.02576
R17950 VDD.n3749 VDD.n3748 0.02576
R17951 VDD.n4007 VDD.n4006 0.02576
R17952 VDD.n4265 VDD.n4264 0.02576
R17953 VDD.n4523 VDD.n4522 0.02576
R17954 VDD.n4781 VDD.n4780 0.02576
R17955 VDD.n5039 VDD.n5038 0.02576
R17956 VDD.n5297 VDD.n5296 0.02576
R17957 VDD.n1315 VDD.n1314 0.0254026
R17958 VDD.n1310 VDD.n1308 0.0249681
R17959 VDD.n1311 VDD.n1310 0.0249681
R17960 VDD.n1453 VDD.n1449 0.0249681
R17961 VDD.n1449 VDD.n1447 0.0249681
R17962 VDD.n1447 VDD.n1443 0.0249681
R17963 VDD.n1443 VDD.n1441 0.0249681
R17964 VDD.n1441 VDD.n1437 0.0249681
R17965 VDD.n1437 VDD.n1433 0.0249681
R17966 VDD.n1331 VDD.n1327 0.0249681
R17967 VDD.n1333 VDD.n1331 0.0249681
R17968 VDD.n1337 VDD.n1333 0.0249681
R17969 VDD.n1339 VDD.n1337 0.0249681
R17970 VDD.n1340 VDD.n1339 0.0249681
R17971 VDD.n1422 VDD.n1418 0.0249681
R17972 VDD.n1418 VDD.n1416 0.0249681
R17973 VDD.n1416 VDD.n1412 0.0249681
R17974 VDD.n1412 VDD.n1410 0.0249681
R17975 VDD.n1393 VDD.n1389 0.0249681
R17976 VDD.n1389 VDD.n1387 0.0249681
R17977 VDD.n1387 VDD.n1383 0.0249681
R17978 VDD.n1383 VDD.n1381 0.0249681
R17979 VDD.n1351 VDD.n1349 0.0249681
R17980 VDD.n1354 VDD.n1351 0.0249681
R17981 VDD.n1356 VDD.n1354 0.0249681
R17982 VDD.n1358 VDD.n1356 0.0249681
R17983 VDD.n1365 VDD.n1363 0.0249681
R17984 VDD.n1525 VDD.n1523 0.0249681
R17985 VDD.n1523 VDD.n1519 0.0249681
R17986 VDD.n1519 VDD.n1517 0.0249681
R17987 VDD.n1517 VDD.n1513 0.0249681
R17988 VDD.n1503 VDD.n1501 0.0249681
R17989 VDD.n1501 VDD.n1497 0.0249681
R17990 VDD.n1497 VDD.n1495 0.0249681
R17991 VDD.n1495 VDD.n1491 0.0249681
R17992 VDD.n1491 VDD.n1489 0.0249681
R17993 VDD.n1489 VDD.n1485 0.0249681
R17994 VDD.n1485 VDD.n1481 0.0249681
R17995 VDD.n1481 VDD.n1479 0.0249681
R17996 VDD.n1479 VDD.n1475 0.0249681
R17997 VDD.n1475 VDD.n1473 0.0249681
R17998 VDD.n1473 VDD.n1469 0.0249681
R17999 VDD.n1469 VDD.n1467 0.0249681
R18000 VDD.n1467 VDD.n1463 0.0249681
R18001 VDD.n1286 VDD.n1285 0.0249681
R18002 VDD.n1285 VDD.n1283 0.0249681
R18003 VDD.n1546 VDD.n1544 0.0243281
R18004 VDD.n1454 VDD.n1453 0.0241145
R18005 VDD.n1882 VDD.n1881 0.0228205
R18006 VDD.n2203 VDD.n2202 0.0228205
R18007 VDD.n2461 VDD.n2460 0.0228205
R18008 VDD.n2719 VDD.n2718 0.0228205
R18009 VDD.n2977 VDD.n2976 0.0228205
R18010 VDD.n3235 VDD.n3234 0.0228205
R18011 VDD.n3493 VDD.n3492 0.0228205
R18012 VDD.n5813 VDD.n5812 0.0228205
R18013 VDD.n5559 VDD.n5558 0.0228205
R18014 VDD.n3751 VDD.n3750 0.0228205
R18015 VDD.n4009 VDD.n4008 0.0228205
R18016 VDD.n4267 VDD.n4266 0.0228205
R18017 VDD.n4525 VDD.n4524 0.0228205
R18018 VDD.n4783 VDD.n4782 0.0228205
R18019 VDD.n5041 VDD.n5040 0.0228205
R18020 VDD.n5299 VDD.n5298 0.0228205
R18021 VDD.n1881 VDD.n1820 0.0223212
R18022 VDD.n2202 VDD.n2141 0.0223212
R18023 VDD.n2460 VDD.n2399 0.0223212
R18024 VDD.n2718 VDD.n2657 0.0223212
R18025 VDD.n2976 VDD.n2915 0.0223212
R18026 VDD.n3234 VDD.n3173 0.0223212
R18027 VDD.n3492 VDD.n3431 0.0223212
R18028 VDD.n5812 VDD.n5751 0.0223212
R18029 VDD.n5558 VDD.n5497 0.0223212
R18030 VDD.n3750 VDD.n3689 0.0223212
R18031 VDD.n4008 VDD.n3947 0.0223212
R18032 VDD.n4266 VDD.n4205 0.0223212
R18033 VDD.n4524 VDD.n4463 0.0223212
R18034 VDD.n4782 VDD.n4721 0.0223212
R18035 VDD.n5040 VDD.n4979 0.0223212
R18036 VDD.n5298 VDD.n5237 0.0223212
R18037 VDD.n1374 VDD.n1346 0.0218724
R18038 VDD.n851 VDD 0.02175
R18039 VDD.n845 VDD 0.02175
R18040 VDD.n839 VDD 0.02175
R18041 VDD.n833 VDD 0.02175
R18042 VDD.n827 VDD 0.02175
R18043 VDD.n1234 VDD 0.02175
R18044 VDD.n1228 VDD 0.02175
R18045 VDD.n1222 VDD 0.02175
R18046 VDD.n1216 VDD 0.02175
R18047 VDD.n1210 VDD 0.02175
R18048 VDD.n1600 VDD 0.0213145
R18049 VDD.n1410 VDD.n1406 0.0212447
R18050 VDD.n1504 VDD.n1503 0.0207128
R18051 VDD.n1622 VDD.n1621 0.0205312
R18052 VDD.n1433 VDD.n1431 0.0198592
R18053 VDD.n1461 VDD.n1460 0.0188511
R18054 VDD.n1946 VDD.n1945 0.0183679
R18055 VDD.n1799 VDD.n1798 0.0182941
R18056 VDD.n2007 VDD.n2006 0.0182941
R18057 VDD.n2378 VDD.n2377 0.0182941
R18058 VDD.n2636 VDD.n2635 0.0182941
R18059 VDD.n2894 VDD.n2893 0.0182941
R18060 VDD.n3152 VDD.n3151 0.0182941
R18061 VDD.n3410 VDD.n3409 0.0182941
R18062 VDD.n5733 VDD.n5732 0.0182941
R18063 VDD.n5479 VDD.n5478 0.0182941
R18064 VDD.n3668 VDD.n3667 0.0182941
R18065 VDD.n3926 VDD.n3925 0.0182941
R18066 VDD.n4184 VDD.n4183 0.0182941
R18067 VDD.n4442 VDD.n4441 0.0182941
R18068 VDD.n4700 VDD.n4699 0.0182941
R18069 VDD.n4958 VDD.n4957 0.0182941
R18070 VDD.n5216 VDD.n5215 0.0182941
R18071 VDD.n1779 VDD.n1777 0.0178611
R18072 VDD.n1987 VDD.n1985 0.0178611
R18073 VDD.n2358 VDD.n2356 0.0178611
R18074 VDD.n2616 VDD.n2614 0.0178611
R18075 VDD.n2874 VDD.n2872 0.0178611
R18076 VDD.n3132 VDD.n3130 0.0178611
R18077 VDD.n3390 VDD.n3388 0.0178611
R18078 VDD.n5713 VDD.n5711 0.0178611
R18079 VDD.n5459 VDD.n5457 0.0178611
R18080 VDD.n3648 VDD.n3646 0.0178611
R18081 VDD.n3906 VDD.n3904 0.0178611
R18082 VDD.n4164 VDD.n4162 0.0178611
R18083 VDD.n4422 VDD.n4420 0.0178611
R18084 VDD.n4680 VDD.n4678 0.0178611
R18085 VDD.n4938 VDD.n4936 0.0178611
R18086 VDD.n5196 VDD.n5194 0.0178611
R18087 VDD.n1808 VDD.n1807 0.0177731
R18088 VDD.n2387 VDD.n2386 0.0177731
R18089 VDD.n2645 VDD.n2644 0.0177731
R18090 VDD.n2903 VDD.n2902 0.0177731
R18091 VDD.n3161 VDD.n3160 0.0177731
R18092 VDD.n3419 VDD.n3418 0.0177731
R18093 VDD.n3677 VDD.n3676 0.0177731
R18094 VDD.n3935 VDD.n3934 0.0177731
R18095 VDD.n4193 VDD.n4192 0.0177731
R18096 VDD.n4451 VDD.n4450 0.0177731
R18097 VDD.n4709 VDD.n4708 0.0177731
R18098 VDD.n4967 VDD.n4966 0.0177731
R18099 VDD.n5225 VDD.n5224 0.0177731
R18100 VDD.n1368 VDD.n1366 0.0172553
R18101 VDD.n810 VDD 0.0171185
R18102 VDD VDD.n799 0.0171185
R18103 VDD.n1193 VDD 0.0171185
R18104 VDD VDD.n1182 0.0171185
R18105 VDD.n1758 VDD.n1757 0.0168386
R18106 VDD.n2107 VDD.n2106 0.0168386
R18107 VDD.n2337 VDD.n2336 0.0168386
R18108 VDD.n2595 VDD.n2594 0.0168386
R18109 VDD.n2853 VDD.n2852 0.0168386
R18110 VDD.n3111 VDD.n3110 0.0168386
R18111 VDD.n3369 VDD.n3368 0.0168386
R18112 VDD.n5692 VDD.n5691 0.0168386
R18113 VDD.n5438 VDD.n5437 0.0168386
R18114 VDD.n3627 VDD.n3626 0.0168386
R18115 VDD.n3885 VDD.n3884 0.0168386
R18116 VDD.n4143 VDD.n4142 0.0168386
R18117 VDD.n4401 VDD.n4400 0.0168386
R18118 VDD.n4659 VDD.n4658 0.0168386
R18119 VDD.n4917 VDD.n4916 0.0168386
R18120 VDD.n5175 VDD.n5174 0.0168386
R18121 VDD.n1710 VDD.n1679 0.0168372
R18122 VDD.n2059 VDD.n2028 0.0168372
R18123 VDD.n2289 VDD.n2258 0.0168372
R18124 VDD.n2547 VDD.n2516 0.0168372
R18125 VDD.n2805 VDD.n2774 0.0168372
R18126 VDD.n3063 VDD.n3032 0.0168372
R18127 VDD.n3321 VDD.n3290 0.0168372
R18128 VDD.n5644 VDD.n5613 0.0168372
R18129 VDD.n5390 VDD.n5359 0.0168372
R18130 VDD.n3579 VDD.n3548 0.0168372
R18131 VDD.n3837 VDD.n3806 0.0168372
R18132 VDD.n4095 VDD.n4064 0.0168372
R18133 VDD.n4353 VDD.n4322 0.0168372
R18134 VDD.n4611 VDD.n4580 0.0168372
R18135 VDD.n4869 VDD.n4838 0.0168372
R18136 VDD.n5127 VDD.n5096 0.0168372
R18137 VDD.n861 VDD.n860 0.0165987
R18138 VDD.n1244 VDD.n1243 0.0165987
R18139 VDD.n1679 VDD.n1669 0.0163404
R18140 VDD.n1758 VDD.n1717 0.0163404
R18141 VDD.n2028 VDD.n2018 0.0163404
R18142 VDD.n2107 VDD.n2066 0.0163404
R18143 VDD.n2258 VDD.n2248 0.0163404
R18144 VDD.n2337 VDD.n2296 0.0163404
R18145 VDD.n2516 VDD.n2506 0.0163404
R18146 VDD.n2595 VDD.n2554 0.0163404
R18147 VDD.n2774 VDD.n2764 0.0163404
R18148 VDD.n2853 VDD.n2812 0.0163404
R18149 VDD.n3032 VDD.n3022 0.0163404
R18150 VDD.n3111 VDD.n3070 0.0163404
R18151 VDD.n3290 VDD.n3280 0.0163404
R18152 VDD.n3369 VDD.n3328 0.0163404
R18153 VDD.n5613 VDD.n5603 0.0163404
R18154 VDD.n5692 VDD.n5651 0.0163404
R18155 VDD.n5359 VDD.n5349 0.0163404
R18156 VDD.n5438 VDD.n5397 0.0163404
R18157 VDD.n3548 VDD.n3538 0.0163404
R18158 VDD.n3627 VDD.n3586 0.0163404
R18159 VDD.n3806 VDD.n3796 0.0163404
R18160 VDD.n3885 VDD.n3844 0.0163404
R18161 VDD.n4064 VDD.n4054 0.0163404
R18162 VDD.n4143 VDD.n4102 0.0163404
R18163 VDD.n4322 VDD.n4312 0.0163404
R18164 VDD.n4401 VDD.n4360 0.0163404
R18165 VDD.n4580 VDD.n4570 0.0163404
R18166 VDD.n4659 VDD.n4618 0.0163404
R18167 VDD.n4838 VDD.n4828 0.0163404
R18168 VDD.n4917 VDD.n4876 0.0163404
R18169 VDD.n5096 VDD.n5086 0.0163404
R18170 VDD.n5175 VDD.n5134 0.0163404
R18171 VDD.n1423 VDD.n1422 0.0161915
R18172 VDD.n855 VDD.n854 0.016125
R18173 VDD.n1238 VDD.n1237 0.016125
R18174 VDD.n1961 VDD.n1941 0.0154506
R18175 VDD.n1969 VDD.n1968 0.015449
R18176 VDD.n1405 VDD.n1401 0.0153936
R18177 VDD.n1513 VDD.n1511 0.0151277
R18178 VDD.n1971 VDD.n1970 0.0150463
R18179 VDD.n1970 VDD.t1043 0.0150463
R18180 VDD.n1963 VDD.n1929 0.0150463
R18181 VDD.t863 VDD.n1963 0.0150463
R18182 VDD.n1961 VDD.n1960 0.0150463
R18183 VDD.n1964 VDD.t863 0.0150463
R18184 VDD.n1968 VDD.n1967 0.0150463
R18185 VDD.n1965 VDD.n1964 0.0150463
R18186 VDD.t1041 VDD.n1951 0.0150463
R18187 VDD.n1951 VDD.n1950 0.0150463
R18188 VDD.n794 VDD.n513 0.015
R18189 VDD.n1839 VDD.n1827 0.0149834
R18190 VDD.n2160 VDD.n2148 0.0149834
R18191 VDD.n2418 VDD.n2406 0.0149834
R18192 VDD.n2676 VDD.n2664 0.0149834
R18193 VDD.n2934 VDD.n2922 0.0149834
R18194 VDD.n3192 VDD.n3180 0.0149834
R18195 VDD.n3450 VDD.n3438 0.0149834
R18196 VDD.n5770 VDD.n5758 0.0149834
R18197 VDD.n5516 VDD.n5504 0.0149834
R18198 VDD.n3708 VDD.n3696 0.0149834
R18199 VDD.n3966 VDD.n3954 0.0149834
R18200 VDD.n4224 VDD.n4212 0.0149834
R18201 VDD.n4482 VDD.n4470 0.0149834
R18202 VDD.n4740 VDD.n4728 0.0149834
R18203 VDD.n4998 VDD.n4986 0.0149834
R18204 VDD.n5256 VDD.n5244 0.0149834
R18205 VDD.n1325 VDD.n1324 0.0148617
R18206 VDD.n676 VDD.n674 0.0146339
R18207 VDD.n1026 VDD.n1024 0.0146339
R18208 VDD.n271 VDD.n269 0.0146339
R18209 VDD.n1394 VDD.n1393 0.0145957
R18210 VDD.n1377 VDD.n1376 0.0145957
R18211 VDD.n1886 VDD.n1817 0.0145797
R18212 VDD.n2207 VDD.n2138 0.0145797
R18213 VDD.n2465 VDD.n2396 0.0145797
R18214 VDD.n2723 VDD.n2654 0.0145797
R18215 VDD.n2981 VDD.n2912 0.0145797
R18216 VDD.n3239 VDD.n3170 0.0145797
R18217 VDD.n3497 VDD.n3428 0.0145797
R18218 VDD.n5817 VDD.n5748 0.0145797
R18219 VDD.n5563 VDD.n5494 0.0145797
R18220 VDD.n3755 VDD.n3686 0.0145797
R18221 VDD.n4013 VDD.n3944 0.0145797
R18222 VDD.n4271 VDD.n4202 0.0145797
R18223 VDD.n4529 VDD.n4460 0.0145797
R18224 VDD.n4787 VDD.n4718 0.0145797
R18225 VDD.n5045 VDD.n4976 0.0145797
R18226 VDD.n5303 VDD.n5234 0.0145797
R18227 VDD.n1721 VDD.n1720 0.0143889
R18228 VDD.n2070 VDD.n2069 0.0143889
R18229 VDD.n2300 VDD.n2299 0.0143889
R18230 VDD.n2558 VDD.n2557 0.0143889
R18231 VDD.n2816 VDD.n2815 0.0143889
R18232 VDD.n3074 VDD.n3073 0.0143889
R18233 VDD.n3332 VDD.n3331 0.0143889
R18234 VDD.n5655 VDD.n5654 0.0143889
R18235 VDD.n5401 VDD.n5400 0.0143889
R18236 VDD.n3590 VDD.n3589 0.0143889
R18237 VDD.n3848 VDD.n3847 0.0143889
R18238 VDD.n4106 VDD.n4105 0.0143889
R18239 VDD.n4364 VDD.n4363 0.0143889
R18240 VDD.n4622 VDD.n4621 0.0143889
R18241 VDD.n4880 VDD.n4879 0.0143889
R18242 VDD.n5138 VDD.n5137 0.0143889
R18243 VDD.n485 VDD.n481 0.0143889
R18244 VDD.n83 VDD.n79 0.0143889
R18245 VDD.n1308 VDD.n1304 0.0143298
R18246 VDD.n1180 VDD.n1179 0.0142984
R18247 VDD.n1979 VDD.n1978 0.0138929
R18248 VDD.n1345 VDD.n1343 0.0137979
R18249 VDD VDD.n1840 0.0131689
R18250 VDD VDD.n2161 0.0131689
R18251 VDD VDD.n2419 0.0131689
R18252 VDD VDD.n2677 0.0131689
R18253 VDD VDD.n2935 0.0131689
R18254 VDD VDD.n3193 0.0131689
R18255 VDD VDD.n3451 0.0131689
R18256 VDD VDD.n5771 0.0131689
R18257 VDD VDD.n5517 0.0131689
R18258 VDD VDD.n3709 0.0131689
R18259 VDD VDD.n3967 0.0131689
R18260 VDD VDD.n4225 0.0131689
R18261 VDD VDD.n4483 0.0131689
R18262 VDD VDD.n4741 0.0131689
R18263 VDD VDD.n4999 0.0131689
R18264 VDD VDD.n5257 0.0131689
R18265 VDD.n447 VDD 0.013
R18266 VDD.n44 VDD 0.013
R18267 VDD.n1314 VDD 0.012734
R18268 VDD.n1349 VDD 0.012734
R18269 VDD.n1261 VDD 0.012734
R18270 VDD.n1544 VDD.n1543 0.0126094
R18271 VDD.n537 VDD.n533 0.0126053
R18272 VDD.n576 VDD.n572 0.0126053
R18273 VDD.n572 VDD.n570 0.0126053
R18274 VDD.n570 VDD.n566 0.0126053
R18275 VDD.n566 VDD.n564 0.0126053
R18276 VDD.n564 VDD.n560 0.0126053
R18277 VDD.n560 VDD.n558 0.0126053
R18278 VDD.n558 VDD.n554 0.0126053
R18279 VDD.n554 VDD.n552 0.0126053
R18280 VDD.n551 VDD.n550 0.0126053
R18281 VDD.n550 VDD.n548 0.0126053
R18282 VDD.n548 VDD.n544 0.0126053
R18283 VDD.n544 VDD.n528 0.0126053
R18284 VDD.n598 VDD.n594 0.0126053
R18285 VDD.n600 VDD.n598 0.0126053
R18286 VDD.n604 VDD.n600 0.0126053
R18287 VDD.n606 VDD.n604 0.0126053
R18288 VDD.n610 VDD.n606 0.0126053
R18289 VDD.n612 VDD.n610 0.0126053
R18290 VDD.n616 VDD.n612 0.0126053
R18291 VDD.n618 VDD.n616 0.0126053
R18292 VDD.n619 VDD.n618 0.0126053
R18293 VDD.n624 VDD.n622 0.0126053
R18294 VDD.n628 VDD.n624 0.0126053
R18295 VDD.n630 VDD.n628 0.0126053
R18296 VDD.n634 VDD.n630 0.0126053
R18297 VDD.n659 VDD.n655 0.0126053
R18298 VDD.n655 VDD.n653 0.0126053
R18299 VDD.n653 VDD.n649 0.0126053
R18300 VDD.n649 VDD.n647 0.0126053
R18301 VDD.n647 VDD.n643 0.0126053
R18302 VDD.n643 VDD.n641 0.0126053
R18303 VDD.n641 VDD.n515 0.0126053
R18304 VDD.n791 VDD.n790 0.0126053
R18305 VDD.n790 VDD.n788 0.0126053
R18306 VDD.n775 VDD.n773 0.0126053
R18307 VDD.n773 VDD.n769 0.0126053
R18308 VDD.n769 VDD.n765 0.0126053
R18309 VDD.n765 VDD.n763 0.0126053
R18310 VDD.n763 VDD.n759 0.0126053
R18311 VDD.n759 VDD.n757 0.0126053
R18312 VDD.n757 VDD.n753 0.0126053
R18313 VDD.n753 VDD.n751 0.0126053
R18314 VDD.n751 VDD.n747 0.0126053
R18315 VDD.n747 VDD.n745 0.0126053
R18316 VDD.n744 VDD.n743 0.0126053
R18317 VDD.n732 VDD.n728 0.0126053
R18318 VDD.n728 VDD.n726 0.0126053
R18319 VDD.n726 VDD.n722 0.0126053
R18320 VDD.n722 VDD.n718 0.0126053
R18321 VDD.n718 VDD.n716 0.0126053
R18322 VDD.n716 VDD.n712 0.0126053
R18323 VDD.n712 VDD.n710 0.0126053
R18324 VDD.n710 VDD.n706 0.0126053
R18325 VDD.n706 VDD.n704 0.0126053
R18326 VDD.n704 VDD.n700 0.0126053
R18327 VDD.n700 VDD.n698 0.0126053
R18328 VDD.n697 VDD.n696 0.0126053
R18329 VDD.n696 VDD.n694 0.0126053
R18330 VDD.n694 VDD.n691 0.0126053
R18331 VDD.n691 VDD.n689 0.0126053
R18332 VDD.n682 VDD.n680 0.0126053
R18333 VDD.n677 VDD.n676 0.0126053
R18334 VDD.n887 VDD.n883 0.0126053
R18335 VDD.n926 VDD.n922 0.0126053
R18336 VDD.n922 VDD.n920 0.0126053
R18337 VDD.n920 VDD.n916 0.0126053
R18338 VDD.n916 VDD.n914 0.0126053
R18339 VDD.n914 VDD.n910 0.0126053
R18340 VDD.n910 VDD.n908 0.0126053
R18341 VDD.n908 VDD.n904 0.0126053
R18342 VDD.n904 VDD.n902 0.0126053
R18343 VDD.n901 VDD.n900 0.0126053
R18344 VDD.n900 VDD.n898 0.0126053
R18345 VDD.n898 VDD.n894 0.0126053
R18346 VDD.n894 VDD.n878 0.0126053
R18347 VDD.n948 VDD.n944 0.0126053
R18348 VDD.n950 VDD.n948 0.0126053
R18349 VDD.n954 VDD.n950 0.0126053
R18350 VDD.n956 VDD.n954 0.0126053
R18351 VDD.n960 VDD.n956 0.0126053
R18352 VDD.n962 VDD.n960 0.0126053
R18353 VDD.n966 VDD.n962 0.0126053
R18354 VDD.n968 VDD.n966 0.0126053
R18355 VDD.n969 VDD.n968 0.0126053
R18356 VDD.n974 VDD.n972 0.0126053
R18357 VDD.n978 VDD.n974 0.0126053
R18358 VDD.n980 VDD.n978 0.0126053
R18359 VDD.n984 VDD.n980 0.0126053
R18360 VDD.n1009 VDD.n1005 0.0126053
R18361 VDD.n1005 VDD.n1003 0.0126053
R18362 VDD.n1003 VDD.n999 0.0126053
R18363 VDD.n999 VDD.n997 0.0126053
R18364 VDD.n997 VDD.n993 0.0126053
R18365 VDD.n993 VDD.n991 0.0126053
R18366 VDD.n991 VDD.n865 0.0126053
R18367 VDD.n1141 VDD.n1140 0.0126053
R18368 VDD.n1140 VDD.n1138 0.0126053
R18369 VDD.n1125 VDD.n1123 0.0126053
R18370 VDD.n1123 VDD.n1119 0.0126053
R18371 VDD.n1119 VDD.n1115 0.0126053
R18372 VDD.n1115 VDD.n1113 0.0126053
R18373 VDD.n1113 VDD.n1109 0.0126053
R18374 VDD.n1109 VDD.n1107 0.0126053
R18375 VDD.n1107 VDD.n1103 0.0126053
R18376 VDD.n1103 VDD.n1101 0.0126053
R18377 VDD.n1101 VDD.n1097 0.0126053
R18378 VDD.n1097 VDD.n1095 0.0126053
R18379 VDD.n1094 VDD.n1093 0.0126053
R18380 VDD.n1082 VDD.n1078 0.0126053
R18381 VDD.n1078 VDD.n1076 0.0126053
R18382 VDD.n1076 VDD.n1072 0.0126053
R18383 VDD.n1072 VDD.n1068 0.0126053
R18384 VDD.n1068 VDD.n1066 0.0126053
R18385 VDD.n1066 VDD.n1062 0.0126053
R18386 VDD.n1062 VDD.n1060 0.0126053
R18387 VDD.n1060 VDD.n1056 0.0126053
R18388 VDD.n1056 VDD.n1054 0.0126053
R18389 VDD.n1054 VDD.n1050 0.0126053
R18390 VDD.n1050 VDD.n1048 0.0126053
R18391 VDD.n1047 VDD.n1046 0.0126053
R18392 VDD.n1046 VDD.n1044 0.0126053
R18393 VDD.n1044 VDD.n1041 0.0126053
R18394 VDD.n1041 VDD.n1039 0.0126053
R18395 VDD.n1032 VDD.n1030 0.0126053
R18396 VDD.n1027 VDD.n1026 0.0126053
R18397 VDD.n136 VDD.n132 0.0126053
R18398 VDD.n175 VDD.n171 0.0126053
R18399 VDD.n171 VDD.n169 0.0126053
R18400 VDD.n169 VDD.n165 0.0126053
R18401 VDD.n165 VDD.n163 0.0126053
R18402 VDD.n163 VDD.n159 0.0126053
R18403 VDD.n159 VDD.n157 0.0126053
R18404 VDD.n157 VDD.n153 0.0126053
R18405 VDD.n153 VDD.n151 0.0126053
R18406 VDD.n150 VDD.n149 0.0126053
R18407 VDD.n149 VDD.n147 0.0126053
R18408 VDD.n147 VDD.n143 0.0126053
R18409 VDD.n143 VDD.n127 0.0126053
R18410 VDD.n197 VDD.n193 0.0126053
R18411 VDD.n199 VDD.n197 0.0126053
R18412 VDD.n203 VDD.n199 0.0126053
R18413 VDD.n205 VDD.n203 0.0126053
R18414 VDD.n209 VDD.n205 0.0126053
R18415 VDD.n211 VDD.n209 0.0126053
R18416 VDD.n215 VDD.n211 0.0126053
R18417 VDD.n217 VDD.n215 0.0126053
R18418 VDD.n218 VDD.n217 0.0126053
R18419 VDD.n223 VDD.n221 0.0126053
R18420 VDD.n227 VDD.n223 0.0126053
R18421 VDD.n229 VDD.n227 0.0126053
R18422 VDD.n233 VDD.n229 0.0126053
R18423 VDD.n254 VDD.n250 0.0126053
R18424 VDD.n250 VDD.n248 0.0126053
R18425 VDD.n248 VDD.n244 0.0126053
R18426 VDD.n244 VDD.n242 0.0126053
R18427 VDD.n242 VDD.n238 0.0126053
R18428 VDD.n238 VDD.n114 0.0126053
R18429 VDD.n389 VDD.n387 0.0126053
R18430 VDD.n386 VDD.n385 0.0126053
R18431 VDD.n385 VDD.n383 0.0126053
R18432 VDD.n370 VDD.n368 0.0126053
R18433 VDD.n368 VDD.n364 0.0126053
R18434 VDD.n364 VDD.n360 0.0126053
R18435 VDD.n360 VDD.n358 0.0126053
R18436 VDD.n358 VDD.n354 0.0126053
R18437 VDD.n354 VDD.n352 0.0126053
R18438 VDD.n352 VDD.n348 0.0126053
R18439 VDD.n348 VDD.n346 0.0126053
R18440 VDD.n346 VDD.n342 0.0126053
R18441 VDD.n342 VDD.n340 0.0126053
R18442 VDD.n339 VDD.n338 0.0126053
R18443 VDD.n327 VDD.n323 0.0126053
R18444 VDD.n323 VDD.n321 0.0126053
R18445 VDD.n321 VDD.n317 0.0126053
R18446 VDD.n317 VDD.n313 0.0126053
R18447 VDD.n313 VDD.n311 0.0126053
R18448 VDD.n311 VDD.n307 0.0126053
R18449 VDD.n307 VDD.n305 0.0126053
R18450 VDD.n305 VDD.n301 0.0126053
R18451 VDD.n301 VDD.n299 0.0126053
R18452 VDD.n299 VDD.n295 0.0126053
R18453 VDD.n295 VDD.n293 0.0126053
R18454 VDD.n292 VDD.n291 0.0126053
R18455 VDD.n291 VDD.n289 0.0126053
R18456 VDD.n289 VDD.n286 0.0126053
R18457 VDD.n286 VDD.n284 0.0126053
R18458 VDD.n277 VDD.n275 0.0126053
R18459 VDD.n272 VDD.n271 0.0126053
R18460 VDD.n474 VDD 0.0125739
R18461 VDD.n72 VDD 0.0125739
R18462 VDD.n1611 VDD.n1609 0.0125192
R18463 VDD.n793 VDD.n792 0.0124737
R18464 VDD.n1143 VDD.n1142 0.0124737
R18465 VDD.n1785 VDD 0.0123056
R18466 VDD.n1993 VDD 0.0123056
R18467 VDD.n2364 VDD 0.0123056
R18468 VDD.n2622 VDD 0.0123056
R18469 VDD.n2880 VDD 0.0123056
R18470 VDD.n3138 VDD 0.0123056
R18471 VDD.n3396 VDD 0.0123056
R18472 VDD.n5719 VDD 0.0123056
R18473 VDD.n5465 VDD 0.0123056
R18474 VDD.n3654 VDD 0.0123056
R18475 VDD.n3912 VDD 0.0123056
R18476 VDD.n4170 VDD 0.0123056
R18477 VDD.n4428 VDD 0.0123056
R18478 VDD.n4686 VDD 0.0123056
R18479 VDD.n4944 VDD 0.0123056
R18480 VDD.n5202 VDD 0.0123056
R18481 VDD VDD.n467 0.0123056
R18482 VDD.n413 VDD 0.0123056
R18483 VDD VDD.n65 0.0123056
R18484 VDD.n1571 VDD 0.0123056
R18485 VDD.n390 VDD.n114 0.0122105
R18486 VDD.n587 VDD.n528 0.0119152
R18487 VDD.n937 VDD.n878 0.0119152
R18488 VDD.n1842 VDD 0.0118881
R18489 VDD.n2163 VDD 0.0118881
R18490 VDD.n2421 VDD 0.0118881
R18491 VDD.n2679 VDD 0.0118881
R18492 VDD.n2937 VDD 0.0118881
R18493 VDD.n3195 VDD 0.0118881
R18494 VDD.n3453 VDD 0.0118881
R18495 VDD.n5773 VDD 0.0118881
R18496 VDD.n5519 VDD 0.0118881
R18497 VDD.n3711 VDD 0.0118881
R18498 VDD.n3969 VDD 0.0118881
R18499 VDD.n4227 VDD 0.0118881
R18500 VDD.n4485 VDD 0.0118881
R18501 VDD.n4743 VDD 0.0118881
R18502 VDD.n5001 VDD 0.0118881
R18503 VDD.n5259 VDD 0.0118881
R18504 VDD.n1255 VDD.n1251 0.0117745
R18505 VDD.n1539 VDD.n1537 0.0117745
R18506 VDD.n1537 VDD.n1533 0.0117745
R18507 VDD.n1533 VDD.n1529 0.0117745
R18508 VDD.n1529 VDD.n1527 0.0117745
R18509 VDD.n1613 VDD.n1611 0.0117367
R18510 VDD.n501 VDD 0.0116111
R18511 VDD.n428 VDD 0.0116111
R18512 VDD.n394 VDD 0.0116111
R18513 VDD.n99 VDD 0.0116111
R18514 VDD.n1586 VDD 0.0116111
R18515 VDD.n1552 VDD 0.0116111
R18516 VDD.n11 VDD 0.0114012
R18517 VDD.n1155 VDD 0.0114012
R18518 VDD.n186 VDD.n127 0.0113889
R18519 VDD.n1875 VDD.n1874 0.0111456
R18520 VDD.n2196 VDD.n2195 0.0111456
R18521 VDD.n2454 VDD.n2453 0.0111456
R18522 VDD.n2712 VDD.n2711 0.0111456
R18523 VDD.n2970 VDD.n2969 0.0111456
R18524 VDD.n3228 VDD.n3227 0.0111456
R18525 VDD.n3486 VDD.n3485 0.0111456
R18526 VDD.n5806 VDD.n5805 0.0111456
R18527 VDD.n5552 VDD.n5551 0.0111456
R18528 VDD.n3744 VDD.n3743 0.0111456
R18529 VDD.n4002 VDD.n4001 0.0111456
R18530 VDD.n4260 VDD.n4259 0.0111456
R18531 VDD.n4518 VDD.n4517 0.0111456
R18532 VDD.n4776 VDD.n4775 0.0111456
R18533 VDD.n5034 VDD.n5033 0.0111456
R18534 VDD.n5292 VDD.n5291 0.0111456
R18535 VDD.n255 VDD.n254 0.0108947
R18536 VDD.n1396 VDD.n1394 0.0108723
R18537 VDD.n1381 VDD.n1377 0.0108723
R18538 VDD.n1957 VDD.n1922 0.0108144
R18539 VDD.n371 VDD.n370 0.0106316
R18540 VDD.n328 VDD.n327 0.0106316
R18541 VDD.n1327 VDD.n1325 0.0106064
R18542 VDD.n538 VDD.n537 0.0103684
R18543 VDD.n660 VDD.n659 0.0103684
R18544 VDD.n888 VDD.n887 0.0103684
R18545 VDD.n1010 VDD.n1009 0.0103684
R18546 VDD.n1426 VDD.n1425 0.0103404
R18547 VDD.n1511 VDD.n1510 0.0103404
R18548 VDD.n1527 VDD.n1526 0.0103039
R18549 VDD.n1696 VDD.n1695 0.0101514
R18550 VDD.n2045 VDD.n2044 0.0101514
R18551 VDD.n2275 VDD.n2274 0.0101514
R18552 VDD.n2533 VDD.n2532 0.0101514
R18553 VDD.n2791 VDD.n2790 0.0101514
R18554 VDD.n3049 VDD.n3048 0.0101514
R18555 VDD.n3307 VDD.n3306 0.0101514
R18556 VDD.n5630 VDD.n5629 0.0101514
R18557 VDD.n5376 VDD.n5375 0.0101514
R18558 VDD.n3565 VDD.n3564 0.0101514
R18559 VDD.n3823 VDD.n3822 0.0101514
R18560 VDD.n4081 VDD.n4080 0.0101514
R18561 VDD.n4339 VDD.n4338 0.0101514
R18562 VDD.n4597 VDD.n4596 0.0101514
R18563 VDD.n4855 VDD.n4854 0.0101514
R18564 VDD.n5113 VDD.n5112 0.0101514
R18565 VDD.n776 VDD.n775 0.0101053
R18566 VDD.n733 VDD.n732 0.0101053
R18567 VDD.n1126 VDD.n1125 0.0101053
R18568 VDD.n1083 VDD.n1082 0.0101053
R18569 VDD.n1883 VDD.n1882 0.0101
R18570 VDD.n2204 VDD.n2203 0.0101
R18571 VDD.n2462 VDD.n2461 0.0101
R18572 VDD.n2720 VDD.n2719 0.0101
R18573 VDD.n2978 VDD.n2977 0.0101
R18574 VDD.n3236 VDD.n3235 0.0101
R18575 VDD.n3494 VDD.n3493 0.0101
R18576 VDD.n5814 VDD.n5813 0.0101
R18577 VDD.n5560 VDD.n5559 0.0101
R18578 VDD.n3752 VDD.n3751 0.0101
R18579 VDD.n4010 VDD.n4009 0.0101
R18580 VDD.n4268 VDD.n4267 0.0101
R18581 VDD.n4526 VDD.n4525 0.0101
R18582 VDD.n4784 VDD.n4783 0.0101
R18583 VDD.n5042 VDD.n5041 0.0101
R18584 VDD.n5300 VDD.n5299 0.0101
R18585 VDD.n1597 VDD.n1181 0.00985484
R18586 VDD.n137 VDD.n136 0.00984211
R18587 VDD.n2129 VDD.n2128 0.00977468
R18588 VDD.n1884 VDD.n1883 0.0096003
R18589 VDD.n1870 VDD.n1869 0.0096003
R18590 VDD.n1869 VDD.t106 0.0096003
R18591 VDD.n2191 VDD.n2190 0.0096003
R18592 VDD.n2190 VDD.t719 0.0096003
R18593 VDD.n2205 VDD.n2204 0.0096003
R18594 VDD.n2449 VDD.n2448 0.0096003
R18595 VDD.n2448 VDD.t485 0.0096003
R18596 VDD.n2463 VDD.n2462 0.0096003
R18597 VDD.n2707 VDD.n2706 0.0096003
R18598 VDD.n2706 VDD.t531 0.0096003
R18599 VDD.n2721 VDD.n2720 0.0096003
R18600 VDD.n2965 VDD.n2964 0.0096003
R18601 VDD.n2964 VDD.t15 0.0096003
R18602 VDD.n2979 VDD.n2978 0.0096003
R18603 VDD.n3223 VDD.n3222 0.0096003
R18604 VDD.n3222 VDD.t412 0.0096003
R18605 VDD.n3237 VDD.n3236 0.0096003
R18606 VDD.n3481 VDD.n3480 0.0096003
R18607 VDD.n3480 VDD.t538 0.0096003
R18608 VDD.n3495 VDD.n3494 0.0096003
R18609 VDD.n5801 VDD.n5800 0.0096003
R18610 VDD.n5800 VDD.t109 0.0096003
R18611 VDD.n5815 VDD.n5814 0.0096003
R18612 VDD.n5547 VDD.n5546 0.0096003
R18613 VDD.n5546 VDD.t186 0.0096003
R18614 VDD.n5561 VDD.n5560 0.0096003
R18615 VDD.n3739 VDD.n3738 0.0096003
R18616 VDD.n3738 VDD.t413 0.0096003
R18617 VDD.n3753 VDD.n3752 0.0096003
R18618 VDD.n3997 VDD.n3996 0.0096003
R18619 VDD.n3996 VDD.t108 0.0096003
R18620 VDD.n4011 VDD.n4010 0.0096003
R18621 VDD.n4255 VDD.n4254 0.0096003
R18622 VDD.n4254 VDD.t0 0.0096003
R18623 VDD.n4269 VDD.n4268 0.0096003
R18624 VDD.n4513 VDD.n4512 0.0096003
R18625 VDD.n4512 VDD.t13 0.0096003
R18626 VDD.n4527 VDD.n4526 0.0096003
R18627 VDD.n4771 VDD.n4770 0.0096003
R18628 VDD.n4770 VDD.t117 0.0096003
R18629 VDD.n4785 VDD.n4784 0.0096003
R18630 VDD.n5029 VDD.n5028 0.0096003
R18631 VDD.n5028 VDD.t651 0.0096003
R18632 VDD.n5043 VDD.n5042 0.0096003
R18633 VDD.n5287 VDD.n5286 0.0096003
R18634 VDD.n5286 VDD.t85 0.0096003
R18635 VDD.n5301 VDD.n5300 0.0096003
R18636 VDD.t28 VDD.n1891 0.00959985
R18637 VDD.n1891 VDD.n1889 0.00959985
R18638 VDD.t103 VDD.n2212 0.00959985
R18639 VDD.n2212 VDD.n2210 0.00959985
R18640 VDD.t471 VDD.n2470 0.00959985
R18641 VDD.n2470 VDD.n2468 0.00959985
R18642 VDD.t184 VDD.n2728 0.00959985
R18643 VDD.n2728 VDD.n2726 0.00959985
R18644 VDD.t488 VDD.n2986 0.00959985
R18645 VDD.n2986 VDD.n2984 0.00959985
R18646 VDD.t234 VDD.n3244 0.00959985
R18647 VDD.n3244 VDD.n3242 0.00959985
R18648 VDD.t18 VDD.n3502 0.00959985
R18649 VDD.n3502 VDD.n3500 0.00959985
R18650 VDD.t746 VDD.n5822 0.00959985
R18651 VDD.n5822 VDD.n5820 0.00959985
R18652 VDD.t88 VDD.n5568 0.00959985
R18653 VDD.n5568 VDD.n5566 0.00959985
R18654 VDD.t82 VDD.n3760 0.00959985
R18655 VDD.n3760 VDD.n3758 0.00959985
R18656 VDD.t409 VDD.n4018 0.00959985
R18657 VDD.n4018 VDD.n4016 0.00959985
R18658 VDD.t727 VDD.n4276 0.00959985
R18659 VDD.n4276 VDD.n4274 0.00959985
R18660 VDD.t122 VDD.n4534 0.00959985
R18661 VDD.n4534 VDD.n4532 0.00959985
R18662 VDD.t484 VDD.n4792 0.00959985
R18663 VDD.n4792 VDD.n4790 0.00959985
R18664 VDD.t14 VDD.n5050 0.00959985
R18665 VDD.n5050 VDD.n5048 0.00959985
R18666 VDD.t119 VDD.n5308 0.00959985
R18667 VDD.n5308 VDD.n5306 0.00959985
R18668 VDD.n1361 VDD 0.00954255
R18669 VDD.n461 VDD.n458 0.0095362
R18670 VDD.n58 VDD.n55 0.0095362
R18671 VDD.n1425 VDD.n1423 0.0092766
R18672 VDD.n489 VDD.n467 0.00906279
R18673 VDD.n87 VDD.n65 0.00906279
R18674 VDD.n176 VDD.n175 0.00905263
R18675 VDD.n1283 VDD.n1282 0.00883333
R18676 VDD.n1282 VDD.n1280 0.00883333
R18677 VDD.n1280 VDD.n1276 0.00883333
R18678 VDD.n1276 VDD.n1274 0.00883333
R18679 VDD.n1274 VDD.n1270 0.00883333
R18680 VDD.n1295 VDD.n1291 0.00883333
R18681 VDD.n1297 VDD.n1295 0.00883333
R18682 VDD.n1301 VDD.n1297 0.00883333
R18683 VDD.n1303 VDD.n1301 0.00883333
R18684 VDD.n788 VDD.n784 0.00878947
R18685 VDD.n743 VDD.n741 0.00878947
R18686 VDD.n685 VDD.n683 0.00878947
R18687 VDD.n1138 VDD.n1134 0.00878947
R18688 VDD.n1093 VDD.n1091 0.00878947
R18689 VDD.n1035 VDD.n1033 0.00878947
R18690 VDD.n1399 VDD.n1396 0.00874468
R18691 VDD.n577 VDD.n576 0.00852632
R18692 VDD.n590 VDD.n589 0.00852632
R18693 VDD.n635 VDD.n634 0.00852632
R18694 VDD.n927 VDD.n926 0.00852632
R18695 VDD.n940 VDD.n939 0.00852632
R18696 VDD.n985 VDD.n984 0.00852632
R18697 VDD.n2128 VDD.n2127 0.00849839
R18698 VDD.n1287 VDD 0.00847872
R18699 VDD.n1742 VDD.n1741 0.0084202
R18700 VDD.n1699 VDD.n1698 0.0084202
R18701 VDD.n1698 VDD.t642 0.0084202
R18702 VDD.n1676 VDD.n1672 0.0084202
R18703 VDD.n1764 VDD.n1676 0.0084202
R18704 VDD.n1766 VDD.n1765 0.0084202
R18705 VDD.n1765 VDD.n1764 0.0084202
R18706 VDD.n2091 VDD.n2090 0.0084202
R18707 VDD.n2048 VDD.n2047 0.0084202
R18708 VDD.n2047 VDD.t243 0.0084202
R18709 VDD.n2025 VDD.n2021 0.0084202
R18710 VDD.n2113 VDD.n2025 0.0084202
R18711 VDD.n2115 VDD.n2114 0.0084202
R18712 VDD.n2114 VDD.n2113 0.0084202
R18713 VDD.n2321 VDD.n2320 0.0084202
R18714 VDD.n2278 VDD.n2277 0.0084202
R18715 VDD.n2277 VDD.t624 0.0084202
R18716 VDD.n2255 VDD.n2251 0.0084202
R18717 VDD.n2343 VDD.n2255 0.0084202
R18718 VDD.n2345 VDD.n2344 0.0084202
R18719 VDD.n2344 VDD.n2343 0.0084202
R18720 VDD.n2579 VDD.n2578 0.0084202
R18721 VDD.n2536 VDD.n2535 0.0084202
R18722 VDD.n2535 VDD.t842 0.0084202
R18723 VDD.n2513 VDD.n2509 0.0084202
R18724 VDD.n2601 VDD.n2513 0.0084202
R18725 VDD.n2603 VDD.n2602 0.0084202
R18726 VDD.n2602 VDD.n2601 0.0084202
R18727 VDD.n2837 VDD.n2836 0.0084202
R18728 VDD.n2794 VDD.n2793 0.0084202
R18729 VDD.n2793 VDD.t134 0.0084202
R18730 VDD.n2771 VDD.n2767 0.0084202
R18731 VDD.n2859 VDD.n2771 0.0084202
R18732 VDD.n2861 VDD.n2860 0.0084202
R18733 VDD.n2860 VDD.n2859 0.0084202
R18734 VDD.n3095 VDD.n3094 0.0084202
R18735 VDD.n3052 VDD.n3051 0.0084202
R18736 VDD.n3051 VDD.t473 0.0084202
R18737 VDD.n3029 VDD.n3025 0.0084202
R18738 VDD.n3117 VDD.n3029 0.0084202
R18739 VDD.n3119 VDD.n3118 0.0084202
R18740 VDD.n3118 VDD.n3117 0.0084202
R18741 VDD.n3353 VDD.n3352 0.0084202
R18742 VDD.n3310 VDD.n3309 0.0084202
R18743 VDD.n3309 VDD.t1331 0.0084202
R18744 VDD.n3287 VDD.n3283 0.0084202
R18745 VDD.n3375 VDD.n3287 0.0084202
R18746 VDD.n3377 VDD.n3376 0.0084202
R18747 VDD.n3376 VDD.n3375 0.0084202
R18748 VDD.n5676 VDD.n5675 0.0084202
R18749 VDD.n5633 VDD.n5632 0.0084202
R18750 VDD.n5632 VDD.t613 0.0084202
R18751 VDD.n5610 VDD.n5606 0.0084202
R18752 VDD.n5698 VDD.n5610 0.0084202
R18753 VDD.n5700 VDD.n5699 0.0084202
R18754 VDD.n5699 VDD.n5698 0.0084202
R18755 VDD.n5422 VDD.n5421 0.0084202
R18756 VDD.n5379 VDD.n5378 0.0084202
R18757 VDD.n5378 VDD.t6 0.0084202
R18758 VDD.n5356 VDD.n5352 0.0084202
R18759 VDD.n5444 VDD.n5356 0.0084202
R18760 VDD.n5446 VDD.n5445 0.0084202
R18761 VDD.n5445 VDD.n5444 0.0084202
R18762 VDD.n3611 VDD.n3610 0.0084202
R18763 VDD.n3568 VDD.n3567 0.0084202
R18764 VDD.n3567 VDD.t631 0.0084202
R18765 VDD.n3545 VDD.n3541 0.0084202
R18766 VDD.n3633 VDD.n3545 0.0084202
R18767 VDD.n3635 VDD.n3634 0.0084202
R18768 VDD.n3634 VDD.n3633 0.0084202
R18769 VDD.n3869 VDD.n3868 0.0084202
R18770 VDD.n3826 VDD.n3825 0.0084202
R18771 VDD.n3825 VDD.t1386 0.0084202
R18772 VDD.n3803 VDD.n3799 0.0084202
R18773 VDD.n3891 VDD.n3803 0.0084202
R18774 VDD.n3893 VDD.n3892 0.0084202
R18775 VDD.n3892 VDD.n3891 0.0084202
R18776 VDD.n4127 VDD.n4126 0.0084202
R18777 VDD.n4084 VDD.n4083 0.0084202
R18778 VDD.n4083 VDD.t888 0.0084202
R18779 VDD.n4061 VDD.n4057 0.0084202
R18780 VDD.n4149 VDD.n4061 0.0084202
R18781 VDD.n4151 VDD.n4150 0.0084202
R18782 VDD.n4150 VDD.n4149 0.0084202
R18783 VDD.n4385 VDD.n4384 0.0084202
R18784 VDD.n4342 VDD.n4341 0.0084202
R18785 VDD.n4341 VDD.t126 0.0084202
R18786 VDD.n4319 VDD.n4315 0.0084202
R18787 VDD.n4407 VDD.n4319 0.0084202
R18788 VDD.n4409 VDD.n4408 0.0084202
R18789 VDD.n4408 VDD.n4407 0.0084202
R18790 VDD.n4643 VDD.n4642 0.0084202
R18791 VDD.n4600 VDD.n4599 0.0084202
R18792 VDD.n4599 VDD.t72 0.0084202
R18793 VDD.n4577 VDD.n4573 0.0084202
R18794 VDD.n4665 VDD.n4577 0.0084202
R18795 VDD.n4667 VDD.n4666 0.0084202
R18796 VDD.n4666 VDD.n4665 0.0084202
R18797 VDD.n4901 VDD.n4900 0.0084202
R18798 VDD.n4858 VDD.n4857 0.0084202
R18799 VDD.n4857 VDD.t783 0.0084202
R18800 VDD.n4835 VDD.n4831 0.0084202
R18801 VDD.n4923 VDD.n4835 0.0084202
R18802 VDD.n4925 VDD.n4924 0.0084202
R18803 VDD.n4924 VDD.n4923 0.0084202
R18804 VDD.n5159 VDD.n5158 0.0084202
R18805 VDD.n5116 VDD.n5115 0.0084202
R18806 VDD.n5115 VDD.t1374 0.0084202
R18807 VDD.n5093 VDD.n5089 0.0084202
R18808 VDD.n5181 VDD.n5093 0.0084202
R18809 VDD.n5183 VDD.n5182 0.0084202
R18810 VDD.n5182 VDD.n5181 0.0084202
R18811 VDD.n1615 VDD.n1614 0.0083125
R18812 VDD.n383 VDD.n379 0.00826316
R18813 VDD.n338 VDD.n336 0.00826316
R18814 VDD.n280 VDD.n278 0.00826316
R18815 VDD.n1366 VDD.n1365 0.00821277
R18816 VDD.n396 VDD.n395 0.00802802
R18817 VDD.n1554 VDD.n1553 0.00802802
R18818 VDD.n189 VDD.n188 0.008
R18819 VDD.n234 VDD.n233 0.008
R18820 VDD.n260 VDD.n259 0.008
R18821 VDD.n424 VDD.n421 0.00775202
R18822 VDD.n403 VDD.n400 0.00775202
R18823 VDD.n1582 VDD.n1579 0.00775202
R18824 VDD.n1561 VDD.n1558 0.00775202
R18825 VDD.n376 VDD.n375 0.00773684
R18826 VDD.n331 VDD.n330 0.00773684
R18827 VDD.n582 VDD.n540 0.00747368
R18828 VDD.n665 VDD.n664 0.00747368
R18829 VDD.n932 VDD.n890 0.00747368
R18830 VDD.n1015 VDD.n1014 0.00747368
R18831 VDD VDD.n1320 0.00741489
R18832 VDD.n781 VDD.n780 0.00721053
R18833 VDD.n736 VDD.n735 0.00721053
R18834 VDD.n1131 VDD.n1130 0.00721053
R18835 VDD.n1086 VDD.n1085 0.00721053
R18836 VDD.n1543 VDD 0.00714063
R18837 VDD.n1743 VDD.n1742 0.00702894
R18838 VDD.n2092 VDD.n2091 0.00702894
R18839 VDD.n2322 VDD.n2321 0.00702894
R18840 VDD.n2580 VDD.n2579 0.00702894
R18841 VDD.n2838 VDD.n2837 0.00702894
R18842 VDD.n3096 VDD.n3095 0.00702894
R18843 VDD.n3354 VDD.n3353 0.00702894
R18844 VDD.n5677 VDD.n5676 0.00702894
R18845 VDD.n5423 VDD.n5422 0.00702894
R18846 VDD.n3612 VDD.n3611 0.00702894
R18847 VDD.n3870 VDD.n3869 0.00702894
R18848 VDD.n4128 VDD.n4127 0.00702894
R18849 VDD.n4386 VDD.n4385 0.00702894
R18850 VDD.n4644 VDD.n4643 0.00702894
R18851 VDD.n4902 VDD.n4901 0.00702894
R18852 VDD.n5160 VDD.n5159 0.00702894
R18853 VDD.n1291 VDD.n1246 0.00702174
R18854 VDD.n816 VDD 0.00700289
R18855 VDD.n1199 VDD 0.00700289
R18856 VDD.n181 VDD.n139 0.00694737
R18857 VDD.n1829 VDD.n1828 0.00693382
R18858 VDD.n2150 VDD.n2149 0.00693382
R18859 VDD.n2408 VDD.n2407 0.00693382
R18860 VDD.n2666 VDD.n2665 0.00693382
R18861 VDD.n2924 VDD.n2923 0.00693382
R18862 VDD.n3182 VDD.n3181 0.00693382
R18863 VDD.n3440 VDD.n3439 0.00693382
R18864 VDD.n5760 VDD.n5759 0.00693382
R18865 VDD.n5506 VDD.n5505 0.00693382
R18866 VDD.n3698 VDD.n3697 0.00693382
R18867 VDD.n3956 VDD.n3955 0.00693382
R18868 VDD.n4214 VDD.n4213 0.00693382
R18869 VDD.n4472 VDD.n4471 0.00693382
R18870 VDD.n4730 VDD.n4729 0.00693382
R18871 VDD.n4988 VDD.n4987 0.00693382
R18872 VDD.n5246 VDD.n5245 0.00693382
R18873 VDD.n1181 VDD.n1180 0.00681452
R18874 VDD.n809 VDD 0.00675
R18875 VDD.n1192 VDD 0.00675
R18876 VDD.n1540 VDD.n1255 0.00662745
R18877 VDD.n1463 VDD.n1461 0.00661702
R18878 VDD VDD.n551 0.00655263
R18879 VDD.n622 VDD 0.00655263
R18880 VDD VDD.n791 0.00655263
R18881 VDD VDD.n744 0.00655263
R18882 VDD VDD.n697 0.00655263
R18883 VDD.n677 VDD 0.00655263
R18884 VDD VDD.n901 0.00655263
R18885 VDD.n972 VDD 0.00655263
R18886 VDD VDD.n1141 0.00655263
R18887 VDD VDD.n1094 0.00655263
R18888 VDD VDD.n1047 0.00655263
R18889 VDD.n1027 VDD 0.00655263
R18890 VDD VDD.n150 0.00655263
R18891 VDD.n221 VDD 0.00655263
R18892 VDD VDD.n386 0.00655263
R18893 VDD VDD.n339 0.00655263
R18894 VDD VDD.n292 0.00655263
R18895 VDD.n272 VDD 0.00655263
R18896 VDD.n794 VDD.n35 0.00638056
R18897 VDD.n181 VDD.n180 0.00615789
R18898 VDD VDD.n808 0.00609211
R18899 VDD VDD.n1191 0.00609211
R18900 VDD.n1739 VDD.n1736 0.00605556
R18901 VDD.n2088 VDD.n2085 0.00605556
R18902 VDD.n2318 VDD.n2315 0.00605556
R18903 VDD.n2576 VDD.n2573 0.00605556
R18904 VDD.n2834 VDD.n2831 0.00605556
R18905 VDD.n3092 VDD.n3089 0.00605556
R18906 VDD.n3350 VDD.n3347 0.00605556
R18907 VDD.n5673 VDD.n5670 0.00605556
R18908 VDD.n5419 VDD.n5416 0.00605556
R18909 VDD.n3608 VDD.n3605 0.00605556
R18910 VDD.n3866 VDD.n3863 0.00605556
R18911 VDD.n4124 VDD.n4121 0.00605556
R18912 VDD.n4382 VDD.n4379 0.00605556
R18913 VDD.n4640 VDD.n4637 0.00605556
R18914 VDD.n4898 VDD.n4895 0.00605556
R18915 VDD.n5156 VDD.n5153 0.00605556
R18916 VDD.n783 VDD.n781 0.00589474
R18917 VDD.n740 VDD.n736 0.00589474
R18918 VDD.n1133 VDD.n1131 0.00589474
R18919 VDD.n1090 VDD.n1086 0.00589474
R18920 VDD.n1343 VDD.n1320 0.00581915
R18921 VDD.n1982 VDD.n1981 0.00573228
R18922 VDD.n1982 VDD.n1980 0.00573228
R18923 VDD.n1540 VDD.n1539 0.00564706
R18924 VDD.n582 VDD.n581 0.00563158
R18925 VDD.n665 VDD.n637 0.00563158
R18926 VDD.n686 VDD 0.00563158
R18927 VDD.n932 VDD.n931 0.00563158
R18928 VDD.n1015 VDD.n987 0.00563158
R18929 VDD.n1036 VDD 0.00563158
R18930 VDD.n1376 VDD.n1374 0.00552129
R18931 VDD.n1603 VDD.n1602 0.00542857
R18932 VDD.n378 VDD.n376 0.00536842
R18933 VDD.n335 VDD.n331 0.00536842
R18934 VDD.n1617 VDD.n1615 0.0051875
R18935 VDD.n193 VDD.n189 0.00510526
R18936 VDD.n236 VDD.n234 0.00510526
R18937 VDD.n260 VDD.n236 0.00510526
R18938 VDD.n281 VDD 0.00510526
R18939 VDD.n1913 VDD.n1912 0.00505015
R18940 VDD.t28 VDD.n1913 0.00505015
R18941 VDD.t28 VDD.n1894 0.00505015
R18942 VDD.n1909 VDD.n1894 0.00505015
R18943 VDD.n1824 VDD.n1823 0.00505015
R18944 VDD.n1861 VDD.n1848 0.00505015
R18945 VDD.t106 VDD.n1848 0.00505015
R18946 VDD.n1868 VDD.n1867 0.00505015
R18947 VDD.t106 VDD.n1868 0.00505015
R18948 VDD.n2182 VDD.n2169 0.00505015
R18949 VDD.t719 VDD.n2169 0.00505015
R18950 VDD.n2189 VDD.n2188 0.00505015
R18951 VDD.t719 VDD.n2189 0.00505015
R18952 VDD.n2145 VDD.n2144 0.00505015
R18953 VDD.n2234 VDD.n2233 0.00505015
R18954 VDD.t103 VDD.n2234 0.00505015
R18955 VDD.t103 VDD.n2215 0.00505015
R18956 VDD.n2230 VDD.n2215 0.00505015
R18957 VDD.n2440 VDD.n2427 0.00505015
R18958 VDD.t485 VDD.n2427 0.00505015
R18959 VDD.n2447 VDD.n2446 0.00505015
R18960 VDD.t485 VDD.n2447 0.00505015
R18961 VDD.n2403 VDD.n2402 0.00505015
R18962 VDD.n2492 VDD.n2491 0.00505015
R18963 VDD.t471 VDD.n2492 0.00505015
R18964 VDD.t471 VDD.n2473 0.00505015
R18965 VDD.n2488 VDD.n2473 0.00505015
R18966 VDD.n2698 VDD.n2685 0.00505015
R18967 VDD.t531 VDD.n2685 0.00505015
R18968 VDD.n2705 VDD.n2704 0.00505015
R18969 VDD.t531 VDD.n2705 0.00505015
R18970 VDD.n2661 VDD.n2660 0.00505015
R18971 VDD.n2750 VDD.n2749 0.00505015
R18972 VDD.t184 VDD.n2750 0.00505015
R18973 VDD.t184 VDD.n2731 0.00505015
R18974 VDD.n2746 VDD.n2731 0.00505015
R18975 VDD.n2956 VDD.n2943 0.00505015
R18976 VDD.t15 VDD.n2943 0.00505015
R18977 VDD.n2963 VDD.n2962 0.00505015
R18978 VDD.t15 VDD.n2963 0.00505015
R18979 VDD.n2919 VDD.n2918 0.00505015
R18980 VDD.n3008 VDD.n3007 0.00505015
R18981 VDD.t488 VDD.n3008 0.00505015
R18982 VDD.t488 VDD.n2989 0.00505015
R18983 VDD.n3004 VDD.n2989 0.00505015
R18984 VDD.n3214 VDD.n3201 0.00505015
R18985 VDD.t412 VDD.n3201 0.00505015
R18986 VDD.n3221 VDD.n3220 0.00505015
R18987 VDD.t412 VDD.n3221 0.00505015
R18988 VDD.n3177 VDD.n3176 0.00505015
R18989 VDD.n3266 VDD.n3265 0.00505015
R18990 VDD.t234 VDD.n3266 0.00505015
R18991 VDD.t234 VDD.n3247 0.00505015
R18992 VDD.n3262 VDD.n3247 0.00505015
R18993 VDD.n3472 VDD.n3459 0.00505015
R18994 VDD.t538 VDD.n3459 0.00505015
R18995 VDD.n3479 VDD.n3478 0.00505015
R18996 VDD.t538 VDD.n3479 0.00505015
R18997 VDD.n3435 VDD.n3434 0.00505015
R18998 VDD.n3524 VDD.n3523 0.00505015
R18999 VDD.t18 VDD.n3524 0.00505015
R19000 VDD.t18 VDD.n3505 0.00505015
R19001 VDD.n3520 VDD.n3505 0.00505015
R19002 VDD.n5792 VDD.n5779 0.00505015
R19003 VDD.t109 VDD.n5779 0.00505015
R19004 VDD.n5799 VDD.n5798 0.00505015
R19005 VDD.t109 VDD.n5799 0.00505015
R19006 VDD.n5755 VDD.n5754 0.00505015
R19007 VDD.n5844 VDD.n5843 0.00505015
R19008 VDD.t746 VDD.n5844 0.00505015
R19009 VDD.t746 VDD.n5825 0.00505015
R19010 VDD.n5840 VDD.n5825 0.00505015
R19011 VDD.n5538 VDD.n5525 0.00505015
R19012 VDD.t186 VDD.n5525 0.00505015
R19013 VDD.n5545 VDD.n5544 0.00505015
R19014 VDD.t186 VDD.n5545 0.00505015
R19015 VDD.n5501 VDD.n5500 0.00505015
R19016 VDD.n5590 VDD.n5589 0.00505015
R19017 VDD.t88 VDD.n5590 0.00505015
R19018 VDD.t88 VDD.n5571 0.00505015
R19019 VDD.n5586 VDD.n5571 0.00505015
R19020 VDD.n3730 VDD.n3717 0.00505015
R19021 VDD.t413 VDD.n3717 0.00505015
R19022 VDD.n3737 VDD.n3736 0.00505015
R19023 VDD.t413 VDD.n3737 0.00505015
R19024 VDD.n3693 VDD.n3692 0.00505015
R19025 VDD.n3782 VDD.n3781 0.00505015
R19026 VDD.t82 VDD.n3782 0.00505015
R19027 VDD.t82 VDD.n3763 0.00505015
R19028 VDD.n3778 VDD.n3763 0.00505015
R19029 VDD.n3988 VDD.n3975 0.00505015
R19030 VDD.t108 VDD.n3975 0.00505015
R19031 VDD.n3995 VDD.n3994 0.00505015
R19032 VDD.t108 VDD.n3995 0.00505015
R19033 VDD.n3951 VDD.n3950 0.00505015
R19034 VDD.n4040 VDD.n4039 0.00505015
R19035 VDD.t409 VDD.n4040 0.00505015
R19036 VDD.t409 VDD.n4021 0.00505015
R19037 VDD.n4036 VDD.n4021 0.00505015
R19038 VDD.n4246 VDD.n4233 0.00505015
R19039 VDD.t0 VDD.n4233 0.00505015
R19040 VDD.n4253 VDD.n4252 0.00505015
R19041 VDD.t0 VDD.n4253 0.00505015
R19042 VDD.n4209 VDD.n4208 0.00505015
R19043 VDD.n4298 VDD.n4297 0.00505015
R19044 VDD.t727 VDD.n4298 0.00505015
R19045 VDD.t727 VDD.n4279 0.00505015
R19046 VDD.n4294 VDD.n4279 0.00505015
R19047 VDD.n4504 VDD.n4491 0.00505015
R19048 VDD.t13 VDD.n4491 0.00505015
R19049 VDD.n4511 VDD.n4510 0.00505015
R19050 VDD.t13 VDD.n4511 0.00505015
R19051 VDD.n4467 VDD.n4466 0.00505015
R19052 VDD.n4556 VDD.n4555 0.00505015
R19053 VDD.t122 VDD.n4556 0.00505015
R19054 VDD.t122 VDD.n4537 0.00505015
R19055 VDD.n4552 VDD.n4537 0.00505015
R19056 VDD.n4762 VDD.n4749 0.00505015
R19057 VDD.t117 VDD.n4749 0.00505015
R19058 VDD.n4769 VDD.n4768 0.00505015
R19059 VDD.t117 VDD.n4769 0.00505015
R19060 VDD.n4725 VDD.n4724 0.00505015
R19061 VDD.n4814 VDD.n4813 0.00505015
R19062 VDD.t484 VDD.n4814 0.00505015
R19063 VDD.t484 VDD.n4795 0.00505015
R19064 VDD.n4810 VDD.n4795 0.00505015
R19065 VDD.n5020 VDD.n5007 0.00505015
R19066 VDD.t651 VDD.n5007 0.00505015
R19067 VDD.n5027 VDD.n5026 0.00505015
R19068 VDD.t651 VDD.n5027 0.00505015
R19069 VDD.n4983 VDD.n4982 0.00505015
R19070 VDD.n5072 VDD.n5071 0.00505015
R19071 VDD.t14 VDD.n5072 0.00505015
R19072 VDD.t14 VDD.n5053 0.00505015
R19073 VDD.n5068 VDD.n5053 0.00505015
R19074 VDD.n5278 VDD.n5265 0.00505015
R19075 VDD.t85 VDD.n5265 0.00505015
R19076 VDD.n5285 VDD.n5284 0.00505015
R19077 VDD.t85 VDD.n5285 0.00505015
R19078 VDD.n5241 VDD.n5240 0.00505015
R19079 VDD.n5330 VDD.n5329 0.00505015
R19080 VDD.t119 VDD.n5330 0.00505015
R19081 VDD.t119 VDD.n5311 0.00505015
R19082 VDD.n5326 VDD.n5311 0.00505015
R19083 VDD.n1311 VDD 0.00502128
R19084 VDD.n1340 VDD 0.00502128
R19085 VDD VDD.n1346 0.00502128
R19086 VDD.n1363 VDD 0.00502128
R19087 VDD.n1510 VDD 0.00502128
R19088 VDD.n379 VDD.n378 0.00484211
R19089 VDD.n336 VDD.n335 0.00484211
R19090 VDD.n278 VDD.n277 0.00484211
R19091 VDD.n1324 VDD.n1319 0.00475532
R19092 VDD VDD.n1509 0.00475532
R19093 VDD.n1504 VDD.n1261 0.00475532
R19094 VDD.n1287 VDD.n1286 0.00475532
R19095 VDD.n1751 VDD.n1722 0.00466667
R19096 VDD.n1703 VDD.n1702 0.00466667
R19097 VDD.n1692 VDD.n1691 0.00466667
R19098 VDD.n2100 VDD.n2071 0.00466667
R19099 VDD.n2052 VDD.n2051 0.00466667
R19100 VDD.n2041 VDD.n2040 0.00466667
R19101 VDD.n2330 VDD.n2301 0.00466667
R19102 VDD.n2282 VDD.n2281 0.00466667
R19103 VDD.n2271 VDD.n2270 0.00466667
R19104 VDD.n2588 VDD.n2559 0.00466667
R19105 VDD.n2540 VDD.n2539 0.00466667
R19106 VDD.n2529 VDD.n2528 0.00466667
R19107 VDD.n2846 VDD.n2817 0.00466667
R19108 VDD.n2798 VDD.n2797 0.00466667
R19109 VDD.n2787 VDD.n2786 0.00466667
R19110 VDD.n3104 VDD.n3075 0.00466667
R19111 VDD.n3056 VDD.n3055 0.00466667
R19112 VDD.n3045 VDD.n3044 0.00466667
R19113 VDD.n3362 VDD.n3333 0.00466667
R19114 VDD.n3314 VDD.n3313 0.00466667
R19115 VDD.n3303 VDD.n3302 0.00466667
R19116 VDD.n5685 VDD.n5656 0.00466667
R19117 VDD.n5637 VDD.n5636 0.00466667
R19118 VDD.n5626 VDD.n5625 0.00466667
R19119 VDD.n5431 VDD.n5402 0.00466667
R19120 VDD.n5383 VDD.n5382 0.00466667
R19121 VDD.n5372 VDD.n5371 0.00466667
R19122 VDD.n3620 VDD.n3591 0.00466667
R19123 VDD.n3572 VDD.n3571 0.00466667
R19124 VDD.n3561 VDD.n3560 0.00466667
R19125 VDD.n3878 VDD.n3849 0.00466667
R19126 VDD.n3830 VDD.n3829 0.00466667
R19127 VDD.n3819 VDD.n3818 0.00466667
R19128 VDD.n4136 VDD.n4107 0.00466667
R19129 VDD.n4088 VDD.n4087 0.00466667
R19130 VDD.n4077 VDD.n4076 0.00466667
R19131 VDD.n4394 VDD.n4365 0.00466667
R19132 VDD.n4346 VDD.n4345 0.00466667
R19133 VDD.n4335 VDD.n4334 0.00466667
R19134 VDD.n4652 VDD.n4623 0.00466667
R19135 VDD.n4604 VDD.n4603 0.00466667
R19136 VDD.n4593 VDD.n4592 0.00466667
R19137 VDD.n4910 VDD.n4881 0.00466667
R19138 VDD.n4862 VDD.n4861 0.00466667
R19139 VDD.n4851 VDD.n4850 0.00466667
R19140 VDD.n5168 VDD.n5139 0.00466667
R19141 VDD.n5120 VDD.n5119 0.00466667
R19142 VDD.n5109 VDD.n5108 0.00466667
R19143 VDD VDD.n35 0.00460833
R19144 VDD.n581 VDD.n577 0.00457895
R19145 VDD.n594 VDD.n590 0.00457895
R19146 VDD.n637 VDD.n635 0.00457895
R19147 VDD.n931 VDD.n927 0.00457895
R19148 VDD.n944 VDD.n940 0.00457895
R19149 VDD.n987 VDD.n985 0.00457895
R19150 VDD.n1547 VDD.n1546 0.00451563
R19151 VDD.n784 VDD.n783 0.00431579
R19152 VDD.n741 VDD.n740 0.00431579
R19153 VDD.n683 VDD.n682 0.00431579
R19154 VDD.n1134 VDD.n1133 0.00431579
R19155 VDD.n1091 VDD.n1090 0.00431579
R19156 VDD.n1033 VDD.n1032 0.00431579
R19157 VDD.n1406 VDD.n1405 0.0042234
R19158 VDD.n1304 VDD.n1303 0.00412319
R19159 VDD VDD.n809 0.00411272
R19160 VDD VDD.n1192 0.00411272
R19161 VDD.n1611 VDD.n1610 0.00410577
R19162 VDD.n180 VDD.n176 0.00405263
R19163 VDD.n512 VDD 0.00400806
R19164 VDD.n2125 VDD.n2013 0.00390318
R19165 VDD.n809 VDD 0.00378947
R19166 VDD.n1192 VDD 0.00378947
R19167 VDD.n1526 VDD.n1525 0.00369149
R19168 VDD.n1816 VDD.n1809 0.00364862
R19169 VDD.n2137 VDD.n2130 0.00364862
R19170 VDD.n2395 VDD.n2388 0.00364862
R19171 VDD.n2653 VDD.n2646 0.00364862
R19172 VDD.n2911 VDD.n2904 0.00364862
R19173 VDD.n3169 VDD.n3162 0.00364862
R19174 VDD.n3427 VDD.n3420 0.00364862
R19175 VDD.n5747 VDD.n5740 0.00364862
R19176 VDD.n5493 VDD.n5486 0.00364862
R19177 VDD.n3685 VDD.n3678 0.00364862
R19178 VDD.n3943 VDD.n3936 0.00364862
R19179 VDD.n4201 VDD.n4194 0.00364862
R19180 VDD.n4459 VDD.n4452 0.00364862
R19181 VDD.n4717 VDD.n4710 0.00364862
R19182 VDD.n4975 VDD.n4968 0.00364862
R19183 VDD.n5233 VDD.n5226 0.00364862
R19184 VDD.n1289 VDD 0.00342553
R19185 VDD.n1609 VDD.n1604 0.00339649
R19186 VDD VDD.n796 0.00330645
R19187 VDD.n139 VDD.n137 0.00326316
R19188 VDD.n1934 VDD.n1926 0.00317113
R19189 VDD.n1955 VDD.n1944 0.00317113
R19190 VDD.n1359 VDD.n1358 0.00315957
R19191 VDD.n1600 VDD 0.00304286
R19192 VDD.n780 VDD.n776 0.003
R19193 VDD.n735 VDD.n733 0.003
R19194 VDD.n1130 VDD.n1126 0.003
R19195 VDD.n1085 VDD.n1083 0.003
R19196 VDD.n1743 VDD.t1359 0.00289124
R19197 VDD.n2092 VDD.t1493 0.00289124
R19198 VDD.n2322 VDD.t222 0.00289124
R19199 VDD.n2580 VDD.t55 0.00289124
R19200 VDD.n2838 VDD.t595 0.00289124
R19201 VDD.n3096 VDD.t41 0.00289124
R19202 VDD.n3354 VDD.t731 0.00289124
R19203 VDD.n5677 VDD.t164 0.00289124
R19204 VDD.n5423 VDD.t517 0.00289124
R19205 VDD.n3612 VDD.t194 0.00289124
R19206 VDD.n3870 VDD.t173 0.00289124
R19207 VDD.n4128 VDD.t92 0.00289124
R19208 VDD.n4386 VDD.t497 0.00289124
R19209 VDD.n4644 VDD.t587 0.00289124
R19210 VDD.n4902 VDD.t579 0.00289124
R19211 VDD.n5160 VDD.t857 0.00289124
R19212 VDD.n540 VDD.n538 0.00273684
R19213 VDD.n552 VDD 0.00273684
R19214 VDD.n619 VDD 0.00273684
R19215 VDD.n664 VDD.n660 0.00273684
R19216 VDD.n792 VDD 0.00273684
R19217 VDD.n745 VDD 0.00273684
R19218 VDD.n698 VDD 0.00273684
R19219 VDD.n680 VDD 0.00273684
R19220 VDD.n890 VDD.n888 0.00273684
R19221 VDD.n902 VDD 0.00273684
R19222 VDD.n969 VDD 0.00273684
R19223 VDD.n1014 VDD.n1010 0.00273684
R19224 VDD.n1142 VDD 0.00273684
R19225 VDD.n1095 VDD 0.00273684
R19226 VDD.n1048 VDD 0.00273684
R19227 VDD.n1030 VDD 0.00273684
R19228 VDD.n151 VDD 0.00273684
R19229 VDD.n218 VDD 0.00273684
R19230 VDD.n387 VDD 0.00273684
R19231 VDD.n340 VDD 0.00273684
R19232 VDD.n293 VDD 0.00273684
R19233 VDD.n275 VDD 0.00273684
R19234 VDD.n188 VDD.n186 0.00271053
R19235 VDD.n1926 VDD.n1925 0.00267116
R19236 VDD.n1956 VDD.n1955 0.00267116
R19237 VDD.n1506 VDD 0.00262766
R19238 VDD.n689 VDD.n688 0.00247368
R19239 VDD.n1039 VDD.n1038 0.00247368
R19240 VDD.n375 VDD.n371 0.00247368
R19241 VDD.n330 VDD.n328 0.00247368
R19242 VDD.n5859 VDD.n5858 0.00240789
R19243 VDD.n1838 VDD.n1837 0.00240766
R19244 VDD.n2159 VDD.n2158 0.00240766
R19245 VDD.n2417 VDD.n2416 0.00240766
R19246 VDD.n2675 VDD.n2674 0.00240766
R19247 VDD.n2933 VDD.n2932 0.00240766
R19248 VDD.n3191 VDD.n3190 0.00240766
R19249 VDD.n3449 VDD.n3448 0.00240766
R19250 VDD.n5769 VDD.n5768 0.00240766
R19251 VDD.n5515 VDD.n5514 0.00240766
R19252 VDD.n3707 VDD.n3706 0.00240766
R19253 VDD.n3965 VDD.n3964 0.00240766
R19254 VDD.n4223 VDD.n4222 0.00240766
R19255 VDD.n4481 VDD.n4480 0.00240766
R19256 VDD.n4739 VDD.n4738 0.00240766
R19257 VDD.n4997 VDD.n4996 0.00240766
R19258 VDD.n5255 VDD.n5254 0.00240766
R19259 VDD.n1601 VDD.n1600 0.00237143
R19260 VDD.n1359 VDD 0.0023617
R19261 VDD.n1369 VDD.n1368 0.0023617
R19262 VDD.n1829 VDD.n1825 0.00233824
R19263 VDD.n1831 VDD 0.00233824
R19264 VDD.n2150 VDD.n2146 0.00233824
R19265 VDD.n2152 VDD 0.00233824
R19266 VDD.n2408 VDD.n2404 0.00233824
R19267 VDD.n2410 VDD 0.00233824
R19268 VDD.n2666 VDD.n2662 0.00233824
R19269 VDD.n2668 VDD 0.00233824
R19270 VDD.n2924 VDD.n2920 0.00233824
R19271 VDD.n2926 VDD 0.00233824
R19272 VDD.n3182 VDD.n3178 0.00233824
R19273 VDD.n3184 VDD 0.00233824
R19274 VDD.n3440 VDD.n3436 0.00233824
R19275 VDD.n3442 VDD 0.00233824
R19276 VDD.n5760 VDD.n5756 0.00233824
R19277 VDD.n5762 VDD 0.00233824
R19278 VDD.n5506 VDD.n5502 0.00233824
R19279 VDD.n5508 VDD 0.00233824
R19280 VDD.n3698 VDD.n3694 0.00233824
R19281 VDD.n3700 VDD 0.00233824
R19282 VDD.n3956 VDD.n3952 0.00233824
R19283 VDD.n3958 VDD 0.00233824
R19284 VDD.n4214 VDD.n4210 0.00233824
R19285 VDD.n4216 VDD 0.00233824
R19286 VDD.n4472 VDD.n4468 0.00233824
R19287 VDD.n4474 VDD 0.00233824
R19288 VDD.n4730 VDD.n4726 0.00233824
R19289 VDD.n4732 VDD 0.00233824
R19290 VDD.n4988 VDD.n4984 0.00233824
R19291 VDD.n4990 VDD 0.00233824
R19292 VDD.n5246 VDD.n5242 0.00233824
R19293 VDD.n5248 VDD 0.00233824
R19294 VDD.n1454 VDD.n1317 0.00232979
R19295 VDD.n1431 VDD.n1319 0.00232979
R19296 VDD.n1879 VDD.t528 0.00231811
R19297 VDD.n2200 VDD.t481 0.00231811
R19298 VDD.n2458 VDD.t118 0.00231811
R19299 VDD.n2716 VDD.t652 0.00231811
R19300 VDD.n2974 VDD.t12 0.00231811
R19301 VDD.n3232 VDD.t718 0.00231811
R19302 VDD.n3490 VDD.t411 0.00231811
R19303 VDD.n5810 VDD.t530 0.00231811
R19304 VDD.n5556 VDD.t482 0.00231811
R19305 VDD.n3748 VDD.t410 0.00231811
R19306 VDD.n4006 VDD.t116 0.00231811
R19307 VDD.n4264 VDD.t489 0.00231811
R19308 VDD.n4522 VDD.t84 0.00231811
R19309 VDD.n4780 VDD.t717 0.00231811
R19310 VDD.n5038 VDD.t1353 0.00231811
R19311 VDD.n5296 VDD.t529 0.00231811
R19312 VDD.n1270 VDD.n1246 0.00231159
R19313 VDD.n1726 VDD.n1724 0.00228571
R19314 VDD.n2075 VDD.n2073 0.00228571
R19315 VDD.n2305 VDD.n2303 0.00228571
R19316 VDD.n2563 VDD.n2561 0.00228571
R19317 VDD.n2821 VDD.n2819 0.00228571
R19318 VDD.n3079 VDD.n3077 0.00228571
R19319 VDD.n3337 VDD.n3335 0.00228571
R19320 VDD.n5660 VDD.n5658 0.00228571
R19321 VDD.n5406 VDD.n5404 0.00228571
R19322 VDD.n3595 VDD.n3593 0.00228571
R19323 VDD.n3853 VDD.n3851 0.00228571
R19324 VDD.n4111 VDD.n4109 0.00228571
R19325 VDD.n4369 VDD.n4367 0.00228571
R19326 VDD.n4627 VDD.n4625 0.00228571
R19327 VDD.n4885 VDD.n4883 0.00228571
R19328 VDD.n5143 VDD.n5141 0.00228571
R19329 VDD.n1694 VDD.n1693 0.00221302
R19330 VDD.n1695 VDD.n1694 0.00221302
R19331 VDD.n2043 VDD.n2042 0.00221302
R19332 VDD.n2044 VDD.n2043 0.00221302
R19333 VDD.n2273 VDD.n2272 0.00221302
R19334 VDD.n2274 VDD.n2273 0.00221302
R19335 VDD.n2531 VDD.n2530 0.00221302
R19336 VDD.n2532 VDD.n2531 0.00221302
R19337 VDD.n2789 VDD.n2788 0.00221302
R19338 VDD.n2790 VDD.n2789 0.00221302
R19339 VDD.n3047 VDD.n3046 0.00221302
R19340 VDD.n3048 VDD.n3047 0.00221302
R19341 VDD.n3305 VDD.n3304 0.00221302
R19342 VDD.n3306 VDD.n3305 0.00221302
R19343 VDD.n5628 VDD.n5627 0.00221302
R19344 VDD.n5629 VDD.n5628 0.00221302
R19345 VDD.n5374 VDD.n5373 0.00221302
R19346 VDD.n5375 VDD.n5374 0.00221302
R19347 VDD.n3563 VDD.n3562 0.00221302
R19348 VDD.n3564 VDD.n3563 0.00221302
R19349 VDD.n3821 VDD.n3820 0.00221302
R19350 VDD.n3822 VDD.n3821 0.00221302
R19351 VDD.n4079 VDD.n4078 0.00221302
R19352 VDD.n4080 VDD.n4079 0.00221302
R19353 VDD.n4337 VDD.n4336 0.00221302
R19354 VDD.n4338 VDD.n4337 0.00221302
R19355 VDD.n4595 VDD.n4594 0.00221302
R19356 VDD.n4596 VDD.n4595 0.00221302
R19357 VDD.n4853 VDD.n4852 0.00221302
R19358 VDD.n4854 VDD.n4853 0.00221302
R19359 VDD.n5111 VDD.n5110 0.00221302
R19360 VDD.n5112 VDD.n5111 0.00221302
R19361 VDD.n1693 VDD.n1692 0.00221271
R19362 VDD.n2042 VDD.n2041 0.00221271
R19363 VDD.n2272 VDD.n2271 0.00221271
R19364 VDD.n2530 VDD.n2529 0.00221271
R19365 VDD.n2788 VDD.n2787 0.00221271
R19366 VDD.n3046 VDD.n3045 0.00221271
R19367 VDD.n3304 VDD.n3303 0.00221271
R19368 VDD.n5627 VDD.n5626 0.00221271
R19369 VDD.n5373 VDD.n5372 0.00221271
R19370 VDD.n3562 VDD.n3561 0.00221271
R19371 VDD.n3820 VDD.n3819 0.00221271
R19372 VDD.n4078 VDD.n4077 0.00221271
R19373 VDD.n4336 VDD.n4335 0.00221271
R19374 VDD.n4594 VDD.n4593 0.00221271
R19375 VDD.n4852 VDD.n4851 0.00221271
R19376 VDD.n5110 VDD.n5109 0.00221271
R19377 VDD.n259 VDD.n255 0.00221053
R19378 VDD.n1732 VDD.n1730 0.00220611
R19379 VDD.n2081 VDD.n2079 0.00220611
R19380 VDD.n2311 VDD.n2309 0.00220611
R19381 VDD.n2569 VDD.n2567 0.00220611
R19382 VDD.n2827 VDD.n2825 0.00220611
R19383 VDD.n3085 VDD.n3083 0.00220611
R19384 VDD.n3343 VDD.n3341 0.00220611
R19385 VDD.n5666 VDD.n5664 0.00220611
R19386 VDD.n5412 VDD.n5410 0.00220611
R19387 VDD.n3601 VDD.n3599 0.00220611
R19388 VDD.n3859 VDD.n3857 0.00220611
R19389 VDD.n4117 VDD.n4115 0.00220611
R19390 VDD.n4375 VDD.n4373 0.00220611
R19391 VDD.n4633 VDD.n4631 0.00220611
R19392 VDD.n4891 VDD.n4889 0.00220611
R19393 VDD.n5149 VDD.n5147 0.00220611
R19394 VDD.n1702 VDD.n1681 0.0022058
R19395 VDD.n2051 VDD.n2030 0.0022058
R19396 VDD.n2281 VDD.n2260 0.0022058
R19397 VDD.n2539 VDD.n2518 0.0022058
R19398 VDD.n2797 VDD.n2776 0.0022058
R19399 VDD.n3055 VDD.n3034 0.0022058
R19400 VDD.n3313 VDD.n3292 0.0022058
R19401 VDD.n5636 VDD.n5615 0.0022058
R19402 VDD.n5382 VDD.n5361 0.0022058
R19403 VDD.n3571 VDD.n3550 0.0022058
R19404 VDD.n3829 VDD.n3808 0.0022058
R19405 VDD.n4087 VDD.n4066 0.0022058
R19406 VDD.n4345 VDD.n4324 0.0022058
R19407 VDD.n4603 VDD.n4582 0.0022058
R19408 VDD.n4861 VDD.n4840 0.0022058
R19409 VDD.n5119 VDD.n5098 0.0022058
R19410 VDD.n1745 VDD.n1724 0.0022058
R19411 VDD.n2094 VDD.n2073 0.0022058
R19412 VDD.n2324 VDD.n2303 0.0022058
R19413 VDD.n2582 VDD.n2561 0.0022058
R19414 VDD.n2840 VDD.n2819 0.0022058
R19415 VDD.n3098 VDD.n3077 0.0022058
R19416 VDD.n3356 VDD.n3335 0.0022058
R19417 VDD.n5679 VDD.n5658 0.0022058
R19418 VDD.n5425 VDD.n5404 0.0022058
R19419 VDD.n3614 VDD.n3593 0.0022058
R19420 VDD.n3872 VDD.n3851 0.0022058
R19421 VDD.n4130 VDD.n4109 0.0022058
R19422 VDD.n4388 VDD.n4367 0.0022058
R19423 VDD.n4646 VDD.n4625 0.0022058
R19424 VDD.n4904 VDD.n4883 0.0022058
R19425 VDD.n5162 VDD.n5141 0.0022058
R19426 VDD.n589 VDD.n587 0.00218421
R19427 VDD.n939 VDD.n937 0.00218421
R19428 VDD.n1745 VDD.n1744 0.00212475
R19429 VDD.n1681 VDD.n1678 0.00212475
R19430 VDD.n1732 VDD.n1712 0.00212475
R19431 VDD.n2094 VDD.n2093 0.00212475
R19432 VDD.n2030 VDD.n2027 0.00212475
R19433 VDD.n2081 VDD.n2061 0.00212475
R19434 VDD.n2324 VDD.n2323 0.00212475
R19435 VDD.n2260 VDD.n2257 0.00212475
R19436 VDD.n2311 VDD.n2291 0.00212475
R19437 VDD.n2582 VDD.n2581 0.00212475
R19438 VDD.n2518 VDD.n2515 0.00212475
R19439 VDD.n2569 VDD.n2549 0.00212475
R19440 VDD.n2840 VDD.n2839 0.00212475
R19441 VDD.n2776 VDD.n2773 0.00212475
R19442 VDD.n2827 VDD.n2807 0.00212475
R19443 VDD.n3098 VDD.n3097 0.00212475
R19444 VDD.n3034 VDD.n3031 0.00212475
R19445 VDD.n3085 VDD.n3065 0.00212475
R19446 VDD.n3356 VDD.n3355 0.00212475
R19447 VDD.n3292 VDD.n3289 0.00212475
R19448 VDD.n3343 VDD.n3323 0.00212475
R19449 VDD.n5679 VDD.n5678 0.00212475
R19450 VDD.n5615 VDD.n5612 0.00212475
R19451 VDD.n5666 VDD.n5646 0.00212475
R19452 VDD.n5425 VDD.n5424 0.00212475
R19453 VDD.n5361 VDD.n5358 0.00212475
R19454 VDD.n5412 VDD.n5392 0.00212475
R19455 VDD.n3614 VDD.n3613 0.00212475
R19456 VDD.n3550 VDD.n3547 0.00212475
R19457 VDD.n3601 VDD.n3581 0.00212475
R19458 VDD.n3872 VDD.n3871 0.00212475
R19459 VDD.n3808 VDD.n3805 0.00212475
R19460 VDD.n3859 VDD.n3839 0.00212475
R19461 VDD.n4130 VDD.n4129 0.00212475
R19462 VDD.n4066 VDD.n4063 0.00212475
R19463 VDD.n4117 VDD.n4097 0.00212475
R19464 VDD.n4388 VDD.n4387 0.00212475
R19465 VDD.n4324 VDD.n4321 0.00212475
R19466 VDD.n4375 VDD.n4355 0.00212475
R19467 VDD.n4646 VDD.n4645 0.00212475
R19468 VDD.n4582 VDD.n4579 0.00212475
R19469 VDD.n4633 VDD.n4613 0.00212475
R19470 VDD.n4904 VDD.n4903 0.00212475
R19471 VDD.n4840 VDD.n4837 0.00212475
R19472 VDD.n4891 VDD.n4871 0.00212475
R19473 VDD.n5162 VDD.n5161 0.00212475
R19474 VDD.n5098 VDD.n5095 0.00212475
R19475 VDD.n5149 VDD.n5129 0.00212475
R19476 VDD VDD.n1599 0.00202016
R19477 VDD.n22 VDD.n3 0.00195349
R19478 VDD.n21 VDD.n4 0.00195349
R19479 VDD.n17 VDD.n16 0.00195349
R19480 VDD.n15 VDD.n14 0.00195349
R19481 VDD.n11 VDD.n10 0.00195349
R19482 VDD.n1166 VDD.n1147 0.00195349
R19483 VDD.n1165 VDD.n1148 0.00195349
R19484 VDD.n1161 VDD.n1160 0.00195349
R19485 VDD.n1159 VDD.n1158 0.00195349
R19486 VDD.n1155 VDD.n1154 0.00195349
R19487 VDD.n284 VDD.n283 0.00194737
R19488 VDD.n281 VDD.n280 0.00194737
R19489 VDD.n1757 VDD.n1756 0.00194704
R19490 VDD.n2106 VDD.n2105 0.00194704
R19491 VDD.n2336 VDD.n2335 0.00194704
R19492 VDD.n2594 VDD.n2593 0.00194704
R19493 VDD.n2852 VDD.n2851 0.00194704
R19494 VDD.n3110 VDD.n3109 0.00194704
R19495 VDD.n3368 VDD.n3367 0.00194704
R19496 VDD.n5691 VDD.n5690 0.00194704
R19497 VDD.n5437 VDD.n5436 0.00194704
R19498 VDD.n3626 VDD.n3625 0.00194704
R19499 VDD.n3884 VDD.n3883 0.00194704
R19500 VDD.n4142 VDD.n4141 0.00194704
R19501 VDD.n4400 VDD.n4399 0.00194704
R19502 VDD.n4658 VDD.n4657 0.00194704
R19503 VDD.n4916 VDD.n4915 0.00194704
R19504 VDD.n5174 VDD.n5173 0.00194704
R19505 VDD.n795 VDD.n794 0.00190323
R19506 VDD.n1735 VDD.n1730 0.00188889
R19507 VDD.n2084 VDD.n2079 0.00188889
R19508 VDD.n2314 VDD.n2309 0.00188889
R19509 VDD.n2572 VDD.n2567 0.00188889
R19510 VDD.n2830 VDD.n2825 0.00188889
R19511 VDD.n3088 VDD.n3083 0.00188889
R19512 VDD.n3346 VDD.n3341 0.00188889
R19513 VDD.n5669 VDD.n5664 0.00188889
R19514 VDD.n5415 VDD.n5410 0.00188889
R19515 VDD.n3604 VDD.n3599 0.00188889
R19516 VDD.n3862 VDD.n3857 0.00188889
R19517 VDD.n4120 VDD.n4115 0.00188889
R19518 VDD.n4378 VDD.n4373 0.00188889
R19519 VDD.n4636 VDD.n4631 0.00188889
R19520 VDD.n4894 VDD.n4889 0.00188889
R19521 VDD.n5152 VDD.n5147 0.00188889
R19522 VDD.n1426 VDD.n1345 0.00182979
R19523 VDD.n1401 VDD.n1399 0.00182979
R19524 VDD.n1369 VDD.n1361 0.00182979
R19525 VDD.n1509 VDD.n1506 0.00182979
R19526 VDD.n1459 VDD.n1289 0.00182979
R19527 VDD.n1599 VDD.n1598 0.00178629
R19528 VDD.n1803 VDD.n1777 0.00175592
R19529 VDD.n1802 VDD.n1777 0.00175592
R19530 VDD.n2011 VDD.n1985 0.00175592
R19531 VDD.n2010 VDD.n1985 0.00175592
R19532 VDD.n2382 VDD.n2356 0.00175592
R19533 VDD.n2381 VDD.n2356 0.00175592
R19534 VDD.n2640 VDD.n2614 0.00175592
R19535 VDD.n2639 VDD.n2614 0.00175592
R19536 VDD.n2898 VDD.n2872 0.00175592
R19537 VDD.n2897 VDD.n2872 0.00175592
R19538 VDD.n3156 VDD.n3130 0.00175592
R19539 VDD.n3155 VDD.n3130 0.00175592
R19540 VDD.n3414 VDD.n3388 0.00175592
R19541 VDD.n3413 VDD.n3388 0.00175592
R19542 VDD.n5737 VDD.n5711 0.00175592
R19543 VDD.n5736 VDD.n5711 0.00175592
R19544 VDD.n5483 VDD.n5457 0.00175592
R19545 VDD.n5482 VDD.n5457 0.00175592
R19546 VDD.n3672 VDD.n3646 0.00175592
R19547 VDD.n3671 VDD.n3646 0.00175592
R19548 VDD.n3930 VDD.n3904 0.00175592
R19549 VDD.n3929 VDD.n3904 0.00175592
R19550 VDD.n4188 VDD.n4162 0.00175592
R19551 VDD.n4187 VDD.n4162 0.00175592
R19552 VDD.n4446 VDD.n4420 0.00175592
R19553 VDD.n4445 VDD.n4420 0.00175592
R19554 VDD.n4704 VDD.n4678 0.00175592
R19555 VDD.n4703 VDD.n4678 0.00175592
R19556 VDD.n4962 VDD.n4936 0.00175592
R19557 VDD.n4961 VDD.n4936 0.00175592
R19558 VDD.n5220 VDD.n5194 0.00175592
R19559 VDD.n5219 VDD.n5194 0.00175592
R19560 VDD.n1838 VDD.n1825 0.00162613
R19561 VDD.n2159 VDD.n2146 0.00162613
R19562 VDD.n2417 VDD.n2404 0.00162613
R19563 VDD.n2675 VDD.n2662 0.00162613
R19564 VDD.n2933 VDD.n2920 0.00162613
R19565 VDD.n3191 VDD.n3178 0.00162613
R19566 VDD.n3449 VDD.n3436 0.00162613
R19567 VDD.n5769 VDD.n5756 0.00162613
R19568 VDD.n5515 VDD.n5502 0.00162613
R19569 VDD.n3707 VDD.n3694 0.00162613
R19570 VDD.n3965 VDD.n3952 0.00162613
R19571 VDD.n4223 VDD.n4210 0.00162613
R19572 VDD.n4481 VDD.n4468 0.00162613
R19573 VDD.n4739 VDD.n4726 0.00162613
R19574 VDD.n4997 VDD.n4984 0.00162613
R19575 VDD.n5255 VDD.n5242 0.00162613
R19576 VDD.n1921 VDD.n1664 0.00162258
R19577 VDD.n2242 VDD.n1983 0.00162258
R19578 VDD.n2500 VDD.n2243 0.00162258
R19579 VDD.n2758 VDD.n2501 0.00162258
R19580 VDD.n3016 VDD.n2759 0.00162258
R19581 VDD.n3274 VDD.n3017 0.00162258
R19582 VDD.n3532 VDD.n3275 0.00162258
R19583 VDD.n3790 VDD.n3533 0.00162258
R19584 VDD.n4048 VDD.n3791 0.00162258
R19585 VDD.n4306 VDD.n4049 0.00162258
R19586 VDD.n4564 VDD.n4307 0.00162258
R19587 VDD.n4822 VDD.n4565 0.00162258
R19588 VDD.n5080 VDD.n4823 0.00162258
R19589 VDD.n5338 VDD.n5081 0.00162258
R19590 VDD.n1815 VDD.n1810 0.00161113
R19591 VDD.n2136 VDD.n2131 0.00161113
R19592 VDD.n2394 VDD.n2389 0.00161113
R19593 VDD.n2652 VDD.n2647 0.00161113
R19594 VDD.n2910 VDD.n2905 0.00161113
R19595 VDD.n3168 VDD.n3163 0.00161113
R19596 VDD.n3426 VDD.n3421 0.00161113
R19597 VDD.n5746 VDD.n5741 0.00161113
R19598 VDD.n5492 VDD.n5487 0.00161113
R19599 VDD.n3684 VDD.n3679 0.00161113
R19600 VDD.n3942 VDD.n3937 0.00161113
R19601 VDD.n4200 VDD.n4195 0.00161113
R19602 VDD.n4458 VDD.n4453 0.00161113
R19603 VDD.n4716 VDD.n4711 0.00161113
R19604 VDD.n4974 VDD.n4969 0.00161113
R19605 VDD.n5232 VDD.n5227 0.00161113
R19606 VDD.n1808 VDD.n1664 0.00160808
R19607 VDD.n2129 VDD.n1983 0.00160808
R19608 VDD.n2387 VDD.n2243 0.00160808
R19609 VDD.n2645 VDD.n2501 0.00160808
R19610 VDD.n2903 VDD.n2759 0.00160808
R19611 VDD.n3161 VDD.n3017 0.00160808
R19612 VDD.n3419 VDD.n3275 0.00160808
R19613 VDD.n3677 VDD.n3533 0.00160808
R19614 VDD.n3935 VDD.n3791 0.00160808
R19615 VDD.n4193 VDD.n4049 0.00160808
R19616 VDD.n4451 VDD.n4307 0.00160808
R19617 VDD.n4709 VDD.n4565 0.00160808
R19618 VDD.n4967 VDD.n4823 0.00160808
R19619 VDD.n5225 VDD.n5081 0.00160808
R19620 VDD.n1949 VDD.n1942 0.00158558
R19621 VDD.n1931 VDD.n1930 0.00158558
R19622 VDD.n1807 VDD.n1775 0.00157581
R19623 VDD.n2127 VDD.n2124 0.00157581
R19624 VDD.n2386 VDD.n2354 0.00157581
R19625 VDD.n2644 VDD.n2612 0.00157581
R19626 VDD.n2902 VDD.n2870 0.00157581
R19627 VDD.n3160 VDD.n3128 0.00157581
R19628 VDD.n3418 VDD.n3386 0.00157581
R19629 VDD.n3676 VDD.n3644 0.00157581
R19630 VDD.n3934 VDD.n3902 0.00157581
R19631 VDD.n4192 VDD.n4160 0.00157581
R19632 VDD.n4450 VDD.n4418 0.00157581
R19633 VDD.n4708 VDD.n4676 0.00157581
R19634 VDD.n4966 VDD.n4934 0.00157581
R19635 VDD.n5224 VDD.n5192 0.00157581
R19636 VDD.n1801 VDD.n1800 0.00151809
R19637 VDD.n2009 VDD.n2008 0.00151809
R19638 VDD.n2380 VDD.n2379 0.00151809
R19639 VDD.n2638 VDD.n2637 0.00151809
R19640 VDD.n2896 VDD.n2895 0.00151809
R19641 VDD.n3154 VDD.n3153 0.00151809
R19642 VDD.n3412 VDD.n3411 0.00151809
R19643 VDD.n5735 VDD.n5734 0.00151809
R19644 VDD.n5481 VDD.n5480 0.00151809
R19645 VDD.n3670 VDD.n3669 0.00151809
R19646 VDD.n3928 VDD.n3927 0.00151809
R19647 VDD.n4186 VDD.n4185 0.00151809
R19648 VDD.n4444 VDD.n4443 0.00151809
R19649 VDD.n4702 VDD.n4701 0.00151809
R19650 VDD.n4960 VDD.n4959 0.00151809
R19651 VDD.n5218 VDD.n5217 0.00151809
R19652 VDD.n1801 VDD.n1777 0.00149567
R19653 VDD.n2009 VDD.n1985 0.00149567
R19654 VDD.n2380 VDD.n2356 0.00149567
R19655 VDD.n2638 VDD.n2614 0.00149567
R19656 VDD.n2896 VDD.n2872 0.00149567
R19657 VDD.n3154 VDD.n3130 0.00149567
R19658 VDD.n3412 VDD.n3388 0.00149567
R19659 VDD.n5735 VDD.n5711 0.00149567
R19660 VDD.n5481 VDD.n5457 0.00149567
R19661 VDD.n3670 VDD.n3646 0.00149567
R19662 VDD.n3928 VDD.n3904 0.00149567
R19663 VDD.n4186 VDD.n4162 0.00149567
R19664 VDD.n4444 VDD.n4420 0.00149567
R19665 VDD.n4702 VDD.n4678 0.00149567
R19666 VDD.n4960 VDD.n4936 0.00149567
R19667 VDD.n5218 VDD.n5194 0.00149567
R19668 VDD.n1917 VDD.n1916 0.00148913
R19669 VDD.n2238 VDD.n2237 0.00148913
R19670 VDD.n2496 VDD.n2495 0.00148913
R19671 VDD.n2754 VDD.n2753 0.00148913
R19672 VDD.n3012 VDD.n3011 0.00148913
R19673 VDD.n3270 VDD.n3269 0.00148913
R19674 VDD.n3528 VDD.n3527 0.00148913
R19675 VDD.n5848 VDD.n5847 0.00148913
R19676 VDD.n5594 VDD.n5593 0.00148913
R19677 VDD.n3786 VDD.n3785 0.00148913
R19678 VDD.n4044 VDD.n4043 0.00148913
R19679 VDD.n4302 VDD.n4301 0.00148913
R19680 VDD.n4560 VDD.n4559 0.00148913
R19681 VDD.n4818 VDD.n4817 0.00148913
R19682 VDD.n5076 VDD.n5075 0.00148913
R19683 VDD.n5334 VDD.n5333 0.00148913
R19684 VDD.n1602 VDD.n1601 0.00147143
R19685 VDD.n1806 VDD.n1805 0.00147065
R19686 VDD.n2126 VDD.n2125 0.00147065
R19687 VDD.n2385 VDD.n2384 0.00147065
R19688 VDD.n2643 VDD.n2642 0.00147065
R19689 VDD.n2901 VDD.n2900 0.00147065
R19690 VDD.n3159 VDD.n3158 0.00147065
R19691 VDD.n3417 VDD.n3416 0.00147065
R19692 VDD.n3675 VDD.n3674 0.00147065
R19693 VDD.n3933 VDD.n3932 0.00147065
R19694 VDD.n4191 VDD.n4190 0.00147065
R19695 VDD.n4449 VDD.n4448 0.00147065
R19696 VDD.n4707 VDD.n4706 0.00147065
R19697 VDD.n4965 VDD.n4964 0.00147065
R19698 VDD.n5223 VDD.n5222 0.00147065
R19699 VDD.n1769 VDD.n1670 0.00145131
R19700 VDD.n1711 VDD.n1670 0.00145131
R19701 VDD.n2118 VDD.n2019 0.00145131
R19702 VDD.n2060 VDD.n2019 0.00145131
R19703 VDD.n2348 VDD.n2249 0.00145131
R19704 VDD.n2290 VDD.n2249 0.00145131
R19705 VDD.n2606 VDD.n2507 0.00145131
R19706 VDD.n2548 VDD.n2507 0.00145131
R19707 VDD.n2864 VDD.n2765 0.00145131
R19708 VDD.n2806 VDD.n2765 0.00145131
R19709 VDD.n3122 VDD.n3023 0.00145131
R19710 VDD.n3064 VDD.n3023 0.00145131
R19711 VDD.n3380 VDD.n3281 0.00145131
R19712 VDD.n3322 VDD.n3281 0.00145131
R19713 VDD.n5703 VDD.n5604 0.00145131
R19714 VDD.n5645 VDD.n5604 0.00145131
R19715 VDD.n5449 VDD.n5350 0.00145131
R19716 VDD.n5391 VDD.n5350 0.00145131
R19717 VDD.n3638 VDD.n3539 0.00145131
R19718 VDD.n3580 VDD.n3539 0.00145131
R19719 VDD.n3896 VDD.n3797 0.00145131
R19720 VDD.n3838 VDD.n3797 0.00145131
R19721 VDD.n4154 VDD.n4055 0.00145131
R19722 VDD.n4096 VDD.n4055 0.00145131
R19723 VDD.n4412 VDD.n4313 0.00145131
R19724 VDD.n4354 VDD.n4313 0.00145131
R19725 VDD.n4670 VDD.n4571 0.00145131
R19726 VDD.n4612 VDD.n4571 0.00145131
R19727 VDD.n4928 VDD.n4829 0.00145131
R19728 VDD.n4870 VDD.n4829 0.00145131
R19729 VDD.n5186 VDD.n5087 0.00145131
R19730 VDD.n5128 VDD.n5087 0.00145131
R19731 VDD.n1770 VDD.n1769 0.00145112
R19732 VDD.n2119 VDD.n2118 0.00145112
R19733 VDD.n2349 VDD.n2348 0.00145112
R19734 VDD.n2607 VDD.n2606 0.00145112
R19735 VDD.n2865 VDD.n2864 0.00145112
R19736 VDD.n3123 VDD.n3122 0.00145112
R19737 VDD.n3381 VDD.n3380 0.00145112
R19738 VDD.n5704 VDD.n5703 0.00145112
R19739 VDD.n5450 VDD.n5449 0.00145112
R19740 VDD.n3639 VDD.n3638 0.00145112
R19741 VDD.n3897 VDD.n3896 0.00145112
R19742 VDD.n4155 VDD.n4154 0.00145112
R19743 VDD.n4413 VDD.n4412 0.00145112
R19744 VDD.n4671 VDD.n4670 0.00145112
R19745 VDD.n4929 VDD.n4928 0.00145112
R19746 VDD.n5187 VDD.n5186 0.00145112
R19747 VDD.n1756 VDD.n1755 0.00144714
R19748 VDD.n2105 VDD.n2104 0.00144714
R19749 VDD.n2335 VDD.n2334 0.00144714
R19750 VDD.n2593 VDD.n2592 0.00144714
R19751 VDD.n2851 VDD.n2850 0.00144714
R19752 VDD.n3109 VDD.n3108 0.00144714
R19753 VDD.n3367 VDD.n3366 0.00144714
R19754 VDD.n5690 VDD.n5689 0.00144714
R19755 VDD.n5436 VDD.n5435 0.00144714
R19756 VDD.n3625 VDD.n3624 0.00144714
R19757 VDD.n3883 VDD.n3882 0.00144714
R19758 VDD.n4141 VDD.n4140 0.00144714
R19759 VDD.n4399 VDD.n4398 0.00144714
R19760 VDD.n4657 VDD.n4656 0.00144714
R19761 VDD.n4915 VDD.n4914 0.00144714
R19762 VDD.n5173 VDD.n5172 0.00144714
R19763 VDD.n1755 VDD.n1754 0.00144695
R19764 VDD.n2104 VDD.n2103 0.00144695
R19765 VDD.n2334 VDD.n2333 0.00144695
R19766 VDD.n2592 VDD.n2591 0.00144695
R19767 VDD.n2850 VDD.n2849 0.00144695
R19768 VDD.n3108 VDD.n3107 0.00144695
R19769 VDD.n3366 VDD.n3365 0.00144695
R19770 VDD.n5689 VDD.n5688 0.00144695
R19771 VDD.n5435 VDD.n5434 0.00144695
R19772 VDD.n3624 VDD.n3623 0.00144695
R19773 VDD.n3882 VDD.n3881 0.00144695
R19774 VDD.n4140 VDD.n4139 0.00144695
R19775 VDD.n4398 VDD.n4397 0.00144695
R19776 VDD.n4656 VDD.n4655 0.00144695
R19777 VDD.n4914 VDD.n4913 0.00144695
R19778 VDD.n5172 VDD.n5171 0.00144695
R19779 VDD.n798 VDD.n797 0.00143548
R19780 VDD.n686 VDD.n685 0.00142105
R19781 VDD.n1036 VDD.n1035 0.00142105
R19782 VDD.n1978 VDD.n1924 0.00139286
R19783 VDD.n1719 VDD.n1668 0.00139286
R19784 VDD.n2068 VDD.n2017 0.00139286
R19785 VDD.n2298 VDD.n2247 0.00139286
R19786 VDD.n2556 VDD.n2505 0.00139286
R19787 VDD.n2814 VDD.n2763 0.00139286
R19788 VDD.n3072 VDD.n3021 0.00139286
R19789 VDD.n3330 VDD.n3279 0.00139286
R19790 VDD.n5653 VDD.n5602 0.00139286
R19791 VDD.n5399 VDD.n5348 0.00139286
R19792 VDD.n3588 VDD.n3537 0.00139286
R19793 VDD.n3846 VDD.n3795 0.00139286
R19794 VDD.n4104 VDD.n4053 0.00139286
R19795 VDD.n4362 VDD.n4311 0.00139286
R19796 VDD.n4620 VDD.n4569 0.00139286
R19797 VDD.n4878 VDD.n4827 0.00139286
R19798 VDD.n5136 VDD.n5085 0.00139286
R19799 VDD.t1041 VDD.n1941 0.00134143
R19800 VDD.n1885 VDD.n1819 0.00133663
R19801 VDD.n1821 VDD.n1819 0.00133663
R19802 VDD.n2206 VDD.n2140 0.00133663
R19803 VDD.n2142 VDD.n2140 0.00133663
R19804 VDD.n2464 VDD.n2398 0.00133663
R19805 VDD.n2400 VDD.n2398 0.00133663
R19806 VDD.n2722 VDD.n2656 0.00133663
R19807 VDD.n2658 VDD.n2656 0.00133663
R19808 VDD.n2980 VDD.n2914 0.00133663
R19809 VDD.n2916 VDD.n2914 0.00133663
R19810 VDD.n3238 VDD.n3172 0.00133663
R19811 VDD.n3174 VDD.n3172 0.00133663
R19812 VDD.n3496 VDD.n3430 0.00133663
R19813 VDD.n3432 VDD.n3430 0.00133663
R19814 VDD.n5816 VDD.n5750 0.00133663
R19815 VDD.n5752 VDD.n5750 0.00133663
R19816 VDD.n5562 VDD.n5496 0.00133663
R19817 VDD.n5498 VDD.n5496 0.00133663
R19818 VDD.n3754 VDD.n3688 0.00133663
R19819 VDD.n3690 VDD.n3688 0.00133663
R19820 VDD.n4012 VDD.n3946 0.00133663
R19821 VDD.n3948 VDD.n3946 0.00133663
R19822 VDD.n4270 VDD.n4204 0.00133663
R19823 VDD.n4206 VDD.n4204 0.00133663
R19824 VDD.n4528 VDD.n4462 0.00133663
R19825 VDD.n4464 VDD.n4462 0.00133663
R19826 VDD.n4786 VDD.n4720 0.00133663
R19827 VDD.n4722 VDD.n4720 0.00133663
R19828 VDD.n5044 VDD.n4978 0.00133663
R19829 VDD.n4980 VDD.n4978 0.00133663
R19830 VDD.n5302 VDD.n5236 0.00133663
R19831 VDD.n5238 VDD.n5236 0.00133663
R19832 VDD.n1981 VDD 0.00130357
R19833 VDD.n283 VDD 0.00128947
R19834 VDD.n1805 VDD.n1775 0.00120516
R19835 VDD.n2125 VDD.n2124 0.00120516
R19836 VDD.n2384 VDD.n2354 0.00120516
R19837 VDD.n2642 VDD.n2612 0.00120516
R19838 VDD.n2900 VDD.n2870 0.00120516
R19839 VDD.n3158 VDD.n3128 0.00120516
R19840 VDD.n3416 VDD.n3386 0.00120516
R19841 VDD.n3674 VDD.n3644 0.00120516
R19842 VDD.n3932 VDD.n3902 0.00120516
R19843 VDD.n4190 VDD.n4160 0.00120516
R19844 VDD.n4448 VDD.n4418 0.00120516
R19845 VDD.n4706 VDD.n4676 0.00120516
R19846 VDD.n4964 VDD.n4934 0.00120516
R19847 VDD.n5222 VDD.n5192 0.00120516
R19848 VDD.n855 VDD.n821 0.00116652
R19849 VDD.n1238 VDD.n1204 0.00116652
R19850 VDD.n859 VDD.n858 0.00114708
R19851 VDD.n858 VDD.n856 0.00114708
R19852 VDD.n1242 VDD.n1241 0.00114708
R19853 VDD.n1241 VDD.n1239 0.00114708
R19854 VDD.n1871 VDD.n1844 0.00114565
R19855 VDD.n1847 VDD.n1844 0.00114565
R19856 VDD.n2192 VDD.n2165 0.00114565
R19857 VDD.n2168 VDD.n2165 0.00114565
R19858 VDD.n2450 VDD.n2423 0.00114565
R19859 VDD.n2426 VDD.n2423 0.00114565
R19860 VDD.n2708 VDD.n2681 0.00114565
R19861 VDD.n2684 VDD.n2681 0.00114565
R19862 VDD.n2966 VDD.n2939 0.00114565
R19863 VDD.n2942 VDD.n2939 0.00114565
R19864 VDD.n3224 VDD.n3197 0.00114565
R19865 VDD.n3200 VDD.n3197 0.00114565
R19866 VDD.n3482 VDD.n3455 0.00114565
R19867 VDD.n3458 VDD.n3455 0.00114565
R19868 VDD.n5802 VDD.n5775 0.00114565
R19869 VDD.n5778 VDD.n5775 0.00114565
R19870 VDD.n5548 VDD.n5521 0.00114565
R19871 VDD.n5524 VDD.n5521 0.00114565
R19872 VDD.n3740 VDD.n3713 0.00114565
R19873 VDD.n3716 VDD.n3713 0.00114565
R19874 VDD.n3998 VDD.n3971 0.00114565
R19875 VDD.n3974 VDD.n3971 0.00114565
R19876 VDD.n4256 VDD.n4229 0.00114565
R19877 VDD.n4232 VDD.n4229 0.00114565
R19878 VDD.n4514 VDD.n4487 0.00114565
R19879 VDD.n4490 VDD.n4487 0.00114565
R19880 VDD.n4772 VDD.n4745 0.00114565
R19881 VDD.n4748 VDD.n4745 0.00114565
R19882 VDD.n5030 VDD.n5003 0.00114565
R19883 VDD.n5006 VDD.n5003 0.00114565
R19884 VDD.n5288 VDD.n5261 0.00114565
R19885 VDD.n5264 VDD.n5261 0.00114565
R19886 VDD.n1739 VDD.n1738 0.00113805
R19887 VDD.n2088 VDD.n2087 0.00113805
R19888 VDD.n2318 VDD.n2317 0.00113805
R19889 VDD.n2576 VDD.n2575 0.00113805
R19890 VDD.n2834 VDD.n2833 0.00113805
R19891 VDD.n3092 VDD.n3091 0.00113805
R19892 VDD.n3350 VDD.n3349 0.00113805
R19893 VDD.n5673 VDD.n5672 0.00113805
R19894 VDD.n5419 VDD.n5418 0.00113805
R19895 VDD.n3608 VDD.n3607 0.00113805
R19896 VDD.n3866 VDD.n3865 0.00113805
R19897 VDD.n4124 VDD.n4123 0.00113805
R19898 VDD.n4382 VDD.n4381 0.00113805
R19899 VDD.n4640 VDD.n4639 0.00113805
R19900 VDD.n4898 VDD.n4897 0.00113805
R19901 VDD.n5156 VDD.n5155 0.00113805
R19902 VDD.n1621 VDD.n1620 0.00111657
R19903 VDD.n1976 VDD.n1975 0.00111635
R19904 VDD.t1043 VDD.n1969 0.0010973
R19905 VDD.n1798 VDD.n1797 0.00108642
R19906 VDD.n2006 VDD.n2005 0.00108642
R19907 VDD.n2377 VDD.n2376 0.00108642
R19908 VDD.n2635 VDD.n2634 0.00108642
R19909 VDD.n2893 VDD.n2892 0.00108642
R19910 VDD.n3151 VDD.n3150 0.00108642
R19911 VDD.n3409 VDD.n3408 0.00108642
R19912 VDD.n5732 VDD.n5731 0.00108642
R19913 VDD.n5478 VDD.n5477 0.00108642
R19914 VDD.n3667 VDD.n3666 0.00108642
R19915 VDD.n3925 VDD.n3924 0.00108642
R19916 VDD.n4183 VDD.n4182 0.00108642
R19917 VDD.n4441 VDD.n4440 0.00108642
R19918 VDD.n4699 VDD.n4698 0.00108642
R19919 VDD.n4957 VDD.n4956 0.00108642
R19920 VDD.n5215 VDD.n5214 0.00108642
R19921 VDD.n860 VDD.n859 0.00107711
R19922 VDD.n1243 VDD.n1242 0.00107711
R19923 VDD.n1642 VDD.n1641 0.00107006
R19924 VDD.n1613 VDD.n1612 0.00106596
R19925 VDD.n1752 VDD.n1720 0.00105202
R19926 VDD.n2101 VDD.n2069 0.00105202
R19927 VDD.n2331 VDD.n2299 0.00105202
R19928 VDD.n2589 VDD.n2557 0.00105202
R19929 VDD.n2847 VDD.n2815 0.00105202
R19930 VDD.n3105 VDD.n3073 0.00105202
R19931 VDD.n3363 VDD.n3331 0.00105202
R19932 VDD.n5686 VDD.n5654 0.00105202
R19933 VDD.n5432 VDD.n5400 0.00105202
R19934 VDD.n3621 VDD.n3589 0.00105202
R19935 VDD.n3879 VDD.n3847 0.00105202
R19936 VDD.n4137 VDD.n4105 0.00105202
R19937 VDD.n4395 VDD.n4363 0.00105202
R19938 VDD.n4653 VDD.n4621 0.00105202
R19939 VDD.n4911 VDD.n4879 0.00105202
R19940 VDD.n5169 VDD.n5137 0.00105202
R19941 VDD.n1431 VDD.n1430 0.00100344
R19942 VDD.n1455 VDD.n1454 0.00100344
R19943 VDD.n1374 VDD.n1373 0.00100342
R19944 VDD.n1711 VDD.n1710 0.00100293
R19945 VDD.n2060 VDD.n2059 0.00100293
R19946 VDD.n2290 VDD.n2289 0.00100293
R19947 VDD.n2548 VDD.n2547 0.00100293
R19948 VDD.n2806 VDD.n2805 0.00100293
R19949 VDD.n3064 VDD.n3063 0.00100293
R19950 VDD.n3322 VDD.n3321 0.00100293
R19951 VDD.n5645 VDD.n5644 0.00100293
R19952 VDD.n5391 VDD.n5390 0.00100293
R19953 VDD.n3580 VDD.n3579 0.00100293
R19954 VDD.n3838 VDD.n3837 0.00100293
R19955 VDD.n4096 VDD.n4095 0.00100293
R19956 VDD.n4354 VDD.n4353 0.00100293
R19957 VDD.n4612 VDD.n4611 0.00100293
R19958 VDD.n4870 VDD.n4869 0.00100293
R19959 VDD.n5128 VDD.n5127 0.00100293
R19960 VDD.n464 VDD.n463 0.00100258
R19961 VDD.n61 VDD.n60 0.00100258
R19962 VDD.n1837 VDD.n1826 0.00100132
R19963 VDD.n2158 VDD.n2147 0.00100132
R19964 VDD.n2416 VDD.n2405 0.00100132
R19965 VDD.n2674 VDD.n2663 0.00100132
R19966 VDD.n2932 VDD.n2921 0.00100132
R19967 VDD.n3190 VDD.n3179 0.00100132
R19968 VDD.n3448 VDD.n3437 0.00100132
R19969 VDD.n5768 VDD.n5757 0.00100132
R19970 VDD.n5514 VDD.n5503 0.00100132
R19971 VDD.n3706 VDD.n3695 0.00100132
R19972 VDD.n3964 VDD.n3953 0.00100132
R19973 VDD.n4222 VDD.n4211 0.00100132
R19974 VDD.n4480 VDD.n4469 0.00100132
R19975 VDD.n4738 VDD.n4727 0.00100132
R19976 VDD.n4996 VDD.n4985 0.00100132
R19977 VDD.n5254 VDD.n5243 0.00100132
R19978 VDD.n587 VDD.n586 0.00100097
R19979 VDD.n937 VDD.n936 0.00100097
R19980 VDD.n186 VDD.n185 0.00100097
R19981 VDD.n1547 VDD.n1541 0.00100097
R19982 VDD.n1620 VDD.n1614 0.00100057
R19983 VDD.n1798 VDD.n1777 0.00100033
R19984 VDD.n2006 VDD.n1985 0.00100033
R19985 VDD.n2377 VDD.n2356 0.00100033
R19986 VDD.n2635 VDD.n2614 0.00100033
R19987 VDD.n2893 VDD.n2872 0.00100033
R19988 VDD.n3151 VDD.n3130 0.00100033
R19989 VDD.n3409 VDD.n3388 0.00100033
R19990 VDD.n5732 VDD.n5711 0.00100033
R19991 VDD.n5478 VDD.n5457 0.00100033
R19992 VDD.n3667 VDD.n3646 0.00100033
R19993 VDD.n3925 VDD.n3904 0.00100033
R19994 VDD.n4183 VDD.n4162 0.00100033
R19995 VDD.n4441 VDD.n4420 0.00100033
R19996 VDD.n4699 VDD.n4678 0.00100033
R19997 VDD.n4957 VDD.n4936 0.00100033
R19998 VDD.n5215 VDD.n5194 0.00100033
R19999 VDD.n1882 VDD.n1821 0.00100021
R20000 VDD.n2203 VDD.n2142 0.00100021
R20001 VDD.n2461 VDD.n2400 0.00100021
R20002 VDD.n2719 VDD.n2658 0.00100021
R20003 VDD.n2977 VDD.n2916 0.00100021
R20004 VDD.n3235 VDD.n3174 0.00100021
R20005 VDD.n3493 VDD.n3432 0.00100021
R20006 VDD.n5813 VDD.n5752 0.00100021
R20007 VDD.n5559 VDD.n5498 0.00100021
R20008 VDD.n3751 VDD.n3690 0.00100021
R20009 VDD.n4009 VDD.n3948 0.00100021
R20010 VDD.n4267 VDD.n4206 0.00100021
R20011 VDD.n4525 VDD.n4464 0.00100021
R20012 VDD.n4783 VDD.n4722 0.00100021
R20013 VDD.n5041 VDD.n4980 0.00100021
R20014 VDD.n5299 VDD.n5238 0.00100021
R20015 VDD.n860 VDD.n855 0.00100013
R20016 VDD.n1243 VDD.n1238 0.00100013
R20017 VDD.n1757 VDD.n1711 0.0010001
R20018 VDD.n2106 VDD.n2060 0.0010001
R20019 VDD.n2336 VDD.n2290 0.0010001
R20020 VDD.n2594 VDD.n2548 0.0010001
R20021 VDD.n2852 VDD.n2806 0.0010001
R20022 VDD.n3110 VDD.n3064 0.0010001
R20023 VDD.n3368 VDD.n3322 0.0010001
R20024 VDD.n5691 VDD.n5645 0.0010001
R20025 VDD.n5437 VDD.n5391 0.0010001
R20026 VDD.n3626 VDD.n3580 0.0010001
R20027 VDD.n3884 VDD.n3838 0.0010001
R20028 VDD.n4142 VDD.n4096 0.0010001
R20029 VDD.n4400 VDD.n4354 0.0010001
R20030 VDD.n4658 VDD.n4612 0.0010001
R20031 VDD.n4916 VDD.n4870 0.0010001
R20032 VDD.n5174 VDD.n5128 0.0010001
R20033 VDD.n1641 VDD.n1640 0.00100008
R20034 VDD.n1952 VDD.n1944 0.00100003
R20035 VDD.n1934 VDD.n1927 0.00100003
R20036 VDD.n1920 VDD.n1808 0.00100002
R20037 VDD.n2241 VDD.n2129 0.00100002
R20038 VDD.n2499 VDD.n2387 0.00100002
R20039 VDD.n2757 VDD.n2645 0.00100002
R20040 VDD.n3015 VDD.n2903 0.00100002
R20041 VDD.n3273 VDD.n3161 0.00100002
R20042 VDD.n3531 VDD.n3419 0.00100002
R20043 VDD.n3789 VDD.n3677 0.00100002
R20044 VDD.n4047 VDD.n3935 0.00100002
R20045 VDD.n4305 VDD.n4193 0.00100002
R20046 VDD.n4563 VDD.n4451 0.00100002
R20047 VDD.n4821 VDD.n4709 0.00100002
R20048 VDD.n5079 VDD.n4967 0.00100002
R20049 VDD.n5337 VDD.n5225 0.00100002
R20050 VDD.n1317 VDD.n1315 0.001
R20051 VDD.n1975 VDD.n1927 0.001
R20052 VDD.n1979 VDD.n1923 0.001
R20053 VDD.n858 VDD.n857 0.001
R20054 VDD.n1241 VDD.n1240 0.001
R20055 VDD.n390 VDD.n389 0.000894737
R20056 VDD.n1640 VDD.n1638 0.000834423
R20057 VDD.n1460 VDD.n1459 0.000765957
R20058 VDD.n688 VDD 0.000763158
R20059 VDD.n1038 VDD 0.000763158
R20060 VDD.n793 VDD.n515 0.000631579
R20061 VDD.n1143 VDD.n865 0.000631579
R20062 VDD.n1621 VDD.n1615 0.000625544
R20063 VDD.n1619 VDD.n1615 0.000625542
R20064 VDD.n1977 VDD.n1976 0.00061635
R20065 VDD.n1978 VDD.n1977 0.000616347
R20066 VDD.n1736 VDD.n1729 0.000594432
R20067 VDD.n2085 VDD.n2078 0.000594432
R20068 VDD.n2315 VDD.n2308 0.000594432
R20069 VDD.n2573 VDD.n2566 0.000594432
R20070 VDD.n2831 VDD.n2824 0.000594432
R20071 VDD.n3089 VDD.n3082 0.000594432
R20072 VDD.n3347 VDD.n3340 0.000594432
R20073 VDD.n5670 VDD.n5663 0.000594432
R20074 VDD.n5416 VDD.n5409 0.000594432
R20075 VDD.n3605 VDD.n3598 0.000594432
R20076 VDD.n3863 VDD.n3856 0.000594432
R20077 VDD.n4121 VDD.n4114 0.000594432
R20078 VDD.n4379 VDD.n4372 0.000594432
R20079 VDD.n4637 VDD.n4630 0.000594432
R20080 VDD.n4895 VDD.n4888 0.000594432
R20081 VDD.n5153 VDD.n5146 0.000594432
R20082 VDD.n1773 VDD.n1772 0.000558569
R20083 VDD.n2122 VDD.n2121 0.000558569
R20084 VDD.n2352 VDD.n2351 0.000558569
R20085 VDD.n2610 VDD.n2609 0.000558569
R20086 VDD.n2868 VDD.n2867 0.000558569
R20087 VDD.n3126 VDD.n3125 0.000558569
R20088 VDD.n3384 VDD.n3383 0.000558569
R20089 VDD.n5707 VDD.n5706 0.000558569
R20090 VDD.n5453 VDD.n5452 0.000558569
R20091 VDD.n3642 VDD.n3641 0.000558569
R20092 VDD.n3900 VDD.n3899 0.000558569
R20093 VDD.n4158 VDD.n4157 0.000558569
R20094 VDD.n4416 VDD.n4415 0.000558569
R20095 VDD.n4674 VDD.n4673 0.000558569
R20096 VDD.n4932 VDD.n4931 0.000558569
R20097 VDD.n5190 VDD.n5189 0.000558569
R20098 VDD.n1740 VDD.n1739 0.000555817
R20099 VDD.n2089 VDD.n2088 0.000555817
R20100 VDD.n2319 VDD.n2318 0.000555817
R20101 VDD.n2577 VDD.n2576 0.000555817
R20102 VDD.n2835 VDD.n2834 0.000555817
R20103 VDD.n3093 VDD.n3092 0.000555817
R20104 VDD.n3351 VDD.n3350 0.000555817
R20105 VDD.n5674 VDD.n5673 0.000555817
R20106 VDD.n5420 VDD.n5419 0.000555817
R20107 VDD.n3609 VDD.n3608 0.000555817
R20108 VDD.n3867 VDD.n3866 0.000555817
R20109 VDD.n4125 VDD.n4124 0.000555817
R20110 VDD.n4383 VDD.n4382 0.000555817
R20111 VDD.n4641 VDD.n4640 0.000555817
R20112 VDD.n4899 VDD.n4898 0.000555817
R20113 VDD.n5157 VDD.n5156 0.000555817
R20114 VDD.n1768 VDD.n1668 0.000534058
R20115 VDD.n2117 VDD.n2017 0.000534058
R20116 VDD.n2347 VDD.n2247 0.000534058
R20117 VDD.n2605 VDD.n2505 0.000534058
R20118 VDD.n2863 VDD.n2763 0.000534058
R20119 VDD.n3121 VDD.n3021 0.000534058
R20120 VDD.n3379 VDD.n3279 0.000534058
R20121 VDD.n5702 VDD.n5602 0.000534058
R20122 VDD.n5448 VDD.n5348 0.000534058
R20123 VDD.n3637 VDD.n3537 0.000534058
R20124 VDD.n3895 VDD.n3795 0.000534058
R20125 VDD.n4153 VDD.n4053 0.000534058
R20126 VDD.n4411 VDD.n4311 0.000534058
R20127 VDD.n4669 VDD.n4569 0.000534058
R20128 VDD.n4927 VDD.n4827 0.000534058
R20129 VDD.n5185 VDD.n5085 0.000534058
R20130 VDD.n1886 VDD.n1885 0.000523376
R20131 VDD.n2207 VDD.n2206 0.000523376
R20132 VDD.n2465 VDD.n2464 0.000523376
R20133 VDD.n2723 VDD.n2722 0.000523376
R20134 VDD.n2981 VDD.n2980 0.000523376
R20135 VDD.n3239 VDD.n3238 0.000523376
R20136 VDD.n3497 VDD.n3496 0.000523376
R20137 VDD.n5817 VDD.n5816 0.000523376
R20138 VDD.n5563 VDD.n5562 0.000523376
R20139 VDD.n3755 VDD.n3754 0.000523376
R20140 VDD.n4013 VDD.n4012 0.000523376
R20141 VDD.n4271 VDD.n4270 0.000523376
R20142 VDD.n4529 VDD.n4528 0.000523376
R20143 VDD.n4787 VDD.n4786 0.000523376
R20144 VDD.n5045 VDD.n5044 0.000523376
R20145 VDD.n5303 VDD.n5302 0.000523376
R20146 VDD.n1704 VDD.n1703 0.000516232
R20147 VDD.n1691 VDD.n1685 0.000516232
R20148 VDD.n2053 VDD.n2052 0.000516232
R20149 VDD.n2040 VDD.n2034 0.000516232
R20150 VDD.n2283 VDD.n2282 0.000516232
R20151 VDD.n2270 VDD.n2264 0.000516232
R20152 VDD.n2541 VDD.n2540 0.000516232
R20153 VDD.n2528 VDD.n2522 0.000516232
R20154 VDD.n2799 VDD.n2798 0.000516232
R20155 VDD.n2786 VDD.n2780 0.000516232
R20156 VDD.n3057 VDD.n3056 0.000516232
R20157 VDD.n3044 VDD.n3038 0.000516232
R20158 VDD.n3315 VDD.n3314 0.000516232
R20159 VDD.n3302 VDD.n3296 0.000516232
R20160 VDD.n5638 VDD.n5637 0.000516232
R20161 VDD.n5625 VDD.n5619 0.000516232
R20162 VDD.n5384 VDD.n5383 0.000516232
R20163 VDD.n5371 VDD.n5365 0.000516232
R20164 VDD.n3573 VDD.n3572 0.000516232
R20165 VDD.n3560 VDD.n3554 0.000516232
R20166 VDD.n3831 VDD.n3830 0.000516232
R20167 VDD.n3818 VDD.n3812 0.000516232
R20168 VDD.n4089 VDD.n4088 0.000516232
R20169 VDD.n4076 VDD.n4070 0.000516232
R20170 VDD.n4347 VDD.n4346 0.000516232
R20171 VDD.n4334 VDD.n4328 0.000516232
R20172 VDD.n4605 VDD.n4604 0.000516232
R20173 VDD.n4592 VDD.n4586 0.000516232
R20174 VDD.n4863 VDD.n4862 0.000516232
R20175 VDD.n4850 VDD.n4844 0.000516232
R20176 VDD.n5121 VDD.n5120 0.000516232
R20177 VDD.n5108 VDD.n5102 0.000516232
R20178 VDD.n1735 VDD.n1734 0.000515622
R20179 VDD.n2084 VDD.n2083 0.000515622
R20180 VDD.n2314 VDD.n2313 0.000515622
R20181 VDD.n2572 VDD.n2571 0.000515622
R20182 VDD.n2830 VDD.n2829 0.000515622
R20183 VDD.n3088 VDD.n3087 0.000515622
R20184 VDD.n3346 VDD.n3345 0.000515622
R20185 VDD.n5669 VDD.n5668 0.000515622
R20186 VDD.n5415 VDD.n5414 0.000515622
R20187 VDD.n3604 VDD.n3603 0.000515622
R20188 VDD.n3862 VDD.n3861 0.000515622
R20189 VDD.n4120 VDD.n4119 0.000515622
R20190 VDD.n4378 VDD.n4377 0.000515622
R20191 VDD.n4636 VDD.n4635 0.000515622
R20192 VDD.n4894 VDD.n4893 0.000515622
R20193 VDD.n5152 VDD.n5151 0.000515622
R20194 VDD.n1876 VDD.n1875 0.000514451
R20195 VDD.n2197 VDD.n2196 0.000514451
R20196 VDD.n2455 VDD.n2454 0.000514451
R20197 VDD.n2713 VDD.n2712 0.000514451
R20198 VDD.n2971 VDD.n2970 0.000514451
R20199 VDD.n3229 VDD.n3228 0.000514451
R20200 VDD.n3487 VDD.n3486 0.000514451
R20201 VDD.n5807 VDD.n5806 0.000514451
R20202 VDD.n5553 VDD.n5552 0.000514451
R20203 VDD.n3745 VDD.n3744 0.000514451
R20204 VDD.n4003 VDD.n4002 0.000514451
R20205 VDD.n4261 VDD.n4260 0.000514451
R20206 VDD.n4519 VDD.n4518 0.000514451
R20207 VDD.n4777 VDD.n4776 0.000514451
R20208 VDD.n5035 VDD.n5034 0.000514451
R20209 VDD.n5293 VDD.n5292 0.000514451
R20210 VDD.n669 VDD.n521 0.000506553
R20211 VDD.n668 VDD.n518 0.000506553
R20212 VDD.n667 VDD.n666 0.000506553
R20213 VDD.n586 VDD.n585 0.000506553
R20214 VDD.n584 VDD.n583 0.000506553
R20215 VDD.n687 VDD.n670 0.000506553
R20216 VDD.n1019 VDD.n871 0.000506553
R20217 VDD.n1018 VDD.n868 0.000506553
R20218 VDD.n1017 VDD.n1016 0.000506553
R20219 VDD.n936 VDD.n935 0.000506553
R20220 VDD.n934 VDD.n933 0.000506553
R20221 VDD.n1037 VDD.n1020 0.000506553
R20222 VDD.n264 VDD.n120 0.000506553
R20223 VDD.n263 VDD.n117 0.000506553
R20224 VDD.n262 VDD.n261 0.000506553
R20225 VDD.n185 VDD.n184 0.000506553
R20226 VDD.n183 VDD.n182 0.000506553
R20227 VDD.n282 VDD.n265 0.000506553
R20228 VDD.n1458 VDD.n1457 0.000506553
R20229 VDD.n1508 VDD.n1507 0.000506553
R20230 VDD.n1456 VDD.n1455 0.000506553
R20231 VDD.n1430 VDD.n1429 0.000506553
R20232 VDD.n1398 VDD.n1397 0.000506553
R20233 VDD.n1373 VDD.n1372 0.000506553
R20234 VDD.n1371 VDD.n1370 0.000506553
R20235 VDD.n1428 VDD.n1427 0.000506553
R20236 VDD.n1726 VDD.n1725 0.000505865
R20237 VDD.n2075 VDD.n2074 0.000505865
R20238 VDD.n2305 VDD.n2304 0.000505865
R20239 VDD.n2563 VDD.n2562 0.000505865
R20240 VDD.n2821 VDD.n2820 0.000505865
R20241 VDD.n3079 VDD.n3078 0.000505865
R20242 VDD.n3337 VDD.n3336 0.000505865
R20243 VDD.n5660 VDD.n5659 0.000505865
R20244 VDD.n5406 VDD.n5405 0.000505865
R20245 VDD.n3595 VDD.n3594 0.000505865
R20246 VDD.n3853 VDD.n3852 0.000505865
R20247 VDD.n4111 VDD.n4110 0.000505865
R20248 VDD.n4369 VDD.n4368 0.000505865
R20249 VDD.n4627 VDD.n4626 0.000505865
R20250 VDD.n4885 VDD.n4884 0.000505865
R20251 VDD.n5143 VDD.n5142 0.000505865
R20252 VDD.n1839 VDD.n1838 0.000504381
R20253 VDD.n2160 VDD.n2159 0.000504381
R20254 VDD.n2418 VDD.n2417 0.000504381
R20255 VDD.n2676 VDD.n2675 0.000504381
R20256 VDD.n2934 VDD.n2933 0.000504381
R20257 VDD.n3192 VDD.n3191 0.000504381
R20258 VDD.n3450 VDD.n3449 0.000504381
R20259 VDD.n5770 VDD.n5769 0.000504381
R20260 VDD.n5516 VDD.n5515 0.000504381
R20261 VDD.n3708 VDD.n3707 0.000504381
R20262 VDD.n3966 VDD.n3965 0.000504381
R20263 VDD.n4224 VDD.n4223 0.000504381
R20264 VDD.n4482 VDD.n4481 0.000504381
R20265 VDD.n4740 VDD.n4739 0.000504381
R20266 VDD.n4998 VDD.n4997 0.000504381
R20267 VDD.n5256 VDD.n5255 0.000504381
R20268 VDD.n1719 VDD.n1671 0.000503792
R20269 VDD.n2068 VDD.n2020 0.000503792
R20270 VDD.n2298 VDD.n2250 0.000503792
R20271 VDD.n2556 VDD.n2508 0.000503792
R20272 VDD.n2814 VDD.n2766 0.000503792
R20273 VDD.n3072 VDD.n3024 0.000503792
R20274 VDD.n3330 VDD.n3282 0.000503792
R20275 VDD.n5653 VDD.n5605 0.000503792
R20276 VDD.n5399 VDD.n5351 0.000503792
R20277 VDD.n3588 VDD.n3540 0.000503792
R20278 VDD.n3846 VDD.n3798 0.000503792
R20279 VDD.n4104 VDD.n4056 0.000503792
R20280 VDD.n4362 VDD.n4314 0.000503792
R20281 VDD.n4620 VDD.n4572 0.000503792
R20282 VDD.n4878 VDD.n4830 0.000503792
R20283 VDD.n5136 VDD.n5088 0.000503792
R20284 VDD.n1427 VDD.n1426 0.000503441
R20285 VDD.n1399 VDD.n1398 0.000503441
R20286 VDD.n1370 VDD.n1369 0.000503441
R20287 VDD.n1459 VDD.n1458 0.000503441
R20288 VDD.n1509 VDD.n1508 0.000503441
R20289 VDD.n1345 VDD.n1344 0.000501258
R20290 VDD.n1319 VDD.n1318 0.000501258
R20291 VDD.n1401 VDD.n1400 0.000501258
R20292 VDD.n1361 VDD.n1360 0.000501258
R20293 VDD.n1289 VDD.n1288 0.000501258
R20294 VDD.n1506 VDD.n1505 0.000501258
R20295 VDD.n1818 VDD.n1817 0.000501164
R20296 VDD.n2139 VDD.n2138 0.000501164
R20297 VDD.n2397 VDD.n2396 0.000501164
R20298 VDD.n2655 VDD.n2654 0.000501164
R20299 VDD.n2913 VDD.n2912 0.000501164
R20300 VDD.n3171 VDD.n3170 0.000501164
R20301 VDD.n3429 VDD.n3428 0.000501164
R20302 VDD.n5749 VDD.n5748 0.000501164
R20303 VDD.n5495 VDD.n5494 0.000501164
R20304 VDD.n3687 VDD.n3686 0.000501164
R20305 VDD.n3945 VDD.n3944 0.000501164
R20306 VDD.n4203 VDD.n4202 0.000501164
R20307 VDD.n4461 VDD.n4460 0.000501164
R20308 VDD.n4719 VDD.n4718 0.000501164
R20309 VDD.n4977 VDD.n4976 0.000501164
R20310 VDD.n5235 VDD.n5234 0.000501164
R20311 VDD.n736 VDD.n521 0.00050097
R20312 VDD.n781 VDD.n518 0.00050097
R20313 VDD.n666 VDD.n665 0.00050097
R20314 VDD.n583 VDD.n582 0.00050097
R20315 VDD.n1086 VDD.n871 0.00050097
R20316 VDD.n1131 VDD.n868 0.00050097
R20317 VDD.n1016 VDD.n1015 0.00050097
R20318 VDD.n933 VDD.n932 0.00050097
R20319 VDD.n331 VDD.n120 0.00050097
R20320 VDD.n376 VDD.n117 0.00050097
R20321 VDD.n261 VDD.n260 0.00050097
R20322 VDD.n182 VDD.n181 0.00050097
R20323 VDD.n687 VDD.n686 0.00050097
R20324 VDD.n1037 VDD.n1036 0.00050097
R20325 VDD.n282 VDD.n281 0.00050097
R20326 VDD.n2193 VDD.n2192 0.000500414
R20327 VDD.n2451 VDD.n2450 0.000500414
R20328 VDD.n2709 VDD.n2708 0.000500414
R20329 VDD.n2967 VDD.n2966 0.000500414
R20330 VDD.n3225 VDD.n3224 0.000500414
R20331 VDD.n3483 VDD.n3482 0.000500414
R20332 VDD.n5803 VDD.n5802 0.000500414
R20333 VDD.n5549 VDD.n5548 0.000500414
R20334 VDD.n3741 VDD.n3740 0.000500414
R20335 VDD.n3999 VDD.n3998 0.000500414
R20336 VDD.n4257 VDD.n4256 0.000500414
R20337 VDD.n4515 VDD.n4514 0.000500414
R20338 VDD.n4773 VDD.n4772 0.000500414
R20339 VDD.n5031 VDD.n5030 0.000500414
R20340 VDD.n5289 VDD.n5288 0.000500414
R20341 VDD.n1872 VDD.n1871 0.000500414
R20342 VDD.n863 VDD.n862 0.000500259
R20343 VDD.n1920 VDD.n1919 0.000500184
R20344 VDD.n2241 VDD.n2240 0.000500184
R20345 VDD.n2499 VDD.n2498 0.000500184
R20346 VDD.n2757 VDD.n2756 0.000500184
R20347 VDD.n3015 VDD.n3014 0.000500184
R20348 VDD.n3273 VDD.n3272 0.000500184
R20349 VDD.n3531 VDD.n3530 0.000500184
R20350 VDD.n3789 VDD.n3788 0.000500184
R20351 VDD.n4047 VDD.n4046 0.000500184
R20352 VDD.n4305 VDD.n4304 0.000500184
R20353 VDD.n4563 VDD.n4562 0.000500184
R20354 VDD.n4821 VDD.n4820 0.000500184
R20355 VDD.n5079 VDD.n5078 0.000500184
R20356 VDD.n5337 VDD.n5336 0.000500184
R20357 VDD.n1775 VDD.n1774 0.000500121
R20358 VDD.n2124 VDD.n2123 0.000500121
R20359 VDD.n2354 VDD.n2353 0.000500121
R20360 VDD.n2612 VDD.n2611 0.000500121
R20361 VDD.n2870 VDD.n2869 0.000500121
R20362 VDD.n3128 VDD.n3127 0.000500121
R20363 VDD.n3386 VDD.n3385 0.000500121
R20364 VDD.n3644 VDD.n3643 0.000500121
R20365 VDD.n3902 VDD.n3901 0.000500121
R20366 VDD.n4160 VDD.n4159 0.000500121
R20367 VDD.n4418 VDD.n4417 0.000500121
R20368 VDD.n4676 VDD.n4675 0.000500121
R20369 VDD.n4934 VDD.n4933 0.000500121
R20370 VDD.n5192 VDD.n5191 0.000500121
R20371 VDD.n2162 VDD.n1983 0.000500117
R20372 VDD.n2420 VDD.n2243 0.000500117
R20373 VDD.n2678 VDD.n2501 0.000500117
R20374 VDD.n2936 VDD.n2759 0.000500117
R20375 VDD.n3194 VDD.n3017 0.000500117
R20376 VDD.n3452 VDD.n3275 0.000500117
R20377 VDD.n5772 VDD.n5709 0.000500117
R20378 VDD.n5518 VDD.n5455 0.000500117
R20379 VDD.n3710 VDD.n3533 0.000500117
R20380 VDD.n3968 VDD.n3791 0.000500117
R20381 VDD.n4226 VDD.n4049 0.000500117
R20382 VDD.n4484 VDD.n4307 0.000500117
R20383 VDD.n4742 VDD.n4565 0.000500117
R20384 VDD.n5000 VDD.n4823 0.000500117
R20385 VDD.n5258 VDD.n5081 0.000500117
R20386 VDD.n1841 VDD.n1664 0.000500117
R20387 VDD.n1602 VDD.n1246 0.000500071
R20388 VDD.n1601 VDD.n1540 0.000500071
R20389 OUT3.n142 OUT3.n140 145.809
R20390 OUT3.n91 OUT3.n89 145.809
R20391 OUT3.n53 OUT3.n51 145.809
R20392 OUT3.n7 OUT3.n5 145.809
R20393 OUT3.n91 OUT3.n90 107.409
R20394 OUT3.n93 OUT3.n92 107.409
R20395 OUT3.n95 OUT3.n94 107.409
R20396 OUT3.n97 OUT3.n96 107.409
R20397 OUT3.n99 OUT3.n98 107.409
R20398 OUT3.n101 OUT3.n100 107.409
R20399 OUT3.n53 OUT3.n52 107.409
R20400 OUT3.n55 OUT3.n54 107.409
R20401 OUT3.n57 OUT3.n56 107.409
R20402 OUT3.n59 OUT3.n58 107.409
R20403 OUT3.n61 OUT3.n60 107.409
R20404 OUT3.n63 OUT3.n62 107.409
R20405 OUT3.n7 OUT3.n6 107.409
R20406 OUT3.n9 OUT3.n8 107.409
R20407 OUT3.n11 OUT3.n10 107.409
R20408 OUT3.n13 OUT3.n12 107.409
R20409 OUT3.n15 OUT3.n14 107.409
R20410 OUT3.n17 OUT3.n16 107.409
R20411 OUT3.n142 OUT3.n141 107.407
R20412 OUT3.n144 OUT3.n143 107.407
R20413 OUT3.n146 OUT3.n145 107.407
R20414 OUT3.n148 OUT3.n147 107.407
R20415 OUT3.n150 OUT3.n149 107.407
R20416 OUT3.n152 OUT3.n151 107.407
R20417 OUT3.n160 OUT3.n158 87.1779
R20418 OUT3.n114 OUT3.n112 87.1779
R20419 OUT3.n72 OUT3.n70 87.1779
R20420 OUT3.n26 OUT3.n24 87.1779
R20421 OUT3.n160 OUT3.n159 52.82
R20422 OUT3.n162 OUT3.n161 52.82
R20423 OUT3.n164 OUT3.n163 52.82
R20424 OUT3.n166 OUT3.n165 52.82
R20425 OUT3.n168 OUT3.n167 52.82
R20426 OUT3.n170 OUT3.n169 52.82
R20427 OUT3.n114 OUT3.n113 52.82
R20428 OUT3.n116 OUT3.n115 52.82
R20429 OUT3.n118 OUT3.n117 52.82
R20430 OUT3.n120 OUT3.n119 52.82
R20431 OUT3.n122 OUT3.n121 52.82
R20432 OUT3.n124 OUT3.n123 52.82
R20433 OUT3.n72 OUT3.n71 52.82
R20434 OUT3.n74 OUT3.n73 52.82
R20435 OUT3.n76 OUT3.n75 52.82
R20436 OUT3.n78 OUT3.n77 52.82
R20437 OUT3.n80 OUT3.n79 52.82
R20438 OUT3.n82 OUT3.n81 52.82
R20439 OUT3.n26 OUT3.n25 52.82
R20440 OUT3.n28 OUT3.n27 52.82
R20441 OUT3.n30 OUT3.n29 52.82
R20442 OUT3.n32 OUT3.n31 52.82
R20443 OUT3.n34 OUT3.n33 52.82
R20444 OUT3.n36 OUT3.n35 52.82
R20445 OUT3.n144 OUT3.n142 38.4005
R20446 OUT3.n146 OUT3.n144 38.4005
R20447 OUT3.n148 OUT3.n146 38.4005
R20448 OUT3.n150 OUT3.n148 38.4005
R20449 OUT3.n152 OUT3.n150 38.4005
R20450 OUT3.n153 OUT3.n152 38.4005
R20451 OUT3.n93 OUT3.n91 38.4005
R20452 OUT3.n95 OUT3.n93 38.4005
R20453 OUT3.n97 OUT3.n95 38.4005
R20454 OUT3.n99 OUT3.n97 38.4005
R20455 OUT3.n101 OUT3.n99 38.4005
R20456 OUT3.n102 OUT3.n101 38.4005
R20457 OUT3.n55 OUT3.n53 38.4005
R20458 OUT3.n57 OUT3.n55 38.4005
R20459 OUT3.n59 OUT3.n57 38.4005
R20460 OUT3.n61 OUT3.n59 38.4005
R20461 OUT3.n63 OUT3.n61 38.4005
R20462 OUT3.n64 OUT3.n63 38.4005
R20463 OUT3.n9 OUT3.n7 38.4005
R20464 OUT3.n11 OUT3.n9 38.4005
R20465 OUT3.n13 OUT3.n11 38.4005
R20466 OUT3.n15 OUT3.n13 38.4005
R20467 OUT3.n17 OUT3.n15 38.4005
R20468 OUT3.n18 OUT3.n17 38.4005
R20469 OUT3.n162 OUT3.n160 34.3584
R20470 OUT3.n164 OUT3.n162 34.3584
R20471 OUT3.n166 OUT3.n164 34.3584
R20472 OUT3.n168 OUT3.n166 34.3584
R20473 OUT3.n170 OUT3.n168 34.3584
R20474 OUT3.n174 OUT3.n170 34.3584
R20475 OUT3.n116 OUT3.n114 34.3584
R20476 OUT3.n118 OUT3.n116 34.3584
R20477 OUT3.n120 OUT3.n118 34.3584
R20478 OUT3.n122 OUT3.n120 34.3584
R20479 OUT3.n124 OUT3.n122 34.3584
R20480 OUT3.n129 OUT3.n124 34.3584
R20481 OUT3.n74 OUT3.n72 34.3584
R20482 OUT3.n76 OUT3.n74 34.3584
R20483 OUT3.n78 OUT3.n76 34.3584
R20484 OUT3.n80 OUT3.n78 34.3584
R20485 OUT3.n82 OUT3.n80 34.3584
R20486 OUT3.n83 OUT3.n82 34.3584
R20487 OUT3.n28 OUT3.n26 34.3584
R20488 OUT3.n30 OUT3.n28 34.3584
R20489 OUT3.n32 OUT3.n30 34.3584
R20490 OUT3.n34 OUT3.n32 34.3584
R20491 OUT3.n36 OUT3.n34 34.3584
R20492 OUT3.n40 OUT3.n36 34.3584
R20493 OUT3.n135 OUT3.t11 26.5955
R20494 OUT3.n135 OUT3.t37 26.5955
R20495 OUT3.n140 OUT3.t21 26.5955
R20496 OUT3.n140 OUT3.t60 26.5955
R20497 OUT3.n141 OUT3.t35 26.5955
R20498 OUT3.n141 OUT3.t8 26.5955
R20499 OUT3.n143 OUT3.t6 26.5955
R20500 OUT3.n143 OUT3.t19 26.5955
R20501 OUT3.n145 OUT3.t27 26.5955
R20502 OUT3.n145 OUT3.t43 26.5955
R20503 OUT3.n147 OUT3.t41 26.5955
R20504 OUT3.n147 OUT3.t63 26.5955
R20505 OUT3.n149 OUT3.t61 26.5955
R20506 OUT3.n149 OUT3.t25 26.5955
R20507 OUT3.n151 OUT3.t52 26.5955
R20508 OUT3.n151 OUT3.t13 26.5955
R20509 OUT3.n89 OUT3.t22 26.5955
R20510 OUT3.n89 OUT3.t48 26.5955
R20511 OUT3.n90 OUT3.t46 26.5955
R20512 OUT3.n90 OUT3.t9 26.5955
R20513 OUT3.n92 OUT3.t0 26.5955
R20514 OUT3.n92 OUT3.t30 26.5955
R20515 OUT3.n94 OUT3.t1 26.5955
R20516 OUT3.n94 OUT3.t17 26.5955
R20517 OUT3.n96 OUT3.t15 26.5955
R20518 OUT3.n96 OUT3.t33 26.5955
R20519 OUT3.n98 OUT3.t40 26.5955
R20520 OUT3.n98 OUT3.t54 26.5955
R20521 OUT3.n100 OUT3.t59 26.5955
R20522 OUT3.n100 OUT3.t24 26.5955
R20523 OUT3.n51 OUT3.t4 26.5955
R20524 OUT3.n51 OUT3.t49 26.5955
R20525 OUT3.n52 OUT3.t20 26.5955
R20526 OUT3.n52 OUT3.t36 26.5955
R20527 OUT3.n54 OUT3.t44 26.5955
R20528 OUT3.n54 OUT3.t7 26.5955
R20529 OUT3.n56 OUT3.t56 26.5955
R20530 OUT3.n56 OUT3.t18 26.5955
R20531 OUT3.n58 OUT3.t26 26.5955
R20532 OUT3.n58 OUT3.t42 26.5955
R20533 OUT3.n60 OUT3.t50 26.5955
R20534 OUT3.n60 OUT3.t62 26.5955
R20535 OUT3.n62 OUT3.t29 26.5955
R20536 OUT3.n62 OUT3.t5 26.5955
R20537 OUT3.n1 OUT3.t58 26.5955
R20538 OUT3.n1 OUT3.t3 26.5955
R20539 OUT3.n5 OUT3.t10 26.5955
R20540 OUT3.n5 OUT3.t23 26.5955
R20541 OUT3.n6 OUT3.t31 26.5955
R20542 OUT3.n6 OUT3.t47 26.5955
R20543 OUT3.n8 OUT3.t45 26.5955
R20544 OUT3.n8 OUT3.t57 26.5955
R20545 OUT3.n10 OUT3.t34 26.5955
R20546 OUT3.n10 OUT3.t28 26.5955
R20547 OUT3.n12 OUT3.t55 26.5955
R20548 OUT3.n12 OUT3.t16 26.5955
R20549 OUT3.n14 OUT3.t14 26.5955
R20550 OUT3.n14 OUT3.t32 26.5955
R20551 OUT3.n16 OUT3.t39 26.5955
R20552 OUT3.n16 OUT3.t53 26.5955
R20553 OUT3.n46 OUT3.t51 25.6105
R20554 OUT3.n171 OUT3.t91 24.9236
R20555 OUT3.n171 OUT3.t117 24.9236
R20556 OUT3.n158 OUT3.t101 24.9236
R20557 OUT3.n158 OUT3.t76 24.9236
R20558 OUT3.n159 OUT3.t115 24.9236
R20559 OUT3.n159 OUT3.t88 24.9236
R20560 OUT3.n161 OUT3.t86 24.9236
R20561 OUT3.n161 OUT3.t99 24.9236
R20562 OUT3.n163 OUT3.t107 24.9236
R20563 OUT3.n163 OUT3.t123 24.9236
R20564 OUT3.n165 OUT3.t121 24.9236
R20565 OUT3.n165 OUT3.t79 24.9236
R20566 OUT3.n167 OUT3.t77 24.9236
R20567 OUT3.n167 OUT3.t105 24.9236
R20568 OUT3.n169 OUT3.t68 24.9236
R20569 OUT3.n169 OUT3.t93 24.9236
R20570 OUT3.n112 OUT3.t102 24.9236
R20571 OUT3.n112 OUT3.t64 24.9236
R20572 OUT3.n113 OUT3.t126 24.9236
R20573 OUT3.n113 OUT3.t89 24.9236
R20574 OUT3.n115 OUT3.t80 24.9236
R20575 OUT3.n115 OUT3.t110 24.9236
R20576 OUT3.n117 OUT3.t81 24.9236
R20577 OUT3.n117 OUT3.t97 24.9236
R20578 OUT3.n119 OUT3.t95 24.9236
R20579 OUT3.n119 OUT3.t113 24.9236
R20580 OUT3.n121 OUT3.t120 24.9236
R20581 OUT3.n121 OUT3.t70 24.9236
R20582 OUT3.n123 OUT3.t75 24.9236
R20583 OUT3.n123 OUT3.t104 24.9236
R20584 OUT3.n70 OUT3.t84 24.9236
R20585 OUT3.n70 OUT3.t65 24.9236
R20586 OUT3.n71 OUT3.t100 24.9236
R20587 OUT3.n71 OUT3.t116 24.9236
R20588 OUT3.n73 OUT3.t124 24.9236
R20589 OUT3.n73 OUT3.t87 24.9236
R20590 OUT3.n75 OUT3.t72 24.9236
R20591 OUT3.n75 OUT3.t98 24.9236
R20592 OUT3.n77 OUT3.t106 24.9236
R20593 OUT3.n77 OUT3.t122 24.9236
R20594 OUT3.n79 OUT3.t66 24.9236
R20595 OUT3.n79 OUT3.t78 24.9236
R20596 OUT3.n81 OUT3.t109 24.9236
R20597 OUT3.n81 OUT3.t85 24.9236
R20598 OUT3.n37 OUT3.t74 24.9236
R20599 OUT3.n37 OUT3.t83 24.9236
R20600 OUT3.n24 OUT3.t90 24.9236
R20601 OUT3.n24 OUT3.t103 24.9236
R20602 OUT3.n25 OUT3.t111 24.9236
R20603 OUT3.n25 OUT3.t127 24.9236
R20604 OUT3.n27 OUT3.t125 24.9236
R20605 OUT3.n27 OUT3.t73 24.9236
R20606 OUT3.n29 OUT3.t114 24.9236
R20607 OUT3.n29 OUT3.t108 24.9236
R20608 OUT3.n31 OUT3.t71 24.9236
R20609 OUT3.n31 OUT3.t96 24.9236
R20610 OUT3.n33 OUT3.t94 24.9236
R20611 OUT3.n33 OUT3.t112 24.9236
R20612 OUT3.n35 OUT3.t119 24.9236
R20613 OUT3.n35 OUT3.t69 24.9236
R20614 OUT3.n68 OUT3.t67 24.7196
R20615 OUT3.n105 OUT3.t2 24.6255
R20616 OUT3.n68 OUT3.t92 23.9564
R20617 OUT3.n127 OUT3.t82 23.1655
R20618 OUT3.n103 OUT3.t38 19.1164
R20619 OUT3.n126 OUT3.n125 13.8467
R20620 OUT3 OUT3.n174 11.4429
R20621 OUT3 OUT3.n129 11.4429
R20622 OUT3 OUT3.n83 11.4429
R20623 OUT3 OUT3.n40 11.4429
R20624 OUT3.n125 OUT3.t118 11.0774
R20625 OUT3.n47 OUT3.t12 10.8355
R20626 OUT3.n106 OUT3.n105 9.3005
R20627 OUT3.n110 OUT3.n109 9.3005
R20628 OUT3.n128 OUT3.n127 8.77252
R20629 OUT3.n136 OUT3.n135 8.76605
R20630 OUT3.n2 OUT3.n1 8.76605
R20631 OUT3.n50 OUT3.n49 8.70762
R20632 OUT3.n49 OUT3.n48 8.69892
R20633 OUT3.n172 OUT3.n171 7.87147
R20634 OUT3.n38 OUT3.n37 7.87147
R20635 OUT3.n48 OUT3.n47 7.77627
R20636 OUT3.n104 OUT3.n103 7.29637
R20637 OUT3.n69 OUT3.n68 6.88889
R20638 OUT3.n85 OUT3.n69 4.758
R20639 OUT3.n128 OUT3.n111 4.6505
R20640 OUT3.n107 OUT3.n106 4.6505
R20641 OUT3.n39 OUT3.n23 4.6505
R20642 OUT3.n20 OUT3.n19 4.6505
R20643 OUT3.n3 OUT3.n2 4.26717
R20644 OUT3.n175 OUT3 3.10353
R20645 OUT3.n130 OUT3 3.10353
R20646 OUT3.n84 OUT3 3.10353
R20647 OUT3.n41 OUT3 3.10353
R20648 OUT3.n173 OUT3.n157 3.1005
R20649 OUT3.n137 OUT3.n136 3.1005
R20650 OUT3.n155 OUT3.n154 3.1005
R20651 OUT3.n66 OUT3.n65 2.75
R20652 OUT3.n154 OUT3.n153 2.71565
R20653 OUT3.n106 OUT3.n102 2.71565
R20654 OUT3.n65 OUT3.n64 2.71565
R20655 OUT3.n19 OUT3.n18 2.71565
R20656 OUT3.n66 OUT3.n50 2.69896
R20657 OUT3.n105 OUT3.n104 1.9705
R20658 OUT3.n174 OUT3 1.74595
R20659 OUT3 OUT3.n173 1.74595
R20660 OUT3.n129 OUT3 1.74595
R20661 OUT3 OUT3.n128 1.74595
R20662 OUT3.n83 OUT3 1.74595
R20663 OUT3.n40 OUT3 1.74595
R20664 OUT3 OUT3.n39 1.74595
R20665 OUT3.n127 OUT3.n126 1.74224
R20666 OUT3.n181 OUT3.n180 0.810582
R20667 OUT3 OUT3.n183 0.597838
R20668 OUT3.n183 OUT3.n182 0.531962
R20669 OUT3.n182 OUT3.n181 0.531962
R20670 OUT3.n182 OUT3.n86 0.475506
R20671 OUT3 OUT3.n69 0.388379
R20672 OUT3.n173 OUT3.n172 0.300854
R20673 OUT3.n39 OUT3.n38 0.300854
R20674 OUT3.n183 OUT3.n45 0.275505
R20675 OUT3.n181 OUT3.n134 0.263005
R20676 OUT3.n180 OUT3.n179 0.1755
R20677 OUT3.n134 OUT3.n133 0.1755
R20678 OUT3.n45 OUT3.n44 0.1755
R20679 OUT3.n176 OUT3.n157 0.11675
R20680 OUT3.n131 OUT3.n111 0.11675
R20681 OUT3.n42 OUT3.n23 0.11675
R20682 OUT3.n132 OUT3.n107 0.10425
R20683 OUT3.n178 OUT3.n155 0.09175
R20684 OUT3.n43 OUT3.n20 0.09175
R20685 OUT3.n86 OUT3.n66 0.0855244
R20686 OUT3.n49 OUT3.n46 0.0578287
R20687 OUT3.n86 OUT3.n85 0.0505
R20688 OUT3.n155 OUT3.n139 0.04425
R20689 OUT3.n20 OUT3.n4 0.04425
R20690 OUT3.n107 OUT3.n88 0.043
R20691 OUT3.n111 OUT3.n110 0.03175
R20692 OUT3.n139 OUT3.n137 0.028
R20693 OUT3.n4 OUT3.n0 0.028
R20694 OUT3.n178 OUT3.n176 0.0255
R20695 OUT3.n157 OUT3.n156 0.0255
R20696 OUT3.n43 OUT3.n42 0.0255
R20697 OUT3.n23 OUT3.n22 0.0255
R20698 OUT3.n132 OUT3.n131 0.013
R20699 OUT3.n88 OUT3.n87 0.00450862
R20700 OUT3.n139 OUT3.n138 0.0025557
R20701 OUT3.n4 OUT3.n3 0.0025557
R20702 OUT3.n176 OUT3.n175 0.00053521
R20703 OUT3.n131 OUT3.n130 0.00053521
R20704 OUT3.n85 OUT3.n84 0.00053521
R20705 OUT3.n42 OUT3.n41 0.00053521
R20706 OUT3.n178 OUT3.n177 0.00050852
R20707 OUT3.n132 OUT3.n108 0.00050852
R20708 OUT3.n86 OUT3.n67 0.00050852
R20709 OUT3.n43 OUT3.n21 0.00050852
R20710 OUT3.n179 OUT3.n178 0.000500999
R20711 OUT3.n133 OUT3.n132 0.000500999
R20712 OUT3.n44 OUT3.n43 0.000500999
R20713 frontAnalog_v0p0p1_15.x63.A.n2 frontAnalog_v0p0p1_15.x63.A.t4 260.322
R20714 frontAnalog_v0p0p1_15.x63.A.n4 frontAnalog_v0p0p1_15.x63.A.t5 233.888
R20715 frontAnalog_v0p0p1_15.x63.A.n2 frontAnalog_v0p0p1_15.x63.A.t6 175.169
R20716 frontAnalog_v0p0p1_15.x63.A.n3 frontAnalog_v0p0p1_15.x63.A.t7 159.725
R20717 frontAnalog_v0p0p1_15.x63.A.n1 frontAnalog_v0p0p1_15.x63.A.t2 17.4109
R20718 frontAnalog_v0p0p1_15.x63.A.n0 frontAnalog_v0p0p1_15.x63.A.n2 9.75129
R20719 frontAnalog_v0p0p1_15.x63.A.n1 frontAnalog_v0p0p1_15.x63.A.t1 9.6037
R20720 frontAnalog_v0p0p1_15.x63.A.n0 frontAnalog_v0p0p1_15.x63.A 2.33338
R20721 frontAnalog_v0p0p1_15.x63.A.n5 frontAnalog_v0p0p1_15.x63.A.t3 8.40929
R20722 frontAnalog_v0p0p1_15.x63.A.n3 frontAnalog_v0p0p1_15.x63.A.t0 8.06629
R20723 frontAnalog_v0p0p1_15.x63.A.n4 frontAnalog_v0p0p1_15.x63.A.n3 1.73501
R20724 frontAnalog_v0p0p1_15.x63.A.n1 frontAnalog_v0p0p1_15.x63.A.n4 0.99025
R20725 frontAnalog_v0p0p1_15.x63.A.n5 frontAnalog_v0p0p1_15.x63.A.n1 0.853186
R20726 frontAnalog_v0p0p1_15.x63.A frontAnalog_v0p0p1_15.x63.A.n0 0.349517
R20727 frontAnalog_v0p0p1_15.x63.A frontAnalog_v0p0p1_15.x63.A.n5 0.24425
R20728 OUT0.n122 OUT0.n120 145.809
R20729 OUT0.n65 OUT0.n63 145.809
R20730 OUT0.n25 OUT0.n23 145.809
R20731 OUT0.n102 OUT0.n100 145.808
R20732 OUT0.n65 OUT0.n64 107.409
R20733 OUT0.n67 OUT0.n66 107.409
R20734 OUT0.n69 OUT0.n68 107.409
R20735 OUT0.n71 OUT0.n70 107.409
R20736 OUT0.n73 OUT0.n72 107.409
R20737 OUT0.n75 OUT0.n74 107.409
R20738 OUT0.n25 OUT0.n24 107.409
R20739 OUT0.n27 OUT0.n26 107.409
R20740 OUT0.n29 OUT0.n28 107.409
R20741 OUT0.n31 OUT0.n30 107.409
R20742 OUT0.n33 OUT0.n32 107.409
R20743 OUT0.n35 OUT0.n34 107.409
R20744 OUT0.n122 OUT0.n121 107.407
R20745 OUT0.n124 OUT0.n123 107.407
R20746 OUT0.n126 OUT0.n125 107.407
R20747 OUT0.n128 OUT0.n127 107.407
R20748 OUT0.n130 OUT0.n129 107.407
R20749 OUT0.n132 OUT0.n131 107.407
R20750 OUT0.n102 OUT0.n101 107.407
R20751 OUT0.n104 OUT0.n103 107.407
R20752 OUT0.n106 OUT0.n105 107.407
R20753 OUT0.n108 OUT0.n107 107.407
R20754 OUT0.n110 OUT0.n109 107.407
R20755 OUT0.n112 OUT0.n111 107.407
R20756 OUT0.n138 OUT0.n136 87.1779
R20757 OUT0.n83 OUT0.n81 87.1779
R20758 OUT0.n44 OUT0.n42 87.1779
R20759 OUT0.n4 OUT0.n2 87.1779
R20760 OUT0.n54 OUT0.n53 52.82
R20761 OUT0.n14 OUT0.n13 52.82
R20762 OUT0.n138 OUT0.n137 52.82
R20763 OUT0.n140 OUT0.n139 52.82
R20764 OUT0.n142 OUT0.n141 52.82
R20765 OUT0.n144 OUT0.n143 52.82
R20766 OUT0.n146 OUT0.n145 52.82
R20767 OUT0.n148 OUT0.n147 52.82
R20768 OUT0.n83 OUT0.n82 52.82
R20769 OUT0.n85 OUT0.n84 52.82
R20770 OUT0.n87 OUT0.n86 52.82
R20771 OUT0.n89 OUT0.n88 52.82
R20772 OUT0.n91 OUT0.n90 52.82
R20773 OUT0.n93 OUT0.n92 52.82
R20774 OUT0.n44 OUT0.n43 52.82
R20775 OUT0.n46 OUT0.n45 52.82
R20776 OUT0.n48 OUT0.n47 52.82
R20777 OUT0.n50 OUT0.n49 52.82
R20778 OUT0.n52 OUT0.n51 52.82
R20779 OUT0.n4 OUT0.n3 52.82
R20780 OUT0.n6 OUT0.n5 52.82
R20781 OUT0.n8 OUT0.n7 52.82
R20782 OUT0.n10 OUT0.n9 52.82
R20783 OUT0.n12 OUT0.n11 52.82
R20784 OUT0 OUT0.n149 51.0745
R20785 OUT0 OUT0.n94 51.0745
R20786 OUT0.n124 OUT0.n122 38.4005
R20787 OUT0.n126 OUT0.n124 38.4005
R20788 OUT0.n128 OUT0.n126 38.4005
R20789 OUT0.n130 OUT0.n128 38.4005
R20790 OUT0.n132 OUT0.n130 38.4005
R20791 OUT0.n133 OUT0.n132 38.4005
R20792 OUT0.n104 OUT0.n102 38.4005
R20793 OUT0.n106 OUT0.n104 38.4005
R20794 OUT0.n108 OUT0.n106 38.4005
R20795 OUT0.n110 OUT0.n108 38.4005
R20796 OUT0.n112 OUT0.n110 38.4005
R20797 OUT0.n113 OUT0.n112 38.4005
R20798 OUT0.n67 OUT0.n65 38.4005
R20799 OUT0.n69 OUT0.n67 38.4005
R20800 OUT0.n71 OUT0.n69 38.4005
R20801 OUT0.n73 OUT0.n71 38.4005
R20802 OUT0.n75 OUT0.n73 38.4005
R20803 OUT0.n76 OUT0.n75 38.4005
R20804 OUT0.n27 OUT0.n25 38.4005
R20805 OUT0.n29 OUT0.n27 38.4005
R20806 OUT0.n31 OUT0.n29 38.4005
R20807 OUT0.n33 OUT0.n31 38.4005
R20808 OUT0.n35 OUT0.n33 38.4005
R20809 OUT0.n36 OUT0.n35 38.4005
R20810 OUT0.n140 OUT0.n138 34.3584
R20811 OUT0.n142 OUT0.n140 34.3584
R20812 OUT0.n144 OUT0.n142 34.3584
R20813 OUT0.n146 OUT0.n144 34.3584
R20814 OUT0.n148 OUT0.n146 34.3584
R20815 OUT0.n150 OUT0.n148 34.3584
R20816 OUT0.n85 OUT0.n83 34.3584
R20817 OUT0.n87 OUT0.n85 34.3584
R20818 OUT0.n89 OUT0.n87 34.3584
R20819 OUT0.n91 OUT0.n89 34.3584
R20820 OUT0.n93 OUT0.n91 34.3584
R20821 OUT0.n95 OUT0.n93 34.3584
R20822 OUT0.n46 OUT0.n44 34.3584
R20823 OUT0.n48 OUT0.n46 34.3584
R20824 OUT0.n50 OUT0.n48 34.3584
R20825 OUT0.n52 OUT0.n50 34.3584
R20826 OUT0.n54 OUT0.n52 34.3584
R20827 OUT0.n58 OUT0.n54 34.3584
R20828 OUT0.n6 OUT0.n4 34.3584
R20829 OUT0.n8 OUT0.n6 34.3584
R20830 OUT0.n10 OUT0.n8 34.3584
R20831 OUT0.n12 OUT0.n10 34.3584
R20832 OUT0.n14 OUT0.n12 34.3584
R20833 OUT0.n18 OUT0.n14 34.3584
R20834 OUT0.n118 OUT0.t41 26.5955
R20835 OUT0.n118 OUT0.t54 26.5955
R20836 OUT0.n120 OUT0.t39 26.5955
R20837 OUT0.n120 OUT0.t11 26.5955
R20838 OUT0.n121 OUT0.t61 26.5955
R20839 OUT0.n121 OUT0.t27 26.5955
R20840 OUT0.n123 OUT0.t6 26.5955
R20841 OUT0.n123 OUT0.t47 26.5955
R20842 OUT0.n125 OUT0.t17 26.5955
R20843 OUT0.n125 OUT0.t35 26.5955
R20844 OUT0.n127 OUT0.t33 26.5955
R20845 OUT0.n127 OUT0.t50 26.5955
R20846 OUT0.n129 OUT0.t56 26.5955
R20847 OUT0.n129 OUT0.t22 26.5955
R20848 OUT0.n131 OUT0.t3 26.5955
R20849 OUT0.n131 OUT0.t43 26.5955
R20850 OUT0.n99 OUT0.t2 26.5955
R20851 OUT0.n99 OUT0.t31 26.5955
R20852 OUT0.n100 OUT0.t21 26.5955
R20853 OUT0.n100 OUT0.t30 26.5955
R20854 OUT0.n101 OUT0.t37 26.5955
R20855 OUT0.n101 OUT0.t10 26.5955
R20856 OUT0.n103 OUT0.t52 26.5955
R20857 OUT0.n103 OUT0.t24 26.5955
R20858 OUT0.n105 OUT0.t23 26.5955
R20859 OUT0.n105 OUT0.t36 26.5955
R20860 OUT0.n107 OUT0.t44 26.5955
R20861 OUT0.n107 OUT0.t58 26.5955
R20862 OUT0.n109 OUT0.t57 26.5955
R20863 OUT0.n109 OUT0.t12 26.5955
R20864 OUT0.n111 OUT0.t46 26.5955
R20865 OUT0.n111 OUT0.t14 26.5955
R20866 OUT0.n62 OUT0.t8 26.5955
R20867 OUT0.n62 OUT0.t42 26.5955
R20868 OUT0.n63 OUT0.t28 26.5955
R20869 OUT0.n63 OUT0.t40 26.5955
R20870 OUT0.n64 OUT0.t38 26.5955
R20871 OUT0.n64 OUT0.t62 26.5955
R20872 OUT0.n66 OUT0.t59 26.5955
R20873 OUT0.n66 OUT0.t25 26.5955
R20874 OUT0.n68 OUT0.t51 26.5955
R20875 OUT0.n68 OUT0.t19 26.5955
R20876 OUT0.n70 OUT0.t15 26.5955
R20877 OUT0.n70 OUT0.t34 26.5955
R20878 OUT0.n72 OUT0.t32 26.5955
R20879 OUT0.n72 OUT0.t49 26.5955
R20880 OUT0.n74 OUT0.t55 26.5955
R20881 OUT0.n74 OUT0.t4 26.5955
R20882 OUT0.n22 OUT0.t7 26.5955
R20883 OUT0.n22 OUT0.t20 26.5955
R20884 OUT0.n23 OUT0.t26 26.5955
R20885 OUT0.n23 OUT0.t48 26.5955
R20886 OUT0.n24 OUT0.t45 26.5955
R20887 OUT0.n24 OUT0.t60 26.5955
R20888 OUT0.n26 OUT0.t1 26.5955
R20889 OUT0.n26 OUT0.t13 26.5955
R20890 OUT0.n28 OUT0.t18 26.5955
R20891 OUT0.n28 OUT0.t53 26.5955
R20892 OUT0.n30 OUT0.t29 26.5955
R20893 OUT0.n30 OUT0.t0 26.5955
R20894 OUT0.n32 OUT0.t5 26.5955
R20895 OUT0.n32 OUT0.t16 26.5955
R20896 OUT0.n34 OUT0.t63 26.5955
R20897 OUT0.n34 OUT0.t9 26.5955
R20898 OUT0.n149 OUT0.t105 24.9236
R20899 OUT0.n149 OUT0.t118 24.9236
R20900 OUT0.n136 OUT0.t103 24.9236
R20901 OUT0.n136 OUT0.t75 24.9236
R20902 OUT0.n137 OUT0.t125 24.9236
R20903 OUT0.n137 OUT0.t91 24.9236
R20904 OUT0.n139 OUT0.t70 24.9236
R20905 OUT0.n139 OUT0.t111 24.9236
R20906 OUT0.n141 OUT0.t81 24.9236
R20907 OUT0.n141 OUT0.t99 24.9236
R20908 OUT0.n143 OUT0.t97 24.9236
R20909 OUT0.n143 OUT0.t114 24.9236
R20910 OUT0.n145 OUT0.t120 24.9236
R20911 OUT0.n145 OUT0.t86 24.9236
R20912 OUT0.n147 OUT0.t67 24.9236
R20913 OUT0.n147 OUT0.t107 24.9236
R20914 OUT0.n94 OUT0.t66 24.9236
R20915 OUT0.n94 OUT0.t95 24.9236
R20916 OUT0.n81 OUT0.t85 24.9236
R20917 OUT0.n81 OUT0.t94 24.9236
R20918 OUT0.n82 OUT0.t101 24.9236
R20919 OUT0.n82 OUT0.t74 24.9236
R20920 OUT0.n84 OUT0.t116 24.9236
R20921 OUT0.n84 OUT0.t88 24.9236
R20922 OUT0.n86 OUT0.t87 24.9236
R20923 OUT0.n86 OUT0.t100 24.9236
R20924 OUT0.n88 OUT0.t108 24.9236
R20925 OUT0.n88 OUT0.t122 24.9236
R20926 OUT0.n90 OUT0.t121 24.9236
R20927 OUT0.n90 OUT0.t76 24.9236
R20928 OUT0.n92 OUT0.t110 24.9236
R20929 OUT0.n92 OUT0.t78 24.9236
R20930 OUT0.n55 OUT0.t72 24.9236
R20931 OUT0.n55 OUT0.t106 24.9236
R20932 OUT0.n42 OUT0.t92 24.9236
R20933 OUT0.n42 OUT0.t104 24.9236
R20934 OUT0.n43 OUT0.t102 24.9236
R20935 OUT0.n43 OUT0.t126 24.9236
R20936 OUT0.n45 OUT0.t123 24.9236
R20937 OUT0.n45 OUT0.t89 24.9236
R20938 OUT0.n47 OUT0.t115 24.9236
R20939 OUT0.n47 OUT0.t83 24.9236
R20940 OUT0.n49 OUT0.t79 24.9236
R20941 OUT0.n49 OUT0.t98 24.9236
R20942 OUT0.n51 OUT0.t96 24.9236
R20943 OUT0.n51 OUT0.t113 24.9236
R20944 OUT0.n53 OUT0.t119 24.9236
R20945 OUT0.n53 OUT0.t68 24.9236
R20946 OUT0.n15 OUT0.t71 24.9236
R20947 OUT0.n15 OUT0.t84 24.9236
R20948 OUT0.n2 OUT0.t90 24.9236
R20949 OUT0.n2 OUT0.t112 24.9236
R20950 OUT0.n3 OUT0.t109 24.9236
R20951 OUT0.n3 OUT0.t124 24.9236
R20952 OUT0.n5 OUT0.t65 24.9236
R20953 OUT0.n5 OUT0.t77 24.9236
R20954 OUT0.n7 OUT0.t82 24.9236
R20955 OUT0.n7 OUT0.t117 24.9236
R20956 OUT0.n9 OUT0.t93 24.9236
R20957 OUT0.n9 OUT0.t64 24.9236
R20958 OUT0.n11 OUT0.t69 24.9236
R20959 OUT0.n11 OUT0.t80 24.9236
R20960 OUT0.n13 OUT0.t127 24.9236
R20961 OUT0.n13 OUT0.t73 24.9236
R20962 OUT0 OUT0.n150 11.4429
R20963 OUT0 OUT0.n95 11.4429
R20964 OUT0 OUT0.n58 11.4429
R20965 OUT0 OUT0.n18 11.4429
R20966 OUT0.n77 OUT0.n62 8.55118
R20967 OUT0.n37 OUT0.n22 8.55118
R20968 OUT0.n114 OUT0.n99 8.55117
R20969 OUT0.n119 OUT0.n118 8.47293
R20970 OUT0.n56 OUT0.n55 7.80093
R20971 OUT0.n16 OUT0.n15 7.80093
R20972 OUT0.n78 OUT0.n77 3.20954
R20973 OUT0.n38 OUT0.n37 3.20953
R20974 OUT0.n115 OUT0.n114 3.20289
R20975 OUT0.n151 OUT0 3.10353
R20976 OUT0.n96 OUT0 3.10353
R20977 OUT0.n59 OUT0 3.10353
R20978 OUT0.n19 OUT0 3.10353
R20979 OUT0.n135 OUT0.n134 3.1005
R20980 OUT0.n57 OUT0.n41 3.1005
R20981 OUT0.n17 OUT0.n1 3.1005
R20982 OUT0.n134 OUT0.n133 2.71565
R20983 OUT0.n114 OUT0.n113 2.13383
R20984 OUT0.n77 OUT0.n76 2.13383
R20985 OUT0.n37 OUT0.n36 2.13383
R20986 OUT0.n150 OUT0 1.74595
R20987 OUT0.n95 OUT0 1.74595
R20988 OUT0.n58 OUT0.n57 1.16414
R20989 OUT0.n18 OUT0.n17 1.16414
R20990 OUT0.n157 OUT0.n156 1.07337
R20991 OUT0.n158 OUT0.n157 0.69375
R20992 OUT0.n159 OUT0.n158 0.68905
R20993 OUT0.n56 OUT0 0.488972
R20994 OUT0.n16 OUT0 0.488972
R20995 OUT0.n158 OUT0.n79 0.414635
R20996 OUT0.n157 OUT0.n116 0.382465
R20997 OUT0.n159 OUT0.n39 0.368576
R20998 OUT0 OUT0.n159 0.281623
R20999 OUT0.n134 OUT0.n119 0.196887
R21000 OUT0.n79 OUT0.n78 0.157252
R21001 OUT0.n39 OUT0.n38 0.139891
R21002 OUT0.n156 OUT0.n155 0.139389
R21003 OUT0.n116 OUT0.n115 0.132946
R21004 OUT0.n60 OUT0.n41 0.113
R21005 OUT0.n20 OUT0.n1 0.113
R21006 OUT0.n154 OUT0.n135 0.101889
R21007 OUT0.n57 OUT0.n56 0.0893205
R21008 OUT0.n17 OUT0.n16 0.0893205
R21009 OUT0.n154 OUT0.n152 0.0282778
R21010 OUT0.n135 OUT0.n117 0.0268889
R21011 OUT0.n98 OUT0.n97 0.0213333
R21012 OUT0.n61 OUT0.n60 0.0143889
R21013 OUT0.n21 OUT0.n20 0.0143889
R21014 OUT0.n115 OUT0.n98 0.00100004
R21015 OUT0.n38 OUT0.n21 0.00100004
R21016 OUT0.n78 OUT0.n61 0.00100004
R21017 OUT0.n152 OUT0.n151 0.000513335
R21018 OUT0.n97 OUT0.n96 0.000513335
R21019 OUT0.n60 OUT0.n59 0.000513218
R21020 OUT0.n20 OUT0.n19 0.000513218
R21021 OUT0.n98 OUT0.n80 0.00050517
R21022 OUT0.n154 OUT0.n153 0.000504838
R21023 OUT0.n61 OUT0.n40 0.000504838
R21024 OUT0.n21 OUT0.n0 0.000504838
R21025 OUT0.n155 OUT0.n154 0.000501713
R21026 frontAnalog_v0p0p1_10.Q.t11 frontAnalog_v0p0p1_10.Q.t13 618.109
R21027 frontAnalog_v0p0p1_10.Q.n12 frontAnalog_v0p0p1_10.Q.t6 259.74
R21028 frontAnalog_v0p0p1_10.Q frontAnalog_v0p0p1_10.Q.t11 253.56
R21029 frontAnalog_v0p0p1_10.Q.n0 frontAnalog_v0p0p1_10.Q.t9 228.899
R21030 frontAnalog_v0p0p1_10.Q.n19 frontAnalog_v0p0p1_10.Q.t7 180.286
R21031 frontAnalog_v0p0p1_10.Q.n0 frontAnalog_v0p0p1_10.Q.t8 159.411
R21032 frontAnalog_v0p0p1_10.Q.n12 frontAnalog_v0p0p1_10.Q.t10 157.083
R21033 frontAnalog_v0p0p1_10.Q.n26 frontAnalog_v0p0p1_10.Q.t5 117.314
R21034 frontAnalog_v0p0p1_10.Q.n20 frontAnalog_v0p0p1_10.Q.t14 111.091
R21035 frontAnalog_v0p0p1_10.Q.n26 frontAnalog_v0p0p1_10.Q.t12 110.853
R21036 frontAnalog_v0p0p1_10.Q.n24 frontAnalog_v0p0p1_10.Q 37.6855
R21037 frontAnalog_v0p0p1_10.Q.n27 frontAnalog_v0p0p1_10.Q.t2 17.6181
R21038 frontAnalog_v0p0p1_10.Q.n29 frontAnalog_v0p0p1_10.Q.t4 14.2865
R21039 frontAnalog_v0p0p1_10.Q.n31 frontAnalog_v0p0p1_10.Q.t1 14.283
R21040 frontAnalog_v0p0p1_10.Q.n31 frontAnalog_v0p0p1_10.Q.t0 14.283
R21041 frontAnalog_v0p0p1_10.Q.n21 frontAnalog_v0p0p1_10.Q.n20 9.3005
R21042 frontAnalog_v0p0p1_10.Q frontAnalog_v0p0p1_10.Q.n11 9.3005
R21043 frontAnalog_v0p0p1_10.Q.n33 frontAnalog_v0p0p1_10.Q.t3 8.77744
R21044 frontAnalog_v0p0p1_10.Q.n22 frontAnalog_v0p0p1_10.Q.n21 7.80966
R21045 frontAnalog_v0p0p1_10.Q.n13 frontAnalog_v0p0p1_10.Q.n12 7.57248
R21046 frontAnalog_v0p0p1_10.Q.n1 frontAnalog_v0p0p1_10.Q.n0 7.36978
R21047 frontAnalog_v0p0p1_10.Q.n20 frontAnalog_v0p0p1_10.Q.n19 6.53562
R21048 frontAnalog_v0p0p1_10.Q.n13 frontAnalog_v0p0p1_10.Q 4.8645
R21049 frontAnalog_v0p0p1_10.Q.n34 frontAnalog_v0p0p1_10.Q.n25 4.31885
R21050 frontAnalog_v0p0p1_10.Q.n3 frontAnalog_v0p0p1_10.Q.n2 3.46717
R21051 frontAnalog_v0p0p1_10.Q.n4 frontAnalog_v0p0p1_10.Q.n3 3.03286
R21052 frontAnalog_v0p0p1_10.Q.n18 frontAnalog_v0p0p1_10.Q.n17 2.32777
R21053 frontAnalog_v0p0p1_10.Q.n22 frontAnalog_v0p0p1_10.Q.n16 2.19001
R21054 frontAnalog_v0p0p1_10.Q.n17 frontAnalog_v0p0p1_10.Q 1.4966
R21055 frontAnalog_v0p0p1_10.Q.n23 frontAnalog_v0p0p1_10.Q.n9 1.36032
R21056 frontAnalog_v0p0p1_10.Q.n33 frontAnalog_v0p0p1_10.Q.n32 1.20426
R21057 frontAnalog_v0p0p1_10.Q.n23 frontAnalog_v0p0p1_10.Q.n22 1.07639
R21058 frontAnalog_v0p0p1_10.Q.n3 frontAnalog_v0p0p1_10.Q.n1 1.06717
R21059 frontAnalog_v0p0p1_10.Q.n2 frontAnalog_v0p0p1_10.Q 1.06717
R21060 frontAnalog_v0p0p1_10.Q.n9 frontAnalog_v0p0p1_10.Q.n8 0.71595
R21061 frontAnalog_v0p0p1_10.Q.n21 frontAnalog_v0p0p1_10.Q.n18 0.499201
R21062 frontAnalog_v0p0p1_10.Q.n25 frontAnalog_v0p0p1_10.Q.n24 0.435179
R21063 frontAnalog_v0p0p1_10.Q.n34 frontAnalog_v0p0p1_10.Q.n33 0.325111
R21064 frontAnalog_v0p0p1_10.Q.n30 frontAnalog_v0p0p1_10.Q.n29 0.301242
R21065 frontAnalog_v0p0p1_10.Q.n9 frontAnalog_v0p0p1_10.Q 0.221483
R21066 frontAnalog_v0p0p1_10.Q.n25 frontAnalog_v0p0p1_10.Q 0.20675
R21067 frontAnalog_v0p0p1_10.Q.n28 frontAnalog_v0p0p1_10.Q.n26 0.159555
R21068 frontAnalog_v0p0p1_10.Q.n32 frontAnalog_v0p0p1_10.Q.n31 0.106617
R21069 frontAnalog_v0p0p1_10.Q.n30 frontAnalog_v0p0p1_10.Q.n28 0.0796167
R21070 frontAnalog_v0p0p1_10.Q.n32 frontAnalog_v0p0p1_10.Q.n30 0.0480595
R21071 frontAnalog_v0p0p1_10.Q frontAnalog_v0p0p1_10.Q.n34 0.0469368
R21072 frontAnalog_v0p0p1_10.Q.n11 frontAnalog_v0p0p1_10.Q.n10 0.0301875
R21073 frontAnalog_v0p0p1_10.Q.n16 frontAnalog_v0p0p1_10.Q.n15 0.0205312
R21074 frontAnalog_v0p0p1_10.Q.n6 frontAnalog_v0p0p1_10.Q.n5 0.00618182
R21075 frontAnalog_v0p0p1_10.Q.n5 frontAnalog_v0p0p1_10.Q.n4 0.00555107
R21076 frontAnalog_v0p0p1_10.Q.n7 frontAnalog_v0p0p1_10.Q.n6 0.00530477
R21077 frontAnalog_v0p0p1_10.Q.n15 frontAnalog_v0p0p1_10.Q.n14 0.00210765
R21078 frontAnalog_v0p0p1_10.Q.n14 frontAnalog_v0p0p1_10.Q.n13 0.00133438
R21079 frontAnalog_v0p0p1_10.Q.n8 frontAnalog_v0p0p1_10.Q.n7 0.00101192
R21080 frontAnalog_v0p0p1_10.Q.n14 frontAnalog_v0p0p1_10.Q.n10 0.00100001
R21081 frontAnalog_v0p0p1_10.Q.n24 frontAnalog_v0p0p1_10.Q.n23 0.000507778
R21082 frontAnalog_v0p0p1_10.Q.n28 frontAnalog_v0p0p1_10.Q.n27 0.000504658
R21083 OUT2.n122 OUT2.n120 145.809
R21084 OUT2.n65 OUT2.n63 145.809
R21085 OUT2.n25 OUT2.n23 145.809
R21086 OUT2.n102 OUT2.n100 145.808
R21087 OUT2.n65 OUT2.n64 107.409
R21088 OUT2.n67 OUT2.n66 107.409
R21089 OUT2.n69 OUT2.n68 107.409
R21090 OUT2.n71 OUT2.n70 107.409
R21091 OUT2.n73 OUT2.n72 107.409
R21092 OUT2.n75 OUT2.n74 107.409
R21093 OUT2.n25 OUT2.n24 107.409
R21094 OUT2.n27 OUT2.n26 107.409
R21095 OUT2.n29 OUT2.n28 107.409
R21096 OUT2.n31 OUT2.n30 107.409
R21097 OUT2.n33 OUT2.n32 107.409
R21098 OUT2.n35 OUT2.n34 107.409
R21099 OUT2.n122 OUT2.n121 107.407
R21100 OUT2.n124 OUT2.n123 107.407
R21101 OUT2.n126 OUT2.n125 107.407
R21102 OUT2.n128 OUT2.n127 107.407
R21103 OUT2.n130 OUT2.n129 107.407
R21104 OUT2.n132 OUT2.n131 107.407
R21105 OUT2.n102 OUT2.n101 107.407
R21106 OUT2.n104 OUT2.n103 107.407
R21107 OUT2.n106 OUT2.n105 107.407
R21108 OUT2.n108 OUT2.n107 107.407
R21109 OUT2.n110 OUT2.n109 107.407
R21110 OUT2.n112 OUT2.n111 107.407
R21111 OUT2.n138 OUT2.n136 87.1779
R21112 OUT2.n83 OUT2.n81 87.1779
R21113 OUT2.n44 OUT2.n42 87.1779
R21114 OUT2.n4 OUT2.n2 87.1779
R21115 OUT2.n54 OUT2.n53 52.82
R21116 OUT2.n14 OUT2.n13 52.82
R21117 OUT2.n138 OUT2.n137 52.82
R21118 OUT2.n140 OUT2.n139 52.82
R21119 OUT2.n142 OUT2.n141 52.82
R21120 OUT2.n144 OUT2.n143 52.82
R21121 OUT2.n146 OUT2.n145 52.82
R21122 OUT2.n148 OUT2.n147 52.82
R21123 OUT2.n83 OUT2.n82 52.82
R21124 OUT2.n85 OUT2.n84 52.82
R21125 OUT2.n87 OUT2.n86 52.82
R21126 OUT2.n89 OUT2.n88 52.82
R21127 OUT2.n91 OUT2.n90 52.82
R21128 OUT2.n93 OUT2.n92 52.82
R21129 OUT2.n44 OUT2.n43 52.82
R21130 OUT2.n46 OUT2.n45 52.82
R21131 OUT2.n48 OUT2.n47 52.82
R21132 OUT2.n50 OUT2.n49 52.82
R21133 OUT2.n52 OUT2.n51 52.82
R21134 OUT2.n4 OUT2.n3 52.82
R21135 OUT2.n6 OUT2.n5 52.82
R21136 OUT2.n8 OUT2.n7 52.82
R21137 OUT2.n10 OUT2.n9 52.82
R21138 OUT2.n12 OUT2.n11 52.82
R21139 OUT2 OUT2.n149 51.0745
R21140 OUT2 OUT2.n94 51.0745
R21141 OUT2.n124 OUT2.n122 38.4005
R21142 OUT2.n126 OUT2.n124 38.4005
R21143 OUT2.n128 OUT2.n126 38.4005
R21144 OUT2.n130 OUT2.n128 38.4005
R21145 OUT2.n132 OUT2.n130 38.4005
R21146 OUT2.n133 OUT2.n132 38.4005
R21147 OUT2.n104 OUT2.n102 38.4005
R21148 OUT2.n106 OUT2.n104 38.4005
R21149 OUT2.n108 OUT2.n106 38.4005
R21150 OUT2.n110 OUT2.n108 38.4005
R21151 OUT2.n112 OUT2.n110 38.4005
R21152 OUT2.n113 OUT2.n112 38.4005
R21153 OUT2.n67 OUT2.n65 38.4005
R21154 OUT2.n69 OUT2.n67 38.4005
R21155 OUT2.n71 OUT2.n69 38.4005
R21156 OUT2.n73 OUT2.n71 38.4005
R21157 OUT2.n75 OUT2.n73 38.4005
R21158 OUT2.n76 OUT2.n75 38.4005
R21159 OUT2.n27 OUT2.n25 38.4005
R21160 OUT2.n29 OUT2.n27 38.4005
R21161 OUT2.n31 OUT2.n29 38.4005
R21162 OUT2.n33 OUT2.n31 38.4005
R21163 OUT2.n35 OUT2.n33 38.4005
R21164 OUT2.n36 OUT2.n35 38.4005
R21165 OUT2.n140 OUT2.n138 34.3584
R21166 OUT2.n142 OUT2.n140 34.3584
R21167 OUT2.n144 OUT2.n142 34.3584
R21168 OUT2.n146 OUT2.n144 34.3584
R21169 OUT2.n148 OUT2.n146 34.3584
R21170 OUT2.n150 OUT2.n148 34.3584
R21171 OUT2.n85 OUT2.n83 34.3584
R21172 OUT2.n87 OUT2.n85 34.3584
R21173 OUT2.n89 OUT2.n87 34.3584
R21174 OUT2.n91 OUT2.n89 34.3584
R21175 OUT2.n93 OUT2.n91 34.3584
R21176 OUT2.n95 OUT2.n93 34.3584
R21177 OUT2.n46 OUT2.n44 34.3584
R21178 OUT2.n48 OUT2.n46 34.3584
R21179 OUT2.n50 OUT2.n48 34.3584
R21180 OUT2.n52 OUT2.n50 34.3584
R21181 OUT2.n54 OUT2.n52 34.3584
R21182 OUT2.n58 OUT2.n54 34.3584
R21183 OUT2.n6 OUT2.n4 34.3584
R21184 OUT2.n8 OUT2.n6 34.3584
R21185 OUT2.n10 OUT2.n8 34.3584
R21186 OUT2.n12 OUT2.n10 34.3584
R21187 OUT2.n14 OUT2.n12 34.3584
R21188 OUT2.n18 OUT2.n14 34.3584
R21189 OUT2.n118 OUT2.t52 26.5955
R21190 OUT2.n118 OUT2.t1 26.5955
R21191 OUT2.n120 OUT2.t50 26.5955
R21192 OUT2.n120 OUT2.t22 26.5955
R21193 OUT2.n121 OUT2.t8 26.5955
R21194 OUT2.n121 OUT2.t38 26.5955
R21195 OUT2.n123 OUT2.t17 26.5955
R21196 OUT2.n123 OUT2.t58 26.5955
R21197 OUT2.n125 OUT2.t28 26.5955
R21198 OUT2.n125 OUT2.t46 26.5955
R21199 OUT2.n127 OUT2.t44 26.5955
R21200 OUT2.n127 OUT2.t61 26.5955
R21201 OUT2.n129 OUT2.t3 26.5955
R21202 OUT2.n129 OUT2.t33 26.5955
R21203 OUT2.n131 OUT2.t14 26.5955
R21204 OUT2.n131 OUT2.t54 26.5955
R21205 OUT2.n99 OUT2.t13 26.5955
R21206 OUT2.n99 OUT2.t42 26.5955
R21207 OUT2.n100 OUT2.t32 26.5955
R21208 OUT2.n100 OUT2.t41 26.5955
R21209 OUT2.n101 OUT2.t48 26.5955
R21210 OUT2.n101 OUT2.t21 26.5955
R21211 OUT2.n103 OUT2.t63 26.5955
R21212 OUT2.n103 OUT2.t35 26.5955
R21213 OUT2.n105 OUT2.t34 26.5955
R21214 OUT2.n105 OUT2.t47 26.5955
R21215 OUT2.n107 OUT2.t55 26.5955
R21216 OUT2.n107 OUT2.t5 26.5955
R21217 OUT2.n109 OUT2.t4 26.5955
R21218 OUT2.n109 OUT2.t23 26.5955
R21219 OUT2.n111 OUT2.t57 26.5955
R21220 OUT2.n111 OUT2.t25 26.5955
R21221 OUT2.n62 OUT2.t19 26.5955
R21222 OUT2.n62 OUT2.t53 26.5955
R21223 OUT2.n63 OUT2.t39 26.5955
R21224 OUT2.n63 OUT2.t51 26.5955
R21225 OUT2.n64 OUT2.t49 26.5955
R21226 OUT2.n64 OUT2.t9 26.5955
R21227 OUT2.n66 OUT2.t6 26.5955
R21228 OUT2.n66 OUT2.t36 26.5955
R21229 OUT2.n68 OUT2.t62 26.5955
R21230 OUT2.n68 OUT2.t30 26.5955
R21231 OUT2.n70 OUT2.t27 26.5955
R21232 OUT2.n70 OUT2.t45 26.5955
R21233 OUT2.n72 OUT2.t43 26.5955
R21234 OUT2.n72 OUT2.t60 26.5955
R21235 OUT2.n74 OUT2.t2 26.5955
R21236 OUT2.n74 OUT2.t15 26.5955
R21237 OUT2.n22 OUT2.t18 26.5955
R21238 OUT2.n22 OUT2.t31 26.5955
R21239 OUT2.n23 OUT2.t37 26.5955
R21240 OUT2.n23 OUT2.t59 26.5955
R21241 OUT2.n24 OUT2.t56 26.5955
R21242 OUT2.n24 OUT2.t7 26.5955
R21243 OUT2.n26 OUT2.t12 26.5955
R21244 OUT2.n26 OUT2.t24 26.5955
R21245 OUT2.n28 OUT2.t29 26.5955
R21246 OUT2.n28 OUT2.t0 26.5955
R21247 OUT2.n30 OUT2.t40 26.5955
R21248 OUT2.n30 OUT2.t11 26.5955
R21249 OUT2.n32 OUT2.t16 26.5955
R21250 OUT2.n32 OUT2.t26 26.5955
R21251 OUT2.n34 OUT2.t10 26.5955
R21252 OUT2.n34 OUT2.t20 26.5955
R21253 OUT2.n149 OUT2.t70 24.9236
R21254 OUT2.n149 OUT2.t83 24.9236
R21255 OUT2.n136 OUT2.t68 24.9236
R21256 OUT2.n136 OUT2.t104 24.9236
R21257 OUT2.n137 OUT2.t90 24.9236
R21258 OUT2.n137 OUT2.t120 24.9236
R21259 OUT2.n139 OUT2.t99 24.9236
R21260 OUT2.n139 OUT2.t76 24.9236
R21261 OUT2.n141 OUT2.t110 24.9236
R21262 OUT2.n141 OUT2.t64 24.9236
R21263 OUT2.n143 OUT2.t126 24.9236
R21264 OUT2.n143 OUT2.t79 24.9236
R21265 OUT2.n145 OUT2.t85 24.9236
R21266 OUT2.n145 OUT2.t115 24.9236
R21267 OUT2.n147 OUT2.t96 24.9236
R21268 OUT2.n147 OUT2.t72 24.9236
R21269 OUT2.n94 OUT2.t95 24.9236
R21270 OUT2.n94 OUT2.t124 24.9236
R21271 OUT2.n81 OUT2.t114 24.9236
R21272 OUT2.n81 OUT2.t123 24.9236
R21273 OUT2.n82 OUT2.t66 24.9236
R21274 OUT2.n82 OUT2.t103 24.9236
R21275 OUT2.n84 OUT2.t81 24.9236
R21276 OUT2.n84 OUT2.t117 24.9236
R21277 OUT2.n86 OUT2.t116 24.9236
R21278 OUT2.n86 OUT2.t65 24.9236
R21279 OUT2.n88 OUT2.t73 24.9236
R21280 OUT2.n88 OUT2.t87 24.9236
R21281 OUT2.n90 OUT2.t86 24.9236
R21282 OUT2.n90 OUT2.t105 24.9236
R21283 OUT2.n92 OUT2.t75 24.9236
R21284 OUT2.n92 OUT2.t107 24.9236
R21285 OUT2.n55 OUT2.t101 24.9236
R21286 OUT2.n55 OUT2.t71 24.9236
R21287 OUT2.n42 OUT2.t121 24.9236
R21288 OUT2.n42 OUT2.t69 24.9236
R21289 OUT2.n43 OUT2.t67 24.9236
R21290 OUT2.n43 OUT2.t91 24.9236
R21291 OUT2.n45 OUT2.t88 24.9236
R21292 OUT2.n45 OUT2.t118 24.9236
R21293 OUT2.n47 OUT2.t80 24.9236
R21294 OUT2.n47 OUT2.t112 24.9236
R21295 OUT2.n49 OUT2.t108 24.9236
R21296 OUT2.n49 OUT2.t127 24.9236
R21297 OUT2.n51 OUT2.t125 24.9236
R21298 OUT2.n51 OUT2.t78 24.9236
R21299 OUT2.n53 OUT2.t84 24.9236
R21300 OUT2.n53 OUT2.t97 24.9236
R21301 OUT2.n15 OUT2.t100 24.9236
R21302 OUT2.n15 OUT2.t113 24.9236
R21303 OUT2.n2 OUT2.t119 24.9236
R21304 OUT2.n2 OUT2.t77 24.9236
R21305 OUT2.n3 OUT2.t74 24.9236
R21306 OUT2.n3 OUT2.t89 24.9236
R21307 OUT2.n5 OUT2.t94 24.9236
R21308 OUT2.n5 OUT2.t106 24.9236
R21309 OUT2.n7 OUT2.t111 24.9236
R21310 OUT2.n7 OUT2.t82 24.9236
R21311 OUT2.n9 OUT2.t122 24.9236
R21312 OUT2.n9 OUT2.t93 24.9236
R21313 OUT2.n11 OUT2.t98 24.9236
R21314 OUT2.n11 OUT2.t109 24.9236
R21315 OUT2.n13 OUT2.t92 24.9236
R21316 OUT2.n13 OUT2.t102 24.9236
R21317 OUT2 OUT2.n150 11.4429
R21318 OUT2 OUT2.n95 11.4429
R21319 OUT2 OUT2.n58 11.4429
R21320 OUT2 OUT2.n18 11.4429
R21321 OUT2.n77 OUT2.n62 8.55118
R21322 OUT2.n37 OUT2.n22 8.55118
R21323 OUT2.n114 OUT2.n99 8.55117
R21324 OUT2.n119 OUT2.n118 8.47293
R21325 OUT2.n56 OUT2.n55 7.80093
R21326 OUT2.n16 OUT2.n15 7.80093
R21327 OUT2.n78 OUT2.n77 3.20954
R21328 OUT2.n38 OUT2.n37 3.20953
R21329 OUT2.n115 OUT2.n114 3.20289
R21330 OUT2.n151 OUT2 3.10353
R21331 OUT2.n96 OUT2 3.10353
R21332 OUT2.n59 OUT2 3.10353
R21333 OUT2.n19 OUT2 3.10353
R21334 OUT2.n135 OUT2.n134 3.1005
R21335 OUT2.n57 OUT2.n41 3.1005
R21336 OUT2.n17 OUT2.n1 3.1005
R21337 OUT2.n134 OUT2.n133 2.71565
R21338 OUT2.n114 OUT2.n113 2.13383
R21339 OUT2.n77 OUT2.n76 2.13383
R21340 OUT2.n37 OUT2.n36 2.13383
R21341 OUT2.n150 OUT2 1.74595
R21342 OUT2.n95 OUT2 1.74595
R21343 OUT2.n58 OUT2.n57 1.16414
R21344 OUT2.n18 OUT2.n17 1.16414
R21345 OUT2.n157 OUT2.n156 1.07337
R21346 OUT2.n158 OUT2.n157 0.69375
R21347 OUT2.n159 OUT2.n158 0.68905
R21348 OUT2.n56 OUT2 0.488972
R21349 OUT2.n16 OUT2 0.488972
R21350 OUT2.n158 OUT2.n79 0.414635
R21351 OUT2.n157 OUT2.n116 0.382465
R21352 OUT2.n159 OUT2.n39 0.368576
R21353 OUT2 OUT2.n159 0.281623
R21354 OUT2.n134 OUT2.n119 0.196887
R21355 OUT2.n79 OUT2.n78 0.157252
R21356 OUT2.n39 OUT2.n38 0.139891
R21357 OUT2.n156 OUT2.n155 0.139389
R21358 OUT2.n116 OUT2.n115 0.132946
R21359 OUT2.n60 OUT2.n41 0.113
R21360 OUT2.n20 OUT2.n1 0.113
R21361 OUT2.n154 OUT2.n135 0.101889
R21362 OUT2.n57 OUT2.n56 0.0893205
R21363 OUT2.n17 OUT2.n16 0.0893205
R21364 OUT2.n154 OUT2.n152 0.0282778
R21365 OUT2.n135 OUT2.n117 0.0268889
R21366 OUT2.n98 OUT2.n97 0.0213333
R21367 OUT2.n61 OUT2.n60 0.0143889
R21368 OUT2.n21 OUT2.n20 0.0143889
R21369 OUT2.n115 OUT2.n98 0.00100004
R21370 OUT2.n38 OUT2.n21 0.00100004
R21371 OUT2.n78 OUT2.n61 0.00100004
R21372 OUT2.n152 OUT2.n151 0.000513335
R21373 OUT2.n97 OUT2.n96 0.000513335
R21374 OUT2.n60 OUT2.n59 0.000513218
R21375 OUT2.n20 OUT2.n19 0.000513218
R21376 OUT2.n98 OUT2.n80 0.00050517
R21377 OUT2.n154 OUT2.n153 0.000504838
R21378 OUT2.n61 OUT2.n40 0.000504838
R21379 OUT2.n21 OUT2.n0 0.000504838
R21380 OUT2.n155 OUT2.n154 0.000501713
R21381 VFS.n3 VFS 0.239679
R21382 VFS.n4 VFS.t2 0.0274553
R21383 VFS.n0 VFS.t7 0.0274553
R21384 VFS.n1 VFS.n0 0.0274531
R21385 VFS.n2 VFS.n1 0.0274531
R21386 VFS.n6 VFS.n5 0.0274531
R21387 VFS.n5 VFS.n4 0.0274531
R21388 VFS VFS.n6 0.014671
R21389 VFS.n3 VFS.n2 0.011546
R21390 VFS VFS.n3 0.00223611
R21391 VFS.n4 VFS.t4 0.000502142
R21392 VFS.n5 VFS.t0 0.000502142
R21393 VFS.n6 VFS.t5 0.000502142
R21394 VFS.n2 VFS.t3 0.000502142
R21395 VFS.n1 VFS.t1 0.000502142
R21396 VFS.n0 VFS.t6 0.000502142
R21397 resistorDivider_v0p0p1_0.V16.n0 resistorDivider_v0p0p1_0.V16.t17 167.365
R21398 resistorDivider_v0p0p1_0.V16.n0 resistorDivider_v0p0p1_0.V16.t16 92.4496
R21399 resistorDivider_v0p0p1_0.V16.n1 resistorDivider_v0p0p1_0.V16.n0 2.07493
R21400 resistorDivider_v0p0p1_0.V16.n15 resistorDivider_v0p0p1_0.V16.n14 0.141409
R21401 resistorDivider_v0p0p1_0.V16.n13 resistorDivider_v0p0p1_0.V16.n12 0.141409
R21402 resistorDivider_v0p0p1_0.V16.n11 resistorDivider_v0p0p1_0.V16.n10 0.141409
R21403 resistorDivider_v0p0p1_0.V16.n9 resistorDivider_v0p0p1_0.V16.n8 0.141409
R21404 resistorDivider_v0p0p1_0.V16.n7 resistorDivider_v0p0p1_0.V16.n6 0.141409
R21405 resistorDivider_v0p0p1_0.V16.n5 resistorDivider_v0p0p1_0.V16.n4 0.141409
R21406 resistorDivider_v0p0p1_0.V16.n3 resistorDivider_v0p0p1_0.V16.n2 0.141409
R21407 resistorDivider_v0p0p1_0.V16.n1 resistorDivider_v0p0p1_0.V16 0.12425
R21408 resistorDivider_v0p0p1_0.V16 resistorDivider_v0p0p1_0.V16.n16 0.105614
R21409 resistorDivider_v0p0p1_0.V16 resistorDivider_v0p0p1_0.V16.n1 0.05
R21410 resistorDivider_v0p0p1_0.V16.n5 resistorDivider_v0p0p1_0.V16.t0 0.00250214
R21411 resistorDivider_v0p0p1_0.V16.n2 resistorDivider_v0p0p1_0.V16.t7 0.000729415
R21412 resistorDivider_v0p0p1_0.V16.n16 resistorDivider_v0p0p1_0.V16.n15 0.000727273
R21413 resistorDivider_v0p0p1_0.V16.n14 resistorDivider_v0p0p1_0.V16.n13 0.000727273
R21414 resistorDivider_v0p0p1_0.V16.n12 resistorDivider_v0p0p1_0.V16.n11 0.000727273
R21415 resistorDivider_v0p0p1_0.V16.n10 resistorDivider_v0p0p1_0.V16.n9 0.000727273
R21416 resistorDivider_v0p0p1_0.V16.n8 resistorDivider_v0p0p1_0.V16.n7 0.000727273
R21417 resistorDivider_v0p0p1_0.V16.n6 resistorDivider_v0p0p1_0.V16.n5 0.000727273
R21418 resistorDivider_v0p0p1_0.V16.n4 resistorDivider_v0p0p1_0.V16.n3 0.000727273
R21419 resistorDivider_v0p0p1_0.V16.n3 resistorDivider_v0p0p1_0.V16.t11 0.000502142
R21420 resistorDivider_v0p0p1_0.V16.n7 resistorDivider_v0p0p1_0.V16.t3 0.000502142
R21421 resistorDivider_v0p0p1_0.V16.n9 resistorDivider_v0p0p1_0.V16.t15 0.000502142
R21422 resistorDivider_v0p0p1_0.V16.n11 resistorDivider_v0p0p1_0.V16.t14 0.000502142
R21423 resistorDivider_v0p0p1_0.V16.n13 resistorDivider_v0p0p1_0.V16.t12 0.000502142
R21424 resistorDivider_v0p0p1_0.V16.n15 resistorDivider_v0p0p1_0.V16.t1 0.000502142
R21425 resistorDivider_v0p0p1_0.V16.n16 resistorDivider_v0p0p1_0.V16.t13 0.000502142
R21426 resistorDivider_v0p0p1_0.V16.n14 resistorDivider_v0p0p1_0.V16.t10 0.000502142
R21427 resistorDivider_v0p0p1_0.V16.n12 resistorDivider_v0p0p1_0.V16.t4 0.000502142
R21428 resistorDivider_v0p0p1_0.V16.n10 resistorDivider_v0p0p1_0.V16.t6 0.000502142
R21429 resistorDivider_v0p0p1_0.V16.n8 resistorDivider_v0p0p1_0.V16.t9 0.000502142
R21430 resistorDivider_v0p0p1_0.V16.n6 resistorDivider_v0p0p1_0.V16.t2 0.000502142
R21431 resistorDivider_v0p0p1_0.V16.n4 resistorDivider_v0p0p1_0.V16.t8 0.000502142
R21432 resistorDivider_v0p0p1_0.V16.n2 resistorDivider_v0p0p1_0.V16.t5 0.000502142
R21433 a_16599_n13205.n12 a_16599_n13205.t21 182.77
R21434 a_16599_n13205.n13 a_16599_n13205.t14 182.77
R21435 a_16599_n13205.n14 a_16599_n13205.t6 182.77
R21436 a_16599_n13205.n15 a_16599_n13205.t10 182.77
R21437 a_16599_n13205.n16 a_16599_n13205.t18 182.77
R21438 a_16599_n13205.n17 a_16599_n13205.t4 182.77
R21439 a_16599_n13205.n18 a_16599_n13205.t19 182.77
R21440 a_16599_n13205.n19 a_16599_n13205.t9 182.77
R21441 a_16599_n13205.n20 a_16599_n13205.t5 182.77
R21442 a_16599_n13205.n21 a_16599_n13205.t0 182.77
R21443 a_16599_n13205.n2 a_16599_n13205.t8 182.77
R21444 a_16599_n13205.n3 a_16599_n13205.t23 182.77
R21445 a_16599_n13205.n4 a_16599_n13205.t12 182.77
R21446 a_16599_n13205.n5 a_16599_n13205.t20 182.77
R21447 a_16599_n13205.n6 a_16599_n13205.t13 182.77
R21448 a_16599_n13205.n7 a_16599_n13205.t7 182.77
R21449 a_16599_n13205.n8 a_16599_n13205.t22 182.77
R21450 a_16599_n13205.n9 a_16599_n13205.t11 182.77
R21451 a_16599_n13205.n10 a_16599_n13205.t16 182.77
R21452 a_16599_n13205.n11 a_16599_n13205.t17 90.7933
R21453 a_16599_n13205.n1 a_16599_n13205.t15 90.7875
R21454 a_16599_n13205.n43 a_16599_n13205.t2 42.4202
R21455 a_16599_n13205.n0 a_16599_n13205.t1 4.35105
R21456 a_16599_n13205.t3 a_16599_n13205.n43 2.70045
R21457 a_16599_n13205.n2 a_16599_n13205.n1 2.03273
R21458 a_16599_n13205.n12 a_16599_n13205.n11 2.02124
R21459 a_16599_n13205.n41 a_16599_n13205.n40 0.835222
R21460 a_16599_n13205.n40 a_16599_n13205.n39 0.835222
R21461 a_16599_n13205.n39 a_16599_n13205.n38 0.835222
R21462 a_16599_n13205.n38 a_16599_n13205.n37 0.835222
R21463 a_16599_n13205.n37 a_16599_n13205.n36 0.835222
R21464 a_16599_n13205.n36 a_16599_n13205.n35 0.835222
R21465 a_16599_n13205.n35 a_16599_n13205.n34 0.835222
R21466 a_16599_n13205.n34 a_16599_n13205.n33 0.835222
R21467 a_16599_n13205.n33 a_16599_n13205.n32 0.835222
R21468 a_16599_n13205.n13 a_16599_n13205.n12 0.835222
R21469 a_16599_n13205.n14 a_16599_n13205.n13 0.835222
R21470 a_16599_n13205.n15 a_16599_n13205.n14 0.835222
R21471 a_16599_n13205.n16 a_16599_n13205.n15 0.835222
R21472 a_16599_n13205.n17 a_16599_n13205.n16 0.835222
R21473 a_16599_n13205.n18 a_16599_n13205.n17 0.835222
R21474 a_16599_n13205.n19 a_16599_n13205.n18 0.835222
R21475 a_16599_n13205.n20 a_16599_n13205.n19 0.835222
R21476 a_16599_n13205.n21 a_16599_n13205.n20 0.835222
R21477 a_16599_n13205.n10 a_16599_n13205.n9 0.835222
R21478 a_16599_n13205.n9 a_16599_n13205.n8 0.835222
R21479 a_16599_n13205.n8 a_16599_n13205.n7 0.835222
R21480 a_16599_n13205.n7 a_16599_n13205.n6 0.835222
R21481 a_16599_n13205.n6 a_16599_n13205.n5 0.835222
R21482 a_16599_n13205.n5 a_16599_n13205.n4 0.835222
R21483 a_16599_n13205.n4 a_16599_n13205.n3 0.835222
R21484 a_16599_n13205.n3 a_16599_n13205.n2 0.835222
R21485 a_16599_n13205.n24 a_16599_n13205.n23 0.835222
R21486 a_16599_n13205.n25 a_16599_n13205.n24 0.835222
R21487 a_16599_n13205.n26 a_16599_n13205.n25 0.835222
R21488 a_16599_n13205.n27 a_16599_n13205.n26 0.835222
R21489 a_16599_n13205.n28 a_16599_n13205.n27 0.835222
R21490 a_16599_n13205.n29 a_16599_n13205.n28 0.835222
R21491 a_16599_n13205.n30 a_16599_n13205.n29 0.835222
R21492 a_16599_n13205.n31 a_16599_n13205.n30 0.835222
R21493 a_16599_n13205.n0 a_16599_n13205.n42 0.750184
R21494 a_16599_n13205.n0 a_16599_n13205.n22 0.715064
R21495 a_16599_n13205.n22 a_16599_n13205.n10 0.553972
R21496 a_16599_n13205.n42 a_16599_n13205.n31 0.553972
R21497 a_16599_n13205.n43 a_16599_n13205.n0 0.403234
R21498 a_16599_n13205.n42 a_16599_n13205.n41 0.233139
R21499 a_16599_n13205.n22 a_16599_n13205.n21 0.233139
R21500 a_16541_n13117.n0 a_16541_n13117.t13 5.73525
R21501 a_16541_n13117.n18 a_16541_n13117.t11 5.34571
R21502 a_16541_n13117.n0 a_16541_n13117.t4 5.18362
R21503 a_16541_n13117.n1 a_16541_n13117.t19 5.18362
R21504 a_16541_n13117.n2 a_16541_n13117.t0 5.18362
R21505 a_16541_n13117.n3 a_16541_n13117.t8 5.18362
R21506 a_16541_n13117.n4 a_16541_n13117.t15 5.18362
R21507 a_16541_n13117.n5 a_16541_n13117.t5 5.18362
R21508 a_16541_n13117.n6 a_16541_n13117.t6 5.18362
R21509 a_16541_n13117.n7 a_16541_n13117.t1 5.18362
R21510 a_16541_n13117.n8 a_16541_n13117.t12 5.18362
R21511 a_16541_n13117.n9 a_16541_n13117.t17 5.18362
R21512 a_16541_n13117.n10 a_16541_n13117.t3 5.18362
R21513 a_16541_n13117.n11 a_16541_n13117.t9 5.18362
R21514 a_16541_n13117.n12 a_16541_n13117.t18 5.18362
R21515 a_16541_n13117.n13 a_16541_n13117.t10 5.18362
R21516 a_16541_n13117.n14 a_16541_n13117.t2 5.18362
R21517 a_16541_n13117.n15 a_16541_n13117.t16 5.18362
R21518 a_16541_n13117.n16 a_16541_n13117.t14 5.18362
R21519 a_16541_n13117.n17 a_16541_n13117.t7 5.18362
R21520 a_16541_n13117.t20 a_16541_n13117.n19 2.79552
R21521 a_16541_n13117.n19 a_16541_n13117.t21 2.38201
R21522 a_16541_n13117.n9 a_16541_n13117.n8 1.10376
R21523 a_16541_n13117.n1 a_16541_n13117.n0 0.55213
R21524 a_16541_n13117.n2 a_16541_n13117.n1 0.55213
R21525 a_16541_n13117.n3 a_16541_n13117.n2 0.55213
R21526 a_16541_n13117.n4 a_16541_n13117.n3 0.55213
R21527 a_16541_n13117.n5 a_16541_n13117.n4 0.55213
R21528 a_16541_n13117.n6 a_16541_n13117.n5 0.55213
R21529 a_16541_n13117.n7 a_16541_n13117.n6 0.55213
R21530 a_16541_n13117.n8 a_16541_n13117.n7 0.55213
R21531 a_16541_n13117.n10 a_16541_n13117.n9 0.55213
R21532 a_16541_n13117.n11 a_16541_n13117.n10 0.55213
R21533 a_16541_n13117.n12 a_16541_n13117.n11 0.55213
R21534 a_16541_n13117.n13 a_16541_n13117.n12 0.55213
R21535 a_16541_n13117.n14 a_16541_n13117.n13 0.55213
R21536 a_16541_n13117.n15 a_16541_n13117.n14 0.55213
R21537 a_16541_n13117.n16 a_16541_n13117.n15 0.55213
R21538 a_16541_n13117.n17 a_16541_n13117.n16 0.512683
R21539 a_16541_n13117.n19 a_16541_n13117.n18 0.168655
R21540 a_16541_n13117.n18 a_16541_n13117.n17 0.0581389
R21541 a_16719_n13117.n15 a_16719_n13117.t24 473.437
R21542 a_16719_n13117.n19 a_16719_n13117.t25 473.332
R21543 a_16719_n13117.n0 a_16719_n13117.t22 473.329
R21544 a_16719_n13117.n18 a_16719_n13117.t20 140.444
R21545 a_16719_n13117.n18 a_16719_n13117.t21 41.6504
R21546 a_16719_n13117.n2 a_16719_n13117.t8 5.95597
R21547 a_16719_n13117.n26 a_16719_n13117.t6 5.95597
R21548 a_16719_n13117.n8 a_16719_n13117.t1 5.32159
R21549 a_16719_n13117.n7 a_16719_n13117.t16 5.32159
R21550 a_16719_n13117.n6 a_16719_n13117.t10 5.32159
R21551 a_16719_n13117.n5 a_16719_n13117.t3 5.32159
R21552 a_16719_n13117.n4 a_16719_n13117.t11 5.32159
R21553 a_16719_n13117.n3 a_16719_n13117.t0 5.32159
R21554 a_16719_n13117.n2 a_16719_n13117.t15 5.32159
R21555 a_16719_n13117.n1 a_16719_n13117.t7 5.32159
R21556 a_16719_n13117.n11 a_16719_n13117.t12 5.32159
R21557 a_16719_n13117.n26 a_16719_n13117.t2 5.32159
R21558 a_16719_n13117.n27 a_16719_n13117.t9 5.32159
R21559 a_16719_n13117.n28 a_16719_n13117.t17 5.32159
R21560 a_16719_n13117.n29 a_16719_n13117.t13 5.32159
R21561 a_16719_n13117.n30 a_16719_n13117.t5 5.32159
R21562 a_16719_n13117.n25 a_16719_n13117.t4 5.32159
R21563 a_16719_n13117.n24 a_16719_n13117.t14 5.32159
R21564 a_16719_n13117.n23 a_16719_n13117.t18 5.32159
R21565 a_16719_n13117.t19 a_16719_n13117.n31 5.32059
R21566 a_16719_n13117.n14 a_16719_n13117.n13 2.75606
R21567 a_16719_n13117.n17 a_16719_n13117.n14 2.75328
R21568 a_16719_n13117.n14 a_16719_n13117.t23 1.50409
R21569 a_16719_n13117.n19 a_16719_n13117.n18 1.23545
R21570 a_16719_n13117.n23 a_16719_n13117.n22 1.02772
R21571 a_16719_n13117.n3 a_16719_n13117.n2 0.634875
R21572 a_16719_n13117.n4 a_16719_n13117.n3 0.634875
R21573 a_16719_n13117.n5 a_16719_n13117.n4 0.634875
R21574 a_16719_n13117.n6 a_16719_n13117.n5 0.634875
R21575 a_16719_n13117.n7 a_16719_n13117.n6 0.634875
R21576 a_16719_n13117.n8 a_16719_n13117.n7 0.634875
R21577 a_16719_n13117.n24 a_16719_n13117.n23 0.634875
R21578 a_16719_n13117.n25 a_16719_n13117.n24 0.634875
R21579 a_16719_n13117.n31 a_16719_n13117.n25 0.634875
R21580 a_16719_n13117.n31 a_16719_n13117.n30 0.634875
R21581 a_16719_n13117.n30 a_16719_n13117.n29 0.634875
R21582 a_16719_n13117.n29 a_16719_n13117.n28 0.634875
R21583 a_16719_n13117.n28 a_16719_n13117.n27 0.634875
R21584 a_16719_n13117.n27 a_16719_n13117.n26 0.634875
R21585 a_16719_n13117.n0 a_16719_n13117.n21 0.376529
R21586 a_16719_n13117.n16 a_16719_n13117.n15 0.271346
R21587 a_16719_n13117.n21 a_16719_n13117.n20 0.253053
R21588 a_16719_n13117.n9 a_16719_n13117.n8 0.202227
R21589 a_16719_n13117.n20 a_16719_n13117.n19 0.124538
R21590 a_16719_n13117.n17 a_16719_n13117.n16 0.119076
R21591 a_16719_n13117.n13 a_16719_n13117.n12 0.113872
R21592 a_16719_n13117.n0 a_16719_n13117.n17 0.10111
R21593 a_16719_n13117.n1 a_16719_n13117.n0 0.0537895
R21594 a_16719_n13117.n10 a_16719_n13117.n9 0.0386579
R21595 a_16719_n13117.n22 a_16719_n13117.n1 0.0360263
R21596 a_16719_n13117.n0 a_16719_n13117.n11 0.035794
R21597 a_16719_n13117.n11 a_16719_n13117.n10 0.0202368
R21598 CLK.t85 CLK.t89 344.122
R21599 CLK.t72 CLK.t34 344.122
R21600 CLK.t60 CLK.t16 344.122
R21601 CLK.t7 CLK.t57 344.122
R21602 CLK.t87 CLK.t36 344.122
R21603 CLK.t28 CLK.t80 344.122
R21604 CLK.t13 CLK.t70 344.122
R21605 CLK.t51 CLK.t6 344.122
R21606 CLK.t39 CLK.t95 344.122
R21607 CLK.t74 CLK.t71 344.122
R21608 CLK.t64 CLK.t18 344.122
R21609 CLK.t47 CLK.t5 344.122
R21610 CLK.t90 CLK.t38 344.122
R21611 CLK.t73 CLK.t27 344.122
R21612 CLK.t14 CLK.t63 344.122
R21613 CLK.t48 CLK.t46 344.122
R21614 CLK.n1 CLK.t50 232.299
R21615 CLK.n114 CLK.t42 232.299
R21616 CLK.n106 CLK.t84 232.299
R21617 CLK.n98 CLK.t67 232.299
R21618 CLK.n90 CLK.t52 232.299
R21619 CLK.n82 CLK.t1 232.299
R21620 CLK.n74 CLK.t75 232.299
R21621 CLK.n66 CLK.t21 232.299
R21622 CLK.n58 CLK.t3 232.299
R21623 CLK.n50 CLK.t43 232.299
R21624 CLK.n42 CLK.t31 232.299
R21625 CLK.n34 CLK.t68 232.299
R21626 CLK.n26 CLK.t55 232.299
R21627 CLK.n18 CLK.t93 232.299
R21628 CLK.n10 CLK.t77 232.299
R21629 CLK.n137 CLK.t22 232.299
R21630 CLK.n5 CLK.t94 182.915
R21631 CLK.n118 CLK.t81 182.915
R21632 CLK.n110 CLK.t61 182.915
R21633 CLK.n102 CLK.t8 182.915
R21634 CLK.n94 CLK.t88 182.915
R21635 CLK.n86 CLK.t29 182.915
R21636 CLK.n78 CLK.t19 182.915
R21637 CLK.n70 CLK.t53 182.915
R21638 CLK.n62 CLK.t40 182.915
R21639 CLK.n54 CLK.t76 182.915
R21640 CLK.n46 CLK.t65 182.915
R21641 CLK.n38 CLK.t10 182.915
R21642 CLK.n30 CLK.t91 182.915
R21643 CLK.n22 CLK.t32 182.915
R21644 CLK.n14 CLK.t15 182.915
R21645 CLK.n140 CLK.t49 182.915
R21646 CLK.n5 CLK.t85 182.91
R21647 CLK.n118 CLK.t72 182.91
R21648 CLK.n110 CLK.t60 182.91
R21649 CLK.n102 CLK.t7 182.91
R21650 CLK.n94 CLK.t87 182.91
R21651 CLK.n86 CLK.t28 182.91
R21652 CLK.n78 CLK.t13 182.91
R21653 CLK.n70 CLK.t51 182.91
R21654 CLK.n62 CLK.t39 182.91
R21655 CLK.n54 CLK.t74 182.91
R21656 CLK.n46 CLK.t64 182.91
R21657 CLK.n38 CLK.t47 182.91
R21658 CLK.n30 CLK.t90 182.91
R21659 CLK.n22 CLK.t73 182.91
R21660 CLK.n14 CLK.t14 182.91
R21661 CLK.n140 CLK.t48 182.91
R21662 CLK.t94 CLK.n4 182.769
R21663 CLK.t81 CLK.n117 182.769
R21664 CLK.t61 CLK.n109 182.769
R21665 CLK.t8 CLK.n101 182.769
R21666 CLK.t88 CLK.n93 182.769
R21667 CLK.t29 CLK.n85 182.769
R21668 CLK.t19 CLK.n77 182.769
R21669 CLK.t53 CLK.n69 182.769
R21670 CLK.t40 CLK.n61 182.769
R21671 CLK.t76 CLK.n53 182.769
R21672 CLK.t65 CLK.n45 182.769
R21673 CLK.t10 CLK.n37 182.769
R21674 CLK.t91 CLK.n29 182.769
R21675 CLK.t32 CLK.n21 182.769
R21676 CLK.t15 CLK.n13 182.769
R21677 CLK.t49 CLK.n139 182.769
R21678 CLK.n2 CLK.t26 161.262
R21679 CLK.n115 CLK.t59 161.262
R21680 CLK.n107 CLK.t37 161.262
R21681 CLK.n99 CLK.t82 161.262
R21682 CLK.n91 CLK.t62 161.262
R21683 CLK.n83 CLK.t9 161.262
R21684 CLK.n75 CLK.t0 161.262
R21685 CLK.n67 CLK.t30 161.262
R21686 CLK.n59 CLK.t20 161.262
R21687 CLK.n51 CLK.t54 161.262
R21688 CLK.n43 CLK.t41 161.262
R21689 CLK.n35 CLK.t83 161.262
R21690 CLK.n27 CLK.t66 161.262
R21691 CLK.n19 CLK.t11 161.262
R21692 CLK.n11 CLK.t92 161.262
R21693 CLK.n135 CLK.t86 161.262
R21694 CLK.n6 CLK.t23 159.958
R21695 CLK.n119 CLK.t24 159.958
R21696 CLK.n111 CLK.t12 159.958
R21697 CLK.n103 CLK.t44 159.958
R21698 CLK.n95 CLK.t33 159.958
R21699 CLK.n87 CLK.t69 159.958
R21700 CLK.n79 CLK.t56 159.958
R21701 CLK.n71 CLK.t2 159.958
R21702 CLK.n63 CLK.t79 159.958
R21703 CLK.n55 CLK.t25 159.958
R21704 CLK.n47 CLK.t4 159.958
R21705 CLK.n39 CLK.t45 159.958
R21706 CLK.n31 CLK.t35 159.958
R21707 CLK.n23 CLK.t17 159.958
R21708 CLK.n15 CLK.t58 159.958
R21709 CLK.n141 CLK.t78 159.958
R21710 CLK.n121 CLK 4.70942
R21711 CLK.n3 CLK.n2 4.5005
R21712 CLK.n116 CLK.n115 4.5005
R21713 CLK.n108 CLK.n107 4.5005
R21714 CLK.n100 CLK.n99 4.5005
R21715 CLK.n92 CLK.n91 4.5005
R21716 CLK.n84 CLK.n83 4.5005
R21717 CLK.n76 CLK.n75 4.5005
R21718 CLK.n68 CLK.n67 4.5005
R21719 CLK.n60 CLK.n59 4.5005
R21720 CLK.n52 CLK.n51 4.5005
R21721 CLK.n44 CLK.n43 4.5005
R21722 CLK.n36 CLK.n35 4.5005
R21723 CLK.n28 CLK.n27 4.5005
R21724 CLK.n20 CLK.n19 4.5005
R21725 CLK.n12 CLK.n11 4.5005
R21726 CLK.n122 CLK 4.19834
R21727 CLK.n124 CLK 4.19834
R21728 CLK.n127 CLK 4.19834
R21729 CLK.n123 CLK 4.18793
R21730 CLK.n126 CLK 4.18793
R21731 CLK.n125 CLK 4.17751
R21732 CLK.n132 CLK 4.17751
R21733 CLK.n128 CLK 4.16709
R21734 CLK.n129 CLK 4.16709
R21735 CLK.n131 CLK 4.16709
R21736 CLK.n133 CLK 4.16709
R21737 CLK CLK.n134 4.16709
R21738 CLK.n8 CLK 4.15668
R21739 CLK.n121 CLK 4.14654
R21740 CLK.n130 CLK 4.12571
R21741 CLK.n8 CLK 0.757091
R21742 CLK.n128 CLK.n127 0.620955
R21743 CLK.n125 CLK.n124 0.618682
R21744 CLK.n134 CLK.n8 0.616409
R21745 CLK.n133 CLK.n132 0.616409
R21746 CLK.n130 CLK.n129 0.616409
R21747 CLK.n123 CLK.n122 0.616409
R21748 CLK.n134 CLK.n133 0.614136
R21749 CLK.n129 CLK.n128 0.614136
R21750 CLK.n132 CLK.n131 0.611864
R21751 CLK.n131 CLK.n130 0.611864
R21752 CLK.n127 CLK.n126 0.611864
R21753 CLK.n126 CLK.n125 0.611864
R21754 CLK.n124 CLK.n123 0.611864
R21755 CLK.n122 CLK.n121 0.609591
R21756 CLK.n6 CLK.n5 0.56781
R21757 CLK.n119 CLK.n118 0.56781
R21758 CLK.n111 CLK.n110 0.56781
R21759 CLK.n103 CLK.n102 0.56781
R21760 CLK.n95 CLK.n94 0.56781
R21761 CLK.n87 CLK.n86 0.56781
R21762 CLK.n79 CLK.n78 0.56781
R21763 CLK.n71 CLK.n70 0.56781
R21764 CLK.n63 CLK.n62 0.56781
R21765 CLK.n55 CLK.n54 0.56781
R21766 CLK.n47 CLK.n46 0.56781
R21767 CLK.n39 CLK.n38 0.56781
R21768 CLK.n31 CLK.n30 0.56781
R21769 CLK.n23 CLK.n22 0.56781
R21770 CLK.n15 CLK.n14 0.56781
R21771 CLK.n141 CLK.n140 0.56781
R21772 CLK.n7 CLK.n6 0.428385
R21773 CLK.n120 CLK.n119 0.428385
R21774 CLK.n112 CLK.n111 0.428385
R21775 CLK.n104 CLK.n103 0.428385
R21776 CLK.n96 CLK.n95 0.428385
R21777 CLK.n88 CLK.n87 0.428385
R21778 CLK.n80 CLK.n79 0.428385
R21779 CLK.n72 CLK.n71 0.428385
R21780 CLK.n64 CLK.n63 0.428385
R21781 CLK.n56 CLK.n55 0.428385
R21782 CLK.n48 CLK.n47 0.428385
R21783 CLK.n40 CLK.n39 0.428385
R21784 CLK.n32 CLK.n31 0.428385
R21785 CLK.n24 CLK.n23 0.428385
R21786 CLK.n16 CLK.n15 0.428385
R21787 CLK.n142 CLK.n141 0.428385
R21788 CLK.n7 CLK 0.0573182
R21789 CLK.n104 CLK 0.0573182
R21790 CLK.n96 CLK 0.0573182
R21791 CLK.n88 CLK 0.0573182
R21792 CLK.n80 CLK 0.0573182
R21793 CLK.n72 CLK 0.0573182
R21794 CLK.n64 CLK 0.0573182
R21795 CLK.n56 CLK 0.0573182
R21796 CLK.n48 CLK 0.0573182
R21797 CLK.n32 CLK 0.0573182
R21798 CLK.n24 CLK 0.0573182
R21799 CLK.n16 CLK 0.0573182
R21800 CLK.n142 CLK 0.0573182
R21801 CLK.n120 CLK 0.0525833
R21802 CLK.n112 CLK 0.0525833
R21803 CLK.n40 CLK 0.0525833
R21804 CLK CLK.n7 0.0436818
R21805 CLK CLK.n104 0.0436818
R21806 CLK CLK.n96 0.0436818
R21807 CLK CLK.n88 0.0436818
R21808 CLK CLK.n80 0.0436818
R21809 CLK CLK.n72 0.0436818
R21810 CLK CLK.n64 0.0436818
R21811 CLK CLK.n56 0.0436818
R21812 CLK CLK.n48 0.0436818
R21813 CLK CLK.n32 0.0436818
R21814 CLK CLK.n24 0.0436818
R21815 CLK CLK.n16 0.0436818
R21816 CLK CLK.n142 0.0436818
R21817 CLK CLK.n120 0.0400833
R21818 CLK CLK.n112 0.0400833
R21819 CLK CLK.n40 0.0400833
R21820 CLK.n1 CLK.n0 0.0211923
R21821 CLK.n114 CLK.n113 0.0211923
R21822 CLK.n106 CLK.n105 0.0211923
R21823 CLK.n98 CLK.n97 0.0211923
R21824 CLK.n90 CLK.n89 0.0211923
R21825 CLK.n82 CLK.n81 0.0211923
R21826 CLK.n74 CLK.n73 0.0211923
R21827 CLK.n66 CLK.n65 0.0211923
R21828 CLK.n58 CLK.n57 0.0211923
R21829 CLK.n50 CLK.n49 0.0211923
R21830 CLK.n42 CLK.n41 0.0211923
R21831 CLK.n34 CLK.n33 0.0211923
R21832 CLK.n26 CLK.n25 0.0211923
R21833 CLK.n18 CLK.n17 0.0211923
R21834 CLK.n10 CLK.n9 0.0211923
R21835 CLK.n2 CLK.n0 0.0178077
R21836 CLK.n115 CLK.n113 0.0178077
R21837 CLK.n107 CLK.n105 0.0178077
R21838 CLK.n99 CLK.n97 0.0178077
R21839 CLK.n91 CLK.n89 0.0178077
R21840 CLK.n83 CLK.n81 0.0178077
R21841 CLK.n75 CLK.n73 0.0178077
R21842 CLK.n67 CLK.n65 0.0178077
R21843 CLK.n59 CLK.n57 0.0178077
R21844 CLK.n51 CLK.n49 0.0178077
R21845 CLK.n43 CLK.n41 0.0178077
R21846 CLK.n35 CLK.n33 0.0178077
R21847 CLK.n27 CLK.n25 0.0178077
R21848 CLK.n19 CLK.n17 0.0178077
R21849 CLK.n11 CLK.n9 0.0178077
R21850 CLK.n136 CLK.n135 0.0178077
R21851 CLK.n4 CLK.n0 0.00531334
R21852 CLK.n117 CLK.n113 0.00531334
R21853 CLK.n109 CLK.n105 0.00531334
R21854 CLK.n101 CLK.n97 0.00531334
R21855 CLK.n93 CLK.n89 0.00531334
R21856 CLK.n85 CLK.n81 0.00531334
R21857 CLK.n77 CLK.n73 0.00531334
R21858 CLK.n69 CLK.n65 0.00531334
R21859 CLK.n61 CLK.n57 0.00531334
R21860 CLK.n53 CLK.n49 0.00531334
R21861 CLK.n45 CLK.n41 0.00531334
R21862 CLK.n37 CLK.n33 0.00531334
R21863 CLK.n29 CLK.n25 0.00531334
R21864 CLK.n21 CLK.n17 0.00531334
R21865 CLK.n13 CLK.n9 0.00531334
R21866 CLK.n139 CLK.n136 0.00531334
R21867 CLK.n4 CLK.n3 0.00224847
R21868 CLK.n117 CLK.n116 0.00224847
R21869 CLK.n109 CLK.n108 0.00224847
R21870 CLK.n101 CLK.n100 0.00224847
R21871 CLK.n93 CLK.n92 0.00224847
R21872 CLK.n85 CLK.n84 0.00224847
R21873 CLK.n77 CLK.n76 0.00224847
R21874 CLK.n69 CLK.n68 0.00224847
R21875 CLK.n61 CLK.n60 0.00224847
R21876 CLK.n53 CLK.n52 0.00224847
R21877 CLK.n45 CLK.n44 0.00224847
R21878 CLK.n37 CLK.n36 0.00224847
R21879 CLK.n29 CLK.n28 0.00224847
R21880 CLK.n21 CLK.n20 0.00224847
R21881 CLK.n13 CLK.n12 0.00224847
R21882 CLK.n139 CLK.n138 0.00224847
R21883 CLK.n3 CLK.n1 0.00100535
R21884 CLK.n116 CLK.n114 0.00100535
R21885 CLK.n108 CLK.n106 0.00100535
R21886 CLK.n100 CLK.n98 0.00100535
R21887 CLK.n92 CLK.n90 0.00100535
R21888 CLK.n84 CLK.n82 0.00100535
R21889 CLK.n76 CLK.n74 0.00100535
R21890 CLK.n68 CLK.n66 0.00100535
R21891 CLK.n60 CLK.n58 0.00100535
R21892 CLK.n52 CLK.n50 0.00100535
R21893 CLK.n44 CLK.n42 0.00100535
R21894 CLK.n36 CLK.n34 0.00100535
R21895 CLK.n28 CLK.n26 0.00100535
R21896 CLK.n20 CLK.n18 0.00100535
R21897 CLK.n12 CLK.n10 0.00100535
R21898 CLK.n138 CLK.n137 0.00100535
R21899 frontAnalog_v0p0p1_10.x65.A.n1 frontAnalog_v0p0p1_10.x65.A.t4 260.322
R21900 frontAnalog_v0p0p1_10.x65.A.n3 frontAnalog_v0p0p1_10.x65.A.t7 233.929
R21901 frontAnalog_v0p0p1_10.x65.A.n1 frontAnalog_v0p0p1_10.x65.A.t6 175.169
R21902 frontAnalog_v0p0p1_10.x65.A.n2 frontAnalog_v0p0p1_10.x65.A.t5 160.416
R21903 frontAnalog_v0p0p1_10.x65.A.n4 frontAnalog_v0p0p1_10.x65.A.t1 17.4109
R21904 frontAnalog_v0p0p1_10.x65.A.n4 frontAnalog_v0p0p1_10.x65.A.t0 10.2053
R21905 frontAnalog_v0p0p1_10.x65.A.n0 frontAnalog_v0p0p1_10.x65.A 2.78715
R21906 frontAnalog_v0p0p1_10.x65.A.n0 frontAnalog_v0p0p1_10.x65.A.n1 9.09103
R21907 frontAnalog_v0p0p1_10.x65.A.n6 frontAnalog_v0p0p1_10.x65.A.t3 7.94569
R21908 frontAnalog_v0p0p1_10.x65.A.n2 frontAnalog_v0p0p1_10.x65.A.t2 7.55846
R21909 frontAnalog_v0p0p1_10.x65.A.n5 frontAnalog_v0p0p1_10.x65.A.n3 1.4614
R21910 frontAnalog_v0p0p1_10.x65.A.n3 frontAnalog_v0p0p1_10.x65.A.n2 1.19626
R21911 frontAnalog_v0p0p1_10.x65.A.n6 frontAnalog_v0p0p1_10.x65.A.n5 0.836961
R21912 frontAnalog_v0p0p1_10.x65.A frontAnalog_v0p0p1_10.x65.A.n0 0.390342
R21913 frontAnalog_v0p0p1_10.x65.A.n5 frontAnalog_v0p0p1_10.x65.A.n4 0.154668
R21914 frontAnalog_v0p0p1_10.x65.A frontAnalog_v0p0p1_10.x65.A.n6 0.08175
R21915 resistorDivider_v0p0p1_0.V4.n0 resistorDivider_v0p0p1_0.V4.t17 167.365
R21916 resistorDivider_v0p0p1_0.V4.n0 resistorDivider_v0p0p1_0.V4.t16 92.4488
R21917 resistorDivider_v0p0p1_0.V4.n1 resistorDivider_v0p0p1_0.V4.n0 2.07493
R21918 resistorDivider_v0p0p1_0.V4.n9 resistorDivider_v0p0p1_0.V4.n8 0.141636
R21919 resistorDivider_v0p0p1_0.V4.n8 resistorDivider_v0p0p1_0.V4.n7 0.141636
R21920 resistorDivider_v0p0p1_0.V4.n7 resistorDivider_v0p0p1_0.V4.n6 0.141636
R21921 resistorDivider_v0p0p1_0.V4.n6 resistorDivider_v0p0p1_0.V4.n5 0.141636
R21922 resistorDivider_v0p0p1_0.V4.n5 resistorDivider_v0p0p1_0.V4.n4 0.141636
R21923 resistorDivider_v0p0p1_0.V4.n4 resistorDivider_v0p0p1_0.V4.n3 0.141636
R21924 resistorDivider_v0p0p1_0.V4.n3 resistorDivider_v0p0p1_0.V4.n2 0.141636
R21925 resistorDivider_v0p0p1_0.V4.n1 resistorDivider_v0p0p1_0.V4 0.12425
R21926 resistorDivider_v0p0p1_0.V4 resistorDivider_v0p0p1_0.V4.n9 0.103284
R21927 resistorDivider_v0p0p1_0.V4 resistorDivider_v0p0p1_0.V4.n1 0.0314375
R21928 resistorDivider_v0p0p1_0.V4.n7 resistorDivider_v0p0p1_0.V4.t0 0.00250214
R21929 resistorDivider_v0p0p1_0.V4.n3 resistorDivider_v0p0p1_0.V4.t15 0.000502142
R21930 resistorDivider_v0p0p1_0.V4.n4 resistorDivider_v0p0p1_0.V4.t2 0.000502142
R21931 resistorDivider_v0p0p1_0.V4.n5 resistorDivider_v0p0p1_0.V4.t6 0.000502142
R21932 resistorDivider_v0p0p1_0.V4.n6 resistorDivider_v0p0p1_0.V4.t9 0.000502142
R21933 resistorDivider_v0p0p1_0.V4.n7 resistorDivider_v0p0p1_0.V4.t11 0.000502142
R21934 resistorDivider_v0p0p1_0.V4.n8 resistorDivider_v0p0p1_0.V4.t7 0.000502142
R21935 resistorDivider_v0p0p1_0.V4.n9 resistorDivider_v0p0p1_0.V4.t3 0.000502142
R21936 resistorDivider_v0p0p1_0.V4.n2 resistorDivider_v0p0p1_0.V4.t1 0.000502142
R21937 resistorDivider_v0p0p1_0.V4.n3 resistorDivider_v0p0p1_0.V4.t4 0.000502142
R21938 resistorDivider_v0p0p1_0.V4.n4 resistorDivider_v0p0p1_0.V4.t14 0.000502142
R21939 resistorDivider_v0p0p1_0.V4.n5 resistorDivider_v0p0p1_0.V4.t12 0.000502142
R21940 resistorDivider_v0p0p1_0.V4.n6 resistorDivider_v0p0p1_0.V4.t8 0.000502142
R21941 resistorDivider_v0p0p1_0.V4.n8 resistorDivider_v0p0p1_0.V4.t10 0.000502142
R21942 resistorDivider_v0p0p1_0.V4.n9 resistorDivider_v0p0p1_0.V4.t5 0.000502142
R21943 resistorDivider_v0p0p1_0.V4.n2 resistorDivider_v0p0p1_0.V4.t13 0.000502142
R21944 resistorDivider_v0p0p1_0.V3.n0 resistorDivider_v0p0p1_0.V3.t17 167.365
R21945 resistorDivider_v0p0p1_0.V3.n0 resistorDivider_v0p0p1_0.V3.t16 92.4488
R21946 resistorDivider_v0p0p1_0.V3.n1 resistorDivider_v0p0p1_0.V3.n0 2.07493
R21947 resistorDivider_v0p0p1_0.V3.n15 resistorDivider_v0p0p1_0.V3.n14 0.141409
R21948 resistorDivider_v0p0p1_0.V3.n13 resistorDivider_v0p0p1_0.V3.n12 0.141409
R21949 resistorDivider_v0p0p1_0.V3.n11 resistorDivider_v0p0p1_0.V3.n10 0.141409
R21950 resistorDivider_v0p0p1_0.V3.n9 resistorDivider_v0p0p1_0.V3.n8 0.141409
R21951 resistorDivider_v0p0p1_0.V3.n7 resistorDivider_v0p0p1_0.V3.n6 0.141409
R21952 resistorDivider_v0p0p1_0.V3.n5 resistorDivider_v0p0p1_0.V3.n4 0.141409
R21953 resistorDivider_v0p0p1_0.V3.n3 resistorDivider_v0p0p1_0.V3.n2 0.141409
R21954 resistorDivider_v0p0p1_0.V3.n1 resistorDivider_v0p0p1_0.V3 0.12425
R21955 resistorDivider_v0p0p1_0.V3 resistorDivider_v0p0p1_0.V3.n16 0.100973
R21956 resistorDivider_v0p0p1_0.V3 resistorDivider_v0p0p1_0.V3.n1 0.0314375
R21957 resistorDivider_v0p0p1_0.V3.n11 resistorDivider_v0p0p1_0.V3.t0 0.00250214
R21958 resistorDivider_v0p0p1_0.V3.n2 resistorDivider_v0p0p1_0.V3.t1 0.000729415
R21959 resistorDivider_v0p0p1_0.V3.n16 resistorDivider_v0p0p1_0.V3.n15 0.000727273
R21960 resistorDivider_v0p0p1_0.V3.n14 resistorDivider_v0p0p1_0.V3.n13 0.000727273
R21961 resistorDivider_v0p0p1_0.V3.n12 resistorDivider_v0p0p1_0.V3.n11 0.000727273
R21962 resistorDivider_v0p0p1_0.V3.n10 resistorDivider_v0p0p1_0.V3.n9 0.000727273
R21963 resistorDivider_v0p0p1_0.V3.n8 resistorDivider_v0p0p1_0.V3.n7 0.000727273
R21964 resistorDivider_v0p0p1_0.V3.n6 resistorDivider_v0p0p1_0.V3.n5 0.000727273
R21965 resistorDivider_v0p0p1_0.V3.n4 resistorDivider_v0p0p1_0.V3.n3 0.000727273
R21966 resistorDivider_v0p0p1_0.V3.n3 resistorDivider_v0p0p1_0.V3.t2 0.000502142
R21967 resistorDivider_v0p0p1_0.V3.n5 resistorDivider_v0p0p1_0.V3.t9 0.000502142
R21968 resistorDivider_v0p0p1_0.V3.n7 resistorDivider_v0p0p1_0.V3.t8 0.000502142
R21969 resistorDivider_v0p0p1_0.V3.n9 resistorDivider_v0p0p1_0.V3.t5 0.000502142
R21970 resistorDivider_v0p0p1_0.V3.n13 resistorDivider_v0p0p1_0.V3.t6 0.000502142
R21971 resistorDivider_v0p0p1_0.V3.n15 resistorDivider_v0p0p1_0.V3.t3 0.000502142
R21972 resistorDivider_v0p0p1_0.V3.n2 resistorDivider_v0p0p1_0.V3.t10 0.000502142
R21973 resistorDivider_v0p0p1_0.V3.n4 resistorDivider_v0p0p1_0.V3.t14 0.000502142
R21974 resistorDivider_v0p0p1_0.V3.n6 resistorDivider_v0p0p1_0.V3.t12 0.000502142
R21975 resistorDivider_v0p0p1_0.V3.n8 resistorDivider_v0p0p1_0.V3.t11 0.000502142
R21976 resistorDivider_v0p0p1_0.V3.n10 resistorDivider_v0p0p1_0.V3.t7 0.000502142
R21977 resistorDivider_v0p0p1_0.V3.n12 resistorDivider_v0p0p1_0.V3.t13 0.000502142
R21978 resistorDivider_v0p0p1_0.V3.n14 resistorDivider_v0p0p1_0.V3.t15 0.000502142
R21979 resistorDivider_v0p0p1_0.V3.n16 resistorDivider_v0p0p1_0.V3.t4 0.000502142
R21980 frontAnalog_v0p0p1_14.x63.A.n2 frontAnalog_v0p0p1_14.x63.A.t7 260.322
R21981 frontAnalog_v0p0p1_14.x63.A.n4 frontAnalog_v0p0p1_14.x63.A.t4 233.888
R21982 frontAnalog_v0p0p1_14.x63.A.n2 frontAnalog_v0p0p1_14.x63.A.t5 175.169
R21983 frontAnalog_v0p0p1_14.x63.A.n3 frontAnalog_v0p0p1_14.x63.A.t6 159.725
R21984 frontAnalog_v0p0p1_14.x63.A.n1 frontAnalog_v0p0p1_14.x63.A.t2 17.4109
R21985 frontAnalog_v0p0p1_14.x63.A.n0 frontAnalog_v0p0p1_14.x63.A.n2 9.75129
R21986 frontAnalog_v0p0p1_14.x63.A.n1 frontAnalog_v0p0p1_14.x63.A.t3 9.6037
R21987 frontAnalog_v0p0p1_14.x63.A.n0 frontAnalog_v0p0p1_14.x63.A 2.33338
R21988 frontAnalog_v0p0p1_14.x63.A.n5 frontAnalog_v0p0p1_14.x63.A.t1 8.40929
R21989 frontAnalog_v0p0p1_14.x63.A.n3 frontAnalog_v0p0p1_14.x63.A.t0 8.06629
R21990 frontAnalog_v0p0p1_14.x63.A.n4 frontAnalog_v0p0p1_14.x63.A.n3 1.73501
R21991 frontAnalog_v0p0p1_14.x63.A.n1 frontAnalog_v0p0p1_14.x63.A.n4 0.99025
R21992 frontAnalog_v0p0p1_14.x63.A.n5 frontAnalog_v0p0p1_14.x63.A.n1 0.853186
R21993 frontAnalog_v0p0p1_14.x63.A frontAnalog_v0p0p1_14.x63.A.n0 0.349517
R21994 frontAnalog_v0p0p1_14.x63.A frontAnalog_v0p0p1_14.x63.A.n5 0.24425
R21995 frontAnalog_v0p0p1_14.x65.A.n1 frontAnalog_v0p0p1_14.x65.A.t7 260.322
R21996 frontAnalog_v0p0p1_14.x65.A.n3 frontAnalog_v0p0p1_14.x65.A.t5 233.929
R21997 frontAnalog_v0p0p1_14.x65.A.n1 frontAnalog_v0p0p1_14.x65.A.t4 175.169
R21998 frontAnalog_v0p0p1_14.x65.A.n2 frontAnalog_v0p0p1_14.x65.A.t6 160.416
R21999 frontAnalog_v0p0p1_14.x65.A.n4 frontAnalog_v0p0p1_14.x65.A.t0 17.4109
R22000 frontAnalog_v0p0p1_14.x65.A.n4 frontAnalog_v0p0p1_14.x65.A.t1 10.2053
R22001 frontAnalog_v0p0p1_14.x65.A.n0 frontAnalog_v0p0p1_14.x65.A 2.78715
R22002 frontAnalog_v0p0p1_14.x65.A.n0 frontAnalog_v0p0p1_14.x65.A.n1 9.09103
R22003 frontAnalog_v0p0p1_14.x65.A.n6 frontAnalog_v0p0p1_14.x65.A.t2 7.94569
R22004 frontAnalog_v0p0p1_14.x65.A.n2 frontAnalog_v0p0p1_14.x65.A.t3 7.55846
R22005 frontAnalog_v0p0p1_14.x65.A.n5 frontAnalog_v0p0p1_14.x65.A.n3 1.4614
R22006 frontAnalog_v0p0p1_14.x65.A.n3 frontAnalog_v0p0p1_14.x65.A.n2 1.19626
R22007 frontAnalog_v0p0p1_14.x65.A.n6 frontAnalog_v0p0p1_14.x65.A.n5 0.836961
R22008 frontAnalog_v0p0p1_14.x65.A frontAnalog_v0p0p1_14.x65.A.n0 0.390342
R22009 frontAnalog_v0p0p1_14.x65.A.n5 frontAnalog_v0p0p1_14.x65.A.n4 0.154668
R22010 frontAnalog_v0p0p1_14.x65.A frontAnalog_v0p0p1_14.x65.A.n6 0.08175
R22011 frontAnalog_v0p0p1_5.RSfetsym_0.QN.n1 frontAnalog_v0p0p1_5.RSfetsym_0.QN.t6 117.511
R22012 frontAnalog_v0p0p1_5.RSfetsym_0.QN.n1 frontAnalog_v0p0p1_5.RSfetsym_0.QN.t5 110.698
R22013 frontAnalog_v0p0p1_5.RSfetsym_0.QN.n4 frontAnalog_v0p0p1_5.RSfetsym_0.QN.t0 19.1963
R22014 frontAnalog_v0p0p1_5.RSfetsym_0.QN.n7 frontAnalog_v0p0p1_5.RSfetsym_0.QN.t4 14.2842
R22015 frontAnalog_v0p0p1_5.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_5.RSfetsym_0.QN.t2 14.283
R22016 frontAnalog_v0p0p1_5.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_5.RSfetsym_0.QN.t1 14.283
R22017 frontAnalog_v0p0p1_5.RSfetsym_0.QN.n11 frontAnalog_v0p0p1_5.RSfetsym_0.QN.t3 9.14075
R22018 frontAnalog_v0p0p1_5.RSfetsym_0.QN.n11 frontAnalog_v0p0p1_5.RSfetsym_0.QN.n10 0.74645
R22019 frontAnalog_v0p0p1_5.RSfetsym_0.QN.n2 frontAnalog_v0p0p1_5.RSfetsym_0.QN.n1 0.688382
R22020 frontAnalog_v0p0p1_5.RSfetsym_0.QN.n10 frontAnalog_v0p0p1_5.RSfetsym_0.QN.n9 0.2402
R22021 frontAnalog_v0p0p1_5.RSfetsym_0.QN.n9 frontAnalog_v0p0p1_5.RSfetsym_0.QN.n8 0.236824
R22022 frontAnalog_v0p0p1_5.RSfetsym_0.QN.n4 frontAnalog_v0p0p1_5.RSfetsym_0.QN.n3 0.132187
R22023 frontAnalog_v0p0p1_5.RSfetsym_0.QN.n9 frontAnalog_v0p0p1_5.RSfetsym_0.QN.n4 0.0968646
R22024 frontAnalog_v0p0p1_5.RSfetsym_0.QN frontAnalog_v0p0p1_5.RSfetsym_0.QN.n11 0.0446535
R22025 frontAnalog_v0p0p1_5.RSfetsym_0.QN.n8 frontAnalog_v0p0p1_5.RSfetsym_0.QN.n6 0.0272538
R22026 frontAnalog_v0p0p1_5.RSfetsym_0.QN.n10 frontAnalog_v0p0p1_5.RSfetsym_0.QN.n0 0.00981499
R22027 frontAnalog_v0p0p1_5.RSfetsym_0.QN.n3 frontAnalog_v0p0p1_5.RSfetsym_0.QN.n2 0.00725433
R22028 frontAnalog_v0p0p1_5.RSfetsym_0.QN.n6 frontAnalog_v0p0p1_5.RSfetsym_0.QN.n5 0.00610579
R22029 frontAnalog_v0p0p1_5.RSfetsym_0.QN.n8 frontAnalog_v0p0p1_5.RSfetsym_0.QN.n7 0.00225341
R22030 resistorDivider_v0p0p1_0.V11.n0 resistorDivider_v0p0p1_0.V11.t17 167.365
R22031 resistorDivider_v0p0p1_0.V11.n0 resistorDivider_v0p0p1_0.V11.t16 92.4496
R22032 resistorDivider_v0p0p1_0.V11.n1 resistorDivider_v0p0p1_0.V11.n0 2.07493
R22033 resistorDivider_v0p0p1_0.V11.n15 resistorDivider_v0p0p1_0.V11.n14 0.141409
R22034 resistorDivider_v0p0p1_0.V11.n13 resistorDivider_v0p0p1_0.V11.n12 0.141409
R22035 resistorDivider_v0p0p1_0.V11.n11 resistorDivider_v0p0p1_0.V11.n10 0.141409
R22036 resistorDivider_v0p0p1_0.V11.n9 resistorDivider_v0p0p1_0.V11.n8 0.141409
R22037 resistorDivider_v0p0p1_0.V11.n7 resistorDivider_v0p0p1_0.V11.n6 0.141409
R22038 resistorDivider_v0p0p1_0.V11.n5 resistorDivider_v0p0p1_0.V11.n4 0.141409
R22039 resistorDivider_v0p0p1_0.V11.n3 resistorDivider_v0p0p1_0.V11.n2 0.141409
R22040 resistorDivider_v0p0p1_0.V11.n1 resistorDivider_v0p0p1_0.V11 0.12425
R22041 resistorDivider_v0p0p1_0.V11 resistorDivider_v0p0p1_0.V11.n16 0.104098
R22042 resistorDivider_v0p0p1_0.V11 resistorDivider_v0p0p1_0.V11.n1 0.0314375
R22043 resistorDivider_v0p0p1_0.V11.n10 resistorDivider_v0p0p1_0.V11.t0 0.00250214
R22044 resistorDivider_v0p0p1_0.V11.n2 resistorDivider_v0p0p1_0.V11.t11 0.000729415
R22045 resistorDivider_v0p0p1_0.V11.n16 resistorDivider_v0p0p1_0.V11.n15 0.000727273
R22046 resistorDivider_v0p0p1_0.V11.n14 resistorDivider_v0p0p1_0.V11.n13 0.000727273
R22047 resistorDivider_v0p0p1_0.V11.n12 resistorDivider_v0p0p1_0.V11.n11 0.000727273
R22048 resistorDivider_v0p0p1_0.V11.n10 resistorDivider_v0p0p1_0.V11.n9 0.000727273
R22049 resistorDivider_v0p0p1_0.V11.n8 resistorDivider_v0p0p1_0.V11.n7 0.000727273
R22050 resistorDivider_v0p0p1_0.V11.n6 resistorDivider_v0p0p1_0.V11.n5 0.000727273
R22051 resistorDivider_v0p0p1_0.V11.n4 resistorDivider_v0p0p1_0.V11.n3 0.000727273
R22052 resistorDivider_v0p0p1_0.V11.n3 resistorDivider_v0p0p1_0.V11.t4 0.000502142
R22053 resistorDivider_v0p0p1_0.V11.n5 resistorDivider_v0p0p1_0.V11.t2 0.000502142
R22054 resistorDivider_v0p0p1_0.V11.n7 resistorDivider_v0p0p1_0.V11.t13 0.000502142
R22055 resistorDivider_v0p0p1_0.V11.n9 resistorDivider_v0p0p1_0.V11.t15 0.000502142
R22056 resistorDivider_v0p0p1_0.V11.n11 resistorDivider_v0p0p1_0.V11.t3 0.000502142
R22057 resistorDivider_v0p0p1_0.V11.n13 resistorDivider_v0p0p1_0.V11.t1 0.000502142
R22058 resistorDivider_v0p0p1_0.V11.n15 resistorDivider_v0p0p1_0.V11.t6 0.000502142
R22059 resistorDivider_v0p0p1_0.V11.n16 resistorDivider_v0p0p1_0.V11.t14 0.000502142
R22060 resistorDivider_v0p0p1_0.V11.n14 resistorDivider_v0p0p1_0.V11.t5 0.000502142
R22061 resistorDivider_v0p0p1_0.V11.n12 resistorDivider_v0p0p1_0.V11.t9 0.000502142
R22062 resistorDivider_v0p0p1_0.V11.n8 resistorDivider_v0p0p1_0.V11.t12 0.000502142
R22063 resistorDivider_v0p0p1_0.V11.n6 resistorDivider_v0p0p1_0.V11.t10 0.000502142
R22064 resistorDivider_v0p0p1_0.V11.n4 resistorDivider_v0p0p1_0.V11.t8 0.000502142
R22065 resistorDivider_v0p0p1_0.V11.n2 resistorDivider_v0p0p1_0.V11.t7 0.000502142
R22066 resistorDivider_v0p0p1_0.V10.n0 resistorDivider_v0p0p1_0.V10.t16 167.365
R22067 resistorDivider_v0p0p1_0.V10.n0 resistorDivider_v0p0p1_0.V10.t17 92.4496
R22068 resistorDivider_v0p0p1_0.V10.n1 resistorDivider_v0p0p1_0.V10.n0 2.07493
R22069 resistorDivider_v0p0p1_0.V10.n9 resistorDivider_v0p0p1_0.V10.n8 0.141636
R22070 resistorDivider_v0p0p1_0.V10.n8 resistorDivider_v0p0p1_0.V10.n7 0.141636
R22071 resistorDivider_v0p0p1_0.V10.n7 resistorDivider_v0p0p1_0.V10.n6 0.141636
R22072 resistorDivider_v0p0p1_0.V10.n6 resistorDivider_v0p0p1_0.V10.n5 0.141636
R22073 resistorDivider_v0p0p1_0.V10.n5 resistorDivider_v0p0p1_0.V10.n4 0.141636
R22074 resistorDivider_v0p0p1_0.V10.n4 resistorDivider_v0p0p1_0.V10.n3 0.141636
R22075 resistorDivider_v0p0p1_0.V10.n3 resistorDivider_v0p0p1_0.V10.n2 0.141636
R22076 resistorDivider_v0p0p1_0.V10.n1 resistorDivider_v0p0p1_0.V10 0.12425
R22077 resistorDivider_v0p0p1_0.V10 resistorDivider_v0p0p1_0.V10.n9 0.104326
R22078 resistorDivider_v0p0p1_0.V10 resistorDivider_v0p0p1_0.V10.n1 0.028
R22079 resistorDivider_v0p0p1_0.V10.n2 resistorDivider_v0p0p1_0.V10.t0 0.00250214
R22080 resistorDivider_v0p0p1_0.V10.n3 resistorDivider_v0p0p1_0.V10.t13 0.000502142
R22081 resistorDivider_v0p0p1_0.V10.n4 resistorDivider_v0p0p1_0.V10.t12 0.000502142
R22082 resistorDivider_v0p0p1_0.V10.n5 resistorDivider_v0p0p1_0.V10.t9 0.000502142
R22083 resistorDivider_v0p0p1_0.V10.n6 resistorDivider_v0p0p1_0.V10.t7 0.000502142
R22084 resistorDivider_v0p0p1_0.V10.n7 resistorDivider_v0p0p1_0.V10.t15 0.000502142
R22085 resistorDivider_v0p0p1_0.V10.n8 resistorDivider_v0p0p1_0.V10.t11 0.000502142
R22086 resistorDivider_v0p0p1_0.V10.n9 resistorDivider_v0p0p1_0.V10.t1 0.000502142
R22087 resistorDivider_v0p0p1_0.V10.n9 resistorDivider_v0p0p1_0.V10.t6 0.000502142
R22088 resistorDivider_v0p0p1_0.V10.n8 resistorDivider_v0p0p1_0.V10.t2 0.000502142
R22089 resistorDivider_v0p0p1_0.V10.n7 resistorDivider_v0p0p1_0.V10.t4 0.000502142
R22090 resistorDivider_v0p0p1_0.V10.n6 resistorDivider_v0p0p1_0.V10.t14 0.000502142
R22091 resistorDivider_v0p0p1_0.V10.n5 resistorDivider_v0p0p1_0.V10.t10 0.000502142
R22092 resistorDivider_v0p0p1_0.V10.n4 resistorDivider_v0p0p1_0.V10.t3 0.000502142
R22093 resistorDivider_v0p0p1_0.V10.n3 resistorDivider_v0p0p1_0.V10.t5 0.000502142
R22094 resistorDivider_v0p0p1_0.V10.n2 resistorDivider_v0p0p1_0.V10.t8 0.000502142
R22095 resistorDivider_v0p0p1_0.V2.n0 resistorDivider_v0p0p1_0.V2.t16 167.365
R22096 resistorDivider_v0p0p1_0.V2.n0 resistorDivider_v0p0p1_0.V2.t17 92.4488
R22097 resistorDivider_v0p0p1_0.V2.n1 resistorDivider_v0p0p1_0.V2.n0 2.07493
R22098 resistorDivider_v0p0p1_0.V2.n15 resistorDivider_v0p0p1_0.V2.n14 0.141409
R22099 resistorDivider_v0p0p1_0.V2.n13 resistorDivider_v0p0p1_0.V2.n12 0.141409
R22100 resistorDivider_v0p0p1_0.V2.n11 resistorDivider_v0p0p1_0.V2.n10 0.141409
R22101 resistorDivider_v0p0p1_0.V2.n9 resistorDivider_v0p0p1_0.V2.n8 0.141409
R22102 resistorDivider_v0p0p1_0.V2.n7 resistorDivider_v0p0p1_0.V2.n6 0.141409
R22103 resistorDivider_v0p0p1_0.V2.n5 resistorDivider_v0p0p1_0.V2.n4 0.141409
R22104 resistorDivider_v0p0p1_0.V2.n3 resistorDivider_v0p0p1_0.V2.n2 0.141409
R22105 resistorDivider_v0p0p1_0.V2.n1 resistorDivider_v0p0p1_0.V2 0.12425
R22106 resistorDivider_v0p0p1_0.V2 resistorDivider_v0p0p1_0.V2.n16 0.0968068
R22107 resistorDivider_v0p0p1_0.V2 resistorDivider_v0p0p1_0.V2.n1 0.028
R22108 resistorDivider_v0p0p1_0.V2.n15 resistorDivider_v0p0p1_0.V2.t0 0.00250214
R22109 resistorDivider_v0p0p1_0.V2.n2 resistorDivider_v0p0p1_0.V2.t5 0.000729415
R22110 resistorDivider_v0p0p1_0.V2.n16 resistorDivider_v0p0p1_0.V2.n15 0.000727273
R22111 resistorDivider_v0p0p1_0.V2.n14 resistorDivider_v0p0p1_0.V2.n13 0.000727273
R22112 resistorDivider_v0p0p1_0.V2.n12 resistorDivider_v0p0p1_0.V2.n11 0.000727273
R22113 resistorDivider_v0p0p1_0.V2.n10 resistorDivider_v0p0p1_0.V2.n9 0.000727273
R22114 resistorDivider_v0p0p1_0.V2.n8 resistorDivider_v0p0p1_0.V2.n7 0.000727273
R22115 resistorDivider_v0p0p1_0.V2.n6 resistorDivider_v0p0p1_0.V2.n5 0.000727273
R22116 resistorDivider_v0p0p1_0.V2.n4 resistorDivider_v0p0p1_0.V2.n3 0.000727273
R22117 resistorDivider_v0p0p1_0.V2.n4 resistorDivider_v0p0p1_0.V2.t14 0.000502142
R22118 resistorDivider_v0p0p1_0.V2.n6 resistorDivider_v0p0p1_0.V2.t12 0.000502142
R22119 resistorDivider_v0p0p1_0.V2.n8 resistorDivider_v0p0p1_0.V2.t10 0.000502142
R22120 resistorDivider_v0p0p1_0.V2.n10 resistorDivider_v0p0p1_0.V2.t6 0.000502142
R22121 resistorDivider_v0p0p1_0.V2.n12 resistorDivider_v0p0p1_0.V2.t13 0.000502142
R22122 resistorDivider_v0p0p1_0.V2.n14 resistorDivider_v0p0p1_0.V2.t15 0.000502142
R22123 resistorDivider_v0p0p1_0.V2.n16 resistorDivider_v0p0p1_0.V2.t2 0.000502142
R22124 resistorDivider_v0p0p1_0.V2.n3 resistorDivider_v0p0p1_0.V2.t3 0.000502142
R22125 resistorDivider_v0p0p1_0.V2.n5 resistorDivider_v0p0p1_0.V2.t8 0.000502142
R22126 resistorDivider_v0p0p1_0.V2.n7 resistorDivider_v0p0p1_0.V2.t4 0.000502142
R22127 resistorDivider_v0p0p1_0.V2.n9 resistorDivider_v0p0p1_0.V2.t7 0.000502142
R22128 resistorDivider_v0p0p1_0.V2.n11 resistorDivider_v0p0p1_0.V2.t1 0.000502142
R22129 resistorDivider_v0p0p1_0.V2.n13 resistorDivider_v0p0p1_0.V2.t11 0.000502142
R22130 resistorDivider_v0p0p1_0.V2.n2 resistorDivider_v0p0p1_0.V2.t9 0.000502142
R22131 resistorDivider_v0p0p1_0.V1.n0 resistorDivider_v0p0p1_0.V1.t17 167.365
R22132 resistorDivider_v0p0p1_0.V1.n0 resistorDivider_v0p0p1_0.V1.t16 92.4488
R22133 resistorDivider_v0p0p1_0.V1.n1 resistorDivider_v0p0p1_0.V1.n0 2.07493
R22134 resistorDivider_v0p0p1_0.V1.n9 resistorDivider_v0p0p1_0.V1.n8 0.141636
R22135 resistorDivider_v0p0p1_0.V1.n8 resistorDivider_v0p0p1_0.V1.n7 0.141636
R22136 resistorDivider_v0p0p1_0.V1.n7 resistorDivider_v0p0p1_0.V1.n6 0.141636
R22137 resistorDivider_v0p0p1_0.V1.n6 resistorDivider_v0p0p1_0.V1.n5 0.141636
R22138 resistorDivider_v0p0p1_0.V1.n5 resistorDivider_v0p0p1_0.V1.n4 0.141636
R22139 resistorDivider_v0p0p1_0.V1.n4 resistorDivider_v0p0p1_0.V1.n3 0.141636
R22140 resistorDivider_v0p0p1_0.V1.n3 resistorDivider_v0p0p1_0.V1.n2 0.141636
R22141 resistorDivider_v0p0p1_0.V1.n1 resistorDivider_v0p0p1_0.V1 0.12425
R22142 resistorDivider_v0p0p1_0.V1 resistorDivider_v0p0p1_0.V1.n9 0.0980758
R22143 resistorDivider_v0p0p1_0.V1 resistorDivider_v0p0p1_0.V1.n1 0.0314375
R22144 resistorDivider_v0p0p1_0.V1.n9 resistorDivider_v0p0p1_0.V1.t0 0.00250214
R22145 resistorDivider_v0p0p1_0.V1.n3 resistorDivider_v0p0p1_0.V1.t3 0.000502142
R22146 resistorDivider_v0p0p1_0.V1.n4 resistorDivider_v0p0p1_0.V1.t12 0.000502142
R22147 resistorDivider_v0p0p1_0.V1.n5 resistorDivider_v0p0p1_0.V1.t5 0.000502142
R22148 resistorDivider_v0p0p1_0.V1.n6 resistorDivider_v0p0p1_0.V1.t11 0.000502142
R22149 resistorDivider_v0p0p1_0.V1.n7 resistorDivider_v0p0p1_0.V1.t1 0.000502142
R22150 resistorDivider_v0p0p1_0.V1.n8 resistorDivider_v0p0p1_0.V1.t14 0.000502142
R22151 resistorDivider_v0p0p1_0.V1.n2 resistorDivider_v0p0p1_0.V1.t9 0.000502142
R22152 resistorDivider_v0p0p1_0.V1.n3 resistorDivider_v0p0p1_0.V1.t7 0.000502142
R22153 resistorDivider_v0p0p1_0.V1.n4 resistorDivider_v0p0p1_0.V1.t4 0.000502142
R22154 resistorDivider_v0p0p1_0.V1.n5 resistorDivider_v0p0p1_0.V1.t6 0.000502142
R22155 resistorDivider_v0p0p1_0.V1.n6 resistorDivider_v0p0p1_0.V1.t15 0.000502142
R22156 resistorDivider_v0p0p1_0.V1.n7 resistorDivider_v0p0p1_0.V1.t13 0.000502142
R22157 resistorDivider_v0p0p1_0.V1.n8 resistorDivider_v0p0p1_0.V1.t10 0.000502142
R22158 resistorDivider_v0p0p1_0.V1.n9 resistorDivider_v0p0p1_0.V1.t2 0.000502142
R22159 resistorDivider_v0p0p1_0.V1.n2 resistorDivider_v0p0p1_0.V1.t8 0.000502142
R22160 frontAnalog_v0p0p1_15.Q.n0 frontAnalog_v0p0p1_15.Q.t5 196.549
R22161 frontAnalog_v0p0p1_15.Q.n0 frontAnalog_v0p0p1_15.Q.t7 148.35
R22162 frontAnalog_v0p0p1_15.Q.n4 frontAnalog_v0p0p1_15.Q.t8 117.314
R22163 frontAnalog_v0p0p1_15.Q.n4 frontAnalog_v0p0p1_15.Q.t6 110.853
R22164 frontAnalog_v0p0p1_15.Q.n5 frontAnalog_v0p0p1_15.Q.t2 17.6181
R22165 frontAnalog_v0p0p1_15.Q.n7 frontAnalog_v0p0p1_15.Q.t0 14.2865
R22166 frontAnalog_v0p0p1_15.Q.n9 frontAnalog_v0p0p1_15.Q.t3 14.283
R22167 frontAnalog_v0p0p1_15.Q.n9 frontAnalog_v0p0p1_15.Q.t4 14.283
R22168 frontAnalog_v0p0p1_15.Q.n12 frontAnalog_v0p0p1_15.Q.n3 10.185
R22169 frontAnalog_v0p0p1_15.Q.n1 frontAnalog_v0p0p1_15.Q.n0 9.49592
R22170 frontAnalog_v0p0p1_15.Q.n11 frontAnalog_v0p0p1_15.Q.t1 8.77744
R22171 frontAnalog_v0p0p1_15.Q.n2 frontAnalog_v0p0p1_15.Q.n1 7.58085
R22172 frontAnalog_v0p0p1_15.Q.n1 frontAnalog_v0p0p1_15.Q 6.44187
R22173 frontAnalog_v0p0p1_15.Q.n3 frontAnalog_v0p0p1_15.Q.n2 2.50858
R22174 frontAnalog_v0p0p1_15.Q.n11 frontAnalog_v0p0p1_15.Q.n10 1.20426
R22175 frontAnalog_v0p0p1_15.Q.n2 frontAnalog_v0p0p1_15.Q 0.88934
R22176 frontAnalog_v0p0p1_15.Q.n12 frontAnalog_v0p0p1_15.Q.n11 0.325111
R22177 frontAnalog_v0p0p1_15.Q.n8 frontAnalog_v0p0p1_15.Q.n7 0.301242
R22178 frontAnalog_v0p0p1_15.Q.n3 frontAnalog_v0p0p1_15.Q 0.2005
R22179 frontAnalog_v0p0p1_15.Q.n6 frontAnalog_v0p0p1_15.Q.n4 0.159555
R22180 frontAnalog_v0p0p1_15.Q.n10 frontAnalog_v0p0p1_15.Q.n9 0.106617
R22181 frontAnalog_v0p0p1_15.Q.n8 frontAnalog_v0p0p1_15.Q.n6 0.0796167
R22182 frontAnalog_v0p0p1_15.Q.n10 frontAnalog_v0p0p1_15.Q.n8 0.0480595
R22183 frontAnalog_v0p0p1_15.Q frontAnalog_v0p0p1_15.Q.n12 0.0469368
R22184 frontAnalog_v0p0p1_15.Q.n6 frontAnalog_v0p0p1_15.Q.n5 0.000504658
R22185 frontAnalog_v0p0p1_12.Q.n6 frontAnalog_v0p0p1_12.Q.t5 323.342
R22186 frontAnalog_v0p0p1_12.Q.n0 frontAnalog_v0p0p1_12.Q.t9 228.927
R22187 frontAnalog_v0p0p1_12.Q.n3 frontAnalog_v0p0p1_12.Q.t7 196.549
R22188 frontAnalog_v0p0p1_12.Q.n6 frontAnalog_v0p0p1_12.Q.t8 194.809
R22189 frontAnalog_v0p0p1_12.Q.n0 frontAnalog_v0p0p1_12.Q.t6 159.391
R22190 frontAnalog_v0p0p1_12.Q.n3 frontAnalog_v0p0p1_12.Q.t11 148.35
R22191 frontAnalog_v0p0p1_12.Q.n10 frontAnalog_v0p0p1_12.Q.t12 117.314
R22192 frontAnalog_v0p0p1_12.Q.n10 frontAnalog_v0p0p1_12.Q.t10 110.853
R22193 frontAnalog_v0p0p1_12.Q.n7 frontAnalog_v0p0p1_12.Q.n6 76.0005
R22194 frontAnalog_v0p0p1_12.Q.n4 frontAnalog_v0p0p1_12.Q.n3 76.0005
R22195 frontAnalog_v0p0p1_12.Q.n8 frontAnalog_v0p0p1_12.Q.n7 29.2624
R22196 frontAnalog_v0p0p1_12.Q.n11 frontAnalog_v0p0p1_12.Q.t1 17.6181
R22197 frontAnalog_v0p0p1_12.Q.n13 frontAnalog_v0p0p1_12.Q.t0 14.2865
R22198 frontAnalog_v0p0p1_12.Q.n15 frontAnalog_v0p0p1_12.Q.t2 14.283
R22199 frontAnalog_v0p0p1_12.Q.n15 frontAnalog_v0p0p1_12.Q.t3 14.283
R22200 frontAnalog_v0p0p1_12.Q.n5 frontAnalog_v0p0p1_12.Q 9.11
R22201 frontAnalog_v0p0p1_12.Q.n17 frontAnalog_v0p0p1_12.Q.t4 8.77744
R22202 frontAnalog_v0p0p1_12.Q.n1 frontAnalog_v0p0p1_12.Q.n0 8.68501
R22203 frontAnalog_v0p0p1_12.Q.n18 frontAnalog_v0p0p1_12.Q.n9 7.84168
R22204 frontAnalog_v0p0p1_12.Q.n4 frontAnalog_v0p0p1_12.Q 5.78114
R22205 frontAnalog_v0p0p1_12.Q.n2 frontAnalog_v0p0p1_12.Q.n1 4.26764
R22206 frontAnalog_v0p0p1_12.Q frontAnalog_v0p0p1_12.Q.n4 3.71663
R22207 frontAnalog_v0p0p1_12.Q.n1 frontAnalog_v0p0p1_12.Q 1.99697
R22208 frontAnalog_v0p0p1_12.Q.n7 frontAnalog_v0p0p1_12.Q 1.92927
R22209 frontAnalog_v0p0p1_12.Q.n8 frontAnalog_v0p0p1_12.Q.n5 1.79514
R22210 frontAnalog_v0p0p1_12.Q.n17 frontAnalog_v0p0p1_12.Q.n16 1.20426
R22211 frontAnalog_v0p0p1_12.Q.n5 frontAnalog_v0p0p1_12.Q.n2 0.570143
R22212 frontAnalog_v0p0p1_12.Q.n18 frontAnalog_v0p0p1_12.Q.n17 0.325111
R22213 frontAnalog_v0p0p1_12.Q.n14 frontAnalog_v0p0p1_12.Q.n13 0.301242
R22214 frontAnalog_v0p0p1_12.Q.n9 frontAnalog_v0p0p1_12.Q.n8 0.226885
R22215 frontAnalog_v0p0p1_12.Q.n2 frontAnalog_v0p0p1_12.Q 0.221483
R22216 frontAnalog_v0p0p1_12.Q.n9 frontAnalog_v0p0p1_12.Q 0.20675
R22217 frontAnalog_v0p0p1_12.Q.n12 frontAnalog_v0p0p1_12.Q.n10 0.159555
R22218 frontAnalog_v0p0p1_12.Q.n16 frontAnalog_v0p0p1_12.Q.n15 0.106617
R22219 frontAnalog_v0p0p1_12.Q.n14 frontAnalog_v0p0p1_12.Q.n12 0.0796167
R22220 frontAnalog_v0p0p1_12.Q.n16 frontAnalog_v0p0p1_12.Q.n14 0.0480595
R22221 frontAnalog_v0p0p1_12.Q frontAnalog_v0p0p1_12.Q.n18 0.0469368
R22222 frontAnalog_v0p0p1_12.Q.n12 frontAnalog_v0p0p1_12.Q.n11 0.000504658
R22223 OUT1.n122 OUT1.n120 145.809
R22224 OUT1.n65 OUT1.n63 145.809
R22225 OUT1.n25 OUT1.n23 145.809
R22226 OUT1.n102 OUT1.n100 145.808
R22227 OUT1.n65 OUT1.n64 107.409
R22228 OUT1.n67 OUT1.n66 107.409
R22229 OUT1.n69 OUT1.n68 107.409
R22230 OUT1.n71 OUT1.n70 107.409
R22231 OUT1.n73 OUT1.n72 107.409
R22232 OUT1.n75 OUT1.n74 107.409
R22233 OUT1.n25 OUT1.n24 107.409
R22234 OUT1.n27 OUT1.n26 107.409
R22235 OUT1.n29 OUT1.n28 107.409
R22236 OUT1.n31 OUT1.n30 107.409
R22237 OUT1.n33 OUT1.n32 107.409
R22238 OUT1.n35 OUT1.n34 107.409
R22239 OUT1.n122 OUT1.n121 107.407
R22240 OUT1.n124 OUT1.n123 107.407
R22241 OUT1.n126 OUT1.n125 107.407
R22242 OUT1.n128 OUT1.n127 107.407
R22243 OUT1.n130 OUT1.n129 107.407
R22244 OUT1.n132 OUT1.n131 107.407
R22245 OUT1.n102 OUT1.n101 107.407
R22246 OUT1.n104 OUT1.n103 107.407
R22247 OUT1.n106 OUT1.n105 107.407
R22248 OUT1.n108 OUT1.n107 107.407
R22249 OUT1.n110 OUT1.n109 107.407
R22250 OUT1.n112 OUT1.n111 107.407
R22251 OUT1.n138 OUT1.n136 87.1779
R22252 OUT1.n83 OUT1.n81 87.1779
R22253 OUT1.n44 OUT1.n42 87.1779
R22254 OUT1.n4 OUT1.n2 87.1779
R22255 OUT1.n54 OUT1.n53 52.82
R22256 OUT1.n14 OUT1.n13 52.82
R22257 OUT1.n138 OUT1.n137 52.82
R22258 OUT1.n140 OUT1.n139 52.82
R22259 OUT1.n142 OUT1.n141 52.82
R22260 OUT1.n144 OUT1.n143 52.82
R22261 OUT1.n146 OUT1.n145 52.82
R22262 OUT1.n148 OUT1.n147 52.82
R22263 OUT1.n83 OUT1.n82 52.82
R22264 OUT1.n85 OUT1.n84 52.82
R22265 OUT1.n87 OUT1.n86 52.82
R22266 OUT1.n89 OUT1.n88 52.82
R22267 OUT1.n91 OUT1.n90 52.82
R22268 OUT1.n93 OUT1.n92 52.82
R22269 OUT1.n44 OUT1.n43 52.82
R22270 OUT1.n46 OUT1.n45 52.82
R22271 OUT1.n48 OUT1.n47 52.82
R22272 OUT1.n50 OUT1.n49 52.82
R22273 OUT1.n52 OUT1.n51 52.82
R22274 OUT1.n4 OUT1.n3 52.82
R22275 OUT1.n6 OUT1.n5 52.82
R22276 OUT1.n8 OUT1.n7 52.82
R22277 OUT1.n10 OUT1.n9 52.82
R22278 OUT1.n12 OUT1.n11 52.82
R22279 OUT1 OUT1.n149 51.0745
R22280 OUT1 OUT1.n94 51.0745
R22281 OUT1.n124 OUT1.n122 38.4005
R22282 OUT1.n126 OUT1.n124 38.4005
R22283 OUT1.n128 OUT1.n126 38.4005
R22284 OUT1.n130 OUT1.n128 38.4005
R22285 OUT1.n132 OUT1.n130 38.4005
R22286 OUT1.n133 OUT1.n132 38.4005
R22287 OUT1.n104 OUT1.n102 38.4005
R22288 OUT1.n106 OUT1.n104 38.4005
R22289 OUT1.n108 OUT1.n106 38.4005
R22290 OUT1.n110 OUT1.n108 38.4005
R22291 OUT1.n112 OUT1.n110 38.4005
R22292 OUT1.n113 OUT1.n112 38.4005
R22293 OUT1.n67 OUT1.n65 38.4005
R22294 OUT1.n69 OUT1.n67 38.4005
R22295 OUT1.n71 OUT1.n69 38.4005
R22296 OUT1.n73 OUT1.n71 38.4005
R22297 OUT1.n75 OUT1.n73 38.4005
R22298 OUT1.n76 OUT1.n75 38.4005
R22299 OUT1.n27 OUT1.n25 38.4005
R22300 OUT1.n29 OUT1.n27 38.4005
R22301 OUT1.n31 OUT1.n29 38.4005
R22302 OUT1.n33 OUT1.n31 38.4005
R22303 OUT1.n35 OUT1.n33 38.4005
R22304 OUT1.n36 OUT1.n35 38.4005
R22305 OUT1.n140 OUT1.n138 34.3584
R22306 OUT1.n142 OUT1.n140 34.3584
R22307 OUT1.n144 OUT1.n142 34.3584
R22308 OUT1.n146 OUT1.n144 34.3584
R22309 OUT1.n148 OUT1.n146 34.3584
R22310 OUT1.n150 OUT1.n148 34.3584
R22311 OUT1.n85 OUT1.n83 34.3584
R22312 OUT1.n87 OUT1.n85 34.3584
R22313 OUT1.n89 OUT1.n87 34.3584
R22314 OUT1.n91 OUT1.n89 34.3584
R22315 OUT1.n93 OUT1.n91 34.3584
R22316 OUT1.n95 OUT1.n93 34.3584
R22317 OUT1.n46 OUT1.n44 34.3584
R22318 OUT1.n48 OUT1.n46 34.3584
R22319 OUT1.n50 OUT1.n48 34.3584
R22320 OUT1.n52 OUT1.n50 34.3584
R22321 OUT1.n54 OUT1.n52 34.3584
R22322 OUT1.n58 OUT1.n54 34.3584
R22323 OUT1.n6 OUT1.n4 34.3584
R22324 OUT1.n8 OUT1.n6 34.3584
R22325 OUT1.n10 OUT1.n8 34.3584
R22326 OUT1.n12 OUT1.n10 34.3584
R22327 OUT1.n14 OUT1.n12 34.3584
R22328 OUT1.n18 OUT1.n14 34.3584
R22329 OUT1.n118 OUT1.t35 26.5955
R22330 OUT1.n118 OUT1.t48 26.5955
R22331 OUT1.n120 OUT1.t33 26.5955
R22332 OUT1.n120 OUT1.t5 26.5955
R22333 OUT1.n121 OUT1.t55 26.5955
R22334 OUT1.n121 OUT1.t21 26.5955
R22335 OUT1.n123 OUT1.t0 26.5955
R22336 OUT1.n123 OUT1.t41 26.5955
R22337 OUT1.n125 OUT1.t11 26.5955
R22338 OUT1.n125 OUT1.t29 26.5955
R22339 OUT1.n127 OUT1.t27 26.5955
R22340 OUT1.n127 OUT1.t44 26.5955
R22341 OUT1.n129 OUT1.t50 26.5955
R22342 OUT1.n129 OUT1.t16 26.5955
R22343 OUT1.n131 OUT1.t61 26.5955
R22344 OUT1.n131 OUT1.t37 26.5955
R22345 OUT1.n99 OUT1.t60 26.5955
R22346 OUT1.n99 OUT1.t25 26.5955
R22347 OUT1.n100 OUT1.t15 26.5955
R22348 OUT1.n100 OUT1.t24 26.5955
R22349 OUT1.n101 OUT1.t31 26.5955
R22350 OUT1.n101 OUT1.t4 26.5955
R22351 OUT1.n103 OUT1.t46 26.5955
R22352 OUT1.n103 OUT1.t18 26.5955
R22353 OUT1.n105 OUT1.t17 26.5955
R22354 OUT1.n105 OUT1.t30 26.5955
R22355 OUT1.n107 OUT1.t38 26.5955
R22356 OUT1.n107 OUT1.t52 26.5955
R22357 OUT1.n109 OUT1.t51 26.5955
R22358 OUT1.n109 OUT1.t6 26.5955
R22359 OUT1.n111 OUT1.t40 26.5955
R22360 OUT1.n111 OUT1.t8 26.5955
R22361 OUT1.n62 OUT1.t2 26.5955
R22362 OUT1.n62 OUT1.t36 26.5955
R22363 OUT1.n63 OUT1.t22 26.5955
R22364 OUT1.n63 OUT1.t34 26.5955
R22365 OUT1.n64 OUT1.t32 26.5955
R22366 OUT1.n64 OUT1.t56 26.5955
R22367 OUT1.n66 OUT1.t53 26.5955
R22368 OUT1.n66 OUT1.t19 26.5955
R22369 OUT1.n68 OUT1.t45 26.5955
R22370 OUT1.n68 OUT1.t12 26.5955
R22371 OUT1.n70 OUT1.t10 26.5955
R22372 OUT1.n70 OUT1.t28 26.5955
R22373 OUT1.n72 OUT1.t26 26.5955
R22374 OUT1.n72 OUT1.t43 26.5955
R22375 OUT1.n74 OUT1.t49 26.5955
R22376 OUT1.n74 OUT1.t62 26.5955
R22377 OUT1.n22 OUT1.t1 26.5955
R22378 OUT1.n22 OUT1.t14 26.5955
R22379 OUT1.n23 OUT1.t20 26.5955
R22380 OUT1.n23 OUT1.t42 26.5955
R22381 OUT1.n24 OUT1.t39 26.5955
R22382 OUT1.n24 OUT1.t54 26.5955
R22383 OUT1.n26 OUT1.t59 26.5955
R22384 OUT1.n26 OUT1.t7 26.5955
R22385 OUT1.n28 OUT1.t13 26.5955
R22386 OUT1.n28 OUT1.t47 26.5955
R22387 OUT1.n30 OUT1.t23 26.5955
R22388 OUT1.n30 OUT1.t58 26.5955
R22389 OUT1.n32 OUT1.t63 26.5955
R22390 OUT1.n32 OUT1.t9 26.5955
R22391 OUT1.n34 OUT1.t57 26.5955
R22392 OUT1.n34 OUT1.t3 26.5955
R22393 OUT1.n149 OUT1.t110 24.9236
R22394 OUT1.n149 OUT1.t123 24.9236
R22395 OUT1.n136 OUT1.t108 24.9236
R22396 OUT1.n136 OUT1.t80 24.9236
R22397 OUT1.n137 OUT1.t66 24.9236
R22398 OUT1.n137 OUT1.t96 24.9236
R22399 OUT1.n139 OUT1.t75 24.9236
R22400 OUT1.n139 OUT1.t116 24.9236
R22401 OUT1.n141 OUT1.t86 24.9236
R22402 OUT1.n141 OUT1.t104 24.9236
R22403 OUT1.n143 OUT1.t102 24.9236
R22404 OUT1.n143 OUT1.t119 24.9236
R22405 OUT1.n145 OUT1.t125 24.9236
R22406 OUT1.n145 OUT1.t91 24.9236
R22407 OUT1.n147 OUT1.t72 24.9236
R22408 OUT1.n147 OUT1.t112 24.9236
R22409 OUT1.n94 OUT1.t71 24.9236
R22410 OUT1.n94 OUT1.t100 24.9236
R22411 OUT1.n81 OUT1.t90 24.9236
R22412 OUT1.n81 OUT1.t99 24.9236
R22413 OUT1.n82 OUT1.t106 24.9236
R22414 OUT1.n82 OUT1.t79 24.9236
R22415 OUT1.n84 OUT1.t121 24.9236
R22416 OUT1.n84 OUT1.t93 24.9236
R22417 OUT1.n86 OUT1.t92 24.9236
R22418 OUT1.n86 OUT1.t105 24.9236
R22419 OUT1.n88 OUT1.t113 24.9236
R22420 OUT1.n88 OUT1.t127 24.9236
R22421 OUT1.n90 OUT1.t126 24.9236
R22422 OUT1.n90 OUT1.t81 24.9236
R22423 OUT1.n92 OUT1.t115 24.9236
R22424 OUT1.n92 OUT1.t83 24.9236
R22425 OUT1.n55 OUT1.t77 24.9236
R22426 OUT1.n55 OUT1.t111 24.9236
R22427 OUT1.n42 OUT1.t97 24.9236
R22428 OUT1.n42 OUT1.t109 24.9236
R22429 OUT1.n43 OUT1.t107 24.9236
R22430 OUT1.n43 OUT1.t67 24.9236
R22431 OUT1.n45 OUT1.t64 24.9236
R22432 OUT1.n45 OUT1.t94 24.9236
R22433 OUT1.n47 OUT1.t120 24.9236
R22434 OUT1.n47 OUT1.t88 24.9236
R22435 OUT1.n49 OUT1.t84 24.9236
R22436 OUT1.n49 OUT1.t103 24.9236
R22437 OUT1.n51 OUT1.t101 24.9236
R22438 OUT1.n51 OUT1.t118 24.9236
R22439 OUT1.n53 OUT1.t124 24.9236
R22440 OUT1.n53 OUT1.t73 24.9236
R22441 OUT1.n15 OUT1.t76 24.9236
R22442 OUT1.n15 OUT1.t89 24.9236
R22443 OUT1.n2 OUT1.t95 24.9236
R22444 OUT1.n2 OUT1.t117 24.9236
R22445 OUT1.n3 OUT1.t114 24.9236
R22446 OUT1.n3 OUT1.t65 24.9236
R22447 OUT1.n5 OUT1.t70 24.9236
R22448 OUT1.n5 OUT1.t82 24.9236
R22449 OUT1.n7 OUT1.t87 24.9236
R22450 OUT1.n7 OUT1.t122 24.9236
R22451 OUT1.n9 OUT1.t98 24.9236
R22452 OUT1.n9 OUT1.t69 24.9236
R22453 OUT1.n11 OUT1.t74 24.9236
R22454 OUT1.n11 OUT1.t85 24.9236
R22455 OUT1.n13 OUT1.t68 24.9236
R22456 OUT1.n13 OUT1.t78 24.9236
R22457 OUT1 OUT1.n150 11.4429
R22458 OUT1 OUT1.n95 11.4429
R22459 OUT1 OUT1.n58 11.4429
R22460 OUT1 OUT1.n18 11.4429
R22461 OUT1.n77 OUT1.n62 8.55024
R22462 OUT1.n37 OUT1.n22 8.55024
R22463 OUT1.n114 OUT1.n99 8.55024
R22464 OUT1.n119 OUT1.n118 8.46262
R22465 OUT1.n56 OUT1.n55 7.77479
R22466 OUT1.n16 OUT1.n15 7.77479
R22467 OUT1.n135 OUT1.n134 4.6505
R22468 OUT1.n151 OUT1 3.29747
R22469 OUT1.n96 OUT1 3.29747
R22470 OUT1.n78 OUT1.n77 3.20821
R22471 OUT1.n38 OUT1.n37 3.2082
R22472 OUT1.n115 OUT1.n114 3.20156
R22473 OUT1.n59 OUT1 3.10353
R22474 OUT1.n19 OUT1 3.10353
R22475 OUT1.n57 OUT1.n41 3.1005
R22476 OUT1.n17 OUT1.n1 3.1005
R22477 OUT1.n134 OUT1.n133 2.71565
R22478 OUT1.n114 OUT1.n113 2.32777
R22479 OUT1.n77 OUT1.n76 2.32777
R22480 OUT1.n37 OUT1.n36 2.32777
R22481 OUT1.n150 OUT1 1.74595
R22482 OUT1.n95 OUT1 1.74595
R22483 OUT1.n157 OUT1.n156 1.07337
R22484 OUT1.n58 OUT1.n57 0.970197
R22485 OUT1.n18 OUT1.n17 0.970197
R22486 OUT1.n158 OUT1.n157 0.69375
R22487 OUT1.n159 OUT1.n158 0.68905
R22488 OUT1.n56 OUT1 0.649449
R22489 OUT1.n16 OUT1 0.649449
R22490 OUT1.n158 OUT1.n79 0.414635
R22491 OUT1.n157 OUT1.n116 0.382465
R22492 OUT1.n159 OUT1.n39 0.368576
R22493 OUT1 OUT1.n159 0.279743
R22494 OUT1.n134 OUT1.n119 0.207197
R22495 OUT1.n79 OUT1.n78 0.157252
R22496 OUT1.n39 OUT1.n38 0.139891
R22497 OUT1.n156 OUT1.n155 0.139389
R22498 OUT1.n116 OUT1.n115 0.132946
R22499 OUT1.n57 OUT1.n56 0.118507
R22500 OUT1.n17 OUT1.n16 0.118507
R22501 OUT1.n60 OUT1.n41 0.111611
R22502 OUT1.n20 OUT1.n1 0.111611
R22503 OUT1.n154 OUT1.n135 0.0991111
R22504 OUT1.n154 OUT1.n152 0.0296667
R22505 OUT1.n135 OUT1.n117 0.0282778
R22506 OUT1.n98 OUT1.n97 0.0227222
R22507 OUT1.n61 OUT1.n60 0.0171667
R22508 OUT1.n21 OUT1.n20 0.0171667
R22509 OUT1.n115 OUT1.n98 0.00100004
R22510 OUT1.n38 OUT1.n21 0.00100004
R22511 OUT1.n78 OUT1.n61 0.00100004
R22512 OUT1.n152 OUT1.n151 0.000513563
R22513 OUT1.n97 OUT1.n96 0.000513563
R22514 OUT1.n60 OUT1.n59 0.000513218
R22515 OUT1.n20 OUT1.n19 0.000513218
R22516 OUT1.n98 OUT1.n80 0.00050517
R22517 OUT1.n154 OUT1.n153 0.000504838
R22518 OUT1.n61 OUT1.n40 0.000504838
R22519 OUT1.n21 OUT1.n0 0.000504838
R22520 OUT1.n155 OUT1.n154 0.000501713
R22521 frontAnalog_v0p0p1_8.RSfetsym_0.QN.n1 frontAnalog_v0p0p1_8.RSfetsym_0.QN.t5 117.511
R22522 frontAnalog_v0p0p1_8.RSfetsym_0.QN.n1 frontAnalog_v0p0p1_8.RSfetsym_0.QN.t6 110.698
R22523 frontAnalog_v0p0p1_8.RSfetsym_0.QN.n4 frontAnalog_v0p0p1_8.RSfetsym_0.QN.t1 19.1963
R22524 frontAnalog_v0p0p1_8.RSfetsym_0.QN.n7 frontAnalog_v0p0p1_8.RSfetsym_0.QN.t4 14.2842
R22525 frontAnalog_v0p0p1_8.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_8.RSfetsym_0.QN.t2 14.283
R22526 frontAnalog_v0p0p1_8.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_8.RSfetsym_0.QN.t3 14.283
R22527 frontAnalog_v0p0p1_8.RSfetsym_0.QN.n11 frontAnalog_v0p0p1_8.RSfetsym_0.QN.t0 9.14075
R22528 frontAnalog_v0p0p1_8.RSfetsym_0.QN.n11 frontAnalog_v0p0p1_8.RSfetsym_0.QN.n10 0.74645
R22529 frontAnalog_v0p0p1_8.RSfetsym_0.QN.n2 frontAnalog_v0p0p1_8.RSfetsym_0.QN.n1 0.688382
R22530 frontAnalog_v0p0p1_8.RSfetsym_0.QN.n10 frontAnalog_v0p0p1_8.RSfetsym_0.QN.n9 0.2402
R22531 frontAnalog_v0p0p1_8.RSfetsym_0.QN.n9 frontAnalog_v0p0p1_8.RSfetsym_0.QN.n8 0.236824
R22532 frontAnalog_v0p0p1_8.RSfetsym_0.QN.n4 frontAnalog_v0p0p1_8.RSfetsym_0.QN.n3 0.132187
R22533 frontAnalog_v0p0p1_8.RSfetsym_0.QN.n9 frontAnalog_v0p0p1_8.RSfetsym_0.QN.n4 0.0968646
R22534 frontAnalog_v0p0p1_8.RSfetsym_0.QN frontAnalog_v0p0p1_8.RSfetsym_0.QN.n11 0.0446535
R22535 frontAnalog_v0p0p1_8.RSfetsym_0.QN.n8 frontAnalog_v0p0p1_8.RSfetsym_0.QN.n6 0.0272538
R22536 frontAnalog_v0p0p1_8.RSfetsym_0.QN.n10 frontAnalog_v0p0p1_8.RSfetsym_0.QN.n0 0.00981499
R22537 frontAnalog_v0p0p1_8.RSfetsym_0.QN.n3 frontAnalog_v0p0p1_8.RSfetsym_0.QN.n2 0.00725433
R22538 frontAnalog_v0p0p1_8.RSfetsym_0.QN.n6 frontAnalog_v0p0p1_8.RSfetsym_0.QN.n5 0.00610579
R22539 frontAnalog_v0p0p1_8.RSfetsym_0.QN.n8 frontAnalog_v0p0p1_8.RSfetsym_0.QN.n7 0.00225341
R22540 resistorDivider_v0p0p1_0.V9.n0 resistorDivider_v0p0p1_0.V9.t17 167.365
R22541 resistorDivider_v0p0p1_0.V9.n0 resistorDivider_v0p0p1_0.V9.t16 92.4496
R22542 resistorDivider_v0p0p1_0.V9.n1 resistorDivider_v0p0p1_0.V9.n0 2.07493
R22543 resistorDivider_v0p0p1_0.V9.n9 resistorDivider_v0p0p1_0.V9.n8 0.141636
R22544 resistorDivider_v0p0p1_0.V9.n8 resistorDivider_v0p0p1_0.V9.n7 0.141636
R22545 resistorDivider_v0p0p1_0.V9.n7 resistorDivider_v0p0p1_0.V9.n6 0.141636
R22546 resistorDivider_v0p0p1_0.V9.n6 resistorDivider_v0p0p1_0.V9.n5 0.141636
R22547 resistorDivider_v0p0p1_0.V9.n5 resistorDivider_v0p0p1_0.V9.n4 0.141636
R22548 resistorDivider_v0p0p1_0.V9.n4 resistorDivider_v0p0p1_0.V9.n3 0.141636
R22549 resistorDivider_v0p0p1_0.V9.n3 resistorDivider_v0p0p1_0.V9.n2 0.141636
R22550 resistorDivider_v0p0p1_0.V9.n1 resistorDivider_v0p0p1_0.V9 0.12425
R22551 resistorDivider_v0p0p1_0.V9 resistorDivider_v0p0p1_0.V9.n9 0.102242
R22552 resistorDivider_v0p0p1_0.V9 resistorDivider_v0p0p1_0.V9.n1 0.0314375
R22553 resistorDivider_v0p0p1_0.V9.n9 resistorDivider_v0p0p1_0.V9.t0 0.00250214
R22554 resistorDivider_v0p0p1_0.V9.n2 resistorDivider_v0p0p1_0.V9.t6 0.000502142
R22555 resistorDivider_v0p0p1_0.V9.n3 resistorDivider_v0p0p1_0.V9.t5 0.000502142
R22556 resistorDivider_v0p0p1_0.V9.n4 resistorDivider_v0p0p1_0.V9.t14 0.000502142
R22557 resistorDivider_v0p0p1_0.V9.n5 resistorDivider_v0p0p1_0.V9.t3 0.000502142
R22558 resistorDivider_v0p0p1_0.V9.n6 resistorDivider_v0p0p1_0.V9.t7 0.000502142
R22559 resistorDivider_v0p0p1_0.V9.n7 resistorDivider_v0p0p1_0.V9.t8 0.000502142
R22560 resistorDivider_v0p0p1_0.V9.n8 resistorDivider_v0p0p1_0.V9.t11 0.000502142
R22561 resistorDivider_v0p0p1_0.V9.n9 resistorDivider_v0p0p1_0.V9.t2 0.000502142
R22562 resistorDivider_v0p0p1_0.V9.n8 resistorDivider_v0p0p1_0.V9.t10 0.000502142
R22563 resistorDivider_v0p0p1_0.V9.n7 resistorDivider_v0p0p1_0.V9.t15 0.000502142
R22564 resistorDivider_v0p0p1_0.V9.n6 resistorDivider_v0p0p1_0.V9.t4 0.000502142
R22565 resistorDivider_v0p0p1_0.V9.n5 resistorDivider_v0p0p1_0.V9.t9 0.000502142
R22566 resistorDivider_v0p0p1_0.V9.n4 resistorDivider_v0p0p1_0.V9.t12 0.000502142
R22567 resistorDivider_v0p0p1_0.V9.n3 resistorDivider_v0p0p1_0.V9.t13 0.000502142
R22568 resistorDivider_v0p0p1_0.V9.n2 resistorDivider_v0p0p1_0.V9.t1 0.000502142
R22569 resistorDivider_v0p0p1_0.V15.n0 resistorDivider_v0p0p1_0.V15.t16 167.365
R22570 resistorDivider_v0p0p1_0.V15.n0 resistorDivider_v0p0p1_0.V15.t17 92.4496
R22571 resistorDivider_v0p0p1_0.V15.n1 resistorDivider_v0p0p1_0.V15.n0 2.07493
R22572 resistorDivider_v0p0p1_0.V15.n9 resistorDivider_v0p0p1_0.V15.n8 0.141636
R22573 resistorDivider_v0p0p1_0.V15.n8 resistorDivider_v0p0p1_0.V15.n7 0.141636
R22574 resistorDivider_v0p0p1_0.V15.n7 resistorDivider_v0p0p1_0.V15.n6 0.141636
R22575 resistorDivider_v0p0p1_0.V15.n6 resistorDivider_v0p0p1_0.V15.n5 0.141636
R22576 resistorDivider_v0p0p1_0.V15.n5 resistorDivider_v0p0p1_0.V15.n4 0.141636
R22577 resistorDivider_v0p0p1_0.V15.n4 resistorDivider_v0p0p1_0.V15.n3 0.141636
R22578 resistorDivider_v0p0p1_0.V15.n3 resistorDivider_v0p0p1_0.V15.n2 0.141636
R22579 resistorDivider_v0p0p1_0.V15.n1 resistorDivider_v0p0p1_0.V15 0.12425
R22580 resistorDivider_v0p0p1_0.V15 resistorDivider_v0p0p1_0.V15.n9 0.100159
R22581 resistorDivider_v0p0p1_0.V15 resistorDivider_v0p0p1_0.V15.n1 0.0358571
R22582 resistorDivider_v0p0p1_0.V15.n5 resistorDivider_v0p0p1_0.V15.t0 0.00250214
R22583 resistorDivider_v0p0p1_0.V15.n2 resistorDivider_v0p0p1_0.V15.t7 0.000502142
R22584 resistorDivider_v0p0p1_0.V15.n3 resistorDivider_v0p0p1_0.V15.t2 0.000502142
R22585 resistorDivider_v0p0p1_0.V15.n4 resistorDivider_v0p0p1_0.V15.t10 0.000502142
R22586 resistorDivider_v0p0p1_0.V15.n6 resistorDivider_v0p0p1_0.V15.t3 0.000502142
R22587 resistorDivider_v0p0p1_0.V15.n7 resistorDivider_v0p0p1_0.V15.t8 0.000502142
R22588 resistorDivider_v0p0p1_0.V15.n8 resistorDivider_v0p0p1_0.V15.t14 0.000502142
R22589 resistorDivider_v0p0p1_0.V15.n9 resistorDivider_v0p0p1_0.V15.t1 0.000502142
R22590 resistorDivider_v0p0p1_0.V15.n9 resistorDivider_v0p0p1_0.V15.t5 0.000502142
R22591 resistorDivider_v0p0p1_0.V15.n8 resistorDivider_v0p0p1_0.V15.t12 0.000502142
R22592 resistorDivider_v0p0p1_0.V15.n7 resistorDivider_v0p0p1_0.V15.t13 0.000502142
R22593 resistorDivider_v0p0p1_0.V15.n6 resistorDivider_v0p0p1_0.V15.t15 0.000502142
R22594 resistorDivider_v0p0p1_0.V15.n5 resistorDivider_v0p0p1_0.V15.t6 0.000502142
R22595 resistorDivider_v0p0p1_0.V15.n4 resistorDivider_v0p0p1_0.V15.t4 0.000502142
R22596 resistorDivider_v0p0p1_0.V15.n3 resistorDivider_v0p0p1_0.V15.t11 0.000502142
R22597 resistorDivider_v0p0p1_0.V15.n2 resistorDivider_v0p0p1_0.V15.t9 0.000502142
R22598 frontAnalog_v0p0p1_2.x63.A.n2 frontAnalog_v0p0p1_2.x63.A.t5 260.322
R22599 frontAnalog_v0p0p1_2.x63.A.n4 frontAnalog_v0p0p1_2.x63.A.t4 233.888
R22600 frontAnalog_v0p0p1_2.x63.A.n2 frontAnalog_v0p0p1_2.x63.A.t6 175.169
R22601 frontAnalog_v0p0p1_2.x63.A.n3 frontAnalog_v0p0p1_2.x63.A.t7 159.725
R22602 frontAnalog_v0p0p1_2.x63.A.n1 frontAnalog_v0p0p1_2.x63.A.t0 17.4109
R22603 frontAnalog_v0p0p1_2.x63.A.n0 frontAnalog_v0p0p1_2.x63.A.n2 9.75129
R22604 frontAnalog_v0p0p1_2.x63.A.n1 frontAnalog_v0p0p1_2.x63.A.t1 9.6027
R22605 frontAnalog_v0p0p1_2.x63.A.n0 frontAnalog_v0p0p1_2.x63.A 2.33338
R22606 frontAnalog_v0p0p1_2.x63.A.n5 frontAnalog_v0p0p1_2.x63.A.t2 8.40929
R22607 frontAnalog_v0p0p1_2.x63.A.n3 frontAnalog_v0p0p1_2.x63.A.t3 8.06629
R22608 frontAnalog_v0p0p1_2.x63.A.n4 frontAnalog_v0p0p1_2.x63.A.n3 1.73501
R22609 frontAnalog_v0p0p1_2.x63.A.n1 frontAnalog_v0p0p1_2.x63.A.n4 0.99025
R22610 frontAnalog_v0p0p1_2.x63.A.n5 frontAnalog_v0p0p1_2.x63.A.n1 0.853186
R22611 frontAnalog_v0p0p1_2.x63.A frontAnalog_v0p0p1_2.x63.A.n0 0.349517
R22612 frontAnalog_v0p0p1_2.x63.A frontAnalog_v0p0p1_2.x63.A.n5 0.24425
R22613 frontAnalog_v0p0p1_2.x65.A.n1 frontAnalog_v0p0p1_2.x65.A.t4 260.322
R22614 frontAnalog_v0p0p1_2.x65.A.n4 frontAnalog_v0p0p1_2.x65.A.t6 233.929
R22615 frontAnalog_v0p0p1_2.x65.A.n1 frontAnalog_v0p0p1_2.x65.A.t5 175.169
R22616 frontAnalog_v0p0p1_2.x65.A.n3 frontAnalog_v0p0p1_2.x65.A.t7 160.416
R22617 frontAnalog_v0p0p1_2.x65.A.n2 frontAnalog_v0p0p1_2.x65.A.t2 17.4109
R22618 frontAnalog_v0p0p1_2.x65.A.n2 frontAnalog_v0p0p1_2.x65.A.t3 10.2053
R22619 frontAnalog_v0p0p1_2.x65.A.n0 frontAnalog_v0p0p1_2.x65.A 2.78715
R22620 frontAnalog_v0p0p1_2.x65.A.n0 frontAnalog_v0p0p1_2.x65.A.n1 9.09103
R22621 frontAnalog_v0p0p1_2.x65.A.n6 frontAnalog_v0p0p1_2.x65.A.t1 7.94569
R22622 frontAnalog_v0p0p1_2.x65.A.n3 frontAnalog_v0p0p1_2.x65.A.t0 7.55846
R22623 frontAnalog_v0p0p1_2.x65.A.n5 frontAnalog_v0p0p1_2.x65.A.n4 1.4614
R22624 frontAnalog_v0p0p1_2.x65.A.n4 frontAnalog_v0p0p1_2.x65.A.n3 1.19626
R22625 frontAnalog_v0p0p1_2.x65.A.n6 frontAnalog_v0p0p1_2.x65.A.n5 0.836961
R22626 frontAnalog_v0p0p1_2.x65.A frontAnalog_v0p0p1_2.x65.A.n0 0.390342
R22627 frontAnalog_v0p0p1_2.x65.A.n5 frontAnalog_v0p0p1_2.x65.A.n2 0.154668
R22628 frontAnalog_v0p0p1_2.x65.A frontAnalog_v0p0p1_2.x65.A.n6 0.08175
R22629 frontAnalog_v0p0p1_15.RSfetsym_0.QN.n1 frontAnalog_v0p0p1_15.RSfetsym_0.QN.t6 117.511
R22630 frontAnalog_v0p0p1_15.RSfetsym_0.QN.n1 frontAnalog_v0p0p1_15.RSfetsym_0.QN.t5 110.698
R22631 frontAnalog_v0p0p1_15.RSfetsym_0.QN.n4 frontAnalog_v0p0p1_15.RSfetsym_0.QN.t4 19.1963
R22632 frontAnalog_v0p0p1_15.RSfetsym_0.QN.n7 frontAnalog_v0p0p1_15.RSfetsym_0.QN.t0 14.2842
R22633 frontAnalog_v0p0p1_15.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_15.RSfetsym_0.QN.t3 14.283
R22634 frontAnalog_v0p0p1_15.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_15.RSfetsym_0.QN.t2 14.283
R22635 frontAnalog_v0p0p1_15.RSfetsym_0.QN.n11 frontAnalog_v0p0p1_15.RSfetsym_0.QN.t1 9.14075
R22636 frontAnalog_v0p0p1_15.RSfetsym_0.QN.n11 frontAnalog_v0p0p1_15.RSfetsym_0.QN.n10 0.74645
R22637 frontAnalog_v0p0p1_15.RSfetsym_0.QN.n2 frontAnalog_v0p0p1_15.RSfetsym_0.QN.n1 0.688382
R22638 frontAnalog_v0p0p1_15.RSfetsym_0.QN.n10 frontAnalog_v0p0p1_15.RSfetsym_0.QN.n9 0.2402
R22639 frontAnalog_v0p0p1_15.RSfetsym_0.QN.n9 frontAnalog_v0p0p1_15.RSfetsym_0.QN.n8 0.236824
R22640 frontAnalog_v0p0p1_15.RSfetsym_0.QN.n4 frontAnalog_v0p0p1_15.RSfetsym_0.QN.n3 0.132187
R22641 frontAnalog_v0p0p1_15.RSfetsym_0.QN.n9 frontAnalog_v0p0p1_15.RSfetsym_0.QN.n4 0.0968646
R22642 frontAnalog_v0p0p1_15.RSfetsym_0.QN frontAnalog_v0p0p1_15.RSfetsym_0.QN.n11 0.0446535
R22643 frontAnalog_v0p0p1_15.RSfetsym_0.QN.n8 frontAnalog_v0p0p1_15.RSfetsym_0.QN.n6 0.0272538
R22644 frontAnalog_v0p0p1_15.RSfetsym_0.QN.n10 frontAnalog_v0p0p1_15.RSfetsym_0.QN.n0 0.00981499
R22645 frontAnalog_v0p0p1_15.RSfetsym_0.QN.n3 frontAnalog_v0p0p1_15.RSfetsym_0.QN.n2 0.00725433
R22646 frontAnalog_v0p0p1_15.RSfetsym_0.QN.n6 frontAnalog_v0p0p1_15.RSfetsym_0.QN.n5 0.00610579
R22647 frontAnalog_v0p0p1_15.RSfetsym_0.QN.n8 frontAnalog_v0p0p1_15.RSfetsym_0.QN.n7 0.00225341
R22648 frontAnalog_v0p0p1_6.Q.n14 frontAnalog_v0p0p1_6.Q.t12 323.342
R22649 frontAnalog_v0p0p1_6.Q.n8 frontAnalog_v0p0p1_6.Q.t11 228.927
R22650 frontAnalog_v0p0p1_6.Q.n11 frontAnalog_v0p0p1_6.Q.t6 196.549
R22651 frontAnalog_v0p0p1_6.Q.n14 frontAnalog_v0p0p1_6.Q.t10 194.809
R22652 frontAnalog_v0p0p1_6.Q.n8 frontAnalog_v0p0p1_6.Q.t8 159.391
R22653 frontAnalog_v0p0p1_6.Q.n11 frontAnalog_v0p0p1_6.Q.t9 148.35
R22654 frontAnalog_v0p0p1_6.Q.n0 frontAnalog_v0p0p1_6.Q.t7 117.314
R22655 frontAnalog_v0p0p1_6.Q.n0 frontAnalog_v0p0p1_6.Q.t5 110.852
R22656 frontAnalog_v0p0p1_6.Q.n15 frontAnalog_v0p0p1_6.Q.n14 76.0005
R22657 frontAnalog_v0p0p1_6.Q.n12 frontAnalog_v0p0p1_6.Q.n11 76.0005
R22658 frontAnalog_v0p0p1_6.Q.n16 frontAnalog_v0p0p1_6.Q.n15 29.3651
R22659 frontAnalog_v0p0p1_6.Q.n1 frontAnalog_v0p0p1_6.Q.t0 17.6181
R22660 frontAnalog_v0p0p1_6.Q.n3 frontAnalog_v0p0p1_6.Q.t3 14.2865
R22661 frontAnalog_v0p0p1_6.Q.n5 frontAnalog_v0p0p1_6.Q.t1 14.283
R22662 frontAnalog_v0p0p1_6.Q.n5 frontAnalog_v0p0p1_6.Q.t2 14.283
R22663 frontAnalog_v0p0p1_6.Q.n13 frontAnalog_v0p0p1_6.Q 9.11
R22664 frontAnalog_v0p0p1_6.Q.n7 frontAnalog_v0p0p1_6.Q.t4 8.77592
R22665 frontAnalog_v0p0p1_6.Q.n9 frontAnalog_v0p0p1_6.Q.n8 8.6846
R22666 frontAnalog_v0p0p1_6.Q.n12 frontAnalog_v0p0p1_6.Q 5.78114
R22667 frontAnalog_v0p0p1_6.Q.n10 frontAnalog_v0p0p1_6.Q.n9 4.26809
R22668 frontAnalog_v0p0p1_6.Q.n18 frontAnalog_v0p0p1_6.Q.n17 3.72735
R22669 frontAnalog_v0p0p1_6.Q frontAnalog_v0p0p1_6.Q.n12 3.71663
R22670 frontAnalog_v0p0p1_6.Q.n9 frontAnalog_v0p0p1_6.Q 1.99652
R22671 frontAnalog_v0p0p1_6.Q.n15 frontAnalog_v0p0p1_6.Q 1.92927
R22672 frontAnalog_v0p0p1_6.Q.n16 frontAnalog_v0p0p1_6.Q.n13 1.69246
R22673 frontAnalog_v0p0p1_6.Q.n7 frontAnalog_v0p0p1_6.Q.n6 1.20426
R22674 frontAnalog_v0p0p1_6.Q.n13 frontAnalog_v0p0p1_6.Q.n10 0.570143
R22675 frontAnalog_v0p0p1_6.Q.n18 frontAnalog_v0p0p1_6.Q.n7 0.336084
R22676 frontAnalog_v0p0p1_6.Q.n4 frontAnalog_v0p0p1_6.Q.n3 0.300242
R22677 frontAnalog_v0p0p1_6.Q.n17 frontAnalog_v0p0p1_6.Q.n16 0.224535
R22678 frontAnalog_v0p0p1_6.Q.n10 frontAnalog_v0p0p1_6.Q 0.221483
R22679 frontAnalog_v0p0p1_6.Q.n17 frontAnalog_v0p0p1_6.Q 0.2005
R22680 frontAnalog_v0p0p1_6.Q.n2 frontAnalog_v0p0p1_6.Q.n0 0.159555
R22681 frontAnalog_v0p0p1_6.Q.n6 frontAnalog_v0p0p1_6.Q.n5 0.106617
R22682 frontAnalog_v0p0p1_6.Q.n4 frontAnalog_v0p0p1_6.Q.n2 0.0796167
R22683 frontAnalog_v0p0p1_6.Q.n6 frontAnalog_v0p0p1_6.Q.n4 0.0480595
R22684 frontAnalog_v0p0p1_6.Q frontAnalog_v0p0p1_6.Q.n18 0.00658123
R22685 frontAnalog_v0p0p1_6.Q.n2 frontAnalog_v0p0p1_6.Q.n1 0.000504658
R22686 frontAnalog_v0p0p1_6.RSfetsym_0.QN.n1 frontAnalog_v0p0p1_6.RSfetsym_0.QN.t6 117.511
R22687 frontAnalog_v0p0p1_6.RSfetsym_0.QN.n1 frontAnalog_v0p0p1_6.RSfetsym_0.QN.t5 110.698
R22688 frontAnalog_v0p0p1_6.RSfetsym_0.QN.n4 frontAnalog_v0p0p1_6.RSfetsym_0.QN.t0 19.1963
R22689 frontAnalog_v0p0p1_6.RSfetsym_0.QN.n7 frontAnalog_v0p0p1_6.RSfetsym_0.QN.t3 14.2842
R22690 frontAnalog_v0p0p1_6.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_6.RSfetsym_0.QN.t1 14.283
R22691 frontAnalog_v0p0p1_6.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_6.RSfetsym_0.QN.t2 14.283
R22692 frontAnalog_v0p0p1_6.RSfetsym_0.QN.n11 frontAnalog_v0p0p1_6.RSfetsym_0.QN.t4 9.14075
R22693 frontAnalog_v0p0p1_6.RSfetsym_0.QN.n11 frontAnalog_v0p0p1_6.RSfetsym_0.QN.n10 0.74645
R22694 frontAnalog_v0p0p1_6.RSfetsym_0.QN.n2 frontAnalog_v0p0p1_6.RSfetsym_0.QN.n1 0.688382
R22695 frontAnalog_v0p0p1_6.RSfetsym_0.QN.n10 frontAnalog_v0p0p1_6.RSfetsym_0.QN.n9 0.2402
R22696 frontAnalog_v0p0p1_6.RSfetsym_0.QN.n9 frontAnalog_v0p0p1_6.RSfetsym_0.QN.n8 0.236824
R22697 frontAnalog_v0p0p1_6.RSfetsym_0.QN.n4 frontAnalog_v0p0p1_6.RSfetsym_0.QN.n3 0.132187
R22698 frontAnalog_v0p0p1_6.RSfetsym_0.QN.n9 frontAnalog_v0p0p1_6.RSfetsym_0.QN.n4 0.0968646
R22699 frontAnalog_v0p0p1_6.RSfetsym_0.QN frontAnalog_v0p0p1_6.RSfetsym_0.QN.n11 0.0446535
R22700 frontAnalog_v0p0p1_6.RSfetsym_0.QN.n8 frontAnalog_v0p0p1_6.RSfetsym_0.QN.n6 0.0272538
R22701 frontAnalog_v0p0p1_6.RSfetsym_0.QN.n10 frontAnalog_v0p0p1_6.RSfetsym_0.QN.n0 0.00981499
R22702 frontAnalog_v0p0p1_6.RSfetsym_0.QN.n3 frontAnalog_v0p0p1_6.RSfetsym_0.QN.n2 0.00725433
R22703 frontAnalog_v0p0p1_6.RSfetsym_0.QN.n6 frontAnalog_v0p0p1_6.RSfetsym_0.QN.n5 0.00610579
R22704 frontAnalog_v0p0p1_6.RSfetsym_0.QN.n8 frontAnalog_v0p0p1_6.RSfetsym_0.QN.n7 0.00225341
R22705 16to4_PriorityEncoder_v0p0p1_0.I13.t9 16to4_PriorityEncoder_v0p0p1_0.I13.t13 618.109
R22706 16to4_PriorityEncoder_v0p0p1_0.I13.n20 16to4_PriorityEncoder_v0p0p1_0.I13.t14 259.74
R22707 16to4_PriorityEncoder_v0p0p1_0.I13 16to4_PriorityEncoder_v0p0p1_0.I13.t9 253.56
R22708 16to4_PriorityEncoder_v0p0p1_0.I13.n8 16to4_PriorityEncoder_v0p0p1_0.I13.t11 228.899
R22709 16to4_PriorityEncoder_v0p0p1_0.I13.n27 16to4_PriorityEncoder_v0p0p1_0.I13.t6 180.286
R22710 16to4_PriorityEncoder_v0p0p1_0.I13.n8 16to4_PriorityEncoder_v0p0p1_0.I13.t10 159.411
R22711 16to4_PriorityEncoder_v0p0p1_0.I13.n20 16to4_PriorityEncoder_v0p0p1_0.I13.t8 157.083
R22712 16to4_PriorityEncoder_v0p0p1_0.I13.n0 16to4_PriorityEncoder_v0p0p1_0.I13.t5 117.314
R22713 16to4_PriorityEncoder_v0p0p1_0.I13.n28 16to4_PriorityEncoder_v0p0p1_0.I13.t7 111.091
R22714 16to4_PriorityEncoder_v0p0p1_0.I13.n0 16to4_PriorityEncoder_v0p0p1_0.I13.t12 110.852
R22715 16to4_PriorityEncoder_v0p0p1_0.I13.n31 16to4_PriorityEncoder_v0p0p1_0.I13 37.7071
R22716 16to4_PriorityEncoder_v0p0p1_0.I13.n1 16to4_PriorityEncoder_v0p0p1_0.I13.t2 17.6181
R22717 16to4_PriorityEncoder_v0p0p1_0.I13.n3 16to4_PriorityEncoder_v0p0p1_0.I13.t4 14.2865
R22718 16to4_PriorityEncoder_v0p0p1_0.I13.n5 16to4_PriorityEncoder_v0p0p1_0.I13.t0 14.283
R22719 16to4_PriorityEncoder_v0p0p1_0.I13.n5 16to4_PriorityEncoder_v0p0p1_0.I13.t1 14.283
R22720 16to4_PriorityEncoder_v0p0p1_0.I13.n29 16to4_PriorityEncoder_v0p0p1_0.I13.n28 9.3005
R22721 16to4_PriorityEncoder_v0p0p1_0.I13 16to4_PriorityEncoder_v0p0p1_0.I13.n19 9.3005
R22722 16to4_PriorityEncoder_v0p0p1_0.I13.n7 16to4_PriorityEncoder_v0p0p1_0.I13.t3 8.77592
R22723 16to4_PriorityEncoder_v0p0p1_0.I13.n30 16to4_PriorityEncoder_v0p0p1_0.I13.n29 7.80966
R22724 16to4_PriorityEncoder_v0p0p1_0.I13.n21 16to4_PriorityEncoder_v0p0p1_0.I13.n20 7.57248
R22725 16to4_PriorityEncoder_v0p0p1_0.I13.n9 16to4_PriorityEncoder_v0p0p1_0.I13.n8 7.36885
R22726 16to4_PriorityEncoder_v0p0p1_0.I13.n34 16to4_PriorityEncoder_v0p0p1_0.I13.n33 6.59722
R22727 16to4_PriorityEncoder_v0p0p1_0.I13.n28 16to4_PriorityEncoder_v0p0p1_0.I13.n27 6.53562
R22728 16to4_PriorityEncoder_v0p0p1_0.I13.n21 16to4_PriorityEncoder_v0p0p1_0.I13 4.8645
R22729 16to4_PriorityEncoder_v0p0p1_0.I13.n11 16to4_PriorityEncoder_v0p0p1_0.I13.n10 3.46717
R22730 16to4_PriorityEncoder_v0p0p1_0.I13.n12 16to4_PriorityEncoder_v0p0p1_0.I13.n11 3.03286
R22731 16to4_PriorityEncoder_v0p0p1_0.I13.n26 16to4_PriorityEncoder_v0p0p1_0.I13.n25 2.32777
R22732 16to4_PriorityEncoder_v0p0p1_0.I13.n30 16to4_PriorityEncoder_v0p0p1_0.I13.n24 2.19001
R22733 16to4_PriorityEncoder_v0p0p1_0.I13.n25 16to4_PriorityEncoder_v0p0p1_0.I13 1.4966
R22734 16to4_PriorityEncoder_v0p0p1_0.I13.n7 16to4_PriorityEncoder_v0p0p1_0.I13.n6 1.20426
R22735 16to4_PriorityEncoder_v0p0p1_0.I13.n32 16to4_PriorityEncoder_v0p0p1_0.I13.n17 1.16836
R22736 16to4_PriorityEncoder_v0p0p1_0.I13.n31 16to4_PriorityEncoder_v0p0p1_0.I13.n30 1.07639
R22737 16to4_PriorityEncoder_v0p0p1_0.I13.n11 16to4_PriorityEncoder_v0p0p1_0.I13.n9 1.06717
R22738 16to4_PriorityEncoder_v0p0p1_0.I13.n10 16to4_PriorityEncoder_v0p0p1_0.I13 1.06717
R22739 16to4_PriorityEncoder_v0p0p1_0.I13.n17 16to4_PriorityEncoder_v0p0p1_0.I13.n16 0.71595
R22740 16to4_PriorityEncoder_v0p0p1_0.I13.n29 16to4_PriorityEncoder_v0p0p1_0.I13.n26 0.499201
R22741 16to4_PriorityEncoder_v0p0p1_0.I13.n33 16to4_PriorityEncoder_v0p0p1_0.I13.n32 0.458555
R22742 16to4_PriorityEncoder_v0p0p1_0.I13.n34 16to4_PriorityEncoder_v0p0p1_0.I13.n7 0.336084
R22743 16to4_PriorityEncoder_v0p0p1_0.I13.n4 16to4_PriorityEncoder_v0p0p1_0.I13.n3 0.300242
R22744 16to4_PriorityEncoder_v0p0p1_0.I13.n17 16to4_PriorityEncoder_v0p0p1_0.I13 0.221483
R22745 16to4_PriorityEncoder_v0p0p1_0.I13.n33 16to4_PriorityEncoder_v0p0p1_0.I13 0.2005
R22746 16to4_PriorityEncoder_v0p0p1_0.I13.n32 16to4_PriorityEncoder_v0p0p1_0.I13.n31 0.192464
R22747 16to4_PriorityEncoder_v0p0p1_0.I13.n2 16to4_PriorityEncoder_v0p0p1_0.I13.n0 0.159555
R22748 16to4_PriorityEncoder_v0p0p1_0.I13.n6 16to4_PriorityEncoder_v0p0p1_0.I13.n5 0.106617
R22749 16to4_PriorityEncoder_v0p0p1_0.I13.n4 16to4_PriorityEncoder_v0p0p1_0.I13.n2 0.0796167
R22750 16to4_PriorityEncoder_v0p0p1_0.I13.n6 16to4_PriorityEncoder_v0p0p1_0.I13.n4 0.0480595
R22751 16to4_PriorityEncoder_v0p0p1_0.I13.n19 16to4_PriorityEncoder_v0p0p1_0.I13.n18 0.0301875
R22752 16to4_PriorityEncoder_v0p0p1_0.I13.n24 16to4_PriorityEncoder_v0p0p1_0.I13.n23 0.0205312
R22753 16to4_PriorityEncoder_v0p0p1_0.I13 16to4_PriorityEncoder_v0p0p1_0.I13.n34 0.00658123
R22754 16to4_PriorityEncoder_v0p0p1_0.I13.n14 16to4_PriorityEncoder_v0p0p1_0.I13.n13 0.00618182
R22755 16to4_PriorityEncoder_v0p0p1_0.I13.n13 16to4_PriorityEncoder_v0p0p1_0.I13.n12 0.00555107
R22756 16to4_PriorityEncoder_v0p0p1_0.I13.n15 16to4_PriorityEncoder_v0p0p1_0.I13.n14 0.00430477
R22757 16to4_PriorityEncoder_v0p0p1_0.I13.n23 16to4_PriorityEncoder_v0p0p1_0.I13.n22 0.00210765
R22758 16to4_PriorityEncoder_v0p0p1_0.I13.n22 16to4_PriorityEncoder_v0p0p1_0.I13.n21 0.00133438
R22759 16to4_PriorityEncoder_v0p0p1_0.I13.n16 16to4_PriorityEncoder_v0p0p1_0.I13.n15 0.00101192
R22760 16to4_PriorityEncoder_v0p0p1_0.I13.n22 16to4_PriorityEncoder_v0p0p1_0.I13.n18 0.00100001
R22761 16to4_PriorityEncoder_v0p0p1_0.I13.n2 16to4_PriorityEncoder_v0p0p1_0.I13.n1 0.000504658
R22762 frontAnalog_v0p0p1_10.IB.n0 frontAnalog_v0p0p1_10.IB.t0 182.794
R22763 frontAnalog_v0p0p1_10.IB.n1 frontAnalog_v0p0p1_10.IB.t12 91.7714
R22764 frontAnalog_v0p0p1_10.IB.n17 frontAnalog_v0p0p1_10.IB.t17 91.7714
R22765 frontAnalog_v0p0p1_10.IB.n16 frontAnalog_v0p0p1_10.IB.t14 91.7714
R22766 frontAnalog_v0p0p1_10.IB.n15 frontAnalog_v0p0p1_10.IB.t27 91.7714
R22767 frontAnalog_v0p0p1_10.IB.n14 frontAnalog_v0p0p1_10.IB.t21 91.7714
R22768 frontAnalog_v0p0p1_10.IB.n13 frontAnalog_v0p0p1_10.IB.t4 91.7714
R22769 frontAnalog_v0p0p1_10.IB.n12 frontAnalog_v0p0p1_10.IB.t31 91.7714
R22770 frontAnalog_v0p0p1_10.IB.n11 frontAnalog_v0p0p1_10.IB.t10 91.7714
R22771 frontAnalog_v0p0p1_10.IB.n10 frontAnalog_v0p0p1_10.IB.t7 91.7714
R22772 frontAnalog_v0p0p1_10.IB.n9 frontAnalog_v0p0p1_10.IB.t18 91.7714
R22773 frontAnalog_v0p0p1_10.IB.n8 frontAnalog_v0p0p1_10.IB.t15 91.7714
R22774 frontAnalog_v0p0p1_10.IB.n7 frontAnalog_v0p0p1_10.IB.t26 91.7714
R22775 frontAnalog_v0p0p1_10.IB.n6 frontAnalog_v0p0p1_10.IB.t22 91.7714
R22776 frontAnalog_v0p0p1_10.IB.n5 frontAnalog_v0p0p1_10.IB.t5 91.7714
R22777 frontAnalog_v0p0p1_10.IB.n4 frontAnalog_v0p0p1_10.IB.t32 91.7714
R22778 frontAnalog_v0p0p1_10.IB.n2 frontAnalog_v0p0p1_10.IB.t3 91.7714
R22779 frontAnalog_v0p0p1_10.IB.n17 frontAnalog_v0p0p1_10.IB.t28 91.3136
R22780 frontAnalog_v0p0p1_10.IB.n16 frontAnalog_v0p0p1_10.IB.t24 91.3136
R22781 frontAnalog_v0p0p1_10.IB.n15 frontAnalog_v0p0p1_10.IB.t6 91.3136
R22782 frontAnalog_v0p0p1_10.IB.n14 frontAnalog_v0p0p1_10.IB.t33 91.3136
R22783 frontAnalog_v0p0p1_10.IB.n13 frontAnalog_v0p0p1_10.IB.t13 91.3136
R22784 frontAnalog_v0p0p1_10.IB.n12 frontAnalog_v0p0p1_10.IB.t8 91.3136
R22785 frontAnalog_v0p0p1_10.IB.n11 frontAnalog_v0p0p1_10.IB.t20 91.3136
R22786 frontAnalog_v0p0p1_10.IB.n10 frontAnalog_v0p0p1_10.IB.t16 91.3136
R22787 frontAnalog_v0p0p1_10.IB.n9 frontAnalog_v0p0p1_10.IB.t30 91.3136
R22788 frontAnalog_v0p0p1_10.IB.n8 frontAnalog_v0p0p1_10.IB.t25 91.3136
R22789 frontAnalog_v0p0p1_10.IB.n7 frontAnalog_v0p0p1_10.IB.t19 91.3136
R22790 frontAnalog_v0p0p1_10.IB.n6 frontAnalog_v0p0p1_10.IB.t34 91.3136
R22791 frontAnalog_v0p0p1_10.IB.n5 frontAnalog_v0p0p1_10.IB.t29 91.3136
R22792 frontAnalog_v0p0p1_10.IB.n4 frontAnalog_v0p0p1_10.IB.t9 91.3136
R22793 frontAnalog_v0p0p1_10.IB.n2 frontAnalog_v0p0p1_10.IB.t11 91.3136
R22794 frontAnalog_v0p0p1_10.IB.n1 frontAnalog_v0p0p1_10.IB.t23 91.3136
R22795 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_10.IB.n17 45.9747
R22796 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_10.IB.n16 45.9747
R22797 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_10.IB.n15 45.9747
R22798 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_10.IB.n14 45.9747
R22799 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_10.IB.n13 45.9747
R22800 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_10.IB.n12 45.9747
R22801 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_10.IB.n11 45.9747
R22802 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_10.IB.n10 45.9747
R22803 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_10.IB.n9 45.9747
R22804 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_10.IB.n8 45.9747
R22805 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_10.IB.n7 45.9747
R22806 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_10.IB.n6 45.9747
R22807 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_10.IB.n5 45.9747
R22808 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_10.IB.n4 45.9747
R22809 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_10.IB.n2 45.9747
R22810 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_10.IB.n1 45.973
R22811 frontAnalog_v0p0p1_10.IB.n34 frontAnalog_v0p0p1_10.IB.t2 5.91044
R22812 frontAnalog_v0p0p1_10.IB.n32 frontAnalog_v0p0p1_10.IB.t1 4.35136
R22813 frontAnalog_v0p0p1_10.IB.n18 frontAnalog_v0p0p1_10.IB 1.53808
R22814 frontAnalog_v0p0p1_10.IB.n34 frontAnalog_v0p0p1_10.IB.n31 1.41054
R22815 frontAnalog_v0p0p1_10.IB.n3 frontAnalog_v0p0p1_10.IB 1.28321
R22816 frontAnalog_v0p0p1_10.IB.n29 frontAnalog_v0p0p1_10.IB 1.15021
R22817 frontAnalog_v0p0p1_10.IB.n28 frontAnalog_v0p0p1_10.IB 1.14904
R22818 frontAnalog_v0p0p1_10.IB.n26 frontAnalog_v0p0p1_10.IB 1.14883
R22819 frontAnalog_v0p0p1_10.IB.n30 frontAnalog_v0p0p1_10.IB 1.14802
R22820 frontAnalog_v0p0p1_10.IB.n19 frontAnalog_v0p0p1_10.IB 1.14536
R22821 frontAnalog_v0p0p1_10.IB.n25 frontAnalog_v0p0p1_10.IB 1.14495
R22822 frontAnalog_v0p0p1_10.IB.n27 frontAnalog_v0p0p1_10.IB 1.14447
R22823 frontAnalog_v0p0p1_10.IB.n21 frontAnalog_v0p0p1_10.IB 1.14439
R22824 frontAnalog_v0p0p1_10.IB.n22 frontAnalog_v0p0p1_10.IB 1.14419
R22825 frontAnalog_v0p0p1_10.IB.n24 frontAnalog_v0p0p1_10.IB 1.14189
R22826 frontAnalog_v0p0p1_10.IB.n23 frontAnalog_v0p0p1_10.IB 1.14114
R22827 frontAnalog_v0p0p1_10.IB.n18 frontAnalog_v0p0p1_10.IB 1.13988
R22828 frontAnalog_v0p0p1_10.IB.n20 frontAnalog_v0p0p1_10.IB 1.13929
R22829 frontAnalog_v0p0p1_10.IB.n3 frontAnalog_v0p0p1_10.IB 0.957022
R22830 frontAnalog_v0p0p1_10.IB.n33 frontAnalog_v0p0p1_10.IB.n32 0.807781
R22831 frontAnalog_v0p0p1_10.IB.n34 frontAnalog_v0p0p1_10.IB.n0 0.504831
R22832 frontAnalog_v0p0p1_10.IB.n30 frontAnalog_v0p0p1_10.IB.n29 0.399765
R22833 frontAnalog_v0p0p1_10.IB.n28 frontAnalog_v0p0p1_10.IB.n27 0.399029
R22834 frontAnalog_v0p0p1_10.IB.n25 frontAnalog_v0p0p1_10.IB.n24 0.399029
R22835 frontAnalog_v0p0p1_10.IB.n23 frontAnalog_v0p0p1_10.IB.n22 0.398294
R22836 frontAnalog_v0p0p1_10.IB.n21 frontAnalog_v0p0p1_10.IB.n20 0.398294
R22837 frontAnalog_v0p0p1_10.IB.n26 frontAnalog_v0p0p1_10.IB.n25 0.397559
R22838 frontAnalog_v0p0p1_10.IB.n22 frontAnalog_v0p0p1_10.IB.n21 0.396824
R22839 frontAnalog_v0p0p1_10.IB.n20 frontAnalog_v0p0p1_10.IB.n19 0.396824
R22840 frontAnalog_v0p0p1_10.IB.n19 frontAnalog_v0p0p1_10.IB.n18 0.396824
R22841 frontAnalog_v0p0p1_10.IB.n27 frontAnalog_v0p0p1_10.IB.n26 0.396088
R22842 frontAnalog_v0p0p1_10.IB.n24 frontAnalog_v0p0p1_10.IB.n23 0.396088
R22843 frontAnalog_v0p0p1_10.IB.n29 frontAnalog_v0p0p1_10.IB.n28 0.395353
R22844 frontAnalog_v0p0p1_10.IB.n31 frontAnalog_v0p0p1_10.IB.n30 0.249029
R22845 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_10.IB.n34 0.168769
R22846 frontAnalog_v0p0p1_10.IB.n31 frontAnalog_v0p0p1_10.IB.n3 0.151971
R22847 frontAnalog_v0p0p1_10.IB.n0 frontAnalog_v0p0p1_10.IB.n33 0.0762967
R22848 resistorDivider_v0p0p1_0.V14.n0 resistorDivider_v0p0p1_0.V14.t17 167.365
R22849 resistorDivider_v0p0p1_0.V14.n0 resistorDivider_v0p0p1_0.V14.t16 92.4496
R22850 resistorDivider_v0p0p1_0.V14.n1 resistorDivider_v0p0p1_0.V14.n0 2.07493
R22851 resistorDivider_v0p0p1_0.V14.n9 resistorDivider_v0p0p1_0.V14.n8 0.141636
R22852 resistorDivider_v0p0p1_0.V14.n8 resistorDivider_v0p0p1_0.V14.n7 0.141636
R22853 resistorDivider_v0p0p1_0.V14.n7 resistorDivider_v0p0p1_0.V14.n6 0.141636
R22854 resistorDivider_v0p0p1_0.V14.n6 resistorDivider_v0p0p1_0.V14.n5 0.141636
R22855 resistorDivider_v0p0p1_0.V14.n5 resistorDivider_v0p0p1_0.V14.n4 0.141636
R22856 resistorDivider_v0p0p1_0.V14.n4 resistorDivider_v0p0p1_0.V14.n3 0.141636
R22857 resistorDivider_v0p0p1_0.V14.n3 resistorDivider_v0p0p1_0.V14.n2 0.141636
R22858 resistorDivider_v0p0p1_0.V14.n1 resistorDivider_v0p0p1_0.V14 0.12425
R22859 resistorDivider_v0p0p1_0.V14 resistorDivider_v0p0p1_0.V14.n9 0.102242
R22860 resistorDivider_v0p0p1_0.V14 resistorDivider_v0p0p1_0.V14.n1 0.0358571
R22861 resistorDivider_v0p0p1_0.V14.n2 resistorDivider_v0p0p1_0.V14.t0 0.00250214
R22862 resistorDivider_v0p0p1_0.V14.n3 resistorDivider_v0p0p1_0.V14.t13 0.000502142
R22863 resistorDivider_v0p0p1_0.V14.n4 resistorDivider_v0p0p1_0.V14.t7 0.000502142
R22864 resistorDivider_v0p0p1_0.V14.n5 resistorDivider_v0p0p1_0.V14.t10 0.000502142
R22865 resistorDivider_v0p0p1_0.V14.n6 resistorDivider_v0p0p1_0.V14.t5 0.000502142
R22866 resistorDivider_v0p0p1_0.V14.n7 resistorDivider_v0p0p1_0.V14.t8 0.000502142
R22867 resistorDivider_v0p0p1_0.V14.n8 resistorDivider_v0p0p1_0.V14.t11 0.000502142
R22868 resistorDivider_v0p0p1_0.V14.n9 resistorDivider_v0p0p1_0.V14.t15 0.000502142
R22869 resistorDivider_v0p0p1_0.V14.n9 resistorDivider_v0p0p1_0.V14.t2 0.000502142
R22870 resistorDivider_v0p0p1_0.V14.n8 resistorDivider_v0p0p1_0.V14.t14 0.000502142
R22871 resistorDivider_v0p0p1_0.V14.n7 resistorDivider_v0p0p1_0.V14.t9 0.000502142
R22872 resistorDivider_v0p0p1_0.V14.n6 resistorDivider_v0p0p1_0.V14.t4 0.000502142
R22873 resistorDivider_v0p0p1_0.V14.n5 resistorDivider_v0p0p1_0.V14.t1 0.000502142
R22874 resistorDivider_v0p0p1_0.V14.n4 resistorDivider_v0p0p1_0.V14.t12 0.000502142
R22875 resistorDivider_v0p0p1_0.V14.n3 resistorDivider_v0p0p1_0.V14.t3 0.000502142
R22876 resistorDivider_v0p0p1_0.V14.n2 resistorDivider_v0p0p1_0.V14.t6 0.000502142
R22877 resistorDivider_v0p0p1_0.V13.n0 resistorDivider_v0p0p1_0.V13.t16 167.365
R22878 resistorDivider_v0p0p1_0.V13.n0 resistorDivider_v0p0p1_0.V13.t17 92.4496
R22879 resistorDivider_v0p0p1_0.V13.n1 resistorDivider_v0p0p1_0.V13.n0 2.07493
R22880 resistorDivider_v0p0p1_0.V13.n9 resistorDivider_v0p0p1_0.V13.n8 0.141636
R22881 resistorDivider_v0p0p1_0.V13.n8 resistorDivider_v0p0p1_0.V13.n7 0.141636
R22882 resistorDivider_v0p0p1_0.V13.n7 resistorDivider_v0p0p1_0.V13.n6 0.141636
R22883 resistorDivider_v0p0p1_0.V13.n6 resistorDivider_v0p0p1_0.V13.n5 0.141636
R22884 resistorDivider_v0p0p1_0.V13.n5 resistorDivider_v0p0p1_0.V13.n4 0.141636
R22885 resistorDivider_v0p0p1_0.V13.n4 resistorDivider_v0p0p1_0.V13.n3 0.141636
R22886 resistorDivider_v0p0p1_0.V13.n3 resistorDivider_v0p0p1_0.V13.n2 0.141636
R22887 resistorDivider_v0p0p1_0.V13.n1 resistorDivider_v0p0p1_0.V13 0.12425
R22888 resistorDivider_v0p0p1_0.V13 resistorDivider_v0p0p1_0.V13.n9 0.0991174
R22889 resistorDivider_v0p0p1_0.V13 resistorDivider_v0p0p1_0.V13.n1 0.0314375
R22890 resistorDivider_v0p0p1_0.V13.n2 resistorDivider_v0p0p1_0.V13.t0 0.00250214
R22891 resistorDivider_v0p0p1_0.V13.n2 resistorDivider_v0p0p1_0.V13.t4 0.000502142
R22892 resistorDivider_v0p0p1_0.V13.n3 resistorDivider_v0p0p1_0.V13.t5 0.000502142
R22893 resistorDivider_v0p0p1_0.V13.n4 resistorDivider_v0p0p1_0.V13.t3 0.000502142
R22894 resistorDivider_v0p0p1_0.V13.n5 resistorDivider_v0p0p1_0.V13.t1 0.000502142
R22895 resistorDivider_v0p0p1_0.V13.n6 resistorDivider_v0p0p1_0.V13.t11 0.000502142
R22896 resistorDivider_v0p0p1_0.V13.n7 resistorDivider_v0p0p1_0.V13.t8 0.000502142
R22897 resistorDivider_v0p0p1_0.V13.n8 resistorDivider_v0p0p1_0.V13.t12 0.000502142
R22898 resistorDivider_v0p0p1_0.V13.n9 resistorDivider_v0p0p1_0.V13.t14 0.000502142
R22899 resistorDivider_v0p0p1_0.V13.n9 resistorDivider_v0p0p1_0.V13.t15 0.000502142
R22900 resistorDivider_v0p0p1_0.V13.n8 resistorDivider_v0p0p1_0.V13.t10 0.000502142
R22901 resistorDivider_v0p0p1_0.V13.n7 resistorDivider_v0p0p1_0.V13.t7 0.000502142
R22902 resistorDivider_v0p0p1_0.V13.n6 resistorDivider_v0p0p1_0.V13.t2 0.000502142
R22903 resistorDivider_v0p0p1_0.V13.n5 resistorDivider_v0p0p1_0.V13.t9 0.000502142
R22904 resistorDivider_v0p0p1_0.V13.n4 resistorDivider_v0p0p1_0.V13.t6 0.000502142
R22905 resistorDivider_v0p0p1_0.V13.n3 resistorDivider_v0p0p1_0.V13.t13 0.000502142
R22906 VIN.n3 VIN.t19 167.326
R22907 VIN.n18 VIN.t11 167.326
R22908 VIN.n17 VIN.t5 167.326
R22909 VIN.n16 VIN.t20 167.326
R22910 VIN.n15 VIN.t15 167.326
R22911 VIN.n14 VIN.t26 167.326
R22912 VIN.n13 VIN.t23 167.326
R22913 VIN.n12 VIN.t1 167.326
R22914 VIN.n11 VIN.t28 167.326
R22915 VIN.n10 VIN.t13 167.326
R22916 VIN.n9 VIN.t6 167.326
R22917 VIN.n8 VIN.t31 167.326
R22918 VIN.n7 VIN.t16 167.326
R22919 VIN.n6 VIN.t10 167.326
R22920 VIN.n5 VIN.t24 167.326
R22921 VIN.n0 VIN.t4 167.326
R22922 VIN.n3 VIN.t17 92.4649
R22923 VIN.n18 VIN.t7 92.4649
R22924 VIN.n17 VIN.t0 92.4649
R22925 VIN.n16 VIN.t18 92.4649
R22926 VIN.n15 VIN.t12 92.4649
R22927 VIN.n14 VIN.t25 92.4649
R22928 VIN.n13 VIN.t21 92.4649
R22929 VIN.n12 VIN.t30 92.4649
R22930 VIN.n11 VIN.t27 92.4649
R22931 VIN.n10 VIN.t9 92.4649
R22932 VIN.n9 VIN.t2 92.4649
R22933 VIN.n8 VIN.t29 92.4649
R22934 VIN.n7 VIN.t14 92.4649
R22935 VIN.n6 VIN.t8 92.4649
R22936 VIN.n5 VIN.t22 92.4649
R22937 VIN.n0 VIN.t3 92.4649
R22938 VIN.n1 VIN 4.6255
R22939 VIN.n2 VIN.n1 1.6255
R22940 VIN VIN.n18 1.49913
R22941 VIN VIN.n17 1.49913
R22942 VIN VIN.n16 1.49913
R22943 VIN VIN.n15 1.49913
R22944 VIN VIN.n14 1.49913
R22945 VIN VIN.n13 1.49913
R22946 VIN VIN.n12 1.49913
R22947 VIN VIN.n11 1.49913
R22948 VIN VIN.n10 1.49913
R22949 VIN VIN.n9 1.49913
R22950 VIN VIN.n8 1.49913
R22951 VIN VIN.n7 1.49913
R22952 VIN VIN.n5 1.49913
R22953 VIN.n1 VIN.n0 1.49913
R22954 VIN VIN.n3 1.46056
R22955 VIN VIN.n6 1.46056
R22956 VIN.n19 VIN 1.04323
R22957 VIN.n32 VIN.n4 0.573417
R22958 VIN.n32 VIN.n31 0.563
R22959 VIN.n31 VIN.n30 0.563
R22960 VIN.n30 VIN.n29 0.563
R22961 VIN.n29 VIN.n28 0.563
R22962 VIN.n28 VIN.n27 0.563
R22963 VIN.n27 VIN.n26 0.563
R22964 VIN.n26 VIN.n25 0.563
R22965 VIN.n25 VIN.n24 0.563
R22966 VIN.n24 VIN.n23 0.563
R22967 VIN.n23 VIN.n22 0.563
R22968 VIN.n22 VIN.n21 0.563
R22969 VIN.n21 VIN.n20 0.563
R22970 VIN.n20 VIN.n19 0.563
R22971 VIN.n4 VIN 0.517333
R22972 VIN.n25 VIN 0.496386
R22973 VIN.n20 VIN 0.484963
R22974 VIN.n22 VIN 0.484963
R22975 VIN.n23 VIN 0.484963
R22976 VIN.n24 VIN 0.484963
R22977 VIN.n26 VIN 0.484963
R22978 VIN.n27 VIN 0.484963
R22979 VIN.n28 VIN 0.484963
R22980 VIN.n21 VIN 0.480732
R22981 VIN.n29 VIN 0.480732
R22982 VIN.n33 VIN.n32 0.47425
R22983 VIN.n19 VIN 0.473007
R22984 VIN.n31 VIN 0.473007
R22985 VIN.n30 VIN 0.45875
R22986 VIN.n2 VIN 0.316289
R22987 VIN.n4 VIN 0.169571
R22988 VIN VIN.n33 0.01
R22989 VIN.n33 VIN.n2 0.00707895
R22990 frontAnalog_v0p0p1_4.x65.A.n1 frontAnalog_v0p0p1_4.x65.A.t4 260.322
R22991 frontAnalog_v0p0p1_4.x65.A.n3 frontAnalog_v0p0p1_4.x65.A.t7 233.929
R22992 frontAnalog_v0p0p1_4.x65.A.n1 frontAnalog_v0p0p1_4.x65.A.t5 175.169
R22993 frontAnalog_v0p0p1_4.x65.A.n2 frontAnalog_v0p0p1_4.x65.A.t6 160.416
R22994 frontAnalog_v0p0p1_4.x65.A.n4 frontAnalog_v0p0p1_4.x65.A.t2 17.4109
R22995 frontAnalog_v0p0p1_4.x65.A.n4 frontAnalog_v0p0p1_4.x65.A.t3 10.2053
R22996 frontAnalog_v0p0p1_4.x65.A.n0 frontAnalog_v0p0p1_4.x65.A 2.78715
R22997 frontAnalog_v0p0p1_4.x65.A.n0 frontAnalog_v0p0p1_4.x65.A.n1 9.09103
R22998 frontAnalog_v0p0p1_4.x65.A.n6 frontAnalog_v0p0p1_4.x65.A.t0 7.94569
R22999 frontAnalog_v0p0p1_4.x65.A.n2 frontAnalog_v0p0p1_4.x65.A.t1 7.55846
R23000 frontAnalog_v0p0p1_4.x65.A.n5 frontAnalog_v0p0p1_4.x65.A.n3 1.4614
R23001 frontAnalog_v0p0p1_4.x65.A.n3 frontAnalog_v0p0p1_4.x65.A.n2 1.19626
R23002 frontAnalog_v0p0p1_4.x65.A.n6 frontAnalog_v0p0p1_4.x65.A.n5 0.836961
R23003 frontAnalog_v0p0p1_4.x65.A frontAnalog_v0p0p1_4.x65.A.n0 0.390342
R23004 frontAnalog_v0p0p1_4.x65.A.n5 frontAnalog_v0p0p1_4.x65.A.n4 0.154668
R23005 frontAnalog_v0p0p1_4.x65.A frontAnalog_v0p0p1_4.x65.A.n6 0.08175
R23006 resistorDivider_v0p0p1_0.V12.n0 resistorDivider_v0p0p1_0.V12.t17 167.365
R23007 resistorDivider_v0p0p1_0.V12.n0 resistorDivider_v0p0p1_0.V12.t16 92.4496
R23008 resistorDivider_v0p0p1_0.V12.n1 resistorDivider_v0p0p1_0.V12.n0 2.07493
R23009 resistorDivider_v0p0p1_0.V12.n15 resistorDivider_v0p0p1_0.V12.n14 0.141409
R23010 resistorDivider_v0p0p1_0.V12.n13 resistorDivider_v0p0p1_0.V12.n12 0.141409
R23011 resistorDivider_v0p0p1_0.V12.n11 resistorDivider_v0p0p1_0.V12.n10 0.141409
R23012 resistorDivider_v0p0p1_0.V12.n9 resistorDivider_v0p0p1_0.V12.n8 0.141409
R23013 resistorDivider_v0p0p1_0.V12.n7 resistorDivider_v0p0p1_0.V12.n6 0.141409
R23014 resistorDivider_v0p0p1_0.V12.n5 resistorDivider_v0p0p1_0.V12.n4 0.141409
R23015 resistorDivider_v0p0p1_0.V12.n3 resistorDivider_v0p0p1_0.V12.n2 0.141409
R23016 resistorDivider_v0p0p1_0.V12.n1 resistorDivider_v0p0p1_0.V12 0.12425
R23017 resistorDivider_v0p0p1_0.V12 resistorDivider_v0p0p1_0.V12.n16 0.100973
R23018 resistorDivider_v0p0p1_0.V12 resistorDivider_v0p0p1_0.V12.n1 0.0314375
R23019 resistorDivider_v0p0p1_0.V12.n7 resistorDivider_v0p0p1_0.V12.t0 0.00250214
R23020 resistorDivider_v0p0p1_0.V12.n2 resistorDivider_v0p0p1_0.V12.t3 0.000729415
R23021 resistorDivider_v0p0p1_0.V12.n16 resistorDivider_v0p0p1_0.V12.n15 0.000727273
R23022 resistorDivider_v0p0p1_0.V12.n14 resistorDivider_v0p0p1_0.V12.n13 0.000727273
R23023 resistorDivider_v0p0p1_0.V12.n12 resistorDivider_v0p0p1_0.V12.n11 0.000727273
R23024 resistorDivider_v0p0p1_0.V12.n10 resistorDivider_v0p0p1_0.V12.n9 0.000727273
R23025 resistorDivider_v0p0p1_0.V12.n8 resistorDivider_v0p0p1_0.V12.n7 0.000727273
R23026 resistorDivider_v0p0p1_0.V12.n6 resistorDivider_v0p0p1_0.V12.n5 0.000727273
R23027 resistorDivider_v0p0p1_0.V12.n4 resistorDivider_v0p0p1_0.V12.n3 0.000727273
R23028 resistorDivider_v0p0p1_0.V12.n2 resistorDivider_v0p0p1_0.V12.t6 0.000502142
R23029 resistorDivider_v0p0p1_0.V12.n4 resistorDivider_v0p0p1_0.V12.t7 0.000502142
R23030 resistorDivider_v0p0p1_0.V12.n6 resistorDivider_v0p0p1_0.V12.t10 0.000502142
R23031 resistorDivider_v0p0p1_0.V12.n8 resistorDivider_v0p0p1_0.V12.t12 0.000502142
R23032 resistorDivider_v0p0p1_0.V12.n10 resistorDivider_v0p0p1_0.V12.t1 0.000502142
R23033 resistorDivider_v0p0p1_0.V12.n12 resistorDivider_v0p0p1_0.V12.t9 0.000502142
R23034 resistorDivider_v0p0p1_0.V12.n14 resistorDivider_v0p0p1_0.V12.t4 0.000502142
R23035 resistorDivider_v0p0p1_0.V12.n16 resistorDivider_v0p0p1_0.V12.t14 0.000502142
R23036 resistorDivider_v0p0p1_0.V12.n15 resistorDivider_v0p0p1_0.V12.t15 0.000502142
R23037 resistorDivider_v0p0p1_0.V12.n13 resistorDivider_v0p0p1_0.V12.t13 0.000502142
R23038 resistorDivider_v0p0p1_0.V12.n11 resistorDivider_v0p0p1_0.V12.t8 0.000502142
R23039 resistorDivider_v0p0p1_0.V12.n9 resistorDivider_v0p0p1_0.V12.t11 0.000502142
R23040 resistorDivider_v0p0p1_0.V12.n5 resistorDivider_v0p0p1_0.V12.t2 0.000502142
R23041 resistorDivider_v0p0p1_0.V12.n3 resistorDivider_v0p0p1_0.V12.t5 0.000502142
R23042 frontAnalog_v0p0p1_9.x63.A.n2 frontAnalog_v0p0p1_9.x63.A.t5 260.322
R23043 frontAnalog_v0p0p1_9.x63.A.n4 frontAnalog_v0p0p1_9.x63.A.t6 233.888
R23044 frontAnalog_v0p0p1_9.x63.A.n2 frontAnalog_v0p0p1_9.x63.A.t7 175.169
R23045 frontAnalog_v0p0p1_9.x63.A.n3 frontAnalog_v0p0p1_9.x63.A.t4 159.725
R23046 frontAnalog_v0p0p1_9.x63.A.n1 frontAnalog_v0p0p1_9.x63.A.t0 17.4109
R23047 frontAnalog_v0p0p1_9.x63.A.n0 frontAnalog_v0p0p1_9.x63.A.n2 9.75129
R23048 frontAnalog_v0p0p1_9.x63.A.n1 frontAnalog_v0p0p1_9.x63.A.t1 9.6027
R23049 frontAnalog_v0p0p1_9.x63.A.n0 frontAnalog_v0p0p1_9.x63.A 2.33338
R23050 frontAnalog_v0p0p1_9.x63.A.n5 frontAnalog_v0p0p1_9.x63.A.t2 8.40929
R23051 frontAnalog_v0p0p1_9.x63.A.n3 frontAnalog_v0p0p1_9.x63.A.t3 8.06629
R23052 frontAnalog_v0p0p1_9.x63.A.n4 frontAnalog_v0p0p1_9.x63.A.n3 1.73501
R23053 frontAnalog_v0p0p1_9.x63.A.n1 frontAnalog_v0p0p1_9.x63.A.n4 0.99025
R23054 frontAnalog_v0p0p1_9.x63.A.n5 frontAnalog_v0p0p1_9.x63.A.n1 0.853186
R23055 frontAnalog_v0p0p1_9.x63.A frontAnalog_v0p0p1_9.x63.A.n0 0.349517
R23056 frontAnalog_v0p0p1_9.x63.A frontAnalog_v0p0p1_9.x63.A.n5 0.24425
R23057 frontAnalog_v0p0p1_9.x65.A.n1 frontAnalog_v0p0p1_9.x65.A.t6 260.322
R23058 frontAnalog_v0p0p1_9.x65.A.n3 frontAnalog_v0p0p1_9.x65.A.t5 233.929
R23059 frontAnalog_v0p0p1_9.x65.A.n1 frontAnalog_v0p0p1_9.x65.A.t4 175.169
R23060 frontAnalog_v0p0p1_9.x65.A.n2 frontAnalog_v0p0p1_9.x65.A.t7 160.416
R23061 frontAnalog_v0p0p1_9.x65.A.n4 frontAnalog_v0p0p1_9.x65.A.t0 17.4109
R23062 frontAnalog_v0p0p1_9.x65.A.n4 frontAnalog_v0p0p1_9.x65.A.t1 10.2053
R23063 frontAnalog_v0p0p1_9.x65.A.n0 frontAnalog_v0p0p1_9.x65.A 2.78715
R23064 frontAnalog_v0p0p1_9.x65.A.n0 frontAnalog_v0p0p1_9.x65.A.n1 9.09103
R23065 frontAnalog_v0p0p1_9.x65.A.n6 frontAnalog_v0p0p1_9.x65.A.t2 7.94569
R23066 frontAnalog_v0p0p1_9.x65.A.n2 frontAnalog_v0p0p1_9.x65.A.t3 7.55846
R23067 frontAnalog_v0p0p1_9.x65.A.n5 frontAnalog_v0p0p1_9.x65.A.n3 1.4614
R23068 frontAnalog_v0p0p1_9.x65.A.n3 frontAnalog_v0p0p1_9.x65.A.n2 1.19626
R23069 frontAnalog_v0p0p1_9.x65.A.n6 frontAnalog_v0p0p1_9.x65.A.n5 0.836961
R23070 frontAnalog_v0p0p1_9.x65.A frontAnalog_v0p0p1_9.x65.A.n0 0.390342
R23071 frontAnalog_v0p0p1_9.x65.A.n5 frontAnalog_v0p0p1_9.x65.A.n4 0.154668
R23072 frontAnalog_v0p0p1_9.x65.A frontAnalog_v0p0p1_9.x65.A.n6 0.08175
R23073 frontAnalog_v0p0p1_14.Q.t8 frontAnalog_v0p0p1_14.Q.t9 618.109
R23074 frontAnalog_v0p0p1_14.Q.n1 frontAnalog_v0p0p1_14.Q.t7 334.723
R23075 frontAnalog_v0p0p1_14.Q frontAnalog_v0p0p1_14.Q.t8 253.56
R23076 frontAnalog_v0p0p1_14.Q.n1 frontAnalog_v0p0p1_14.Q.t6 206.19
R23077 frontAnalog_v0p0p1_14.Q.n5 frontAnalog_v0p0p1_14.Q.t10 117.314
R23078 frontAnalog_v0p0p1_14.Q.n5 frontAnalog_v0p0p1_14.Q.t5 110.853
R23079 frontAnalog_v0p0p1_14.Q frontAnalog_v0p0p1_14.Q.n1 90.4462
R23080 frontAnalog_v0p0p1_14.Q.n0 frontAnalog_v0p0p1_14.Q 39.0702
R23081 frontAnalog_v0p0p1_14.Q.n6 frontAnalog_v0p0p1_14.Q.t0 17.6181
R23082 frontAnalog_v0p0p1_14.Q.n8 frontAnalog_v0p0p1_14.Q.t3 14.2865
R23083 frontAnalog_v0p0p1_14.Q.n10 frontAnalog_v0p0p1_14.Q.t1 14.283
R23084 frontAnalog_v0p0p1_14.Q.n10 frontAnalog_v0p0p1_14.Q.t2 14.283
R23085 frontAnalog_v0p0p1_14.Q.n13 frontAnalog_v0p0p1_14.Q.n4 9.01335
R23086 frontAnalog_v0p0p1_14.Q.n12 frontAnalog_v0p0p1_14.Q.t4 8.77744
R23087 frontAnalog_v0p0p1_14.Q.n2 frontAnalog_v0p0p1_14.Q 7.13193
R23088 frontAnalog_v0p0p1_14.Q.n2 frontAnalog_v0p0p1_14.Q 5.30336
R23089 frontAnalog_v0p0p1_14.Q.n3 frontAnalog_v0p0p1_14.Q.n2 5.16688
R23090 frontAnalog_v0p0p1_14.Q.n3 frontAnalog_v0p0p1_14.Q.n0 2.29514
R23091 frontAnalog_v0p0p1_14.Q.n12 frontAnalog_v0p0p1_14.Q.n11 1.20426
R23092 frontAnalog_v0p0p1_14.Q.n0 frontAnalog_v0p0p1_14.Q 0.692911
R23093 frontAnalog_v0p0p1_14.Q.n13 frontAnalog_v0p0p1_14.Q.n12 0.325111
R23094 frontAnalog_v0p0p1_14.Q.n9 frontAnalog_v0p0p1_14.Q.n8 0.301242
R23095 frontAnalog_v0p0p1_14.Q.n4 frontAnalog_v0p0p1_14.Q 0.20675
R23096 frontAnalog_v0p0p1_14.Q.n7 frontAnalog_v0p0p1_14.Q.n5 0.159555
R23097 frontAnalog_v0p0p1_14.Q.n4 frontAnalog_v0p0p1_14.Q.n3 0.153447
R23098 frontAnalog_v0p0p1_14.Q.n11 frontAnalog_v0p0p1_14.Q.n10 0.106617
R23099 frontAnalog_v0p0p1_14.Q.n9 frontAnalog_v0p0p1_14.Q.n7 0.0796167
R23100 frontAnalog_v0p0p1_14.Q.n11 frontAnalog_v0p0p1_14.Q.n9 0.0480595
R23101 frontAnalog_v0p0p1_14.Q frontAnalog_v0p0p1_14.Q.n13 0.0469368
R23102 frontAnalog_v0p0p1_14.Q.n7 frontAnalog_v0p0p1_14.Q.n6 0.000504658
R23103 frontAnalog_v0p0p1_9.RSfetsym_0.QN.n1 frontAnalog_v0p0p1_9.RSfetsym_0.QN.t6 117.511
R23104 frontAnalog_v0p0p1_9.RSfetsym_0.QN.n1 frontAnalog_v0p0p1_9.RSfetsym_0.QN.t5 110.698
R23105 frontAnalog_v0p0p1_9.RSfetsym_0.QN.n4 frontAnalog_v0p0p1_9.RSfetsym_0.QN.t3 19.1963
R23106 frontAnalog_v0p0p1_9.RSfetsym_0.QN.n7 frontAnalog_v0p0p1_9.RSfetsym_0.QN.t4 14.2842
R23107 frontAnalog_v0p0p1_9.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_9.RSfetsym_0.QN.t1 14.283
R23108 frontAnalog_v0p0p1_9.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_9.RSfetsym_0.QN.t2 14.283
R23109 frontAnalog_v0p0p1_9.RSfetsym_0.QN.n11 frontAnalog_v0p0p1_9.RSfetsym_0.QN.t0 9.14075
R23110 frontAnalog_v0p0p1_9.RSfetsym_0.QN.n11 frontAnalog_v0p0p1_9.RSfetsym_0.QN.n10 0.74645
R23111 frontAnalog_v0p0p1_9.RSfetsym_0.QN.n2 frontAnalog_v0p0p1_9.RSfetsym_0.QN.n1 0.688382
R23112 frontAnalog_v0p0p1_9.RSfetsym_0.QN.n10 frontAnalog_v0p0p1_9.RSfetsym_0.QN.n9 0.2402
R23113 frontAnalog_v0p0p1_9.RSfetsym_0.QN.n9 frontAnalog_v0p0p1_9.RSfetsym_0.QN.n8 0.236824
R23114 frontAnalog_v0p0p1_9.RSfetsym_0.QN.n4 frontAnalog_v0p0p1_9.RSfetsym_0.QN.n3 0.132187
R23115 frontAnalog_v0p0p1_9.RSfetsym_0.QN.n9 frontAnalog_v0p0p1_9.RSfetsym_0.QN.n4 0.0968646
R23116 frontAnalog_v0p0p1_9.RSfetsym_0.QN frontAnalog_v0p0p1_9.RSfetsym_0.QN.n11 0.0446535
R23117 frontAnalog_v0p0p1_9.RSfetsym_0.QN.n8 frontAnalog_v0p0p1_9.RSfetsym_0.QN.n6 0.0272538
R23118 frontAnalog_v0p0p1_9.RSfetsym_0.QN.n10 frontAnalog_v0p0p1_9.RSfetsym_0.QN.n0 0.00981499
R23119 frontAnalog_v0p0p1_9.RSfetsym_0.QN.n3 frontAnalog_v0p0p1_9.RSfetsym_0.QN.n2 0.00725433
R23120 frontAnalog_v0p0p1_9.RSfetsym_0.QN.n6 frontAnalog_v0p0p1_9.RSfetsym_0.QN.n5 0.00610579
R23121 frontAnalog_v0p0p1_9.RSfetsym_0.QN.n8 frontAnalog_v0p0p1_9.RSfetsym_0.QN.n7 0.00225341
R23122 frontAnalog_v0p0p1_9.Q.n17 frontAnalog_v0p0p1_9.Q.t6 260.435
R23123 frontAnalog_v0p0p1_9.Q.n2 frontAnalog_v0p0p1_9.Q.t10 229.433
R23124 frontAnalog_v0p0p1_9.Q.n12 frontAnalog_v0p0p1_9.Q.t11 196.549
R23125 frontAnalog_v0p0p1_9.Q.n2 frontAnalog_v0p0p1_9.Q.t7 158.885
R23126 frontAnalog_v0p0p1_9.Q.n17 frontAnalog_v0p0p1_9.Q.t8 156.403
R23127 frontAnalog_v0p0p1_9.Q.n12 frontAnalog_v0p0p1_9.Q.t12 148.35
R23128 frontAnalog_v0p0p1_9.Q.n25 frontAnalog_v0p0p1_9.Q.t9 117.314
R23129 frontAnalog_v0p0p1_9.Q.n25 frontAnalog_v0p0p1_9.Q.t5 110.853
R23130 frontAnalog_v0p0p1_9.Q.n13 frontAnalog_v0p0p1_9.Q.n12 76.0005
R23131 frontAnalog_v0p0p1_9.Q.n26 frontAnalog_v0p0p1_9.Q.t2 17.6181
R23132 frontAnalog_v0p0p1_9.Q.n28 frontAnalog_v0p0p1_9.Q.t3 14.2865
R23133 frontAnalog_v0p0p1_9.Q.n30 frontAnalog_v0p0p1_9.Q.t0 14.283
R23134 frontAnalog_v0p0p1_9.Q.n30 frontAnalog_v0p0p1_9.Q.t1 14.283
R23135 frontAnalog_v0p0p1_9.Q frontAnalog_v0p0p1_9.Q.n16 9.3005
R23136 frontAnalog_v0p0p1_9.Q.n32 frontAnalog_v0p0p1_9.Q.t4 8.77744
R23137 frontAnalog_v0p0p1_9.Q.n18 frontAnalog_v0p0p1_9.Q.n17 7.60183
R23138 frontAnalog_v0p0p1_9.Q.n3 frontAnalog_v0p0p1_9.Q.n2 7.39171
R23139 frontAnalog_v0p0p1_9.Q.n22 frontAnalog_v0p0p1_9.Q.n14 6.24391
R23140 frontAnalog_v0p0p1_9.Q.n13 frontAnalog_v0p0p1_9.Q 5.78114
R23141 frontAnalog_v0p0p1_9.Q.n18 frontAnalog_v0p0p1_9.Q 4.8645
R23142 frontAnalog_v0p0p1_9.Q.n6 frontAnalog_v0p0p1_9.Q.n5 4.5005
R23143 frontAnalog_v0p0p1_9.Q.n22 frontAnalog_v0p0p1_9.Q.n21 3.53643
R23144 frontAnalog_v0p0p1_9.Q.n14 frontAnalog_v0p0p1_9.Q.n13 3.51018
R23145 frontAnalog_v0p0p1_9.Q.n5 frontAnalog_v0p0p1_9.Q.n4 3.46717
R23146 frontAnalog_v0p0p1_9.Q.n33 frontAnalog_v0p0p1_9.Q.n24 3.13935
R23147 frontAnalog_v0p0p1_9.Q.n32 frontAnalog_v0p0p1_9.Q.n31 1.20426
R23148 frontAnalog_v0p0p1_9.Q.n11 frontAnalog_v0p0p1_9.Q.n10 1.11384
R23149 frontAnalog_v0p0p1_9.Q.n5 frontAnalog_v0p0p1_9.Q.n3 1.06717
R23150 frontAnalog_v0p0p1_9.Q.n4 frontAnalog_v0p0p1_9.Q 1.06717
R23151 frontAnalog_v0p0p1_9.Q.n23 frontAnalog_v0p0p1_9.Q.n11 0.874607
R23152 frontAnalog_v0p0p1_9.Q.n24 frontAnalog_v0p0p1_9.Q.n23 0.520635
R23153 frontAnalog_v0p0p1_9.Q.n11 frontAnalog_v0p0p1_9.Q 0.372375
R23154 frontAnalog_v0p0p1_9.Q.n33 frontAnalog_v0p0p1_9.Q.n32 0.325111
R23155 frontAnalog_v0p0p1_9.Q.n29 frontAnalog_v0p0p1_9.Q.n28 0.301242
R23156 frontAnalog_v0p0p1_9.Q.n23 frontAnalog_v0p0p1_9.Q.n22 0.214786
R23157 frontAnalog_v0p0p1_9.Q.n14 frontAnalog_v0p0p1_9.Q 0.206952
R23158 frontAnalog_v0p0p1_9.Q.n24 frontAnalog_v0p0p1_9.Q 0.20675
R23159 frontAnalog_v0p0p1_9.Q.n27 frontAnalog_v0p0p1_9.Q.n25 0.159555
R23160 frontAnalog_v0p0p1_9.Q.n31 frontAnalog_v0p0p1_9.Q.n30 0.106617
R23161 frontAnalog_v0p0p1_9.Q.n29 frontAnalog_v0p0p1_9.Q.n27 0.0796167
R23162 frontAnalog_v0p0p1_9.Q.n31 frontAnalog_v0p0p1_9.Q.n29 0.0480595
R23163 frontAnalog_v0p0p1_9.Q frontAnalog_v0p0p1_9.Q.n33 0.0469368
R23164 frontAnalog_v0p0p1_9.Q.n20 frontAnalog_v0p0p1_9.Q.n16 0.0344286
R23165 frontAnalog_v0p0p1_9.Q.n10 frontAnalog_v0p0p1_9.Q.n9 0.028
R23166 frontAnalog_v0p0p1_9.Q.n8 frontAnalog_v0p0p1_9.Q.n7 0.0142363
R23167 frontAnalog_v0p0p1_9.Q.n8 frontAnalog_v0p0p1_9.Q.n6 0.00599451
R23168 frontAnalog_v0p0p1_9.Q.n1 frontAnalog_v0p0p1_9.Q.n0 0.00484776
R23169 frontAnalog_v0p0p1_9.Q.n6 frontAnalog_v0p0p1_9.Q.n1 0.00226981
R23170 frontAnalog_v0p0p1_9.Q.n21 frontAnalog_v0p0p1_9.Q.n15 0.00182856
R23171 frontAnalog_v0p0p1_9.Q.n21 frontAnalog_v0p0p1_9.Q.n20 0.00149885
R23172 frontAnalog_v0p0p1_9.Q.n19 frontAnalog_v0p0p1_9.Q.n18 0.00133362
R23173 frontAnalog_v0p0p1_9.Q.n20 frontAnalog_v0p0p1_9.Q.n19 0.00100077
R23174 frontAnalog_v0p0p1_9.Q.n9 frontAnalog_v0p0p1_9.Q.n8 0.000617139
R23175 frontAnalog_v0p0p1_9.Q.n27 frontAnalog_v0p0p1_9.Q.n26 0.000504658
R23176 frontAnalog_v0p0p1_13.RSfetsym_0.QN.n1 frontAnalog_v0p0p1_13.RSfetsym_0.QN.t6 117.511
R23177 frontAnalog_v0p0p1_13.RSfetsym_0.QN.n1 frontAnalog_v0p0p1_13.RSfetsym_0.QN.t5 110.698
R23178 frontAnalog_v0p0p1_13.RSfetsym_0.QN.n4 frontAnalog_v0p0p1_13.RSfetsym_0.QN.t2 19.1963
R23179 frontAnalog_v0p0p1_13.RSfetsym_0.QN.n7 frontAnalog_v0p0p1_13.RSfetsym_0.QN.t4 14.2842
R23180 frontAnalog_v0p0p1_13.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_13.RSfetsym_0.QN.t1 14.283
R23181 frontAnalog_v0p0p1_13.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_13.RSfetsym_0.QN.t0 14.283
R23182 frontAnalog_v0p0p1_13.RSfetsym_0.QN.n11 frontAnalog_v0p0p1_13.RSfetsym_0.QN.t3 9.14075
R23183 frontAnalog_v0p0p1_13.RSfetsym_0.QN.n11 frontAnalog_v0p0p1_13.RSfetsym_0.QN.n10 0.74645
R23184 frontAnalog_v0p0p1_13.RSfetsym_0.QN.n2 frontAnalog_v0p0p1_13.RSfetsym_0.QN.n1 0.688382
R23185 frontAnalog_v0p0p1_13.RSfetsym_0.QN.n10 frontAnalog_v0p0p1_13.RSfetsym_0.QN.n9 0.2402
R23186 frontAnalog_v0p0p1_13.RSfetsym_0.QN.n9 frontAnalog_v0p0p1_13.RSfetsym_0.QN.n8 0.236824
R23187 frontAnalog_v0p0p1_13.RSfetsym_0.QN.n4 frontAnalog_v0p0p1_13.RSfetsym_0.QN.n3 0.132187
R23188 frontAnalog_v0p0p1_13.RSfetsym_0.QN.n9 frontAnalog_v0p0p1_13.RSfetsym_0.QN.n4 0.0968646
R23189 frontAnalog_v0p0p1_13.RSfetsym_0.QN frontAnalog_v0p0p1_13.RSfetsym_0.QN.n11 0.0446535
R23190 frontAnalog_v0p0p1_13.RSfetsym_0.QN.n8 frontAnalog_v0p0p1_13.RSfetsym_0.QN.n6 0.0272538
R23191 frontAnalog_v0p0p1_13.RSfetsym_0.QN.n10 frontAnalog_v0p0p1_13.RSfetsym_0.QN.n0 0.00981499
R23192 frontAnalog_v0p0p1_13.RSfetsym_0.QN.n3 frontAnalog_v0p0p1_13.RSfetsym_0.QN.n2 0.00725433
R23193 frontAnalog_v0p0p1_13.RSfetsym_0.QN.n6 frontAnalog_v0p0p1_13.RSfetsym_0.QN.n5 0.00610579
R23194 frontAnalog_v0p0p1_13.RSfetsym_0.QN.n8 frontAnalog_v0p0p1_13.RSfetsym_0.QN.n7 0.00225341
R23195 frontAnalog_v0p0p1_7.x65.A.n1 frontAnalog_v0p0p1_7.x65.A.t7 260.322
R23196 frontAnalog_v0p0p1_7.x65.A.n3 frontAnalog_v0p0p1_7.x65.A.t6 233.929
R23197 frontAnalog_v0p0p1_7.x65.A.n1 frontAnalog_v0p0p1_7.x65.A.t5 175.169
R23198 frontAnalog_v0p0p1_7.x65.A.n2 frontAnalog_v0p0p1_7.x65.A.t4 160.416
R23199 frontAnalog_v0p0p1_7.x65.A.n4 frontAnalog_v0p0p1_7.x65.A.t3 17.4109
R23200 frontAnalog_v0p0p1_7.x65.A.n4 frontAnalog_v0p0p1_7.x65.A.t2 10.2053
R23201 frontAnalog_v0p0p1_7.x65.A.n0 frontAnalog_v0p0p1_7.x65.A 2.78715
R23202 frontAnalog_v0p0p1_7.x65.A.n0 frontAnalog_v0p0p1_7.x65.A.n1 9.09103
R23203 frontAnalog_v0p0p1_7.x65.A.n6 frontAnalog_v0p0p1_7.x65.A.t0 7.94569
R23204 frontAnalog_v0p0p1_7.x65.A.n2 frontAnalog_v0p0p1_7.x65.A.t1 7.55846
R23205 frontAnalog_v0p0p1_7.x65.A.n5 frontAnalog_v0p0p1_7.x65.A.n3 1.4614
R23206 frontAnalog_v0p0p1_7.x65.A.n3 frontAnalog_v0p0p1_7.x65.A.n2 1.19626
R23207 frontAnalog_v0p0p1_7.x65.A.n6 frontAnalog_v0p0p1_7.x65.A.n5 0.836961
R23208 frontAnalog_v0p0p1_7.x65.A frontAnalog_v0p0p1_7.x65.A.n0 0.390342
R23209 frontAnalog_v0p0p1_7.x65.A.n5 frontAnalog_v0p0p1_7.x65.A.n4 0.154668
R23210 frontAnalog_v0p0p1_7.x65.A frontAnalog_v0p0p1_7.x65.A.n6 0.08175
R23211 frontAnalog_v0p0p1_7.x63.A.n2 frontAnalog_v0p0p1_7.x63.A.t6 260.322
R23212 frontAnalog_v0p0p1_7.x63.A.n4 frontAnalog_v0p0p1_7.x63.A.t7 233.888
R23213 frontAnalog_v0p0p1_7.x63.A.n2 frontAnalog_v0p0p1_7.x63.A.t4 175.169
R23214 frontAnalog_v0p0p1_7.x63.A.n3 frontAnalog_v0p0p1_7.x63.A.t5 159.725
R23215 frontAnalog_v0p0p1_7.x63.A.n1 frontAnalog_v0p0p1_7.x63.A.t2 17.4109
R23216 frontAnalog_v0p0p1_7.x63.A.n0 frontAnalog_v0p0p1_7.x63.A.n2 9.75129
R23217 frontAnalog_v0p0p1_7.x63.A.n1 frontAnalog_v0p0p1_7.x63.A.t3 9.6037
R23218 frontAnalog_v0p0p1_7.x63.A.n0 frontAnalog_v0p0p1_7.x63.A 2.33338
R23219 frontAnalog_v0p0p1_7.x63.A.n5 frontAnalog_v0p0p1_7.x63.A.t1 8.40929
R23220 frontAnalog_v0p0p1_7.x63.A.n3 frontAnalog_v0p0p1_7.x63.A.t0 8.06629
R23221 frontAnalog_v0p0p1_7.x63.A.n4 frontAnalog_v0p0p1_7.x63.A.n3 1.73501
R23222 frontAnalog_v0p0p1_7.x63.A.n1 frontAnalog_v0p0p1_7.x63.A.n4 0.99025
R23223 frontAnalog_v0p0p1_7.x63.A.n5 frontAnalog_v0p0p1_7.x63.A.n1 0.853186
R23224 frontAnalog_v0p0p1_7.x63.A frontAnalog_v0p0p1_7.x63.A.n0 0.349517
R23225 frontAnalog_v0p0p1_7.x63.A frontAnalog_v0p0p1_7.x63.A.n5 0.24425
R23226 frontAnalog_v0p0p1_7.Q.t7 frontAnalog_v0p0p1_7.Q.t9 618.109
R23227 frontAnalog_v0p0p1_7.Q.n0 frontAnalog_v0p0p1_7.Q.t8 334.723
R23228 frontAnalog_v0p0p1_7.Q frontAnalog_v0p0p1_7.Q.t7 253.56
R23229 frontAnalog_v0p0p1_7.Q.n0 frontAnalog_v0p0p1_7.Q.t5 206.19
R23230 frontAnalog_v0p0p1_7.Q.n2 frontAnalog_v0p0p1_7.Q.t10 117.314
R23231 frontAnalog_v0p0p1_7.Q.n2 frontAnalog_v0p0p1_7.Q.t6 110.852
R23232 frontAnalog_v0p0p1_7.Q frontAnalog_v0p0p1_7.Q.n0 90.4462
R23233 frontAnalog_v0p0p1_7.Q frontAnalog_v0p0p1_7.Q.n13 39.0702
R23234 frontAnalog_v0p0p1_7.Q.n4 frontAnalog_v0p0p1_7.Q.t3 17.6181
R23235 frontAnalog_v0p0p1_7.Q.n5 frontAnalog_v0p0p1_7.Q.t0 14.2865
R23236 frontAnalog_v0p0p1_7.Q.n7 frontAnalog_v0p0p1_7.Q.t1 14.283
R23237 frontAnalog_v0p0p1_7.Q.n7 frontAnalog_v0p0p1_7.Q.t2 14.283
R23238 frontAnalog_v0p0p1_7.Q.n9 frontAnalog_v0p0p1_7.Q.t4 8.77592
R23239 frontAnalog_v0p0p1_7.Q.n1 frontAnalog_v0p0p1_7.Q 7.13193
R23240 frontAnalog_v0p0p1_7.Q.n1 frontAnalog_v0p0p1_7.Q 5.30336
R23241 frontAnalog_v0p0p1_7.Q.n12 frontAnalog_v0p0p1_7.Q.n1 5.27402
R23242 frontAnalog_v0p0p1_7.Q.n11 frontAnalog_v0p0p1_7.Q.n10 3.52037
R23243 frontAnalog_v0p0p1_7.Q.n13 frontAnalog_v0p0p1_7.Q.n12 2.188
R23244 frontAnalog_v0p0p1_7.Q.n9 frontAnalog_v0p0p1_7.Q.n8 1.20426
R23245 frontAnalog_v0p0p1_7.Q.n13 frontAnalog_v0p0p1_7.Q 0.692911
R23246 frontAnalog_v0p0p1_7.Q.n10 frontAnalog_v0p0p1_7.Q.n9 0.338241
R23247 frontAnalog_v0p0p1_7.Q.n5 frontAnalog_v0p0p1_7.Q.n4 0.313689
R23248 frontAnalog_v0p0p1_7.Q.n6 frontAnalog_v0p0p1_7.Q.n5 0.300242
R23249 frontAnalog_v0p0p1_7.Q.n11 frontAnalog_v0p0p1_7.Q 0.2005
R23250 frontAnalog_v0p0p1_7.Q.n12 frontAnalog_v0p0p1_7.Q.n11 0.166764
R23251 frontAnalog_v0p0p1_7.Q.n3 frontAnalog_v0p0p1_7.Q.n2 0.159555
R23252 frontAnalog_v0p0p1_7.Q.n8 frontAnalog_v0p0p1_7.Q.n7 0.106617
R23253 frontAnalog_v0p0p1_7.Q.n6 frontAnalog_v0p0p1_7.Q.n3 0.0796167
R23254 frontAnalog_v0p0p1_7.Q.n8 frontAnalog_v0p0p1_7.Q.n6 0.0480595
R23255 frontAnalog_v0p0p1_7.Q.n10 frontAnalog_v0p0p1_7.Q 0.00440792
R23256 frontAnalog_v0p0p1_7.Q.n4 frontAnalog_v0p0p1_7.Q.n3 0.000504658
R23257 resistorDivider_v0p0p1_0.V7.n0 resistorDivider_v0p0p1_0.V7.t16 167.365
R23258 resistorDivider_v0p0p1_0.V7.n0 resistorDivider_v0p0p1_0.V7.t17 92.4488
R23259 resistorDivider_v0p0p1_0.V7.n1 resistorDivider_v0p0p1_0.V7.n0 2.07493
R23260 resistorDivider_v0p0p1_0.V7.n9 resistorDivider_v0p0p1_0.V7.n8 0.141636
R23261 resistorDivider_v0p0p1_0.V7.n8 resistorDivider_v0p0p1_0.V7.n7 0.141636
R23262 resistorDivider_v0p0p1_0.V7.n7 resistorDivider_v0p0p1_0.V7.n6 0.141636
R23263 resistorDivider_v0p0p1_0.V7.n6 resistorDivider_v0p0p1_0.V7.n5 0.141636
R23264 resistorDivider_v0p0p1_0.V7.n5 resistorDivider_v0p0p1_0.V7.n4 0.141636
R23265 resistorDivider_v0p0p1_0.V7.n4 resistorDivider_v0p0p1_0.V7.n3 0.141636
R23266 resistorDivider_v0p0p1_0.V7.n3 resistorDivider_v0p0p1_0.V7.n2 0.141636
R23267 resistorDivider_v0p0p1_0.V7.n1 resistorDivider_v0p0p1_0.V7 0.12425
R23268 resistorDivider_v0p0p1_0.V7 resistorDivider_v0p0p1_0.V7.n9 0.101201
R23269 resistorDivider_v0p0p1_0.V7 resistorDivider_v0p0p1_0.V7.n1 0.028
R23270 resistorDivider_v0p0p1_0.V7.n9 resistorDivider_v0p0p1_0.V7.t0 0.00250214
R23271 resistorDivider_v0p0p1_0.V7.n3 resistorDivider_v0p0p1_0.V7.t3 0.000502142
R23272 resistorDivider_v0p0p1_0.V7.n4 resistorDivider_v0p0p1_0.V7.t10 0.000502142
R23273 resistorDivider_v0p0p1_0.V7.n5 resistorDivider_v0p0p1_0.V7.t8 0.000502142
R23274 resistorDivider_v0p0p1_0.V7.n6 resistorDivider_v0p0p1_0.V7.t1 0.000502142
R23275 resistorDivider_v0p0p1_0.V7.n7 resistorDivider_v0p0p1_0.V7.t15 0.000502142
R23276 resistorDivider_v0p0p1_0.V7.n8 resistorDivider_v0p0p1_0.V7.t6 0.000502142
R23277 resistorDivider_v0p0p1_0.V7.n2 resistorDivider_v0p0p1_0.V7.t2 0.000502142
R23278 resistorDivider_v0p0p1_0.V7.n3 resistorDivider_v0p0p1_0.V7.t7 0.000502142
R23279 resistorDivider_v0p0p1_0.V7.n4 resistorDivider_v0p0p1_0.V7.t11 0.000502142
R23280 resistorDivider_v0p0p1_0.V7.n5 resistorDivider_v0p0p1_0.V7.t12 0.000502142
R23281 resistorDivider_v0p0p1_0.V7.n6 resistorDivider_v0p0p1_0.V7.t9 0.000502142
R23282 resistorDivider_v0p0p1_0.V7.n7 resistorDivider_v0p0p1_0.V7.t14 0.000502142
R23283 resistorDivider_v0p0p1_0.V7.n8 resistorDivider_v0p0p1_0.V7.t4 0.000502142
R23284 resistorDivider_v0p0p1_0.V7.n9 resistorDivider_v0p0p1_0.V7.t13 0.000502142
R23285 resistorDivider_v0p0p1_0.V7.n2 resistorDivider_v0p0p1_0.V7.t5 0.000502142
R23286 resistorDivider_v0p0p1_0.V6.n0 resistorDivider_v0p0p1_0.V6.t17 167.365
R23287 resistorDivider_v0p0p1_0.V6.n0 resistorDivider_v0p0p1_0.V6.t16 92.4488
R23288 resistorDivider_v0p0p1_0.V6.n1 resistorDivider_v0p0p1_0.V6.n0 2.07493
R23289 resistorDivider_v0p0p1_0.V6.n15 resistorDivider_v0p0p1_0.V6.n14 0.141409
R23290 resistorDivider_v0p0p1_0.V6.n13 resistorDivider_v0p0p1_0.V6.n12 0.141409
R23291 resistorDivider_v0p0p1_0.V6.n11 resistorDivider_v0p0p1_0.V6.n10 0.141409
R23292 resistorDivider_v0p0p1_0.V6.n9 resistorDivider_v0p0p1_0.V6.n8 0.141409
R23293 resistorDivider_v0p0p1_0.V6.n7 resistorDivider_v0p0p1_0.V6.n6 0.141409
R23294 resistorDivider_v0p0p1_0.V6.n5 resistorDivider_v0p0p1_0.V6.n4 0.141409
R23295 resistorDivider_v0p0p1_0.V6.n3 resistorDivider_v0p0p1_0.V6.n2 0.141409
R23296 resistorDivider_v0p0p1_0.V6.n1 resistorDivider_v0p0p1_0.V6 0.12425
R23297 resistorDivider_v0p0p1_0.V6 resistorDivider_v0p0p1_0.V6.n16 0.0988902
R23298 resistorDivider_v0p0p1_0.V6 resistorDivider_v0p0p1_0.V6.n1 0.0314375
R23299 resistorDivider_v0p0p1_0.V6.n2 resistorDivider_v0p0p1_0.V6.t0 0.000729415
R23300 resistorDivider_v0p0p1_0.V6.n16 resistorDivider_v0p0p1_0.V6.n15 0.000727273
R23301 resistorDivider_v0p0p1_0.V6.n14 resistorDivider_v0p0p1_0.V6.n13 0.000727273
R23302 resistorDivider_v0p0p1_0.V6.n12 resistorDivider_v0p0p1_0.V6.n11 0.000727273
R23303 resistorDivider_v0p0p1_0.V6.n10 resistorDivider_v0p0p1_0.V6.n9 0.000727273
R23304 resistorDivider_v0p0p1_0.V6.n8 resistorDivider_v0p0p1_0.V6.n7 0.000727273
R23305 resistorDivider_v0p0p1_0.V6.n6 resistorDivider_v0p0p1_0.V6.n5 0.000727273
R23306 resistorDivider_v0p0p1_0.V6.n4 resistorDivider_v0p0p1_0.V6.n3 0.000727273
R23307 resistorDivider_v0p0p1_0.V6.n3 resistorDivider_v0p0p1_0.V6.t4 0.000502142
R23308 resistorDivider_v0p0p1_0.V6.n5 resistorDivider_v0p0p1_0.V6.t7 0.000502142
R23309 resistorDivider_v0p0p1_0.V6.n7 resistorDivider_v0p0p1_0.V6.t10 0.000502142
R23310 resistorDivider_v0p0p1_0.V6.n9 resistorDivider_v0p0p1_0.V6.t5 0.000502142
R23311 resistorDivider_v0p0p1_0.V6.n11 resistorDivider_v0p0p1_0.V6.t14 0.000502142
R23312 resistorDivider_v0p0p1_0.V6.n13 resistorDivider_v0p0p1_0.V6.t3 0.000502142
R23313 resistorDivider_v0p0p1_0.V6.n15 resistorDivider_v0p0p1_0.V6.t11 0.000502142
R23314 resistorDivider_v0p0p1_0.V6.n2 resistorDivider_v0p0p1_0.V6.t13 0.000502142
R23315 resistorDivider_v0p0p1_0.V6.n4 resistorDivider_v0p0p1_0.V6.t12 0.000502142
R23316 resistorDivider_v0p0p1_0.V6.n6 resistorDivider_v0p0p1_0.V6.t15 0.000502142
R23317 resistorDivider_v0p0p1_0.V6.n8 resistorDivider_v0p0p1_0.V6.t8 0.000502142
R23318 resistorDivider_v0p0p1_0.V6.n10 resistorDivider_v0p0p1_0.V6.t9 0.000502142
R23319 resistorDivider_v0p0p1_0.V6.n12 resistorDivider_v0p0p1_0.V6.t1 0.000502142
R23320 resistorDivider_v0p0p1_0.V6.n14 resistorDivider_v0p0p1_0.V6.t6 0.000502142
R23321 resistorDivider_v0p0p1_0.V6.n16 resistorDivider_v0p0p1_0.V6.t2 0.000502142
R23322 resistorDivider_v0p0p1_0.V5.n0 resistorDivider_v0p0p1_0.V5.t17 167.365
R23323 resistorDivider_v0p0p1_0.V5.n0 resistorDivider_v0p0p1_0.V5.t16 92.4488
R23324 resistorDivider_v0p0p1_0.V5.n1 resistorDivider_v0p0p1_0.V5.n0 2.07493
R23325 resistorDivider_v0p0p1_0.V5.n15 resistorDivider_v0p0p1_0.V5.n14 0.141409
R23326 resistorDivider_v0p0p1_0.V5.n13 resistorDivider_v0p0p1_0.V5.n12 0.141409
R23327 resistorDivider_v0p0p1_0.V5.n11 resistorDivider_v0p0p1_0.V5.n10 0.141409
R23328 resistorDivider_v0p0p1_0.V5.n9 resistorDivider_v0p0p1_0.V5.n8 0.141409
R23329 resistorDivider_v0p0p1_0.V5.n7 resistorDivider_v0p0p1_0.V5.n6 0.141409
R23330 resistorDivider_v0p0p1_0.V5.n5 resistorDivider_v0p0p1_0.V5.n4 0.141409
R23331 resistorDivider_v0p0p1_0.V5.n3 resistorDivider_v0p0p1_0.V5.n2 0.141409
R23332 resistorDivider_v0p0p1_0.V5.n1 resistorDivider_v0p0p1_0.V5 0.12425
R23333 resistorDivider_v0p0p1_0.V5 resistorDivider_v0p0p1_0.V5.n16 0.103057
R23334 resistorDivider_v0p0p1_0.V5 resistorDivider_v0p0p1_0.V5.n1 0.0314375
R23335 resistorDivider_v0p0p1_0.V5.n5 resistorDivider_v0p0p1_0.V5.t0 0.00250214
R23336 resistorDivider_v0p0p1_0.V5.n2 resistorDivider_v0p0p1_0.V5.t8 0.000729415
R23337 resistorDivider_v0p0p1_0.V5.n16 resistorDivider_v0p0p1_0.V5.n15 0.000727273
R23338 resistorDivider_v0p0p1_0.V5.n14 resistorDivider_v0p0p1_0.V5.n13 0.000727273
R23339 resistorDivider_v0p0p1_0.V5.n12 resistorDivider_v0p0p1_0.V5.n11 0.000727273
R23340 resistorDivider_v0p0p1_0.V5.n10 resistorDivider_v0p0p1_0.V5.n9 0.000727273
R23341 resistorDivider_v0p0p1_0.V5.n8 resistorDivider_v0p0p1_0.V5.n7 0.000727273
R23342 resistorDivider_v0p0p1_0.V5.n6 resistorDivider_v0p0p1_0.V5.n5 0.000727273
R23343 resistorDivider_v0p0p1_0.V5.n4 resistorDivider_v0p0p1_0.V5.n3 0.000727273
R23344 resistorDivider_v0p0p1_0.V5.n4 resistorDivider_v0p0p1_0.V5.t13 0.000502142
R23345 resistorDivider_v0p0p1_0.V5.n6 resistorDivider_v0p0p1_0.V5.t15 0.000502142
R23346 resistorDivider_v0p0p1_0.V5.n8 resistorDivider_v0p0p1_0.V5.t10 0.000502142
R23347 resistorDivider_v0p0p1_0.V5.n10 resistorDivider_v0p0p1_0.V5.t11 0.000502142
R23348 resistorDivider_v0p0p1_0.V5.n12 resistorDivider_v0p0p1_0.V5.t2 0.000502142
R23349 resistorDivider_v0p0p1_0.V5.n14 resistorDivider_v0p0p1_0.V5.t9 0.000502142
R23350 resistorDivider_v0p0p1_0.V5.n16 resistorDivider_v0p0p1_0.V5.t3 0.000502142
R23351 resistorDivider_v0p0p1_0.V5.n3 resistorDivider_v0p0p1_0.V5.t12 0.000502142
R23352 resistorDivider_v0p0p1_0.V5.n7 resistorDivider_v0p0p1_0.V5.t4 0.000502142
R23353 resistorDivider_v0p0p1_0.V5.n9 resistorDivider_v0p0p1_0.V5.t6 0.000502142
R23354 resistorDivider_v0p0p1_0.V5.n11 resistorDivider_v0p0p1_0.V5.t7 0.000502142
R23355 resistorDivider_v0p0p1_0.V5.n13 resistorDivider_v0p0p1_0.V5.t5 0.000502142
R23356 resistorDivider_v0p0p1_0.V5.n15 resistorDivider_v0p0p1_0.V5.t1 0.000502142
R23357 resistorDivider_v0p0p1_0.V5.n2 resistorDivider_v0p0p1_0.V5.t14 0.000502142
R23358 frontAnalog_v0p0p1_13.x63.A.n2 frontAnalog_v0p0p1_13.x63.A.t4 260.322
R23359 frontAnalog_v0p0p1_13.x63.A.n4 frontAnalog_v0p0p1_13.x63.A.t5 233.888
R23360 frontAnalog_v0p0p1_13.x63.A.n2 frontAnalog_v0p0p1_13.x63.A.t6 175.169
R23361 frontAnalog_v0p0p1_13.x63.A.n3 frontAnalog_v0p0p1_13.x63.A.t7 159.725
R23362 frontAnalog_v0p0p1_13.x63.A.n1 frontAnalog_v0p0p1_13.x63.A.t0 17.4109
R23363 frontAnalog_v0p0p1_13.x63.A.n0 frontAnalog_v0p0p1_13.x63.A.n2 9.75129
R23364 frontAnalog_v0p0p1_13.x63.A.n1 frontAnalog_v0p0p1_13.x63.A.t3 9.6037
R23365 frontAnalog_v0p0p1_13.x63.A.n0 frontAnalog_v0p0p1_13.x63.A 2.33338
R23366 frontAnalog_v0p0p1_13.x63.A.n5 frontAnalog_v0p0p1_13.x63.A.t1 8.40929
R23367 frontAnalog_v0p0p1_13.x63.A.n3 frontAnalog_v0p0p1_13.x63.A.t2 8.06629
R23368 frontAnalog_v0p0p1_13.x63.A.n4 frontAnalog_v0p0p1_13.x63.A.n3 1.73501
R23369 frontAnalog_v0p0p1_13.x63.A.n1 frontAnalog_v0p0p1_13.x63.A.n4 0.99025
R23370 frontAnalog_v0p0p1_13.x63.A.n5 frontAnalog_v0p0p1_13.x63.A.n1 0.853186
R23371 frontAnalog_v0p0p1_13.x63.A frontAnalog_v0p0p1_13.x63.A.n0 0.349517
R23372 frontAnalog_v0p0p1_13.x63.A frontAnalog_v0p0p1_13.x63.A.n5 0.24425
R23373 frontAnalog_v0p0p1_10.x63.A.n2 frontAnalog_v0p0p1_10.x63.A.t5 260.322
R23374 frontAnalog_v0p0p1_10.x63.A.n4 frontAnalog_v0p0p1_10.x63.A.t6 233.888
R23375 frontAnalog_v0p0p1_10.x63.A.n2 frontAnalog_v0p0p1_10.x63.A.t7 175.169
R23376 frontAnalog_v0p0p1_10.x63.A.n3 frontAnalog_v0p0p1_10.x63.A.t4 159.725
R23377 frontAnalog_v0p0p1_10.x63.A.n1 frontAnalog_v0p0p1_10.x63.A.t3 17.4109
R23378 frontAnalog_v0p0p1_10.x63.A.n0 frontAnalog_v0p0p1_10.x63.A.n2 9.75129
R23379 frontAnalog_v0p0p1_10.x63.A.n1 frontAnalog_v0p0p1_10.x63.A.t2 9.6037
R23380 frontAnalog_v0p0p1_10.x63.A.n0 frontAnalog_v0p0p1_10.x63.A 2.33338
R23381 frontAnalog_v0p0p1_10.x63.A.n5 frontAnalog_v0p0p1_10.x63.A.t1 8.40929
R23382 frontAnalog_v0p0p1_10.x63.A.n3 frontAnalog_v0p0p1_10.x63.A.t0 8.06629
R23383 frontAnalog_v0p0p1_10.x63.A.n4 frontAnalog_v0p0p1_10.x63.A.n3 1.73501
R23384 frontAnalog_v0p0p1_10.x63.A.n1 frontAnalog_v0p0p1_10.x63.A.n4 0.99025
R23385 frontAnalog_v0p0p1_10.x63.A.n5 frontAnalog_v0p0p1_10.x63.A.n1 0.853186
R23386 frontAnalog_v0p0p1_10.x63.A frontAnalog_v0p0p1_10.x63.A.n0 0.349517
R23387 frontAnalog_v0p0p1_10.x63.A frontAnalog_v0p0p1_10.x63.A.n5 0.24425
R23388 frontAnalog_v0p0p1_5.x63.A.n2 frontAnalog_v0p0p1_5.x63.A.t4 260.322
R23389 frontAnalog_v0p0p1_5.x63.A.n4 frontAnalog_v0p0p1_5.x63.A.t5 233.888
R23390 frontAnalog_v0p0p1_5.x63.A.n2 frontAnalog_v0p0p1_5.x63.A.t6 175.169
R23391 frontAnalog_v0p0p1_5.x63.A.n3 frontAnalog_v0p0p1_5.x63.A.t7 159.725
R23392 frontAnalog_v0p0p1_5.x63.A.n1 frontAnalog_v0p0p1_5.x63.A.t0 17.4109
R23393 frontAnalog_v0p0p1_5.x63.A.n0 frontAnalog_v0p0p1_5.x63.A.n2 9.75129
R23394 frontAnalog_v0p0p1_5.x63.A.n1 frontAnalog_v0p0p1_5.x63.A.t3 9.6037
R23395 frontAnalog_v0p0p1_5.x63.A.n0 frontAnalog_v0p0p1_5.x63.A 2.33338
R23396 frontAnalog_v0p0p1_5.x63.A.n5 frontAnalog_v0p0p1_5.x63.A.t1 8.40929
R23397 frontAnalog_v0p0p1_5.x63.A.n3 frontAnalog_v0p0p1_5.x63.A.t2 8.06629
R23398 frontAnalog_v0p0p1_5.x63.A.n4 frontAnalog_v0p0p1_5.x63.A.n3 1.73501
R23399 frontAnalog_v0p0p1_5.x63.A.n1 frontAnalog_v0p0p1_5.x63.A.n4 0.99025
R23400 frontAnalog_v0p0p1_5.x63.A.n5 frontAnalog_v0p0p1_5.x63.A.n1 0.853186
R23401 frontAnalog_v0p0p1_5.x63.A frontAnalog_v0p0p1_5.x63.A.n0 0.349517
R23402 frontAnalog_v0p0p1_5.x63.A frontAnalog_v0p0p1_5.x63.A.n5 0.24425
R23403 frontAnalog_v0p0p1_3.x63.A.n2 frontAnalog_v0p0p1_3.x63.A.t5 260.322
R23404 frontAnalog_v0p0p1_3.x63.A.n4 frontAnalog_v0p0p1_3.x63.A.t6 233.888
R23405 frontAnalog_v0p0p1_3.x63.A.n2 frontAnalog_v0p0p1_3.x63.A.t7 175.169
R23406 frontAnalog_v0p0p1_3.x63.A.n3 frontAnalog_v0p0p1_3.x63.A.t4 159.725
R23407 frontAnalog_v0p0p1_3.x63.A.n1 frontAnalog_v0p0p1_3.x63.A.t3 17.4109
R23408 frontAnalog_v0p0p1_3.x63.A.n0 frontAnalog_v0p0p1_3.x63.A.n2 9.75129
R23409 frontAnalog_v0p0p1_3.x63.A.n1 frontAnalog_v0p0p1_3.x63.A.t2 9.6037
R23410 frontAnalog_v0p0p1_3.x63.A.n0 frontAnalog_v0p0p1_3.x63.A 2.33338
R23411 frontAnalog_v0p0p1_3.x63.A.n5 frontAnalog_v0p0p1_3.x63.A.t1 8.40929
R23412 frontAnalog_v0p0p1_3.x63.A.n3 frontAnalog_v0p0p1_3.x63.A.t0 8.06629
R23413 frontAnalog_v0p0p1_3.x63.A.n4 frontAnalog_v0p0p1_3.x63.A.n3 1.73501
R23414 frontAnalog_v0p0p1_3.x63.A.n1 frontAnalog_v0p0p1_3.x63.A.n4 0.99025
R23415 frontAnalog_v0p0p1_3.x63.A.n5 frontAnalog_v0p0p1_3.x63.A.n1 0.853186
R23416 frontAnalog_v0p0p1_3.x63.A frontAnalog_v0p0p1_3.x63.A.n0 0.349517
R23417 frontAnalog_v0p0p1_3.x63.A frontAnalog_v0p0p1_3.x63.A.n5 0.24425
R23418 frontAnalog_v0p0p1_3.x65.A.n1 frontAnalog_v0p0p1_3.x65.A.t4 260.322
R23419 frontAnalog_v0p0p1_3.x65.A.n3 frontAnalog_v0p0p1_3.x65.A.t7 233.929
R23420 frontAnalog_v0p0p1_3.x65.A.n1 frontAnalog_v0p0p1_3.x65.A.t6 175.169
R23421 frontAnalog_v0p0p1_3.x65.A.n2 frontAnalog_v0p0p1_3.x65.A.t5 160.416
R23422 frontAnalog_v0p0p1_3.x65.A.n4 frontAnalog_v0p0p1_3.x65.A.t3 17.4109
R23423 frontAnalog_v0p0p1_3.x65.A.n4 frontAnalog_v0p0p1_3.x65.A.t2 10.2053
R23424 frontAnalog_v0p0p1_3.x65.A.n0 frontAnalog_v0p0p1_3.x65.A 2.78715
R23425 frontAnalog_v0p0p1_3.x65.A.n0 frontAnalog_v0p0p1_3.x65.A.n1 9.09103
R23426 frontAnalog_v0p0p1_3.x65.A.n6 frontAnalog_v0p0p1_3.x65.A.t0 7.94569
R23427 frontAnalog_v0p0p1_3.x65.A.n2 frontAnalog_v0p0p1_3.x65.A.t1 7.55846
R23428 frontAnalog_v0p0p1_3.x65.A.n5 frontAnalog_v0p0p1_3.x65.A.n3 1.4614
R23429 frontAnalog_v0p0p1_3.x65.A.n3 frontAnalog_v0p0p1_3.x65.A.n2 1.19626
R23430 frontAnalog_v0p0p1_3.x65.A.n6 frontAnalog_v0p0p1_3.x65.A.n5 0.836961
R23431 frontAnalog_v0p0p1_3.x65.A frontAnalog_v0p0p1_3.x65.A.n0 0.390342
R23432 frontAnalog_v0p0p1_3.x65.A.n5 frontAnalog_v0p0p1_3.x65.A.n4 0.154668
R23433 frontAnalog_v0p0p1_3.x65.A frontAnalog_v0p0p1_3.x65.A.n6 0.08175
R23434 frontAnalog_v0p0p1_15.x65.A.n1 frontAnalog_v0p0p1_15.x65.A.t4 260.322
R23435 frontAnalog_v0p0p1_15.x65.A.n3 frontAnalog_v0p0p1_15.x65.A.t7 233.929
R23436 frontAnalog_v0p0p1_15.x65.A.n1 frontAnalog_v0p0p1_15.x65.A.t6 175.169
R23437 frontAnalog_v0p0p1_15.x65.A.n2 frontAnalog_v0p0p1_15.x65.A.t5 160.416
R23438 frontAnalog_v0p0p1_15.x65.A.n4 frontAnalog_v0p0p1_15.x65.A.t0 17.4109
R23439 frontAnalog_v0p0p1_15.x65.A.n4 frontAnalog_v0p0p1_15.x65.A.t1 10.2053
R23440 frontAnalog_v0p0p1_15.x65.A.n0 frontAnalog_v0p0p1_15.x65.A 2.78715
R23441 frontAnalog_v0p0p1_15.x65.A.n0 frontAnalog_v0p0p1_15.x65.A.n1 9.09103
R23442 frontAnalog_v0p0p1_15.x65.A.n6 frontAnalog_v0p0p1_15.x65.A.t3 7.94569
R23443 frontAnalog_v0p0p1_15.x65.A.n2 frontAnalog_v0p0p1_15.x65.A.t2 7.55846
R23444 frontAnalog_v0p0p1_15.x65.A.n5 frontAnalog_v0p0p1_15.x65.A.n3 1.4614
R23445 frontAnalog_v0p0p1_15.x65.A.n3 frontAnalog_v0p0p1_15.x65.A.n2 1.19626
R23446 frontAnalog_v0p0p1_15.x65.A.n6 frontAnalog_v0p0p1_15.x65.A.n5 0.836961
R23447 frontAnalog_v0p0p1_15.x65.A frontAnalog_v0p0p1_15.x65.A.n0 0.390342
R23448 frontAnalog_v0p0p1_15.x65.A.n5 frontAnalog_v0p0p1_15.x65.A.n4 0.154668
R23449 frontAnalog_v0p0p1_15.x65.A frontAnalog_v0p0p1_15.x65.A.n6 0.08175
R23450 frontAnalog_v0p0p1_4.x63.A.n2 frontAnalog_v0p0p1_4.x63.A.t6 260.322
R23451 frontAnalog_v0p0p1_4.x63.A.n4 frontAnalog_v0p0p1_4.x63.A.t4 233.888
R23452 frontAnalog_v0p0p1_4.x63.A.n2 frontAnalog_v0p0p1_4.x63.A.t5 175.169
R23453 frontAnalog_v0p0p1_4.x63.A.n3 frontAnalog_v0p0p1_4.x63.A.t7 159.725
R23454 frontAnalog_v0p0p1_4.x63.A.n1 frontAnalog_v0p0p1_4.x63.A.t0 17.4109
R23455 frontAnalog_v0p0p1_4.x63.A.n0 frontAnalog_v0p0p1_4.x63.A.n2 9.75129
R23456 frontAnalog_v0p0p1_4.x63.A.n1 frontAnalog_v0p0p1_4.x63.A.t1 9.6027
R23457 frontAnalog_v0p0p1_4.x63.A.n0 frontAnalog_v0p0p1_4.x63.A 2.33338
R23458 frontAnalog_v0p0p1_4.x63.A.n5 frontAnalog_v0p0p1_4.x63.A.t2 8.40929
R23459 frontAnalog_v0p0p1_4.x63.A.n3 frontAnalog_v0p0p1_4.x63.A.t3 8.06629
R23460 frontAnalog_v0p0p1_4.x63.A.n4 frontAnalog_v0p0p1_4.x63.A.n3 1.73501
R23461 frontAnalog_v0p0p1_4.x63.A.n1 frontAnalog_v0p0p1_4.x63.A.n4 0.99025
R23462 frontAnalog_v0p0p1_4.x63.A.n5 frontAnalog_v0p0p1_4.x63.A.n1 0.853186
R23463 frontAnalog_v0p0p1_4.x63.A frontAnalog_v0p0p1_4.x63.A.n0 0.349517
R23464 frontAnalog_v0p0p1_4.x63.A frontAnalog_v0p0p1_4.x63.A.n5 0.24425
R23465 frontAnalog_v0p0p1_1.x65.A.n1 frontAnalog_v0p0p1_1.x65.A.t4 260.322
R23466 frontAnalog_v0p0p1_1.x65.A.n3 frontAnalog_v0p0p1_1.x65.A.t7 233.929
R23467 frontAnalog_v0p0p1_1.x65.A.n1 frontAnalog_v0p0p1_1.x65.A.t6 175.169
R23468 frontAnalog_v0p0p1_1.x65.A.n2 frontAnalog_v0p0p1_1.x65.A.t5 160.416
R23469 frontAnalog_v0p0p1_1.x65.A.n4 frontAnalog_v0p0p1_1.x65.A.t2 17.4109
R23470 frontAnalog_v0p0p1_1.x65.A.n4 frontAnalog_v0p0p1_1.x65.A.t3 10.2053
R23471 frontAnalog_v0p0p1_1.x65.A.n0 frontAnalog_v0p0p1_1.x65.A 2.78715
R23472 frontAnalog_v0p0p1_1.x65.A.n0 frontAnalog_v0p0p1_1.x65.A.n1 9.09103
R23473 frontAnalog_v0p0p1_1.x65.A.n6 frontAnalog_v0p0p1_1.x65.A.t0 7.94569
R23474 frontAnalog_v0p0p1_1.x65.A.n2 frontAnalog_v0p0p1_1.x65.A.t1 7.55846
R23475 frontAnalog_v0p0p1_1.x65.A.n5 frontAnalog_v0p0p1_1.x65.A.n3 1.4614
R23476 frontAnalog_v0p0p1_1.x65.A.n3 frontAnalog_v0p0p1_1.x65.A.n2 1.19626
R23477 frontAnalog_v0p0p1_1.x65.A.n6 frontAnalog_v0p0p1_1.x65.A.n5 0.836961
R23478 frontAnalog_v0p0p1_1.x65.A frontAnalog_v0p0p1_1.x65.A.n0 0.390342
R23479 frontAnalog_v0p0p1_1.x65.A.n5 frontAnalog_v0p0p1_1.x65.A.n4 0.154668
R23480 frontAnalog_v0p0p1_1.x65.A frontAnalog_v0p0p1_1.x65.A.n6 0.08175
R23481 frontAnalog_v0p0p1_10.RSfetsym_0.QN.n1 frontAnalog_v0p0p1_10.RSfetsym_0.QN.t6 117.511
R23482 frontAnalog_v0p0p1_10.RSfetsym_0.QN.n1 frontAnalog_v0p0p1_10.RSfetsym_0.QN.t5 110.698
R23483 frontAnalog_v0p0p1_10.RSfetsym_0.QN.n4 frontAnalog_v0p0p1_10.RSfetsym_0.QN.t1 19.1963
R23484 frontAnalog_v0p0p1_10.RSfetsym_0.QN.n7 frontAnalog_v0p0p1_10.RSfetsym_0.QN.t0 14.2842
R23485 frontAnalog_v0p0p1_10.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_10.RSfetsym_0.QN.t2 14.283
R23486 frontAnalog_v0p0p1_10.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_10.RSfetsym_0.QN.t3 14.283
R23487 frontAnalog_v0p0p1_10.RSfetsym_0.QN.n11 frontAnalog_v0p0p1_10.RSfetsym_0.QN.t4 9.14075
R23488 frontAnalog_v0p0p1_10.RSfetsym_0.QN.n11 frontAnalog_v0p0p1_10.RSfetsym_0.QN.n10 0.74645
R23489 frontAnalog_v0p0p1_10.RSfetsym_0.QN.n2 frontAnalog_v0p0p1_10.RSfetsym_0.QN.n1 0.688382
R23490 frontAnalog_v0p0p1_10.RSfetsym_0.QN.n10 frontAnalog_v0p0p1_10.RSfetsym_0.QN.n9 0.2402
R23491 frontAnalog_v0p0p1_10.RSfetsym_0.QN.n9 frontAnalog_v0p0p1_10.RSfetsym_0.QN.n8 0.236824
R23492 frontAnalog_v0p0p1_10.RSfetsym_0.QN.n4 frontAnalog_v0p0p1_10.RSfetsym_0.QN.n3 0.132187
R23493 frontAnalog_v0p0p1_10.RSfetsym_0.QN.n9 frontAnalog_v0p0p1_10.RSfetsym_0.QN.n4 0.0968646
R23494 frontAnalog_v0p0p1_10.RSfetsym_0.QN frontAnalog_v0p0p1_10.RSfetsym_0.QN.n11 0.0446535
R23495 frontAnalog_v0p0p1_10.RSfetsym_0.QN.n8 frontAnalog_v0p0p1_10.RSfetsym_0.QN.n6 0.0272538
R23496 frontAnalog_v0p0p1_10.RSfetsym_0.QN.n10 frontAnalog_v0p0p1_10.RSfetsym_0.QN.n0 0.00981499
R23497 frontAnalog_v0p0p1_10.RSfetsym_0.QN.n3 frontAnalog_v0p0p1_10.RSfetsym_0.QN.n2 0.00725433
R23498 frontAnalog_v0p0p1_10.RSfetsym_0.QN.n6 frontAnalog_v0p0p1_10.RSfetsym_0.QN.n5 0.00610579
R23499 frontAnalog_v0p0p1_10.RSfetsym_0.QN.n8 frontAnalog_v0p0p1_10.RSfetsym_0.QN.n7 0.00225341
R23500 frontAnalog_v0p0p1_11.Q.n2 frontAnalog_v0p0p1_11.Q.t5 260.435
R23501 frontAnalog_v0p0p1_11.Q.n7 frontAnalog_v0p0p1_11.Q.t11 230.576
R23502 frontAnalog_v0p0p1_11.Q.n10 frontAnalog_v0p0p1_11.Q.t7 196.549
R23503 frontAnalog_v0p0p1_11.Q.n7 frontAnalog_v0p0p1_11.Q.t8 158.275
R23504 frontAnalog_v0p0p1_11.Q.n2 frontAnalog_v0p0p1_11.Q.t10 156.403
R23505 frontAnalog_v0p0p1_11.Q.n10 frontAnalog_v0p0p1_11.Q.t9 148.35
R23506 frontAnalog_v0p0p1_11.Q.n15 frontAnalog_v0p0p1_11.Q.t6 117.314
R23507 frontAnalog_v0p0p1_11.Q.n15 frontAnalog_v0p0p1_11.Q.t12 110.853
R23508 frontAnalog_v0p0p1_11.Q.n16 frontAnalog_v0p0p1_11.Q.t0 17.6181
R23509 frontAnalog_v0p0p1_11.Q.n18 frontAnalog_v0p0p1_11.Q.t3 14.2865
R23510 frontAnalog_v0p0p1_11.Q.n20 frontAnalog_v0p0p1_11.Q.t2 14.283
R23511 frontAnalog_v0p0p1_11.Q.n20 frontAnalog_v0p0p1_11.Q.t1 14.283
R23512 frontAnalog_v0p0p1_11.Q.n11 frontAnalog_v0p0p1_11.Q.n10 9.49829
R23513 frontAnalog_v0p0p1_11.Q frontAnalog_v0p0p1_11.Q.n1 9.3005
R23514 frontAnalog_v0p0p1_11.Q.n22 frontAnalog_v0p0p1_11.Q.t4 8.77744
R23515 frontAnalog_v0p0p1_11.Q.n8 frontAnalog_v0p0p1_11.Q.n7 8.76429
R23516 frontAnalog_v0p0p1_11.Q.n12 frontAnalog_v0p0p1_11.Q.n11 7.9582
R23517 frontAnalog_v0p0p1_11.Q.n9 frontAnalog_v0p0p1_11.Q.n8 7.74345
R23518 frontAnalog_v0p0p1_11.Q.n3 frontAnalog_v0p0p1_11.Q.n2 7.60183
R23519 frontAnalog_v0p0p1_11.Q.n8 frontAnalog_v0p0p1_11.Q 6.66717
R23520 frontAnalog_v0p0p1_11.Q.n11 frontAnalog_v0p0p1_11.Q 6.44139
R23521 frontAnalog_v0p0p1_11.Q.n23 frontAnalog_v0p0p1_11.Q.n14 5.49051
R23522 frontAnalog_v0p0p1_11.Q.n3 frontAnalog_v0p0p1_11.Q 4.8645
R23523 frontAnalog_v0p0p1_11.Q.n13 frontAnalog_v0p0p1_11.Q.n6 2.33148
R23524 frontAnalog_v0p0p1_11.Q.n22 frontAnalog_v0p0p1_11.Q.n21 1.20426
R23525 frontAnalog_v0p0p1_11.Q.n12 frontAnalog_v0p0p1_11.Q.n9 1.0005
R23526 frontAnalog_v0p0p1_11.Q.n13 frontAnalog_v0p0p1_11.Q.n12 0.446956
R23527 frontAnalog_v0p0p1_11.Q.n9 frontAnalog_v0p0p1_11.Q 0.380411
R23528 frontAnalog_v0p0p1_11.Q.n14 frontAnalog_v0p0p1_11.Q.n13 0.368862
R23529 frontAnalog_v0p0p1_11.Q.n23 frontAnalog_v0p0p1_11.Q.n22 0.325111
R23530 frontAnalog_v0p0p1_11.Q.n19 frontAnalog_v0p0p1_11.Q.n18 0.301242
R23531 frontAnalog_v0p0p1_11.Q.n14 frontAnalog_v0p0p1_11.Q 0.20675
R23532 frontAnalog_v0p0p1_11.Q.n17 frontAnalog_v0p0p1_11.Q.n15 0.159555
R23533 frontAnalog_v0p0p1_11.Q.n21 frontAnalog_v0p0p1_11.Q.n20 0.106617
R23534 frontAnalog_v0p0p1_11.Q.n19 frontAnalog_v0p0p1_11.Q.n17 0.0796167
R23535 frontAnalog_v0p0p1_11.Q.n21 frontAnalog_v0p0p1_11.Q.n19 0.0480595
R23536 frontAnalog_v0p0p1_11.Q frontAnalog_v0p0p1_11.Q.n23 0.0469368
R23537 frontAnalog_v0p0p1_11.Q.n5 frontAnalog_v0p0p1_11.Q.n1 0.0344286
R23538 frontAnalog_v0p0p1_11.Q.n6 frontAnalog_v0p0p1_11.Q.n0 0.00182856
R23539 frontAnalog_v0p0p1_11.Q.n6 frontAnalog_v0p0p1_11.Q.n5 0.00149885
R23540 frontAnalog_v0p0p1_11.Q.n4 frontAnalog_v0p0p1_11.Q.n3 0.00133362
R23541 frontAnalog_v0p0p1_11.Q.n5 frontAnalog_v0p0p1_11.Q.n4 0.00100077
R23542 frontAnalog_v0p0p1_11.Q.n17 frontAnalog_v0p0p1_11.Q.n16 0.000504658
R23543 frontAnalog_v0p0p1_3.RSfetsym_0.QN.n1 frontAnalog_v0p0p1_3.RSfetsym_0.QN.t6 117.511
R23544 frontAnalog_v0p0p1_3.RSfetsym_0.QN.n1 frontAnalog_v0p0p1_3.RSfetsym_0.QN.t5 110.698
R23545 frontAnalog_v0p0p1_3.RSfetsym_0.QN.n4 frontAnalog_v0p0p1_3.RSfetsym_0.QN.t1 19.1963
R23546 frontAnalog_v0p0p1_3.RSfetsym_0.QN.n7 frontAnalog_v0p0p1_3.RSfetsym_0.QN.t4 14.2842
R23547 frontAnalog_v0p0p1_3.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_3.RSfetsym_0.QN.t2 14.283
R23548 frontAnalog_v0p0p1_3.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_3.RSfetsym_0.QN.t3 14.283
R23549 frontAnalog_v0p0p1_3.RSfetsym_0.QN.n11 frontAnalog_v0p0p1_3.RSfetsym_0.QN.t0 9.14075
R23550 frontAnalog_v0p0p1_3.RSfetsym_0.QN.n11 frontAnalog_v0p0p1_3.RSfetsym_0.QN.n10 0.74645
R23551 frontAnalog_v0p0p1_3.RSfetsym_0.QN.n2 frontAnalog_v0p0p1_3.RSfetsym_0.QN.n1 0.688382
R23552 frontAnalog_v0p0p1_3.RSfetsym_0.QN.n10 frontAnalog_v0p0p1_3.RSfetsym_0.QN.n9 0.2402
R23553 frontAnalog_v0p0p1_3.RSfetsym_0.QN.n9 frontAnalog_v0p0p1_3.RSfetsym_0.QN.n8 0.236824
R23554 frontAnalog_v0p0p1_3.RSfetsym_0.QN.n4 frontAnalog_v0p0p1_3.RSfetsym_0.QN.n3 0.132187
R23555 frontAnalog_v0p0p1_3.RSfetsym_0.QN.n9 frontAnalog_v0p0p1_3.RSfetsym_0.QN.n4 0.0968646
R23556 frontAnalog_v0p0p1_3.RSfetsym_0.QN frontAnalog_v0p0p1_3.RSfetsym_0.QN.n11 0.0446535
R23557 frontAnalog_v0p0p1_3.RSfetsym_0.QN.n8 frontAnalog_v0p0p1_3.RSfetsym_0.QN.n6 0.0272538
R23558 frontAnalog_v0p0p1_3.RSfetsym_0.QN.n10 frontAnalog_v0p0p1_3.RSfetsym_0.QN.n0 0.00981499
R23559 frontAnalog_v0p0p1_3.RSfetsym_0.QN.n3 frontAnalog_v0p0p1_3.RSfetsym_0.QN.n2 0.00725433
R23560 frontAnalog_v0p0p1_3.RSfetsym_0.QN.n6 frontAnalog_v0p0p1_3.RSfetsym_0.QN.n5 0.00610579
R23561 frontAnalog_v0p0p1_3.RSfetsym_0.QN.n8 frontAnalog_v0p0p1_3.RSfetsym_0.QN.n7 0.00225341
R23562 frontAnalog_v0p0p1_6.x63.A.n2 frontAnalog_v0p0p1_6.x63.A.t4 260.322
R23563 frontAnalog_v0p0p1_6.x63.A.n4 frontAnalog_v0p0p1_6.x63.A.t7 233.888
R23564 frontAnalog_v0p0p1_6.x63.A.n2 frontAnalog_v0p0p1_6.x63.A.t6 175.169
R23565 frontAnalog_v0p0p1_6.x63.A.n3 frontAnalog_v0p0p1_6.x63.A.t5 159.725
R23566 frontAnalog_v0p0p1_6.x63.A.n1 frontAnalog_v0p0p1_6.x63.A.t1 17.4109
R23567 frontAnalog_v0p0p1_6.x63.A.n0 frontAnalog_v0p0p1_6.x63.A.n2 9.75129
R23568 frontAnalog_v0p0p1_6.x63.A.n1 frontAnalog_v0p0p1_6.x63.A.t0 9.6027
R23569 frontAnalog_v0p0p1_6.x63.A.n0 frontAnalog_v0p0p1_6.x63.A 2.33338
R23570 frontAnalog_v0p0p1_6.x63.A.n5 frontAnalog_v0p0p1_6.x63.A.t2 8.40929
R23571 frontAnalog_v0p0p1_6.x63.A.n3 frontAnalog_v0p0p1_6.x63.A.t3 8.06629
R23572 frontAnalog_v0p0p1_6.x63.A.n4 frontAnalog_v0p0p1_6.x63.A.n3 1.73501
R23573 frontAnalog_v0p0p1_6.x63.A.n1 frontAnalog_v0p0p1_6.x63.A.n4 0.99025
R23574 frontAnalog_v0p0p1_6.x63.A.n5 frontAnalog_v0p0p1_6.x63.A.n1 0.853186
R23575 frontAnalog_v0p0p1_6.x63.A frontAnalog_v0p0p1_6.x63.A.n0 0.349517
R23576 frontAnalog_v0p0p1_6.x63.A frontAnalog_v0p0p1_6.x63.A.n5 0.24425
R23577 frontAnalog_v0p0p1_12.RSfetsym_0.QN.n1 frontAnalog_v0p0p1_12.RSfetsym_0.QN.t6 117.511
R23578 frontAnalog_v0p0p1_12.RSfetsym_0.QN.n1 frontAnalog_v0p0p1_12.RSfetsym_0.QN.t5 110.698
R23579 frontAnalog_v0p0p1_12.RSfetsym_0.QN.n4 frontAnalog_v0p0p1_12.RSfetsym_0.QN.t2 19.1963
R23580 frontAnalog_v0p0p1_12.RSfetsym_0.QN.n7 frontAnalog_v0p0p1_12.RSfetsym_0.QN.t3 14.2842
R23581 frontAnalog_v0p0p1_12.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_12.RSfetsym_0.QN.t1 14.283
R23582 frontAnalog_v0p0p1_12.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_12.RSfetsym_0.QN.t0 14.283
R23583 frontAnalog_v0p0p1_12.RSfetsym_0.QN.n11 frontAnalog_v0p0p1_12.RSfetsym_0.QN.t4 9.14075
R23584 frontAnalog_v0p0p1_12.RSfetsym_0.QN.n11 frontAnalog_v0p0p1_12.RSfetsym_0.QN.n10 0.74645
R23585 frontAnalog_v0p0p1_12.RSfetsym_0.QN.n2 frontAnalog_v0p0p1_12.RSfetsym_0.QN.n1 0.688382
R23586 frontAnalog_v0p0p1_12.RSfetsym_0.QN.n10 frontAnalog_v0p0p1_12.RSfetsym_0.QN.n9 0.2402
R23587 frontAnalog_v0p0p1_12.RSfetsym_0.QN.n9 frontAnalog_v0p0p1_12.RSfetsym_0.QN.n8 0.236824
R23588 frontAnalog_v0p0p1_12.RSfetsym_0.QN.n4 frontAnalog_v0p0p1_12.RSfetsym_0.QN.n3 0.132187
R23589 frontAnalog_v0p0p1_12.RSfetsym_0.QN.n9 frontAnalog_v0p0p1_12.RSfetsym_0.QN.n4 0.0968646
R23590 frontAnalog_v0p0p1_12.RSfetsym_0.QN frontAnalog_v0p0p1_12.RSfetsym_0.QN.n11 0.0446535
R23591 frontAnalog_v0p0p1_12.RSfetsym_0.QN.n8 frontAnalog_v0p0p1_12.RSfetsym_0.QN.n6 0.0272538
R23592 frontAnalog_v0p0p1_12.RSfetsym_0.QN.n10 frontAnalog_v0p0p1_12.RSfetsym_0.QN.n0 0.00981499
R23593 frontAnalog_v0p0p1_12.RSfetsym_0.QN.n3 frontAnalog_v0p0p1_12.RSfetsym_0.QN.n2 0.00725433
R23594 frontAnalog_v0p0p1_12.RSfetsym_0.QN.n6 frontAnalog_v0p0p1_12.RSfetsym_0.QN.n5 0.00610579
R23595 frontAnalog_v0p0p1_12.RSfetsym_0.QN.n8 frontAnalog_v0p0p1_12.RSfetsym_0.QN.n7 0.00225341
R23596 VL.n6 VL 0.23241
R23597 VL.n3 VL.t4 0.0203551
R23598 VL.n0 VL.t0 0.0203551
R23599 VL.n1 VL.n0 0.0203529
R23600 VL.n2 VL.n1 0.0203529
R23601 VL.n5 VL.n4 0.0203529
R23602 VL.n4 VL.n3 0.0203529
R23603 VL VL.n2 0.0111618
R23604 VL VL.n6 0.00913171
R23605 VL.n6 VL.n5 0.00105946
R23606 VL.n3 VL.t3 0.000502142
R23607 VL.n4 VL.t1 0.000502142
R23608 VL.n5 VL.t2 0.000502142
R23609 VL.n2 VL.t7 0.000502142
R23610 VL.n1 VL.t6 0.000502142
R23611 VL.n0 VL.t5 0.000502142
R23612 frontAnalog_v0p0p1_11.x65.A.n1 frontAnalog_v0p0p1_11.x65.A.t4 260.322
R23613 frontAnalog_v0p0p1_11.x65.A.n3 frontAnalog_v0p0p1_11.x65.A.t7 233.929
R23614 frontAnalog_v0p0p1_11.x65.A.n1 frontAnalog_v0p0p1_11.x65.A.t6 175.169
R23615 frontAnalog_v0p0p1_11.x65.A.n2 frontAnalog_v0p0p1_11.x65.A.t5 160.416
R23616 frontAnalog_v0p0p1_11.x65.A.n4 frontAnalog_v0p0p1_11.x65.A.t3 17.4109
R23617 frontAnalog_v0p0p1_11.x65.A.n4 frontAnalog_v0p0p1_11.x65.A.t0 10.2053
R23618 frontAnalog_v0p0p1_11.x65.A.n0 frontAnalog_v0p0p1_11.x65.A 2.78715
R23619 frontAnalog_v0p0p1_11.x65.A.n0 frontAnalog_v0p0p1_11.x65.A.n1 9.09103
R23620 frontAnalog_v0p0p1_11.x65.A.n6 frontAnalog_v0p0p1_11.x65.A.t1 7.94569
R23621 frontAnalog_v0p0p1_11.x65.A.n2 frontAnalog_v0p0p1_11.x65.A.t2 7.55846
R23622 frontAnalog_v0p0p1_11.x65.A.n5 frontAnalog_v0p0p1_11.x65.A.n3 1.4614
R23623 frontAnalog_v0p0p1_11.x65.A.n3 frontAnalog_v0p0p1_11.x65.A.n2 1.19626
R23624 frontAnalog_v0p0p1_11.x65.A.n6 frontAnalog_v0p0p1_11.x65.A.n5 0.836961
R23625 frontAnalog_v0p0p1_11.x65.A frontAnalog_v0p0p1_11.x65.A.n0 0.390342
R23626 frontAnalog_v0p0p1_11.x65.A.n5 frontAnalog_v0p0p1_11.x65.A.n4 0.154668
R23627 frontAnalog_v0p0p1_11.x65.A frontAnalog_v0p0p1_11.x65.A.n6 0.08175
R23628 resistorDivider_v0p0p1_0.V8.n0 resistorDivider_v0p0p1_0.V8.t17 167.365
R23629 resistorDivider_v0p0p1_0.V8.n0 resistorDivider_v0p0p1_0.V8.t16 92.4488
R23630 resistorDivider_v0p0p1_0.V8.n1 resistorDivider_v0p0p1_0.V8.n0 2.07493
R23631 resistorDivider_v0p0p1_0.V8.n9 resistorDivider_v0p0p1_0.V8.n8 0.141636
R23632 resistorDivider_v0p0p1_0.V8.n8 resistorDivider_v0p0p1_0.V8.n7 0.141636
R23633 resistorDivider_v0p0p1_0.V8.n7 resistorDivider_v0p0p1_0.V8.n6 0.141636
R23634 resistorDivider_v0p0p1_0.V8.n6 resistorDivider_v0p0p1_0.V8.n5 0.141636
R23635 resistorDivider_v0p0p1_0.V8.n5 resistorDivider_v0p0p1_0.V8.n4 0.141636
R23636 resistorDivider_v0p0p1_0.V8.n4 resistorDivider_v0p0p1_0.V8.n3 0.141636
R23637 resistorDivider_v0p0p1_0.V8.n3 resistorDivider_v0p0p1_0.V8.n2 0.141636
R23638 resistorDivider_v0p0p1_0.V8.n1 resistorDivider_v0p0p1_0.V8 0.12425
R23639 resistorDivider_v0p0p1_0.V8 resistorDivider_v0p0p1_0.V8.n9 0.100159
R23640 resistorDivider_v0p0p1_0.V8 resistorDivider_v0p0p1_0.V8.n1 0.0314375
R23641 resistorDivider_v0p0p1_0.V8.n9 resistorDivider_v0p0p1_0.V8.t0 0.00250214
R23642 resistorDivider_v0p0p1_0.V8.n3 resistorDivider_v0p0p1_0.V8.t8 0.000502142
R23643 resistorDivider_v0p0p1_0.V8.n4 resistorDivider_v0p0p1_0.V8.t14 0.000502142
R23644 resistorDivider_v0p0p1_0.V8.n5 resistorDivider_v0p0p1_0.V8.t7 0.000502142
R23645 resistorDivider_v0p0p1_0.V8.n6 resistorDivider_v0p0p1_0.V8.t11 0.000502142
R23646 resistorDivider_v0p0p1_0.V8.n7 resistorDivider_v0p0p1_0.V8.t12 0.000502142
R23647 resistorDivider_v0p0p1_0.V8.n8 resistorDivider_v0p0p1_0.V8.t13 0.000502142
R23648 resistorDivider_v0p0p1_0.V8.n9 resistorDivider_v0p0p1_0.V8.t2 0.000502142
R23649 resistorDivider_v0p0p1_0.V8.n2 resistorDivider_v0p0p1_0.V8.t4 0.000502142
R23650 resistorDivider_v0p0p1_0.V8.n3 resistorDivider_v0p0p1_0.V8.t3 0.000502142
R23651 resistorDivider_v0p0p1_0.V8.n4 resistorDivider_v0p0p1_0.V8.t10 0.000502142
R23652 resistorDivider_v0p0p1_0.V8.n5 resistorDivider_v0p0p1_0.V8.t6 0.000502142
R23653 resistorDivider_v0p0p1_0.V8.n6 resistorDivider_v0p0p1_0.V8.t1 0.000502142
R23654 resistorDivider_v0p0p1_0.V8.n7 resistorDivider_v0p0p1_0.V8.t15 0.000502142
R23655 resistorDivider_v0p0p1_0.V8.n8 resistorDivider_v0p0p1_0.V8.t5 0.000502142
R23656 resistorDivider_v0p0p1_0.V8.n2 resistorDivider_v0p0p1_0.V8.t9 0.000502142
R23657 16to4_PriorityEncoder_v0p0p1_0.I12.n10 16to4_PriorityEncoder_v0p0p1_0.I12.t11 260.435
R23658 16to4_PriorityEncoder_v0p0p1_0.I12.n15 16to4_PriorityEncoder_v0p0p1_0.I12.t12 230.576
R23659 16to4_PriorityEncoder_v0p0p1_0.I12.n18 16to4_PriorityEncoder_v0p0p1_0.I12.t6 196.549
R23660 16to4_PriorityEncoder_v0p0p1_0.I12.n15 16to4_PriorityEncoder_v0p0p1_0.I12.t9 158.275
R23661 16to4_PriorityEncoder_v0p0p1_0.I12.n10 16to4_PriorityEncoder_v0p0p1_0.I12.t8 156.403
R23662 16to4_PriorityEncoder_v0p0p1_0.I12.n18 16to4_PriorityEncoder_v0p0p1_0.I12.t5 148.35
R23663 16to4_PriorityEncoder_v0p0p1_0.I12.n0 16to4_PriorityEncoder_v0p0p1_0.I12.t10 117.314
R23664 16to4_PriorityEncoder_v0p0p1_0.I12.n0 16to4_PriorityEncoder_v0p0p1_0.I12.t7 110.852
R23665 16to4_PriorityEncoder_v0p0p1_0.I12.n1 16to4_PriorityEncoder_v0p0p1_0.I12.t2 17.6181
R23666 16to4_PriorityEncoder_v0p0p1_0.I12.n3 16to4_PriorityEncoder_v0p0p1_0.I12.t4 14.2865
R23667 16to4_PriorityEncoder_v0p0p1_0.I12.n5 16to4_PriorityEncoder_v0p0p1_0.I12.t1 14.283
R23668 16to4_PriorityEncoder_v0p0p1_0.I12.n5 16to4_PriorityEncoder_v0p0p1_0.I12.t0 14.283
R23669 16to4_PriorityEncoder_v0p0p1_0.I12.n19 16to4_PriorityEncoder_v0p0p1_0.I12.n18 9.49829
R23670 16to4_PriorityEncoder_v0p0p1_0.I12 16to4_PriorityEncoder_v0p0p1_0.I12.n9 9.3005
R23671 16to4_PriorityEncoder_v0p0p1_0.I12.n7 16to4_PriorityEncoder_v0p0p1_0.I12.t3 8.77592
R23672 16to4_PriorityEncoder_v0p0p1_0.I12.n16 16to4_PriorityEncoder_v0p0p1_0.I12.n15 8.76429
R23673 16to4_PriorityEncoder_v0p0p1_0.I12.n20 16to4_PriorityEncoder_v0p0p1_0.I12.n19 7.9582
R23674 16to4_PriorityEncoder_v0p0p1_0.I12.n17 16to4_PriorityEncoder_v0p0p1_0.I12.n16 7.74345
R23675 16to4_PriorityEncoder_v0p0p1_0.I12.n11 16to4_PriorityEncoder_v0p0p1_0.I12.n10 7.60183
R23676 16to4_PriorityEncoder_v0p0p1_0.I12.n16 16to4_PriorityEncoder_v0p0p1_0.I12 6.66717
R23677 16to4_PriorityEncoder_v0p0p1_0.I12.n19 16to4_PriorityEncoder_v0p0p1_0.I12 6.44139
R23678 16to4_PriorityEncoder_v0p0p1_0.I12.n23 16to4_PriorityEncoder_v0p0p1_0.I12.n22 5.87984
R23679 16to4_PriorityEncoder_v0p0p1_0.I12.n11 16to4_PriorityEncoder_v0p0p1_0.I12 4.8645
R23680 16to4_PriorityEncoder_v0p0p1_0.I12.n21 16to4_PriorityEncoder_v0p0p1_0.I12.n14 2.33638
R23681 16to4_PriorityEncoder_v0p0p1_0.I12.n7 16to4_PriorityEncoder_v0p0p1_0.I12.n6 1.20426
R23682 16to4_PriorityEncoder_v0p0p1_0.I12.n20 16to4_PriorityEncoder_v0p0p1_0.I12.n17 1.0005
R23683 16to4_PriorityEncoder_v0p0p1_0.I12.n21 16to4_PriorityEncoder_v0p0p1_0.I12.n20 0.446956
R23684 16to4_PriorityEncoder_v0p0p1_0.I12.n22 16to4_PriorityEncoder_v0p0p1_0.I12.n21 0.385117
R23685 16to4_PriorityEncoder_v0p0p1_0.I12.n17 16to4_PriorityEncoder_v0p0p1_0.I12 0.380411
R23686 16to4_PriorityEncoder_v0p0p1_0.I12.n23 16to4_PriorityEncoder_v0p0p1_0.I12.n7 0.336084
R23687 16to4_PriorityEncoder_v0p0p1_0.I12.n4 16to4_PriorityEncoder_v0p0p1_0.I12.n3 0.300242
R23688 16to4_PriorityEncoder_v0p0p1_0.I12.n22 16to4_PriorityEncoder_v0p0p1_0.I12 0.2005
R23689 16to4_PriorityEncoder_v0p0p1_0.I12.n2 16to4_PriorityEncoder_v0p0p1_0.I12.n0 0.159555
R23690 16to4_PriorityEncoder_v0p0p1_0.I12.n6 16to4_PriorityEncoder_v0p0p1_0.I12.n5 0.106617
R23691 16to4_PriorityEncoder_v0p0p1_0.I12.n4 16to4_PriorityEncoder_v0p0p1_0.I12.n2 0.0796167
R23692 16to4_PriorityEncoder_v0p0p1_0.I12.n6 16to4_PriorityEncoder_v0p0p1_0.I12.n4 0.0480595
R23693 16to4_PriorityEncoder_v0p0p1_0.I12.n13 16to4_PriorityEncoder_v0p0p1_0.I12.n9 0.0344286
R23694 16to4_PriorityEncoder_v0p0p1_0.I12 16to4_PriorityEncoder_v0p0p1_0.I12.n23 0.00658123
R23695 16to4_PriorityEncoder_v0p0p1_0.I12.n14 16to4_PriorityEncoder_v0p0p1_0.I12.n8 0.00182856
R23696 16to4_PriorityEncoder_v0p0p1_0.I12.n14 16to4_PriorityEncoder_v0p0p1_0.I12.n13 0.00149885
R23697 16to4_PriorityEncoder_v0p0p1_0.I12.n12 16to4_PriorityEncoder_v0p0p1_0.I12.n11 0.00133362
R23698 16to4_PriorityEncoder_v0p0p1_0.I12.n13 16to4_PriorityEncoder_v0p0p1_0.I12.n12 0.00100077
R23699 16to4_PriorityEncoder_v0p0p1_0.I12.n2 16to4_PriorityEncoder_v0p0p1_0.I12.n1 0.000504658
R23700 frontAnalog_v0p0p1_1.x63.A.n2 frontAnalog_v0p0p1_1.x63.A.t7 260.322
R23701 frontAnalog_v0p0p1_1.x63.A.n4 frontAnalog_v0p0p1_1.x63.A.t4 233.888
R23702 frontAnalog_v0p0p1_1.x63.A.n2 frontAnalog_v0p0p1_1.x63.A.t6 175.169
R23703 frontAnalog_v0p0p1_1.x63.A.n3 frontAnalog_v0p0p1_1.x63.A.t5 159.725
R23704 frontAnalog_v0p0p1_1.x63.A.n1 frontAnalog_v0p0p1_1.x63.A.t1 17.4109
R23705 frontAnalog_v0p0p1_1.x63.A.n0 frontAnalog_v0p0p1_1.x63.A.n2 9.75129
R23706 frontAnalog_v0p0p1_1.x63.A.n1 frontAnalog_v0p0p1_1.x63.A.t0 9.6027
R23707 frontAnalog_v0p0p1_1.x63.A.n0 frontAnalog_v0p0p1_1.x63.A 2.33338
R23708 frontAnalog_v0p0p1_1.x63.A.n5 frontAnalog_v0p0p1_1.x63.A.t2 8.40929
R23709 frontAnalog_v0p0p1_1.x63.A.n3 frontAnalog_v0p0p1_1.x63.A.t3 8.06629
R23710 frontAnalog_v0p0p1_1.x63.A.n4 frontAnalog_v0p0p1_1.x63.A.n3 1.73501
R23711 frontAnalog_v0p0p1_1.x63.A.n1 frontAnalog_v0p0p1_1.x63.A.n4 0.99025
R23712 frontAnalog_v0p0p1_1.x63.A.n5 frontAnalog_v0p0p1_1.x63.A.n1 0.853186
R23713 frontAnalog_v0p0p1_1.x63.A frontAnalog_v0p0p1_1.x63.A.n0 0.349517
R23714 frontAnalog_v0p0p1_1.x63.A frontAnalog_v0p0p1_1.x63.A.n5 0.24425
R23715 frontAnalog_v0p0p1_5.x65.A.n1 frontAnalog_v0p0p1_5.x65.A.t4 260.322
R23716 frontAnalog_v0p0p1_5.x65.A.n3 frontAnalog_v0p0p1_5.x65.A.t7 233.929
R23717 frontAnalog_v0p0p1_5.x65.A.n1 frontAnalog_v0p0p1_5.x65.A.t6 175.169
R23718 frontAnalog_v0p0p1_5.x65.A.n2 frontAnalog_v0p0p1_5.x65.A.t5 160.416
R23719 frontAnalog_v0p0p1_5.x65.A.n4 frontAnalog_v0p0p1_5.x65.A.t0 17.4109
R23720 frontAnalog_v0p0p1_5.x65.A.n4 frontAnalog_v0p0p1_5.x65.A.t1 10.2053
R23721 frontAnalog_v0p0p1_5.x65.A.n0 frontAnalog_v0p0p1_5.x65.A 2.78715
R23722 frontAnalog_v0p0p1_5.x65.A.n0 frontAnalog_v0p0p1_5.x65.A.n1 9.09103
R23723 frontAnalog_v0p0p1_5.x65.A.n6 frontAnalog_v0p0p1_5.x65.A.t2 7.94569
R23724 frontAnalog_v0p0p1_5.x65.A.n2 frontAnalog_v0p0p1_5.x65.A.t3 7.55846
R23725 frontAnalog_v0p0p1_5.x65.A.n5 frontAnalog_v0p0p1_5.x65.A.n3 1.4614
R23726 frontAnalog_v0p0p1_5.x65.A.n3 frontAnalog_v0p0p1_5.x65.A.n2 1.19626
R23727 frontAnalog_v0p0p1_5.x65.A.n6 frontAnalog_v0p0p1_5.x65.A.n5 0.836961
R23728 frontAnalog_v0p0p1_5.x65.A frontAnalog_v0p0p1_5.x65.A.n0 0.390342
R23729 frontAnalog_v0p0p1_5.x65.A.n5 frontAnalog_v0p0p1_5.x65.A.n4 0.154668
R23730 frontAnalog_v0p0p1_5.x65.A frontAnalog_v0p0p1_5.x65.A.n6 0.08175
R23731 frontAnalog_v0p0p1_14.RSfetsym_0.QN.n1 frontAnalog_v0p0p1_14.RSfetsym_0.QN.t6 117.511
R23732 frontAnalog_v0p0p1_14.RSfetsym_0.QN.n1 frontAnalog_v0p0p1_14.RSfetsym_0.QN.t5 110.698
R23733 frontAnalog_v0p0p1_14.RSfetsym_0.QN.n4 frontAnalog_v0p0p1_14.RSfetsym_0.QN.t0 19.1963
R23734 frontAnalog_v0p0p1_14.RSfetsym_0.QN.n7 frontAnalog_v0p0p1_14.RSfetsym_0.QN.t4 14.2842
R23735 frontAnalog_v0p0p1_14.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_14.RSfetsym_0.QN.t1 14.283
R23736 frontAnalog_v0p0p1_14.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_14.RSfetsym_0.QN.t2 14.283
R23737 frontAnalog_v0p0p1_14.RSfetsym_0.QN.n11 frontAnalog_v0p0p1_14.RSfetsym_0.QN.t3 9.14075
R23738 frontAnalog_v0p0p1_14.RSfetsym_0.QN.n11 frontAnalog_v0p0p1_14.RSfetsym_0.QN.n10 0.74645
R23739 frontAnalog_v0p0p1_14.RSfetsym_0.QN.n2 frontAnalog_v0p0p1_14.RSfetsym_0.QN.n1 0.688382
R23740 frontAnalog_v0p0p1_14.RSfetsym_0.QN.n10 frontAnalog_v0p0p1_14.RSfetsym_0.QN.n9 0.2402
R23741 frontAnalog_v0p0p1_14.RSfetsym_0.QN.n9 frontAnalog_v0p0p1_14.RSfetsym_0.QN.n8 0.236824
R23742 frontAnalog_v0p0p1_14.RSfetsym_0.QN.n4 frontAnalog_v0p0p1_14.RSfetsym_0.QN.n3 0.132187
R23743 frontAnalog_v0p0p1_14.RSfetsym_0.QN.n9 frontAnalog_v0p0p1_14.RSfetsym_0.QN.n4 0.0968646
R23744 frontAnalog_v0p0p1_14.RSfetsym_0.QN frontAnalog_v0p0p1_14.RSfetsym_0.QN.n11 0.0446535
R23745 frontAnalog_v0p0p1_14.RSfetsym_0.QN.n8 frontAnalog_v0p0p1_14.RSfetsym_0.QN.n6 0.0272538
R23746 frontAnalog_v0p0p1_14.RSfetsym_0.QN.n10 frontAnalog_v0p0p1_14.RSfetsym_0.QN.n0 0.00981499
R23747 frontAnalog_v0p0p1_14.RSfetsym_0.QN.n3 frontAnalog_v0p0p1_14.RSfetsym_0.QN.n2 0.00725433
R23748 frontAnalog_v0p0p1_14.RSfetsym_0.QN.n6 frontAnalog_v0p0p1_14.RSfetsym_0.QN.n5 0.00610579
R23749 frontAnalog_v0p0p1_14.RSfetsym_0.QN.n8 frontAnalog_v0p0p1_14.RSfetsym_0.QN.n7 0.00225341
R23750 frontAnalog_v0p0p1_7.RSfetsym_0.QN.n1 frontAnalog_v0p0p1_7.RSfetsym_0.QN.t6 117.511
R23751 frontAnalog_v0p0p1_7.RSfetsym_0.QN.n1 frontAnalog_v0p0p1_7.RSfetsym_0.QN.t5 110.698
R23752 frontAnalog_v0p0p1_7.RSfetsym_0.QN.n4 frontAnalog_v0p0p1_7.RSfetsym_0.QN.t3 19.1963
R23753 frontAnalog_v0p0p1_7.RSfetsym_0.QN.n7 frontAnalog_v0p0p1_7.RSfetsym_0.QN.t4 14.2842
R23754 frontAnalog_v0p0p1_7.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_7.RSfetsym_0.QN.t1 14.283
R23755 frontAnalog_v0p0p1_7.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_7.RSfetsym_0.QN.t2 14.283
R23756 frontAnalog_v0p0p1_7.RSfetsym_0.QN.n11 frontAnalog_v0p0p1_7.RSfetsym_0.QN.t0 9.14075
R23757 frontAnalog_v0p0p1_7.RSfetsym_0.QN.n11 frontAnalog_v0p0p1_7.RSfetsym_0.QN.n10 0.74645
R23758 frontAnalog_v0p0p1_7.RSfetsym_0.QN.n2 frontAnalog_v0p0p1_7.RSfetsym_0.QN.n1 0.688382
R23759 frontAnalog_v0p0p1_7.RSfetsym_0.QN.n10 frontAnalog_v0p0p1_7.RSfetsym_0.QN.n9 0.2402
R23760 frontAnalog_v0p0p1_7.RSfetsym_0.QN.n9 frontAnalog_v0p0p1_7.RSfetsym_0.QN.n8 0.236824
R23761 frontAnalog_v0p0p1_7.RSfetsym_0.QN.n4 frontAnalog_v0p0p1_7.RSfetsym_0.QN.n3 0.132187
R23762 frontAnalog_v0p0p1_7.RSfetsym_0.QN.n9 frontAnalog_v0p0p1_7.RSfetsym_0.QN.n4 0.0968646
R23763 frontAnalog_v0p0p1_7.RSfetsym_0.QN frontAnalog_v0p0p1_7.RSfetsym_0.QN.n11 0.0446535
R23764 frontAnalog_v0p0p1_7.RSfetsym_0.QN.n8 frontAnalog_v0p0p1_7.RSfetsym_0.QN.n6 0.0272538
R23765 frontAnalog_v0p0p1_7.RSfetsym_0.QN.n10 frontAnalog_v0p0p1_7.RSfetsym_0.QN.n0 0.00981499
R23766 frontAnalog_v0p0p1_7.RSfetsym_0.QN.n3 frontAnalog_v0p0p1_7.RSfetsym_0.QN.n2 0.00725433
R23767 frontAnalog_v0p0p1_7.RSfetsym_0.QN.n6 frontAnalog_v0p0p1_7.RSfetsym_0.QN.n5 0.00610579
R23768 frontAnalog_v0p0p1_7.RSfetsym_0.QN.n8 frontAnalog_v0p0p1_7.RSfetsym_0.QN.n7 0.00225341
R23769 frontAnalog_v0p0p1_0.RSfetsym_0.QN.n1 frontAnalog_v0p0p1_0.RSfetsym_0.QN.t5 117.511
R23770 frontAnalog_v0p0p1_0.RSfetsym_0.QN.n1 frontAnalog_v0p0p1_0.RSfetsym_0.QN.t6 110.698
R23771 frontAnalog_v0p0p1_0.RSfetsym_0.QN.n4 frontAnalog_v0p0p1_0.RSfetsym_0.QN.t1 19.1963
R23772 frontAnalog_v0p0p1_0.RSfetsym_0.QN.n7 frontAnalog_v0p0p1_0.RSfetsym_0.QN.t0 14.2842
R23773 frontAnalog_v0p0p1_0.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_0.RSfetsym_0.QN.t3 14.283
R23774 frontAnalog_v0p0p1_0.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_0.RSfetsym_0.QN.t2 14.283
R23775 frontAnalog_v0p0p1_0.RSfetsym_0.QN.n11 frontAnalog_v0p0p1_0.RSfetsym_0.QN.t4 9.14075
R23776 frontAnalog_v0p0p1_0.RSfetsym_0.QN.n11 frontAnalog_v0p0p1_0.RSfetsym_0.QN.n10 0.74645
R23777 frontAnalog_v0p0p1_0.RSfetsym_0.QN.n2 frontAnalog_v0p0p1_0.RSfetsym_0.QN.n1 0.688382
R23778 frontAnalog_v0p0p1_0.RSfetsym_0.QN.n10 frontAnalog_v0p0p1_0.RSfetsym_0.QN.n9 0.2402
R23779 frontAnalog_v0p0p1_0.RSfetsym_0.QN.n9 frontAnalog_v0p0p1_0.RSfetsym_0.QN.n8 0.236824
R23780 frontAnalog_v0p0p1_0.RSfetsym_0.QN.n4 frontAnalog_v0p0p1_0.RSfetsym_0.QN.n3 0.132187
R23781 frontAnalog_v0p0p1_0.RSfetsym_0.QN.n9 frontAnalog_v0p0p1_0.RSfetsym_0.QN.n4 0.0968646
R23782 frontAnalog_v0p0p1_0.RSfetsym_0.QN frontAnalog_v0p0p1_0.RSfetsym_0.QN.n11 0.0446535
R23783 frontAnalog_v0p0p1_0.RSfetsym_0.QN.n8 frontAnalog_v0p0p1_0.RSfetsym_0.QN.n6 0.0272538
R23784 frontAnalog_v0p0p1_0.RSfetsym_0.QN.n10 frontAnalog_v0p0p1_0.RSfetsym_0.QN.n0 0.00981499
R23785 frontAnalog_v0p0p1_0.RSfetsym_0.QN.n3 frontAnalog_v0p0p1_0.RSfetsym_0.QN.n2 0.00725433
R23786 frontAnalog_v0p0p1_0.RSfetsym_0.QN.n6 frontAnalog_v0p0p1_0.RSfetsym_0.QN.n5 0.00610579
R23787 frontAnalog_v0p0p1_0.RSfetsym_0.QN.n8 frontAnalog_v0p0p1_0.RSfetsym_0.QN.n7 0.00225341
R23788 frontAnalog_v0p0p1_1.Q.n8 frontAnalog_v0p0p1_1.Q.t8 196.549
R23789 frontAnalog_v0p0p1_1.Q.n8 frontAnalog_v0p0p1_1.Q.t6 148.35
R23790 frontAnalog_v0p0p1_1.Q.n0 frontAnalog_v0p0p1_1.Q.t7 117.314
R23791 frontAnalog_v0p0p1_1.Q.n0 frontAnalog_v0p0p1_1.Q.t5 110.853
R23792 frontAnalog_v0p0p1_1.Q.n1 frontAnalog_v0p0p1_1.Q.t2 17.6181
R23793 frontAnalog_v0p0p1_1.Q.n3 frontAnalog_v0p0p1_1.Q.t4 14.2865
R23794 frontAnalog_v0p0p1_1.Q.n5 frontAnalog_v0p0p1_1.Q.t0 14.283
R23795 frontAnalog_v0p0p1_1.Q.n5 frontAnalog_v0p0p1_1.Q.t1 14.283
R23796 frontAnalog_v0p0p1_1.Q.n9 frontAnalog_v0p0p1_1.Q.n8 9.49592
R23797 frontAnalog_v0p0p1_1.Q.n7 frontAnalog_v0p0p1_1.Q.t3 8.77744
R23798 frontAnalog_v0p0p1_1.Q.n10 frontAnalog_v0p0p1_1.Q.n9 7.58085
R23799 frontAnalog_v0p0p1_1.Q.n9 frontAnalog_v0p0p1_1.Q 6.44187
R23800 frontAnalog_v0p0p1_1.Q.n11 frontAnalog_v0p0p1_1.Q.n10 2.34543
R23801 frontAnalog_v0p0p1_1.Q.n7 frontAnalog_v0p0p1_1.Q.n6 1.20426
R23802 frontAnalog_v0p0p1_1.Q.n10 frontAnalog_v0p0p1_1.Q 0.88934
R23803 frontAnalog_v0p0p1_1.Q frontAnalog_v0p0p1_1.Q.n11 0.699808
R23804 frontAnalog_v0p0p1_1.Q frontAnalog_v0p0p1_1.Q.n7 0.357737
R23805 frontAnalog_v0p0p1_1.Q.n4 frontAnalog_v0p0p1_1.Q.n3 0.301242
R23806 frontAnalog_v0p0p1_1.Q.n11 frontAnalog_v0p0p1_1.Q 0.200892
R23807 frontAnalog_v0p0p1_1.Q.n2 frontAnalog_v0p0p1_1.Q.n0 0.159555
R23808 frontAnalog_v0p0p1_1.Q.n6 frontAnalog_v0p0p1_1.Q.n5 0.106617
R23809 frontAnalog_v0p0p1_1.Q.n4 frontAnalog_v0p0p1_1.Q.n2 0.0796167
R23810 frontAnalog_v0p0p1_1.Q.n6 frontAnalog_v0p0p1_1.Q.n4 0.0480595
R23811 frontAnalog_v0p0p1_1.Q.n2 frontAnalog_v0p0p1_1.Q.n1 0.000504658
R23812 frontAnalog_v0p0p1_13.x65.A.n1 frontAnalog_v0p0p1_13.x65.A.t4 260.322
R23813 frontAnalog_v0p0p1_13.x65.A.n4 frontAnalog_v0p0p1_13.x65.A.t7 233.929
R23814 frontAnalog_v0p0p1_13.x65.A.n1 frontAnalog_v0p0p1_13.x65.A.t6 175.169
R23815 frontAnalog_v0p0p1_13.x65.A.n3 frontAnalog_v0p0p1_13.x65.A.t5 160.416
R23816 frontAnalog_v0p0p1_13.x65.A.n2 frontAnalog_v0p0p1_13.x65.A.t2 17.4109
R23817 frontAnalog_v0p0p1_13.x65.A.n2 frontAnalog_v0p0p1_13.x65.A.t3 10.2053
R23818 frontAnalog_v0p0p1_13.x65.A.n0 frontAnalog_v0p0p1_13.x65.A 2.78715
R23819 frontAnalog_v0p0p1_13.x65.A.n0 frontAnalog_v0p0p1_13.x65.A.n1 9.09103
R23820 frontAnalog_v0p0p1_13.x65.A.n6 frontAnalog_v0p0p1_13.x65.A.t1 7.94569
R23821 frontAnalog_v0p0p1_13.x65.A.n3 frontAnalog_v0p0p1_13.x65.A.t0 7.55846
R23822 frontAnalog_v0p0p1_13.x65.A.n5 frontAnalog_v0p0p1_13.x65.A.n4 1.4614
R23823 frontAnalog_v0p0p1_13.x65.A.n4 frontAnalog_v0p0p1_13.x65.A.n3 1.19626
R23824 frontAnalog_v0p0p1_13.x65.A.n6 frontAnalog_v0p0p1_13.x65.A.n5 0.836961
R23825 frontAnalog_v0p0p1_13.x65.A frontAnalog_v0p0p1_13.x65.A.n0 0.390342
R23826 frontAnalog_v0p0p1_13.x65.A.n5 frontAnalog_v0p0p1_13.x65.A.n2 0.154668
R23827 frontAnalog_v0p0p1_13.x65.A frontAnalog_v0p0p1_13.x65.A.n6 0.08175
R23828 frontAnalog_v0p0p1_11.RSfetsym_0.QN.n1 frontAnalog_v0p0p1_11.RSfetsym_0.QN.t6 117.511
R23829 frontAnalog_v0p0p1_11.RSfetsym_0.QN.n1 frontAnalog_v0p0p1_11.RSfetsym_0.QN.t5 110.698
R23830 frontAnalog_v0p0p1_11.RSfetsym_0.QN.n4 frontAnalog_v0p0p1_11.RSfetsym_0.QN.t1 19.1963
R23831 frontAnalog_v0p0p1_11.RSfetsym_0.QN.n7 frontAnalog_v0p0p1_11.RSfetsym_0.QN.t4 14.2842
R23832 frontAnalog_v0p0p1_11.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_11.RSfetsym_0.QN.t2 14.283
R23833 frontAnalog_v0p0p1_11.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_11.RSfetsym_0.QN.t3 14.283
R23834 frontAnalog_v0p0p1_11.RSfetsym_0.QN.n11 frontAnalog_v0p0p1_11.RSfetsym_0.QN.t0 9.14075
R23835 frontAnalog_v0p0p1_11.RSfetsym_0.QN.n11 frontAnalog_v0p0p1_11.RSfetsym_0.QN.n10 0.74645
R23836 frontAnalog_v0p0p1_11.RSfetsym_0.QN.n2 frontAnalog_v0p0p1_11.RSfetsym_0.QN.n1 0.688382
R23837 frontAnalog_v0p0p1_11.RSfetsym_0.QN.n10 frontAnalog_v0p0p1_11.RSfetsym_0.QN.n9 0.2402
R23838 frontAnalog_v0p0p1_11.RSfetsym_0.QN.n9 frontAnalog_v0p0p1_11.RSfetsym_0.QN.n8 0.236824
R23839 frontAnalog_v0p0p1_11.RSfetsym_0.QN.n4 frontAnalog_v0p0p1_11.RSfetsym_0.QN.n3 0.132187
R23840 frontAnalog_v0p0p1_11.RSfetsym_0.QN.n9 frontAnalog_v0p0p1_11.RSfetsym_0.QN.n4 0.0968646
R23841 frontAnalog_v0p0p1_11.RSfetsym_0.QN frontAnalog_v0p0p1_11.RSfetsym_0.QN.n11 0.0446535
R23842 frontAnalog_v0p0p1_11.RSfetsym_0.QN.n8 frontAnalog_v0p0p1_11.RSfetsym_0.QN.n6 0.0272538
R23843 frontAnalog_v0p0p1_11.RSfetsym_0.QN.n10 frontAnalog_v0p0p1_11.RSfetsym_0.QN.n0 0.00981499
R23844 frontAnalog_v0p0p1_11.RSfetsym_0.QN.n3 frontAnalog_v0p0p1_11.RSfetsym_0.QN.n2 0.00725433
R23845 frontAnalog_v0p0p1_11.RSfetsym_0.QN.n6 frontAnalog_v0p0p1_11.RSfetsym_0.QN.n5 0.00610579
R23846 frontAnalog_v0p0p1_11.RSfetsym_0.QN.n8 frontAnalog_v0p0p1_11.RSfetsym_0.QN.n7 0.00225341
R23847 frontAnalog_v0p0p1_12.x63.A.n2 frontAnalog_v0p0p1_12.x63.A.t4 260.322
R23848 frontAnalog_v0p0p1_12.x63.A.n4 frontAnalog_v0p0p1_12.x63.A.t5 233.888
R23849 frontAnalog_v0p0p1_12.x63.A.n2 frontAnalog_v0p0p1_12.x63.A.t6 175.169
R23850 frontAnalog_v0p0p1_12.x63.A.n3 frontAnalog_v0p0p1_12.x63.A.t7 159.725
R23851 frontAnalog_v0p0p1_12.x63.A.n1 frontAnalog_v0p0p1_12.x63.A.t2 17.4109
R23852 frontAnalog_v0p0p1_12.x63.A.n0 frontAnalog_v0p0p1_12.x63.A.n2 9.75129
R23853 frontAnalog_v0p0p1_12.x63.A.n1 frontAnalog_v0p0p1_12.x63.A.t3 9.6037
R23854 frontAnalog_v0p0p1_12.x63.A.n0 frontAnalog_v0p0p1_12.x63.A 2.33338
R23855 frontAnalog_v0p0p1_12.x63.A.n5 frontAnalog_v0p0p1_12.x63.A.t1 8.40929
R23856 frontAnalog_v0p0p1_12.x63.A.n3 frontAnalog_v0p0p1_12.x63.A.t0 8.06629
R23857 frontAnalog_v0p0p1_12.x63.A.n4 frontAnalog_v0p0p1_12.x63.A.n3 1.73501
R23858 frontAnalog_v0p0p1_12.x63.A.n1 frontAnalog_v0p0p1_12.x63.A.n4 0.99025
R23859 frontAnalog_v0p0p1_12.x63.A.n5 frontAnalog_v0p0p1_12.x63.A.n1 0.853186
R23860 frontAnalog_v0p0p1_12.x63.A frontAnalog_v0p0p1_12.x63.A.n0 0.349517
R23861 frontAnalog_v0p0p1_12.x63.A frontAnalog_v0p0p1_12.x63.A.n5 0.24425
R23862 frontAnalog_v0p0p1_4.RSfetsym_0.QN.n1 frontAnalog_v0p0p1_4.RSfetsym_0.QN.t6 117.511
R23863 frontAnalog_v0p0p1_4.RSfetsym_0.QN.n1 frontAnalog_v0p0p1_4.RSfetsym_0.QN.t5 110.698
R23864 frontAnalog_v0p0p1_4.RSfetsym_0.QN.n4 frontAnalog_v0p0p1_4.RSfetsym_0.QN.t0 19.1963
R23865 frontAnalog_v0p0p1_4.RSfetsym_0.QN.n7 frontAnalog_v0p0p1_4.RSfetsym_0.QN.t4 14.2842
R23866 frontAnalog_v0p0p1_4.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_4.RSfetsym_0.QN.t1 14.283
R23867 frontAnalog_v0p0p1_4.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_4.RSfetsym_0.QN.t2 14.283
R23868 frontAnalog_v0p0p1_4.RSfetsym_0.QN.n11 frontAnalog_v0p0p1_4.RSfetsym_0.QN.t3 9.14075
R23869 frontAnalog_v0p0p1_4.RSfetsym_0.QN.n11 frontAnalog_v0p0p1_4.RSfetsym_0.QN.n10 0.74645
R23870 frontAnalog_v0p0p1_4.RSfetsym_0.QN.n2 frontAnalog_v0p0p1_4.RSfetsym_0.QN.n1 0.688382
R23871 frontAnalog_v0p0p1_4.RSfetsym_0.QN.n10 frontAnalog_v0p0p1_4.RSfetsym_0.QN.n9 0.2402
R23872 frontAnalog_v0p0p1_4.RSfetsym_0.QN.n9 frontAnalog_v0p0p1_4.RSfetsym_0.QN.n8 0.236824
R23873 frontAnalog_v0p0p1_4.RSfetsym_0.QN.n4 frontAnalog_v0p0p1_4.RSfetsym_0.QN.n3 0.132187
R23874 frontAnalog_v0p0p1_4.RSfetsym_0.QN.n9 frontAnalog_v0p0p1_4.RSfetsym_0.QN.n4 0.0968646
R23875 frontAnalog_v0p0p1_4.RSfetsym_0.QN frontAnalog_v0p0p1_4.RSfetsym_0.QN.n11 0.0446535
R23876 frontAnalog_v0p0p1_4.RSfetsym_0.QN.n8 frontAnalog_v0p0p1_4.RSfetsym_0.QN.n6 0.0272538
R23877 frontAnalog_v0p0p1_4.RSfetsym_0.QN.n10 frontAnalog_v0p0p1_4.RSfetsym_0.QN.n0 0.00981499
R23878 frontAnalog_v0p0p1_4.RSfetsym_0.QN.n3 frontAnalog_v0p0p1_4.RSfetsym_0.QN.n2 0.00725433
R23879 frontAnalog_v0p0p1_4.RSfetsym_0.QN.n6 frontAnalog_v0p0p1_4.RSfetsym_0.QN.n5 0.00610579
R23880 frontAnalog_v0p0p1_4.RSfetsym_0.QN.n8 frontAnalog_v0p0p1_4.RSfetsym_0.QN.n7 0.00225341
R23881 frontAnalog_v0p0p1_8.Q.n3 frontAnalog_v0p0p1_8.Q.t5 261.116
R23882 frontAnalog_v0p0p1_8.Q.n0 frontAnalog_v0p0p1_8.Q.t7 186.03
R23883 frontAnalog_v0p0p1_8.Q.n3 frontAnalog_v0p0p1_8.Q.t10 155.746
R23884 frontAnalog_v0p0p1_8.Q.n0 frontAnalog_v0p0p1_8.Q.t8 137.829
R23885 frontAnalog_v0p0p1_8.Q.n12 frontAnalog_v0p0p1_8.Q.t6 117.314
R23886 frontAnalog_v0p0p1_8.Q.n12 frontAnalog_v0p0p1_8.Q.t9 110.852
R23887 frontAnalog_v0p0p1_8.Q frontAnalog_v0p0p1_8.Q.n0 78.5605
R23888 frontAnalog_v0p0p1_8.Q.n9 frontAnalog_v0p0p1_8.Q 47.2619
R23889 frontAnalog_v0p0p1_8.Q.n13 frontAnalog_v0p0p1_8.Q.t3 17.6181
R23890 frontAnalog_v0p0p1_8.Q.n15 frontAnalog_v0p0p1_8.Q.t0 14.2865
R23891 frontAnalog_v0p0p1_8.Q.n17 frontAnalog_v0p0p1_8.Q.t2 14.283
R23892 frontAnalog_v0p0p1_8.Q.n17 frontAnalog_v0p0p1_8.Q.t1 14.283
R23893 frontAnalog_v0p0p1_8.Q.n19 frontAnalog_v0p0p1_8.Q.t4 8.77592
R23894 frontAnalog_v0p0p1_8.Q.n4 frontAnalog_v0p0p1_8.Q.n3 7.65549
R23895 frontAnalog_v0p0p1_8.Q.n9 frontAnalog_v0p0p1_8.Q.n8 4.04922
R23896 frontAnalog_v0p0p1_8.Q.n5 frontAnalog_v0p0p1_8.Q 2.46419
R23897 frontAnalog_v0p0p1_8.Q.n20 frontAnalog_v0p0p1_8.Q.n11 1.98646
R23898 frontAnalog_v0p0p1_8.Q.n19 frontAnalog_v0p0p1_8.Q.n18 1.20426
R23899 frontAnalog_v0p0p1_8.Q.n10 frontAnalog_v0p0p1_8.Q 0.808983
R23900 frontAnalog_v0p0p1_8.Q.n5 frontAnalog_v0p0p1_8.Q.n4 0.754023
R23901 frontAnalog_v0p0p1_8.Q.n11 frontAnalog_v0p0p1_8.Q.n10 0.674526
R23902 frontAnalog_v0p0p1_8.Q.n10 frontAnalog_v0p0p1_8.Q.n9 0.478179
R23903 frontAnalog_v0p0p1_8.Q.n20 frontAnalog_v0p0p1_8.Q.n19 0.325111
R23904 frontAnalog_v0p0p1_8.Q.n16 frontAnalog_v0p0p1_8.Q.n15 0.300242
R23905 frontAnalog_v0p0p1_8.Q.n11 frontAnalog_v0p0p1_8.Q 0.20675
R23906 frontAnalog_v0p0p1_8.Q.n14 frontAnalog_v0p0p1_8.Q.n12 0.159555
R23907 frontAnalog_v0p0p1_8.Q.n18 frontAnalog_v0p0p1_8.Q.n17 0.106617
R23908 frontAnalog_v0p0p1_8.Q.n16 frontAnalog_v0p0p1_8.Q.n14 0.0796167
R23909 frontAnalog_v0p0p1_8.Q.n18 frontAnalog_v0p0p1_8.Q.n16 0.0480595
R23910 frontAnalog_v0p0p1_8.Q frontAnalog_v0p0p1_8.Q.n20 0.0469368
R23911 frontAnalog_v0p0p1_8.Q.n7 frontAnalog_v0p0p1_8.Q.n6 0.0326429
R23912 frontAnalog_v0p0p1_8.Q.n7 frontAnalog_v0p0p1_8.Q.n2 0.0197253
R23913 frontAnalog_v0p0p1_8.Q.n8 frontAnalog_v0p0p1_8.Q.n1 0.00182856
R23914 frontAnalog_v0p0p1_8.Q.n8 frontAnalog_v0p0p1_8.Q.n7 0.00149885
R23915 frontAnalog_v0p0p1_8.Q.n7 frontAnalog_v0p0p1_8.Q.n5 0.00125261
R23916 frontAnalog_v0p0p1_8.Q.n14 frontAnalog_v0p0p1_8.Q.n13 0.000504658
R23917 frontAnalog_v0p0p1_11.x63.A.n2 frontAnalog_v0p0p1_11.x63.A.t5 260.322
R23918 frontAnalog_v0p0p1_11.x63.A.n4 frontAnalog_v0p0p1_11.x63.A.t6 233.888
R23919 frontAnalog_v0p0p1_11.x63.A.n2 frontAnalog_v0p0p1_11.x63.A.t7 175.169
R23920 frontAnalog_v0p0p1_11.x63.A.n3 frontAnalog_v0p0p1_11.x63.A.t4 159.725
R23921 frontAnalog_v0p0p1_11.x63.A.n1 frontAnalog_v0p0p1_11.x63.A.t2 17.4109
R23922 frontAnalog_v0p0p1_11.x63.A.n0 frontAnalog_v0p0p1_11.x63.A.n2 9.75129
R23923 frontAnalog_v0p0p1_11.x63.A.n1 frontAnalog_v0p0p1_11.x63.A.t3 9.6037
R23924 frontAnalog_v0p0p1_11.x63.A.n0 frontAnalog_v0p0p1_11.x63.A 2.33338
R23925 frontAnalog_v0p0p1_11.x63.A.n5 frontAnalog_v0p0p1_11.x63.A.t1 8.40929
R23926 frontAnalog_v0p0p1_11.x63.A.n3 frontAnalog_v0p0p1_11.x63.A.t0 8.06629
R23927 frontAnalog_v0p0p1_11.x63.A.n4 frontAnalog_v0p0p1_11.x63.A.n3 1.73501
R23928 frontAnalog_v0p0p1_11.x63.A.n1 frontAnalog_v0p0p1_11.x63.A.n4 0.99025
R23929 frontAnalog_v0p0p1_11.x63.A.n5 frontAnalog_v0p0p1_11.x63.A.n1 0.853186
R23930 frontAnalog_v0p0p1_11.x63.A frontAnalog_v0p0p1_11.x63.A.n0 0.349517
R23931 frontAnalog_v0p0p1_11.x63.A frontAnalog_v0p0p1_11.x63.A.n5 0.24425
R23932 frontAnalog_v0p0p1_8.x65.A.n1 frontAnalog_v0p0p1_8.x65.A.t4 260.322
R23933 frontAnalog_v0p0p1_8.x65.A.n3 frontAnalog_v0p0p1_8.x65.A.t7 233.929
R23934 frontAnalog_v0p0p1_8.x65.A.n1 frontAnalog_v0p0p1_8.x65.A.t6 175.169
R23935 frontAnalog_v0p0p1_8.x65.A.n2 frontAnalog_v0p0p1_8.x65.A.t5 160.416
R23936 frontAnalog_v0p0p1_8.x65.A.n4 frontAnalog_v0p0p1_8.x65.A.t0 17.4109
R23937 frontAnalog_v0p0p1_8.x65.A.n4 frontAnalog_v0p0p1_8.x65.A.t1 10.2053
R23938 frontAnalog_v0p0p1_8.x65.A.n0 frontAnalog_v0p0p1_8.x65.A 2.78715
R23939 frontAnalog_v0p0p1_8.x65.A.n0 frontAnalog_v0p0p1_8.x65.A.n1 9.09103
R23940 frontAnalog_v0p0p1_8.x65.A.n6 frontAnalog_v0p0p1_8.x65.A.t2 7.94569
R23941 frontAnalog_v0p0p1_8.x65.A.n2 frontAnalog_v0p0p1_8.x65.A.t3 7.55846
R23942 frontAnalog_v0p0p1_8.x65.A.n5 frontAnalog_v0p0p1_8.x65.A.n3 1.4614
R23943 frontAnalog_v0p0p1_8.x65.A.n3 frontAnalog_v0p0p1_8.x65.A.n2 1.19626
R23944 frontAnalog_v0p0p1_8.x65.A.n6 frontAnalog_v0p0p1_8.x65.A.n5 0.836961
R23945 frontAnalog_v0p0p1_8.x65.A frontAnalog_v0p0p1_8.x65.A.n0 0.390342
R23946 frontAnalog_v0p0p1_8.x65.A.n5 frontAnalog_v0p0p1_8.x65.A.n4 0.154668
R23947 frontAnalog_v0p0p1_8.x65.A frontAnalog_v0p0p1_8.x65.A.n6 0.08175
R23948 16to4_PriorityEncoder_v0p0p1_0.I14.n25 16to4_PriorityEncoder_v0p0p1_0.I14.t11 260.435
R23949 16to4_PriorityEncoder_v0p0p1_0.I14.n10 16to4_PriorityEncoder_v0p0p1_0.I14.t12 229.433
R23950 16to4_PriorityEncoder_v0p0p1_0.I14.n20 16to4_PriorityEncoder_v0p0p1_0.I14.t9 196.549
R23951 16to4_PriorityEncoder_v0p0p1_0.I14.n10 16to4_PriorityEncoder_v0p0p1_0.I14.t6 158.886
R23952 16to4_PriorityEncoder_v0p0p1_0.I14.n25 16to4_PriorityEncoder_v0p0p1_0.I14.t5 156.403
R23953 16to4_PriorityEncoder_v0p0p1_0.I14.n20 16to4_PriorityEncoder_v0p0p1_0.I14.t7 148.35
R23954 16to4_PriorityEncoder_v0p0p1_0.I14.n0 16to4_PriorityEncoder_v0p0p1_0.I14.t10 117.314
R23955 16to4_PriorityEncoder_v0p0p1_0.I14.n0 16to4_PriorityEncoder_v0p0p1_0.I14.t8 110.852
R23956 16to4_PriorityEncoder_v0p0p1_0.I14.n21 16to4_PriorityEncoder_v0p0p1_0.I14.n20 76.0005
R23957 16to4_PriorityEncoder_v0p0p1_0.I14.n1 16to4_PriorityEncoder_v0p0p1_0.I14.t4 17.6181
R23958 16to4_PriorityEncoder_v0p0p1_0.I14.n3 16to4_PriorityEncoder_v0p0p1_0.I14.t0 14.2865
R23959 16to4_PriorityEncoder_v0p0p1_0.I14.n5 16to4_PriorityEncoder_v0p0p1_0.I14.t2 14.283
R23960 16to4_PriorityEncoder_v0p0p1_0.I14.n5 16to4_PriorityEncoder_v0p0p1_0.I14.t3 14.283
R23961 16to4_PriorityEncoder_v0p0p1_0.I14 16to4_PriorityEncoder_v0p0p1_0.I14.n24 9.3005
R23962 16to4_PriorityEncoder_v0p0p1_0.I14.n7 16to4_PriorityEncoder_v0p0p1_0.I14.t1 8.77592
R23963 16to4_PriorityEncoder_v0p0p1_0.I14.n26 16to4_PriorityEncoder_v0p0p1_0.I14.n25 7.60183
R23964 16to4_PriorityEncoder_v0p0p1_0.I14.n11 16to4_PriorityEncoder_v0p0p1_0.I14.n10 7.39078
R23965 16to4_PriorityEncoder_v0p0p1_0.I14 16to4_PriorityEncoder_v0p0p1_0.I14.n32 7.21371
R23966 16to4_PriorityEncoder_v0p0p1_0.I14.n30 16to4_PriorityEncoder_v0p0p1_0.I14.n22 6.24391
R23967 16to4_PriorityEncoder_v0p0p1_0.I14.n21 16to4_PriorityEncoder_v0p0p1_0.I14 5.78114
R23968 16to4_PriorityEncoder_v0p0p1_0.I14.n26 16to4_PriorityEncoder_v0p0p1_0.I14 4.8645
R23969 16to4_PriorityEncoder_v0p0p1_0.I14.n14 16to4_PriorityEncoder_v0p0p1_0.I14.n13 4.5005
R23970 16to4_PriorityEncoder_v0p0p1_0.I14.n30 16to4_PriorityEncoder_v0p0p1_0.I14.n29 3.53643
R23971 16to4_PriorityEncoder_v0p0p1_0.I14.n22 16to4_PriorityEncoder_v0p0p1_0.I14.n21 3.51018
R23972 16to4_PriorityEncoder_v0p0p1_0.I14.n13 16to4_PriorityEncoder_v0p0p1_0.I14.n12 3.46717
R23973 16to4_PriorityEncoder_v0p0p1_0.I14.n7 16to4_PriorityEncoder_v0p0p1_0.I14.n6 1.20426
R23974 16to4_PriorityEncoder_v0p0p1_0.I14.n19 16to4_PriorityEncoder_v0p0p1_0.I14.n18 1.11384
R23975 16to4_PriorityEncoder_v0p0p1_0.I14.n13 16to4_PriorityEncoder_v0p0p1_0.I14.n11 1.06717
R23976 16to4_PriorityEncoder_v0p0p1_0.I14.n12 16to4_PriorityEncoder_v0p0p1_0.I14 1.06717
R23977 16to4_PriorityEncoder_v0p0p1_0.I14.n31 16to4_PriorityEncoder_v0p0p1_0.I14.n19 0.767464
R23978 16to4_PriorityEncoder_v0p0p1_0.I14.n32 16to4_PriorityEncoder_v0p0p1_0.I14.n31 0.531993
R23979 16to4_PriorityEncoder_v0p0p1_0.I14.n19 16to4_PriorityEncoder_v0p0p1_0.I14 0.372375
R23980 16to4_PriorityEncoder_v0p0p1_0.I14 16to4_PriorityEncoder_v0p0p1_0.I14.n7 0.370547
R23981 16to4_PriorityEncoder_v0p0p1_0.I14.n31 16to4_PriorityEncoder_v0p0p1_0.I14.n30 0.321929
R23982 16to4_PriorityEncoder_v0p0p1_0.I14.n4 16to4_PriorityEncoder_v0p0p1_0.I14.n3 0.300242
R23983 16to4_PriorityEncoder_v0p0p1_0.I14.n22 16to4_PriorityEncoder_v0p0p1_0.I14 0.206952
R23984 16to4_PriorityEncoder_v0p0p1_0.I14.n32 16to4_PriorityEncoder_v0p0p1_0.I14 0.2005
R23985 16to4_PriorityEncoder_v0p0p1_0.I14.n2 16to4_PriorityEncoder_v0p0p1_0.I14.n0 0.159555
R23986 16to4_PriorityEncoder_v0p0p1_0.I14.n6 16to4_PriorityEncoder_v0p0p1_0.I14.n5 0.106617
R23987 16to4_PriorityEncoder_v0p0p1_0.I14.n4 16to4_PriorityEncoder_v0p0p1_0.I14.n2 0.0796167
R23988 16to4_PriorityEncoder_v0p0p1_0.I14.n6 16to4_PriorityEncoder_v0p0p1_0.I14.n4 0.0480595
R23989 16to4_PriorityEncoder_v0p0p1_0.I14.n28 16to4_PriorityEncoder_v0p0p1_0.I14.n24 0.0344286
R23990 16to4_PriorityEncoder_v0p0p1_0.I14.n18 16to4_PriorityEncoder_v0p0p1_0.I14.n17 0.028
R23991 16to4_PriorityEncoder_v0p0p1_0.I14.n16 16to4_PriorityEncoder_v0p0p1_0.I14.n15 0.0142363
R23992 16to4_PriorityEncoder_v0p0p1_0.I14.n16 16to4_PriorityEncoder_v0p0p1_0.I14.n14 0.00599451
R23993 16to4_PriorityEncoder_v0p0p1_0.I14.n9 16to4_PriorityEncoder_v0p0p1_0.I14.n8 0.00409723
R23994 16to4_PriorityEncoder_v0p0p1_0.I14.n14 16to4_PriorityEncoder_v0p0p1_0.I14.n9 0.00202085
R23995 16to4_PriorityEncoder_v0p0p1_0.I14.n29 16to4_PriorityEncoder_v0p0p1_0.I14.n23 0.00182856
R23996 16to4_PriorityEncoder_v0p0p1_0.I14.n29 16to4_PriorityEncoder_v0p0p1_0.I14.n28 0.00149885
R23997 16to4_PriorityEncoder_v0p0p1_0.I14.n27 16to4_PriorityEncoder_v0p0p1_0.I14.n26 0.00133362
R23998 16to4_PriorityEncoder_v0p0p1_0.I14.n28 16to4_PriorityEncoder_v0p0p1_0.I14.n27 0.00100077
R23999 16to4_PriorityEncoder_v0p0p1_0.I14.n17 16to4_PriorityEncoder_v0p0p1_0.I14.n16 0.000617139
R24000 16to4_PriorityEncoder_v0p0p1_0.I14.n2 16to4_PriorityEncoder_v0p0p1_0.I14.n1 0.000504658
R24001 16to4_PriorityEncoder_v0p0p1_0.I15.n11 16to4_PriorityEncoder_v0p0p1_0.I15.t5 261.116
R24002 16to4_PriorityEncoder_v0p0p1_0.I15.n8 16to4_PriorityEncoder_v0p0p1_0.I15.t7 186.03
R24003 16to4_PriorityEncoder_v0p0p1_0.I15.n11 16to4_PriorityEncoder_v0p0p1_0.I15.t9 155.746
R24004 16to4_PriorityEncoder_v0p0p1_0.I15.n8 16to4_PriorityEncoder_v0p0p1_0.I15.t6 137.829
R24005 16to4_PriorityEncoder_v0p0p1_0.I15.n0 16to4_PriorityEncoder_v0p0p1_0.I15.t10 117.314
R24006 16to4_PriorityEncoder_v0p0p1_0.I15.n0 16to4_PriorityEncoder_v0p0p1_0.I15.t8 110.852
R24007 16to4_PriorityEncoder_v0p0p1_0.I15 16to4_PriorityEncoder_v0p0p1_0.I15.n8 78.5605
R24008 16to4_PriorityEncoder_v0p0p1_0.I15.n17 16to4_PriorityEncoder_v0p0p1_0.I15 47.2619
R24009 16to4_PriorityEncoder_v0p0p1_0.I15.n1 16to4_PriorityEncoder_v0p0p1_0.I15.t1 17.6181
R24010 16to4_PriorityEncoder_v0p0p1_0.I15.n3 16to4_PriorityEncoder_v0p0p1_0.I15.t0 14.2865
R24011 16to4_PriorityEncoder_v0p0p1_0.I15.n5 16to4_PriorityEncoder_v0p0p1_0.I15.t3 14.283
R24012 16to4_PriorityEncoder_v0p0p1_0.I15.n5 16to4_PriorityEncoder_v0p0p1_0.I15.t2 14.283
R24013 16to4_PriorityEncoder_v0p0p1_0.I15.n7 16to4_PriorityEncoder_v0p0p1_0.I15.t4 8.77592
R24014 16to4_PriorityEncoder_v0p0p1_0.I15 16to4_PriorityEncoder_v0p0p1_0.I15.n19 8.02299
R24015 16to4_PriorityEncoder_v0p0p1_0.I15.n12 16to4_PriorityEncoder_v0p0p1_0.I15.n11 7.65549
R24016 16to4_PriorityEncoder_v0p0p1_0.I15.n17 16to4_PriorityEncoder_v0p0p1_0.I15.n16 4.04922
R24017 16to4_PriorityEncoder_v0p0p1_0.I15.n13 16to4_PriorityEncoder_v0p0p1_0.I15 2.46419
R24018 16to4_PriorityEncoder_v0p0p1_0.I15.n7 16to4_PriorityEncoder_v0p0p1_0.I15.n6 1.20426
R24019 16to4_PriorityEncoder_v0p0p1_0.I15.n13 16to4_PriorityEncoder_v0p0p1_0.I15.n12 0.754023
R24020 16to4_PriorityEncoder_v0p0p1_0.I15.n18 16to4_PriorityEncoder_v0p0p1_0.I15 0.70184
R24021 16to4_PriorityEncoder_v0p0p1_0.I15.n19 16to4_PriorityEncoder_v0p0p1_0.I15.n18 0.691178
R24022 16to4_PriorityEncoder_v0p0p1_0.I15.n18 16to4_PriorityEncoder_v0p0p1_0.I15.n17 0.585321
R24023 16to4_PriorityEncoder_v0p0p1_0.I15 16to4_PriorityEncoder_v0p0p1_0.I15.n7 0.370547
R24024 16to4_PriorityEncoder_v0p0p1_0.I15.n4 16to4_PriorityEncoder_v0p0p1_0.I15.n3 0.300242
R24025 16to4_PriorityEncoder_v0p0p1_0.I15.n19 16to4_PriorityEncoder_v0p0p1_0.I15 0.2005
R24026 16to4_PriorityEncoder_v0p0p1_0.I15.n2 16to4_PriorityEncoder_v0p0p1_0.I15.n0 0.159555
R24027 16to4_PriorityEncoder_v0p0p1_0.I15.n6 16to4_PriorityEncoder_v0p0p1_0.I15.n5 0.106617
R24028 16to4_PriorityEncoder_v0p0p1_0.I15.n4 16to4_PriorityEncoder_v0p0p1_0.I15.n2 0.0796167
R24029 16to4_PriorityEncoder_v0p0p1_0.I15.n6 16to4_PriorityEncoder_v0p0p1_0.I15.n4 0.0480595
R24030 16to4_PriorityEncoder_v0p0p1_0.I15.n15 16to4_PriorityEncoder_v0p0p1_0.I15.n14 0.0326429
R24031 16to4_PriorityEncoder_v0p0p1_0.I15.n15 16to4_PriorityEncoder_v0p0p1_0.I15.n10 0.0197253
R24032 16to4_PriorityEncoder_v0p0p1_0.I15.n16 16to4_PriorityEncoder_v0p0p1_0.I15.n9 0.00182856
R24033 16to4_PriorityEncoder_v0p0p1_0.I15.n16 16to4_PriorityEncoder_v0p0p1_0.I15.n15 0.00149885
R24034 16to4_PriorityEncoder_v0p0p1_0.I15.n15 16to4_PriorityEncoder_v0p0p1_0.I15.n13 0.00125261
R24035 16to4_PriorityEncoder_v0p0p1_0.I15.n2 16to4_PriorityEncoder_v0p0p1_0.I15.n1 0.000504658
R24036 frontAnalog_v0p0p1_13.Q.n4 frontAnalog_v0p0p1_13.Q.t7 334.723
R24037 frontAnalog_v0p0p1_13.Q.n3 frontAnalog_v0p0p1_13.Q.t10 323.342
R24038 frontAnalog_v0p0p1_13.Q.n4 frontAnalog_v0p0p1_13.Q.t9 206.19
R24039 frontAnalog_v0p0p1_13.Q.n3 frontAnalog_v0p0p1_13.Q.t6 194.809
R24040 frontAnalog_v0p0p1_13.Q.n0 frontAnalog_v0p0p1_13.Q.t5 186.03
R24041 frontAnalog_v0p0p1_13.Q.n0 frontAnalog_v0p0p1_13.Q.t11 137.829
R24042 frontAnalog_v0p0p1_13.Q.n8 frontAnalog_v0p0p1_13.Q.t12 117.314
R24043 frontAnalog_v0p0p1_13.Q.n8 frontAnalog_v0p0p1_13.Q.t8 110.853
R24044 frontAnalog_v0p0p1_13.Q frontAnalog_v0p0p1_13.Q.n4 84.2291
R24045 frontAnalog_v0p0p1_13.Q frontAnalog_v0p0p1_13.Q.n3 82.1338
R24046 frontAnalog_v0p0p1_13.Q.n1 frontAnalog_v0p0p1_13.Q.n0 76.0005
R24047 frontAnalog_v0p0p1_13.Q.n2 frontAnalog_v0p0p1_13.Q 66.7187
R24048 frontAnalog_v0p0p1_13.Q.n5 frontAnalog_v0p0p1_13.Q 26.4877
R24049 frontAnalog_v0p0p1_13.Q.n9 frontAnalog_v0p0p1_13.Q.t1 17.6181
R24050 frontAnalog_v0p0p1_13.Q.n11 frontAnalog_v0p0p1_13.Q.t0 14.2865
R24051 frontAnalog_v0p0p1_13.Q.n13 frontAnalog_v0p0p1_13.Q.t2 14.283
R24052 frontAnalog_v0p0p1_13.Q.n13 frontAnalog_v0p0p1_13.Q.t3 14.283
R24053 frontAnalog_v0p0p1_13.Q.n15 frontAnalog_v0p0p1_13.Q.t4 8.77744
R24054 frontAnalog_v0p0p1_13.Q.n1 frontAnalog_v0p0p1_13.Q 7.31479
R24055 frontAnalog_v0p0p1_13.Q.n16 frontAnalog_v0p0p1_13.Q.n7 6.66218
R24056 frontAnalog_v0p0p1_13.Q.n5 frontAnalog_v0p0p1_13.Q 4.36044
R24057 frontAnalog_v0p0p1_13.Q frontAnalog_v0p0p1_13.Q.n1 4.02336
R24058 frontAnalog_v0p0p1_13.Q.n6 frontAnalog_v0p0p1_13.Q.n5 2.61211
R24059 frontAnalog_v0p0p1_13.Q.n6 frontAnalog_v0p0p1_13.Q.n2 1.25943
R24060 frontAnalog_v0p0p1_13.Q.n15 frontAnalog_v0p0p1_13.Q.n14 1.20426
R24061 frontAnalog_v0p0p1_13.Q.n2 frontAnalog_v0p0p1_13.Q 0.969697
R24062 frontAnalog_v0p0p1_13.Q.n16 frontAnalog_v0p0p1_13.Q.n15 0.325111
R24063 frontAnalog_v0p0p1_13.Q.n12 frontAnalog_v0p0p1_13.Q.n11 0.301242
R24064 frontAnalog_v0p0p1_13.Q.n7 frontAnalog_v0p0p1_13.Q.n6 0.300322
R24065 frontAnalog_v0p0p1_13.Q.n7 frontAnalog_v0p0p1_13.Q 0.20675
R24066 frontAnalog_v0p0p1_13.Q.n10 frontAnalog_v0p0p1_13.Q.n8 0.159555
R24067 frontAnalog_v0p0p1_13.Q.n14 frontAnalog_v0p0p1_13.Q.n13 0.106617
R24068 frontAnalog_v0p0p1_13.Q.n12 frontAnalog_v0p0p1_13.Q.n10 0.0796167
R24069 frontAnalog_v0p0p1_13.Q.n14 frontAnalog_v0p0p1_13.Q.n12 0.0480595
R24070 frontAnalog_v0p0p1_13.Q frontAnalog_v0p0p1_13.Q.n16 0.0469368
R24071 frontAnalog_v0p0p1_13.Q.n10 frontAnalog_v0p0p1_13.Q.n9 0.000504658
R24072 frontAnalog_v0p0p1_1.RSfetsym_0.QN.n1 frontAnalog_v0p0p1_1.RSfetsym_0.QN.t6 117.511
R24073 frontAnalog_v0p0p1_1.RSfetsym_0.QN.n1 frontAnalog_v0p0p1_1.RSfetsym_0.QN.t5 110.698
R24074 frontAnalog_v0p0p1_1.RSfetsym_0.QN.n4 frontAnalog_v0p0p1_1.RSfetsym_0.QN.t1 19.1963
R24075 frontAnalog_v0p0p1_1.RSfetsym_0.QN.n7 frontAnalog_v0p0p1_1.RSfetsym_0.QN.t4 14.2842
R24076 frontAnalog_v0p0p1_1.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_1.RSfetsym_0.QN.t3 14.283
R24077 frontAnalog_v0p0p1_1.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_1.RSfetsym_0.QN.t2 14.283
R24078 frontAnalog_v0p0p1_1.RSfetsym_0.QN.n11 frontAnalog_v0p0p1_1.RSfetsym_0.QN.t0 9.14075
R24079 frontAnalog_v0p0p1_1.RSfetsym_0.QN.n11 frontAnalog_v0p0p1_1.RSfetsym_0.QN.n10 0.74645
R24080 frontAnalog_v0p0p1_1.RSfetsym_0.QN.n2 frontAnalog_v0p0p1_1.RSfetsym_0.QN.n1 0.688382
R24081 frontAnalog_v0p0p1_1.RSfetsym_0.QN.n10 frontAnalog_v0p0p1_1.RSfetsym_0.QN.n9 0.2402
R24082 frontAnalog_v0p0p1_1.RSfetsym_0.QN.n9 frontAnalog_v0p0p1_1.RSfetsym_0.QN.n8 0.236824
R24083 frontAnalog_v0p0p1_1.RSfetsym_0.QN.n4 frontAnalog_v0p0p1_1.RSfetsym_0.QN.n3 0.132187
R24084 frontAnalog_v0p0p1_1.RSfetsym_0.QN.n9 frontAnalog_v0p0p1_1.RSfetsym_0.QN.n4 0.0968646
R24085 frontAnalog_v0p0p1_1.RSfetsym_0.QN frontAnalog_v0p0p1_1.RSfetsym_0.QN.n11 0.0446535
R24086 frontAnalog_v0p0p1_1.RSfetsym_0.QN.n8 frontAnalog_v0p0p1_1.RSfetsym_0.QN.n6 0.0272538
R24087 frontAnalog_v0p0p1_1.RSfetsym_0.QN.n10 frontAnalog_v0p0p1_1.RSfetsym_0.QN.n0 0.00981499
R24088 frontAnalog_v0p0p1_1.RSfetsym_0.QN.n3 frontAnalog_v0p0p1_1.RSfetsym_0.QN.n2 0.00725433
R24089 frontAnalog_v0p0p1_1.RSfetsym_0.QN.n6 frontAnalog_v0p0p1_1.RSfetsym_0.QN.n5 0.00610579
R24090 frontAnalog_v0p0p1_1.RSfetsym_0.QN.n8 frontAnalog_v0p0p1_1.RSfetsym_0.QN.n7 0.00225341
R24091 16to4_PriorityEncoder_v0p0p1_0.I11.n12 16to4_PriorityEncoder_v0p0p1_0.I11.t7 334.723
R24092 16to4_PriorityEncoder_v0p0p1_0.I11.n11 16to4_PriorityEncoder_v0p0p1_0.I11.t9 323.342
R24093 16to4_PriorityEncoder_v0p0p1_0.I11.n12 16to4_PriorityEncoder_v0p0p1_0.I11.t11 206.19
R24094 16to4_PriorityEncoder_v0p0p1_0.I11.n11 16to4_PriorityEncoder_v0p0p1_0.I11.t6 194.809
R24095 16to4_PriorityEncoder_v0p0p1_0.I11.n8 16to4_PriorityEncoder_v0p0p1_0.I11.t5 186.03
R24096 16to4_PriorityEncoder_v0p0p1_0.I11.n8 16to4_PriorityEncoder_v0p0p1_0.I11.t10 137.829
R24097 16to4_PriorityEncoder_v0p0p1_0.I11.n0 16to4_PriorityEncoder_v0p0p1_0.I11.t12 117.314
R24098 16to4_PriorityEncoder_v0p0p1_0.I11.n0 16to4_PriorityEncoder_v0p0p1_0.I11.t8 110.852
R24099 16to4_PriorityEncoder_v0p0p1_0.I11 16to4_PriorityEncoder_v0p0p1_0.I11.n12 84.2291
R24100 16to4_PriorityEncoder_v0p0p1_0.I11 16to4_PriorityEncoder_v0p0p1_0.I11.n11 82.1338
R24101 16to4_PriorityEncoder_v0p0p1_0.I11.n9 16to4_PriorityEncoder_v0p0p1_0.I11.n8 76.0005
R24102 16to4_PriorityEncoder_v0p0p1_0.I11.n10 16to4_PriorityEncoder_v0p0p1_0.I11 66.7187
R24103 16to4_PriorityEncoder_v0p0p1_0.I11.n13 16to4_PriorityEncoder_v0p0p1_0.I11 26.4877
R24104 16to4_PriorityEncoder_v0p0p1_0.I11.n1 16to4_PriorityEncoder_v0p0p1_0.I11.t0 17.6181
R24105 16to4_PriorityEncoder_v0p0p1_0.I11.n3 16to4_PriorityEncoder_v0p0p1_0.I11.t3 14.2865
R24106 16to4_PriorityEncoder_v0p0p1_0.I11.n5 16to4_PriorityEncoder_v0p0p1_0.I11.t1 14.283
R24107 16to4_PriorityEncoder_v0p0p1_0.I11.n5 16to4_PriorityEncoder_v0p0p1_0.I11.t2 14.283
R24108 16to4_PriorityEncoder_v0p0p1_0.I11.n7 16to4_PriorityEncoder_v0p0p1_0.I11.t4 8.77592
R24109 16to4_PriorityEncoder_v0p0p1_0.I11.n9 16to4_PriorityEncoder_v0p0p1_0.I11 7.31479
R24110 16to4_PriorityEncoder_v0p0p1_0.I11.n16 16to4_PriorityEncoder_v0p0p1_0.I11.n15 5.58999
R24111 16to4_PriorityEncoder_v0p0p1_0.I11.n13 16to4_PriorityEncoder_v0p0p1_0.I11 4.36044
R24112 16to4_PriorityEncoder_v0p0p1_0.I11 16to4_PriorityEncoder_v0p0p1_0.I11.n9 4.02336
R24113 16to4_PriorityEncoder_v0p0p1_0.I11.n14 16to4_PriorityEncoder_v0p0p1_0.I11.n13 2.71925
R24114 16to4_PriorityEncoder_v0p0p1_0.I11.n7 16to4_PriorityEncoder_v0p0p1_0.I11.n6 1.20426
R24115 16to4_PriorityEncoder_v0p0p1_0.I11.n14 16to4_PriorityEncoder_v0p0p1_0.I11.n10 1.15229
R24116 16to4_PriorityEncoder_v0p0p1_0.I11.n10 16to4_PriorityEncoder_v0p0p1_0.I11 0.969697
R24117 16to4_PriorityEncoder_v0p0p1_0.I11.n16 16to4_PriorityEncoder_v0p0p1_0.I11.n7 0.33431
R24118 16to4_PriorityEncoder_v0p0p1_0.I11.n15 16to4_PriorityEncoder_v0p0p1_0.I11.n14 0.31168
R24119 16to4_PriorityEncoder_v0p0p1_0.I11.n4 16to4_PriorityEncoder_v0p0p1_0.I11.n3 0.300242
R24120 16to4_PriorityEncoder_v0p0p1_0.I11.n15 16to4_PriorityEncoder_v0p0p1_0.I11 0.2005
R24121 16to4_PriorityEncoder_v0p0p1_0.I11.n2 16to4_PriorityEncoder_v0p0p1_0.I11.n0 0.159555
R24122 16to4_PriorityEncoder_v0p0p1_0.I11.n6 16to4_PriorityEncoder_v0p0p1_0.I11.n5 0.106617
R24123 16to4_PriorityEncoder_v0p0p1_0.I11.n4 16to4_PriorityEncoder_v0p0p1_0.I11.n2 0.0796167
R24124 16to4_PriorityEncoder_v0p0p1_0.I11.n6 16to4_PriorityEncoder_v0p0p1_0.I11.n4 0.0480595
R24125 16to4_PriorityEncoder_v0p0p1_0.I11 16to4_PriorityEncoder_v0p0p1_0.I11.n16 0.0087668
R24126 16to4_PriorityEncoder_v0p0p1_0.I11.n2 16to4_PriorityEncoder_v0p0p1_0.I11.n1 0.000504658
R24127 frontAnalog_v0p0p1_8.x63.A.n2 frontAnalog_v0p0p1_8.x63.A.t5 260.322
R24128 frontAnalog_v0p0p1_8.x63.A.n4 frontAnalog_v0p0p1_8.x63.A.t6 233.888
R24129 frontAnalog_v0p0p1_8.x63.A.n2 frontAnalog_v0p0p1_8.x63.A.t7 175.169
R24130 frontAnalog_v0p0p1_8.x63.A.n3 frontAnalog_v0p0p1_8.x63.A.t4 159.725
R24131 frontAnalog_v0p0p1_8.x63.A.n1 frontAnalog_v0p0p1_8.x63.A.t2 17.4109
R24132 frontAnalog_v0p0p1_8.x63.A.n0 frontAnalog_v0p0p1_8.x63.A.n2 9.75129
R24133 frontAnalog_v0p0p1_8.x63.A.n1 frontAnalog_v0p0p1_8.x63.A.t3 9.6037
R24134 frontAnalog_v0p0p1_8.x63.A.n0 frontAnalog_v0p0p1_8.x63.A 2.33338
R24135 frontAnalog_v0p0p1_8.x63.A.n5 frontAnalog_v0p0p1_8.x63.A.t0 8.40929
R24136 frontAnalog_v0p0p1_8.x63.A.n3 frontAnalog_v0p0p1_8.x63.A.t1 8.06629
R24137 frontAnalog_v0p0p1_8.x63.A.n4 frontAnalog_v0p0p1_8.x63.A.n3 1.73501
R24138 frontAnalog_v0p0p1_8.x63.A.n1 frontAnalog_v0p0p1_8.x63.A.n4 0.99025
R24139 frontAnalog_v0p0p1_8.x63.A.n5 frontAnalog_v0p0p1_8.x63.A.n1 0.853186
R24140 frontAnalog_v0p0p1_8.x63.A frontAnalog_v0p0p1_8.x63.A.n0 0.349517
R24141 frontAnalog_v0p0p1_8.x63.A frontAnalog_v0p0p1_8.x63.A.n5 0.24425
R24142 frontAnalog_v0p0p1_2.RSfetsym_0.QN.n1 frontAnalog_v0p0p1_2.RSfetsym_0.QN.t5 117.511
R24143 frontAnalog_v0p0p1_2.RSfetsym_0.QN.n1 frontAnalog_v0p0p1_2.RSfetsym_0.QN.t6 110.698
R24144 frontAnalog_v0p0p1_2.RSfetsym_0.QN.n4 frontAnalog_v0p0p1_2.RSfetsym_0.QN.t4 19.1963
R24145 frontAnalog_v0p0p1_2.RSfetsym_0.QN.n7 frontAnalog_v0p0p1_2.RSfetsym_0.QN.t1 14.2842
R24146 frontAnalog_v0p0p1_2.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_2.RSfetsym_0.QN.t2 14.283
R24147 frontAnalog_v0p0p1_2.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_2.RSfetsym_0.QN.t3 14.283
R24148 frontAnalog_v0p0p1_2.RSfetsym_0.QN.n11 frontAnalog_v0p0p1_2.RSfetsym_0.QN.t0 9.14075
R24149 frontAnalog_v0p0p1_2.RSfetsym_0.QN.n11 frontAnalog_v0p0p1_2.RSfetsym_0.QN.n10 0.74645
R24150 frontAnalog_v0p0p1_2.RSfetsym_0.QN.n2 frontAnalog_v0p0p1_2.RSfetsym_0.QN.n1 0.688382
R24151 frontAnalog_v0p0p1_2.RSfetsym_0.QN.n10 frontAnalog_v0p0p1_2.RSfetsym_0.QN.n9 0.2402
R24152 frontAnalog_v0p0p1_2.RSfetsym_0.QN.n9 frontAnalog_v0p0p1_2.RSfetsym_0.QN.n8 0.236824
R24153 frontAnalog_v0p0p1_2.RSfetsym_0.QN.n4 frontAnalog_v0p0p1_2.RSfetsym_0.QN.n3 0.132187
R24154 frontAnalog_v0p0p1_2.RSfetsym_0.QN.n9 frontAnalog_v0p0p1_2.RSfetsym_0.QN.n4 0.0968646
R24155 frontAnalog_v0p0p1_2.RSfetsym_0.QN frontAnalog_v0p0p1_2.RSfetsym_0.QN.n11 0.0446535
R24156 frontAnalog_v0p0p1_2.RSfetsym_0.QN.n8 frontAnalog_v0p0p1_2.RSfetsym_0.QN.n6 0.0272538
R24157 frontAnalog_v0p0p1_2.RSfetsym_0.QN.n10 frontAnalog_v0p0p1_2.RSfetsym_0.QN.n0 0.00981499
R24158 frontAnalog_v0p0p1_2.RSfetsym_0.QN.n3 frontAnalog_v0p0p1_2.RSfetsym_0.QN.n2 0.00725433
R24159 frontAnalog_v0p0p1_2.RSfetsym_0.QN.n6 frontAnalog_v0p0p1_2.RSfetsym_0.QN.n5 0.00610579
R24160 frontAnalog_v0p0p1_2.RSfetsym_0.QN.n8 frontAnalog_v0p0p1_2.RSfetsym_0.QN.n7 0.00225341
R24161 frontAnalog_v0p0p1_12.x65.A.n1 frontAnalog_v0p0p1_12.x65.A.t4 260.322
R24162 frontAnalog_v0p0p1_12.x65.A.n4 frontAnalog_v0p0p1_12.x65.A.t7 233.929
R24163 frontAnalog_v0p0p1_12.x65.A.n1 frontAnalog_v0p0p1_12.x65.A.t6 175.169
R24164 frontAnalog_v0p0p1_12.x65.A.n3 frontAnalog_v0p0p1_12.x65.A.t5 160.416
R24165 frontAnalog_v0p0p1_12.x65.A.n2 frontAnalog_v0p0p1_12.x65.A.t2 17.4109
R24166 frontAnalog_v0p0p1_12.x65.A.n2 frontAnalog_v0p0p1_12.x65.A.t3 10.2053
R24167 frontAnalog_v0p0p1_12.x65.A.n0 frontAnalog_v0p0p1_12.x65.A 2.78715
R24168 frontAnalog_v0p0p1_12.x65.A.n0 frontAnalog_v0p0p1_12.x65.A.n1 9.09103
R24169 frontAnalog_v0p0p1_12.x65.A.n6 frontAnalog_v0p0p1_12.x65.A.t1 7.94569
R24170 frontAnalog_v0p0p1_12.x65.A.n3 frontAnalog_v0p0p1_12.x65.A.t0 7.55846
R24171 frontAnalog_v0p0p1_12.x65.A.n5 frontAnalog_v0p0p1_12.x65.A.n4 1.4614
R24172 frontAnalog_v0p0p1_12.x65.A.n4 frontAnalog_v0p0p1_12.x65.A.n3 1.19626
R24173 frontAnalog_v0p0p1_12.x65.A.n6 frontAnalog_v0p0p1_12.x65.A.n5 0.836961
R24174 frontAnalog_v0p0p1_12.x65.A frontAnalog_v0p0p1_12.x65.A.n0 0.390342
R24175 frontAnalog_v0p0p1_12.x65.A.n5 frontAnalog_v0p0p1_12.x65.A.n2 0.154668
R24176 frontAnalog_v0p0p1_12.x65.A frontAnalog_v0p0p1_12.x65.A.n6 0.08175
R24177 frontAnalog_v0p0p1_6.x65.A.n1 frontAnalog_v0p0p1_6.x65.A.t6 260.322
R24178 frontAnalog_v0p0p1_6.x65.A.n4 frontAnalog_v0p0p1_6.x65.A.t5 233.929
R24179 frontAnalog_v0p0p1_6.x65.A.n1 frontAnalog_v0p0p1_6.x65.A.t7 175.169
R24180 frontAnalog_v0p0p1_6.x65.A.n3 frontAnalog_v0p0p1_6.x65.A.t4 160.416
R24181 frontAnalog_v0p0p1_6.x65.A.n2 frontAnalog_v0p0p1_6.x65.A.t3 17.4109
R24182 frontAnalog_v0p0p1_6.x65.A.n2 frontAnalog_v0p0p1_6.x65.A.t2 10.2053
R24183 frontAnalog_v0p0p1_6.x65.A.n0 frontAnalog_v0p0p1_6.x65.A 2.78715
R24184 frontAnalog_v0p0p1_6.x65.A.n0 frontAnalog_v0p0p1_6.x65.A.n1 9.09103
R24185 frontAnalog_v0p0p1_6.x65.A.n6 frontAnalog_v0p0p1_6.x65.A.t1 7.94569
R24186 frontAnalog_v0p0p1_6.x65.A.n3 frontAnalog_v0p0p1_6.x65.A.t0 7.55846
R24187 frontAnalog_v0p0p1_6.x65.A.n5 frontAnalog_v0p0p1_6.x65.A.n4 1.4614
R24188 frontAnalog_v0p0p1_6.x65.A.n4 frontAnalog_v0p0p1_6.x65.A.n3 1.19626
R24189 frontAnalog_v0p0p1_6.x65.A.n6 frontAnalog_v0p0p1_6.x65.A.n5 0.836961
R24190 frontAnalog_v0p0p1_6.x65.A frontAnalog_v0p0p1_6.x65.A.n0 0.390342
R24191 frontAnalog_v0p0p1_6.x65.A.n5 frontAnalog_v0p0p1_6.x65.A.n2 0.154668
R24192 frontAnalog_v0p0p1_6.x65.A frontAnalog_v0p0p1_6.x65.A.n6 0.08175
R24193 frontAnalog_v0p0p1_0.x65.A.n1 frontAnalog_v0p0p1_0.x65.A.t5 260.322
R24194 frontAnalog_v0p0p1_0.x65.A.n4 frontAnalog_v0p0p1_0.x65.A.t7 233.929
R24195 frontAnalog_v0p0p1_0.x65.A.n1 frontAnalog_v0p0p1_0.x65.A.t6 175.169
R24196 frontAnalog_v0p0p1_0.x65.A.n3 frontAnalog_v0p0p1_0.x65.A.t4 160.416
R24197 frontAnalog_v0p0p1_0.x65.A.n2 frontAnalog_v0p0p1_0.x65.A.t3 17.4109
R24198 frontAnalog_v0p0p1_0.x65.A.n2 frontAnalog_v0p0p1_0.x65.A.t2 10.2053
R24199 frontAnalog_v0p0p1_0.x65.A.n0 frontAnalog_v0p0p1_0.x65.A 2.78715
R24200 frontAnalog_v0p0p1_0.x65.A.n0 frontAnalog_v0p0p1_0.x65.A.n1 9.09103
R24201 frontAnalog_v0p0p1_0.x65.A.n6 frontAnalog_v0p0p1_0.x65.A.t1 7.94569
R24202 frontAnalog_v0p0p1_0.x65.A.n3 frontAnalog_v0p0p1_0.x65.A.t0 7.55846
R24203 frontAnalog_v0p0p1_0.x65.A.n5 frontAnalog_v0p0p1_0.x65.A.n4 1.4614
R24204 frontAnalog_v0p0p1_0.x65.A.n4 frontAnalog_v0p0p1_0.x65.A.n3 1.19626
R24205 frontAnalog_v0p0p1_0.x65.A.n6 frontAnalog_v0p0p1_0.x65.A.n5 0.836961
R24206 frontAnalog_v0p0p1_0.x65.A frontAnalog_v0p0p1_0.x65.A.n0 0.390342
R24207 frontAnalog_v0p0p1_0.x65.A.n5 frontAnalog_v0p0p1_0.x65.A.n2 0.154668
R24208 frontAnalog_v0p0p1_0.x65.A frontAnalog_v0p0p1_0.x65.A.n6 0.08175
R24209 frontAnalog_v0p0p1_0.x63.A.n2 frontAnalog_v0p0p1_0.x63.A.t5 260.322
R24210 frontAnalog_v0p0p1_0.x63.A.n4 frontAnalog_v0p0p1_0.x63.A.t4 233.888
R24211 frontAnalog_v0p0p1_0.x63.A.n2 frontAnalog_v0p0p1_0.x63.A.t6 175.169
R24212 frontAnalog_v0p0p1_0.x63.A.n3 frontAnalog_v0p0p1_0.x63.A.t7 159.725
R24213 frontAnalog_v0p0p1_0.x63.A.n1 frontAnalog_v0p0p1_0.x63.A.t2 17.4109
R24214 frontAnalog_v0p0p1_0.x63.A.n0 frontAnalog_v0p0p1_0.x63.A.n2 9.75129
R24215 frontAnalog_v0p0p1_0.x63.A.n1 frontAnalog_v0p0p1_0.x63.A.t3 9.6037
R24216 frontAnalog_v0p0p1_0.x63.A.n0 frontAnalog_v0p0p1_0.x63.A 2.33338
R24217 frontAnalog_v0p0p1_0.x63.A.n5 frontAnalog_v0p0p1_0.x63.A.t1 8.40929
R24218 frontAnalog_v0p0p1_0.x63.A.n3 frontAnalog_v0p0p1_0.x63.A.t0 8.06629
R24219 frontAnalog_v0p0p1_0.x63.A.n4 frontAnalog_v0p0p1_0.x63.A.n3 1.73501
R24220 frontAnalog_v0p0p1_0.x63.A.n1 frontAnalog_v0p0p1_0.x63.A.n4 0.99025
R24221 frontAnalog_v0p0p1_0.x63.A.n5 frontAnalog_v0p0p1_0.x63.A.n1 0.853186
R24222 frontAnalog_v0p0p1_0.x63.A frontAnalog_v0p0p1_0.x63.A.n0 0.349517
R24223 frontAnalog_v0p0p1_0.x63.A frontAnalog_v0p0p1_0.x63.A.n5 0.24425
C0 16to4_PriorityEncoder_v0p0p1_0.x3.EI a_77605_n52819# 0.175f
C1 a_77639_n50381# VDD 0.23f
C2 w_55000_n62950# resistorDivider_v0p0p1_0.V5 0.751f
C3 w_55000_n84550# VDD 0.829f
C4 frontAnalog_v0p0p1_12.x65.A VIN 0.655f
C5 16to4_PriorityEncoder_v0p0p1_0.x3.EI a_77639_n50381# 0.088f
C6 16to4_PriorityEncoder_v0p0p1_0.x3.x18.C 16to4_PriorityEncoder_v0p0p1_0.x3.x20.B 0.491f
C7 a_53630_n14796# VDD 0.134f
C8 16to4_PriorityEncoder_v0p0p1_0.x5.x19.C a_77605_n43545# 0.176f
C9 a_59578_n56970# VDD 0.0213f
C10 16to4_PriorityEncoder_v0p0p1_0.I12 a_59577_n19683# 0.29f
C11 frontAnalog_v0p0p1_14.RSfetsym_0.x1.Y VDD 0.733f
C12 16to4_PriorityEncoder_v0p0p1_0.I11 frontAnalog_v0p0p1_5.RSfetsym_0.x2.Y 0.198f
C13 a_78159_n47589# 16to4_PriorityEncoder_v0p0p1_0.x3.EO 0.128f
C14 frontAnalog_v0p0p1_14.x65.A a_55268_n79536# 0.461f
C15 m3_58396_n31350# VDD 1.3f
C16 a_53630_n79596# CLK 0.0136f
C17 frontAnalog_v0p0p1_11.x63.A a_55268_n63336# 1.24f
C18 a_77637_n48817# VDD 0.23f
C19 16to4_PriorityEncoder_v0p0p1_0.x3.x19.C 16to4_PriorityEncoder_v0p0p1_0.x3.x16.C 1.95f
C20 frontAnalog_v0p0p1_4.x63.X a_59577_n19683# 0.28f
C21 16to4_PriorityEncoder_v0p0p1_0.x28.A VDD 0.538f
C22 frontAnalog_v0p0p1_6.x65.X a_59578_n29970# 0.436f
C23 w_55000_n46128# frontAnalog_v0p0p1_8.x63.A 0.0792f
C24 frontAnalog_v0p0p1_9.RSfetsym_0.x1.Y frontAnalog_v0p0p1_9.x63.X 0.883f
C25 16to4_PriorityEncoder_v0p0p1_0.x3.x19.C a_77605_n52567# 0.157f
C26 frontAnalog_v0p0p1_0.x63.A VDD 3.67f
C27 a_53630_n9396# a_55268_n9336# 0.015f
C28 16to4_PriorityEncoder_v0p0p1_0.x3.EI a_77637_n48817# 0.0883f
C29 w_55000_n40728# CLK 0.571f
C30 frontAnalog_v0p0p1_5.x63.X frontAnalog_v0p0p1_5.RSfetsym_0.x2.Y 0.0923f
C31 a_53630_n9396# VIN 0.265f
C32 frontAnalog_v0p0p1_13.x65.X VDD 3.55f
C33 resistorDivider_v0p0p1_0.V16 CLK 4.89f
C34 16to4_PriorityEncoder_v0p0p1_0.x5.x21.B a_77605_n44779# 0.0141f
C35 w_55000_n8950# VDD 0.829f
C36 w_55000_n29928# a_53630_n30996# 0.359f
C37 a_57123_n79679# VDD 0.222f
C38 16to4_PriorityEncoder_v0p0p1_0.x43.A 16to4_PriorityEncoder_v0p0p1_0.x43.Y 1.52f
C39 frontAnalog_v0p0p1_5.RSfetsym_0.QN a_59577_n25083# 0.418f
C40 16to4_PriorityEncoder_v0p0p1_0.I12 m3_58396_n20550# 0.0416f
C41 a_53630_n84996# VIN 0.265f
C42 w_55000_n19128# frontAnalog_v0p0p1_4.x63.A 0.0792f
C43 w_55000_n25150# frontAnalog_v0p0p1_10.IB 0.0217f
C44 w_55000_n62328# frontAnalog_v0p0p1_11.x65.A 0.658f
C45 16to4_PriorityEncoder_v0p0p1_0.x5.x17.A 16to4_PriorityEncoder_v0p0p1_0.x5.x17.D 0.0198f
C46 16to4_PriorityEncoder_v0p0p1_0.x5.x22.A a_77605_n43295# 0.0116f
C47 frontAnalog_v0p0p1_10.RSfetsym_0.x1.Y VDD 0.733f
C48 frontAnalog_v0p0p1_14.RSfetsym_0.QN VDD 2.56f
C49 a_53630_n84996# a_55268_n84936# 0.015f
C50 16to4_PriorityEncoder_v0p0p1_0.x3.x22.A a_78065_n49349# 0.077f
C51 resistorDivider_v0p0p1_0.V7 a_53630_n52596# 0.28f
C52 frontAnalog_v0p0p1_13.x65.A a_55268_n68736# 0.461f
C53 frontAnalog_v0p0p1_4.x63.X m3_58396_n20550# 0.139f
C54 a_53630_n57996# CLK 0.0136f
C55 frontAnalog_v0p0p1_13.x63.X VDD 3.16f
C56 a_53630_n36396# VIN 0.265f
C57 w_55000_n62950# frontAnalog_v0p0p1_11.x63.A 0.659f
C58 frontAnalog_v0p0p1_6.x65.X frontAnalog_v0p0p1_6.RSfetsym_0.x1.Y 0.182f
C59 w_55000_n78528# a_55268_n79536# 0.149f
C60 w_55000_n79150# a_53630_n79596# 0.394f
C61 frontAnalog_v0p0p1_9.x65.X VDD 3.55f
C62 frontAnalog_v0p0p1_6.x65.A a_55268_n30936# 0.461f
C63 resistorDivider_v0p0p1_0.V11 VIN 2.52f
C64 w_55000_n19750# VIN 0.737f
C65 frontAnalog_v0p0p1_15.x65.A a_57123_n83559# 0.214f
C66 frontAnalog_v0p0p1_2.RSfetsym_0.QN a_59578_n2970# 0.255f
C67 frontAnalog_v0p0p1_10.IB resistorDivider_v0p0p1_0.V15 4.34f
C68 16to4_PriorityEncoder_v0p0p1_0.I11 a_77605_n44779# 0.15f
C69 frontAnalog_v0p0p1_2.x65.X 16to4_PriorityEncoder_v0p0p1_0.I15 0.445f
C70 16to4_PriorityEncoder_v0p0p1_0.x5.x17.D VDD 0.556f
C71 a_53630_n41796# VIN 0.265f
C72 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_6.x65.A 0.0352f
C73 a_57123_n58079# VDD 0.222f
C74 16to4_PriorityEncoder_v0p0p1_0.x1.X VDD 0.347f
C75 frontAnalog_v0p0p1_6.x65.X frontAnalog_v0p0p1_6.RSfetsym_0.QN 2.28f
C76 a_57123_n45759# frontAnalog_v0p0p1_8.x65.X 0.119f
C77 resistorDivider_v0p0p1_0.V6 resistorDivider_v0p0p1_0.V5 4.54f
C78 w_55000_n79150# CLK 0.535f
C79 16to4_PriorityEncoder_v0p0p1_0.x3.x20.B a_77605_n52819# 0.148f
C80 frontAnalog_v0p0p1_14.RSfetsym_0.x2.Y VDD 0.926f
C81 a_53630_n63396# VIN 0.265f
C82 frontAnalog_v0p0p1_10.IB resistorDivider_v0p0p1_0.V2 3.69f
C83 16to4_PriorityEncoder_v0p0p1_0.x3.x18.C a_77605_n52567# 0.117f
C84 resistorDivider_v0p0p1_0.V8 a_53630_n47196# 0.28f
C85 w_55000_n51528# VDD 0.854f
C86 a_53630_n36396# a_55268_n36336# 0.015f
C87 frontAnalog_v0p0p1_10.RSfetsym_0.QN VDD 2.56f
C88 a_53630_n74196# a_55268_n74136# 0.015f
C89 frontAnalog_v0p0p1_10.IB a_53630_n20196# 0.473f
C90 w_55000_n25150# resistorDivider_v0p0p1_0.V12 0.751f
C91 a_55268_n25536# VDD 0.565f
C92 w_55000_n67728# frontAnalog_v0p0p1_10.IB 0.0216f
C93 resistorDivider_v0p0p1_0.V1 frontAnalog_v0p0p1_15.x63.A 0.587f
C94 frontAnalog_v0p0p1_2.x65.X frontAnalog_v0p0p1_2.x63.X 0.136f
C95 16to4_PriorityEncoder_v0p0p1_0.x2.A 16to4_PriorityEncoder_v0p0p1_0.x3.GS 0.0652f
C96 16to4_PriorityEncoder_v0p0p1_0.x5.x17.A 16to4_PriorityEncoder_v0p0p1_0.x5.x17.C 0.0789f
C97 resistorDivider_v0p0p1_0.V3 resistorDivider_v0p0p1_0.V2 4.95f
C98 frontAnalog_v0p0p1_9.x63.A CLK 1.81f
C99 a_53630_n30996# VDD 0.134f
C100 frontAnalog_v0p0p1_12.x65.A a_57123_n72759# 0.214f
C101 frontAnalog_v0p0p1_10.IB resistorDivider_v0p0p1_0.V10 3.7f
C102 a_55268_n68736# CLK 0.236f
C103 frontAnalog_v0p0p1_10.IB resistorDivider_v0p0p1_0.V8 3.7f
C104 frontAnalog_v0p0p1_15.x63.A frontAnalog_v0p0p1_15.x63.X 0.0301f
C105 16to4_PriorityEncoder_v0p0p1_0.x3.x14.B a_78065_n49349# 0.202f
C106 w_55000_n3550# resistorDivider_v0p0p1_0.V16 0.751f
C107 w_55000_n3550# CLK 0.535f
C108 frontAnalog_v0p0p1_2.RSfetsym_0.QN frontAnalog_v0p0p1_2.RSfetsym_0.x1.Y 0.17f
C109 frontAnalog_v0p0p1_6.RSfetsym_0.x1.Y frontAnalog_v0p0p1_6.x63.X 0.883f
C110 frontAnalog_v0p0p1_10.RSfetsym_0.x2.Y VDD 0.926f
C111 a_53630_n41796# a_55268_n41736# 0.015f
C112 w_55000_n62328# VIN 0.866f
C113 16to4_PriorityEncoder_v0p0p1_0.I15 16to4_PriorityEncoder_v0p0p1_0.x5.x4.C 0.0129f
C114 16to4_PriorityEncoder_v0p0p1_0.x3.x22.A 16to4_PriorityEncoder_v0p0p1_0.x3.x17.A 1.27f
C115 a_77637_n49127# 16to4_PriorityEncoder_v0p0p1_0.x3.x22.A 0.0288f
C116 frontAnalog_v0p0p1_2.x65.A VDD 3.45f
C117 w_55000_n40728# frontAnalog_v0p0p1_1.x65.A 0.658f
C118 frontAnalog_v0p0p1_14.x63.A a_57123_n79679# 0.212f
C119 a_59577_n68283# VDD 0.0173f
C120 frontAnalog_v0p0p1_6.x65.X frontAnalog_v0p0p1_6.RSfetsym_0.x2.Y 0.526f
C121 a_55268_n74136# VIN 0.177f
C122 16to4_PriorityEncoder_v0p0p1_0.x5.x22.A 16to4_PriorityEncoder_v0p0p1_0.x5.x17.D 0.0732f
C123 a_53630_n63396# a_55268_n63336# 0.015f
C124 16to4_PriorityEncoder_v0p0p1_0.x5.x17.C VDD 0.272f
C125 frontAnalog_v0p0p1_6.RSfetsym_0.QN frontAnalog_v0p0p1_6.x63.X 0.378f
C126 frontAnalog_v0p0p1_1.x65.A CLK 2.61f
C127 a_78349_n51085# VDD 0.164f
C128 resistorDivider_v0p0p1_0.V6 frontAnalog_v0p0p1_10.x65.A 0.253f
C129 16to4_PriorityEncoder_v0p0p1_0.x3.x22.A 16to4_PriorityEncoder_v0p0p1_0.x3.x21.B 0.064f
C130 16to4_PriorityEncoder_v0p0p1_0.x3.x22.D VDD 0.242f
C131 w_55000_n41350# frontAnalog_v0p0p1_1.x63.A 0.659f
C132 16to4_PriorityEncoder_v0p0p1_0.I15 frontAnalog_v0p0p1_2.x63.X 1.78f
C133 resistorDivider_v0p0p1_0.V7 frontAnalog_v0p0p1_9.x65.A 0.252f
C134 a_55268_n52536# CLK 0.236f
C135 frontAnalog_v0p0p1_6.x63.X a_57123_n31079# 0.121f
C136 frontAnalog_v0p0p1_11.x65.A a_57123_n61959# 0.214f
C137 a_57123_n13359# VDD 0.224f
C138 frontAnalog_v0p0p1_4.x63.A VIN 0.194f
C139 w_55000_n56928# resistorDivider_v0p0p1_0.V6 0.798f
C140 frontAnalog_v0p0p1_12.x63.A frontAnalog_v0p0p1_12.x63.X 0.0301f
C141 16to4_PriorityEncoder_v0p0p1_0.x3.EI 16to4_PriorityEncoder_v0p0p1_0.x3.x22.D 0.208f
C142 frontAnalog_v0p0p1_6.x63.A resistorDivider_v0p0p1_0.V11 0.587f
C143 frontAnalog_v0p0p1_2.x63.A a_55268_n3936# 1.24f
C144 w_55000_n46750# frontAnalog_v0p0p1_8.x65.A 0.0988f
C145 16to4_PriorityEncoder_v0p0p1_0.x42.A 16to4_PriorityEncoder_v0p0p1_0.x43.A 0.392f
C146 frontAnalog_v0p0p1_14.x65.A frontAnalog_v0p0p1_14.x65.X 0.0236f
C147 w_55000_n19128# a_53630_n20196# 0.359f
C148 resistorDivider_v0p0p1_0.V5 VDD 4.19f
C149 m3_58396_n42150# VDD 1.3f
C150 16to4_PriorityEncoder_v0p0p1_0.I11 a_77605_n39305# 0.0597f
C151 w_55000_n46128# CLK 0.571f
C152 frontAnalog_v0p0p1_13.x63.A a_57123_n68879# 0.212f
C153 frontAnalog_v0p0p1_8.x63.X a_59577_n46683# 0.28f
C154 16to4_PriorityEncoder_v0p0p1_0.x3.A2 VDD 1.79f
C155 w_55000_n62950# a_53630_n63396# 0.394f
C156 w_55000_n19750# frontAnalog_v0p0p1_4.x65.A 0.0988f
C157 w_55000_n62328# a_55268_n63336# 0.149f
C158 16to4_PriorityEncoder_v0p0p1_0.x3.x18.C 16to4_PriorityEncoder_v0p0p1_0.x3.x19.C 2.6f
C159 w_55000_n14350# VDD 0.829f
C160 w_55000_n30550# a_55268_n30936# 0.12f
C161 16to4_PriorityEncoder_v0p0p1_0.x2.A 16to4_PriorityEncoder_v0p0p1_0.x3.EO 0.02f
C162 frontAnalog_v0p0p1_9.RSfetsym_0.QN frontAnalog_v0p0p1_9.RSfetsym_0.x2.Y 0.018f
C163 frontAnalog_v0p0p1_15.x63.A VDD 3.67f
C164 16to4_PriorityEncoder_v0p0p1_0.x5.x21.B 16to4_PriorityEncoder_v0p0p1_0.x5.x22.D 0.0561f
C165 16to4_PriorityEncoder_v0p0p1_0.x3.x14.B 16to4_PriorityEncoder_v0p0p1_0.x3.x17.A 0.125f
C166 a_77637_n49127# 16to4_PriorityEncoder_v0p0p1_0.x3.x14.B 0.109f
C167 w_55000_n30550# frontAnalog_v0p0p1_10.IB 0.0217f
C168 frontAnalog_v0p0p1_2.RSfetsym_0.x1.Y frontAnalog_v0p0p1_2.RSfetsym_0.x2.Y 0.0254f
C169 frontAnalog_v0p0p1_11.x63.A frontAnalog_v0p0p1_11.x63.X 0.0301f
C170 16to4_PriorityEncoder_v0p0p1_0.x5.x4.B 16to4_PriorityEncoder_v0p0p1_0.x5.x4.C 0.129f
C171 frontAnalog_v0p0p1_2.RSfetsym_0.QN frontAnalog_v0p0p1_2.RSfetsym_0.x2.Y 0.018f
C172 frontAnalog_v0p0p1_6.x63.X frontAnalog_v0p0p1_6.RSfetsym_0.x2.Y 0.0923f
C173 a_59578_n13770# VDD 0.0213f
C174 frontAnalog_v0p0p1_8.x65.X frontAnalog_v0p0p1_8.RSfetsym_0.QN 2.28f
C175 16to4_PriorityEncoder_v0p0p1_0.I14 frontAnalog_v0p0p1_3.RSfetsym_0.QN 0.0554f
C176 frontAnalog_v0p0p1_5.x65.A CLK 2.61f
C177 16to4_PriorityEncoder_v0p0p1_0.x5.x22.A 16to4_PriorityEncoder_v0p0p1_0.x5.x17.C 0.209f
C178 frontAnalog_v0p0p1_10.IB resistorDivider_v0p0p1_0.V9 3.69f
C179 frontAnalog_v0p0p1_13.x65.A frontAnalog_v0p0p1_13.x65.X 0.0236f
C180 16to4_PriorityEncoder_v0p0p1_0.x5.A2 16to4_PriorityEncoder_v0p0p1_0.x1.A 0.38f
C181 frontAnalog_v0p0p1_6.RSfetsym_0.QN a_59577_n30483# 0.418f
C182 frontAnalog_v0p0p1_6.x63.A a_57123_n31079# 0.212f
C183 frontAnalog_v0p0p1_9.RSfetsym_0.QN a_59577_n52083# 0.418f
C184 frontAnalog_v0p0p1_6.x65.A frontAnalog_v0p0p1_6.x65.X 0.0236f
C185 w_55000_n25150# VIN 0.737f
C186 16to4_PriorityEncoder_v0p0p1_0.I14 16to4_PriorityEncoder_v0p0p1_0.I11 0.782f
C187 a_77605_n53805# VDD 0.201f
C188 resistorDivider_v0p0p1_0.V1 a_53630_n84996# 0.28f
C189 w_55000_n62328# w_55000_n62950# 0.327f
C190 16to4_PriorityEncoder_v0p0p1_0.x5.x4.C 16to4_PriorityEncoder_v0p0p1_0.x5.EO 0.0749f
C191 16to4_PriorityEncoder_v0p0p1_0.I15 a_59577_n3483# 0.29f
C192 frontAnalog_v0p0p1_9.x63.A a_55268_n52536# 1.24f
C193 resistorDivider_v0p0p1_0.V14 VDD 4.05f
C194 frontAnalog_v0p0p1_11.x63.A VDD 3.67f
C195 16to4_PriorityEncoder_v0p0p1_0.x3.EI a_77605_n53805# 0.343f
C196 w_55000_n84550# CLK 0.535f
C197 frontAnalog_v0p0p1_10.x65.A VDD 3.45f
C198 w_55000_n68350# resistorDivider_v0p0p1_0.V4 0.751f
C199 16to4_PriorityEncoder_v0p0p1_0.x3.x22.B VDD 0.501f
C200 16to4_PriorityEncoder_v0p0p1_0.x5.GS 16to4_PriorityEncoder_v0p0p1_0.x43.A 0.0166f
C201 a_53630_n14796# CLK 0.0136f
C202 a_77637_n48817# 16to4_PriorityEncoder_v0p0p1_0.x3.x14.A 0.135f
C203 frontAnalog_v0p0p1_3.RSfetsym_0.x1.Y VDD 0.733f
C204 w_55000_n56928# VDD 0.854f
C205 a_55268_n47136# VDD 0.565f
C206 a_55268_n9336# resistorDivider_v0p0p1_0.V15 0.215f
C207 frontAnalog_v0p0p1_5.x65.X VDD 3.55f
C208 16to4_PriorityEncoder_v0p0p1_0.x3.A0 16to4_PriorityEncoder_v0p0p1_0.x3.x22.D 0.0149f
C209 16to4_PriorityEncoder_v0p0p1_0.x5.x21.B VDD 0.923f
C210 w_55000_n73128# frontAnalog_v0p0p1_10.IB 0.0216f
C211 16to4_PriorityEncoder_v0p0p1_0.I13 a_77605_n40069# 0.16f
C212 resistorDivider_v0p0p1_0.V15 VIN 2.56f
C213 frontAnalog_v0p0p1_6.x65.A VIN 0.655f
C214 resistorDivider_v0p0p1_0.V4 VDD 4.13f
C215 frontAnalog_v0p0p1_0.x63.A CLK 1.8f
C216 frontAnalog_v0p0p1_2.x63.X a_59577_n3483# 0.28f
C217 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3 7.92f
C218 a_57123_n29559# VDD 0.224f
C219 16to4_PriorityEncoder_v0p0p1_0.x5.x9.Y 16to4_PriorityEncoder_v0p0p1_0.x5.x4.C 0.125f
C220 resistorDivider_v0p0p1_0.V2 VIN 2.58f
C221 w_55000_n29928# resistorDivider_v0p0p1_0.V11 0.798f
C222 w_55000_n24528# w_55000_n25150# 0.327f
C223 16to4_PriorityEncoder_v0p0p1_0.x3.x19.C a_77605_n52819# 0.102f
C224 16to4_PriorityEncoder_v0p0p1_0.x3.x17.A a_77637_n50057# 0.14f
C225 frontAnalog_v0p0p1_13.x65.X CLK 0.0407f
C226 frontAnalog_v0p0p1_4.x63.A frontAnalog_v0p0p1_4.x65.A 3.16f
C227 w_55000_n73128# frontAnalog_v0p0p1_12.x63.A 0.0792f
C228 frontAnalog_v0p0p1_12.x65.A VDD 3.45f
C229 w_55000_n8950# CLK 0.535f
C230 a_57123_n14879# VDD 0.222f
C231 frontAnalog_v0p0p1_3.RSfetsym_0.QN VDD 2.56f
C232 a_53630_n20196# VIN 0.265f
C233 frontAnalog_v0p0p1_10.IB a_55268_n3936# 0.0848f
C234 w_55000_n67728# VIN 0.866f
C235 a_59578_n51570# VDD 0.0213f
C236 w_55000_n73128# resistorDivider_v0p0p1_0.V3 0.798f
C237 16to4_PriorityEncoder_v0p0p1_0.x5.x21.B 16to4_PriorityEncoder_v0p0p1_0.x5.x22.B 0.0197f
C238 frontAnalog_v0p0p1_1.x63.X a_59577_n41283# 0.28f
C239 16to4_PriorityEncoder_v0p0p1_0.x3.x14.B 16to4_PriorityEncoder_v0p0p1_0.x3.x22.A 0.0936f
C240 16to4_PriorityEncoder_v0p0p1_0.x3.x22.C VDD 0.892f
C241 resistorDivider_v0p0p1_0.V10 VIN 2.56f
C242 resistorDivider_v0p0p1_0.V8 VIN 2.62f
C243 frontAnalog_v0p0p1_9.RSfetsym_0.x1.Y frontAnalog_v0p0p1_9.RSfetsym_0.x2.Y 0.0254f
C244 16to4_PriorityEncoder_v0p0p1_0.x29.A 16to4_PriorityEncoder_v0p0p1_0.x29.Y 1.51f
C245 frontAnalog_v0p0p1_2.x65.A a_57123_n2559# 0.214f
C246 16to4_PriorityEncoder_v0p0p1_0.x3.EI 16to4_PriorityEncoder_v0p0p1_0.x3.x22.C 0.0149f
C247 frontAnalog_v0p0p1_13.x63.X CLK 0.785f
C248 a_53630_n9396# VDD 0.134f
C249 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_7.x65.A 0.0352f
C250 16to4_PriorityEncoder_v0p0p1_0.I11 VDD 9.88f
C251 16to4_PriorityEncoder_v0p0p1_0.x3.x4.B 16to4_PriorityEncoder_v0p0p1_0.x3.x4.C 0.129f
C252 16to4_PriorityEncoder_v0p0p1_0.x5.GS 16to4_PriorityEncoder_v0p0p1_0.x42.A 0.098f
C253 frontAnalog_v0p0p1_9.x65.X CLK 0.0407f
C254 frontAnalog_v0p0p1_1.x65.X a_59578_n40770# 0.436f
C255 frontAnalog_v0p0p1_3.x65.A a_55268_n14736# 0.461f
C256 a_53630_n84996# VDD 0.134f
C257 frontAnalog_v0p0p1_5.x63.X VDD 3.16f
C258 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_13.x63.A 0.0926f
C259 16to4_PriorityEncoder_v0p0p1_0.x5.x22.A 16to4_PriorityEncoder_v0p0p1_0.x5.x21.B 0.064f
C260 frontAnalog_v0p0p1_3.RSfetsym_0.x2.Y VDD 0.926f
C261 w_55000_n19750# a_55268_n20136# 0.12f
C262 w_55000_n2928# frontAnalog_v0p0p1_2.x63.A 0.0792f
C263 a_59578_n29970# VDD 0.0213f
C264 m3_58396_n52950# VDD 1.3f
C265 a_55268_n36336# resistorDivider_v0p0p1_0.V10 0.215f
C266 16to4_PriorityEncoder_v0p0p1_0.x5.x9.Y 16to4_PriorityEncoder_v0p0p1_0.x5.x4.B 0.118f
C267 16to4_PriorityEncoder_v0p0p1_0.x3.x20.B a_77605_n53805# 0.0838f
C268 w_55000_n51528# CLK 0.571f
C269 frontAnalog_v0p0p1_10.IB resistorDivider_v0p0p1_0.V13 3.7f
C270 frontAnalog_v0p0p1_8.x63.A a_55268_n47136# 1.24f
C271 16to4_PriorityEncoder_v0p0p1_0.x3.x4.C 16to4_PriorityEncoder_v0p0p1_0.x3.EO 0.0749f
C272 a_57123_n7959# frontAnalog_v0p0p1_0.x65.X 0.119f
C273 a_53630_n36396# VDD 0.134f
C274 a_55268_n25536# CLK 0.236f
C275 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_8.x65.A 0.0352f
C276 w_55000_n13728# frontAnalog_v0p0p1_3.x65.A 0.658f
C277 resistorDivider_v0p0p1_0.V11 VDD 4.38f
C278 w_55000_n19750# VDD 0.829f
C279 16to4_PriorityEncoder_v0p0p1_0.x3.EO 16to4_PriorityEncoder_v0p0p1_0.x3.GS 0.9f
C280 frontAnalog_v0p0p1_6.x63.A frontAnalog_v0p0p1_6.x65.A 3.16f
C281 a_53630_n30996# CLK 0.0136f
C282 w_55000_n35950# frontAnalog_v0p0p1_10.IB 0.0217f
C283 16to4_PriorityEncoder_v0p0p1_0.I15 16to4_PriorityEncoder_v0p0p1_0.x5.x20.B 0.244f
C284 a_53630_n41796# VDD 0.134f
C285 16to4_PriorityEncoder_v0p0p1_0.x5.EO 16to4_PriorityEncoder_v0p0p1_0.x5.GS 0.927f
C286 16to4_PriorityEncoder_v0p0p1_0.x3.x17.A 16to4_PriorityEncoder_v0p0p1_0.x3.x17.D 0.0198f
C287 16to4_PriorityEncoder_v0p0p1_0.x5.x9.Y 16to4_PriorityEncoder_v0p0p1_0.x5.EO 0.0491f
C288 a_53630_n63396# VDD 0.134f
C289 16to4_PriorityEncoder_v0p0p1_0.x5.x20.B 16to4_PriorityEncoder_v0p0p1_0.x5.x4.C 0.014f
C290 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_14.x65.A 0.0352f
C291 w_55000_n14350# frontAnalog_v0p0p1_3.x63.A 0.659f
C292 a_57123_n83559# frontAnalog_v0p0p1_15.x65.X 0.119f
C293 frontAnalog_v0p0p1_9.x65.A a_57123_n51159# 0.214f
C294 16to4_PriorityEncoder_v0p0p1_0.x3.x17.D 16to4_PriorityEncoder_v0p0p1_0.x3.x21.B 0.0218f
C295 frontAnalog_v0p0p1_6.RSfetsym_0.x1.Y VDD 0.733f
C296 frontAnalog_v0p0p1_2.x65.A resistorDivider_v0p0p1_0.V16 0.252f
C297 16to4_PriorityEncoder_v0p0p1_0.x3.A1 a_78349_n51085# 0.151f
C298 a_59578_n40770# VDD 0.0213f
C299 frontAnalog_v0p0p1_2.x65.A CLK 2.61f
C300 w_55000_n30550# VIN 0.737f
C301 a_78525_n53555# VDD 0.151f
C302 resistorDivider_v0p0p1_0.V9 VIN 2.55f
C303 frontAnalog_v0p0p1_8.x65.X frontAnalog_v0p0p1_8.RSfetsym_0.x1.Y 0.182f
C304 resistorDivider_v0p0p1_0.V13 resistorDivider_v0p0p1_0.V12 4.41f
C305 frontAnalog_v0p0p1_2.x63.A frontAnalog_v0p0p1_2.x63.X 0.0301f
C306 frontAnalog_v0p0p1_6.RSfetsym_0.QN VDD 2.56f
C307 w_55000_n52150# resistorDivider_v0p0p1_0.V7 0.751f
C308 a_59577_n25083# VDD 0.0173f
C309 16to4_PriorityEncoder_v0p0p1_0.x3.x20.B 16to4_PriorityEncoder_v0p0p1_0.x3.x22.C 0.0195f
C310 frontAnalog_v0p0p1_0.x65.X a_59578_n8370# 0.436f
C311 w_55000_n73128# a_53630_n74196# 0.359f
C312 frontAnalog_v0p0p1_15.x65.X a_59578_n83970# 0.436f
C313 w_55000_n19128# resistorDivider_v0p0p1_0.V13 0.798f
C314 16to4_PriorityEncoder_v0p0p1_0.x3.A0 16to4_PriorityEncoder_v0p0p1_0.x3.x22.C 0.0123f
C315 a_77605_n43545# VDD 0.571f
C316 frontAnalog_v0p0p1_3.x63.A resistorDivider_v0p0p1_0.V14 0.587f
C317 a_57123_n31079# VDD 0.222f
C318 w_55000_n62328# VDD 0.854f
C319 frontAnalog_v0p0p1_8.x65.X VDD 3.55f
C320 16to4_PriorityEncoder_v0p0p1_0.x3.x22.A a_77605_n51335# 0.0116f
C321 a_57123_n34959# frontAnalog_v0p0p1_7.x65.X 0.119f
C322 a_57123_n72759# frontAnalog_v0p0p1_12.x65.X 0.119f
C323 16to4_PriorityEncoder_v0p0p1_0.x3.A2 16to4_PriorityEncoder_v0p0p1_0.x3.x14.A 0.074f
C324 w_55000_n51528# frontAnalog_v0p0p1_9.x63.A 0.0792f
C325 resistorDivider_v0p0p1_0.V5 CLK 5.47f
C326 w_55000_n78528# frontAnalog_v0p0p1_10.IB 0.0216f
C327 w_55000_n73750# frontAnalog_v0p0p1_12.x65.A 0.0988f
C328 frontAnalog_v0p0p1_4.x63.A a_55268_n20136# 1.24f
C329 w_55000_n35328# a_53630_n36396# 0.359f
C330 a_55268_n74136# VDD 0.565f
C331 16to4_PriorityEncoder_v0p0p1_0.x3.A2 16to4_PriorityEncoder_v0p0p1_0.x3.A1 0.787f
C332 16to4_PriorityEncoder_v0p0p1_0.x3.x17.A 16to4_PriorityEncoder_v0p0p1_0.x3.x17.C 0.0789f
C333 a_78097_n45737# 16to4_PriorityEncoder_v0p0p1_0.x5.x22.D 0.137f
C334 frontAnalog_v0p0p1_10.IB resistorDivider_v0p0p1_0.V7 3.69f
C335 16to4_PriorityEncoder_v0p0p1_0.x28.A 16to4_PriorityEncoder_v0p0p1_0.x29.A 0.392f
C336 16to4_PriorityEncoder_v0p0p1_0.x5.x14.A 16to4_PriorityEncoder_v0p0p1_0.x5.A2 0.074f
C337 16to4_PriorityEncoder_v0p0p1_0.I15 16to4_PriorityEncoder_v0p0p1_0.x5.x16.C 0.26f
C338 w_55000_n14350# CLK 0.535f
C339 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_3.x65.A 0.0352f
C340 frontAnalog_v0p0p1_15.x63.A CLK 1.81f
C341 frontAnalog_v0p0p1_1.RSfetsym_0.QN a_59578_n40770# 0.255f
C342 frontAnalog_v0p0p1_4.x63.A VDD 3.67f
C343 a_55268_n41736# resistorDivider_v0p0p1_0.V9 0.215f
C344 w_55000_n73128# VIN 0.866f
C345 a_57123_n40359# frontAnalog_v0p0p1_1.x65.X 0.119f
C346 frontAnalog_v0p0p1_12.x65.X a_59578_n73170# 0.436f
C347 16to4_PriorityEncoder_v0p0p1_0.I14 a_59578_n8370# 0.42f
C348 frontAnalog_v0p0p1_15.x65.X frontAnalog_v0p0p1_15.RSfetsym_0.x1.Y 0.182f
C349 frontAnalog_v0p0p1_0.x65.X frontAnalog_v0p0p1_0.RSfetsym_0.x1.Y 0.182f
C350 resistorDivider_v0p0p1_0.V4 frontAnalog_v0p0p1_13.x65.A 0.253f
C351 frontAnalog_v0p0p1_10.IB a_53630_n68796# 0.473f
C352 16to4_PriorityEncoder_v0p0p1_0.x1.A 16to4_PriorityEncoder_v0p0p1_0.x2.A 0.304f
C353 w_55000_n2928# frontAnalog_v0p0p1_10.IB 0.0216f
C354 frontAnalog_v0p0p1_3.x63.A a_57123_n14879# 0.212f
C355 frontAnalog_v0p0p1_11.x63.X m3_58396_n63750# 0.139f
C356 frontAnalog_v0p0p1_9.x63.X VDD 3.16f
C357 16to4_PriorityEncoder_v0p0p1_0.x3.x22.A 16to4_PriorityEncoder_v0p0p1_0.x3.x17.D 0.0732f
C358 a_57123_n61959# frontAnalog_v0p0p1_11.x65.X 0.119f
C359 frontAnalog_v0p0p1_6.RSfetsym_0.x2.Y VDD 0.926f
C360 resistorDivider_v0p0p1_0.V2 resistorDivider_v0p0p1_0.V1 4.46f
C361 a_57123_n7959# VDD 0.224f
C362 w_55000_n52150# a_53630_n52596# 0.394f
C363 w_55000_n29928# frontAnalog_v0p0p1_6.x65.A 0.658f
C364 w_55000_n51528# a_55268_n52536# 0.149f
C365 frontAnalog_v0p0p1_0.x65.X frontAnalog_v0p0p1_0.RSfetsym_0.QN 2.28f
C366 frontAnalog_v0p0p1_14.RSfetsym_0.QN a_59578_n78570# 0.255f
C367 16to4_PriorityEncoder_v0p0p1_0.x5.x21.B 16to4_PriorityEncoder_v0p0p1_0.x5.x22.C 0.262f
C368 w_55000_n3550# frontAnalog_v0p0p1_2.x65.A 0.0988f
C369 a_55268_n3936# VIN 0.177f
C370 frontAnalog_v0p0p1_3.x65.A frontAnalog_v0p0p1_3.x65.X 0.0236f
C371 w_55000_n30550# frontAnalog_v0p0p1_6.x63.A 0.659f
C372 frontAnalog_v0p0p1_15.RSfetsym_0.x1.Y frontAnalog_v0p0p1_15.x63.X 0.883f
C373 a_57123_n83559# VDD 0.224f
C374 frontAnalog_v0p0p1_8.x65.A a_57123_n45759# 0.214f
C375 resistorDivider_v0p0p1_0.V14 CLK 6.32f
C376 frontAnalog_v0p0p1_11.x63.A CLK 1.81f
C377 frontAnalog_v0p0p1_10.x65.A CLK 2.61f
C378 frontAnalog_v0p0p1_7.x65.X a_59578_n35370# 0.436f
C379 frontAnalog_v0p0p1_11.x65.X a_59578_n62370# 0.436f
C380 m3_58396_n63750# VDD 1.3f
C381 a_78097_n45737# VDD 0.332f
C382 frontAnalog_v0p0p1_7.x65.A VIN 0.655f
C383 16to4_PriorityEncoder_v0p0p1_0.I12 16to4_PriorityEncoder_v0p0p1_0.I11 5.01f
C384 frontAnalog_v0p0p1_10.IB a_53630_n52596# 0.473f
C385 frontAnalog_v0p0p1_12.x65.X frontAnalog_v0p0p1_12.RSfetsym_0.x1.Y 0.182f
C386 16to4_PriorityEncoder_v0p0p1_0.I14 frontAnalog_v0p0p1_0.RSfetsym_0.x1.Y 0.0432f
C387 16to4_PriorityEncoder_v0p0p1_0.x5.x20.B 16to4_PriorityEncoder_v0p0p1_0.x5.x9.Y 0.0516f
C388 w_55000_n56928# CLK 0.571f
C389 frontAnalog_v0p0p1_15.x65.X frontAnalog_v0p0p1_15.RSfetsym_0.QN 2.28f
C390 w_55000_n8328# frontAnalog_v0p0p1_0.x65.A 0.658f
C391 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_1.x63.A 0.0926f
C392 16to4_PriorityEncoder_v0p0p1_0.x3.A0 a_78525_n53555# 0.149f
C393 a_55268_n47136# CLK 0.236f
C394 a_57123_n34959# VDD 0.224f
C395 frontAnalog_v0p0p1_14.x65.X frontAnalog_v0p0p1_14.x63.X 0.136f
C396 frontAnalog_v0p0p1_5.x65.X CLK 0.0398f
C397 frontAnalog_v0p0p1_10.IB a_55268_n79536# 0.0848f
C398 w_55000_n25150# VDD 0.829f
C399 resistorDivider_v0p0p1_0.V4 CLK 5.72f
C400 frontAnalog_v0p0p1_13.x63.A VIN 0.188f
C401 a_59578_n83970# VDD 0.0213f
C402 frontAnalog_v0p0p1_15.x63.X a_57123_n85079# 0.121f
C403 frontAnalog_v0p0p1_0.RSfetsym_0.x1.Y frontAnalog_v0p0p1_0.x63.X 0.883f
C404 frontAnalog_v0p0p1_13.RSfetsym_0.QN a_59578_n67770# 0.255f
C405 w_55000_n8950# frontAnalog_v0p0p1_0.x63.A 0.659f
C406 frontAnalog_v0p0p1_0.RSfetsym_0.QN 16to4_PriorityEncoder_v0p0p1_0.I14 2.02f
C407 a_57123_n40359# VDD 0.224f
C408 w_55000_n41350# frontAnalog_v0p0p1_10.IB 0.0217f
C409 frontAnalog_v0p0p1_14.RSfetsym_0.QN frontAnalog_v0p0p1_14.RSfetsym_0.x1.Y 0.17f
C410 a_78097_n45737# 16to4_PriorityEncoder_v0p0p1_0.x5.x22.B 0.109f
C411 frontAnalog_v0p0p1_3.x63.X m3_58396_n15150# 0.139f
C412 a_77605_n43295# 16to4_PriorityEncoder_v0p0p1_0.x5.x17.D 0.0121f
C413 16to4_PriorityEncoder_v0p0p1_0.x3.x22.A 16to4_PriorityEncoder_v0p0p1_0.x3.x17.C 0.209f
C414 frontAnalog_v0p0p1_12.RSfetsym_0.x1.Y frontAnalog_v0p0p1_12.x63.X 0.883f
C415 16to4_PriorityEncoder_v0p0p1_0.I13 m3_58396_n15150# 0.0416f
C416 a_57123_n61959# VDD 0.224f
C417 frontAnalog_v0p0p1_5.x65.A a_55268_n25536# 0.461f
C418 w_55000_n56928# a_53630_n57996# 0.359f
C419 resistorDivider_v0p0p1_0.V13 VIN 2.58f
C420 a_59578_n8370# VDD 0.0213f
C421 a_78065_n41309# 16to4_PriorityEncoder_v0p0p1_0.x5.A2 0.144f
C422 frontAnalog_v0p0p1_12.x65.A CLK 2.61f
C423 frontAnalog_v0p0p1_0.x65.X frontAnalog_v0p0p1_0.RSfetsym_0.x2.Y 0.526f
C424 frontAnalog_v0p0p1_0.RSfetsym_0.QN frontAnalog_v0p0p1_0.x63.X 0.378f
C425 frontAnalog_v0p0p1_15.x65.X frontAnalog_v0p0p1_15.RSfetsym_0.x2.Y 0.526f
C426 frontAnalog_v0p0p1_7.x65.A a_55268_n36336# 0.461f
C427 frontAnalog_v0p0p1_15.RSfetsym_0.QN frontAnalog_v0p0p1_15.x63.X 0.378f
C428 frontAnalog_v0p0p1_10.x63.A a_55268_n57936# 1.24f
C429 frontAnalog_v0p0p1_8.x63.X m3_58396_n47550# 0.139f
C430 frontAnalog_v0p0p1_8.x65.A VIN 0.654f
C431 frontAnalog_v0p0p1_11.x65.X frontAnalog_v0p0p1_11.RSfetsym_0.x1.Y 0.182f
C432 frontAnalog_v0p0p1_7.x65.X frontAnalog_v0p0p1_7.RSfetsym_0.QN 2.28f
C433 frontAnalog_v0p0p1_7.x65.X frontAnalog_v0p0p1_7.RSfetsym_0.x1.Y 0.182f
C434 frontAnalog_v0p0p1_12.x65.X frontAnalog_v0p0p1_12.RSfetsym_0.QN 2.28f
C435 frontAnalog_v0p0p1_6.x65.A VDD 3.45f
C436 frontAnalog_v0p0p1_0.x63.X a_57123_n9479# 0.121f
C437 resistorDivider_v0p0p1_0.V15 VDD 4.05f
C438 a_53630_n20196# a_55268_n20136# 0.015f
C439 w_55000_n35950# VIN 0.737f
C440 frontAnalog_v0p0p1_13.x65.X frontAnalog_v0p0p1_13.x63.X 0.136f
C441 frontAnalog_v0p0p1_14.RSfetsym_0.x1.Y frontAnalog_v0p0p1_14.RSfetsym_0.x2.Y 0.0254f
C442 resistorDivider_v0p0p1_0.V2 VDD 4.22f
C443 w_55000_n67728# w_55000_n68350# 0.327f
C444 16to4_PriorityEncoder_v0p0p1_0.I15 16to4_PriorityEncoder_v0p0p1_0.x5.x19.C 0.239f
C445 a_53630_n9396# CLK 0.0136f
C446 frontAnalog_v0p0p1_10.IB a_55268_n57936# 0.0848f
C447 frontAnalog_v0p0p1_14.x65.A VIN 0.655f
C448 a_59578_n62370# VDD 0.0213f
C449 16to4_PriorityEncoder_v0p0p1_0.I11 CLK 0.01f
C450 frontAnalog_v0p0p1_12.x63.X a_57123_n74279# 0.121f
C451 frontAnalog_v0p0p1_15.RSfetsym_0.x1.Y VDD 0.733f
C452 a_59577_n41283# VDD 0.0173f
C453 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_5.x63.A 0.0926f
C454 frontAnalog_v0p0p1_15.x63.X frontAnalog_v0p0p1_15.RSfetsym_0.x2.Y 0.0923f
C455 frontAnalog_v0p0p1_10.RSfetsym_0.QN a_59578_n56970# 0.255f
C456 16to4_PriorityEncoder_v0p0p1_0.x1.X 16to4_PriorityEncoder_v0p0p1_0.x28.A 0.0747f
C457 w_55000_n73750# a_55268_n74136# 0.12f
C458 w_55000_n52150# frontAnalog_v0p0p1_9.x65.A 0.0988f
C459 frontAnalog_v0p0p1_4.x65.A a_57123_n18759# 0.214f
C460 frontAnalog_v0p0p1_13.RSfetsym_0.QN frontAnalog_v0p0p1_13.RSfetsym_0.x1.Y 0.17f
C461 a_53630_n84996# CLK 0.0136f
C462 16to4_PriorityEncoder_v0p0p1_0.I14 a_77605_n40069# 0.214f
C463 a_53630_n20196# VDD 0.134f
C464 frontAnalog_v0p0p1_5.x63.X CLK 0.785f
C465 frontAnalog_v0p0p1_11.RSfetsym_0.x1.Y frontAnalog_v0p0p1_11.x63.X 0.883f
C466 w_55000_n67728# VDD 0.854f
C467 frontAnalog_v0p0p1_12.RSfetsym_0.QN frontAnalog_v0p0p1_12.x63.X 0.378f
C468 frontAnalog_v0p0p1_12.x65.X frontAnalog_v0p0p1_12.RSfetsym_0.x2.Y 0.526f
C469 frontAnalog_v0p0p1_0.RSfetsym_0.x1.Y VDD 0.733f
C470 16to4_PriorityEncoder_v0p0p1_0.I15 16to4_PriorityEncoder_v0p0p1_0.I13 1.14f
C471 16to4_PriorityEncoder_v0p0p1_0.I14 frontAnalog_v0p0p1_0.RSfetsym_0.x2.Y 0.195f
C472 a_59578_n35370# VDD 0.0213f
C473 w_55000_n83928# frontAnalog_v0p0p1_10.IB 0.0216f
C474 resistorDivider_v0p0p1_0.V10 VDD 4.56f
C475 w_55000_n35950# a_55268_n36336# 0.12f
C476 frontAnalog_v0p0p1_12.x65.X VDD 3.55f
C477 16to4_PriorityEncoder_v0p0p1_0.x3.x21.B a_78097_n53777# 0.186f
C478 resistorDivider_v0p0p1_0.V8 VDD 4.18f
C479 a_77605_n43295# 16to4_PriorityEncoder_v0p0p1_0.x5.x17.C 0.0951f
C480 frontAnalog_v0p0p1_11.x65.X frontAnalog_v0p0p1_11.RSfetsym_0.QN 2.28f
C481 w_55000_n29928# w_55000_n30550# 0.327f
C482 a_53630_n36396# CLK 0.0136f
C483 a_57123_n85079# VDD 0.222f
C484 frontAnalog_v0p0p1_0.x63.X frontAnalog_v0p0p1_0.RSfetsym_0.x2.Y 0.0923f
C485 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_9.x65.A 0.0352f
C486 frontAnalog_v0p0p1_10.x65.X frontAnalog_v0p0p1_10.x63.X 0.136f
C487 frontAnalog_v0p0p1_0.RSfetsym_0.QN VDD 2.56f
C488 frontAnalog_v0p0p1_13.RSfetsym_0.x1.Y frontAnalog_v0p0p1_13.RSfetsym_0.x2.Y 0.0254f
C489 resistorDivider_v0p0p1_0.V4 a_55268_n68736# 0.215f
C490 resistorDivider_v0p0p1_0.V11 CLK 6.86f
C491 w_55000_n19750# CLK 0.535f
C492 w_55000_n40728# a_53630_n41796# 0.359f
C493 frontAnalog_v0p0p1_11.x63.X a_57123_n63479# 0.121f
C494 frontAnalog_v0p0p1_14.RSfetsym_0.QN frontAnalog_v0p0p1_14.RSfetsym_0.x2.Y 0.018f
C495 frontAnalog_v0p0p1_11.RSfetsym_0.x1.Y VDD 0.733f
C496 frontAnalog_v0p0p1_12.x63.X frontAnalog_v0p0p1_12.RSfetsym_0.x2.Y 0.0923f
C497 a_53630_n41796# CLK 0.0136f
C498 a_82906_n51645# VDD 0.18f
C499 frontAnalog_v0p0p1_15.RSfetsym_0.QN VDD 2.56f
C500 16to4_PriorityEncoder_v0p0p1_0.x5.x17.A 16to4_PriorityEncoder_v0p0p1_0.x5.A2 0.047f
C501 a_57123_n9479# VDD 0.222f
C502 w_55000_n78528# VIN 0.866f
C503 frontAnalog_v0p0p1_10.RSfetsym_0.QN frontAnalog_v0p0p1_10.RSfetsym_0.x1.Y 0.17f
C504 frontAnalog_v0p0p1_0.RSfetsym_0.QN a_59577_n8883# 0.418f
C505 frontAnalog_v0p0p1_15.RSfetsym_0.QN a_59577_n84483# 0.418f
C506 frontAnalog_v0p0p1_14.x63.X a_59577_n79083# 0.28f
C507 a_53630_n63396# CLK 0.0136f
C508 frontAnalog_v0p0p1_12.x63.X VDD 3.16f
C509 16to4_PriorityEncoder_v0p0p1_0.I15 16to4_PriorityEncoder_v0p0p1_0.x5.x18.C 0.229f
C510 resistorDivider_v0p0p1_0.V7 VIN 2.61f
C511 frontAnalog_v0p0p1_1.RSfetsym_0.QN a_59577_n41283# 0.418f
C512 w_55000_n8328# frontAnalog_v0p0p1_10.IB 0.0216f
C513 frontAnalog_v0p0p1_11.x65.X frontAnalog_v0p0p1_11.RSfetsym_0.x2.Y 0.526f
C514 frontAnalog_v0p0p1_8.x65.X a_59578_n46170# 0.436f
C515 frontAnalog_v0p0p1_7.RSfetsym_0.x1.Y frontAnalog_v0p0p1_7.x63.X 0.883f
C516 frontAnalog_v0p0p1_11.RSfetsym_0.QN frontAnalog_v0p0p1_11.x63.X 0.378f
C517 frontAnalog_v0p0p1_7.RSfetsym_0.QN frontAnalog_v0p0p1_7.x63.X 0.378f
C518 frontAnalog_v0p0p1_5.x63.A resistorDivider_v0p0p1_0.V12 0.587f
C519 frontAnalog_v0p0p1_7.x65.X frontAnalog_v0p0p1_7.RSfetsym_0.x2.Y 0.526f
C520 a_78159_n39549# VDD 0.155f
C521 a_82906_n51645# 16to4_PriorityEncoder_v0p0p1_0.x2.X 0.12f
C522 frontAnalog_v0p0p1_7.x63.A resistorDivider_v0p0p1_0.V10 0.587f
C523 frontAnalog_v0p0p1_3.x65.A VIN 0.655f
C524 frontAnalog_v0p0p1_7.RSfetsym_0.QN VDD 2.56f
C525 frontAnalog_v0p0p1_7.RSfetsym_0.x1.Y VDD 0.733f
C526 a_57123_n63479# VDD 0.222f
C527 w_55000_n83928# frontAnalog_v0p0p1_15.x65.A 0.658f
C528 16to4_PriorityEncoder_v0p0p1_0.x5.A2 VDD 3.08f
C529 frontAnalog_v0p0p1_15.RSfetsym_0.x2.Y VDD 0.926f
C530 frontAnalog_v0p0p1_10.RSfetsym_0.x1.Y frontAnalog_v0p0p1_10.RSfetsym_0.x2.Y 0.0254f
C531 a_53630_n68796# VIN 0.265f
C532 frontAnalog_v0p0p1_4.x65.A resistorDivider_v0p0p1_0.V13 0.253f
C533 frontAnalog_v0p0p1_4.x63.A frontAnalog_v0p0p1_4.x63.X 0.0301f
C534 a_77605_n51335# 16to4_PriorityEncoder_v0p0p1_0.x3.x17.D 0.0121f
C535 w_55000_n2928# VIN 0.867f
C536 frontAnalog_v0p0p1_13.RSfetsym_0.QN frontAnalog_v0p0p1_13.RSfetsym_0.x2.Y 0.018f
C537 a_77605_n40069# VDD 0.156f
C538 16to4_PriorityEncoder_v0p0p1_0.x3.EI 16to4_PriorityEncoder_v0p0p1_0.x5.A2 0.507f
C539 frontAnalog_v0p0p1_7.x63.X a_57123_n36479# 0.121f
C540 frontAnalog_v0p0p1_11.x63.X frontAnalog_v0p0p1_11.RSfetsym_0.x2.Y 0.0923f
C541 frontAnalog_v0p0p1_11.RSfetsym_0.QN VDD 2.56f
C542 m3_58396_n74550# VDD 1.3f
C543 w_55000_n46128# a_55268_n47136# 0.149f
C544 frontAnalog_v0p0p1_12.RSfetsym_0.QN a_59577_n73683# 0.418f
C545 w_55000_n84550# frontAnalog_v0p0p1_15.x63.A 0.659f
C546 w_55000_n46750# a_53630_n47196# 0.394f
C547 w_55000_n13728# a_55268_n14736# 0.149f
C548 w_55000_n14350# a_53630_n14796# 0.394f
C549 frontAnalog_v0p0p1_0.RSfetsym_0.x2.Y VDD 0.926f
C550 resistorDivider_v0p0p1_0.V2 frontAnalog_v0p0p1_14.x63.A 0.587f
C551 w_55000_n62328# CLK 0.571f
C552 frontAnalog_v0p0p1_13.x63.X a_59577_n68283# 0.28f
C553 w_55000_n35328# resistorDivider_v0p0p1_0.V10 0.798f
C554 a_57123_n36479# VDD 0.222f
C555 frontAnalog_v0p0p1_8.x65.X CLK 0.0393f
C556 resistorDivider_v0p0p1_0.V8 frontAnalog_v0p0p1_8.x63.A 0.587f
C557 w_55000_n30550# VDD 0.829f
C558 a_55268_n74136# CLK 0.236f
C559 resistorDivider_v0p0p1_0.V9 VDD 4.76f
C560 16to4_PriorityEncoder_v0p0p1_0.x5.x16.C 16to4_PriorityEncoder_v0p0p1_0.x5.x20.B 1.24f
C561 frontAnalog_v0p0p1_10.x65.A a_57123_n56559# 0.214f
C562 w_55000_n46750# frontAnalog_v0p0p1_10.IB 0.0217f
C563 a_53630_n52596# VIN 0.265f
C564 frontAnalog_v0p0p1_5.x63.A a_57123_n25679# 0.212f
C565 frontAnalog_v0p0p1_11.RSfetsym_0.x2.Y VDD 0.926f
C566 16to4_PriorityEncoder_v0p0p1_0.x5.x17.C 16to4_PriorityEncoder_v0p0p1_0.x5.x17.D 0.253f
C567 frontAnalog_v0p0p1_5.x65.A frontAnalog_v0p0p1_5.x65.X 0.0236f
C568 w_55000_n57550# a_55268_n57936# 0.12f
C569 frontAnalog_v0p0p1_10.IB a_53630_n25596# 0.473f
C570 frontAnalog_v0p0p1_4.x63.A CLK 1.81f
C571 frontAnalog_v0p0p1_1.x63.A VIN 0.187f
C572 frontAnalog_v0p0p1_7.x65.A frontAnalog_v0p0p1_7.x65.X 0.0236f
C573 frontAnalog_v0p0p1_10.RSfetsym_0.QN frontAnalog_v0p0p1_10.RSfetsym_0.x2.Y 0.018f
C574 a_78159_n47589# VDD 0.152f
C575 a_59577_n73683# VDD 0.0173f
C576 16to4_PriorityEncoder_v0p0p1_0.x3.x9.Y a_78159_n47589# 0.299f
C577 frontAnalog_v0p0p1_11.RSfetsym_0.QN a_59577_n62883# 0.418f
C578 a_55268_n79536# VIN 0.177f
C579 frontAnalog_v0p0p1_7.x63.X frontAnalog_v0p0p1_7.RSfetsym_0.x2.Y 0.0923f
C580 frontAnalog_v0p0p1_7.RSfetsym_0.QN a_59577_n35883# 0.418f
C581 a_53630_n14796# resistorDivider_v0p0p1_0.V14 0.28f
C582 a_57123_n52679# VDD 0.222f
C583 frontAnalog_v0p0p1_1.x63.A frontAnalog_v0p0p1_1.x63.X 0.0301f
C584 frontAnalog_v0p0p1_10.x63.X a_59577_n57483# 0.28f
C585 frontAnalog_v0p0p1_7.x63.A a_57123_n36479# 0.212f
C586 w_55000_n41350# VIN 0.737f
C587 16to4_PriorityEncoder_v0p0p1_0.x5.x22.A 16to4_PriorityEncoder_v0p0p1_0.x5.A2 0.0408f
C588 frontAnalog_v0p0p1_7.RSfetsym_0.x2.Y VDD 0.926f
C589 a_77605_n51335# 16to4_PriorityEncoder_v0p0p1_0.x3.x17.C 0.0951f
C590 frontAnalog_v0p0p1_9.x63.X CLK 0.785f
C591 16to4_PriorityEncoder_v0p0p1_0.x5.x20.B a_77605_n44527# 0.14f
C592 16to4_PriorityEncoder_v0p0p1_0.x5.A2 16to4_PriorityEncoder_v0p0p1_0.x35.A 0.0138f
C593 a_82906_n51645# 16to4_PriorityEncoder_v0p0p1_0.x3.A0 0.119f
C594 16to4_PriorityEncoder_v0p0p1_0.x1.A a_82906_n47995# 0.206f
C595 16to4_PriorityEncoder_v0p0p1_0.I13 16to4_PriorityEncoder_v0p0p1_0.x5.x9.Y 0.0107f
C596 frontAnalog_v0p0p1_10.x63.A frontAnalog_v0p0p1_10.x63.X 0.0301f
C597 w_55000_n73128# VDD 0.854f
C598 a_82906_n43855# VDD 0.181f
C599 a_57123_n18759# VDD 0.224f
C600 frontAnalog_v0p0p1_15.x63.X m3_58396_n85350# 0.139f
C601 frontAnalog_v0p0p1_2.x63.A frontAnalog_v0p0p1_10.IB 0.0784f
C602 frontAnalog_v0p0p1_1.x63.A a_55268_n41736# 1.24f
C603 a_77605_n52819# 16to4_PriorityEncoder_v0p0p1_0.x3.x22.C 0.0873f
C604 a_55268_n57936# VIN 0.177f
C605 frontAnalog_v0p0p1_10.IB a_55268_n14736# 0.0848f
C606 frontAnalog_v0p0p1_8.x65.X frontAnalog_v0p0p1_8.RSfetsym_0.x2.Y 0.526f
C607 frontAnalog_v0p0p1_8.RSfetsym_0.QN frontAnalog_v0p0p1_8.x63.X 0.378f
C608 frontAnalog_v0p0p1_5.x63.A VIN 0.188f
C609 a_53630_n25596# resistorDivider_v0p0p1_0.V12 0.28f
C610 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_0.x65.A 0.0352f
C611 frontAnalog_v0p0p1_9.RSfetsym_0.x2.Y VDD 0.926f
C612 m3_58396_n4350# VDD 1.3f
C613 16to4_PriorityEncoder_v0p0p1_0.x3.x17.C 16to4_PriorityEncoder_v0p0p1_0.x3.x17.D 0.253f
C614 w_55000_n41350# a_55268_n41736# 0.12f
C615 a_55268_n3936# VDD 0.565f
C616 w_55000_n25150# CLK 0.535f
C617 w_55000_n67728# frontAnalog_v0p0p1_13.x65.A 0.658f
C618 w_55000_n83928# VIN 0.866f
C619 a_53630_n3996# a_55268_n3936# 0.015f
C620 w_55000_n68350# frontAnalog_v0p0p1_13.x63.A 0.659f
C621 frontAnalog_v0p0p1_7.x65.A VDD 3.45f
C622 a_78525_n45515# 16to4_PriorityEncoder_v0p0p1_0.x2.A 0.148f
C623 16to4_PriorityEncoder_v0p0p1_0.x5.A2 16to4_PriorityEncoder_v0p0p1_0.x34.A 0.0422f
C624 frontAnalog_v0p0p1_9.x65.A VIN 0.655f
C625 a_78349_n43045# 16to4_PriorityEncoder_v0p0p1_0.x1.A 0.151f
C626 w_55000_n13728# frontAnalog_v0p0p1_10.IB 0.0216f
C627 a_59577_n52083# VDD 0.0173f
C628 w_55000_n83928# a_55268_n84936# 0.149f
C629 w_55000_n84550# a_53630_n84996# 0.394f
C630 frontAnalog_v0p0p1_1.x63.A a_57123_n41879# 0.212f
C631 resistorDivider_v0p0p1_0.V2 a_53630_n79596# 0.28f
C632 a_55268_n20136# resistorDivider_v0p0p1_0.V13 0.215f
C633 16to4_PriorityEncoder_v0p0p1_0.x5.x19.C 16to4_PriorityEncoder_v0p0p1_0.x5.x20.B 0.996f
C634 frontAnalog_v0p0p1_9.x63.A frontAnalog_v0p0p1_9.x63.X 0.0301f
C635 w_55000_n24528# frontAnalog_v0p0p1_5.x63.A 0.0792f
C636 resistorDivider_v0p0p1_0.V16 resistorDivider_v0p0p1_0.V15 4.68f
C637 resistorDivider_v0p0p1_0.V15 CLK 6.32f
C638 a_59578_n19170# VDD 0.0213f
C639 frontAnalog_v0p0p1_6.x65.A CLK 2.62f
C640 frontAnalog_v0p0p1_13.x63.A VDD 3.67f
C641 resistorDivider_v0p0p1_0.V2 CLK 6.06f
C642 16to4_PriorityEncoder_v0p0p1_0.x5.x17.D 16to4_PriorityEncoder_v0p0p1_0.x5.x21.B 0.0218f
C643 w_55000_n8950# a_53630_n9396# 0.394f
C644 w_55000_n8328# a_55268_n9336# 0.149f
C645 frontAnalog_v0p0p1_9.RSfetsym_0.QN frontAnalog_v0p0p1_9.RSfetsym_0.x1.Y 0.17f
C646 w_55000_n8328# VIN 0.866f
C647 resistorDivider_v0p0p1_0.V7 resistorDivider_v0p0p1_0.V6 4.01f
C648 resistorDivider_v0p0p1_0.V13 VDD 4.13f
C649 16to4_PriorityEncoder_v0p0p1_0.x5.x22.D 16to4_PriorityEncoder_v0p0p1_0.x2.A 0.0148f
C650 m3_58396_n85350# VDD 1.3f
C651 16to4_PriorityEncoder_v0p0p1_0.I13 16to4_PriorityEncoder_v0p0p1_0.x5.x20.B 0.551f
C652 a_53630_n20196# CLK 0.0136f
C653 frontAnalog_v0p0p1_8.x65.A VDD 3.45f
C654 w_55000_n67728# CLK 0.571f
C655 frontAnalog_v0p0p1_9.x65.X a_59578_n51570# 0.436f
C656 frontAnalog_v0p0p1_7.x63.A frontAnalog_v0p0p1_7.x65.A 3.16f
C657 frontAnalog_v0p0p1_8.RSfetsym_0.QN a_59577_n46683# 0.418f
C658 16to4_PriorityEncoder_v0p0p1_0.x2.A 16to4_PriorityEncoder_v0p0p1_0.x21.A 0.0121f
C659 resistorDivider_v0p0p1_0.V10 CLK 6.39f
C660 w_55000_n35950# VDD 0.829f
C661 frontAnalog_v0p0p1_12.x65.X CLK 0.0402f
C662 resistorDivider_v0p0p1_0.V8 CLK 5.47f
C663 16to4_PriorityEncoder_v0p0p1_0.I12 a_77605_n40069# 0.208f
C664 frontAnalog_v0p0p1_14.x65.A VDD 3.45f
C665 frontAnalog_v0p0p1_4.RSfetsym_0.x1.Y VDD 0.733f
C666 w_55000_n52150# frontAnalog_v0p0p1_10.IB 0.0217f
C667 a_78065_n49349# VDD 0.156f
C668 frontAnalog_v0p0p1_10.IB a_53630_n47196# 0.473f
C669 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_10.x63.A 0.0926f
C670 a_77605_n39305# 16to4_PriorityEncoder_v0p0p1_0.x5.x4.C 0.0313f
C671 a_77605_n53805# 16to4_PriorityEncoder_v0p0p1_0.x3.x22.D 0.0895f
C672 16to4_PriorityEncoder_v0p0p1_0.I11 16to4_PriorityEncoder_v0p0p1_0.x5.x17.D 0.0148f
C673 w_55000_n79150# resistorDivider_v0p0p1_0.V2 0.751f
C674 16to4_PriorityEncoder_v0p0p1_0.x5.x18.C 16to4_PriorityEncoder_v0p0p1_0.x5.x20.B 0.491f
C675 frontAnalog_v0p0p1_4.RSfetsym_0.QN VDD 2.56f
C676 w_55000_n35328# frontAnalog_v0p0p1_7.x65.A 0.658f
C677 frontAnalog_v0p0p1_10.IB a_55268_n30936# 0.0848f
C678 16to4_PriorityEncoder_v0p0p1_0.x3.x22.D 16to4_PriorityEncoder_v0p0p1_0.x3.x22.B 0.122f
C679 frontAnalog_v0p0p1_12.x63.X CLK 0.785f
C680 w_55000_n46750# VIN 0.737f
C681 a_57123_n18759# frontAnalog_v0p0p1_4.x65.X 0.119f
C682 a_57123_n20279# VDD 0.222f
C683 16to4_PriorityEncoder_v0p0p1_0.x5.x19.C 16to4_PriorityEncoder_v0p0p1_0.x5.x16.C 1.95f
C684 a_82906_n43855# 16to4_PriorityEncoder_v0p0p1_0.x34.A 0.12f
C685 w_55000_n73128# w_55000_n73750# 0.327f
C686 w_55000_n35950# frontAnalog_v0p0p1_7.x63.A 0.659f
C687 16to4_PriorityEncoder_v0p0p1_0.x2.A VDD 1.89f
C688 a_53630_n25596# VIN 0.265f
C689 resistorDivider_v0p0p1_0.V5 frontAnalog_v0p0p1_11.x63.A 0.587f
C690 16to4_PriorityEncoder_v0p0p1_0.x3.EI 16to4_PriorityEncoder_v0p0p1_0.x2.A 0.645f
C691 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_12.x63.A 0.0926f
C692 frontAnalog_v0p0p1_1.x65.A a_57123_n40359# 0.214f
C693 16to4_PriorityEncoder_v0p0p1_0.I15 16to4_PriorityEncoder_v0p0p1_0.I14 5.72f
C694 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD 11.4f
C695 w_55000_n78528# VDD 0.854f
C696 16to4_PriorityEncoder_v0p0p1_0.x2.A 16to4_PriorityEncoder_v0p0p1_0.x2.X 0.0402f
C697 w_55000_n14350# resistorDivider_v0p0p1_0.V14 0.751f
C698 16to4_PriorityEncoder_v0p0p1_0.I14 16to4_PriorityEncoder_v0p0p1_0.x5.x4.C 0.0177f
C699 16to4_PriorityEncoder_v0p0p1_0.I13 16to4_PriorityEncoder_v0p0p1_0.x5.x16.C 0.415f
C700 frontAnalog_v0p0p1_10.IB resistorDivider_v0p0p1_0.V3 3.7f
C701 resistorDivider_v0p0p1_0.V7 VDD 4.76f
C702 resistorDivider_v0p0p1_0.V5 resistorDivider_v0p0p1_0.V4 5.09f
C703 w_55000_n67728# a_55268_n68736# 0.149f
C704 w_55000_n68350# a_53630_n68796# 0.394f
C705 16to4_PriorityEncoder_v0p0p1_0.x5.x19.C a_77605_n44527# 0.157f
C706 frontAnalog_v0p0p1_8.x63.A frontAnalog_v0p0p1_8.x65.A 3.16f
C707 w_55000_n35328# w_55000_n35950# 0.327f
C708 a_77605_n39305# 16to4_PriorityEncoder_v0p0p1_0.x5.x4.B 0.0991f
C709 frontAnalog_v0p0p1_3.x65.A VDD 3.45f
C710 m3_58396_n15150# VDD 1.3f
C711 resistorDivider_v0p0p1_0.V3 frontAnalog_v0p0p1_12.x63.A 0.587f
C712 16to4_PriorityEncoder_v0p0p1_0.x3.x22.C 16to4_PriorityEncoder_v0p0p1_0.x3.x22.D 0.145f
C713 w_55000_n40728# resistorDivider_v0p0p1_0.V9 0.798f
C714 frontAnalog_v0p0p1_2.x65.X VDD 3.55f
C715 w_55000_n30550# CLK 0.535f
C716 frontAnalog_v0p0p1_4.RSfetsym_0.x2.Y VDD 0.926f
C717 w_55000_n24528# a_53630_n25596# 0.359f
C718 16to4_PriorityEncoder_v0p0p1_0.x3.x17.A VDD 1.34f
C719 a_53630_n68796# VDD 0.134f
C720 a_77637_n49127# VDD 0.218f
C721 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_15.x65.A 0.0352f
C722 resistorDivider_v0p0p1_0.V9 CLK 6.38f
C723 frontAnalog_v0p0p1_10.IB resistorDivider_v0p0p1_0.V12 3.69f
C724 a_53630_n30996# resistorDivider_v0p0p1_0.V11 0.28f
C725 w_55000_n2928# VDD 0.854f
C726 frontAnalog_v0p0p1_2.x63.A VIN 0.187f
C727 16to4_PriorityEncoder_v0p0p1_0.x3.EI 16to4_PriorityEncoder_v0p0p1_0.x3.x17.A 0.02f
C728 frontAnalog_v0p0p1_4.x65.X a_59578_n19170# 0.436f
C729 resistorDivider_v0p0p1_0.V6 a_55268_n57936# 0.215f
C730 a_55268_n14736# VIN 0.177f
C731 16to4_PriorityEncoder_v0p0p1_0.x3.EI a_77637_n49127# 0.0829f
C732 frontAnalog_v0p0p1_0.x65.A a_55268_n9336# 0.461f
C733 w_55000_n25150# frontAnalog_v0p0p1_5.x65.A 0.0988f
C734 w_55000_n2928# a_53630_n3996# 0.359f
C735 frontAnalog_v0p0p1_8.RSfetsym_0.x1.Y frontAnalog_v0p0p1_8.x63.X 0.883f
C736 frontAnalog_v0p0p1_0.x65.A VIN 0.655f
C737 16to4_PriorityEncoder_v0p0p1_0.x3.x21.B VDD 0.721f
C738 w_55000_n19128# frontAnalog_v0p0p1_10.IB 0.0216f
C739 16to4_PriorityEncoder_v0p0p1_0.x5.x22.A 16to4_PriorityEncoder_v0p0p1_0.x2.A 0.132f
C740 frontAnalog_v0p0p1_14.x63.A frontAnalog_v0p0p1_14.x65.A 3.16f
C741 16to4_PriorityEncoder_v0p0p1_0.x5.x20.B a_77605_n45765# 0.0838f
C742 16to4_PriorityEncoder_v0p0p1_0.x3.EI 16to4_PriorityEncoder_v0p0p1_0.x3.x21.B 0.187f
C743 frontAnalog_v0p0p1_3.RSfetsym_0.QN a_59578_n13770# 0.255f
C744 frontAnalog_v0p0p1_8.x63.X VDD 3.16f
C745 16to4_PriorityEncoder_v0p0p1_0.x43.A VDD 1.46f
C746 16to4_PriorityEncoder_v0p0p1_0.x5.x17.D a_77605_n43545# 0.102f
C747 frontAnalog_v0p0p1_10.x63.X m3_58396_n58350# 0.139f
C748 16to4_PriorityEncoder_v0p0p1_0.x3.x17.D a_77605_n51585# 0.102f
C749 w_55000_n83928# resistorDivider_v0p0p1_0.V1 0.798f
C750 w_55000_n56928# frontAnalog_v0p0p1_10.x65.A 0.658f
C751 a_53630_n52596# VDD 0.134f
C752 w_55000_n13728# VIN 0.866f
C753 16to4_PriorityEncoder_v0p0p1_0.I15 VDD 9.55f
C754 16to4_PriorityEncoder_v0p0p1_0.x5.x20.B a_77605_n44779# 0.148f
C755 16to4_PriorityEncoder_v0p0p1_0.x5.x18.C a_77605_n44527# 0.117f
C756 a_77605_n47345# 16to4_PriorityEncoder_v0p0p1_0.x3.x4.C 0.0313f
C757 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_11.x65.A 0.0352f
C758 frontAnalog_v0p0p1_1.x63.A VDD 3.67f
C759 16to4_PriorityEncoder_v0p0p1_0.x5.x4.C VDD 0.367f
C760 16to4_PriorityEncoder_v0p0p1_0.I12 a_59578_n19170# 0.42f
C761 16to4_PriorityEncoder_v0p0p1_0.x5.x9.Y a_77605_n39305# 0.0112f
C762 w_55000_n57550# frontAnalog_v0p0p1_10.x63.A 0.659f
C763 frontAnalog_v0p0p1_4.x65.X frontAnalog_v0p0p1_4.RSfetsym_0.x1.Y 0.182f
C764 w_55000_n73128# CLK 0.571f
C765 a_55268_n79536# VDD 0.565f
C766 w_55000_n46128# resistorDivider_v0p0p1_0.V8 0.798f
C767 16to4_PriorityEncoder_v0p0p1_0.x2.A 16to4_PriorityEncoder_v0p0p1_0.x3.A0 0.398f
C768 frontAnalog_v0p0p1_3.x65.X frontAnalog_v0p0p1_3.x63.X 0.136f
C769 frontAnalog_v0p0p1_13.x63.A frontAnalog_v0p0p1_13.x65.A 3.16f
C770 frontAnalog_v0p0p1_3.x65.X 16to4_PriorityEncoder_v0p0p1_0.I13 0.446f
C771 w_55000_n41350# VDD 0.829f
C772 frontAnalog_v0p0p1_9.x65.X frontAnalog_v0p0p1_9.x63.X 0.136f
C773 w_55000_n78528# frontAnalog_v0p0p1_14.x63.A 0.0792f
C774 frontAnalog_v0p0p1_2.x63.X VDD 3.16f
C775 frontAnalog_v0p0p1_4.x65.X frontAnalog_v0p0p1_4.RSfetsym_0.QN 2.28f
C776 w_55000_n57550# frontAnalog_v0p0p1_10.IB 0.0217f
C777 frontAnalog_v0p0p1_3.RSfetsym_0.QN frontAnalog_v0p0p1_3.RSfetsym_0.x1.Y 0.17f
C778 resistorDivider_v0p0p1_0.V5 a_53630_n63396# 0.28f
C779 a_55268_n3936# resistorDivider_v0p0p1_0.V16 0.214f
C780 16to4_PriorityEncoder_v0p0p1_0.I13 16to4_PriorityEncoder_v0p0p1_0.x5.x19.C 0.407f
C781 a_55268_n3936# CLK 0.236f
C782 a_78525_n53555# 16to4_PriorityEncoder_v0p0p1_0.x3.x22.D 0.0765f
C783 16to4_PriorityEncoder_v0p0p1_0.x3.x22.C 16to4_PriorityEncoder_v0p0p1_0.x3.x22.B 0.131f
C784 frontAnalog_v0p0p1_10.IB a_53630_n74196# 0.473f
C785 16to4_PriorityEncoder_v0p0p1_0.x42.A VDD 0.536f
C786 frontAnalog_v0p0p1_5.RSfetsym_0.QN a_59578_n24570# 0.255f
C787 16to4_PriorityEncoder_v0p0p1_0.x3.x22.A VDD 3.23f
C788 16to4_PriorityEncoder_v0p0p1_0.I12 frontAnalog_v0p0p1_4.RSfetsym_0.x1.Y 0.0436f
C789 16to4_PriorityEncoder_v0p0p1_0.x3.x4.C VDD 0.371f
C790 a_55268_n57936# VDD 0.565f
C791 frontAnalog_v0p0p1_7.x65.A CLK 2.61f
C792 w_55000_n52150# VIN 0.737f
C793 16to4_PriorityEncoder_v0p0p1_0.x3.EI 16to4_PriorityEncoder_v0p0p1_0.x3.x22.A 0.0483f
C794 frontAnalog_v0p0p1_9.x63.A a_57123_n52679# 0.212f
C795 frontAnalog_v0p0p1_0.x63.A resistorDivider_v0p0p1_0.V15 0.587f
C796 a_53630_n47196# VIN 0.265f
C797 frontAnalog_v0p0p1_5.x63.A VDD 3.67f
C798 16to4_PriorityEncoder_v0p0p1_0.I15 16to4_PriorityEncoder_v0p0p1_0.x5.x22.A 0.0853f
C799 frontAnalog_v0p0p1_10.x63.A VIN 0.187f
C800 16to4_PriorityEncoder_v0p0p1_0.I13 frontAnalog_v0p0p1_3.x63.X 1.85f
C801 a_59577_n46683# VDD 0.0173f
C802 frontAnalog_v0p0p1_5.x65.X 16to4_PriorityEncoder_v0p0p1_0.I11 0.446f
C803 16to4_PriorityEncoder_v0p0p1_0.x3.x9.Y 16to4_PriorityEncoder_v0p0p1_0.x3.x4.C 0.125f
C804 a_77605_n47345# 16to4_PriorityEncoder_v0p0p1_0.x3.x4.B 0.0991f
C805 16to4_PriorityEncoder_v0p0p1_0.I11 16to4_PriorityEncoder_v0p0p1_0.x5.x21.B 0.0112f
C806 16to4_PriorityEncoder_v0p0p1_0.x5.x4.B VDD 0.39f
C807 resistorDivider_v0p0p1_0.V3 a_53630_n74196# 0.28f
C808 frontAnalog_v0p0p1_8.x63.A frontAnalog_v0p0p1_8.x63.X 0.0301f
C809 frontAnalog_v0p0p1_1.x65.A resistorDivider_v0p0p1_0.V9 0.253f
C810 frontAnalog_v0p0p1_4.RSfetsym_0.x1.Y frontAnalog_v0p0p1_4.x63.X 0.883f
C811 16to4_PriorityEncoder_v0p0p1_0.x3.GS VDD 0.608f
C812 frontAnalog_v0p0p1_4.RSfetsym_0.QN 16to4_PriorityEncoder_v0p0p1_0.I12 2.02f
C813 16to4_PriorityEncoder_v0p0p1_0.x3.x20.B 16to4_PriorityEncoder_v0p0p1_0.x3.x21.B 0.151f
C814 frontAnalog_v0p0p1_13.x63.A CLK 1.81f
C815 w_55000_n8950# resistorDivider_v0p0p1_0.V15 0.751f
C816 a_55268_n30936# VIN 0.177f
C817 16to4_PriorityEncoder_v0p0p1_0.x5.x18.C 16to4_PriorityEncoder_v0p0p1_0.x5.x19.C 2.6f
C818 frontAnalog_v0p0p1_3.RSfetsym_0.x1.Y frontAnalog_v0p0p1_3.RSfetsym_0.x2.Y 0.0254f
C819 frontAnalog_v0p0p1_5.x65.X frontAnalog_v0p0p1_5.x63.X 0.136f
C820 16to4_PriorityEncoder_v0p0p1_0.x3.EI 16to4_PriorityEncoder_v0p0p1_0.x3.GS 0.123f
C821 w_55000_n83928# VDD 0.854f
C822 w_55000_n62328# resistorDivider_v0p0p1_0.V5 0.798f
C823 frontAnalog_v0p0p1_10.IB VIN 32.9f
C824 frontAnalog_v0p0p1_10.IB a_55268_n9336# 0.0848f
C825 resistorDivider_v0p0p1_0.V13 CLK 6.01f
C826 frontAnalog_v0p0p1_4.RSfetsym_0.QN frontAnalog_v0p0p1_4.x63.X 0.378f
C827 frontAnalog_v0p0p1_4.x65.X frontAnalog_v0p0p1_4.RSfetsym_0.x2.Y 0.526f
C828 frontAnalog_v0p0p1_9.x65.A VDD 3.45f
C829 frontAnalog_v0p0p1_5.RSfetsym_0.QN frontAnalog_v0p0p1_5.RSfetsym_0.x1.Y 0.17f
C830 frontAnalog_v0p0p1_8.x65.A CLK 2.61f
C831 16to4_PriorityEncoder_v0p0p1_0.x5.EO VDD 1.06f
C832 frontAnalog_v0p0p1_10.IB a_55268_n84936# 0.0848f
C833 m3_58396_n25950# VDD 1.3f
C834 frontAnalog_v0p0p1_12.x63.A VIN 0.187f
C835 16to4_PriorityEncoder_v0p0p1_0.I13 16to4_PriorityEncoder_v0p0p1_0.x5.x18.C 0.3f
C836 frontAnalog_v0p0p1_4.x63.X a_57123_n20279# 0.121f
C837 a_59577_n3483# VDD 0.0173f
C838 16to4_PriorityEncoder_v0p0p1_0.x5.EO 16to4_PriorityEncoder_v0p0p1_0.x3.EI 0.644f
C839 w_55000_n35950# CLK 0.535f
C840 16to4_PriorityEncoder_v0p0p1_0.x3.x14.A a_78065_n49349# 0.197f
C841 w_55000_n25150# a_55268_n25536# 0.12f
C842 frontAnalog_v0p0p1_3.RSfetsym_0.QN frontAnalog_v0p0p1_3.RSfetsym_0.x2.Y 0.018f
C843 resistorDivider_v0p0p1_0.V3 VIN 2.63f
C844 a_57123_n67359# VDD 0.224f
C845 frontAnalog_v0p0p1_14.x63.A a_55268_n79536# 1.24f
C846 16to4_PriorityEncoder_v0p0p1_0.x3.x14.B VDD 0.507f
C847 frontAnalog_v0p0p1_14.x65.A CLK 2.62f
C848 a_57123_n2559# frontAnalog_v0p0p1_2.x65.X 0.119f
C849 w_55000_n8328# VDD 0.854f
C850 frontAnalog_v0p0p1_3.x63.A frontAnalog_v0p0p1_3.x65.A 3.16f
C851 frontAnalog_v0p0p1_10.IB a_55268_n36336# 0.0848f
C852 16to4_PriorityEncoder_v0p0p1_0.x5.x22.C 16to4_PriorityEncoder_v0p0p1_0.x2.A 0.0122f
C853 16to4_PriorityEncoder_v0p0p1_0.x3.x4.B VDD 0.393f
C854 frontAnalog_v0p0p1_0.x63.A a_57123_n9479# 0.212f
C855 frontAnalog_v0p0p1_0.x65.A frontAnalog_v0p0p1_0.x65.X 0.0236f
C856 16to4_PriorityEncoder_v0p0p1_0.I11 frontAnalog_v0p0p1_5.x63.X 1.93f
C857 w_55000_n3550# a_55268_n3936# 0.12f
C858 16to4_PriorityEncoder_v0p0p1_0.x5.GS VDD 0.771f
C859 w_55000_n24528# frontAnalog_v0p0p1_10.IB 0.0216f
C860 16to4_PriorityEncoder_v0p0p1_0.x3.x9.Y 16to4_PriorityEncoder_v0p0p1_0.x3.x4.B 0.118f
C861 a_78649_n39527# 16to4_PriorityEncoder_v0p0p1_0.x5.EO 0.135f
C862 16to4_PriorityEncoder_v0p0p1_0.x5.x9.Y VDD 1.92f
C863 a_78525_n53555# 16to4_PriorityEncoder_v0p0p1_0.x3.x22.B 0.202f
C864 16to4_PriorityEncoder_v0p0p1_0.I12 frontAnalog_v0p0p1_4.RSfetsym_0.x2.Y 0.196f
C865 frontAnalog_v0p0p1_10.IB a_55268_n41736# 0.0848f
C866 frontAnalog_v0p0p1_3.x63.X a_59577_n14283# 0.28f
C867 16to4_PriorityEncoder_v0p0p1_0.I13 a_59577_n14283# 0.29f
C868 frontAnalog_v0p0p1_10.IB a_55268_n63336# 0.0848f
C869 frontAnalog_v0p0p1_15.x65.A VIN 0.655f
C870 a_59578_n67770# VDD 0.0213f
C871 resistorDivider_v0p0p1_0.V12 VIN 2.55f
C872 16to4_PriorityEncoder_v0p0p1_0.x2.A 16to4_PriorityEncoder_v0p0p1_0.x3.A1 1.21f
C873 w_55000_n62328# frontAnalog_v0p0p1_11.x63.A 0.0792f
C874 w_55000_n78528# a_53630_n79596# 0.359f
C875 frontAnalog_v0p0p1_4.x63.X frontAnalog_v0p0p1_4.RSfetsym_0.x2.Y 0.0923f
C876 16to4_PriorityEncoder_v0p0p1_0.x3.EO VDD 0.761f
C877 16to4_PriorityEncoder_v0p0p1_0.I14 16to4_PriorityEncoder_v0p0p1_0.x5.x20.B 0.464f
C878 16to4_PriorityEncoder_v0p0p1_0.x3.x20.B 16to4_PriorityEncoder_v0p0p1_0.x3.x22.A 0.0292f
C879 a_57123_n51159# VDD 0.224f
C880 w_55000_n19128# VIN 0.868f
C881 frontAnalog_v0p0p1_15.x65.A a_55268_n84936# 0.461f
C882 frontAnalog_v0p0p1_5.RSfetsym_0.x1.Y frontAnalog_v0p0p1_5.RSfetsym_0.x2.Y 0.0254f
C883 frontAnalog_v0p0p1_13.x63.A a_55268_n68736# 1.24f
C884 16to4_PriorityEncoder_v0p0p1_0.x3.EI 16to4_PriorityEncoder_v0p0p1_0.x3.EO 0.187f
C885 16to4_PriorityEncoder_v0p0p1_0.x3.x9.Y 16to4_PriorityEncoder_v0p0p1_0.x3.EO 0.0491f
C886 16to4_PriorityEncoder_v0p0p1_0.x3.x22.A 16to4_PriorityEncoder_v0p0p1_0.x3.A0 0.132f
C887 16to4_PriorityEncoder_v0p0p1_0.x3.x20.B 16to4_PriorityEncoder_v0p0p1_0.x3.x4.C 0.014f
C888 a_77605_n52567# 16to4_PriorityEncoder_v0p0p1_0.x3.x21.B 0.116f
C889 a_78649_n39527# 16to4_PriorityEncoder_v0p0p1_0.x5.GS 0.136f
C890 frontAnalog_v0p0p1_4.RSfetsym_0.QN a_59577_n19683# 0.418f
C891 w_55000_n79150# frontAnalog_v0p0p1_14.x65.A 0.0988f
C892 a_82906_n47995# VDD 0.179f
C893 w_55000_n78528# CLK 0.571f
C894 frontAnalog_v0p0p1_6.x63.A a_55268_n30936# 1.24f
C895 frontAnalog_v0p0p1_14.x65.X VDD 3.55f
C896 a_78649_n47567# 16to4_PriorityEncoder_v0p0p1_0.x3.GS 0.136f
C897 frontAnalog_v0p0p1_5.RSfetsym_0.QN frontAnalog_v0p0p1_5.RSfetsym_0.x2.Y 0.018f
C898 resistorDivider_v0p0p1_0.V7 CLK 5.72f
C899 w_55000_n46750# VDD 0.829f
C900 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_6.x63.A 0.0926f
C901 16to4_PriorityEncoder_v0p0p1_0.I15 16to4_PriorityEncoder_v0p0p1_0.I12 0.786f
C902 16to4_PriorityEncoder_v0p0p1_0.x3.x22.C a_78525_n53555# 0.193f
C903 w_55000_n24528# resistorDivider_v0p0p1_0.V12 0.798f
C904 frontAnalog_v0p0p1_11.x65.A VIN 0.655f
C905 16to4_PriorityEncoder_v0p0p1_0.I12 16to4_PriorityEncoder_v0p0p1_0.x5.x4.C 0.0262f
C906 frontAnalog_v0p0p1_3.x65.A CLK 2.61f
C907 16to4_PriorityEncoder_v0p0p1_0.x3.x14.A 16to4_PriorityEncoder_v0p0p1_0.x3.x17.A 0.105f
C908 w_55000_n62950# frontAnalog_v0p0p1_10.IB 0.0217f
C909 a_53630_n25596# VDD 0.134f
C910 a_77637_n50057# VDD 0.234f
C911 16to4_PriorityEncoder_v0p0p1_0.x5.x19.C a_77605_n44779# 0.102f
C912 16to4_PriorityEncoder_v0p0p1_0.x3.A1 16to4_PriorityEncoder_v0p0p1_0.x3.x17.A 0.115f
C913 frontAnalog_v0p0p1_13.RSfetsym_0.x1.Y VDD 0.733f
C914 16to4_PriorityEncoder_v0p0p1_0.I13 a_77605_n45765# 0.193f
C915 frontAnalog_v0p0p1_2.x65.X a_59578_n2970# 0.436f
C916 16to4_PriorityEncoder_v0p0p1_0.x5.x17.A a_78349_n43045# 0.213f
C917 frontAnalog_v0p0p1_2.x65.X CLK 0.0302f
C918 frontAnalog_v0p0p1_12.x65.A a_55268_n74136# 0.461f
C919 16to4_PriorityEncoder_v0p0p1_0.x3.EI a_77637_n50057# 0.0878f
C920 a_53630_n68796# CLK 0.0136f
C921 frontAnalog_v0p0p1_14.x63.X VDD 3.16f
C922 16to4_PriorityEncoder_v0p0p1_0.I11 frontAnalog_v0p0p1_6.RSfetsym_0.QN 0.0512f
C923 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_4.x65.A 0.0352f
C924 w_55000_n2928# resistorDivider_v0p0p1_0.V16 0.798f
C925 w_55000_n2928# CLK 0.57f
C926 16to4_PriorityEncoder_v0p0p1_0.I11 a_59577_n25083# 0.29f
C927 w_55000_n57550# VIN 0.737f
C928 16to4_PriorityEncoder_v0p0p1_0.I11 a_77605_n43545# 0.162f
C929 VDD OUT3 7.1f
C930 frontAnalog_v0p0p1_10.x65.X VDD 3.55f
C931 w_55000_n78528# w_55000_n79150# 0.327f
C932 frontAnalog_v0p0p1_5.x63.X a_59577_n25083# 0.28f
C933 a_57123_n68879# VDD 0.222f
C934 frontAnalog_v0p0p1_6.RSfetsym_0.QN a_59578_n29970# 0.255f
C935 a_78349_n43045# VDD 0.164f
C936 a_53630_n74196# VIN 0.265f
C937 16to4_PriorityEncoder_v0p0p1_0.x5.x20.B VDD 3.27f
C938 a_77605_n51335# VDD 0.435f
C939 frontAnalog_v0p0p1_8.x63.X CLK 0.785f
C940 16to4_PriorityEncoder_v0p0p1_0.I14 16to4_PriorityEncoder_v0p0p1_0.x5.x16.C 0.491f
C941 frontAnalog_v0p0p1_13.RSfetsym_0.QN VDD 2.56f
C942 frontAnalog_v0p0p1_2.x63.A VDD 3.67f
C943 16to4_PriorityEncoder_v0p0p1_0.x3.EI a_77605_n51335# 0.122f
C944 a_53630_n79596# a_55268_n79536# 0.015f
C945 16to4_PriorityEncoder_v0p0p1_0.I15 a_59578_n2970# 0.42f
C946 w_55000_n40728# frontAnalog_v0p0p1_1.x63.A 0.0792f
C947 a_53630_n52596# CLK 0.0136f
C948 frontAnalog_v0p0p1_2.x65.X frontAnalog_v0p0p1_2.RSfetsym_0.QN 2.28f
C949 a_55268_n14736# VDD 0.565f
C950 frontAnalog_v0p0p1_11.x65.A a_55268_n63336# 0.461f
C951 frontAnalog_v0p0p1_2.x65.X frontAnalog_v0p0p1_2.RSfetsym_0.x1.Y 0.182f
C952 16to4_PriorityEncoder_v0p0p1_0.I15 CLK 0.01f
C953 frontAnalog_v0p0p1_10.x63.X VDD 3.16f
C954 w_55000_n46128# frontAnalog_v0p0p1_8.x65.A 0.658f
C955 frontAnalog_v0p0p1_0.x65.A VDD 3.45f
C956 frontAnalog_v0p0p1_7.x63.X m3_58396_n36750# 0.139f
C957 16to4_PriorityEncoder_v0p0p1_0.x5.x21.B a_78097_n45737# 0.186f
C958 frontAnalog_v0p0p1_1.x63.A CLK 1.81f
C959 frontAnalog_v0p0p1_1.RSfetsym_0.x1.Y frontAnalog_v0p0p1_1.x63.X 0.883f
C960 a_78649_n47567# 16to4_PriorityEncoder_v0p0p1_0.x3.EO 0.135f
C961 resistorDivider_v0p0p1_0.V6 frontAnalog_v0p0p1_10.x63.A 0.587f
C962 frontAnalog_v0p0p1_14.x65.A a_57123_n78159# 0.214f
C963 resistorDivider_v0p0p1_0.V7 frontAnalog_v0p0p1_9.x63.A 0.587f
C964 m3_58396_n36750# VDD 1.3f
C965 a_55268_n79536# CLK 0.236f
C966 w_55000_n40728# w_55000_n41350# 0.327f
C967 frontAnalog_v0p0p1_6.x65.X frontAnalog_v0p0p1_6.x63.X 0.136f
C968 w_55000_n46750# frontAnalog_v0p0p1_8.x63.A 0.659f
C969 frontAnalog_v0p0p1_14.x63.X m3_58396_n79950# 0.139f
C970 16to4_PriorityEncoder_v0p0p1_0.x3.x19.C 16to4_PriorityEncoder_v0p0p1_0.x3.x21.B 0.0127f
C971 w_55000_n41350# CLK 0.535f
C972 frontAnalog_v0p0p1_8.x63.X a_57123_n47279# 0.121f
C973 a_77637_n40777# 16to4_PriorityEncoder_v0p0p1_0.x5.x14.A 0.135f
C974 a_55268_n9336# VIN 0.177f
C975 resistorDivider_v0p0p1_0.V16 VFS 4.16f
C976 frontAnalog_v0p0p1_13.RSfetsym_0.x2.Y VDD 0.926f
C977 w_55000_n19128# frontAnalog_v0p0p1_4.x65.A 0.658f
C978 w_55000_n62328# a_53630_n63396# 0.359f
C979 frontAnalog_v0p0p1_10.IB resistorDivider_v0p0p1_0.V6 3.7f
C980 frontAnalog_v0p0p1_2.x63.X CLK 0.785f
C981 w_55000_n30550# a_53630_n30996# 0.394f
C982 frontAnalog_v0p0p1_6.RSfetsym_0.QN frontAnalog_v0p0p1_6.RSfetsym_0.x1.Y 0.17f
C983 w_55000_n29928# a_55268_n30936# 0.149f
C984 frontAnalog_v0p0p1_10.IB resistorDivider_v0p0p1_0.V1 0.0595f
C985 resistorDivider_v0p0p1_0.V15 resistorDivider_v0p0p1_0.V14 5.48f
C986 w_55000_n13728# VDD 0.854f
C987 16to4_PriorityEncoder_v0p0p1_0.x3.x17.D VDD 0.505f
C988 a_59577_n79083# VDD 0.0173f
C989 frontAnalog_v0p0p1_15.x63.A a_57123_n85079# 0.212f
C990 frontAnalog_v0p0p1_9.RSfetsym_0.QN VDD 2.56f
C991 16to4_PriorityEncoder_v0p0p1_0.I15 a_77639_n42341# 0.192f
C992 a_53630_n68796# a_55268_n68736# 0.015f
C993 a_55268_n84936# VIN 0.177f
C994 w_55000_n29928# frontAnalog_v0p0p1_10.IB 0.0216f
C995 16to4_PriorityEncoder_v0p0p1_0.x3.x14.A 16to4_PriorityEncoder_v0p0p1_0.x3.x22.A 0.0179f
C996 w_55000_n19750# frontAnalog_v0p0p1_4.x63.A 0.659f
C997 16to4_PriorityEncoder_v0p0p1_0.x3.EI 16to4_PriorityEncoder_v0p0p1_0.x3.x17.D 0.076f
C998 16to4_PriorityEncoder_v0p0p1_0.x3.A1 16to4_PriorityEncoder_v0p0p1_0.x3.x22.A 0.519f
C999 frontAnalog_v0p0p1_9.x63.X m3_58396_n52950# 0.139f
C1000 frontAnalog_v0p0p1_2.RSfetsym_0.QN 16to4_PriorityEncoder_v0p0p1_0.I15 2.02f
C1001 16to4_PriorityEncoder_v0p0p1_0.I15 frontAnalog_v0p0p1_2.RSfetsym_0.x1.Y 0.0432f
C1002 w_55000_n62950# frontAnalog_v0p0p1_11.x65.A 0.0988f
C1003 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2 8.68f
C1004 16to4_PriorityEncoder_v0p0p1_0.x5.x22.A a_78349_n43045# 0.17f
C1005 w_55000_n2928# w_55000_n3550# 0.327f
C1006 16to4_PriorityEncoder_v0p0p1_0.x5.x20.B 16to4_PriorityEncoder_v0p0p1_0.x5.x22.A 0.0292f
C1007 resistorDivider_v0p0p1_0.V7 a_55268_n52536# 0.215f
C1008 frontAnalog_v0p0p1_13.x65.A a_57123_n67359# 0.214f
C1009 frontAnalog_v0p0p1_14.x63.A frontAnalog_v0p0p1_14.x63.X 0.0301f
C1010 a_55268_n57936# CLK 0.236f
C1011 a_55268_n36336# VIN 0.177f
C1012 frontAnalog_v0p0p1_5.x63.A CLK 1.81f
C1013 w_55000_n79150# a_55268_n79536# 0.12f
C1014 16to4_PriorityEncoder_v0p0p1_0.x5.x16.C VDD 2.83f
C1015 frontAnalog_v0p0p1_9.x65.X frontAnalog_v0p0p1_9.RSfetsym_0.x2.Y 0.526f
C1016 frontAnalog_v0p0p1_6.x65.A a_57123_n29559# 0.214f
C1017 frontAnalog_v0p0p1_15.x65.A frontAnalog_v0p0p1_15.x65.X 0.0236f
C1018 w_55000_n24528# VIN 0.866f
C1019 16to4_PriorityEncoder_v0p0p1_0.x5.A2 16to4_PriorityEncoder_v0p0p1_0.x3.A2 0.358f
C1020 frontAnalog_v0p0p1_8.x63.X frontAnalog_v0p0p1_8.RSfetsym_0.x2.Y 0.0923f
C1021 frontAnalog_v0p0p1_2.RSfetsym_0.QN frontAnalog_v0p0p1_2.x63.X 0.378f
C1022 frontAnalog_v0p0p1_2.x65.X frontAnalog_v0p0p1_2.RSfetsym_0.x2.Y 0.526f
C1023 frontAnalog_v0p0p1_2.RSfetsym_0.x1.Y frontAnalog_v0p0p1_2.x63.X 0.883f
C1024 a_55268_n41736# VIN 0.177f
C1025 a_59577_n57483# VDD 0.0173f
C1026 frontAnalog_v0p0p1_12.x63.A a_57123_n74279# 0.212f
C1027 w_55000_n83928# CLK 0.571f
C1028 16to4_PriorityEncoder_v0p0p1_0.x3.x18.C 16to4_PriorityEncoder_v0p0p1_0.x3.x21.B 0.014f
C1029 a_55268_n63336# VIN 0.177f
C1030 a_53630_n57996# a_55268_n57936# 0.015f
C1031 w_55000_n67728# resistorDivider_v0p0p1_0.V4 0.798f
C1032 resistorDivider_v0p0p1_0.V8 a_55268_n47136# 0.215f
C1033 resistorDivider_v0p0p1_0.V1 frontAnalog_v0p0p1_15.x65.A 0.252f
C1034 frontAnalog_v0p0p1_6.RSfetsym_0.x1.Y frontAnalog_v0p0p1_6.RSfetsym_0.x2.Y 0.0254f
C1035 frontAnalog_v0p0p1_9.x65.A CLK 2.61f
C1036 w_55000_n52150# VDD 0.829f
C1037 a_53630_n47196# VDD 0.134f
C1038 16to4_PriorityEncoder_v0p0p1_0.x3.x17.C VDD 0.26f
C1039 VDD OUT2 6.68f
C1040 16to4_PriorityEncoder_v0p0p1_0.I14 16to4_PriorityEncoder_v0p0p1_0.x5.x19.C 0.305f
C1041 frontAnalog_v0p0p1_10.IB a_55268_n20136# 0.0848f
C1042 frontAnalog_v0p0p1_10.x63.A VDD 3.67f
C1043 a_77605_n44527# VDD 0.439f
C1044 a_53630_n9396# resistorDivider_v0p0p1_0.V15 0.28f
C1045 frontAnalog_v0p0p1_13.x63.A frontAnalog_v0p0p1_13.x63.X 0.0301f
C1046 a_57123_n24159# VDD 0.224f
C1047 w_55000_n68350# frontAnalog_v0p0p1_10.IB 0.0217f
C1048 16to4_PriorityEncoder_v0p0p1_0.x3.x14.A 16to4_PriorityEncoder_v0p0p1_0.x3.x14.B 0.0721f
C1049 frontAnalog_v0p0p1_2.x63.X a_57123_n4079# 0.121f
C1050 16to4_PriorityEncoder_v0p0p1_0.x3.EI 16to4_PriorityEncoder_v0p0p1_0.x3.x17.C 0.0245f
C1051 frontAnalog_v0p0p1_6.RSfetsym_0.QN frontAnalog_v0p0p1_6.RSfetsym_0.x2.Y 0.018f
C1052 a_55268_n30936# VDD 0.565f
C1053 frontAnalog_v0p0p1_12.x65.A frontAnalog_v0p0p1_12.x65.X 0.0236f
C1054 frontAnalog_v0p0p1_1.x63.A frontAnalog_v0p0p1_1.x65.A 3.16f
C1055 a_53630_n52596# a_55268_n52536# 0.015f
C1056 w_55000_n8328# CLK 0.571f
C1057 frontAnalog_v0p0p1_6.x63.A VIN 0.187f
C1058 16to4_PriorityEncoder_v0p0p1_0.I15 frontAnalog_v0p0p1_2.RSfetsym_0.x2.Y 0.194f
C1059 frontAnalog_v0p0p1_10.IB VDD 47.1f
C1060 frontAnalog_v0p0p1_11.x63.A a_57123_n63479# 0.212f
C1061 16to4_PriorityEncoder_v0p0p1_0.I14 16to4_PriorityEncoder_v0p0p1_0.I13 10.5f
C1062 w_55000_n62950# VIN 0.737f
C1063 frontAnalog_v0p0p1_10.IB a_53630_n3996# 0.472f
C1064 frontAnalog_v0p0p1_1.RSfetsym_0.x1.Y frontAnalog_v0p0p1_1.RSfetsym_0.x2.Y 0.0254f
C1065 frontAnalog_v0p0p1_1.x63.X a_57123_n41879# 0.121f
C1066 w_55000_n41350# frontAnalog_v0p0p1_1.x65.A 0.0988f
C1067 frontAnalog_v0p0p1_12.x63.A VDD 3.67f
C1068 16to4_PriorityEncoder_v0p0p1_0.x5.x17.A 16to4_PriorityEncoder_v0p0p1_0.x1.A 0.115f
C1069 frontAnalog_v0p0p1_4.x65.A VIN 0.657f
C1070 frontAnalog_v0p0p1_2.x65.A a_55268_n3936# 0.461f
C1071 frontAnalog_v0p0p1_6.x63.A frontAnalog_v0p0p1_6.x63.X 0.0301f
C1072 frontAnalog_v0p0p1_6.x65.A resistorDivider_v0p0p1_0.V11 0.253f
C1073 frontAnalog_v0p0p1_9.RSfetsym_0.x1.Y VDD 0.733f
C1074 resistorDivider_v0p0p1_0.V3 VDD 4.13f
C1075 frontAnalog_v0p0p1_2.x63.X frontAnalog_v0p0p1_2.RSfetsym_0.x2.Y 0.0923f
C1076 frontAnalog_v0p0p1_6.x63.X a_59577_n30483# 0.28f
C1077 frontAnalog_v0p0p1_2.RSfetsym_0.QN a_59577_n3483# 0.418f
C1078 frontAnalog_v0p0p1_3.x65.X VDD 3.55f
C1079 frontAnalog_v0p0p1_11.x65.A frontAnalog_v0p0p1_11.x65.X 0.0236f
C1080 w_55000_n57550# resistorDivider_v0p0p1_0.V6 0.751f
C1081 a_82906_n47995# 16to4_PriorityEncoder_v0p0p1_0.x3.A1 0.121f
C1082 a_82906_n43855# 16to4_PriorityEncoder_v0p0p1_0.x3.A2 0.119f
C1083 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_7.x63.A 0.0926f
C1084 a_59578_n24570# VDD 0.0213f
C1085 16to4_PriorityEncoder_v0p0p1_0.I14 16to4_PriorityEncoder_v0p0p1_0.x5.x18.C 0.301f
C1086 16to4_PriorityEncoder_v0p0p1_0.x3.x21.B a_77605_n52819# 0.0141f
C1087 w_55000_n19750# a_53630_n20196# 0.394f
C1088 16to4_PriorityEncoder_v0p0p1_0.I12 16to4_PriorityEncoder_v0p0p1_0.x5.x20.B 0.206f
C1089 w_55000_n19128# a_55268_n20136# 0.149f
C1090 16to4_PriorityEncoder_v0p0p1_0.x1.A VDD 2.17f
C1091 16to4_PriorityEncoder_v0p0p1_0.x3.x16.C a_77605_n51335# 0.0949f
C1092 frontAnalog_v0p0p1_3.x63.A a_55268_n14736# 1.24f
C1093 frontAnalog_v0p0p1_14.x65.X CLK 0.0415f
C1094 m3_58396_n47550# VDD 1.3f
C1095 frontAnalog_v0p0p1_9.x63.A frontAnalog_v0p0p1_9.x65.A 3.16f
C1096 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0 8.68f
C1097 16to4_PriorityEncoder_v0p0p1_0.I13 a_77637_n41087# 0.194f
C1098 a_53630_n36396# resistorDivider_v0p0p1_0.V10 0.28f
C1099 16to4_PriorityEncoder_v0p0p1_0.x5.x19.C VDD 2.86f
C1100 frontAnalog_v0p0p1_15.x65.A VDD 3.45f
C1101 16to4_PriorityEncoder_v0p0p1_0.x3.EI 16to4_PriorityEncoder_v0p0p1_0.x1.A 0.534f
C1102 resistorDivider_v0p0p1_0.V12 VDD 4.13f
C1103 w_55000_n46750# CLK 0.535f
C1104 resistorDivider_v0p0p1_0.V11 resistorDivider_v0p0p1_0.V10 3.38f
C1105 frontAnalog_v0p0p1_1.x63.X frontAnalog_v0p0p1_1.RSfetsym_0.x2.Y 0.0923f
C1106 w_55000_n62950# a_55268_n63336# 0.12f
C1107 a_53630_n25596# CLK 0.0136f
C1108 w_55000_n19128# VDD 0.854f
C1109 16to4_PriorityEncoder_v0p0p1_0.x3.x4.C a_77605_n48109# 0.134f
C1110 16to4_PriorityEncoder_v0p0p1_0.x5.x20.B 16to4_PriorityEncoder_v0p0p1_0.x5.x22.C 0.0195f
C1111 w_55000_n35328# frontAnalog_v0p0p1_10.IB 0.0216f
C1112 frontAnalog_v0p0p1_1.x65.X frontAnalog_v0p0p1_1.RSfetsym_0.x1.Y 0.182f
C1113 frontAnalog_v0p0p1_3.x63.X VDD 3.16f
C1114 frontAnalog_v0p0p1_14.x63.X CLK 0.785f
C1115 16to4_PriorityEncoder_v0p0p1_0.I13 VDD 12.2f
C1116 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_8.x63.A 0.0926f
C1117 w_55000_n13728# frontAnalog_v0p0p1_3.x63.A 0.0792f
C1118 frontAnalog_v0p0p1_5.RSfetsym_0.x1.Y VDD 0.733f
C1119 resistorDivider_v0p0p1_0.V6 VIN 2.58f
C1120 frontAnalog_v0p0p1_10.x65.X CLK 0.0402f
C1121 16to4_PriorityEncoder_v0p0p1_0.x3.x16.C 16to4_PriorityEncoder_v0p0p1_0.x3.x17.D 0.07f
C1122 resistorDivider_v0p0p1_0.V1 VIN 2.01f
C1123 frontAnalog_v0p0p1_9.x65.A a_55268_n52536# 0.461f
C1124 frontAnalog_v0p0p1_11.x65.A VDD 3.45f
C1125 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_14.x63.A 0.0926f
C1126 VDD OUT1 6.71f
C1127 a_77637_n40777# VDD 0.318f
C1128 w_55000_n29928# VIN 0.866f
C1129 frontAnalog_v0p0p1_5.RSfetsym_0.QN VDD 2.56f
C1130 a_78097_n53777# VDD 0.219f
C1131 resistorDivider_v0p0p1_0.V1 a_55268_n84936# 0.214f
C1132 16to4_PriorityEncoder_v0p0p1_0.x5.x22.A 16to4_PriorityEncoder_v0p0p1_0.x1.A 0.492f
C1133 frontAnalog_v0p0p1_5.x63.A frontAnalog_v0p0p1_5.x65.A 3.16f
C1134 w_55000_n51528# resistorDivider_v0p0p1_0.V7 0.798f
C1135 a_57123_n25679# VDD 0.222f
C1136 16to4_PriorityEncoder_v0p0p1_0.x5.x18.C VDD 2.22f
C1137 16to4_PriorityEncoder_v0p0p1_0.x3.EI a_78097_n53777# 0.106f
C1138 frontAnalog_v0p0p1_2.x63.A resistorDivider_v0p0p1_0.V16 0.587f
C1139 frontAnalog_v0p0p1_2.x63.A CLK 1.8f
C1140 a_55268_n14736# CLK 0.236f
C1141 frontAnalog_v0p0p1_10.x63.X CLK 0.785f
C1142 16to4_PriorityEncoder_v0p0p1_0.I12 16to4_PriorityEncoder_v0p0p1_0.x5.x16.C 0.202f
C1143 frontAnalog_v0p0p1_0.x65.A CLK 2.61f
C1144 frontAnalog_v0p0p1_1.x65.X frontAnalog_v0p0p1_1.x63.X 0.136f
C1145 w_55000_n57550# VDD 0.829f
C1146 a_57123_n45759# VDD 0.224f
C1147 16to4_PriorityEncoder_v0p0p1_0.x3.x22.A a_77639_n50381# 0.155f
C1148 w_55000_n73750# frontAnalog_v0p0p1_10.IB 0.0217f
C1149 w_55000_n73128# frontAnalog_v0p0p1_12.x65.A 0.658f
C1150 a_53630_n74196# VDD 0.134f
C1151 a_77605_n45765# 16to4_PriorityEncoder_v0p0p1_0.x5.x22.D 0.0895f
C1152 frontAnalog_v0p0p1_6.x65.X VDD 3.55f
C1153 w_55000_n30550# resistorDivider_v0p0p1_0.V11 0.751f
C1154 16to4_PriorityEncoder_v0p0p1_0.I13 16to4_PriorityEncoder_v0p0p1_0.x5.x22.A 0.066f
C1155 16to4_PriorityEncoder_v0p0p1_0.x3.A1 16to4_PriorityEncoder_v0p0p1_0.x3.x17.D 0.0159f
C1156 16to4_PriorityEncoder_v0p0p1_0.x3.A2 a_78065_n49349# 0.144f
C1157 16to4_PriorityEncoder_v0p0p1_0.x5.x14.A a_78065_n41309# 0.197f
C1158 frontAnalog_v0p0p1_1.RSfetsym_0.x1.Y VDD 0.733f
C1159 w_55000_n73750# frontAnalog_v0p0p1_12.x63.A 0.659f
C1160 w_55000_n13728# CLK 0.571f
C1161 16to4_PriorityEncoder_v0p0p1_0.x3.x19.C a_77605_n51335# 0.173f
C1162 16to4_PriorityEncoder_v0p0p1_0.x3.x16.C 16to4_PriorityEncoder_v0p0p1_0.x3.x17.C 0.0319f
C1163 a_59577_n14283# VDD 0.0173f
C1164 a_55268_n20136# VIN 0.177f
C1165 a_53630_n41796# resistorDivider_v0p0p1_0.V9 0.28f
C1166 w_55000_n68350# VIN 0.737f
C1167 frontAnalog_v0p0p1_5.RSfetsym_0.x2.Y VDD 0.926f
C1168 w_55000_n73750# resistorDivider_v0p0p1_0.V3 0.751f
C1169 w_55000_n83928# w_55000_n84550# 0.327f
C1170 resistorDivider_v0p0p1_0.V14 resistorDivider_v0p0p1_0.V13 4.07f
C1171 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_3.x63.A 0.0926f
C1172 a_77605_n51585# VDD 0.432f
C1173 16to4_PriorityEncoder_v0p0p1_0.x22.A 16to4_PriorityEncoder_v0p0p1_0.x22.Y 1.51f
C1174 a_55268_n9336# VDD 0.565f
C1175 w_55000_n51528# a_53630_n52596# 0.359f
C1176 frontAnalog_v0p0p1_2.x65.A frontAnalog_v0p0p1_2.x65.X 0.0236f
C1177 VDD VIN 32.7f
C1178 resistorDivider_v0p0p1_0.V4 frontAnalog_v0p0p1_13.x63.A 0.587f
C1179 16to4_PriorityEncoder_v0p0p1_0.x3.A2 16to4_PriorityEncoder_v0p0p1_0.x2.A 0.401f
C1180 16to4_PriorityEncoder_v0p0p1_0.x3.EI a_77605_n51585# 0.14f
C1181 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_13.x65.A 0.0352f
C1182 a_57123_n78159# frontAnalog_v0p0p1_14.x65.X 0.119f
C1183 w_55000_n2928# frontAnalog_v0p0p1_2.x65.A 0.658f
C1184 16to4_PriorityEncoder_v0p0p1_0.x3.x17.A a_78349_n51085# 0.213f
C1185 a_53630_n3996# VIN 0.265f
C1186 frontAnalog_v0p0p1_3.x65.A a_57123_n13359# 0.214f
C1187 frontAnalog_v0p0p1_2.x63.A a_57123_n4079# 0.212f
C1188 w_55000_n29928# frontAnalog_v0p0p1_6.x63.A 0.0792f
C1189 a_55268_n84936# VDD 0.565f
C1190 frontAnalog_v0p0p1_1.x63.X VDD 3.16f
C1191 frontAnalog_v0p0p1_8.x65.A a_55268_n47136# 0.461f
C1192 frontAnalog_v0p0p1_1.RSfetsym_0.QN frontAnalog_v0p0p1_1.RSfetsym_0.x1.Y 0.17f
C1193 w_55000_n3550# frontAnalog_v0p0p1_2.x63.A 0.659f
C1194 w_55000_n46128# w_55000_n46750# 0.327f
C1195 m3_58396_n58350# VDD 1.3f
C1196 frontAnalog_v0p0p1_6.x63.X VDD 3.16f
C1197 a_77605_n45765# VDD 0.552f
C1198 16to4_PriorityEncoder_v0p0p1_0.I13 16to4_PriorityEncoder_v0p0p1_0.x5.x14.B 0.0201f
C1199 16to4_PriorityEncoder_v0p0p1_0.x3.A1 16to4_PriorityEncoder_v0p0p1_0.x3.x17.C 0.0206f
C1200 w_55000_n52150# CLK 0.535f
C1201 16to4_PriorityEncoder_v0p0p1_0.x3.x21.B 16to4_PriorityEncoder_v0p0p1_0.x3.x22.D 0.0561f
C1202 a_53630_n47196# CLK 0.0136f
C1203 a_55268_n36336# VDD 0.565f
C1204 frontAnalog_v0p0p1_10.x63.A CLK 1.81f
C1205 frontAnalog_v0p0p1_14.x65.X a_59578_n78570# 0.436f
C1206 w_55000_n14350# frontAnalog_v0p0p1_3.x65.A 0.0988f
C1207 frontAnalog_v0p0p1_7.x63.A VIN 0.187f
C1208 w_55000_n24528# VDD 0.854f
C1209 frontAnalog_v0p0p1_10.IB a_53630_n79596# 0.473f
C1210 VDD OUT0 6.72f
C1211 16to4_PriorityEncoder_v0p0p1_0.x5.x14.A 16to4_PriorityEncoder_v0p0p1_0.x5.x17.A 0.105f
C1212 16to4_PriorityEncoder_v0p0p1_0.x3.A2 16to4_PriorityEncoder_v0p0p1_0.x3.x17.A 0.047f
C1213 w_55000_n8328# frontAnalog_v0p0p1_0.x63.A 0.0792f
C1214 a_77605_n44779# VDD 0.614f
C1215 a_55268_n41736# VDD 0.565f
C1216 a_57123_n67359# frontAnalog_v0p0p1_13.x65.X 0.119f
C1217 a_55268_n30936# CLK 0.236f
C1218 w_55000_n40728# frontAnalog_v0p0p1_10.IB 0.0216f
C1219 16to4_PriorityEncoder_v0p0p1_0.I12 16to4_PriorityEncoder_v0p0p1_0.x5.x19.C 0.405f
C1220 a_55268_n63336# VDD 0.565f
C1221 frontAnalog_v0p0p1_8.RSfetsym_0.QN frontAnalog_v0p0p1_8.RSfetsym_0.x1.Y 0.17f
C1222 w_55000_n8328# w_55000_n8950# 0.327f
C1223 frontAnalog_v0p0p1_10.IB resistorDivider_v0p0p1_0.V16 6.01f
C1224 frontAnalog_v0p0p1_10.IB CLK 33.4f
C1225 frontAnalog_v0p0p1_15.RSfetsym_0.QN a_59578_n83970# 0.255f
C1226 frontAnalog_v0p0p1_0.RSfetsym_0.QN a_59578_n8370# 0.255f
C1227 frontAnalog_v0p0p1_1.RSfetsym_0.QN frontAnalog_v0p0p1_1.x63.X 0.378f
C1228 frontAnalog_v0p0p1_1.x65.X frontAnalog_v0p0p1_1.RSfetsym_0.x2.Y 0.526f
C1229 frontAnalog_v0p0p1_9.x65.A frontAnalog_v0p0p1_9.x65.X 0.0236f
C1230 frontAnalog_v0p0p1_3.x63.A frontAnalog_v0p0p1_3.x63.X 0.0301f
C1231 frontAnalog_v0p0p1_5.x63.A a_55268_n25536# 1.24f
C1232 frontAnalog_v0p0p1_8.RSfetsym_0.QN VDD 2.56f
C1233 frontAnalog_v0p0p1_12.x63.A CLK 1.81f
C1234 16to4_PriorityEncoder_v0p0p1_0.x5.x14.A VDD 0.487f
C1235 frontAnalog_v0p0p1_7.x63.A a_55268_n36336# 1.24f
C1236 frontAnalog_v0p0p1_0.x65.X 16to4_PriorityEncoder_v0p0p1_0.I14 0.445f
C1237 w_55000_n35328# VIN 0.866f
C1238 frontAnalog_v0p0p1_13.x65.X a_59578_n67770# 0.436f
C1239 resistorDivider_v0p0p1_0.V1 VL 1.96f
C1240 16to4_PriorityEncoder_v0p0p1_0.I13 16to4_PriorityEncoder_v0p0p1_0.I12 7.14f
C1241 frontAnalog_v0p0p1_8.x63.A VIN 0.186f
C1242 frontAnalog_v0p0p1_14.x65.X frontAnalog_v0p0p1_14.RSfetsym_0.x1.Y 0.182f
C1243 frontAnalog_v0p0p1_10.IB a_53630_n57996# 0.473f
C1244 16to4_PriorityEncoder_v0p0p1_0.x3.EI 16to4_PriorityEncoder_v0p0p1_0.x5.x14.A 0.0145f
C1245 frontAnalog_v0p0p1_3.x65.A resistorDivider_v0p0p1_0.V14 0.253f
C1246 resistorDivider_v0p0p1_0.V3 CLK 5.47f
C1247 a_57123_n41879# VDD 0.222f
C1248 frontAnalog_v0p0p1_6.x63.A VDD 3.67f
C1249 w_55000_n73128# a_55268_n74136# 0.149f
C1250 frontAnalog_v0p0p1_15.x65.X frontAnalog_v0p0p1_15.x63.X 0.136f
C1251 w_55000_n73750# a_53630_n74196# 0.394f
C1252 frontAnalog_v0p0p1_0.x65.X frontAnalog_v0p0p1_0.x63.X 0.136f
C1253 w_55000_n51528# frontAnalog_v0p0p1_9.x65.A 0.658f
C1254 a_57123_n56559# frontAnalog_v0p0p1_10.x65.X 0.119f
C1255 frontAnalog_v0p0p1_4.x65.A a_55268_n20136# 0.461f
C1256 frontAnalog_v0p0p1_3.x65.X CLK 0.0393f
C1257 w_55000_n19750# resistorDivider_v0p0p1_0.V13 0.751f
C1258 frontAnalog_v0p0p1_14.x63.A VIN 0.19f
C1259 a_59577_n30483# VDD 0.0173f
C1260 w_55000_n62950# VDD 0.829f
C1261 frontAnalog_v0p0p1_9.x63.X a_57123_n52679# 0.121f
C1262 16to4_PriorityEncoder_v0p0p1_0.I12 a_77637_n40777# 0.188f
C1263 16to4_PriorityEncoder_v0p0p1_0.x1.A 16to4_PriorityEncoder_v0p0p1_0.x3.A1 0.426f
C1264 frontAnalog_v0p0p1_12.RSfetsym_0.QN a_59578_n73170# 0.255f
C1265 16to4_PriorityEncoder_v0p0p1_0.x3.x22.A a_78349_n51085# 0.17f
C1266 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD 17f
C1267 frontAnalog_v0p0p1_15.RSfetsym_0.QN frontAnalog_v0p0p1_15.RSfetsym_0.x1.Y 0.17f
C1268 w_55000_n52150# frontAnalog_v0p0p1_9.x63.A 0.659f
C1269 frontAnalog_v0p0p1_0.RSfetsym_0.QN frontAnalog_v0p0p1_0.RSfetsym_0.x1.Y 0.17f
C1270 w_55000_n79150# frontAnalog_v0p0p1_10.IB 0.0217f
C1271 w_55000_n35950# a_53630_n36396# 0.394f
C1272 w_55000_n35328# a_55268_n36336# 0.149f
C1273 a_57123_n72759# VDD 0.224f
C1274 frontAnalog_v0p0p1_14.RSfetsym_0.x1.Y frontAnalog_v0p0p1_14.x63.X 0.883f
C1275 frontAnalog_v0p0p1_15.x65.A CLK 2.62f
C1276 frontAnalog_v0p0p1_4.x65.A VDD 3.45f
C1277 resistorDivider_v0p0p1_0.V12 CLK 6.38f
C1278 16to4_PriorityEncoder_v0p0p1_0.I12 16to4_PriorityEncoder_v0p0p1_0.x5.x18.C 0.432f
C1279 a_78525_n45515# 16to4_PriorityEncoder_v0p0p1_0.x5.x22.D 0.0765f
C1280 16to4_PriorityEncoder_v0p0p1_0.x21.A 16to4_PriorityEncoder_v0p0p1_0.x22.A 0.392f
C1281 16to4_PriorityEncoder_v0p0p1_0.x3.x21.B 16to4_PriorityEncoder_v0p0p1_0.x3.x22.B 0.0197f
C1282 frontAnalog_v0p0p1_10.x65.X a_59578_n56970# 0.436f
C1283 resistorDivider_v0p0p1_0.V4 a_53630_n68796# 0.28f
C1284 frontAnalog_v0p0p1_13.x65.X frontAnalog_v0p0p1_13.RSfetsym_0.x1.Y 0.182f
C1285 w_55000_n19128# CLK 0.571f
C1286 a_57123_n51159# frontAnalog_v0p0p1_9.x65.X 0.119f
C1287 frontAnalog_v0p0p1_14.x65.X frontAnalog_v0p0p1_14.RSfetsym_0.QN 2.28f
C1288 frontAnalog_v0p0p1_12.x65.X frontAnalog_v0p0p1_12.x63.X 0.136f
C1289 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_9.x63.A 0.0926f
C1290 w_55000_n73750# VIN 0.737f
C1291 16to4_PriorityEncoder_v0p0p1_0.x5.x17.A a_78065_n41309# 0.2f
C1292 frontAnalog_v0p0p1_3.x63.X CLK 0.785f
C1293 frontAnalog_v0p0p1_1.RSfetsym_0.x2.Y VDD 0.926f
C1294 16to4_PriorityEncoder_v0p0p1_0.x3.A2 16to4_PriorityEncoder_v0p0p1_0.x3.x22.A 0.0408f
C1295 frontAnalog_v0p0p1_15.RSfetsym_0.x1.Y frontAnalog_v0p0p1_15.RSfetsym_0.x2.Y 0.0254f
C1296 16to4_PriorityEncoder_v0p0p1_0.I14 frontAnalog_v0p0p1_0.x63.X 1.78f
C1297 16to4_PriorityEncoder_v0p0p1_0.x5.x14.A 16to4_PriorityEncoder_v0p0p1_0.x5.x22.A 0.0179f
C1298 frontAnalog_v0p0p1_10.IB a_55268_n68736# 0.0848f
C1299 16to4_PriorityEncoder_v0p0p1_0.I13 CLK 0.01f
C1300 frontAnalog_v0p0p1_14.x63.X a_57123_n79679# 0.121f
C1301 a_59578_n73170# VDD 0.0213f
C1302 frontAnalog_v0p0p1_11.RSfetsym_0.QN a_59578_n62370# 0.255f
C1303 w_55000_n3550# frontAnalog_v0p0p1_10.IB 0.0217f
C1304 a_53630_n14796# a_55268_n14736# 0.015f
C1305 frontAnalog_v0p0p1_7.RSfetsym_0.QN a_59578_n35370# 0.255f
C1306 frontAnalog_v0p0p1_9.x63.X frontAnalog_v0p0p1_9.RSfetsym_0.x2.Y 0.0923f
C1307 frontAnalog_v0p0p1_12.RSfetsym_0.QN frontAnalog_v0p0p1_12.RSfetsym_0.x1.Y 0.17f
C1308 a_77605_n39305# VDD 0.149f
C1309 a_82906_n47995# 16to4_PriorityEncoder_v0p0p1_0.x1.X 0.12f
C1310 frontAnalog_v0p0p1_0.x65.X VDD 3.55f
C1311 w_55000_n52150# a_55268_n52536# 0.12f
C1312 w_55000_n30550# frontAnalog_v0p0p1_6.x65.A 0.0988f
C1313 frontAnalog_v0p0p1_13.RSfetsym_0.x1.Y frontAnalog_v0p0p1_13.x63.X 0.883f
C1314 frontAnalog_v0p0p1_11.x65.A CLK 2.61f
C1315 frontAnalog_v0p0p1_14.x65.X frontAnalog_v0p0p1_14.RSfetsym_0.x2.Y 0.526f
C1316 frontAnalog_v0p0p1_14.RSfetsym_0.QN frontAnalog_v0p0p1_14.x63.X 0.378f
C1317 a_78065_n41309# VDD 0.161f
C1318 16to4_PriorityEncoder_v0p0p1_0.x22.A VDD 1.52f
C1319 frontAnalog_v0p0p1_0.RSfetsym_0.x1.Y frontAnalog_v0p0p1_0.RSfetsym_0.x2.Y 0.0254f
C1320 16to4_PriorityEncoder_v0p0p1_0.I14 16to4_PriorityEncoder_v0p0p1_0.x5.x17.A 0.0474f
C1321 frontAnalog_v0p0p1_15.x65.X VDD 3.55f
C1322 frontAnalog_v0p0p1_10.x65.X frontAnalog_v0p0p1_10.RSfetsym_0.x1.Y 0.182f
C1323 frontAnalog_v0p0p1_3.x63.A VIN 0.19f
C1324 frontAnalog_v0p0p1_8.x65.A frontAnalog_v0p0p1_8.x65.X 0.0236f
C1325 16to4_PriorityEncoder_v0p0p1_0.x3.x16.C a_77605_n51585# 0.0677f
C1326 frontAnalog_v0p0p1_13.x65.X frontAnalog_v0p0p1_13.RSfetsym_0.QN 2.28f
C1327 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_1.x65.A 0.0352f
C1328 16to4_PriorityEncoder_v0p0p1_0.x3.x21.B 16to4_PriorityEncoder_v0p0p1_0.x3.x22.C 0.262f
C1329 frontAnalog_v0p0p1_0.x63.A frontAnalog_v0p0p1_0.x65.A 3.16f
C1330 m3_58396_n69150# VDD 1.3f
C1331 frontAnalog_v0p0p1_7.x65.X frontAnalog_v0p0p1_7.x63.X 0.136f
C1332 frontAnalog_v0p0p1_11.x65.X frontAnalog_v0p0p1_11.x63.X 0.136f
C1333 frontAnalog_v0p0p1_9.x63.X a_59577_n52083# 0.28f
C1334 w_55000_n13728# a_53630_n14796# 0.359f
C1335 w_55000_n46128# a_53630_n47196# 0.359f
C1336 frontAnalog_v0p0p1_10.IB a_55268_n52536# 0.0848f
C1337 a_78525_n45515# VDD 0.165f
C1338 frontAnalog_v0p0p1_12.RSfetsym_0.x1.Y frontAnalog_v0p0p1_12.RSfetsym_0.x2.Y 0.0254f
C1339 w_55000_n83928# frontAnalog_v0p0p1_15.x63.A 0.0792f
C1340 frontAnalog_v0p0p1_13.x65.A VIN 0.655f
C1341 resistorDivider_v0p0p1_0.V6 VDD 4.67f
C1342 w_55000_n57550# CLK 0.535f
C1343 frontAnalog_v0p0p1_15.RSfetsym_0.QN frontAnalog_v0p0p1_15.RSfetsym_0.x2.Y 0.018f
C1344 frontAnalog_v0p0p1_0.RSfetsym_0.QN frontAnalog_v0p0p1_0.RSfetsym_0.x2.Y 0.018f
C1345 frontAnalog_v0p0p1_13.x63.X a_57123_n68879# 0.121f
C1346 frontAnalog_v0p0p1_4.x63.A resistorDivider_v0p0p1_0.V13 0.587f
C1347 w_55000_n8950# frontAnalog_v0p0p1_0.x65.A 0.0988f
C1348 resistorDivider_v0p0p1_0.V1 VDD 2.06f
C1349 frontAnalog_v0p0p1_7.x65.X VDD 3.55f
C1350 frontAnalog_v0p0p1_14.x63.X frontAnalog_v0p0p1_14.RSfetsym_0.x2.Y 0.0923f
C1351 frontAnalog_v0p0p1_12.RSfetsym_0.x1.Y VDD 0.733f
C1352 frontAnalog_v0p0p1_1.RSfetsym_0.QN frontAnalog_v0p0p1_1.RSfetsym_0.x2.Y 0.018f
C1353 frontAnalog_v0p0p1_11.RSfetsym_0.QN frontAnalog_v0p0p1_11.RSfetsym_0.x1.Y 0.17f
C1354 frontAnalog_v0p0p1_7.RSfetsym_0.QN frontAnalog_v0p0p1_7.RSfetsym_0.x1.Y 0.17f
C1355 resistorDivider_v0p0p1_0.V10 resistorDivider_v0p0p1_0.V9 2.78f
C1356 a_53630_n25596# a_55268_n25536# 0.015f
C1357 resistorDivider_v0p0p1_0.V9 resistorDivider_v0p0p1_0.V8 3.01f
C1358 w_55000_n29928# VDD 0.854f
C1359 a_53630_n74196# CLK 0.0136f
C1360 16to4_PriorityEncoder_v0p0p1_0.I14 VDD 7.96f
C1361 frontAnalog_v0p0p1_10.RSfetsym_0.x1.Y frontAnalog_v0p0p1_10.x63.X 0.883f
C1362 frontAnalog_v0p0p1_15.x63.X VDD 3.16f
C1363 frontAnalog_v0p0p1_15.x63.X a_59577_n84483# 0.28f
C1364 16to4_PriorityEncoder_v0p0p1_0.x5.x16.C a_77605_n43295# 0.0949f
C1365 16to4_PriorityEncoder_v0p0p1_0.x3.x22.A 16to4_PriorityEncoder_v0p0p1_0.x3.x22.B 0.0749f
C1366 frontAnalog_v0p0p1_12.x63.X m3_58396_n74550# 0.139f
C1367 16to4_PriorityEncoder_v0p0p1_0.x5.x14.A 16to4_PriorityEncoder_v0p0p1_0.x5.x14.B 0.0721f
C1368 frontAnalog_v0p0p1_10.x65.A a_55268_n57936# 0.461f
C1369 frontAnalog_v0p0p1_13.RSfetsym_0.QN frontAnalog_v0p0p1_13.x63.X 0.378f
C1370 frontAnalog_v0p0p1_13.x65.X frontAnalog_v0p0p1_13.RSfetsym_0.x2.Y 0.526f
C1371 w_55000_n46128# frontAnalog_v0p0p1_10.IB 0.0216f
C1372 frontAnalog_v0p0p1_6.x65.X CLK 0.0402f
C1373 frontAnalog_v0p0p1_1.x65.X VDD 3.55f
C1374 a_78525_n45515# 16to4_PriorityEncoder_v0p0p1_0.x5.x22.B 0.202f
C1375 16to4_PriorityEncoder_v0p0p1_0.I15 16to4_PriorityEncoder_v0p0p1_0.I11 1.03f
C1376 a_78349_n43045# 16to4_PriorityEncoder_v0p0p1_0.x5.x17.D 0.0673f
C1377 w_55000_n57550# a_53630_n57996# 0.394f
C1378 16to4_PriorityEncoder_v0p0p1_0.x5.x22.D VDD 0.473f
C1379 frontAnalog_v0p0p1_11.x65.X VDD 3.55f
C1380 frontAnalog_v0p0p1_5.x65.A a_57123_n24159# 0.214f
C1381 w_55000_n56928# a_55268_n57936# 0.149f
C1382 frontAnalog_v0p0p1_0.x63.X VDD 3.16f
C1383 frontAnalog_v0p0p1_7.x65.A a_57123_n34959# 0.214f
C1384 frontAnalog_v0p0p1_10.x65.X frontAnalog_v0p0p1_10.RSfetsym_0.QN 2.28f
C1385 16to4_PriorityEncoder_v0p0p1_0.I14 a_59577_n8883# 0.29f
C1386 a_77605_n47345# VDD 0.152f
C1387 a_57123_n74279# VDD 0.222f
C1388 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD 16.6f
C1389 frontAnalog_v0p0p1_11.RSfetsym_0.x1.Y frontAnalog_v0p0p1_11.RSfetsym_0.x2.Y 0.0254f
C1390 16to4_PriorityEncoder_v0p0p1_0.x3.x9.Y a_77605_n47345# 0.0112f
C1391 a_53630_n79596# VIN 0.265f
C1392 frontAnalog_v0p0p1_10.x63.X a_57123_n58079# 0.121f
C1393 frontAnalog_v0p0p1_12.RSfetsym_0.QN frontAnalog_v0p0p1_12.RSfetsym_0.x2.Y 0.018f
C1394 16to4_PriorityEncoder_v0p0p1_0.x21.A VDD 0.539f
C1395 frontAnalog_v0p0p1_0.x63.X a_59577_n8883# 0.28f
C1396 16to4_PriorityEncoder_v0p0p1_0.x5.x22.A a_78065_n41309# 0.077f
C1397 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_5.x65.A 0.0352f
C1398 w_55000_n40728# VIN 0.866f
C1399 16to4_PriorityEncoder_v0p0p1_0.x36.A 16to4_PriorityEncoder_v0p0p1_0.x36.Y 1.51f
C1400 frontAnalog_v0p0p1_13.x63.X frontAnalog_v0p0p1_13.RSfetsym_0.x2.Y 0.0923f
C1401 frontAnalog_v0p0p1_12.RSfetsym_0.QN VDD 2.56f
C1402 16to4_PriorityEncoder_v0p0p1_0.x3.A2 16to4_PriorityEncoder_v0p0p1_0.x3.EO 0.162f
C1403 frontAnalog_v0p0p1_14.RSfetsym_0.QN a_59577_n79083# 0.418f
C1404 16to4_PriorityEncoder_v0p0p1_0.x5.x22.D 16to4_PriorityEncoder_v0p0p1_0.x5.x22.B 0.122f
C1405 resistorDivider_v0p0p1_0.V16 VIN 2.34f
C1406 CLK VIN 46f
C1407 a_55268_n9336# CLK 0.236f
C1408 frontAnalog_v0p0p1_11.x63.X VDD 3.16f
C1409 frontAnalog_v0p0p1_12.x63.X a_59577_n73683# 0.28f
C1410 16to4_PriorityEncoder_v0p0p1_0.x5.x17.A VDD 1.36f
C1411 16to4_PriorityEncoder_v0p0p1_0.x5.x22.A a_78525_n45515# 0.209f
C1412 16to4_PriorityEncoder_v0p0p1_0.x2.X 16to4_PriorityEncoder_v0p0p1_0.x21.A 0.0749f
C1413 frontAnalog_v0p0p1_10.RSfetsym_0.QN frontAnalog_v0p0p1_10.x63.X 0.378f
C1414 frontAnalog_v0p0p1_10.x65.X frontAnalog_v0p0p1_10.RSfetsym_0.x2.Y 0.526f
C1415 a_77637_n41087# VDD 0.307f
C1416 frontAnalog_v0p0p1_4.x63.A a_57123_n20279# 0.212f
C1417 frontAnalog_v0p0p1_4.x65.A frontAnalog_v0p0p1_4.x65.X 0.0236f
C1418 16to4_PriorityEncoder_v0p0p1_0.x3.x22.A 16to4_PriorityEncoder_v0p0p1_0.x3.x22.C 0.418f
C1419 16to4_PriorityEncoder_v0p0p1_0.x3.EI 16to4_PriorityEncoder_v0p0p1_0.x5.x17.A 0.0296f
C1420 frontAnalog_v0p0p1_9.x65.X frontAnalog_v0p0p1_9.RSfetsym_0.QN 2.28f
C1421 a_77605_n44779# 16to4_PriorityEncoder_v0p0p1_0.x5.x22.C 0.0873f
C1422 w_55000_n68350# VDD 0.829f
C1423 a_55268_n84936# CLK 0.236f
C1424 frontAnalog_v0p0p1_1.x63.X CLK 0.785f
C1425 a_55268_n20136# VDD 0.565f
C1426 frontAnalog_v0p0p1_8.RSfetsym_0.x1.Y VDD 0.733f
C1427 16to4_PriorityEncoder_v0p0p1_0.I12 16to4_PriorityEncoder_v0p0p1_0.x5.x14.A 0.0493f
C1428 frontAnalog_v0p0p1_1.x65.X frontAnalog_v0p0p1_1.RSfetsym_0.QN 2.28f
C1429 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1 8.67f
C1430 16to4_PriorityEncoder_v0p0p1_0.I14 16to4_PriorityEncoder_v0p0p1_0.x5.x22.A 0.0536f
C1431 w_55000_n84550# frontAnalog_v0p0p1_10.IB 0.0217f
C1432 frontAnalog_v0p0p1_12.RSfetsym_0.x2.Y VDD 0.926f
C1433 frontAnalog_v0p0p1_6.x63.X CLK 0.785f
C1434 frontAnalog_v0p0p1_7.x63.X VDD 3.16f
C1435 a_53630_n57996# VIN 0.265f
C1436 frontAnalog_v0p0p1_10.IB a_53630_n14796# 0.473f
C1437 frontAnalog_v0p0p1_8.RSfetsym_0.QN a_59578_n46170# 0.255f
C1438 frontAnalog_v0p0p1_7.RSfetsym_0.x1.Y frontAnalog_v0p0p1_7.RSfetsym_0.x2.Y 0.0254f
C1439 a_78349_n43045# 16to4_PriorityEncoder_v0p0p1_0.x5.x17.C 0.219f
C1440 frontAnalog_v0p0p1_7.RSfetsym_0.QN frontAnalog_v0p0p1_7.RSfetsym_0.x2.Y 0.018f
C1441 frontAnalog_v0p0p1_11.RSfetsym_0.QN frontAnalog_v0p0p1_11.RSfetsym_0.x2.Y 0.018f
C1442 a_55268_n36336# CLK 0.236f
C1443 a_59577_n84483# VDD 0.0173f
C1444 frontAnalog_v0p0p1_10.x63.X frontAnalog_v0p0p1_10.RSfetsym_0.x2.Y 0.0923f
C1445 16to4_PriorityEncoder_v0p0p1_0.x3.x9.Y VDD 1.55f
C1446 frontAnalog_v0p0p1_2.x63.A frontAnalog_v0p0p1_2.x65.A 3.16f
C1447 frontAnalog_v0p0p1_13.RSfetsym_0.QN a_59577_n68283# 0.418f
C1448 a_53630_n3996# VDD 0.134f
C1449 w_55000_n40728# a_55268_n41736# 0.149f
C1450 w_55000_n24528# CLK 0.571f
C1451 16to4_PriorityEncoder_v0p0p1_0.x3.x19.C a_77605_n51585# 0.176f
C1452 w_55000_n41350# a_53630_n41796# 0.394f
C1453 16to4_PriorityEncoder_v0p0p1_0.x3.EI VDD 7.86f
C1454 frontAnalog_v0p0p1_11.x63.X a_59577_n62883# 0.28f
C1455 16to4_PriorityEncoder_v0p0p1_0.x36.A VDD 1.52f
C1456 frontAnalog_v0p0p1_5.x63.A frontAnalog_v0p0p1_5.x63.X 0.0301f
C1457 frontAnalog_v0p0p1_5.x65.A resistorDivider_v0p0p1_0.V12 0.253f
C1458 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_0.x63.A 0.0858f
C1459 16to4_PriorityEncoder_v0p0p1_0.x3.EI 16to4_PriorityEncoder_v0p0p1_0.x3.x9.Y 0.547f
C1460 w_55000_n79150# VIN 0.737f
C1461 16to4_PriorityEncoder_v0p0p1_0.x5.x16.C 16to4_PriorityEncoder_v0p0p1_0.x5.x17.D 0.07f
C1462 a_59577_n8883# VDD 0.0173f
C1463 a_55268_n41736# CLK 0.236f
C1464 16to4_PriorityEncoder_v0p0p1_0.x2.X VDD 0.351f
C1465 frontAnalog_v0p0p1_7.x65.A resistorDivider_v0p0p1_0.V10 0.252f
C1466 16to4_PriorityEncoder_v0p0p1_0.x5.x14.B a_78065_n41309# 0.202f
C1467 a_55268_n63336# CLK 0.236f
C1468 w_55000_n67728# frontAnalog_v0p0p1_13.x63.A 0.0792f
C1469 frontAnalog_v0p0p1_8.x65.X frontAnalog_v0p0p1_8.x63.X 0.136f
C1470 16to4_PriorityEncoder_v0p0p1_0.x5.A2 a_82906_n43855# 0.208f
C1471 w_55000_n8950# frontAnalog_v0p0p1_10.IB 0.0217f
C1472 16to4_PriorityEncoder_v0p0p1_0.x5.x22.B VDD 0.514f
C1473 w_55000_n83928# a_53630_n84996# 0.359f
C1474 frontAnalog_v0p0p1_7.x63.A frontAnalog_v0p0p1_7.x63.X 0.0301f
C1475 a_78649_n39527# VDD 0.414f
C1476 a_77637_n41087# 16to4_PriorityEncoder_v0p0p1_0.x5.x22.A 0.0288f
C1477 16to4_PriorityEncoder_v0p0p1_0.x5.x19.C a_77605_n43295# 0.173f
C1478 16to4_PriorityEncoder_v0p0p1_0.x5.x22.A 16to4_PriorityEncoder_v0p0p1_0.x5.x17.A 1.27f
C1479 a_53630_n20196# resistorDivider_v0p0p1_0.V13 0.28f
C1480 16to4_PriorityEncoder_v0p0p1_0.I11 m3_58396_n25950# 0.0416f
C1481 frontAnalog_v0p0p1_7.x63.A VDD 3.67f
C1482 frontAnalog_v0p0p1_9.x63.A VIN 0.187f
C1483 a_59577_n62883# VDD 0.0173f
C1484 w_55000_n84550# frontAnalog_v0p0p1_15.x65.A 0.0988f
C1485 resistorDivider_v0p0p1_0.V2 frontAnalog_v0p0p1_14.x65.A 0.253f
C1486 a_55268_n68736# VIN 0.177f
C1487 frontAnalog_v0p0p1_10.RSfetsym_0.QN a_59577_n57483# 0.418f
C1488 16to4_PriorityEncoder_v0p0p1_0.I14 a_77637_n42017# 0.186f
C1489 w_55000_n8328# a_53630_n9396# 0.359f
C1490 frontAnalog_v0p0p1_5.x63.X m3_58396_n25950# 0.139f
C1491 frontAnalog_v0p0p1_10.x63.A a_57123_n58079# 0.212f
C1492 w_55000_n3550# VIN 0.735f
C1493 a_78349_n51085# 16to4_PriorityEncoder_v0p0p1_0.x3.x17.D 0.0673f
C1494 frontAnalog_v0p0p1_1.RSfetsym_0.QN VDD 2.56f
C1495 frontAnalog_v0p0p1_7.x63.X a_59577_n35883# 0.28f
C1496 frontAnalog_v0p0p1_6.x63.A CLK 1.81f
C1497 w_55000_n51528# w_55000_n52150# 0.327f
C1498 16to4_PriorityEncoder_v0p0p1_0.x1.A 16to4_PriorityEncoder_v0p0p1_0.x28.A 0.0126f
C1499 m3_58396_n79950# VDD 1.3f
C1500 w_55000_n46750# a_55268_n47136# 0.12f
C1501 w_55000_n14350# a_55268_n14736# 0.12f
C1502 resistorDivider_v0p0p1_0.V8 frontAnalog_v0p0p1_8.x65.A 0.253f
C1503 16to4_PriorityEncoder_v0p0p1_0.x5.x22.A VDD 3.25f
C1504 a_59577_n35883# VDD 0.0173f
C1505 w_55000_n62950# CLK 0.535f
C1506 w_55000_n35950# resistorDivider_v0p0p1_0.V10 0.751f
C1507 16to4_PriorityEncoder_v0p0p1_0.x3.x22.A a_78525_n53555# 0.209f
C1508 16to4_PriorityEncoder_v0p0p1_0.I11 16to4_PriorityEncoder_v0p0p1_0.x5.x9.Y 0.0406f
C1509 16to4_PriorityEncoder_v0p0p1_0.x3.EI 16to4_PriorityEncoder_v0p0p1_0.x5.x22.A 0.208f
C1510 16to4_PriorityEncoder_v0p0p1_0.x35.A VDD 0.539f
C1511 w_55000_n35328# VDD 0.854f
C1512 frontAnalog_v0p0p1_1.x65.A VIN 0.655f
C1513 16to4_PriorityEncoder_v0p0p1_0.x5.x16.C 16to4_PriorityEncoder_v0p0p1_0.x5.x17.C 0.0319f
C1514 16to4_PriorityEncoder_v0p0p1_0.I14 m3_58396_n9750# 0.0416f
C1515 frontAnalog_v0p0p1_4.x65.A CLK 2.61f
C1516 frontAnalog_v0p0p1_10.x65.A frontAnalog_v0p0p1_10.x65.X 0.0236f
C1517 16to4_PriorityEncoder_v0p0p1_0.x35.A 16to4_PriorityEncoder_v0p0p1_0.x36.A 0.392f
C1518 frontAnalog_v0p0p1_8.x63.A VDD 3.67f
C1519 w_55000_n51528# frontAnalog_v0p0p1_10.IB 0.0216f
C1520 frontAnalog_v0p0p1_9.x65.X frontAnalog_v0p0p1_9.RSfetsym_0.x1.Y 0.182f
C1521 a_55268_n52536# VIN 0.177f
C1522 16to4_PriorityEncoder_v0p0p1_0.x5.x22.A 16to4_PriorityEncoder_v0p0p1_0.x5.x22.B 0.0749f
C1523 w_55000_n13728# w_55000_n14350# 0.327f
C1524 16to4_PriorityEncoder_v0p0p1_0.x5.x17.A a_77637_n42017# 0.14f
C1525 frontAnalog_v0p0p1_10.IB a_55268_n25536# 0.0848f
C1526 frontAnalog_v0p0p1_0.x63.X m3_58396_n9750# 0.139f
C1527 a_53630_n30996# a_55268_n30936# 0.015f
C1528 16to4_PriorityEncoder_v0p0p1_0.x5.x14.B 16to4_PriorityEncoder_v0p0p1_0.x5.x17.A 0.125f
C1529 a_77637_n41087# 16to4_PriorityEncoder_v0p0p1_0.x5.x14.B 0.109f
C1530 a_78649_n47567# VDD 0.235f
C1531 w_55000_n78528# resistorDivider_v0p0p1_0.V2 0.798f
C1532 frontAnalog_v0p0p1_14.x63.A VDD 3.67f
C1533 16to4_PriorityEncoder_v0p0p1_0.x3.x20.B VDD 1.32f
C1534 frontAnalog_v0p0p1_10.IB a_53630_n30996# 0.473f
C1535 a_55268_n14736# resistorDivider_v0p0p1_0.V14 0.215f
C1536 16to4_PriorityEncoder_v0p0p1_0.I14 16to4_PriorityEncoder_v0p0p1_0.I12 2.36f
C1537 16to4_PriorityEncoder_v0p0p1_0.x3.EI 16to4_PriorityEncoder_v0p0p1_0.x3.x20.B 1.93f
C1538 16to4_PriorityEncoder_v0p0p1_0.x3.EI a_78649_n47567# 0.181f
C1539 16to4_PriorityEncoder_v0p0p1_0.x3.A0 VDD 0.829f
C1540 16to4_PriorityEncoder_v0p0p1_0.x3.x20.B 16to4_PriorityEncoder_v0p0p1_0.x3.x9.Y 0.0516f
C1541 w_55000_n46128# VIN 0.866f
C1542 16to4_PriorityEncoder_v0p0p1_0.x5.x22.C a_78525_n45515# 0.193f
C1543 a_78349_n51085# 16to4_PriorityEncoder_v0p0p1_0.x3.x17.C 0.219f
C1544 w_55000_n35328# frontAnalog_v0p0p1_7.x63.A 0.0792f
C1545 16to4_PriorityEncoder_v0p0p1_0.x5.x20.B 16to4_PriorityEncoder_v0p0p1_0.x5.x21.B 0.151f
C1546 frontAnalog_v0p0p1_8.RSfetsym_0.QN frontAnalog_v0p0p1_8.RSfetsym_0.x2.Y 0.018f
C1547 frontAnalog_v0p0p1_0.x65.X CLK 0.0389f
C1548 16to4_PriorityEncoder_v0p0p1_0.x5.x17.D 16to4_PriorityEncoder_v0p0p1_0.x1.A 0.0159f
C1549 16to4_PriorityEncoder_v0p0p1_0.x1.A 16to4_PriorityEncoder_v0p0p1_0.x1.X 0.0412f
C1550 a_77637_n42017# VDD 0.322f
C1551 16to4_PriorityEncoder_v0p0p1_0.x5.x14.B VDD 0.514f
C1552 frontAnalog_v0p0p1_2.x65.A frontAnalog_v0p0p1_10.IB 0.0352f
C1553 frontAnalog_v0p0p1_1.x65.A a_55268_n41736# 0.461f
C1554 frontAnalog_v0p0p1_15.x65.X CLK 0.0406f
C1555 frontAnalog_v0p0p1_4.x65.X VDD 3.55f
C1556 16to4_PriorityEncoder_v0p0p1_0.x34.A VDD 0.347f
C1557 w_55000_n73750# VDD 0.829f
C1558 frontAnalog_v0p0p1_5.x65.A VIN 0.655f
C1559 16to4_PriorityEncoder_v0p0p1_0.x2.A a_82906_n51645# 0.207f
C1560 resistorDivider_v0p0p1_0.V8 resistorDivider_v0p0p1_0.V7 3.46f
C1561 w_55000_n13728# resistorDivider_v0p0p1_0.V14 0.798f
C1562 16to4_PriorityEncoder_v0p0p1_0.x5.x22.C 16to4_PriorityEncoder_v0p0p1_0.x5.x22.D 0.145f
C1563 w_55000_n67728# a_53630_n68796# 0.359f
C1564 resistorDivider_v0p0p1_0.V6 CLK 6.01f
C1565 a_55268_n25536# resistorDivider_v0p0p1_0.V12 0.215f
C1566 resistorDivider_v0p0p1_0.V1 CLK 5.44f
C1567 frontAnalog_v0p0p1_7.x65.X CLK 0.0389f
C1568 m3_58396_n9750# VDD 1.3f
C1569 16to4_PriorityEncoder_v0p0p1_0.I11 16to4_PriorityEncoder_v0p0p1_0.x5.x20.B 1.27f
C1570 a_57123_n2559# VDD 0.224f
C1571 w_55000_n29928# CLK 0.571f
C1572 w_55000_n68350# frontAnalog_v0p0p1_13.x65.A 0.0988f
C1573 frontAnalog_v0p0p1_15.x63.X CLK 0.785f
C1574 frontAnalog_v0p0p1_10.IB resistorDivider_v0p0p1_0.V5 3.69f
C1575 16to4_PriorityEncoder_v0p0p1_0.I14 CLK 0.01f
C1576 frontAnalog_v0p0p1_3.x63.A VDD 3.67f
C1577 frontAnalog_v0p0p1_1.x65.X CLK 0.0393f
C1578 w_55000_n84550# VIN 0.737f
C1579 a_53630_n14796# VIN 0.265f
C1580 resistorDivider_v0p0p1_0.V6 a_53630_n57996# 0.28f
C1581 frontAnalog_v0p0p1_11.x65.X CLK 0.0398f
C1582 w_55000_n24528# frontAnalog_v0p0p1_5.x65.A 0.658f
C1583 16to4_PriorityEncoder_v0p0p1_0.x3.x16.C VDD 0.834f
C1584 16to4_PriorityEncoder_v0p0p1_0.I12 VDD 11.6f
C1585 frontAnalog_v0p0p1_0.x63.X CLK 0.785f
C1586 frontAnalog_v0p0p1_13.x65.A VDD 3.45f
C1587 w_55000_n14350# frontAnalog_v0p0p1_10.IB 0.0217f
C1588 16to4_PriorityEncoder_v0p0p1_0.x5.x17.C 16to4_PriorityEncoder_v0p0p1_0.x1.A 0.0206f
C1589 16to4_PriorityEncoder_v0p0p1_0.x43.Y 16to4_PriorityEncoder_v0p0p1_0.x5.A2 0.0114f
C1590 a_57123_n13359# frontAnalog_v0p0p1_3.x65.X 0.119f
C1591 w_55000_n84550# a_55268_n84936# 0.12f
C1592 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_15.x63.A 0.0926f
C1593 a_77605_n52567# VDD 0.432f
C1594 resistorDivider_v0p0p1_0.V2 a_55268_n79536# 0.215f
C1595 16to4_PriorityEncoder_v0p0p1_0.x3.EI 16to4_PriorityEncoder_v0p0p1_0.x3.x16.C 2.08f
C1596 16to4_PriorityEncoder_v0p0p1_0.x5.x14.B 16to4_PriorityEncoder_v0p0p1_0.x5.x22.A 0.0936f
C1597 frontAnalog_v0p0p1_9.RSfetsym_0.QN a_59578_n51570# 0.255f
C1598 w_55000_n25150# frontAnalog_v0p0p1_5.x63.A 0.659f
C1599 frontAnalog_v0p0p1_0.x63.A VIN 0.19f
C1600 frontAnalog_v0p0p1_0.x63.A a_55268_n9336# 1.24f
C1601 frontAnalog_v0p0p1_4.x63.X VDD 3.16f
C1602 a_59578_n46170# VDD 0.0213f
C1603 16to4_PriorityEncoder_v0p0p1_0.x5.x22.C VDD 0.938f
C1604 w_55000_n8950# a_55268_n9336# 0.12f
C1605 w_55000_n8950# VIN 0.737f
C1606 frontAnalog_v0p0p1_11.x63.X CLK 0.785f
C1607 16to4_PriorityEncoder_v0p0p1_0.x34.A 16to4_PriorityEncoder_v0p0p1_0.x35.A 0.0737f
C1608 frontAnalog_v0p0p1_10.x63.A frontAnalog_v0p0p1_10.x65.A 3.16f
C1609 16to4_PriorityEncoder_v0p0p1_0.I15 frontAnalog_v0p0p1_0.RSfetsym_0.QN 0.0512f
C1610 frontAnalog_v0p0p1_6.x63.X m3_58396_n31350# 0.139f
C1611 a_55268_n20136# CLK 0.236f
C1612 a_53630_n47196# a_55268_n47136# 0.015f
C1613 w_55000_n56928# frontAnalog_v0p0p1_10.x63.A 0.0792f
C1614 w_55000_n68350# CLK 0.535f
C1615 16to4_PriorityEncoder_v0p0p1_0.x1.A 16to4_PriorityEncoder_v0p0p1_0.x3.A2 1.46f
C1616 a_53630_n79596# VDD 0.134f
C1617 frontAnalog_v0p0p1_10.IB resistorDivider_v0p0p1_0.V14 3.7f
C1618 frontAnalog_v0p0p1_3.x65.X a_59578_n13770# 0.436f
C1619 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_11.x63.A 0.0926f
C1620 16to4_PriorityEncoder_v0p0p1_0.x3.x14.A VDD 0.462f
C1621 a_57123_n24159# frontAnalog_v0p0p1_5.x65.X 0.119f
C1622 frontAnalog_v0p0p1_7.x63.X CLK 0.785f
C1623 w_55000_n40728# VDD 0.854f
C1624 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_10.x65.A 0.0352f
C1625 16to4_PriorityEncoder_v0p0p1_0.x3.A1 VDD 1.93f
C1626 a_77605_n44527# 16to4_PriorityEncoder_v0p0p1_0.x5.x21.B 0.116f
C1627 16to4_PriorityEncoder_v0p0p1_0.x5.x22.C 16to4_PriorityEncoder_v0p0p1_0.x5.x22.B 0.131f
C1628 a_59578_n2970# VDD 0.0213f
C1629 16to4_PriorityEncoder_v0p0p1_0.x3.EI 16to4_PriorityEncoder_v0p0p1_0.x3.x14.A 0.0111f
C1630 w_55000_n56928# frontAnalog_v0p0p1_10.IB 0.0216f
C1631 resistorDivider_v0p0p1_0.V16 VDD 4.5f
C1632 VDD CLK 73.4f
C1633 frontAnalog_v0p0p1_15.x63.A frontAnalog_v0p0p1_15.x65.A 3.16f
C1634 16to4_PriorityEncoder_v0p0p1_0.I11 16to4_PriorityEncoder_v0p0p1_0.x5.x16.C 0.132f
C1635 frontAnalog_v0p0p1_10.IB a_55268_n47136# 0.0848f
C1636 a_53630_n3996# resistorDivider_v0p0p1_0.V16 0.28f
C1637 a_78159_n39549# 16to4_PriorityEncoder_v0p0p1_0.x5.x4.C 0.121f
C1638 a_53630_n3996# CLK 0.0136f
C1639 a_78097_n53777# 16to4_PriorityEncoder_v0p0p1_0.x3.x22.D 0.137f
C1640 frontAnalog_v0p0p1_10.IB resistorDivider_v0p0p1_0.V4 3.7f
C1641 w_55000_n35950# frontAnalog_v0p0p1_7.x65.A 0.0988f
C1642 16to4_PriorityEncoder_v0p0p1_0.I15 a_77605_n40069# 0.0614f
C1643 resistorDivider_v0p0p1_0.V5 frontAnalog_v0p0p1_11.x65.A 0.253f
C1644 w_55000_n51528# VIN 0.866f
C1645 a_53630_n57996# VDD 0.134f
C1646 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_12.x65.A 0.0352f
C1647 16to4_PriorityEncoder_v0p0p1_0.x5.x22.A 16to4_PriorityEncoder_v0p0p1_0.x5.x22.C 0.418f
C1648 16to4_PriorityEncoder_v0p0p1_0.x5.x4.C a_77605_n40069# 0.134f
C1649 a_59577_n19683# VDD 0.0173f
C1650 16to4_PriorityEncoder_v0p0p1_0.I13 a_59578_n13770# 0.42f
C1651 a_57123_n47279# VDD 0.222f
C1652 frontAnalog_v0p0p1_3.x65.X frontAnalog_v0p0p1_3.RSfetsym_0.x1.Y 0.182f
C1653 a_55268_n25536# VIN 0.177f
C1654 16to4_PriorityEncoder_v0p0p1_0.x3.x16.C 16to4_PriorityEncoder_v0p0p1_0.x3.x20.B 1.24f
C1655 a_77639_n42341# VDD 0.318f
C1656 resistorDivider_v0p0p1_0.V4 resistorDivider_v0p0p1_0.V3 5.64f
C1657 frontAnalog_v0p0p1_7.x63.A CLK 1.81f
C1658 w_55000_n8328# resistorDivider_v0p0p1_0.V15 0.798f
C1659 16to4_PriorityEncoder_v0p0p1_0.x3.x20.B a_77605_n52567# 0.14f
C1660 frontAnalog_v0p0p1_12.x63.A frontAnalog_v0p0p1_12.x65.A 3.16f
C1661 frontAnalog_v0p0p1_1.x65.A frontAnalog_v0p0p1_1.x65.X 0.0236f
C1662 frontAnalog_v0p0p1_2.RSfetsym_0.QN VDD 2.56f
C1663 frontAnalog_v0p0p1_2.RSfetsym_0.x1.Y VDD 0.733f
C1664 a_53630_n30996# VIN 0.265f
C1665 16to4_PriorityEncoder_v0p0p1_0.x3.x19.C VDD 1.19f
C1666 frontAnalog_v0p0p1_5.x65.X a_59578_n24570# 0.436f
C1667 w_55000_n79150# VDD 0.829f
C1668 resistorDivider_v0p0p1_0.V3 frontAnalog_v0p0p1_12.x65.A 0.253f
C1669 frontAnalog_v0p0p1_10.IB a_53630_n9396# 0.473f
C1670 16to4_PriorityEncoder_v0p0p1_0.x3.EI 16to4_PriorityEncoder_v0p0p1_0.x3.x19.C 1.71f
C1671 frontAnalog_v0p0p1_1.x63.A resistorDivider_v0p0p1_0.V9 0.587f
C1672 frontAnalog_v0p0p1_4.RSfetsym_0.QN a_59578_n19170# 0.255f
C1673 w_55000_n68350# a_55268_n68736# 0.12f
C1674 frontAnalog_v0p0p1_8.RSfetsym_0.x1.Y frontAnalog_v0p0p1_8.RSfetsym_0.x2.Y 0.0254f
C1675 16to4_PriorityEncoder_v0p0p1_0.x5.x19.C 16to4_PriorityEncoder_v0p0p1_0.x5.x21.B 0.0127f
C1676 frontAnalog_v0p0p1_3.x65.X frontAnalog_v0p0p1_3.RSfetsym_0.QN 2.28f
C1677 m3_58396_n20550# VDD 1.3f
C1678 a_78159_n39549# 16to4_PriorityEncoder_v0p0p1_0.x5.x4.B 0.192f
C1679 frontAnalog_v0p0p1_10.IB a_53630_n84996# 0.473f
C1680 frontAnalog_v0p0p1_2.x65.A VIN 0.653f
C1681 frontAnalog_v0p0p1_4.x65.X 16to4_PriorityEncoder_v0p0p1_0.I12 0.446f
C1682 w_55000_n41350# resistorDivider_v0p0p1_0.V9 0.751f
C1683 a_57123_n4079# VDD 0.222f
C1684 w_55000_n35328# CLK 0.571f
C1685 w_55000_n24528# a_55268_n25536# 0.149f
C1686 w_55000_n25150# a_53630_n25596# 0.394f
C1687 frontAnalog_v0p0p1_9.x63.A VDD 3.67f
C1688 frontAnalog_v0p0p1_3.RSfetsym_0.x1.Y frontAnalog_v0p0p1_3.x63.X 0.883f
C1689 16to4_PriorityEncoder_v0p0p1_0.I13 frontAnalog_v0p0p1_3.RSfetsym_0.x1.Y 0.0436f
C1690 a_55268_n68736# VDD 0.565f
C1691 frontAnalog_v0p0p1_8.RSfetsym_0.x2.Y VDD 0.926f
C1692 frontAnalog_v0p0p1_8.x63.A CLK 1.81f
C1693 w_55000_n3550# VDD 0.829f
C1694 frontAnalog_v0p0p1_11.x63.A frontAnalog_v0p0p1_11.x65.A 3.16f
C1695 a_55268_n30936# resistorDivider_v0p0p1_0.V11 0.215f
C1696 frontAnalog_v0p0p1_4.x65.X frontAnalog_v0p0p1_4.x63.X 0.136f
C1697 frontAnalog_v0p0p1_10.IB a_53630_n36396# 0.473f
C1698 frontAnalog_v0p0p1_0.x65.A a_57123_n7959# 0.214f
C1699 w_55000_n2928# a_55268_n3936# 0.149f
C1700 16to4_PriorityEncoder_v0p0p1_0.I11 a_59578_n24570# 0.42f
C1701 w_55000_n3550# a_53630_n3996# 0.394f
C1702 frontAnalog_v0p0p1_10.IB resistorDivider_v0p0p1_0.V11 3.7f
C1703 w_55000_n19750# frontAnalog_v0p0p1_10.IB 0.0217f
C1704 frontAnalog_v0p0p1_5.x65.X frontAnalog_v0p0p1_5.RSfetsym_0.x1.Y 0.182f
C1705 a_78159_n39549# 16to4_PriorityEncoder_v0p0p1_0.x5.EO 0.128f
C1706 16to4_PriorityEncoder_v0p0p1_0.x5.x16.C a_77605_n43545# 0.0677f
C1707 frontAnalog_v0p0p1_14.x63.A CLK 1.81f
C1708 16to4_PriorityEncoder_v0p0p1_0.x5.x22.A a_77639_n42341# 0.155f
C1709 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD 16.6f
C1710 a_78097_n53777# 16to4_PriorityEncoder_v0p0p1_0.x3.x22.B 0.109f
C1711 frontAnalog_v0p0p1_4.RSfetsym_0.QN frontAnalog_v0p0p1_4.RSfetsym_0.x1.Y 0.17f
C1712 frontAnalog_v0p0p1_10.IB a_53630_n41796# 0.473f
C1713 resistorDivider_v0p0p1_0.V5 VIN 2.63f
C1714 16to4_PriorityEncoder_v0p0p1_0.x3.x18.C VDD 0.691f
C1715 frontAnalog_v0p0p1_10.IB a_53630_n63396# 0.473f
C1716 frontAnalog_v0p0p1_3.x63.X a_57123_n14879# 0.121f
C1717 16to4_PriorityEncoder_v0p0p1_0.I11 16to4_PriorityEncoder_v0p0p1_0.x5.x19.C 0.921f
C1718 frontAnalog_v0p0p1_3.RSfetsym_0.QN frontAnalog_v0p0p1_3.x63.X 0.378f
C1719 frontAnalog_v0p0p1_3.RSfetsym_0.QN 16to4_PriorityEncoder_v0p0p1_0.I13 2.02f
C1720 frontAnalog_v0p0p1_3.x65.X frontAnalog_v0p0p1_3.RSfetsym_0.x2.Y 0.526f
C1721 16to4_PriorityEncoder_v0p0p1_0.x5.EO 16to4_PriorityEncoder_v0p0p1_0.x5.A2 0.136f
C1722 frontAnalog_v0p0p1_1.x65.A VDD 3.45f
C1723 frontAnalog_v0p0p1_5.x65.X frontAnalog_v0p0p1_5.RSfetsym_0.QN 2.28f
C1724 16to4_PriorityEncoder_v0p0p1_0.x3.EI 16to4_PriorityEncoder_v0p0p1_0.x3.x18.C 1.56f
C1725 w_55000_n84550# resistorDivider_v0p0p1_0.V1 0.751f
C1726 w_55000_n57550# frontAnalog_v0p0p1_10.x65.A 0.0988f
C1727 frontAnalog_v0p0p1_1.x63.X m3_58396_n42150# 0.139f
C1728 frontAnalog_v0p0p1_8.x63.A a_57123_n47279# 0.212f
C1729 a_55268_n52536# VDD 0.565f
C1730 frontAnalog_v0p0p1_9.RSfetsym_0.QN frontAnalog_v0p0p1_9.x63.X 0.378f
C1731 frontAnalog_v0p0p1_2.RSfetsym_0.x2.Y VDD 0.926f
C1732 w_55000_n14350# VIN 0.737f
C1733 16to4_PriorityEncoder_v0p0p1_0.I15 m3_58396_n4350# 0.0416f
C1734 frontAnalog_v0p0p1_15.x63.A VIN 0.188f
C1735 w_55000_n56928# w_55000_n57550# 0.327f
C1736 16to4_PriorityEncoder_v0p0p1_0.x5.x18.C 16to4_PriorityEncoder_v0p0p1_0.x5.x21.B 0.014f
C1737 a_78159_n47589# 16to4_PriorityEncoder_v0p0p1_0.x3.x4.C 0.121f
C1738 16to4_PriorityEncoder_v0p0p1_0.x5.x9.Y a_78159_n39549# 0.299f
C1739 w_55000_n78528# frontAnalog_v0p0p1_14.x65.A 0.658f
C1740 16to4_PriorityEncoder_v0p0p1_0.I12 frontAnalog_v0p0p1_4.x63.X 1.85f
C1741 frontAnalog_v0p0p1_4.x65.X CLK 0.0393f
C1742 a_77605_n48109# VDD 0.154f
C1743 w_55000_n73750# CLK 0.535f
C1744 16to4_PriorityEncoder_v0p0p1_0.I13 16to4_PriorityEncoder_v0p0p1_0.I11 1.27f
C1745 a_57123_n78159# VDD 0.224f
C1746 frontAnalog_v0p0p1_15.x63.A a_55268_n84936# 1.24f
C1747 w_55000_n46750# resistorDivider_v0p0p1_0.V8 0.751f
C1748 16to4_PriorityEncoder_v0p0p1_0.I11 frontAnalog_v0p0p1_5.RSfetsym_0.x1.Y 0.0436f
C1749 16to4_PriorityEncoder_v0p0p1_0.x3.x19.C 16to4_PriorityEncoder_v0p0p1_0.x3.x20.B 0.996f
C1750 w_55000_n46128# VDD 0.854f
C1751 w_55000_n79150# frontAnalog_v0p0p1_14.x63.A 0.659f
C1752 resistorDivider_v0p0p1_0.V12 resistorDivider_v0p0p1_0.V11 3.43f
C1753 w_55000_n62328# frontAnalog_v0p0p1_10.IB 0.0216f
C1754 frontAnalog_v0p0p1_2.x63.X m3_58396_n4350# 0.139f
C1755 frontAnalog_v0p0p1_5.RSfetsym_0.x1.Y frontAnalog_v0p0p1_5.x63.X 0.883f
C1756 frontAnalog_v0p0p1_3.x63.X frontAnalog_v0p0p1_3.RSfetsym_0.x2.Y 0.0923f
C1757 16to4_PriorityEncoder_v0p0p1_0.I13 frontAnalog_v0p0p1_3.RSfetsym_0.x2.Y 0.196f
C1758 frontAnalog_v0p0p1_5.RSfetsym_0.QN 16to4_PriorityEncoder_v0p0p1_0.I11 2.02f
C1759 resistorDivider_v0p0p1_0.V5 a_55268_n63336# 0.215f
C1760 w_55000_n19128# w_55000_n19750# 0.327f
C1761 16to4_PriorityEncoder_v0p0p1_0.x29.A VDD 1.52f
C1762 frontAnalog_v0p0p1_4.RSfetsym_0.x1.Y frontAnalog_v0p0p1_4.RSfetsym_0.x2.Y 0.0254f
C1763 resistorDivider_v0p0p1_0.V14 VIN 2.56f
C1764 a_57123_n29559# frontAnalog_v0p0p1_6.x65.X 0.119f
C1765 frontAnalog_v0p0p1_10.IB a_55268_n74136# 0.0848f
C1766 a_59578_n78570# VDD 0.0213f
C1767 frontAnalog_v0p0p1_11.x63.A VIN 0.187f
C1768 frontAnalog_v0p0p1_5.x65.A VDD 3.45f
C1769 frontAnalog_v0p0p1_0.x65.A resistorDivider_v0p0p1_0.V15 0.253f
C1770 16to4_PriorityEncoder_v0p0p1_0.x3.x17.A a_78065_n49349# 0.2f
C1771 frontAnalog_v0p0p1_0.x63.A frontAnalog_v0p0p1_0.x63.X 0.0301f
C1772 frontAnalog_v0p0p1_3.x63.A CLK 1.81f
C1773 16to4_PriorityEncoder_v0p0p1_0.I11 16to4_PriorityEncoder_v0p0p1_0.x5.x18.C 0.251f
C1774 frontAnalog_v0p0p1_10.x65.A VIN 0.655f
C1775 frontAnalog_v0p0p1_13.x63.X m3_58396_n69150# 0.139f
C1776 frontAnalog_v0p0p1_5.x65.X frontAnalog_v0p0p1_5.RSfetsym_0.x2.Y 0.526f
C1777 frontAnalog_v0p0p1_5.RSfetsym_0.QN frontAnalog_v0p0p1_5.x63.X 0.378f
C1778 frontAnalog_v0p0p1_4.RSfetsym_0.QN frontAnalog_v0p0p1_4.RSfetsym_0.x2.Y 0.018f
C1779 frontAnalog_v0p0p1_12.x63.A a_55268_n74136# 1.24f
C1780 a_57123_n56559# VDD 0.224f
C1781 w_55000_n56928# VIN 0.866f
C1782 16to4_PriorityEncoder_v0p0p1_0.I12 CLK 0.01f
C1783 frontAnalog_v0p0p1_13.x65.A CLK 2.61f
C1784 a_55268_n47136# VIN 0.177f
C1785 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_4.x63.A 0.0926f
C1786 frontAnalog_v0p0p1_5.x63.X a_57123_n25679# 0.121f
C1787 a_77605_n52819# VDD 0.435f
C1788 frontAnalog_v0p0p1_3.RSfetsym_0.QN a_59577_n14283# 0.418f
C1789 a_78159_n47589# 16to4_PriorityEncoder_v0p0p1_0.x3.x4.B 0.192f
C1790 frontAnalog_v0p0p1_4.x63.X CLK 0.785f
C1791 resistorDivider_v0p0p1_0.V3 a_55268_n74136# 0.215f
C1792 resistorDivider_v0p0p1_0.V4 VIN 2.6f
C1793 a_77605_n43295# VDD 0.551f
C1794 VL GND 0.131p
C1795 OUT0 GND 30.2f
C1796 OUT1 GND 30.3f
C1797 OUT2 GND 30.2f
C1798 OUT3 GND 31.9f
C1799 VFS GND 0.114p
C1800 VIN GND 0.208p
C1801 CLK GND 0.279p
C1802 VDD GND 2.19p
C1803 m3_58396_n85350# GND 0.216f $ **FLOATING
C1804 m3_58396_n79950# GND 0.216f $ **FLOATING
C1805 m3_58396_n74550# GND 0.216f $ **FLOATING
C1806 m3_58396_n69150# GND 0.216f $ **FLOATING
C1807 m3_58396_n63750# GND 0.216f $ **FLOATING
C1808 m3_58396_n58350# GND 0.216f $ **FLOATING
C1809 m3_58396_n52950# GND 0.216f $ **FLOATING
C1810 m3_58396_n47550# GND 0.216f $ **FLOATING
C1811 m3_58396_n42150# GND 0.216f $ **FLOATING
C1812 m3_58396_n36750# GND 0.216f $ **FLOATING
C1813 m3_58396_n31350# GND 0.216f $ **FLOATING
C1814 m3_58396_n25950# GND 0.216f $ **FLOATING
C1815 m3_58396_n20550# GND 0.216f $ **FLOATING
C1816 m3_58396_n15150# GND 0.216f $ **FLOATING
C1817 m3_58396_n9750# GND 0.216f $ **FLOATING
C1818 m3_58396_n4350# GND 0.216f $ **FLOATING
C1819 a_59577_n84483# GND 0.561f
C1820 a_57123_n85079# GND 0.319f
C1821 frontAnalog_v0p0p1_15.RSfetsym_0.x2.Y GND 1.53f
C1822 frontAnalog_v0p0p1_15.x63.X GND 5.15f
C1823 a_59578_n83970# GND 0.555f
C1824 frontAnalog_v0p0p1_15.RSfetsym_0.x1.Y GND 1.93f
C1825 frontAnalog_v0p0p1_15.RSfetsym_0.QN GND 3.84f
C1826 frontAnalog_v0p0p1_15.x65.X GND 5.07f
C1827 a_57123_n83559# GND 0.318f
C1828 a_55268_n84936# GND 1.17f
C1829 a_53630_n84996# GND 2.61f
C1830 frontAnalog_v0p0p1_15.x65.A GND 2.63f
C1831 frontAnalog_v0p0p1_15.x63.A GND 2.46f
C1832 a_59577_n79083# GND 0.561f
C1833 a_57123_n79679# GND 0.319f
C1834 frontAnalog_v0p0p1_14.RSfetsym_0.x2.Y GND 1.53f
C1835 frontAnalog_v0p0p1_14.x63.X GND 5.15f
C1836 a_59578_n78570# GND 0.555f
C1837 frontAnalog_v0p0p1_14.RSfetsym_0.x1.Y GND 1.93f
C1838 frontAnalog_v0p0p1_14.RSfetsym_0.QN GND 3.84f
C1839 frontAnalog_v0p0p1_14.x65.X GND 5.07f
C1840 a_57123_n78159# GND 0.318f
C1841 a_55268_n79536# GND 1.17f
C1842 a_53630_n79596# GND 2.61f
C1843 frontAnalog_v0p0p1_14.x65.A GND 2.63f
C1844 frontAnalog_v0p0p1_14.x63.A GND 2.46f
C1845 a_59577_n73683# GND 0.561f
C1846 a_57123_n74279# GND 0.319f
C1847 frontAnalog_v0p0p1_12.RSfetsym_0.x2.Y GND 1.53f
C1848 frontAnalog_v0p0p1_12.x63.X GND 5.15f
C1849 a_59578_n73170# GND 0.555f
C1850 frontAnalog_v0p0p1_12.RSfetsym_0.x1.Y GND 1.93f
C1851 frontAnalog_v0p0p1_12.RSfetsym_0.QN GND 3.84f
C1852 frontAnalog_v0p0p1_12.x65.X GND 5.07f
C1853 a_57123_n72759# GND 0.318f
C1854 a_55268_n74136# GND 1.17f
C1855 a_53630_n74196# GND 2.61f
C1856 frontAnalog_v0p0p1_12.x65.A GND 2.64f
C1857 frontAnalog_v0p0p1_12.x63.A GND 2.46f
C1858 a_59577_n68283# GND 0.561f
C1859 a_57123_n68879# GND 0.319f
C1860 frontAnalog_v0p0p1_13.RSfetsym_0.x2.Y GND 1.53f
C1861 frontAnalog_v0p0p1_13.x63.X GND 5.15f
C1862 a_59578_n67770# GND 0.555f
C1863 frontAnalog_v0p0p1_13.RSfetsym_0.x1.Y GND 1.93f
C1864 frontAnalog_v0p0p1_13.RSfetsym_0.QN GND 3.84f
C1865 frontAnalog_v0p0p1_13.x65.X GND 5.07f
C1866 a_57123_n67359# GND 0.318f
C1867 a_55268_n68736# GND 1.17f
C1868 a_53630_n68796# GND 2.61f
C1869 frontAnalog_v0p0p1_13.x65.A GND 2.64f
C1870 frontAnalog_v0p0p1_13.x63.A GND 2.46f
C1871 a_59577_n62883# GND 0.561f
C1872 a_57123_n63479# GND 0.319f
C1873 frontAnalog_v0p0p1_11.RSfetsym_0.x2.Y GND 1.53f
C1874 frontAnalog_v0p0p1_11.x63.X GND 5.15f
C1875 a_59578_n62370# GND 0.555f
C1876 frontAnalog_v0p0p1_11.RSfetsym_0.x1.Y GND 1.93f
C1877 frontAnalog_v0p0p1_11.RSfetsym_0.QN GND 3.84f
C1878 frontAnalog_v0p0p1_11.x65.X GND 5.07f
C1879 a_57123_n61959# GND 0.318f
C1880 a_55268_n63336# GND 1.17f
C1881 a_53630_n63396# GND 2.61f
C1882 frontAnalog_v0p0p1_11.x65.A GND 2.64f
C1883 frontAnalog_v0p0p1_11.x63.A GND 2.46f
C1884 a_59577_n57483# GND 0.561f
C1885 a_57123_n58079# GND 0.319f
C1886 frontAnalog_v0p0p1_10.RSfetsym_0.x2.Y GND 1.53f
C1887 frontAnalog_v0p0p1_10.x63.X GND 5.15f
C1888 a_59578_n56970# GND 0.555f
C1889 frontAnalog_v0p0p1_10.RSfetsym_0.x1.Y GND 1.93f
C1890 frontAnalog_v0p0p1_10.RSfetsym_0.QN GND 3.84f
C1891 frontAnalog_v0p0p1_10.x65.X GND 5.07f
C1892 a_57123_n56559# GND 0.318f
C1893 a_55268_n57936# GND 1.17f
C1894 a_53630_n57996# GND 2.61f
C1895 frontAnalog_v0p0p1_10.x65.A GND 2.64f
C1896 frontAnalog_v0p0p1_10.x63.A GND 2.46f
C1897 resistorDivider_v0p0p1_0.V1 GND 72.9f
C1898 16to4_PriorityEncoder_v0p0p1_0.x3.x22.B GND 0.245f
C1899 16to4_PriorityEncoder_v0p0p1_0.x3.x22.D GND 0.69f
C1900 resistorDivider_v0p0p1_0.V2 GND 83f
C1901 a_78525_n53555# GND 0.366f
C1902 a_78097_n53777# GND 0.22f
C1903 a_77605_n53805# GND 0.296f
C1904 16to4_PriorityEncoder_v0p0p1_0.x3.x22.C GND 0.443f
C1905 a_77605_n52819# GND 0.295f
C1906 16to4_PriorityEncoder_v0p0p1_0.x3.x21.B GND 0.662f
C1907 a_77605_n52567# GND 0.295f
C1908 a_59577_n52083# GND 0.561f
C1909 16to4_PriorityEncoder_v0p0p1_0.x3.A0 GND 7.55f
C1910 a_57123_n52679# GND 0.319f
C1911 frontAnalog_v0p0p1_9.RSfetsym_0.x2.Y GND 1.53f
C1912 frontAnalog_v0p0p1_9.x63.X GND 5.15f
C1913 a_77605_n51585# GND 0.297f
C1914 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND 9.85f
C1915 16to4_PriorityEncoder_v0p0p1_0.x22.A GND 2.13f
C1916 16to4_PriorityEncoder_v0p0p1_0.x21.A GND 0.663f
C1917 16to4_PriorityEncoder_v0p0p1_0.x2.X GND 0.382f
C1918 a_82906_n51645# GND 0.263f
C1919 a_59578_n51570# GND 0.555f
C1920 16to4_PriorityEncoder_v0p0p1_0.x3.x17.D GND 0.871f
C1921 16to4_PriorityEncoder_v0p0p1_0.x3.x17.C GND 0.334f
C1922 frontAnalog_v0p0p1_9.RSfetsym_0.x1.Y GND 1.93f
C1923 a_78349_n51085# GND 0.369f
C1924 a_77605_n51335# GND 0.296f
C1925 frontAnalog_v0p0p1_9.RSfetsym_0.QN GND 3.84f
C1926 frontAnalog_v0p0p1_9.x65.X GND 5.07f
C1927 a_57123_n51159# GND 0.318f
C1928 a_55268_n52536# GND 1.17f
C1929 a_53630_n52596# GND 2.61f
C1930 resistorDivider_v0p0p1_0.V3 GND 78.4f
C1931 a_77639_n50381# GND 0.286f
C1932 frontAnalog_v0p0p1_9.x65.A GND 2.64f
C1933 frontAnalog_v0p0p1_9.x63.A GND 2.46f
C1934 resistorDivider_v0p0p1_0.V4 GND 74.3f
C1935 a_77637_n50057# GND 0.288f
C1936 a_78065_n49349# GND 0.367f
C1937 16to4_PriorityEncoder_v0p0p1_0.x3.x17.A GND 0.917f
C1938 16to4_PriorityEncoder_v0p0p1_0.x3.x22.A GND 2.02f
C1939 16to4_PriorityEncoder_v0p0p1_0.x3.x14.B GND 0.263f
C1940 a_77637_n49127# GND 0.28f
C1941 16to4_PriorityEncoder_v0p0p1_0.x3.x14.A GND 0.978f
C1942 resistorDivider_v0p0p1_0.V5 GND 73.2f
C1943 a_77637_n48817# GND 0.289f
C1944 16to4_PriorityEncoder_v0p0p1_0.x3.A1 GND 5.12f
C1945 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND 9.86f
C1946 16to4_PriorityEncoder_v0p0p1_0.x29.A GND 2.13f
C1947 16to4_PriorityEncoder_v0p0p1_0.x28.A GND 0.665f
C1948 16to4_PriorityEncoder_v0p0p1_0.x1.X GND 0.383f
C1949 a_82906_n47995# GND 0.265f
C1950 a_77605_n48109# GND 0.388f
C1951 16to4_PriorityEncoder_v0p0p1_0.x3.GS GND 2.06f
C1952 16to4_PriorityEncoder_v0p0p1_0.x3.EO GND 2.32f
C1953 16to4_PriorityEncoder_v0p0p1_0.x3.x4.C GND 0.676f
C1954 16to4_PriorityEncoder_v0p0p1_0.x3.x4.B GND 0.162f
C1955 a_78649_n47567# GND 0.258f
C1956 a_78159_n47589# GND 0.343f
C1957 a_77605_n47345# GND 0.379f
C1958 16to4_PriorityEncoder_v0p0p1_0.x3.x9.Y GND 1.07f
C1959 16to4_PriorityEncoder_v0p0p1_0.x3.x20.B GND 4.1f
C1960 16to4_PriorityEncoder_v0p0p1_0.x3.x16.C GND 1.84f
C1961 16to4_PriorityEncoder_v0p0p1_0.x3.x19.C GND 4.41f
C1962 16to4_PriorityEncoder_v0p0p1_0.x3.x18.C GND 1.88f
C1963 a_59577_n46683# GND 0.561f
C1964 a_57123_n47279# GND 0.319f
C1965 frontAnalog_v0p0p1_8.RSfetsym_0.x2.Y GND 1.53f
C1966 frontAnalog_v0p0p1_8.x63.X GND 5.15f
C1967 a_59578_n46170# GND 0.555f
C1968 16to4_PriorityEncoder_v0p0p1_0.x2.A GND 6.65f
C1969 16to4_PriorityEncoder_v0p0p1_0.x5.x22.B GND 0.242f
C1970 16to4_PriorityEncoder_v0p0p1_0.x5.x22.D GND 0.684f
C1971 frontAnalog_v0p0p1_8.RSfetsym_0.x1.Y GND 1.93f
C1972 a_78525_n45515# GND 0.364f
C1973 a_78097_n45737# GND 0.217f
C1974 a_77605_n45765# GND 0.291f
C1975 frontAnalog_v0p0p1_8.RSfetsym_0.QN GND 3.81f
C1976 frontAnalog_v0p0p1_8.x65.X GND 5.03f
C1977 a_57123_n45759# GND 0.318f
C1978 a_55268_n47136# GND 1.17f
C1979 a_53630_n47196# GND 2.61f
C1980 resistorDivider_v0p0p1_0.V6 GND 71.3f
C1981 resistorDivider_v0p0p1_0.V7 GND 68.6f
C1982 16to4_PriorityEncoder_v0p0p1_0.x5.x22.C GND 0.434f
C1983 frontAnalog_v0p0p1_8.x65.A GND 2.64f
C1984 frontAnalog_v0p0p1_8.x63.A GND 2.46f
C1985 a_77605_n44779# GND 0.293f
C1986 16to4_PriorityEncoder_v0p0p1_0.x5.x21.B GND 0.652f
C1987 a_77605_n44527# GND 0.295f
C1988 16to4_PriorityEncoder_v0p0p1_0.x3.A2 GND 7.64f
C1989 resistorDivider_v0p0p1_0.V8 GND 65.6f
C1990 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND 9.83f
C1991 16to4_PriorityEncoder_v0p0p1_0.x36.A GND 2.12f
C1992 16to4_PriorityEncoder_v0p0p1_0.x35.A GND 0.662f
C1993 16to4_PriorityEncoder_v0p0p1_0.x34.A GND 0.379f
C1994 a_82906_n43855# GND 0.263f
C1995 a_77605_n43545# GND 0.297f
C1996 16to4_PriorityEncoder_v0p0p1_0.x1.A GND 5.67f
C1997 16to4_PriorityEncoder_v0p0p1_0.x5.x17.D GND 0.871f
C1998 16to4_PriorityEncoder_v0p0p1_0.x5.x17.C GND 0.334f
C1999 a_78349_n43045# GND 0.369f
C2000 a_77605_n43295# GND 0.296f
C2001 a_77639_n42341# GND 0.286f
C2002 a_77637_n42017# GND 0.288f
C2003 16to4_PriorityEncoder_v0p0p1_0.x5.A2 GND 5.29f
C2004 a_78065_n41309# GND 0.367f
C2005 16to4_PriorityEncoder_v0p0p1_0.x5.x17.A GND 0.876f
C2006 16to4_PriorityEncoder_v0p0p1_0.x5.x22.A GND 1.77f
C2007 16to4_PriorityEncoder_v0p0p1_0.x5.x14.B GND 0.263f
C2008 a_77637_n41087# GND 0.28f
C2009 a_59577_n41283# GND 0.561f
C2010 a_57123_n41879# GND 0.319f
C2011 frontAnalog_v0p0p1_1.RSfetsym_0.x2.Y GND 1.51f
C2012 frontAnalog_v0p0p1_1.x63.X GND 5.14f
C2013 16to4_PriorityEncoder_v0p0p1_0.x5.x14.A GND 0.958f
C2014 a_59578_n40770# GND 0.555f
C2015 a_77637_n40777# GND 0.289f
C2016 frontAnalog_v0p0p1_1.RSfetsym_0.x1.Y GND 1.92f
C2017 resistorDivider_v0p0p1_0.V9 GND 62.3f
C2018 16to4_PriorityEncoder_v0p0p1_0.x3.EI GND 18.6f
C2019 frontAnalog_v0p0p1_1.RSfetsym_0.QN GND 3.91f
C2020 a_77605_n40069# GND 0.391f
C2021 frontAnalog_v0p0p1_1.x65.X GND 5f
C2022 a_57123_n40359# GND 0.318f
C2023 a_55268_n41736# GND 1.17f
C2024 a_53630_n41796# GND 2.61f
C2025 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND 9.88f
C2026 16to4_PriorityEncoder_v0p0p1_0.x43.A GND 2.02f
C2027 16to4_PriorityEncoder_v0p0p1_0.x42.A GND 0.633f
C2028 16to4_PriorityEncoder_v0p0p1_0.x5.GS GND 2.51f
C2029 frontAnalog_v0p0p1_1.x65.A GND 2.64f
C2030 frontAnalog_v0p0p1_1.x63.A GND 2.46f
C2031 16to4_PriorityEncoder_v0p0p1_0.x5.EO GND 2.62f
C2032 16to4_PriorityEncoder_v0p0p1_0.x5.x4.C GND 0.684f
C2033 16to4_PriorityEncoder_v0p0p1_0.x5.x4.B GND 0.167f
C2034 a_78649_n39527# GND 0.262f
C2035 a_78159_n39549# GND 0.347f
C2036 a_77605_n39305# GND 0.384f
C2037 16to4_PriorityEncoder_v0p0p1_0.x5.x9.Y GND 1.5f
C2038 16to4_PriorityEncoder_v0p0p1_0.x5.x20.B GND 4.1f
C2039 16to4_PriorityEncoder_v0p0p1_0.x5.x16.C GND 1.85f
C2040 16to4_PriorityEncoder_v0p0p1_0.x5.x19.C GND 4.42f
C2041 16to4_PriorityEncoder_v0p0p1_0.x5.x18.C GND 1.89f
C2042 a_59577_n35883# GND 0.561f
C2043 a_57123_n36479# GND 0.319f
C2044 frontAnalog_v0p0p1_7.RSfetsym_0.x2.Y GND 1.53f
C2045 frontAnalog_v0p0p1_7.x63.X GND 5.23f
C2046 a_59578_n35370# GND 0.555f
C2047 frontAnalog_v0p0p1_7.RSfetsym_0.x1.Y GND 1.93f
C2048 resistorDivider_v0p0p1_0.V10 GND 65.4f
C2049 frontAnalog_v0p0p1_7.RSfetsym_0.QN GND 3.91f
C2050 frontAnalog_v0p0p1_7.x65.X GND 5.07f
C2051 a_57123_n34959# GND 0.318f
C2052 a_55268_n36336# GND 1.17f
C2053 a_53630_n36396# GND 2.61f
C2054 frontAnalog_v0p0p1_7.x65.A GND 2.64f
C2055 frontAnalog_v0p0p1_7.x63.A GND 2.46f
C2056 a_59577_n30483# GND 0.561f
C2057 a_57123_n31079# GND 0.319f
C2058 frontAnalog_v0p0p1_6.RSfetsym_0.x2.Y GND 1.53f
C2059 frontAnalog_v0p0p1_6.x63.X GND 5.17f
C2060 a_59578_n29970# GND 0.555f
C2061 frontAnalog_v0p0p1_6.RSfetsym_0.x1.Y GND 1.93f
C2062 resistorDivider_v0p0p1_0.V11 GND 69.9f
C2063 frontAnalog_v0p0p1_6.RSfetsym_0.QN GND 3.84f
C2064 frontAnalog_v0p0p1_6.x65.X GND 5.07f
C2065 a_57123_n29559# GND 0.318f
C2066 a_55268_n30936# GND 1.17f
C2067 a_53630_n30996# GND 2.61f
C2068 frontAnalog_v0p0p1_6.x65.A GND 2.63f
C2069 frontAnalog_v0p0p1_6.x63.A GND 2.46f
C2070 a_59577_n25083# GND 0.561f
C2071 a_57123_n25679# GND 0.319f
C2072 frontAnalog_v0p0p1_5.RSfetsym_0.x2.Y GND 1.53f
C2073 frontAnalog_v0p0p1_5.x63.X GND 5.13f
C2074 a_59578_n24570# GND 0.555f
C2075 frontAnalog_v0p0p1_5.RSfetsym_0.x1.Y GND 1.93f
C2076 16to4_PriorityEncoder_v0p0p1_0.I11 GND 24.7f
C2077 resistorDivider_v0p0p1_0.V12 GND 74.9f
C2078 frontAnalog_v0p0p1_5.RSfetsym_0.QN GND 3.91f
C2079 frontAnalog_v0p0p1_5.x65.X GND 5.07f
C2080 a_57123_n24159# GND 0.318f
C2081 a_55268_n25536# GND 1.17f
C2082 a_53630_n25596# GND 2.61f
C2083 frontAnalog_v0p0p1_5.x65.A GND 2.64f
C2084 frontAnalog_v0p0p1_5.x63.A GND 2.46f
C2085 a_59577_n19683# GND 0.561f
C2086 a_57123_n20279# GND 0.319f
C2087 frontAnalog_v0p0p1_4.RSfetsym_0.x2.Y GND 1.53f
C2088 frontAnalog_v0p0p1_4.x63.X GND 5.17f
C2089 a_59578_n19170# GND 0.555f
C2090 frontAnalog_v0p0p1_4.RSfetsym_0.x1.Y GND 1.93f
C2091 16to4_PriorityEncoder_v0p0p1_0.I12 GND 25.3f
C2092 resistorDivider_v0p0p1_0.V13 GND 76.5f
C2093 frontAnalog_v0p0p1_4.RSfetsym_0.QN GND 3.91f
C2094 frontAnalog_v0p0p1_4.x65.X GND 5.07f
C2095 a_57123_n18759# GND 0.318f
C2096 a_55268_n20136# GND 1.17f
C2097 a_53630_n20196# GND 2.61f
C2098 frontAnalog_v0p0p1_4.x65.A GND 2.63f
C2099 frontAnalog_v0p0p1_4.x63.A GND 2.46f
C2100 a_59577_n14283# GND 0.561f
C2101 a_57123_n14879# GND 0.319f
C2102 frontAnalog_v0p0p1_3.RSfetsym_0.x2.Y GND 1.53f
C2103 frontAnalog_v0p0p1_3.x63.X GND 5.17f
C2104 a_59578_n13770# GND 0.555f
C2105 frontAnalog_v0p0p1_3.RSfetsym_0.x1.Y GND 1.93f
C2106 16to4_PriorityEncoder_v0p0p1_0.I13 GND 30.8f
C2107 resistorDivider_v0p0p1_0.V14 GND 75.9f
C2108 frontAnalog_v0p0p1_3.RSfetsym_0.QN GND 3.84f
C2109 frontAnalog_v0p0p1_3.x65.X GND 5.07f
C2110 a_57123_n13359# GND 0.318f
C2111 a_55268_n14736# GND 1.17f
C2112 a_53630_n14796# GND 2.61f
C2113 frontAnalog_v0p0p1_3.x65.A GND 2.64f
C2114 frontAnalog_v0p0p1_3.x63.A GND 2.46f
C2115 a_59577_n8883# GND 0.561f
C2116 a_57123_n9479# GND 0.319f
C2117 frontAnalog_v0p0p1_0.RSfetsym_0.x2.Y GND 1.53f
C2118 frontAnalog_v0p0p1_0.x63.X GND 5.18f
C2119 a_59578_n8370# GND 0.555f
C2120 frontAnalog_v0p0p1_0.RSfetsym_0.x1.Y GND 1.93f
C2121 16to4_PriorityEncoder_v0p0p1_0.I14 GND 59.3f
C2122 resistorDivider_v0p0p1_0.V15 GND 76f
C2123 frontAnalog_v0p0p1_0.RSfetsym_0.QN GND 3.84f
C2124 frontAnalog_v0p0p1_0.x65.X GND 5.07f
C2125 a_57123_n7959# GND 0.318f
C2126 a_55268_n9336# GND 1.17f
C2127 a_53630_n9396# GND 2.61f
C2128 frontAnalog_v0p0p1_0.x65.A GND 2.64f
C2129 frontAnalog_v0p0p1_0.x63.A GND 2.46f
C2130 a_59577_n3483# GND 0.561f
C2131 a_57123_n4079# GND 0.319f
C2132 frontAnalog_v0p0p1_2.RSfetsym_0.x2.Y GND 1.53f
C2133 frontAnalog_v0p0p1_2.x63.X GND 5.18f
C2134 a_59578_n2970# GND 0.555f
C2135 frontAnalog_v0p0p1_2.RSfetsym_0.x1.Y GND 1.93f
C2136 16to4_PriorityEncoder_v0p0p1_0.I15 GND 66.8f
C2137 resistorDivider_v0p0p1_0.V16 GND 79.6f
C2138 frontAnalog_v0p0p1_2.RSfetsym_0.QN GND 3.91f
C2139 frontAnalog_v0p0p1_2.x65.X GND 5.07f
C2140 a_57123_n2559# GND 0.318f
C2141 a_55268_n3936# GND 1.17f
C2142 a_53630_n3996# GND 2.61f
C2143 frontAnalog_v0p0p1_10.IB GND 0.288p
C2144 frontAnalog_v0p0p1_2.x65.A GND 2.63f
C2145 frontAnalog_v0p0p1_2.x63.A GND 2.46f
C2146 w_55000_n84550# GND 2.69f
C2147 w_55000_n83928# GND 2.69f
C2148 w_55000_n79150# GND 2.69f
C2149 w_55000_n78528# GND 2.69f
C2150 w_55000_n73750# GND 2.69f
C2151 w_55000_n73128# GND 2.69f
C2152 w_55000_n68350# GND 2.69f
C2153 w_55000_n67728# GND 2.69f
C2154 w_55000_n62950# GND 2.69f
C2155 w_55000_n62328# GND 2.69f
C2156 w_55000_n57550# GND 2.69f
C2157 w_55000_n56928# GND 2.69f
C2158 w_55000_n52150# GND 2.69f
C2159 w_55000_n51528# GND 2.69f
C2160 w_55000_n46750# GND 2.69f
C2161 w_55000_n46128# GND 2.69f
C2162 w_55000_n41350# GND 2.69f
C2163 w_55000_n40728# GND 2.69f
C2164 w_55000_n35950# GND 2.69f
C2165 w_55000_n35328# GND 2.69f
C2166 w_55000_n30550# GND 2.69f
C2167 w_55000_n29928# GND 2.69f
C2168 w_55000_n25150# GND 2.69f
C2169 w_55000_n24528# GND 2.69f
C2170 w_55000_n19750# GND 2.69f
C2171 w_55000_n19128# GND 2.68f
C2172 w_55000_n14350# GND 2.69f
C2173 w_55000_n13728# GND 2.69f
C2174 w_55000_n8950# GND 2.69f
C2175 w_55000_n8328# GND 2.69f
C2176 w_55000_n3550# GND 2.69f
C2177 w_55000_n2928# GND 2.68f
C2178 frontAnalog_v0p0p1_0.x63.A.n0 GND 0.12f
C2179 frontAnalog_v0p0p1_0.x63.A.n1 GND 2.22f
C2180 frontAnalog_v0p0p1_0.x63.A.t6 GND 0.014f
C2181 frontAnalog_v0p0p1_0.x63.A.t5 GND 0.0225f
C2182 frontAnalog_v0p0p1_0.x63.A.n2 GND 0.0465f
C2183 frontAnalog_v0p0p1_0.x63.A.t1 GND 0.151f
C2184 frontAnalog_v0p0p1_0.x63.A.t2 GND 0.0156f
C2185 frontAnalog_v0p0p1_0.x63.A.t3 GND 0.335f
C2186 frontAnalog_v0p0p1_0.x63.A.t4 GND 0.0256f
C2187 frontAnalog_v0p0p1_0.x63.A.t0 GND 0.173f
C2188 frontAnalog_v0p0p1_0.x63.A.t7 GND 0.175f
C2189 frontAnalog_v0p0p1_0.x63.A.n3 GND 1f
C2190 frontAnalog_v0p0p1_0.x63.A.n4 GND 0.953f
C2191 frontAnalog_v0p0p1_0.x63.A.n5 GND 1.25f
C2192 frontAnalog_v0p0p1_0.x65.A.n0 GND 0.139f
C2193 frontAnalog_v0p0p1_0.x65.A.t5 GND 0.028f
C2194 frontAnalog_v0p0p1_0.x65.A.t6 GND 0.0175f
C2195 frontAnalog_v0p0p1_0.x65.A.n1 GND 0.0568f
C2196 frontAnalog_v0p0p1_0.x65.A.t1 GND 0.149f
C2197 frontAnalog_v0p0p1_0.x65.A.t2 GND 0.463f
C2198 frontAnalog_v0p0p1_0.x65.A.t3 GND 0.0194f
C2199 frontAnalog_v0p0p1_0.x65.A.n2 GND 1.6f
C2200 frontAnalog_v0p0p1_0.x65.A.t7 GND 0.0318f
C2201 frontAnalog_v0p0p1_0.x65.A.t0 GND 0.141f
C2202 frontAnalog_v0p0p1_0.x65.A.t4 GND 0.219f
C2203 frontAnalog_v0p0p1_0.x65.A.n3 GND 1.37f
C2204 frontAnalog_v0p0p1_0.x65.A.n4 GND 0.898f
C2205 frontAnalog_v0p0p1_0.x65.A.n5 GND 2.01f
C2206 frontAnalog_v0p0p1_0.x65.A.n6 GND 1.72f
C2207 frontAnalog_v0p0p1_6.x65.A.n0 GND 0.139f
C2208 frontAnalog_v0p0p1_6.x65.A.t6 GND 0.028f
C2209 frontAnalog_v0p0p1_6.x65.A.t7 GND 0.0175f
C2210 frontAnalog_v0p0p1_6.x65.A.n1 GND 0.0568f
C2211 frontAnalog_v0p0p1_6.x65.A.t1 GND 0.149f
C2212 frontAnalog_v0p0p1_6.x65.A.t2 GND 0.463f
C2213 frontAnalog_v0p0p1_6.x65.A.t3 GND 0.0194f
C2214 frontAnalog_v0p0p1_6.x65.A.n2 GND 1.6f
C2215 frontAnalog_v0p0p1_6.x65.A.t5 GND 0.0318f
C2216 frontAnalog_v0p0p1_6.x65.A.t0 GND 0.141f
C2217 frontAnalog_v0p0p1_6.x65.A.t4 GND 0.219f
C2218 frontAnalog_v0p0p1_6.x65.A.n3 GND 1.37f
C2219 frontAnalog_v0p0p1_6.x65.A.n4 GND 0.898f
C2220 frontAnalog_v0p0p1_6.x65.A.n5 GND 2.01f
C2221 frontAnalog_v0p0p1_6.x65.A.n6 GND 1.72f
C2222 frontAnalog_v0p0p1_12.x65.A.n0 GND 0.139f
C2223 frontAnalog_v0p0p1_12.x65.A.t4 GND 0.028f
C2224 frontAnalog_v0p0p1_12.x65.A.t6 GND 0.0175f
C2225 frontAnalog_v0p0p1_12.x65.A.n1 GND 0.0568f
C2226 frontAnalog_v0p0p1_12.x65.A.t1 GND 0.149f
C2227 frontAnalog_v0p0p1_12.x65.A.t3 GND 0.463f
C2228 frontAnalog_v0p0p1_12.x65.A.t2 GND 0.0194f
C2229 frontAnalog_v0p0p1_12.x65.A.n2 GND 1.6f
C2230 frontAnalog_v0p0p1_12.x65.A.t7 GND 0.0318f
C2231 frontAnalog_v0p0p1_12.x65.A.t0 GND 0.141f
C2232 frontAnalog_v0p0p1_12.x65.A.t5 GND 0.219f
C2233 frontAnalog_v0p0p1_12.x65.A.n3 GND 1.37f
C2234 frontAnalog_v0p0p1_12.x65.A.n4 GND 0.898f
C2235 frontAnalog_v0p0p1_12.x65.A.n5 GND 2.01f
C2236 frontAnalog_v0p0p1_12.x65.A.n6 GND 1.72f
C2237 frontAnalog_v0p0p1_2.RSfetsym_0.QN.t2 GND 0.0322f
C2238 frontAnalog_v0p0p1_2.RSfetsym_0.QN.t3 GND 0.0322f
C2239 frontAnalog_v0p0p1_2.RSfetsym_0.QN.n0 GND 0.136f
C2240 frontAnalog_v0p0p1_2.RSfetsym_0.QN.t5 GND 0.0321f
C2241 frontAnalog_v0p0p1_2.RSfetsym_0.QN.t6 GND 0.0947f
C2242 frontAnalog_v0p0p1_2.RSfetsym_0.QN.n1 GND 1.46f
C2243 frontAnalog_v0p0p1_2.RSfetsym_0.QN.n2 GND 0.0784f
C2244 frontAnalog_v0p0p1_2.RSfetsym_0.QN.n3 GND 0.102f
C2245 frontAnalog_v0p0p1_2.RSfetsym_0.QN.n4 GND 0.445f
C2246 frontAnalog_v0p0p1_2.RSfetsym_0.QN.n5 GND 0.0126f
C2247 frontAnalog_v0p0p1_2.RSfetsym_0.QN.n6 GND 0.0341f
C2248 frontAnalog_v0p0p1_2.RSfetsym_0.QN.t1 GND 0.0322f
C2249 frontAnalog_v0p0p1_2.RSfetsym_0.QN.n7 GND 0.107f
C2250 frontAnalog_v0p0p1_2.RSfetsym_0.QN.n8 GND 0.131f
C2251 frontAnalog_v0p0p1_2.RSfetsym_0.QN.n9 GND 0.351f
C2252 frontAnalog_v0p0p1_2.RSfetsym_0.QN.n10 GND 0.871f
C2253 frontAnalog_v0p0p1_2.RSfetsym_0.QN.t0 GND 0.0566f
C2254 frontAnalog_v0p0p1_2.RSfetsym_0.QN.n11 GND 2.48f
C2255 frontAnalog_v0p0p1_8.x63.A.n0 GND 0.12f
C2256 frontAnalog_v0p0p1_8.x63.A.n1 GND 2.22f
C2257 frontAnalog_v0p0p1_8.x63.A.t7 GND 0.014f
C2258 frontAnalog_v0p0p1_8.x63.A.t5 GND 0.0225f
C2259 frontAnalog_v0p0p1_8.x63.A.n2 GND 0.0465f
C2260 frontAnalog_v0p0p1_8.x63.A.t6 GND 0.0256f
C2261 frontAnalog_v0p0p1_8.x63.A.t1 GND 0.173f
C2262 frontAnalog_v0p0p1_8.x63.A.t4 GND 0.175f
C2263 frontAnalog_v0p0p1_8.x63.A.n3 GND 1f
C2264 frontAnalog_v0p0p1_8.x63.A.n4 GND 0.953f
C2265 frontAnalog_v0p0p1_8.x63.A.t2 GND 0.0156f
C2266 frontAnalog_v0p0p1_8.x63.A.t3 GND 0.335f
C2267 frontAnalog_v0p0p1_8.x63.A.t0 GND 0.151f
C2268 frontAnalog_v0p0p1_8.x63.A.n5 GND 1.25f
C2269 16to4_PriorityEncoder_v0p0p1_0.I11.t8 GND 0.0238f
C2270 16to4_PriorityEncoder_v0p0p1_0.I11.n0 GND 0.373f
C2271 16to4_PriorityEncoder_v0p0p1_0.I11.n1 GND 0.112f
C2272 16to4_PriorityEncoder_v0p0p1_0.I11.n2 GND 0.0495f
C2273 16to4_PriorityEncoder_v0p0p1_0.I11.n3 GND 0.0744f
C2274 16to4_PriorityEncoder_v0p0p1_0.I11.n4 GND 0.0795f
C2275 16to4_PriorityEncoder_v0p0p1_0.I11.n5 GND 0.11f
C2276 16to4_PriorityEncoder_v0p0p1_0.I11.n6 GND 0.104f
C2277 16to4_PriorityEncoder_v0p0p1_0.I11.n7 GND 0.25f
C2278 16to4_PriorityEncoder_v0p0p1_0.I11.n8 GND 0.0104f
C2279 16to4_PriorityEncoder_v0p0p1_0.I11.n10 GND 0.656f
C2280 16to4_PriorityEncoder_v0p0p1_0.I11.n11 GND 0.0139f
C2281 16to4_PriorityEncoder_v0p0p1_0.I11.n12 GND 0.0107f
C2282 16to4_PriorityEncoder_v0p0p1_0.I11.n13 GND 1.18f
C2283 16to4_PriorityEncoder_v0p0p1_0.I11.n14 GND 0.552f
C2284 16to4_PriorityEncoder_v0p0p1_0.I11.n15 GND 6f
C2285 16to4_PriorityEncoder_v0p0p1_0.I11.n16 GND 13.9f
C2286 frontAnalog_v0p0p1_1.RSfetsym_0.QN.t3 GND 0.0322f
C2287 frontAnalog_v0p0p1_1.RSfetsym_0.QN.t2 GND 0.0322f
C2288 frontAnalog_v0p0p1_1.RSfetsym_0.QN.n0 GND 0.136f
C2289 frontAnalog_v0p0p1_1.RSfetsym_0.QN.t6 GND 0.0321f
C2290 frontAnalog_v0p0p1_1.RSfetsym_0.QN.t5 GND 0.0947f
C2291 frontAnalog_v0p0p1_1.RSfetsym_0.QN.n1 GND 1.46f
C2292 frontAnalog_v0p0p1_1.RSfetsym_0.QN.n2 GND 0.0784f
C2293 frontAnalog_v0p0p1_1.RSfetsym_0.QN.n3 GND 0.102f
C2294 frontAnalog_v0p0p1_1.RSfetsym_0.QN.n4 GND 0.445f
C2295 frontAnalog_v0p0p1_1.RSfetsym_0.QN.n5 GND 0.0126f
C2296 frontAnalog_v0p0p1_1.RSfetsym_0.QN.n6 GND 0.0341f
C2297 frontAnalog_v0p0p1_1.RSfetsym_0.QN.t4 GND 0.0322f
C2298 frontAnalog_v0p0p1_1.RSfetsym_0.QN.n7 GND 0.107f
C2299 frontAnalog_v0p0p1_1.RSfetsym_0.QN.n8 GND 0.131f
C2300 frontAnalog_v0p0p1_1.RSfetsym_0.QN.n9 GND 0.351f
C2301 frontAnalog_v0p0p1_1.RSfetsym_0.QN.n10 GND 0.871f
C2302 frontAnalog_v0p0p1_1.RSfetsym_0.QN.t0 GND 0.0566f
C2303 frontAnalog_v0p0p1_1.RSfetsym_0.QN.n11 GND 2.48f
C2304 frontAnalog_v0p0p1_13.Q.n2 GND 0.415f
C2305 frontAnalog_v0p0p1_13.Q.n5 GND 0.725f
C2306 frontAnalog_v0p0p1_13.Q.n6 GND 0.341f
C2307 frontAnalog_v0p0p1_13.Q.n7 GND 6.16f
C2308 frontAnalog_v0p0p1_13.Q.t8 GND 0.0148f
C2309 frontAnalog_v0p0p1_13.Q.n8 GND 0.232f
C2310 frontAnalog_v0p0p1_13.Q.n9 GND 0.0697f
C2311 frontAnalog_v0p0p1_13.Q.n10 GND 0.0307f
C2312 frontAnalog_v0p0p1_13.Q.n11 GND 0.0462f
C2313 frontAnalog_v0p0p1_13.Q.n12 GND 0.0494f
C2314 frontAnalog_v0p0p1_13.Q.n13 GND 0.0681f
C2315 frontAnalog_v0p0p1_13.Q.n14 GND 0.0644f
C2316 frontAnalog_v0p0p1_13.Q.n15 GND 0.148f
C2317 frontAnalog_v0p0p1_13.Q.n16 GND 9.39f
C2318 16to4_PriorityEncoder_v0p0p1_0.I15.n0 GND 0.14f
C2319 16to4_PriorityEncoder_v0p0p1_0.I15.n1 GND 0.0419f
C2320 16to4_PriorityEncoder_v0p0p1_0.I15.n2 GND 0.0185f
C2321 16to4_PriorityEncoder_v0p0p1_0.I15.n3 GND 0.0278f
C2322 16to4_PriorityEncoder_v0p0p1_0.I15.n4 GND 0.0297f
C2323 16to4_PriorityEncoder_v0p0p1_0.I15.n5 GND 0.041f
C2324 16to4_PriorityEncoder_v0p0p1_0.I15.n6 GND 0.0388f
C2325 16to4_PriorityEncoder_v0p0p1_0.I15.n7 GND 0.101f
C2326 16to4_PriorityEncoder_v0p0p1_0.I15.n16 GND 0.145f
C2327 16to4_PriorityEncoder_v0p0p1_0.I15.n17 GND 0.314f
C2328 16to4_PriorityEncoder_v0p0p1_0.I15.n18 GND 0.134f
C2329 16to4_PriorityEncoder_v0p0p1_0.I15.n19 GND 6.69f
C2330 16to4_PriorityEncoder_v0p0p1_0.I14.t8 GND 0.0161f
C2331 16to4_PriorityEncoder_v0p0p1_0.I14.n0 GND 0.253f
C2332 16to4_PriorityEncoder_v0p0p1_0.I14.n1 GND 0.076f
C2333 16to4_PriorityEncoder_v0p0p1_0.I14.n2 GND 0.0335f
C2334 16to4_PriorityEncoder_v0p0p1_0.I14.n3 GND 0.0504f
C2335 16to4_PriorityEncoder_v0p0p1_0.I14.n4 GND 0.0539f
C2336 16to4_PriorityEncoder_v0p0p1_0.I14.n5 GND 0.0742f
C2337 16to4_PriorityEncoder_v0p0p1_0.I14.n6 GND 0.0703f
C2338 16to4_PriorityEncoder_v0p0p1_0.I14.n7 GND 0.184f
C2339 16to4_PriorityEncoder_v0p0p1_0.I14.n18 GND 0.0698f
C2340 16to4_PriorityEncoder_v0p0p1_0.I14.n19 GND 0.169f
C2341 16to4_PriorityEncoder_v0p0p1_0.I14.n22 GND 0.0912f
C2342 16to4_PriorityEncoder_v0p0p1_0.I14.n29 GND 0.219f
C2343 16to4_PriorityEncoder_v0p0p1_0.I14.n30 GND 0.364f
C2344 16to4_PriorityEncoder_v0p0p1_0.I14.n31 GND 0.226f
C2345 16to4_PriorityEncoder_v0p0p1_0.I14.n32 GND 9.99f
C2346 frontAnalog_v0p0p1_8.x65.A.n0 GND 0.139f
C2347 frontAnalog_v0p0p1_8.x65.A.t4 GND 0.028f
C2348 frontAnalog_v0p0p1_8.x65.A.t6 GND 0.0175f
C2349 frontAnalog_v0p0p1_8.x65.A.n1 GND 0.0568f
C2350 frontAnalog_v0p0p1_8.x65.A.t2 GND 0.149f
C2351 frontAnalog_v0p0p1_8.x65.A.t7 GND 0.0318f
C2352 frontAnalog_v0p0p1_8.x65.A.t3 GND 0.141f
C2353 frontAnalog_v0p0p1_8.x65.A.t5 GND 0.219f
C2354 frontAnalog_v0p0p1_8.x65.A.n2 GND 1.37f
C2355 frontAnalog_v0p0p1_8.x65.A.n3 GND 0.898f
C2356 frontAnalog_v0p0p1_8.x65.A.t1 GND 0.463f
C2357 frontAnalog_v0p0p1_8.x65.A.t0 GND 0.0194f
C2358 frontAnalog_v0p0p1_8.x65.A.n4 GND 1.6f
C2359 frontAnalog_v0p0p1_8.x65.A.n5 GND 2.01f
C2360 frontAnalog_v0p0p1_8.x65.A.n6 GND 1.72f
C2361 frontAnalog_v0p0p1_11.x63.A.n0 GND 0.12f
C2362 frontAnalog_v0p0p1_11.x63.A.n1 GND 2.22f
C2363 frontAnalog_v0p0p1_11.x63.A.t7 GND 0.014f
C2364 frontAnalog_v0p0p1_11.x63.A.t5 GND 0.0225f
C2365 frontAnalog_v0p0p1_11.x63.A.n2 GND 0.0465f
C2366 frontAnalog_v0p0p1_11.x63.A.t1 GND 0.151f
C2367 frontAnalog_v0p0p1_11.x63.A.t2 GND 0.0156f
C2368 frontAnalog_v0p0p1_11.x63.A.t3 GND 0.335f
C2369 frontAnalog_v0p0p1_11.x63.A.t6 GND 0.0256f
C2370 frontAnalog_v0p0p1_11.x63.A.t0 GND 0.173f
C2371 frontAnalog_v0p0p1_11.x63.A.t4 GND 0.175f
C2372 frontAnalog_v0p0p1_11.x63.A.n3 GND 1f
C2373 frontAnalog_v0p0p1_11.x63.A.n4 GND 0.953f
C2374 frontAnalog_v0p0p1_11.x63.A.n5 GND 1.25f
C2375 frontAnalog_v0p0p1_8.Q.n0 GND 0.0144f
C2376 frontAnalog_v0p0p1_8.Q.n3 GND 0.0134f
C2377 frontAnalog_v0p0p1_8.Q.n8 GND 0.524f
C2378 frontAnalog_v0p0p1_8.Q.n9 GND 1.12f
C2379 frontAnalog_v0p0p1_8.Q.n10 GND 0.477f
C2380 frontAnalog_v0p0p1_8.Q.n11 GND 4.5f
C2381 frontAnalog_v0p0p1_8.Q.t6 GND 0.0105f
C2382 frontAnalog_v0p0p1_8.Q.t9 GND 0.0322f
C2383 frontAnalog_v0p0p1_8.Q.n12 GND 0.505f
C2384 frontAnalog_v0p0p1_8.Q.n13 GND 0.152f
C2385 frontAnalog_v0p0p1_8.Q.n14 GND 0.0669f
C2386 frontAnalog_v0p0p1_8.Q.t0 GND 0.0108f
C2387 frontAnalog_v0p0p1_8.Q.n15 GND 0.101f
C2388 frontAnalog_v0p0p1_8.Q.n16 GND 0.108f
C2389 frontAnalog_v0p0p1_8.Q.t2 GND 0.0108f
C2390 frontAnalog_v0p0p1_8.Q.t1 GND 0.0108f
C2391 frontAnalog_v0p0p1_8.Q.n17 GND 0.148f
C2392 frontAnalog_v0p0p1_8.Q.n18 GND 0.14f
C2393 frontAnalog_v0p0p1_8.Q.t4 GND 0.0119f
C2394 frontAnalog_v0p0p1_8.Q.n19 GND 0.323f
C2395 frontAnalog_v0p0p1_8.Q.n20 GND 8.86f
C2396 frontAnalog_v0p0p1_4.RSfetsym_0.QN.t1 GND 0.0322f
C2397 frontAnalog_v0p0p1_4.RSfetsym_0.QN.t2 GND 0.0322f
C2398 frontAnalog_v0p0p1_4.RSfetsym_0.QN.n0 GND 0.136f
C2399 frontAnalog_v0p0p1_4.RSfetsym_0.QN.t6 GND 0.0321f
C2400 frontAnalog_v0p0p1_4.RSfetsym_0.QN.t5 GND 0.0947f
C2401 frontAnalog_v0p0p1_4.RSfetsym_0.QN.n1 GND 1.46f
C2402 frontAnalog_v0p0p1_4.RSfetsym_0.QN.n2 GND 0.0784f
C2403 frontAnalog_v0p0p1_4.RSfetsym_0.QN.n3 GND 0.102f
C2404 frontAnalog_v0p0p1_4.RSfetsym_0.QN.n4 GND 0.445f
C2405 frontAnalog_v0p0p1_4.RSfetsym_0.QN.n5 GND 0.0126f
C2406 frontAnalog_v0p0p1_4.RSfetsym_0.QN.n6 GND 0.0341f
C2407 frontAnalog_v0p0p1_4.RSfetsym_0.QN.t4 GND 0.0322f
C2408 frontAnalog_v0p0p1_4.RSfetsym_0.QN.n7 GND 0.107f
C2409 frontAnalog_v0p0p1_4.RSfetsym_0.QN.n8 GND 0.131f
C2410 frontAnalog_v0p0p1_4.RSfetsym_0.QN.n9 GND 0.351f
C2411 frontAnalog_v0p0p1_4.RSfetsym_0.QN.n10 GND 0.871f
C2412 frontAnalog_v0p0p1_4.RSfetsym_0.QN.t3 GND 0.0566f
C2413 frontAnalog_v0p0p1_4.RSfetsym_0.QN.n11 GND 2.48f
C2414 frontAnalog_v0p0p1_12.x63.A.n0 GND 0.12f
C2415 frontAnalog_v0p0p1_12.x63.A.n1 GND 2.22f
C2416 frontAnalog_v0p0p1_12.x63.A.t6 GND 0.014f
C2417 frontAnalog_v0p0p1_12.x63.A.t4 GND 0.0225f
C2418 frontAnalog_v0p0p1_12.x63.A.n2 GND 0.0465f
C2419 frontAnalog_v0p0p1_12.x63.A.t1 GND 0.151f
C2420 frontAnalog_v0p0p1_12.x63.A.t2 GND 0.0156f
C2421 frontAnalog_v0p0p1_12.x63.A.t3 GND 0.335f
C2422 frontAnalog_v0p0p1_12.x63.A.t5 GND 0.0256f
C2423 frontAnalog_v0p0p1_12.x63.A.t0 GND 0.173f
C2424 frontAnalog_v0p0p1_12.x63.A.t7 GND 0.175f
C2425 frontAnalog_v0p0p1_12.x63.A.n3 GND 1f
C2426 frontAnalog_v0p0p1_12.x63.A.n4 GND 0.953f
C2427 frontAnalog_v0p0p1_12.x63.A.n5 GND 1.25f
C2428 frontAnalog_v0p0p1_11.RSfetsym_0.QN.t2 GND 0.0322f
C2429 frontAnalog_v0p0p1_11.RSfetsym_0.QN.t3 GND 0.0322f
C2430 frontAnalog_v0p0p1_11.RSfetsym_0.QN.n0 GND 0.136f
C2431 frontAnalog_v0p0p1_11.RSfetsym_0.QN.t6 GND 0.0321f
C2432 frontAnalog_v0p0p1_11.RSfetsym_0.QN.t5 GND 0.0947f
C2433 frontAnalog_v0p0p1_11.RSfetsym_0.QN.n1 GND 1.46f
C2434 frontAnalog_v0p0p1_11.RSfetsym_0.QN.n2 GND 0.0784f
C2435 frontAnalog_v0p0p1_11.RSfetsym_0.QN.n3 GND 0.102f
C2436 frontAnalog_v0p0p1_11.RSfetsym_0.QN.n4 GND 0.445f
C2437 frontAnalog_v0p0p1_11.RSfetsym_0.QN.n5 GND 0.0126f
C2438 frontAnalog_v0p0p1_11.RSfetsym_0.QN.n6 GND 0.0341f
C2439 frontAnalog_v0p0p1_11.RSfetsym_0.QN.t4 GND 0.0322f
C2440 frontAnalog_v0p0p1_11.RSfetsym_0.QN.n7 GND 0.107f
C2441 frontAnalog_v0p0p1_11.RSfetsym_0.QN.n8 GND 0.131f
C2442 frontAnalog_v0p0p1_11.RSfetsym_0.QN.n9 GND 0.351f
C2443 frontAnalog_v0p0p1_11.RSfetsym_0.QN.n10 GND 0.871f
C2444 frontAnalog_v0p0p1_11.RSfetsym_0.QN.t0 GND 0.0566f
C2445 frontAnalog_v0p0p1_11.RSfetsym_0.QN.n11 GND 2.48f
C2446 frontAnalog_v0p0p1_13.x65.A.n0 GND 0.139f
C2447 frontAnalog_v0p0p1_13.x65.A.t4 GND 0.028f
C2448 frontAnalog_v0p0p1_13.x65.A.t6 GND 0.0175f
C2449 frontAnalog_v0p0p1_13.x65.A.n1 GND 0.0568f
C2450 frontAnalog_v0p0p1_13.x65.A.t1 GND 0.149f
C2451 frontAnalog_v0p0p1_13.x65.A.t3 GND 0.463f
C2452 frontAnalog_v0p0p1_13.x65.A.t2 GND 0.0194f
C2453 frontAnalog_v0p0p1_13.x65.A.n2 GND 1.6f
C2454 frontAnalog_v0p0p1_13.x65.A.t7 GND 0.0318f
C2455 frontAnalog_v0p0p1_13.x65.A.t0 GND 0.141f
C2456 frontAnalog_v0p0p1_13.x65.A.t5 GND 0.219f
C2457 frontAnalog_v0p0p1_13.x65.A.n3 GND 1.37f
C2458 frontAnalog_v0p0p1_13.x65.A.n4 GND 0.898f
C2459 frontAnalog_v0p0p1_13.x65.A.n5 GND 2.01f
C2460 frontAnalog_v0p0p1_13.x65.A.n6 GND 1.72f
C2461 frontAnalog_v0p0p1_1.Q.t5 GND 0.0145f
C2462 frontAnalog_v0p0p1_1.Q.n0 GND 0.228f
C2463 frontAnalog_v0p0p1_1.Q.n1 GND 0.0684f
C2464 frontAnalog_v0p0p1_1.Q.n2 GND 0.0302f
C2465 frontAnalog_v0p0p1_1.Q.n3 GND 0.0454f
C2466 frontAnalog_v0p0p1_1.Q.n4 GND 0.0485f
C2467 frontAnalog_v0p0p1_1.Q.n5 GND 0.0668f
C2468 frontAnalog_v0p0p1_1.Q.n6 GND 0.0632f
C2469 frontAnalog_v0p0p1_1.Q.n7 GND 0.165f
C2470 frontAnalog_v0p0p1_1.Q.n9 GND 0.148f
C2471 frontAnalog_v0p0p1_1.Q.n10 GND 0.382f
C2472 frontAnalog_v0p0p1_1.Q.n11 GND 6.35f
C2473 frontAnalog_v0p0p1_0.RSfetsym_0.QN.t3 GND 0.0322f
C2474 frontAnalog_v0p0p1_0.RSfetsym_0.QN.t2 GND 0.0322f
C2475 frontAnalog_v0p0p1_0.RSfetsym_0.QN.n0 GND 0.136f
C2476 frontAnalog_v0p0p1_0.RSfetsym_0.QN.t5 GND 0.0321f
C2477 frontAnalog_v0p0p1_0.RSfetsym_0.QN.t6 GND 0.0947f
C2478 frontAnalog_v0p0p1_0.RSfetsym_0.QN.n1 GND 1.46f
C2479 frontAnalog_v0p0p1_0.RSfetsym_0.QN.n2 GND 0.0784f
C2480 frontAnalog_v0p0p1_0.RSfetsym_0.QN.n3 GND 0.102f
C2481 frontAnalog_v0p0p1_0.RSfetsym_0.QN.n4 GND 0.445f
C2482 frontAnalog_v0p0p1_0.RSfetsym_0.QN.n5 GND 0.0126f
C2483 frontAnalog_v0p0p1_0.RSfetsym_0.QN.n6 GND 0.0341f
C2484 frontAnalog_v0p0p1_0.RSfetsym_0.QN.t0 GND 0.0322f
C2485 frontAnalog_v0p0p1_0.RSfetsym_0.QN.n7 GND 0.107f
C2486 frontAnalog_v0p0p1_0.RSfetsym_0.QN.n8 GND 0.131f
C2487 frontAnalog_v0p0p1_0.RSfetsym_0.QN.n9 GND 0.351f
C2488 frontAnalog_v0p0p1_0.RSfetsym_0.QN.n10 GND 0.871f
C2489 frontAnalog_v0p0p1_0.RSfetsym_0.QN.t4 GND 0.0566f
C2490 frontAnalog_v0p0p1_0.RSfetsym_0.QN.n11 GND 2.48f
C2491 frontAnalog_v0p0p1_7.RSfetsym_0.QN.t1 GND 0.0322f
C2492 frontAnalog_v0p0p1_7.RSfetsym_0.QN.t2 GND 0.0322f
C2493 frontAnalog_v0p0p1_7.RSfetsym_0.QN.n0 GND 0.136f
C2494 frontAnalog_v0p0p1_7.RSfetsym_0.QN.t6 GND 0.0321f
C2495 frontAnalog_v0p0p1_7.RSfetsym_0.QN.t5 GND 0.0947f
C2496 frontAnalog_v0p0p1_7.RSfetsym_0.QN.n1 GND 1.46f
C2497 frontAnalog_v0p0p1_7.RSfetsym_0.QN.n2 GND 0.0784f
C2498 frontAnalog_v0p0p1_7.RSfetsym_0.QN.n3 GND 0.102f
C2499 frontAnalog_v0p0p1_7.RSfetsym_0.QN.n4 GND 0.445f
C2500 frontAnalog_v0p0p1_7.RSfetsym_0.QN.n5 GND 0.0126f
C2501 frontAnalog_v0p0p1_7.RSfetsym_0.QN.n6 GND 0.0341f
C2502 frontAnalog_v0p0p1_7.RSfetsym_0.QN.t4 GND 0.0322f
C2503 frontAnalog_v0p0p1_7.RSfetsym_0.QN.n7 GND 0.107f
C2504 frontAnalog_v0p0p1_7.RSfetsym_0.QN.n8 GND 0.131f
C2505 frontAnalog_v0p0p1_7.RSfetsym_0.QN.n9 GND 0.351f
C2506 frontAnalog_v0p0p1_7.RSfetsym_0.QN.n10 GND 0.871f
C2507 frontAnalog_v0p0p1_7.RSfetsym_0.QN.t0 GND 0.0566f
C2508 frontAnalog_v0p0p1_7.RSfetsym_0.QN.n11 GND 2.48f
C2509 frontAnalog_v0p0p1_14.RSfetsym_0.QN.t1 GND 0.0322f
C2510 frontAnalog_v0p0p1_14.RSfetsym_0.QN.t2 GND 0.0322f
C2511 frontAnalog_v0p0p1_14.RSfetsym_0.QN.n0 GND 0.136f
C2512 frontAnalog_v0p0p1_14.RSfetsym_0.QN.t6 GND 0.0321f
C2513 frontAnalog_v0p0p1_14.RSfetsym_0.QN.t5 GND 0.0947f
C2514 frontAnalog_v0p0p1_14.RSfetsym_0.QN.n1 GND 1.46f
C2515 frontAnalog_v0p0p1_14.RSfetsym_0.QN.n2 GND 0.0784f
C2516 frontAnalog_v0p0p1_14.RSfetsym_0.QN.n3 GND 0.102f
C2517 frontAnalog_v0p0p1_14.RSfetsym_0.QN.n4 GND 0.445f
C2518 frontAnalog_v0p0p1_14.RSfetsym_0.QN.n5 GND 0.0126f
C2519 frontAnalog_v0p0p1_14.RSfetsym_0.QN.n6 GND 0.0341f
C2520 frontAnalog_v0p0p1_14.RSfetsym_0.QN.t4 GND 0.0322f
C2521 frontAnalog_v0p0p1_14.RSfetsym_0.QN.n7 GND 0.107f
C2522 frontAnalog_v0p0p1_14.RSfetsym_0.QN.n8 GND 0.131f
C2523 frontAnalog_v0p0p1_14.RSfetsym_0.QN.n9 GND 0.351f
C2524 frontAnalog_v0p0p1_14.RSfetsym_0.QN.n10 GND 0.871f
C2525 frontAnalog_v0p0p1_14.RSfetsym_0.QN.t3 GND 0.0566f
C2526 frontAnalog_v0p0p1_14.RSfetsym_0.QN.n11 GND 2.48f
C2527 frontAnalog_v0p0p1_5.x65.A.n0 GND 0.139f
C2528 frontAnalog_v0p0p1_5.x65.A.t4 GND 0.028f
C2529 frontAnalog_v0p0p1_5.x65.A.t6 GND 0.0175f
C2530 frontAnalog_v0p0p1_5.x65.A.n1 GND 0.0568f
C2531 frontAnalog_v0p0p1_5.x65.A.t2 GND 0.149f
C2532 frontAnalog_v0p0p1_5.x65.A.t7 GND 0.0318f
C2533 frontAnalog_v0p0p1_5.x65.A.t3 GND 0.141f
C2534 frontAnalog_v0p0p1_5.x65.A.t5 GND 0.219f
C2535 frontAnalog_v0p0p1_5.x65.A.n2 GND 1.37f
C2536 frontAnalog_v0p0p1_5.x65.A.n3 GND 0.898f
C2537 frontAnalog_v0p0p1_5.x65.A.t1 GND 0.463f
C2538 frontAnalog_v0p0p1_5.x65.A.t0 GND 0.0194f
C2539 frontAnalog_v0p0p1_5.x65.A.n4 GND 1.6f
C2540 frontAnalog_v0p0p1_5.x65.A.n5 GND 2.01f
C2541 frontAnalog_v0p0p1_5.x65.A.n6 GND 1.72f
C2542 frontAnalog_v0p0p1_1.x63.A.n0 GND 0.12f
C2543 frontAnalog_v0p0p1_1.x63.A.n1 GND 2.22f
C2544 frontAnalog_v0p0p1_1.x63.A.t6 GND 0.014f
C2545 frontAnalog_v0p0p1_1.x63.A.t7 GND 0.0225f
C2546 frontAnalog_v0p0p1_1.x63.A.n2 GND 0.0465f
C2547 frontAnalog_v0p0p1_1.x63.A.t2 GND 0.151f
C2548 frontAnalog_v0p0p1_1.x63.A.t4 GND 0.0256f
C2549 frontAnalog_v0p0p1_1.x63.A.t3 GND 0.173f
C2550 frontAnalog_v0p0p1_1.x63.A.t5 GND 0.175f
C2551 frontAnalog_v0p0p1_1.x63.A.n3 GND 1f
C2552 frontAnalog_v0p0p1_1.x63.A.n4 GND 0.953f
C2553 frontAnalog_v0p0p1_1.x63.A.t1 GND 0.0156f
C2554 frontAnalog_v0p0p1_1.x63.A.t0 GND 0.334f
C2555 frontAnalog_v0p0p1_1.x63.A.n5 GND 1.25f
C2556 16to4_PriorityEncoder_v0p0p1_0.I12.t7 GND 0.0226f
C2557 16to4_PriorityEncoder_v0p0p1_0.I12.n0 GND 0.355f
C2558 16to4_PriorityEncoder_v0p0p1_0.I12.n1 GND 0.107f
C2559 16to4_PriorityEncoder_v0p0p1_0.I12.n2 GND 0.047f
C2560 16to4_PriorityEncoder_v0p0p1_0.I12.n3 GND 0.0707f
C2561 16to4_PriorityEncoder_v0p0p1_0.I12.n4 GND 0.0756f
C2562 16to4_PriorityEncoder_v0p0p1_0.I12.n5 GND 0.104f
C2563 16to4_PriorityEncoder_v0p0p1_0.I12.n6 GND 0.0986f
C2564 16to4_PriorityEncoder_v0p0p1_0.I12.n7 GND 0.237f
C2565 16to4_PriorityEncoder_v0p0p1_0.I12.n14 GND 0.186f
C2566 16to4_PriorityEncoder_v0p0p1_0.I12.n15 GND 0.011f
C2567 16to4_PriorityEncoder_v0p0p1_0.I12.n16 GND 0.0301f
C2568 16to4_PriorityEncoder_v0p0p1_0.I12.n17 GND 0.327f
C2569 16to4_PriorityEncoder_v0p0p1_0.I12.n19 GND 0.142f
C2570 16to4_PriorityEncoder_v0p0p1_0.I12.n20 GND 0.303f
C2571 16to4_PriorityEncoder_v0p0p1_0.I12.n21 GND 0.41f
C2572 16to4_PriorityEncoder_v0p0p1_0.I12.n22 GND 8.85f
C2573 16to4_PriorityEncoder_v0p0p1_0.I12.n23 GND 16.3f
C2574 resistorDivider_v0p0p1_0.V8.t16 GND 0.022f
C2575 resistorDivider_v0p0p1_0.V8.n0 GND 0.18f
C2576 resistorDivider_v0p0p1_0.V8.n1 GND 0.0872f
C2577 resistorDivider_v0p0p1_0.V8.t13 GND 0.288f
C2578 resistorDivider_v0p0p1_0.V8.t5 GND 0.288f
C2579 resistorDivider_v0p0p1_0.V8.t12 GND 0.288f
C2580 resistorDivider_v0p0p1_0.V8.t15 GND 0.288f
C2581 resistorDivider_v0p0p1_0.V8.t11 GND 0.288f
C2582 resistorDivider_v0p0p1_0.V8.t1 GND 0.288f
C2583 resistorDivider_v0p0p1_0.V8.t7 GND 0.288f
C2584 resistorDivider_v0p0p1_0.V8.t6 GND 0.288f
C2585 resistorDivider_v0p0p1_0.V8.t14 GND 0.288f
C2586 resistorDivider_v0p0p1_0.V8.t10 GND 0.288f
C2587 resistorDivider_v0p0p1_0.V8.t8 GND 0.288f
C2588 resistorDivider_v0p0p1_0.V8.t3 GND 0.288f
C2589 resistorDivider_v0p0p1_0.V8.t4 GND 0.288f
C2590 resistorDivider_v0p0p1_0.V8.t9 GND 0.288f
C2591 resistorDivider_v0p0p1_0.V8.n2 GND 0.688f
C2592 resistorDivider_v0p0p1_0.V8.n3 GND 0.707f
C2593 resistorDivider_v0p0p1_0.V8.n4 GND 0.707f
C2594 resistorDivider_v0p0p1_0.V8.n5 GND 0.707f
C2595 resistorDivider_v0p0p1_0.V8.n6 GND 0.707f
C2596 resistorDivider_v0p0p1_0.V8.n7 GND 0.707f
C2597 resistorDivider_v0p0p1_0.V8.n8 GND 0.707f
C2598 resistorDivider_v0p0p1_0.V8.t2 GND 0.288f
C2599 resistorDivider_v0p0p1_0.V8.t0 GND 0.157f
C2600 resistorDivider_v0p0p1_0.V8.n9 GND 0.761f
C2601 frontAnalog_v0p0p1_11.x65.A.n0 GND 0.139f
C2602 frontAnalog_v0p0p1_11.x65.A.t4 GND 0.028f
C2603 frontAnalog_v0p0p1_11.x65.A.t6 GND 0.0175f
C2604 frontAnalog_v0p0p1_11.x65.A.n1 GND 0.0568f
C2605 frontAnalog_v0p0p1_11.x65.A.t1 GND 0.149f
C2606 frontAnalog_v0p0p1_11.x65.A.t7 GND 0.0318f
C2607 frontAnalog_v0p0p1_11.x65.A.t2 GND 0.141f
C2608 frontAnalog_v0p0p1_11.x65.A.t5 GND 0.219f
C2609 frontAnalog_v0p0p1_11.x65.A.n2 GND 1.37f
C2610 frontAnalog_v0p0p1_11.x65.A.n3 GND 0.898f
C2611 frontAnalog_v0p0p1_11.x65.A.t0 GND 0.463f
C2612 frontAnalog_v0p0p1_11.x65.A.t3 GND 0.0194f
C2613 frontAnalog_v0p0p1_11.x65.A.n4 GND 1.6f
C2614 frontAnalog_v0p0p1_11.x65.A.n5 GND 2.01f
C2615 frontAnalog_v0p0p1_11.x65.A.n6 GND 1.72f
C2616 frontAnalog_v0p0p1_12.RSfetsym_0.QN.t1 GND 0.0322f
C2617 frontAnalog_v0p0p1_12.RSfetsym_0.QN.t0 GND 0.0322f
C2618 frontAnalog_v0p0p1_12.RSfetsym_0.QN.n0 GND 0.136f
C2619 frontAnalog_v0p0p1_12.RSfetsym_0.QN.t6 GND 0.0321f
C2620 frontAnalog_v0p0p1_12.RSfetsym_0.QN.t5 GND 0.0947f
C2621 frontAnalog_v0p0p1_12.RSfetsym_0.QN.n1 GND 1.46f
C2622 frontAnalog_v0p0p1_12.RSfetsym_0.QN.n2 GND 0.0784f
C2623 frontAnalog_v0p0p1_12.RSfetsym_0.QN.n3 GND 0.102f
C2624 frontAnalog_v0p0p1_12.RSfetsym_0.QN.n4 GND 0.445f
C2625 frontAnalog_v0p0p1_12.RSfetsym_0.QN.n5 GND 0.0126f
C2626 frontAnalog_v0p0p1_12.RSfetsym_0.QN.n6 GND 0.0341f
C2627 frontAnalog_v0p0p1_12.RSfetsym_0.QN.t3 GND 0.0322f
C2628 frontAnalog_v0p0p1_12.RSfetsym_0.QN.n7 GND 0.107f
C2629 frontAnalog_v0p0p1_12.RSfetsym_0.QN.n8 GND 0.131f
C2630 frontAnalog_v0p0p1_12.RSfetsym_0.QN.n9 GND 0.351f
C2631 frontAnalog_v0p0p1_12.RSfetsym_0.QN.n10 GND 0.871f
C2632 frontAnalog_v0p0p1_12.RSfetsym_0.QN.t4 GND 0.0566f
C2633 frontAnalog_v0p0p1_12.RSfetsym_0.QN.n11 GND 2.48f
C2634 frontAnalog_v0p0p1_6.x63.A.n0 GND 0.12f
C2635 frontAnalog_v0p0p1_6.x63.A.n1 GND 2.22f
C2636 frontAnalog_v0p0p1_6.x63.A.t6 GND 0.014f
C2637 frontAnalog_v0p0p1_6.x63.A.t4 GND 0.0225f
C2638 frontAnalog_v0p0p1_6.x63.A.n2 GND 0.0465f
C2639 frontAnalog_v0p0p1_6.x63.A.t2 GND 0.151f
C2640 frontAnalog_v0p0p1_6.x63.A.t7 GND 0.0256f
C2641 frontAnalog_v0p0p1_6.x63.A.t3 GND 0.173f
C2642 frontAnalog_v0p0p1_6.x63.A.t5 GND 0.175f
C2643 frontAnalog_v0p0p1_6.x63.A.n3 GND 1f
C2644 frontAnalog_v0p0p1_6.x63.A.n4 GND 0.953f
C2645 frontAnalog_v0p0p1_6.x63.A.t1 GND 0.0156f
C2646 frontAnalog_v0p0p1_6.x63.A.t0 GND 0.334f
C2647 frontAnalog_v0p0p1_6.x63.A.n5 GND 1.25f
C2648 frontAnalog_v0p0p1_3.RSfetsym_0.QN.t2 GND 0.0322f
C2649 frontAnalog_v0p0p1_3.RSfetsym_0.QN.t3 GND 0.0322f
C2650 frontAnalog_v0p0p1_3.RSfetsym_0.QN.n0 GND 0.136f
C2651 frontAnalog_v0p0p1_3.RSfetsym_0.QN.t6 GND 0.0321f
C2652 frontAnalog_v0p0p1_3.RSfetsym_0.QN.t5 GND 0.0947f
C2653 frontAnalog_v0p0p1_3.RSfetsym_0.QN.n1 GND 1.46f
C2654 frontAnalog_v0p0p1_3.RSfetsym_0.QN.n2 GND 0.0784f
C2655 frontAnalog_v0p0p1_3.RSfetsym_0.QN.n3 GND 0.102f
C2656 frontAnalog_v0p0p1_3.RSfetsym_0.QN.n4 GND 0.445f
C2657 frontAnalog_v0p0p1_3.RSfetsym_0.QN.n5 GND 0.0126f
C2658 frontAnalog_v0p0p1_3.RSfetsym_0.QN.n6 GND 0.0341f
C2659 frontAnalog_v0p0p1_3.RSfetsym_0.QN.t4 GND 0.0322f
C2660 frontAnalog_v0p0p1_3.RSfetsym_0.QN.n7 GND 0.107f
C2661 frontAnalog_v0p0p1_3.RSfetsym_0.QN.n8 GND 0.131f
C2662 frontAnalog_v0p0p1_3.RSfetsym_0.QN.n9 GND 0.351f
C2663 frontAnalog_v0p0p1_3.RSfetsym_0.QN.n10 GND 0.871f
C2664 frontAnalog_v0p0p1_3.RSfetsym_0.QN.t0 GND 0.0566f
C2665 frontAnalog_v0p0p1_3.RSfetsym_0.QN.n11 GND 2.48f
C2666 frontAnalog_v0p0p1_11.Q.n6 GND 0.166f
C2667 frontAnalog_v0p0p1_11.Q.n8 GND 0.0269f
C2668 frontAnalog_v0p0p1_11.Q.n9 GND 0.292f
C2669 frontAnalog_v0p0p1_11.Q.n11 GND 0.127f
C2670 frontAnalog_v0p0p1_11.Q.n12 GND 0.271f
C2671 frontAnalog_v0p0p1_11.Q.n13 GND 0.373f
C2672 frontAnalog_v0p0p1_11.Q.n14 GND 7.04f
C2673 frontAnalog_v0p0p1_11.Q.t12 GND 0.0202f
C2674 frontAnalog_v0p0p1_11.Q.n15 GND 0.317f
C2675 frontAnalog_v0p0p1_11.Q.n16 GND 0.0953f
C2676 frontAnalog_v0p0p1_11.Q.n17 GND 0.042f
C2677 frontAnalog_v0p0p1_11.Q.n18 GND 0.0632f
C2678 frontAnalog_v0p0p1_11.Q.n19 GND 0.0676f
C2679 frontAnalog_v0p0p1_11.Q.n20 GND 0.0931f
C2680 frontAnalog_v0p0p1_11.Q.n21 GND 0.0881f
C2681 frontAnalog_v0p0p1_11.Q.n22 GND 0.203f
C2682 frontAnalog_v0p0p1_11.Q.n23 GND 11f
C2683 frontAnalog_v0p0p1_10.RSfetsym_0.QN.t2 GND 0.0322f
C2684 frontAnalog_v0p0p1_10.RSfetsym_0.QN.t3 GND 0.0322f
C2685 frontAnalog_v0p0p1_10.RSfetsym_0.QN.n0 GND 0.136f
C2686 frontAnalog_v0p0p1_10.RSfetsym_0.QN.t6 GND 0.0321f
C2687 frontAnalog_v0p0p1_10.RSfetsym_0.QN.t5 GND 0.0947f
C2688 frontAnalog_v0p0p1_10.RSfetsym_0.QN.n1 GND 1.46f
C2689 frontAnalog_v0p0p1_10.RSfetsym_0.QN.n2 GND 0.0784f
C2690 frontAnalog_v0p0p1_10.RSfetsym_0.QN.n3 GND 0.102f
C2691 frontAnalog_v0p0p1_10.RSfetsym_0.QN.n4 GND 0.445f
C2692 frontAnalog_v0p0p1_10.RSfetsym_0.QN.n5 GND 0.0126f
C2693 frontAnalog_v0p0p1_10.RSfetsym_0.QN.n6 GND 0.0341f
C2694 frontAnalog_v0p0p1_10.RSfetsym_0.QN.t0 GND 0.0322f
C2695 frontAnalog_v0p0p1_10.RSfetsym_0.QN.n7 GND 0.107f
C2696 frontAnalog_v0p0p1_10.RSfetsym_0.QN.n8 GND 0.131f
C2697 frontAnalog_v0p0p1_10.RSfetsym_0.QN.n9 GND 0.351f
C2698 frontAnalog_v0p0p1_10.RSfetsym_0.QN.n10 GND 0.871f
C2699 frontAnalog_v0p0p1_10.RSfetsym_0.QN.t4 GND 0.0566f
C2700 frontAnalog_v0p0p1_10.RSfetsym_0.QN.n11 GND 2.48f
C2701 frontAnalog_v0p0p1_1.x65.A.n0 GND 0.139f
C2702 frontAnalog_v0p0p1_1.x65.A.t4 GND 0.028f
C2703 frontAnalog_v0p0p1_1.x65.A.t6 GND 0.0175f
C2704 frontAnalog_v0p0p1_1.x65.A.n1 GND 0.0568f
C2705 frontAnalog_v0p0p1_1.x65.A.t7 GND 0.0318f
C2706 frontAnalog_v0p0p1_1.x65.A.t1 GND 0.141f
C2707 frontAnalog_v0p0p1_1.x65.A.t5 GND 0.219f
C2708 frontAnalog_v0p0p1_1.x65.A.n2 GND 1.37f
C2709 frontAnalog_v0p0p1_1.x65.A.n3 GND 0.898f
C2710 frontAnalog_v0p0p1_1.x65.A.t3 GND 0.463f
C2711 frontAnalog_v0p0p1_1.x65.A.t2 GND 0.0194f
C2712 frontAnalog_v0p0p1_1.x65.A.n4 GND 1.6f
C2713 frontAnalog_v0p0p1_1.x65.A.n5 GND 2.01f
C2714 frontAnalog_v0p0p1_1.x65.A.t0 GND 0.149f
C2715 frontAnalog_v0p0p1_1.x65.A.n6 GND 1.72f
C2716 frontAnalog_v0p0p1_4.x63.A.n0 GND 0.12f
C2717 frontAnalog_v0p0p1_4.x63.A.n1 GND 2.22f
C2718 frontAnalog_v0p0p1_4.x63.A.t5 GND 0.014f
C2719 frontAnalog_v0p0p1_4.x63.A.t6 GND 0.0225f
C2720 frontAnalog_v0p0p1_4.x63.A.n2 GND 0.0465f
C2721 frontAnalog_v0p0p1_4.x63.A.t2 GND 0.151f
C2722 frontAnalog_v0p0p1_4.x63.A.t4 GND 0.0256f
C2723 frontAnalog_v0p0p1_4.x63.A.t3 GND 0.173f
C2724 frontAnalog_v0p0p1_4.x63.A.t7 GND 0.175f
C2725 frontAnalog_v0p0p1_4.x63.A.n3 GND 1f
C2726 frontAnalog_v0p0p1_4.x63.A.n4 GND 0.953f
C2727 frontAnalog_v0p0p1_4.x63.A.t0 GND 0.0156f
C2728 frontAnalog_v0p0p1_4.x63.A.t1 GND 0.334f
C2729 frontAnalog_v0p0p1_4.x63.A.n5 GND 1.25f
C2730 frontAnalog_v0p0p1_15.x65.A.n0 GND 0.139f
C2731 frontAnalog_v0p0p1_15.x65.A.t4 GND 0.028f
C2732 frontAnalog_v0p0p1_15.x65.A.t6 GND 0.0175f
C2733 frontAnalog_v0p0p1_15.x65.A.n1 GND 0.0568f
C2734 frontAnalog_v0p0p1_15.x65.A.t3 GND 0.149f
C2735 frontAnalog_v0p0p1_15.x65.A.t7 GND 0.0318f
C2736 frontAnalog_v0p0p1_15.x65.A.t2 GND 0.141f
C2737 frontAnalog_v0p0p1_15.x65.A.t5 GND 0.219f
C2738 frontAnalog_v0p0p1_15.x65.A.n2 GND 1.37f
C2739 frontAnalog_v0p0p1_15.x65.A.n3 GND 0.898f
C2740 frontAnalog_v0p0p1_15.x65.A.t1 GND 0.463f
C2741 frontAnalog_v0p0p1_15.x65.A.t0 GND 0.0194f
C2742 frontAnalog_v0p0p1_15.x65.A.n4 GND 1.6f
C2743 frontAnalog_v0p0p1_15.x65.A.n5 GND 2.01f
C2744 frontAnalog_v0p0p1_15.x65.A.n6 GND 1.72f
C2745 frontAnalog_v0p0p1_3.x65.A.n0 GND 0.139f
C2746 frontAnalog_v0p0p1_3.x65.A.t4 GND 0.028f
C2747 frontAnalog_v0p0p1_3.x65.A.t6 GND 0.0175f
C2748 frontAnalog_v0p0p1_3.x65.A.n1 GND 0.0568f
C2749 frontAnalog_v0p0p1_3.x65.A.t7 GND 0.0318f
C2750 frontAnalog_v0p0p1_3.x65.A.t1 GND 0.141f
C2751 frontAnalog_v0p0p1_3.x65.A.t5 GND 0.219f
C2752 frontAnalog_v0p0p1_3.x65.A.n2 GND 1.37f
C2753 frontAnalog_v0p0p1_3.x65.A.n3 GND 0.898f
C2754 frontAnalog_v0p0p1_3.x65.A.t2 GND 0.463f
C2755 frontAnalog_v0p0p1_3.x65.A.t3 GND 0.0194f
C2756 frontAnalog_v0p0p1_3.x65.A.n4 GND 1.6f
C2757 frontAnalog_v0p0p1_3.x65.A.n5 GND 2.01f
C2758 frontAnalog_v0p0p1_3.x65.A.t0 GND 0.149f
C2759 frontAnalog_v0p0p1_3.x65.A.n6 GND 1.72f
C2760 frontAnalog_v0p0p1_3.x63.A.n0 GND 0.12f
C2761 frontAnalog_v0p0p1_3.x63.A.n1 GND 2.22f
C2762 frontAnalog_v0p0p1_3.x63.A.t7 GND 0.014f
C2763 frontAnalog_v0p0p1_3.x63.A.t5 GND 0.0225f
C2764 frontAnalog_v0p0p1_3.x63.A.n2 GND 0.0465f
C2765 frontAnalog_v0p0p1_3.x63.A.t1 GND 0.151f
C2766 frontAnalog_v0p0p1_3.x63.A.t3 GND 0.0156f
C2767 frontAnalog_v0p0p1_3.x63.A.t2 GND 0.335f
C2768 frontAnalog_v0p0p1_3.x63.A.t6 GND 0.0256f
C2769 frontAnalog_v0p0p1_3.x63.A.t0 GND 0.173f
C2770 frontAnalog_v0p0p1_3.x63.A.t4 GND 0.175f
C2771 frontAnalog_v0p0p1_3.x63.A.n3 GND 1f
C2772 frontAnalog_v0p0p1_3.x63.A.n4 GND 0.953f
C2773 frontAnalog_v0p0p1_3.x63.A.n5 GND 1.25f
C2774 frontAnalog_v0p0p1_5.x63.A.n0 GND 0.12f
C2775 frontAnalog_v0p0p1_5.x63.A.n1 GND 2.22f
C2776 frontAnalog_v0p0p1_5.x63.A.t6 GND 0.014f
C2777 frontAnalog_v0p0p1_5.x63.A.t4 GND 0.0225f
C2778 frontAnalog_v0p0p1_5.x63.A.n2 GND 0.0465f
C2779 frontAnalog_v0p0p1_5.x63.A.t5 GND 0.0256f
C2780 frontAnalog_v0p0p1_5.x63.A.t2 GND 0.173f
C2781 frontAnalog_v0p0p1_5.x63.A.t7 GND 0.175f
C2782 frontAnalog_v0p0p1_5.x63.A.n3 GND 1f
C2783 frontAnalog_v0p0p1_5.x63.A.n4 GND 0.953f
C2784 frontAnalog_v0p0p1_5.x63.A.t0 GND 0.0156f
C2785 frontAnalog_v0p0p1_5.x63.A.t3 GND 0.335f
C2786 frontAnalog_v0p0p1_5.x63.A.t1 GND 0.151f
C2787 frontAnalog_v0p0p1_5.x63.A.n5 GND 1.25f
C2788 frontAnalog_v0p0p1_10.x63.A.n0 GND 0.12f
C2789 frontAnalog_v0p0p1_10.x63.A.n1 GND 2.22f
C2790 frontAnalog_v0p0p1_10.x63.A.t7 GND 0.014f
C2791 frontAnalog_v0p0p1_10.x63.A.t5 GND 0.0225f
C2792 frontAnalog_v0p0p1_10.x63.A.n2 GND 0.0465f
C2793 frontAnalog_v0p0p1_10.x63.A.t1 GND 0.151f
C2794 frontAnalog_v0p0p1_10.x63.A.t3 GND 0.0156f
C2795 frontAnalog_v0p0p1_10.x63.A.t2 GND 0.335f
C2796 frontAnalog_v0p0p1_10.x63.A.t6 GND 0.0256f
C2797 frontAnalog_v0p0p1_10.x63.A.t0 GND 0.173f
C2798 frontAnalog_v0p0p1_10.x63.A.t4 GND 0.175f
C2799 frontAnalog_v0p0p1_10.x63.A.n3 GND 1f
C2800 frontAnalog_v0p0p1_10.x63.A.n4 GND 0.953f
C2801 frontAnalog_v0p0p1_10.x63.A.n5 GND 1.25f
C2802 frontAnalog_v0p0p1_13.x63.A.n0 GND 0.12f
C2803 frontAnalog_v0p0p1_13.x63.A.n1 GND 2.22f
C2804 frontAnalog_v0p0p1_13.x63.A.t6 GND 0.014f
C2805 frontAnalog_v0p0p1_13.x63.A.t4 GND 0.0225f
C2806 frontAnalog_v0p0p1_13.x63.A.n2 GND 0.0465f
C2807 frontAnalog_v0p0p1_13.x63.A.t5 GND 0.0256f
C2808 frontAnalog_v0p0p1_13.x63.A.t2 GND 0.173f
C2809 frontAnalog_v0p0p1_13.x63.A.t7 GND 0.175f
C2810 frontAnalog_v0p0p1_13.x63.A.n3 GND 1f
C2811 frontAnalog_v0p0p1_13.x63.A.n4 GND 0.953f
C2812 frontAnalog_v0p0p1_13.x63.A.t0 GND 0.0156f
C2813 frontAnalog_v0p0p1_13.x63.A.t3 GND 0.335f
C2814 frontAnalog_v0p0p1_13.x63.A.t1 GND 0.151f
C2815 frontAnalog_v0p0p1_13.x63.A.n5 GND 1.25f
C2816 resistorDivider_v0p0p1_0.V5.t16 GND 0.0238f
C2817 resistorDivider_v0p0p1_0.V5.n0 GND 0.195f
C2818 resistorDivider_v0p0p1_0.V5.n1 GND 0.0942f
C2819 resistorDivider_v0p0p1_0.V5.t3 GND 0.311f
C2820 resistorDivider_v0p0p1_0.V5.t1 GND 0.311f
C2821 resistorDivider_v0p0p1_0.V5.t9 GND 0.311f
C2822 resistorDivider_v0p0p1_0.V5.t5 GND 0.311f
C2823 resistorDivider_v0p0p1_0.V5.t2 GND 0.311f
C2824 resistorDivider_v0p0p1_0.V5.t7 GND 0.311f
C2825 resistorDivider_v0p0p1_0.V5.t11 GND 0.311f
C2826 resistorDivider_v0p0p1_0.V5.t6 GND 0.311f
C2827 resistorDivider_v0p0p1_0.V5.t10 GND 0.311f
C2828 resistorDivider_v0p0p1_0.V5.t4 GND 0.311f
C2829 resistorDivider_v0p0p1_0.V5.t15 GND 0.311f
C2830 resistorDivider_v0p0p1_0.V5.t13 GND 0.311f
C2831 resistorDivider_v0p0p1_0.V5.t12 GND 0.311f
C2832 resistorDivider_v0p0p1_0.V5.t8 GND 0.67f
C2833 resistorDivider_v0p0p1_0.V5.t14 GND 0.311f
C2834 resistorDivider_v0p0p1_0.V5.n2 GND 0.385f
C2835 resistorDivider_v0p0p1_0.V5.n3 GND 0.382f
C2836 resistorDivider_v0p0p1_0.V5.n4 GND 0.382f
C2837 resistorDivider_v0p0p1_0.V5.t0 GND 0.17f
C2838 resistorDivider_v0p0p1_0.V5.n5 GND 0.523f
C2839 resistorDivider_v0p0p1_0.V5.n6 GND 0.382f
C2840 resistorDivider_v0p0p1_0.V5.n7 GND 0.382f
C2841 resistorDivider_v0p0p1_0.V5.n8 GND 0.382f
C2842 resistorDivider_v0p0p1_0.V5.n9 GND 0.382f
C2843 resistorDivider_v0p0p1_0.V5.n10 GND 0.382f
C2844 resistorDivider_v0p0p1_0.V5.n11 GND 0.382f
C2845 resistorDivider_v0p0p1_0.V5.n12 GND 0.382f
C2846 resistorDivider_v0p0p1_0.V5.n13 GND 0.382f
C2847 resistorDivider_v0p0p1_0.V5.n14 GND 0.382f
C2848 resistorDivider_v0p0p1_0.V5.n15 GND 0.382f
C2849 resistorDivider_v0p0p1_0.V5.n16 GND 0.306f
C2850 resistorDivider_v0p0p1_0.V6.t16 GND 0.0241f
C2851 resistorDivider_v0p0p1_0.V6.n0 GND 0.197f
C2852 resistorDivider_v0p0p1_0.V6.n1 GND 0.0955f
C2853 resistorDivider_v0p0p1_0.V6.t2 GND 0.315f
C2854 resistorDivider_v0p0p1_0.V6.t11 GND 0.315f
C2855 resistorDivider_v0p0p1_0.V6.t6 GND 0.315f
C2856 resistorDivider_v0p0p1_0.V6.t3 GND 0.315f
C2857 resistorDivider_v0p0p1_0.V6.t1 GND 0.315f
C2858 resistorDivider_v0p0p1_0.V6.t14 GND 0.315f
C2859 resistorDivider_v0p0p1_0.V6.t9 GND 0.315f
C2860 resistorDivider_v0p0p1_0.V6.t5 GND 0.315f
C2861 resistorDivider_v0p0p1_0.V6.t8 GND 0.315f
C2862 resistorDivider_v0p0p1_0.V6.t10 GND 0.315f
C2863 resistorDivider_v0p0p1_0.V6.t15 GND 0.315f
C2864 resistorDivider_v0p0p1_0.V6.t7 GND 0.315f
C2865 resistorDivider_v0p0p1_0.V6.t12 GND 0.315f
C2866 resistorDivider_v0p0p1_0.V6.t4 GND 0.315f
C2867 resistorDivider_v0p0p1_0.V6.t13 GND 0.315f
C2868 resistorDivider_v0p0p1_0.V6.t0 GND 0.679f
C2869 resistorDivider_v0p0p1_0.V6.n2 GND 0.39f
C2870 resistorDivider_v0p0p1_0.V6.n3 GND 0.387f
C2871 resistorDivider_v0p0p1_0.V6.n4 GND 0.387f
C2872 resistorDivider_v0p0p1_0.V6.n5 GND 0.387f
C2873 resistorDivider_v0p0p1_0.V6.n6 GND 0.387f
C2874 resistorDivider_v0p0p1_0.V6.n7 GND 0.387f
C2875 resistorDivider_v0p0p1_0.V6.n8 GND 0.387f
C2876 resistorDivider_v0p0p1_0.V6.n9 GND 0.387f
C2877 resistorDivider_v0p0p1_0.V6.n10 GND 0.387f
C2878 resistorDivider_v0p0p1_0.V6.n11 GND 0.387f
C2879 resistorDivider_v0p0p1_0.V6.n12 GND 0.387f
C2880 resistorDivider_v0p0p1_0.V6.n13 GND 0.387f
C2881 resistorDivider_v0p0p1_0.V6.n14 GND 0.387f
C2882 resistorDivider_v0p0p1_0.V6.n15 GND 0.387f
C2883 resistorDivider_v0p0p1_0.V6.n16 GND 0.301f
C2884 resistorDivider_v0p0p1_0.V7.t17 GND 0.0233f
C2885 resistorDivider_v0p0p1_0.V7.n0 GND 0.191f
C2886 resistorDivider_v0p0p1_0.V7.n1 GND 0.0964f
C2887 resistorDivider_v0p0p1_0.V7.t13 GND 0.305f
C2888 resistorDivider_v0p0p1_0.V7.t6 GND 0.305f
C2889 resistorDivider_v0p0p1_0.V7.t4 GND 0.305f
C2890 resistorDivider_v0p0p1_0.V7.t15 GND 0.305f
C2891 resistorDivider_v0p0p1_0.V7.t14 GND 0.305f
C2892 resistorDivider_v0p0p1_0.V7.t1 GND 0.305f
C2893 resistorDivider_v0p0p1_0.V7.t9 GND 0.305f
C2894 resistorDivider_v0p0p1_0.V7.t8 GND 0.305f
C2895 resistorDivider_v0p0p1_0.V7.t12 GND 0.305f
C2896 resistorDivider_v0p0p1_0.V7.t10 GND 0.305f
C2897 resistorDivider_v0p0p1_0.V7.t11 GND 0.305f
C2898 resistorDivider_v0p0p1_0.V7.t3 GND 0.305f
C2899 resistorDivider_v0p0p1_0.V7.t7 GND 0.305f
C2900 resistorDivider_v0p0p1_0.V7.t2 GND 0.305f
C2901 resistorDivider_v0p0p1_0.V7.t5 GND 0.305f
C2902 resistorDivider_v0p0p1_0.V7.n2 GND 0.73f
C2903 resistorDivider_v0p0p1_0.V7.n3 GND 0.749f
C2904 resistorDivider_v0p0p1_0.V7.n4 GND 0.749f
C2905 resistorDivider_v0p0p1_0.V7.n5 GND 0.749f
C2906 resistorDivider_v0p0p1_0.V7.n6 GND 0.749f
C2907 resistorDivider_v0p0p1_0.V7.n7 GND 0.749f
C2908 resistorDivider_v0p0p1_0.V7.n8 GND 0.749f
C2909 resistorDivider_v0p0p1_0.V7.t0 GND 0.167f
C2910 resistorDivider_v0p0p1_0.V7.n9 GND 0.808f
C2911 frontAnalog_v0p0p1_7.Q.t7 GND 0.0147f
C2912 frontAnalog_v0p0p1_7.Q.n0 GND 0.0157f
C2913 frontAnalog_v0p0p1_7.Q.n1 GND 0.674f
C2914 frontAnalog_v0p0p1_7.Q.t10 GND 0.0108f
C2915 frontAnalog_v0p0p1_7.Q.t6 GND 0.0331f
C2916 frontAnalog_v0p0p1_7.Q.n2 GND 0.519f
C2917 frontAnalog_v0p0p1_7.Q.n3 GND 0.0687f
C2918 frontAnalog_v0p0p1_7.Q.n4 GND 0.156f
C2919 frontAnalog_v0p0p1_7.Q.t0 GND 0.0111f
C2920 frontAnalog_v0p0p1_7.Q.n5 GND 0.103f
C2921 frontAnalog_v0p0p1_7.Q.n6 GND 0.11f
C2922 frontAnalog_v0p0p1_7.Q.t1 GND 0.0111f
C2923 frontAnalog_v0p0p1_7.Q.t2 GND 0.0111f
C2924 frontAnalog_v0p0p1_7.Q.n7 GND 0.152f
C2925 frontAnalog_v0p0p1_7.Q.n8 GND 0.144f
C2926 frontAnalog_v0p0p1_7.Q.t4 GND 0.0122f
C2927 frontAnalog_v0p0p1_7.Q.n9 GND 0.345f
C2928 frontAnalog_v0p0p1_7.Q.n10 GND 9.94f
C2929 frontAnalog_v0p0p1_7.Q.n11 GND 4.4f
C2930 frontAnalog_v0p0p1_7.Q.n12 GND 1.18f
C2931 frontAnalog_v0p0p1_7.Q.n13 GND 0.872f
C2932 frontAnalog_v0p0p1_7.x63.A.n0 GND 0.12f
C2933 frontAnalog_v0p0p1_7.x63.A.n1 GND 2.22f
C2934 frontAnalog_v0p0p1_7.x63.A.t4 GND 0.014f
C2935 frontAnalog_v0p0p1_7.x63.A.t6 GND 0.0225f
C2936 frontAnalog_v0p0p1_7.x63.A.n2 GND 0.0465f
C2937 frontAnalog_v0p0p1_7.x63.A.t1 GND 0.151f
C2938 frontAnalog_v0p0p1_7.x63.A.t2 GND 0.0156f
C2939 frontAnalog_v0p0p1_7.x63.A.t3 GND 0.335f
C2940 frontAnalog_v0p0p1_7.x63.A.t7 GND 0.0256f
C2941 frontAnalog_v0p0p1_7.x63.A.t0 GND 0.173f
C2942 frontAnalog_v0p0p1_7.x63.A.t5 GND 0.175f
C2943 frontAnalog_v0p0p1_7.x63.A.n3 GND 1f
C2944 frontAnalog_v0p0p1_7.x63.A.n4 GND 0.953f
C2945 frontAnalog_v0p0p1_7.x63.A.n5 GND 1.25f
C2946 frontAnalog_v0p0p1_7.x65.A.n0 GND 0.139f
C2947 frontAnalog_v0p0p1_7.x65.A.t7 GND 0.028f
C2948 frontAnalog_v0p0p1_7.x65.A.t5 GND 0.0175f
C2949 frontAnalog_v0p0p1_7.x65.A.n1 GND 0.0568f
C2950 frontAnalog_v0p0p1_7.x65.A.t6 GND 0.0318f
C2951 frontAnalog_v0p0p1_7.x65.A.t1 GND 0.141f
C2952 frontAnalog_v0p0p1_7.x65.A.t4 GND 0.219f
C2953 frontAnalog_v0p0p1_7.x65.A.n2 GND 1.37f
C2954 frontAnalog_v0p0p1_7.x65.A.n3 GND 0.898f
C2955 frontAnalog_v0p0p1_7.x65.A.t2 GND 0.463f
C2956 frontAnalog_v0p0p1_7.x65.A.t3 GND 0.0194f
C2957 frontAnalog_v0p0p1_7.x65.A.n4 GND 1.6f
C2958 frontAnalog_v0p0p1_7.x65.A.n5 GND 2.01f
C2959 frontAnalog_v0p0p1_7.x65.A.t0 GND 0.149f
C2960 frontAnalog_v0p0p1_7.x65.A.n6 GND 1.72f
C2961 frontAnalog_v0p0p1_13.RSfetsym_0.QN.t1 GND 0.0322f
C2962 frontAnalog_v0p0p1_13.RSfetsym_0.QN.t0 GND 0.0322f
C2963 frontAnalog_v0p0p1_13.RSfetsym_0.QN.n0 GND 0.136f
C2964 frontAnalog_v0p0p1_13.RSfetsym_0.QN.t6 GND 0.0321f
C2965 frontAnalog_v0p0p1_13.RSfetsym_0.QN.t5 GND 0.0947f
C2966 frontAnalog_v0p0p1_13.RSfetsym_0.QN.n1 GND 1.46f
C2967 frontAnalog_v0p0p1_13.RSfetsym_0.QN.n2 GND 0.0784f
C2968 frontAnalog_v0p0p1_13.RSfetsym_0.QN.n3 GND 0.102f
C2969 frontAnalog_v0p0p1_13.RSfetsym_0.QN.n4 GND 0.445f
C2970 frontAnalog_v0p0p1_13.RSfetsym_0.QN.n5 GND 0.0126f
C2971 frontAnalog_v0p0p1_13.RSfetsym_0.QN.n6 GND 0.0341f
C2972 frontAnalog_v0p0p1_13.RSfetsym_0.QN.t4 GND 0.0322f
C2973 frontAnalog_v0p0p1_13.RSfetsym_0.QN.n7 GND 0.107f
C2974 frontAnalog_v0p0p1_13.RSfetsym_0.QN.n8 GND 0.131f
C2975 frontAnalog_v0p0p1_13.RSfetsym_0.QN.n9 GND 0.351f
C2976 frontAnalog_v0p0p1_13.RSfetsym_0.QN.n10 GND 0.871f
C2977 frontAnalog_v0p0p1_13.RSfetsym_0.QN.t3 GND 0.0566f
C2978 frontAnalog_v0p0p1_13.RSfetsym_0.QN.n11 GND 2.48f
C2979 frontAnalog_v0p0p1_9.Q.n2 GND 0.0175f
C2980 frontAnalog_v0p0p1_9.Q.n9 GND 0.0126f
C2981 frontAnalog_v0p0p1_9.Q.n10 GND 0.155f
C2982 frontAnalog_v0p0p1_9.Q.n11 GND 0.393f
C2983 frontAnalog_v0p0p1_9.Q.n12 GND 0.0114f
C2984 frontAnalog_v0p0p1_9.Q.n13 GND 0.0116f
C2985 frontAnalog_v0p0p1_9.Q.n14 GND 0.203f
C2986 frontAnalog_v0p0p1_9.Q.n17 GND 0.0149f
C2987 frontAnalog_v0p0p1_9.Q.n21 GND 0.487f
C2988 frontAnalog_v0p0p1_9.Q.n22 GND 0.793f
C2989 frontAnalog_v0p0p1_9.Q.n23 GND 0.497f
C2990 frontAnalog_v0p0p1_9.Q.n24 GND 7.52f
C2991 frontAnalog_v0p0p1_9.Q.t9 GND 0.0117f
C2992 frontAnalog_v0p0p1_9.Q.t5 GND 0.0359f
C2993 frontAnalog_v0p0p1_9.Q.n25 GND 0.563f
C2994 frontAnalog_v0p0p1_9.Q.n26 GND 0.169f
C2995 frontAnalog_v0p0p1_9.Q.n27 GND 0.0746f
C2996 frontAnalog_v0p0p1_9.Q.t3 GND 0.0121f
C2997 frontAnalog_v0p0p1_9.Q.n28 GND 0.112f
C2998 frontAnalog_v0p0p1_9.Q.n29 GND 0.12f
C2999 frontAnalog_v0p0p1_9.Q.t0 GND 0.0121f
C3000 frontAnalog_v0p0p1_9.Q.t1 GND 0.0121f
C3001 frontAnalog_v0p0p1_9.Q.n30 GND 0.165f
C3002 frontAnalog_v0p0p1_9.Q.n31 GND 0.156f
C3003 frontAnalog_v0p0p1_9.Q.t4 GND 0.0132f
C3004 frontAnalog_v0p0p1_9.Q.n32 GND 0.36f
C3005 frontAnalog_v0p0p1_9.Q.n33 GND 12.9f
C3006 frontAnalog_v0p0p1_9.RSfetsym_0.QN.t1 GND 0.0322f
C3007 frontAnalog_v0p0p1_9.RSfetsym_0.QN.t2 GND 0.0322f
C3008 frontAnalog_v0p0p1_9.RSfetsym_0.QN.n0 GND 0.136f
C3009 frontAnalog_v0p0p1_9.RSfetsym_0.QN.t6 GND 0.0321f
C3010 frontAnalog_v0p0p1_9.RSfetsym_0.QN.t5 GND 0.0947f
C3011 frontAnalog_v0p0p1_9.RSfetsym_0.QN.n1 GND 1.46f
C3012 frontAnalog_v0p0p1_9.RSfetsym_0.QN.n2 GND 0.0784f
C3013 frontAnalog_v0p0p1_9.RSfetsym_0.QN.n3 GND 0.102f
C3014 frontAnalog_v0p0p1_9.RSfetsym_0.QN.n4 GND 0.445f
C3015 frontAnalog_v0p0p1_9.RSfetsym_0.QN.n5 GND 0.0126f
C3016 frontAnalog_v0p0p1_9.RSfetsym_0.QN.n6 GND 0.0341f
C3017 frontAnalog_v0p0p1_9.RSfetsym_0.QN.t4 GND 0.0322f
C3018 frontAnalog_v0p0p1_9.RSfetsym_0.QN.n7 GND 0.107f
C3019 frontAnalog_v0p0p1_9.RSfetsym_0.QN.n8 GND 0.131f
C3020 frontAnalog_v0p0p1_9.RSfetsym_0.QN.n9 GND 0.351f
C3021 frontAnalog_v0p0p1_9.RSfetsym_0.QN.n10 GND 0.871f
C3022 frontAnalog_v0p0p1_9.RSfetsym_0.QN.t0 GND 0.0566f
C3023 frontAnalog_v0p0p1_9.RSfetsym_0.QN.n11 GND 2.48f
C3024 frontAnalog_v0p0p1_14.Q.n0 GND 0.369f
C3025 frontAnalog_v0p0p1_14.Q.n2 GND 0.274f
C3026 frontAnalog_v0p0p1_14.Q.n3 GND 0.487f
C3027 frontAnalog_v0p0p1_14.Q.n4 GND 7.62f
C3028 frontAnalog_v0p0p1_14.Q.t5 GND 0.0138f
C3029 frontAnalog_v0p0p1_14.Q.n5 GND 0.216f
C3030 frontAnalog_v0p0p1_14.Q.n6 GND 0.0648f
C3031 frontAnalog_v0p0p1_14.Q.n7 GND 0.0286f
C3032 frontAnalog_v0p0p1_14.Q.n8 GND 0.043f
C3033 frontAnalog_v0p0p1_14.Q.n9 GND 0.046f
C3034 frontAnalog_v0p0p1_14.Q.n10 GND 0.0634f
C3035 frontAnalog_v0p0p1_14.Q.n11 GND 0.0599f
C3036 frontAnalog_v0p0p1_14.Q.n12 GND 0.138f
C3037 frontAnalog_v0p0p1_14.Q.n13 GND 11.3f
C3038 frontAnalog_v0p0p1_9.x65.A.n0 GND 0.139f
C3039 frontAnalog_v0p0p1_9.x65.A.t6 GND 0.028f
C3040 frontAnalog_v0p0p1_9.x65.A.t4 GND 0.0175f
C3041 frontAnalog_v0p0p1_9.x65.A.n1 GND 0.0568f
C3042 frontAnalog_v0p0p1_9.x65.A.t2 GND 0.149f
C3043 frontAnalog_v0p0p1_9.x65.A.t5 GND 0.0318f
C3044 frontAnalog_v0p0p1_9.x65.A.t3 GND 0.141f
C3045 frontAnalog_v0p0p1_9.x65.A.t7 GND 0.219f
C3046 frontAnalog_v0p0p1_9.x65.A.n2 GND 1.37f
C3047 frontAnalog_v0p0p1_9.x65.A.n3 GND 0.898f
C3048 frontAnalog_v0p0p1_9.x65.A.t1 GND 0.463f
C3049 frontAnalog_v0p0p1_9.x65.A.t0 GND 0.0194f
C3050 frontAnalog_v0p0p1_9.x65.A.n4 GND 1.6f
C3051 frontAnalog_v0p0p1_9.x65.A.n5 GND 2.01f
C3052 frontAnalog_v0p0p1_9.x65.A.n6 GND 1.72f
C3053 frontAnalog_v0p0p1_9.x63.A.n0 GND 0.12f
C3054 frontAnalog_v0p0p1_9.x63.A.n1 GND 2.22f
C3055 frontAnalog_v0p0p1_9.x63.A.t7 GND 0.014f
C3056 frontAnalog_v0p0p1_9.x63.A.t5 GND 0.0225f
C3057 frontAnalog_v0p0p1_9.x63.A.n2 GND 0.0465f
C3058 frontAnalog_v0p0p1_9.x63.A.t2 GND 0.151f
C3059 frontAnalog_v0p0p1_9.x63.A.t6 GND 0.0256f
C3060 frontAnalog_v0p0p1_9.x63.A.t3 GND 0.173f
C3061 frontAnalog_v0p0p1_9.x63.A.t4 GND 0.175f
C3062 frontAnalog_v0p0p1_9.x63.A.n3 GND 1f
C3063 frontAnalog_v0p0p1_9.x63.A.n4 GND 0.953f
C3064 frontAnalog_v0p0p1_9.x63.A.t0 GND 0.0156f
C3065 frontAnalog_v0p0p1_9.x63.A.t1 GND 0.334f
C3066 frontAnalog_v0p0p1_9.x63.A.n5 GND 1.25f
C3067 resistorDivider_v0p0p1_0.V12.t16 GND 0.0235f
C3068 resistorDivider_v0p0p1_0.V12.n0 GND 0.193f
C3069 resistorDivider_v0p0p1_0.V12.n1 GND 0.0932f
C3070 resistorDivider_v0p0p1_0.V12.t14 GND 0.308f
C3071 resistorDivider_v0p0p1_0.V12.t15 GND 0.308f
C3072 resistorDivider_v0p0p1_0.V12.t4 GND 0.308f
C3073 resistorDivider_v0p0p1_0.V12.t13 GND 0.308f
C3074 resistorDivider_v0p0p1_0.V12.t9 GND 0.308f
C3075 resistorDivider_v0p0p1_0.V12.t8 GND 0.308f
C3076 resistorDivider_v0p0p1_0.V12.t1 GND 0.308f
C3077 resistorDivider_v0p0p1_0.V12.t11 GND 0.308f
C3078 resistorDivider_v0p0p1_0.V12.t12 GND 0.308f
C3079 resistorDivider_v0p0p1_0.V12.t10 GND 0.308f
C3080 resistorDivider_v0p0p1_0.V12.t2 GND 0.308f
C3081 resistorDivider_v0p0p1_0.V12.t7 GND 0.308f
C3082 resistorDivider_v0p0p1_0.V12.t5 GND 0.308f
C3083 resistorDivider_v0p0p1_0.V12.t6 GND 0.308f
C3084 resistorDivider_v0p0p1_0.V12.t3 GND 0.664f
C3085 resistorDivider_v0p0p1_0.V12.n2 GND 0.381f
C3086 resistorDivider_v0p0p1_0.V12.n3 GND 0.378f
C3087 resistorDivider_v0p0p1_0.V12.n4 GND 0.378f
C3088 resistorDivider_v0p0p1_0.V12.n5 GND 0.378f
C3089 resistorDivider_v0p0p1_0.V12.n6 GND 0.378f
C3090 resistorDivider_v0p0p1_0.V12.t0 GND 0.168f
C3091 resistorDivider_v0p0p1_0.V12.n7 GND 0.517f
C3092 resistorDivider_v0p0p1_0.V12.n8 GND 0.378f
C3093 resistorDivider_v0p0p1_0.V12.n9 GND 0.378f
C3094 resistorDivider_v0p0p1_0.V12.n10 GND 0.378f
C3095 resistorDivider_v0p0p1_0.V12.n11 GND 0.378f
C3096 resistorDivider_v0p0p1_0.V12.n12 GND 0.378f
C3097 resistorDivider_v0p0p1_0.V12.n13 GND 0.378f
C3098 resistorDivider_v0p0p1_0.V12.n14 GND 0.378f
C3099 resistorDivider_v0p0p1_0.V12.n15 GND 0.378f
C3100 resistorDivider_v0p0p1_0.V12.n16 GND 0.298f
C3101 frontAnalog_v0p0p1_4.x65.A.n0 GND 0.139f
C3102 frontAnalog_v0p0p1_4.x65.A.t4 GND 0.028f
C3103 frontAnalog_v0p0p1_4.x65.A.t5 GND 0.0175f
C3104 frontAnalog_v0p0p1_4.x65.A.n1 GND 0.0568f
C3105 frontAnalog_v0p0p1_4.x65.A.t7 GND 0.0318f
C3106 frontAnalog_v0p0p1_4.x65.A.t1 GND 0.141f
C3107 frontAnalog_v0p0p1_4.x65.A.t6 GND 0.219f
C3108 frontAnalog_v0p0p1_4.x65.A.n2 GND 1.37f
C3109 frontAnalog_v0p0p1_4.x65.A.n3 GND 0.898f
C3110 frontAnalog_v0p0p1_4.x65.A.t3 GND 0.463f
C3111 frontAnalog_v0p0p1_4.x65.A.t2 GND 0.0194f
C3112 frontAnalog_v0p0p1_4.x65.A.n4 GND 1.6f
C3113 frontAnalog_v0p0p1_4.x65.A.n5 GND 2.01f
C3114 frontAnalog_v0p0p1_4.x65.A.t0 GND 0.149f
C3115 frontAnalog_v0p0p1_4.x65.A.n6 GND 1.72f
C3116 VIN.t3 GND 0.0561f
C3117 VIN.n0 GND 0.453f
C3118 VIN.n1 GND 0.127f
C3119 VIN.t17 GND 0.0561f
C3120 VIN.n3 GND 0.45f
C3121 VIN.n4 GND 5.68f
C3122 VIN.t22 GND 0.0561f
C3123 VIN.n5 GND 0.453f
C3124 VIN.t8 GND 0.0561f
C3125 VIN.n6 GND 0.45f
C3126 VIN.t14 GND 0.0561f
C3127 VIN.n7 GND 0.453f
C3128 VIN.t29 GND 0.0561f
C3129 VIN.n8 GND 0.453f
C3130 VIN.t2 GND 0.0561f
C3131 VIN.n9 GND 0.453f
C3132 VIN.t9 GND 0.0561f
C3133 VIN.n10 GND 0.453f
C3134 VIN.t27 GND 0.0561f
C3135 VIN.n11 GND 0.453f
C3136 VIN.t30 GND 0.0561f
C3137 VIN.n12 GND 0.453f
C3138 VIN.t21 GND 0.0561f
C3139 VIN.n13 GND 0.453f
C3140 VIN.t25 GND 0.0561f
C3141 VIN.n14 GND 0.453f
C3142 VIN.t12 GND 0.0561f
C3143 VIN.n15 GND 0.453f
C3144 VIN.t18 GND 0.0561f
C3145 VIN.n16 GND 0.453f
C3146 VIN.t0 GND 0.0561f
C3147 VIN.n17 GND 0.453f
C3148 VIN.t7 GND 0.0561f
C3149 VIN.n18 GND 0.453f
C3150 VIN.n19 GND 11.9f
C3151 VIN.n20 GND 7.41f
C3152 VIN.n21 GND 7.41f
C3153 VIN.n22 GND 7.41f
C3154 VIN.n23 GND 7.41f
C3155 VIN.n24 GND 7.41f
C3156 VIN.n25 GND 7.42f
C3157 VIN.n26 GND 7.41f
C3158 VIN.n27 GND 7.41f
C3159 VIN.n28 GND 7.41f
C3160 VIN.n29 GND 7.41f
C3161 VIN.n30 GND 7.38f
C3162 VIN.n31 GND 7.41f
C3163 VIN.n32 GND 7.49f
C3164 VIN.n33 GND 1.18f
C3165 resistorDivider_v0p0p1_0.V13.t17 GND 0.024f
C3166 resistorDivider_v0p0p1_0.V13.n0 GND 0.196f
C3167 resistorDivider_v0p0p1_0.V13.n1 GND 0.095f
C3168 resistorDivider_v0p0p1_0.V13.t14 GND 0.313f
C3169 resistorDivider_v0p0p1_0.V13.t15 GND 0.313f
C3170 resistorDivider_v0p0p1_0.V13.t12 GND 0.313f
C3171 resistorDivider_v0p0p1_0.V13.t10 GND 0.313f
C3172 resistorDivider_v0p0p1_0.V13.t8 GND 0.313f
C3173 resistorDivider_v0p0p1_0.V13.t7 GND 0.313f
C3174 resistorDivider_v0p0p1_0.V13.t11 GND 0.313f
C3175 resistorDivider_v0p0p1_0.V13.t2 GND 0.313f
C3176 resistorDivider_v0p0p1_0.V13.t1 GND 0.313f
C3177 resistorDivider_v0p0p1_0.V13.t9 GND 0.313f
C3178 resistorDivider_v0p0p1_0.V13.t3 GND 0.313f
C3179 resistorDivider_v0p0p1_0.V13.t6 GND 0.313f
C3180 resistorDivider_v0p0p1_0.V13.t5 GND 0.313f
C3181 resistorDivider_v0p0p1_0.V13.t13 GND 0.313f
C3182 resistorDivider_v0p0p1_0.V13.t4 GND 0.313f
C3183 resistorDivider_v0p0p1_0.V13.t0 GND 0.171f
C3184 resistorDivider_v0p0p1_0.V13.n2 GND 0.892f
C3185 resistorDivider_v0p0p1_0.V13.n3 GND 0.77f
C3186 resistorDivider_v0p0p1_0.V13.n4 GND 0.77f
C3187 resistorDivider_v0p0p1_0.V13.n5 GND 0.77f
C3188 resistorDivider_v0p0p1_0.V13.n6 GND 0.77f
C3189 resistorDivider_v0p0p1_0.V13.n7 GND 0.77f
C3190 resistorDivider_v0p0p1_0.V13.n8 GND 0.77f
C3191 resistorDivider_v0p0p1_0.V13.n9 GND 0.684f
C3192 resistorDivider_v0p0p1_0.V14.t16 GND 0.0249f
C3193 resistorDivider_v0p0p1_0.V14.n0 GND 0.204f
C3194 resistorDivider_v0p0p1_0.V14.n1 GND 0.0945f
C3195 resistorDivider_v0p0p1_0.V14.t15 GND 0.326f
C3196 resistorDivider_v0p0p1_0.V14.t2 GND 0.326f
C3197 resistorDivider_v0p0p1_0.V14.t11 GND 0.326f
C3198 resistorDivider_v0p0p1_0.V14.t14 GND 0.326f
C3199 resistorDivider_v0p0p1_0.V14.t8 GND 0.326f
C3200 resistorDivider_v0p0p1_0.V14.t9 GND 0.326f
C3201 resistorDivider_v0p0p1_0.V14.t5 GND 0.326f
C3202 resistorDivider_v0p0p1_0.V14.t4 GND 0.326f
C3203 resistorDivider_v0p0p1_0.V14.t10 GND 0.326f
C3204 resistorDivider_v0p0p1_0.V14.t1 GND 0.326f
C3205 resistorDivider_v0p0p1_0.V14.t7 GND 0.326f
C3206 resistorDivider_v0p0p1_0.V14.t12 GND 0.326f
C3207 resistorDivider_v0p0p1_0.V14.t13 GND 0.326f
C3208 resistorDivider_v0p0p1_0.V14.t3 GND 0.326f
C3209 resistorDivider_v0p0p1_0.V14.t6 GND 0.326f
C3210 resistorDivider_v0p0p1_0.V14.t0 GND 0.178f
C3211 resistorDivider_v0p0p1_0.V14.n2 GND 0.929f
C3212 resistorDivider_v0p0p1_0.V14.n3 GND 0.801f
C3213 resistorDivider_v0p0p1_0.V14.n4 GND 0.801f
C3214 resistorDivider_v0p0p1_0.V14.n5 GND 0.801f
C3215 resistorDivider_v0p0p1_0.V14.n6 GND 0.801f
C3216 resistorDivider_v0p0p1_0.V14.n7 GND 0.801f
C3217 resistorDivider_v0p0p1_0.V14.n8 GND 0.801f
C3218 resistorDivider_v0p0p1_0.V14.n9 GND 0.719f
C3219 frontAnalog_v0p0p1_10.IB.n0 GND 0.0726f
C3220 frontAnalog_v0p0p1_10.IB.t12 GND 0.0832f
C3221 frontAnalog_v0p0p1_10.IB.t23 GND 0.0823f
C3222 frontAnalog_v0p0p1_10.IB.t3 GND 0.0832f
C3223 frontAnalog_v0p0p1_10.IB.t11 GND 0.0823f
C3224 frontAnalog_v0p0p1_10.IB.n3 GND 8.18f
C3225 frontAnalog_v0p0p1_10.IB.t32 GND 0.0832f
C3226 frontAnalog_v0p0p1_10.IB.t9 GND 0.0823f
C3227 frontAnalog_v0p0p1_10.IB.t5 GND 0.0832f
C3228 frontAnalog_v0p0p1_10.IB.t29 GND 0.0823f
C3229 frontAnalog_v0p0p1_10.IB.t22 GND 0.0832f
C3230 frontAnalog_v0p0p1_10.IB.t34 GND 0.0823f
C3231 frontAnalog_v0p0p1_10.IB.t26 GND 0.0832f
C3232 frontAnalog_v0p0p1_10.IB.t19 GND 0.0823f
C3233 frontAnalog_v0p0p1_10.IB.t15 GND 0.0832f
C3234 frontAnalog_v0p0p1_10.IB.t25 GND 0.0823f
C3235 frontAnalog_v0p0p1_10.IB.t18 GND 0.0832f
C3236 frontAnalog_v0p0p1_10.IB.t30 GND 0.0823f
C3237 frontAnalog_v0p0p1_10.IB.t7 GND 0.0832f
C3238 frontAnalog_v0p0p1_10.IB.t16 GND 0.0823f
C3239 frontAnalog_v0p0p1_10.IB.t10 GND 0.0832f
C3240 frontAnalog_v0p0p1_10.IB.t20 GND 0.0823f
C3241 frontAnalog_v0p0p1_10.IB.t31 GND 0.0832f
C3242 frontAnalog_v0p0p1_10.IB.t8 GND 0.0823f
C3243 frontAnalog_v0p0p1_10.IB.t4 GND 0.0832f
C3244 frontAnalog_v0p0p1_10.IB.t13 GND 0.0823f
C3245 frontAnalog_v0p0p1_10.IB.t21 GND 0.0832f
C3246 frontAnalog_v0p0p1_10.IB.t33 GND 0.0823f
C3247 frontAnalog_v0p0p1_10.IB.t27 GND 0.0832f
C3248 frontAnalog_v0p0p1_10.IB.t6 GND 0.0823f
C3249 frontAnalog_v0p0p1_10.IB.t14 GND 0.0832f
C3250 frontAnalog_v0p0p1_10.IB.t24 GND 0.0823f
C3251 frontAnalog_v0p0p1_10.IB.t17 GND 0.0832f
C3252 frontAnalog_v0p0p1_10.IB.t28 GND 0.0823f
C3253 frontAnalog_v0p0p1_10.IB.n18 GND 12.2f
C3254 frontAnalog_v0p0p1_10.IB.n19 GND 8.47f
C3255 frontAnalog_v0p0p1_10.IB.n20 GND 8.42f
C3256 frontAnalog_v0p0p1_10.IB.n21 GND 8.53f
C3257 frontAnalog_v0p0p1_10.IB.n22 GND 8.42f
C3258 frontAnalog_v0p0p1_10.IB.n23 GND 8.48f
C3259 frontAnalog_v0p0p1_10.IB.n24 GND 8.43f
C3260 frontAnalog_v0p0p1_10.IB.n25 GND 8.47f
C3261 frontAnalog_v0p0p1_10.IB.n26 GND 8.42f
C3262 frontAnalog_v0p0p1_10.IB.n27 GND 8.43f
C3263 frontAnalog_v0p0p1_10.IB.n28 GND 8.48f
C3264 frontAnalog_v0p0p1_10.IB.n29 GND 8.53f
C3265 frontAnalog_v0p0p1_10.IB.n30 GND 7.05f
C3266 frontAnalog_v0p0p1_10.IB.n31 GND 14.7f
C3267 frontAnalog_v0p0p1_10.IB.t0 GND 0.0463f
C3268 frontAnalog_v0p0p1_10.IB.n32 GND 0.124f
C3269 frontAnalog_v0p0p1_10.IB.n33 GND 0.0147f
C3270 frontAnalog_v0p0p1_10.IB.t2 GND 0.634f
C3271 frontAnalog_v0p0p1_10.IB.n34 GND 10.9f
C3272 16to4_PriorityEncoder_v0p0p1_0.I13.t12 GND 0.0207f
C3273 16to4_PriorityEncoder_v0p0p1_0.I13.n0 GND 0.325f
C3274 16to4_PriorityEncoder_v0p0p1_0.I13.n1 GND 0.0975f
C3275 16to4_PriorityEncoder_v0p0p1_0.I13.n2 GND 0.043f
C3276 16to4_PriorityEncoder_v0p0p1_0.I13.n3 GND 0.0647f
C3277 16to4_PriorityEncoder_v0p0p1_0.I13.n4 GND 0.0691f
C3278 16to4_PriorityEncoder_v0p0p1_0.I13.n5 GND 0.0953f
C3279 16to4_PriorityEncoder_v0p0p1_0.I13.n6 GND 0.0902f
C3280 16to4_PriorityEncoder_v0p0p1_0.I13.n7 GND 0.217f
C3281 16to4_PriorityEncoder_v0p0p1_0.I13.n8 GND 0.0101f
C3282 16to4_PriorityEncoder_v0p0p1_0.I13.n16 GND 0.113f
C3283 16to4_PriorityEncoder_v0p0p1_0.I13.n17 GND 0.263f
C3284 16to4_PriorityEncoder_v0p0p1_0.I13.n24 GND 0.16f
C3285 16to4_PriorityEncoder_v0p0p1_0.I13.n29 GND 0.425f
C3286 16to4_PriorityEncoder_v0p0p1_0.I13.n30 GND 1.01f
C3287 16to4_PriorityEncoder_v0p0p1_0.I13.n31 GND 0.47f
C3288 16to4_PriorityEncoder_v0p0p1_0.I13.n32 GND 0.292f
C3289 16to4_PriorityEncoder_v0p0p1_0.I13.n33 GND 10.5f
C3290 16to4_PriorityEncoder_v0p0p1_0.I13.n34 GND 17.1f
C3291 frontAnalog_v0p0p1_6.RSfetsym_0.QN.t1 GND 0.0322f
C3292 frontAnalog_v0p0p1_6.RSfetsym_0.QN.t2 GND 0.0322f
C3293 frontAnalog_v0p0p1_6.RSfetsym_0.QN.n0 GND 0.136f
C3294 frontAnalog_v0p0p1_6.RSfetsym_0.QN.t6 GND 0.0321f
C3295 frontAnalog_v0p0p1_6.RSfetsym_0.QN.t5 GND 0.0947f
C3296 frontAnalog_v0p0p1_6.RSfetsym_0.QN.n1 GND 1.46f
C3297 frontAnalog_v0p0p1_6.RSfetsym_0.QN.n2 GND 0.0784f
C3298 frontAnalog_v0p0p1_6.RSfetsym_0.QN.n3 GND 0.102f
C3299 frontAnalog_v0p0p1_6.RSfetsym_0.QN.n4 GND 0.445f
C3300 frontAnalog_v0p0p1_6.RSfetsym_0.QN.n5 GND 0.0126f
C3301 frontAnalog_v0p0p1_6.RSfetsym_0.QN.n6 GND 0.0341f
C3302 frontAnalog_v0p0p1_6.RSfetsym_0.QN.t3 GND 0.0322f
C3303 frontAnalog_v0p0p1_6.RSfetsym_0.QN.n7 GND 0.107f
C3304 frontAnalog_v0p0p1_6.RSfetsym_0.QN.n8 GND 0.131f
C3305 frontAnalog_v0p0p1_6.RSfetsym_0.QN.n9 GND 0.351f
C3306 frontAnalog_v0p0p1_6.RSfetsym_0.QN.n10 GND 0.871f
C3307 frontAnalog_v0p0p1_6.RSfetsym_0.QN.t4 GND 0.0566f
C3308 frontAnalog_v0p0p1_6.RSfetsym_0.QN.n11 GND 2.48f
C3309 frontAnalog_v0p0p1_6.Q.t7 GND 0.0109f
C3310 frontAnalog_v0p0p1_6.Q.t5 GND 0.0333f
C3311 frontAnalog_v0p0p1_6.Q.n0 GND 0.522f
C3312 frontAnalog_v0p0p1_6.Q.n1 GND 0.157f
C3313 frontAnalog_v0p0p1_6.Q.n2 GND 0.0691f
C3314 frontAnalog_v0p0p1_6.Q.t3 GND 0.0112f
C3315 frontAnalog_v0p0p1_6.Q.n3 GND 0.104f
C3316 frontAnalog_v0p0p1_6.Q.n4 GND 0.111f
C3317 frontAnalog_v0p0p1_6.Q.t1 GND 0.0112f
C3318 frontAnalog_v0p0p1_6.Q.t2 GND 0.0112f
C3319 frontAnalog_v0p0p1_6.Q.n5 GND 0.153f
C3320 frontAnalog_v0p0p1_6.Q.n6 GND 0.145f
C3321 frontAnalog_v0p0p1_6.Q.t4 GND 0.0123f
C3322 frontAnalog_v0p0p1_6.Q.n7 GND 0.349f
C3323 frontAnalog_v0p0p1_6.Q.n8 GND 0.0165f
C3324 frontAnalog_v0p0p1_6.Q.n9 GND 0.119f
C3325 frontAnalog_v0p0p1_6.Q.n10 GND 0.243f
C3326 frontAnalog_v0p0p1_6.Q.n11 GND 0.0105f
C3327 frontAnalog_v0p0p1_6.Q.n12 GND 0.011f
C3328 frontAnalog_v0p0p1_6.Q.n13 GND 0.603f
C3329 frontAnalog_v0p0p1_6.Q.n14 GND 0.0188f
C3330 frontAnalog_v0p0p1_6.Q.n15 GND 0.0877f
C3331 frontAnalog_v0p0p1_6.Q.n16 GND 1.47f
C3332 frontAnalog_v0p0p1_6.Q.n17 GND 9.05f
C3333 frontAnalog_v0p0p1_6.Q.n18 GND 13.6f
C3334 frontAnalog_v0p0p1_15.RSfetsym_0.QN.t3 GND 0.0322f
C3335 frontAnalog_v0p0p1_15.RSfetsym_0.QN.t2 GND 0.0322f
C3336 frontAnalog_v0p0p1_15.RSfetsym_0.QN.n0 GND 0.136f
C3337 frontAnalog_v0p0p1_15.RSfetsym_0.QN.t6 GND 0.0321f
C3338 frontAnalog_v0p0p1_15.RSfetsym_0.QN.t5 GND 0.0947f
C3339 frontAnalog_v0p0p1_15.RSfetsym_0.QN.n1 GND 1.46f
C3340 frontAnalog_v0p0p1_15.RSfetsym_0.QN.n2 GND 0.0784f
C3341 frontAnalog_v0p0p1_15.RSfetsym_0.QN.n3 GND 0.102f
C3342 frontAnalog_v0p0p1_15.RSfetsym_0.QN.n4 GND 0.445f
C3343 frontAnalog_v0p0p1_15.RSfetsym_0.QN.n5 GND 0.0126f
C3344 frontAnalog_v0p0p1_15.RSfetsym_0.QN.n6 GND 0.0341f
C3345 frontAnalog_v0p0p1_15.RSfetsym_0.QN.t0 GND 0.0322f
C3346 frontAnalog_v0p0p1_15.RSfetsym_0.QN.n7 GND 0.107f
C3347 frontAnalog_v0p0p1_15.RSfetsym_0.QN.n8 GND 0.131f
C3348 frontAnalog_v0p0p1_15.RSfetsym_0.QN.n9 GND 0.351f
C3349 frontAnalog_v0p0p1_15.RSfetsym_0.QN.n10 GND 0.871f
C3350 frontAnalog_v0p0p1_15.RSfetsym_0.QN.t1 GND 0.0566f
C3351 frontAnalog_v0p0p1_15.RSfetsym_0.QN.n11 GND 2.48f
C3352 frontAnalog_v0p0p1_2.x65.A.n0 GND 0.139f
C3353 frontAnalog_v0p0p1_2.x65.A.t4 GND 0.028f
C3354 frontAnalog_v0p0p1_2.x65.A.t5 GND 0.0175f
C3355 frontAnalog_v0p0p1_2.x65.A.n1 GND 0.0568f
C3356 frontAnalog_v0p0p1_2.x65.A.t1 GND 0.149f
C3357 frontAnalog_v0p0p1_2.x65.A.t3 GND 0.463f
C3358 frontAnalog_v0p0p1_2.x65.A.t2 GND 0.0194f
C3359 frontAnalog_v0p0p1_2.x65.A.n2 GND 1.6f
C3360 frontAnalog_v0p0p1_2.x65.A.t6 GND 0.0318f
C3361 frontAnalog_v0p0p1_2.x65.A.t0 GND 0.141f
C3362 frontAnalog_v0p0p1_2.x65.A.t7 GND 0.219f
C3363 frontAnalog_v0p0p1_2.x65.A.n3 GND 1.37f
C3364 frontAnalog_v0p0p1_2.x65.A.n4 GND 0.898f
C3365 frontAnalog_v0p0p1_2.x65.A.n5 GND 2.01f
C3366 frontAnalog_v0p0p1_2.x65.A.n6 GND 1.72f
C3367 frontAnalog_v0p0p1_2.x63.A.n0 GND 0.12f
C3368 frontAnalog_v0p0p1_2.x63.A.n1 GND 2.22f
C3369 frontAnalog_v0p0p1_2.x63.A.t6 GND 0.014f
C3370 frontAnalog_v0p0p1_2.x63.A.t5 GND 0.0225f
C3371 frontAnalog_v0p0p1_2.x63.A.n2 GND 0.0465f
C3372 frontAnalog_v0p0p1_2.x63.A.t2 GND 0.151f
C3373 frontAnalog_v0p0p1_2.x63.A.t4 GND 0.0256f
C3374 frontAnalog_v0p0p1_2.x63.A.t3 GND 0.173f
C3375 frontAnalog_v0p0p1_2.x63.A.t7 GND 0.175f
C3376 frontAnalog_v0p0p1_2.x63.A.n3 GND 1f
C3377 frontAnalog_v0p0p1_2.x63.A.n4 GND 0.953f
C3378 frontAnalog_v0p0p1_2.x63.A.t0 GND 0.0156f
C3379 frontAnalog_v0p0p1_2.x63.A.t1 GND 0.334f
C3380 frontAnalog_v0p0p1_2.x63.A.n5 GND 1.25f
C3381 resistorDivider_v0p0p1_0.V15.t17 GND 0.0258f
C3382 resistorDivider_v0p0p1_0.V15.n0 GND 0.212f
C3383 resistorDivider_v0p0p1_0.V15.n1 GND 0.0979f
C3384 resistorDivider_v0p0p1_0.V15.t1 GND 0.338f
C3385 resistorDivider_v0p0p1_0.V15.t5 GND 0.338f
C3386 resistorDivider_v0p0p1_0.V15.t14 GND 0.338f
C3387 resistorDivider_v0p0p1_0.V15.t12 GND 0.338f
C3388 resistorDivider_v0p0p1_0.V15.t8 GND 0.338f
C3389 resistorDivider_v0p0p1_0.V15.t13 GND 0.338f
C3390 resistorDivider_v0p0p1_0.V15.t3 GND 0.338f
C3391 resistorDivider_v0p0p1_0.V15.t15 GND 0.338f
C3392 resistorDivider_v0p0p1_0.V15.t6 GND 0.338f
C3393 resistorDivider_v0p0p1_0.V15.t10 GND 0.338f
C3394 resistorDivider_v0p0p1_0.V15.t4 GND 0.338f
C3395 resistorDivider_v0p0p1_0.V15.t2 GND 0.338f
C3396 resistorDivider_v0p0p1_0.V15.t11 GND 0.338f
C3397 resistorDivider_v0p0p1_0.V15.t7 GND 0.338f
C3398 resistorDivider_v0p0p1_0.V15.t9 GND 0.338f
C3399 resistorDivider_v0p0p1_0.V15.n2 GND 0.808f
C3400 resistorDivider_v0p0p1_0.V15.n3 GND 0.829f
C3401 resistorDivider_v0p0p1_0.V15.n4 GND 0.829f
C3402 resistorDivider_v0p0p1_0.V15.t0 GND 0.185f
C3403 resistorDivider_v0p0p1_0.V15.n5 GND 0.982f
C3404 resistorDivider_v0p0p1_0.V15.n6 GND 0.829f
C3405 resistorDivider_v0p0p1_0.V15.n7 GND 0.829f
C3406 resistorDivider_v0p0p1_0.V15.n8 GND 0.829f
C3407 resistorDivider_v0p0p1_0.V15.n9 GND 0.74f
C3408 resistorDivider_v0p0p1_0.V9.t16 GND 0.0231f
C3409 resistorDivider_v0p0p1_0.V9.n0 GND 0.189f
C3410 resistorDivider_v0p0p1_0.V9.n1 GND 0.0915f
C3411 resistorDivider_v0p0p1_0.V9.t2 GND 0.302f
C3412 resistorDivider_v0p0p1_0.V9.t11 GND 0.302f
C3413 resistorDivider_v0p0p1_0.V9.t10 GND 0.302f
C3414 resistorDivider_v0p0p1_0.V9.t8 GND 0.302f
C3415 resistorDivider_v0p0p1_0.V9.t15 GND 0.302f
C3416 resistorDivider_v0p0p1_0.V9.t7 GND 0.302f
C3417 resistorDivider_v0p0p1_0.V9.t4 GND 0.302f
C3418 resistorDivider_v0p0p1_0.V9.t3 GND 0.302f
C3419 resistorDivider_v0p0p1_0.V9.t9 GND 0.302f
C3420 resistorDivider_v0p0p1_0.V9.t14 GND 0.302f
C3421 resistorDivider_v0p0p1_0.V9.t12 GND 0.302f
C3422 resistorDivider_v0p0p1_0.V9.t5 GND 0.302f
C3423 resistorDivider_v0p0p1_0.V9.t13 GND 0.302f
C3424 resistorDivider_v0p0p1_0.V9.t6 GND 0.302f
C3425 resistorDivider_v0p0p1_0.V9.t1 GND 0.302f
C3426 resistorDivider_v0p0p1_0.V9.n2 GND 0.723f
C3427 resistorDivider_v0p0p1_0.V9.n3 GND 0.742f
C3428 resistorDivider_v0p0p1_0.V9.n4 GND 0.742f
C3429 resistorDivider_v0p0p1_0.V9.n5 GND 0.742f
C3430 resistorDivider_v0p0p1_0.V9.n6 GND 0.742f
C3431 resistorDivider_v0p0p1_0.V9.n7 GND 0.742f
C3432 resistorDivider_v0p0p1_0.V9.n8 GND 0.742f
C3433 resistorDivider_v0p0p1_0.V9.t0 GND 0.165f
C3434 resistorDivider_v0p0p1_0.V9.n9 GND 0.803f
C3435 frontAnalog_v0p0p1_8.RSfetsym_0.QN.t2 GND 0.0322f
C3436 frontAnalog_v0p0p1_8.RSfetsym_0.QN.t3 GND 0.0322f
C3437 frontAnalog_v0p0p1_8.RSfetsym_0.QN.n0 GND 0.136f
C3438 frontAnalog_v0p0p1_8.RSfetsym_0.QN.t5 GND 0.0321f
C3439 frontAnalog_v0p0p1_8.RSfetsym_0.QN.t6 GND 0.0947f
C3440 frontAnalog_v0p0p1_8.RSfetsym_0.QN.n1 GND 1.46f
C3441 frontAnalog_v0p0p1_8.RSfetsym_0.QN.n2 GND 0.0784f
C3442 frontAnalog_v0p0p1_8.RSfetsym_0.QN.n3 GND 0.102f
C3443 frontAnalog_v0p0p1_8.RSfetsym_0.QN.n4 GND 0.445f
C3444 frontAnalog_v0p0p1_8.RSfetsym_0.QN.n5 GND 0.0126f
C3445 frontAnalog_v0p0p1_8.RSfetsym_0.QN.n6 GND 0.0341f
C3446 frontAnalog_v0p0p1_8.RSfetsym_0.QN.t4 GND 0.0322f
C3447 frontAnalog_v0p0p1_8.RSfetsym_0.QN.n7 GND 0.107f
C3448 frontAnalog_v0p0p1_8.RSfetsym_0.QN.n8 GND 0.131f
C3449 frontAnalog_v0p0p1_8.RSfetsym_0.QN.n9 GND 0.351f
C3450 frontAnalog_v0p0p1_8.RSfetsym_0.QN.n10 GND 0.871f
C3451 frontAnalog_v0p0p1_8.RSfetsym_0.QN.t0 GND 0.0566f
C3452 frontAnalog_v0p0p1_8.RSfetsym_0.QN.n11 GND 2.48f
C3453 OUT1.n2 GND 0.0114f
C3454 OUT1.n4 GND 0.0242f
C3455 OUT1.n6 GND 0.0161f
C3456 OUT1.n8 GND 0.0161f
C3457 OUT1.n10 GND 0.0161f
C3458 OUT1.n12 GND 0.0161f
C3459 OUT1.n14 GND 0.0161f
C3460 OUT1.n23 GND 0.014f
C3461 OUT1.n25 GND 0.0348f
C3462 OUT1.n27 GND 0.021f
C3463 OUT1.n29 GND 0.021f
C3464 OUT1.n31 GND 0.021f
C3465 OUT1.n33 GND 0.021f
C3466 OUT1.n35 GND 0.021f
C3467 OUT1.n37 GND 0.0147f
C3468 OUT1.n38 GND 0.0297f
C3469 OUT1.n39 GND 0.0229f
C3470 OUT1.n42 GND 0.0114f
C3471 OUT1.n44 GND 0.0242f
C3472 OUT1.n46 GND 0.0161f
C3473 OUT1.n48 GND 0.0161f
C3474 OUT1.n50 GND 0.0161f
C3475 OUT1.n52 GND 0.0161f
C3476 OUT1.n54 GND 0.0161f
C3477 OUT1.n63 GND 0.014f
C3478 OUT1.n65 GND 0.0348f
C3479 OUT1.n67 GND 0.021f
C3480 OUT1.n69 GND 0.021f
C3481 OUT1.n71 GND 0.021f
C3482 OUT1.n73 GND 0.021f
C3483 OUT1.n75 GND 0.021f
C3484 OUT1.n77 GND 0.0147f
C3485 OUT1.n78 GND 0.0274f
C3486 OUT1.n79 GND 0.0203f
C3487 OUT1.n81 GND 0.0114f
C3488 OUT1.n83 GND 0.0242f
C3489 OUT1.n85 GND 0.0161f
C3490 OUT1.n87 GND 0.0161f
C3491 OUT1.n89 GND 0.0161f
C3492 OUT1.n91 GND 0.0161f
C3493 OUT1.n93 GND 0.0161f
C3494 OUT1.n97 GND 0.0126f
C3495 OUT1.n100 GND 0.014f
C3496 OUT1.n102 GND 0.0348f
C3497 OUT1.n104 GND 0.021f
C3498 OUT1.n106 GND 0.021f
C3499 OUT1.n108 GND 0.021f
C3500 OUT1.n110 GND 0.021f
C3501 OUT1.n112 GND 0.021f
C3502 OUT1.n114 GND 0.0147f
C3503 OUT1.n115 GND 0.0284f
C3504 OUT1.n116 GND 0.0234f
C3505 OUT1.n120 GND 0.014f
C3506 OUT1.n122 GND 0.0348f
C3507 OUT1.n124 GND 0.021f
C3508 OUT1.n126 GND 0.021f
C3509 OUT1.n128 GND 0.021f
C3510 OUT1.n130 GND 0.021f
C3511 OUT1.n132 GND 0.021f
C3512 OUT1.n136 GND 0.0114f
C3513 OUT1.n138 GND 0.0242f
C3514 OUT1.n140 GND 0.0161f
C3515 OUT1.n142 GND 0.0161f
C3516 OUT1.n144 GND 0.0161f
C3517 OUT1.n146 GND 0.0161f
C3518 OUT1.n148 GND 0.0161f
C3519 OUT1.n152 GND 0.0129f
C3520 OUT1.n155 GND 0.0204f
C3521 OUT1.n156 GND 0.108f
C3522 OUT1.n157 GND 0.275f
C3523 OUT1.n158 GND 0.224f
C3524 OUT1.n159 GND 0.228f
C3525 frontAnalog_v0p0p1_12.Q.n1 GND 0.0619f
C3526 frontAnalog_v0p0p1_12.Q.n2 GND 0.126f
C3527 frontAnalog_v0p0p1_12.Q.n5 GND 0.321f
C3528 frontAnalog_v0p0p1_12.Q.n7 GND 0.0436f
C3529 frontAnalog_v0p0p1_12.Q.n8 GND 0.762f
C3530 frontAnalog_v0p0p1_12.Q.n9 GND 8.38f
C3531 frontAnalog_v0p0p1_12.Q.t10 GND 0.0173f
C3532 frontAnalog_v0p0p1_12.Q.n10 GND 0.271f
C3533 frontAnalog_v0p0p1_12.Q.n11 GND 0.0814f
C3534 frontAnalog_v0p0p1_12.Q.n12 GND 0.0359f
C3535 frontAnalog_v0p0p1_12.Q.n13 GND 0.054f
C3536 frontAnalog_v0p0p1_12.Q.n14 GND 0.0577f
C3537 frontAnalog_v0p0p1_12.Q.n15 GND 0.0795f
C3538 frontAnalog_v0p0p1_12.Q.n16 GND 0.0752f
C3539 frontAnalog_v0p0p1_12.Q.n17 GND 0.173f
C3540 frontAnalog_v0p0p1_12.Q.n18 GND 12.5f
C3541 frontAnalog_v0p0p1_15.Q.n1 GND 0.0912f
C3542 frontAnalog_v0p0p1_15.Q.n2 GND 0.243f
C3543 frontAnalog_v0p0p1_15.Q.n3 GND 5.7f
C3544 frontAnalog_v0p0p1_15.Q.n4 GND 0.141f
C3545 frontAnalog_v0p0p1_15.Q.n5 GND 0.0422f
C3546 frontAnalog_v0p0p1_15.Q.n6 GND 0.0186f
C3547 frontAnalog_v0p0p1_15.Q.n7 GND 0.028f
C3548 frontAnalog_v0p0p1_15.Q.n8 GND 0.0299f
C3549 frontAnalog_v0p0p1_15.Q.n9 GND 0.0413f
C3550 frontAnalog_v0p0p1_15.Q.n10 GND 0.039f
C3551 frontAnalog_v0p0p1_15.Q.n11 GND 0.0899f
C3552 frontAnalog_v0p0p1_15.Q.n12 GND 8.16f
C3553 resistorDivider_v0p0p1_0.V1.t16 GND 0.0127f
C3554 resistorDivider_v0p0p1_0.V1.n0 GND 0.104f
C3555 resistorDivider_v0p0p1_0.V1.n1 GND 0.0503f
C3556 resistorDivider_v0p0p1_0.V1.t2 GND 0.166f
C3557 resistorDivider_v0p0p1_0.V1.t14 GND 0.166f
C3558 resistorDivider_v0p0p1_0.V1.t10 GND 0.166f
C3559 resistorDivider_v0p0p1_0.V1.t1 GND 0.166f
C3560 resistorDivider_v0p0p1_0.V1.t13 GND 0.166f
C3561 resistorDivider_v0p0p1_0.V1.t11 GND 0.166f
C3562 resistorDivider_v0p0p1_0.V1.t15 GND 0.166f
C3563 resistorDivider_v0p0p1_0.V1.t5 GND 0.166f
C3564 resistorDivider_v0p0p1_0.V1.t6 GND 0.166f
C3565 resistorDivider_v0p0p1_0.V1.t12 GND 0.166f
C3566 resistorDivider_v0p0p1_0.V1.t4 GND 0.166f
C3567 resistorDivider_v0p0p1_0.V1.t3 GND 0.166f
C3568 resistorDivider_v0p0p1_0.V1.t7 GND 0.166f
C3569 resistorDivider_v0p0p1_0.V1.t9 GND 0.166f
C3570 resistorDivider_v0p0p1_0.V1.t8 GND 0.166f
C3571 resistorDivider_v0p0p1_0.V1.n2 GND 0.398f
C3572 resistorDivider_v0p0p1_0.V1.n3 GND 0.408f
C3573 resistorDivider_v0p0p1_0.V1.n4 GND 0.408f
C3574 resistorDivider_v0p0p1_0.V1.n5 GND 0.408f
C3575 resistorDivider_v0p0p1_0.V1.n6 GND 0.408f
C3576 resistorDivider_v0p0p1_0.V1.n7 GND 0.408f
C3577 resistorDivider_v0p0p1_0.V1.n8 GND 0.408f
C3578 resistorDivider_v0p0p1_0.V1.t0 GND 0.0908f
C3579 resistorDivider_v0p0p1_0.V1.n9 GND 0.437f
C3580 resistorDivider_v0p0p1_0.V2.t17 GND 0.023f
C3581 resistorDivider_v0p0p1_0.V2.n0 GND 0.188f
C3582 resistorDivider_v0p0p1_0.V2.n1 GND 0.0951f
C3583 resistorDivider_v0p0p1_0.V2.t2 GND 0.301f
C3584 resistorDivider_v0p0p1_0.V2.t15 GND 0.301f
C3585 resistorDivider_v0p0p1_0.V2.t11 GND 0.301f
C3586 resistorDivider_v0p0p1_0.V2.t13 GND 0.301f
C3587 resistorDivider_v0p0p1_0.V2.t1 GND 0.301f
C3588 resistorDivider_v0p0p1_0.V2.t6 GND 0.301f
C3589 resistorDivider_v0p0p1_0.V2.t7 GND 0.301f
C3590 resistorDivider_v0p0p1_0.V2.t10 GND 0.301f
C3591 resistorDivider_v0p0p1_0.V2.t4 GND 0.301f
C3592 resistorDivider_v0p0p1_0.V2.t12 GND 0.301f
C3593 resistorDivider_v0p0p1_0.V2.t8 GND 0.301f
C3594 resistorDivider_v0p0p1_0.V2.t14 GND 0.301f
C3595 resistorDivider_v0p0p1_0.V2.t3 GND 0.301f
C3596 resistorDivider_v0p0p1_0.V2.t5 GND 0.648f
C3597 resistorDivider_v0p0p1_0.V2.t9 GND 0.301f
C3598 resistorDivider_v0p0p1_0.V2.n2 GND 0.372f
C3599 resistorDivider_v0p0p1_0.V2.n3 GND 0.369f
C3600 resistorDivider_v0p0p1_0.V2.n4 GND 0.369f
C3601 resistorDivider_v0p0p1_0.V2.n5 GND 0.369f
C3602 resistorDivider_v0p0p1_0.V2.n6 GND 0.369f
C3603 resistorDivider_v0p0p1_0.V2.n7 GND 0.369f
C3604 resistorDivider_v0p0p1_0.V2.n8 GND 0.369f
C3605 resistorDivider_v0p0p1_0.V2.n9 GND 0.369f
C3606 resistorDivider_v0p0p1_0.V2.n10 GND 0.369f
C3607 resistorDivider_v0p0p1_0.V2.n11 GND 0.369f
C3608 resistorDivider_v0p0p1_0.V2.n12 GND 0.369f
C3609 resistorDivider_v0p0p1_0.V2.n13 GND 0.369f
C3610 resistorDivider_v0p0p1_0.V2.n14 GND 0.369f
C3611 resistorDivider_v0p0p1_0.V2.t0 GND 0.164f
C3612 resistorDivider_v0p0p1_0.V2.n15 GND 0.505f
C3613 resistorDivider_v0p0p1_0.V2.n16 GND 0.283f
C3614 resistorDivider_v0p0p1_0.V10.t17 GND 0.0223f
C3615 resistorDivider_v0p0p1_0.V10.n0 GND 0.183f
C3616 resistorDivider_v0p0p1_0.V10.n1 GND 0.0923f
C3617 resistorDivider_v0p0p1_0.V10.t1 GND 0.292f
C3618 resistorDivider_v0p0p1_0.V10.t6 GND 0.292f
C3619 resistorDivider_v0p0p1_0.V10.t11 GND 0.292f
C3620 resistorDivider_v0p0p1_0.V10.t2 GND 0.292f
C3621 resistorDivider_v0p0p1_0.V10.t15 GND 0.292f
C3622 resistorDivider_v0p0p1_0.V10.t4 GND 0.292f
C3623 resistorDivider_v0p0p1_0.V10.t7 GND 0.292f
C3624 resistorDivider_v0p0p1_0.V10.t14 GND 0.292f
C3625 resistorDivider_v0p0p1_0.V10.t9 GND 0.292f
C3626 resistorDivider_v0p0p1_0.V10.t10 GND 0.292f
C3627 resistorDivider_v0p0p1_0.V10.t12 GND 0.292f
C3628 resistorDivider_v0p0p1_0.V10.t3 GND 0.292f
C3629 resistorDivider_v0p0p1_0.V10.t13 GND 0.292f
C3630 resistorDivider_v0p0p1_0.V10.t5 GND 0.292f
C3631 resistorDivider_v0p0p1_0.V10.t8 GND 0.292f
C3632 resistorDivider_v0p0p1_0.V10.t0 GND 0.16f
C3633 resistorDivider_v0p0p1_0.V10.n2 GND 0.831f
C3634 resistorDivider_v0p0p1_0.V10.n3 GND 0.717f
C3635 resistorDivider_v0p0p1_0.V10.n4 GND 0.717f
C3636 resistorDivider_v0p0p1_0.V10.n5 GND 0.717f
C3637 resistorDivider_v0p0p1_0.V10.n6 GND 0.717f
C3638 resistorDivider_v0p0p1_0.V10.n7 GND 0.717f
C3639 resistorDivider_v0p0p1_0.V10.n8 GND 0.717f
C3640 resistorDivider_v0p0p1_0.V10.n9 GND 0.648f
C3641 resistorDivider_v0p0p1_0.V11.t16 GND 0.0237f
C3642 resistorDivider_v0p0p1_0.V11.n0 GND 0.194f
C3643 resistorDivider_v0p0p1_0.V11.n1 GND 0.0938f
C3644 resistorDivider_v0p0p1_0.V11.t14 GND 0.309f
C3645 resistorDivider_v0p0p1_0.V11.t6 GND 0.309f
C3646 resistorDivider_v0p0p1_0.V11.t5 GND 0.309f
C3647 resistorDivider_v0p0p1_0.V11.t1 GND 0.309f
C3648 resistorDivider_v0p0p1_0.V11.t9 GND 0.309f
C3649 resistorDivider_v0p0p1_0.V11.t3 GND 0.309f
C3650 resistorDivider_v0p0p1_0.V11.t15 GND 0.309f
C3651 resistorDivider_v0p0p1_0.V11.t12 GND 0.309f
C3652 resistorDivider_v0p0p1_0.V11.t13 GND 0.309f
C3653 resistorDivider_v0p0p1_0.V11.t10 GND 0.309f
C3654 resistorDivider_v0p0p1_0.V11.t2 GND 0.309f
C3655 resistorDivider_v0p0p1_0.V11.t8 GND 0.309f
C3656 resistorDivider_v0p0p1_0.V11.t4 GND 0.309f
C3657 resistorDivider_v0p0p1_0.V11.t7 GND 0.309f
C3658 resistorDivider_v0p0p1_0.V11.t11 GND 0.666f
C3659 resistorDivider_v0p0p1_0.V11.n2 GND 0.383f
C3660 resistorDivider_v0p0p1_0.V11.n3 GND 0.38f
C3661 resistorDivider_v0p0p1_0.V11.n4 GND 0.38f
C3662 resistorDivider_v0p0p1_0.V11.n5 GND 0.38f
C3663 resistorDivider_v0p0p1_0.V11.n6 GND 0.38f
C3664 resistorDivider_v0p0p1_0.V11.n7 GND 0.38f
C3665 resistorDivider_v0p0p1_0.V11.n8 GND 0.38f
C3666 resistorDivider_v0p0p1_0.V11.n9 GND 0.38f
C3667 resistorDivider_v0p0p1_0.V11.t0 GND 0.169f
C3668 resistorDivider_v0p0p1_0.V11.n10 GND 0.52f
C3669 resistorDivider_v0p0p1_0.V11.n11 GND 0.38f
C3670 resistorDivider_v0p0p1_0.V11.n12 GND 0.38f
C3671 resistorDivider_v0p0p1_0.V11.n13 GND 0.38f
C3672 resistorDivider_v0p0p1_0.V11.n14 GND 0.38f
C3673 resistorDivider_v0p0p1_0.V11.n15 GND 0.38f
C3674 resistorDivider_v0p0p1_0.V11.n16 GND 0.307f
C3675 frontAnalog_v0p0p1_5.RSfetsym_0.QN.t2 GND 0.0322f
C3676 frontAnalog_v0p0p1_5.RSfetsym_0.QN.t1 GND 0.0322f
C3677 frontAnalog_v0p0p1_5.RSfetsym_0.QN.n0 GND 0.136f
C3678 frontAnalog_v0p0p1_5.RSfetsym_0.QN.t6 GND 0.0321f
C3679 frontAnalog_v0p0p1_5.RSfetsym_0.QN.t5 GND 0.0947f
C3680 frontAnalog_v0p0p1_5.RSfetsym_0.QN.n1 GND 1.46f
C3681 frontAnalog_v0p0p1_5.RSfetsym_0.QN.n2 GND 0.0784f
C3682 frontAnalog_v0p0p1_5.RSfetsym_0.QN.n3 GND 0.102f
C3683 frontAnalog_v0p0p1_5.RSfetsym_0.QN.n4 GND 0.445f
C3684 frontAnalog_v0p0p1_5.RSfetsym_0.QN.n5 GND 0.0126f
C3685 frontAnalog_v0p0p1_5.RSfetsym_0.QN.n6 GND 0.0341f
C3686 frontAnalog_v0p0p1_5.RSfetsym_0.QN.t4 GND 0.0322f
C3687 frontAnalog_v0p0p1_5.RSfetsym_0.QN.n7 GND 0.107f
C3688 frontAnalog_v0p0p1_5.RSfetsym_0.QN.n8 GND 0.131f
C3689 frontAnalog_v0p0p1_5.RSfetsym_0.QN.n9 GND 0.351f
C3690 frontAnalog_v0p0p1_5.RSfetsym_0.QN.n10 GND 0.871f
C3691 frontAnalog_v0p0p1_5.RSfetsym_0.QN.t3 GND 0.0566f
C3692 frontAnalog_v0p0p1_5.RSfetsym_0.QN.n11 GND 2.48f
C3693 frontAnalog_v0p0p1_14.x65.A.n0 GND 0.139f
C3694 frontAnalog_v0p0p1_14.x65.A.t7 GND 0.028f
C3695 frontAnalog_v0p0p1_14.x65.A.t4 GND 0.0175f
C3696 frontAnalog_v0p0p1_14.x65.A.n1 GND 0.0568f
C3697 frontAnalog_v0p0p1_14.x65.A.t2 GND 0.149f
C3698 frontAnalog_v0p0p1_14.x65.A.t5 GND 0.0318f
C3699 frontAnalog_v0p0p1_14.x65.A.t3 GND 0.141f
C3700 frontAnalog_v0p0p1_14.x65.A.t6 GND 0.219f
C3701 frontAnalog_v0p0p1_14.x65.A.n2 GND 1.37f
C3702 frontAnalog_v0p0p1_14.x65.A.n3 GND 0.898f
C3703 frontAnalog_v0p0p1_14.x65.A.t1 GND 0.463f
C3704 frontAnalog_v0p0p1_14.x65.A.t0 GND 0.0194f
C3705 frontAnalog_v0p0p1_14.x65.A.n4 GND 1.6f
C3706 frontAnalog_v0p0p1_14.x65.A.n5 GND 2.01f
C3707 frontAnalog_v0p0p1_14.x65.A.n6 GND 1.72f
C3708 frontAnalog_v0p0p1_14.x63.A.n0 GND 0.12f
C3709 frontAnalog_v0p0p1_14.x63.A.n1 GND 2.22f
C3710 frontAnalog_v0p0p1_14.x63.A.t5 GND 0.014f
C3711 frontAnalog_v0p0p1_14.x63.A.t7 GND 0.0225f
C3712 frontAnalog_v0p0p1_14.x63.A.n2 GND 0.0465f
C3713 frontAnalog_v0p0p1_14.x63.A.t1 GND 0.151f
C3714 frontAnalog_v0p0p1_14.x63.A.t2 GND 0.0156f
C3715 frontAnalog_v0p0p1_14.x63.A.t3 GND 0.335f
C3716 frontAnalog_v0p0p1_14.x63.A.t4 GND 0.0256f
C3717 frontAnalog_v0p0p1_14.x63.A.t0 GND 0.173f
C3718 frontAnalog_v0p0p1_14.x63.A.t6 GND 0.175f
C3719 frontAnalog_v0p0p1_14.x63.A.n3 GND 1f
C3720 frontAnalog_v0p0p1_14.x63.A.n4 GND 0.953f
C3721 frontAnalog_v0p0p1_14.x63.A.n5 GND 1.25f
C3722 resistorDivider_v0p0p1_0.V3.t16 GND 0.0237f
C3723 resistorDivider_v0p0p1_0.V3.n0 GND 0.194f
C3724 resistorDivider_v0p0p1_0.V3.n1 GND 0.094f
C3725 resistorDivider_v0p0p1_0.V3.t4 GND 0.31f
C3726 resistorDivider_v0p0p1_0.V3.t3 GND 0.31f
C3727 resistorDivider_v0p0p1_0.V3.t15 GND 0.31f
C3728 resistorDivider_v0p0p1_0.V3.t6 GND 0.31f
C3729 resistorDivider_v0p0p1_0.V3.t13 GND 0.31f
C3730 resistorDivider_v0p0p1_0.V3.t7 GND 0.31f
C3731 resistorDivider_v0p0p1_0.V3.t5 GND 0.31f
C3732 resistorDivider_v0p0p1_0.V3.t11 GND 0.31f
C3733 resistorDivider_v0p0p1_0.V3.t8 GND 0.31f
C3734 resistorDivider_v0p0p1_0.V3.t12 GND 0.31f
C3735 resistorDivider_v0p0p1_0.V3.t9 GND 0.31f
C3736 resistorDivider_v0p0p1_0.V3.t14 GND 0.31f
C3737 resistorDivider_v0p0p1_0.V3.t2 GND 0.31f
C3738 resistorDivider_v0p0p1_0.V3.t10 GND 0.31f
C3739 resistorDivider_v0p0p1_0.V3.t1 GND 0.669f
C3740 resistorDivider_v0p0p1_0.V3.n2 GND 0.384f
C3741 resistorDivider_v0p0p1_0.V3.n3 GND 0.381f
C3742 resistorDivider_v0p0p1_0.V3.n4 GND 0.381f
C3743 resistorDivider_v0p0p1_0.V3.n5 GND 0.381f
C3744 resistorDivider_v0p0p1_0.V3.n6 GND 0.381f
C3745 resistorDivider_v0p0p1_0.V3.n7 GND 0.381f
C3746 resistorDivider_v0p0p1_0.V3.n8 GND 0.381f
C3747 resistorDivider_v0p0p1_0.V3.n9 GND 0.381f
C3748 resistorDivider_v0p0p1_0.V3.n10 GND 0.381f
C3749 resistorDivider_v0p0p1_0.V3.t0 GND 0.17f
C3750 resistorDivider_v0p0p1_0.V3.n11 GND 0.521f
C3751 resistorDivider_v0p0p1_0.V3.n12 GND 0.381f
C3752 resistorDivider_v0p0p1_0.V3.n13 GND 0.381f
C3753 resistorDivider_v0p0p1_0.V3.n14 GND 0.381f
C3754 resistorDivider_v0p0p1_0.V3.n15 GND 0.381f
C3755 resistorDivider_v0p0p1_0.V3.n16 GND 0.301f
C3756 resistorDivider_v0p0p1_0.V4.t16 GND 0.0245f
C3757 resistorDivider_v0p0p1_0.V4.n0 GND 0.201f
C3758 resistorDivider_v0p0p1_0.V4.n1 GND 0.097f
C3759 resistorDivider_v0p0p1_0.V4.t3 GND 0.32f
C3760 resistorDivider_v0p0p1_0.V4.t5 GND 0.32f
C3761 resistorDivider_v0p0p1_0.V4.t7 GND 0.32f
C3762 resistorDivider_v0p0p1_0.V4.t10 GND 0.32f
C3763 resistorDivider_v0p0p1_0.V4.t9 GND 0.32f
C3764 resistorDivider_v0p0p1_0.V4.t8 GND 0.32f
C3765 resistorDivider_v0p0p1_0.V4.t6 GND 0.32f
C3766 resistorDivider_v0p0p1_0.V4.t12 GND 0.32f
C3767 resistorDivider_v0p0p1_0.V4.t2 GND 0.32f
C3768 resistorDivider_v0p0p1_0.V4.t14 GND 0.32f
C3769 resistorDivider_v0p0p1_0.V4.t15 GND 0.32f
C3770 resistorDivider_v0p0p1_0.V4.t4 GND 0.32f
C3771 resistorDivider_v0p0p1_0.V4.t1 GND 0.32f
C3772 resistorDivider_v0p0p1_0.V4.t13 GND 0.32f
C3773 resistorDivider_v0p0p1_0.V4.n2 GND 0.766f
C3774 resistorDivider_v0p0p1_0.V4.n3 GND 0.786f
C3775 resistorDivider_v0p0p1_0.V4.n4 GND 0.786f
C3776 resistorDivider_v0p0p1_0.V4.n5 GND 0.786f
C3777 resistorDivider_v0p0p1_0.V4.n6 GND 0.786f
C3778 resistorDivider_v0p0p1_0.V4.t11 GND 0.32f
C3779 resistorDivider_v0p0p1_0.V4.t0 GND 0.175f
C3780 resistorDivider_v0p0p1_0.V4.n7 GND 0.931f
C3781 resistorDivider_v0p0p1_0.V4.n8 GND 0.786f
C3782 resistorDivider_v0p0p1_0.V4.n9 GND 0.708f
C3783 frontAnalog_v0p0p1_10.x65.A.n0 GND 0.139f
C3784 frontAnalog_v0p0p1_10.x65.A.t4 GND 0.028f
C3785 frontAnalog_v0p0p1_10.x65.A.t6 GND 0.0175f
C3786 frontAnalog_v0p0p1_10.x65.A.n1 GND 0.0568f
C3787 frontAnalog_v0p0p1_10.x65.A.t3 GND 0.149f
C3788 frontAnalog_v0p0p1_10.x65.A.t7 GND 0.0318f
C3789 frontAnalog_v0p0p1_10.x65.A.t2 GND 0.141f
C3790 frontAnalog_v0p0p1_10.x65.A.t5 GND 0.219f
C3791 frontAnalog_v0p0p1_10.x65.A.n2 GND 1.37f
C3792 frontAnalog_v0p0p1_10.x65.A.n3 GND 0.898f
C3793 frontAnalog_v0p0p1_10.x65.A.t0 GND 0.463f
C3794 frontAnalog_v0p0p1_10.x65.A.t1 GND 0.0194f
C3795 frontAnalog_v0p0p1_10.x65.A.n4 GND 1.6f
C3796 frontAnalog_v0p0p1_10.x65.A.n5 GND 2.01f
C3797 frontAnalog_v0p0p1_10.x65.A.n6 GND 1.72f
C3798 CLK.t23 GND 0.0562f
C3799 CLK.t89 GND 0.325f
C3800 CLK.t85 GND 0.329f
C3801 CLK.n1 GND 0.286f
C3802 CLK.t26 GND 0.0592f
C3803 CLK.n2 GND 0.463f
C3804 CLK.n4 GND 0.0676f
C3805 CLK.t94 GND 0.0942f
C3806 CLK.n5 GND 0.395f
C3807 CLK.n6 GND 0.36f
C3808 CLK.n7 GND 0.1f
C3809 CLK.n8 GND 14.1f
C3810 CLK.t58 GND 0.0562f
C3811 CLK.t63 GND 0.325f
C3812 CLK.t14 GND 0.329f
C3813 CLK.n10 GND 0.286f
C3814 CLK.t92 GND 0.0592f
C3815 CLK.n11 GND 0.463f
C3816 CLK.n13 GND 0.0676f
C3817 CLK.t15 GND 0.0942f
C3818 CLK.n14 GND 0.395f
C3819 CLK.n15 GND 0.36f
C3820 CLK.n16 GND 0.1f
C3821 CLK.t17 GND 0.0562f
C3822 CLK.t27 GND 0.325f
C3823 CLK.t73 GND 0.329f
C3824 CLK.n18 GND 0.286f
C3825 CLK.t11 GND 0.0592f
C3826 CLK.n19 GND 0.463f
C3827 CLK.n21 GND 0.0676f
C3828 CLK.t32 GND 0.0942f
C3829 CLK.n22 GND 0.395f
C3830 CLK.n23 GND 0.36f
C3831 CLK.n24 GND 0.1f
C3832 CLK.t35 GND 0.0562f
C3833 CLK.t38 GND 0.325f
C3834 CLK.t90 GND 0.329f
C3835 CLK.n26 GND 0.286f
C3836 CLK.t66 GND 0.0592f
C3837 CLK.n27 GND 0.463f
C3838 CLK.n29 GND 0.0676f
C3839 CLK.t91 GND 0.0942f
C3840 CLK.n30 GND 0.395f
C3841 CLK.n31 GND 0.36f
C3842 CLK.n32 GND 0.1f
C3843 CLK.t45 GND 0.0562f
C3844 CLK.t5 GND 0.325f
C3845 CLK.t47 GND 0.329f
C3846 CLK.n34 GND 0.286f
C3847 CLK.t83 GND 0.0592f
C3848 CLK.n35 GND 0.463f
C3849 CLK.n37 GND 0.0676f
C3850 CLK.t10 GND 0.0942f
C3851 CLK.n38 GND 0.395f
C3852 CLK.n39 GND 0.36f
C3853 CLK.n40 GND 0.104f
C3854 CLK.t4 GND 0.0562f
C3855 CLK.t18 GND 0.325f
C3856 CLK.t64 GND 0.329f
C3857 CLK.n42 GND 0.286f
C3858 CLK.t41 GND 0.0592f
C3859 CLK.n43 GND 0.463f
C3860 CLK.n45 GND 0.0676f
C3861 CLK.t65 GND 0.0942f
C3862 CLK.n46 GND 0.395f
C3863 CLK.n47 GND 0.36f
C3864 CLK.n48 GND 0.1f
C3865 CLK.t25 GND 0.0562f
C3866 CLK.t71 GND 0.325f
C3867 CLK.t74 GND 0.329f
C3868 CLK.n50 GND 0.286f
C3869 CLK.t54 GND 0.0592f
C3870 CLK.n51 GND 0.463f
C3871 CLK.n53 GND 0.0676f
C3872 CLK.t76 GND 0.0942f
C3873 CLK.n54 GND 0.395f
C3874 CLK.n55 GND 0.36f
C3875 CLK.n56 GND 0.1f
C3876 CLK.t79 GND 0.0562f
C3877 CLK.t95 GND 0.325f
C3878 CLK.t39 GND 0.329f
C3879 CLK.n58 GND 0.286f
C3880 CLK.t20 GND 0.0592f
C3881 CLK.n59 GND 0.463f
C3882 CLK.n61 GND 0.0676f
C3883 CLK.t40 GND 0.0942f
C3884 CLK.n62 GND 0.395f
C3885 CLK.n63 GND 0.36f
C3886 CLK.n64 GND 0.1f
C3887 CLK.t2 GND 0.0562f
C3888 CLK.t6 GND 0.325f
C3889 CLK.t51 GND 0.329f
C3890 CLK.n66 GND 0.286f
C3891 CLK.t30 GND 0.0592f
C3892 CLK.n67 GND 0.463f
C3893 CLK.n69 GND 0.0676f
C3894 CLK.t53 GND 0.0942f
C3895 CLK.n70 GND 0.395f
C3896 CLK.n71 GND 0.36f
C3897 CLK.n72 GND 0.1f
C3898 CLK.t56 GND 0.0562f
C3899 CLK.t70 GND 0.325f
C3900 CLK.t13 GND 0.329f
C3901 CLK.n74 GND 0.286f
C3902 CLK.t0 GND 0.0592f
C3903 CLK.n75 GND 0.463f
C3904 CLK.n77 GND 0.0676f
C3905 CLK.t19 GND 0.0942f
C3906 CLK.n78 GND 0.395f
C3907 CLK.n79 GND 0.36f
C3908 CLK.n80 GND 0.1f
C3909 CLK.t69 GND 0.0562f
C3910 CLK.t80 GND 0.325f
C3911 CLK.t28 GND 0.329f
C3912 CLK.n82 GND 0.286f
C3913 CLK.t9 GND 0.0592f
C3914 CLK.n83 GND 0.463f
C3915 CLK.n85 GND 0.0676f
C3916 CLK.t29 GND 0.0942f
C3917 CLK.n86 GND 0.395f
C3918 CLK.n87 GND 0.36f
C3919 CLK.n88 GND 0.1f
C3920 CLK.t33 GND 0.0562f
C3921 CLK.t36 GND 0.325f
C3922 CLK.t87 GND 0.329f
C3923 CLK.n90 GND 0.286f
C3924 CLK.t62 GND 0.0592f
C3925 CLK.n91 GND 0.463f
C3926 CLK.n93 GND 0.0676f
C3927 CLK.t88 GND 0.0942f
C3928 CLK.n94 GND 0.395f
C3929 CLK.n95 GND 0.36f
C3930 CLK.n96 GND 0.1f
C3931 CLK.t44 GND 0.0562f
C3932 CLK.t57 GND 0.325f
C3933 CLK.t7 GND 0.329f
C3934 CLK.n98 GND 0.286f
C3935 CLK.t82 GND 0.0592f
C3936 CLK.n99 GND 0.463f
C3937 CLK.n101 GND 0.0676f
C3938 CLK.t8 GND 0.0942f
C3939 CLK.n102 GND 0.395f
C3940 CLK.n103 GND 0.36f
C3941 CLK.n104 GND 0.1f
C3942 CLK.t12 GND 0.0562f
C3943 CLK.t16 GND 0.325f
C3944 CLK.t60 GND 0.329f
C3945 CLK.n106 GND 0.286f
C3946 CLK.t37 GND 0.0592f
C3947 CLK.n107 GND 0.463f
C3948 CLK.n109 GND 0.0676f
C3949 CLK.t61 GND 0.0942f
C3950 CLK.n110 GND 0.395f
C3951 CLK.n111 GND 0.36f
C3952 CLK.n112 GND 0.104f
C3953 CLK.t24 GND 0.0562f
C3954 CLK.t34 GND 0.325f
C3955 CLK.t72 GND 0.329f
C3956 CLK.n114 GND 0.286f
C3957 CLK.t59 GND 0.0592f
C3958 CLK.n115 GND 0.463f
C3959 CLK.n117 GND 0.0676f
C3960 CLK.t81 GND 0.0942f
C3961 CLK.n118 GND 0.395f
C3962 CLK.n119 GND 0.36f
C3963 CLK.n120 GND 0.104f
C3964 CLK.n121 GND 19.3f
C3965 CLK.n122 GND 12.7f
C3966 CLK.n123 GND 12.8f
C3967 CLK.n124 GND 12.8f
C3968 CLK.n125 GND 12.8f
C3969 CLK.n126 GND 12.7f
C3970 CLK.n127 GND 12.8f
C3971 CLK.n128 GND 12.8f
C3972 CLK.n129 GND 12.8f
C3973 CLK.n130 GND 12.7f
C3974 CLK.n131 GND 12.7f
C3975 CLK.n132 GND 12.8f
C3976 CLK.n133 GND 12.8f
C3977 CLK.n134 GND 12.8f
C3978 CLK.t78 GND 0.0562f
C3979 CLK.t46 GND 0.325f
C3980 CLK.t48 GND 0.329f
C3981 CLK.t86 GND 0.0592f
C3982 CLK.n135 GND 0.463f
C3983 CLK.n137 GND 0.286f
C3984 CLK.n139 GND 0.0676f
C3985 CLK.t49 GND 0.0942f
C3986 CLK.n140 GND 0.395f
C3987 CLK.n141 GND 0.36f
C3988 CLK.n142 GND 0.1f
C3989 a_16719_n13117.n0 GND 1.47f
C3990 a_16719_n13117.n1 GND 1.14f
C3991 a_16719_n13117.t4 GND 0.177f
C3992 a_16719_n13117.t14 GND 0.177f
C3993 a_16719_n13117.t18 GND 0.177f
C3994 a_16719_n13117.t7 GND 0.177f
C3995 a_16719_n13117.t12 GND 0.177f
C3996 a_16719_n13117.t1 GND 0.177f
C3997 a_16719_n13117.t16 GND 0.177f
C3998 a_16719_n13117.t10 GND 0.177f
C3999 a_16719_n13117.t3 GND 0.177f
C4000 a_16719_n13117.t11 GND 0.177f
C4001 a_16719_n13117.t0 GND 0.177f
C4002 a_16719_n13117.t15 GND 0.177f
C4003 a_16719_n13117.t8 GND 0.252f
C4004 a_16719_n13117.n2 GND 1.4f
C4005 a_16719_n13117.n3 GND 0.768f
C4006 a_16719_n13117.n4 GND 0.768f
C4007 a_16719_n13117.n5 GND 0.768f
C4008 a_16719_n13117.n6 GND 0.768f
C4009 a_16719_n13117.n7 GND 0.768f
C4010 a_16719_n13117.n8 GND 0.72f
C4011 a_16719_n13117.n9 GND 0.273f
C4012 a_16719_n13117.n10 GND 0.325f
C4013 a_16719_n13117.n11 GND 0.912f
C4014 a_16719_n13117.n12 GND 2.03f
C4015 a_16719_n13117.n13 GND 1.47f
C4016 a_16719_n13117.t23 GND 0.238f
C4017 a_16719_n13117.n14 GND 2.05f
C4018 a_16719_n13117.t24 GND 1.7f
C4019 a_16719_n13117.n15 GND 0.991f
C4020 a_16719_n13117.n16 GND 0.0433f
C4021 a_16719_n13117.n17 GND 0.426f
C4022 a_16719_n13117.t22 GND 1.7f
C4023 a_16719_n13117.t20 GND 0.0103f
C4024 a_16719_n13117.n18 GND 0.213f
C4025 a_16719_n13117.t25 GND 1.7f
C4026 a_16719_n13117.n19 GND 1.05f
C4027 a_16719_n13117.n20 GND 0.0503f
C4028 a_16719_n13117.n21 GND 0.0699f
C4029 a_16719_n13117.n22 GND 0.308f
C4030 a_16719_n13117.n23 GND 0.811f
C4031 a_16719_n13117.n24 GND 0.768f
C4032 a_16719_n13117.n25 GND 0.768f
C4033 a_16719_n13117.t5 GND 0.177f
C4034 a_16719_n13117.t13 GND 0.177f
C4035 a_16719_n13117.t17 GND 0.177f
C4036 a_16719_n13117.t9 GND 0.177f
C4037 a_16719_n13117.t2 GND 0.177f
C4038 a_16719_n13117.t6 GND 0.252f
C4039 a_16719_n13117.n26 GND 1.4f
C4040 a_16719_n13117.n27 GND 0.768f
C4041 a_16719_n13117.n28 GND 0.768f
C4042 a_16719_n13117.n29 GND 0.768f
C4043 a_16719_n13117.n30 GND 0.768f
C4044 a_16719_n13117.n31 GND 0.768f
C4045 a_16719_n13117.t19 GND 0.177f
C4046 a_16541_n13117.t7 GND 0.112f
C4047 a_16541_n13117.t14 GND 0.112f
C4048 a_16541_n13117.t16 GND 0.112f
C4049 a_16541_n13117.t2 GND 0.112f
C4050 a_16541_n13117.t10 GND 0.112f
C4051 a_16541_n13117.t18 GND 0.112f
C4052 a_16541_n13117.t9 GND 0.112f
C4053 a_16541_n13117.t3 GND 0.112f
C4054 a_16541_n13117.t17 GND 0.112f
C4055 a_16541_n13117.t12 GND 0.112f
C4056 a_16541_n13117.t1 GND 0.112f
C4057 a_16541_n13117.t6 GND 0.112f
C4058 a_16541_n13117.t5 GND 0.112f
C4059 a_16541_n13117.t15 GND 0.112f
C4060 a_16541_n13117.t8 GND 0.112f
C4061 a_16541_n13117.t0 GND 0.112f
C4062 a_16541_n13117.t19 GND 0.112f
C4063 a_16541_n13117.t4 GND 0.112f
C4064 a_16541_n13117.t13 GND 0.161f
C4065 a_16541_n13117.n0 GND 1.02f
C4066 a_16541_n13117.n1 GND 0.558f
C4067 a_16541_n13117.n2 GND 0.558f
C4068 a_16541_n13117.n3 GND 0.558f
C4069 a_16541_n13117.n4 GND 0.558f
C4070 a_16541_n13117.n5 GND 0.558f
C4071 a_16541_n13117.n6 GND 0.558f
C4072 a_16541_n13117.n7 GND 0.558f
C4073 a_16541_n13117.n8 GND 0.614f
C4074 a_16541_n13117.n9 GND 0.614f
C4075 a_16541_n13117.n10 GND 0.558f
C4076 a_16541_n13117.n11 GND 0.558f
C4077 a_16541_n13117.n12 GND 0.558f
C4078 a_16541_n13117.n13 GND 0.558f
C4079 a_16541_n13117.n14 GND 0.558f
C4080 a_16541_n13117.n15 GND 0.558f
C4081 a_16541_n13117.n16 GND 0.554f
C4082 a_16541_n13117.n17 GND 0.627f
C4083 a_16541_n13117.t11 GND 0.127f
C4084 a_16541_n13117.n18 GND 1.13f
C4085 a_16541_n13117.t21 GND 0.376f
C4086 a_16541_n13117.n19 GND 10.1f
C4087 a_16541_n13117.t20 GND 1.21f
C4088 a_16599_n13205.n0 GND 0.681f
C4089 a_16599_n13205.t15 GND 0.179f
C4090 a_16599_n13205.n1 GND 0.251f
C4091 a_16599_n13205.t8 GND 0.179f
C4092 a_16599_n13205.n2 GND 0.378f
C4093 a_16599_n13205.t23 GND 0.179f
C4094 a_16599_n13205.n3 GND 0.197f
C4095 a_16599_n13205.t12 GND 0.179f
C4096 a_16599_n13205.n4 GND 0.197f
C4097 a_16599_n13205.t20 GND 0.179f
C4098 a_16599_n13205.n5 GND 0.197f
C4099 a_16599_n13205.t13 GND 0.179f
C4100 a_16599_n13205.n6 GND 0.197f
C4101 a_16599_n13205.t7 GND 0.179f
C4102 a_16599_n13205.n7 GND 0.197f
C4103 a_16599_n13205.t22 GND 0.179f
C4104 a_16599_n13205.n8 GND 0.197f
C4105 a_16599_n13205.t11 GND 0.179f
C4106 a_16599_n13205.n9 GND 0.197f
C4107 a_16599_n13205.t16 GND 0.179f
C4108 a_16599_n13205.n10 GND 0.184f
C4109 a_16599_n13205.t0 GND 0.179f
C4110 a_16599_n13205.t5 GND 0.179f
C4111 a_16599_n13205.t9 GND 0.179f
C4112 a_16599_n13205.t19 GND 0.179f
C4113 a_16599_n13205.t4 GND 0.179f
C4114 a_16599_n13205.t18 GND 0.179f
C4115 a_16599_n13205.t10 GND 0.179f
C4116 a_16599_n13205.t6 GND 0.179f
C4117 a_16599_n13205.t14 GND 0.179f
C4118 a_16599_n13205.t21 GND 0.179f
C4119 a_16599_n13205.t17 GND 0.179f
C4120 a_16599_n13205.n11 GND 0.252f
C4121 a_16599_n13205.n12 GND 0.376f
C4122 a_16599_n13205.n13 GND 0.197f
C4123 a_16599_n13205.n14 GND 0.197f
C4124 a_16599_n13205.n15 GND 0.197f
C4125 a_16599_n13205.n16 GND 0.197f
C4126 a_16599_n13205.n17 GND 0.197f
C4127 a_16599_n13205.n18 GND 0.197f
C4128 a_16599_n13205.n19 GND 0.197f
C4129 a_16599_n13205.n20 GND 0.197f
C4130 a_16599_n13205.n21 GND 0.169f
C4131 a_16599_n13205.n22 GND 0.102f
C4132 a_16599_n13205.n23 GND 0.377f
C4133 a_16599_n13205.n24 GND 0.197f
C4134 a_16599_n13205.n25 GND 0.197f
C4135 a_16599_n13205.n26 GND 0.197f
C4136 a_16599_n13205.n27 GND 0.197f
C4137 a_16599_n13205.n28 GND 0.197f
C4138 a_16599_n13205.n29 GND 0.197f
C4139 a_16599_n13205.n30 GND 0.197f
C4140 a_16599_n13205.n31 GND 0.184f
C4141 a_16599_n13205.n32 GND 0.376f
C4142 a_16599_n13205.n33 GND 0.197f
C4143 a_16599_n13205.n34 GND 0.197f
C4144 a_16599_n13205.n35 GND 0.197f
C4145 a_16599_n13205.n36 GND 0.197f
C4146 a_16599_n13205.n37 GND 0.197f
C4147 a_16599_n13205.n38 GND 0.197f
C4148 a_16599_n13205.n39 GND 0.197f
C4149 a_16599_n13205.n40 GND 0.197f
C4150 a_16599_n13205.n41 GND 0.169f
C4151 a_16599_n13205.n42 GND 0.108f
C4152 a_16599_n13205.t1 GND 0.0381f
C4153 a_16599_n13205.n43 GND 2.83f
C4154 a_16599_n13205.t3 GND 1.94f
C4155 resistorDivider_v0p0p1_0.V16.t16 GND 0.0223f
C4156 resistorDivider_v0p0p1_0.V16.n0 GND 0.183f
C4157 resistorDivider_v0p0p1_0.V16.n1 GND 0.077f
C4158 resistorDivider_v0p0p1_0.V16.t13 GND 0.292f
C4159 resistorDivider_v0p0p1_0.V16.t1 GND 0.292f
C4160 resistorDivider_v0p0p1_0.V16.t10 GND 0.292f
C4161 resistorDivider_v0p0p1_0.V16.t12 GND 0.292f
C4162 resistorDivider_v0p0p1_0.V16.t4 GND 0.292f
C4163 resistorDivider_v0p0p1_0.V16.t14 GND 0.292f
C4164 resistorDivider_v0p0p1_0.V16.t6 GND 0.292f
C4165 resistorDivider_v0p0p1_0.V16.t15 GND 0.292f
C4166 resistorDivider_v0p0p1_0.V16.t9 GND 0.292f
C4167 resistorDivider_v0p0p1_0.V16.t3 GND 0.292f
C4168 resistorDivider_v0p0p1_0.V16.t2 GND 0.292f
C4169 resistorDivider_v0p0p1_0.V16.t8 GND 0.292f
C4170 resistorDivider_v0p0p1_0.V16.t11 GND 0.292f
C4171 resistorDivider_v0p0p1_0.V16.t5 GND 0.292f
C4172 resistorDivider_v0p0p1_0.V16.t7 GND 0.629f
C4173 resistorDivider_v0p0p1_0.V16.n2 GND 0.362f
C4174 resistorDivider_v0p0p1_0.V16.n3 GND 0.359f
C4175 resistorDivider_v0p0p1_0.V16.n4 GND 0.359f
C4176 resistorDivider_v0p0p1_0.V16.t0 GND 0.16f
C4177 resistorDivider_v0p0p1_0.V16.n5 GND 0.491f
C4178 resistorDivider_v0p0p1_0.V16.n6 GND 0.359f
C4179 resistorDivider_v0p0p1_0.V16.n7 GND 0.359f
C4180 resistorDivider_v0p0p1_0.V16.n8 GND 0.359f
C4181 resistorDivider_v0p0p1_0.V16.n9 GND 0.359f
C4182 resistorDivider_v0p0p1_0.V16.n10 GND 0.359f
C4183 resistorDivider_v0p0p1_0.V16.n11 GND 0.359f
C4184 resistorDivider_v0p0p1_0.V16.n12 GND 0.359f
C4185 resistorDivider_v0p0p1_0.V16.n13 GND 0.359f
C4186 resistorDivider_v0p0p1_0.V16.n14 GND 0.359f
C4187 resistorDivider_v0p0p1_0.V16.n15 GND 0.359f
C4188 resistorDivider_v0p0p1_0.V16.n16 GND 0.291f
C4189 VFS.t7 GND 0.108f
C4190 VFS.n0 GND 0.0961f
C4191 VFS.n1 GND 0.0961f
C4192 VFS.n2 GND 0.0687f
C4193 VFS.n3 GND 2.49f
C4194 VFS.t2 GND 0.0898f
C4195 VFS.n4 GND 0.0961f
C4196 VFS.n5 GND 0.0961f
C4197 VFS.n6 GND 0.0741f
C4198 OUT2.n2 GND 0.0114f
C4199 OUT2.n4 GND 0.0241f
C4200 OUT2.n6 GND 0.0161f
C4201 OUT2.n8 GND 0.0161f
C4202 OUT2.n10 GND 0.0161f
C4203 OUT2.n12 GND 0.0161f
C4204 OUT2.n14 GND 0.0161f
C4205 OUT2.n23 GND 0.014f
C4206 OUT2.n25 GND 0.0348f
C4207 OUT2.n27 GND 0.021f
C4208 OUT2.n29 GND 0.021f
C4209 OUT2.n31 GND 0.021f
C4210 OUT2.n33 GND 0.021f
C4211 OUT2.n35 GND 0.021f
C4212 OUT2.n37 GND 0.0147f
C4213 OUT2.n38 GND 0.0296f
C4214 OUT2.n39 GND 0.0229f
C4215 OUT2.n42 GND 0.0114f
C4216 OUT2.n44 GND 0.0241f
C4217 OUT2.n46 GND 0.0161f
C4218 OUT2.n48 GND 0.0161f
C4219 OUT2.n50 GND 0.0161f
C4220 OUT2.n52 GND 0.0161f
C4221 OUT2.n54 GND 0.0161f
C4222 OUT2.n63 GND 0.014f
C4223 OUT2.n65 GND 0.0348f
C4224 OUT2.n67 GND 0.021f
C4225 OUT2.n69 GND 0.021f
C4226 OUT2.n71 GND 0.021f
C4227 OUT2.n73 GND 0.021f
C4228 OUT2.n75 GND 0.021f
C4229 OUT2.n77 GND 0.0147f
C4230 OUT2.n78 GND 0.0273f
C4231 OUT2.n79 GND 0.0203f
C4232 OUT2.n81 GND 0.0114f
C4233 OUT2.n83 GND 0.0241f
C4234 OUT2.n85 GND 0.0161f
C4235 OUT2.n87 GND 0.0161f
C4236 OUT2.n89 GND 0.0161f
C4237 OUT2.n91 GND 0.0161f
C4238 OUT2.n93 GND 0.0161f
C4239 OUT2.n97 GND 0.0126f
C4240 OUT2.n100 GND 0.014f
C4241 OUT2.n102 GND 0.0348f
C4242 OUT2.n104 GND 0.021f
C4243 OUT2.n106 GND 0.021f
C4244 OUT2.n108 GND 0.021f
C4245 OUT2.n110 GND 0.021f
C4246 OUT2.n112 GND 0.021f
C4247 OUT2.n114 GND 0.0147f
C4248 OUT2.n115 GND 0.0284f
C4249 OUT2.n116 GND 0.0234f
C4250 OUT2.n120 GND 0.014f
C4251 OUT2.n122 GND 0.0348f
C4252 OUT2.n124 GND 0.021f
C4253 OUT2.n126 GND 0.021f
C4254 OUT2.n128 GND 0.021f
C4255 OUT2.n130 GND 0.021f
C4256 OUT2.n132 GND 0.021f
C4257 OUT2.n136 GND 0.0114f
C4258 OUT2.n138 GND 0.0241f
C4259 OUT2.n140 GND 0.0161f
C4260 OUT2.n142 GND 0.0161f
C4261 OUT2.n144 GND 0.0161f
C4262 OUT2.n146 GND 0.0161f
C4263 OUT2.n148 GND 0.0161f
C4264 OUT2.n152 GND 0.013f
C4265 OUT2.n155 GND 0.0204f
C4266 OUT2.n156 GND 0.108f
C4267 OUT2.n157 GND 0.275f
C4268 OUT2.n158 GND 0.224f
C4269 OUT2.n159 GND 0.228f
C4270 frontAnalog_v0p0p1_10.Q.t11 GND 0.0123f
C4271 frontAnalog_v0p0p1_10.Q.n0 GND 0.0135f
C4272 frontAnalog_v0p0p1_10.Q.n8 GND 0.15f
C4273 frontAnalog_v0p0p1_10.Q.n9 GND 0.374f
C4274 frontAnalog_v0p0p1_10.Q.n12 GND 0.0114f
C4275 frontAnalog_v0p0p1_10.Q.n16 GND 0.213f
C4276 frontAnalog_v0p0p1_10.Q.n21 GND 0.567f
C4277 frontAnalog_v0p0p1_10.Q.n22 GND 1.34f
C4278 frontAnalog_v0p0p1_10.Q.n23 GND 0.305f
C4279 frontAnalog_v0p0p1_10.Q.n24 GND 0.686f
C4280 frontAnalog_v0p0p1_10.Q.n25 GND 7.69f
C4281 frontAnalog_v0p0p1_10.Q.t12 GND 0.0276f
C4282 frontAnalog_v0p0p1_10.Q.n26 GND 0.432f
C4283 frontAnalog_v0p0p1_10.Q.n27 GND 0.13f
C4284 frontAnalog_v0p0p1_10.Q.n28 GND 0.0573f
C4285 frontAnalog_v0p0p1_10.Q.n29 GND 0.0862f
C4286 frontAnalog_v0p0p1_10.Q.n30 GND 0.0921f
C4287 frontAnalog_v0p0p1_10.Q.n31 GND 0.127f
C4288 frontAnalog_v0p0p1_10.Q.n32 GND 0.12f
C4289 frontAnalog_v0p0p1_10.Q.t3 GND 0.0102f
C4290 frontAnalog_v0p0p1_10.Q.n33 GND 0.276f
C4291 frontAnalog_v0p0p1_10.Q.n34 GND 12.4f
C4292 OUT0.n2 GND 0.0114f
C4293 OUT0.n4 GND 0.0241f
C4294 OUT0.n6 GND 0.0161f
C4295 OUT0.n8 GND 0.0161f
C4296 OUT0.n10 GND 0.0161f
C4297 OUT0.n12 GND 0.0161f
C4298 OUT0.n14 GND 0.0161f
C4299 OUT0.n23 GND 0.014f
C4300 OUT0.n25 GND 0.0348f
C4301 OUT0.n27 GND 0.021f
C4302 OUT0.n29 GND 0.021f
C4303 OUT0.n31 GND 0.021f
C4304 OUT0.n33 GND 0.021f
C4305 OUT0.n35 GND 0.021f
C4306 OUT0.n37 GND 0.0147f
C4307 OUT0.n38 GND 0.0296f
C4308 OUT0.n39 GND 0.0229f
C4309 OUT0.n42 GND 0.0114f
C4310 OUT0.n44 GND 0.0241f
C4311 OUT0.n46 GND 0.0161f
C4312 OUT0.n48 GND 0.0161f
C4313 OUT0.n50 GND 0.0161f
C4314 OUT0.n52 GND 0.0161f
C4315 OUT0.n54 GND 0.0161f
C4316 OUT0.n63 GND 0.014f
C4317 OUT0.n65 GND 0.0348f
C4318 OUT0.n67 GND 0.021f
C4319 OUT0.n69 GND 0.021f
C4320 OUT0.n71 GND 0.021f
C4321 OUT0.n73 GND 0.021f
C4322 OUT0.n75 GND 0.021f
C4323 OUT0.n77 GND 0.0147f
C4324 OUT0.n78 GND 0.0273f
C4325 OUT0.n79 GND 0.0203f
C4326 OUT0.n81 GND 0.0114f
C4327 OUT0.n83 GND 0.0241f
C4328 OUT0.n85 GND 0.0161f
C4329 OUT0.n87 GND 0.0161f
C4330 OUT0.n89 GND 0.0161f
C4331 OUT0.n91 GND 0.0161f
C4332 OUT0.n93 GND 0.0161f
C4333 OUT0.n97 GND 0.0126f
C4334 OUT0.n100 GND 0.014f
C4335 OUT0.n102 GND 0.0348f
C4336 OUT0.n104 GND 0.021f
C4337 OUT0.n106 GND 0.021f
C4338 OUT0.n108 GND 0.021f
C4339 OUT0.n110 GND 0.021f
C4340 OUT0.n112 GND 0.021f
C4341 OUT0.n114 GND 0.0147f
C4342 OUT0.n115 GND 0.0284f
C4343 OUT0.n116 GND 0.0234f
C4344 OUT0.n120 GND 0.014f
C4345 OUT0.n122 GND 0.0348f
C4346 OUT0.n124 GND 0.021f
C4347 OUT0.n126 GND 0.021f
C4348 OUT0.n128 GND 0.021f
C4349 OUT0.n130 GND 0.021f
C4350 OUT0.n132 GND 0.021f
C4351 OUT0.n136 GND 0.0114f
C4352 OUT0.n138 GND 0.0241f
C4353 OUT0.n140 GND 0.0161f
C4354 OUT0.n142 GND 0.0161f
C4355 OUT0.n144 GND 0.0161f
C4356 OUT0.n146 GND 0.0161f
C4357 OUT0.n148 GND 0.0161f
C4358 OUT0.n152 GND 0.013f
C4359 OUT0.n155 GND 0.0204f
C4360 OUT0.n156 GND 0.108f
C4361 OUT0.n157 GND 0.275f
C4362 OUT0.n158 GND 0.224f
C4363 OUT0.n159 GND 0.228f
C4364 frontAnalog_v0p0p1_15.x63.A.n0 GND 0.12f
C4365 frontAnalog_v0p0p1_15.x63.A.n1 GND 2.22f
C4366 frontAnalog_v0p0p1_15.x63.A.t6 GND 0.014f
C4367 frontAnalog_v0p0p1_15.x63.A.t4 GND 0.0225f
C4368 frontAnalog_v0p0p1_15.x63.A.n2 GND 0.0465f
C4369 frontAnalog_v0p0p1_15.x63.A.t3 GND 0.151f
C4370 frontAnalog_v0p0p1_15.x63.A.t2 GND 0.0156f
C4371 frontAnalog_v0p0p1_15.x63.A.t1 GND 0.335f
C4372 frontAnalog_v0p0p1_15.x63.A.t5 GND 0.0256f
C4373 frontAnalog_v0p0p1_15.x63.A.t0 GND 0.173f
C4374 frontAnalog_v0p0p1_15.x63.A.t7 GND 0.175f
C4375 frontAnalog_v0p0p1_15.x63.A.n3 GND 1f
C4376 frontAnalog_v0p0p1_15.x63.A.n4 GND 0.953f
C4377 frontAnalog_v0p0p1_15.x63.A.n5 GND 1.25f
C4378 OUT3.n5 GND 0.0122f
C4379 OUT3.n7 GND 0.0305f
C4380 OUT3.n9 GND 0.0184f
C4381 OUT3.n11 GND 0.0184f
C4382 OUT3.n13 GND 0.0184f
C4383 OUT3.n15 GND 0.0184f
C4384 OUT3.n17 GND 0.0184f
C4385 OUT3.n26 GND 0.0212f
C4386 OUT3.n28 GND 0.0141f
C4387 OUT3.n30 GND 0.0141f
C4388 OUT3.n32 GND 0.0141f
C4389 OUT3.n34 GND 0.0141f
C4390 OUT3.n36 GND 0.0141f
C4391 OUT3.n44 GND 0.027f
C4392 OUT3.n45 GND 0.0219f
C4393 OUT3.n51 GND 0.0122f
C4394 OUT3.n53 GND 0.0305f
C4395 OUT3.n55 GND 0.0184f
C4396 OUT3.n57 GND 0.0184f
C4397 OUT3.n59 GND 0.0184f
C4398 OUT3.n61 GND 0.0184f
C4399 OUT3.n63 GND 0.0184f
C4400 OUT3.n66 GND 0.0157f
C4401 OUT3.n72 GND 0.0212f
C4402 OUT3.n74 GND 0.0141f
C4403 OUT3.n76 GND 0.0141f
C4404 OUT3.n78 GND 0.0141f
C4405 OUT3.n80 GND 0.0141f
C4406 OUT3.n82 GND 0.0141f
C4407 OUT3.n85 GND 0.015f
C4408 OUT3.n86 GND 0.0477f
C4409 OUT3.n87 GND 0.0111f
C4410 OUT3.n89 GND 0.0122f
C4411 OUT3.n91 GND 0.0305f
C4412 OUT3.n93 GND 0.0184f
C4413 OUT3.n95 GND 0.0184f
C4414 OUT3.n97 GND 0.0184f
C4415 OUT3.n99 GND 0.0184f
C4416 OUT3.n101 GND 0.0184f
C4417 OUT3.n114 GND 0.0212f
C4418 OUT3.n116 GND 0.0141f
C4419 OUT3.n118 GND 0.0141f
C4420 OUT3.n120 GND 0.0141f
C4421 OUT3.n122 GND 0.0141f
C4422 OUT3.n124 GND 0.0141f
C4423 OUT3.n133 GND 0.0282f
C4424 OUT3.n134 GND 0.0213f
C4425 OUT3.n140 GND 0.0122f
C4426 OUT3.n142 GND 0.0305f
C4427 OUT3.n144 GND 0.0184f
C4428 OUT3.n146 GND 0.0184f
C4429 OUT3.n148 GND 0.0184f
C4430 OUT3.n150 GND 0.0184f
C4431 OUT3.n152 GND 0.0184f
C4432 OUT3.n160 GND 0.0212f
C4433 OUT3.n162 GND 0.0141f
C4434 OUT3.n164 GND 0.0141f
C4435 OUT3.n166 GND 0.0141f
C4436 OUT3.n168 GND 0.0141f
C4437 OUT3.n170 GND 0.0141f
C4438 OUT3.n179 GND 0.027f
C4439 OUT3.n180 GND 0.119f
C4440 OUT3.n181 GND 0.304f
C4441 OUT3.n182 GND 0.264f
C4442 OUT3.n183 GND 0.577f
C4443 VDD.t216 GND 0.0126f
C4444 VDD.t808 GND 0.0124f
C4445 VDD.t699 GND 0.0104f
C4446 VDD.t232 GND 0.0129f
C4447 VDD.t150 GND 0.0134f
C4448 VDD.t1381 GND 0.0107f
C4449 VDD.t810 GND 0.0281f
C4450 VDD.t139 GND 0.0485f
C4451 VDD.t1339 GND 0.0199f
C4452 VDD.t205 GND 0.0209f
C4453 VDD.t867 GND 0.0209f
C4454 VDD.t157 GND 0.0241f
C4455 VDD.t820 GND 0.0392f
C4456 VDD.n0 GND 0.0192f
C4457 VDD.n26 GND 0.0309f
C4458 VDD.n28 GND 0.013f
C4459 VDD.n33 GND 0.0119f
C4460 VDD.n34 GND 0.119f
C4461 VDD.n35 GND 0.374f
C4462 VDD.n59 GND 0.0109f
C4463 VDD.t155 GND 0.115f
C4464 VDD.t145 GND 0.0557f
C4465 VDD.t159 GND 0.117f
C4466 VDD.t33 GND 0.0441f
C4467 VDD.n60 GND 0.0473f
C4468 VDD.n61 GND 0.0681f
C4469 VDD.n62 GND 0.734f
C4470 VDD.t415 GND 0.0191f
C4471 VDD.t850 GND 0.0128f
C4472 VDD.t206 GND 0.0119f
C4473 VDD.t754 GND 0.0133f
C4474 VDD.t143 GND 0.0122f
C4475 VDD.t791 GND 0.011f
C4476 VDD.t853 GND 0.0158f
C4477 VDD.t747 GND 0.0129f
C4478 VDD.t770 GND 0.0159f
C4479 VDD.t1484 GND 0.0246f
C4480 VDD.t751 GND 0.0353f
C4481 VDD.t161 GND 0.0205f
C4482 VDD.t152 GND 0.0215f
C4483 VDD.t839 GND 0.0215f
C4484 VDD.t553 GND 0.0248f
C4485 VDD.t606 GND 0.0409f
C4486 VDD.n79 GND 0.0137f
C4487 VDD.n108 GND 0.0126f
C4488 VDD.n109 GND 0.0861f
C4489 VDD.n110 GND 0.734f
C4490 VDD.n114 GND 0.0334f
C4491 VDD.n117 GND 0.0144f
C4492 VDD.n120 GND 0.0144f
C4493 VDD.t265 GND 0.0109f
C4494 VDD.n127 GND 0.0327f
C4495 VDD.t255 GND 0.0428f
C4496 VDD.t281 GND 0.0183f
C4497 VDD.t367 GND 0.0183f
C4498 VDD.t259 GND 0.0183f
C4499 VDD.t379 GND 0.0183f
C4500 VDD.t271 GND 0.0124f
C4501 VDD.n130 GND 0.0218f
C4502 VDD.n132 GND 0.136f
C4503 VDD.n136 GND 0.03f
C4504 VDD.n137 GND 0.0182f
C4505 VDD.n139 GND 0.0129f
C4506 VDD.n143 GND 0.0339f
C4507 VDD.n147 GND 0.0339f
C4508 VDD.n149 GND 0.0339f
C4509 VDD.n150 GND 0.0254f
C4510 VDD.n151 GND 0.0201f
C4511 VDD.n153 GND 0.0339f
C4512 VDD.n157 GND 0.0339f
C4513 VDD.n159 GND 0.0339f
C4514 VDD.n163 GND 0.0339f
C4515 VDD.n165 GND 0.0339f
C4516 VDD.n169 GND 0.0339f
C4517 VDD.n171 GND 0.0339f
C4518 VDD.n175 GND 0.0289f
C4519 VDD.n176 GND 0.0182f
C4520 VDD.n180 GND 0.0129f
C4521 VDD.n181 GND 0.017f
C4522 VDD.n182 GND 0.0144f
C4523 VDD.n183 GND 0.0147f
C4524 VDD.t299 GND 0.015f
C4525 VDD.t369 GND 0.0183f
C4526 VDD.t279 GND 0.0183f
C4527 VDD.t347 GND 0.0183f
C4528 VDD.t371 GND 0.0183f
C4529 VDD.t267 GND 0.0183f
C4530 VDD.t331 GND 0.0183f
C4531 VDD.t361 GND 0.0183f
C4532 VDD.t293 GND 0.0183f
C4533 VDD.t337 GND 0.0176f
C4534 VDD.t257 GND 0.0237f
C4535 VDD.t325 GND 0.0183f
C4536 VDD.t351 GND 0.0183f
C4537 VDD.t377 GND 0.0183f
C4538 VDD.t305 GND 0.0148f
C4539 VDD.t355 GND 0.0183f
C4540 VDD.t269 GND 0.0183f
C4541 VDD.t333 GND 0.0183f
C4542 VDD.t303 GND 0.0183f
C4543 VDD.t373 GND 0.0237f
C4544 VDD.t321 GND 0.0176f
C4545 VDD.t297 GND 0.0183f
C4546 VDD.t365 GND 0.0183f
C4547 VDD.t317 GND 0.0183f
C4548 VDD.t291 GND 0.0183f
C4549 VDD.t359 GND 0.0183f
C4550 VDD.t277 GND 0.0183f
C4551 VDD.t343 GND 0.0183f
C4552 VDD.t309 GND 0.0183f
C4553 VDD.t273 GND 0.0183f
C4554 VDD.t339 GND 0.0126f
C4555 VDD.n184 GND 0.0147f
C4556 VDD.n185 GND 0.0144f
C4557 VDD.n186 GND 0.0136f
C4558 VDD.n188 GND 0.0164f
C4559 VDD.n189 GND 0.0182f
C4560 VDD.n193 GND 0.0234f
C4561 VDD.n197 GND 0.0339f
C4562 VDD.n199 GND 0.0339f
C4563 VDD.n203 GND 0.0339f
C4564 VDD.n205 GND 0.0339f
C4565 VDD.n209 GND 0.0339f
C4566 VDD.n211 GND 0.0339f
C4567 VDD.n215 GND 0.0339f
C4568 VDD.n217 GND 0.0339f
C4569 VDD.n218 GND 0.0201f
C4570 VDD.n221 GND 0.0254f
C4571 VDD.n223 GND 0.0339f
C4572 VDD.n227 GND 0.0339f
C4573 VDD.n229 GND 0.0339f
C4574 VDD.n233 GND 0.0275f
C4575 VDD.n234 GND 0.0182f
C4576 VDD.n236 GND 0.0129f
C4577 VDD.n238 GND 0.0339f
C4578 VDD.n242 GND 0.0339f
C4579 VDD.n244 GND 0.0339f
C4580 VDD.n248 GND 0.0339f
C4581 VDD.n250 GND 0.0339f
C4582 VDD.n254 GND 0.0315f
C4583 VDD.n255 GND 0.0182f
C4584 VDD.n259 GND 0.0129f
C4585 VDD.n260 GND 0.017f
C4586 VDD.n261 GND 0.0144f
C4587 VDD.n262 GND 0.0147f
C4588 VDD.t329 GND 0.0165f
C4589 VDD.t357 GND 0.0183f
C4590 VDD.t287 GND 0.0183f
C4591 VDD.t313 GND 0.0183f
C4592 VDD.t345 GND 0.0183f
C4593 VDD.t289 GND 0.0183f
C4594 VDD.t315 GND 0.0183f
C4595 VDD.t261 GND 0.0183f
C4596 VDD.t283 GND 0.0183f
C4597 VDD.t301 GND 0.0176f
C4598 VDD.t323 GND 0.0237f
C4599 VDD.t349 GND 0.0183f
C4600 VDD.t375 GND 0.0183f
C4601 VDD.n263 GND 0.0147f
C4602 VDD.t353 GND 0.018f
C4603 VDD.t285 GND 0.0183f
C4604 VDD.t307 GND 0.0183f
C4605 VDD.t341 GND 0.0183f
C4606 VDD.t275 GND 0.0183f
C4607 VDD.t311 GND 0.0183f
C4608 VDD.t253 GND 0.0183f
C4609 VDD.t335 GND 0.0183f
C4610 VDD.t363 GND 0.0183f
C4611 VDD.t295 GND 0.0183f
C4612 VDD.t319 GND 0.0183f
C4613 VDD.t263 GND 0.0176f
C4614 VDD.t437 GND 0.0237f
C4615 VDD.t451 GND 0.0176f
C4616 VDD.n264 GND 0.0147f
C4617 VDD.t439 GND 0.0183f
C4618 VDD.t449 GND 0.0183f
C4619 VDD.t445 GND 0.0183f
C4620 VDD.t453 GND 0.0183f
C4621 VDD.t433 GND 0.0183f
C4622 VDD.t447 GND 0.0183f
C4623 VDD.t455 GND 0.0183f
C4624 VDD.t435 GND 0.0183f
C4625 VDD.t441 GND 0.0183f
C4626 VDD.t425 GND 0.0183f
C4627 VDD.t429 GND 0.0183f
C4628 VDD.t443 GND 0.0183f
C4629 VDD.t427 GND 0.0176f
C4630 VDD.t64 GND 0.0236f
C4631 VDD.t66 GND 0.0183f
C4632 VDD.t68 GND 0.0183f
C4633 VDD.t70 GND 0.0173f
C4634 VDD.t1343 GND 0.0193f
C4635 VDD.t398 GND 0.0184f
C4636 VDD.t705 GND 0.0306f
C4637 VDD.t830 GND 0.023f
C4638 VDD.n265 GND 0.0241f
C4639 VDD.n269 GND 0.0507f
C4640 VDD.n271 GND 0.0395f
C4641 VDD.n272 GND 0.0254f
C4642 VDD.n275 GND 0.0201f
C4643 VDD.n277 GND 0.023f
C4644 VDD.n278 GND 0.0182f
C4645 VDD.n280 GND 0.0129f
C4646 VDD.n282 GND 0.0144f
C4647 VDD.n284 GND 0.019f
C4648 VDD.n286 GND 0.0339f
C4649 VDD.n289 GND 0.0339f
C4650 VDD.n291 GND 0.0339f
C4651 VDD.n292 GND 0.0254f
C4652 VDD.n293 GND 0.0201f
C4653 VDD.n295 GND 0.0339f
C4654 VDD.n299 GND 0.0339f
C4655 VDD.n301 GND 0.0339f
C4656 VDD.n305 GND 0.0339f
C4657 VDD.n307 GND 0.0339f
C4658 VDD.n311 GND 0.0339f
C4659 VDD.n313 GND 0.0339f
C4660 VDD.n317 GND 0.0339f
C4661 VDD.n321 GND 0.0339f
C4662 VDD.n323 GND 0.0339f
C4663 VDD.n327 GND 0.0312f
C4664 VDD.n328 GND 0.0182f
C4665 VDD.n330 GND 0.0129f
C4666 VDD.n331 GND 0.017f
C4667 VDD.n335 GND 0.0129f
C4668 VDD.n336 GND 0.0182f
C4669 VDD.n338 GND 0.0278f
C4670 VDD.n339 GND 0.0254f
C4671 VDD.n340 GND 0.0201f
C4672 VDD.n342 GND 0.0339f
C4673 VDD.n346 GND 0.0339f
C4674 VDD.n348 GND 0.0339f
C4675 VDD.n352 GND 0.0339f
C4676 VDD.n354 GND 0.0339f
C4677 VDD.n358 GND 0.0339f
C4678 VDD.n360 GND 0.0339f
C4679 VDD.n364 GND 0.0339f
C4680 VDD.n368 GND 0.0339f
C4681 VDD.n370 GND 0.0312f
C4682 VDD.n371 GND 0.0182f
C4683 VDD.n375 GND 0.0129f
C4684 VDD.n376 GND 0.017f
C4685 VDD.n378 GND 0.0129f
C4686 VDD.n379 GND 0.0182f
C4687 VDD.n383 GND 0.0278f
C4688 VDD.n385 GND 0.0339f
C4689 VDD.n386 GND 0.0254f
C4690 VDD.n387 GND 0.0201f
C4691 VDD.n389 GND 0.0175f
C4692 VDD.n390 GND 11.9f
C4693 VDD.t737 GND 0.0126f
C4694 VDD.t797 GND 0.0121f
C4695 VDD.t1342 GND 0.0106f
C4696 VDD.t552 GND 0.0134f
C4697 VDD.t506 GND 0.0121f
C4698 VDD.t419 GND 0.0169f
C4699 VDD.t629 GND 0.0465f
C4700 VDD.n406 GND 0.0153f
C4701 VDD.n407 GND 0.257f
C4702 VDD.t63 GND 0.0452f
C4703 VDD.t386 GND 0.0156f
C4704 VDD.t546 GND 0.0346f
C4705 VDD.t210 GND 0.0646f
C4706 VDD.t37 GND 0.0274f
C4707 VDD.n408 GND 0.0207f
C4708 VDD.n437 GND 0.0116f
C4709 VDD.n438 GND 0.16f
C4710 VDD.n462 GND 0.0109f
C4711 VDD.t462 GND 0.115f
C4712 VDD.t148 GND 0.0557f
C4713 VDD.t404 GND 0.117f
C4714 VDD.t114 GND 0.0441f
C4715 VDD.n463 GND 0.0473f
C4716 VDD.n464 GND 0.0681f
C4717 VDD.t548 GND 0.0191f
C4718 VDD.t490 GND 0.0128f
C4719 VDD.t1029 GND 0.0119f
C4720 VDD.t795 GND 0.0133f
C4721 VDD.t701 GND 0.0122f
C4722 VDD.t508 GND 0.011f
C4723 VDD.t492 GND 0.0158f
C4724 VDD.t711 GND 0.0129f
C4725 VDD.t801 GND 0.0159f
C4726 VDD.t526 GND 0.0246f
C4727 VDD.t21 GND 0.0353f
C4728 VDD.t620 GND 0.0205f
C4729 VDD.t574 GND 0.0215f
C4730 VDD.t385 GND 0.0215f
C4731 VDD.t865 GND 0.0248f
C4732 VDD.t1430 GND 0.0409f
C4733 VDD.n481 GND 0.0137f
C4734 VDD.n510 GND 0.0126f
C4735 VDD.n511 GND 0.0861f
C4736 VDD.n512 GND 0.467f
C4737 VDD.n513 GND 0.589f
C4738 VDD.n515 GND 0.0171f
C4739 VDD.n518 GND 0.0144f
C4740 VDD.n521 GND 0.0144f
C4741 VDD.t1071 GND 0.0113f
C4742 VDD.n528 GND 0.0334f
C4743 VDD.t1061 GND 0.0419f
C4744 VDD.t1087 GND 0.0183f
C4745 VDD.t1173 GND 0.0183f
C4746 VDD.t1065 GND 0.0183f
C4747 VDD.t1057 GND 0.0183f
C4748 VDD.t1079 GND 0.0128f
C4749 VDD.n531 GND 0.0216f
C4750 VDD.n533 GND 0.135f
C4751 VDD.n537 GND 0.0308f
C4752 VDD.n538 GND 0.0182f
C4753 VDD.n540 GND 0.0129f
C4754 VDD.n544 GND 0.0339f
C4755 VDD.n548 GND 0.0339f
C4756 VDD.n550 GND 0.0339f
C4757 VDD.n551 GND 0.0254f
C4758 VDD.n552 GND 0.0201f
C4759 VDD.n554 GND 0.0339f
C4760 VDD.n558 GND 0.0339f
C4761 VDD.n560 GND 0.0339f
C4762 VDD.n564 GND 0.0339f
C4763 VDD.n566 GND 0.0339f
C4764 VDD.n570 GND 0.0339f
C4765 VDD.n572 GND 0.0339f
C4766 VDD.n576 GND 0.0282f
C4767 VDD.n577 GND 0.0182f
C4768 VDD.n581 GND 0.0129f
C4769 VDD.n582 GND 0.017f
C4770 VDD.n583 GND 0.0144f
C4771 VDD.n584 GND 0.0147f
C4772 VDD.t1105 GND 0.0146f
C4773 VDD.t1047 GND 0.0183f
C4774 VDD.t1083 GND 0.0183f
C4775 VDD.t1153 GND 0.0183f
C4776 VDD.t1049 GND 0.0183f
C4777 VDD.t1073 GND 0.0183f
C4778 VDD.t1137 GND 0.0183f
C4779 VDD.t1167 GND 0.0183f
C4780 VDD.t1099 GND 0.0183f
C4781 VDD.t1143 GND 0.0176f
C4782 VDD.t1063 GND 0.0237f
C4783 VDD.t1131 GND 0.0183f
C4784 VDD.t1157 GND 0.0183f
C4785 VDD.t1055 GND 0.0183f
C4786 VDD.t1111 GND 0.0152f
C4787 VDD.t1161 GND 0.0183f
C4788 VDD.t1075 GND 0.0183f
C4789 VDD.t1139 GND 0.0183f
C4790 VDD.t1109 GND 0.0183f
C4791 VDD.t1051 GND 0.0237f
C4792 VDD.t1127 GND 0.0176f
C4793 VDD.t1103 GND 0.0183f
C4794 VDD.t1171 GND 0.0183f
C4795 VDD.t1123 GND 0.0183f
C4796 VDD.t1097 GND 0.0183f
C4797 VDD.t1165 GND 0.0183f
C4798 VDD.t1085 GND 0.0183f
C4799 VDD.t1149 GND 0.0183f
C4800 VDD.t1115 GND 0.0183f
C4801 VDD.t1077 GND 0.0183f
C4802 VDD.t1145 GND 0.0122f
C4803 VDD.n585 GND 0.0147f
C4804 VDD.n586 GND 0.0144f
C4805 VDD.n587 GND 0.0127f
C4806 VDD.n589 GND 0.0172f
C4807 VDD.n590 GND 0.0182f
C4808 VDD.n594 GND 0.0227f
C4809 VDD.n598 GND 0.0339f
C4810 VDD.n600 GND 0.0339f
C4811 VDD.n604 GND 0.0339f
C4812 VDD.n606 GND 0.0339f
C4813 VDD.n610 GND 0.0339f
C4814 VDD.n612 GND 0.0339f
C4815 VDD.n616 GND 0.0339f
C4816 VDD.n618 GND 0.0339f
C4817 VDD.n619 GND 0.0201f
C4818 VDD.n622 GND 0.0254f
C4819 VDD.n624 GND 0.0339f
C4820 VDD.n628 GND 0.0339f
C4821 VDD.n630 GND 0.0339f
C4822 VDD.n634 GND 0.0282f
C4823 VDD.n635 GND 0.0182f
C4824 VDD.n637 GND 0.0129f
C4825 VDD.n641 GND 0.0339f
C4826 VDD.n643 GND 0.0339f
C4827 VDD.n647 GND 0.0339f
C4828 VDD.n649 GND 0.0339f
C4829 VDD.n653 GND 0.0339f
C4830 VDD.n655 GND 0.0339f
C4831 VDD.n659 GND 0.0308f
C4832 VDD.n660 GND 0.0182f
C4833 VDD.n664 GND 0.0129f
C4834 VDD.n665 GND 0.017f
C4835 VDD.n666 GND 0.0144f
C4836 VDD.n667 GND 0.0147f
C4837 VDD.t1135 GND 0.0161f
C4838 VDD.t1163 GND 0.0183f
C4839 VDD.t1093 GND 0.0183f
C4840 VDD.t1119 GND 0.0183f
C4841 VDD.t1151 GND 0.0183f
C4842 VDD.t1095 GND 0.0183f
C4843 VDD.t1121 GND 0.0183f
C4844 VDD.t1067 GND 0.0183f
C4845 VDD.t1089 GND 0.0183f
C4846 VDD.t1107 GND 0.0176f
C4847 VDD.t1129 GND 0.0237f
C4848 VDD.t1155 GND 0.0183f
C4849 VDD.t1053 GND 0.0183f
C4850 VDD.n668 GND 0.0147f
C4851 VDD.t1159 GND 0.0176f
C4852 VDD.t1091 GND 0.0183f
C4853 VDD.t1113 GND 0.0183f
C4854 VDD.t1147 GND 0.0183f
C4855 VDD.t1081 GND 0.0183f
C4856 VDD.t1117 GND 0.0183f
C4857 VDD.t1059 GND 0.0183f
C4858 VDD.t1141 GND 0.0183f
C4859 VDD.t1169 GND 0.0183f
C4860 VDD.t1101 GND 0.0183f
C4861 VDD.t1125 GND 0.0183f
C4862 VDD.t1069 GND 0.0176f
C4863 VDD.t1462 GND 0.0237f
C4864 VDD.t1476 GND 0.018f
C4865 VDD.n669 GND 0.0147f
C4866 VDD.t1464 GND 0.0183f
C4867 VDD.t1474 GND 0.0183f
C4868 VDD.t1470 GND 0.0183f
C4869 VDD.t1478 GND 0.0183f
C4870 VDD.t1458 GND 0.0183f
C4871 VDD.t1472 GND 0.0183f
C4872 VDD.t1480 GND 0.0183f
C4873 VDD.t1460 GND 0.0183f
C4874 VDD.t1466 GND 0.0183f
C4875 VDD.t1450 GND 0.0183f
C4876 VDD.t1454 GND 0.0183f
C4877 VDD.t1468 GND 0.0183f
C4878 VDD.t1452 GND 0.0176f
C4879 VDD.t566 GND 0.0236f
C4880 VDD.t568 GND 0.0183f
C4881 VDD.t570 GND 0.0183f
C4882 VDD.t564 GND 0.0173f
C4883 VDD.t826 GND 0.0193f
C4884 VDD.t251 GND 0.0184f
C4885 VDD.t218 GND 0.0306f
C4886 VDD.t512 GND 0.0226f
C4887 VDD.n670 GND 0.0241f
C4888 VDD.n674 GND 0.0507f
C4889 VDD.n676 GND 0.0395f
C4890 VDD.n677 GND 0.0254f
C4891 VDD.n680 GND 0.0201f
C4892 VDD.n682 GND 0.0223f
C4893 VDD.n683 GND 0.0182f
C4894 VDD.n685 GND 0.0129f
C4895 VDD.n687 GND 0.0144f
C4896 VDD.n689 GND 0.0197f
C4897 VDD.n691 GND 0.0339f
C4898 VDD.n694 GND 0.0339f
C4899 VDD.n696 GND 0.0339f
C4900 VDD.n697 GND 0.0254f
C4901 VDD.n698 GND 0.0201f
C4902 VDD.n700 GND 0.0339f
C4903 VDD.n704 GND 0.0339f
C4904 VDD.n706 GND 0.0339f
C4905 VDD.n710 GND 0.0339f
C4906 VDD.n712 GND 0.0339f
C4907 VDD.n716 GND 0.0339f
C4908 VDD.n718 GND 0.0339f
C4909 VDD.n722 GND 0.0339f
C4910 VDD.n726 GND 0.0339f
C4911 VDD.n728 GND 0.0339f
C4912 VDD.n732 GND 0.0304f
C4913 VDD.n733 GND 0.0182f
C4914 VDD.n735 GND 0.0129f
C4915 VDD.n736 GND 0.017f
C4916 VDD.n740 GND 0.0129f
C4917 VDD.n741 GND 0.0182f
C4918 VDD.n743 GND 0.0286f
C4919 VDD.n744 GND 0.0254f
C4920 VDD.n745 GND 0.0201f
C4921 VDD.n747 GND 0.0339f
C4922 VDD.n751 GND 0.0339f
C4923 VDD.n753 GND 0.0339f
C4924 VDD.n757 GND 0.0339f
C4925 VDD.n759 GND 0.0339f
C4926 VDD.n763 GND 0.0339f
C4927 VDD.n765 GND 0.0339f
C4928 VDD.n769 GND 0.0339f
C4929 VDD.n773 GND 0.0339f
C4930 VDD.n775 GND 0.0304f
C4931 VDD.n776 GND 0.0182f
C4932 VDD.n780 GND 0.0129f
C4933 VDD.n781 GND 0.017f
C4934 VDD.n783 GND 0.0129f
C4935 VDD.n784 GND 0.0182f
C4936 VDD.n788 GND 0.0286f
C4937 VDD.n790 GND 0.0339f
C4938 VDD.n791 GND 0.0254f
C4939 VDD.n792 GND 0.0199f
C4940 VDD.n793 GND 11.9f
C4941 VDD.n794 GND 3.73f
C4942 VDD.n795 GND 0.519f
C4943 VDD.n796 GND 0.596f
C4944 VDD.n797 GND 2.81f
C4945 VDD.n798 GND 1.01f
C4946 VDD.n799 GND 0.0114f
C4947 VDD.n802 GND 0.0124f
C4948 VDD.n807 GND 0.0138f
C4949 VDD.n808 GND 0.056f
C4950 VDD.n814 GND 0.0124f
C4951 VDD.n815 GND 0.0124f
C4952 VDD.n820 GND 0.0323f
C4953 VDD.n853 GND 0.0239f
C4954 VDD.t559 GND 0.0103f
C4955 VDD.t806 GND 0.0257f
C4956 VDD.t1037 GND 0.0248f
C4957 VDD.t1039 GND 0.0302f
C4958 VDD.t201 GND 0.026f
C4959 VDD.t563 GND 0.0225f
C4960 VDD.t1200 GND 0.0188f
C4961 VDD.t468 GND 0.0298f
C4962 VDD.t383 GND 0.026f
C4963 VDD.t535 GND 0.0225f
C4964 VDD.t1394 GND 0.0225f
C4965 VDD.t1034 GND 0.0215f
C4966 VDD.t1391 GND 0.0231f
C4967 VDD.t421 GND 0.0229f
C4968 VDD.t550 GND 0.0231f
C4969 VDD.t1340 GND 0.0231f
C4970 VDD.t804 GND 0.0291f
C4971 VDD.n857 GND 0.0704f
C4972 VDD.n861 GND 0.0196f
C4973 VDD.n862 GND 0.0687f
C4974 VDD.n863 GND 4.84f
C4975 VDD.n865 GND 0.0171f
C4976 VDD.n868 GND 0.0144f
C4977 VDD.n871 GND 0.0144f
C4978 VDD.t942 GND 0.0113f
C4979 VDD.n878 GND 0.0334f
C4980 VDD.t932 GND 0.0419f
C4981 VDD.t958 GND 0.0183f
C4982 VDD.t916 GND 0.0183f
C4983 VDD.t936 GND 0.0183f
C4984 VDD.t928 GND 0.0183f
C4985 VDD.t948 GND 0.0128f
C4986 VDD.n881 GND 0.0216f
C4987 VDD.n883 GND 0.135f
C4988 VDD.n887 GND 0.0308f
C4989 VDD.n888 GND 0.0182f
C4990 VDD.n890 GND 0.0129f
C4991 VDD.n894 GND 0.0339f
C4992 VDD.n898 GND 0.0339f
C4993 VDD.n900 GND 0.0339f
C4994 VDD.n901 GND 0.0254f
C4995 VDD.n902 GND 0.0201f
C4996 VDD.n904 GND 0.0339f
C4997 VDD.n908 GND 0.0339f
C4998 VDD.n910 GND 0.0339f
C4999 VDD.n914 GND 0.0339f
C5000 VDD.n916 GND 0.0339f
C5001 VDD.n920 GND 0.0339f
C5002 VDD.n922 GND 0.0339f
C5003 VDD.n926 GND 0.0282f
C5004 VDD.n927 GND 0.0182f
C5005 VDD.n931 GND 0.0129f
C5006 VDD.n932 GND 0.017f
C5007 VDD.n933 GND 0.0144f
C5008 VDD.n934 GND 0.0147f
C5009 VDD.t976 GND 0.0146f
C5010 VDD.t918 GND 0.0183f
C5011 VDD.t954 GND 0.0183f
C5012 VDD.t896 GND 0.0183f
C5013 VDD.t920 GND 0.0183f
C5014 VDD.t944 GND 0.0183f
C5015 VDD.t1008 GND 0.0183f
C5016 VDD.t910 GND 0.0183f
C5017 VDD.t970 GND 0.0183f
C5018 VDD.t1014 GND 0.0176f
C5019 VDD.t934 GND 0.0237f
C5020 VDD.t982 GND 0.0183f
C5021 VDD.t900 GND 0.0183f
C5022 VDD.t926 GND 0.0183f
C5023 VDD.t984 GND 0.0152f
C5024 VDD.t904 GND 0.0183f
C5025 VDD.t946 GND 0.0183f
C5026 VDD.t1010 GND 0.0183f
C5027 VDD.t980 GND 0.0183f
C5028 VDD.t922 GND 0.0237f
C5029 VDD.t1000 GND 0.0176f
C5030 VDD.t974 GND 0.0183f
C5031 VDD.t914 GND 0.0183f
C5032 VDD.t996 GND 0.0183f
C5033 VDD.t968 GND 0.0183f
C5034 VDD.t908 GND 0.0183f
C5035 VDD.t956 GND 0.0183f
C5036 VDD.t1020 GND 0.0183f
C5037 VDD.t988 GND 0.0183f
C5038 VDD.t950 GND 0.0183f
C5039 VDD.t1016 GND 0.0122f
C5040 VDD.n935 GND 0.0147f
C5041 VDD.n936 GND 0.0144f
C5042 VDD.n937 GND 0.0127f
C5043 VDD.n939 GND 0.0172f
C5044 VDD.n940 GND 0.0182f
C5045 VDD.n944 GND 0.0227f
C5046 VDD.n948 GND 0.0339f
C5047 VDD.n950 GND 0.0339f
C5048 VDD.n954 GND 0.0339f
C5049 VDD.n956 GND 0.0339f
C5050 VDD.n960 GND 0.0339f
C5051 VDD.n962 GND 0.0339f
C5052 VDD.n966 GND 0.0339f
C5053 VDD.n968 GND 0.0339f
C5054 VDD.n969 GND 0.0201f
C5055 VDD.n972 GND 0.0254f
C5056 VDD.n974 GND 0.0339f
C5057 VDD.n978 GND 0.0339f
C5058 VDD.n980 GND 0.0339f
C5059 VDD.n984 GND 0.0282f
C5060 VDD.n985 GND 0.0182f
C5061 VDD.n987 GND 0.0129f
C5062 VDD.n991 GND 0.0339f
C5063 VDD.n993 GND 0.0339f
C5064 VDD.n997 GND 0.0339f
C5065 VDD.n999 GND 0.0339f
C5066 VDD.n1003 GND 0.0339f
C5067 VDD.n1005 GND 0.0339f
C5068 VDD.n1009 GND 0.0308f
C5069 VDD.n1010 GND 0.0182f
C5070 VDD.n1014 GND 0.0129f
C5071 VDD.n1015 GND 0.017f
C5072 VDD.n1016 GND 0.0144f
C5073 VDD.n1017 GND 0.0147f
C5074 VDD.t1006 GND 0.0161f
C5075 VDD.t906 GND 0.0183f
C5076 VDD.t960 GND 0.0183f
C5077 VDD.t992 GND 0.0183f
C5078 VDD.t1022 GND 0.0183f
C5079 VDD.t966 GND 0.0183f
C5080 VDD.t994 GND 0.0183f
C5081 VDD.t938 GND 0.0183f
C5082 VDD.t962 GND 0.0183f
C5083 VDD.t978 GND 0.0176f
C5084 VDD.t1002 GND 0.0237f
C5085 VDD.t898 GND 0.0183f
C5086 VDD.t924 GND 0.0183f
C5087 VDD.n1018 GND 0.0147f
C5088 VDD.t902 GND 0.0176f
C5089 VDD.t964 GND 0.0183f
C5090 VDD.t986 GND 0.0183f
C5091 VDD.t1018 GND 0.0183f
C5092 VDD.t952 GND 0.0183f
C5093 VDD.t990 GND 0.0183f
C5094 VDD.t930 GND 0.0183f
C5095 VDD.t1012 GND 0.0183f
C5096 VDD.t912 GND 0.0183f
C5097 VDD.t972 GND 0.0183f
C5098 VDD.t998 GND 0.0183f
C5099 VDD.t940 GND 0.0176f
C5100 VDD.t1416 GND 0.0237f
C5101 VDD.t1398 GND 0.018f
C5102 VDD.n1019 GND 0.0147f
C5103 VDD.t1418 GND 0.0183f
C5104 VDD.t1428 GND 0.0183f
C5105 VDD.t1424 GND 0.0183f
C5106 VDD.t1400 GND 0.0183f
C5107 VDD.t1412 GND 0.0183f
C5108 VDD.t1426 GND 0.0183f
C5109 VDD.t1402 GND 0.0183f
C5110 VDD.t1414 GND 0.0183f
C5111 VDD.t1420 GND 0.0183f
C5112 VDD.t1404 GND 0.0183f
C5113 VDD.t1408 GND 0.0183f
C5114 VDD.t1422 GND 0.0183f
C5115 VDD.t1406 GND 0.0176f
C5116 VDD.t51 GND 0.0236f
C5117 VDD.t53 GND 0.0183f
C5118 VDD.t47 GND 0.0183f
C5119 VDD.t49 GND 0.0173f
C5120 VDD.t603 GND 0.0193f
C5121 VDD.t822 GND 0.0184f
C5122 VDD.t1367 GND 0.0306f
C5123 VDD.t396 GND 0.0226f
C5124 VDD.n1020 GND 0.0241f
C5125 VDD.n1024 GND 0.0507f
C5126 VDD.n1026 GND 0.0395f
C5127 VDD.n1027 GND 0.0254f
C5128 VDD.n1030 GND 0.0201f
C5129 VDD.n1032 GND 0.0223f
C5130 VDD.n1033 GND 0.0182f
C5131 VDD.n1035 GND 0.0129f
C5132 VDD.n1037 GND 0.0144f
C5133 VDD.n1039 GND 0.0197f
C5134 VDD.n1041 GND 0.0339f
C5135 VDD.n1044 GND 0.0339f
C5136 VDD.n1046 GND 0.0339f
C5137 VDD.n1047 GND 0.0254f
C5138 VDD.n1048 GND 0.0201f
C5139 VDD.n1050 GND 0.0339f
C5140 VDD.n1054 GND 0.0339f
C5141 VDD.n1056 GND 0.0339f
C5142 VDD.n1060 GND 0.0339f
C5143 VDD.n1062 GND 0.0339f
C5144 VDD.n1066 GND 0.0339f
C5145 VDD.n1068 GND 0.0339f
C5146 VDD.n1072 GND 0.0339f
C5147 VDD.n1076 GND 0.0339f
C5148 VDD.n1078 GND 0.0339f
C5149 VDD.n1082 GND 0.0304f
C5150 VDD.n1083 GND 0.0182f
C5151 VDD.n1085 GND 0.0129f
C5152 VDD.n1086 GND 0.017f
C5153 VDD.n1090 GND 0.0129f
C5154 VDD.n1091 GND 0.0182f
C5155 VDD.n1093 GND 0.0286f
C5156 VDD.n1094 GND 0.0254f
C5157 VDD.n1095 GND 0.0201f
C5158 VDD.n1097 GND 0.0339f
C5159 VDD.n1101 GND 0.0339f
C5160 VDD.n1103 GND 0.0339f
C5161 VDD.n1107 GND 0.0339f
C5162 VDD.n1109 GND 0.0339f
C5163 VDD.n1113 GND 0.0339f
C5164 VDD.n1115 GND 0.0339f
C5165 VDD.n1119 GND 0.0339f
C5166 VDD.n1123 GND 0.0339f
C5167 VDD.n1125 GND 0.0304f
C5168 VDD.n1126 GND 0.0182f
C5169 VDD.n1130 GND 0.0129f
C5170 VDD.n1131 GND 0.017f
C5171 VDD.n1133 GND 0.0129f
C5172 VDD.n1134 GND 0.0182f
C5173 VDD.n1138 GND 0.0286f
C5174 VDD.n1140 GND 0.0339f
C5175 VDD.n1141 GND 0.0254f
C5176 VDD.n1142 GND 0.0199f
C5177 VDD.n1143 GND 13.2f
C5178 VDD.t880 GND 0.0126f
C5179 VDD.t778 GND 0.0124f
C5180 VDD.t141 GND 0.0104f
C5181 VDD.t1177 GND 0.0129f
C5182 VDD.t504 GND 0.0134f
C5183 VDD.t572 GND 0.0107f
C5184 VDD.t781 GND 0.0281f
C5185 VDD.t392 GND 0.0485f
C5186 VDD.t464 GND 0.0199f
C5187 VDD.t242 GND 0.0209f
C5188 VDD.t555 GND 0.0209f
C5189 VDD.t1437 GND 0.0241f
C5190 VDD.t1439 GND 0.0392f
C5191 VDD.n1144 GND 0.0192f
C5192 VDD.n1170 GND 0.0309f
C5193 VDD.n1172 GND 0.013f
C5194 VDD.n1177 GND 0.0119f
C5195 VDD.n1178 GND 0.119f
C5196 VDD.n1179 GND 0.593f
C5197 VDD.n1180 GND 3.2f
C5198 VDD.n1181 GND 4.94f
C5199 VDD.n1182 GND 0.0114f
C5200 VDD.n1185 GND 0.0124f
C5201 VDD.n1190 GND 0.0138f
C5202 VDD.n1191 GND 0.056f
C5203 VDD.n1197 GND 0.0124f
C5204 VDD.n1198 GND 0.0124f
C5205 VDD.n1203 GND 0.0323f
C5206 VDD.n1236 GND 0.0239f
C5207 VDD.t19 GND 0.0103f
C5208 VDD.t775 GND 0.0257f
C5209 VDD.t832 GND 0.0248f
C5210 VDD.t203 GND 0.0302f
C5211 VDD.t465 GND 0.026f
C5212 VDD.t838 GND 0.0225f
C5213 VDD.t716 GND 0.0188f
C5214 VDD.t510 GND 0.0298f
C5215 VDD.t400 GND 0.026f
C5216 VDD.t32 GND 0.0225f
C5217 VDD.t467 GND 0.0225f
C5218 VDD.t1199 GND 0.0215f
C5219 VDD.t878 GND 0.0231f
C5220 VDD.t824 GND 0.0229f
C5221 VDD.t179 GND 0.0231f
C5222 VDD.t741 GND 0.0231f
C5223 VDD.t767 GND 0.0291f
C5224 VDD.n1240 GND 0.0704f
C5225 VDD.n1244 GND 0.0196f
C5226 VDD.n1245 GND 0.599f
C5227 VDD.n1246 GND 0.414f
C5228 VDD.n1249 GND 0.0195f
C5229 VDD.n1251 GND 0.133f
C5230 VDD.n1255 GND 0.0281f
C5231 VDD.n1270 GND 0.03f
C5232 VDD.n1274 GND 0.0493f
C5233 VDD.n1276 GND 0.0493f
C5234 VDD.n1280 GND 0.0493f
C5235 VDD.n1282 GND 0.0493f
C5236 VDD.n1283 GND 0.146f
C5237 VDD.n1285 GND 0.0168f
C5238 VDD.t1315 GND 0.0238f
C5239 VDD.t1239 GND 0.0238f
C5240 VDD.t1291 GND 0.0238f
C5241 VDD.t1217 GND 0.0238f
C5242 VDD.t1243 GND 0.0238f
C5243 VDD.t1275 GND 0.0238f
C5244 VDD.t1211 GND 0.0238f
C5245 VDD.t1301 GND 0.0207f
C5246 VDD.n1291 GND 0.0439f
C5247 VDD.n1295 GND 0.0493f
C5248 VDD.n1297 GND 0.0493f
C5249 VDD.n1301 GND 0.0493f
C5250 VDD.n1303 GND 0.0353f
C5251 VDD.n1304 GND 0.091f
C5252 VDD.n1308 GND 0.0131f
C5253 VDD.n1310 GND 0.0168f
C5254 VDD.n1314 GND 0.0154f
C5255 VDD.t1253 GND 0.0238f
C5256 VDD.t1285 GND 0.0238f
C5257 VDD.t1329 GND 0.0238f
C5258 VDD.t1257 GND 0.0227f
C5259 VDD.t685 GND 0.0238f
C5260 VDD.t675 GND 0.0238f
C5261 VDD.t697 GND 0.0238f
C5262 VDD.t691 GND 0.0125f
C5263 VDD.n1325 GND 0.012f
C5264 VDD.n1327 GND 0.0119f
C5265 VDD.n1331 GND 0.0168f
C5266 VDD.n1333 GND 0.0168f
C5267 VDD.n1337 GND 0.0168f
C5268 VDD.n1339 GND 0.0168f
C5269 VDD.n1346 GND 0.0124f
C5270 VDD.t671 GND 0.0238f
C5271 VDD.t681 GND 0.0238f
C5272 VDD.t689 GND 0.0218f
C5273 VDD.n1349 GND 0.0126f
C5274 VDD.n1351 GND 0.0168f
C5275 VDD.n1354 GND 0.0168f
C5276 VDD.n1356 GND 0.0168f
C5277 VDD.n1363 GND 0.0104f
C5278 VDD.n1365 GND 0.011f
C5279 VDD.n1370 GND 0.0105f
C5280 VDD.t1498 GND 0.0295f
C5281 VDD.n1371 GND 0.03f
C5282 VDD.t661 GND 0.0225f
C5283 VDD.t657 GND 0.0238f
C5284 VDD.t655 GND 0.0238f
C5285 VDD.t659 GND 0.0307f
C5286 VDD.t669 GND 0.013f
C5287 VDD.n1372 GND 0.0178f
C5288 VDD.n1373 GND 0.0105f
C5289 VDD.n1374 GND 0.0101f
C5290 VDD.n1381 GND 0.0119f
C5291 VDD.n1383 GND 0.0168f
C5292 VDD.n1387 GND 0.0168f
C5293 VDD.n1389 GND 0.0168f
C5294 VDD.n1393 GND 0.0132f
C5295 VDD.t695 GND 0.0238f
C5296 VDD.t677 GND 0.0238f
C5297 VDD.t687 GND 0.0238f
C5298 VDD.t667 GND 0.0201f
C5299 VDD.t693 GND 0.0238f
C5300 VDD.t679 GND 0.0238f
C5301 VDD.t683 GND 0.0238f
C5302 VDD.t673 GND 0.0156f
C5303 VDD.n1397 GND 0.0178f
C5304 VDD.n1398 GND 0.0105f
C5305 VDD.n1406 GND 0.012f
C5306 VDD.n1410 GND 0.0155f
C5307 VDD.n1412 GND 0.0168f
C5308 VDD.n1416 GND 0.0168f
C5309 VDD.n1418 GND 0.0168f
C5310 VDD.n1422 GND 0.0138f
C5311 VDD.n1427 GND 0.0105f
C5312 VDD.n1428 GND 0.0249f
C5313 VDD.t1323 GND 0.0229f
C5314 VDD.t1245 GND 0.0238f
C5315 VDD.t1219 GND 0.0238f
C5316 VDD.t1273 GND 0.0238f
C5317 VDD.t1241 GND 0.0238f
C5318 VDD.t1215 GND 0.0238f
C5319 VDD.t1289 GND 0.013f
C5320 VDD.n1429 GND 0.0178f
C5321 VDD.n1430 GND 0.0105f
C5322 VDD.n1433 GND 0.016f
C5323 VDD.n1437 GND 0.0168f
C5324 VDD.n1441 GND 0.0168f
C5325 VDD.n1443 GND 0.0168f
C5326 VDD.n1447 GND 0.0168f
C5327 VDD.n1449 GND 0.0168f
C5328 VDD.n1453 GND 0.0173f
C5329 VDD.n1455 GND 0.0105f
C5330 VDD.t1325 GND 0.0238f
C5331 VDD.t1229 GND 0.0238f
C5332 VDD.t1307 GND 0.0238f
C5333 VDD.t1277 GND 0.0184f
C5334 VDD.n1456 GND 0.0178f
C5335 VDD.t1225 GND 0.0244f
C5336 VDD.t1299 GND 0.0229f
C5337 VDD.t1247 GND 0.0238f
C5338 VDD.t1221 GND 0.0365f
C5339 VDD.t1295 GND 0.0522f
C5340 VDD.t1263 GND 0.0528f
C5341 VDD.t1203 GND 0.0528f
C5342 VDD.t1237 GND 0.0528f
C5343 VDD.t1205 GND 0.0528f
C5344 VDD.t1269 GND 0.0528f
C5345 VDD.t1233 GND 0.0528f
C5346 VDD.t1311 GND 0.0528f
C5347 VDD.t1283 GND 0.0528f
C5348 VDD.t1251 GND 0.0528f
C5349 VDD.t1321 GND 0.053f
C5350 VDD.t1279 GND 0.0239f
C5351 VDD.t1207 GND 0.0309f
C5352 VDD.n1457 GND 0.017f
C5353 VDD.n1458 GND 0.0105f
C5354 VDD.n1463 GND 0.0105f
C5355 VDD.n1467 GND 0.0168f
C5356 VDD.n1469 GND 0.0168f
C5357 VDD.n1473 GND 0.0168f
C5358 VDD.n1475 GND 0.0168f
C5359 VDD.n1479 GND 0.0168f
C5360 VDD.n1481 GND 0.0168f
C5361 VDD.n1485 GND 0.0168f
C5362 VDD.n1489 GND 0.0168f
C5363 VDD.n1491 GND 0.0168f
C5364 VDD.n1495 GND 0.0168f
C5365 VDD.n1497 GND 0.0168f
C5366 VDD.n1501 GND 0.0168f
C5367 VDD.n1503 GND 0.0153f
C5368 VDD.n1504 GND 0.012f
C5369 VDD.t1319 GND 0.0547f
C5370 VDD.t1209 GND 0.0238f
C5371 VDD.t1281 GND 0.0238f
C5372 VDD.t1309 GND 0.0238f
C5373 VDD.t1231 GND 0.0238f
C5374 VDD.t1267 GND 0.0238f
C5375 VDD.t1313 GND 0.0238f
C5376 VDD.t1235 GND 0.0238f
C5377 VDD.t1271 GND 0.0238f
C5378 VDD.t1259 GND 0.0238f
C5379 VDD.t1293 GND 0.0238f
C5380 VDD.t1317 GND 0.0238f
C5381 VDD.t1265 GND 0.0238f
C5382 VDD.t1297 GND 0.0238f
C5383 VDD.t1223 GND 0.0238f
C5384 VDD.t1249 GND 0.0229f
C5385 VDD.t1287 GND 0.0238f
C5386 VDD.t1255 GND 0.0238f
C5387 VDD.t1327 GND 0.0238f
C5388 VDD.t1303 GND 0.0238f
C5389 VDD.t1213 GND 0.0238f
C5390 VDD.t1261 GND 0.0238f
C5391 VDD.t1227 GND 0.0238f
C5392 VDD.t1305 GND 0.0286f
C5393 VDD.n1507 GND 0.0249f
C5394 VDD.n1508 GND 0.0105f
C5395 VDD.n1513 GND 0.0134f
C5396 VDD.n1517 GND 0.0168f
C5397 VDD.n1519 GND 0.0168f
C5398 VDD.n1523 GND 0.0168f
C5399 VDD.n1526 GND 0.119f
C5400 VDD.n1527 GND 0.034f
C5401 VDD.n1529 GND 0.0364f
C5402 VDD.n1533 GND 0.0364f
C5403 VDD.n1537 GND 0.0364f
C5404 VDD.n1539 GND 0.0265f
C5405 VDD.n1540 GND 0.407f
C5406 VDD.t834 GND 0.0326f
C5407 VDD.n1541 GND 0.047f
C5408 VDD.n1548 GND 0.116f
C5409 VDD.t1396 GND 0.0126f
C5410 VDD.t757 GND 0.0121f
C5411 VDD.t25 GND 0.0106f
C5412 VDD.t414 GND 0.0134f
C5413 VDD.t212 GND 0.0121f
C5414 VDD.t1192 GND 0.0169f
C5415 VDD.t557 GND 0.0465f
C5416 VDD.n1564 GND 0.0153f
C5417 VDD.n1565 GND 0.257f
C5418 VDD.t556 GND 0.0452f
C5419 VDD.t100 GND 0.0156f
C5420 VDD.t230 GND 0.0346f
C5421 VDD.t876 GND 0.0646f
C5422 VDD.t764 GND 0.0274f
C5423 VDD.n1566 GND 0.0207f
C5424 VDD.n1595 GND 0.0116f
C5425 VDD.n1596 GND 0.16f
C5426 VDD.n1597 GND 0.6f
C5427 VDD.n1598 GND 0.58f
C5428 VDD.n1599 GND 0.445f
C5429 VDD.n1600 GND 3.26f
C5430 VDD.n1601 GND 2.59f
C5431 VDD.n1602 GND 4.7f
C5432 VDD.n1603 GND 13.5f
C5433 VDD.n1613 GND 0.0244f
C5434 VDD.n1622 GND 0.0743f
C5435 VDD.n1623 GND 0.0594f
C5436 VDD.n1642 GND 0.0459f
C5437 VDD.n1646 GND 0.0396f
C5438 VDD.n1652 GND 0.035f
C5439 VDD.n1653 GND 0.156f
C5440 VDD.n1654 GND 0.13f
C5441 VDD.n1655 GND 0.0932f
C5442 VDD.n1656 GND 0.12f
C5443 VDD.n1657 GND 0.148f
C5444 VDD.n1658 GND 0.146f
C5445 VDD.n1659 GND 0.133f
C5446 VDD.n1660 GND 0.152f
C5447 VDD.n1661 GND 0.114f
C5448 VDD.n1662 GND 0.299f
C5449 VDD.n1663 GND 11.5f
C5450 VDD.n1664 GND 0.274f
C5451 VDD.n1665 GND 0.0237f
C5452 VDD.n1666 GND 0.0462f
C5453 VDD.t642 GND 0.0597f
C5454 VDD.n1678 GND 0.035f
C5455 VDD.n1686 GND 0.0437f
C5456 VDD.n1687 GND 0.0152f
C5457 VDD.n1688 GND 0.0128f
C5458 VDD.n1695 GND 0.0504f
C5459 VDD.n1711 GND 0.0735f
C5460 VDD.t1359 GND 0.0597f
C5461 VDD.n1712 GND 0.035f
C5462 VDD.n1721 GND 0.0491f
C5463 VDD.n1723 GND 0.0135f
C5464 VDD.n1737 GND 0.0484f
C5465 VDD.n1738 GND 0.0582f
C5466 VDD.n1744 GND 0.0583f
C5467 VDD.n1748 GND 0.0134f
C5468 VDD.n1749 GND 0.047f
C5469 VDD.n1753 GND 0.0289f
C5470 VDD.n1754 GND 0.0135f
C5471 VDD.t388 GND 0.169f
C5472 VDD.n1764 GND 0.0735f
C5473 VDD.n1770 GND 0.0135f
C5474 VDD.n1771 GND 0.0287f
C5475 VDD.n1773 GND 0.0248f
C5476 VDD.n1774 GND 0.13f
C5477 VDD.n1775 GND 0.427f
C5478 VDD.n1801 GND 0.0443f
C5479 VDD.t1361 GND 0.0187f
C5480 VDD.n1802 GND 0.0194f
C5481 VDD.n1803 GND 0.0239f
C5482 VDD.t639 GND 0.0185f
C5483 VDD.n1804 GND 0.16f
C5484 VDD.n1805 GND 0.966f
C5485 VDD.n1806 GND 0.102f
C5486 VDD.n1807 GND 1.15f
C5487 VDD.n1808 GND 0.921f
C5488 VDD.t1357 GND 0.0383f
C5489 VDD.t608 GND 0.0134f
C5490 VDD.n1809 GND 0.0699f
C5491 VDD.n1816 GND 0.0579f
C5492 VDD.n1817 GND 0.0223f
C5493 VDD.n1821 GND 0.0682f
C5494 VDD.n1823 GND 0.0779f
C5495 VDD.n1825 GND 0.0106f
C5496 VDD.t208 GND 0.0288f
C5497 VDD.t26 GND 0.0109f
C5498 VDD.n1836 GND 0.0397f
C5499 VDD.n1839 GND 0.0201f
C5500 VDD.n1840 GND 0.0133f
C5501 VDD.n1841 GND 0.114f
C5502 VDD.n1842 GND 0.0382f
C5503 VDD.n1847 GND 0.0681f
C5504 VDD.n1849 GND 0.0898f
C5505 VDD.n1857 GND 0.0865f
C5506 VDD.n1858 GND 0.0386f
C5507 VDD.n1863 GND 0.0419f
C5508 VDD.t106 GND 0.0681f
C5509 VDD.n1872 GND 0.294f
C5510 VDD.n1873 GND 0.165f
C5511 VDD.n1874 GND 0.0664f
C5512 VDD.n1875 GND 0.0215f
C5513 VDD.t528 GND 0.0855f
C5514 VDD.n1886 GND 0.0455f
C5515 VDD.n1887 GND 0.112f
C5516 VDD.n1889 GND 0.0121f
C5517 VDD.n1892 GND 0.0857f
C5518 VDD.n1893 GND 0.0898f
C5519 VDD.n1901 GND 0.0427f
C5520 VDD.n1905 GND 0.0386f
C5521 VDD.t28 GND 0.0681f
C5522 VDD.n1914 GND 0.0681f
C5523 VDD.n1916 GND 0.0875f
C5524 VDD.n1917 GND 0.28f
C5525 VDD.n1918 GND 0.166f
C5526 VDD.n1919 GND 0.196f
C5527 VDD.n1920 GND 0.0783f
C5528 VDD.n1921 GND 6.11f
C5529 VDD.n1922 GND 0.159f
C5530 VDD.n1923 GND 0.138f
C5531 VDD.t864 GND 0.0214f
C5532 VDD.t1044 GND 0.0214f
C5533 VDD.n1924 GND 0.326f
C5534 VDD.n1925 GND 0.0174f
C5535 VDD.n1926 GND 0.0127f
C5536 VDD.n1927 GND 0.4f
C5537 VDD.n1930 GND 0.0303f
C5538 VDD.n1931 GND 0.317f
C5539 VDD.n1933 GND 0.127f
C5540 VDD.n1935 GND 0.0135f
C5541 VDD.n1939 GND 0.2f
C5542 VDD.n1940 GND 0.0135f
C5543 VDD.n1942 GND 0.0303f
C5544 VDD.n1943 GND 0.0181f
C5545 VDD.t1042 GND 0.0214f
C5546 VDD.n1945 GND 0.163f
C5547 VDD.n1946 GND 0.0851f
C5548 VDD.n1948 GND 0.0135f
C5549 VDD.n1949 GND 0.317f
C5550 VDD.n1950 GND 0.0169f
C5551 VDD.n1951 GND 0.0169f
C5552 VDD.t1041 GND 0.399f
C5553 VDD.n1952 GND 0.014f
C5554 VDD.n1953 GND 0.2f
C5555 VDD.n1954 GND 0.0127f
C5556 VDD.n1955 GND 0.0127f
C5557 VDD.n1957 GND 0.0884f
C5558 VDD.n1960 GND 0.0169f
C5559 VDD.n1961 GND 0.0169f
C5560 VDD.t863 GND 0.387f
C5561 VDD.n1967 GND 0.0169f
C5562 VDD.n1968 GND 0.0169f
C5563 VDD.t1043 GND 0.4f
C5564 VDD.n1970 GND 0.0169f
C5565 VDD.n1971 GND 0.0169f
C5566 VDD.n1974 GND 0.0135f
C5567 VDD.n1976 GND 0.0127f
C5568 VDD.n1979 GND 0.202f
C5569 VDD.n1980 GND 0.127f
C5570 VDD.n1981 GND 0.0329f
C5571 VDD.n1982 GND 9.56f
C5572 VDD.n1983 GND 0.274f
C5573 VDD.n2009 GND 0.0443f
C5574 VDD.t1490 GND 0.0187f
C5575 VDD.n2010 GND 0.0194f
C5576 VDD.n2011 GND 0.0239f
C5577 VDD.t245 GND 0.0185f
C5578 VDD.n2012 GND 0.611f
C5579 VDD.n2013 GND 0.461f
C5580 VDD.n2014 GND 0.0237f
C5581 VDD.n2015 GND 0.0462f
C5582 VDD.t243 GND 0.0597f
C5583 VDD.n2027 GND 0.035f
C5584 VDD.n2035 GND 0.0437f
C5585 VDD.n2036 GND 0.0152f
C5586 VDD.n2037 GND 0.0128f
C5587 VDD.n2044 GND 0.0504f
C5588 VDD.n2060 GND 0.0735f
C5589 VDD.t1493 GND 0.0597f
C5590 VDD.n2061 GND 0.035f
C5591 VDD.n2070 GND 0.0491f
C5592 VDD.n2072 GND 0.0135f
C5593 VDD.n2086 GND 0.0484f
C5594 VDD.n2087 GND 0.0582f
C5595 VDD.n2093 GND 0.0583f
C5596 VDD.n2097 GND 0.0134f
C5597 VDD.n2098 GND 0.047f
C5598 VDD.n2102 GND 0.0289f
C5599 VDD.n2103 GND 0.0135f
C5600 VDD.t228 GND 0.169f
C5601 VDD.n2113 GND 0.0735f
C5602 VDD.n2119 GND 0.0135f
C5603 VDD.n2120 GND 0.0287f
C5604 VDD.n2122 GND 0.0248f
C5605 VDD.n2123 GND 0.13f
C5606 VDD.n2124 GND 0.427f
C5607 VDD.n2125 GND 0.0484f
C5608 VDD.n2126 GND 0.102f
C5609 VDD.n2127 GND 0.583f
C5610 VDD.n2128 GND 1.1f
C5611 VDD.n2129 GND 0.436f
C5612 VDD.t815 GND 0.0383f
C5613 VDD.t1175 GND 0.0134f
C5614 VDD.n2130 GND 0.0699f
C5615 VDD.n2137 GND 0.0579f
C5616 VDD.n2138 GND 0.0223f
C5617 VDD.n2142 GND 0.0682f
C5618 VDD.n2144 GND 0.0779f
C5619 VDD.n2146 GND 0.0106f
C5620 VDD.t836 GND 0.0288f
C5621 VDD.t1182 GND 0.0109f
C5622 VDD.n2157 GND 0.0397f
C5623 VDD.n2160 GND 0.0201f
C5624 VDD.n2161 GND 0.0133f
C5625 VDD.n2162 GND 0.114f
C5626 VDD.n2163 GND 0.0382f
C5627 VDD.n2168 GND 0.0681f
C5628 VDD.n2170 GND 0.0898f
C5629 VDD.n2178 GND 0.0865f
C5630 VDD.n2179 GND 0.0386f
C5631 VDD.n2184 GND 0.0419f
C5632 VDD.t719 GND 0.0681f
C5633 VDD.n2193 GND 0.295f
C5634 VDD.n2194 GND 0.165f
C5635 VDD.n2195 GND 0.0664f
C5636 VDD.n2196 GND 0.0215f
C5637 VDD.t481 GND 0.0855f
C5638 VDD.n2207 GND 0.0455f
C5639 VDD.n2208 GND 0.112f
C5640 VDD.n2210 GND 0.0121f
C5641 VDD.n2213 GND 0.0857f
C5642 VDD.n2214 GND 0.0898f
C5643 VDD.n2222 GND 0.0427f
C5644 VDD.n2226 GND 0.0386f
C5645 VDD.t103 GND 0.0681f
C5646 VDD.n2235 GND 0.0681f
C5647 VDD.n2237 GND 0.0875f
C5648 VDD.n2238 GND 0.28f
C5649 VDD.n2239 GND 0.166f
C5650 VDD.n2240 GND 0.196f
C5651 VDD.n2241 GND 0.0783f
C5652 VDD.n2242 GND 6.11f
C5653 VDD.n2243 GND 0.274f
C5654 VDD.n2244 GND 0.0237f
C5655 VDD.n2245 GND 0.0462f
C5656 VDD.t624 GND 0.0597f
C5657 VDD.n2257 GND 0.035f
C5658 VDD.n2265 GND 0.0437f
C5659 VDD.n2266 GND 0.0152f
C5660 VDD.n2267 GND 0.0128f
C5661 VDD.n2274 GND 0.0504f
C5662 VDD.n2290 GND 0.0735f
C5663 VDD.t222 GND 0.0597f
C5664 VDD.n2291 GND 0.035f
C5665 VDD.n2300 GND 0.0491f
C5666 VDD.n2302 GND 0.0135f
C5667 VDD.n2316 GND 0.0484f
C5668 VDD.n2317 GND 0.0582f
C5669 VDD.n2323 GND 0.0583f
C5670 VDD.n2327 GND 0.0134f
C5671 VDD.n2328 GND 0.047f
C5672 VDD.n2332 GND 0.0289f
C5673 VDD.n2333 GND 0.0135f
C5674 VDD.t181 GND 0.169f
C5675 VDD.n2343 GND 0.0735f
C5676 VDD.n2349 GND 0.0135f
C5677 VDD.n2350 GND 0.0287f
C5678 VDD.n2352 GND 0.0248f
C5679 VDD.n2353 GND 0.13f
C5680 VDD.n2354 GND 0.427f
C5681 VDD.n2380 GND 0.0443f
C5682 VDD.t220 GND 0.0187f
C5683 VDD.n2381 GND 0.0194f
C5684 VDD.n2382 GND 0.0239f
C5685 VDD.t621 GND 0.0185f
C5686 VDD.n2383 GND 0.16f
C5687 VDD.n2384 GND 0.966f
C5688 VDD.n2385 GND 0.102f
C5689 VDD.n2386 GND 1.15f
C5690 VDD.n2387 GND 0.921f
C5691 VDD.t1379 GND 0.0383f
C5692 VDD.t818 GND 0.0134f
C5693 VDD.n2388 GND 0.0699f
C5694 VDD.n2395 GND 0.0579f
C5695 VDD.n2396 GND 0.0223f
C5696 VDD.n2400 GND 0.0682f
C5697 VDD.n2402 GND 0.0779f
C5698 VDD.n2404 GND 0.0106f
C5699 VDD.t1500 GND 0.0288f
C5700 VDD.t722 GND 0.0109f
C5701 VDD.n2415 GND 0.0397f
C5702 VDD.n2418 GND 0.0201f
C5703 VDD.n2419 GND 0.0133f
C5704 VDD.n2420 GND 0.114f
C5705 VDD.n2421 GND 0.0382f
C5706 VDD.n2426 GND 0.0681f
C5707 VDD.n2428 GND 0.0898f
C5708 VDD.n2436 GND 0.0865f
C5709 VDD.n2437 GND 0.0386f
C5710 VDD.n2442 GND 0.0419f
C5711 VDD.t485 GND 0.0681f
C5712 VDD.n2451 GND 0.295f
C5713 VDD.n2452 GND 0.165f
C5714 VDD.n2453 GND 0.0664f
C5715 VDD.n2454 GND 0.0215f
C5716 VDD.t118 GND 0.0855f
C5717 VDD.n2465 GND 0.0455f
C5718 VDD.n2466 GND 0.112f
C5719 VDD.n2468 GND 0.0121f
C5720 VDD.n2471 GND 0.0857f
C5721 VDD.n2472 GND 0.0898f
C5722 VDD.n2480 GND 0.0427f
C5723 VDD.n2484 GND 0.0386f
C5724 VDD.t471 GND 0.0681f
C5725 VDD.n2493 GND 0.0681f
C5726 VDD.n2495 GND 0.0875f
C5727 VDD.n2496 GND 0.28f
C5728 VDD.n2497 GND 0.166f
C5729 VDD.n2498 GND 0.196f
C5730 VDD.n2499 GND 0.0783f
C5731 VDD.n2500 GND 6.11f
C5732 VDD.n2501 GND 0.274f
C5733 VDD.n2502 GND 0.0237f
C5734 VDD.n2503 GND 0.0462f
C5735 VDD.t842 GND 0.0597f
C5736 VDD.n2515 GND 0.035f
C5737 VDD.n2523 GND 0.0437f
C5738 VDD.n2524 GND 0.0152f
C5739 VDD.n2525 GND 0.0128f
C5740 VDD.n2532 GND 0.0504f
C5741 VDD.n2548 GND 0.0735f
C5742 VDD.t55 GND 0.0597f
C5743 VDD.n2549 GND 0.035f
C5744 VDD.n2558 GND 0.0491f
C5745 VDD.n2560 GND 0.0135f
C5746 VDD.n2574 GND 0.0484f
C5747 VDD.n2575 GND 0.0582f
C5748 VDD.n2581 GND 0.0583f
C5749 VDD.n2585 GND 0.0134f
C5750 VDD.n2586 GND 0.047f
C5751 VDD.n2590 GND 0.0289f
C5752 VDD.n2591 GND 0.0135f
C5753 VDD.t713 GND 0.169f
C5754 VDD.n2601 GND 0.0735f
C5755 VDD.n2607 GND 0.0135f
C5756 VDD.n2608 GND 0.0287f
C5757 VDD.n2610 GND 0.0248f
C5758 VDD.n2611 GND 0.13f
C5759 VDD.n2612 GND 0.427f
C5760 VDD.n2638 GND 0.0443f
C5761 VDD.t57 GND 0.0187f
C5762 VDD.n2639 GND 0.0194f
C5763 VDD.n2640 GND 0.0239f
C5764 VDD.t844 GND 0.0185f
C5765 VDD.n2641 GND 0.16f
C5766 VDD.n2642 GND 0.966f
C5767 VDD.n2643 GND 0.102f
C5768 VDD.n2644 GND 1.15f
C5769 VDD.n2645 GND 0.921f
C5770 VDD.t872 GND 0.0383f
C5771 VDD.t1189 GND 0.0134f
C5772 VDD.n2646 GND 0.0699f
C5773 VDD.n2653 GND 0.0579f
C5774 VDD.n2654 GND 0.0223f
C5775 VDD.n2658 GND 0.0682f
C5776 VDD.n2660 GND 0.0779f
C5777 VDD.n2662 GND 0.0106f
C5778 VDD.t665 GND 0.0288f
C5779 VDD.t601 GND 0.0109f
C5780 VDD.n2673 GND 0.0397f
C5781 VDD.n2676 GND 0.0201f
C5782 VDD.n2677 GND 0.0133f
C5783 VDD.n2678 GND 0.114f
C5784 VDD.n2679 GND 0.0382f
C5785 VDD.n2684 GND 0.0681f
C5786 VDD.n2686 GND 0.0898f
C5787 VDD.n2694 GND 0.0865f
C5788 VDD.n2695 GND 0.0386f
C5789 VDD.n2700 GND 0.0419f
C5790 VDD.t531 GND 0.0681f
C5791 VDD.n2709 GND 0.295f
C5792 VDD.n2710 GND 0.165f
C5793 VDD.n2711 GND 0.0664f
C5794 VDD.n2712 GND 0.0215f
C5795 VDD.t652 GND 0.0855f
C5796 VDD.n2723 GND 0.0455f
C5797 VDD.n2724 GND 0.112f
C5798 VDD.n2726 GND 0.0121f
C5799 VDD.n2729 GND 0.0857f
C5800 VDD.n2730 GND 0.0898f
C5801 VDD.n2738 GND 0.0427f
C5802 VDD.n2742 GND 0.0386f
C5803 VDD.t184 GND 0.0681f
C5804 VDD.n2751 GND 0.0681f
C5805 VDD.n2753 GND 0.0875f
C5806 VDD.n2754 GND 0.28f
C5807 VDD.n2755 GND 0.166f
C5808 VDD.n2756 GND 0.196f
C5809 VDD.n2757 GND 0.0783f
C5810 VDD.n2758 GND 6.11f
C5811 VDD.n2759 GND 0.274f
C5812 VDD.n2760 GND 0.0237f
C5813 VDD.n2761 GND 0.0462f
C5814 VDD.t134 GND 0.0597f
C5815 VDD.n2773 GND 0.035f
C5816 VDD.n2781 GND 0.0437f
C5817 VDD.n2782 GND 0.0152f
C5818 VDD.n2783 GND 0.0128f
C5819 VDD.n2790 GND 0.0504f
C5820 VDD.n2806 GND 0.0735f
C5821 VDD.t595 GND 0.0597f
C5822 VDD.n2807 GND 0.035f
C5823 VDD.n2816 GND 0.0491f
C5824 VDD.n2818 GND 0.0135f
C5825 VDD.n2832 GND 0.0484f
C5826 VDD.n2833 GND 0.0582f
C5827 VDD.n2839 GND 0.0583f
C5828 VDD.n2843 GND 0.0134f
C5829 VDD.n2844 GND 0.047f
C5830 VDD.n2848 GND 0.0289f
C5831 VDD.n2849 GND 0.0135f
C5832 VDD.t542 GND 0.169f
C5833 VDD.n2859 GND 0.0735f
C5834 VDD.n2865 GND 0.0135f
C5835 VDD.n2866 GND 0.0287f
C5836 VDD.n2868 GND 0.0248f
C5837 VDD.n2869 GND 0.13f
C5838 VDD.n2870 GND 0.427f
C5839 VDD.n2896 GND 0.0443f
C5840 VDD.t593 GND 0.0187f
C5841 VDD.n2897 GND 0.0194f
C5842 VDD.n2898 GND 0.0239f
C5843 VDD.t131 GND 0.0185f
C5844 VDD.n2899 GND 0.16f
C5845 VDD.n2900 GND 0.966f
C5846 VDD.n2901 GND 0.102f
C5847 VDD.n2902 GND 1.15f
C5848 VDD.n2903 GND 0.921f
C5849 VDD.t394 GND 0.0383f
C5850 VDD.t406 GND 0.0134f
C5851 VDD.n2904 GND 0.0699f
C5852 VDD.n2911 GND 0.0579f
C5853 VDD.n2912 GND 0.0223f
C5854 VDD.n2916 GND 0.0682f
C5855 VDD.n2918 GND 0.0779f
C5856 VDD.n2920 GND 0.0106f
C5857 VDD.t561 GND 0.0288f
C5858 VDD.t1024 GND 0.0109f
C5859 VDD.n2931 GND 0.0397f
C5860 VDD.n2934 GND 0.0201f
C5861 VDD.n2935 GND 0.0133f
C5862 VDD.n2936 GND 0.114f
C5863 VDD.n2937 GND 0.0382f
C5864 VDD.n2942 GND 0.0681f
C5865 VDD.n2944 GND 0.0898f
C5866 VDD.n2952 GND 0.0865f
C5867 VDD.n2953 GND 0.0386f
C5868 VDD.n2958 GND 0.0419f
C5869 VDD.t15 GND 0.0681f
C5870 VDD.n2967 GND 0.295f
C5871 VDD.n2968 GND 0.165f
C5872 VDD.n2969 GND 0.0664f
C5873 VDD.n2970 GND 0.0215f
C5874 VDD.t12 GND 0.0855f
C5875 VDD.n2981 GND 0.0455f
C5876 VDD.n2982 GND 0.112f
C5877 VDD.n2984 GND 0.0121f
C5878 VDD.n2987 GND 0.0857f
C5879 VDD.n2988 GND 0.0898f
C5880 VDD.n2996 GND 0.0427f
C5881 VDD.n3000 GND 0.0386f
C5882 VDD.t488 GND 0.0681f
C5883 VDD.n3009 GND 0.0681f
C5884 VDD.n3011 GND 0.0875f
C5885 VDD.n3012 GND 0.28f
C5886 VDD.n3013 GND 0.166f
C5887 VDD.n3014 GND 0.196f
C5888 VDD.n3015 GND 0.0783f
C5889 VDD.n3016 GND 6.11f
C5890 VDD.n3017 GND 0.274f
C5891 VDD.n3018 GND 0.0237f
C5892 VDD.n3019 GND 0.0462f
C5893 VDD.t473 GND 0.0597f
C5894 VDD.n3031 GND 0.035f
C5895 VDD.n3039 GND 0.0437f
C5896 VDD.n3040 GND 0.0152f
C5897 VDD.n3041 GND 0.0128f
C5898 VDD.n3048 GND 0.0504f
C5899 VDD.n3064 GND 0.0735f
C5900 VDD.t41 GND 0.0597f
C5901 VDD.n3065 GND 0.035f
C5902 VDD.n3074 GND 0.0491f
C5903 VDD.n3076 GND 0.0135f
C5904 VDD.n3090 GND 0.0484f
C5905 VDD.n3091 GND 0.0582f
C5906 VDD.n3097 GND 0.0583f
C5907 VDD.n3101 GND 0.0134f
C5908 VDD.n3102 GND 0.047f
C5909 VDD.n3106 GND 0.0289f
C5910 VDD.n3107 GND 0.0135f
C5911 VDD.t647 GND 0.169f
C5912 VDD.n3117 GND 0.0735f
C5913 VDD.n3123 GND 0.0135f
C5914 VDD.n3124 GND 0.0287f
C5915 VDD.n3126 GND 0.0248f
C5916 VDD.n3127 GND 0.13f
C5917 VDD.n3128 GND 0.427f
C5918 VDD.n3154 GND 0.0443f
C5919 VDD.t39 GND 0.0187f
C5920 VDD.n3155 GND 0.0194f
C5921 VDD.n3156 GND 0.0239f
C5922 VDD.t475 GND 0.0185f
C5923 VDD.n3157 GND 0.16f
C5924 VDD.n3158 GND 0.966f
C5925 VDD.n3159 GND 0.102f
C5926 VDD.n3160 GND 1.15f
C5927 VDD.n3161 GND 0.921f
C5928 VDD.t544 GND 0.0383f
C5929 VDD.t827 GND 0.0134f
C5930 VDD.n3162 GND 0.0699f
C5931 VDD.n3169 GND 0.0579f
C5932 VDD.n3170 GND 0.0223f
C5933 VDD.n3174 GND 0.0682f
C5934 VDD.n3176 GND 0.0779f
C5935 VDD.n3178 GND 0.0106f
C5936 VDD.t840 GND 0.0288f
C5937 VDD.t1482 GND 0.0109f
C5938 VDD.n3189 GND 0.0397f
C5939 VDD.n3192 GND 0.0201f
C5940 VDD.n3193 GND 0.0133f
C5941 VDD.n3194 GND 0.114f
C5942 VDD.n3195 GND 0.0382f
C5943 VDD.n3200 GND 0.0681f
C5944 VDD.n3202 GND 0.0898f
C5945 VDD.n3210 GND 0.0865f
C5946 VDD.n3211 GND 0.0386f
C5947 VDD.n3216 GND 0.0419f
C5948 VDD.t412 GND 0.0681f
C5949 VDD.n3225 GND 0.295f
C5950 VDD.n3226 GND 0.165f
C5951 VDD.n3227 GND 0.0664f
C5952 VDD.n3228 GND 0.0215f
C5953 VDD.t718 GND 0.0855f
C5954 VDD.n3239 GND 0.0455f
C5955 VDD.n3240 GND 0.112f
C5956 VDD.n3242 GND 0.0121f
C5957 VDD.n3245 GND 0.0857f
C5958 VDD.n3246 GND 0.0898f
C5959 VDD.n3254 GND 0.0427f
C5960 VDD.n3258 GND 0.0386f
C5961 VDD.t234 GND 0.0681f
C5962 VDD.n3267 GND 0.0681f
C5963 VDD.n3269 GND 0.0875f
C5964 VDD.n3270 GND 0.28f
C5965 VDD.n3271 GND 0.166f
C5966 VDD.n3272 GND 0.196f
C5967 VDD.n3273 GND 0.0783f
C5968 VDD.n3274 GND 6.11f
C5969 VDD.n3275 GND 0.274f
C5970 VDD.n3276 GND 0.0237f
C5971 VDD.n3277 GND 0.0462f
C5972 VDD.t1331 GND 0.0597f
C5973 VDD.n3289 GND 0.035f
C5974 VDD.n3297 GND 0.0437f
C5975 VDD.n3298 GND 0.0152f
C5976 VDD.n3299 GND 0.0128f
C5977 VDD.n3306 GND 0.0504f
C5978 VDD.n3322 GND 0.0735f
C5979 VDD.t731 GND 0.0597f
C5980 VDD.n3323 GND 0.035f
C5981 VDD.n3332 GND 0.0491f
C5982 VDD.n3334 GND 0.0135f
C5983 VDD.n3348 GND 0.0484f
C5984 VDD.n3349 GND 0.0582f
C5985 VDD.n3355 GND 0.0583f
C5986 VDD.n3359 GND 0.0134f
C5987 VDD.n3360 GND 0.047f
C5988 VDD.n3364 GND 0.0289f
C5989 VDD.n3365 GND 0.0135f
C5990 VDD.t30 GND 0.169f
C5991 VDD.n3375 GND 0.0735f
C5992 VDD.n3381 GND 0.0135f
C5993 VDD.n3382 GND 0.0287f
C5994 VDD.n3384 GND 0.0248f
C5995 VDD.n3385 GND 0.13f
C5996 VDD.n3386 GND 0.427f
C5997 VDD.n3412 GND 0.0443f
C5998 VDD.t729 GND 0.0187f
C5999 VDD.n3413 GND 0.0194f
C6000 VDD.n3414 GND 0.0239f
C6001 VDD.t1333 GND 0.0185f
C6002 VDD.n3415 GND 0.16f
C6003 VDD.n3416 GND 0.966f
C6004 VDD.n3417 GND 0.102f
C6005 VDD.n3418 GND 1.15f
C6006 VDD.n3419 GND 0.921f
C6007 VDD.t618 GND 0.0383f
C6008 VDD.t663 GND 0.0134f
C6009 VDD.n3420 GND 0.0699f
C6010 VDD.n3427 GND 0.0579f
C6011 VDD.n3428 GND 0.0223f
C6012 VDD.n3432 GND 0.0682f
C6013 VDD.n3434 GND 0.0779f
C6014 VDD.n3436 GND 0.0106f
C6015 VDD.t1355 GND 0.0288f
C6016 VDD.t1447 GND 0.0109f
C6017 VDD.n3447 GND 0.0397f
C6018 VDD.n3450 GND 0.0201f
C6019 VDD.n3451 GND 0.0133f
C6020 VDD.n3452 GND 0.114f
C6021 VDD.n3453 GND 0.0382f
C6022 VDD.n3458 GND 0.0681f
C6023 VDD.n3460 GND 0.0898f
C6024 VDD.n3468 GND 0.0865f
C6025 VDD.n3469 GND 0.0386f
C6026 VDD.n3474 GND 0.0419f
C6027 VDD.t538 GND 0.0681f
C6028 VDD.n3483 GND 0.295f
C6029 VDD.n3484 GND 0.165f
C6030 VDD.n3485 GND 0.0664f
C6031 VDD.n3486 GND 0.0215f
C6032 VDD.t411 GND 0.0855f
C6033 VDD.n3497 GND 0.0455f
C6034 VDD.n3498 GND 0.112f
C6035 VDD.n3500 GND 0.0121f
C6036 VDD.n3503 GND 0.0857f
C6037 VDD.n3504 GND 0.0898f
C6038 VDD.n3512 GND 0.0427f
C6039 VDD.n3516 GND 0.0386f
C6040 VDD.t18 GND 0.0681f
C6041 VDD.n3525 GND 0.0681f
C6042 VDD.n3527 GND 0.0875f
C6043 VDD.n3528 GND 0.28f
C6044 VDD.n3529 GND 0.166f
C6045 VDD.n3530 GND 0.196f
C6046 VDD.n3531 GND 0.0783f
C6047 VDD.n3532 GND 6.11f
C6048 VDD.n3533 GND 0.274f
C6049 VDD.n3534 GND 0.0237f
C6050 VDD.n3535 GND 0.0462f
C6051 VDD.t631 GND 0.0597f
C6052 VDD.n3547 GND 0.035f
C6053 VDD.n3555 GND 0.0437f
C6054 VDD.n3556 GND 0.0152f
C6055 VDD.n3557 GND 0.0128f
C6056 VDD.n3564 GND 0.0504f
C6057 VDD.n3580 GND 0.0735f
C6058 VDD.t194 GND 0.0597f
C6059 VDD.n3581 GND 0.035f
C6060 VDD.n3590 GND 0.0491f
C6061 VDD.n3592 GND 0.0135f
C6062 VDD.n3606 GND 0.0484f
C6063 VDD.n3607 GND 0.0582f
C6064 VDD.n3613 GND 0.0583f
C6065 VDD.n3617 GND 0.0134f
C6066 VDD.n3618 GND 0.047f
C6067 VDD.n3622 GND 0.0289f
C6068 VDD.n3623 GND 0.0135f
C6069 VDD.t214 GND 0.169f
C6070 VDD.n3633 GND 0.0735f
C6071 VDD.n3639 GND 0.0135f
C6072 VDD.n3640 GND 0.0287f
C6073 VDD.n3642 GND 0.0248f
C6074 VDD.n3643 GND 0.13f
C6075 VDD.n3644 GND 0.427f
C6076 VDD.n3670 GND 0.0443f
C6077 VDD.t191 GND 0.0187f
C6078 VDD.n3671 GND 0.0194f
C6079 VDD.n3672 GND 0.0239f
C6080 VDD.t633 GND 0.0185f
C6081 VDD.n3673 GND 0.16f
C6082 VDD.n3674 GND 0.966f
C6083 VDD.n3675 GND 0.102f
C6084 VDD.n3676 GND 1.15f
C6085 VDD.n3677 GND 0.921f
C6086 VDD.t515 GND 0.0383f
C6087 VDD.t1345 GND 0.0134f
C6088 VDD.n3678 GND 0.0699f
C6089 VDD.n3685 GND 0.0579f
C6090 VDD.n3686 GND 0.0223f
C6091 VDD.n3690 GND 0.0682f
C6092 VDD.n3692 GND 0.0779f
C6093 VDD.n3694 GND 0.0106f
C6094 VDD.t390 GND 0.0288f
C6095 VDD.t457 GND 0.0109f
C6096 VDD.n3705 GND 0.0397f
C6097 VDD.n3708 GND 0.0201f
C6098 VDD.n3709 GND 0.0133f
C6099 VDD.n3710 GND 0.114f
C6100 VDD.n3711 GND 0.0382f
C6101 VDD.n3716 GND 0.0681f
C6102 VDD.n3718 GND 0.0898f
C6103 VDD.n3726 GND 0.0865f
C6104 VDD.n3727 GND 0.0386f
C6105 VDD.n3732 GND 0.0419f
C6106 VDD.t413 GND 0.0681f
C6107 VDD.n3741 GND 0.295f
C6108 VDD.n3742 GND 0.165f
C6109 VDD.n3743 GND 0.0664f
C6110 VDD.n3744 GND 0.0215f
C6111 VDD.t410 GND 0.0855f
C6112 VDD.n3755 GND 0.0455f
C6113 VDD.n3756 GND 0.112f
C6114 VDD.n3758 GND 0.0121f
C6115 VDD.n3761 GND 0.0857f
C6116 VDD.n3762 GND 0.0898f
C6117 VDD.n3770 GND 0.0427f
C6118 VDD.n3774 GND 0.0386f
C6119 VDD.t82 GND 0.0681f
C6120 VDD.n3783 GND 0.0681f
C6121 VDD.n3785 GND 0.0875f
C6122 VDD.n3786 GND 0.28f
C6123 VDD.n3787 GND 0.166f
C6124 VDD.n3788 GND 0.196f
C6125 VDD.n3789 GND 0.0783f
C6126 VDD.n3790 GND 6.11f
C6127 VDD.n3791 GND 0.274f
C6128 VDD.n3792 GND 0.0237f
C6129 VDD.n3793 GND 0.0462f
C6130 VDD.t1386 GND 0.0597f
C6131 VDD.n3805 GND 0.035f
C6132 VDD.n3813 GND 0.0437f
C6133 VDD.n3814 GND 0.0152f
C6134 VDD.n3815 GND 0.0128f
C6135 VDD.n3822 GND 0.0504f
C6136 VDD.n3838 GND 0.0735f
C6137 VDD.t173 GND 0.0597f
C6138 VDD.n3839 GND 0.035f
C6139 VDD.n3848 GND 0.0491f
C6140 VDD.n3850 GND 0.0135f
C6141 VDD.n3864 GND 0.0484f
C6142 VDD.n3865 GND 0.0582f
C6143 VDD.n3871 GND 0.0583f
C6144 VDD.n3875 GND 0.0134f
C6145 VDD.n3876 GND 0.047f
C6146 VDD.n3880 GND 0.0289f
C6147 VDD.n3881 GND 0.0135f
C6148 VDD.t1027 GND 0.169f
C6149 VDD.n3891 GND 0.0735f
C6150 VDD.n3897 GND 0.0135f
C6151 VDD.n3898 GND 0.0287f
C6152 VDD.n3900 GND 0.0248f
C6153 VDD.n3901 GND 0.13f
C6154 VDD.n3902 GND 0.427f
C6155 VDD.n3928 GND 0.0443f
C6156 VDD.t171 GND 0.0187f
C6157 VDD.n3929 GND 0.0194f
C6158 VDD.n3930 GND 0.0239f
C6159 VDD.t1383 GND 0.0185f
C6160 VDD.n3931 GND 0.16f
C6161 VDD.n3932 GND 0.966f
C6162 VDD.n3933 GND 0.102f
C6163 VDD.n3934 GND 1.15f
C6164 VDD.n3935 GND 0.921f
C6165 VDD.t460 GND 0.0383f
C6166 VDD.t240 GND 0.0134f
C6167 VDD.n3936 GND 0.0699f
C6168 VDD.n3943 GND 0.0579f
C6169 VDD.n3944 GND 0.0223f
C6170 VDD.n3948 GND 0.0682f
C6171 VDD.n3950 GND 0.0779f
C6172 VDD.n3952 GND 0.0106f
C6173 VDD.t868 GND 0.0288f
C6174 VDD.t1441 GND 0.0109f
C6175 VDD.n3963 GND 0.0397f
C6176 VDD.n3966 GND 0.0201f
C6177 VDD.n3967 GND 0.0133f
C6178 VDD.n3968 GND 0.114f
C6179 VDD.n3969 GND 0.0382f
C6180 VDD.n3974 GND 0.0681f
C6181 VDD.n3976 GND 0.0898f
C6182 VDD.n3984 GND 0.0865f
C6183 VDD.n3985 GND 0.0386f
C6184 VDD.n3990 GND 0.0419f
C6185 VDD.t108 GND 0.0681f
C6186 VDD.n3999 GND 0.295f
C6187 VDD.n4000 GND 0.165f
C6188 VDD.n4001 GND 0.0664f
C6189 VDD.n4002 GND 0.0215f
C6190 VDD.t116 GND 0.0855f
C6191 VDD.n4013 GND 0.0455f
C6192 VDD.n4014 GND 0.112f
C6193 VDD.n4016 GND 0.0121f
C6194 VDD.n4019 GND 0.0857f
C6195 VDD.n4020 GND 0.0898f
C6196 VDD.n4028 GND 0.0427f
C6197 VDD.n4032 GND 0.0386f
C6198 VDD.t409 GND 0.0681f
C6199 VDD.n4041 GND 0.0681f
C6200 VDD.n4043 GND 0.0875f
C6201 VDD.n4044 GND 0.28f
C6202 VDD.n4045 GND 0.166f
C6203 VDD.n4046 GND 0.196f
C6204 VDD.n4047 GND 0.0783f
C6205 VDD.n4048 GND 6.11f
C6206 VDD.n4049 GND 0.274f
C6207 VDD.n4050 GND 0.0237f
C6208 VDD.n4051 GND 0.0462f
C6209 VDD.t888 GND 0.0597f
C6210 VDD.n4063 GND 0.035f
C6211 VDD.n4071 GND 0.0437f
C6212 VDD.n4072 GND 0.0152f
C6213 VDD.n4073 GND 0.0128f
C6214 VDD.n4080 GND 0.0504f
C6215 VDD.n4096 GND 0.0735f
C6216 VDD.t92 GND 0.0597f
C6217 VDD.n4097 GND 0.035f
C6218 VDD.n4106 GND 0.0491f
C6219 VDD.n4108 GND 0.0135f
C6220 VDD.n4122 GND 0.0484f
C6221 VDD.n4123 GND 0.0582f
C6222 VDD.n4129 GND 0.0583f
C6223 VDD.n4133 GND 0.0134f
C6224 VDD.n4134 GND 0.047f
C6225 VDD.n4138 GND 0.0289f
C6226 VDD.n4139 GND 0.0135f
C6227 VDD.t423 GND 0.169f
C6228 VDD.n4149 GND 0.0735f
C6229 VDD.n4155 GND 0.0135f
C6230 VDD.n4156 GND 0.0287f
C6231 VDD.n4158 GND 0.0248f
C6232 VDD.n4159 GND 0.13f
C6233 VDD.n4160 GND 0.427f
C6234 VDD.n4186 GND 0.0443f
C6235 VDD.t94 GND 0.0187f
C6236 VDD.n4187 GND 0.0194f
C6237 VDD.n4188 GND 0.0239f
C6238 VDD.t885 GND 0.0185f
C6239 VDD.n4189 GND 0.16f
C6240 VDD.n4190 GND 0.966f
C6241 VDD.n4191 GND 0.102f
C6242 VDD.n4192 GND 1.15f
C6243 VDD.n4193 GND 0.921f
C6244 VDD.t894 GND 0.0383f
C6245 VDD.t2 GND 0.0134f
C6246 VDD.n4194 GND 0.0699f
C6247 VDD.n4201 GND 0.0579f
C6248 VDD.n4202 GND 0.0223f
C6249 VDD.n4206 GND 0.0682f
C6250 VDD.n4208 GND 0.0779f
C6251 VDD.n4210 GND 0.0106f
C6252 VDD.t604 GND 0.0288f
C6253 VDD.t725 GND 0.0109f
C6254 VDD.n4221 GND 0.0397f
C6255 VDD.n4224 GND 0.0201f
C6256 VDD.n4225 GND 0.0133f
C6257 VDD.n4226 GND 0.114f
C6258 VDD.n4227 GND 0.0382f
C6259 VDD.n4232 GND 0.0681f
C6260 VDD.n4234 GND 0.0898f
C6261 VDD.n4242 GND 0.0865f
C6262 VDD.n4243 GND 0.0386f
C6263 VDD.n4248 GND 0.0419f
C6264 VDD.t0 GND 0.0681f
C6265 VDD.n4257 GND 0.295f
C6266 VDD.n4258 GND 0.165f
C6267 VDD.n4259 GND 0.0664f
C6268 VDD.n4260 GND 0.0215f
C6269 VDD.t489 GND 0.0855f
C6270 VDD.n4271 GND 0.0455f
C6271 VDD.n4272 GND 0.112f
C6272 VDD.n4274 GND 0.0121f
C6273 VDD.n4277 GND 0.0857f
C6274 VDD.n4278 GND 0.0898f
C6275 VDD.n4286 GND 0.0427f
C6276 VDD.n4290 GND 0.0386f
C6277 VDD.t727 GND 0.0681f
C6278 VDD.n4299 GND 0.0681f
C6279 VDD.n4301 GND 0.0875f
C6280 VDD.n4302 GND 0.28f
C6281 VDD.n4303 GND 0.166f
C6282 VDD.n4304 GND 0.196f
C6283 VDD.n4305 GND 0.0783f
C6284 VDD.n4306 GND 6.11f
C6285 VDD.n4307 GND 0.274f
C6286 VDD.n4308 GND 0.0237f
C6287 VDD.n4309 GND 0.0462f
C6288 VDD.t126 GND 0.0597f
C6289 VDD.n4321 GND 0.035f
C6290 VDD.n4329 GND 0.0437f
C6291 VDD.n4330 GND 0.0152f
C6292 VDD.n4331 GND 0.0128f
C6293 VDD.n4338 GND 0.0504f
C6294 VDD.n4354 GND 0.0735f
C6295 VDD.t497 GND 0.0597f
C6296 VDD.n4355 GND 0.035f
C6297 VDD.n4364 GND 0.0491f
C6298 VDD.n4366 GND 0.0135f
C6299 VDD.n4380 GND 0.0484f
C6300 VDD.n4381 GND 0.0582f
C6301 VDD.n4387 GND 0.0583f
C6302 VDD.n4391 GND 0.0134f
C6303 VDD.n4392 GND 0.047f
C6304 VDD.n4396 GND 0.0289f
C6305 VDD.n4397 GND 0.0135f
C6306 VDD.t1031 GND 0.169f
C6307 VDD.n4407 GND 0.0735f
C6308 VDD.n4413 GND 0.0135f
C6309 VDD.n4414 GND 0.0287f
C6310 VDD.n4416 GND 0.0248f
C6311 VDD.n4417 GND 0.13f
C6312 VDD.n4418 GND 0.427f
C6313 VDD.n4444 GND 0.0443f
C6314 VDD.t495 GND 0.0187f
C6315 VDD.n4445 GND 0.0194f
C6316 VDD.n4446 GND 0.0239f
C6317 VDD.t123 GND 0.0185f
C6318 VDD.n4447 GND 0.16f
C6319 VDD.n4448 GND 0.966f
C6320 VDD.n4449 GND 0.102f
C6321 VDD.n4450 GND 1.15f
C6322 VDD.n4451 GND 0.921f
C6323 VDD.t793 GND 0.0383f
C6324 VDD.t1186 GND 0.0134f
C6325 VDD.n4452 GND 0.0699f
C6326 VDD.n4459 GND 0.0579f
C6327 VDD.n4460 GND 0.0223f
C6328 VDD.n4464 GND 0.0682f
C6329 VDD.n4466 GND 0.0779f
C6330 VDD.n4468 GND 0.0106f
C6331 VDD.t1433 GND 0.0288f
C6332 VDD.t882 GND 0.0109f
C6333 VDD.n4479 GND 0.0397f
C6334 VDD.n4482 GND 0.0201f
C6335 VDD.n4483 GND 0.0133f
C6336 VDD.n4484 GND 0.114f
C6337 VDD.n4485 GND 0.0382f
C6338 VDD.n4490 GND 0.0681f
C6339 VDD.n4492 GND 0.0898f
C6340 VDD.n4500 GND 0.0865f
C6341 VDD.n4501 GND 0.0386f
C6342 VDD.n4506 GND 0.0419f
C6343 VDD.t13 GND 0.0681f
C6344 VDD.n4515 GND 0.295f
C6345 VDD.n4516 GND 0.165f
C6346 VDD.n4517 GND 0.0664f
C6347 VDD.n4518 GND 0.0215f
C6348 VDD.t84 GND 0.0855f
C6349 VDD.n4529 GND 0.0455f
C6350 VDD.n4530 GND 0.112f
C6351 VDD.n4532 GND 0.0121f
C6352 VDD.n4535 GND 0.0857f
C6353 VDD.n4536 GND 0.0898f
C6354 VDD.n4544 GND 0.0427f
C6355 VDD.n4548 GND 0.0386f
C6356 VDD.t122 GND 0.0681f
C6357 VDD.n4557 GND 0.0681f
C6358 VDD.n4559 GND 0.0875f
C6359 VDD.n4560 GND 0.28f
C6360 VDD.n4561 GND 0.166f
C6361 VDD.n4562 GND 0.196f
C6362 VDD.n4563 GND 0.0783f
C6363 VDD.n4564 GND 6.11f
C6364 VDD.n4565 GND 0.274f
C6365 VDD.n4566 GND 0.0237f
C6366 VDD.n4567 GND 0.0462f
C6367 VDD.t72 GND 0.0597f
C6368 VDD.n4579 GND 0.035f
C6369 VDD.n4587 GND 0.0437f
C6370 VDD.n4588 GND 0.0152f
C6371 VDD.n4589 GND 0.0128f
C6372 VDD.n4596 GND 0.0504f
C6373 VDD.n4612 GND 0.0735f
C6374 VDD.t587 GND 0.0597f
C6375 VDD.n4613 GND 0.035f
C6376 VDD.n4622 GND 0.0491f
C6377 VDD.n4624 GND 0.0135f
C6378 VDD.n4638 GND 0.0484f
C6379 VDD.n4639 GND 0.0582f
C6380 VDD.n4645 GND 0.0583f
C6381 VDD.n4649 GND 0.0134f
C6382 VDD.n4650 GND 0.047f
C6383 VDD.n4654 GND 0.0289f
C6384 VDD.n4655 GND 0.0135f
C6385 VDD.t402 GND 0.169f
C6386 VDD.n4665 GND 0.0735f
C6387 VDD.n4671 GND 0.0135f
C6388 VDD.n4672 GND 0.0287f
C6389 VDD.n4674 GND 0.0248f
C6390 VDD.n4675 GND 0.13f
C6391 VDD.n4676 GND 0.427f
C6392 VDD.n4702 GND 0.0443f
C6393 VDD.t585 GND 0.0187f
C6394 VDD.n4703 GND 0.0194f
C6395 VDD.n4704 GND 0.0239f
C6396 VDD.t74 GND 0.0185f
C6397 VDD.n4705 GND 0.16f
C6398 VDD.n4706 GND 0.966f
C6399 VDD.n4707 GND 0.102f
C6400 VDD.n4708 GND 1.15f
C6401 VDD.n4709 GND 0.921f
C6402 VDD.t23 GND 0.0383f
C6403 VDD.t1369 GND 0.0134f
C6404 VDD.n4710 GND 0.0699f
C6405 VDD.n4717 GND 0.0579f
C6406 VDD.n4718 GND 0.0223f
C6407 VDD.n4722 GND 0.0682f
C6408 VDD.n4724 GND 0.0779f
C6409 VDD.n4726 GND 0.0106f
C6410 VDD.t874 GND 0.0288f
C6411 VDD.t1347 GND 0.0109f
C6412 VDD.n4737 GND 0.0397f
C6413 VDD.n4740 GND 0.0201f
C6414 VDD.n4741 GND 0.0133f
C6415 VDD.n4742 GND 0.114f
C6416 VDD.n4743 GND 0.0382f
C6417 VDD.n4748 GND 0.0681f
C6418 VDD.n4750 GND 0.0898f
C6419 VDD.n4758 GND 0.0865f
C6420 VDD.n4759 GND 0.0386f
C6421 VDD.n4764 GND 0.0419f
C6422 VDD.t117 GND 0.0681f
C6423 VDD.n4773 GND 0.295f
C6424 VDD.n4774 GND 0.165f
C6425 VDD.n4775 GND 0.0664f
C6426 VDD.n4776 GND 0.0215f
C6427 VDD.t717 GND 0.0855f
C6428 VDD.n4787 GND 0.0455f
C6429 VDD.n4788 GND 0.112f
C6430 VDD.n4790 GND 0.0121f
C6431 VDD.n4793 GND 0.0857f
C6432 VDD.n4794 GND 0.0898f
C6433 VDD.n4802 GND 0.0427f
C6434 VDD.n4806 GND 0.0386f
C6435 VDD.t484 GND 0.0681f
C6436 VDD.n4815 GND 0.0681f
C6437 VDD.n4817 GND 0.0875f
C6438 VDD.n4818 GND 0.28f
C6439 VDD.n4819 GND 0.166f
C6440 VDD.n4820 GND 0.196f
C6441 VDD.n4821 GND 0.0783f
C6442 VDD.n4822 GND 6.11f
C6443 VDD.n4823 GND 0.274f
C6444 VDD.n4824 GND 0.0237f
C6445 VDD.n4825 GND 0.0462f
C6446 VDD.t783 GND 0.0597f
C6447 VDD.n4837 GND 0.035f
C6448 VDD.n4845 GND 0.0437f
C6449 VDD.n4846 GND 0.0152f
C6450 VDD.n4847 GND 0.0128f
C6451 VDD.n4854 GND 0.0504f
C6452 VDD.n4870 GND 0.0735f
C6453 VDD.t579 GND 0.0597f
C6454 VDD.n4871 GND 0.035f
C6455 VDD.n4880 GND 0.0491f
C6456 VDD.n4882 GND 0.0135f
C6457 VDD.n4896 GND 0.0484f
C6458 VDD.n4897 GND 0.0582f
C6459 VDD.n4903 GND 0.0583f
C6460 VDD.n4907 GND 0.0134f
C6461 VDD.n4908 GND 0.047f
C6462 VDD.n4912 GND 0.0289f
C6463 VDD.n4913 GND 0.0135f
C6464 VDD.t532 GND 0.169f
C6465 VDD.n4923 GND 0.0735f
C6466 VDD.n4929 GND 0.0135f
C6467 VDD.n4930 GND 0.0287f
C6468 VDD.n4932 GND 0.0248f
C6469 VDD.n4933 GND 0.13f
C6470 VDD.n4934 GND 0.427f
C6471 VDD.n4960 GND 0.0443f
C6472 VDD.t577 GND 0.0187f
C6473 VDD.n4961 GND 0.0194f
C6474 VDD.n4962 GND 0.0239f
C6475 VDD.t785 GND 0.0185f
C6476 VDD.n4963 GND 0.16f
C6477 VDD.n4964 GND 0.966f
C6478 VDD.n4965 GND 0.102f
C6479 VDD.n4966 GND 1.15f
C6480 VDD.n4967 GND 0.921f
C6481 VDD.t707 GND 0.0383f
C6482 VDD.t540 GND 0.0134f
C6483 VDD.n4968 GND 0.0699f
C6484 VDD.n4975 GND 0.0579f
C6485 VDD.n4976 GND 0.0223f
C6486 VDD.n4980 GND 0.0682f
C6487 VDD.n4982 GND 0.0779f
C6488 VDD.n4984 GND 0.0106f
C6489 VDD.t1435 GND 0.0288f
C6490 VDD.t739 GND 0.0109f
C6491 VDD.n4995 GND 0.0397f
C6492 VDD.n4998 GND 0.0201f
C6493 VDD.n4999 GND 0.0133f
C6494 VDD.n5000 GND 0.114f
C6495 VDD.n5001 GND 0.0382f
C6496 VDD.n5006 GND 0.0681f
C6497 VDD.n5008 GND 0.0898f
C6498 VDD.n5016 GND 0.0865f
C6499 VDD.n5017 GND 0.0386f
C6500 VDD.n5022 GND 0.0419f
C6501 VDD.t651 GND 0.0681f
C6502 VDD.n5031 GND 0.295f
C6503 VDD.n5032 GND 0.165f
C6504 VDD.n5033 GND 0.0664f
C6505 VDD.n5034 GND 0.0215f
C6506 VDD.t1353 GND 0.0855f
C6507 VDD.n5045 GND 0.0455f
C6508 VDD.n5046 GND 0.112f
C6509 VDD.n5048 GND 0.0121f
C6510 VDD.n5051 GND 0.0857f
C6511 VDD.n5052 GND 0.0898f
C6512 VDD.n5060 GND 0.0427f
C6513 VDD.n5064 GND 0.0386f
C6514 VDD.t14 GND 0.0681f
C6515 VDD.n5073 GND 0.0681f
C6516 VDD.n5075 GND 0.0875f
C6517 VDD.n5076 GND 0.28f
C6518 VDD.n5077 GND 0.166f
C6519 VDD.n5078 GND 0.196f
C6520 VDD.n5079 GND 0.0783f
C6521 VDD.n5080 GND 6.11f
C6522 VDD.n5081 GND 0.274f
C6523 VDD.n5082 GND 0.0237f
C6524 VDD.n5083 GND 0.0462f
C6525 VDD.t1374 GND 0.0597f
C6526 VDD.n5095 GND 0.035f
C6527 VDD.n5103 GND 0.0437f
C6528 VDD.n5104 GND 0.0152f
C6529 VDD.n5105 GND 0.0128f
C6530 VDD.n5112 GND 0.0504f
C6531 VDD.n5128 GND 0.0735f
C6532 VDD.t857 GND 0.0597f
C6533 VDD.n5129 GND 0.035f
C6534 VDD.n5138 GND 0.0491f
C6535 VDD.n5140 GND 0.0135f
C6536 VDD.n5154 GND 0.0484f
C6537 VDD.n5155 GND 0.0582f
C6538 VDD.n5161 GND 0.0583f
C6539 VDD.n5165 GND 0.0134f
C6540 VDD.n5166 GND 0.047f
C6541 VDD.n5170 GND 0.0289f
C6542 VDD.n5171 GND 0.0135f
C6543 VDD.t381 GND 0.169f
C6544 VDD.n5181 GND 0.0735f
C6545 VDD.n5187 GND 0.0135f
C6546 VDD.n5188 GND 0.0287f
C6547 VDD.n5190 GND 0.0248f
C6548 VDD.n5191 GND 0.13f
C6549 VDD.n5192 GND 0.427f
C6550 VDD.n5218 GND 0.0443f
C6551 VDD.t855 GND 0.0187f
C6552 VDD.n5219 GND 0.0194f
C6553 VDD.n5220 GND 0.0239f
C6554 VDD.t1371 GND 0.0185f
C6555 VDD.n5221 GND 0.16f
C6556 VDD.n5222 GND 0.966f
C6557 VDD.n5223 GND 0.102f
C6558 VDD.n5224 GND 1.15f
C6559 VDD.n5225 GND 0.921f
C6560 VDD.t199 GND 0.0383f
C6561 VDD.t1184 GND 0.0134f
C6562 VDD.n5226 GND 0.0699f
C6563 VDD.n5233 GND 0.0579f
C6564 VDD.n5234 GND 0.0223f
C6565 VDD.n5238 GND 0.0682f
C6566 VDD.n5240 GND 0.0779f
C6567 VDD.n5242 GND 0.0106f
C6568 VDD.t153 GND 0.0288f
C6569 VDD.t236 GND 0.0109f
C6570 VDD.n5253 GND 0.0397f
C6571 VDD.n5256 GND 0.0201f
C6572 VDD.n5257 GND 0.0133f
C6573 VDD.n5258 GND 0.114f
C6574 VDD.n5259 GND 0.0382f
C6575 VDD.n5264 GND 0.0681f
C6576 VDD.n5266 GND 0.0898f
C6577 VDD.n5274 GND 0.0865f
C6578 VDD.n5275 GND 0.0386f
C6579 VDD.n5280 GND 0.0419f
C6580 VDD.t85 GND 0.0681f
C6581 VDD.n5289 GND 0.295f
C6582 VDD.n5290 GND 0.165f
C6583 VDD.n5291 GND 0.0664f
C6584 VDD.n5292 GND 0.0215f
C6585 VDD.t529 GND 0.0855f
C6586 VDD.n5303 GND 0.0455f
C6587 VDD.n5304 GND 0.112f
C6588 VDD.n5306 GND 0.0121f
C6589 VDD.n5309 GND 0.0857f
C6590 VDD.n5310 GND 0.0898f
C6591 VDD.n5318 GND 0.0427f
C6592 VDD.n5322 GND 0.0386f
C6593 VDD.t119 GND 0.0681f
C6594 VDD.n5331 GND 0.0681f
C6595 VDD.n5333 GND 0.0875f
C6596 VDD.n5334 GND 0.28f
C6597 VDD.n5335 GND 0.166f
C6598 VDD.n5336 GND 0.196f
C6599 VDD.n5337 GND 0.0783f
C6600 VDD.n5338 GND 9.87f
C6601 VDD.n5339 GND 22.6f
C6602 VDD.n5340 GND 14f
C6603 VDD.n5341 GND 14f
C6604 VDD.n5342 GND 14f
C6605 VDD.n5343 GND 14f
C6606 VDD.n5344 GND 14.5f
C6607 VDD.n5345 GND 0.0237f
C6608 VDD.n5346 GND 0.0462f
C6609 VDD.t6 GND 0.0597f
C6610 VDD.n5358 GND 0.035f
C6611 VDD.n5366 GND 0.0437f
C6612 VDD.n5367 GND 0.0152f
C6613 VDD.n5368 GND 0.0128f
C6614 VDD.n5375 GND 0.0504f
C6615 VDD.n5391 GND 0.0735f
C6616 VDD.t517 GND 0.0597f
C6617 VDD.n5392 GND 0.035f
C6618 VDD.n5401 GND 0.0491f
C6619 VDD.n5403 GND 0.0135f
C6620 VDD.n5417 GND 0.0484f
C6621 VDD.n5418 GND 0.0582f
C6622 VDD.n5424 GND 0.0583f
C6623 VDD.n5428 GND 0.0134f
C6624 VDD.n5429 GND 0.047f
C6625 VDD.n5433 GND 0.0289f
C6626 VDD.n5434 GND 0.0135f
C6627 VDD.t709 GND 0.169f
C6628 VDD.n5444 GND 0.0735f
C6629 VDD.n5450 GND 0.0135f
C6630 VDD.n5451 GND 0.0287f
C6631 VDD.n5453 GND 0.0248f
C6632 VDD.n5454 GND 0.926f
C6633 VDD.n5455 GND 1.67f
C6634 VDD.n5481 GND 0.0443f
C6635 VDD.t519 GND 0.0187f
C6636 VDD.n5482 GND 0.0194f
C6637 VDD.n5483 GND 0.0239f
C6638 VDD.t4 GND 0.0185f
C6639 VDD.n5484 GND 0.169f
C6640 VDD.n5485 GND 1.7f
C6641 VDD.t1486 GND 0.0383f
C6642 VDD.t188 GND 0.0134f
C6643 VDD.n5486 GND 0.0699f
C6644 VDD.n5493 GND 0.0579f
C6645 VDD.n5494 GND 0.0223f
C6646 VDD.n5498 GND 0.0682f
C6647 VDD.n5500 GND 0.0779f
C6648 VDD.n5502 GND 0.0106f
C6649 VDD.t813 GND 0.0288f
C6650 VDD.t86 GND 0.0109f
C6651 VDD.n5513 GND 0.0397f
C6652 VDD.n5516 GND 0.0201f
C6653 VDD.n5517 GND 0.0133f
C6654 VDD.n5518 GND 0.114f
C6655 VDD.n5519 GND 0.0382f
C6656 VDD.n5524 GND 0.0681f
C6657 VDD.n5526 GND 0.0898f
C6658 VDD.n5534 GND 0.0865f
C6659 VDD.n5535 GND 0.0386f
C6660 VDD.n5540 GND 0.0419f
C6661 VDD.t186 GND 0.0681f
C6662 VDD.n5549 GND 0.295f
C6663 VDD.n5550 GND 0.165f
C6664 VDD.n5551 GND 0.0664f
C6665 VDD.n5552 GND 0.0215f
C6666 VDD.t482 GND 0.0855f
C6667 VDD.n5563 GND 0.0455f
C6668 VDD.n5564 GND 0.112f
C6669 VDD.n5566 GND 0.0121f
C6670 VDD.n5569 GND 0.0857f
C6671 VDD.n5570 GND 0.0898f
C6672 VDD.n5578 GND 0.0427f
C6673 VDD.n5582 GND 0.0386f
C6674 VDD.t88 GND 0.0681f
C6675 VDD.n5591 GND 0.0681f
C6676 VDD.n5593 GND 0.0875f
C6677 VDD.n5594 GND 0.28f
C6678 VDD.n5595 GND 0.166f
C6679 VDD.n5596 GND 1.98f
C6680 VDD.n5597 GND 6.4f
C6681 VDD.n5598 GND 11.2f
C6682 VDD.n5599 GND 0.0237f
C6683 VDD.n5600 GND 0.0462f
C6684 VDD.t613 GND 0.0597f
C6685 VDD.n5612 GND 0.035f
C6686 VDD.n5620 GND 0.0437f
C6687 VDD.n5621 GND 0.0152f
C6688 VDD.n5622 GND 0.0128f
C6689 VDD.n5629 GND 0.0504f
C6690 VDD.n5645 GND 0.0735f
C6691 VDD.t164 GND 0.0597f
C6692 VDD.n5646 GND 0.035f
C6693 VDD.n5655 GND 0.0491f
C6694 VDD.n5657 GND 0.0135f
C6695 VDD.n5671 GND 0.0484f
C6696 VDD.n5672 GND 0.0582f
C6697 VDD.n5678 GND 0.0583f
C6698 VDD.n5682 GND 0.0134f
C6699 VDD.n5683 GND 0.047f
C6700 VDD.n5687 GND 0.0289f
C6701 VDD.n5688 GND 0.0135f
C6702 VDD.t870 GND 0.169f
C6703 VDD.n5698 GND 0.0735f
C6704 VDD.n5704 GND 0.0135f
C6705 VDD.n5705 GND 0.0287f
C6706 VDD.n5707 GND 0.0248f
C6707 VDD.n5708 GND 0.926f
C6708 VDD.n5709 GND 1.67f
C6709 VDD.n5735 GND 0.0443f
C6710 VDD.t162 GND 0.0187f
C6711 VDD.n5736 GND 0.0194f
C6712 VDD.n5737 GND 0.0239f
C6713 VDD.t610 GND 0.0185f
C6714 VDD.n5738 GND 0.169f
C6715 VDD.n5739 GND 1.7f
C6716 VDD.t575 GND 0.0383f
C6717 VDD.t90 GND 0.0134f
C6718 VDD.n5740 GND 0.0699f
C6719 VDD.n5747 GND 0.0579f
C6720 VDD.n5748 GND 0.0223f
C6721 VDD.n5752 GND 0.0682f
C6722 VDD.n5754 GND 0.0779f
C6723 VDD.n5756 GND 0.0106f
C6724 VDD.t417 GND 0.0288f
C6725 VDD.t1195 GND 0.0109f
C6726 VDD.n5767 GND 0.0397f
C6727 VDD.n5770 GND 0.0201f
C6728 VDD.n5771 GND 0.0133f
C6729 VDD.n5772 GND 0.114f
C6730 VDD.n5773 GND 0.0382f
C6731 VDD.n5778 GND 0.0681f
C6732 VDD.n5780 GND 0.0898f
C6733 VDD.n5788 GND 0.0865f
C6734 VDD.n5789 GND 0.0386f
C6735 VDD.n5794 GND 0.0419f
C6736 VDD.t109 GND 0.0681f
C6737 VDD.n5803 GND 0.295f
C6738 VDD.n5804 GND 0.165f
C6739 VDD.n5805 GND 0.0664f
C6740 VDD.n5806 GND 0.0215f
C6741 VDD.t530 GND 0.0855f
C6742 VDD.n5817 GND 0.0455f
C6743 VDD.n5818 GND 0.112f
C6744 VDD.n5820 GND 0.0121f
C6745 VDD.n5823 GND 0.0857f
C6746 VDD.n5824 GND 0.0898f
C6747 VDD.n5832 GND 0.0427f
C6748 VDD.n5836 GND 0.0386f
C6749 VDD.t746 GND 0.0681f
C6750 VDD.n5845 GND 0.0681f
C6751 VDD.n5847 GND 0.0875f
C6752 VDD.n5848 GND 0.28f
C6753 VDD.n5849 GND 0.166f
C6754 VDD.n5850 GND 1.98f
C6755 VDD.n5851 GND 6.4f
C6756 VDD.n5852 GND 11.2f
C6757 VDD.n5853 GND 14.5f
C6758 VDD.n5854 GND 14f
C6759 VDD.n5855 GND 14f
C6760 VDD.n5856 GND 14f
C6761 VDD.n5857 GND 14f
C6762 VDD.n5858 GND 10.2f
C6763 VDD.n5859 GND 7.31f
C6764 VDD.n5860 GND 20.4f
C6765 VDD.n5861 GND 34.2f
C6766 VDD.n5862 GND 10.2f
C6767 VDD.n5863 GND 14.2f
.ends

