magic
tech sky130A
magscale 1 2
timestamp 1714790421
<< error_p >>
rect -573 34 573 36
<< pwell >>
rect -739 -632 739 632
<< psubdiff >>
rect -703 562 -607 596
rect 607 562 703 596
rect -703 500 -669 562
rect 669 500 703 562
rect -703 -562 -669 -500
rect 669 -562 703 -500
rect -703 -596 -607 -562
rect 607 -596 703 -562
<< psubdiffcont >>
rect -607 562 607 596
rect -703 -500 -669 500
rect 669 -500 703 500
rect -607 -596 607 -562
<< xpolycontact >>
rect -573 34 573 466
rect -573 -466 573 -34
<< xpolyres >>
rect -573 -34 573 34
<< locali >>
rect -703 562 -607 596
rect 607 562 703 596
rect -703 500 -669 562
rect 669 500 703 562
rect -703 -562 -669 -500
rect 669 -562 703 -500
rect -703 -596 -607 -562
rect 607 -596 703 -562
<< viali >>
rect -557 51 557 448
rect -557 -448 557 -51
<< metal1 >>
rect -569 448 569 454
rect -569 51 -557 448
rect 557 51 569 448
rect -569 45 569 51
rect -569 -51 569 -45
rect -569 -448 -557 -51
rect 557 -448 569 -51
rect -569 -454 569 -448
<< properties >>
string FIXED_BBOX -686 -579 686 579
string gencell sky130_fd_pr__res_xhigh_po_5p73
string library sky130
string parameters w 5.73 l 0.5 m 1 nx 1 wmin 5.730 lmin 0.50 rho 2000 val 240.209 dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 5.730 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
