magic
tech sky130A
magscale 1 2
timestamp 1682173151
<< nwell >>
rect 42138 689988 48798 694738
rect 41638 681839 49308 683080
rect 41660 681838 49278 681839
<< pwell >>
rect 38335 692595 41531 695533
rect 49405 692595 52601 695533
rect 44757 688449 46197 689869
rect 44757 686929 46197 688349
rect 43758 685408 47188 686828
rect 43502 683888 47448 685308
rect 44434 681048 46508 681640
rect 44650 680523 46288 681015
rect 41713 679898 49223 680490
rect 42178 673578 48758 678890
rect 42188 666076 48758 673578
<< nmos >>
rect 44953 688659 45053 689659
rect 45111 688659 45211 689659
rect 45269 688659 45369 689659
rect 45427 688659 45527 689659
rect 45585 688659 45685 689659
rect 45743 688659 45843 689659
rect 45901 688659 46001 689659
rect 44953 687139 45053 688139
rect 45111 687139 45211 688139
rect 45269 687139 45369 688139
rect 45427 687139 45527 688139
rect 45585 687139 45685 688139
rect 45743 687139 45843 688139
rect 45901 687139 46001 688139
rect 43954 685618 44154 686618
rect 44212 685618 44412 686618
rect 44470 685618 44670 686618
rect 44728 685618 44928 686618
rect 44986 685618 45186 686618
rect 45244 685618 45444 686618
rect 45502 685618 45702 686618
rect 45760 685618 45960 686618
rect 46018 685618 46218 686618
rect 46276 685618 46476 686618
rect 46534 685618 46734 686618
rect 46792 685618 46992 686618
rect 43698 684098 43898 685098
rect 43956 684098 44156 685098
rect 44214 684098 44414 685098
rect 44472 684098 44672 685098
rect 44730 684098 44930 685098
rect 44988 684098 45188 685098
rect 45246 684098 45446 685098
rect 45504 684098 45704 685098
rect 45762 684098 45962 685098
rect 46020 684098 46220 685098
rect 46278 684098 46478 685098
rect 46536 684098 46736 685098
rect 46794 684098 46994 685098
rect 47052 684098 47252 685098
rect 44644 681244 44894 681444
rect 45112 681244 45362 681444
rect 45580 681244 45830 681444
rect 46048 681244 46298 681444
rect 44860 680719 45360 680819
rect 45578 680719 46078 680819
rect 41923 680094 42923 680294
rect 43141 680094 44141 680294
rect 44359 680094 45359 680294
rect 45577 680094 46577 680294
rect 46795 680094 47795 680294
rect 48013 680094 49013 680294
<< pmos >>
rect 42340 693437 42440 694437
rect 42498 693437 42598 694437
rect 42656 693437 42756 694437
rect 42814 693437 42914 694437
rect 42972 693437 43072 694437
rect 43130 693437 43230 694437
rect 43288 693437 43388 694437
rect 43446 693437 43546 694437
rect 43604 693437 43704 694437
rect 43762 693437 43862 694437
rect 43920 693437 44020 694437
rect 44078 693437 44178 694437
rect 44236 693437 44336 694437
rect 44394 693437 44494 694437
rect 44552 693437 44652 694437
rect 44710 693437 44810 694437
rect 44868 693437 44968 694437
rect 45026 693437 45126 694437
rect 45184 693437 45284 694437
rect 45342 693437 45442 694437
rect 45500 693437 45600 694437
rect 45658 693437 45758 694437
rect 45816 693437 45916 694437
rect 45974 693437 46074 694437
rect 46132 693437 46232 694437
rect 46290 693437 46390 694437
rect 46448 693437 46548 694437
rect 46606 693437 46706 694437
rect 46764 693437 46864 694437
rect 46922 693437 47022 694437
rect 47080 693437 47180 694437
rect 47238 693437 47338 694437
rect 47396 693437 47496 694437
rect 47554 693437 47654 694437
rect 47712 693437 47812 694437
rect 47870 693437 47970 694437
rect 48028 693437 48128 694437
rect 48186 693437 48286 694437
rect 48344 693437 48444 694437
rect 48502 693437 48602 694437
rect 43842 691767 43942 692767
rect 44000 691767 44100 692767
rect 44158 691767 44258 692767
rect 44316 691767 44416 692767
rect 44474 691767 44574 692767
rect 44632 691767 44732 692767
rect 44790 691767 44890 692767
rect 44948 691767 45048 692767
rect 45106 691767 45206 692767
rect 45264 691767 45364 692767
rect 45422 691767 45522 692767
rect 45580 691767 45680 692767
rect 45738 691767 45838 692767
rect 45896 691767 45996 692767
rect 46054 691767 46154 692767
rect 46212 691767 46312 692767
rect 46370 691767 46470 692767
rect 46528 691767 46628 692767
rect 46686 691767 46786 692767
rect 46844 691767 46944 692767
rect 47002 691767 47102 692767
rect 43842 690227 43942 691227
rect 44000 690227 44100 691227
rect 44158 690227 44258 691227
rect 44316 690227 44416 691227
rect 44474 690227 44574 691227
rect 44632 690227 44732 691227
rect 44790 690227 44890 691227
rect 44948 690227 45048 691227
rect 45106 690227 45206 691227
rect 45264 690227 45364 691227
rect 45422 690227 45522 691227
rect 45580 690227 45680 691227
rect 45738 690227 45838 691227
rect 45896 690227 45996 691227
rect 46054 690227 46154 691227
rect 46212 690227 46312 691227
rect 46370 690227 46470 691227
rect 46528 690227 46628 691227
rect 46686 690227 46786 691227
rect 46844 690227 46944 691227
rect 47002 690227 47102 691227
rect 41879 682624 42879 682824
rect 43115 682624 44115 682824
rect 44351 682624 45351 682824
rect 45587 682624 46587 682824
rect 46823 682624 47823 682824
rect 48059 682624 49059 682824
rect 41879 682034 42879 682234
rect 43115 682034 44115 682234
rect 44351 682034 45351 682234
rect 45587 682034 46587 682234
rect 46823 682034 47823 682234
rect 48059 682034 49059 682234
<< ndiff >>
rect 44895 689647 44953 689659
rect 44895 688671 44907 689647
rect 44941 688671 44953 689647
rect 44895 688659 44953 688671
rect 45053 689647 45111 689659
rect 45053 688671 45065 689647
rect 45099 688671 45111 689647
rect 45053 688659 45111 688671
rect 45211 689647 45269 689659
rect 45211 688671 45223 689647
rect 45257 688671 45269 689647
rect 45211 688659 45269 688671
rect 45369 689647 45427 689659
rect 45369 688671 45381 689647
rect 45415 688671 45427 689647
rect 45369 688659 45427 688671
rect 45527 689647 45585 689659
rect 45527 688671 45539 689647
rect 45573 688671 45585 689647
rect 45527 688659 45585 688671
rect 45685 689647 45743 689659
rect 45685 688671 45697 689647
rect 45731 688671 45743 689647
rect 45685 688659 45743 688671
rect 45843 689647 45901 689659
rect 45843 688671 45855 689647
rect 45889 688671 45901 689647
rect 45843 688659 45901 688671
rect 46001 689647 46059 689659
rect 46001 688671 46013 689647
rect 46047 688671 46059 689647
rect 46001 688659 46059 688671
rect 44895 688127 44953 688139
rect 44895 687151 44907 688127
rect 44941 687151 44953 688127
rect 44895 687139 44953 687151
rect 45053 688127 45111 688139
rect 45053 687151 45065 688127
rect 45099 687151 45111 688127
rect 45053 687139 45111 687151
rect 45211 688127 45269 688139
rect 45211 687151 45223 688127
rect 45257 687151 45269 688127
rect 45211 687139 45269 687151
rect 45369 688127 45427 688139
rect 45369 687151 45381 688127
rect 45415 687151 45427 688127
rect 45369 687139 45427 687151
rect 45527 688127 45585 688139
rect 45527 687151 45539 688127
rect 45573 687151 45585 688127
rect 45527 687139 45585 687151
rect 45685 688127 45743 688139
rect 45685 687151 45697 688127
rect 45731 687151 45743 688127
rect 45685 687139 45743 687151
rect 45843 688127 45901 688139
rect 45843 687151 45855 688127
rect 45889 687151 45901 688127
rect 45843 687139 45901 687151
rect 46001 688127 46059 688139
rect 46001 687151 46013 688127
rect 46047 687151 46059 688127
rect 46001 687139 46059 687151
rect 43896 686606 43954 686618
rect 43896 685630 43908 686606
rect 43942 685630 43954 686606
rect 43896 685618 43954 685630
rect 44154 686606 44212 686618
rect 44154 685630 44166 686606
rect 44200 685630 44212 686606
rect 44154 685618 44212 685630
rect 44412 686606 44470 686618
rect 44412 685630 44424 686606
rect 44458 685630 44470 686606
rect 44412 685618 44470 685630
rect 44670 686606 44728 686618
rect 44670 685630 44682 686606
rect 44716 685630 44728 686606
rect 44670 685618 44728 685630
rect 44928 686606 44986 686618
rect 44928 685630 44940 686606
rect 44974 685630 44986 686606
rect 44928 685618 44986 685630
rect 45186 686606 45244 686618
rect 45186 685630 45198 686606
rect 45232 685630 45244 686606
rect 45186 685618 45244 685630
rect 45444 686606 45502 686618
rect 45444 685630 45456 686606
rect 45490 685630 45502 686606
rect 45444 685618 45502 685630
rect 45702 686606 45760 686618
rect 45702 685630 45714 686606
rect 45748 685630 45760 686606
rect 45702 685618 45760 685630
rect 45960 686606 46018 686618
rect 45960 685630 45972 686606
rect 46006 685630 46018 686606
rect 45960 685618 46018 685630
rect 46218 686606 46276 686618
rect 46218 685630 46230 686606
rect 46264 685630 46276 686606
rect 46218 685618 46276 685630
rect 46476 686606 46534 686618
rect 46476 685630 46488 686606
rect 46522 685630 46534 686606
rect 46476 685618 46534 685630
rect 46734 686606 46792 686618
rect 46734 685630 46746 686606
rect 46780 685630 46792 686606
rect 46734 685618 46792 685630
rect 46992 686606 47050 686618
rect 46992 685630 47004 686606
rect 47038 685630 47050 686606
rect 46992 685618 47050 685630
rect 43640 685086 43698 685098
rect 43640 684110 43652 685086
rect 43686 684110 43698 685086
rect 43640 684098 43698 684110
rect 43898 685086 43956 685098
rect 43898 684110 43910 685086
rect 43944 684110 43956 685086
rect 43898 684098 43956 684110
rect 44156 685086 44214 685098
rect 44156 684110 44168 685086
rect 44202 684110 44214 685086
rect 44156 684098 44214 684110
rect 44414 685086 44472 685098
rect 44414 684110 44426 685086
rect 44460 684110 44472 685086
rect 44414 684098 44472 684110
rect 44672 685086 44730 685098
rect 44672 684110 44684 685086
rect 44718 684110 44730 685086
rect 44672 684098 44730 684110
rect 44930 685086 44988 685098
rect 44930 684110 44942 685086
rect 44976 684110 44988 685086
rect 44930 684098 44988 684110
rect 45188 685086 45246 685098
rect 45188 684110 45200 685086
rect 45234 684110 45246 685086
rect 45188 684098 45246 684110
rect 45446 685086 45504 685098
rect 45446 684110 45458 685086
rect 45492 684110 45504 685086
rect 45446 684098 45504 684110
rect 45704 685086 45762 685098
rect 45704 684110 45716 685086
rect 45750 684110 45762 685086
rect 45704 684098 45762 684110
rect 45962 685086 46020 685098
rect 45962 684110 45974 685086
rect 46008 684110 46020 685086
rect 45962 684098 46020 684110
rect 46220 685086 46278 685098
rect 46220 684110 46232 685086
rect 46266 684110 46278 685086
rect 46220 684098 46278 684110
rect 46478 685086 46536 685098
rect 46478 684110 46490 685086
rect 46524 684110 46536 685086
rect 46478 684098 46536 684110
rect 46736 685086 46794 685098
rect 46736 684110 46748 685086
rect 46782 684110 46794 685086
rect 46736 684098 46794 684110
rect 46994 685086 47052 685098
rect 46994 684110 47006 685086
rect 47040 684110 47052 685086
rect 46994 684098 47052 684110
rect 47252 685086 47310 685098
rect 47252 684110 47264 685086
rect 47298 684110 47310 685086
rect 47252 684098 47310 684110
rect 44644 681490 44894 681502
rect 44644 681456 44656 681490
rect 44882 681456 44894 681490
rect 44644 681444 44894 681456
rect 45112 681490 45362 681502
rect 45112 681456 45124 681490
rect 45350 681456 45362 681490
rect 45112 681444 45362 681456
rect 45580 681490 45830 681502
rect 45580 681456 45592 681490
rect 45818 681456 45830 681490
rect 45580 681444 45830 681456
rect 46048 681490 46298 681502
rect 46048 681456 46060 681490
rect 46286 681456 46298 681490
rect 46048 681444 46298 681456
rect 44644 681232 44894 681244
rect 44644 681198 44656 681232
rect 44882 681198 44894 681232
rect 44644 681186 44894 681198
rect 45112 681232 45362 681244
rect 45112 681198 45124 681232
rect 45350 681198 45362 681232
rect 45112 681186 45362 681198
rect 45580 681232 45830 681244
rect 45580 681198 45592 681232
rect 45818 681198 45830 681232
rect 45580 681186 45830 681198
rect 46048 681232 46298 681244
rect 46048 681198 46060 681232
rect 46286 681198 46298 681232
rect 46048 681186 46298 681198
rect 44860 680865 45360 680877
rect 44860 680831 44872 680865
rect 45348 680831 45360 680865
rect 44860 680819 45360 680831
rect 45578 680865 46078 680877
rect 45578 680831 45590 680865
rect 46066 680831 46078 680865
rect 45578 680819 46078 680831
rect 44860 680707 45360 680719
rect 44860 680673 44872 680707
rect 45348 680673 45360 680707
rect 44860 680661 45360 680673
rect 45578 680707 46078 680719
rect 45578 680673 45590 680707
rect 46066 680673 46078 680707
rect 45578 680661 46078 680673
rect 41923 680340 42923 680352
rect 41923 680306 41935 680340
rect 42911 680306 42923 680340
rect 41923 680294 42923 680306
rect 43141 680340 44141 680352
rect 43141 680306 43153 680340
rect 44129 680306 44141 680340
rect 43141 680294 44141 680306
rect 44359 680340 45359 680352
rect 44359 680306 44371 680340
rect 45347 680306 45359 680340
rect 44359 680294 45359 680306
rect 45577 680340 46577 680352
rect 45577 680306 45589 680340
rect 46565 680306 46577 680340
rect 45577 680294 46577 680306
rect 46795 680340 47795 680352
rect 46795 680306 46807 680340
rect 47783 680306 47795 680340
rect 46795 680294 47795 680306
rect 48013 680340 49013 680352
rect 48013 680306 48025 680340
rect 49001 680306 49013 680340
rect 48013 680294 49013 680306
rect 41923 680082 42923 680094
rect 41923 680048 41935 680082
rect 42911 680048 42923 680082
rect 41923 680036 42923 680048
rect 43141 680082 44141 680094
rect 43141 680048 43153 680082
rect 44129 680048 44141 680082
rect 43141 680036 44141 680048
rect 44359 680082 45359 680094
rect 44359 680048 44371 680082
rect 45347 680048 45359 680082
rect 44359 680036 45359 680048
rect 45577 680082 46577 680094
rect 45577 680048 45589 680082
rect 46565 680048 46577 680082
rect 45577 680036 46577 680048
rect 46795 680082 47795 680094
rect 46795 680048 46807 680082
rect 47783 680048 47795 680082
rect 46795 680036 47795 680048
rect 48013 680082 49013 680094
rect 48013 680048 48025 680082
rect 49001 680048 49013 680082
rect 48013 680036 49013 680048
<< pdiff >>
rect 42282 694425 42340 694437
rect 42282 693449 42294 694425
rect 42328 693449 42340 694425
rect 42282 693437 42340 693449
rect 42440 694425 42498 694437
rect 42440 693449 42452 694425
rect 42486 693449 42498 694425
rect 42440 693437 42498 693449
rect 42598 694425 42656 694437
rect 42598 693449 42610 694425
rect 42644 693449 42656 694425
rect 42598 693437 42656 693449
rect 42756 694425 42814 694437
rect 42756 693449 42768 694425
rect 42802 693449 42814 694425
rect 42756 693437 42814 693449
rect 42914 694425 42972 694437
rect 42914 693449 42926 694425
rect 42960 693449 42972 694425
rect 42914 693437 42972 693449
rect 43072 694425 43130 694437
rect 43072 693449 43084 694425
rect 43118 693449 43130 694425
rect 43072 693437 43130 693449
rect 43230 694425 43288 694437
rect 43230 693449 43242 694425
rect 43276 693449 43288 694425
rect 43230 693437 43288 693449
rect 43388 694425 43446 694437
rect 43388 693449 43400 694425
rect 43434 693449 43446 694425
rect 43388 693437 43446 693449
rect 43546 694425 43604 694437
rect 43546 693449 43558 694425
rect 43592 693449 43604 694425
rect 43546 693437 43604 693449
rect 43704 694425 43762 694437
rect 43704 693449 43716 694425
rect 43750 693449 43762 694425
rect 43704 693437 43762 693449
rect 43862 694425 43920 694437
rect 43862 693449 43874 694425
rect 43908 693449 43920 694425
rect 43862 693437 43920 693449
rect 44020 694425 44078 694437
rect 44020 693449 44032 694425
rect 44066 693449 44078 694425
rect 44020 693437 44078 693449
rect 44178 694425 44236 694437
rect 44178 693449 44190 694425
rect 44224 693449 44236 694425
rect 44178 693437 44236 693449
rect 44336 694425 44394 694437
rect 44336 693449 44348 694425
rect 44382 693449 44394 694425
rect 44336 693437 44394 693449
rect 44494 694425 44552 694437
rect 44494 693449 44506 694425
rect 44540 693449 44552 694425
rect 44494 693437 44552 693449
rect 44652 694425 44710 694437
rect 44652 693449 44664 694425
rect 44698 693449 44710 694425
rect 44652 693437 44710 693449
rect 44810 694425 44868 694437
rect 44810 693449 44822 694425
rect 44856 693449 44868 694425
rect 44810 693437 44868 693449
rect 44968 694425 45026 694437
rect 44968 693449 44980 694425
rect 45014 693449 45026 694425
rect 44968 693437 45026 693449
rect 45126 694425 45184 694437
rect 45126 693449 45138 694425
rect 45172 693449 45184 694425
rect 45126 693437 45184 693449
rect 45284 694425 45342 694437
rect 45284 693449 45296 694425
rect 45330 693449 45342 694425
rect 45284 693437 45342 693449
rect 45442 694425 45500 694437
rect 45442 693449 45454 694425
rect 45488 693449 45500 694425
rect 45442 693437 45500 693449
rect 45600 694425 45658 694437
rect 45600 693449 45612 694425
rect 45646 693449 45658 694425
rect 45600 693437 45658 693449
rect 45758 694425 45816 694437
rect 45758 693449 45770 694425
rect 45804 693449 45816 694425
rect 45758 693437 45816 693449
rect 45916 694425 45974 694437
rect 45916 693449 45928 694425
rect 45962 693449 45974 694425
rect 45916 693437 45974 693449
rect 46074 694425 46132 694437
rect 46074 693449 46086 694425
rect 46120 693449 46132 694425
rect 46074 693437 46132 693449
rect 46232 694425 46290 694437
rect 46232 693449 46244 694425
rect 46278 693449 46290 694425
rect 46232 693437 46290 693449
rect 46390 694425 46448 694437
rect 46390 693449 46402 694425
rect 46436 693449 46448 694425
rect 46390 693437 46448 693449
rect 46548 694425 46606 694437
rect 46548 693449 46560 694425
rect 46594 693449 46606 694425
rect 46548 693437 46606 693449
rect 46706 694425 46764 694437
rect 46706 693449 46718 694425
rect 46752 693449 46764 694425
rect 46706 693437 46764 693449
rect 46864 694425 46922 694437
rect 46864 693449 46876 694425
rect 46910 693449 46922 694425
rect 46864 693437 46922 693449
rect 47022 694425 47080 694437
rect 47022 693449 47034 694425
rect 47068 693449 47080 694425
rect 47022 693437 47080 693449
rect 47180 694425 47238 694437
rect 47180 693449 47192 694425
rect 47226 693449 47238 694425
rect 47180 693437 47238 693449
rect 47338 694425 47396 694437
rect 47338 693449 47350 694425
rect 47384 693449 47396 694425
rect 47338 693437 47396 693449
rect 47496 694425 47554 694437
rect 47496 693449 47508 694425
rect 47542 693449 47554 694425
rect 47496 693437 47554 693449
rect 47654 694425 47712 694437
rect 47654 693449 47666 694425
rect 47700 693449 47712 694425
rect 47654 693437 47712 693449
rect 47812 694425 47870 694437
rect 47812 693449 47824 694425
rect 47858 693449 47870 694425
rect 47812 693437 47870 693449
rect 47970 694425 48028 694437
rect 47970 693449 47982 694425
rect 48016 693449 48028 694425
rect 47970 693437 48028 693449
rect 48128 694425 48186 694437
rect 48128 693449 48140 694425
rect 48174 693449 48186 694425
rect 48128 693437 48186 693449
rect 48286 694425 48344 694437
rect 48286 693449 48298 694425
rect 48332 693449 48344 694425
rect 48286 693437 48344 693449
rect 48444 694425 48502 694437
rect 48444 693449 48456 694425
rect 48490 693449 48502 694425
rect 48444 693437 48502 693449
rect 48602 694425 48660 694437
rect 48602 693449 48614 694425
rect 48648 693449 48660 694425
rect 48602 693437 48660 693449
rect 43784 692755 43842 692767
rect 43784 691779 43796 692755
rect 43830 691779 43842 692755
rect 43784 691767 43842 691779
rect 43942 692755 44000 692767
rect 43942 691779 43954 692755
rect 43988 691779 44000 692755
rect 43942 691767 44000 691779
rect 44100 692755 44158 692767
rect 44100 691779 44112 692755
rect 44146 691779 44158 692755
rect 44100 691767 44158 691779
rect 44258 692755 44316 692767
rect 44258 691779 44270 692755
rect 44304 691779 44316 692755
rect 44258 691767 44316 691779
rect 44416 692755 44474 692767
rect 44416 691779 44428 692755
rect 44462 691779 44474 692755
rect 44416 691767 44474 691779
rect 44574 692755 44632 692767
rect 44574 691779 44586 692755
rect 44620 691779 44632 692755
rect 44574 691767 44632 691779
rect 44732 692755 44790 692767
rect 44732 691779 44744 692755
rect 44778 691779 44790 692755
rect 44732 691767 44790 691779
rect 44890 692755 44948 692767
rect 44890 691779 44902 692755
rect 44936 691779 44948 692755
rect 44890 691767 44948 691779
rect 45048 692755 45106 692767
rect 45048 691779 45060 692755
rect 45094 691779 45106 692755
rect 45048 691767 45106 691779
rect 45206 692755 45264 692767
rect 45206 691779 45218 692755
rect 45252 691779 45264 692755
rect 45206 691767 45264 691779
rect 45364 692755 45422 692767
rect 45364 691779 45376 692755
rect 45410 691779 45422 692755
rect 45364 691767 45422 691779
rect 45522 692755 45580 692767
rect 45522 691779 45534 692755
rect 45568 691779 45580 692755
rect 45522 691767 45580 691779
rect 45680 692755 45738 692767
rect 45680 691779 45692 692755
rect 45726 691779 45738 692755
rect 45680 691767 45738 691779
rect 45838 692755 45896 692767
rect 45838 691779 45850 692755
rect 45884 691779 45896 692755
rect 45838 691767 45896 691779
rect 45996 692755 46054 692767
rect 45996 691779 46008 692755
rect 46042 691779 46054 692755
rect 45996 691767 46054 691779
rect 46154 692755 46212 692767
rect 46154 691779 46166 692755
rect 46200 691779 46212 692755
rect 46154 691767 46212 691779
rect 46312 692755 46370 692767
rect 46312 691779 46324 692755
rect 46358 691779 46370 692755
rect 46312 691767 46370 691779
rect 46470 692755 46528 692767
rect 46470 691779 46482 692755
rect 46516 691779 46528 692755
rect 46470 691767 46528 691779
rect 46628 692755 46686 692767
rect 46628 691779 46640 692755
rect 46674 691779 46686 692755
rect 46628 691767 46686 691779
rect 46786 692755 46844 692767
rect 46786 691779 46798 692755
rect 46832 691779 46844 692755
rect 46786 691767 46844 691779
rect 46944 692755 47002 692767
rect 46944 691779 46956 692755
rect 46990 691779 47002 692755
rect 46944 691767 47002 691779
rect 47102 692755 47160 692767
rect 47102 691779 47114 692755
rect 47148 691779 47160 692755
rect 47102 691767 47160 691779
rect 43784 691215 43842 691227
rect 43784 690239 43796 691215
rect 43830 690239 43842 691215
rect 43784 690227 43842 690239
rect 43942 691215 44000 691227
rect 43942 690239 43954 691215
rect 43988 690239 44000 691215
rect 43942 690227 44000 690239
rect 44100 691215 44158 691227
rect 44100 690239 44112 691215
rect 44146 690239 44158 691215
rect 44100 690227 44158 690239
rect 44258 691215 44316 691227
rect 44258 690239 44270 691215
rect 44304 690239 44316 691215
rect 44258 690227 44316 690239
rect 44416 691215 44474 691227
rect 44416 690239 44428 691215
rect 44462 690239 44474 691215
rect 44416 690227 44474 690239
rect 44574 691215 44632 691227
rect 44574 690239 44586 691215
rect 44620 690239 44632 691215
rect 44574 690227 44632 690239
rect 44732 691215 44790 691227
rect 44732 690239 44744 691215
rect 44778 690239 44790 691215
rect 44732 690227 44790 690239
rect 44890 691215 44948 691227
rect 44890 690239 44902 691215
rect 44936 690239 44948 691215
rect 44890 690227 44948 690239
rect 45048 691215 45106 691227
rect 45048 690239 45060 691215
rect 45094 690239 45106 691215
rect 45048 690227 45106 690239
rect 45206 691215 45264 691227
rect 45206 690239 45218 691215
rect 45252 690239 45264 691215
rect 45206 690227 45264 690239
rect 45364 691215 45422 691227
rect 45364 690239 45376 691215
rect 45410 690239 45422 691215
rect 45364 690227 45422 690239
rect 45522 691215 45580 691227
rect 45522 690239 45534 691215
rect 45568 690239 45580 691215
rect 45522 690227 45580 690239
rect 45680 691215 45738 691227
rect 45680 690239 45692 691215
rect 45726 690239 45738 691215
rect 45680 690227 45738 690239
rect 45838 691215 45896 691227
rect 45838 690239 45850 691215
rect 45884 690239 45896 691215
rect 45838 690227 45896 690239
rect 45996 691215 46054 691227
rect 45996 690239 46008 691215
rect 46042 690239 46054 691215
rect 45996 690227 46054 690239
rect 46154 691215 46212 691227
rect 46154 690239 46166 691215
rect 46200 690239 46212 691215
rect 46154 690227 46212 690239
rect 46312 691215 46370 691227
rect 46312 690239 46324 691215
rect 46358 690239 46370 691215
rect 46312 690227 46370 690239
rect 46470 691215 46528 691227
rect 46470 690239 46482 691215
rect 46516 690239 46528 691215
rect 46470 690227 46528 690239
rect 46628 691215 46686 691227
rect 46628 690239 46640 691215
rect 46674 690239 46686 691215
rect 46628 690227 46686 690239
rect 46786 691215 46844 691227
rect 46786 690239 46798 691215
rect 46832 690239 46844 691215
rect 46786 690227 46844 690239
rect 46944 691215 47002 691227
rect 46944 690239 46956 691215
rect 46990 690239 47002 691215
rect 46944 690227 47002 690239
rect 47102 691215 47160 691227
rect 47102 690239 47114 691215
rect 47148 690239 47160 691215
rect 47102 690227 47160 690239
rect 41879 682870 42879 682882
rect 41879 682836 41891 682870
rect 42867 682836 42879 682870
rect 41879 682824 42879 682836
rect 43115 682870 44115 682882
rect 43115 682836 43127 682870
rect 44103 682836 44115 682870
rect 43115 682824 44115 682836
rect 44351 682870 45351 682882
rect 44351 682836 44363 682870
rect 45339 682836 45351 682870
rect 44351 682824 45351 682836
rect 45587 682870 46587 682882
rect 45587 682836 45599 682870
rect 46575 682836 46587 682870
rect 45587 682824 46587 682836
rect 46823 682870 47823 682882
rect 46823 682836 46835 682870
rect 47811 682836 47823 682870
rect 46823 682824 47823 682836
rect 48059 682870 49059 682882
rect 48059 682836 48071 682870
rect 49047 682836 49059 682870
rect 48059 682824 49059 682836
rect 41879 682612 42879 682624
rect 41879 682578 41891 682612
rect 42867 682578 42879 682612
rect 41879 682566 42879 682578
rect 43115 682612 44115 682624
rect 43115 682578 43127 682612
rect 44103 682578 44115 682612
rect 43115 682566 44115 682578
rect 44351 682612 45351 682624
rect 44351 682578 44363 682612
rect 45339 682578 45351 682612
rect 44351 682566 45351 682578
rect 45587 682612 46587 682624
rect 45587 682578 45599 682612
rect 46575 682578 46587 682612
rect 45587 682566 46587 682578
rect 46823 682612 47823 682624
rect 46823 682578 46835 682612
rect 47811 682578 47823 682612
rect 46823 682566 47823 682578
rect 48059 682612 49059 682624
rect 48059 682578 48071 682612
rect 49047 682578 49059 682612
rect 48059 682566 49059 682578
rect 41879 682280 42879 682292
rect 41879 682246 41891 682280
rect 42867 682246 42879 682280
rect 41879 682234 42879 682246
rect 43115 682280 44115 682292
rect 43115 682246 43127 682280
rect 44103 682246 44115 682280
rect 43115 682234 44115 682246
rect 44351 682280 45351 682292
rect 44351 682246 44363 682280
rect 45339 682246 45351 682280
rect 44351 682234 45351 682246
rect 45587 682280 46587 682292
rect 45587 682246 45599 682280
rect 46575 682246 46587 682280
rect 45587 682234 46587 682246
rect 46823 682280 47823 682292
rect 46823 682246 46835 682280
rect 47811 682246 47823 682280
rect 46823 682234 47823 682246
rect 48059 682280 49059 682292
rect 48059 682246 48071 682280
rect 49047 682246 49059 682280
rect 48059 682234 49059 682246
rect 41879 682022 42879 682034
rect 41879 681988 41891 682022
rect 42867 681988 42879 682022
rect 41879 681976 42879 681988
rect 43115 682022 44115 682034
rect 43115 681988 43127 682022
rect 44103 681988 44115 682022
rect 43115 681976 44115 681988
rect 44351 682022 45351 682034
rect 44351 681988 44363 682022
rect 45339 681988 45351 682022
rect 44351 681976 45351 681988
rect 45587 682022 46587 682034
rect 45587 681988 45599 682022
rect 46575 681988 46587 682022
rect 45587 681976 46587 681988
rect 46823 682022 47823 682034
rect 46823 681988 46835 682022
rect 47811 681988 47823 682022
rect 46823 681976 47823 681988
rect 48059 682022 49059 682034
rect 48059 681988 48071 682022
rect 49047 681988 49059 682022
rect 48059 681976 49059 681988
<< ndiffc >>
rect 44907 688671 44941 689647
rect 45065 688671 45099 689647
rect 45223 688671 45257 689647
rect 45381 688671 45415 689647
rect 45539 688671 45573 689647
rect 45697 688671 45731 689647
rect 45855 688671 45889 689647
rect 46013 688671 46047 689647
rect 44907 687151 44941 688127
rect 45065 687151 45099 688127
rect 45223 687151 45257 688127
rect 45381 687151 45415 688127
rect 45539 687151 45573 688127
rect 45697 687151 45731 688127
rect 45855 687151 45889 688127
rect 46013 687151 46047 688127
rect 43908 685630 43942 686606
rect 44166 685630 44200 686606
rect 44424 685630 44458 686606
rect 44682 685630 44716 686606
rect 44940 685630 44974 686606
rect 45198 685630 45232 686606
rect 45456 685630 45490 686606
rect 45714 685630 45748 686606
rect 45972 685630 46006 686606
rect 46230 685630 46264 686606
rect 46488 685630 46522 686606
rect 46746 685630 46780 686606
rect 47004 685630 47038 686606
rect 43652 684110 43686 685086
rect 43910 684110 43944 685086
rect 44168 684110 44202 685086
rect 44426 684110 44460 685086
rect 44684 684110 44718 685086
rect 44942 684110 44976 685086
rect 45200 684110 45234 685086
rect 45458 684110 45492 685086
rect 45716 684110 45750 685086
rect 45974 684110 46008 685086
rect 46232 684110 46266 685086
rect 46490 684110 46524 685086
rect 46748 684110 46782 685086
rect 47006 684110 47040 685086
rect 47264 684110 47298 685086
rect 44656 681456 44882 681490
rect 45124 681456 45350 681490
rect 45592 681456 45818 681490
rect 46060 681456 46286 681490
rect 44656 681198 44882 681232
rect 45124 681198 45350 681232
rect 45592 681198 45818 681232
rect 46060 681198 46286 681232
rect 44872 680831 45348 680865
rect 45590 680831 46066 680865
rect 44872 680673 45348 680707
rect 45590 680673 46066 680707
rect 41935 680306 42911 680340
rect 43153 680306 44129 680340
rect 44371 680306 45347 680340
rect 45589 680306 46565 680340
rect 46807 680306 47783 680340
rect 48025 680306 49001 680340
rect 41935 680048 42911 680082
rect 43153 680048 44129 680082
rect 44371 680048 45347 680082
rect 45589 680048 46565 680082
rect 46807 680048 47783 680082
rect 48025 680048 49001 680082
<< pdiffc >>
rect 42294 693449 42328 694425
rect 42452 693449 42486 694425
rect 42610 693449 42644 694425
rect 42768 693449 42802 694425
rect 42926 693449 42960 694425
rect 43084 693449 43118 694425
rect 43242 693449 43276 694425
rect 43400 693449 43434 694425
rect 43558 693449 43592 694425
rect 43716 693449 43750 694425
rect 43874 693449 43908 694425
rect 44032 693449 44066 694425
rect 44190 693449 44224 694425
rect 44348 693449 44382 694425
rect 44506 693449 44540 694425
rect 44664 693449 44698 694425
rect 44822 693449 44856 694425
rect 44980 693449 45014 694425
rect 45138 693449 45172 694425
rect 45296 693449 45330 694425
rect 45454 693449 45488 694425
rect 45612 693449 45646 694425
rect 45770 693449 45804 694425
rect 45928 693449 45962 694425
rect 46086 693449 46120 694425
rect 46244 693449 46278 694425
rect 46402 693449 46436 694425
rect 46560 693449 46594 694425
rect 46718 693449 46752 694425
rect 46876 693449 46910 694425
rect 47034 693449 47068 694425
rect 47192 693449 47226 694425
rect 47350 693449 47384 694425
rect 47508 693449 47542 694425
rect 47666 693449 47700 694425
rect 47824 693449 47858 694425
rect 47982 693449 48016 694425
rect 48140 693449 48174 694425
rect 48298 693449 48332 694425
rect 48456 693449 48490 694425
rect 48614 693449 48648 694425
rect 43796 691779 43830 692755
rect 43954 691779 43988 692755
rect 44112 691779 44146 692755
rect 44270 691779 44304 692755
rect 44428 691779 44462 692755
rect 44586 691779 44620 692755
rect 44744 691779 44778 692755
rect 44902 691779 44936 692755
rect 45060 691779 45094 692755
rect 45218 691779 45252 692755
rect 45376 691779 45410 692755
rect 45534 691779 45568 692755
rect 45692 691779 45726 692755
rect 45850 691779 45884 692755
rect 46008 691779 46042 692755
rect 46166 691779 46200 692755
rect 46324 691779 46358 692755
rect 46482 691779 46516 692755
rect 46640 691779 46674 692755
rect 46798 691779 46832 692755
rect 46956 691779 46990 692755
rect 47114 691779 47148 692755
rect 43796 690239 43830 691215
rect 43954 690239 43988 691215
rect 44112 690239 44146 691215
rect 44270 690239 44304 691215
rect 44428 690239 44462 691215
rect 44586 690239 44620 691215
rect 44744 690239 44778 691215
rect 44902 690239 44936 691215
rect 45060 690239 45094 691215
rect 45218 690239 45252 691215
rect 45376 690239 45410 691215
rect 45534 690239 45568 691215
rect 45692 690239 45726 691215
rect 45850 690239 45884 691215
rect 46008 690239 46042 691215
rect 46166 690239 46200 691215
rect 46324 690239 46358 691215
rect 46482 690239 46516 691215
rect 46640 690239 46674 691215
rect 46798 690239 46832 691215
rect 46956 690239 46990 691215
rect 47114 690239 47148 691215
rect 41891 682836 42867 682870
rect 43127 682836 44103 682870
rect 44363 682836 45339 682870
rect 45599 682836 46575 682870
rect 46835 682836 47811 682870
rect 48071 682836 49047 682870
rect 41891 682578 42867 682612
rect 43127 682578 44103 682612
rect 44363 682578 45339 682612
rect 45599 682578 46575 682612
rect 46835 682578 47811 682612
rect 48071 682578 49047 682612
rect 41891 682246 42867 682280
rect 43127 682246 44103 682280
rect 44363 682246 45339 682280
rect 45599 682246 46575 682280
rect 46835 682246 47811 682280
rect 48071 682246 49047 682280
rect 41891 681988 42867 682022
rect 43127 681988 44103 682022
rect 44363 681988 45339 682022
rect 45599 681988 46575 682022
rect 46835 681988 47811 682022
rect 48071 681988 49047 682022
<< psubdiff >>
rect 38371 695463 38467 695497
rect 41399 695463 41495 695497
rect 38371 695401 38405 695463
rect 41461 695401 41495 695463
rect 38371 694125 38405 694187
rect 49441 695463 49537 695497
rect 52469 695463 52565 695497
rect 49441 695401 49475 695463
rect 41461 694125 41495 694187
rect 38371 694091 38467 694125
rect 41399 694091 41495 694125
rect 38371 694003 38467 694037
rect 41399 694003 41495 694037
rect 38371 693941 38405 694003
rect 41461 693941 41495 694003
rect 38371 692665 38405 692727
rect 52531 695401 52565 695463
rect 49441 694125 49475 694187
rect 52531 694125 52565 694187
rect 49441 694091 49537 694125
rect 52469 694091 52565 694125
rect 49441 694003 49537 694037
rect 52469 694003 52565 694037
rect 49441 693941 49475 694003
rect 41461 692665 41495 692727
rect 38371 692631 38467 692665
rect 41399 692631 41495 692665
rect 52531 693941 52565 694003
rect 49441 692665 49475 692727
rect 52531 692665 52565 692727
rect 49441 692631 49537 692665
rect 52469 692631 52565 692665
rect 44793 689799 44889 689833
rect 46065 689799 46161 689833
rect 44793 689737 44827 689799
rect 46127 689737 46161 689799
rect 44793 688519 44827 688581
rect 46127 688519 46161 688581
rect 44793 688485 44889 688519
rect 46065 688485 46161 688519
rect 44793 688279 44889 688313
rect 46065 688279 46161 688313
rect 44793 688217 44827 688279
rect 46127 688217 46161 688279
rect 44793 686999 44827 687061
rect 46127 686999 46161 687061
rect 44793 686965 44889 686999
rect 46065 686965 46161 686999
rect 43794 686758 43890 686792
rect 47056 686758 47152 686792
rect 43794 686696 43828 686758
rect 47118 686696 47152 686758
rect 43794 685478 43828 685540
rect 47118 685478 47152 685540
rect 43794 685444 43890 685478
rect 47056 685444 47152 685478
rect 43538 685238 43634 685272
rect 47316 685238 47412 685272
rect 43538 685176 43572 685238
rect 47378 685176 47412 685238
rect 43538 683958 43572 684020
rect 47378 683958 47412 684020
rect 43538 683924 43634 683958
rect 47316 683924 47412 683958
rect 44470 681570 44566 681604
rect 46376 681570 46472 681604
rect 44470 681508 44504 681570
rect 46438 681508 46472 681570
rect 44470 681118 44504 681180
rect 46438 681118 46472 681180
rect 44470 681084 44566 681118
rect 46376 681084 46472 681118
rect 44686 680945 44782 680979
rect 46156 680945 46252 680979
rect 44686 680883 44720 680945
rect 46218 680883 46252 680945
rect 44686 680593 44720 680655
rect 46218 680593 46252 680655
rect 44686 680559 44782 680593
rect 46156 680559 46252 680593
rect 41749 680420 41845 680454
rect 49091 680420 49187 680454
rect 41749 680358 41783 680420
rect 49153 680358 49187 680420
rect 41749 679968 41783 680030
rect 49153 679968 49187 680030
rect 41749 679934 41845 679968
rect 49091 679934 49187 679968
rect 42218 678658 42338 678682
rect 42218 678514 42338 678538
rect 42218 675658 42338 675682
rect 42218 675514 42338 675538
rect 42218 672658 42338 672682
rect 42218 672514 42338 672538
rect 42218 669658 42338 669682
rect 42218 669514 42338 669538
rect 42218 666658 42338 666682
rect 42218 666514 42338 666538
rect 48588 678658 48708 678682
rect 48588 678514 48708 678538
rect 48588 675658 48708 675682
rect 48588 675514 48708 675538
rect 48588 672658 48708 672682
rect 48588 672514 48708 672538
rect 48588 669658 48708 669682
rect 48588 669514 48708 669538
rect 48588 666658 48708 666682
rect 48588 666514 48708 666538
<< nsubdiff >>
rect 42180 694586 42276 694620
rect 48666 694586 48762 694620
rect 42180 694524 42214 694586
rect 48728 694524 48762 694586
rect 42180 693288 42214 693350
rect 48728 693288 48762 693350
rect 42180 693254 42276 693288
rect 48666 693254 48762 693288
rect 43682 692916 43778 692950
rect 47166 692916 47262 692950
rect 43682 692854 43716 692916
rect 47228 692854 47262 692916
rect 43682 691618 43716 691680
rect 47228 691618 47262 691680
rect 43682 691584 43778 691618
rect 47166 691584 47262 691618
rect 43682 691376 43778 691410
rect 47166 691376 47262 691410
rect 43682 691314 43716 691376
rect 47228 691314 47262 691376
rect 43682 690078 43716 690140
rect 47228 690078 47262 690140
rect 43682 690044 43778 690078
rect 47166 690044 47262 690078
rect 41696 682950 41792 682984
rect 49146 682950 49242 682984
rect 41696 682888 41730 682950
rect 49208 682888 49242 682950
rect 41696 682498 41730 682560
rect 49208 682498 49242 682560
rect 41696 682464 41792 682498
rect 49146 682464 49242 682498
rect 41696 682360 41792 682394
rect 49146 682360 49242 682394
rect 41696 682298 41730 682360
rect 49208 682298 49242 682360
rect 41696 681908 41730 681970
rect 49208 681908 49242 681970
rect 41696 681874 41792 681908
rect 49146 681874 49242 681908
<< psubdiffcont >>
rect 38467 695463 41399 695497
rect 38371 694187 38405 695401
rect 41461 694187 41495 695401
rect 49537 695463 52469 695497
rect 38467 694091 41399 694125
rect 38467 694003 41399 694037
rect 38371 692727 38405 693941
rect 41461 692727 41495 693941
rect 49441 694187 49475 695401
rect 52531 694187 52565 695401
rect 49537 694091 52469 694125
rect 49537 694003 52469 694037
rect 38467 692631 41399 692665
rect 49441 692727 49475 693941
rect 52531 692727 52565 693941
rect 49537 692631 52469 692665
rect 44889 689799 46065 689833
rect 44793 688581 44827 689737
rect 46127 688581 46161 689737
rect 44889 688485 46065 688519
rect 44889 688279 46065 688313
rect 44793 687061 44827 688217
rect 46127 687061 46161 688217
rect 44889 686965 46065 686999
rect 43890 686758 47056 686792
rect 43794 685540 43828 686696
rect 47118 685540 47152 686696
rect 43890 685444 47056 685478
rect 43634 685238 47316 685272
rect 43538 684020 43572 685176
rect 47378 684020 47412 685176
rect 43634 683924 47316 683958
rect 44566 681570 46376 681604
rect 44470 681180 44504 681508
rect 46438 681180 46472 681508
rect 44566 681084 46376 681118
rect 44782 680945 46156 680979
rect 44686 680655 44720 680883
rect 46218 680655 46252 680883
rect 44782 680559 46156 680593
rect 41845 680420 49091 680454
rect 41749 680030 41783 680358
rect 49153 680030 49187 680358
rect 41845 679934 49091 679968
rect 42218 678538 42338 678658
rect 42218 675538 42338 675658
rect 42218 672538 42338 672658
rect 42218 669538 42338 669658
rect 42218 666538 42338 666658
rect 48588 678538 48708 678658
rect 48588 675538 48708 675658
rect 48588 672538 48708 672658
rect 48588 669538 48708 669658
rect 48588 666538 48708 666658
<< nsubdiffcont >>
rect 42276 694586 48666 694620
rect 42180 693350 42214 694524
rect 48728 693350 48762 694524
rect 42276 693254 48666 693288
rect 43778 692916 47166 692950
rect 43682 691680 43716 692854
rect 47228 691680 47262 692854
rect 43778 691584 47166 691618
rect 43778 691376 47166 691410
rect 43682 690140 43716 691314
rect 47228 690140 47262 691314
rect 43778 690044 47166 690078
rect 41792 682950 49146 682984
rect 41696 682560 41730 682888
rect 49208 682560 49242 682888
rect 41792 682464 49146 682498
rect 41792 682360 49146 682394
rect 41696 681970 41730 682298
rect 49208 681970 49242 682298
rect 41792 681874 49146 681908
<< poly >>
rect 42340 694518 42440 694534
rect 42340 694484 42356 694518
rect 42424 694484 42440 694518
rect 42340 694437 42440 694484
rect 42498 694518 42598 694534
rect 42498 694484 42514 694518
rect 42582 694484 42598 694518
rect 42498 694437 42598 694484
rect 42656 694518 42756 694534
rect 42656 694484 42672 694518
rect 42740 694484 42756 694518
rect 42656 694437 42756 694484
rect 42814 694518 42914 694534
rect 42814 694484 42830 694518
rect 42898 694484 42914 694518
rect 42814 694437 42914 694484
rect 42972 694518 43072 694534
rect 42972 694484 42988 694518
rect 43056 694484 43072 694518
rect 42972 694437 43072 694484
rect 43130 694518 43230 694534
rect 43130 694484 43146 694518
rect 43214 694484 43230 694518
rect 43130 694437 43230 694484
rect 43288 694518 43388 694534
rect 43288 694484 43304 694518
rect 43372 694484 43388 694518
rect 43288 694437 43388 694484
rect 43446 694518 43546 694534
rect 43446 694484 43462 694518
rect 43530 694484 43546 694518
rect 43446 694437 43546 694484
rect 43604 694518 43704 694534
rect 43604 694484 43620 694518
rect 43688 694484 43704 694518
rect 43604 694437 43704 694484
rect 43762 694518 43862 694534
rect 43762 694484 43778 694518
rect 43846 694484 43862 694518
rect 43762 694437 43862 694484
rect 43920 694518 44020 694534
rect 43920 694484 43936 694518
rect 44004 694484 44020 694518
rect 43920 694437 44020 694484
rect 44078 694518 44178 694534
rect 44078 694484 44094 694518
rect 44162 694484 44178 694518
rect 44078 694437 44178 694484
rect 44236 694518 44336 694534
rect 44236 694484 44252 694518
rect 44320 694484 44336 694518
rect 44236 694437 44336 694484
rect 44394 694518 44494 694534
rect 44394 694484 44410 694518
rect 44478 694484 44494 694518
rect 44394 694437 44494 694484
rect 44552 694518 44652 694534
rect 44552 694484 44568 694518
rect 44636 694484 44652 694518
rect 44552 694437 44652 694484
rect 44710 694518 44810 694534
rect 44710 694484 44726 694518
rect 44794 694484 44810 694518
rect 44710 694437 44810 694484
rect 44868 694518 44968 694534
rect 44868 694484 44884 694518
rect 44952 694484 44968 694518
rect 44868 694437 44968 694484
rect 45026 694518 45126 694534
rect 45026 694484 45042 694518
rect 45110 694484 45126 694518
rect 45026 694437 45126 694484
rect 45184 694518 45284 694534
rect 45184 694484 45200 694518
rect 45268 694484 45284 694518
rect 45184 694437 45284 694484
rect 45342 694518 45442 694534
rect 45342 694484 45358 694518
rect 45426 694484 45442 694518
rect 45342 694437 45442 694484
rect 45500 694518 45600 694534
rect 45500 694484 45516 694518
rect 45584 694484 45600 694518
rect 45500 694437 45600 694484
rect 45658 694518 45758 694534
rect 45658 694484 45674 694518
rect 45742 694484 45758 694518
rect 45658 694437 45758 694484
rect 45816 694518 45916 694534
rect 45816 694484 45832 694518
rect 45900 694484 45916 694518
rect 45816 694437 45916 694484
rect 45974 694518 46074 694534
rect 45974 694484 45990 694518
rect 46058 694484 46074 694518
rect 45974 694437 46074 694484
rect 46132 694518 46232 694534
rect 46132 694484 46148 694518
rect 46216 694484 46232 694518
rect 46132 694437 46232 694484
rect 46290 694518 46390 694534
rect 46290 694484 46306 694518
rect 46374 694484 46390 694518
rect 46290 694437 46390 694484
rect 46448 694518 46548 694534
rect 46448 694484 46464 694518
rect 46532 694484 46548 694518
rect 46448 694437 46548 694484
rect 46606 694518 46706 694534
rect 46606 694484 46622 694518
rect 46690 694484 46706 694518
rect 46606 694437 46706 694484
rect 46764 694518 46864 694534
rect 46764 694484 46780 694518
rect 46848 694484 46864 694518
rect 46764 694437 46864 694484
rect 46922 694518 47022 694534
rect 46922 694484 46938 694518
rect 47006 694484 47022 694518
rect 46922 694437 47022 694484
rect 47080 694518 47180 694534
rect 47080 694484 47096 694518
rect 47164 694484 47180 694518
rect 47080 694437 47180 694484
rect 47238 694518 47338 694534
rect 47238 694484 47254 694518
rect 47322 694484 47338 694518
rect 47238 694437 47338 694484
rect 47396 694518 47496 694534
rect 47396 694484 47412 694518
rect 47480 694484 47496 694518
rect 47396 694437 47496 694484
rect 47554 694518 47654 694534
rect 47554 694484 47570 694518
rect 47638 694484 47654 694518
rect 47554 694437 47654 694484
rect 47712 694518 47812 694534
rect 47712 694484 47728 694518
rect 47796 694484 47812 694518
rect 47712 694437 47812 694484
rect 47870 694518 47970 694534
rect 47870 694484 47886 694518
rect 47954 694484 47970 694518
rect 47870 694437 47970 694484
rect 48028 694518 48128 694534
rect 48028 694484 48044 694518
rect 48112 694484 48128 694518
rect 48028 694437 48128 694484
rect 48186 694518 48286 694534
rect 48186 694484 48202 694518
rect 48270 694484 48286 694518
rect 48186 694437 48286 694484
rect 48344 694518 48444 694534
rect 48344 694484 48360 694518
rect 48428 694484 48444 694518
rect 48344 694437 48444 694484
rect 48502 694518 48602 694534
rect 48502 694484 48518 694518
rect 48586 694484 48602 694518
rect 48502 694437 48602 694484
rect 42340 693390 42440 693437
rect 42340 693356 42356 693390
rect 42424 693356 42440 693390
rect 42340 693340 42440 693356
rect 42498 693390 42598 693437
rect 42498 693356 42514 693390
rect 42582 693356 42598 693390
rect 42498 693340 42598 693356
rect 42656 693390 42756 693437
rect 42656 693356 42672 693390
rect 42740 693356 42756 693390
rect 42656 693340 42756 693356
rect 42814 693390 42914 693437
rect 42814 693356 42830 693390
rect 42898 693356 42914 693390
rect 42814 693340 42914 693356
rect 42972 693390 43072 693437
rect 42972 693356 42988 693390
rect 43056 693356 43072 693390
rect 42972 693340 43072 693356
rect 43130 693390 43230 693437
rect 43130 693356 43146 693390
rect 43214 693356 43230 693390
rect 43130 693340 43230 693356
rect 43288 693390 43388 693437
rect 43288 693356 43304 693390
rect 43372 693356 43388 693390
rect 43288 693340 43388 693356
rect 43446 693390 43546 693437
rect 43446 693356 43462 693390
rect 43530 693356 43546 693390
rect 43446 693340 43546 693356
rect 43604 693390 43704 693437
rect 43604 693356 43620 693390
rect 43688 693356 43704 693390
rect 43604 693340 43704 693356
rect 43762 693390 43862 693437
rect 43762 693356 43778 693390
rect 43846 693356 43862 693390
rect 43762 693340 43862 693356
rect 43920 693390 44020 693437
rect 43920 693356 43936 693390
rect 44004 693356 44020 693390
rect 43920 693340 44020 693356
rect 44078 693390 44178 693437
rect 44078 693356 44094 693390
rect 44162 693356 44178 693390
rect 44078 693340 44178 693356
rect 44236 693390 44336 693437
rect 44236 693356 44252 693390
rect 44320 693356 44336 693390
rect 44236 693340 44336 693356
rect 44394 693390 44494 693437
rect 44394 693356 44410 693390
rect 44478 693356 44494 693390
rect 44394 693340 44494 693356
rect 44552 693390 44652 693437
rect 44552 693356 44568 693390
rect 44636 693356 44652 693390
rect 44552 693340 44652 693356
rect 44710 693390 44810 693437
rect 44710 693356 44726 693390
rect 44794 693356 44810 693390
rect 44710 693340 44810 693356
rect 44868 693390 44968 693437
rect 44868 693356 44884 693390
rect 44952 693356 44968 693390
rect 44868 693340 44968 693356
rect 45026 693390 45126 693437
rect 45026 693356 45042 693390
rect 45110 693356 45126 693390
rect 45026 693340 45126 693356
rect 45184 693390 45284 693437
rect 45184 693356 45200 693390
rect 45268 693356 45284 693390
rect 45184 693340 45284 693356
rect 45342 693390 45442 693437
rect 45342 693356 45358 693390
rect 45426 693356 45442 693390
rect 45342 693340 45442 693356
rect 45500 693390 45600 693437
rect 45500 693356 45516 693390
rect 45584 693356 45600 693390
rect 45500 693340 45600 693356
rect 45658 693390 45758 693437
rect 45658 693356 45674 693390
rect 45742 693356 45758 693390
rect 45658 693340 45758 693356
rect 45816 693390 45916 693437
rect 45816 693356 45832 693390
rect 45900 693356 45916 693390
rect 45816 693340 45916 693356
rect 45974 693390 46074 693437
rect 45974 693356 45990 693390
rect 46058 693356 46074 693390
rect 45974 693340 46074 693356
rect 46132 693390 46232 693437
rect 46132 693356 46148 693390
rect 46216 693356 46232 693390
rect 46132 693340 46232 693356
rect 46290 693390 46390 693437
rect 46290 693356 46306 693390
rect 46374 693356 46390 693390
rect 46290 693340 46390 693356
rect 46448 693390 46548 693437
rect 46448 693356 46464 693390
rect 46532 693356 46548 693390
rect 46448 693340 46548 693356
rect 46606 693390 46706 693437
rect 46606 693356 46622 693390
rect 46690 693356 46706 693390
rect 46606 693340 46706 693356
rect 46764 693390 46864 693437
rect 46764 693356 46780 693390
rect 46848 693356 46864 693390
rect 46764 693340 46864 693356
rect 46922 693390 47022 693437
rect 46922 693356 46938 693390
rect 47006 693356 47022 693390
rect 46922 693340 47022 693356
rect 47080 693390 47180 693437
rect 47080 693356 47096 693390
rect 47164 693356 47180 693390
rect 47080 693340 47180 693356
rect 47238 693390 47338 693437
rect 47238 693356 47254 693390
rect 47322 693356 47338 693390
rect 47238 693340 47338 693356
rect 47396 693390 47496 693437
rect 47396 693356 47412 693390
rect 47480 693356 47496 693390
rect 47396 693340 47496 693356
rect 47554 693390 47654 693437
rect 47554 693356 47570 693390
rect 47638 693356 47654 693390
rect 47554 693340 47654 693356
rect 47712 693390 47812 693437
rect 47712 693356 47728 693390
rect 47796 693356 47812 693390
rect 47712 693340 47812 693356
rect 47870 693390 47970 693437
rect 47870 693356 47886 693390
rect 47954 693356 47970 693390
rect 47870 693340 47970 693356
rect 48028 693390 48128 693437
rect 48028 693356 48044 693390
rect 48112 693356 48128 693390
rect 48028 693340 48128 693356
rect 48186 693390 48286 693437
rect 48186 693356 48202 693390
rect 48270 693356 48286 693390
rect 48186 693340 48286 693356
rect 48344 693390 48444 693437
rect 48344 693356 48360 693390
rect 48428 693356 48444 693390
rect 48344 693340 48444 693356
rect 48502 693390 48602 693437
rect 48502 693356 48518 693390
rect 48586 693356 48602 693390
rect 48502 693340 48602 693356
rect 43842 692848 43942 692864
rect 43842 692814 43858 692848
rect 43926 692814 43942 692848
rect 43842 692767 43942 692814
rect 44000 692848 44100 692864
rect 44000 692814 44016 692848
rect 44084 692814 44100 692848
rect 44000 692767 44100 692814
rect 44158 692848 44258 692864
rect 44158 692814 44174 692848
rect 44242 692814 44258 692848
rect 44158 692767 44258 692814
rect 44316 692848 44416 692864
rect 44316 692814 44332 692848
rect 44400 692814 44416 692848
rect 44316 692767 44416 692814
rect 44474 692848 44574 692864
rect 44474 692814 44490 692848
rect 44558 692814 44574 692848
rect 44474 692767 44574 692814
rect 44632 692848 44732 692864
rect 44632 692814 44648 692848
rect 44716 692814 44732 692848
rect 44632 692767 44732 692814
rect 44790 692848 44890 692864
rect 44790 692814 44806 692848
rect 44874 692814 44890 692848
rect 44790 692767 44890 692814
rect 44948 692848 45048 692864
rect 44948 692814 44964 692848
rect 45032 692814 45048 692848
rect 44948 692767 45048 692814
rect 45106 692848 45206 692864
rect 45106 692814 45122 692848
rect 45190 692814 45206 692848
rect 45106 692767 45206 692814
rect 45264 692848 45364 692864
rect 45264 692814 45280 692848
rect 45348 692814 45364 692848
rect 45264 692767 45364 692814
rect 45422 692848 45522 692864
rect 45422 692814 45438 692848
rect 45506 692814 45522 692848
rect 45422 692767 45522 692814
rect 45580 692848 45680 692864
rect 45580 692814 45596 692848
rect 45664 692814 45680 692848
rect 45580 692767 45680 692814
rect 45738 692848 45838 692864
rect 45738 692814 45754 692848
rect 45822 692814 45838 692848
rect 45738 692767 45838 692814
rect 45896 692848 45996 692864
rect 45896 692814 45912 692848
rect 45980 692814 45996 692848
rect 45896 692767 45996 692814
rect 46054 692848 46154 692864
rect 46054 692814 46070 692848
rect 46138 692814 46154 692848
rect 46054 692767 46154 692814
rect 46212 692848 46312 692864
rect 46212 692814 46228 692848
rect 46296 692814 46312 692848
rect 46212 692767 46312 692814
rect 46370 692848 46470 692864
rect 46370 692814 46386 692848
rect 46454 692814 46470 692848
rect 46370 692767 46470 692814
rect 46528 692848 46628 692864
rect 46528 692814 46544 692848
rect 46612 692814 46628 692848
rect 46528 692767 46628 692814
rect 46686 692848 46786 692864
rect 46686 692814 46702 692848
rect 46770 692814 46786 692848
rect 46686 692767 46786 692814
rect 46844 692848 46944 692864
rect 46844 692814 46860 692848
rect 46928 692814 46944 692848
rect 46844 692767 46944 692814
rect 47002 692848 47102 692864
rect 47002 692814 47018 692848
rect 47086 692814 47102 692848
rect 47002 692767 47102 692814
rect 43842 691720 43942 691767
rect 43842 691686 43858 691720
rect 43926 691686 43942 691720
rect 43842 691670 43942 691686
rect 44000 691720 44100 691767
rect 44000 691686 44016 691720
rect 44084 691686 44100 691720
rect 44000 691670 44100 691686
rect 44158 691720 44258 691767
rect 44158 691686 44174 691720
rect 44242 691686 44258 691720
rect 44158 691670 44258 691686
rect 44316 691720 44416 691767
rect 44316 691686 44332 691720
rect 44400 691686 44416 691720
rect 44316 691670 44416 691686
rect 44474 691720 44574 691767
rect 44474 691686 44490 691720
rect 44558 691686 44574 691720
rect 44474 691670 44574 691686
rect 44632 691720 44732 691767
rect 44632 691686 44648 691720
rect 44716 691686 44732 691720
rect 44632 691670 44732 691686
rect 44790 691720 44890 691767
rect 44790 691686 44806 691720
rect 44874 691686 44890 691720
rect 44790 691670 44890 691686
rect 44948 691720 45048 691767
rect 44948 691686 44964 691720
rect 45032 691686 45048 691720
rect 44948 691670 45048 691686
rect 45106 691720 45206 691767
rect 45106 691686 45122 691720
rect 45190 691686 45206 691720
rect 45106 691670 45206 691686
rect 45264 691720 45364 691767
rect 45264 691686 45280 691720
rect 45348 691686 45364 691720
rect 45264 691670 45364 691686
rect 45422 691720 45522 691767
rect 45422 691686 45438 691720
rect 45506 691686 45522 691720
rect 45422 691670 45522 691686
rect 45580 691720 45680 691767
rect 45580 691686 45596 691720
rect 45664 691686 45680 691720
rect 45580 691670 45680 691686
rect 45738 691720 45838 691767
rect 45738 691686 45754 691720
rect 45822 691686 45838 691720
rect 45738 691670 45838 691686
rect 45896 691720 45996 691767
rect 45896 691686 45912 691720
rect 45980 691686 45996 691720
rect 45896 691670 45996 691686
rect 46054 691720 46154 691767
rect 46054 691686 46070 691720
rect 46138 691686 46154 691720
rect 46054 691670 46154 691686
rect 46212 691720 46312 691767
rect 46212 691686 46228 691720
rect 46296 691686 46312 691720
rect 46212 691670 46312 691686
rect 46370 691720 46470 691767
rect 46370 691686 46386 691720
rect 46454 691686 46470 691720
rect 46370 691670 46470 691686
rect 46528 691720 46628 691767
rect 46528 691686 46544 691720
rect 46612 691686 46628 691720
rect 46528 691670 46628 691686
rect 46686 691720 46786 691767
rect 46686 691686 46702 691720
rect 46770 691686 46786 691720
rect 46686 691670 46786 691686
rect 46844 691720 46944 691767
rect 46844 691686 46860 691720
rect 46928 691686 46944 691720
rect 46844 691670 46944 691686
rect 47002 691720 47102 691767
rect 47002 691686 47018 691720
rect 47086 691686 47102 691720
rect 47002 691670 47102 691686
rect 43842 691308 43942 691324
rect 43842 691274 43858 691308
rect 43926 691274 43942 691308
rect 43842 691227 43942 691274
rect 44000 691308 44100 691324
rect 44000 691274 44016 691308
rect 44084 691274 44100 691308
rect 44000 691227 44100 691274
rect 44158 691308 44258 691324
rect 44158 691274 44174 691308
rect 44242 691274 44258 691308
rect 44158 691227 44258 691274
rect 44316 691308 44416 691324
rect 44316 691274 44332 691308
rect 44400 691274 44416 691308
rect 44316 691227 44416 691274
rect 44474 691308 44574 691324
rect 44474 691274 44490 691308
rect 44558 691274 44574 691308
rect 44474 691227 44574 691274
rect 44632 691308 44732 691324
rect 44632 691274 44648 691308
rect 44716 691274 44732 691308
rect 44632 691227 44732 691274
rect 44790 691308 44890 691324
rect 44790 691274 44806 691308
rect 44874 691274 44890 691308
rect 44790 691227 44890 691274
rect 44948 691308 45048 691324
rect 44948 691274 44964 691308
rect 45032 691274 45048 691308
rect 44948 691227 45048 691274
rect 45106 691308 45206 691324
rect 45106 691274 45122 691308
rect 45190 691274 45206 691308
rect 45106 691227 45206 691274
rect 45264 691308 45364 691324
rect 45264 691274 45280 691308
rect 45348 691274 45364 691308
rect 45264 691227 45364 691274
rect 45422 691308 45522 691324
rect 45422 691274 45438 691308
rect 45506 691274 45522 691308
rect 45422 691227 45522 691274
rect 45580 691308 45680 691324
rect 45580 691274 45596 691308
rect 45664 691274 45680 691308
rect 45580 691227 45680 691274
rect 45738 691308 45838 691324
rect 45738 691274 45754 691308
rect 45822 691274 45838 691308
rect 45738 691227 45838 691274
rect 45896 691308 45996 691324
rect 45896 691274 45912 691308
rect 45980 691274 45996 691308
rect 45896 691227 45996 691274
rect 46054 691308 46154 691324
rect 46054 691274 46070 691308
rect 46138 691274 46154 691308
rect 46054 691227 46154 691274
rect 46212 691308 46312 691324
rect 46212 691274 46228 691308
rect 46296 691274 46312 691308
rect 46212 691227 46312 691274
rect 46370 691308 46470 691324
rect 46370 691274 46386 691308
rect 46454 691274 46470 691308
rect 46370 691227 46470 691274
rect 46528 691308 46628 691324
rect 46528 691274 46544 691308
rect 46612 691274 46628 691308
rect 46528 691227 46628 691274
rect 46686 691308 46786 691324
rect 46686 691274 46702 691308
rect 46770 691274 46786 691308
rect 46686 691227 46786 691274
rect 46844 691308 46944 691324
rect 46844 691274 46860 691308
rect 46928 691274 46944 691308
rect 46844 691227 46944 691274
rect 47002 691308 47102 691324
rect 47002 691274 47018 691308
rect 47086 691274 47102 691308
rect 47002 691227 47102 691274
rect 43842 690180 43942 690227
rect 43842 690146 43858 690180
rect 43926 690146 43942 690180
rect 43842 690130 43942 690146
rect 44000 690180 44100 690227
rect 44000 690146 44016 690180
rect 44084 690146 44100 690180
rect 44000 690130 44100 690146
rect 44158 690180 44258 690227
rect 44158 690146 44174 690180
rect 44242 690146 44258 690180
rect 44158 690130 44258 690146
rect 44316 690180 44416 690227
rect 44316 690146 44332 690180
rect 44400 690146 44416 690180
rect 44316 690130 44416 690146
rect 44474 690180 44574 690227
rect 44474 690146 44490 690180
rect 44558 690146 44574 690180
rect 44474 690130 44574 690146
rect 44632 690180 44732 690227
rect 44632 690146 44648 690180
rect 44716 690146 44732 690180
rect 44632 690130 44732 690146
rect 44790 690180 44890 690227
rect 44790 690146 44806 690180
rect 44874 690146 44890 690180
rect 44790 690130 44890 690146
rect 44948 690180 45048 690227
rect 44948 690146 44964 690180
rect 45032 690146 45048 690180
rect 44948 690130 45048 690146
rect 45106 690180 45206 690227
rect 45106 690146 45122 690180
rect 45190 690146 45206 690180
rect 45106 690130 45206 690146
rect 45264 690180 45364 690227
rect 45264 690146 45280 690180
rect 45348 690146 45364 690180
rect 45264 690130 45364 690146
rect 45422 690180 45522 690227
rect 45422 690146 45438 690180
rect 45506 690146 45522 690180
rect 45422 690130 45522 690146
rect 45580 690180 45680 690227
rect 45580 690146 45596 690180
rect 45664 690146 45680 690180
rect 45580 690130 45680 690146
rect 45738 690180 45838 690227
rect 45738 690146 45754 690180
rect 45822 690146 45838 690180
rect 45738 690130 45838 690146
rect 45896 690180 45996 690227
rect 45896 690146 45912 690180
rect 45980 690146 45996 690180
rect 45896 690130 45996 690146
rect 46054 690180 46154 690227
rect 46054 690146 46070 690180
rect 46138 690146 46154 690180
rect 46054 690130 46154 690146
rect 46212 690180 46312 690227
rect 46212 690146 46228 690180
rect 46296 690146 46312 690180
rect 46212 690130 46312 690146
rect 46370 690180 46470 690227
rect 46370 690146 46386 690180
rect 46454 690146 46470 690180
rect 46370 690130 46470 690146
rect 46528 690180 46628 690227
rect 46528 690146 46544 690180
rect 46612 690146 46628 690180
rect 46528 690130 46628 690146
rect 46686 690180 46786 690227
rect 46686 690146 46702 690180
rect 46770 690146 46786 690180
rect 46686 690130 46786 690146
rect 46844 690180 46944 690227
rect 46844 690146 46860 690180
rect 46928 690146 46944 690180
rect 46844 690130 46944 690146
rect 47002 690180 47102 690227
rect 47002 690146 47018 690180
rect 47086 690146 47102 690180
rect 47002 690130 47102 690146
rect 44953 689731 45053 689747
rect 44953 689697 44969 689731
rect 45037 689697 45053 689731
rect 44953 689659 45053 689697
rect 45111 689731 45211 689747
rect 45111 689697 45127 689731
rect 45195 689697 45211 689731
rect 45111 689659 45211 689697
rect 45269 689731 45369 689747
rect 45269 689697 45285 689731
rect 45353 689697 45369 689731
rect 45269 689659 45369 689697
rect 45427 689731 45527 689747
rect 45427 689697 45443 689731
rect 45511 689697 45527 689731
rect 45427 689659 45527 689697
rect 45585 689731 45685 689747
rect 45585 689697 45601 689731
rect 45669 689697 45685 689731
rect 45585 689659 45685 689697
rect 45743 689731 45843 689747
rect 45743 689697 45759 689731
rect 45827 689697 45843 689731
rect 45743 689659 45843 689697
rect 45901 689731 46001 689747
rect 45901 689697 45917 689731
rect 45985 689697 46001 689731
rect 45901 689659 46001 689697
rect 44953 688621 45053 688659
rect 44953 688587 44969 688621
rect 45037 688587 45053 688621
rect 44953 688571 45053 688587
rect 45111 688621 45211 688659
rect 45111 688587 45127 688621
rect 45195 688587 45211 688621
rect 45111 688571 45211 688587
rect 45269 688621 45369 688659
rect 45269 688587 45285 688621
rect 45353 688587 45369 688621
rect 45269 688571 45369 688587
rect 45427 688621 45527 688659
rect 45427 688587 45443 688621
rect 45511 688587 45527 688621
rect 45427 688571 45527 688587
rect 45585 688621 45685 688659
rect 45585 688587 45601 688621
rect 45669 688587 45685 688621
rect 45585 688571 45685 688587
rect 45743 688621 45843 688659
rect 45743 688587 45759 688621
rect 45827 688587 45843 688621
rect 45743 688571 45843 688587
rect 45901 688621 46001 688659
rect 45901 688587 45917 688621
rect 45985 688587 46001 688621
rect 45901 688571 46001 688587
rect 44953 688211 45053 688227
rect 44953 688177 44969 688211
rect 45037 688177 45053 688211
rect 44953 688139 45053 688177
rect 45111 688211 45211 688227
rect 45111 688177 45127 688211
rect 45195 688177 45211 688211
rect 45111 688139 45211 688177
rect 45269 688211 45369 688227
rect 45269 688177 45285 688211
rect 45353 688177 45369 688211
rect 45269 688139 45369 688177
rect 45427 688211 45527 688227
rect 45427 688177 45443 688211
rect 45511 688177 45527 688211
rect 45427 688139 45527 688177
rect 45585 688211 45685 688227
rect 45585 688177 45601 688211
rect 45669 688177 45685 688211
rect 45585 688139 45685 688177
rect 45743 688211 45843 688227
rect 45743 688177 45759 688211
rect 45827 688177 45843 688211
rect 45743 688139 45843 688177
rect 45901 688211 46001 688227
rect 45901 688177 45917 688211
rect 45985 688177 46001 688211
rect 45901 688139 46001 688177
rect 44953 687101 45053 687139
rect 44953 687067 44969 687101
rect 45037 687067 45053 687101
rect 44953 687051 45053 687067
rect 45111 687101 45211 687139
rect 45111 687067 45127 687101
rect 45195 687067 45211 687101
rect 45111 687051 45211 687067
rect 45269 687101 45369 687139
rect 45269 687067 45285 687101
rect 45353 687067 45369 687101
rect 45269 687051 45369 687067
rect 45427 687101 45527 687139
rect 45427 687067 45443 687101
rect 45511 687067 45527 687101
rect 45427 687051 45527 687067
rect 45585 687101 45685 687139
rect 45585 687067 45601 687101
rect 45669 687067 45685 687101
rect 45585 687051 45685 687067
rect 45743 687101 45843 687139
rect 45743 687067 45759 687101
rect 45827 687067 45843 687101
rect 45743 687051 45843 687067
rect 45901 687101 46001 687139
rect 45901 687067 45917 687101
rect 45985 687067 46001 687101
rect 45901 687051 46001 687067
rect 43954 686690 44154 686706
rect 43954 686656 43970 686690
rect 44138 686656 44154 686690
rect 43954 686618 44154 686656
rect 44212 686690 44412 686706
rect 44212 686656 44228 686690
rect 44396 686656 44412 686690
rect 44212 686618 44412 686656
rect 44470 686690 44670 686706
rect 44470 686656 44486 686690
rect 44654 686656 44670 686690
rect 44470 686618 44670 686656
rect 44728 686690 44928 686706
rect 44728 686656 44744 686690
rect 44912 686656 44928 686690
rect 44728 686618 44928 686656
rect 44986 686690 45186 686706
rect 44986 686656 45002 686690
rect 45170 686656 45186 686690
rect 44986 686618 45186 686656
rect 45244 686690 45444 686706
rect 45244 686656 45260 686690
rect 45428 686656 45444 686690
rect 45244 686618 45444 686656
rect 45502 686690 45702 686706
rect 45502 686656 45518 686690
rect 45686 686656 45702 686690
rect 45502 686618 45702 686656
rect 45760 686690 45960 686706
rect 45760 686656 45776 686690
rect 45944 686656 45960 686690
rect 45760 686618 45960 686656
rect 46018 686690 46218 686706
rect 46018 686656 46034 686690
rect 46202 686656 46218 686690
rect 46018 686618 46218 686656
rect 46276 686690 46476 686706
rect 46276 686656 46292 686690
rect 46460 686656 46476 686690
rect 46276 686618 46476 686656
rect 46534 686690 46734 686706
rect 46534 686656 46550 686690
rect 46718 686656 46734 686690
rect 46534 686618 46734 686656
rect 46792 686690 46992 686706
rect 46792 686656 46808 686690
rect 46976 686656 46992 686690
rect 46792 686618 46992 686656
rect 43954 685580 44154 685618
rect 43954 685546 43970 685580
rect 44138 685546 44154 685580
rect 43954 685530 44154 685546
rect 44212 685580 44412 685618
rect 44212 685546 44228 685580
rect 44396 685546 44412 685580
rect 44212 685530 44412 685546
rect 44470 685580 44670 685618
rect 44470 685546 44486 685580
rect 44654 685546 44670 685580
rect 44470 685530 44670 685546
rect 44728 685580 44928 685618
rect 44728 685546 44744 685580
rect 44912 685546 44928 685580
rect 44728 685530 44928 685546
rect 44986 685580 45186 685618
rect 44986 685546 45002 685580
rect 45170 685546 45186 685580
rect 44986 685530 45186 685546
rect 45244 685580 45444 685618
rect 45244 685546 45260 685580
rect 45428 685546 45444 685580
rect 45244 685530 45444 685546
rect 45502 685580 45702 685618
rect 45502 685546 45518 685580
rect 45686 685546 45702 685580
rect 45502 685530 45702 685546
rect 45760 685580 45960 685618
rect 45760 685546 45776 685580
rect 45944 685546 45960 685580
rect 45760 685530 45960 685546
rect 46018 685580 46218 685618
rect 46018 685546 46034 685580
rect 46202 685546 46218 685580
rect 46018 685530 46218 685546
rect 46276 685580 46476 685618
rect 46276 685546 46292 685580
rect 46460 685546 46476 685580
rect 46276 685530 46476 685546
rect 46534 685580 46734 685618
rect 46534 685546 46550 685580
rect 46718 685546 46734 685580
rect 46534 685530 46734 685546
rect 46792 685580 46992 685618
rect 46792 685546 46808 685580
rect 46976 685546 46992 685580
rect 46792 685530 46992 685546
rect 43698 685170 43898 685186
rect 43698 685136 43714 685170
rect 43882 685136 43898 685170
rect 43698 685098 43898 685136
rect 43956 685170 44156 685186
rect 43956 685136 43972 685170
rect 44140 685136 44156 685170
rect 43956 685098 44156 685136
rect 44214 685170 44414 685186
rect 44214 685136 44230 685170
rect 44398 685136 44414 685170
rect 44214 685098 44414 685136
rect 44472 685170 44672 685186
rect 44472 685136 44488 685170
rect 44656 685136 44672 685170
rect 44472 685098 44672 685136
rect 44730 685170 44930 685186
rect 44730 685136 44746 685170
rect 44914 685136 44930 685170
rect 44730 685098 44930 685136
rect 44988 685170 45188 685186
rect 44988 685136 45004 685170
rect 45172 685136 45188 685170
rect 44988 685098 45188 685136
rect 45246 685170 45446 685186
rect 45246 685136 45262 685170
rect 45430 685136 45446 685170
rect 45246 685098 45446 685136
rect 45504 685170 45704 685186
rect 45504 685136 45520 685170
rect 45688 685136 45704 685170
rect 45504 685098 45704 685136
rect 45762 685170 45962 685186
rect 45762 685136 45778 685170
rect 45946 685136 45962 685170
rect 45762 685098 45962 685136
rect 46020 685170 46220 685186
rect 46020 685136 46036 685170
rect 46204 685136 46220 685170
rect 46020 685098 46220 685136
rect 46278 685170 46478 685186
rect 46278 685136 46294 685170
rect 46462 685136 46478 685170
rect 46278 685098 46478 685136
rect 46536 685170 46736 685186
rect 46536 685136 46552 685170
rect 46720 685136 46736 685170
rect 46536 685098 46736 685136
rect 46794 685170 46994 685186
rect 46794 685136 46810 685170
rect 46978 685136 46994 685170
rect 46794 685098 46994 685136
rect 47052 685170 47252 685186
rect 47052 685136 47068 685170
rect 47236 685136 47252 685170
rect 47052 685098 47252 685136
rect 43698 684060 43898 684098
rect 43698 684026 43714 684060
rect 43882 684026 43898 684060
rect 43698 684010 43898 684026
rect 43956 684060 44156 684098
rect 43956 684026 43972 684060
rect 44140 684026 44156 684060
rect 43956 684010 44156 684026
rect 44214 684060 44414 684098
rect 44214 684026 44230 684060
rect 44398 684026 44414 684060
rect 44214 684010 44414 684026
rect 44472 684060 44672 684098
rect 44472 684026 44488 684060
rect 44656 684026 44672 684060
rect 44472 684010 44672 684026
rect 44730 684060 44930 684098
rect 44730 684026 44746 684060
rect 44914 684026 44930 684060
rect 44730 684010 44930 684026
rect 44988 684060 45188 684098
rect 44988 684026 45004 684060
rect 45172 684026 45188 684060
rect 44988 684010 45188 684026
rect 45246 684060 45446 684098
rect 45246 684026 45262 684060
rect 45430 684026 45446 684060
rect 45246 684010 45446 684026
rect 45504 684060 45704 684098
rect 45504 684026 45520 684060
rect 45688 684026 45704 684060
rect 45504 684010 45704 684026
rect 45762 684060 45962 684098
rect 45762 684026 45778 684060
rect 45946 684026 45962 684060
rect 45762 684010 45962 684026
rect 46020 684060 46220 684098
rect 46020 684026 46036 684060
rect 46204 684026 46220 684060
rect 46020 684010 46220 684026
rect 46278 684060 46478 684098
rect 46278 684026 46294 684060
rect 46462 684026 46478 684060
rect 46278 684010 46478 684026
rect 46536 684060 46736 684098
rect 46536 684026 46552 684060
rect 46720 684026 46736 684060
rect 46536 684010 46736 684026
rect 46794 684060 46994 684098
rect 46794 684026 46810 684060
rect 46978 684026 46994 684060
rect 46794 684010 46994 684026
rect 47052 684060 47252 684098
rect 47052 684026 47068 684060
rect 47236 684026 47252 684060
rect 47052 684010 47252 684026
rect 41782 682808 41879 682824
rect 41782 682640 41798 682808
rect 41832 682640 41879 682808
rect 41782 682624 41879 682640
rect 42879 682808 42976 682824
rect 42879 682640 42926 682808
rect 42960 682640 42976 682808
rect 42879 682624 42976 682640
rect 43018 682808 43115 682824
rect 43018 682640 43034 682808
rect 43068 682640 43115 682808
rect 43018 682624 43115 682640
rect 44115 682808 44212 682824
rect 44115 682640 44162 682808
rect 44196 682640 44212 682808
rect 44115 682624 44212 682640
rect 44254 682808 44351 682824
rect 44254 682640 44270 682808
rect 44304 682640 44351 682808
rect 44254 682624 44351 682640
rect 45351 682808 45448 682824
rect 45351 682640 45398 682808
rect 45432 682640 45448 682808
rect 45351 682624 45448 682640
rect 45490 682808 45587 682824
rect 45490 682640 45506 682808
rect 45540 682640 45587 682808
rect 45490 682624 45587 682640
rect 46587 682808 46684 682824
rect 46587 682640 46634 682808
rect 46668 682640 46684 682808
rect 46587 682624 46684 682640
rect 46726 682808 46823 682824
rect 46726 682640 46742 682808
rect 46776 682640 46823 682808
rect 46726 682624 46823 682640
rect 47823 682808 47920 682824
rect 47823 682640 47870 682808
rect 47904 682640 47920 682808
rect 47823 682624 47920 682640
rect 47962 682808 48059 682824
rect 47962 682640 47978 682808
rect 48012 682640 48059 682808
rect 47962 682624 48059 682640
rect 49059 682808 49156 682824
rect 49059 682640 49106 682808
rect 49140 682640 49156 682808
rect 49059 682624 49156 682640
rect 41782 682218 41879 682234
rect 41782 682050 41798 682218
rect 41832 682050 41879 682218
rect 41782 682034 41879 682050
rect 42879 682218 42976 682234
rect 42879 682050 42926 682218
rect 42960 682050 42976 682218
rect 42879 682034 42976 682050
rect 43018 682218 43115 682234
rect 43018 682050 43034 682218
rect 43068 682050 43115 682218
rect 43018 682034 43115 682050
rect 44115 682218 44212 682234
rect 44115 682050 44162 682218
rect 44196 682050 44212 682218
rect 44115 682034 44212 682050
rect 44254 682218 44351 682234
rect 44254 682050 44270 682218
rect 44304 682050 44351 682218
rect 44254 682034 44351 682050
rect 45351 682218 45448 682234
rect 45351 682050 45398 682218
rect 45432 682050 45448 682218
rect 45351 682034 45448 682050
rect 45490 682218 45587 682234
rect 45490 682050 45506 682218
rect 45540 682050 45587 682218
rect 45490 682034 45587 682050
rect 46587 682218 46684 682234
rect 46587 682050 46634 682218
rect 46668 682050 46684 682218
rect 46587 682034 46684 682050
rect 46726 682218 46823 682234
rect 46726 682050 46742 682218
rect 46776 682050 46823 682218
rect 46726 682034 46823 682050
rect 47823 682218 47920 682234
rect 47823 682050 47870 682218
rect 47904 682050 47920 682218
rect 47823 682034 47920 682050
rect 47962 682218 48059 682234
rect 47962 682050 47978 682218
rect 48012 682050 48059 682218
rect 47962 682034 48059 682050
rect 49059 682218 49156 682234
rect 49059 682050 49106 682218
rect 49140 682050 49156 682218
rect 49059 682034 49156 682050
rect 44556 681428 44644 681444
rect 44556 681260 44572 681428
rect 44606 681260 44644 681428
rect 44556 681244 44644 681260
rect 44894 681428 44982 681444
rect 44894 681260 44932 681428
rect 44966 681260 44982 681428
rect 44894 681244 44982 681260
rect 45024 681428 45112 681444
rect 45024 681260 45040 681428
rect 45074 681260 45112 681428
rect 45024 681244 45112 681260
rect 45362 681428 45450 681444
rect 45362 681260 45400 681428
rect 45434 681260 45450 681428
rect 45362 681244 45450 681260
rect 45492 681428 45580 681444
rect 45492 681260 45508 681428
rect 45542 681260 45580 681428
rect 45492 681244 45580 681260
rect 45830 681428 45918 681444
rect 45830 681260 45868 681428
rect 45902 681260 45918 681428
rect 45830 681244 45918 681260
rect 45960 681428 46048 681444
rect 45960 681260 45976 681428
rect 46010 681260 46048 681428
rect 45960 681244 46048 681260
rect 46298 681428 46386 681444
rect 46298 681260 46336 681428
rect 46370 681260 46386 681428
rect 46298 681244 46386 681260
rect 44772 680803 44860 680819
rect 44772 680735 44788 680803
rect 44822 680735 44860 680803
rect 44772 680719 44860 680735
rect 45360 680803 45448 680819
rect 45360 680735 45398 680803
rect 45432 680735 45448 680803
rect 45360 680719 45448 680735
rect 45490 680803 45578 680819
rect 45490 680735 45506 680803
rect 45540 680735 45578 680803
rect 45490 680719 45578 680735
rect 46078 680803 46166 680819
rect 46078 680735 46116 680803
rect 46150 680735 46166 680803
rect 46078 680719 46166 680735
rect 41835 680278 41923 680294
rect 41835 680110 41851 680278
rect 41885 680110 41923 680278
rect 41835 680094 41923 680110
rect 42923 680278 43011 680294
rect 42923 680110 42961 680278
rect 42995 680110 43011 680278
rect 42923 680094 43011 680110
rect 43053 680278 43141 680294
rect 43053 680110 43069 680278
rect 43103 680110 43141 680278
rect 43053 680094 43141 680110
rect 44141 680278 44229 680294
rect 44141 680110 44179 680278
rect 44213 680110 44229 680278
rect 44141 680094 44229 680110
rect 44271 680278 44359 680294
rect 44271 680110 44287 680278
rect 44321 680110 44359 680278
rect 44271 680094 44359 680110
rect 45359 680278 45447 680294
rect 45359 680110 45397 680278
rect 45431 680110 45447 680278
rect 45359 680094 45447 680110
rect 45489 680278 45577 680294
rect 45489 680110 45505 680278
rect 45539 680110 45577 680278
rect 45489 680094 45577 680110
rect 46577 680278 46665 680294
rect 46577 680110 46615 680278
rect 46649 680110 46665 680278
rect 46577 680094 46665 680110
rect 46707 680278 46795 680294
rect 46707 680110 46723 680278
rect 46757 680110 46795 680278
rect 46707 680094 46795 680110
rect 47795 680278 47883 680294
rect 47795 680110 47833 680278
rect 47867 680110 47883 680278
rect 47795 680094 47883 680110
rect 47925 680278 48013 680294
rect 47925 680110 47941 680278
rect 47975 680110 48013 680278
rect 47925 680094 48013 680110
rect 49013 680278 49101 680294
rect 49013 680110 49051 680278
rect 49085 680110 49101 680278
rect 49013 680094 49101 680110
<< polycont >>
rect 42356 694484 42424 694518
rect 42514 694484 42582 694518
rect 42672 694484 42740 694518
rect 42830 694484 42898 694518
rect 42988 694484 43056 694518
rect 43146 694484 43214 694518
rect 43304 694484 43372 694518
rect 43462 694484 43530 694518
rect 43620 694484 43688 694518
rect 43778 694484 43846 694518
rect 43936 694484 44004 694518
rect 44094 694484 44162 694518
rect 44252 694484 44320 694518
rect 44410 694484 44478 694518
rect 44568 694484 44636 694518
rect 44726 694484 44794 694518
rect 44884 694484 44952 694518
rect 45042 694484 45110 694518
rect 45200 694484 45268 694518
rect 45358 694484 45426 694518
rect 45516 694484 45584 694518
rect 45674 694484 45742 694518
rect 45832 694484 45900 694518
rect 45990 694484 46058 694518
rect 46148 694484 46216 694518
rect 46306 694484 46374 694518
rect 46464 694484 46532 694518
rect 46622 694484 46690 694518
rect 46780 694484 46848 694518
rect 46938 694484 47006 694518
rect 47096 694484 47164 694518
rect 47254 694484 47322 694518
rect 47412 694484 47480 694518
rect 47570 694484 47638 694518
rect 47728 694484 47796 694518
rect 47886 694484 47954 694518
rect 48044 694484 48112 694518
rect 48202 694484 48270 694518
rect 48360 694484 48428 694518
rect 48518 694484 48586 694518
rect 42356 693356 42424 693390
rect 42514 693356 42582 693390
rect 42672 693356 42740 693390
rect 42830 693356 42898 693390
rect 42988 693356 43056 693390
rect 43146 693356 43214 693390
rect 43304 693356 43372 693390
rect 43462 693356 43530 693390
rect 43620 693356 43688 693390
rect 43778 693356 43846 693390
rect 43936 693356 44004 693390
rect 44094 693356 44162 693390
rect 44252 693356 44320 693390
rect 44410 693356 44478 693390
rect 44568 693356 44636 693390
rect 44726 693356 44794 693390
rect 44884 693356 44952 693390
rect 45042 693356 45110 693390
rect 45200 693356 45268 693390
rect 45358 693356 45426 693390
rect 45516 693356 45584 693390
rect 45674 693356 45742 693390
rect 45832 693356 45900 693390
rect 45990 693356 46058 693390
rect 46148 693356 46216 693390
rect 46306 693356 46374 693390
rect 46464 693356 46532 693390
rect 46622 693356 46690 693390
rect 46780 693356 46848 693390
rect 46938 693356 47006 693390
rect 47096 693356 47164 693390
rect 47254 693356 47322 693390
rect 47412 693356 47480 693390
rect 47570 693356 47638 693390
rect 47728 693356 47796 693390
rect 47886 693356 47954 693390
rect 48044 693356 48112 693390
rect 48202 693356 48270 693390
rect 48360 693356 48428 693390
rect 48518 693356 48586 693390
rect 43858 692814 43926 692848
rect 44016 692814 44084 692848
rect 44174 692814 44242 692848
rect 44332 692814 44400 692848
rect 44490 692814 44558 692848
rect 44648 692814 44716 692848
rect 44806 692814 44874 692848
rect 44964 692814 45032 692848
rect 45122 692814 45190 692848
rect 45280 692814 45348 692848
rect 45438 692814 45506 692848
rect 45596 692814 45664 692848
rect 45754 692814 45822 692848
rect 45912 692814 45980 692848
rect 46070 692814 46138 692848
rect 46228 692814 46296 692848
rect 46386 692814 46454 692848
rect 46544 692814 46612 692848
rect 46702 692814 46770 692848
rect 46860 692814 46928 692848
rect 47018 692814 47086 692848
rect 43858 691686 43926 691720
rect 44016 691686 44084 691720
rect 44174 691686 44242 691720
rect 44332 691686 44400 691720
rect 44490 691686 44558 691720
rect 44648 691686 44716 691720
rect 44806 691686 44874 691720
rect 44964 691686 45032 691720
rect 45122 691686 45190 691720
rect 45280 691686 45348 691720
rect 45438 691686 45506 691720
rect 45596 691686 45664 691720
rect 45754 691686 45822 691720
rect 45912 691686 45980 691720
rect 46070 691686 46138 691720
rect 46228 691686 46296 691720
rect 46386 691686 46454 691720
rect 46544 691686 46612 691720
rect 46702 691686 46770 691720
rect 46860 691686 46928 691720
rect 47018 691686 47086 691720
rect 43858 691274 43926 691308
rect 44016 691274 44084 691308
rect 44174 691274 44242 691308
rect 44332 691274 44400 691308
rect 44490 691274 44558 691308
rect 44648 691274 44716 691308
rect 44806 691274 44874 691308
rect 44964 691274 45032 691308
rect 45122 691274 45190 691308
rect 45280 691274 45348 691308
rect 45438 691274 45506 691308
rect 45596 691274 45664 691308
rect 45754 691274 45822 691308
rect 45912 691274 45980 691308
rect 46070 691274 46138 691308
rect 46228 691274 46296 691308
rect 46386 691274 46454 691308
rect 46544 691274 46612 691308
rect 46702 691274 46770 691308
rect 46860 691274 46928 691308
rect 47018 691274 47086 691308
rect 43858 690146 43926 690180
rect 44016 690146 44084 690180
rect 44174 690146 44242 690180
rect 44332 690146 44400 690180
rect 44490 690146 44558 690180
rect 44648 690146 44716 690180
rect 44806 690146 44874 690180
rect 44964 690146 45032 690180
rect 45122 690146 45190 690180
rect 45280 690146 45348 690180
rect 45438 690146 45506 690180
rect 45596 690146 45664 690180
rect 45754 690146 45822 690180
rect 45912 690146 45980 690180
rect 46070 690146 46138 690180
rect 46228 690146 46296 690180
rect 46386 690146 46454 690180
rect 46544 690146 46612 690180
rect 46702 690146 46770 690180
rect 46860 690146 46928 690180
rect 47018 690146 47086 690180
rect 44969 689697 45037 689731
rect 45127 689697 45195 689731
rect 45285 689697 45353 689731
rect 45443 689697 45511 689731
rect 45601 689697 45669 689731
rect 45759 689697 45827 689731
rect 45917 689697 45985 689731
rect 44969 688587 45037 688621
rect 45127 688587 45195 688621
rect 45285 688587 45353 688621
rect 45443 688587 45511 688621
rect 45601 688587 45669 688621
rect 45759 688587 45827 688621
rect 45917 688587 45985 688621
rect 44969 688177 45037 688211
rect 45127 688177 45195 688211
rect 45285 688177 45353 688211
rect 45443 688177 45511 688211
rect 45601 688177 45669 688211
rect 45759 688177 45827 688211
rect 45917 688177 45985 688211
rect 44969 687067 45037 687101
rect 45127 687067 45195 687101
rect 45285 687067 45353 687101
rect 45443 687067 45511 687101
rect 45601 687067 45669 687101
rect 45759 687067 45827 687101
rect 45917 687067 45985 687101
rect 43970 686656 44138 686690
rect 44228 686656 44396 686690
rect 44486 686656 44654 686690
rect 44744 686656 44912 686690
rect 45002 686656 45170 686690
rect 45260 686656 45428 686690
rect 45518 686656 45686 686690
rect 45776 686656 45944 686690
rect 46034 686656 46202 686690
rect 46292 686656 46460 686690
rect 46550 686656 46718 686690
rect 46808 686656 46976 686690
rect 43970 685546 44138 685580
rect 44228 685546 44396 685580
rect 44486 685546 44654 685580
rect 44744 685546 44912 685580
rect 45002 685546 45170 685580
rect 45260 685546 45428 685580
rect 45518 685546 45686 685580
rect 45776 685546 45944 685580
rect 46034 685546 46202 685580
rect 46292 685546 46460 685580
rect 46550 685546 46718 685580
rect 46808 685546 46976 685580
rect 43714 685136 43882 685170
rect 43972 685136 44140 685170
rect 44230 685136 44398 685170
rect 44488 685136 44656 685170
rect 44746 685136 44914 685170
rect 45004 685136 45172 685170
rect 45262 685136 45430 685170
rect 45520 685136 45688 685170
rect 45778 685136 45946 685170
rect 46036 685136 46204 685170
rect 46294 685136 46462 685170
rect 46552 685136 46720 685170
rect 46810 685136 46978 685170
rect 47068 685136 47236 685170
rect 43714 684026 43882 684060
rect 43972 684026 44140 684060
rect 44230 684026 44398 684060
rect 44488 684026 44656 684060
rect 44746 684026 44914 684060
rect 45004 684026 45172 684060
rect 45262 684026 45430 684060
rect 45520 684026 45688 684060
rect 45778 684026 45946 684060
rect 46036 684026 46204 684060
rect 46294 684026 46462 684060
rect 46552 684026 46720 684060
rect 46810 684026 46978 684060
rect 47068 684026 47236 684060
rect 41798 682640 41832 682808
rect 42926 682640 42960 682808
rect 43034 682640 43068 682808
rect 44162 682640 44196 682808
rect 44270 682640 44304 682808
rect 45398 682640 45432 682808
rect 45506 682640 45540 682808
rect 46634 682640 46668 682808
rect 46742 682640 46776 682808
rect 47870 682640 47904 682808
rect 47978 682640 48012 682808
rect 49106 682640 49140 682808
rect 41798 682050 41832 682218
rect 42926 682050 42960 682218
rect 43034 682050 43068 682218
rect 44162 682050 44196 682218
rect 44270 682050 44304 682218
rect 45398 682050 45432 682218
rect 45506 682050 45540 682218
rect 46634 682050 46668 682218
rect 46742 682050 46776 682218
rect 47870 682050 47904 682218
rect 47978 682050 48012 682218
rect 49106 682050 49140 682218
rect 44572 681260 44606 681428
rect 44932 681260 44966 681428
rect 45040 681260 45074 681428
rect 45400 681260 45434 681428
rect 45508 681260 45542 681428
rect 45868 681260 45902 681428
rect 45976 681260 46010 681428
rect 46336 681260 46370 681428
rect 44788 680735 44822 680803
rect 45398 680735 45432 680803
rect 45506 680735 45540 680803
rect 46116 680735 46150 680803
rect 41851 680110 41885 680278
rect 42961 680110 42995 680278
rect 43069 680110 43103 680278
rect 44179 680110 44213 680278
rect 44287 680110 44321 680278
rect 45397 680110 45431 680278
rect 45505 680110 45539 680278
rect 46615 680110 46649 680278
rect 46723 680110 46757 680278
rect 47833 680110 47867 680278
rect 47941 680110 47975 680278
rect 49051 680110 49085 680278
<< xpolycontact >>
rect 38501 694221 38933 695367
rect 40933 694221 41365 695367
rect 38501 692761 38933 693907
rect 40933 692761 41365 693907
rect 49571 694221 50003 695367
rect 52003 694221 52435 695367
rect 49571 692761 50003 693907
rect 52003 692761 52435 693907
rect 42625 679176 43771 679608
rect 42625 664944 43771 665376
rect 44135 679176 45281 679608
rect 44135 664944 45281 665376
rect 45645 679170 46791 679602
rect 45645 664938 46791 665370
rect 47165 679170 48311 679602
rect 47165 664938 48311 665370
<< xpolyres >>
rect 38933 694221 40933 695367
rect 38933 692761 40933 693907
rect 50003 694221 52003 695367
rect 50003 692761 52003 693907
rect 42625 665376 43771 679176
rect 44135 665376 45281 679176
rect 45645 665370 46791 679170
rect 47165 665370 48311 679170
<< locali >>
rect 38371 695463 38467 695497
rect 41399 695463 41495 695497
rect 38371 695401 38405 695463
rect 41461 695401 41495 695463
rect 38371 694125 38405 694187
rect 49441 695463 49537 695497
rect 52469 695463 52565 695497
rect 49441 695401 49475 695463
rect 39548 694125 40208 694128
rect 41461 694125 41495 694187
rect 38371 694091 38467 694125
rect 41399 694091 41495 694125
rect 42180 694586 42276 694620
rect 48666 694586 48762 694620
rect 42180 694524 42214 694586
rect 39548 694037 40208 694091
rect 38371 694003 38467 694037
rect 41399 694003 41495 694037
rect 38371 693941 38405 694003
rect 41461 693941 41495 694003
rect 38371 692665 38405 692727
rect 48728 694524 48762 694586
rect 42340 694484 42356 694518
rect 42424 694484 42440 694518
rect 42498 694484 42514 694518
rect 42582 694484 42598 694518
rect 42656 694484 42672 694518
rect 42740 694484 42756 694518
rect 42814 694484 42830 694518
rect 42898 694484 42914 694518
rect 42972 694484 42988 694518
rect 43056 694484 43072 694518
rect 43130 694484 43146 694518
rect 43214 694484 43230 694518
rect 43288 694484 43304 694518
rect 43372 694484 43388 694518
rect 43446 694484 43462 694518
rect 43530 694484 43546 694518
rect 43604 694484 43620 694518
rect 43688 694484 43704 694518
rect 43762 694484 43778 694518
rect 43846 694484 43862 694518
rect 43920 694484 43936 694518
rect 44004 694484 44020 694518
rect 44078 694484 44094 694518
rect 44162 694484 44178 694518
rect 44236 694484 44252 694518
rect 44320 694484 44336 694518
rect 44394 694484 44410 694518
rect 44478 694484 44494 694518
rect 44552 694484 44568 694518
rect 44636 694484 44652 694518
rect 44710 694484 44726 694518
rect 44794 694484 44810 694518
rect 44868 694484 44884 694518
rect 44952 694484 44968 694518
rect 45026 694484 45042 694518
rect 45110 694484 45126 694518
rect 45184 694484 45200 694518
rect 45268 694484 45284 694518
rect 45342 694484 45358 694518
rect 45426 694484 45442 694518
rect 45500 694484 45516 694518
rect 45584 694484 45600 694518
rect 45658 694484 45674 694518
rect 45742 694484 45758 694518
rect 45816 694484 45832 694518
rect 45900 694484 45916 694518
rect 45974 694484 45990 694518
rect 46058 694484 46074 694518
rect 46132 694484 46148 694518
rect 46216 694484 46232 694518
rect 46290 694484 46306 694518
rect 46374 694484 46390 694518
rect 46448 694484 46464 694518
rect 46532 694484 46548 694518
rect 46606 694484 46622 694518
rect 46690 694484 46706 694518
rect 46764 694484 46780 694518
rect 46848 694484 46864 694518
rect 46922 694484 46938 694518
rect 47006 694484 47022 694518
rect 47080 694484 47096 694518
rect 47164 694484 47180 694518
rect 47238 694484 47254 694518
rect 47322 694484 47338 694518
rect 47396 694484 47412 694518
rect 47480 694484 47496 694518
rect 47554 694484 47570 694518
rect 47638 694484 47654 694518
rect 47712 694484 47728 694518
rect 47796 694484 47812 694518
rect 47870 694484 47886 694518
rect 47954 694484 47970 694518
rect 48028 694484 48044 694518
rect 48112 694484 48128 694518
rect 48186 694484 48202 694518
rect 48270 694484 48286 694518
rect 48344 694484 48360 694518
rect 48428 694484 48444 694518
rect 48502 694484 48518 694518
rect 48586 694484 48602 694518
rect 42294 694425 42328 694441
rect 42294 693433 42328 693449
rect 42452 694425 42486 694441
rect 42452 693433 42486 693449
rect 42610 694425 42644 694441
rect 42610 693433 42644 693449
rect 42768 694425 42802 694441
rect 42768 693433 42802 693449
rect 42926 694425 42960 694441
rect 42926 693433 42960 693449
rect 43084 694425 43118 694441
rect 43084 693433 43118 693449
rect 43242 694425 43276 694441
rect 43242 693433 43276 693449
rect 43400 694425 43434 694441
rect 43400 693433 43434 693449
rect 43558 694425 43592 694441
rect 43558 693433 43592 693449
rect 43716 694425 43750 694441
rect 43716 693433 43750 693449
rect 43874 694425 43908 694441
rect 43874 693433 43908 693449
rect 44032 694425 44066 694441
rect 44032 693433 44066 693449
rect 44190 694425 44224 694441
rect 44190 693433 44224 693449
rect 44348 694425 44382 694441
rect 44348 693433 44382 693449
rect 44506 694425 44540 694441
rect 44506 693433 44540 693449
rect 44664 694425 44698 694441
rect 44664 693433 44698 693449
rect 44822 694425 44856 694441
rect 44822 693433 44856 693449
rect 44980 694425 45014 694441
rect 44980 693433 45014 693449
rect 45138 694425 45172 694441
rect 45138 693433 45172 693449
rect 45296 694425 45330 694441
rect 45296 693433 45330 693449
rect 45454 694425 45488 694441
rect 45454 693433 45488 693449
rect 45612 694425 45646 694441
rect 45612 693433 45646 693449
rect 45770 694425 45804 694441
rect 45770 693433 45804 693449
rect 45928 694425 45962 694441
rect 45928 693433 45962 693449
rect 46086 694425 46120 694441
rect 46086 693433 46120 693449
rect 46244 694425 46278 694441
rect 46244 693433 46278 693449
rect 46402 694425 46436 694441
rect 46402 693433 46436 693449
rect 46560 694425 46594 694441
rect 46560 693433 46594 693449
rect 46718 694425 46752 694441
rect 46718 693433 46752 693449
rect 46876 694425 46910 694441
rect 46876 693433 46910 693449
rect 47034 694425 47068 694441
rect 47034 693433 47068 693449
rect 47192 694425 47226 694441
rect 47192 693433 47226 693449
rect 47350 694425 47384 694441
rect 47350 693433 47384 693449
rect 47508 694425 47542 694441
rect 47508 693433 47542 693449
rect 47666 694425 47700 694441
rect 47666 693433 47700 693449
rect 47824 694425 47858 694441
rect 47824 693433 47858 693449
rect 47982 694425 48016 694441
rect 47982 693433 48016 693449
rect 48140 694425 48174 694441
rect 48140 693433 48174 693449
rect 48298 694425 48332 694441
rect 48298 693433 48332 693449
rect 48456 694425 48490 694441
rect 48456 693433 48490 693449
rect 48614 694425 48648 694441
rect 48614 693433 48648 693449
rect 42340 693356 42356 693390
rect 42424 693356 42440 693390
rect 42498 693356 42514 693390
rect 42582 693356 42598 693390
rect 42656 693356 42672 693390
rect 42740 693356 42756 693390
rect 42814 693356 42830 693390
rect 42898 693356 42914 693390
rect 42972 693356 42988 693390
rect 43056 693356 43072 693390
rect 43130 693356 43146 693390
rect 43214 693356 43230 693390
rect 43288 693356 43304 693390
rect 43372 693356 43388 693390
rect 43446 693356 43462 693390
rect 43530 693356 43546 693390
rect 43604 693356 43620 693390
rect 43688 693356 43704 693390
rect 43762 693356 43778 693390
rect 43846 693356 43862 693390
rect 43920 693356 43936 693390
rect 44004 693356 44020 693390
rect 44078 693356 44094 693390
rect 44162 693356 44178 693390
rect 44236 693356 44252 693390
rect 44320 693356 44336 693390
rect 44394 693356 44410 693390
rect 44478 693356 44494 693390
rect 44552 693356 44568 693390
rect 44636 693356 44652 693390
rect 44710 693356 44726 693390
rect 44794 693356 44810 693390
rect 44868 693356 44884 693390
rect 44952 693356 44968 693390
rect 45026 693356 45042 693390
rect 45110 693356 45126 693390
rect 45184 693356 45200 693390
rect 45268 693356 45284 693390
rect 45342 693356 45358 693390
rect 45426 693356 45442 693390
rect 45500 693356 45516 693390
rect 45584 693356 45600 693390
rect 45658 693356 45674 693390
rect 45742 693356 45758 693390
rect 45816 693356 45832 693390
rect 45900 693356 45916 693390
rect 45974 693356 45990 693390
rect 46058 693356 46074 693390
rect 46132 693356 46148 693390
rect 46216 693356 46232 693390
rect 46290 693356 46306 693390
rect 46374 693356 46390 693390
rect 46448 693356 46464 693390
rect 46532 693356 46548 693390
rect 46606 693356 46622 693390
rect 46690 693356 46706 693390
rect 46764 693356 46780 693390
rect 46848 693356 46864 693390
rect 46922 693356 46938 693390
rect 47006 693356 47022 693390
rect 47080 693356 47096 693390
rect 47164 693356 47180 693390
rect 47238 693356 47254 693390
rect 47322 693356 47338 693390
rect 47396 693356 47412 693390
rect 47480 693356 47496 693390
rect 47554 693356 47570 693390
rect 47638 693356 47654 693390
rect 47712 693356 47728 693390
rect 47796 693356 47812 693390
rect 47870 693356 47886 693390
rect 47954 693356 47970 693390
rect 48028 693356 48044 693390
rect 48112 693356 48128 693390
rect 48186 693356 48202 693390
rect 48270 693356 48286 693390
rect 48344 693356 48360 693390
rect 48428 693356 48444 693390
rect 48502 693356 48518 693390
rect 48586 693356 48602 693390
rect 42180 693288 42214 693350
rect 52531 695401 52565 695463
rect 49441 694125 49475 694187
rect 50798 694125 51458 694128
rect 52531 694125 52565 694187
rect 49441 694091 49537 694125
rect 52469 694091 52565 694125
rect 50798 694037 51458 694091
rect 48728 693288 48762 693350
rect 42180 693254 42276 693288
rect 48666 693254 48762 693288
rect 49441 694003 49537 694037
rect 52469 694003 52565 694037
rect 49441 693941 49475 694003
rect 41461 692665 41495 692727
rect 38371 692631 38467 692665
rect 41399 692631 41495 692665
rect 43682 692916 43778 692950
rect 47166 692916 47262 692950
rect 43682 692854 43716 692916
rect 47228 692854 47262 692916
rect 43842 692814 43858 692848
rect 43926 692814 43942 692848
rect 44000 692814 44016 692848
rect 44084 692814 44100 692848
rect 44158 692814 44174 692848
rect 44242 692814 44258 692848
rect 44316 692814 44332 692848
rect 44400 692814 44416 692848
rect 44474 692814 44490 692848
rect 44558 692814 44574 692848
rect 44632 692814 44648 692848
rect 44716 692814 44732 692848
rect 44790 692814 44806 692848
rect 44874 692814 44890 692848
rect 44948 692814 44964 692848
rect 45032 692814 45048 692848
rect 45106 692814 45122 692848
rect 45190 692814 45206 692848
rect 45264 692814 45280 692848
rect 45348 692814 45364 692848
rect 45422 692814 45438 692848
rect 45506 692814 45522 692848
rect 45580 692814 45596 692848
rect 45664 692814 45680 692848
rect 45738 692814 45754 692848
rect 45822 692814 45838 692848
rect 45896 692814 45912 692848
rect 45980 692814 45996 692848
rect 46054 692814 46070 692848
rect 46138 692814 46154 692848
rect 46212 692814 46228 692848
rect 46296 692814 46312 692848
rect 46370 692814 46386 692848
rect 46454 692814 46470 692848
rect 46528 692814 46544 692848
rect 46612 692814 46628 692848
rect 46686 692814 46702 692848
rect 46770 692814 46786 692848
rect 46844 692814 46860 692848
rect 46928 692814 46944 692848
rect 47002 692814 47018 692848
rect 47086 692814 47102 692848
rect 43796 692755 43830 692771
rect 43796 691763 43830 691779
rect 43954 692755 43988 692771
rect 43954 691763 43988 691779
rect 44112 692755 44146 692771
rect 44112 691763 44146 691779
rect 44270 692755 44304 692771
rect 44270 691763 44304 691779
rect 44428 692755 44462 692771
rect 44428 691763 44462 691779
rect 44586 692755 44620 692771
rect 44586 691763 44620 691779
rect 44744 692755 44778 692771
rect 44744 691763 44778 691779
rect 44902 692755 44936 692771
rect 44902 691763 44936 691779
rect 45060 692755 45094 692771
rect 45060 691763 45094 691779
rect 45218 692755 45252 692771
rect 45218 691763 45252 691779
rect 45376 692755 45410 692771
rect 45376 691763 45410 691779
rect 45534 692755 45568 692771
rect 45534 691763 45568 691779
rect 45692 692755 45726 692771
rect 45692 691763 45726 691779
rect 45850 692755 45884 692771
rect 45850 691763 45884 691779
rect 46008 692755 46042 692771
rect 46008 691763 46042 691779
rect 46166 692755 46200 692771
rect 46166 691763 46200 691779
rect 46324 692755 46358 692771
rect 46324 691763 46358 691779
rect 46482 692755 46516 692771
rect 46482 691763 46516 691779
rect 46640 692755 46674 692771
rect 46640 691763 46674 691779
rect 46798 692755 46832 692771
rect 46798 691763 46832 691779
rect 46956 692755 46990 692771
rect 46956 691763 46990 691779
rect 47114 692755 47148 692771
rect 47114 691763 47148 691779
rect 43842 691686 43858 691720
rect 43926 691686 43942 691720
rect 44000 691686 44016 691720
rect 44084 691686 44100 691720
rect 44158 691686 44174 691720
rect 44242 691686 44258 691720
rect 44316 691686 44332 691720
rect 44400 691686 44416 691720
rect 44474 691686 44490 691720
rect 44558 691686 44574 691720
rect 44632 691686 44648 691720
rect 44716 691686 44732 691720
rect 44790 691686 44806 691720
rect 44874 691686 44890 691720
rect 44948 691686 44964 691720
rect 45032 691686 45048 691720
rect 45106 691686 45122 691720
rect 45190 691686 45206 691720
rect 45264 691686 45280 691720
rect 45348 691686 45364 691720
rect 45422 691686 45438 691720
rect 45506 691686 45522 691720
rect 45580 691686 45596 691720
rect 45664 691686 45680 691720
rect 45738 691686 45754 691720
rect 45822 691686 45838 691720
rect 45896 691686 45912 691720
rect 45980 691686 45996 691720
rect 46054 691686 46070 691720
rect 46138 691686 46154 691720
rect 46212 691686 46228 691720
rect 46296 691686 46312 691720
rect 46370 691686 46386 691720
rect 46454 691686 46470 691720
rect 46528 691686 46544 691720
rect 46612 691686 46628 691720
rect 46686 691686 46702 691720
rect 46770 691686 46786 691720
rect 46844 691686 46860 691720
rect 46928 691686 46944 691720
rect 47002 691686 47018 691720
rect 47086 691686 47102 691720
rect 43682 691618 43716 691680
rect 52531 693941 52565 694003
rect 49441 692665 49475 692727
rect 52531 692665 52565 692727
rect 49441 692631 49537 692665
rect 52469 692631 52565 692665
rect 47228 691618 47262 691680
rect 43682 691584 43778 691618
rect 47166 691584 47262 691618
rect 43682 691376 43778 691410
rect 47166 691376 47262 691410
rect 43682 691314 43716 691376
rect 47228 691314 47262 691376
rect 43842 691274 43858 691308
rect 43926 691274 43942 691308
rect 44000 691274 44016 691308
rect 44084 691274 44100 691308
rect 44158 691274 44174 691308
rect 44242 691274 44258 691308
rect 44316 691274 44332 691308
rect 44400 691274 44416 691308
rect 44474 691274 44490 691308
rect 44558 691274 44574 691308
rect 44632 691274 44648 691308
rect 44716 691274 44732 691308
rect 44790 691274 44806 691308
rect 44874 691274 44890 691308
rect 44948 691274 44964 691308
rect 45032 691274 45048 691308
rect 45106 691274 45122 691308
rect 45190 691274 45206 691308
rect 45264 691274 45280 691308
rect 45348 691274 45364 691308
rect 45422 691274 45438 691308
rect 45506 691274 45522 691308
rect 45580 691274 45596 691308
rect 45664 691274 45680 691308
rect 45738 691274 45754 691308
rect 45822 691274 45838 691308
rect 45896 691274 45912 691308
rect 45980 691274 45996 691308
rect 46054 691274 46070 691308
rect 46138 691274 46154 691308
rect 46212 691274 46228 691308
rect 46296 691274 46312 691308
rect 46370 691274 46386 691308
rect 46454 691274 46470 691308
rect 46528 691274 46544 691308
rect 46612 691274 46628 691308
rect 46686 691274 46702 691308
rect 46770 691274 46786 691308
rect 46844 691274 46860 691308
rect 46928 691274 46944 691308
rect 47002 691274 47018 691308
rect 47086 691274 47102 691308
rect 43796 691215 43830 691231
rect 43796 690223 43830 690239
rect 43954 691215 43988 691231
rect 43954 690223 43988 690239
rect 44112 691215 44146 691231
rect 44112 690223 44146 690239
rect 44270 691215 44304 691231
rect 44270 690223 44304 690239
rect 44428 691215 44462 691231
rect 44428 690223 44462 690239
rect 44586 691215 44620 691231
rect 44586 690223 44620 690239
rect 44744 691215 44778 691231
rect 44744 690223 44778 690239
rect 44902 691215 44936 691231
rect 44902 690223 44936 690239
rect 45060 691215 45094 691231
rect 45060 690223 45094 690239
rect 45218 691215 45252 691231
rect 45218 690223 45252 690239
rect 45376 691215 45410 691231
rect 45376 690223 45410 690239
rect 45534 691215 45568 691231
rect 45534 690223 45568 690239
rect 45692 691215 45726 691231
rect 45692 690223 45726 690239
rect 45850 691215 45884 691231
rect 45850 690223 45884 690239
rect 46008 691215 46042 691231
rect 46008 690223 46042 690239
rect 46166 691215 46200 691231
rect 46166 690223 46200 690239
rect 46324 691215 46358 691231
rect 46324 690223 46358 690239
rect 46482 691215 46516 691231
rect 46482 690223 46516 690239
rect 46640 691215 46674 691231
rect 46640 690223 46674 690239
rect 46798 691215 46832 691231
rect 46798 690223 46832 690239
rect 46956 691215 46990 691231
rect 46956 690223 46990 690239
rect 47114 691215 47148 691231
rect 47114 690223 47148 690239
rect 43842 690146 43858 690180
rect 43926 690146 43942 690180
rect 44000 690146 44016 690180
rect 44084 690146 44100 690180
rect 44158 690146 44174 690180
rect 44242 690146 44258 690180
rect 44316 690146 44332 690180
rect 44400 690146 44416 690180
rect 44474 690146 44490 690180
rect 44558 690146 44574 690180
rect 44632 690146 44648 690180
rect 44716 690146 44732 690180
rect 44790 690146 44806 690180
rect 44874 690146 44890 690180
rect 44948 690146 44964 690180
rect 45032 690146 45048 690180
rect 45106 690146 45122 690180
rect 45190 690146 45206 690180
rect 45264 690146 45280 690180
rect 45348 690146 45364 690180
rect 45422 690146 45438 690180
rect 45506 690146 45522 690180
rect 45580 690146 45596 690180
rect 45664 690146 45680 690180
rect 45738 690146 45754 690180
rect 45822 690146 45838 690180
rect 45896 690146 45912 690180
rect 45980 690146 45996 690180
rect 46054 690146 46070 690180
rect 46138 690146 46154 690180
rect 46212 690146 46228 690180
rect 46296 690146 46312 690180
rect 46370 690146 46386 690180
rect 46454 690146 46470 690180
rect 46528 690146 46544 690180
rect 46612 690146 46628 690180
rect 46686 690146 46702 690180
rect 46770 690146 46786 690180
rect 46844 690146 46860 690180
rect 46928 690146 46944 690180
rect 47002 690146 47018 690180
rect 47086 690146 47102 690180
rect 43682 690078 43716 690140
rect 47228 690078 47262 690140
rect 43682 690044 43778 690078
rect 47166 690044 47262 690078
rect 44793 689799 44889 689833
rect 46065 689799 46161 689833
rect 44793 689737 44827 689799
rect 46127 689737 46161 689799
rect 44953 689697 44969 689731
rect 45037 689697 45053 689731
rect 45111 689697 45127 689731
rect 45195 689697 45211 689731
rect 45269 689697 45285 689731
rect 45353 689697 45369 689731
rect 45427 689697 45443 689731
rect 45511 689697 45527 689731
rect 45585 689697 45601 689731
rect 45669 689697 45685 689731
rect 45743 689697 45759 689731
rect 45827 689697 45843 689731
rect 45901 689697 45917 689731
rect 45985 689697 46001 689731
rect 44907 689647 44941 689663
rect 44907 688655 44941 688671
rect 45065 689647 45099 689663
rect 45065 688655 45099 688671
rect 45223 689647 45257 689663
rect 45223 688655 45257 688671
rect 45381 689647 45415 689663
rect 45381 688655 45415 688671
rect 45539 689647 45573 689663
rect 45539 688655 45573 688671
rect 45697 689647 45731 689663
rect 45697 688655 45731 688671
rect 45855 689647 45889 689663
rect 45855 688655 45889 688671
rect 46013 689647 46047 689663
rect 46013 688655 46047 688671
rect 44953 688587 44969 688621
rect 45037 688587 45053 688621
rect 45111 688587 45127 688621
rect 45195 688587 45211 688621
rect 45269 688587 45285 688621
rect 45353 688587 45369 688621
rect 45427 688587 45443 688621
rect 45511 688587 45527 688621
rect 45585 688587 45601 688621
rect 45669 688587 45685 688621
rect 45743 688587 45759 688621
rect 45827 688587 45843 688621
rect 45901 688587 45917 688621
rect 45985 688587 46001 688621
rect 44793 688519 44827 688581
rect 46127 688519 46161 688581
rect 44793 688485 44889 688519
rect 46065 688485 46161 688519
rect 44793 688279 44889 688313
rect 46065 688279 46161 688313
rect 44793 688217 44827 688279
rect 46127 688217 46161 688279
rect 44953 688177 44969 688211
rect 45037 688177 45053 688211
rect 45111 688177 45127 688211
rect 45195 688177 45211 688211
rect 45269 688177 45285 688211
rect 45353 688177 45369 688211
rect 45427 688177 45443 688211
rect 45511 688177 45527 688211
rect 45585 688177 45601 688211
rect 45669 688177 45685 688211
rect 45743 688177 45759 688211
rect 45827 688177 45843 688211
rect 45901 688177 45917 688211
rect 45985 688177 46001 688211
rect 44907 688127 44941 688143
rect 44907 687135 44941 687151
rect 45065 688127 45099 688143
rect 45065 687135 45099 687151
rect 45223 688127 45257 688143
rect 45223 687135 45257 687151
rect 45381 688127 45415 688143
rect 45381 687135 45415 687151
rect 45539 688127 45573 688143
rect 45539 687135 45573 687151
rect 45697 688127 45731 688143
rect 45697 687135 45731 687151
rect 45855 688127 45889 688143
rect 45855 687135 45889 687151
rect 46013 688127 46047 688143
rect 46013 687135 46047 687151
rect 44953 687067 44969 687101
rect 45037 687067 45053 687101
rect 45111 687067 45127 687101
rect 45195 687067 45211 687101
rect 45269 687067 45285 687101
rect 45353 687067 45369 687101
rect 45427 687067 45443 687101
rect 45511 687067 45527 687101
rect 45585 687067 45601 687101
rect 45669 687067 45685 687101
rect 45743 687067 45759 687101
rect 45827 687067 45843 687101
rect 45901 687067 45917 687101
rect 45985 687067 46001 687101
rect 44793 686999 44827 687061
rect 46127 686999 46161 687061
rect 44793 686965 44889 686999
rect 46065 686965 46161 686999
rect 43794 686758 43890 686792
rect 47056 686758 47152 686792
rect 43794 686696 43828 686758
rect 47118 686696 47152 686758
rect 43954 686656 43970 686690
rect 44138 686656 44154 686690
rect 44212 686656 44228 686690
rect 44396 686656 44412 686690
rect 44470 686656 44486 686690
rect 44654 686656 44670 686690
rect 44728 686656 44744 686690
rect 44912 686656 44928 686690
rect 44986 686656 45002 686690
rect 45170 686656 45186 686690
rect 45244 686656 45260 686690
rect 45428 686656 45444 686690
rect 45502 686656 45518 686690
rect 45686 686656 45702 686690
rect 45760 686656 45776 686690
rect 45944 686656 45960 686690
rect 46018 686656 46034 686690
rect 46202 686656 46218 686690
rect 46276 686656 46292 686690
rect 46460 686656 46476 686690
rect 46534 686656 46550 686690
rect 46718 686656 46734 686690
rect 46792 686656 46808 686690
rect 46976 686656 46992 686690
rect 43908 686606 43942 686622
rect 43908 685614 43942 685630
rect 44166 686606 44200 686622
rect 44166 685614 44200 685630
rect 44424 686606 44458 686622
rect 44424 685614 44458 685630
rect 44682 686606 44716 686622
rect 44682 685614 44716 685630
rect 44940 686606 44974 686622
rect 44940 685614 44974 685630
rect 45198 686606 45232 686622
rect 45198 685614 45232 685630
rect 45456 686606 45490 686622
rect 45456 685614 45490 685630
rect 45714 686606 45748 686622
rect 45714 685614 45748 685630
rect 45972 686606 46006 686622
rect 45972 685614 46006 685630
rect 46230 686606 46264 686622
rect 46230 685614 46264 685630
rect 46488 686606 46522 686622
rect 46488 685614 46522 685630
rect 46746 686606 46780 686622
rect 46746 685614 46780 685630
rect 47004 686606 47038 686622
rect 47004 685614 47038 685630
rect 43954 685546 43970 685580
rect 44138 685546 44154 685580
rect 44212 685546 44228 685580
rect 44396 685546 44412 685580
rect 44470 685546 44486 685580
rect 44654 685546 44670 685580
rect 44728 685546 44744 685580
rect 44912 685546 44928 685580
rect 44986 685546 45002 685580
rect 45170 685546 45186 685580
rect 45244 685546 45260 685580
rect 45428 685546 45444 685580
rect 45502 685546 45518 685580
rect 45686 685546 45702 685580
rect 45760 685546 45776 685580
rect 45944 685546 45960 685580
rect 46018 685546 46034 685580
rect 46202 685546 46218 685580
rect 46276 685546 46292 685580
rect 46460 685546 46476 685580
rect 46534 685546 46550 685580
rect 46718 685546 46734 685580
rect 46792 685546 46808 685580
rect 46976 685546 46992 685580
rect 43794 685478 43828 685540
rect 47118 685478 47152 685540
rect 43794 685444 43890 685478
rect 47056 685444 47152 685478
rect 43538 685238 43634 685272
rect 47316 685238 47412 685272
rect 43538 685176 43572 685238
rect 47378 685176 47412 685238
rect 43698 685136 43714 685170
rect 43882 685136 43898 685170
rect 43956 685136 43972 685170
rect 44140 685136 44156 685170
rect 44214 685136 44230 685170
rect 44398 685136 44414 685170
rect 44472 685136 44488 685170
rect 44656 685136 44672 685170
rect 44730 685136 44746 685170
rect 44914 685136 44930 685170
rect 44988 685136 45004 685170
rect 45172 685136 45188 685170
rect 45246 685136 45262 685170
rect 45430 685136 45446 685170
rect 45504 685136 45520 685170
rect 45688 685136 45704 685170
rect 45762 685136 45778 685170
rect 45946 685136 45962 685170
rect 46020 685136 46036 685170
rect 46204 685136 46220 685170
rect 46278 685136 46294 685170
rect 46462 685136 46478 685170
rect 46536 685136 46552 685170
rect 46720 685136 46736 685170
rect 46794 685136 46810 685170
rect 46978 685136 46994 685170
rect 47052 685136 47068 685170
rect 47236 685136 47252 685170
rect 43652 685086 43686 685102
rect 43652 684094 43686 684110
rect 43910 685086 43944 685102
rect 43910 684094 43944 684110
rect 44168 685086 44202 685102
rect 44168 684094 44202 684110
rect 44426 685086 44460 685102
rect 44426 684094 44460 684110
rect 44684 685086 44718 685102
rect 44684 684094 44718 684110
rect 44942 685086 44976 685102
rect 44942 684094 44976 684110
rect 45200 685086 45234 685102
rect 45200 684094 45234 684110
rect 45458 685086 45492 685102
rect 45458 684094 45492 684110
rect 45716 685086 45750 685102
rect 45716 684094 45750 684110
rect 45974 685086 46008 685102
rect 45974 684094 46008 684110
rect 46232 685086 46266 685102
rect 46232 684094 46266 684110
rect 46490 685086 46524 685102
rect 46490 684094 46524 684110
rect 46748 685086 46782 685102
rect 46748 684094 46782 684110
rect 47006 685086 47040 685102
rect 47006 684094 47040 684110
rect 47264 685086 47298 685102
rect 47264 684094 47298 684110
rect 43698 684026 43714 684060
rect 43882 684026 43898 684060
rect 43956 684026 43972 684060
rect 44140 684026 44156 684060
rect 44214 684026 44230 684060
rect 44398 684026 44414 684060
rect 44472 684026 44488 684060
rect 44656 684026 44672 684060
rect 44730 684026 44746 684060
rect 44914 684026 44930 684060
rect 44988 684026 45004 684060
rect 45172 684026 45188 684060
rect 45246 684026 45262 684060
rect 45430 684026 45446 684060
rect 45504 684026 45520 684060
rect 45688 684026 45704 684060
rect 45762 684026 45778 684060
rect 45946 684026 45962 684060
rect 46020 684026 46036 684060
rect 46204 684026 46220 684060
rect 46278 684026 46294 684060
rect 46462 684026 46478 684060
rect 46536 684026 46552 684060
rect 46720 684026 46736 684060
rect 46794 684026 46810 684060
rect 46978 684026 46994 684060
rect 47052 684026 47068 684060
rect 47236 684026 47252 684060
rect 43538 683958 43572 684020
rect 47378 683958 47412 684020
rect 43538 683924 43634 683958
rect 47316 683924 47412 683958
rect 41696 682950 41792 682984
rect 49146 682950 49242 682984
rect 41696 682888 41730 682950
rect 49208 682888 49242 682950
rect 41875 682836 41891 682870
rect 42867 682836 42883 682870
rect 43111 682836 43127 682870
rect 44103 682836 44119 682870
rect 44347 682836 44363 682870
rect 45339 682836 45355 682870
rect 45583 682836 45599 682870
rect 46575 682836 46591 682870
rect 46819 682836 46835 682870
rect 47811 682836 47827 682870
rect 48055 682836 48071 682870
rect 49047 682836 49063 682870
rect 41798 682808 41832 682824
rect 41798 682624 41832 682640
rect 42926 682808 42960 682824
rect 42926 682624 42960 682640
rect 43034 682808 43068 682824
rect 43034 682624 43068 682640
rect 44162 682808 44196 682824
rect 44162 682624 44196 682640
rect 44270 682808 44304 682824
rect 44270 682624 44304 682640
rect 45398 682808 45432 682824
rect 45398 682624 45432 682640
rect 45506 682808 45540 682824
rect 45506 682624 45540 682640
rect 46634 682808 46668 682824
rect 46634 682624 46668 682640
rect 46742 682808 46776 682824
rect 46742 682624 46776 682640
rect 47870 682808 47904 682824
rect 47870 682624 47904 682640
rect 47978 682808 48012 682824
rect 47978 682624 48012 682640
rect 49106 682808 49140 682824
rect 49106 682624 49140 682640
rect 41875 682578 41891 682612
rect 42867 682578 42883 682612
rect 43111 682578 43127 682612
rect 44103 682578 44119 682612
rect 44347 682578 44363 682612
rect 45339 682578 45355 682612
rect 45583 682578 45599 682612
rect 46575 682578 46591 682612
rect 46819 682578 46835 682612
rect 47811 682578 47827 682612
rect 48055 682578 48071 682612
rect 49047 682578 49063 682612
rect 41696 682498 41730 682560
rect 49208 682498 49242 682560
rect 41696 682464 41792 682498
rect 49146 682464 49242 682498
rect 41696 682360 41792 682394
rect 49146 682360 49242 682394
rect 41696 682298 41730 682360
rect 49208 682298 49242 682360
rect 41875 682246 41891 682280
rect 42867 682246 42883 682280
rect 43111 682246 43127 682280
rect 44103 682246 44119 682280
rect 44347 682246 44363 682280
rect 45339 682246 45355 682280
rect 45583 682246 45599 682280
rect 46575 682246 46591 682280
rect 46819 682246 46835 682280
rect 47811 682246 47827 682280
rect 48055 682246 48071 682280
rect 49047 682246 49063 682280
rect 41798 682218 41832 682234
rect 41798 682034 41832 682050
rect 42926 682218 42960 682234
rect 42926 682034 42960 682050
rect 43034 682218 43068 682234
rect 43034 682034 43068 682050
rect 44162 682218 44196 682234
rect 44162 682034 44196 682050
rect 44270 682218 44304 682234
rect 44270 682034 44304 682050
rect 45398 682218 45432 682234
rect 45398 682034 45432 682050
rect 45506 682218 45540 682234
rect 45506 682034 45540 682050
rect 46634 682218 46668 682234
rect 46634 682034 46668 682050
rect 46742 682218 46776 682234
rect 46742 682034 46776 682050
rect 47870 682218 47904 682234
rect 47870 682034 47904 682050
rect 47978 682218 48012 682234
rect 47978 682034 48012 682050
rect 49106 682218 49140 682234
rect 49106 682034 49140 682050
rect 41875 681988 41891 682022
rect 42867 681988 42883 682022
rect 43111 681988 43127 682022
rect 44103 681988 44119 682022
rect 44347 681988 44363 682022
rect 45339 681988 45355 682022
rect 45583 681988 45599 682022
rect 46575 681988 46591 682022
rect 46819 681988 46835 682022
rect 47811 681988 47827 682022
rect 48055 681988 48071 682022
rect 49047 681988 49063 682022
rect 41696 681908 41730 681970
rect 49208 681908 49242 681970
rect 41696 681874 41792 681908
rect 49146 681874 49242 681908
rect 44470 681570 44566 681604
rect 46376 681570 46472 681604
rect 44470 681508 44504 681570
rect 46438 681508 46472 681570
rect 44640 681456 44656 681490
rect 44882 681456 44898 681490
rect 45108 681456 45124 681490
rect 45350 681456 45366 681490
rect 45576 681456 45592 681490
rect 45818 681456 45834 681490
rect 46044 681456 46060 681490
rect 46286 681456 46302 681490
rect 44572 681428 44606 681444
rect 44572 681244 44606 681260
rect 44932 681428 44966 681444
rect 44932 681244 44966 681260
rect 45040 681428 45074 681444
rect 45040 681244 45074 681260
rect 45400 681428 45434 681444
rect 45400 681244 45434 681260
rect 45508 681428 45542 681444
rect 45508 681244 45542 681260
rect 45868 681428 45902 681444
rect 45868 681244 45902 681260
rect 45976 681428 46010 681444
rect 45976 681244 46010 681260
rect 46336 681428 46370 681444
rect 46336 681244 46370 681260
rect 44640 681198 44656 681232
rect 44882 681198 44898 681232
rect 45108 681198 45124 681232
rect 45350 681198 45366 681232
rect 45576 681198 45592 681232
rect 45818 681198 45834 681232
rect 46044 681198 46060 681232
rect 46286 681198 46302 681232
rect 44470 681118 44504 681180
rect 46438 681118 46472 681180
rect 44470 681084 44566 681118
rect 46376 681084 46472 681118
rect 44686 680945 44782 680968
rect 46156 680945 46252 680968
rect 44686 680883 44720 680945
rect 46218 680883 46252 680945
rect 44856 680831 44872 680865
rect 45348 680831 45364 680865
rect 45574 680831 45590 680865
rect 46066 680831 46082 680865
rect 44788 680803 44822 680819
rect 44788 680719 44822 680735
rect 45398 680803 45432 680819
rect 45398 680719 45432 680735
rect 45506 680803 45540 680819
rect 45506 680719 45540 680735
rect 46116 680803 46150 680819
rect 46116 680719 46150 680735
rect 44856 680673 44872 680707
rect 45348 680673 45364 680707
rect 45574 680673 45590 680707
rect 46066 680673 46082 680707
rect 44686 680593 44720 680655
rect 46218 680593 46252 680655
rect 44686 680559 44782 680593
rect 46156 680559 46252 680593
rect 41749 680420 41845 680454
rect 49091 680420 49187 680454
rect 41749 680358 41783 680420
rect 49153 680358 49187 680420
rect 41919 680306 41935 680340
rect 42911 680306 42927 680340
rect 43137 680306 43153 680340
rect 44129 680306 44145 680340
rect 44355 680306 44371 680340
rect 45347 680306 45363 680340
rect 45573 680306 45589 680340
rect 46565 680306 46581 680340
rect 46791 680306 46807 680340
rect 47783 680306 47799 680340
rect 48009 680306 48025 680340
rect 49001 680306 49017 680340
rect 41851 680278 41885 680294
rect 41851 680094 41885 680110
rect 42961 680278 42995 680294
rect 42961 680094 42995 680110
rect 43069 680278 43103 680294
rect 43069 680094 43103 680110
rect 44179 680278 44213 680294
rect 44179 680094 44213 680110
rect 44287 680278 44321 680294
rect 44287 680094 44321 680110
rect 45397 680278 45431 680294
rect 45397 680094 45431 680110
rect 45505 680278 45539 680294
rect 45505 680094 45539 680110
rect 46615 680278 46649 680294
rect 46615 680094 46649 680110
rect 46723 680278 46757 680294
rect 46723 680094 46757 680110
rect 47833 680278 47867 680294
rect 47833 680094 47867 680110
rect 47941 680278 47975 680294
rect 47941 680094 47975 680110
rect 49051 680278 49085 680294
rect 49051 680094 49085 680110
rect 41919 680048 41935 680082
rect 42911 680048 42927 680082
rect 43137 680048 43153 680082
rect 44129 680048 44145 680082
rect 44355 680048 44371 680082
rect 45347 680048 45363 680082
rect 45573 680048 45589 680082
rect 46565 680048 46581 680082
rect 46791 680048 46807 680082
rect 47783 680048 47799 680082
rect 48009 680048 48025 680082
rect 49001 680048 49017 680082
rect 41749 679968 41783 680030
rect 49153 679968 49187 680030
rect 41749 679934 41845 679968
rect 49091 679934 49187 679968
rect 42218 678658 42338 678674
rect 42218 678522 42338 678538
rect 48588 678658 48708 678674
rect 48588 678522 48708 678538
rect 42218 675658 42338 675674
rect 42218 675522 42338 675538
rect 48588 675658 48708 675674
rect 48588 675522 48708 675538
rect 42218 672658 42338 672674
rect 42218 672522 42338 672538
rect 48588 672658 48708 672674
rect 48588 672522 48708 672538
rect 42218 669658 42338 669674
rect 42218 669522 42338 669538
rect 48588 669658 48708 669674
rect 48588 669522 48708 669538
rect 42218 666658 42338 666674
rect 42218 666522 42338 666538
rect 48588 666658 48708 666674
rect 48588 666522 48708 666538
<< viali >>
rect 38519 694237 38916 695351
rect 40950 694237 41347 695351
rect 43843 694586 47099 694620
rect 38519 692777 38916 693891
rect 40950 692777 41347 693891
rect 42356 694484 42424 694518
rect 42514 694484 42582 694518
rect 42672 694484 42740 694518
rect 42830 694484 42898 694518
rect 42988 694484 43056 694518
rect 43146 694484 43214 694518
rect 43304 694484 43372 694518
rect 43462 694484 43530 694518
rect 43620 694484 43688 694518
rect 43778 694484 43846 694518
rect 43936 694484 44004 694518
rect 44094 694484 44162 694518
rect 44252 694484 44320 694518
rect 44410 694484 44478 694518
rect 44568 694484 44636 694518
rect 44726 694484 44794 694518
rect 44884 694484 44952 694518
rect 45042 694484 45110 694518
rect 45200 694484 45268 694518
rect 45358 694484 45426 694518
rect 45516 694484 45584 694518
rect 45674 694484 45742 694518
rect 45832 694484 45900 694518
rect 45990 694484 46058 694518
rect 46148 694484 46216 694518
rect 46306 694484 46374 694518
rect 46464 694484 46532 694518
rect 46622 694484 46690 694518
rect 46780 694484 46848 694518
rect 46938 694484 47006 694518
rect 47096 694484 47164 694518
rect 47254 694484 47322 694518
rect 47412 694484 47480 694518
rect 47570 694484 47638 694518
rect 47728 694484 47796 694518
rect 47886 694484 47954 694518
rect 48044 694484 48112 694518
rect 48202 694484 48270 694518
rect 48360 694484 48428 694518
rect 48518 694484 48586 694518
rect 42294 693449 42328 694425
rect 42452 693449 42486 694425
rect 42610 693449 42644 694425
rect 42768 693449 42802 694425
rect 42926 693449 42960 694425
rect 43084 693449 43118 694425
rect 43242 693449 43276 694425
rect 43400 693449 43434 694425
rect 43558 693449 43592 694425
rect 43716 693449 43750 694425
rect 43874 693449 43908 694425
rect 44032 693449 44066 694425
rect 44190 693449 44224 694425
rect 44348 693449 44382 694425
rect 44506 693449 44540 694425
rect 44664 693449 44698 694425
rect 44822 693449 44856 694425
rect 44980 693449 45014 694425
rect 45138 693449 45172 694425
rect 45296 693449 45330 694425
rect 45454 693449 45488 694425
rect 45612 693449 45646 694425
rect 45770 693449 45804 694425
rect 45928 693449 45962 694425
rect 46086 693449 46120 694425
rect 46244 693449 46278 694425
rect 46402 693449 46436 694425
rect 46560 693449 46594 694425
rect 46718 693449 46752 694425
rect 46876 693449 46910 694425
rect 47034 693449 47068 694425
rect 47192 693449 47226 694425
rect 47350 693449 47384 694425
rect 47508 693449 47542 694425
rect 47666 693449 47700 694425
rect 47824 693449 47858 694425
rect 47982 693449 48016 694425
rect 48140 693449 48174 694425
rect 48298 693449 48332 694425
rect 48456 693449 48490 694425
rect 48614 693449 48648 694425
rect 42356 693356 42424 693390
rect 42514 693356 42582 693390
rect 42672 693356 42740 693390
rect 42830 693356 42898 693390
rect 42988 693356 43056 693390
rect 43146 693356 43214 693390
rect 43304 693356 43372 693390
rect 43462 693356 43530 693390
rect 43620 693356 43688 693390
rect 43778 693356 43846 693390
rect 43936 693356 44004 693390
rect 44094 693356 44162 693390
rect 44252 693356 44320 693390
rect 44410 693356 44478 693390
rect 44568 693356 44636 693390
rect 44726 693356 44794 693390
rect 44884 693356 44952 693390
rect 45042 693356 45110 693390
rect 45200 693356 45268 693390
rect 45358 693356 45426 693390
rect 45516 693356 45584 693390
rect 45674 693356 45742 693390
rect 45832 693356 45900 693390
rect 45990 693356 46058 693390
rect 46148 693356 46216 693390
rect 46306 693356 46374 693390
rect 46464 693356 46532 693390
rect 46622 693356 46690 693390
rect 46780 693356 46848 693390
rect 46938 693356 47006 693390
rect 47096 693356 47164 693390
rect 47254 693356 47322 693390
rect 47412 693356 47480 693390
rect 47570 693356 47638 693390
rect 47728 693356 47796 693390
rect 47886 693356 47954 693390
rect 48044 693356 48112 693390
rect 48202 693356 48270 693390
rect 48360 693356 48428 693390
rect 48518 693356 48586 693390
rect 49589 694237 49986 695351
rect 52020 694237 52417 695351
rect 43843 693254 47099 693288
rect 39578 692665 39758 692698
rect 39998 692665 40178 692698
rect 39578 692631 39758 692665
rect 39998 692631 40178 692665
rect 44594 692916 46350 692950
rect 39578 692598 39758 692631
rect 39998 692598 40178 692631
rect 43858 692814 43926 692848
rect 44016 692814 44084 692848
rect 44174 692814 44242 692848
rect 44332 692814 44400 692848
rect 44490 692814 44558 692848
rect 44648 692814 44716 692848
rect 44806 692814 44874 692848
rect 44964 692814 45032 692848
rect 45122 692814 45190 692848
rect 45280 692814 45348 692848
rect 45438 692814 45506 692848
rect 45596 692814 45664 692848
rect 45754 692814 45822 692848
rect 45912 692814 45980 692848
rect 46070 692814 46138 692848
rect 46228 692814 46296 692848
rect 46386 692814 46454 692848
rect 46544 692814 46612 692848
rect 46702 692814 46770 692848
rect 46860 692814 46928 692848
rect 47018 692814 47086 692848
rect 43796 691779 43830 692755
rect 43954 691779 43988 692755
rect 44112 691779 44146 692755
rect 44270 691779 44304 692755
rect 44428 691779 44462 692755
rect 44586 691779 44620 692755
rect 44744 691779 44778 692755
rect 44902 691779 44936 692755
rect 45060 691779 45094 692755
rect 45218 691779 45252 692755
rect 45376 691779 45410 692755
rect 45534 691779 45568 692755
rect 45692 691779 45726 692755
rect 45850 691779 45884 692755
rect 46008 691779 46042 692755
rect 46166 691779 46200 692755
rect 46324 691779 46358 692755
rect 46482 691779 46516 692755
rect 46640 691779 46674 692755
rect 46798 691779 46832 692755
rect 46956 691779 46990 692755
rect 47114 691779 47148 692755
rect 43858 691686 43926 691720
rect 44016 691686 44084 691720
rect 44174 691686 44242 691720
rect 44332 691686 44400 691720
rect 44490 691686 44558 691720
rect 44648 691686 44716 691720
rect 44806 691686 44874 691720
rect 44964 691686 45032 691720
rect 45122 691686 45190 691720
rect 45280 691686 45348 691720
rect 45438 691686 45506 691720
rect 45596 691686 45664 691720
rect 45754 691686 45822 691720
rect 45912 691686 45980 691720
rect 46070 691686 46138 691720
rect 46228 691686 46296 691720
rect 46386 691686 46454 691720
rect 46544 691686 46612 691720
rect 46702 691686 46770 691720
rect 46860 691686 46928 691720
rect 47018 691686 47086 691720
rect 49589 692777 49986 693891
rect 52020 692777 52417 693891
rect 50828 692665 51008 692698
rect 51248 692665 51428 692698
rect 50828 692631 51008 692665
rect 51248 692631 51428 692665
rect 50828 692598 51008 692631
rect 51248 692598 51428 692631
rect 44448 691584 45018 691618
rect 45918 691584 46488 691618
rect 44448 691410 45018 691584
rect 45918 691410 46488 691584
rect 44448 691378 45018 691410
rect 45918 691378 46488 691410
rect 43858 691274 43926 691308
rect 44016 691274 44084 691308
rect 44174 691274 44242 691308
rect 44332 691274 44400 691308
rect 44490 691274 44558 691308
rect 44648 691274 44716 691308
rect 44806 691274 44874 691308
rect 44964 691274 45032 691308
rect 45122 691274 45190 691308
rect 45280 691274 45348 691308
rect 45438 691274 45506 691308
rect 45596 691274 45664 691308
rect 45754 691274 45822 691308
rect 45912 691274 45980 691308
rect 46070 691274 46138 691308
rect 46228 691274 46296 691308
rect 46386 691274 46454 691308
rect 46544 691274 46612 691308
rect 46702 691274 46770 691308
rect 46860 691274 46928 691308
rect 47018 691274 47086 691308
rect 43796 690239 43830 691215
rect 43954 690239 43988 691215
rect 44112 690239 44146 691215
rect 44270 690239 44304 691215
rect 44428 690239 44462 691215
rect 44586 690239 44620 691215
rect 44744 690239 44778 691215
rect 44902 690239 44936 691215
rect 45060 690239 45094 691215
rect 45218 690239 45252 691215
rect 45376 690239 45410 691215
rect 45534 690239 45568 691215
rect 45692 690239 45726 691215
rect 45850 690239 45884 691215
rect 46008 690239 46042 691215
rect 46166 690239 46200 691215
rect 46324 690239 46358 691215
rect 46482 690239 46516 691215
rect 46640 690239 46674 691215
rect 46798 690239 46832 691215
rect 46956 690239 46990 691215
rect 47114 690239 47148 691215
rect 43858 690146 43926 690180
rect 44016 690146 44084 690180
rect 44174 690146 44242 690180
rect 44332 690146 44400 690180
rect 44490 690146 44558 690180
rect 44648 690146 44716 690180
rect 44806 690146 44874 690180
rect 44964 690146 45032 690180
rect 45122 690146 45190 690180
rect 45280 690146 45348 690180
rect 45438 690146 45506 690180
rect 45596 690146 45664 690180
rect 45754 690146 45822 690180
rect 45912 690146 45980 690180
rect 46070 690146 46138 690180
rect 46228 690146 46296 690180
rect 46386 690146 46454 690180
rect 46544 690146 46612 690180
rect 46702 690146 46770 690180
rect 46860 690146 46928 690180
rect 47018 690146 47086 690180
rect 45152 689799 45802 689833
rect 44969 689697 45037 689731
rect 45127 689697 45195 689731
rect 45285 689697 45353 689731
rect 45443 689697 45511 689731
rect 45601 689697 45669 689731
rect 45759 689697 45827 689731
rect 45917 689697 45985 689731
rect 44907 688671 44941 689647
rect 45065 688671 45099 689647
rect 45223 688671 45257 689647
rect 45381 688671 45415 689647
rect 45539 688671 45573 689647
rect 45697 688671 45731 689647
rect 45855 688671 45889 689647
rect 46013 688671 46047 689647
rect 44969 688587 45037 688621
rect 45127 688587 45195 688621
rect 45285 688587 45353 688621
rect 45443 688587 45511 688621
rect 45601 688587 45669 688621
rect 45759 688587 45827 688621
rect 45917 688587 45985 688621
rect 45152 688485 45802 688519
rect 45152 688279 45802 688313
rect 44969 688177 45037 688211
rect 45127 688177 45195 688211
rect 45285 688177 45353 688211
rect 45443 688177 45511 688211
rect 45601 688177 45669 688211
rect 45759 688177 45827 688211
rect 45917 688177 45985 688211
rect 44907 687151 44941 688127
rect 45065 687151 45099 688127
rect 45223 687151 45257 688127
rect 45381 687151 45415 688127
rect 45539 687151 45573 688127
rect 45697 687151 45731 688127
rect 45855 687151 45889 688127
rect 46013 687151 46047 688127
rect 44969 687067 45037 687101
rect 45127 687067 45195 687101
rect 45285 687067 45353 687101
rect 45443 687067 45511 687101
rect 45601 687067 45669 687101
rect 45759 687067 45827 687101
rect 45917 687067 45985 687101
rect 45152 686965 45802 686999
rect 44651 686758 46295 686792
rect 43970 686656 44138 686690
rect 44228 686656 44396 686690
rect 44486 686656 44654 686690
rect 44744 686656 44912 686690
rect 45002 686656 45170 686690
rect 45260 686656 45428 686690
rect 45518 686656 45686 686690
rect 45776 686656 45944 686690
rect 46034 686656 46202 686690
rect 46292 686656 46460 686690
rect 46550 686656 46718 686690
rect 46808 686656 46976 686690
rect 43908 685630 43942 686606
rect 44166 685630 44200 686606
rect 44424 685630 44458 686606
rect 44682 685630 44716 686606
rect 44940 685630 44974 686606
rect 45198 685630 45232 686606
rect 45456 685630 45490 686606
rect 45714 685630 45748 686606
rect 45972 685630 46006 686606
rect 46230 685630 46264 686606
rect 46488 685630 46522 686606
rect 46746 685630 46780 686606
rect 47004 685630 47038 686606
rect 43970 685546 44138 685580
rect 44228 685546 44396 685580
rect 44486 685546 44654 685580
rect 44744 685546 44912 685580
rect 45002 685546 45170 685580
rect 45260 685546 45428 685580
rect 45518 685546 45686 685580
rect 45776 685546 45944 685580
rect 46034 685546 46202 685580
rect 46292 685546 46460 685580
rect 46550 685546 46718 685580
rect 46808 685546 46976 685580
rect 44651 685444 46295 685478
rect 44524 685238 46426 685272
rect 43714 685136 43882 685170
rect 43972 685136 44140 685170
rect 44230 685136 44398 685170
rect 44488 685136 44656 685170
rect 44746 685136 44914 685170
rect 45004 685136 45172 685170
rect 45262 685136 45430 685170
rect 45520 685136 45688 685170
rect 45778 685136 45946 685170
rect 46036 685136 46204 685170
rect 46294 685136 46462 685170
rect 46552 685136 46720 685170
rect 46810 685136 46978 685170
rect 47068 685136 47236 685170
rect 43652 684110 43686 685086
rect 43910 684110 43944 685086
rect 44168 684110 44202 685086
rect 44426 684110 44460 685086
rect 44684 684110 44718 685086
rect 44942 684110 44976 685086
rect 45200 684110 45234 685086
rect 45458 684110 45492 685086
rect 45716 684110 45750 685086
rect 45974 684110 46008 685086
rect 46232 684110 46266 685086
rect 46490 684110 46524 685086
rect 46748 684110 46782 685086
rect 47006 684110 47040 685086
rect 47264 684110 47298 685086
rect 43714 684026 43882 684060
rect 43972 684026 44140 684060
rect 44230 684026 44398 684060
rect 44488 684026 44656 684060
rect 44746 684026 44914 684060
rect 45004 684026 45172 684060
rect 45262 684026 45430 684060
rect 45520 684026 45688 684060
rect 45778 684026 45946 684060
rect 46036 684026 46204 684060
rect 46294 684026 46462 684060
rect 46552 684026 46720 684060
rect 46810 684026 46978 684060
rect 47068 684026 47236 684060
rect 44524 683924 46426 683958
rect 42308 682984 42468 683078
rect 43308 682984 43468 683078
rect 44788 682984 44948 683078
rect 46008 682984 46168 683078
rect 47468 682984 47628 683078
rect 48528 682984 48688 683078
rect 42308 682950 42468 682984
rect 43308 682950 43468 682984
rect 44788 682950 44948 682984
rect 46008 682950 46168 682984
rect 47468 682950 47628 682984
rect 48528 682950 48688 682984
rect 42308 682918 42468 682950
rect 43308 682918 43468 682950
rect 44788 682918 44948 682950
rect 46008 682918 46168 682950
rect 47468 682918 47628 682950
rect 48528 682918 48688 682950
rect 41891 682836 42867 682870
rect 43127 682836 44103 682870
rect 44363 682836 45339 682870
rect 45599 682836 46575 682870
rect 46835 682836 47811 682870
rect 48071 682836 49047 682870
rect 41798 682640 41832 682808
rect 42926 682640 42960 682808
rect 43034 682640 43068 682808
rect 44162 682640 44196 682808
rect 44270 682640 44304 682808
rect 45398 682640 45432 682808
rect 45506 682640 45540 682808
rect 46634 682640 46668 682808
rect 46742 682640 46776 682808
rect 47870 682640 47904 682808
rect 47978 682640 48012 682808
rect 49106 682640 49140 682808
rect 41891 682578 42867 682612
rect 43127 682578 44103 682612
rect 44363 682578 45339 682612
rect 45599 682578 46575 682612
rect 46835 682578 47811 682612
rect 48071 682578 49047 682612
rect 42308 682464 42468 682498
rect 43308 682464 43468 682498
rect 44788 682464 44948 682498
rect 46008 682464 46168 682498
rect 47468 682464 47628 682498
rect 48528 682464 48688 682498
rect 42308 682394 42468 682464
rect 43308 682394 43468 682464
rect 44788 682394 44948 682464
rect 46008 682394 46168 682464
rect 47468 682394 47628 682464
rect 48528 682394 48688 682464
rect 42308 682360 42468 682394
rect 43308 682360 43468 682394
rect 44788 682360 44948 682394
rect 46008 682360 46168 682394
rect 47468 682360 47628 682394
rect 48528 682360 48688 682394
rect 42308 682338 42468 682360
rect 43308 682338 43468 682360
rect 44788 682338 44948 682360
rect 46008 682338 46168 682360
rect 47468 682338 47628 682360
rect 48528 682338 48688 682360
rect 41891 682246 42867 682280
rect 43127 682246 44103 682280
rect 44363 682246 45339 682280
rect 45599 682246 46575 682280
rect 46835 682246 47811 682280
rect 48071 682246 49047 682280
rect 41798 682050 41832 682218
rect 42926 682050 42960 682218
rect 43034 682050 43068 682218
rect 44162 682050 44196 682218
rect 44270 682050 44304 682218
rect 45398 682050 45432 682218
rect 45506 682050 45540 682218
rect 46634 682050 46668 682218
rect 46742 682050 46776 682218
rect 47870 682050 47904 682218
rect 47978 682050 48012 682218
rect 49106 682050 49140 682218
rect 41891 681988 42867 682022
rect 43127 681988 44103 682022
rect 44363 681988 45339 682022
rect 45599 681988 46575 682022
rect 46835 681988 47811 682022
rect 48071 681988 49047 682022
rect 44656 681456 44882 681490
rect 45124 681456 45350 681490
rect 45592 681456 45818 681490
rect 46060 681456 46286 681490
rect 44572 681260 44606 681428
rect 44932 681260 44966 681428
rect 45040 681260 45074 681428
rect 45400 681260 45434 681428
rect 45508 681260 45542 681428
rect 45868 681260 45902 681428
rect 45976 681260 46010 681428
rect 46336 681260 46370 681428
rect 44656 681198 44882 681232
rect 45124 681198 45350 681232
rect 45592 681198 45818 681232
rect 46060 681198 46286 681232
rect 44598 681084 44818 681118
rect 45148 681084 45368 681118
rect 45568 681084 45788 681118
rect 46088 681084 46308 681118
rect 44598 680979 44818 681084
rect 45148 680979 45368 681084
rect 45568 680979 45788 681084
rect 46088 680979 46308 681084
rect 44598 680968 44782 680979
rect 44782 680968 44818 680979
rect 45148 680968 45368 680979
rect 45568 680968 45788 680979
rect 46088 680968 46156 680979
rect 46156 680968 46308 680979
rect 44872 680831 45348 680865
rect 45590 680831 46066 680865
rect 44788 680735 44822 680803
rect 45398 680735 45432 680803
rect 45506 680735 45540 680803
rect 46116 680735 46150 680803
rect 44872 680673 45348 680707
rect 45590 680673 46066 680707
rect 42368 680454 42548 680568
rect 43368 680454 43548 680568
rect 45158 680559 45338 680568
rect 45598 680559 45778 680568
rect 44438 680454 44618 680558
rect 45158 680454 45338 680559
rect 45598 680454 45778 680559
rect 46368 680454 46548 680568
rect 47348 680454 47528 680558
rect 48488 680454 48668 680558
rect 42368 680438 42548 680454
rect 43368 680438 43548 680454
rect 44438 680428 44618 680454
rect 45158 680438 45338 680454
rect 45598 680438 45778 680454
rect 46368 680438 46548 680454
rect 47348 680428 47528 680454
rect 48488 680428 48668 680454
rect 41935 680306 42911 680340
rect 43153 680306 44129 680340
rect 44371 680306 45347 680340
rect 45589 680306 46565 680340
rect 46807 680306 47783 680340
rect 48025 680306 49001 680340
rect 41851 680110 41885 680278
rect 42961 680110 42995 680278
rect 43069 680110 43103 680278
rect 44179 680110 44213 680278
rect 44287 680110 44321 680278
rect 45397 680110 45431 680278
rect 45505 680110 45539 680278
rect 46615 680110 46649 680278
rect 46723 680110 46757 680278
rect 47833 680110 47867 680278
rect 47941 680110 47975 680278
rect 49051 680110 49085 680278
rect 41935 680048 42911 680082
rect 43153 680048 44129 680082
rect 44371 680048 45347 680082
rect 45589 680048 46565 680082
rect 46807 680048 47783 680082
rect 48025 680048 49001 680082
rect 42641 679193 43755 679590
rect 44151 679193 45265 679590
rect 45661 679187 46775 679584
rect 47181 679187 48295 679584
rect 42218 678538 42338 678658
rect 48588 678538 48708 678658
rect 42218 675538 42338 675658
rect 48588 675538 48708 675658
rect 42218 672538 42338 672658
rect 48588 672538 48708 672658
rect 42218 669538 42338 669658
rect 48588 669538 48708 669658
rect 42218 666538 42338 666658
rect 48588 666538 48708 666658
rect 42641 664962 43755 665359
rect 44151 664962 45265 665359
rect 45661 664956 46775 665353
rect 47181 664956 48295 665353
<< metal1 >>
rect 38498 695351 38938 695368
rect 38498 694237 38519 695351
rect 38916 694237 38938 695351
rect 38498 694178 38938 694237
rect 37608 694158 38938 694178
rect 37608 694088 37738 694158
rect 37808 694088 38938 694158
rect 37608 694048 38938 694088
rect 37608 693978 37628 694048
rect 37698 693978 38938 694048
rect 37608 693958 38938 693978
rect 38498 693891 38938 693958
rect 38498 692777 38519 693891
rect 38916 692777 38938 693891
rect 38498 692758 38938 692777
rect 40938 695351 41368 695368
rect 40938 694237 40950 695351
rect 41347 694237 41368 695351
rect 49568 695351 50008 695378
rect 44768 694878 46148 694928
rect 44768 694626 44798 694878
rect 43831 694620 44798 694626
rect 45068 694620 45848 694878
rect 46118 694626 46148 694878
rect 46118 694620 47111 694626
rect 43831 694586 43843 694620
rect 47099 694586 47111 694620
rect 43831 694580 47111 694586
rect 40938 694098 41368 694237
rect 42138 694518 48798 694528
rect 42138 694484 42356 694518
rect 42424 694484 42514 694518
rect 42582 694484 42672 694518
rect 42740 694484 42830 694518
rect 42898 694484 42988 694518
rect 43056 694484 43146 694518
rect 43214 694484 43304 694518
rect 43372 694484 43462 694518
rect 43530 694484 43620 694518
rect 43688 694484 43778 694518
rect 43846 694484 43936 694518
rect 44004 694484 44094 694518
rect 44162 694484 44252 694518
rect 44320 694484 44410 694518
rect 44478 694484 44568 694518
rect 44636 694484 44726 694518
rect 44794 694484 44884 694518
rect 44952 694484 45042 694518
rect 45110 694484 45200 694518
rect 45268 694484 45358 694518
rect 45426 694484 45516 694518
rect 45584 694484 45674 694518
rect 45742 694484 45832 694518
rect 45900 694484 45990 694518
rect 46058 694484 46148 694518
rect 46216 694484 46306 694518
rect 46374 694484 46464 694518
rect 46532 694484 46622 694518
rect 46690 694484 46780 694518
rect 46848 694484 46938 694518
rect 47006 694484 47096 694518
rect 47164 694484 47254 694518
rect 47322 694484 47412 694518
rect 47480 694484 47570 694518
rect 47638 694484 47728 694518
rect 47796 694484 47886 694518
rect 47954 694484 48044 694518
rect 48112 694484 48202 694518
rect 48270 694484 48360 694518
rect 48428 694484 48518 694518
rect 48586 694484 48798 694518
rect 42138 694478 48798 694484
rect 42138 694098 42218 694478
rect 42288 694425 42334 694437
rect 42288 694398 42294 694425
rect 42328 694398 42334 694425
rect 42446 694425 42492 694437
rect 42268 694328 42278 694398
rect 42348 694328 42358 694398
rect 42288 694158 42294 694328
rect 42328 694158 42334 694328
rect 40938 693891 42218 694098
rect 42268 694088 42278 694158
rect 42348 694088 42358 694158
rect 40938 692777 40950 693891
rect 41347 693808 42218 693891
rect 41347 692777 41368 693808
rect 42138 693398 42218 693808
rect 42288 693449 42294 694088
rect 42328 693449 42334 694088
rect 42446 693788 42452 694425
rect 42486 693788 42492 694425
rect 42604 694425 42650 694437
rect 42604 694398 42610 694425
rect 42644 694398 42650 694425
rect 42762 694425 42808 694437
rect 42578 694328 42588 694398
rect 42658 694328 42668 694398
rect 42604 694158 42610 694328
rect 42644 694158 42650 694328
rect 42578 694088 42588 694158
rect 42658 694088 42668 694158
rect 42418 693718 42428 693788
rect 42498 693718 42508 693788
rect 42446 693548 42452 693718
rect 42486 693548 42492 693718
rect 42418 693478 42428 693548
rect 42498 693478 42508 693548
rect 42288 693437 42334 693449
rect 42446 693449 42452 693478
rect 42486 693449 42492 693478
rect 42446 693437 42492 693449
rect 42604 693449 42610 694088
rect 42644 693449 42650 694088
rect 42762 693788 42768 694425
rect 42802 693788 42808 694425
rect 42920 694425 42966 694437
rect 42920 694398 42926 694425
rect 42960 694398 42966 694425
rect 43078 694425 43124 694437
rect 42898 694328 42908 694398
rect 42978 694328 42988 694398
rect 42920 694158 42926 694328
rect 42960 694158 42966 694328
rect 42898 694088 42908 694158
rect 42978 694088 42988 694158
rect 42738 693718 42748 693788
rect 42818 693718 42828 693788
rect 42762 693548 42768 693718
rect 42802 693548 42808 693718
rect 42738 693478 42748 693548
rect 42818 693478 42828 693548
rect 42604 693437 42650 693449
rect 42762 693449 42768 693478
rect 42802 693449 42808 693478
rect 42762 693437 42808 693449
rect 42920 693449 42926 694088
rect 42960 693449 42966 694088
rect 43078 693788 43084 694425
rect 43118 693788 43124 694425
rect 43236 694425 43282 694437
rect 43236 694398 43242 694425
rect 43276 694398 43282 694425
rect 43394 694425 43440 694437
rect 43218 694328 43228 694398
rect 43298 694328 43308 694398
rect 43236 694158 43242 694328
rect 43276 694158 43282 694328
rect 43218 694088 43228 694158
rect 43298 694088 43308 694158
rect 43058 693718 43068 693788
rect 43138 693718 43148 693788
rect 43078 693548 43084 693718
rect 43118 693548 43124 693718
rect 43058 693478 43068 693548
rect 43138 693478 43148 693548
rect 42920 693437 42966 693449
rect 43078 693449 43084 693478
rect 43118 693449 43124 693478
rect 43078 693437 43124 693449
rect 43236 693449 43242 694088
rect 43276 693449 43282 694088
rect 43394 693788 43400 694425
rect 43434 693788 43440 694425
rect 43552 694425 43598 694437
rect 43552 694398 43558 694425
rect 43592 694398 43598 694425
rect 43710 694425 43756 694437
rect 43528 694328 43538 694398
rect 43608 694328 43618 694398
rect 43552 694158 43558 694328
rect 43592 694158 43598 694328
rect 43528 694088 43538 694158
rect 43608 694088 43618 694158
rect 43368 693718 43378 693788
rect 43448 693718 43458 693788
rect 43394 693548 43400 693718
rect 43434 693548 43440 693718
rect 43368 693478 43378 693548
rect 43448 693478 43458 693548
rect 43236 693437 43282 693449
rect 43394 693449 43400 693478
rect 43434 693449 43440 693478
rect 43394 693437 43440 693449
rect 43552 693449 43558 694088
rect 43592 693449 43598 694088
rect 43710 693788 43716 694425
rect 43750 693788 43756 694425
rect 43868 694425 43914 694437
rect 43868 694398 43874 694425
rect 43908 694398 43914 694425
rect 44026 694425 44072 694437
rect 43848 694328 43858 694398
rect 43928 694328 43938 694398
rect 43868 694158 43874 694328
rect 43908 694158 43914 694328
rect 43848 694088 43858 694158
rect 43928 694088 43938 694158
rect 43688 693718 43698 693788
rect 43768 693718 43778 693788
rect 43710 693548 43716 693718
rect 43750 693548 43756 693718
rect 43688 693478 43698 693548
rect 43768 693478 43778 693548
rect 43552 693437 43598 693449
rect 43710 693449 43716 693478
rect 43750 693449 43756 693478
rect 43710 693437 43756 693449
rect 43868 693449 43874 694088
rect 43908 693449 43914 694088
rect 44026 693788 44032 694425
rect 44066 693788 44072 694425
rect 44184 694425 44230 694437
rect 44184 694398 44190 694425
rect 44224 694398 44230 694425
rect 44342 694425 44388 694437
rect 44158 694328 44168 694398
rect 44238 694328 44248 694398
rect 44184 694158 44190 694328
rect 44224 694158 44230 694328
rect 44158 694088 44168 694158
rect 44238 694088 44248 694158
rect 44008 693718 44018 693788
rect 44088 693718 44098 693788
rect 44026 693548 44032 693718
rect 44066 693548 44072 693718
rect 44008 693478 44018 693548
rect 44088 693478 44098 693548
rect 43868 693437 43914 693449
rect 44026 693449 44032 693478
rect 44066 693449 44072 693478
rect 44026 693437 44072 693449
rect 44184 693449 44190 694088
rect 44224 693449 44230 694088
rect 44342 693788 44348 694425
rect 44382 693788 44388 694425
rect 44500 694425 44546 694437
rect 44500 694398 44506 694425
rect 44540 694398 44546 694425
rect 44658 694425 44704 694437
rect 44478 694328 44488 694398
rect 44558 694328 44568 694398
rect 44500 694158 44506 694328
rect 44540 694158 44546 694328
rect 44478 694088 44488 694158
rect 44558 694088 44568 694158
rect 44318 693718 44328 693788
rect 44398 693718 44408 693788
rect 44342 693548 44348 693718
rect 44382 693548 44388 693718
rect 44318 693478 44328 693548
rect 44398 693478 44408 693548
rect 44184 693437 44230 693449
rect 44342 693449 44348 693478
rect 44382 693449 44388 693478
rect 44342 693437 44388 693449
rect 44500 693449 44506 694088
rect 44540 693449 44546 694088
rect 44658 693788 44664 694425
rect 44698 693788 44704 694425
rect 44816 694425 44862 694437
rect 44816 694398 44822 694425
rect 44856 694398 44862 694425
rect 44974 694425 45020 694437
rect 44798 694328 44808 694398
rect 44878 694328 44888 694398
rect 44816 694158 44822 694328
rect 44856 694158 44862 694328
rect 44798 694088 44808 694158
rect 44878 694088 44888 694158
rect 44638 693718 44648 693788
rect 44718 693718 44728 693788
rect 44658 693548 44664 693718
rect 44698 693548 44704 693718
rect 44638 693478 44648 693548
rect 44718 693478 44728 693548
rect 44500 693437 44546 693449
rect 44658 693449 44664 693478
rect 44698 693449 44704 693478
rect 44658 693437 44704 693449
rect 44816 693449 44822 694088
rect 44856 693449 44862 694088
rect 44974 693788 44980 694425
rect 45014 693788 45020 694425
rect 45132 694425 45178 694437
rect 45132 694398 45138 694425
rect 45172 694398 45178 694425
rect 45290 694425 45336 694437
rect 45108 694328 45118 694398
rect 45188 694328 45198 694398
rect 45132 694158 45138 694328
rect 45172 694158 45178 694328
rect 45108 694088 45118 694158
rect 45188 694088 45198 694158
rect 44948 693718 44958 693788
rect 45028 693718 45038 693788
rect 44974 693548 44980 693718
rect 45014 693548 45020 693718
rect 44948 693478 44958 693548
rect 45028 693478 45038 693548
rect 44816 693437 44862 693449
rect 44974 693449 44980 693478
rect 45014 693449 45020 693478
rect 44974 693437 45020 693449
rect 45132 693449 45138 694088
rect 45172 693449 45178 694088
rect 45290 693788 45296 694425
rect 45330 693788 45336 694425
rect 45448 694425 45494 694437
rect 45448 694398 45454 694425
rect 45488 694398 45494 694425
rect 45606 694425 45652 694437
rect 45428 694328 45438 694398
rect 45508 694328 45518 694398
rect 45448 694158 45454 694328
rect 45488 694158 45494 694328
rect 45428 694088 45438 694158
rect 45508 694088 45518 694158
rect 45268 693718 45278 693788
rect 45348 693718 45358 693788
rect 45290 693548 45296 693718
rect 45330 693548 45336 693718
rect 45268 693478 45278 693548
rect 45348 693478 45358 693548
rect 45132 693437 45178 693449
rect 45290 693449 45296 693478
rect 45330 693449 45336 693478
rect 45290 693437 45336 693449
rect 45448 693449 45454 694088
rect 45488 693449 45494 694088
rect 45606 693788 45612 694425
rect 45646 693788 45652 694425
rect 45764 694425 45810 694437
rect 45764 694398 45770 694425
rect 45804 694398 45810 694425
rect 45922 694425 45968 694437
rect 45738 694328 45748 694398
rect 45818 694328 45828 694398
rect 45764 694158 45770 694328
rect 45804 694158 45810 694328
rect 45738 694088 45748 694158
rect 45818 694088 45828 694158
rect 45588 693718 45598 693788
rect 45668 693718 45678 693788
rect 45606 693548 45612 693718
rect 45646 693548 45652 693718
rect 45588 693478 45598 693548
rect 45668 693478 45678 693548
rect 45448 693437 45494 693449
rect 45606 693449 45612 693478
rect 45646 693449 45652 693478
rect 45606 693437 45652 693449
rect 45764 693449 45770 694088
rect 45804 693449 45810 694088
rect 45922 693788 45928 694425
rect 45962 693788 45968 694425
rect 46080 694425 46126 694437
rect 46080 694398 46086 694425
rect 46120 694398 46126 694425
rect 46238 694425 46284 694437
rect 46058 694328 46068 694398
rect 46138 694328 46148 694398
rect 46080 694158 46086 694328
rect 46120 694158 46126 694328
rect 46058 694088 46068 694158
rect 46138 694088 46148 694158
rect 45898 693718 45908 693788
rect 45978 693718 45988 693788
rect 45922 693548 45928 693718
rect 45962 693548 45968 693718
rect 45898 693478 45908 693548
rect 45978 693478 45988 693548
rect 45764 693437 45810 693449
rect 45922 693449 45928 693478
rect 45962 693449 45968 693478
rect 45922 693437 45968 693449
rect 46080 693449 46086 694088
rect 46120 693449 46126 694088
rect 46238 693788 46244 694425
rect 46278 693788 46284 694425
rect 46396 694425 46442 694437
rect 46396 694398 46402 694425
rect 46436 694398 46442 694425
rect 46554 694425 46600 694437
rect 46378 694328 46388 694398
rect 46458 694328 46468 694398
rect 46396 694158 46402 694328
rect 46436 694158 46442 694328
rect 46378 694088 46388 694158
rect 46458 694088 46468 694158
rect 46218 693718 46228 693788
rect 46298 693718 46308 693788
rect 46238 693548 46244 693718
rect 46278 693548 46284 693718
rect 46218 693478 46228 693548
rect 46298 693478 46308 693548
rect 46080 693437 46126 693449
rect 46238 693449 46244 693478
rect 46278 693449 46284 693478
rect 46238 693437 46284 693449
rect 46396 693449 46402 694088
rect 46436 693449 46442 694088
rect 46554 693788 46560 694425
rect 46594 693788 46600 694425
rect 46712 694425 46758 694437
rect 46712 694398 46718 694425
rect 46752 694398 46758 694425
rect 46870 694425 46916 694437
rect 46688 694328 46698 694398
rect 46768 694328 46778 694398
rect 46712 694158 46718 694328
rect 46752 694158 46758 694328
rect 46688 694088 46698 694158
rect 46768 694088 46778 694158
rect 46538 693718 46548 693788
rect 46618 693718 46628 693788
rect 46554 693548 46560 693718
rect 46594 693548 46600 693718
rect 46538 693478 46548 693548
rect 46618 693478 46628 693548
rect 46396 693437 46442 693449
rect 46554 693449 46560 693478
rect 46594 693449 46600 693478
rect 46554 693437 46600 693449
rect 46712 693449 46718 694088
rect 46752 693449 46758 694088
rect 46870 693788 46876 694425
rect 46910 693788 46916 694425
rect 47028 694425 47074 694437
rect 47028 694398 47034 694425
rect 47068 694398 47074 694425
rect 47186 694425 47232 694437
rect 47008 694328 47018 694398
rect 47088 694328 47098 694398
rect 47028 694158 47034 694328
rect 47068 694158 47074 694328
rect 47008 694088 47018 694158
rect 47088 694088 47098 694158
rect 46848 693718 46858 693788
rect 46928 693718 46938 693788
rect 46870 693548 46876 693718
rect 46910 693548 46916 693718
rect 46848 693478 46858 693548
rect 46928 693478 46938 693548
rect 46712 693437 46758 693449
rect 46870 693449 46876 693478
rect 46910 693449 46916 693478
rect 46870 693437 46916 693449
rect 47028 693449 47034 694088
rect 47068 693449 47074 694088
rect 47186 693788 47192 694425
rect 47226 693788 47232 694425
rect 47344 694425 47390 694437
rect 47344 694398 47350 694425
rect 47384 694398 47390 694425
rect 47502 694425 47548 694437
rect 47328 694328 47338 694398
rect 47408 694328 47418 694398
rect 47344 694158 47350 694328
rect 47384 694158 47390 694328
rect 47328 694088 47338 694158
rect 47408 694088 47418 694158
rect 47168 693718 47178 693788
rect 47248 693718 47258 693788
rect 47186 693548 47192 693718
rect 47226 693548 47232 693718
rect 47168 693478 47178 693548
rect 47248 693478 47258 693548
rect 47028 693437 47074 693449
rect 47186 693449 47192 693478
rect 47226 693449 47232 693478
rect 47186 693437 47232 693449
rect 47344 693449 47350 694088
rect 47384 693449 47390 694088
rect 47502 693788 47508 694425
rect 47542 693788 47548 694425
rect 47660 694425 47706 694437
rect 47660 694398 47666 694425
rect 47700 694398 47706 694425
rect 47818 694425 47864 694437
rect 47638 694328 47648 694398
rect 47718 694328 47728 694398
rect 47660 694158 47666 694328
rect 47700 694158 47706 694328
rect 47638 694088 47648 694158
rect 47718 694088 47728 694158
rect 47478 693718 47488 693788
rect 47558 693718 47568 693788
rect 47502 693548 47508 693718
rect 47542 693548 47548 693718
rect 47478 693478 47488 693548
rect 47558 693478 47568 693548
rect 47344 693437 47390 693449
rect 47502 693449 47508 693478
rect 47542 693449 47548 693478
rect 47502 693437 47548 693449
rect 47660 693449 47666 694088
rect 47700 693449 47706 694088
rect 47818 693788 47824 694425
rect 47858 693788 47864 694425
rect 47976 694425 48022 694437
rect 47976 694398 47982 694425
rect 48016 694398 48022 694425
rect 48134 694425 48180 694437
rect 47958 694328 47968 694398
rect 48038 694328 48048 694398
rect 47976 694158 47982 694328
rect 48016 694158 48022 694328
rect 47958 694088 47968 694158
rect 48038 694088 48048 694158
rect 47798 693718 47808 693788
rect 47878 693718 47888 693788
rect 47818 693548 47824 693718
rect 47858 693548 47864 693718
rect 47798 693478 47808 693548
rect 47878 693478 47888 693548
rect 47660 693437 47706 693449
rect 47818 693449 47824 693478
rect 47858 693449 47864 693478
rect 47818 693437 47864 693449
rect 47976 693449 47982 694088
rect 48016 693449 48022 694088
rect 48134 693788 48140 694425
rect 48174 693788 48180 694425
rect 48292 694425 48338 694437
rect 48292 694398 48298 694425
rect 48332 694398 48338 694425
rect 48450 694425 48496 694437
rect 48268 694328 48278 694398
rect 48348 694328 48358 694398
rect 48292 694158 48298 694328
rect 48332 694158 48338 694328
rect 48268 694088 48278 694158
rect 48348 694088 48358 694158
rect 48118 693718 48128 693788
rect 48198 693718 48208 693788
rect 48134 693548 48140 693718
rect 48174 693548 48180 693718
rect 48118 693478 48128 693548
rect 48198 693478 48208 693548
rect 47976 693437 48022 693449
rect 48134 693449 48140 693478
rect 48174 693449 48180 693478
rect 48134 693437 48180 693449
rect 48292 693449 48298 694088
rect 48332 693449 48338 694088
rect 48450 693788 48456 694425
rect 48490 693788 48496 694425
rect 48608 694425 48654 694437
rect 48608 694398 48614 694425
rect 48648 694398 48654 694425
rect 48588 694328 48598 694398
rect 48668 694328 48678 694398
rect 48608 694158 48614 694328
rect 48648 694158 48654 694328
rect 48588 694088 48598 694158
rect 48668 694088 48678 694158
rect 48718 694098 48798 694478
rect 49568 694237 49589 695351
rect 49986 694237 50008 695351
rect 49568 694098 50008 694237
rect 48428 693718 48438 693788
rect 48508 693718 48518 693788
rect 48450 693556 48456 693718
rect 48428 693474 48456 693556
rect 48292 693437 48338 693449
rect 48450 693449 48456 693474
rect 48490 693556 48496 693718
rect 48490 693474 48520 693556
rect 48490 693449 48496 693474
rect 48450 693437 48496 693449
rect 48608 693449 48614 694088
rect 48648 693449 48654 694088
rect 48608 693437 48654 693449
rect 48718 693891 50008 694098
rect 48718 693808 49589 693891
rect 48718 693398 48798 693808
rect 42138 693390 48798 693398
rect 42138 693356 42356 693390
rect 42424 693356 42514 693390
rect 42582 693356 42672 693390
rect 42740 693356 42830 693390
rect 42898 693356 42988 693390
rect 43056 693356 43146 693390
rect 43214 693356 43304 693390
rect 43372 693378 43462 693390
rect 43372 693356 43408 693378
rect 43530 693356 43620 693390
rect 43688 693356 43778 693390
rect 43846 693356 43936 693390
rect 44004 693356 44094 693390
rect 44162 693356 44252 693390
rect 44320 693356 44410 693390
rect 44478 693356 44568 693390
rect 44636 693356 44726 693390
rect 44794 693356 44884 693390
rect 44952 693356 45042 693390
rect 45110 693356 45200 693390
rect 45268 693356 45358 693390
rect 45426 693356 45516 693390
rect 45584 693356 45674 693390
rect 45742 693356 45832 693390
rect 45900 693356 45990 693390
rect 46058 693356 46148 693390
rect 46216 693356 46306 693390
rect 46374 693356 46464 693390
rect 46532 693356 46622 693390
rect 46690 693356 46780 693390
rect 46848 693356 46938 693390
rect 47006 693356 47096 693390
rect 47164 693356 47254 693390
rect 47322 693356 47412 693390
rect 47480 693378 47570 693390
rect 47548 693356 47570 693378
rect 47638 693356 47728 693390
rect 47796 693356 47886 693390
rect 47954 693356 48044 693390
rect 48112 693356 48202 693390
rect 48270 693356 48360 693390
rect 48428 693356 48518 693390
rect 48586 693356 48798 693390
rect 42138 693348 43408 693356
rect 43368 693298 43408 693348
rect 43488 693348 47468 693356
rect 43488 693298 43528 693348
rect 47428 693298 47468 693348
rect 47548 693348 48798 693356
rect 47548 693298 47588 693348
rect 43368 693288 43528 693298
rect 44578 693294 46368 693298
rect 43831 693288 47111 693294
rect 47428 693288 47588 693298
rect 43831 693254 43843 693288
rect 47099 693254 47111 693288
rect 43831 693248 47111 693254
rect 44578 693238 46368 693248
rect 44578 692968 44798 693238
rect 45068 692968 45848 693238
rect 46118 692968 46368 693238
rect 44578 692950 46368 692968
rect 44578 692916 44594 692950
rect 46350 692916 46368 692950
rect 44578 692908 46368 692916
rect 40938 692758 41368 692777
rect 43648 692848 47298 692858
rect 43648 692814 43858 692848
rect 43926 692814 44016 692848
rect 44084 692814 44174 692848
rect 44242 692814 44332 692848
rect 44400 692814 44490 692848
rect 44558 692814 44648 692848
rect 44716 692814 44806 692848
rect 44874 692814 44964 692848
rect 45032 692814 45122 692848
rect 45190 692814 45280 692848
rect 45348 692814 45438 692848
rect 45506 692814 45596 692848
rect 45664 692814 45754 692848
rect 45822 692814 45912 692848
rect 45980 692814 46070 692848
rect 46138 692814 46228 692848
rect 46296 692814 46386 692848
rect 46454 692814 46544 692848
rect 46612 692814 46702 692848
rect 46770 692814 46860 692848
rect 46928 692814 47018 692848
rect 47086 692814 47298 692848
rect 43648 692808 47298 692814
rect 39566 692698 39770 692704
rect 39566 692598 39578 692698
rect 39758 692598 39770 692698
rect 39566 692592 39770 692598
rect 39986 692698 40190 692704
rect 39986 692598 39998 692698
rect 40178 692598 40190 692698
rect 39986 692592 40190 692598
rect 43648 692440 43728 692808
rect 43790 692755 43836 692767
rect 43648 692282 43730 692440
rect 43648 691728 43728 692282
rect 43790 692088 43796 692755
rect 43830 692088 43836 692755
rect 43948 692755 43994 692767
rect 43948 692728 43954 692755
rect 43988 692728 43994 692755
rect 44106 692755 44152 692767
rect 43928 692658 43938 692728
rect 44008 692658 44018 692728
rect 43948 692518 43954 692658
rect 43988 692518 43994 692658
rect 43928 692448 43938 692518
rect 44008 692448 44018 692518
rect 43768 692018 43778 692088
rect 43848 692018 43858 692088
rect 43790 691878 43796 692018
rect 43830 691878 43836 692018
rect 43768 691808 43778 691878
rect 43848 691808 43858 691878
rect 43790 691779 43796 691808
rect 43830 691779 43836 691808
rect 43790 691767 43836 691779
rect 43948 691779 43954 692448
rect 43988 691779 43994 692448
rect 44106 692088 44112 692755
rect 44146 692088 44152 692755
rect 44264 692755 44310 692767
rect 44264 692728 44270 692755
rect 44304 692728 44310 692755
rect 44422 692755 44468 692767
rect 44238 692658 44248 692728
rect 44318 692658 44328 692728
rect 44264 692518 44270 692658
rect 44304 692518 44310 692658
rect 44238 692448 44248 692518
rect 44318 692448 44328 692518
rect 44078 692018 44088 692088
rect 44158 692018 44168 692088
rect 44106 691878 44112 692018
rect 44146 691878 44152 692018
rect 44078 691808 44088 691878
rect 44158 691808 44168 691878
rect 43948 691767 43994 691779
rect 44106 691779 44112 691808
rect 44146 691779 44152 691808
rect 44106 691767 44152 691779
rect 44264 691779 44270 692448
rect 44304 691779 44310 692448
rect 44422 692088 44428 692755
rect 44462 692088 44468 692755
rect 44580 692755 44626 692767
rect 44580 692728 44586 692755
rect 44620 692728 44626 692755
rect 44738 692755 44784 692767
rect 44558 692658 44568 692728
rect 44638 692658 44648 692728
rect 44580 692518 44586 692658
rect 44620 692518 44626 692658
rect 44558 692448 44568 692518
rect 44638 692448 44648 692518
rect 44398 692018 44408 692088
rect 44478 692018 44488 692088
rect 44422 691878 44428 692018
rect 44462 691878 44468 692018
rect 44398 691808 44408 691878
rect 44478 691808 44488 691878
rect 44264 691767 44310 691779
rect 44422 691779 44428 691808
rect 44462 691779 44468 691808
rect 44422 691767 44468 691779
rect 44580 691779 44586 692448
rect 44620 691779 44626 692448
rect 44738 692088 44744 692755
rect 44778 692088 44784 692755
rect 44896 692755 44942 692767
rect 44896 692728 44902 692755
rect 44936 692728 44942 692755
rect 45054 692755 45100 692767
rect 44868 692658 44878 692728
rect 44948 692658 44958 692728
rect 44896 692518 44902 692658
rect 44936 692518 44942 692658
rect 44868 692448 44878 692518
rect 44948 692448 44958 692518
rect 44718 692018 44728 692088
rect 44798 692018 44808 692088
rect 44738 691878 44744 692018
rect 44778 691878 44784 692018
rect 44718 691808 44728 691878
rect 44798 691808 44808 691878
rect 44580 691767 44626 691779
rect 44738 691779 44744 691808
rect 44778 691779 44784 691808
rect 44738 691767 44784 691779
rect 44896 691779 44902 692448
rect 44936 691779 44942 692448
rect 45054 692088 45060 692755
rect 45094 692088 45100 692755
rect 45212 692755 45258 692767
rect 45212 692728 45218 692755
rect 45252 692728 45258 692755
rect 45370 692755 45416 692767
rect 45188 692658 45198 692728
rect 45268 692658 45278 692728
rect 45212 692518 45218 692658
rect 45252 692518 45258 692658
rect 45188 692448 45198 692518
rect 45268 692448 45278 692518
rect 45028 692018 45038 692088
rect 45108 692018 45118 692088
rect 45054 691878 45060 692018
rect 45094 691878 45100 692018
rect 45028 691808 45038 691878
rect 45108 691808 45118 691878
rect 44896 691767 44942 691779
rect 45054 691779 45060 691808
rect 45094 691779 45100 691808
rect 45054 691767 45100 691779
rect 45212 691779 45218 692448
rect 45252 691779 45258 692448
rect 45370 692088 45376 692755
rect 45410 692088 45416 692755
rect 45528 692755 45574 692767
rect 45528 692728 45534 692755
rect 45568 692728 45574 692755
rect 45686 692755 45732 692767
rect 45508 692658 45518 692728
rect 45588 692658 45598 692728
rect 45528 692518 45534 692658
rect 45568 692518 45574 692658
rect 45508 692448 45518 692518
rect 45588 692448 45598 692518
rect 45348 692018 45358 692088
rect 45428 692018 45438 692088
rect 45370 691878 45376 692018
rect 45410 691878 45416 692018
rect 45348 691808 45358 691878
rect 45428 691808 45438 691878
rect 45212 691767 45258 691779
rect 45370 691779 45376 691808
rect 45410 691779 45416 691808
rect 45370 691767 45416 691779
rect 45528 691779 45534 692448
rect 45568 691779 45574 692448
rect 45686 692088 45692 692755
rect 45726 692088 45732 692755
rect 45844 692755 45890 692767
rect 45844 692728 45850 692755
rect 45884 692728 45890 692755
rect 46002 692755 46048 692767
rect 45818 692658 45828 692728
rect 45898 692658 45908 692728
rect 45844 692518 45850 692658
rect 45884 692518 45890 692658
rect 45818 692448 45828 692518
rect 45898 692448 45908 692518
rect 45658 692018 45668 692088
rect 45738 692018 45748 692088
rect 45686 691878 45692 692018
rect 45726 691878 45732 692018
rect 45658 691808 45668 691878
rect 45738 691808 45748 691878
rect 45528 691767 45574 691779
rect 45686 691779 45692 691808
rect 45726 691779 45732 691808
rect 45686 691767 45732 691779
rect 45844 691779 45850 692448
rect 45884 691779 45890 692448
rect 46002 692088 46008 692755
rect 46042 692088 46048 692755
rect 46160 692755 46206 692767
rect 46160 692728 46166 692755
rect 46200 692728 46206 692755
rect 46318 692755 46364 692767
rect 46138 692658 46148 692728
rect 46218 692658 46228 692728
rect 46160 692518 46166 692658
rect 46200 692518 46206 692658
rect 46138 692448 46148 692518
rect 46218 692448 46228 692518
rect 45978 692018 45988 692088
rect 46058 692018 46068 692088
rect 46002 691878 46008 692018
rect 46042 691878 46048 692018
rect 45978 691808 45988 691878
rect 46058 691808 46068 691878
rect 45844 691767 45890 691779
rect 46002 691779 46008 691808
rect 46042 691779 46048 691808
rect 46002 691767 46048 691779
rect 46160 691779 46166 692448
rect 46200 691779 46206 692448
rect 46318 692088 46324 692755
rect 46358 692088 46364 692755
rect 46476 692755 46522 692767
rect 46476 692728 46482 692755
rect 46516 692728 46522 692755
rect 46634 692755 46680 692767
rect 46458 692658 46468 692728
rect 46538 692658 46548 692728
rect 46476 692518 46482 692658
rect 46516 692518 46522 692658
rect 46458 692448 46468 692518
rect 46538 692448 46548 692518
rect 46298 692018 46308 692088
rect 46378 692018 46388 692088
rect 46318 691878 46324 692018
rect 46358 691878 46364 692018
rect 46298 691808 46308 691878
rect 46378 691808 46388 691878
rect 46160 691767 46206 691779
rect 46318 691779 46324 691808
rect 46358 691779 46364 691808
rect 46318 691767 46364 691779
rect 46476 691779 46482 692448
rect 46516 691779 46522 692448
rect 46634 692088 46640 692755
rect 46674 692088 46680 692755
rect 46792 692755 46838 692767
rect 46792 692728 46798 692755
rect 46832 692728 46838 692755
rect 46950 692755 46996 692767
rect 46768 692658 46778 692728
rect 46848 692658 46858 692728
rect 46792 692518 46798 692658
rect 46832 692518 46838 692658
rect 46768 692448 46778 692518
rect 46848 692448 46858 692518
rect 46608 692018 46618 692088
rect 46688 692018 46698 692088
rect 46634 691878 46640 692018
rect 46674 691878 46680 692018
rect 46608 691808 46618 691878
rect 46688 691808 46698 691878
rect 46476 691767 46522 691779
rect 46634 691779 46640 691808
rect 46674 691779 46680 691808
rect 46634 691767 46680 691779
rect 46792 691779 46798 692448
rect 46832 691779 46838 692448
rect 46950 692088 46956 692755
rect 46990 692088 46996 692755
rect 47108 692755 47154 692767
rect 47108 692728 47114 692755
rect 47148 692728 47154 692755
rect 47088 692658 47098 692728
rect 47168 692658 47178 692728
rect 47108 692518 47114 692658
rect 47148 692518 47154 692658
rect 47088 692448 47098 692518
rect 47168 692448 47178 692518
rect 46928 692018 46938 692088
rect 47008 692018 47018 692088
rect 46950 691878 46956 692018
rect 46990 691878 46996 692018
rect 46928 691808 46938 691878
rect 47008 691808 47018 691878
rect 46792 691767 46838 691779
rect 46950 691779 46956 691808
rect 46990 691779 46996 691808
rect 46950 691767 46996 691779
rect 47108 691779 47114 692448
rect 47148 691779 47154 692448
rect 47108 691767 47154 691779
rect 47218 691728 47298 692808
rect 49568 692777 49589 693808
rect 49986 692777 50008 693891
rect 49568 692758 50008 692777
rect 51998 695351 52438 695368
rect 51998 694237 52020 695351
rect 52417 694237 52438 695351
rect 51998 694178 52438 694237
rect 51998 694158 53328 694178
rect 51998 694088 53128 694158
rect 53198 694088 53328 694158
rect 51998 694048 53328 694088
rect 51998 693978 53238 694048
rect 53308 693978 53328 694048
rect 51998 693958 53328 693978
rect 51998 693891 52438 693958
rect 51998 692777 52020 693891
rect 52417 692777 52438 693891
rect 51998 692758 52438 692777
rect 50816 692698 51020 692704
rect 50816 692598 50828 692698
rect 51008 692598 51020 692698
rect 50816 692592 51020 692598
rect 51236 692698 51440 692704
rect 51236 692598 51248 692698
rect 51428 692598 51440 692698
rect 51236 692592 51440 692598
rect 43648 691720 47298 691728
rect 43648 691686 43858 691720
rect 43926 691686 44016 691720
rect 44084 691686 44174 691720
rect 44242 691686 44332 691720
rect 44400 691686 44490 691720
rect 44558 691686 44648 691720
rect 44716 691686 44806 691720
rect 44874 691686 44964 691720
rect 45032 691686 45122 691720
rect 45190 691686 45280 691720
rect 45348 691686 45438 691720
rect 45506 691686 45596 691720
rect 45664 691686 45754 691720
rect 45822 691686 45912 691720
rect 45980 691686 46070 691720
rect 46138 691686 46228 691720
rect 46296 691686 46386 691720
rect 46454 691686 46544 691720
rect 46612 691686 46702 691720
rect 46770 691686 46860 691720
rect 46928 691686 47018 691720
rect 47086 691686 47298 691720
rect 43648 691678 47298 691686
rect 43838 691318 44108 691678
rect 44578 691624 44588 691628
rect 44436 691618 44588 691624
rect 44848 691624 44858 691628
rect 44848 691618 45030 691624
rect 44436 691378 44448 691618
rect 45018 691378 45030 691618
rect 44436 691372 44588 691378
rect 44578 691368 44588 691372
rect 44848 691372 45030 691378
rect 44848 691368 44858 691372
rect 45338 691318 45608 691678
rect 46078 691624 46088 691628
rect 45906 691618 46088 691624
rect 46348 691624 46358 691628
rect 46348 691618 46500 691624
rect 45906 691378 45918 691618
rect 46488 691378 46500 691618
rect 45906 691372 46088 691378
rect 46078 691368 46088 691372
rect 46348 691372 46500 691378
rect 46348 691368 46358 691372
rect 46838 691318 47108 691678
rect 43838 691308 47108 691318
rect 43838 691274 43858 691308
rect 43926 691274 44016 691308
rect 44084 691274 44174 691308
rect 44242 691274 44332 691308
rect 44400 691274 44490 691308
rect 44558 691274 44648 691308
rect 44716 691274 44806 691308
rect 44874 691274 44964 691308
rect 45032 691274 45122 691308
rect 45190 691274 45280 691308
rect 45348 691274 45438 691308
rect 45506 691274 45596 691308
rect 45664 691274 45754 691308
rect 45822 691274 45912 691308
rect 45980 691274 46070 691308
rect 46138 691274 46228 691308
rect 46296 691274 46386 691308
rect 46454 691274 46544 691308
rect 46612 691274 46702 691308
rect 46770 691274 46860 691308
rect 46928 691274 47018 691308
rect 47086 691274 47108 691308
rect 43838 691268 47108 691274
rect 43790 691215 43836 691227
rect 43790 690548 43796 691215
rect 43830 690548 43836 691215
rect 43948 691215 43994 691227
rect 43948 691178 43954 691215
rect 43988 691178 43994 691215
rect 44098 691215 44158 691268
rect 43928 691108 43938 691178
rect 44008 691108 44018 691178
rect 43948 690968 43954 691108
rect 43988 690968 43994 691108
rect 43928 690898 43938 690968
rect 44008 690898 44018 690968
rect 43768 690478 43778 690548
rect 43848 690478 43858 690548
rect 43790 690338 43796 690478
rect 43830 690338 43836 690478
rect 43768 690268 43778 690338
rect 43848 690268 43858 690338
rect 43790 690239 43796 690268
rect 43830 690239 43836 690268
rect 43790 690227 43836 690239
rect 43948 690239 43954 690898
rect 43988 690239 43994 690898
rect 44098 690548 44112 691215
rect 44146 690548 44158 691215
rect 44264 691215 44310 691227
rect 44264 691178 44270 691215
rect 44304 691178 44310 691215
rect 44418 691215 44478 691268
rect 44238 691108 44248 691178
rect 44318 691108 44328 691178
rect 44264 690968 44270 691108
rect 44304 690968 44310 691108
rect 44238 690898 44248 690968
rect 44318 690898 44328 690968
rect 44088 690478 44098 690548
rect 44168 690478 44178 690548
rect 44098 690338 44112 690478
rect 44146 690338 44158 690478
rect 44088 690268 44098 690338
rect 44168 690268 44178 690338
rect 43948 690227 43994 690239
rect 44098 690239 44112 690268
rect 44146 690239 44158 690268
rect 44098 690188 44158 690239
rect 44264 690239 44270 690898
rect 44304 690239 44310 690898
rect 44418 690548 44428 691215
rect 44462 690548 44478 691215
rect 44580 691215 44626 691227
rect 44580 691178 44586 691215
rect 44620 691178 44626 691215
rect 44738 691215 44784 691227
rect 44558 691108 44568 691178
rect 44638 691108 44648 691178
rect 44580 690968 44586 691108
rect 44620 690968 44626 691108
rect 44558 690898 44568 690968
rect 44638 690898 44648 690968
rect 44398 690478 44408 690548
rect 44478 690478 44488 690548
rect 44418 690338 44428 690478
rect 44462 690338 44478 690478
rect 44398 690268 44408 690338
rect 44478 690268 44488 690338
rect 44264 690227 44310 690239
rect 44418 690239 44428 690268
rect 44462 690239 44478 690268
rect 44418 690188 44478 690239
rect 44580 690239 44586 690898
rect 44620 690239 44626 690898
rect 44738 690548 44744 691215
rect 44778 690548 44784 691215
rect 44896 691215 44942 691227
rect 44896 691178 44902 691215
rect 44936 691178 44942 691215
rect 45054 691215 45100 691227
rect 44878 691108 44888 691178
rect 44958 691108 44968 691178
rect 44896 690968 44902 691108
rect 44936 690968 44942 691108
rect 44878 690898 44888 690968
rect 44958 690898 44968 690968
rect 44718 690478 44728 690548
rect 44798 690478 44808 690548
rect 44738 690338 44744 690478
rect 44778 690338 44784 690478
rect 44718 690268 44728 690338
rect 44798 690268 44808 690338
rect 44580 690227 44626 690239
rect 44738 690239 44744 690268
rect 44778 690239 44784 690268
rect 44738 690227 44784 690239
rect 44896 690239 44902 690898
rect 44936 690239 44942 690898
rect 45054 690548 45060 691215
rect 45094 690548 45100 691215
rect 45212 691215 45258 691227
rect 45212 691178 45218 691215
rect 45252 691178 45258 691215
rect 45370 691215 45416 691227
rect 45188 691108 45198 691178
rect 45268 691108 45278 691178
rect 45212 690968 45218 691108
rect 45252 690968 45258 691108
rect 45188 690898 45198 690968
rect 45268 690898 45278 690968
rect 45028 690478 45038 690548
rect 45108 690478 45118 690548
rect 45054 690338 45060 690478
rect 45094 690338 45100 690478
rect 45028 690268 45038 690338
rect 45108 690268 45118 690338
rect 44896 690227 44942 690239
rect 45054 690239 45060 690268
rect 45094 690239 45100 690268
rect 45054 690227 45100 690239
rect 45212 690239 45218 690898
rect 45252 690239 45258 690898
rect 45370 690548 45376 691215
rect 45410 690548 45416 691215
rect 45528 691215 45574 691227
rect 45528 691178 45534 691215
rect 45568 691178 45574 691215
rect 45686 691215 45732 691227
rect 45508 691108 45518 691178
rect 45588 691108 45598 691178
rect 45528 690968 45534 691108
rect 45568 690968 45574 691108
rect 45508 690898 45518 690968
rect 45588 690898 45598 690968
rect 45348 690478 45358 690548
rect 45428 690478 45438 690548
rect 45370 690338 45376 690478
rect 45410 690338 45416 690478
rect 45348 690268 45358 690338
rect 45428 690268 45438 690338
rect 45212 690227 45258 690239
rect 45370 690239 45376 690268
rect 45410 690239 45416 690268
rect 45370 690227 45416 690239
rect 45528 690239 45534 690898
rect 45568 690239 45574 690898
rect 45686 690548 45692 691215
rect 45726 690548 45732 691215
rect 45844 691215 45890 691227
rect 45844 691178 45850 691215
rect 45884 691178 45890 691215
rect 46002 691215 46048 691227
rect 45818 691108 45828 691178
rect 45898 691108 45908 691178
rect 45844 690968 45850 691108
rect 45884 690968 45890 691108
rect 45818 690898 45828 690968
rect 45898 690898 45908 690968
rect 45668 690478 45678 690548
rect 45748 690478 45758 690548
rect 45686 690338 45692 690478
rect 45726 690338 45732 690478
rect 45668 690268 45678 690338
rect 45748 690268 45758 690338
rect 45528 690227 45574 690239
rect 45686 690239 45692 690268
rect 45726 690239 45732 690268
rect 45686 690227 45732 690239
rect 45844 690239 45850 690898
rect 45884 690239 45890 690898
rect 46002 690548 46008 691215
rect 46042 690548 46048 691215
rect 46160 691215 46206 691227
rect 46160 691178 46166 691215
rect 46200 691178 46206 691215
rect 46308 691215 46368 691268
rect 46138 691108 46148 691178
rect 46218 691108 46228 691178
rect 46160 690968 46166 691108
rect 46200 690968 46206 691108
rect 46138 690898 46148 690968
rect 46218 690898 46228 690968
rect 45978 690478 45988 690548
rect 46058 690478 46068 690548
rect 46002 690338 46008 690478
rect 46042 690338 46048 690478
rect 45978 690268 45988 690338
rect 46058 690268 46068 690338
rect 45844 690227 45890 690239
rect 46002 690239 46008 690268
rect 46042 690239 46048 690268
rect 46002 690227 46048 690239
rect 46160 690239 46166 690898
rect 46200 690239 46206 690898
rect 46308 690548 46324 691215
rect 46358 690548 46368 691215
rect 46476 691215 46522 691227
rect 46476 691178 46482 691215
rect 46516 691178 46522 691215
rect 46628 691215 46688 691268
rect 46458 691108 46468 691178
rect 46538 691108 46548 691178
rect 46476 690968 46482 691108
rect 46516 690968 46522 691108
rect 46458 690898 46468 690968
rect 46538 690898 46548 690968
rect 46298 690478 46308 690548
rect 46378 690478 46388 690548
rect 46308 690338 46324 690478
rect 46358 690338 46368 690478
rect 46298 690268 46308 690338
rect 46378 690268 46388 690338
rect 46160 690227 46206 690239
rect 46308 690239 46324 690268
rect 46358 690239 46368 690268
rect 46308 690188 46368 690239
rect 46476 690239 46482 690898
rect 46516 690239 46522 690898
rect 46628 690548 46640 691215
rect 46674 690548 46688 691215
rect 46792 691215 46838 691227
rect 46792 691178 46798 691215
rect 46832 691178 46838 691215
rect 46950 691215 46996 691227
rect 46768 691108 46778 691178
rect 46848 691108 46858 691178
rect 46792 690968 46798 691108
rect 46832 690968 46838 691108
rect 46768 690898 46778 690968
rect 46848 690898 46858 690968
rect 46608 690478 46618 690548
rect 46688 690478 46698 690548
rect 46628 690338 46640 690478
rect 46674 690338 46688 690478
rect 46608 690268 46618 690338
rect 46688 690268 46698 690338
rect 46476 690227 46522 690239
rect 46628 690239 46640 690268
rect 46674 690239 46688 690268
rect 46628 690188 46688 690239
rect 46792 690239 46798 690898
rect 46832 690239 46838 690898
rect 46950 690548 46956 691215
rect 46990 690548 46996 691215
rect 47108 691215 47154 691227
rect 47108 691178 47114 691215
rect 47148 691178 47154 691215
rect 47088 691108 47098 691178
rect 47168 691108 47178 691178
rect 47108 690968 47114 691108
rect 47148 690968 47154 691108
rect 47088 690898 47098 690968
rect 47168 690898 47178 690968
rect 46928 690478 46938 690548
rect 47008 690478 47018 690548
rect 46950 690338 46956 690478
rect 46990 690338 46996 690478
rect 46928 690268 46938 690338
rect 47008 690268 47018 690338
rect 46792 690227 46838 690239
rect 46950 690239 46956 690268
rect 46990 690239 46996 690268
rect 46950 690227 46996 690239
rect 47108 690239 47114 690898
rect 47148 690239 47154 690898
rect 47108 690227 47154 690239
rect 43838 690180 47108 690188
rect 43838 690146 43858 690180
rect 43926 690146 44016 690180
rect 44084 690146 44174 690180
rect 44242 690146 44332 690180
rect 44400 690146 44490 690180
rect 44558 690146 44648 690180
rect 44716 690146 44806 690180
rect 44874 690146 44964 690180
rect 45032 690146 45122 690180
rect 45190 690146 45280 690180
rect 45348 690146 45438 690180
rect 45506 690146 45596 690180
rect 45664 690146 45754 690180
rect 45822 690146 45912 690180
rect 45980 690146 46070 690180
rect 46138 690146 46228 690180
rect 46296 690146 46386 690180
rect 46454 690146 46544 690180
rect 46612 690146 46702 690180
rect 46770 690146 46860 690180
rect 46928 690146 47018 690180
rect 47086 690146 47108 690180
rect 43838 690138 47108 690146
rect 45140 689833 45814 689839
rect 45140 689799 45152 689833
rect 45802 689799 45814 689833
rect 45140 689793 45814 689799
rect 44698 689731 46258 689738
rect 44698 689697 44969 689731
rect 45037 689697 45127 689731
rect 45195 689697 45285 689731
rect 45353 689697 45443 689731
rect 45511 689697 45601 689731
rect 45669 689697 45759 689731
rect 45827 689697 45917 689731
rect 45985 689697 46258 689731
rect 44698 689688 46258 689697
rect 44698 688628 44778 689688
rect 44901 689647 44947 689659
rect 44901 689058 44907 689647
rect 44941 689058 44947 689647
rect 45059 689647 45105 689659
rect 45059 689618 45065 689647
rect 45099 689618 45105 689647
rect 45217 689647 45263 689659
rect 45038 689548 45048 689618
rect 45118 689548 45128 689618
rect 45059 689328 45065 689548
rect 45099 689328 45105 689548
rect 45038 689258 45048 689328
rect 45118 689258 45128 689328
rect 44878 688988 44888 689058
rect 44958 688988 44968 689058
rect 44901 688768 44907 688988
rect 44941 688768 44947 688988
rect 44878 688698 44888 688768
rect 44958 688698 44968 688768
rect 44901 688671 44907 688698
rect 44941 688671 44947 688698
rect 44901 688659 44947 688671
rect 45059 688671 45065 689258
rect 45099 688671 45105 689258
rect 45217 689058 45223 689647
rect 45257 689058 45263 689647
rect 45375 689647 45421 689659
rect 45375 689618 45381 689647
rect 45415 689618 45421 689647
rect 45533 689647 45579 689659
rect 45358 689548 45368 689618
rect 45438 689548 45448 689618
rect 45375 689328 45381 689548
rect 45415 689328 45421 689548
rect 45358 689258 45368 689328
rect 45438 689258 45448 689328
rect 45198 688988 45208 689058
rect 45278 688988 45288 689058
rect 45217 688768 45223 688988
rect 45257 688768 45263 688988
rect 45198 688698 45208 688768
rect 45278 688698 45288 688768
rect 45059 688659 45105 688671
rect 45217 688671 45223 688698
rect 45257 688671 45263 688698
rect 45217 688659 45263 688671
rect 45375 688671 45381 689258
rect 45415 688671 45421 689258
rect 45533 689058 45539 689647
rect 45573 689058 45579 689647
rect 45691 689647 45737 689659
rect 45691 689618 45697 689647
rect 45731 689618 45737 689647
rect 45849 689647 45895 689659
rect 45668 689548 45678 689618
rect 45748 689548 45758 689618
rect 45691 689328 45697 689548
rect 45731 689328 45737 689548
rect 45668 689258 45678 689328
rect 45748 689258 45758 689328
rect 45518 688988 45528 689058
rect 45598 688988 45608 689058
rect 45533 688768 45539 688988
rect 45573 688768 45579 688988
rect 45518 688698 45528 688768
rect 45598 688698 45608 688768
rect 45375 688659 45421 688671
rect 45533 688671 45539 688698
rect 45573 688671 45579 688698
rect 45533 688659 45579 688671
rect 45691 688671 45697 689258
rect 45731 688671 45737 689258
rect 45849 689058 45855 689647
rect 45889 689058 45895 689647
rect 46007 689647 46053 689659
rect 46007 689618 46013 689647
rect 46047 689618 46053 689647
rect 45988 689548 45998 689618
rect 46068 689548 46078 689618
rect 46007 689328 46013 689548
rect 46047 689328 46053 689548
rect 45988 689258 45998 689328
rect 46068 689258 46078 689328
rect 46178 689280 46258 689688
rect 47940 689280 48120 689400
rect 45828 688988 45838 689058
rect 45908 688988 45918 689058
rect 45849 688768 45855 688988
rect 45889 688768 45895 688988
rect 45828 688698 45838 688768
rect 45908 688698 45918 688768
rect 45691 688659 45737 688671
rect 45849 688671 45855 688698
rect 45889 688671 45895 688698
rect 45849 688659 45895 688671
rect 46007 688671 46013 689258
rect 46047 688671 46053 689258
rect 46007 688659 46053 688671
rect 46178 689220 48120 689280
rect 46178 689100 47960 689220
rect 48100 689100 48120 689220
rect 46178 689040 48120 689100
rect 46178 688628 46258 689040
rect 47940 688900 48120 689040
rect 44698 688621 46258 688628
rect 44698 688587 44969 688621
rect 45037 688587 45127 688621
rect 45195 688587 45285 688621
rect 45353 688587 45443 688621
rect 45511 688587 45601 688621
rect 45669 688587 45759 688621
rect 45827 688587 45917 688621
rect 45985 688587 46258 688621
rect 44698 688578 46258 688587
rect 45338 688525 45348 688528
rect 45140 688519 45348 688525
rect 45608 688525 45618 688528
rect 45608 688519 45814 688525
rect 45140 688485 45152 688519
rect 45802 688485 45814 688519
rect 45140 688479 45348 688485
rect 45338 688319 45348 688479
rect 45140 688313 45348 688319
rect 45608 688479 45814 688485
rect 45608 688319 45618 688479
rect 45608 688313 45814 688319
rect 45140 688279 45152 688313
rect 45802 688279 45814 688313
rect 45140 688273 45348 688279
rect 45338 688268 45348 688273
rect 45608 688273 45814 688279
rect 45608 688268 45618 688273
rect 44698 688211 46258 688218
rect 44698 688177 44969 688211
rect 45037 688177 45127 688211
rect 45195 688177 45285 688211
rect 45353 688177 45443 688211
rect 45511 688177 45601 688211
rect 45669 688177 45759 688211
rect 45827 688177 45917 688211
rect 45985 688177 46258 688211
rect 44698 688168 46258 688177
rect 44698 687920 44778 688168
rect 44901 688127 44947 688139
rect 43320 687720 44780 687920
rect 43320 687560 43340 687720
rect 43460 687560 44780 687720
rect 43320 687520 44780 687560
rect 44901 687538 44907 688127
rect 44941 687538 44947 688127
rect 45059 688127 45105 688139
rect 45059 688098 45065 688127
rect 45099 688098 45105 688127
rect 45217 688127 45263 688139
rect 45038 688028 45048 688098
rect 45118 688028 45128 688098
rect 45059 687808 45065 688028
rect 45099 687808 45105 688028
rect 45038 687738 45048 687808
rect 45118 687738 45128 687808
rect 44698 687108 44778 687520
rect 44878 687468 44888 687538
rect 44958 687468 44968 687538
rect 44901 687248 44907 687468
rect 44941 687248 44947 687468
rect 44878 687178 44888 687248
rect 44958 687178 44968 687248
rect 44901 687151 44907 687178
rect 44941 687151 44947 687178
rect 44901 687139 44947 687151
rect 45059 687151 45065 687738
rect 45099 687151 45105 687738
rect 45217 687538 45223 688127
rect 45257 687538 45263 688127
rect 45375 688127 45421 688139
rect 45375 688098 45381 688127
rect 45415 688098 45421 688127
rect 45533 688127 45579 688139
rect 45358 688028 45368 688098
rect 45438 688028 45448 688098
rect 45375 687808 45381 688028
rect 45415 687808 45421 688028
rect 45358 687738 45368 687808
rect 45438 687738 45448 687808
rect 45198 687468 45208 687538
rect 45278 687468 45288 687538
rect 45217 687248 45223 687468
rect 45257 687248 45263 687468
rect 45198 687178 45208 687248
rect 45278 687178 45288 687248
rect 45059 687139 45105 687151
rect 45217 687151 45223 687178
rect 45257 687151 45263 687178
rect 45217 687139 45263 687151
rect 45375 687151 45381 687738
rect 45415 687151 45421 687738
rect 45533 687538 45539 688127
rect 45573 687538 45579 688127
rect 45691 688127 45737 688139
rect 45691 688098 45697 688127
rect 45731 688098 45737 688127
rect 45849 688127 45895 688139
rect 45668 688028 45678 688098
rect 45748 688028 45758 688098
rect 45691 687808 45697 688028
rect 45731 687808 45737 688028
rect 45668 687738 45678 687808
rect 45748 687738 45758 687808
rect 45518 687468 45528 687538
rect 45598 687468 45608 687538
rect 45533 687248 45539 687468
rect 45573 687248 45579 687468
rect 45518 687178 45528 687248
rect 45598 687178 45608 687248
rect 45375 687139 45421 687151
rect 45533 687151 45539 687178
rect 45573 687151 45579 687178
rect 45533 687139 45579 687151
rect 45691 687151 45697 687738
rect 45731 687151 45737 687738
rect 45849 687538 45855 688127
rect 45889 687538 45895 688127
rect 46007 688127 46053 688139
rect 46007 688098 46013 688127
rect 46047 688098 46053 688127
rect 45988 688028 45998 688098
rect 46068 688028 46078 688098
rect 46007 687808 46013 688028
rect 46047 687808 46053 688028
rect 45988 687738 45998 687808
rect 46068 687738 46078 687808
rect 45828 687468 45838 687538
rect 45908 687468 45918 687538
rect 45849 687248 45855 687468
rect 45889 687248 45895 687468
rect 45828 687178 45838 687248
rect 45908 687178 45918 687248
rect 45691 687139 45737 687151
rect 45849 687151 45855 687178
rect 45889 687151 45895 687178
rect 45849 687139 45895 687151
rect 46007 687151 46013 687738
rect 46047 687151 46053 687738
rect 46007 687139 46053 687151
rect 46178 687108 46258 688168
rect 44698 687101 46258 687108
rect 44698 687067 44969 687101
rect 45037 687067 45127 687101
rect 45195 687067 45285 687101
rect 45353 687067 45443 687101
rect 45511 687067 45601 687101
rect 45669 687067 45759 687101
rect 45827 687067 45917 687101
rect 45985 687067 46258 687101
rect 44698 687058 46258 687067
rect 45338 687005 45348 687008
rect 45140 686999 45348 687005
rect 45608 687005 45618 687008
rect 45608 686999 45814 687005
rect 45140 686965 45152 686999
rect 45802 686965 45814 686999
rect 45140 686959 45348 686965
rect 45338 686798 45348 686959
rect 44639 686792 45348 686798
rect 45608 686959 45814 686965
rect 45608 686798 45618 686959
rect 45608 686792 46307 686798
rect 44639 686758 44651 686792
rect 46295 686758 46307 686792
rect 44639 686752 45348 686758
rect 45338 686748 45348 686752
rect 45608 686752 46307 686758
rect 45608 686748 45618 686752
rect 43098 686698 43108 686728
rect 43088 686648 43108 686698
rect 43098 686618 43108 686648
rect 43218 686698 43228 686728
rect 43348 686698 43358 686728
rect 43218 686648 43358 686698
rect 43218 686618 43228 686648
rect 43348 686618 43358 686648
rect 43468 686698 43478 686728
rect 47498 686698 47508 686728
rect 43468 686690 47508 686698
rect 43468 686656 43970 686690
rect 44138 686656 44228 686690
rect 44396 686656 44486 686690
rect 44654 686656 44744 686690
rect 44912 686656 45002 686690
rect 45170 686656 45260 686690
rect 45428 686656 45518 686690
rect 45686 686656 45776 686690
rect 45944 686656 46034 686690
rect 46202 686656 46292 686690
rect 46460 686656 46550 686690
rect 46718 686656 46808 686690
rect 46976 686656 47508 686690
rect 43468 686648 47508 686656
rect 43468 686618 43478 686648
rect 47498 686618 47508 686648
rect 47618 686698 47628 686728
rect 47748 686698 47758 686728
rect 47618 686648 47758 686698
rect 47618 686618 47628 686648
rect 47748 686618 47758 686648
rect 47868 686698 47878 686728
rect 47868 686648 47888 686698
rect 47868 686618 47878 686648
rect 43902 686606 43948 686618
rect 43902 686578 43908 686606
rect 43942 686578 43948 686606
rect 44160 686606 44206 686618
rect 43878 686508 43888 686578
rect 43958 686508 43968 686578
rect 43902 686398 43908 686508
rect 43942 686398 43948 686508
rect 43878 686328 43888 686398
rect 43958 686328 43968 686398
rect 43902 685630 43908 686328
rect 43942 685630 43948 686328
rect 44160 685908 44166 686606
rect 44200 685908 44206 686606
rect 44418 686606 44464 686618
rect 44418 686578 44424 686606
rect 44458 686578 44464 686606
rect 44676 686606 44722 686618
rect 44398 686508 44408 686578
rect 44478 686508 44488 686578
rect 44418 686398 44424 686508
rect 44458 686398 44464 686508
rect 44398 686328 44408 686398
rect 44478 686328 44488 686398
rect 44138 685838 44148 685908
rect 44218 685838 44228 685908
rect 44160 685728 44166 685838
rect 44200 685728 44206 685838
rect 44138 685658 44148 685728
rect 44218 685658 44228 685728
rect 43902 685618 43948 685630
rect 44160 685630 44166 685658
rect 44200 685630 44206 685658
rect 44160 685618 44206 685630
rect 44418 685630 44424 686328
rect 44458 685630 44464 686328
rect 44676 685908 44682 686606
rect 44716 685908 44722 686606
rect 44934 686606 44980 686618
rect 44934 686578 44940 686606
rect 44974 686578 44980 686606
rect 45192 686606 45238 686618
rect 44918 686508 44928 686578
rect 44998 686508 45008 686578
rect 44934 686398 44940 686508
rect 44974 686398 44980 686508
rect 44918 686328 44928 686398
rect 44998 686328 45008 686398
rect 44658 685838 44668 685908
rect 44738 685838 44748 685908
rect 44676 685728 44682 685838
rect 44716 685728 44722 685838
rect 44658 685658 44668 685728
rect 44738 685658 44748 685728
rect 44418 685618 44464 685630
rect 44676 685630 44682 685658
rect 44716 685630 44722 685658
rect 44676 685618 44722 685630
rect 44934 685630 44940 686328
rect 44974 685630 44980 686328
rect 45192 685908 45198 686606
rect 45232 685908 45238 686606
rect 45450 686606 45496 686618
rect 45450 686578 45456 686606
rect 45490 686578 45496 686606
rect 45708 686606 45754 686618
rect 45428 686508 45438 686578
rect 45508 686508 45518 686578
rect 45450 686398 45456 686508
rect 45490 686398 45496 686508
rect 45428 686328 45438 686398
rect 45508 686328 45518 686398
rect 45168 685838 45178 685908
rect 45248 685838 45258 685908
rect 45192 685728 45198 685838
rect 45232 685728 45238 685838
rect 45168 685658 45178 685728
rect 45248 685658 45258 685728
rect 44934 685618 44980 685630
rect 45192 685630 45198 685658
rect 45232 685630 45238 685658
rect 45192 685618 45238 685630
rect 45450 685630 45456 686328
rect 45490 685630 45496 686328
rect 45708 685908 45714 686606
rect 45748 685908 45754 686606
rect 45966 686606 46012 686618
rect 45966 686578 45972 686606
rect 46006 686578 46012 686606
rect 46224 686606 46270 686618
rect 45948 686508 45958 686578
rect 46028 686508 46038 686578
rect 45966 686398 45972 686508
rect 46006 686398 46012 686508
rect 45948 686328 45958 686398
rect 46028 686328 46038 686398
rect 45688 685838 45698 685908
rect 45768 685838 45778 685908
rect 45708 685728 45714 685838
rect 45748 685728 45754 685838
rect 45688 685658 45698 685728
rect 45768 685658 45778 685728
rect 45450 685618 45496 685630
rect 45708 685630 45714 685658
rect 45748 685630 45754 685658
rect 45708 685618 45754 685630
rect 45966 685630 45972 686328
rect 46006 685630 46012 686328
rect 46224 685908 46230 686606
rect 46264 685908 46270 686606
rect 46482 686606 46528 686618
rect 46482 686578 46488 686606
rect 46522 686578 46528 686606
rect 46740 686606 46786 686618
rect 46458 686508 46468 686578
rect 46538 686508 46548 686578
rect 46482 686398 46488 686508
rect 46522 686398 46528 686508
rect 46458 686328 46468 686398
rect 46538 686328 46548 686398
rect 46208 685838 46218 685908
rect 46288 685838 46298 685908
rect 46224 685728 46230 685838
rect 46264 685728 46270 685838
rect 46208 685658 46218 685728
rect 46288 685658 46298 685728
rect 45966 685618 46012 685630
rect 46224 685630 46230 685658
rect 46264 685630 46270 685658
rect 46224 685618 46270 685630
rect 46482 685630 46488 686328
rect 46522 685630 46528 686328
rect 46740 685908 46746 686606
rect 46780 685908 46786 686606
rect 46998 686606 47044 686618
rect 46998 686578 47004 686606
rect 47038 686578 47044 686606
rect 46978 686508 46988 686578
rect 47058 686508 47068 686578
rect 46998 686398 47004 686508
rect 47038 686398 47044 686508
rect 46978 686328 46988 686398
rect 47058 686328 47068 686398
rect 46718 685838 46728 685908
rect 46798 685838 46808 685908
rect 46740 685728 46746 685838
rect 46780 685728 46786 685838
rect 46718 685658 46728 685728
rect 46798 685658 46808 685728
rect 46482 685618 46528 685630
rect 46740 685630 46746 685658
rect 46780 685630 46786 685658
rect 46740 685618 46786 685630
rect 46998 685630 47004 686328
rect 47038 685630 47044 686328
rect 46998 685618 47044 685630
rect 43098 685588 43108 685618
rect 43088 685538 43108 685588
rect 43098 685508 43108 685538
rect 43218 685588 43228 685618
rect 43348 685588 43358 685618
rect 43218 685538 43358 685588
rect 43218 685508 43228 685538
rect 43348 685508 43358 685538
rect 43468 685588 43478 685618
rect 47498 685588 47508 685618
rect 43468 685580 47508 685588
rect 43468 685546 43970 685580
rect 44138 685546 44228 685580
rect 44396 685546 44486 685580
rect 44654 685546 44744 685580
rect 44912 685546 45002 685580
rect 45170 685546 45260 685580
rect 45428 685546 45518 685580
rect 45686 685546 45776 685580
rect 45944 685546 46034 685580
rect 46202 685546 46292 685580
rect 46460 685546 46550 685580
rect 46718 685546 46808 685580
rect 46976 685546 47508 685580
rect 43468 685538 47508 685546
rect 43468 685508 43478 685538
rect 47498 685508 47508 685538
rect 47618 685588 47628 685618
rect 47748 685588 47758 685618
rect 47618 685538 47758 685588
rect 47618 685508 47628 685538
rect 47748 685508 47758 685538
rect 47868 685588 47878 685618
rect 47868 685538 47888 685588
rect 47868 685508 47878 685538
rect 45338 685484 45348 685488
rect 44639 685478 45348 685484
rect 45598 685484 45608 685488
rect 45598 685478 46307 685484
rect 44639 685444 44651 685478
rect 46295 685444 46307 685478
rect 44639 685438 45348 685444
rect 45338 685278 45348 685438
rect 44512 685272 45348 685278
rect 45598 685438 46307 685444
rect 45598 685278 45608 685438
rect 45598 685272 46438 685278
rect 44512 685238 44524 685272
rect 46426 685238 46438 685272
rect 44512 685232 46438 685238
rect 45338 685228 45608 685232
rect 43098 685178 43108 685208
rect 43088 685128 43108 685178
rect 43098 685098 43108 685128
rect 43218 685178 43228 685208
rect 43348 685178 43358 685208
rect 43218 685128 43358 685178
rect 43218 685098 43228 685128
rect 43348 685098 43358 685128
rect 43468 685178 43478 685208
rect 47498 685178 47508 685208
rect 43468 685170 47508 685178
rect 43468 685136 43714 685170
rect 43882 685136 43972 685170
rect 44140 685136 44230 685170
rect 44398 685136 44488 685170
rect 44656 685136 44746 685170
rect 44914 685136 45004 685170
rect 45172 685136 45262 685170
rect 45430 685136 45520 685170
rect 45688 685136 45778 685170
rect 45946 685136 46036 685170
rect 46204 685136 46294 685170
rect 46462 685136 46552 685170
rect 46720 685136 46810 685170
rect 46978 685136 47068 685170
rect 47236 685136 47508 685170
rect 43468 685128 47508 685136
rect 43468 685098 43478 685128
rect 47498 685098 47508 685128
rect 47618 685178 47628 685208
rect 47748 685178 47758 685208
rect 47618 685128 47758 685178
rect 47618 685098 47628 685128
rect 47748 685098 47758 685128
rect 47868 685178 47878 685208
rect 47868 685128 47888 685178
rect 47868 685098 47878 685128
rect 43646 685086 43692 685098
rect 43646 685058 43652 685086
rect 43686 685058 43692 685086
rect 43904 685086 43950 685098
rect 43628 684988 43638 685058
rect 43708 684988 43718 685058
rect 43646 684878 43652 684988
rect 43686 684878 43692 684988
rect 43628 684808 43638 684878
rect 43708 684808 43718 684878
rect 43646 684110 43652 684808
rect 43686 684110 43692 684808
rect 43904 684388 43910 685086
rect 43944 684388 43950 685086
rect 44162 685086 44208 685098
rect 44162 685058 44168 685086
rect 44202 685058 44208 685086
rect 44420 685086 44466 685098
rect 44138 684988 44148 685058
rect 44218 684988 44228 685058
rect 44162 684878 44168 684988
rect 44202 684878 44208 684988
rect 44138 684808 44148 684878
rect 44218 684808 44228 684878
rect 43888 684318 43898 684388
rect 43968 684318 43978 684388
rect 43904 684208 43910 684318
rect 43944 684208 43950 684318
rect 43888 684138 43898 684208
rect 43968 684138 43978 684208
rect 43646 684098 43692 684110
rect 43904 684110 43910 684138
rect 43944 684110 43950 684138
rect 43904 684098 43950 684110
rect 44162 684110 44168 684808
rect 44202 684110 44208 684808
rect 44420 684388 44426 685086
rect 44460 684388 44466 685086
rect 44678 685086 44724 685098
rect 44678 685058 44684 685086
rect 44718 685058 44724 685086
rect 44936 685086 44982 685098
rect 44658 684988 44668 685058
rect 44738 684988 44748 685058
rect 44678 684878 44684 684988
rect 44718 684878 44724 684988
rect 44658 684808 44668 684878
rect 44738 684808 44748 684878
rect 44398 684318 44408 684388
rect 44478 684318 44488 684388
rect 44420 684208 44426 684318
rect 44460 684208 44466 684318
rect 44398 684138 44408 684208
rect 44478 684138 44488 684208
rect 44162 684098 44208 684110
rect 44420 684110 44426 684138
rect 44460 684110 44466 684138
rect 44420 684098 44466 684110
rect 44678 684110 44684 684808
rect 44718 684110 44724 684808
rect 44936 684388 44942 685086
rect 44976 684388 44982 685086
rect 45194 685086 45240 685098
rect 45194 685058 45200 685086
rect 45234 685058 45240 685086
rect 45452 685086 45498 685098
rect 45178 684988 45188 685058
rect 45258 684988 45268 685058
rect 45194 684878 45200 684988
rect 45234 684878 45240 684988
rect 45178 684808 45188 684878
rect 45258 684808 45268 684878
rect 44918 684318 44928 684388
rect 44998 684318 45008 684388
rect 44936 684208 44942 684318
rect 44976 684208 44982 684318
rect 44918 684138 44928 684208
rect 44998 684138 45008 684208
rect 44678 684098 44724 684110
rect 44936 684110 44942 684138
rect 44976 684110 44982 684138
rect 44936 684098 44982 684110
rect 45194 684110 45200 684808
rect 45234 684110 45240 684808
rect 45452 684388 45458 685086
rect 45492 684388 45498 685086
rect 45710 685086 45756 685098
rect 45710 685058 45716 685086
rect 45750 685058 45756 685086
rect 45968 685086 46014 685098
rect 45688 684988 45698 685058
rect 45768 684988 45778 685058
rect 45710 684878 45716 684988
rect 45750 684878 45756 684988
rect 45688 684808 45698 684878
rect 45768 684808 45778 684878
rect 45428 684318 45438 684388
rect 45508 684318 45518 684388
rect 45452 684208 45458 684318
rect 45492 684208 45498 684318
rect 45428 684138 45438 684208
rect 45508 684138 45518 684208
rect 45194 684098 45240 684110
rect 45452 684110 45458 684138
rect 45492 684110 45498 684138
rect 45452 684098 45498 684110
rect 45710 684110 45716 684808
rect 45750 684110 45756 684808
rect 45968 684388 45974 685086
rect 46008 684388 46014 685086
rect 46226 685086 46272 685098
rect 46226 685058 46232 685086
rect 46266 685058 46272 685086
rect 46484 685086 46530 685098
rect 46208 684988 46218 685058
rect 46288 684988 46298 685058
rect 46226 684878 46232 684988
rect 46266 684878 46272 684988
rect 46208 684808 46218 684878
rect 46288 684808 46298 684878
rect 45948 684318 45958 684388
rect 46028 684318 46038 684388
rect 45968 684208 45974 684318
rect 46008 684208 46014 684318
rect 45948 684138 45958 684208
rect 46028 684138 46038 684208
rect 45710 684098 45756 684110
rect 45968 684110 45974 684138
rect 46008 684110 46014 684138
rect 45968 684098 46014 684110
rect 46226 684110 46232 684808
rect 46266 684110 46272 684808
rect 46484 684388 46490 685086
rect 46524 684388 46530 685086
rect 46742 685086 46788 685098
rect 46742 685058 46748 685086
rect 46782 685058 46788 685086
rect 47000 685086 47046 685098
rect 46718 684988 46728 685058
rect 46798 684988 46808 685058
rect 46742 684878 46748 684988
rect 46782 684878 46788 684988
rect 46718 684808 46728 684878
rect 46798 684808 46808 684878
rect 46468 684318 46478 684388
rect 46548 684318 46558 684388
rect 46484 684208 46490 684318
rect 46524 684208 46530 684318
rect 46468 684138 46478 684208
rect 46548 684138 46558 684208
rect 46226 684098 46272 684110
rect 46484 684110 46490 684138
rect 46524 684110 46530 684138
rect 46484 684098 46530 684110
rect 46742 684110 46748 684808
rect 46782 684110 46788 684808
rect 47000 684388 47006 685086
rect 47040 684388 47046 685086
rect 47258 685086 47304 685098
rect 47258 685058 47264 685086
rect 47298 685058 47304 685086
rect 47238 684988 47248 685058
rect 47318 684988 47328 685058
rect 47258 684878 47264 684988
rect 47298 684878 47304 684988
rect 47238 684808 47248 684878
rect 47318 684808 47328 684878
rect 46978 684318 46988 684388
rect 47058 684318 47068 684388
rect 47000 684208 47006 684318
rect 47040 684208 47046 684318
rect 46978 684138 46988 684208
rect 47058 684138 47068 684208
rect 46742 684098 46788 684110
rect 47000 684110 47006 684138
rect 47040 684110 47046 684138
rect 47000 684098 47046 684110
rect 47258 684110 47264 684808
rect 47298 684110 47304 684808
rect 47258 684098 47304 684110
rect 43098 684068 43108 684098
rect 43088 684018 43108 684068
rect 43098 683988 43108 684018
rect 43218 684068 43228 684098
rect 43348 684068 43358 684098
rect 43218 684018 43358 684068
rect 43218 683988 43228 684018
rect 43348 683988 43358 684018
rect 43468 684068 43478 684098
rect 47498 684068 47508 684098
rect 43468 684060 47508 684068
rect 43468 684026 43714 684060
rect 43882 684026 43972 684060
rect 44140 684026 44230 684060
rect 44398 684026 44488 684060
rect 44656 684026 44746 684060
rect 44914 684026 45004 684060
rect 45172 684026 45262 684060
rect 45430 684026 45520 684060
rect 45688 684026 45778 684060
rect 45946 684026 46036 684060
rect 46204 684026 46294 684060
rect 46462 684026 46552 684060
rect 46720 684026 46810 684060
rect 46978 684026 47068 684060
rect 47236 684026 47508 684060
rect 43468 684018 47508 684026
rect 43468 683988 43478 684018
rect 47498 683988 47508 684018
rect 47618 684068 47628 684098
rect 47748 684068 47758 684098
rect 47618 684018 47758 684068
rect 47618 683988 47628 684018
rect 47748 683988 47758 684018
rect 47868 684068 47878 684098
rect 47868 684018 47888 684068
rect 47868 683988 47878 684018
rect 44512 683958 46438 683964
rect 44512 683924 44524 683958
rect 46426 683924 46438 683958
rect 44512 683918 45348 683924
rect 45338 683708 45348 683918
rect 45598 683918 46438 683924
rect 45598 683708 45608 683918
rect 42296 683078 42480 683084
rect 43296 683078 43480 683084
rect 44776 683078 44960 683084
rect 45996 683078 46180 683084
rect 47456 683078 47640 683084
rect 48516 683078 48700 683084
rect 41868 682918 42308 683078
rect 42468 682918 43308 683078
rect 43468 682918 44788 683078
rect 44948 682918 46008 683078
rect 46168 682918 47468 683078
rect 47628 682918 48528 683078
rect 48688 682918 49068 683078
rect 41868 682870 49068 682918
rect 41868 682836 41891 682870
rect 42867 682858 43127 682870
rect 42867 682836 42888 682858
rect 41792 682808 41838 682820
rect 41868 682818 42888 682836
rect 43108 682836 43127 682858
rect 44103 682858 44363 682870
rect 44103 682836 44128 682858
rect 41792 682640 41798 682808
rect 41832 682768 41838 682808
rect 42920 682808 42966 682820
rect 42920 682768 42926 682808
rect 41832 682640 42926 682768
rect 42960 682768 42966 682808
rect 43028 682808 43074 682820
rect 43108 682818 44128 682836
rect 44348 682836 44363 682858
rect 45339 682858 45599 682870
rect 45339 682836 45351 682858
rect 44348 682830 45351 682836
rect 45587 682836 45599 682858
rect 46575 682858 46835 682870
rect 46575 682836 46588 682858
rect 45587 682830 46588 682836
rect 46823 682836 46835 682858
rect 47811 682858 48071 682870
rect 47811 682836 47828 682858
rect 46823 682830 47828 682836
rect 43028 682768 43034 682808
rect 42960 682640 43034 682768
rect 43068 682768 43074 682808
rect 44156 682808 44202 682820
rect 44156 682768 44162 682808
rect 43068 682758 44162 682768
rect 43068 682688 43698 682758
rect 43768 682688 43938 682758
rect 44008 682688 44162 682758
rect 43068 682640 44162 682688
rect 44196 682768 44202 682808
rect 44264 682808 44310 682820
rect 44348 682818 45348 682830
rect 44264 682768 44270 682808
rect 44196 682640 44270 682768
rect 44304 682768 44310 682808
rect 45392 682808 45438 682820
rect 45392 682768 45398 682808
rect 44304 682640 45398 682768
rect 45432 682768 45438 682808
rect 45500 682808 45546 682820
rect 45588 682818 46588 682830
rect 45500 682768 45506 682808
rect 45432 682640 45506 682768
rect 45540 682768 45546 682808
rect 46628 682808 46674 682820
rect 46628 682768 46634 682808
rect 45540 682640 46634 682768
rect 46668 682768 46674 682808
rect 46736 682808 46782 682820
rect 46828 682818 47828 682830
rect 48048 682836 48071 682858
rect 49047 682836 49068 682870
rect 46736 682768 46742 682808
rect 46668 682640 46742 682768
rect 46776 682768 46782 682808
rect 47864 682808 47910 682820
rect 47864 682768 47870 682808
rect 46776 682758 47870 682768
rect 46776 682688 46898 682758
rect 46968 682688 47118 682758
rect 47188 682688 47870 682758
rect 46776 682640 47870 682688
rect 47904 682768 47910 682808
rect 47972 682808 48018 682820
rect 48048 682818 49068 682836
rect 47972 682768 47978 682808
rect 47904 682640 47978 682768
rect 48012 682768 48018 682808
rect 49100 682808 49146 682820
rect 49100 682768 49106 682808
rect 48012 682640 49106 682768
rect 49140 682640 49146 682808
rect 41792 682628 49146 682640
rect 41798 682612 49146 682628
rect 41798 682578 41891 682612
rect 42867 682578 43127 682612
rect 44103 682578 44363 682612
rect 45339 682578 45599 682612
rect 46575 682578 46835 682612
rect 47811 682578 48071 682612
rect 49047 682578 49146 682612
rect 41798 682556 49146 682578
rect 42296 682498 42480 682504
rect 43296 682498 43480 682504
rect 44776 682498 44960 682504
rect 45996 682498 46180 682504
rect 47456 682498 47640 682504
rect 48516 682498 48700 682504
rect 41868 682338 42308 682498
rect 42468 682338 43308 682498
rect 43468 682338 44788 682498
rect 44948 682338 46008 682498
rect 46168 682338 47468 682498
rect 47628 682338 48528 682498
rect 48688 682338 49068 682498
rect 41868 682280 49068 682338
rect 41868 682258 41891 682280
rect 41879 682246 41891 682258
rect 42867 682268 43127 682280
rect 42867 682246 42879 682268
rect 41879 682240 42879 682246
rect 43115 682246 43127 682268
rect 44103 682268 44363 682280
rect 44103 682246 44115 682268
rect 43115 682240 44115 682246
rect 44351 682246 44363 682268
rect 45339 682268 45599 682280
rect 45339 682246 45351 682268
rect 44351 682240 45351 682246
rect 45587 682246 45599 682268
rect 46575 682268 46835 682280
rect 46575 682246 46587 682268
rect 45587 682240 46587 682246
rect 46823 682246 46835 682268
rect 47811 682268 48071 682280
rect 47811 682246 47823 682268
rect 46823 682240 47823 682246
rect 48059 682246 48071 682268
rect 49047 682258 49068 682280
rect 49047 682246 49059 682258
rect 48059 682240 49059 682246
rect 41792 682218 41838 682230
rect 41792 682050 41798 682218
rect 41832 682178 41838 682218
rect 42920 682218 42966 682230
rect 42920 682178 42926 682218
rect 41832 682088 42926 682178
rect 41832 682050 41838 682088
rect 41792 682038 41838 682050
rect 42920 682050 42926 682088
rect 42960 682178 42966 682218
rect 43028 682218 43074 682230
rect 43028 682178 43034 682218
rect 42960 682088 43034 682178
rect 42960 682050 42966 682088
rect 42920 682038 42966 682050
rect 43028 682050 43034 682088
rect 43068 682178 43074 682218
rect 44156 682218 44202 682230
rect 44156 682178 44162 682218
rect 43068 682168 44162 682178
rect 43068 682098 43698 682168
rect 43768 682098 43938 682168
rect 44008 682098 44162 682168
rect 43068 682088 44162 682098
rect 43068 682050 43074 682088
rect 43028 682038 43074 682050
rect 44156 682050 44162 682088
rect 44196 682178 44202 682218
rect 44264 682218 44310 682230
rect 44264 682178 44270 682218
rect 44196 682088 44270 682178
rect 44196 682050 44202 682088
rect 44156 682038 44202 682050
rect 44264 682050 44270 682088
rect 44304 682178 44310 682218
rect 45392 682218 45438 682230
rect 45392 682178 45398 682218
rect 44304 682088 45398 682178
rect 44304 682050 44310 682088
rect 44264 682038 44310 682050
rect 45392 682050 45398 682088
rect 45432 682178 45438 682218
rect 45500 682218 45546 682230
rect 45500 682178 45506 682218
rect 45432 682088 45506 682178
rect 45432 682050 45438 682088
rect 45392 682038 45438 682050
rect 45500 682050 45506 682088
rect 45540 682178 45546 682218
rect 46628 682218 46674 682230
rect 46628 682178 46634 682218
rect 45540 682088 46634 682178
rect 45540 682050 45546 682088
rect 45500 682038 45546 682050
rect 46628 682050 46634 682088
rect 46668 682178 46674 682218
rect 46736 682218 46782 682230
rect 46736 682178 46742 682218
rect 46668 682088 46742 682178
rect 46668 682050 46674 682088
rect 46628 682038 46674 682050
rect 46736 682050 46742 682088
rect 46776 682178 46782 682218
rect 47864 682218 47910 682230
rect 47864 682178 47870 682218
rect 46776 682168 47870 682178
rect 46776 682098 46898 682168
rect 46968 682098 47118 682168
rect 47188 682098 47870 682168
rect 46776 682088 47870 682098
rect 46776 682050 46782 682088
rect 46736 682038 46782 682050
rect 47864 682050 47870 682088
rect 47904 682178 47910 682218
rect 47972 682218 48018 682230
rect 47972 682178 47978 682218
rect 47904 682088 47978 682178
rect 47904 682050 47910 682088
rect 47864 682038 47910 682050
rect 47972 682050 47978 682088
rect 48012 682178 48018 682218
rect 49100 682218 49146 682230
rect 49100 682178 49106 682218
rect 48012 682088 49106 682178
rect 48012 682050 48018 682088
rect 47972 682038 48018 682050
rect 49100 682050 49106 682088
rect 49140 682178 49146 682218
rect 49140 682088 49148 682178
rect 49140 682050 49146 682088
rect 49100 682038 49146 682050
rect 41874 682022 42879 682028
rect 41874 681988 41891 682022
rect 42867 682008 42879 682022
rect 43115 682022 44115 682028
rect 43115 682008 43127 682022
rect 42867 681988 43127 682008
rect 44103 682008 44115 682022
rect 44351 682022 45351 682028
rect 44351 682008 44363 682022
rect 45339 682008 45351 682022
rect 45587 682022 46587 682028
rect 45587 682008 45599 682022
rect 46575 682008 46587 682022
rect 46823 682022 47823 682028
rect 46823 682008 46835 682022
rect 44103 681988 44363 682008
rect 45339 681988 45599 682008
rect 46575 681988 46835 682008
rect 47811 682008 47823 682022
rect 48059 682022 49068 682028
rect 48059 682008 48071 682022
rect 47811 681988 48071 682008
rect 49047 681988 49068 682022
rect 41874 681938 44908 681988
rect 44978 681938 45018 681988
rect 45088 681938 45848 681988
rect 45918 681938 45958 681988
rect 46028 681938 49068 681988
rect 41874 681928 49068 681938
rect 44568 681490 46388 681518
rect 44568 681456 44656 681490
rect 44882 681456 45124 681490
rect 45350 681456 45592 681490
rect 45818 681456 46060 681490
rect 46286 681456 46388 681490
rect 44568 681448 46388 681456
rect 44568 681440 44908 681448
rect 44566 681428 44908 681440
rect 44566 681260 44572 681428
rect 44606 681378 44908 681428
rect 44978 681378 45018 681448
rect 45088 681438 46388 681448
rect 45088 681428 45848 681438
rect 45088 681378 45400 681428
rect 44606 681288 44932 681378
rect 44606 681260 44612 681288
rect 44566 681248 44612 681260
rect 44923 681260 44932 681288
rect 44966 681260 45040 681378
rect 45074 681288 45400 681378
rect 45074 681260 45080 681288
rect 44923 681248 45080 681260
rect 45393 681260 45400 681288
rect 45434 681260 45508 681428
rect 45542 681368 45848 681428
rect 45918 681368 45958 681438
rect 46028 681428 46388 681438
rect 46028 681368 46336 681428
rect 45542 681288 45868 681368
rect 45542 681260 45548 681288
rect 45393 681248 45548 681260
rect 45858 681260 45868 681288
rect 45902 681260 45976 681368
rect 46010 681288 46336 681368
rect 46010 681260 46018 681288
rect 45858 681248 46018 681260
rect 46330 681260 46336 681288
rect 46370 681368 46388 681428
rect 46370 681260 46376 681368
rect 46330 681248 46376 681260
rect 44644 681232 44894 681238
rect 44644 681218 44656 681232
rect 44638 681198 44656 681218
rect 44882 681218 44894 681232
rect 45112 681232 45362 681238
rect 45112 681218 45124 681232
rect 44882 681198 45124 681218
rect 45350 681218 45362 681232
rect 45580 681232 45830 681238
rect 45580 681218 45592 681232
rect 45350 681198 45592 681218
rect 45818 681218 45830 681232
rect 46048 681232 46298 681238
rect 46048 681218 46060 681232
rect 45818 681198 46060 681218
rect 46286 681218 46298 681232
rect 46286 681198 46308 681218
rect 44638 681178 46308 681198
rect 44598 681124 46308 681178
rect 44586 681118 46320 681124
rect 44586 680968 44598 681118
rect 44818 681108 45148 681118
rect 44818 680968 44830 681108
rect 44586 680962 44830 680968
rect 45136 680968 45148 681108
rect 45368 681108 45568 681118
rect 45368 680968 45380 681108
rect 45136 680962 45380 680968
rect 45556 680968 45568 681108
rect 45788 681108 46088 681118
rect 45788 680968 45800 681108
rect 45556 680962 45800 680968
rect 46076 680968 46088 681108
rect 46308 680968 46320 681118
rect 46076 680962 46320 680968
rect 43678 680928 44028 680948
rect 43678 680858 43698 680928
rect 43768 680858 43938 680928
rect 44008 680908 47208 680928
rect 44008 680865 46908 680908
rect 44008 680858 44872 680865
rect 43678 680838 44872 680858
rect 43678 680768 43698 680838
rect 43768 680768 43938 680838
rect 44008 680831 44872 680838
rect 45348 680831 45590 680865
rect 46066 680838 46908 680865
rect 46978 680838 47118 680908
rect 47188 680838 47208 680908
rect 46066 680831 47208 680838
rect 44008 680818 47208 680831
rect 44008 680803 46908 680818
rect 44008 680768 44788 680803
rect 43678 680748 44788 680768
rect 44782 680735 44788 680748
rect 44822 680748 45398 680803
rect 44822 680735 44828 680748
rect 44782 680723 44828 680735
rect 45392 680735 45398 680748
rect 45432 680748 45506 680803
rect 45432 680735 45438 680748
rect 45392 680723 45438 680735
rect 45500 680735 45506 680748
rect 45540 680748 46116 680803
rect 45540 680735 45546 680748
rect 45500 680723 45546 680735
rect 46110 680735 46116 680748
rect 46150 680748 46908 680803
rect 46978 680748 47118 680818
rect 47188 680748 47208 680818
rect 46150 680735 46156 680748
rect 46110 680723 46156 680735
rect 46878 680718 47208 680748
rect 44860 680707 45360 680713
rect 44860 680693 44872 680707
rect 44848 680678 44872 680693
rect 45348 680693 45360 680707
rect 45578 680707 46078 680713
rect 45578 680693 45590 680707
rect 44838 680673 44872 680678
rect 45348 680673 45590 680693
rect 46066 680693 46078 680707
rect 46066 680678 46083 680693
rect 46066 680673 46088 680678
rect 44838 680618 44908 680673
rect 44978 680618 45018 680673
rect 45088 680618 45848 680673
rect 45918 680618 45958 680673
rect 46028 680618 46088 680673
rect 44838 680608 46088 680618
rect 42356 680568 42560 680574
rect 42356 680438 42368 680568
rect 42548 680438 42560 680568
rect 42356 680432 42560 680438
rect 43356 680568 43560 680574
rect 43356 680438 43368 680568
rect 43548 680438 43560 680568
rect 45146 680568 45350 680574
rect 43356 680432 43560 680438
rect 44426 680558 44630 680564
rect 44426 680428 44438 680558
rect 44618 680428 44630 680558
rect 45146 680438 45158 680568
rect 45338 680438 45350 680568
rect 45146 680432 45350 680438
rect 45586 680568 45790 680574
rect 45586 680438 45598 680568
rect 45778 680438 45790 680568
rect 45586 680432 45790 680438
rect 46356 680568 46560 680574
rect 46356 680438 46368 680568
rect 46548 680438 46560 680568
rect 46356 680432 46560 680438
rect 47336 680558 47540 680564
rect 44426 680422 44630 680428
rect 47336 680428 47348 680558
rect 47528 680428 47540 680558
rect 47336 680422 47540 680428
rect 48476 680558 48680 680564
rect 48476 680428 48488 680558
rect 48668 680428 48680 680558
rect 48476 680422 48680 680428
rect 41928 680388 49018 680393
rect 41928 680346 43698 680388
rect 41923 680340 43698 680346
rect 43768 680340 43938 680388
rect 44008 680340 46898 680388
rect 46968 680340 47118 680388
rect 47188 680340 49018 680388
rect 41923 680306 41935 680340
rect 42911 680318 43153 680340
rect 44129 680318 44371 680340
rect 42911 680306 42923 680318
rect 41923 680300 42923 680306
rect 43141 680306 43153 680318
rect 44129 680306 44141 680318
rect 43141 680300 44141 680306
rect 44359 680306 44371 680318
rect 45347 680318 45589 680340
rect 45347 680306 45359 680318
rect 44359 680300 45359 680306
rect 45577 680306 45589 680318
rect 46565 680318 46807 680340
rect 47783 680318 48025 680340
rect 46565 680306 46577 680318
rect 45577 680300 46577 680306
rect 46795 680306 46807 680318
rect 47783 680306 47795 680318
rect 46795 680300 47795 680306
rect 48013 680306 48025 680318
rect 49001 680318 49018 680340
rect 49001 680306 49013 680318
rect 48013 680300 49013 680306
rect 41845 680278 41891 680290
rect 41845 680110 41851 680278
rect 41885 680243 41891 680278
rect 42955 680278 43001 680290
rect 42955 680243 42961 680278
rect 41885 680158 42961 680243
rect 41885 680110 41891 680158
rect 41845 680098 41891 680110
rect 42955 680110 42961 680158
rect 42995 680243 43001 680278
rect 43063 680278 43109 680290
rect 43063 680243 43069 680278
rect 42995 680158 43069 680243
rect 42995 680110 43001 680158
rect 42955 680098 43001 680110
rect 43063 680110 43069 680158
rect 43103 680243 43109 680278
rect 44173 680278 44219 680290
rect 44173 680243 44179 680278
rect 43103 680158 44179 680243
rect 43103 680110 43109 680158
rect 43063 680098 43109 680110
rect 44173 680110 44179 680158
rect 44213 680243 44219 680278
rect 44281 680278 44327 680290
rect 44281 680243 44287 680278
rect 44213 680158 44287 680243
rect 44213 680110 44219 680158
rect 44173 680098 44219 680110
rect 44281 680110 44287 680158
rect 44321 680243 44327 680278
rect 45391 680278 45437 680290
rect 45391 680243 45397 680278
rect 44321 680238 45397 680243
rect 44321 680168 44908 680238
rect 44978 680168 45018 680238
rect 45088 680168 45397 680238
rect 44321 680158 45397 680168
rect 44321 680110 44327 680158
rect 44281 680098 44327 680110
rect 45391 680110 45397 680158
rect 45431 680243 45437 680278
rect 45499 680278 45545 680290
rect 45499 680243 45505 680278
rect 45431 680158 45505 680243
rect 45431 680110 45437 680158
rect 45391 680098 45437 680110
rect 45499 680110 45505 680158
rect 45539 680243 45545 680278
rect 46609 680278 46655 680290
rect 46609 680243 46615 680278
rect 45539 680238 46615 680243
rect 45539 680168 45848 680238
rect 45918 680168 45958 680238
rect 46028 680168 46615 680238
rect 45539 680158 46615 680168
rect 45539 680110 45545 680158
rect 45499 680098 45545 680110
rect 46609 680110 46615 680158
rect 46649 680243 46655 680278
rect 46717 680278 46763 680290
rect 46717 680243 46723 680278
rect 46649 680158 46723 680243
rect 46649 680110 46655 680158
rect 46609 680098 46655 680110
rect 46717 680110 46723 680158
rect 46757 680243 46763 680278
rect 47827 680278 47873 680290
rect 47827 680243 47833 680278
rect 46757 680158 47833 680243
rect 46757 680110 46763 680158
rect 46717 680098 46763 680110
rect 47827 680110 47833 680158
rect 47867 680243 47873 680278
rect 47935 680278 47981 680290
rect 47935 680243 47941 680278
rect 47867 680158 47941 680243
rect 47867 680110 47873 680158
rect 47827 680098 47873 680110
rect 47935 680110 47941 680158
rect 47975 680243 47981 680278
rect 49045 680278 49091 680290
rect 49045 680243 49051 680278
rect 47975 680158 49051 680243
rect 47975 680110 47981 680158
rect 47935 680098 47981 680110
rect 49045 680110 49051 680158
rect 49085 680110 49091 680278
rect 49045 680098 49091 680110
rect 41923 680082 42923 680088
rect 41923 680048 41935 680082
rect 42911 680068 42923 680082
rect 43141 680082 44141 680088
rect 43141 680068 43153 680082
rect 42911 680048 43153 680068
rect 44129 680068 44141 680082
rect 44359 680082 45359 680088
rect 44359 680068 44371 680082
rect 44129 680048 44371 680068
rect 45347 680068 45359 680082
rect 45577 680082 46577 680088
rect 45577 680068 45589 680082
rect 45347 680048 45589 680068
rect 46565 680068 46577 680082
rect 46795 680082 47795 680088
rect 46795 680068 46807 680082
rect 46565 680048 46807 680068
rect 47783 680068 47795 680082
rect 48013 680082 49013 680088
rect 48013 680068 48025 680082
rect 47783 680048 48025 680068
rect 49001 680068 49013 680082
rect 49001 680048 49018 680068
rect 41923 680042 49018 680048
rect 41928 679993 49018 680042
rect 43268 679698 43678 679993
rect 44568 679698 44968 679993
rect 45868 679698 46268 679993
rect 47268 679698 47668 679993
rect 42468 679590 48468 679698
rect 42468 679193 42641 679590
rect 43755 679193 44151 679590
rect 45265 679584 48468 679590
rect 45265 679193 45661 679584
rect 42468 679187 45661 679193
rect 46775 679187 47181 679584
rect 48295 679187 48468 679584
rect 42468 679098 48468 679187
rect 42206 678658 42350 678664
rect 42206 678538 42218 678658
rect 42338 678538 42350 678658
rect 42206 678532 42350 678538
rect 48576 678658 48720 678664
rect 48576 678538 48588 678658
rect 48708 678538 48720 678658
rect 48576 678532 48720 678538
rect 42206 675658 42350 675664
rect 42206 675538 42218 675658
rect 42338 675538 42350 675658
rect 42206 675532 42350 675538
rect 48576 675658 48720 675664
rect 48576 675538 48588 675658
rect 48708 675538 48720 675658
rect 48576 675532 48720 675538
rect 42206 672658 42350 672664
rect 42206 672538 42218 672658
rect 42338 672538 42350 672658
rect 42206 672532 42350 672538
rect 48576 672658 48720 672664
rect 48576 672538 48588 672658
rect 48708 672538 48720 672658
rect 48576 672532 48720 672538
rect 42206 669658 42350 669664
rect 42206 669538 42218 669658
rect 42338 669538 42350 669658
rect 42206 669532 42350 669538
rect 48576 669658 48720 669664
rect 48576 669538 48588 669658
rect 48708 669538 48720 669658
rect 48576 669532 48720 669538
rect 42206 666658 42350 666664
rect 42206 666538 42218 666658
rect 42338 666538 42350 666658
rect 42206 666532 42350 666538
rect 48576 666658 48720 666664
rect 48576 666538 48588 666658
rect 48708 666538 48720 666658
rect 48576 666532 48720 666538
rect 42468 665359 48468 665398
rect 42468 665338 42641 665359
rect 43755 665338 44151 665359
rect 42468 664928 42608 665338
rect 43778 665328 44151 665338
rect 45265 665353 48468 665359
rect 45265 665328 45661 665353
rect 46775 665328 47181 665353
rect 48295 665328 48468 665353
rect 43778 664928 44128 665328
rect 42468 664918 44128 664928
rect 45298 664918 45648 665328
rect 46818 664918 47158 665328
rect 48328 664918 48468 665328
rect 42468 664898 48468 664918
<< via1 >>
rect 37738 694088 37808 694158
rect 37628 693978 37698 694048
rect 44798 694620 45068 694878
rect 45848 694620 46118 694878
rect 44798 694608 45068 694620
rect 45848 694608 46118 694620
rect 42278 694328 42294 694398
rect 42294 694328 42328 694398
rect 42328 694328 42348 694398
rect 42278 694088 42294 694158
rect 42294 694088 42328 694158
rect 42328 694088 42348 694158
rect 42588 694328 42610 694398
rect 42610 694328 42644 694398
rect 42644 694328 42658 694398
rect 42588 694088 42610 694158
rect 42610 694088 42644 694158
rect 42644 694088 42658 694158
rect 42428 693718 42452 693788
rect 42452 693718 42486 693788
rect 42486 693718 42498 693788
rect 42428 693478 42452 693548
rect 42452 693478 42486 693548
rect 42486 693478 42498 693548
rect 42908 694328 42926 694398
rect 42926 694328 42960 694398
rect 42960 694328 42978 694398
rect 42908 694088 42926 694158
rect 42926 694088 42960 694158
rect 42960 694088 42978 694158
rect 42748 693718 42768 693788
rect 42768 693718 42802 693788
rect 42802 693718 42818 693788
rect 42748 693478 42768 693548
rect 42768 693478 42802 693548
rect 42802 693478 42818 693548
rect 43228 694328 43242 694398
rect 43242 694328 43276 694398
rect 43276 694328 43298 694398
rect 43228 694088 43242 694158
rect 43242 694088 43276 694158
rect 43276 694088 43298 694158
rect 43068 693718 43084 693788
rect 43084 693718 43118 693788
rect 43118 693718 43138 693788
rect 43068 693478 43084 693548
rect 43084 693478 43118 693548
rect 43118 693478 43138 693548
rect 43538 694328 43558 694398
rect 43558 694328 43592 694398
rect 43592 694328 43608 694398
rect 43538 694088 43558 694158
rect 43558 694088 43592 694158
rect 43592 694088 43608 694158
rect 43378 693718 43400 693788
rect 43400 693718 43434 693788
rect 43434 693718 43448 693788
rect 43378 693478 43400 693548
rect 43400 693478 43434 693548
rect 43434 693478 43448 693548
rect 43858 694328 43874 694398
rect 43874 694328 43908 694398
rect 43908 694328 43928 694398
rect 43858 694088 43874 694158
rect 43874 694088 43908 694158
rect 43908 694088 43928 694158
rect 43698 693718 43716 693788
rect 43716 693718 43750 693788
rect 43750 693718 43768 693788
rect 43698 693478 43716 693548
rect 43716 693478 43750 693548
rect 43750 693478 43768 693548
rect 44168 694328 44190 694398
rect 44190 694328 44224 694398
rect 44224 694328 44238 694398
rect 44168 694088 44190 694158
rect 44190 694088 44224 694158
rect 44224 694088 44238 694158
rect 44018 693718 44032 693788
rect 44032 693718 44066 693788
rect 44066 693718 44088 693788
rect 44018 693478 44032 693548
rect 44032 693478 44066 693548
rect 44066 693478 44088 693548
rect 44488 694328 44506 694398
rect 44506 694328 44540 694398
rect 44540 694328 44558 694398
rect 44488 694088 44506 694158
rect 44506 694088 44540 694158
rect 44540 694088 44558 694158
rect 44328 693718 44348 693788
rect 44348 693718 44382 693788
rect 44382 693718 44398 693788
rect 44328 693478 44348 693548
rect 44348 693478 44382 693548
rect 44382 693478 44398 693548
rect 44808 694328 44822 694398
rect 44822 694328 44856 694398
rect 44856 694328 44878 694398
rect 44808 694088 44822 694158
rect 44822 694088 44856 694158
rect 44856 694088 44878 694158
rect 44648 693718 44664 693788
rect 44664 693718 44698 693788
rect 44698 693718 44718 693788
rect 44648 693478 44664 693548
rect 44664 693478 44698 693548
rect 44698 693478 44718 693548
rect 45118 694328 45138 694398
rect 45138 694328 45172 694398
rect 45172 694328 45188 694398
rect 45118 694088 45138 694158
rect 45138 694088 45172 694158
rect 45172 694088 45188 694158
rect 44958 693718 44980 693788
rect 44980 693718 45014 693788
rect 45014 693718 45028 693788
rect 44958 693478 44980 693548
rect 44980 693478 45014 693548
rect 45014 693478 45028 693548
rect 45438 694328 45454 694398
rect 45454 694328 45488 694398
rect 45488 694328 45508 694398
rect 45438 694088 45454 694158
rect 45454 694088 45488 694158
rect 45488 694088 45508 694158
rect 45278 693718 45296 693788
rect 45296 693718 45330 693788
rect 45330 693718 45348 693788
rect 45278 693478 45296 693548
rect 45296 693478 45330 693548
rect 45330 693478 45348 693548
rect 45748 694328 45770 694398
rect 45770 694328 45804 694398
rect 45804 694328 45818 694398
rect 45748 694088 45770 694158
rect 45770 694088 45804 694158
rect 45804 694088 45818 694158
rect 45598 693718 45612 693788
rect 45612 693718 45646 693788
rect 45646 693718 45668 693788
rect 45598 693478 45612 693548
rect 45612 693478 45646 693548
rect 45646 693478 45668 693548
rect 46068 694328 46086 694398
rect 46086 694328 46120 694398
rect 46120 694328 46138 694398
rect 46068 694088 46086 694158
rect 46086 694088 46120 694158
rect 46120 694088 46138 694158
rect 45908 693718 45928 693788
rect 45928 693718 45962 693788
rect 45962 693718 45978 693788
rect 45908 693478 45928 693548
rect 45928 693478 45962 693548
rect 45962 693478 45978 693548
rect 46388 694328 46402 694398
rect 46402 694328 46436 694398
rect 46436 694328 46458 694398
rect 46388 694088 46402 694158
rect 46402 694088 46436 694158
rect 46436 694088 46458 694158
rect 46228 693718 46244 693788
rect 46244 693718 46278 693788
rect 46278 693718 46298 693788
rect 46228 693478 46244 693548
rect 46244 693478 46278 693548
rect 46278 693478 46298 693548
rect 46698 694328 46718 694398
rect 46718 694328 46752 694398
rect 46752 694328 46768 694398
rect 46698 694088 46718 694158
rect 46718 694088 46752 694158
rect 46752 694088 46768 694158
rect 46548 693718 46560 693788
rect 46560 693718 46594 693788
rect 46594 693718 46618 693788
rect 46548 693478 46560 693548
rect 46560 693478 46594 693548
rect 46594 693478 46618 693548
rect 47018 694328 47034 694398
rect 47034 694328 47068 694398
rect 47068 694328 47088 694398
rect 47018 694088 47034 694158
rect 47034 694088 47068 694158
rect 47068 694088 47088 694158
rect 46858 693718 46876 693788
rect 46876 693718 46910 693788
rect 46910 693718 46928 693788
rect 46858 693478 46876 693548
rect 46876 693478 46910 693548
rect 46910 693478 46928 693548
rect 47338 694328 47350 694398
rect 47350 694328 47384 694398
rect 47384 694328 47408 694398
rect 47338 694088 47350 694158
rect 47350 694088 47384 694158
rect 47384 694088 47408 694158
rect 47178 693718 47192 693788
rect 47192 693718 47226 693788
rect 47226 693718 47248 693788
rect 47178 693478 47192 693548
rect 47192 693478 47226 693548
rect 47226 693478 47248 693548
rect 47648 694328 47666 694398
rect 47666 694328 47700 694398
rect 47700 694328 47718 694398
rect 47648 694088 47666 694158
rect 47666 694088 47700 694158
rect 47700 694088 47718 694158
rect 47488 693718 47508 693788
rect 47508 693718 47542 693788
rect 47542 693718 47558 693788
rect 47488 693478 47508 693548
rect 47508 693478 47542 693548
rect 47542 693478 47558 693548
rect 47968 694328 47982 694398
rect 47982 694328 48016 694398
rect 48016 694328 48038 694398
rect 47968 694088 47982 694158
rect 47982 694088 48016 694158
rect 48016 694088 48038 694158
rect 47808 693718 47824 693788
rect 47824 693718 47858 693788
rect 47858 693718 47878 693788
rect 47808 693478 47824 693548
rect 47824 693478 47858 693548
rect 47858 693478 47878 693548
rect 48278 694328 48298 694398
rect 48298 694328 48332 694398
rect 48332 694328 48348 694398
rect 48278 694088 48298 694158
rect 48298 694088 48332 694158
rect 48332 694088 48348 694158
rect 48128 693718 48140 693788
rect 48140 693718 48174 693788
rect 48174 693718 48198 693788
rect 48128 693478 48140 693548
rect 48140 693478 48174 693548
rect 48174 693478 48198 693548
rect 48598 694328 48614 694398
rect 48614 694328 48648 694398
rect 48648 694328 48668 694398
rect 48598 694088 48614 694158
rect 48614 694088 48648 694158
rect 48648 694088 48668 694158
rect 48438 693718 48456 693788
rect 48456 693718 48490 693788
rect 48490 693718 48508 693788
rect 43408 693356 43462 693378
rect 43462 693356 43488 693378
rect 47468 693356 47480 693378
rect 47480 693356 47548 693378
rect 43408 693298 43488 693356
rect 47468 693298 47548 693356
rect 44798 692968 45068 693238
rect 45848 692968 46118 693238
rect 39578 692598 39758 692698
rect 39998 692598 40178 692698
rect 43938 692658 43954 692728
rect 43954 692658 43988 692728
rect 43988 692658 44008 692728
rect 43938 692448 43954 692518
rect 43954 692448 43988 692518
rect 43988 692448 44008 692518
rect 43778 692018 43796 692088
rect 43796 692018 43830 692088
rect 43830 692018 43848 692088
rect 43778 691808 43796 691878
rect 43796 691808 43830 691878
rect 43830 691808 43848 691878
rect 44248 692658 44270 692728
rect 44270 692658 44304 692728
rect 44304 692658 44318 692728
rect 44248 692448 44270 692518
rect 44270 692448 44304 692518
rect 44304 692448 44318 692518
rect 44088 692018 44112 692088
rect 44112 692018 44146 692088
rect 44146 692018 44158 692088
rect 44088 691808 44112 691878
rect 44112 691808 44146 691878
rect 44146 691808 44158 691878
rect 44568 692658 44586 692728
rect 44586 692658 44620 692728
rect 44620 692658 44638 692728
rect 44568 692448 44586 692518
rect 44586 692448 44620 692518
rect 44620 692448 44638 692518
rect 44408 692018 44428 692088
rect 44428 692018 44462 692088
rect 44462 692018 44478 692088
rect 44408 691808 44428 691878
rect 44428 691808 44462 691878
rect 44462 691808 44478 691878
rect 44878 692658 44902 692728
rect 44902 692658 44936 692728
rect 44936 692658 44948 692728
rect 44878 692448 44902 692518
rect 44902 692448 44936 692518
rect 44936 692448 44948 692518
rect 44728 692018 44744 692088
rect 44744 692018 44778 692088
rect 44778 692018 44798 692088
rect 44728 691808 44744 691878
rect 44744 691808 44778 691878
rect 44778 691808 44798 691878
rect 45198 692658 45218 692728
rect 45218 692658 45252 692728
rect 45252 692658 45268 692728
rect 45198 692448 45218 692518
rect 45218 692448 45252 692518
rect 45252 692448 45268 692518
rect 45038 692018 45060 692088
rect 45060 692018 45094 692088
rect 45094 692018 45108 692088
rect 45038 691808 45060 691878
rect 45060 691808 45094 691878
rect 45094 691808 45108 691878
rect 45518 692658 45534 692728
rect 45534 692658 45568 692728
rect 45568 692658 45588 692728
rect 45518 692448 45534 692518
rect 45534 692448 45568 692518
rect 45568 692448 45588 692518
rect 45358 692018 45376 692088
rect 45376 692018 45410 692088
rect 45410 692018 45428 692088
rect 45358 691808 45376 691878
rect 45376 691808 45410 691878
rect 45410 691808 45428 691878
rect 45828 692658 45850 692728
rect 45850 692658 45884 692728
rect 45884 692658 45898 692728
rect 45828 692448 45850 692518
rect 45850 692448 45884 692518
rect 45884 692448 45898 692518
rect 45668 692018 45692 692088
rect 45692 692018 45726 692088
rect 45726 692018 45738 692088
rect 45668 691808 45692 691878
rect 45692 691808 45726 691878
rect 45726 691808 45738 691878
rect 46148 692658 46166 692728
rect 46166 692658 46200 692728
rect 46200 692658 46218 692728
rect 46148 692448 46166 692518
rect 46166 692448 46200 692518
rect 46200 692448 46218 692518
rect 45988 692018 46008 692088
rect 46008 692018 46042 692088
rect 46042 692018 46058 692088
rect 45988 691808 46008 691878
rect 46008 691808 46042 691878
rect 46042 691808 46058 691878
rect 46468 692658 46482 692728
rect 46482 692658 46516 692728
rect 46516 692658 46538 692728
rect 46468 692448 46482 692518
rect 46482 692448 46516 692518
rect 46516 692448 46538 692518
rect 46308 692018 46324 692088
rect 46324 692018 46358 692088
rect 46358 692018 46378 692088
rect 46308 691808 46324 691878
rect 46324 691808 46358 691878
rect 46358 691808 46378 691878
rect 46778 692658 46798 692728
rect 46798 692658 46832 692728
rect 46832 692658 46848 692728
rect 46778 692448 46798 692518
rect 46798 692448 46832 692518
rect 46832 692448 46848 692518
rect 46618 692018 46640 692088
rect 46640 692018 46674 692088
rect 46674 692018 46688 692088
rect 46618 691808 46640 691878
rect 46640 691808 46674 691878
rect 46674 691808 46688 691878
rect 47098 692658 47114 692728
rect 47114 692658 47148 692728
rect 47148 692658 47168 692728
rect 47098 692448 47114 692518
rect 47114 692448 47148 692518
rect 47148 692448 47168 692518
rect 46938 692018 46956 692088
rect 46956 692018 46990 692088
rect 46990 692018 47008 692088
rect 46938 691808 46956 691878
rect 46956 691808 46990 691878
rect 46990 691808 47008 691878
rect 53128 694088 53198 694158
rect 53238 693978 53308 694048
rect 50828 692598 51008 692698
rect 51248 692598 51428 692698
rect 44588 691618 44848 691628
rect 44588 691378 44848 691618
rect 44588 691368 44848 691378
rect 46088 691618 46348 691628
rect 46088 691378 46348 691618
rect 46088 691368 46348 691378
rect 43938 691108 43954 691178
rect 43954 691108 43988 691178
rect 43988 691108 44008 691178
rect 43938 690898 43954 690968
rect 43954 690898 43988 690968
rect 43988 690898 44008 690968
rect 43778 690478 43796 690548
rect 43796 690478 43830 690548
rect 43830 690478 43848 690548
rect 43778 690268 43796 690338
rect 43796 690268 43830 690338
rect 43830 690268 43848 690338
rect 44248 691108 44270 691178
rect 44270 691108 44304 691178
rect 44304 691108 44318 691178
rect 44248 690898 44270 690968
rect 44270 690898 44304 690968
rect 44304 690898 44318 690968
rect 44098 690478 44112 690548
rect 44112 690478 44146 690548
rect 44146 690478 44168 690548
rect 44098 690268 44112 690338
rect 44112 690268 44146 690338
rect 44146 690268 44168 690338
rect 44568 691108 44586 691178
rect 44586 691108 44620 691178
rect 44620 691108 44638 691178
rect 44568 690898 44586 690968
rect 44586 690898 44620 690968
rect 44620 690898 44638 690968
rect 44408 690478 44428 690548
rect 44428 690478 44462 690548
rect 44462 690478 44478 690548
rect 44408 690268 44428 690338
rect 44428 690268 44462 690338
rect 44462 690268 44478 690338
rect 44888 691108 44902 691178
rect 44902 691108 44936 691178
rect 44936 691108 44958 691178
rect 44888 690898 44902 690968
rect 44902 690898 44936 690968
rect 44936 690898 44958 690968
rect 44728 690478 44744 690548
rect 44744 690478 44778 690548
rect 44778 690478 44798 690548
rect 44728 690268 44744 690338
rect 44744 690268 44778 690338
rect 44778 690268 44798 690338
rect 45198 691108 45218 691178
rect 45218 691108 45252 691178
rect 45252 691108 45268 691178
rect 45198 690898 45218 690968
rect 45218 690898 45252 690968
rect 45252 690898 45268 690968
rect 45038 690478 45060 690548
rect 45060 690478 45094 690548
rect 45094 690478 45108 690548
rect 45038 690268 45060 690338
rect 45060 690268 45094 690338
rect 45094 690268 45108 690338
rect 45518 691108 45534 691178
rect 45534 691108 45568 691178
rect 45568 691108 45588 691178
rect 45518 690898 45534 690968
rect 45534 690898 45568 690968
rect 45568 690898 45588 690968
rect 45358 690478 45376 690548
rect 45376 690478 45410 690548
rect 45410 690478 45428 690548
rect 45358 690268 45376 690338
rect 45376 690268 45410 690338
rect 45410 690268 45428 690338
rect 45828 691108 45850 691178
rect 45850 691108 45884 691178
rect 45884 691108 45898 691178
rect 45828 690898 45850 690968
rect 45850 690898 45884 690968
rect 45884 690898 45898 690968
rect 45678 690478 45692 690548
rect 45692 690478 45726 690548
rect 45726 690478 45748 690548
rect 45678 690268 45692 690338
rect 45692 690268 45726 690338
rect 45726 690268 45748 690338
rect 46148 691108 46166 691178
rect 46166 691108 46200 691178
rect 46200 691108 46218 691178
rect 46148 690898 46166 690968
rect 46166 690898 46200 690968
rect 46200 690898 46218 690968
rect 45988 690478 46008 690548
rect 46008 690478 46042 690548
rect 46042 690478 46058 690548
rect 45988 690268 46008 690338
rect 46008 690268 46042 690338
rect 46042 690268 46058 690338
rect 46468 691108 46482 691178
rect 46482 691108 46516 691178
rect 46516 691108 46538 691178
rect 46468 690898 46482 690968
rect 46482 690898 46516 690968
rect 46516 690898 46538 690968
rect 46308 690478 46324 690548
rect 46324 690478 46358 690548
rect 46358 690478 46378 690548
rect 46308 690268 46324 690338
rect 46324 690268 46358 690338
rect 46358 690268 46378 690338
rect 46778 691108 46798 691178
rect 46798 691108 46832 691178
rect 46832 691108 46848 691178
rect 46778 690898 46798 690968
rect 46798 690898 46832 690968
rect 46832 690898 46848 690968
rect 46618 690478 46640 690548
rect 46640 690478 46674 690548
rect 46674 690478 46688 690548
rect 46618 690268 46640 690338
rect 46640 690268 46674 690338
rect 46674 690268 46688 690338
rect 47098 691108 47114 691178
rect 47114 691108 47148 691178
rect 47148 691108 47168 691178
rect 47098 690898 47114 690968
rect 47114 690898 47148 690968
rect 47148 690898 47168 690968
rect 46938 690478 46956 690548
rect 46956 690478 46990 690548
rect 46990 690478 47008 690548
rect 46938 690268 46956 690338
rect 46956 690268 46990 690338
rect 46990 690268 47008 690338
rect 45048 689548 45065 689618
rect 45065 689548 45099 689618
rect 45099 689548 45118 689618
rect 45048 689258 45065 689328
rect 45065 689258 45099 689328
rect 45099 689258 45118 689328
rect 44888 688988 44907 689058
rect 44907 688988 44941 689058
rect 44941 688988 44958 689058
rect 44888 688698 44907 688768
rect 44907 688698 44941 688768
rect 44941 688698 44958 688768
rect 45368 689548 45381 689618
rect 45381 689548 45415 689618
rect 45415 689548 45438 689618
rect 45368 689258 45381 689328
rect 45381 689258 45415 689328
rect 45415 689258 45438 689328
rect 45208 688988 45223 689058
rect 45223 688988 45257 689058
rect 45257 688988 45278 689058
rect 45208 688698 45223 688768
rect 45223 688698 45257 688768
rect 45257 688698 45278 688768
rect 45678 689548 45697 689618
rect 45697 689548 45731 689618
rect 45731 689548 45748 689618
rect 45678 689258 45697 689328
rect 45697 689258 45731 689328
rect 45731 689258 45748 689328
rect 45528 688988 45539 689058
rect 45539 688988 45573 689058
rect 45573 688988 45598 689058
rect 45528 688698 45539 688768
rect 45539 688698 45573 688768
rect 45573 688698 45598 688768
rect 45998 689548 46013 689618
rect 46013 689548 46047 689618
rect 46047 689548 46068 689618
rect 45998 689258 46013 689328
rect 46013 689258 46047 689328
rect 46047 689258 46068 689328
rect 45838 688988 45855 689058
rect 45855 688988 45889 689058
rect 45889 688988 45908 689058
rect 45838 688698 45855 688768
rect 45855 688698 45889 688768
rect 45889 688698 45908 688768
rect 47960 689100 48100 689220
rect 45348 688519 45608 688528
rect 45348 688485 45608 688519
rect 45348 688313 45608 688485
rect 45348 688279 45608 688313
rect 45348 688268 45608 688279
rect 43340 687560 43460 687720
rect 45048 688028 45065 688098
rect 45065 688028 45099 688098
rect 45099 688028 45118 688098
rect 45048 687738 45065 687808
rect 45065 687738 45099 687808
rect 45099 687738 45118 687808
rect 44888 687468 44907 687538
rect 44907 687468 44941 687538
rect 44941 687468 44958 687538
rect 44888 687178 44907 687248
rect 44907 687178 44941 687248
rect 44941 687178 44958 687248
rect 45368 688028 45381 688098
rect 45381 688028 45415 688098
rect 45415 688028 45438 688098
rect 45368 687738 45381 687808
rect 45381 687738 45415 687808
rect 45415 687738 45438 687808
rect 45208 687468 45223 687538
rect 45223 687468 45257 687538
rect 45257 687468 45278 687538
rect 45208 687178 45223 687248
rect 45223 687178 45257 687248
rect 45257 687178 45278 687248
rect 45678 688028 45697 688098
rect 45697 688028 45731 688098
rect 45731 688028 45748 688098
rect 45678 687738 45697 687808
rect 45697 687738 45731 687808
rect 45731 687738 45748 687808
rect 45528 687468 45539 687538
rect 45539 687468 45573 687538
rect 45573 687468 45598 687538
rect 45528 687178 45539 687248
rect 45539 687178 45573 687248
rect 45573 687178 45598 687248
rect 45998 688028 46013 688098
rect 46013 688028 46047 688098
rect 46047 688028 46068 688098
rect 45998 687738 46013 687808
rect 46013 687738 46047 687808
rect 46047 687738 46068 687808
rect 45838 687468 45855 687538
rect 45855 687468 45889 687538
rect 45889 687468 45908 687538
rect 45838 687178 45855 687248
rect 45855 687178 45889 687248
rect 45889 687178 45908 687248
rect 45348 686999 45608 687008
rect 45348 686965 45608 686999
rect 45348 686792 45608 686965
rect 45348 686758 45608 686792
rect 45348 686748 45608 686758
rect 43108 686618 43218 686728
rect 43358 686618 43468 686728
rect 47508 686618 47618 686728
rect 47758 686618 47868 686728
rect 43888 686508 43908 686578
rect 43908 686508 43942 686578
rect 43942 686508 43958 686578
rect 43888 686328 43908 686398
rect 43908 686328 43942 686398
rect 43942 686328 43958 686398
rect 44408 686508 44424 686578
rect 44424 686508 44458 686578
rect 44458 686508 44478 686578
rect 44408 686328 44424 686398
rect 44424 686328 44458 686398
rect 44458 686328 44478 686398
rect 44148 685838 44166 685908
rect 44166 685838 44200 685908
rect 44200 685838 44218 685908
rect 44148 685658 44166 685728
rect 44166 685658 44200 685728
rect 44200 685658 44218 685728
rect 44928 686508 44940 686578
rect 44940 686508 44974 686578
rect 44974 686508 44998 686578
rect 44928 686328 44940 686398
rect 44940 686328 44974 686398
rect 44974 686328 44998 686398
rect 44668 685838 44682 685908
rect 44682 685838 44716 685908
rect 44716 685838 44738 685908
rect 44668 685658 44682 685728
rect 44682 685658 44716 685728
rect 44716 685658 44738 685728
rect 45438 686508 45456 686578
rect 45456 686508 45490 686578
rect 45490 686508 45508 686578
rect 45438 686328 45456 686398
rect 45456 686328 45490 686398
rect 45490 686328 45508 686398
rect 45178 685838 45198 685908
rect 45198 685838 45232 685908
rect 45232 685838 45248 685908
rect 45178 685658 45198 685728
rect 45198 685658 45232 685728
rect 45232 685658 45248 685728
rect 45958 686508 45972 686578
rect 45972 686508 46006 686578
rect 46006 686508 46028 686578
rect 45958 686328 45972 686398
rect 45972 686328 46006 686398
rect 46006 686328 46028 686398
rect 45698 685838 45714 685908
rect 45714 685838 45748 685908
rect 45748 685838 45768 685908
rect 45698 685658 45714 685728
rect 45714 685658 45748 685728
rect 45748 685658 45768 685728
rect 46468 686508 46488 686578
rect 46488 686508 46522 686578
rect 46522 686508 46538 686578
rect 46468 686328 46488 686398
rect 46488 686328 46522 686398
rect 46522 686328 46538 686398
rect 46218 685838 46230 685908
rect 46230 685838 46264 685908
rect 46264 685838 46288 685908
rect 46218 685658 46230 685728
rect 46230 685658 46264 685728
rect 46264 685658 46288 685728
rect 46988 686508 47004 686578
rect 47004 686508 47038 686578
rect 47038 686508 47058 686578
rect 46988 686328 47004 686398
rect 47004 686328 47038 686398
rect 47038 686328 47058 686398
rect 46728 685838 46746 685908
rect 46746 685838 46780 685908
rect 46780 685838 46798 685908
rect 46728 685658 46746 685728
rect 46746 685658 46780 685728
rect 46780 685658 46798 685728
rect 43108 685508 43218 685618
rect 43358 685508 43468 685618
rect 47508 685508 47618 685618
rect 47758 685508 47868 685618
rect 45348 685478 45598 685488
rect 45348 685444 45598 685478
rect 45348 685272 45598 685444
rect 45348 685238 45598 685272
rect 43108 685098 43218 685208
rect 43358 685098 43468 685208
rect 47508 685098 47618 685208
rect 47758 685098 47868 685208
rect 43638 684988 43652 685058
rect 43652 684988 43686 685058
rect 43686 684988 43708 685058
rect 43638 684808 43652 684878
rect 43652 684808 43686 684878
rect 43686 684808 43708 684878
rect 44148 684988 44168 685058
rect 44168 684988 44202 685058
rect 44202 684988 44218 685058
rect 44148 684808 44168 684878
rect 44168 684808 44202 684878
rect 44202 684808 44218 684878
rect 43898 684318 43910 684388
rect 43910 684318 43944 684388
rect 43944 684318 43968 684388
rect 43898 684138 43910 684208
rect 43910 684138 43944 684208
rect 43944 684138 43968 684208
rect 44668 684988 44684 685058
rect 44684 684988 44718 685058
rect 44718 684988 44738 685058
rect 44668 684808 44684 684878
rect 44684 684808 44718 684878
rect 44718 684808 44738 684878
rect 44408 684318 44426 684388
rect 44426 684318 44460 684388
rect 44460 684318 44478 684388
rect 44408 684138 44426 684208
rect 44426 684138 44460 684208
rect 44460 684138 44478 684208
rect 45188 684988 45200 685058
rect 45200 684988 45234 685058
rect 45234 684988 45258 685058
rect 45188 684808 45200 684878
rect 45200 684808 45234 684878
rect 45234 684808 45258 684878
rect 44928 684318 44942 684388
rect 44942 684318 44976 684388
rect 44976 684318 44998 684388
rect 44928 684138 44942 684208
rect 44942 684138 44976 684208
rect 44976 684138 44998 684208
rect 45698 684988 45716 685058
rect 45716 684988 45750 685058
rect 45750 684988 45768 685058
rect 45698 684808 45716 684878
rect 45716 684808 45750 684878
rect 45750 684808 45768 684878
rect 45438 684318 45458 684388
rect 45458 684318 45492 684388
rect 45492 684318 45508 684388
rect 45438 684138 45458 684208
rect 45458 684138 45492 684208
rect 45492 684138 45508 684208
rect 46218 684988 46232 685058
rect 46232 684988 46266 685058
rect 46266 684988 46288 685058
rect 46218 684808 46232 684878
rect 46232 684808 46266 684878
rect 46266 684808 46288 684878
rect 45958 684318 45974 684388
rect 45974 684318 46008 684388
rect 46008 684318 46028 684388
rect 45958 684138 45974 684208
rect 45974 684138 46008 684208
rect 46008 684138 46028 684208
rect 46728 684988 46748 685058
rect 46748 684988 46782 685058
rect 46782 684988 46798 685058
rect 46728 684808 46748 684878
rect 46748 684808 46782 684878
rect 46782 684808 46798 684878
rect 46478 684318 46490 684388
rect 46490 684318 46524 684388
rect 46524 684318 46548 684388
rect 46478 684138 46490 684208
rect 46490 684138 46524 684208
rect 46524 684138 46548 684208
rect 47248 684988 47264 685058
rect 47264 684988 47298 685058
rect 47298 684988 47318 685058
rect 47248 684808 47264 684878
rect 47264 684808 47298 684878
rect 47298 684808 47318 684878
rect 46988 684318 47006 684388
rect 47006 684318 47040 684388
rect 47040 684318 47058 684388
rect 46988 684138 47006 684208
rect 47006 684138 47040 684208
rect 47040 684138 47058 684208
rect 43108 683988 43218 684098
rect 43358 683988 43468 684098
rect 47508 683988 47618 684098
rect 47758 683988 47868 684098
rect 45348 683924 45598 683958
rect 45348 683708 45598 683924
rect 42308 682918 42468 683078
rect 43308 682918 43468 683078
rect 44788 682918 44948 683078
rect 46008 682918 46168 683078
rect 47468 682918 47628 683078
rect 48528 682918 48688 683078
rect 43698 682688 43768 682758
rect 43938 682688 44008 682758
rect 46898 682688 46968 682758
rect 47118 682688 47188 682758
rect 42308 682338 42468 682498
rect 43308 682338 43468 682498
rect 44788 682338 44948 682498
rect 46008 682338 46168 682498
rect 47468 682338 47628 682498
rect 48528 682338 48688 682498
rect 43698 682098 43768 682168
rect 43938 682098 44008 682168
rect 46898 682098 46968 682168
rect 47118 682098 47188 682168
rect 44908 681988 44978 682008
rect 45018 681988 45088 682008
rect 45848 681988 45918 682008
rect 45958 681988 46028 682008
rect 44908 681938 44978 681988
rect 45018 681938 45088 681988
rect 45848 681938 45918 681988
rect 45958 681938 46028 681988
rect 44908 681428 44978 681448
rect 44908 681378 44932 681428
rect 44932 681378 44966 681428
rect 44966 681378 44978 681428
rect 45018 681428 45088 681448
rect 45848 681428 45918 681438
rect 45018 681378 45040 681428
rect 45040 681378 45074 681428
rect 45074 681378 45088 681428
rect 45848 681368 45868 681428
rect 45868 681368 45902 681428
rect 45902 681368 45918 681428
rect 45958 681428 46028 681438
rect 45958 681368 45976 681428
rect 45976 681368 46010 681428
rect 46010 681368 46028 681428
rect 44598 680968 44818 681118
rect 46088 680968 46308 681118
rect 43698 680858 43768 680928
rect 43938 680858 44008 680928
rect 43698 680768 43768 680838
rect 43938 680768 44008 680838
rect 46908 680838 46978 680908
rect 47118 680838 47188 680908
rect 46908 680748 46978 680818
rect 47118 680748 47188 680818
rect 44908 680673 44978 680688
rect 45018 680673 45088 680688
rect 45848 680673 45918 680688
rect 45958 680673 46028 680688
rect 44908 680618 44978 680673
rect 45018 680618 45088 680673
rect 45848 680618 45918 680673
rect 45958 680618 46028 680673
rect 42368 680438 42548 680568
rect 43368 680438 43548 680568
rect 44438 680428 44618 680558
rect 45158 680438 45338 680568
rect 45598 680438 45778 680568
rect 46368 680438 46548 680568
rect 47348 680428 47528 680558
rect 48488 680428 48668 680558
rect 43698 680340 43768 680388
rect 43938 680340 44008 680388
rect 46898 680340 46968 680388
rect 47118 680340 47188 680388
rect 43698 680318 43768 680340
rect 43938 680318 44008 680340
rect 46898 680318 46968 680340
rect 47118 680318 47188 680340
rect 44908 680168 44978 680238
rect 45018 680168 45088 680238
rect 45848 680168 45918 680238
rect 45958 680168 46028 680238
rect 42218 678538 42338 678658
rect 48588 678538 48708 678658
rect 42218 675538 42338 675658
rect 48588 675538 48708 675658
rect 42218 672538 42338 672658
rect 48588 672538 48708 672658
rect 42218 669538 42338 669658
rect 48588 669538 48708 669658
rect 42218 666538 42338 666658
rect 48588 666538 48708 666658
rect 42608 664962 42641 665338
rect 42641 664962 43755 665338
rect 43755 664962 43778 665338
rect 42608 664928 43778 664962
rect 44128 664962 44151 665328
rect 44151 664962 45265 665328
rect 45265 664962 45298 665328
rect 44128 664918 45298 664962
rect 45648 664956 45661 665328
rect 45661 664956 46775 665328
rect 46775 664956 46818 665328
rect 45648 664918 46818 664956
rect 47158 664956 47181 665328
rect 47181 664956 48295 665328
rect 48295 664956 48328 665328
rect 47158 664918 48328 664956
<< metal2 >>
rect 44798 694878 45068 694888
rect 44798 694598 45068 694608
rect 45848 694878 46118 694888
rect 45848 694598 46118 694608
rect 42278 694398 42348 694408
rect 42278 694318 42348 694328
rect 42588 694398 42658 694408
rect 42588 694318 42658 694328
rect 42908 694398 42978 694408
rect 42908 694318 42978 694328
rect 43228 694398 43298 694408
rect 43228 694318 43298 694328
rect 43538 694398 43608 694408
rect 43538 694318 43608 694328
rect 43858 694398 43928 694408
rect 43858 694318 43928 694328
rect 44168 694398 44238 694408
rect 44168 694318 44238 694328
rect 44488 694398 44558 694408
rect 44488 694318 44558 694328
rect 44808 694398 44878 694408
rect 44808 694318 44878 694328
rect 45118 694398 45188 694408
rect 45118 694318 45188 694328
rect 45438 694398 45508 694408
rect 45438 694318 45508 694328
rect 45748 694398 45818 694408
rect 45748 694318 45818 694328
rect 46068 694398 46138 694408
rect 46068 694318 46138 694328
rect 46388 694398 46458 694408
rect 46388 694318 46458 694328
rect 46698 694398 46768 694408
rect 46698 694318 46768 694328
rect 47018 694398 47088 694408
rect 47018 694318 47088 694328
rect 47338 694398 47408 694408
rect 47338 694318 47408 694328
rect 47648 694398 47718 694408
rect 47648 694318 47718 694328
rect 47968 694398 48038 694408
rect 47968 694318 48038 694328
rect 48278 694398 48348 694408
rect 48278 694318 48348 694328
rect 48598 694398 48668 694408
rect 48598 694318 48668 694328
rect 37608 694158 37828 694178
rect 37608 694088 37738 694158
rect 37808 694088 37828 694158
rect 37608 694048 37828 694088
rect 42278 694158 42348 694168
rect 42278 694078 42348 694088
rect 42588 694158 42658 694168
rect 42588 694078 42658 694088
rect 42908 694158 42978 694168
rect 42908 694078 42978 694088
rect 43228 694158 43298 694168
rect 43228 694078 43298 694088
rect 43538 694158 43608 694168
rect 43538 694078 43608 694088
rect 43858 694158 43928 694168
rect 43858 694078 43928 694088
rect 44168 694158 44238 694168
rect 44168 694078 44238 694088
rect 44488 694158 44558 694168
rect 44488 694078 44558 694088
rect 44808 694158 44878 694168
rect 44808 694078 44878 694088
rect 45118 694158 45188 694168
rect 45118 694078 45188 694088
rect 45438 694158 45508 694168
rect 45438 694078 45508 694088
rect 45748 694158 45818 694168
rect 45748 694078 45818 694088
rect 46068 694158 46138 694168
rect 46068 694078 46138 694088
rect 46388 694158 46458 694168
rect 46388 694078 46458 694088
rect 46698 694158 46768 694168
rect 46698 694078 46768 694088
rect 47018 694158 47088 694168
rect 47018 694078 47088 694088
rect 47338 694158 47408 694168
rect 47338 694078 47408 694088
rect 47648 694158 47718 694168
rect 47648 694078 47718 694088
rect 47968 694158 48038 694168
rect 47968 694078 48038 694088
rect 48278 694158 48348 694168
rect 48278 694078 48348 694088
rect 48598 694158 48668 694168
rect 48598 694078 48668 694088
rect 53108 694158 53328 694178
rect 53108 694088 53128 694158
rect 53198 694088 53328 694158
rect 37608 693978 37628 694048
rect 37698 693978 37828 694048
rect 37608 693958 37828 693978
rect 53108 694048 53328 694088
rect 53108 693978 53238 694048
rect 53308 693978 53328 694048
rect 53108 693958 53328 693978
rect 42398 693788 42528 693798
rect 42398 693718 42428 693788
rect 42498 693718 42528 693788
rect 42398 693548 42528 693718
rect 42748 693788 42818 693798
rect 42748 693708 42818 693718
rect 43068 693788 43138 693798
rect 43068 693708 43138 693718
rect 43378 693788 43448 693798
rect 43378 693708 43448 693718
rect 43698 693788 43768 693798
rect 43698 693708 43768 693718
rect 44018 693788 44088 693798
rect 44018 693708 44088 693718
rect 44328 693788 44398 693798
rect 44328 693708 44398 693718
rect 44648 693788 44718 693798
rect 44648 693708 44718 693718
rect 44958 693788 45028 693798
rect 44958 693708 45028 693718
rect 45278 693788 45348 693798
rect 45278 693708 45348 693718
rect 45598 693788 45668 693798
rect 45598 693708 45668 693718
rect 45908 693788 45978 693798
rect 45908 693708 45978 693718
rect 46228 693788 46298 693798
rect 46228 693708 46298 693718
rect 46548 693788 46618 693798
rect 46548 693708 46618 693718
rect 46858 693788 46928 693798
rect 46858 693708 46928 693718
rect 47178 693788 47248 693798
rect 47178 693708 47248 693718
rect 47488 693788 47558 693798
rect 47488 693708 47558 693718
rect 47808 693788 47878 693798
rect 47808 693708 47878 693718
rect 48128 693788 48198 693798
rect 48128 693708 48198 693718
rect 48408 693788 48538 693798
rect 48408 693718 48438 693788
rect 48508 693718 48538 693788
rect 42398 693478 42428 693548
rect 42498 693478 42528 693548
rect 42398 693178 42528 693478
rect 42748 693548 42818 693558
rect 42748 693468 42818 693478
rect 43068 693548 43138 693558
rect 43068 693468 43138 693478
rect 43378 693548 43448 693558
rect 43378 693468 43448 693478
rect 43698 693548 43768 693558
rect 43698 693468 43768 693478
rect 44018 693548 44088 693558
rect 44018 693468 44088 693478
rect 44328 693548 44398 693558
rect 44328 693468 44398 693478
rect 44648 693548 44718 693558
rect 44648 693468 44718 693478
rect 44958 693548 45028 693558
rect 44958 693468 45028 693478
rect 45278 693548 45348 693558
rect 45278 693468 45348 693478
rect 45598 693548 45668 693558
rect 45598 693468 45668 693478
rect 45908 693548 45978 693558
rect 45908 693468 45978 693478
rect 46228 693548 46298 693558
rect 46228 693468 46298 693478
rect 46548 693548 46618 693558
rect 46548 693468 46618 693478
rect 46858 693548 46928 693558
rect 46858 693468 46928 693478
rect 47178 693548 47248 693558
rect 47178 693468 47248 693478
rect 47488 693548 47558 693558
rect 47488 693468 47558 693478
rect 47808 693548 47878 693558
rect 47808 693468 47878 693478
rect 48128 693548 48198 693558
rect 48128 693468 48198 693478
rect 42398 693108 42428 693178
rect 42498 693108 42528 693178
rect 39578 692698 39758 692708
rect 39578 692588 39758 692598
rect 39998 692698 40178 692708
rect 39998 692588 40178 692598
rect 42398 686568 42528 693108
rect 43368 693378 43528 693398
rect 43368 693298 43408 693378
rect 43488 693298 43528 693378
rect 43368 692078 43528 693298
rect 47428 693378 47588 693398
rect 47428 693298 47468 693378
rect 47548 693298 47588 693378
rect 44798 693238 45068 693248
rect 44798 692958 45068 692968
rect 45848 693238 46118 693248
rect 45848 692958 46118 692968
rect 43938 692728 44008 692738
rect 43938 692648 44008 692658
rect 44248 692728 44318 692738
rect 44248 692648 44318 692658
rect 44568 692728 44638 692738
rect 44568 692648 44638 692658
rect 44878 692728 44948 692738
rect 44878 692648 44948 692658
rect 45198 692728 45268 692738
rect 45198 692648 45268 692658
rect 45518 692728 45588 692738
rect 45518 692648 45588 692658
rect 45828 692728 45898 692738
rect 45828 692648 45898 692658
rect 46148 692728 46218 692738
rect 46148 692648 46218 692658
rect 46468 692728 46538 692738
rect 46468 692648 46538 692658
rect 46778 692728 46848 692738
rect 46778 692648 46848 692658
rect 47098 692728 47168 692738
rect 47098 692648 47168 692658
rect 43938 692518 44008 692528
rect 43938 692438 44008 692448
rect 44248 692518 44318 692528
rect 44248 692438 44318 692448
rect 44568 692518 44638 692528
rect 44568 692438 44638 692448
rect 44878 692518 44948 692528
rect 44878 692438 44948 692448
rect 45198 692518 45268 692528
rect 45198 692438 45268 692448
rect 45518 692518 45588 692528
rect 45518 692438 45588 692448
rect 45828 692518 45898 692528
rect 45828 692438 45898 692448
rect 46148 692518 46218 692528
rect 46148 692438 46218 692448
rect 46468 692518 46538 692528
rect 46468 692438 46538 692448
rect 46778 692518 46848 692528
rect 46778 692438 46848 692448
rect 47098 692518 47168 692528
rect 47098 692438 47168 692448
rect 43368 691998 43408 692078
rect 43488 691998 43528 692078
rect 43778 692088 43848 692098
rect 43778 692008 43848 692018
rect 44088 692088 44158 692098
rect 44088 692008 44158 692018
rect 44408 692088 44478 692098
rect 44408 692008 44478 692018
rect 44728 692088 44798 692098
rect 44728 692008 44798 692018
rect 45038 692088 45108 692098
rect 45038 692008 45108 692018
rect 45358 692088 45428 692098
rect 45358 692008 45428 692018
rect 45668 692088 45738 692098
rect 45668 692008 45738 692018
rect 45988 692088 46058 692098
rect 45988 692008 46058 692018
rect 46308 692088 46378 692098
rect 46308 692008 46378 692018
rect 46618 692088 46688 692098
rect 46618 692008 46688 692018
rect 46938 692088 47008 692098
rect 46938 692008 47008 692018
rect 47428 692078 47588 693298
rect 43368 691898 43528 691998
rect 43368 691818 43408 691898
rect 43488 691818 43528 691898
rect 47428 691998 47468 692078
rect 47548 691998 47588 692078
rect 47428 691898 47588 691998
rect 43368 689608 43528 691818
rect 43778 691878 43848 691888
rect 43778 691798 43848 691808
rect 44088 691878 44158 691888
rect 44088 691798 44158 691808
rect 44408 691878 44478 691888
rect 44408 691798 44478 691808
rect 44728 691878 44798 691888
rect 44728 691798 44798 691808
rect 45038 691878 45108 691888
rect 45038 691798 45108 691808
rect 45358 691878 45428 691888
rect 45358 691798 45428 691808
rect 45668 691878 45738 691888
rect 45668 691798 45738 691808
rect 45988 691878 46058 691888
rect 45988 691798 46058 691808
rect 46308 691878 46378 691888
rect 46308 691798 46378 691808
rect 46618 691878 46688 691888
rect 46618 691798 46688 691808
rect 46938 691878 47008 691888
rect 46938 691798 47008 691808
rect 47428 691818 47468 691898
rect 47548 691818 47588 691898
rect 44588 691628 44848 691638
rect 44588 691358 44848 691368
rect 46088 691628 46348 691638
rect 46088 691358 46348 691368
rect 43938 691178 44008 691188
rect 43938 691098 44008 691108
rect 44248 691178 44318 691188
rect 44248 691098 44318 691108
rect 44568 691178 44638 691188
rect 44568 691098 44638 691108
rect 44888 691178 44958 691188
rect 44888 691098 44958 691108
rect 45198 691178 45268 691188
rect 45198 691098 45268 691108
rect 45518 691178 45588 691188
rect 45518 691098 45588 691108
rect 45828 691178 45898 691188
rect 45828 691098 45898 691108
rect 46148 691178 46218 691188
rect 46148 691098 46218 691108
rect 46468 691178 46538 691188
rect 46468 691098 46538 691108
rect 46778 691178 46848 691188
rect 46778 691098 46848 691108
rect 47098 691178 47168 691188
rect 47098 691098 47168 691108
rect 43938 690968 44008 690978
rect 43938 690888 44008 690898
rect 44248 690968 44318 690978
rect 44248 690888 44318 690898
rect 44568 690968 44638 690978
rect 44568 690888 44638 690898
rect 44888 690968 44958 690978
rect 44888 690888 44958 690898
rect 45198 690968 45268 690978
rect 45198 690888 45268 690898
rect 45518 690968 45588 690978
rect 45518 690888 45588 690898
rect 45828 690968 45898 690978
rect 45828 690888 45898 690898
rect 46148 690968 46218 690978
rect 46148 690888 46218 690898
rect 46468 690968 46538 690978
rect 46468 690888 46538 690898
rect 46778 690968 46848 690978
rect 46778 690888 46848 690898
rect 47098 690968 47168 690978
rect 47098 690888 47168 690898
rect 43778 690548 43848 690558
rect 43778 690468 43848 690478
rect 44068 690548 44198 690558
rect 44068 690478 44098 690548
rect 44168 690478 44198 690548
rect 43778 690338 43848 690348
rect 43778 690258 43848 690268
rect 44068 690338 44198 690478
rect 44408 690548 44478 690558
rect 44408 690468 44478 690478
rect 44728 690548 44798 690558
rect 44728 690468 44798 690478
rect 45038 690548 45108 690558
rect 45038 690468 45108 690478
rect 45358 690548 45428 690558
rect 45358 690468 45428 690478
rect 45678 690548 45748 690558
rect 45678 690468 45748 690478
rect 45988 690548 46058 690558
rect 45988 690468 46058 690478
rect 46308 690548 46378 690558
rect 46308 690468 46378 690478
rect 46588 690548 46718 690558
rect 46588 690478 46618 690548
rect 46688 690478 46718 690548
rect 44068 690268 44098 690338
rect 44168 690268 44198 690338
rect 43368 689488 43388 689608
rect 43508 689488 43528 689608
rect 43368 689388 43528 689488
rect 43368 689268 43388 689388
rect 43508 689268 43528 689388
rect 43368 689248 43528 689268
rect 43608 689048 43768 689068
rect 43608 688928 43628 689048
rect 43748 688928 43768 689048
rect 43608 688828 43768 688928
rect 43608 688708 43628 688828
rect 43748 688708 43768 688828
rect 43608 688088 43768 688708
rect 43608 687968 43628 688088
rect 43748 687968 43768 688088
rect 43300 687920 43480 687960
rect 43300 687760 43340 687920
rect 43460 687760 43480 687920
rect 43300 687720 43480 687760
rect 43300 687560 43340 687720
rect 43460 687560 43480 687720
rect 43300 687520 43480 687560
rect 43608 687868 43768 687968
rect 43608 687748 43628 687868
rect 43748 687748 43768 687868
rect 42398 686498 42428 686568
rect 42498 686498 42528 686568
rect 42398 686408 42528 686498
rect 42398 686338 42428 686408
rect 42498 686338 42528 686408
rect 42398 686318 42528 686338
rect 43088 686728 43488 686848
rect 43088 686618 43108 686728
rect 43218 686618 43358 686728
rect 43468 686618 43488 686728
rect 43088 685618 43488 686618
rect 43088 685508 43108 685618
rect 43218 685508 43358 685618
rect 43468 685508 43488 685618
rect 43088 685208 43488 685508
rect 43088 685098 43108 685208
rect 43218 685098 43358 685208
rect 43468 685098 43488 685208
rect 43088 684098 43488 685098
rect 43608 685058 43768 687748
rect 44068 687518 44198 690268
rect 44408 690338 44478 690348
rect 44408 690258 44478 690268
rect 44728 690338 44798 690348
rect 44728 690258 44798 690268
rect 45038 690338 45108 690348
rect 45038 690258 45108 690268
rect 45358 690338 45428 690348
rect 45358 690258 45428 690268
rect 45678 690338 45748 690348
rect 45678 690258 45748 690268
rect 45988 690338 46058 690348
rect 45988 690258 46058 690268
rect 46308 690338 46378 690348
rect 46308 690258 46378 690268
rect 46588 690338 46718 690478
rect 46938 690548 47008 690558
rect 46938 690468 47008 690478
rect 46588 690268 46618 690338
rect 46688 690268 46718 690338
rect 45048 689618 45118 689628
rect 45048 689538 45118 689548
rect 45368 689618 45438 689628
rect 45368 689538 45438 689548
rect 45678 689618 45748 689628
rect 45678 689538 45748 689548
rect 45998 689618 46068 689628
rect 45998 689538 46068 689548
rect 45048 689328 45118 689338
rect 45048 689248 45118 689258
rect 45368 689328 45438 689338
rect 45368 689248 45438 689258
rect 45678 689328 45748 689338
rect 45678 689248 45748 689258
rect 45998 689328 46068 689338
rect 45998 689248 46068 689258
rect 44888 689058 44958 689068
rect 44888 688978 44958 688988
rect 45208 689058 45278 689068
rect 45208 688978 45278 688988
rect 45528 689058 45598 689068
rect 45528 688978 45598 688988
rect 45838 689058 45908 689068
rect 45838 688978 45908 688988
rect 44888 688768 44958 688778
rect 44888 688688 44958 688698
rect 45208 688768 45278 688778
rect 45208 688688 45278 688698
rect 45528 688768 45598 688778
rect 45528 688688 45598 688698
rect 45838 688768 45908 688778
rect 45838 688688 45908 688698
rect 45348 688528 45608 688538
rect 45348 688258 45608 688268
rect 45048 688098 45118 688108
rect 45048 688018 45118 688028
rect 45368 688098 45438 688108
rect 45368 688018 45438 688028
rect 45678 688098 45748 688108
rect 45678 688018 45748 688028
rect 45998 688098 46068 688108
rect 45998 688018 46068 688028
rect 45048 687808 45118 687818
rect 45048 687728 45118 687738
rect 45368 687808 45438 687818
rect 45368 687728 45438 687738
rect 45678 687808 45748 687818
rect 45678 687728 45748 687738
rect 45998 687808 46068 687818
rect 45998 687728 46068 687738
rect 44068 687448 44098 687518
rect 44168 687448 44198 687518
rect 44888 687538 44958 687548
rect 44888 687458 44958 687468
rect 45208 687538 45278 687548
rect 45208 687458 45278 687468
rect 45528 687538 45598 687548
rect 45528 687458 45598 687468
rect 45838 687538 45908 687548
rect 45838 687458 45908 687468
rect 46588 687518 46718 690268
rect 46938 690338 47008 690348
rect 46938 690258 47008 690268
rect 47428 689608 47588 691818
rect 47428 689488 47448 689608
rect 47568 689488 47588 689608
rect 47428 689388 47588 689488
rect 48408 693178 48538 693718
rect 48408 693108 48438 693178
rect 48508 693108 48538 693178
rect 47428 689268 47448 689388
rect 47568 689268 47588 689388
rect 47428 689248 47588 689268
rect 47940 689380 48120 689400
rect 47940 689260 47960 689380
rect 48100 689260 48120 689380
rect 47940 689220 48120 689260
rect 47940 689100 47960 689220
rect 48100 689100 48120 689220
rect 44068 687268 44198 687448
rect 44068 687198 44098 687268
rect 44168 687198 44198 687268
rect 46588 687448 46618 687518
rect 46688 687448 46718 687518
rect 46588 687268 46718 687448
rect 44068 687168 44198 687198
rect 44888 687248 44958 687258
rect 44888 687168 44958 687178
rect 45208 687248 45278 687258
rect 45208 687168 45278 687178
rect 45528 687248 45598 687258
rect 45528 687168 45598 687178
rect 45838 687248 45908 687258
rect 45838 687168 45908 687178
rect 46588 687198 46618 687268
rect 46688 687198 46718 687268
rect 46588 687168 46718 687198
rect 47188 689048 47348 689068
rect 47188 688928 47208 689048
rect 47328 688928 47348 689048
rect 47188 688828 47348 688928
rect 47940 689040 48120 689100
rect 47940 688920 47960 689040
rect 48100 688920 48120 689040
rect 47940 688900 48120 688920
rect 47188 688708 47208 688828
rect 47328 688708 47348 688828
rect 47188 688088 47348 688708
rect 47188 687968 47208 688088
rect 47328 687968 47348 688088
rect 47188 687868 47348 687968
rect 47188 687748 47208 687868
rect 47328 687748 47348 687868
rect 45348 687008 45608 687018
rect 45348 686738 45608 686748
rect 43888 686578 43958 686588
rect 43888 686498 43958 686508
rect 44408 686578 44478 686588
rect 44408 686498 44478 686508
rect 44928 686578 44998 686588
rect 44928 686498 44998 686508
rect 45438 686578 45508 686588
rect 45438 686498 45508 686508
rect 45958 686578 46028 686588
rect 45958 686498 46028 686508
rect 46468 686578 46538 686588
rect 46468 686498 46538 686508
rect 46988 686578 47058 686588
rect 46988 686498 47058 686508
rect 43888 686398 43958 686408
rect 43888 686318 43958 686328
rect 44408 686398 44478 686408
rect 44408 686318 44478 686328
rect 44928 686398 44998 686408
rect 44928 686318 44998 686328
rect 45438 686398 45508 686408
rect 45438 686318 45508 686328
rect 45958 686398 46028 686408
rect 45958 686318 46028 686328
rect 46468 686398 46538 686408
rect 46468 686318 46538 686328
rect 46988 686398 47058 686408
rect 46988 686318 47058 686328
rect 44148 685908 44218 685918
rect 44148 685828 44218 685838
rect 44668 685908 44738 685918
rect 44668 685828 44738 685838
rect 45178 685908 45248 685918
rect 45178 685828 45248 685838
rect 45698 685908 45768 685918
rect 45698 685828 45768 685838
rect 46218 685908 46288 685918
rect 46218 685828 46288 685838
rect 46728 685908 46798 685918
rect 46728 685828 46798 685838
rect 44148 685728 44218 685738
rect 44148 685648 44218 685658
rect 44668 685728 44738 685738
rect 44668 685648 44738 685658
rect 45178 685728 45248 685738
rect 45178 685648 45248 685658
rect 45698 685728 45768 685738
rect 45698 685648 45768 685658
rect 46218 685728 46288 685738
rect 46218 685648 46288 685658
rect 46728 685728 46798 685738
rect 46728 685648 46798 685658
rect 45348 685488 45598 685498
rect 45348 685228 45598 685238
rect 43608 684988 43638 685058
rect 43708 684988 43768 685058
rect 43608 684878 43768 684988
rect 44148 685058 44218 685068
rect 44148 684978 44218 684988
rect 44668 685058 44738 685068
rect 44668 684978 44738 684988
rect 45188 685058 45258 685068
rect 45188 684978 45258 684988
rect 45698 685058 45768 685068
rect 45698 684978 45768 684988
rect 46218 685058 46288 685068
rect 46218 684978 46288 684988
rect 46728 685058 46798 685068
rect 46728 684978 46798 684988
rect 47188 685058 47348 687748
rect 47188 684988 47248 685058
rect 47318 684988 47348 685058
rect 43608 684808 43638 684878
rect 43708 684808 43768 684878
rect 43608 684798 43768 684808
rect 44148 684878 44218 684888
rect 44148 684798 44218 684808
rect 44668 684878 44738 684888
rect 44668 684798 44738 684808
rect 45188 684878 45258 684888
rect 45188 684798 45258 684808
rect 45698 684878 45768 684888
rect 45698 684798 45768 684808
rect 46218 684878 46288 684888
rect 46218 684798 46288 684808
rect 46728 684878 46798 684888
rect 46728 684798 46798 684808
rect 47188 684878 47348 684988
rect 47188 684808 47248 684878
rect 47318 684808 47348 684878
rect 47188 684798 47348 684808
rect 47488 686728 47888 686848
rect 47488 686618 47508 686728
rect 47618 686618 47758 686728
rect 47868 686618 47888 686728
rect 47488 685618 47888 686618
rect 48408 686568 48538 693108
rect 50828 692698 51008 692708
rect 50828 692588 51008 692598
rect 51248 692698 51428 692708
rect 51248 692588 51428 692598
rect 48408 686498 48438 686568
rect 48508 686498 48538 686568
rect 48408 686408 48538 686498
rect 48408 686338 48438 686408
rect 48508 686338 48538 686408
rect 48408 686318 48538 686338
rect 47488 685508 47508 685618
rect 47618 685508 47758 685618
rect 47868 685508 47888 685618
rect 47488 685208 47888 685508
rect 47488 685098 47508 685208
rect 47618 685098 47758 685208
rect 47868 685098 47888 685208
rect 43898 684388 43968 684398
rect 43898 684308 43968 684318
rect 44408 684388 44478 684398
rect 44408 684308 44478 684318
rect 44928 684388 44998 684398
rect 44928 684308 44998 684318
rect 45438 684388 45508 684398
rect 45438 684308 45508 684318
rect 45958 684388 46028 684398
rect 45958 684308 46028 684318
rect 46478 684388 46548 684398
rect 46478 684308 46548 684318
rect 46988 684388 47058 684398
rect 46988 684308 47058 684318
rect 43898 684208 43968 684218
rect 43898 684128 43968 684138
rect 44408 684208 44478 684218
rect 44408 684128 44478 684138
rect 44928 684208 44998 684218
rect 44928 684128 44998 684138
rect 45438 684208 45508 684218
rect 45438 684128 45508 684138
rect 45958 684208 46028 684218
rect 45958 684128 46028 684138
rect 46478 684208 46548 684218
rect 46478 684128 46548 684138
rect 46988 684208 47058 684218
rect 46988 684128 47058 684138
rect 43088 683988 43108 684098
rect 43218 683988 43358 684098
rect 43468 683988 43488 684098
rect 43088 683808 43488 683988
rect 47488 684098 47888 685098
rect 47488 683988 47508 684098
rect 47618 683988 47758 684098
rect 47868 683988 47888 684098
rect 45348 683958 45598 683968
rect 43088 683608 45138 683808
rect 47488 683808 47888 683988
rect 45348 683698 45598 683708
rect 42308 683078 42468 683088
rect 42308 682908 42468 682918
rect 43308 683078 43468 683088
rect 43308 682908 43468 682918
rect 44788 683078 44948 683088
rect 44788 682908 44948 682918
rect 43678 682758 44028 682768
rect 43678 682688 43698 682758
rect 43768 682688 43938 682758
rect 44008 682688 44028 682758
rect 42308 682498 42468 682508
rect 42308 682328 42468 682338
rect 43308 682498 43468 682508
rect 43308 682328 43468 682338
rect 43678 682168 44028 682688
rect 44788 682498 44948 682508
rect 44788 682328 44948 682338
rect 44988 682268 45138 683608
rect 45798 683608 47888 683808
rect 45798 682268 45948 683608
rect 46008 683078 46168 683088
rect 46008 682908 46168 682918
rect 47468 683078 47628 683088
rect 47468 682908 47628 682918
rect 48528 683078 48688 683088
rect 48528 682908 48688 682918
rect 46878 682688 46898 682758
rect 46968 682688 47118 682758
rect 47188 682688 47208 682758
rect 46008 682498 46168 682508
rect 46008 682328 46168 682338
rect 43678 682098 43698 682168
rect 43768 682098 43938 682168
rect 44008 682098 44028 682168
rect 43678 680928 44028 682098
rect 44888 682008 45108 682268
rect 44888 681938 44908 682008
rect 44978 681938 45018 682008
rect 45088 681938 45108 682008
rect 44888 681448 45108 681938
rect 44888 681378 44908 681448
rect 44978 681378 45018 681448
rect 45088 681378 45108 681448
rect 44598 681118 44818 681128
rect 44598 680958 44818 680968
rect 43678 680858 43698 680928
rect 43768 680858 43938 680928
rect 44008 680858 44028 680928
rect 43678 680838 44028 680858
rect 43678 680768 43698 680838
rect 43768 680768 43938 680838
rect 44008 680768 44028 680838
rect 42368 680568 42548 680578
rect 42368 680428 42548 680438
rect 43368 680568 43548 680578
rect 43368 680428 43548 680438
rect 43678 680388 44028 680768
rect 44888 680688 45108 681378
rect 44888 680618 44908 680688
rect 44978 680618 45018 680688
rect 45088 680618 45108 680688
rect 44438 680558 44618 680568
rect 44438 680418 44618 680428
rect 43678 680318 43698 680388
rect 43768 680318 43938 680388
rect 44008 680318 44028 680388
rect 43678 680288 44028 680318
rect 44888 680238 45108 680618
rect 45828 682008 46048 682268
rect 45828 681938 45848 682008
rect 45918 681938 45958 682008
rect 46028 681938 46048 682008
rect 45828 681438 46048 681938
rect 45828 681368 45848 681438
rect 45918 681368 45958 681438
rect 46028 681368 46048 681438
rect 45828 680688 46048 681368
rect 46878 682168 47208 682688
rect 47468 682498 47628 682508
rect 47468 682328 47628 682338
rect 48528 682498 48688 682508
rect 48528 682328 48688 682338
rect 46878 682098 46898 682168
rect 46968 682098 47118 682168
rect 47188 682098 47208 682168
rect 46088 681118 46308 681128
rect 46088 680958 46308 680968
rect 45828 680618 45848 680688
rect 45918 680618 45958 680688
rect 46028 680618 46048 680688
rect 45158 680568 45338 680578
rect 45158 680428 45338 680438
rect 45598 680568 45778 680578
rect 45598 680428 45778 680438
rect 44888 680168 44908 680238
rect 44978 680168 45018 680238
rect 45088 680168 45108 680238
rect 44888 680108 45108 680168
rect 45828 680238 46048 680618
rect 46878 680908 47208 682098
rect 46878 680838 46908 680908
rect 46978 680838 47118 680908
rect 47188 680838 47208 680908
rect 46878 680818 47208 680838
rect 46878 680748 46908 680818
rect 46978 680748 47118 680818
rect 47188 680748 47208 680818
rect 46368 680568 46548 680578
rect 46368 680428 46548 680438
rect 46878 680388 47208 680748
rect 47348 680558 47528 680568
rect 47348 680418 47528 680428
rect 48488 680558 48668 680568
rect 48488 680418 48668 680428
rect 46878 680318 46898 680388
rect 46968 680318 47118 680388
rect 47188 680318 47208 680388
rect 46878 680308 47208 680318
rect 45828 680168 45848 680238
rect 45918 680168 45958 680238
rect 46028 680168 46048 680238
rect 45828 680098 46048 680168
rect 42218 678658 42338 678668
rect 42218 678528 42338 678538
rect 48588 678658 48708 678668
rect 48588 678528 48708 678538
rect 42218 675658 42338 675668
rect 42218 675528 42338 675538
rect 48588 675658 48708 675668
rect 48588 675528 48708 675538
rect 42218 672658 42338 672668
rect 42218 672528 42338 672538
rect 48588 672658 48708 672668
rect 48588 672528 48708 672538
rect 42218 669658 42338 669668
rect 42218 669528 42338 669538
rect 48588 669658 48708 669668
rect 48588 669528 48708 669538
rect 42218 666658 42338 666668
rect 42218 666528 42338 666538
rect 48588 666658 48708 666668
rect 48588 666528 48708 666538
rect 42608 665338 43778 665348
rect 42608 664918 43778 664928
rect 44128 665328 45298 665338
rect 44128 664908 45298 664918
rect 45648 665328 46818 665338
rect 45648 664908 46818 664918
rect 47158 665328 48328 665338
rect 47158 664908 48328 664918
rect 524 -800 636 480
rect 1706 -800 1818 480
rect 2888 -800 3000 480
rect 4070 -800 4182 480
rect 5252 -800 5364 480
rect 6434 -800 6546 480
rect 7616 -800 7728 480
rect 8798 -800 8910 480
rect 9980 -800 10092 480
rect 11162 -800 11274 480
rect 12344 -800 12456 480
rect 13526 -800 13638 480
rect 14708 -800 14820 480
rect 15890 -800 16002 480
rect 17072 -800 17184 480
rect 18254 -800 18366 480
rect 19436 -800 19548 480
rect 20618 -800 20730 480
rect 21800 -800 21912 480
rect 22982 -800 23094 480
rect 24164 -800 24276 480
rect 25346 -800 25458 480
rect 26528 -800 26640 480
rect 27710 -800 27822 480
rect 28892 -800 29004 480
rect 30074 -800 30186 480
rect 31256 -800 31368 480
rect 32438 -800 32550 480
rect 33620 -800 33732 480
rect 34802 -800 34914 480
rect 35984 -800 36096 480
rect 37166 -800 37278 480
rect 38348 -800 38460 480
rect 39530 -800 39642 480
rect 40712 -800 40824 480
rect 41894 -800 42006 480
rect 43076 -800 43188 480
rect 44258 -800 44370 480
rect 45440 -800 45552 480
rect 46622 -800 46734 480
rect 47804 -800 47916 480
rect 48986 -800 49098 480
rect 50168 -800 50280 480
rect 51350 -800 51462 480
rect 52532 -800 52644 480
rect 53714 -800 53826 480
rect 54896 -800 55008 480
rect 56078 -800 56190 480
rect 57260 -800 57372 480
rect 58442 -800 58554 480
rect 59624 -800 59736 480
rect 60806 -800 60918 480
rect 61988 -800 62100 480
rect 63170 -800 63282 480
rect 64352 -800 64464 480
rect 65534 -800 65646 480
rect 66716 -800 66828 480
rect 67898 -800 68010 480
rect 69080 -800 69192 480
rect 70262 -800 70374 480
rect 71444 -800 71556 480
rect 72626 -800 72738 480
rect 73808 -800 73920 480
rect 74990 -800 75102 480
rect 76172 -800 76284 480
rect 77354 -800 77466 480
rect 78536 -800 78648 480
rect 79718 -800 79830 480
rect 80900 -800 81012 480
rect 82082 -800 82194 480
rect 83264 -800 83376 480
rect 84446 -800 84558 480
rect 85628 -800 85740 480
rect 86810 -800 86922 480
rect 87992 -800 88104 480
rect 89174 -800 89286 480
rect 90356 -800 90468 480
rect 91538 -800 91650 480
rect 92720 -800 92832 480
rect 93902 -800 94014 480
rect 95084 -800 95196 480
rect 96266 -800 96378 480
rect 97448 -800 97560 480
rect 98630 -800 98742 480
rect 99812 -800 99924 480
rect 100994 -800 101106 480
rect 102176 -800 102288 480
rect 103358 -800 103470 480
rect 104540 -800 104652 480
rect 105722 -800 105834 480
rect 106904 -800 107016 480
rect 108086 -800 108198 480
rect 109268 -800 109380 480
rect 110450 -800 110562 480
rect 111632 -800 111744 480
rect 112814 -800 112926 480
rect 113996 -800 114108 480
rect 115178 -800 115290 480
rect 116360 -800 116472 480
rect 117542 -800 117654 480
rect 118724 -800 118836 480
rect 119906 -800 120018 480
rect 121088 -800 121200 480
rect 122270 -800 122382 480
rect 123452 -800 123564 480
rect 124634 -800 124746 480
rect 125816 -800 125928 480
rect 126998 -800 127110 480
rect 128180 -800 128292 480
rect 129362 -800 129474 480
rect 130544 -800 130656 480
rect 131726 -800 131838 480
rect 132908 -800 133020 480
rect 134090 -800 134202 480
rect 135272 -800 135384 480
rect 136454 -800 136566 480
rect 137636 -800 137748 480
rect 138818 -800 138930 480
rect 140000 -800 140112 480
rect 141182 -800 141294 480
rect 142364 -800 142476 480
rect 143546 -800 143658 480
rect 144728 -800 144840 480
rect 145910 -800 146022 480
rect 147092 -800 147204 480
rect 148274 -800 148386 480
rect 149456 -800 149568 480
rect 150638 -800 150750 480
rect 151820 -800 151932 480
rect 153002 -800 153114 480
rect 154184 -800 154296 480
rect 155366 -800 155478 480
rect 156548 -800 156660 480
rect 157730 -800 157842 480
rect 158912 -800 159024 480
rect 160094 -800 160206 480
rect 161276 -800 161388 480
rect 162458 -800 162570 480
rect 163640 -800 163752 480
rect 164822 -800 164934 480
rect 166004 -800 166116 480
rect 167186 -800 167298 480
rect 168368 -800 168480 480
rect 169550 -800 169662 480
rect 170732 -800 170844 480
rect 171914 -800 172026 480
rect 173096 -800 173208 480
rect 174278 -800 174390 480
rect 175460 -800 175572 480
rect 176642 -800 176754 480
rect 177824 -800 177936 480
rect 179006 -800 179118 480
rect 180188 -800 180300 480
rect 181370 -800 181482 480
rect 182552 -800 182664 480
rect 183734 -800 183846 480
rect 184916 -800 185028 480
rect 186098 -800 186210 480
rect 187280 -800 187392 480
rect 188462 -800 188574 480
rect 189644 -800 189756 480
rect 190826 -800 190938 480
rect 192008 -800 192120 480
rect 193190 -800 193302 480
rect 194372 -800 194484 480
rect 195554 -800 195666 480
rect 196736 -800 196848 480
rect 197918 -800 198030 480
rect 199100 -800 199212 480
rect 200282 -800 200394 480
rect 201464 -800 201576 480
rect 202646 -800 202758 480
rect 203828 -800 203940 480
rect 205010 -800 205122 480
rect 206192 -800 206304 480
rect 207374 -800 207486 480
rect 208556 -800 208668 480
rect 209738 -800 209850 480
rect 210920 -800 211032 480
rect 212102 -800 212214 480
rect 213284 -800 213396 480
rect 214466 -800 214578 480
rect 215648 -800 215760 480
rect 216830 -800 216942 480
rect 218012 -800 218124 480
rect 219194 -800 219306 480
rect 220376 -800 220488 480
rect 221558 -800 221670 480
rect 222740 -800 222852 480
rect 223922 -800 224034 480
rect 225104 -800 225216 480
rect 226286 -800 226398 480
rect 227468 -800 227580 480
rect 228650 -800 228762 480
rect 229832 -800 229944 480
rect 231014 -800 231126 480
rect 232196 -800 232308 480
rect 233378 -800 233490 480
rect 234560 -800 234672 480
rect 235742 -800 235854 480
rect 236924 -800 237036 480
rect 238106 -800 238218 480
rect 239288 -800 239400 480
rect 240470 -800 240582 480
rect 241652 -800 241764 480
rect 242834 -800 242946 480
rect 244016 -800 244128 480
rect 245198 -800 245310 480
rect 246380 -800 246492 480
rect 247562 -800 247674 480
rect 248744 -800 248856 480
rect 249926 -800 250038 480
rect 251108 -800 251220 480
rect 252290 -800 252402 480
rect 253472 -800 253584 480
rect 254654 -800 254766 480
rect 255836 -800 255948 480
rect 257018 -800 257130 480
rect 258200 -800 258312 480
rect 259382 -800 259494 480
rect 260564 -800 260676 480
rect 261746 -800 261858 480
rect 262928 -800 263040 480
rect 264110 -800 264222 480
rect 265292 -800 265404 480
rect 266474 -800 266586 480
rect 267656 -800 267768 480
rect 268838 -800 268950 480
rect 270020 -800 270132 480
rect 271202 -800 271314 480
rect 272384 -800 272496 480
rect 273566 -800 273678 480
rect 274748 -800 274860 480
rect 275930 -800 276042 480
rect 277112 -800 277224 480
rect 278294 -800 278406 480
rect 279476 -800 279588 480
rect 280658 -800 280770 480
rect 281840 -800 281952 480
rect 283022 -800 283134 480
rect 284204 -800 284316 480
rect 285386 -800 285498 480
rect 286568 -800 286680 480
rect 287750 -800 287862 480
rect 288932 -800 289044 480
rect 290114 -800 290226 480
rect 291296 -800 291408 480
rect 292478 -800 292590 480
rect 293660 -800 293772 480
rect 294842 -800 294954 480
rect 296024 -800 296136 480
rect 297206 -800 297318 480
rect 298388 -800 298500 480
rect 299570 -800 299682 480
rect 300752 -800 300864 480
rect 301934 -800 302046 480
rect 303116 -800 303228 480
rect 304298 -800 304410 480
rect 305480 -800 305592 480
rect 306662 -800 306774 480
rect 307844 -800 307956 480
rect 309026 -800 309138 480
rect 310208 -800 310320 480
rect 311390 -800 311502 480
rect 312572 -800 312684 480
rect 313754 -800 313866 480
rect 314936 -800 315048 480
rect 316118 -800 316230 480
rect 317300 -800 317412 480
rect 318482 -800 318594 480
rect 319664 -800 319776 480
rect 320846 -800 320958 480
rect 322028 -800 322140 480
rect 323210 -800 323322 480
rect 324392 -800 324504 480
rect 325574 -800 325686 480
rect 326756 -800 326868 480
rect 327938 -800 328050 480
rect 329120 -800 329232 480
rect 330302 -800 330414 480
rect 331484 -800 331596 480
rect 332666 -800 332778 480
rect 333848 -800 333960 480
rect 335030 -800 335142 480
rect 336212 -800 336324 480
rect 337394 -800 337506 480
rect 338576 -800 338688 480
rect 339758 -800 339870 480
rect 340940 -800 341052 480
rect 342122 -800 342234 480
rect 343304 -800 343416 480
rect 344486 -800 344598 480
rect 345668 -800 345780 480
rect 346850 -800 346962 480
rect 348032 -800 348144 480
rect 349214 -800 349326 480
rect 350396 -800 350508 480
rect 351578 -800 351690 480
rect 352760 -800 352872 480
rect 353942 -800 354054 480
rect 355124 -800 355236 480
rect 356306 -800 356418 480
rect 357488 -800 357600 480
rect 358670 -800 358782 480
rect 359852 -800 359964 480
rect 361034 -800 361146 480
rect 362216 -800 362328 480
rect 363398 -800 363510 480
rect 364580 -800 364692 480
rect 365762 -800 365874 480
rect 366944 -800 367056 480
rect 368126 -800 368238 480
rect 369308 -800 369420 480
rect 370490 -800 370602 480
rect 371672 -800 371784 480
rect 372854 -800 372966 480
rect 374036 -800 374148 480
rect 375218 -800 375330 480
rect 376400 -800 376512 480
rect 377582 -800 377694 480
rect 378764 -800 378876 480
rect 379946 -800 380058 480
rect 381128 -800 381240 480
rect 382310 -800 382422 480
rect 383492 -800 383604 480
rect 384674 -800 384786 480
rect 385856 -800 385968 480
rect 387038 -800 387150 480
rect 388220 -800 388332 480
rect 389402 -800 389514 480
rect 390584 -800 390696 480
rect 391766 -800 391878 480
rect 392948 -800 393060 480
rect 394130 -800 394242 480
rect 395312 -800 395424 480
rect 396494 -800 396606 480
rect 397676 -800 397788 480
rect 398858 -800 398970 480
rect 400040 -800 400152 480
rect 401222 -800 401334 480
rect 402404 -800 402516 480
rect 403586 -800 403698 480
rect 404768 -800 404880 480
rect 405950 -800 406062 480
rect 407132 -800 407244 480
rect 408314 -800 408426 480
rect 409496 -800 409608 480
rect 410678 -800 410790 480
rect 411860 -800 411972 480
rect 413042 -800 413154 480
rect 414224 -800 414336 480
rect 415406 -800 415518 480
rect 416588 -800 416700 480
rect 417770 -800 417882 480
rect 418952 -800 419064 480
rect 420134 -800 420246 480
rect 421316 -800 421428 480
rect 422498 -800 422610 480
rect 423680 -800 423792 480
rect 424862 -800 424974 480
rect 426044 -800 426156 480
rect 427226 -800 427338 480
rect 428408 -800 428520 480
rect 429590 -800 429702 480
rect 430772 -800 430884 480
rect 431954 -800 432066 480
rect 433136 -800 433248 480
rect 434318 -800 434430 480
rect 435500 -800 435612 480
rect 436682 -800 436794 480
rect 437864 -800 437976 480
rect 439046 -800 439158 480
rect 440228 -800 440340 480
rect 441410 -800 441522 480
rect 442592 -800 442704 480
rect 443774 -800 443886 480
rect 444956 -800 445068 480
rect 446138 -800 446250 480
rect 447320 -800 447432 480
rect 448502 -800 448614 480
rect 449684 -800 449796 480
rect 450866 -800 450978 480
rect 452048 -800 452160 480
rect 453230 -800 453342 480
rect 454412 -800 454524 480
rect 455594 -800 455706 480
rect 456776 -800 456888 480
rect 457958 -800 458070 480
rect 459140 -800 459252 480
rect 460322 -800 460434 480
rect 461504 -800 461616 480
rect 462686 -800 462798 480
rect 463868 -800 463980 480
rect 465050 -800 465162 480
rect 466232 -800 466344 480
rect 467414 -800 467526 480
rect 468596 -800 468708 480
rect 469778 -800 469890 480
rect 470960 -800 471072 480
rect 472142 -800 472254 480
rect 473324 -800 473436 480
rect 474506 -800 474618 480
rect 475688 -800 475800 480
rect 476870 -800 476982 480
rect 478052 -800 478164 480
rect 479234 -800 479346 480
rect 480416 -800 480528 480
rect 481598 -800 481710 480
rect 482780 -800 482892 480
rect 483962 -800 484074 480
rect 485144 -800 485256 480
rect 486326 -800 486438 480
rect 487508 -800 487620 480
rect 488690 -800 488802 480
rect 489872 -800 489984 480
rect 491054 -800 491166 480
rect 492236 -800 492348 480
rect 493418 -800 493530 480
rect 494600 -800 494712 480
rect 495782 -800 495894 480
rect 496964 -800 497076 480
rect 498146 -800 498258 480
rect 499328 -800 499440 480
rect 500510 -800 500622 480
rect 501692 -800 501804 480
rect 502874 -800 502986 480
rect 504056 -800 504168 480
rect 505238 -800 505350 480
rect 506420 -800 506532 480
rect 507602 -800 507714 480
rect 508784 -800 508896 480
rect 509966 -800 510078 480
rect 511148 -800 511260 480
rect 512330 -800 512442 480
rect 513512 -800 513624 480
rect 514694 -800 514806 480
rect 515876 -800 515988 480
rect 517058 -800 517170 480
rect 518240 -800 518352 480
rect 519422 -800 519534 480
rect 520604 -800 520716 480
rect 521786 -800 521898 480
rect 522968 -800 523080 480
rect 524150 -800 524262 480
rect 525332 -800 525444 480
rect 526514 -800 526626 480
rect 527696 -800 527808 480
rect 528878 -800 528990 480
rect 530060 -800 530172 480
rect 531242 -800 531354 480
rect 532424 -800 532536 480
rect 533606 -800 533718 480
rect 534788 -800 534900 480
rect 535970 -800 536082 480
rect 537152 -800 537264 480
rect 538334 -800 538446 480
rect 539516 -800 539628 480
rect 540698 -800 540810 480
rect 541880 -800 541992 480
rect 543062 -800 543174 480
rect 544244 -800 544356 480
rect 545426 -800 545538 480
rect 546608 -800 546720 480
rect 547790 -800 547902 480
rect 548972 -800 549084 480
rect 550154 -800 550266 480
rect 551336 -800 551448 480
rect 552518 -800 552630 480
rect 553700 -800 553812 480
rect 554882 -800 554994 480
rect 556064 -800 556176 480
rect 557246 -800 557358 480
rect 558428 -800 558540 480
rect 559610 -800 559722 480
rect 560792 -800 560904 480
rect 561974 -800 562086 480
rect 563156 -800 563268 480
rect 564338 -800 564450 480
rect 565520 -800 565632 480
rect 566702 -800 566814 480
rect 567884 -800 567996 480
rect 569066 -800 569178 480
rect 570248 -800 570360 480
rect 571430 -800 571542 480
rect 572612 -800 572724 480
rect 573794 -800 573906 480
rect 574976 -800 575088 480
rect 576158 -800 576270 480
rect 577340 -800 577452 480
rect 578522 -800 578634 480
rect 579704 -800 579816 480
rect 580886 -800 580998 480
rect 582068 -800 582180 480
rect 583250 -800 583362 480
<< via2 >>
rect 44798 694608 45068 694878
rect 45848 694608 46118 694878
rect 42278 694328 42348 694398
rect 42588 694328 42658 694398
rect 42908 694328 42978 694398
rect 43228 694328 43298 694398
rect 43538 694328 43608 694398
rect 43858 694328 43928 694398
rect 44168 694328 44238 694398
rect 44488 694328 44558 694398
rect 44808 694328 44878 694398
rect 45118 694328 45188 694398
rect 45438 694328 45508 694398
rect 45748 694328 45818 694398
rect 46068 694328 46138 694398
rect 46388 694328 46458 694398
rect 46698 694328 46768 694398
rect 47018 694328 47088 694398
rect 47338 694328 47408 694398
rect 47648 694328 47718 694398
rect 47968 694328 48038 694398
rect 48278 694328 48348 694398
rect 48598 694328 48668 694398
rect 37738 694088 37808 694158
rect 42278 694088 42348 694158
rect 42588 694088 42658 694158
rect 42908 694088 42978 694158
rect 43228 694088 43298 694158
rect 43538 694088 43608 694158
rect 43858 694088 43928 694158
rect 44168 694088 44238 694158
rect 44488 694088 44558 694158
rect 44808 694088 44878 694158
rect 45118 694088 45188 694158
rect 45438 694088 45508 694158
rect 45748 694088 45818 694158
rect 46068 694088 46138 694158
rect 46388 694088 46458 694158
rect 46698 694088 46768 694158
rect 47018 694088 47088 694158
rect 47338 694088 47408 694158
rect 47648 694088 47718 694158
rect 47968 694088 48038 694158
rect 48278 694088 48348 694158
rect 48598 694088 48668 694158
rect 53128 694088 53198 694158
rect 37628 693978 37698 694048
rect 53238 693978 53308 694048
rect 42428 693718 42498 693788
rect 42748 693718 42818 693788
rect 43068 693718 43138 693788
rect 43378 693718 43448 693788
rect 43698 693718 43768 693788
rect 44018 693718 44088 693788
rect 44328 693718 44398 693788
rect 44648 693718 44718 693788
rect 44958 693718 45028 693788
rect 45278 693718 45348 693788
rect 45598 693718 45668 693788
rect 45908 693718 45978 693788
rect 46228 693718 46298 693788
rect 46548 693718 46618 693788
rect 46858 693718 46928 693788
rect 47178 693718 47248 693788
rect 47488 693718 47558 693788
rect 47808 693718 47878 693788
rect 48128 693718 48198 693788
rect 48438 693718 48508 693788
rect 42428 693478 42498 693548
rect 42748 693478 42818 693548
rect 43068 693478 43138 693548
rect 43378 693478 43448 693548
rect 43698 693478 43768 693548
rect 44018 693478 44088 693548
rect 44328 693478 44398 693548
rect 44648 693478 44718 693548
rect 44958 693478 45028 693548
rect 45278 693478 45348 693548
rect 45598 693478 45668 693548
rect 45908 693478 45978 693548
rect 46228 693478 46298 693548
rect 46548 693478 46618 693548
rect 46858 693478 46928 693548
rect 47178 693478 47248 693548
rect 47488 693478 47558 693548
rect 47808 693478 47878 693548
rect 48128 693478 48198 693548
rect 42428 693108 42498 693178
rect 39578 692598 39758 692698
rect 39998 692598 40178 692698
rect 44798 692968 45068 693238
rect 45848 692968 46118 693238
rect 43938 692658 44008 692728
rect 44248 692658 44318 692728
rect 44568 692658 44638 692728
rect 44878 692658 44948 692728
rect 45198 692658 45268 692728
rect 45518 692658 45588 692728
rect 45828 692658 45898 692728
rect 46148 692658 46218 692728
rect 46468 692658 46538 692728
rect 46778 692658 46848 692728
rect 47098 692658 47168 692728
rect 43938 692448 44008 692518
rect 44248 692448 44318 692518
rect 44568 692448 44638 692518
rect 44878 692448 44948 692518
rect 45198 692448 45268 692518
rect 45518 692448 45588 692518
rect 45828 692448 45898 692518
rect 46148 692448 46218 692518
rect 46468 692448 46538 692518
rect 46778 692448 46848 692518
rect 47098 692448 47168 692518
rect 43408 691998 43488 692078
rect 43778 692018 43848 692088
rect 44088 692018 44158 692088
rect 44408 692018 44478 692088
rect 44728 692018 44798 692088
rect 45038 692018 45108 692088
rect 45358 692018 45428 692088
rect 45668 692018 45738 692088
rect 45988 692018 46058 692088
rect 46308 692018 46378 692088
rect 46618 692018 46688 692088
rect 46938 692018 47008 692088
rect 43408 691818 43488 691898
rect 47468 691998 47548 692078
rect 43778 691808 43848 691878
rect 44088 691808 44158 691878
rect 44408 691808 44478 691878
rect 44728 691808 44798 691878
rect 45038 691808 45108 691878
rect 45358 691808 45428 691878
rect 45668 691808 45738 691878
rect 45988 691808 46058 691878
rect 46308 691808 46378 691878
rect 46618 691808 46688 691878
rect 46938 691808 47008 691878
rect 47468 691818 47548 691898
rect 44588 691368 44848 691628
rect 46088 691368 46348 691628
rect 43938 691108 44008 691178
rect 44248 691108 44318 691178
rect 44568 691108 44638 691178
rect 44888 691108 44958 691178
rect 45198 691108 45268 691178
rect 45518 691108 45588 691178
rect 45828 691108 45898 691178
rect 46148 691108 46218 691178
rect 46468 691108 46538 691178
rect 46778 691108 46848 691178
rect 47098 691108 47168 691178
rect 43938 690898 44008 690968
rect 44248 690898 44318 690968
rect 44568 690898 44638 690968
rect 44888 690898 44958 690968
rect 45198 690898 45268 690968
rect 45518 690898 45588 690968
rect 45828 690898 45898 690968
rect 46148 690898 46218 690968
rect 46468 690898 46538 690968
rect 46778 690898 46848 690968
rect 47098 690898 47168 690968
rect 43778 690478 43848 690548
rect 44098 690478 44168 690548
rect 43778 690268 43848 690338
rect 44408 690478 44478 690548
rect 44728 690478 44798 690548
rect 45038 690478 45108 690548
rect 45358 690478 45428 690548
rect 45678 690478 45748 690548
rect 45988 690478 46058 690548
rect 46308 690478 46378 690548
rect 46618 690478 46688 690548
rect 44098 690268 44168 690338
rect 43388 689488 43508 689608
rect 43388 689268 43508 689388
rect 43628 688928 43748 689048
rect 43628 688708 43748 688828
rect 43628 687968 43748 688088
rect 43340 687760 43460 687920
rect 43340 687560 43460 687720
rect 43628 687748 43748 687868
rect 42428 686498 42498 686568
rect 42428 686338 42498 686408
rect 44408 690268 44478 690338
rect 44728 690268 44798 690338
rect 45038 690268 45108 690338
rect 45358 690268 45428 690338
rect 45678 690268 45748 690338
rect 45988 690268 46058 690338
rect 46308 690268 46378 690338
rect 46938 690478 47008 690548
rect 46618 690268 46688 690338
rect 45048 689548 45118 689618
rect 45368 689548 45438 689618
rect 45678 689548 45748 689618
rect 45998 689548 46068 689618
rect 45048 689258 45118 689328
rect 45368 689258 45438 689328
rect 45678 689258 45748 689328
rect 45998 689258 46068 689328
rect 44888 688988 44958 689058
rect 45208 688988 45278 689058
rect 45528 688988 45598 689058
rect 45838 688988 45908 689058
rect 44888 688698 44958 688768
rect 45208 688698 45278 688768
rect 45528 688698 45598 688768
rect 45838 688698 45908 688768
rect 45348 688268 45608 688528
rect 45048 688028 45118 688098
rect 45368 688028 45438 688098
rect 45678 688028 45748 688098
rect 45998 688028 46068 688098
rect 45048 687738 45118 687808
rect 45368 687738 45438 687808
rect 45678 687738 45748 687808
rect 45998 687738 46068 687808
rect 44098 687448 44168 687518
rect 44888 687468 44958 687538
rect 45208 687468 45278 687538
rect 45528 687468 45598 687538
rect 45838 687468 45908 687538
rect 46938 690268 47008 690338
rect 47448 689488 47568 689608
rect 48438 693108 48508 693178
rect 47448 689268 47568 689388
rect 47960 689260 48100 689380
rect 47960 689100 48100 689220
rect 44098 687198 44168 687268
rect 46618 687448 46688 687518
rect 44888 687178 44958 687248
rect 45208 687178 45278 687248
rect 45528 687178 45598 687248
rect 45838 687178 45908 687248
rect 46618 687198 46688 687268
rect 47208 688928 47328 689048
rect 47960 688920 48100 689040
rect 47208 688708 47328 688828
rect 47208 687968 47328 688088
rect 47208 687748 47328 687868
rect 45348 686748 45608 687008
rect 43888 686508 43958 686578
rect 44408 686508 44478 686578
rect 44928 686508 44998 686578
rect 45438 686508 45508 686578
rect 45958 686508 46028 686578
rect 46468 686508 46538 686578
rect 46988 686508 47058 686578
rect 43888 686328 43958 686398
rect 44408 686328 44478 686398
rect 44928 686328 44998 686398
rect 45438 686328 45508 686398
rect 45958 686328 46028 686398
rect 46468 686328 46538 686398
rect 46988 686328 47058 686398
rect 44148 685838 44218 685908
rect 44668 685838 44738 685908
rect 45178 685838 45248 685908
rect 45698 685838 45768 685908
rect 46218 685838 46288 685908
rect 46728 685838 46798 685908
rect 44148 685658 44218 685728
rect 44668 685658 44738 685728
rect 45178 685658 45248 685728
rect 45698 685658 45768 685728
rect 46218 685658 46288 685728
rect 46728 685658 46798 685728
rect 45348 685238 45598 685488
rect 43638 684988 43708 685058
rect 44148 684988 44218 685058
rect 44668 684988 44738 685058
rect 45188 684988 45258 685058
rect 45698 684988 45768 685058
rect 46218 684988 46288 685058
rect 46728 684988 46798 685058
rect 47248 684988 47318 685058
rect 43638 684808 43708 684878
rect 44148 684808 44218 684878
rect 44668 684808 44738 684878
rect 45188 684808 45258 684878
rect 45698 684808 45768 684878
rect 46218 684808 46288 684878
rect 46728 684808 46798 684878
rect 47248 684808 47318 684878
rect 50828 692598 51008 692698
rect 51248 692598 51428 692698
rect 48438 686498 48508 686568
rect 48438 686338 48508 686408
rect 43898 684318 43968 684388
rect 44408 684318 44478 684388
rect 44928 684318 44998 684388
rect 45438 684318 45508 684388
rect 45958 684318 46028 684388
rect 46478 684318 46548 684388
rect 46988 684318 47058 684388
rect 43898 684138 43968 684208
rect 44408 684138 44478 684208
rect 44928 684138 44998 684208
rect 45438 684138 45508 684208
rect 45958 684138 46028 684208
rect 46478 684138 46548 684208
rect 46988 684138 47058 684208
rect 45348 683708 45598 683958
rect 42308 682918 42468 683078
rect 43308 682918 43468 683078
rect 44788 682918 44948 683078
rect 42308 682338 42468 682498
rect 43308 682338 43468 682498
rect 44788 682338 44948 682498
rect 46008 682918 46168 683078
rect 47468 682918 47628 683078
rect 48528 682918 48688 683078
rect 46008 682338 46168 682498
rect 44598 680968 44818 681118
rect 42368 680438 42548 680568
rect 43368 680438 43548 680568
rect 44438 680428 44618 680558
rect 47468 682338 47628 682498
rect 48528 682338 48688 682498
rect 46088 680968 46308 681118
rect 45158 680438 45338 680568
rect 45598 680438 45778 680568
rect 46368 680438 46548 680568
rect 47348 680428 47528 680558
rect 48488 680428 48668 680558
rect 42218 678538 42338 678658
rect 48588 678538 48708 678658
rect 42218 675538 42338 675658
rect 48588 675538 48708 675658
rect 42218 672538 42338 672658
rect 48588 672538 48708 672658
rect 42218 669538 42338 669658
rect 48588 669538 48708 669658
rect 42218 666538 42338 666658
rect 48588 666538 48708 666658
rect 42608 664928 43778 665338
rect 44128 664918 45298 665328
rect 45648 664918 46818 665328
rect 47158 664918 48328 665328
<< metal3 >>
rect 16194 703000 21194 704800
rect 16194 702740 18100 703000
rect 18340 702740 18520 703000
rect 18760 702740 18940 703000
rect 19180 702740 21194 703000
rect 16194 702600 21194 702740
rect 16194 702340 18100 702600
rect 18340 702340 18520 702600
rect 18760 702340 18940 702600
rect 19180 702340 21194 702600
rect 16194 702300 21194 702340
rect 68194 702880 73194 704800
rect 68194 702660 70220 702880
rect 70440 702660 70640 702880
rect 70860 702660 71080 702880
rect 71300 702660 73194 702880
rect 68194 702560 73194 702660
rect 68194 702340 70220 702560
rect 70440 702340 70640 702560
rect 70860 702340 71080 702560
rect 71300 702340 73194 702560
rect 68194 702300 73194 702340
rect 120194 702300 125194 704800
rect 165594 702300 170594 704800
rect 170894 702300 173094 704800
rect 173394 702300 175594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 222594 702300 224794 704800
rect 225094 702300 227294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 324294 702300 326494 704800
rect 326794 702300 328994 704800
rect 329294 702300 334294 704800
rect 413394 702300 418394 704800
rect 465394 702300 470394 704800
rect 510594 702500 515394 704800
rect 510594 702340 515400 702500
rect 520594 702400 525394 704800
rect 520594 702340 525400 702400
rect 38078 700347 41478 700367
rect 38078 700283 38106 700347
rect 41450 700283 41478 700347
rect 38078 696868 41478 700283
rect 41878 700347 45278 700367
rect 41878 700283 41906 700347
rect 45250 700283 45278 700347
rect 41878 696868 45278 700283
rect 45678 700347 49078 700367
rect 45678 700283 45706 700347
rect 49050 700283 49078 700347
rect 45678 696868 49078 700283
rect 49478 700347 52878 700367
rect 49478 700283 49506 700347
rect 52850 700283 52878 700347
rect 49478 696868 52878 700283
rect 465520 698972 470020 702300
rect 510600 700384 515400 702340
rect 520600 700384 525400 702340
rect 566594 702300 571594 704800
rect 568220 700736 569760 702300
rect 1600 696380 49440 696400
rect 1600 696200 41600 696380
rect 41800 696360 49440 696380
rect 41800 696200 49180 696360
rect 1600 696180 49180 696200
rect 49380 696180 49440 696360
rect 1600 695920 49440 696180
rect 1600 695900 49180 695920
rect 1600 695720 41600 695900
rect 41800 695740 49180 695900
rect 49380 695740 49440 695920
rect 41800 695720 49440 695740
rect 1600 695700 49440 695720
rect 1600 689400 4500 695700
rect 44788 694878 45078 694883
rect 44788 694608 44798 694878
rect 45068 694608 45078 694878
rect 44788 694603 45078 694608
rect 45838 694878 46128 694883
rect 45838 694608 45848 694878
rect 46118 694608 46128 694878
rect 45838 694603 46128 694608
rect 42278 694403 48668 694408
rect 42268 694398 48678 694403
rect 42268 694328 42278 694398
rect 42348 694328 42588 694398
rect 42658 694368 42908 694398
rect 42268 694323 42658 694328
rect 37608 694158 37828 694178
rect 42278 694163 42658 694323
rect 37608 694088 37738 694158
rect 37808 694088 37828 694158
rect 37608 694048 37828 694088
rect 42268 694158 42658 694163
rect 42268 694088 42278 694158
rect 42348 694088 42588 694158
rect 42978 694328 43228 694398
rect 43298 694328 43538 694398
rect 43608 694328 43858 694398
rect 43928 694328 44168 694398
rect 44238 694328 44488 694398
rect 44558 694368 44808 694398
rect 42908 694158 44558 694328
rect 42658 694088 42908 694118
rect 42978 694088 43228 694158
rect 43298 694088 43538 694158
rect 43608 694088 43858 694158
rect 43928 694088 44168 694158
rect 44238 694088 44488 694158
rect 44878 694328 45118 694398
rect 45188 694328 45438 694398
rect 45508 694328 45748 694398
rect 45818 694328 46068 694398
rect 46138 694368 46388 694398
rect 44808 694158 46138 694328
rect 44558 694088 44808 694118
rect 44878 694088 45118 694158
rect 45188 694088 45438 694158
rect 45508 694088 45748 694158
rect 45818 694088 46068 694158
rect 46458 694328 46698 694398
rect 46768 694328 47018 694398
rect 47088 694328 47338 694398
rect 47408 694328 47648 694398
rect 47718 694328 47968 694398
rect 48038 694378 48278 694398
rect 48348 694328 48598 694398
rect 48668 694328 48678 694398
rect 46388 694158 48038 694328
rect 48288 694323 48678 694328
rect 48288 694163 48668 694323
rect 48288 694158 48678 694163
rect 46138 694088 46388 694118
rect 46458 694088 46698 694158
rect 46768 694088 47018 694158
rect 47088 694088 47338 694158
rect 47408 694088 47648 694158
rect 47718 694088 47968 694158
rect 48038 694088 48278 694128
rect 48348 694088 48598 694158
rect 48668 694088 48678 694158
rect 42268 694083 48678 694088
rect 53108 694158 53328 694178
rect 53108 694088 53128 694158
rect 53198 694088 53328 694158
rect 42278 694078 48668 694083
rect 37608 693978 37628 694048
rect 37698 693978 37828 694048
rect 37608 693958 37828 693978
rect 53108 694048 53328 694088
rect 53108 693978 53238 694048
rect 53308 693978 53328 694048
rect 53108 693958 53328 693978
rect 42278 693788 48668 693798
rect 42278 693718 42428 693788
rect 42498 693718 42748 693788
rect 42818 693718 43068 693788
rect 43138 693718 43378 693788
rect 43448 693718 43698 693788
rect 43768 693718 44018 693788
rect 44088 693718 44328 693788
rect 44398 693718 44648 693788
rect 44718 693718 44958 693788
rect 45028 693718 45278 693788
rect 45348 693718 45598 693788
rect 45668 693718 45908 693788
rect 45978 693718 46228 693788
rect 46298 693718 46548 693788
rect 46618 693718 46858 693788
rect 46928 693718 47178 693788
rect 47248 693718 47488 693788
rect 47558 693718 47808 693788
rect 47878 693718 48128 693788
rect 48198 693718 48438 693788
rect 48508 693718 48668 693788
rect 42278 693548 48668 693718
rect 42278 693478 42428 693548
rect 42498 693478 42748 693548
rect 42818 693478 43068 693548
rect 43138 693478 43378 693548
rect 43448 693478 43698 693548
rect 43768 693478 44018 693548
rect 44088 693478 44328 693548
rect 44398 693478 44648 693548
rect 44718 693478 44958 693548
rect 45028 693478 45278 693548
rect 45348 693478 45598 693548
rect 45668 693478 45908 693548
rect 45978 693478 46228 693548
rect 46298 693478 46548 693548
rect 46618 693478 46858 693548
rect 46928 693478 47178 693548
rect 47248 693478 47488 693548
rect 47558 693478 47808 693548
rect 47878 693478 48128 693548
rect 48198 693478 48668 693548
rect 42278 693468 48668 693478
rect 44788 693238 45078 693243
rect 41508 693198 42528 693218
rect 41508 693098 41528 693198
rect 41618 693098 41718 693198
rect 41808 693178 42528 693198
rect 41808 693108 42428 693178
rect 42498 693108 42528 693178
rect 41808 693098 42528 693108
rect 41508 693078 42528 693098
rect 44788 692968 44798 693238
rect 45068 692968 45078 693238
rect 44788 692963 45078 692968
rect 45838 693238 46128 693243
rect 45838 692968 45848 693238
rect 46118 692968 46128 693238
rect 48408 693198 49438 693218
rect 48408 693178 49138 693198
rect 48408 693108 48438 693178
rect 48508 693108 49138 693178
rect 48408 693098 49138 693108
rect 49228 693098 49328 693198
rect 49418 693098 49438 693198
rect 48408 693078 49438 693098
rect 45838 692963 46128 692968
rect 43778 692733 47168 692738
rect 43778 692728 47178 692733
rect 39568 692698 39768 692703
rect 39568 692598 39578 692698
rect 39758 692598 39768 692698
rect 39568 692593 39768 692598
rect 39988 692698 40188 692703
rect 39988 692598 39998 692698
rect 40178 692598 40188 692698
rect 39988 692593 40188 692598
rect 43778 692658 43938 692728
rect 44008 692718 44248 692728
rect 44318 692658 44568 692728
rect 44638 692658 44878 692728
rect 44948 692658 45198 692728
rect 45268 692718 45518 692728
rect 45588 692658 45828 692728
rect 45898 692658 46148 692728
rect 46218 692658 46468 692728
rect 46538 692718 46778 692728
rect 46848 692658 47098 692728
rect 47168 692658 47178 692728
rect 43778 692518 43998 692658
rect 44258 692518 45258 692658
rect 45518 692518 46528 692658
rect 46788 692653 47178 692658
rect 50818 692698 51018 692703
rect 46788 692523 47168 692653
rect 50818 692598 50828 692698
rect 51008 692598 51018 692698
rect 50818 692593 51018 692598
rect 51238 692698 51438 692703
rect 51238 692598 51248 692698
rect 51428 692598 51438 692698
rect 51238 692593 51438 692598
rect 46788 692518 47178 692523
rect 43778 692448 43938 692518
rect 44008 692448 44248 692458
rect 44318 692448 44568 692518
rect 44638 692448 44878 692518
rect 44948 692448 45198 692518
rect 45268 692448 45518 692458
rect 45588 692448 45828 692518
rect 45898 692448 46148 692518
rect 46218 692448 46468 692518
rect 46538 692448 46778 692458
rect 46848 692448 47098 692518
rect 47168 692448 47178 692518
rect 43778 692443 47178 692448
rect 43778 692438 47168 692443
rect 43368 692088 47588 692098
rect 43368 692078 43778 692088
rect 43368 691998 43408 692078
rect 43488 692018 43778 692078
rect 43848 692018 44088 692088
rect 44158 692018 44408 692088
rect 44478 692018 44728 692088
rect 44798 692018 45038 692088
rect 45108 692018 45358 692088
rect 45428 692018 45668 692088
rect 45738 692018 45988 692088
rect 46058 692018 46308 692088
rect 46378 692018 46618 692088
rect 46688 692018 46938 692088
rect 47008 692078 47588 692088
rect 47008 692018 47468 692078
rect 43488 691998 47468 692018
rect 47548 691998 47588 692078
rect 43368 691898 47588 691998
rect 43368 691818 43408 691898
rect 43488 691878 47468 691898
rect 43488 691818 43778 691878
rect 43368 691808 43778 691818
rect 43848 691808 44088 691878
rect 44158 691808 44408 691878
rect 44478 691808 44728 691878
rect 44798 691808 45038 691878
rect 45108 691808 45358 691878
rect 45428 691808 45668 691878
rect 45738 691808 45988 691878
rect 46058 691808 46308 691878
rect 46378 691808 46618 691878
rect 46688 691808 46938 691878
rect 47008 691818 47468 691878
rect 47548 691818 47588 691898
rect 47008 691808 47588 691818
rect 43368 691798 47588 691808
rect 44578 691628 44858 691633
rect 44578 691368 44588 691628
rect 44848 691368 44858 691628
rect 44578 691363 44858 691368
rect 46078 691628 46358 691633
rect 46078 691368 46088 691628
rect 46348 691368 46358 691628
rect 46078 691363 46358 691368
rect 43778 691183 47168 691188
rect 43778 691178 47178 691183
rect 43778 691108 43938 691178
rect 44008 691168 44248 691178
rect 44318 691108 44568 691178
rect 44638 691108 44888 691178
rect 44958 691108 45198 691178
rect 45268 691168 45518 691178
rect 45588 691108 45828 691178
rect 45898 691108 46148 691178
rect 46218 691108 46468 691178
rect 46538 691168 46778 691178
rect 46848 691108 47098 691178
rect 47168 691108 47178 691178
rect 43778 690968 43998 691108
rect 44258 690968 45258 691108
rect 45518 690968 46528 691108
rect 46788 691103 47178 691108
rect 46788 690973 47168 691103
rect 46788 690968 47178 690973
rect 43778 690898 43938 690968
rect 44008 690898 44248 690908
rect 44318 690898 44568 690968
rect 44638 690898 44888 690968
rect 44958 690898 45198 690968
rect 45268 690898 45518 690908
rect 45588 690898 45828 690968
rect 45898 690898 46148 690968
rect 46218 690898 46468 690968
rect 46538 690898 46778 690908
rect 46848 690898 47098 690968
rect 47168 690898 47178 690968
rect 43778 690893 47178 690898
rect 43778 690888 47168 690893
rect 43778 690553 47168 690558
rect 43768 690548 47168 690553
rect 43768 690478 43778 690548
rect 43848 690478 44098 690548
rect 44168 690478 44408 690548
rect 44478 690478 44728 690548
rect 44798 690478 45038 690548
rect 45108 690478 45358 690548
rect 45428 690478 45678 690548
rect 45748 690478 45988 690548
rect 46058 690478 46308 690548
rect 46378 690478 46618 690548
rect 46688 690478 46938 690548
rect 47008 690478 47168 690548
rect 43768 690473 47168 690478
rect 43778 690343 47168 690473
rect 43768 690338 47168 690343
rect 43768 690268 43778 690338
rect 43848 690268 44098 690338
rect 44168 690268 44408 690338
rect 44478 690268 44728 690338
rect 44798 690268 45038 690338
rect 45108 690268 45358 690338
rect 45428 690268 45678 690338
rect 45748 690268 45988 690338
rect 46058 690268 46308 690338
rect 46378 690268 46618 690338
rect 46688 690268 46938 690338
rect 47008 690268 47168 690338
rect 43768 690263 47168 690268
rect 43778 690258 47168 690263
rect 1640 687800 4500 689400
rect 43368 689618 47588 689628
rect 43368 689608 45048 689618
rect 43368 689488 43388 689608
rect 43508 689548 45048 689608
rect 45118 689548 45368 689618
rect 45438 689548 45678 689618
rect 45748 689548 45998 689618
rect 46068 689608 47588 689618
rect 46068 689548 47448 689608
rect 43508 689488 47448 689548
rect 47568 689488 47588 689608
rect 43368 689388 47588 689488
rect 70180 689540 71340 689560
rect 70180 689400 70240 689540
rect 43368 689268 43388 689388
rect 43508 689328 47448 689388
rect 43508 689268 45048 689328
rect 43368 689258 45048 689268
rect 45118 689258 45368 689328
rect 45438 689258 45678 689328
rect 45748 689258 45998 689328
rect 46068 689268 47448 689328
rect 47568 689268 47588 689388
rect 46068 689258 47588 689268
rect 43368 689248 47588 689258
rect 47940 689380 70240 689400
rect 47940 689260 47960 689380
rect 48100 689320 70240 689380
rect 70460 689320 70640 689540
rect 70860 689320 71060 689540
rect 71280 689320 71340 689540
rect 48100 689280 71340 689320
rect 48100 689260 70240 689280
rect 47940 689220 70240 689260
rect 47940 689100 47960 689220
rect 48100 689100 70240 689220
rect 43608 689058 47348 689068
rect 43608 689048 44888 689058
rect 43608 688928 43628 689048
rect 43748 688988 44888 689048
rect 44958 688988 45208 689058
rect 45278 688988 45528 689058
rect 45598 688988 45838 689058
rect 45908 689048 47348 689058
rect 45908 688988 47208 689048
rect 43748 688928 47208 688988
rect 47328 688928 47348 689048
rect 43608 688828 47348 688928
rect 47940 689060 70240 689100
rect 70460 689060 70640 689280
rect 70860 689060 71060 689280
rect 71280 689060 71340 689280
rect 47940 689040 71340 689060
rect 47940 688920 47960 689040
rect 48100 688940 71340 689040
rect 48100 688920 48120 688940
rect 47940 688900 48120 688920
rect 43608 688708 43628 688828
rect 43748 688768 47208 688828
rect 43748 688708 44888 688768
rect 43608 688698 44888 688708
rect 44958 688698 45208 688768
rect 45278 688698 45528 688768
rect 45598 688698 45838 688768
rect 45908 688708 47208 688768
rect 47328 688708 47348 688828
rect 45908 688698 47348 688708
rect 43608 688688 47348 688698
rect 45338 688528 45618 688533
rect 45338 688268 45348 688528
rect 45608 688268 45618 688528
rect 45338 688263 45618 688268
rect 43608 688098 47348 688108
rect 43608 688088 45048 688098
rect 43608 687968 43628 688088
rect 43748 688028 45048 688088
rect 45118 688028 45368 688098
rect 45438 688028 45678 688098
rect 45748 688028 45998 688098
rect 46068 688088 47348 688098
rect 46068 688028 47208 688088
rect 43748 687968 47208 688028
rect 47328 687968 47348 688088
rect 18060 687920 43480 687960
rect 1640 685242 4522 687800
rect 18060 687760 18100 687920
rect 18240 687760 18440 687920
rect 18580 687760 18620 687920
rect 18760 687760 19000 687920
rect 19140 687760 43340 687920
rect 43460 687760 43480 687920
rect 18060 687720 43480 687760
rect 43608 687868 47348 687968
rect 43608 687748 43628 687868
rect 43748 687808 47208 687868
rect 43748 687748 45048 687808
rect 43608 687738 45048 687748
rect 45118 687738 45368 687808
rect 45438 687738 45678 687808
rect 45748 687738 45998 687808
rect 46068 687748 47208 687808
rect 47328 687748 47348 687868
rect 46068 687738 47348 687748
rect 43608 687728 47348 687738
rect 18060 687560 18100 687720
rect 18240 687560 18440 687720
rect 18580 687560 18620 687720
rect 18760 687560 19000 687720
rect 19140 687560 43340 687720
rect 43460 687560 43480 687720
rect 18060 687480 43480 687560
rect 44068 687538 46718 687548
rect 44068 687518 44888 687538
rect 44068 687448 44098 687518
rect 44168 687468 44888 687518
rect 44958 687468 45208 687538
rect 45278 687468 45528 687538
rect 45598 687468 45838 687538
rect 45908 687518 46718 687538
rect 45908 687468 46618 687518
rect 44168 687448 46618 687468
rect 46688 687448 46718 687518
rect 44068 687268 46718 687448
rect 44068 687198 44098 687268
rect 44168 687248 46618 687268
rect 44168 687198 44888 687248
rect 44068 687178 44888 687198
rect 44958 687178 45208 687248
rect 45278 687178 45528 687248
rect 45598 687178 45838 687248
rect 45908 687198 46618 687248
rect 46688 687198 46718 687268
rect 45908 687178 46718 687198
rect 44068 687168 46718 687178
rect 45338 687008 45618 687013
rect 45338 686748 45348 687008
rect 45608 686748 45618 687008
rect 45338 686743 45618 686748
rect 42398 686578 48538 686588
rect 42398 686568 43888 686578
rect 42398 686498 42428 686568
rect 42498 686508 43888 686568
rect 43958 686508 44408 686578
rect 44478 686508 44928 686578
rect 44998 686508 45438 686578
rect 45508 686508 45958 686578
rect 46028 686508 46468 686578
rect 46538 686508 46988 686578
rect 47058 686568 48538 686578
rect 47058 686508 48438 686568
rect 42498 686498 48438 686508
rect 48508 686498 48538 686568
rect 42398 686408 48538 686498
rect 42398 686338 42428 686408
rect 42498 686398 48438 686408
rect 42498 686338 43888 686398
rect 42398 686328 43888 686338
rect 43958 686328 44408 686398
rect 44478 686328 44928 686398
rect 44998 686328 45438 686398
rect 45508 686328 45958 686398
rect 46028 686328 46468 686398
rect 46538 686328 46988 686398
rect 47058 686338 48438 686398
rect 48508 686338 48538 686408
rect 47058 686328 48538 686338
rect 42398 686318 48538 686328
rect 43888 685908 47058 685918
rect 43888 685838 44148 685908
rect 44218 685838 44318 685908
rect 43888 685728 44318 685838
rect 43888 685658 44148 685728
rect 44218 685658 44318 685728
rect 44568 685838 44668 685908
rect 44738 685838 45178 685908
rect 45248 685838 45698 685908
rect 45768 685838 46218 685908
rect 46288 685838 46378 685908
rect 44568 685728 46378 685838
rect 44568 685658 44668 685728
rect 44738 685658 45178 685728
rect 45248 685658 45698 685728
rect 45768 685658 46218 685728
rect 46288 685658 46378 685728
rect 46628 685838 46728 685908
rect 46798 685838 47058 685908
rect 46628 685728 47058 685838
rect 46628 685658 46728 685728
rect 46798 685658 47058 685728
rect 43888 685648 47058 685658
rect -800 680242 4522 685242
rect 45338 685488 45608 685493
rect 45338 685238 45348 685488
rect 45598 685238 45608 685488
rect 45338 685233 45608 685238
rect 43638 685063 47318 685068
rect 43628 685058 47328 685063
rect 43628 684988 43638 685058
rect 43708 684988 44148 685058
rect 44218 684988 44668 685058
rect 44738 684988 45188 685058
rect 45258 684988 45698 685058
rect 45768 684988 46218 685058
rect 46288 684988 46728 685058
rect 46798 684988 47248 685058
rect 47318 684988 47328 685058
rect 43628 684983 47328 684988
rect 43638 684883 47318 684983
rect 43628 684878 47328 684883
rect 43628 684808 43638 684878
rect 43708 684808 44148 684878
rect 44218 684808 44668 684878
rect 44738 684808 45188 684878
rect 45258 684808 45698 684878
rect 45768 684808 46218 684878
rect 46288 684808 46728 684878
rect 46798 684808 47248 684878
rect 47318 684808 47328 684878
rect 43628 684803 47328 684808
rect 43638 684798 47318 684803
rect 43638 684388 47318 684398
rect 43638 684318 43898 684388
rect 43968 684318 44058 684388
rect 43638 684208 44058 684318
rect 43638 684138 43898 684208
rect 43968 684138 44058 684208
rect 44308 684318 44408 684388
rect 44478 684318 44928 684388
rect 44998 684318 45438 684388
rect 45508 684318 45958 684388
rect 46028 684318 46478 684388
rect 46548 684318 46638 684388
rect 44308 684208 46638 684318
rect 44308 684138 44408 684208
rect 44478 684138 44928 684208
rect 44998 684138 45438 684208
rect 45508 684138 45958 684208
rect 46028 684138 46478 684208
rect 46548 684138 46638 684208
rect 46888 684318 46988 684388
rect 47058 684318 47318 684388
rect 46888 684208 47318 684318
rect 46888 684138 46988 684208
rect 47058 684138 47318 684208
rect 43638 684128 47318 684138
rect 45338 683958 45608 683963
rect 45338 683708 45348 683958
rect 45598 683708 45608 683958
rect 45338 683703 45608 683708
rect 1642 680232 4522 680242
rect 9500 683380 11600 683400
rect 9500 683240 38760 683380
rect 9500 682240 9960 683240
rect 10960 683100 38760 683240
rect 10960 682240 38220 683100
rect 9500 682020 38220 682240
rect 9500 681020 9960 682020
rect 10960 681860 38220 682020
rect 38620 681860 38760 683100
rect 42268 683078 48728 683198
rect 42268 682918 42308 683078
rect 42468 682918 43308 683078
rect 43468 682918 44788 683078
rect 44948 682918 46008 683078
rect 46168 682918 47468 683078
rect 47628 682918 48528 683078
rect 48688 682918 48728 683078
rect 42268 682838 48728 682918
rect 42268 682538 42568 682838
rect 42868 682538 44068 682838
rect 44368 682538 46568 682838
rect 46868 682538 48168 682838
rect 48468 682538 48728 682838
rect 42268 682498 48728 682538
rect 42268 682338 42308 682498
rect 42468 682338 43308 682498
rect 43468 682338 44788 682498
rect 44948 682338 46008 682498
rect 46168 682338 47468 682498
rect 47628 682338 48528 682498
rect 48688 682338 48728 682498
rect 42268 682318 48728 682338
rect 10960 681020 38760 681860
rect 582300 681700 584800 682984
rect 9500 680840 38760 681020
rect 9500 679840 9960 680840
rect 10960 679840 38760 680840
rect 9500 679640 38760 679840
rect 42158 681118 48778 681158
rect 42158 680968 44598 681118
rect 44818 680968 46088 681118
rect 46308 680968 48778 681118
rect 42158 680938 48778 680968
rect 42158 680638 42368 680938
rect 42668 680638 43268 680938
rect 43568 680638 44168 680938
rect 44468 680638 46468 680938
rect 46768 680638 47368 680938
rect 47668 680638 48268 680938
rect 48568 680638 48778 680938
rect 42158 680568 48778 680638
rect 42158 680438 42368 680568
rect 42548 680438 43368 680568
rect 43548 680558 45158 680568
rect 43548 680438 44438 680558
rect 42158 680428 44438 680438
rect 44618 680438 45158 680558
rect 45338 680438 45598 680568
rect 45778 680438 46368 680568
rect 46548 680558 48778 680568
rect 46548 680438 47348 680558
rect 44618 680428 47348 680438
rect 47528 680428 48488 680558
rect 48668 680428 48778 680558
rect 42158 680398 48778 680428
rect 9500 679600 11600 679640
rect 42158 678658 42478 680398
rect 42158 678538 42218 678658
rect 42338 678538 42478 678658
rect 42158 675658 42478 678538
rect 42158 675538 42218 675658
rect 42338 675538 42478 675658
rect 42158 672658 42478 675538
rect 42158 672538 42218 672658
rect 42338 672538 42478 672658
rect 42158 669658 42478 672538
rect 42158 669538 42218 669658
rect 42338 669538 42478 669658
rect 42158 666658 42478 669538
rect 42158 666538 42218 666658
rect 42338 666538 42478 666658
rect 42158 665358 42478 666538
rect 48458 678658 48778 680398
rect 580590 679600 584800 681700
rect 48458 678538 48588 678658
rect 48708 678538 48778 678658
rect 48458 675658 48778 678538
rect 582300 677984 584800 679600
rect 48458 675538 48588 675658
rect 48708 675538 48778 675658
rect 48458 672658 48778 675538
rect 48458 672538 48588 672658
rect 48708 672538 48778 672658
rect 48458 669658 48778 672538
rect 48458 669538 48588 669658
rect 48708 669538 48778 669658
rect 48458 666658 48778 669538
rect 48458 666538 48588 666658
rect 48708 666538 48778 666658
rect 48458 665358 48778 666538
rect 42158 665338 48778 665358
rect 42158 664928 42608 665338
rect 43778 665328 48778 665338
rect 43778 664928 44128 665328
rect 42158 664918 44128 664928
rect 45298 664918 45648 665328
rect 46818 664918 47158 665328
rect 48328 664918 48778 665328
rect 42158 664878 48778 664918
rect 1800 648660 11600 648700
rect 460 648642 11600 648660
rect -800 648500 11600 648642
rect -800 648100 9700 648500
rect 10100 648100 10200 648500
rect 10600 648100 10700 648500
rect 11100 648100 11600 648500
rect -800 647700 11600 648100
rect -800 647660 10700 647700
rect -800 647260 9700 647660
rect 10100 647260 10180 647660
rect 10580 647300 10700 647660
rect 11100 647300 11600 647700
rect 10580 647260 11600 647300
rect -800 645240 11600 647260
rect -800 644840 9700 645240
rect 10100 644840 10200 645240
rect 10600 645200 11600 645240
rect 10600 644840 10700 645200
rect -800 644800 10700 644840
rect 11100 644800 11600 645200
rect -800 644400 11600 644800
rect -800 644000 9700 644400
rect 10100 644000 10200 644400
rect 10600 644000 10700 644400
rect 11100 644000 11600 644400
rect -800 643842 11600 644000
rect 460 643840 11600 643842
rect 1800 643800 11600 643840
rect 577414 644584 582400 644600
rect 577414 639800 584800 644584
rect 582340 639784 584800 639800
rect -800 638640 1660 638642
rect 1800 638640 11600 638700
rect -800 638500 11600 638640
rect -800 638100 9700 638500
rect 10100 638100 10200 638500
rect 10600 638100 10700 638500
rect 11100 638100 11600 638500
rect -800 637600 11600 638100
rect -800 637200 9700 637600
rect 10100 637200 10200 637600
rect 10600 637200 10700 637600
rect 11100 637200 11600 637600
rect -800 636700 11600 637200
rect -800 636300 9700 636700
rect 10100 636300 10200 636700
rect 10600 636300 10700 636700
rect 11100 636300 11600 636700
rect -800 636000 11600 636300
rect -800 635600 9700 636000
rect 10100 635600 10200 636000
rect 10600 635600 10700 636000
rect 11100 635600 11600 636000
rect -800 635300 11600 635600
rect -800 634900 9700 635300
rect 10100 634900 10200 635300
rect 10600 634900 10700 635300
rect 11100 634900 11600 635300
rect -800 634400 11600 634900
rect -800 634000 9700 634400
rect 10100 634000 10200 634400
rect 10600 634000 10700 634400
rect 11100 634000 11600 634400
rect -800 633842 11600 634000
rect 380 633820 11600 633842
rect 1800 633800 11600 633820
rect 577414 634584 582400 634600
rect 577414 629800 584800 634584
rect 582340 629784 584800 629800
rect 583520 589472 584800 589584
rect 583520 588290 584800 588402
rect 583520 587108 584800 587220
rect 583520 585926 584800 586038
rect 583520 584744 584800 584856
rect 583520 583562 584800 583674
rect 1180 564260 7080 564280
rect 34900 564260 41200 564300
rect 1180 564242 41200 564260
rect -800 563900 41200 564242
rect -800 562900 35400 563900
rect 36400 562900 36800 563900
rect 37800 562900 38200 563900
rect 39200 562900 39600 563900
rect 40600 562900 41200 563900
rect -800 562400 41200 562900
rect -800 561400 35400 562400
rect 36400 561400 36800 562400
rect 37800 561400 38200 562400
rect 39200 561400 39600 562400
rect 40600 561400 41200 562400
rect -800 560800 41200 561400
rect -800 559800 35400 560800
rect 36400 559800 36800 560800
rect 37800 559800 38200 560800
rect 39200 559800 39600 560800
rect 40600 559800 41200 560800
rect -800 559442 41200 559800
rect 1180 559440 41200 559442
rect 34900 559400 41200 559440
rect 34900 554280 41200 554300
rect 1380 554242 41200 554280
rect -800 553900 41200 554242
rect -800 552900 35400 553900
rect 36400 552900 36800 553900
rect 37800 552900 38200 553900
rect 39200 552900 39700 553900
rect 40700 552900 41200 553900
rect -800 552400 41200 552900
rect -800 551400 35400 552400
rect 36400 551400 36800 552400
rect 37800 551400 38200 552400
rect 39200 551400 39700 552400
rect 40700 551400 41200 552400
rect -800 550800 41200 551400
rect -800 549800 35400 550800
rect 36400 549800 36800 550800
rect 37800 549800 38200 550800
rect 39200 549800 39700 550800
rect 40700 549800 41200 550800
rect 582340 550562 584800 555362
rect -800 549442 41200 549800
rect 1380 549440 41200 549442
rect 6680 549420 41200 549440
rect 34900 549400 41200 549420
rect 582340 540562 584800 545362
rect -800 511530 480 511642
rect -800 510348 480 510460
rect -800 509166 480 509278
rect -800 507984 480 508096
rect -800 506802 480 506914
rect -800 505620 480 505732
rect 583520 500050 584800 500162
rect 583520 498868 584800 498980
rect 583520 497686 584800 497798
rect 583520 496504 584800 496616
rect 583520 495322 584800 495434
rect 583520 494140 584800 494252
rect -800 468308 480 468420
rect -800 467126 480 467238
rect -800 465944 480 466056
rect -800 464762 480 464874
rect -800 463580 480 463692
rect -800 462398 480 462510
rect 583520 455628 584800 455740
rect 583520 454446 584800 454558
rect 583520 453264 584800 453376
rect 583520 452082 584800 452194
rect 583520 450900 584800 451012
rect 583520 449718 584800 449830
rect -800 425086 480 425198
rect -800 423904 480 424016
rect -800 422722 480 422834
rect -800 421540 480 421652
rect -800 420358 480 420470
rect -800 419176 480 419288
rect 583520 411206 584800 411318
rect 583520 410024 584800 410136
rect 583520 408842 584800 408954
rect 583520 407660 584800 407772
rect 583520 406478 584800 406590
rect 583520 405296 584800 405408
rect -800 381864 480 381976
rect -800 380682 480 380794
rect -800 379500 480 379612
rect -800 378318 480 378430
rect -800 377136 480 377248
rect -800 375954 480 376066
rect 583520 364784 584800 364896
rect 583520 363602 584800 363714
rect 583520 362420 584800 362532
rect 583520 361238 584800 361350
rect 583520 360056 584800 360168
rect 583520 358874 584800 358986
rect -800 338642 480 338754
rect -800 337460 480 337572
rect -800 336278 480 336390
rect -800 335096 480 335208
rect -800 333914 480 334026
rect -800 332732 480 332844
rect 583520 319562 584800 319674
rect 583520 318380 584800 318492
rect 583520 317198 584800 317310
rect 583520 316016 584800 316128
rect 583520 314834 584800 314946
rect 583520 313652 584800 313764
rect -800 295420 480 295532
rect -800 294238 480 294350
rect -800 293056 480 293168
rect -800 291874 480 291986
rect -800 290692 480 290804
rect -800 289510 480 289622
rect 583520 275140 584800 275252
rect 583520 273958 584800 274070
rect 583520 272776 584800 272888
rect 583520 271594 584800 271706
rect 583520 270412 584800 270524
rect 583520 269230 584800 269342
rect -800 252398 480 252510
rect -800 251216 480 251328
rect -800 250034 480 250146
rect -800 248852 480 248964
rect -800 247670 480 247782
rect -800 246488 480 246600
rect 582340 235230 584800 240030
rect 582340 225230 584800 230030
rect -800 214888 1660 219688
rect -800 204888 1660 209688
rect 582340 191430 584800 196230
rect 582340 181430 584800 186230
rect -800 172888 1660 177688
rect -800 162888 1660 167688
rect 582340 146830 584800 151630
rect 582340 136830 584800 141630
rect -800 124776 480 124888
rect -800 123594 480 123706
rect -800 122412 480 122524
rect -800 121230 480 121342
rect -800 120048 480 120160
rect -800 118866 480 118978
rect 583520 95118 584800 95230
rect 583520 93936 584800 94048
rect 583520 92754 584800 92866
rect 583520 91572 584800 91684
rect -800 81554 480 81666
rect -800 80372 480 80484
rect -800 79190 480 79302
rect -800 78008 480 78120
rect -800 76826 480 76938
rect -800 75644 480 75756
rect 583520 50460 584800 50572
rect 583520 49278 584800 49390
rect 583520 48096 584800 48208
rect 583520 46914 584800 47026
rect -800 38332 480 38444
rect -800 37150 480 37262
rect -800 35968 480 36080
rect -800 34786 480 34898
rect -800 33604 480 33716
rect -800 32422 480 32534
rect 583520 24002 584800 24114
rect 583520 22820 584800 22932
rect 583520 21638 584800 21750
rect 583520 20456 584800 20568
rect 583520 19274 584800 19386
rect 583520 18092 584800 18204
rect -800 16910 480 17022
rect 583520 16910 584800 17022
rect -800 15728 480 15840
rect 583520 15728 584800 15840
rect -800 14546 480 14658
rect 583520 14546 584800 14658
rect -800 13364 480 13476
rect 583520 13364 584800 13476
rect -800 12182 480 12294
rect 583520 12182 584800 12294
rect -800 11000 480 11112
rect 583520 11000 584800 11112
rect -800 9818 480 9930
rect 583520 9818 584800 9930
rect -800 8636 480 8748
rect 583520 8636 584800 8748
rect -800 7454 480 7566
rect 583520 7454 584800 7566
rect -800 6272 480 6384
rect 583520 6272 584800 6384
rect -800 5090 480 5202
rect 583520 5090 584800 5202
rect -800 3908 480 4020
rect 583520 3908 584800 4020
rect -800 2726 480 2838
rect 583520 2726 584800 2838
rect -800 1544 480 1656
rect 583520 1544 584800 1656
<< via3 >>
rect 18100 702740 18340 703000
rect 18520 702740 18760 703000
rect 18940 702740 19180 703000
rect 18100 702340 18340 702600
rect 18520 702340 18760 702600
rect 18940 702340 19180 702600
rect 70220 702660 70440 702880
rect 70640 702660 70860 702880
rect 71080 702660 71300 702880
rect 70220 702340 70440 702560
rect 70640 702340 70860 702560
rect 71080 702340 71300 702560
rect 38106 700283 41450 700347
rect 41906 700283 45250 700347
rect 45706 700283 49050 700347
rect 49506 700283 52850 700347
rect 41600 696200 41800 696380
rect 49180 696180 49380 696360
rect 41600 695720 41800 695900
rect 49180 695740 49380 695920
rect 44798 694608 45068 694878
rect 45848 694608 46118 694878
rect 37738 694088 37808 694158
rect 42658 694118 42908 694368
rect 44558 694118 44808 694368
rect 46138 694118 46388 694368
rect 48038 694328 48278 694378
rect 48278 694328 48288 694378
rect 48038 694158 48288 694328
rect 48038 694128 48278 694158
rect 48278 694128 48288 694158
rect 53128 694088 53198 694158
rect 37628 693978 37698 694048
rect 53238 693978 53308 694048
rect 41528 693098 41618 693198
rect 41718 693098 41808 693198
rect 44798 692968 45068 693238
rect 45848 692968 46118 693238
rect 49138 693098 49228 693198
rect 49328 693098 49418 693198
rect 39578 692598 39758 692698
rect 39998 692598 40178 692698
rect 43998 692658 44008 692718
rect 44008 692658 44248 692718
rect 44248 692658 44258 692718
rect 45258 692658 45268 692718
rect 45268 692658 45518 692718
rect 46528 692658 46538 692718
rect 46538 692658 46778 692718
rect 46778 692658 46788 692718
rect 43998 692518 44258 692658
rect 45258 692518 45518 692658
rect 46528 692518 46788 692658
rect 50828 692598 51008 692698
rect 51248 692598 51428 692698
rect 43998 692458 44008 692518
rect 44008 692458 44248 692518
rect 44248 692458 44258 692518
rect 45258 692458 45268 692518
rect 45268 692458 45518 692518
rect 46528 692458 46538 692518
rect 46538 692458 46778 692518
rect 46778 692458 46788 692518
rect 44588 691368 44848 691628
rect 46088 691368 46348 691628
rect 43998 691108 44008 691168
rect 44008 691108 44248 691168
rect 44248 691108 44258 691168
rect 45258 691108 45268 691168
rect 45268 691108 45518 691168
rect 46528 691108 46538 691168
rect 46538 691108 46778 691168
rect 46778 691108 46788 691168
rect 43998 690968 44258 691108
rect 45258 690968 45518 691108
rect 46528 690968 46788 691108
rect 43998 690908 44008 690968
rect 44008 690908 44248 690968
rect 44248 690908 44258 690968
rect 45258 690908 45268 690968
rect 45268 690908 45518 690968
rect 46528 690908 46538 690968
rect 46538 690908 46778 690968
rect 46778 690908 46788 690968
rect 70240 689320 70460 689540
rect 70640 689320 70860 689540
rect 71060 689320 71280 689540
rect 70240 689060 70460 689280
rect 70640 689060 70860 689280
rect 71060 689060 71280 689280
rect 45348 688268 45608 688528
rect 18100 687760 18240 687920
rect 18440 687760 18580 687920
rect 18620 687760 18760 687920
rect 19000 687760 19140 687920
rect 18100 687560 18240 687720
rect 18440 687560 18580 687720
rect 18620 687560 18760 687720
rect 19000 687560 19140 687720
rect 45348 686748 45608 687008
rect 44318 685658 44568 685908
rect 46378 685658 46628 685908
rect 45348 685238 45598 685488
rect 44058 684138 44308 684388
rect 46638 684138 46888 684388
rect 45348 683708 45598 683958
rect 9960 682240 10960 683240
rect 9960 681020 10960 682020
rect 38220 681860 38620 683100
rect 42568 682538 42868 682838
rect 44068 682538 44368 682838
rect 46568 682538 46868 682838
rect 48168 682538 48468 682838
rect 9960 679840 10960 680840
rect 42368 680638 42668 680938
rect 43268 680638 43568 680938
rect 44168 680638 44468 680938
rect 46468 680638 46768 680938
rect 47368 680638 47668 680938
rect 48268 680638 48568 680938
rect 9700 648100 10100 648500
rect 10200 648100 10600 648500
rect 10700 648100 11100 648500
rect 9700 647260 10100 647660
rect 10180 647260 10580 647660
rect 10700 647300 11100 647700
rect 9700 644840 10100 645240
rect 10200 644840 10600 645240
rect 10700 644800 11100 645200
rect 9700 644000 10100 644400
rect 10200 644000 10600 644400
rect 10700 644000 11100 644400
rect 9700 638100 10100 638500
rect 10200 638100 10600 638500
rect 10700 638100 11100 638500
rect 9700 637200 10100 637600
rect 10200 637200 10600 637600
rect 10700 637200 11100 637600
rect 9700 636300 10100 636700
rect 10200 636300 10600 636700
rect 10700 636300 11100 636700
rect 9700 635600 10100 636000
rect 10200 635600 10600 636000
rect 10700 635600 11100 636000
rect 9700 634900 10100 635300
rect 10200 634900 10600 635300
rect 10700 634900 11100 635300
rect 9700 634000 10100 634400
rect 10200 634000 10600 634400
rect 10700 634000 11100 634400
rect 35400 562900 36400 563900
rect 36800 562900 37800 563900
rect 38200 562900 39200 563900
rect 39600 562900 40600 563900
rect 35400 561400 36400 562400
rect 36800 561400 37800 562400
rect 38200 561400 39200 562400
rect 39600 561400 40600 562400
rect 35400 559800 36400 560800
rect 36800 559800 37800 560800
rect 38200 559800 39200 560800
rect 39600 559800 40600 560800
rect 35400 552900 36400 553900
rect 36800 552900 37800 553900
rect 38200 552900 39200 553900
rect 39700 552900 40700 553900
rect 35400 551400 36400 552400
rect 36800 551400 37800 552400
rect 38200 551400 39200 552400
rect 39700 551400 40700 552400
rect 35400 549800 36400 550800
rect 36800 549800 37800 550800
rect 38200 549800 39200 550800
rect 39700 549800 40700 550800
<< mimcap >>
rect 38178 700128 41378 700168
rect 38178 697008 38218 700128
rect 41338 697008 41378 700128
rect 38178 696968 41378 697008
rect 41978 700128 45178 700168
rect 41978 697008 42018 700128
rect 45138 697008 45178 700128
rect 41978 696968 45178 697008
rect 45778 700128 48978 700168
rect 45778 697008 45818 700128
rect 48938 697008 48978 700128
rect 45778 696968 48978 697008
rect 49578 700128 52778 700168
rect 49578 697008 49618 700128
rect 52738 697008 52778 700128
rect 49578 696968 52778 697008
<< mimcapcontact >>
rect 38218 697008 41338 700128
rect 42018 697008 45138 700128
rect 45818 697008 48938 700128
rect 49618 697008 52738 700128
<< metal4 >>
rect 17780 703000 19500 703040
rect 17780 702740 18100 703000
rect 18340 702740 18520 703000
rect 18760 702740 18940 703000
rect 19180 702740 19500 703000
rect 17780 702600 19500 702740
rect 17780 702340 18100 702600
rect 18340 702340 18520 702600
rect 18760 702340 18940 702600
rect 19180 702340 19500 702600
rect 17780 702300 19500 702340
rect 69940 702880 71660 702920
rect 69940 702660 70220 702880
rect 70440 702660 70640 702880
rect 70860 702660 71080 702880
rect 71300 702660 71660 702880
rect 69940 702560 71660 702660
rect 69940 702340 70220 702560
rect 70440 702340 70640 702560
rect 70860 702340 71080 702560
rect 71300 702340 71660 702560
rect 69940 702300 71660 702340
rect 165594 702300 170594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 329294 702300 334294 704800
rect 18060 687920 19220 702300
rect 37608 700347 53328 700498
rect 37608 700283 38106 700347
rect 41450 700283 41906 700347
rect 45250 700283 45706 700347
rect 49050 700283 49506 700347
rect 52850 700283 53328 700347
rect 37608 700258 53328 700283
rect 37608 694158 37828 700258
rect 38217 700128 41339 700129
rect 38217 697008 38218 700128
rect 41338 698788 41339 700128
rect 42017 700128 45139 700129
rect 42017 698788 42018 700128
rect 41338 698428 42018 698788
rect 41338 697008 41339 698428
rect 38217 697007 41339 697008
rect 37608 694088 37738 694158
rect 37808 694088 37828 694158
rect 37608 694048 37828 694088
rect 37608 693978 37628 694048
rect 37698 693978 37828 694048
rect 37608 693958 37828 693978
rect 41508 696380 41828 698428
rect 42017 697008 42018 698428
rect 45138 698788 45139 700128
rect 45817 700128 48939 700129
rect 45817 698788 45818 700128
rect 45138 698428 45818 698788
rect 45138 697008 45139 698428
rect 42017 697007 45139 697008
rect 45817 697008 45818 698428
rect 48938 698788 48939 700128
rect 49617 700128 52739 700129
rect 49617 698788 49618 700128
rect 48938 698428 49618 698788
rect 48938 697008 48939 698428
rect 45817 697007 48939 697008
rect 41508 696200 41600 696380
rect 41800 696200 41828 696380
rect 41508 695900 41828 696200
rect 41508 695720 41600 695900
rect 41800 695720 41828 695900
rect 41508 693198 41828 695720
rect 49118 696360 49438 698428
rect 49617 697008 49618 698428
rect 52738 697008 52739 700128
rect 49617 697007 52739 697008
rect 49118 696180 49180 696360
rect 49380 696180 49438 696360
rect 49118 695920 49438 696180
rect 49118 695740 49180 695920
rect 49380 695740 49438 695920
rect 44797 694878 45069 694879
rect 44797 694608 44798 694878
rect 45068 694608 45069 694878
rect 44797 694607 45069 694608
rect 45847 694878 46119 694879
rect 45847 694608 45848 694878
rect 46118 694608 46119 694878
rect 45847 694607 46119 694608
rect 48037 694378 48289 694379
rect 42657 694368 42909 694369
rect 42657 694118 42658 694368
rect 42908 694118 42909 694368
rect 42657 694117 42909 694118
rect 44557 694368 44809 694369
rect 44557 694118 44558 694368
rect 44808 694118 44809 694368
rect 44557 694117 44809 694118
rect 46137 694368 46389 694369
rect 46137 694118 46138 694368
rect 46388 694118 46389 694368
rect 48037 694128 48038 694378
rect 48288 694128 48289 694378
rect 48037 694127 48289 694128
rect 46137 694117 46389 694118
rect 41508 693098 41528 693198
rect 41618 693098 41718 693198
rect 41808 693098 41828 693198
rect 41508 693078 41828 693098
rect 44797 693238 45069 693239
rect 44797 692968 44798 693238
rect 45068 692968 45069 693238
rect 44797 692967 45069 692968
rect 45847 693238 46119 693239
rect 45847 692968 45848 693238
rect 46118 692968 46119 693238
rect 49118 693198 49438 695740
rect 53108 694158 53328 700258
rect 53108 694088 53128 694158
rect 53198 694088 53328 694158
rect 53108 694048 53328 694088
rect 53108 693978 53238 694048
rect 53308 693978 53328 694048
rect 53108 693958 53328 693978
rect 49118 693098 49138 693198
rect 49228 693098 49328 693198
rect 49418 693098 49438 693198
rect 49118 693078 49438 693098
rect 45847 692967 46119 692968
rect 39548 692700 40208 692728
rect 43997 692718 44259 692719
rect 39500 692698 40400 692700
rect 39500 692598 39578 692698
rect 39758 692598 39998 692698
rect 40178 692598 40400 692698
rect 18060 687760 18100 687920
rect 18240 687760 18440 687920
rect 18580 687760 18620 687920
rect 18760 687760 19000 687920
rect 19140 687760 19220 687920
rect 18060 687720 19220 687760
rect 18060 687560 18100 687720
rect 18240 687560 18440 687720
rect 18580 687560 18620 687720
rect 18760 687560 19000 687720
rect 19140 687560 19220 687720
rect 18060 687520 19220 687560
rect 38088 691778 38758 691808
rect 38088 691538 38118 691778
rect 38358 691538 38488 691778
rect 38728 691538 38758 691778
rect 38088 691108 38758 691538
rect 38088 690868 38118 691108
rect 38358 690868 38488 691108
rect 38728 690868 38758 691108
rect 8500 683240 12600 683500
rect 8500 682240 9960 683240
rect 10960 682240 12600 683240
rect 8500 682020 12600 682240
rect 8500 681020 9960 682020
rect 10960 681020 12600 682020
rect 38088 683208 38758 690868
rect 38088 682968 38118 683208
rect 38358 683100 38488 683208
rect 38728 682968 38758 683208
rect 38088 682008 38220 682968
rect 38620 682008 38758 682968
rect 38088 681768 38118 682008
rect 38358 681768 38488 681860
rect 38728 681768 38758 682008
rect 38088 681738 38758 681768
rect 39500 685258 40400 692598
rect 43997 692458 43998 692718
rect 44258 692458 44259 692718
rect 43997 692457 44259 692458
rect 45257 692718 45519 692719
rect 45257 692458 45258 692718
rect 45518 692458 45519 692718
rect 45257 692457 45519 692458
rect 46527 692718 46789 692719
rect 46527 692458 46528 692718
rect 46788 692458 46789 692718
rect 46527 692457 46789 692458
rect 50798 692698 51458 692728
rect 50798 692598 50828 692698
rect 51008 692598 51248 692698
rect 51428 692598 51458 692698
rect 44587 691628 44849 691629
rect 44587 691368 44588 691628
rect 44848 691368 44849 691628
rect 44587 691367 44849 691368
rect 46087 691628 46349 691629
rect 46087 691368 46088 691628
rect 46348 691368 46349 691628
rect 46087 691367 46349 691368
rect 43997 691168 44259 691169
rect 43997 690908 43998 691168
rect 44258 690908 44259 691168
rect 43997 690907 44259 690908
rect 45257 691168 45519 691169
rect 45257 690908 45258 691168
rect 45518 690908 45519 691168
rect 45257 690907 45519 690908
rect 46527 691168 46789 691169
rect 46527 690908 46528 691168
rect 46788 690908 46789 691168
rect 46527 690907 46789 690908
rect 45347 688528 45609 688529
rect 45347 688268 45348 688528
rect 45608 688268 45609 688528
rect 45347 688267 45609 688268
rect 45347 687008 45609 687009
rect 45347 686748 45348 687008
rect 45608 686748 45609 687008
rect 45347 686747 45609 686748
rect 44317 685908 44569 685909
rect 44317 685658 44318 685908
rect 44568 685658 44569 685908
rect 44317 685657 44569 685658
rect 46377 685908 46629 685909
rect 46377 685658 46378 685908
rect 46628 685658 46629 685908
rect 46377 685657 46629 685658
rect 39500 685018 39578 685258
rect 39818 685018 39938 685258
rect 40178 685018 40400 685258
rect 45347 685488 45599 685489
rect 45347 685238 45348 685488
rect 45598 685238 45599 685488
rect 45347 685237 45599 685238
rect 50798 685258 51458 692598
rect 39500 684918 40400 685018
rect 39500 684678 39578 684918
rect 39818 684678 39938 684918
rect 40178 684678 40400 684918
rect 8500 680840 12600 681020
rect 8500 679840 9960 680840
rect 10960 679840 12600 680840
rect 39500 681108 40400 684678
rect 50798 685018 50828 685258
rect 51068 685018 51188 685258
rect 51428 685018 51458 685258
rect 50798 684918 51458 685018
rect 50798 684678 50828 684918
rect 51068 684678 51188 684918
rect 51428 684678 51458 684918
rect 44057 684388 44309 684389
rect 44057 684138 44058 684388
rect 44308 684138 44309 684388
rect 44057 684137 44309 684138
rect 46637 684388 46889 684389
rect 46637 684138 46638 684388
rect 46888 684138 46889 684388
rect 46637 684137 46889 684138
rect 45347 683958 45599 683959
rect 45347 683708 45348 683958
rect 45598 683708 45599 683958
rect 45347 683707 45599 683708
rect 42567 682838 42869 682839
rect 42567 682538 42568 682838
rect 42868 682538 42869 682838
rect 42567 682537 42869 682538
rect 44067 682838 44369 682839
rect 44067 682538 44068 682838
rect 44368 682538 44369 682838
rect 44067 682537 44369 682538
rect 46567 682838 46869 682839
rect 46567 682538 46568 682838
rect 46868 682538 46869 682838
rect 46567 682537 46869 682538
rect 48167 682838 48469 682839
rect 48167 682538 48168 682838
rect 48468 682538 48469 682838
rect 48167 682537 48469 682538
rect 39500 680868 39578 681108
rect 39818 680868 39938 681108
rect 40178 680868 40400 681108
rect 50798 681108 51458 684678
rect 52248 691678 52918 691708
rect 52248 691438 52278 691678
rect 52518 691438 52648 691678
rect 52888 691438 52918 691678
rect 52248 691108 52918 691438
rect 52248 690868 52278 691108
rect 52518 690868 52648 691108
rect 52888 690868 52918 691108
rect 52248 683208 52918 690868
rect 70180 689540 71340 702300
rect 70180 689320 70240 689540
rect 70460 689320 70640 689540
rect 70860 689320 71060 689540
rect 71280 689320 71340 689540
rect 70180 689280 71340 689320
rect 70180 689060 70240 689280
rect 70460 689060 70640 689280
rect 70860 689060 71060 689280
rect 71280 689060 71340 689280
rect 70180 689020 71340 689060
rect 52248 682968 52278 683208
rect 52518 682968 52648 683208
rect 52888 682968 52918 683208
rect 52248 682008 52918 682968
rect 52248 681768 52278 682008
rect 52518 681768 52648 682008
rect 52888 681768 52918 682008
rect 52248 681738 52918 681768
rect 39500 679840 40400 680868
rect 42367 680938 42669 680939
rect 42367 680638 42368 680938
rect 42668 680638 42669 680938
rect 42367 680637 42669 680638
rect 43267 680938 43569 680939
rect 43267 680638 43268 680938
rect 43568 680638 43569 680938
rect 43267 680637 43569 680638
rect 44167 680938 44469 680939
rect 44167 680638 44168 680938
rect 44468 680638 44469 680938
rect 44167 680637 44469 680638
rect 46467 680938 46769 680939
rect 46467 680638 46468 680938
rect 46768 680638 46769 680938
rect 46467 680637 46769 680638
rect 47367 680938 47669 680939
rect 47367 680638 47368 680938
rect 47668 680638 47669 680938
rect 47367 680637 47669 680638
rect 48267 680938 48569 680939
rect 48267 680638 48268 680938
rect 48568 680638 48569 680938
rect 48267 680637 48569 680638
rect 50798 680868 50828 681108
rect 51068 680868 51188 681108
rect 51428 680868 51458 681108
rect 8500 648500 12600 679840
rect 8500 648100 9700 648500
rect 10100 648100 10200 648500
rect 10600 648100 10700 648500
rect 11100 648100 12600 648500
rect 8500 647700 12600 648100
rect 8500 647660 10700 647700
rect 8500 647260 9700 647660
rect 10100 647260 10180 647660
rect 10580 647300 10700 647660
rect 11100 647300 12600 647700
rect 10580 647260 12600 647300
rect 8500 645240 12600 647260
rect 8500 644840 9700 645240
rect 10100 644840 10200 645240
rect 10600 645200 12600 645240
rect 10600 644840 10700 645200
rect 8500 644800 10700 644840
rect 11100 644800 12600 645200
rect 8500 644400 12600 644800
rect 8500 644000 9700 644400
rect 10100 644000 10200 644400
rect 10600 644000 10700 644400
rect 11100 644000 12600 644400
rect 8500 638500 12600 644000
rect 8500 638100 9700 638500
rect 10100 638100 10200 638500
rect 10600 638100 10700 638500
rect 11100 638100 12600 638500
rect 8500 637600 12600 638100
rect 8500 637200 9700 637600
rect 10100 637200 10200 637600
rect 10600 637200 10700 637600
rect 11100 637200 12600 637600
rect 8500 636700 12600 637200
rect 8500 636300 9700 636700
rect 10100 636300 10200 636700
rect 10600 636300 10700 636700
rect 11100 636300 12600 636700
rect 8500 636000 12600 636300
rect 8500 635600 9700 636000
rect 10100 635600 10200 636000
rect 10600 635600 10700 636000
rect 11100 635600 12600 636000
rect 8500 635300 12600 635600
rect 8500 634900 9700 635300
rect 10100 634900 10200 635300
rect 10600 634900 10700 635300
rect 11100 634900 12600 635300
rect 8500 634400 12600 634900
rect 8500 634000 9700 634400
rect 10100 634000 10200 634400
rect 10600 634000 10700 634400
rect 11100 634000 12600 634400
rect 8500 633800 12600 634000
rect 34940 679808 41060 679840
rect 34940 679568 39578 679808
rect 39818 679568 39938 679808
rect 40178 679568 41060 679808
rect 34940 565100 41060 679568
rect 50798 679808 51458 680868
rect 50798 679568 50828 679808
rect 51068 679568 51188 679808
rect 51428 679568 51458 679808
rect 50798 679538 51458 679568
rect 34940 564300 41100 565100
rect 35000 563900 41100 564300
rect 35000 562900 35400 563900
rect 36400 562900 36800 563900
rect 37800 562900 38200 563900
rect 39200 562900 39600 563900
rect 40600 562900 41100 563900
rect 35000 562400 41100 562900
rect 35000 561400 35400 562400
rect 36400 561400 36800 562400
rect 37800 561400 38200 562400
rect 39200 561400 39600 562400
rect 40600 561400 41100 562400
rect 35000 560800 41100 561400
rect 35000 559800 35400 560800
rect 36400 559800 36800 560800
rect 37800 559800 38200 560800
rect 39200 559800 39600 560800
rect 40600 559800 41100 560800
rect 35000 553900 41100 559800
rect 35000 552900 35400 553900
rect 36400 552900 36800 553900
rect 37800 552900 38200 553900
rect 39200 552900 39700 553900
rect 40700 552900 41100 553900
rect 35000 552400 41100 552900
rect 35000 551400 35400 552400
rect 36400 551400 36800 552400
rect 37800 551400 38200 552400
rect 39200 551400 39700 552400
rect 40700 551400 41100 552400
rect 35000 550800 41100 551400
rect 35000 549800 35400 550800
rect 36400 549800 36800 550800
rect 37800 549800 38200 550800
rect 39200 549800 39700 550800
rect 40700 549800 41100 550800
rect 35000 549400 41100 549800
<< via4 >>
rect 44798 694608 45068 694878
rect 45848 694608 46118 694878
rect 42658 694118 42908 694368
rect 44558 694118 44808 694368
rect 46138 694118 46388 694368
rect 48038 694128 48288 694378
rect 44798 692968 45068 693238
rect 45848 692968 46118 693238
rect 38118 691538 38358 691778
rect 38488 691538 38728 691778
rect 38118 690868 38358 691108
rect 38488 690868 38728 691108
rect 38118 683100 38358 683208
rect 38488 683100 38728 683208
rect 38118 682968 38220 683100
rect 38220 682968 38358 683100
rect 38488 682968 38620 683100
rect 38620 682968 38728 683100
rect 38118 681860 38220 682008
rect 38220 681860 38358 682008
rect 38488 681860 38620 682008
rect 38620 681860 38728 682008
rect 38118 681768 38358 681860
rect 38488 681768 38728 681860
rect 43998 692458 44258 692718
rect 45258 692458 45518 692718
rect 46528 692458 46788 692718
rect 44588 691368 44848 691628
rect 46088 691368 46348 691628
rect 43998 690908 44258 691168
rect 45258 690908 45518 691168
rect 46528 690908 46788 691168
rect 45348 688268 45608 688528
rect 45348 686748 45608 687008
rect 44318 685658 44568 685908
rect 46378 685658 46628 685908
rect 39578 685018 39818 685258
rect 39938 685018 40178 685258
rect 45348 685238 45598 685488
rect 39578 684678 39818 684918
rect 39938 684678 40178 684918
rect 50828 685018 51068 685258
rect 51188 685018 51428 685258
rect 50828 684678 51068 684918
rect 51188 684678 51428 684918
rect 44058 684138 44308 684388
rect 46638 684138 46888 684388
rect 45348 683708 45598 683958
rect 42568 682538 42868 682838
rect 44068 682538 44368 682838
rect 46568 682538 46868 682838
rect 48168 682538 48468 682838
rect 39578 680868 39818 681108
rect 39938 680868 40178 681108
rect 52278 691438 52518 691678
rect 52648 691438 52888 691678
rect 52278 690868 52518 691108
rect 52648 690868 52888 691108
rect 52278 682968 52518 683208
rect 52648 682968 52888 683208
rect 52278 681768 52518 682008
rect 52648 681768 52888 682008
rect 42368 680638 42668 680938
rect 43268 680638 43568 680938
rect 44168 680638 44468 680938
rect 46468 680638 46768 680938
rect 47368 680638 47668 680938
rect 48268 680638 48568 680938
rect 50828 680868 51068 681108
rect 51188 680868 51428 681108
rect 39578 679568 39818 679808
rect 39938 679568 40178 679808
rect 50828 679568 51068 679808
rect 51188 679568 51428 679808
<< metal5 >>
rect 165594 702300 170594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 329294 702300 334294 704800
rect 36568 694878 53768 694938
rect 36568 694608 44798 694878
rect 45068 694608 45848 694878
rect 46118 694608 53768 694878
rect 36568 694378 53768 694608
rect 36568 694368 48038 694378
rect 36568 694118 42658 694368
rect 42908 694118 44558 694368
rect 44808 694118 46138 694368
rect 46388 694128 48038 694368
rect 48288 694128 53768 694378
rect 46388 694118 53768 694128
rect 36568 693238 53768 694118
rect 36568 692968 44798 693238
rect 45068 692968 45848 693238
rect 46118 692968 53768 693238
rect 36568 692718 53768 692968
rect 36568 692458 43998 692718
rect 44258 692458 45258 692718
rect 45518 692458 46528 692718
rect 46788 692458 53768 692718
rect 36568 691778 53768 692458
rect 36568 691538 38118 691778
rect 38358 691538 38488 691778
rect 38728 691678 53768 691778
rect 38728 691628 52278 691678
rect 38728 691538 44588 691628
rect 36568 691368 44588 691538
rect 44848 691368 46088 691628
rect 46348 691438 52278 691628
rect 52518 691438 52648 691678
rect 52888 691438 53768 691678
rect 46348 691368 53768 691438
rect 36568 691168 53768 691368
rect 36568 691108 43998 691168
rect 36568 690868 38118 691108
rect 38358 690868 38488 691108
rect 38728 690908 43998 691108
rect 44258 690908 45258 691168
rect 45518 690908 46528 691168
rect 46788 691108 53768 691168
rect 46788 690908 52278 691108
rect 38728 690868 52278 690908
rect 52518 690868 52648 691108
rect 52888 690868 53768 691108
rect 36568 690838 53768 690868
rect 45258 688528 45698 688568
rect 45258 688268 45348 688528
rect 45608 688268 45698 688528
rect 45258 687008 45698 688268
rect 45258 686748 45348 687008
rect 45608 686748 45698 687008
rect 45258 685958 45698 686748
rect 38088 685908 53168 685958
rect 38088 685658 44318 685908
rect 44568 685658 46378 685908
rect 46628 685658 53168 685908
rect 38088 685488 53168 685658
rect 38088 685258 45348 685488
rect 38088 685018 39578 685258
rect 39818 685018 39938 685258
rect 40178 685238 45348 685258
rect 45598 685258 53168 685488
rect 45598 685238 50828 685258
rect 40178 685018 50828 685238
rect 51068 685018 51188 685258
rect 51428 685018 53168 685258
rect 38088 684918 53168 685018
rect 38088 684678 39578 684918
rect 39818 684678 39938 684918
rect 40178 684678 50828 684918
rect 51068 684678 51188 684918
rect 51428 684678 53168 684918
rect 38088 684388 53168 684678
rect 38088 684138 44058 684388
rect 44308 684138 46638 684388
rect 46888 684138 53168 684388
rect 38088 684098 53168 684138
rect 45248 683958 45688 684098
rect 45248 683708 45348 683958
rect 45598 683708 45688 683958
rect 45248 683638 45688 683708
rect 38088 683208 53168 683238
rect 38088 682968 38118 683208
rect 38358 682968 38488 683208
rect 38728 682968 52278 683208
rect 52518 682968 52648 683208
rect 52888 682968 53168 683208
rect 38088 682838 53168 682968
rect 38088 682538 42568 682838
rect 42868 682538 44068 682838
rect 44368 682538 46568 682838
rect 46868 682538 48168 682838
rect 48468 682538 53168 682838
rect 38088 682008 53168 682538
rect 38088 681768 38118 682008
rect 38358 681768 38488 682008
rect 38728 681768 52278 682008
rect 52518 681768 52648 682008
rect 52888 681768 53168 682008
rect 38088 681738 53168 681768
rect 38088 681108 53168 681138
rect 38088 680868 39578 681108
rect 39818 680868 39938 681108
rect 40178 680938 50828 681108
rect 40178 680868 42368 680938
rect 38088 680638 42368 680868
rect 42668 680638 43268 680938
rect 43568 680638 44168 680938
rect 44468 680638 46468 680938
rect 46768 680638 47368 680938
rect 47668 680638 48268 680938
rect 48568 680868 50828 680938
rect 51068 680868 51188 681108
rect 51428 680868 53168 681108
rect 48568 680638 53168 680868
rect 38088 679808 53168 680638
rect 38088 679568 39578 679808
rect 39818 679568 39938 679808
rect 40178 679568 50828 679808
rect 51068 679568 51188 679808
rect 51428 679568 53168 679808
rect 38088 679538 53168 679568
<< comment >>
rect -100 704000 584100 704100
rect -100 0 0 704000
rect 584000 0 584100 704000
rect -100 -100 584100 0
<< res5p73 >>
rect 38931 694219 40935 695369
rect 50001 694219 52005 695369
rect 38931 692759 40935 693909
rect 50001 692759 52005 693909
rect 42623 665374 43773 679178
rect 44133 665374 45283 679178
rect 45643 665368 46793 679172
rect 47163 665368 48313 679172
<< labels >>
flabel metal3 s 583520 269230 584800 269342 0 FreeSans 1120 0 0 0 gpio_analog[0]
port 624 nsew signal bidirectional
flabel metal3 s -800 381864 480 381976 0 FreeSans 1120 0 0 0 gpio_analog[10]
port 614 nsew signal bidirectional
flabel metal3 s -800 338642 480 338754 0 FreeSans 1120 0 0 0 gpio_analog[11]
port 613 nsew signal bidirectional
flabel metal3 s -800 295420 480 295532 0 FreeSans 1120 0 0 0 gpio_analog[12]
port 612 nsew signal bidirectional
flabel metal3 s -800 252398 480 252510 0 FreeSans 1120 0 0 0 gpio_analog[13]
port 611 nsew signal bidirectional
flabel metal3 s -800 124776 480 124888 0 FreeSans 1120 0 0 0 gpio_analog[14]
port 610 nsew signal bidirectional
flabel metal3 s -800 81554 480 81666 0 FreeSans 1120 0 0 0 gpio_analog[15]
port 609 nsew signal bidirectional
flabel metal3 s -800 38332 480 38444 0 FreeSans 1120 0 0 0 gpio_analog[16]
port 608 nsew signal bidirectional
flabel metal3 s -800 16910 480 17022 0 FreeSans 1120 0 0 0 gpio_analog[17]
port 607 nsew signal bidirectional
flabel metal3 s 583520 313652 584800 313764 0 FreeSans 1120 0 0 0 gpio_analog[1]
port 623 nsew signal bidirectional
flabel metal3 s 583520 358874 584800 358986 0 FreeSans 1120 0 0 0 gpio_analog[2]
port 622 nsew signal bidirectional
flabel metal3 s 583520 405296 584800 405408 0 FreeSans 1120 0 0 0 gpio_analog[3]
port 621 nsew signal bidirectional
flabel metal3 s 583520 449718 584800 449830 0 FreeSans 1120 0 0 0 gpio_analog[4]
port 620 nsew signal bidirectional
flabel metal3 s 583520 494140 584800 494252 0 FreeSans 1120 0 0 0 gpio_analog[5]
port 619 nsew signal bidirectional
flabel metal3 s 583520 583562 584800 583674 0 FreeSans 1120 0 0 0 gpio_analog[6]
port 618 nsew signal bidirectional
flabel metal3 s -800 468308 480 468420 0 FreeSans 1120 0 0 0 gpio_analog[8]
port 616 nsew signal bidirectional
flabel metal3 s -800 425086 480 425198 0 FreeSans 1120 0 0 0 gpio_analog[9]
port 615 nsew signal bidirectional
flabel metal3 s 583520 270412 584800 270524 0 FreeSans 1120 0 0 0 gpio_noesd[0]
port 642 nsew signal bidirectional
flabel metal3 s -800 380682 480 380794 0 FreeSans 1120 0 0 0 gpio_noesd[10]
port 632 nsew signal bidirectional
flabel metal3 s -800 337460 480 337572 0 FreeSans 1120 0 0 0 gpio_noesd[11]
port 631 nsew signal bidirectional
flabel metal3 s -800 294238 480 294350 0 FreeSans 1120 0 0 0 gpio_noesd[12]
port 630 nsew signal bidirectional
flabel metal3 s -800 251216 480 251328 0 FreeSans 1120 0 0 0 gpio_noesd[13]
port 629 nsew signal bidirectional
flabel metal3 s -800 123594 480 123706 0 FreeSans 1120 0 0 0 gpio_noesd[14]
port 628 nsew signal bidirectional
flabel metal3 s -800 80372 480 80484 0 FreeSans 1120 0 0 0 gpio_noesd[15]
port 627 nsew signal bidirectional
flabel metal3 s -800 37150 480 37262 0 FreeSans 1120 0 0 0 gpio_noesd[16]
port 626 nsew signal bidirectional
flabel metal3 s -800 15728 480 15840 0 FreeSans 1120 0 0 0 gpio_noesd[17]
port 625 nsew signal bidirectional
flabel metal3 s 583520 314834 584800 314946 0 FreeSans 1120 0 0 0 gpio_noesd[1]
port 641 nsew signal bidirectional
flabel metal3 s 583520 360056 584800 360168 0 FreeSans 1120 0 0 0 gpio_noesd[2]
port 640 nsew signal bidirectional
flabel metal3 s 583520 406478 584800 406590 0 FreeSans 1120 0 0 0 gpio_noesd[3]
port 639 nsew signal bidirectional
flabel metal3 s 583520 450900 584800 451012 0 FreeSans 1120 0 0 0 gpio_noesd[4]
port 638 nsew signal bidirectional
flabel metal3 s 583520 495322 584800 495434 0 FreeSans 1120 0 0 0 gpio_noesd[5]
port 637 nsew signal bidirectional
flabel metal3 s 583520 584744 584800 584856 0 FreeSans 1120 0 0 0 gpio_noesd[6]
port 636 nsew signal bidirectional
flabel metal3 s -800 467126 480 467238 0 FreeSans 1120 0 0 0 gpio_noesd[8]
port 634 nsew signal bidirectional
flabel metal3 s -800 423904 480 424016 0 FreeSans 1120 0 0 0 gpio_noesd[9]
port 633 nsew signal bidirectional
flabel metal3 s 582300 677984 584800 682984 0 FreeSans 1120 0 0 0 io_analog[0]
port 653 nsew signal bidirectional
flabel metal3 s 566594 702300 571594 704800 0 FreeSans 1920 180 0 0 io_analog[1]
port 652 nsew signal bidirectional
flabel metal3 s 465394 702300 470394 704800 0 FreeSans 1920 180 0 0 io_analog[2]
port 651 nsew signal bidirectional
flabel metal3 s 413394 702300 418394 704800 0 FreeSans 1920 180 0 0 io_analog[3]
port 650 nsew signal bidirectional
flabel metal5 s 329294 702300 334294 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 649 nsew signal bidirectional
flabel metal5 s 227594 702300 232594 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 648 nsew signal bidirectional
flabel metal5 s 175894 702300 180894 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 647 nsew signal bidirectional
flabel metal5 s 318994 702300 323994 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 649 nsew signal bidirectional
flabel metal5 s 217294 702300 222294 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 648 nsew signal bidirectional
flabel metal5 s 165594 702300 170594 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 647 nsew signal bidirectional
flabel metal3 s 583520 2726 584800 2838 0 FreeSans 1120 0 0 0 io_in[0]
port 525 nsew signal input
flabel metal3 s 583520 408842 584800 408954 0 FreeSans 1120 0 0 0 io_in[10]
port 515 nsew signal input
flabel metal3 s 583520 453264 584800 453376 0 FreeSans 1120 0 0 0 io_in[11]
port 514 nsew signal input
flabel metal3 s 583520 497686 584800 497798 0 FreeSans 1120 0 0 0 io_in[12]
port 513 nsew signal input
flabel metal3 s 583520 587108 584800 587220 0 FreeSans 1120 0 0 0 io_in[13]
port 512 nsew signal input
flabel metal3 s -800 464762 480 464874 0 FreeSans 1120 0 0 0 io_in[15]
port 510 nsew signal input
flabel metal3 s -800 421540 480 421652 0 FreeSans 1120 0 0 0 io_in[16]
port 509 nsew signal input
flabel metal3 s -800 378318 480 378430 0 FreeSans 1120 0 0 0 io_in[17]
port 508 nsew signal input
flabel metal3 s -800 335096 480 335208 0 FreeSans 1120 0 0 0 io_in[18]
port 507 nsew signal input
flabel metal3 s -800 291874 480 291986 0 FreeSans 1120 0 0 0 io_in[19]
port 506 nsew signal input
flabel metal3 s 583520 7454 584800 7566 0 FreeSans 1120 0 0 0 io_in[1]
port 524 nsew signal input
flabel metal3 s -800 248852 480 248964 0 FreeSans 1120 0 0 0 io_in[20]
port 505 nsew signal input
flabel metal3 s -800 121230 480 121342 0 FreeSans 1120 0 0 0 io_in[21]
port 504 nsew signal input
flabel metal3 s -800 78008 480 78120 0 FreeSans 1120 0 0 0 io_in[22]
port 503 nsew signal input
flabel metal3 s -800 34786 480 34898 0 FreeSans 1120 0 0 0 io_in[23]
port 502 nsew signal input
flabel metal3 s -800 13364 480 13476 0 FreeSans 1120 0 0 0 io_in[24]
port 501 nsew signal input
flabel metal3 s -800 8636 480 8748 0 FreeSans 1120 0 0 0 io_in[25]
port 500 nsew signal input
flabel metal3 s -800 3908 480 4020 0 FreeSans 1120 0 0 0 io_in[26]
port 499 nsew signal input
flabel metal3 s 583520 12182 584800 12294 0 FreeSans 1120 0 0 0 io_in[2]
port 523 nsew signal input
flabel metal3 s 583520 16910 584800 17022 0 FreeSans 1120 0 0 0 io_in[3]
port 522 nsew signal input
flabel metal3 s 583520 21638 584800 21750 0 FreeSans 1120 0 0 0 io_in[4]
port 521 nsew signal input
flabel metal3 s 583520 48096 584800 48208 0 FreeSans 1120 0 0 0 io_in[5]
port 520 nsew signal input
flabel metal3 s 583520 92754 584800 92866 0 FreeSans 1120 0 0 0 io_in[6]
port 519 nsew signal input
flabel metal3 s 583520 272776 584800 272888 0 FreeSans 1120 0 0 0 io_in[7]
port 518 nsew signal input
flabel metal3 s 583520 317198 584800 317310 0 FreeSans 1120 0 0 0 io_in[8]
port 517 nsew signal input
flabel metal3 s 583520 362420 584800 362532 0 FreeSans 1120 0 0 0 io_in[9]
port 516 nsew signal input
flabel metal3 s 583520 1544 584800 1656 0 FreeSans 1120 0 0 0 io_in_3v3[0]
port 552 nsew signal input
flabel metal3 s 583520 407660 584800 407772 0 FreeSans 1120 0 0 0 io_in_3v3[10]
port 542 nsew signal input
flabel metal3 s 583520 452082 584800 452194 0 FreeSans 1120 0 0 0 io_in_3v3[11]
port 541 nsew signal input
flabel metal3 s 583520 496504 584800 496616 0 FreeSans 1120 0 0 0 io_in_3v3[12]
port 540 nsew signal input
flabel metal3 s 583520 585926 584800 586038 0 FreeSans 1120 0 0 0 io_in_3v3[13]
port 539 nsew signal input
flabel metal3 s -800 465944 480 466056 0 FreeSans 1120 0 0 0 io_in_3v3[15]
port 537 nsew signal input
flabel metal3 s -800 422722 480 422834 0 FreeSans 1120 0 0 0 io_in_3v3[16]
port 536 nsew signal input
flabel metal3 s -800 379500 480 379612 0 FreeSans 1120 0 0 0 io_in_3v3[17]
port 535 nsew signal input
flabel metal3 s -800 336278 480 336390 0 FreeSans 1120 0 0 0 io_in_3v3[18]
port 534 nsew signal input
flabel metal3 s -800 293056 480 293168 0 FreeSans 1120 0 0 0 io_in_3v3[19]
port 533 nsew signal input
flabel metal3 s 583520 6272 584800 6384 0 FreeSans 1120 0 0 0 io_in_3v3[1]
port 551 nsew signal input
flabel metal3 s -800 250034 480 250146 0 FreeSans 1120 0 0 0 io_in_3v3[20]
port 532 nsew signal input
flabel metal3 s -800 122412 480 122524 0 FreeSans 1120 0 0 0 io_in_3v3[21]
port 531 nsew signal input
flabel metal3 s -800 79190 480 79302 0 FreeSans 1120 0 0 0 io_in_3v3[22]
port 530 nsew signal input
flabel metal3 s -800 35968 480 36080 0 FreeSans 1120 0 0 0 io_in_3v3[23]
port 529 nsew signal input
flabel metal3 s -800 14546 480 14658 0 FreeSans 1120 0 0 0 io_in_3v3[24]
port 528 nsew signal input
flabel metal3 s -800 9818 480 9930 0 FreeSans 1120 0 0 0 io_in_3v3[25]
port 527 nsew signal input
flabel metal3 s -800 5090 480 5202 0 FreeSans 1120 0 0 0 io_in_3v3[26]
port 526 nsew signal input
flabel metal3 s 583520 11000 584800 11112 0 FreeSans 1120 0 0 0 io_in_3v3[2]
port 550 nsew signal input
flabel metal3 s 583520 15728 584800 15840 0 FreeSans 1120 0 0 0 io_in_3v3[3]
port 549 nsew signal input
flabel metal3 s 583520 20456 584800 20568 0 FreeSans 1120 0 0 0 io_in_3v3[4]
port 548 nsew signal input
flabel metal3 s 583520 46914 584800 47026 0 FreeSans 1120 0 0 0 io_in_3v3[5]
port 547 nsew signal input
flabel metal3 s 583520 91572 584800 91684 0 FreeSans 1120 0 0 0 io_in_3v3[6]
port 546 nsew signal input
flabel metal3 s 583520 271594 584800 271706 0 FreeSans 1120 0 0 0 io_in_3v3[7]
port 545 nsew signal input
flabel metal3 s 583520 316016 584800 316128 0 FreeSans 1120 0 0 0 io_in_3v3[8]
port 544 nsew signal input
flabel metal3 s 583520 361238 584800 361350 0 FreeSans 1120 0 0 0 io_in_3v3[9]
port 543 nsew signal input
flabel metal3 s 583520 5090 584800 5202 0 FreeSans 1120 0 0 0 io_oeb[0]
port 606 nsew signal tristate
flabel metal3 s 583520 411206 584800 411318 0 FreeSans 1120 0 0 0 io_oeb[10]
port 596 nsew signal tristate
flabel metal3 s 583520 455628 584800 455740 0 FreeSans 1120 0 0 0 io_oeb[11]
port 595 nsew signal tristate
flabel metal3 s 583520 500050 584800 500162 0 FreeSans 1120 0 0 0 io_oeb[12]
port 594 nsew signal tristate
flabel metal3 s 583520 589472 584800 589584 0 FreeSans 1120 0 0 0 io_oeb[13]
port 593 nsew signal tristate
flabel metal3 s -800 462398 480 462510 0 FreeSans 1120 0 0 0 io_oeb[15]
port 591 nsew signal tristate
flabel metal3 s -800 419176 480 419288 0 FreeSans 1120 0 0 0 io_oeb[16]
port 590 nsew signal tristate
flabel metal3 s -800 375954 480 376066 0 FreeSans 1120 0 0 0 io_oeb[17]
port 589 nsew signal tristate
flabel metal3 s -800 332732 480 332844 0 FreeSans 1120 0 0 0 io_oeb[18]
port 588 nsew signal tristate
flabel metal3 s -800 289510 480 289622 0 FreeSans 1120 0 0 0 io_oeb[19]
port 587 nsew signal tristate
flabel metal3 s 583520 9818 584800 9930 0 FreeSans 1120 0 0 0 io_oeb[1]
port 605 nsew signal tristate
flabel metal3 s -800 246488 480 246600 0 FreeSans 1120 0 0 0 io_oeb[20]
port 586 nsew signal tristate
flabel metal3 s -800 118866 480 118978 0 FreeSans 1120 0 0 0 io_oeb[21]
port 585 nsew signal tristate
flabel metal3 s -800 75644 480 75756 0 FreeSans 1120 0 0 0 io_oeb[22]
port 584 nsew signal tristate
flabel metal3 s -800 32422 480 32534 0 FreeSans 1120 0 0 0 io_oeb[23]
port 583 nsew signal tristate
flabel metal3 s -800 11000 480 11112 0 FreeSans 1120 0 0 0 io_oeb[24]
port 582 nsew signal tristate
flabel metal3 s -800 6272 480 6384 0 FreeSans 1120 0 0 0 io_oeb[25]
port 581 nsew signal tristate
flabel metal3 s -800 1544 480 1656 0 FreeSans 1120 0 0 0 io_oeb[26]
port 580 nsew signal tristate
flabel metal3 s 583520 14546 584800 14658 0 FreeSans 1120 0 0 0 io_oeb[2]
port 604 nsew signal tristate
flabel metal3 s 583520 19274 584800 19386 0 FreeSans 1120 0 0 0 io_oeb[3]
port 603 nsew signal tristate
flabel metal3 s 583520 24002 584800 24114 0 FreeSans 1120 0 0 0 io_oeb[4]
port 602 nsew signal tristate
flabel metal3 s 583520 50460 584800 50572 0 FreeSans 1120 0 0 0 io_oeb[5]
port 601 nsew signal tristate
flabel metal3 s 583520 95118 584800 95230 0 FreeSans 1120 0 0 0 io_oeb[6]
port 600 nsew signal tristate
flabel metal3 s 583520 275140 584800 275252 0 FreeSans 1120 0 0 0 io_oeb[7]
port 599 nsew signal tristate
flabel metal3 s 583520 319562 584800 319674 0 FreeSans 1120 0 0 0 io_oeb[8]
port 598 nsew signal tristate
flabel metal3 s 583520 364784 584800 364896 0 FreeSans 1120 0 0 0 io_oeb[9]
port 597 nsew signal tristate
flabel metal3 s 583520 3908 584800 4020 0 FreeSans 1120 0 0 0 io_out[0]
port 579 nsew signal tristate
flabel metal3 s 583520 410024 584800 410136 0 FreeSans 1120 0 0 0 io_out[10]
port 569 nsew signal tristate
flabel metal3 s 583520 454446 584800 454558 0 FreeSans 1120 0 0 0 io_out[11]
port 568 nsew signal tristate
flabel metal3 s 583520 498868 584800 498980 0 FreeSans 1120 0 0 0 io_out[12]
port 567 nsew signal tristate
flabel metal3 s 583520 588290 584800 588402 0 FreeSans 1120 0 0 0 io_out[13]
port 566 nsew signal tristate
flabel metal3 s -800 463580 480 463692 0 FreeSans 1120 0 0 0 io_out[15]
port 564 nsew signal tristate
flabel metal3 s -800 420358 480 420470 0 FreeSans 1120 0 0 0 io_out[16]
port 563 nsew signal tristate
flabel metal3 s -800 377136 480 377248 0 FreeSans 1120 0 0 0 io_out[17]
port 562 nsew signal tristate
flabel metal3 s -800 333914 480 334026 0 FreeSans 1120 0 0 0 io_out[18]
port 561 nsew signal tristate
flabel metal3 s -800 290692 480 290804 0 FreeSans 1120 0 0 0 io_out[19]
port 560 nsew signal tristate
flabel metal3 s 583520 8636 584800 8748 0 FreeSans 1120 0 0 0 io_out[1]
port 578 nsew signal tristate
flabel metal3 s -800 247670 480 247782 0 FreeSans 1120 0 0 0 io_out[20]
port 559 nsew signal tristate
flabel metal3 s -800 120048 480 120160 0 FreeSans 1120 0 0 0 io_out[21]
port 558 nsew signal tristate
flabel metal3 s -800 76826 480 76938 0 FreeSans 1120 0 0 0 io_out[22]
port 557 nsew signal tristate
flabel metal3 s -800 33604 480 33716 0 FreeSans 1120 0 0 0 io_out[23]
port 556 nsew signal tristate
flabel metal3 s -800 12182 480 12294 0 FreeSans 1120 0 0 0 io_out[24]
port 555 nsew signal tristate
flabel metal3 s -800 7454 480 7566 0 FreeSans 1120 0 0 0 io_out[25]
port 554 nsew signal tristate
flabel metal3 s -800 2726 480 2838 0 FreeSans 1120 0 0 0 io_out[26]
port 553 nsew signal tristate
flabel metal3 s 583520 13364 584800 13476 0 FreeSans 1120 0 0 0 io_out[2]
port 577 nsew signal tristate
flabel metal3 s 583520 18092 584800 18204 0 FreeSans 1120 0 0 0 io_out[3]
port 576 nsew signal tristate
flabel metal3 s 583520 22820 584800 22932 0 FreeSans 1120 0 0 0 io_out[4]
port 575 nsew signal tristate
flabel metal3 s 583520 49278 584800 49390 0 FreeSans 1120 0 0 0 io_out[5]
port 574 nsew signal tristate
flabel metal3 s 583520 93936 584800 94048 0 FreeSans 1120 0 0 0 io_out[6]
port 573 nsew signal tristate
flabel metal3 s 583520 273958 584800 274070 0 FreeSans 1120 0 0 0 io_out[7]
port 572 nsew signal tristate
flabel metal3 s 583520 318380 584800 318492 0 FreeSans 1120 0 0 0 io_out[8]
port 571 nsew signal tristate
flabel metal3 s 583520 363602 584800 363714 0 FreeSans 1120 0 0 0 io_out[9]
port 570 nsew signal tristate
flabel metal2 s 125816 -800 125928 480 0 FreeSans 1120 90 0 0 la_data_in[0]
port 242 nsew signal input
flabel metal2 s 480416 -800 480528 480 0 FreeSans 1120 90 0 0 la_data_in[100]
port 142 nsew signal input
flabel metal2 s 483962 -800 484074 480 0 FreeSans 1120 90 0 0 la_data_in[101]
port 141 nsew signal input
flabel metal2 s 487508 -800 487620 480 0 FreeSans 1120 90 0 0 la_data_in[102]
port 140 nsew signal input
flabel metal2 s 491054 -800 491166 480 0 FreeSans 1120 90 0 0 la_data_in[103]
port 139 nsew signal input
flabel metal2 s 494600 -800 494712 480 0 FreeSans 1120 90 0 0 la_data_in[104]
port 138 nsew signal input
flabel metal2 s 498146 -800 498258 480 0 FreeSans 1120 90 0 0 la_data_in[105]
port 137 nsew signal input
flabel metal2 s 501692 -800 501804 480 0 FreeSans 1120 90 0 0 la_data_in[106]
port 136 nsew signal input
flabel metal2 s 505238 -800 505350 480 0 FreeSans 1120 90 0 0 la_data_in[107]
port 135 nsew signal input
flabel metal2 s 508784 -800 508896 480 0 FreeSans 1120 90 0 0 la_data_in[108]
port 134 nsew signal input
flabel metal2 s 512330 -800 512442 480 0 FreeSans 1120 90 0 0 la_data_in[109]
port 133 nsew signal input
flabel metal2 s 161276 -800 161388 480 0 FreeSans 1120 90 0 0 la_data_in[10]
port 232 nsew signal input
flabel metal2 s 515876 -800 515988 480 0 FreeSans 1120 90 0 0 la_data_in[110]
port 132 nsew signal input
flabel metal2 s 519422 -800 519534 480 0 FreeSans 1120 90 0 0 la_data_in[111]
port 131 nsew signal input
flabel metal2 s 522968 -800 523080 480 0 FreeSans 1120 90 0 0 la_data_in[112]
port 130 nsew signal input
flabel metal2 s 526514 -800 526626 480 0 FreeSans 1120 90 0 0 la_data_in[113]
port 129 nsew signal input
flabel metal2 s 530060 -800 530172 480 0 FreeSans 1120 90 0 0 la_data_in[114]
port 128 nsew signal input
flabel metal2 s 533606 -800 533718 480 0 FreeSans 1120 90 0 0 la_data_in[115]
port 127 nsew signal input
flabel metal2 s 537152 -800 537264 480 0 FreeSans 1120 90 0 0 la_data_in[116]
port 126 nsew signal input
flabel metal2 s 540698 -800 540810 480 0 FreeSans 1120 90 0 0 la_data_in[117]
port 125 nsew signal input
flabel metal2 s 544244 -800 544356 480 0 FreeSans 1120 90 0 0 la_data_in[118]
port 124 nsew signal input
flabel metal2 s 547790 -800 547902 480 0 FreeSans 1120 90 0 0 la_data_in[119]
port 123 nsew signal input
flabel metal2 s 164822 -800 164934 480 0 FreeSans 1120 90 0 0 la_data_in[11]
port 231 nsew signal input
flabel metal2 s 551336 -800 551448 480 0 FreeSans 1120 90 0 0 la_data_in[120]
port 122 nsew signal input
flabel metal2 s 554882 -800 554994 480 0 FreeSans 1120 90 0 0 la_data_in[121]
port 121 nsew signal input
flabel metal2 s 558428 -800 558540 480 0 FreeSans 1120 90 0 0 la_data_in[122]
port 120 nsew signal input
flabel metal2 s 561974 -800 562086 480 0 FreeSans 1120 90 0 0 la_data_in[123]
port 119 nsew signal input
flabel metal2 s 565520 -800 565632 480 0 FreeSans 1120 90 0 0 la_data_in[124]
port 118 nsew signal input
flabel metal2 s 569066 -800 569178 480 0 FreeSans 1120 90 0 0 la_data_in[125]
port 117 nsew signal input
flabel metal2 s 572612 -800 572724 480 0 FreeSans 1120 90 0 0 la_data_in[126]
port 116 nsew signal input
flabel metal2 s 576158 -800 576270 480 0 FreeSans 1120 90 0 0 la_data_in[127]
port 115 nsew signal input
flabel metal2 s 168368 -800 168480 480 0 FreeSans 1120 90 0 0 la_data_in[12]
port 230 nsew signal input
flabel metal2 s 171914 -800 172026 480 0 FreeSans 1120 90 0 0 la_data_in[13]
port 229 nsew signal input
flabel metal2 s 175460 -800 175572 480 0 FreeSans 1120 90 0 0 la_data_in[14]
port 228 nsew signal input
flabel metal2 s 179006 -800 179118 480 0 FreeSans 1120 90 0 0 la_data_in[15]
port 227 nsew signal input
flabel metal2 s 182552 -800 182664 480 0 FreeSans 1120 90 0 0 la_data_in[16]
port 226 nsew signal input
flabel metal2 s 186098 -800 186210 480 0 FreeSans 1120 90 0 0 la_data_in[17]
port 225 nsew signal input
flabel metal2 s 189644 -800 189756 480 0 FreeSans 1120 90 0 0 la_data_in[18]
port 224 nsew signal input
flabel metal2 s 193190 -800 193302 480 0 FreeSans 1120 90 0 0 la_data_in[19]
port 223 nsew signal input
flabel metal2 s 129362 -800 129474 480 0 FreeSans 1120 90 0 0 la_data_in[1]
port 241 nsew signal input
flabel metal2 s 196736 -800 196848 480 0 FreeSans 1120 90 0 0 la_data_in[20]
port 222 nsew signal input
flabel metal2 s 200282 -800 200394 480 0 FreeSans 1120 90 0 0 la_data_in[21]
port 221 nsew signal input
flabel metal2 s 203828 -800 203940 480 0 FreeSans 1120 90 0 0 la_data_in[22]
port 220 nsew signal input
flabel metal2 s 207374 -800 207486 480 0 FreeSans 1120 90 0 0 la_data_in[23]
port 219 nsew signal input
flabel metal2 s 210920 -800 211032 480 0 FreeSans 1120 90 0 0 la_data_in[24]
port 218 nsew signal input
flabel metal2 s 214466 -800 214578 480 0 FreeSans 1120 90 0 0 la_data_in[25]
port 217 nsew signal input
flabel metal2 s 218012 -800 218124 480 0 FreeSans 1120 90 0 0 la_data_in[26]
port 216 nsew signal input
flabel metal2 s 221558 -800 221670 480 0 FreeSans 1120 90 0 0 la_data_in[27]
port 215 nsew signal input
flabel metal2 s 225104 -800 225216 480 0 FreeSans 1120 90 0 0 la_data_in[28]
port 214 nsew signal input
flabel metal2 s 228650 -800 228762 480 0 FreeSans 1120 90 0 0 la_data_in[29]
port 213 nsew signal input
flabel metal2 s 132908 -800 133020 480 0 FreeSans 1120 90 0 0 la_data_in[2]
port 240 nsew signal input
flabel metal2 s 232196 -800 232308 480 0 FreeSans 1120 90 0 0 la_data_in[30]
port 212 nsew signal input
flabel metal2 s 235742 -800 235854 480 0 FreeSans 1120 90 0 0 la_data_in[31]
port 211 nsew signal input
flabel metal2 s 239288 -800 239400 480 0 FreeSans 1120 90 0 0 la_data_in[32]
port 210 nsew signal input
flabel metal2 s 242834 -800 242946 480 0 FreeSans 1120 90 0 0 la_data_in[33]
port 209 nsew signal input
flabel metal2 s 246380 -800 246492 480 0 FreeSans 1120 90 0 0 la_data_in[34]
port 208 nsew signal input
flabel metal2 s 249926 -800 250038 480 0 FreeSans 1120 90 0 0 la_data_in[35]
port 207 nsew signal input
flabel metal2 s 253472 -800 253584 480 0 FreeSans 1120 90 0 0 la_data_in[36]
port 206 nsew signal input
flabel metal2 s 257018 -800 257130 480 0 FreeSans 1120 90 0 0 la_data_in[37]
port 205 nsew signal input
flabel metal2 s 260564 -800 260676 480 0 FreeSans 1120 90 0 0 la_data_in[38]
port 204 nsew signal input
flabel metal2 s 264110 -800 264222 480 0 FreeSans 1120 90 0 0 la_data_in[39]
port 203 nsew signal input
flabel metal2 s 136454 -800 136566 480 0 FreeSans 1120 90 0 0 la_data_in[3]
port 239 nsew signal input
flabel metal2 s 267656 -800 267768 480 0 FreeSans 1120 90 0 0 la_data_in[40]
port 202 nsew signal input
flabel metal2 s 271202 -800 271314 480 0 FreeSans 1120 90 0 0 la_data_in[41]
port 201 nsew signal input
flabel metal2 s 274748 -800 274860 480 0 FreeSans 1120 90 0 0 la_data_in[42]
port 200 nsew signal input
flabel metal2 s 278294 -800 278406 480 0 FreeSans 1120 90 0 0 la_data_in[43]
port 199 nsew signal input
flabel metal2 s 281840 -800 281952 480 0 FreeSans 1120 90 0 0 la_data_in[44]
port 198 nsew signal input
flabel metal2 s 285386 -800 285498 480 0 FreeSans 1120 90 0 0 la_data_in[45]
port 197 nsew signal input
flabel metal2 s 288932 -800 289044 480 0 FreeSans 1120 90 0 0 la_data_in[46]
port 196 nsew signal input
flabel metal2 s 292478 -800 292590 480 0 FreeSans 1120 90 0 0 la_data_in[47]
port 195 nsew signal input
flabel metal2 s 296024 -800 296136 480 0 FreeSans 1120 90 0 0 la_data_in[48]
port 194 nsew signal input
flabel metal2 s 299570 -800 299682 480 0 FreeSans 1120 90 0 0 la_data_in[49]
port 193 nsew signal input
flabel metal2 s 140000 -800 140112 480 0 FreeSans 1120 90 0 0 la_data_in[4]
port 238 nsew signal input
flabel metal2 s 303116 -800 303228 480 0 FreeSans 1120 90 0 0 la_data_in[50]
port 192 nsew signal input
flabel metal2 s 306662 -800 306774 480 0 FreeSans 1120 90 0 0 la_data_in[51]
port 191 nsew signal input
flabel metal2 s 310208 -800 310320 480 0 FreeSans 1120 90 0 0 la_data_in[52]
port 190 nsew signal input
flabel metal2 s 313754 -800 313866 480 0 FreeSans 1120 90 0 0 la_data_in[53]
port 189 nsew signal input
flabel metal2 s 317300 -800 317412 480 0 FreeSans 1120 90 0 0 la_data_in[54]
port 188 nsew signal input
flabel metal2 s 320846 -800 320958 480 0 FreeSans 1120 90 0 0 la_data_in[55]
port 187 nsew signal input
flabel metal2 s 324392 -800 324504 480 0 FreeSans 1120 90 0 0 la_data_in[56]
port 186 nsew signal input
flabel metal2 s 327938 -800 328050 480 0 FreeSans 1120 90 0 0 la_data_in[57]
port 185 nsew signal input
flabel metal2 s 331484 -800 331596 480 0 FreeSans 1120 90 0 0 la_data_in[58]
port 184 nsew signal input
flabel metal2 s 335030 -800 335142 480 0 FreeSans 1120 90 0 0 la_data_in[59]
port 183 nsew signal input
flabel metal2 s 143546 -800 143658 480 0 FreeSans 1120 90 0 0 la_data_in[5]
port 237 nsew signal input
flabel metal2 s 338576 -800 338688 480 0 FreeSans 1120 90 0 0 la_data_in[60]
port 182 nsew signal input
flabel metal2 s 342122 -800 342234 480 0 FreeSans 1120 90 0 0 la_data_in[61]
port 181 nsew signal input
flabel metal2 s 345668 -800 345780 480 0 FreeSans 1120 90 0 0 la_data_in[62]
port 180 nsew signal input
flabel metal2 s 349214 -800 349326 480 0 FreeSans 1120 90 0 0 la_data_in[63]
port 179 nsew signal input
flabel metal2 s 352760 -800 352872 480 0 FreeSans 1120 90 0 0 la_data_in[64]
port 178 nsew signal input
flabel metal2 s 356306 -800 356418 480 0 FreeSans 1120 90 0 0 la_data_in[65]
port 177 nsew signal input
flabel metal2 s 359852 -800 359964 480 0 FreeSans 1120 90 0 0 la_data_in[66]
port 176 nsew signal input
flabel metal2 s 363398 -800 363510 480 0 FreeSans 1120 90 0 0 la_data_in[67]
port 175 nsew signal input
flabel metal2 s 366944 -800 367056 480 0 FreeSans 1120 90 0 0 la_data_in[68]
port 174 nsew signal input
flabel metal2 s 370490 -800 370602 480 0 FreeSans 1120 90 0 0 la_data_in[69]
port 173 nsew signal input
flabel metal2 s 147092 -800 147204 480 0 FreeSans 1120 90 0 0 la_data_in[6]
port 236 nsew signal input
flabel metal2 s 374036 -800 374148 480 0 FreeSans 1120 90 0 0 la_data_in[70]
port 172 nsew signal input
flabel metal2 s 377582 -800 377694 480 0 FreeSans 1120 90 0 0 la_data_in[71]
port 171 nsew signal input
flabel metal2 s 381128 -800 381240 480 0 FreeSans 1120 90 0 0 la_data_in[72]
port 170 nsew signal input
flabel metal2 s 384674 -800 384786 480 0 FreeSans 1120 90 0 0 la_data_in[73]
port 169 nsew signal input
flabel metal2 s 388220 -800 388332 480 0 FreeSans 1120 90 0 0 la_data_in[74]
port 168 nsew signal input
flabel metal2 s 391766 -800 391878 480 0 FreeSans 1120 90 0 0 la_data_in[75]
port 167 nsew signal input
flabel metal2 s 395312 -800 395424 480 0 FreeSans 1120 90 0 0 la_data_in[76]
port 166 nsew signal input
flabel metal2 s 398858 -800 398970 480 0 FreeSans 1120 90 0 0 la_data_in[77]
port 165 nsew signal input
flabel metal2 s 402404 -800 402516 480 0 FreeSans 1120 90 0 0 la_data_in[78]
port 164 nsew signal input
flabel metal2 s 405950 -800 406062 480 0 FreeSans 1120 90 0 0 la_data_in[79]
port 163 nsew signal input
flabel metal2 s 150638 -800 150750 480 0 FreeSans 1120 90 0 0 la_data_in[7]
port 235 nsew signal input
flabel metal2 s 409496 -800 409608 480 0 FreeSans 1120 90 0 0 la_data_in[80]
port 162 nsew signal input
flabel metal2 s 413042 -800 413154 480 0 FreeSans 1120 90 0 0 la_data_in[81]
port 161 nsew signal input
flabel metal2 s 416588 -800 416700 480 0 FreeSans 1120 90 0 0 la_data_in[82]
port 160 nsew signal input
flabel metal2 s 420134 -800 420246 480 0 FreeSans 1120 90 0 0 la_data_in[83]
port 159 nsew signal input
flabel metal2 s 423680 -800 423792 480 0 FreeSans 1120 90 0 0 la_data_in[84]
port 158 nsew signal input
flabel metal2 s 427226 -800 427338 480 0 FreeSans 1120 90 0 0 la_data_in[85]
port 157 nsew signal input
flabel metal2 s 430772 -800 430884 480 0 FreeSans 1120 90 0 0 la_data_in[86]
port 156 nsew signal input
flabel metal2 s 434318 -800 434430 480 0 FreeSans 1120 90 0 0 la_data_in[87]
port 155 nsew signal input
flabel metal2 s 437864 -800 437976 480 0 FreeSans 1120 90 0 0 la_data_in[88]
port 154 nsew signal input
flabel metal2 s 441410 -800 441522 480 0 FreeSans 1120 90 0 0 la_data_in[89]
port 153 nsew signal input
flabel metal2 s 154184 -800 154296 480 0 FreeSans 1120 90 0 0 la_data_in[8]
port 234 nsew signal input
flabel metal2 s 444956 -800 445068 480 0 FreeSans 1120 90 0 0 la_data_in[90]
port 152 nsew signal input
flabel metal2 s 448502 -800 448614 480 0 FreeSans 1120 90 0 0 la_data_in[91]
port 151 nsew signal input
flabel metal2 s 452048 -800 452160 480 0 FreeSans 1120 90 0 0 la_data_in[92]
port 150 nsew signal input
flabel metal2 s 455594 -800 455706 480 0 FreeSans 1120 90 0 0 la_data_in[93]
port 149 nsew signal input
flabel metal2 s 459140 -800 459252 480 0 FreeSans 1120 90 0 0 la_data_in[94]
port 148 nsew signal input
flabel metal2 s 462686 -800 462798 480 0 FreeSans 1120 90 0 0 la_data_in[95]
port 147 nsew signal input
flabel metal2 s 466232 -800 466344 480 0 FreeSans 1120 90 0 0 la_data_in[96]
port 146 nsew signal input
flabel metal2 s 469778 -800 469890 480 0 FreeSans 1120 90 0 0 la_data_in[97]
port 145 nsew signal input
flabel metal2 s 473324 -800 473436 480 0 FreeSans 1120 90 0 0 la_data_in[98]
port 144 nsew signal input
flabel metal2 s 476870 -800 476982 480 0 FreeSans 1120 90 0 0 la_data_in[99]
port 143 nsew signal input
flabel metal2 s 157730 -800 157842 480 0 FreeSans 1120 90 0 0 la_data_in[9]
port 233 nsew signal input
flabel metal2 s 126998 -800 127110 480 0 FreeSans 1120 90 0 0 la_data_out[0]
port 370 nsew signal tristate
flabel metal2 s 481598 -800 481710 480 0 FreeSans 1120 90 0 0 la_data_out[100]
port 270 nsew signal tristate
flabel metal2 s 485144 -800 485256 480 0 FreeSans 1120 90 0 0 la_data_out[101]
port 269 nsew signal tristate
flabel metal2 s 488690 -800 488802 480 0 FreeSans 1120 90 0 0 la_data_out[102]
port 268 nsew signal tristate
flabel metal2 s 492236 -800 492348 480 0 FreeSans 1120 90 0 0 la_data_out[103]
port 267 nsew signal tristate
flabel metal2 s 495782 -800 495894 480 0 FreeSans 1120 90 0 0 la_data_out[104]
port 266 nsew signal tristate
flabel metal2 s 499328 -800 499440 480 0 FreeSans 1120 90 0 0 la_data_out[105]
port 265 nsew signal tristate
flabel metal2 s 502874 -800 502986 480 0 FreeSans 1120 90 0 0 la_data_out[106]
port 264 nsew signal tristate
flabel metal2 s 506420 -800 506532 480 0 FreeSans 1120 90 0 0 la_data_out[107]
port 263 nsew signal tristate
flabel metal2 s 509966 -800 510078 480 0 FreeSans 1120 90 0 0 la_data_out[108]
port 262 nsew signal tristate
flabel metal2 s 513512 -800 513624 480 0 FreeSans 1120 90 0 0 la_data_out[109]
port 261 nsew signal tristate
flabel metal2 s 162458 -800 162570 480 0 FreeSans 1120 90 0 0 la_data_out[10]
port 360 nsew signal tristate
flabel metal2 s 517058 -800 517170 480 0 FreeSans 1120 90 0 0 la_data_out[110]
port 260 nsew signal tristate
flabel metal2 s 520604 -800 520716 480 0 FreeSans 1120 90 0 0 la_data_out[111]
port 259 nsew signal tristate
flabel metal2 s 524150 -800 524262 480 0 FreeSans 1120 90 0 0 la_data_out[112]
port 258 nsew signal tristate
flabel metal2 s 527696 -800 527808 480 0 FreeSans 1120 90 0 0 la_data_out[113]
port 257 nsew signal tristate
flabel metal2 s 531242 -800 531354 480 0 FreeSans 1120 90 0 0 la_data_out[114]
port 256 nsew signal tristate
flabel metal2 s 534788 -800 534900 480 0 FreeSans 1120 90 0 0 la_data_out[115]
port 255 nsew signal tristate
flabel metal2 s 538334 -800 538446 480 0 FreeSans 1120 90 0 0 la_data_out[116]
port 254 nsew signal tristate
flabel metal2 s 541880 -800 541992 480 0 FreeSans 1120 90 0 0 la_data_out[117]
port 253 nsew signal tristate
flabel metal2 s 545426 -800 545538 480 0 FreeSans 1120 90 0 0 la_data_out[118]
port 252 nsew signal tristate
flabel metal2 s 548972 -800 549084 480 0 FreeSans 1120 90 0 0 la_data_out[119]
port 251 nsew signal tristate
flabel metal2 s 166004 -800 166116 480 0 FreeSans 1120 90 0 0 la_data_out[11]
port 359 nsew signal tristate
flabel metal2 s 552518 -800 552630 480 0 FreeSans 1120 90 0 0 la_data_out[120]
port 250 nsew signal tristate
flabel metal2 s 556064 -800 556176 480 0 FreeSans 1120 90 0 0 la_data_out[121]
port 249 nsew signal tristate
flabel metal2 s 559610 -800 559722 480 0 FreeSans 1120 90 0 0 la_data_out[122]
port 248 nsew signal tristate
flabel metal2 s 563156 -800 563268 480 0 FreeSans 1120 90 0 0 la_data_out[123]
port 247 nsew signal tristate
flabel metal2 s 566702 -800 566814 480 0 FreeSans 1120 90 0 0 la_data_out[124]
port 246 nsew signal tristate
flabel metal2 s 570248 -800 570360 480 0 FreeSans 1120 90 0 0 la_data_out[125]
port 245 nsew signal tristate
flabel metal2 s 573794 -800 573906 480 0 FreeSans 1120 90 0 0 la_data_out[126]
port 244 nsew signal tristate
flabel metal2 s 577340 -800 577452 480 0 FreeSans 1120 90 0 0 la_data_out[127]
port 243 nsew signal tristate
flabel metal2 s 169550 -800 169662 480 0 FreeSans 1120 90 0 0 la_data_out[12]
port 358 nsew signal tristate
flabel metal2 s 173096 -800 173208 480 0 FreeSans 1120 90 0 0 la_data_out[13]
port 357 nsew signal tristate
flabel metal2 s 176642 -800 176754 480 0 FreeSans 1120 90 0 0 la_data_out[14]
port 356 nsew signal tristate
flabel metal2 s 180188 -800 180300 480 0 FreeSans 1120 90 0 0 la_data_out[15]
port 355 nsew signal tristate
flabel metal2 s 183734 -800 183846 480 0 FreeSans 1120 90 0 0 la_data_out[16]
port 354 nsew signal tristate
flabel metal2 s 187280 -800 187392 480 0 FreeSans 1120 90 0 0 la_data_out[17]
port 353 nsew signal tristate
flabel metal2 s 190826 -800 190938 480 0 FreeSans 1120 90 0 0 la_data_out[18]
port 352 nsew signal tristate
flabel metal2 s 194372 -800 194484 480 0 FreeSans 1120 90 0 0 la_data_out[19]
port 351 nsew signal tristate
flabel metal2 s 130544 -800 130656 480 0 FreeSans 1120 90 0 0 la_data_out[1]
port 369 nsew signal tristate
flabel metal2 s 197918 -800 198030 480 0 FreeSans 1120 90 0 0 la_data_out[20]
port 350 nsew signal tristate
flabel metal2 s 201464 -800 201576 480 0 FreeSans 1120 90 0 0 la_data_out[21]
port 349 nsew signal tristate
flabel metal2 s 205010 -800 205122 480 0 FreeSans 1120 90 0 0 la_data_out[22]
port 348 nsew signal tristate
flabel metal2 s 208556 -800 208668 480 0 FreeSans 1120 90 0 0 la_data_out[23]
port 347 nsew signal tristate
flabel metal2 s 212102 -800 212214 480 0 FreeSans 1120 90 0 0 la_data_out[24]
port 346 nsew signal tristate
flabel metal2 s 215648 -800 215760 480 0 FreeSans 1120 90 0 0 la_data_out[25]
port 345 nsew signal tristate
flabel metal2 s 219194 -800 219306 480 0 FreeSans 1120 90 0 0 la_data_out[26]
port 344 nsew signal tristate
flabel metal2 s 222740 -800 222852 480 0 FreeSans 1120 90 0 0 la_data_out[27]
port 343 nsew signal tristate
flabel metal2 s 226286 -800 226398 480 0 FreeSans 1120 90 0 0 la_data_out[28]
port 342 nsew signal tristate
flabel metal2 s 229832 -800 229944 480 0 FreeSans 1120 90 0 0 la_data_out[29]
port 341 nsew signal tristate
flabel metal2 s 134090 -800 134202 480 0 FreeSans 1120 90 0 0 la_data_out[2]
port 368 nsew signal tristate
flabel metal2 s 233378 -800 233490 480 0 FreeSans 1120 90 0 0 la_data_out[30]
port 340 nsew signal tristate
flabel metal2 s 236924 -800 237036 480 0 FreeSans 1120 90 0 0 la_data_out[31]
port 339 nsew signal tristate
flabel metal2 s 240470 -800 240582 480 0 FreeSans 1120 90 0 0 la_data_out[32]
port 338 nsew signal tristate
flabel metal2 s 244016 -800 244128 480 0 FreeSans 1120 90 0 0 la_data_out[33]
port 337 nsew signal tristate
flabel metal2 s 247562 -800 247674 480 0 FreeSans 1120 90 0 0 la_data_out[34]
port 336 nsew signal tristate
flabel metal2 s 251108 -800 251220 480 0 FreeSans 1120 90 0 0 la_data_out[35]
port 335 nsew signal tristate
flabel metal2 s 254654 -800 254766 480 0 FreeSans 1120 90 0 0 la_data_out[36]
port 334 nsew signal tristate
flabel metal2 s 258200 -800 258312 480 0 FreeSans 1120 90 0 0 la_data_out[37]
port 333 nsew signal tristate
flabel metal2 s 261746 -800 261858 480 0 FreeSans 1120 90 0 0 la_data_out[38]
port 332 nsew signal tristate
flabel metal2 s 265292 -800 265404 480 0 FreeSans 1120 90 0 0 la_data_out[39]
port 331 nsew signal tristate
flabel metal2 s 137636 -800 137748 480 0 FreeSans 1120 90 0 0 la_data_out[3]
port 367 nsew signal tristate
flabel metal2 s 268838 -800 268950 480 0 FreeSans 1120 90 0 0 la_data_out[40]
port 330 nsew signal tristate
flabel metal2 s 272384 -800 272496 480 0 FreeSans 1120 90 0 0 la_data_out[41]
port 329 nsew signal tristate
flabel metal2 s 275930 -800 276042 480 0 FreeSans 1120 90 0 0 la_data_out[42]
port 328 nsew signal tristate
flabel metal2 s 279476 -800 279588 480 0 FreeSans 1120 90 0 0 la_data_out[43]
port 327 nsew signal tristate
flabel metal2 s 283022 -800 283134 480 0 FreeSans 1120 90 0 0 la_data_out[44]
port 326 nsew signal tristate
flabel metal2 s 286568 -800 286680 480 0 FreeSans 1120 90 0 0 la_data_out[45]
port 325 nsew signal tristate
flabel metal2 s 290114 -800 290226 480 0 FreeSans 1120 90 0 0 la_data_out[46]
port 324 nsew signal tristate
flabel metal2 s 293660 -800 293772 480 0 FreeSans 1120 90 0 0 la_data_out[47]
port 323 nsew signal tristate
flabel metal2 s 297206 -800 297318 480 0 FreeSans 1120 90 0 0 la_data_out[48]
port 322 nsew signal tristate
flabel metal2 s 300752 -800 300864 480 0 FreeSans 1120 90 0 0 la_data_out[49]
port 321 nsew signal tristate
flabel metal2 s 141182 -800 141294 480 0 FreeSans 1120 90 0 0 la_data_out[4]
port 366 nsew signal tristate
flabel metal2 s 304298 -800 304410 480 0 FreeSans 1120 90 0 0 la_data_out[50]
port 320 nsew signal tristate
flabel metal2 s 307844 -800 307956 480 0 FreeSans 1120 90 0 0 la_data_out[51]
port 319 nsew signal tristate
flabel metal2 s 311390 -800 311502 480 0 FreeSans 1120 90 0 0 la_data_out[52]
port 318 nsew signal tristate
flabel metal2 s 314936 -800 315048 480 0 FreeSans 1120 90 0 0 la_data_out[53]
port 317 nsew signal tristate
flabel metal2 s 318482 -800 318594 480 0 FreeSans 1120 90 0 0 la_data_out[54]
port 316 nsew signal tristate
flabel metal2 s 322028 -800 322140 480 0 FreeSans 1120 90 0 0 la_data_out[55]
port 315 nsew signal tristate
flabel metal2 s 325574 -800 325686 480 0 FreeSans 1120 90 0 0 la_data_out[56]
port 314 nsew signal tristate
flabel metal2 s 329120 -800 329232 480 0 FreeSans 1120 90 0 0 la_data_out[57]
port 313 nsew signal tristate
flabel metal2 s 332666 -800 332778 480 0 FreeSans 1120 90 0 0 la_data_out[58]
port 312 nsew signal tristate
flabel metal2 s 336212 -800 336324 480 0 FreeSans 1120 90 0 0 la_data_out[59]
port 311 nsew signal tristate
flabel metal2 s 144728 -800 144840 480 0 FreeSans 1120 90 0 0 la_data_out[5]
port 365 nsew signal tristate
flabel metal2 s 339758 -800 339870 480 0 FreeSans 1120 90 0 0 la_data_out[60]
port 310 nsew signal tristate
flabel metal2 s 343304 -800 343416 480 0 FreeSans 1120 90 0 0 la_data_out[61]
port 309 nsew signal tristate
flabel metal2 s 346850 -800 346962 480 0 FreeSans 1120 90 0 0 la_data_out[62]
port 308 nsew signal tristate
flabel metal2 s 350396 -800 350508 480 0 FreeSans 1120 90 0 0 la_data_out[63]
port 307 nsew signal tristate
flabel metal2 s 353942 -800 354054 480 0 FreeSans 1120 90 0 0 la_data_out[64]
port 306 nsew signal tristate
flabel metal2 s 357488 -800 357600 480 0 FreeSans 1120 90 0 0 la_data_out[65]
port 305 nsew signal tristate
flabel metal2 s 361034 -800 361146 480 0 FreeSans 1120 90 0 0 la_data_out[66]
port 304 nsew signal tristate
flabel metal2 s 364580 -800 364692 480 0 FreeSans 1120 90 0 0 la_data_out[67]
port 303 nsew signal tristate
flabel metal2 s 368126 -800 368238 480 0 FreeSans 1120 90 0 0 la_data_out[68]
port 302 nsew signal tristate
flabel metal2 s 371672 -800 371784 480 0 FreeSans 1120 90 0 0 la_data_out[69]
port 301 nsew signal tristate
flabel metal2 s 148274 -800 148386 480 0 FreeSans 1120 90 0 0 la_data_out[6]
port 364 nsew signal tristate
flabel metal2 s 375218 -800 375330 480 0 FreeSans 1120 90 0 0 la_data_out[70]
port 300 nsew signal tristate
flabel metal2 s 378764 -800 378876 480 0 FreeSans 1120 90 0 0 la_data_out[71]
port 299 nsew signal tristate
flabel metal2 s 382310 -800 382422 480 0 FreeSans 1120 90 0 0 la_data_out[72]
port 298 nsew signal tristate
flabel metal2 s 385856 -800 385968 480 0 FreeSans 1120 90 0 0 la_data_out[73]
port 297 nsew signal tristate
flabel metal2 s 389402 -800 389514 480 0 FreeSans 1120 90 0 0 la_data_out[74]
port 296 nsew signal tristate
flabel metal2 s 392948 -800 393060 480 0 FreeSans 1120 90 0 0 la_data_out[75]
port 295 nsew signal tristate
flabel metal2 s 396494 -800 396606 480 0 FreeSans 1120 90 0 0 la_data_out[76]
port 294 nsew signal tristate
flabel metal2 s 400040 -800 400152 480 0 FreeSans 1120 90 0 0 la_data_out[77]
port 293 nsew signal tristate
flabel metal2 s 403586 -800 403698 480 0 FreeSans 1120 90 0 0 la_data_out[78]
port 292 nsew signal tristate
flabel metal2 s 407132 -800 407244 480 0 FreeSans 1120 90 0 0 la_data_out[79]
port 291 nsew signal tristate
flabel metal2 s 151820 -800 151932 480 0 FreeSans 1120 90 0 0 la_data_out[7]
port 363 nsew signal tristate
flabel metal2 s 410678 -800 410790 480 0 FreeSans 1120 90 0 0 la_data_out[80]
port 290 nsew signal tristate
flabel metal2 s 414224 -800 414336 480 0 FreeSans 1120 90 0 0 la_data_out[81]
port 289 nsew signal tristate
flabel metal2 s 417770 -800 417882 480 0 FreeSans 1120 90 0 0 la_data_out[82]
port 288 nsew signal tristate
flabel metal2 s 421316 -800 421428 480 0 FreeSans 1120 90 0 0 la_data_out[83]
port 287 nsew signal tristate
flabel metal2 s 424862 -800 424974 480 0 FreeSans 1120 90 0 0 la_data_out[84]
port 286 nsew signal tristate
flabel metal2 s 428408 -800 428520 480 0 FreeSans 1120 90 0 0 la_data_out[85]
port 285 nsew signal tristate
flabel metal2 s 431954 -800 432066 480 0 FreeSans 1120 90 0 0 la_data_out[86]
port 284 nsew signal tristate
flabel metal2 s 435500 -800 435612 480 0 FreeSans 1120 90 0 0 la_data_out[87]
port 283 nsew signal tristate
flabel metal2 s 439046 -800 439158 480 0 FreeSans 1120 90 0 0 la_data_out[88]
port 282 nsew signal tristate
flabel metal2 s 442592 -800 442704 480 0 FreeSans 1120 90 0 0 la_data_out[89]
port 281 nsew signal tristate
flabel metal2 s 155366 -800 155478 480 0 FreeSans 1120 90 0 0 la_data_out[8]
port 362 nsew signal tristate
flabel metal2 s 446138 -800 446250 480 0 FreeSans 1120 90 0 0 la_data_out[90]
port 280 nsew signal tristate
flabel metal2 s 449684 -800 449796 480 0 FreeSans 1120 90 0 0 la_data_out[91]
port 279 nsew signal tristate
flabel metal2 s 453230 -800 453342 480 0 FreeSans 1120 90 0 0 la_data_out[92]
port 278 nsew signal tristate
flabel metal2 s 456776 -800 456888 480 0 FreeSans 1120 90 0 0 la_data_out[93]
port 277 nsew signal tristate
flabel metal2 s 460322 -800 460434 480 0 FreeSans 1120 90 0 0 la_data_out[94]
port 276 nsew signal tristate
flabel metal2 s 463868 -800 463980 480 0 FreeSans 1120 90 0 0 la_data_out[95]
port 275 nsew signal tristate
flabel metal2 s 467414 -800 467526 480 0 FreeSans 1120 90 0 0 la_data_out[96]
port 274 nsew signal tristate
flabel metal2 s 470960 -800 471072 480 0 FreeSans 1120 90 0 0 la_data_out[97]
port 273 nsew signal tristate
flabel metal2 s 474506 -800 474618 480 0 FreeSans 1120 90 0 0 la_data_out[98]
port 272 nsew signal tristate
flabel metal2 s 478052 -800 478164 480 0 FreeSans 1120 90 0 0 la_data_out[99]
port 271 nsew signal tristate
flabel metal2 s 158912 -800 159024 480 0 FreeSans 1120 90 0 0 la_data_out[9]
port 361 nsew signal tristate
flabel metal2 s 128180 -800 128292 480 0 FreeSans 1120 90 0 0 la_oenb[0]
port 498 nsew signal input
flabel metal2 s 482780 -800 482892 480 0 FreeSans 1120 90 0 0 la_oenb[100]
port 398 nsew signal input
flabel metal2 s 486326 -800 486438 480 0 FreeSans 1120 90 0 0 la_oenb[101]
port 397 nsew signal input
flabel metal2 s 489872 -800 489984 480 0 FreeSans 1120 90 0 0 la_oenb[102]
port 396 nsew signal input
flabel metal2 s 493418 -800 493530 480 0 FreeSans 1120 90 0 0 la_oenb[103]
port 395 nsew signal input
flabel metal2 s 496964 -800 497076 480 0 FreeSans 1120 90 0 0 la_oenb[104]
port 394 nsew signal input
flabel metal2 s 500510 -800 500622 480 0 FreeSans 1120 90 0 0 la_oenb[105]
port 393 nsew signal input
flabel metal2 s 504056 -800 504168 480 0 FreeSans 1120 90 0 0 la_oenb[106]
port 392 nsew signal input
flabel metal2 s 507602 -800 507714 480 0 FreeSans 1120 90 0 0 la_oenb[107]
port 391 nsew signal input
flabel metal2 s 511148 -800 511260 480 0 FreeSans 1120 90 0 0 la_oenb[108]
port 390 nsew signal input
flabel metal2 s 514694 -800 514806 480 0 FreeSans 1120 90 0 0 la_oenb[109]
port 389 nsew signal input
flabel metal2 s 163640 -800 163752 480 0 FreeSans 1120 90 0 0 la_oenb[10]
port 488 nsew signal input
flabel metal2 s 518240 -800 518352 480 0 FreeSans 1120 90 0 0 la_oenb[110]
port 388 nsew signal input
flabel metal2 s 521786 -800 521898 480 0 FreeSans 1120 90 0 0 la_oenb[111]
port 387 nsew signal input
flabel metal2 s 525332 -800 525444 480 0 FreeSans 1120 90 0 0 la_oenb[112]
port 386 nsew signal input
flabel metal2 s 528878 -800 528990 480 0 FreeSans 1120 90 0 0 la_oenb[113]
port 385 nsew signal input
flabel metal2 s 532424 -800 532536 480 0 FreeSans 1120 90 0 0 la_oenb[114]
port 384 nsew signal input
flabel metal2 s 535970 -800 536082 480 0 FreeSans 1120 90 0 0 la_oenb[115]
port 383 nsew signal input
flabel metal2 s 539516 -800 539628 480 0 FreeSans 1120 90 0 0 la_oenb[116]
port 382 nsew signal input
flabel metal2 s 543062 -800 543174 480 0 FreeSans 1120 90 0 0 la_oenb[117]
port 381 nsew signal input
flabel metal2 s 546608 -800 546720 480 0 FreeSans 1120 90 0 0 la_oenb[118]
port 380 nsew signal input
flabel metal2 s 550154 -800 550266 480 0 FreeSans 1120 90 0 0 la_oenb[119]
port 379 nsew signal input
flabel metal2 s 167186 -800 167298 480 0 FreeSans 1120 90 0 0 la_oenb[11]
port 487 nsew signal input
flabel metal2 s 553700 -800 553812 480 0 FreeSans 1120 90 0 0 la_oenb[120]
port 378 nsew signal input
flabel metal2 s 557246 -800 557358 480 0 FreeSans 1120 90 0 0 la_oenb[121]
port 377 nsew signal input
flabel metal2 s 560792 -800 560904 480 0 FreeSans 1120 90 0 0 la_oenb[122]
port 376 nsew signal input
flabel metal2 s 564338 -800 564450 480 0 FreeSans 1120 90 0 0 la_oenb[123]
port 375 nsew signal input
flabel metal2 s 567884 -800 567996 480 0 FreeSans 1120 90 0 0 la_oenb[124]
port 374 nsew signal input
flabel metal2 s 571430 -800 571542 480 0 FreeSans 1120 90 0 0 la_oenb[125]
port 373 nsew signal input
flabel metal2 s 574976 -800 575088 480 0 FreeSans 1120 90 0 0 la_oenb[126]
port 372 nsew signal input
flabel metal2 s 578522 -800 578634 480 0 FreeSans 1120 90 0 0 la_oenb[127]
port 371 nsew signal input
flabel metal2 s 170732 -800 170844 480 0 FreeSans 1120 90 0 0 la_oenb[12]
port 486 nsew signal input
flabel metal2 s 174278 -800 174390 480 0 FreeSans 1120 90 0 0 la_oenb[13]
port 485 nsew signal input
flabel metal2 s 177824 -800 177936 480 0 FreeSans 1120 90 0 0 la_oenb[14]
port 484 nsew signal input
flabel metal2 s 181370 -800 181482 480 0 FreeSans 1120 90 0 0 la_oenb[15]
port 483 nsew signal input
flabel metal2 s 184916 -800 185028 480 0 FreeSans 1120 90 0 0 la_oenb[16]
port 482 nsew signal input
flabel metal2 s 188462 -800 188574 480 0 FreeSans 1120 90 0 0 la_oenb[17]
port 481 nsew signal input
flabel metal2 s 192008 -800 192120 480 0 FreeSans 1120 90 0 0 la_oenb[18]
port 480 nsew signal input
flabel metal2 s 195554 -800 195666 480 0 FreeSans 1120 90 0 0 la_oenb[19]
port 479 nsew signal input
flabel metal2 s 131726 -800 131838 480 0 FreeSans 1120 90 0 0 la_oenb[1]
port 497 nsew signal input
flabel metal2 s 199100 -800 199212 480 0 FreeSans 1120 90 0 0 la_oenb[20]
port 478 nsew signal input
flabel metal2 s 202646 -800 202758 480 0 FreeSans 1120 90 0 0 la_oenb[21]
port 477 nsew signal input
flabel metal2 s 206192 -800 206304 480 0 FreeSans 1120 90 0 0 la_oenb[22]
port 476 nsew signal input
flabel metal2 s 209738 -800 209850 480 0 FreeSans 1120 90 0 0 la_oenb[23]
port 475 nsew signal input
flabel metal2 s 213284 -800 213396 480 0 FreeSans 1120 90 0 0 la_oenb[24]
port 474 nsew signal input
flabel metal2 s 216830 -800 216942 480 0 FreeSans 1120 90 0 0 la_oenb[25]
port 473 nsew signal input
flabel metal2 s 220376 -800 220488 480 0 FreeSans 1120 90 0 0 la_oenb[26]
port 472 nsew signal input
flabel metal2 s 223922 -800 224034 480 0 FreeSans 1120 90 0 0 la_oenb[27]
port 471 nsew signal input
flabel metal2 s 227468 -800 227580 480 0 FreeSans 1120 90 0 0 la_oenb[28]
port 470 nsew signal input
flabel metal2 s 231014 -800 231126 480 0 FreeSans 1120 90 0 0 la_oenb[29]
port 469 nsew signal input
flabel metal2 s 135272 -800 135384 480 0 FreeSans 1120 90 0 0 la_oenb[2]
port 496 nsew signal input
flabel metal2 s 234560 -800 234672 480 0 FreeSans 1120 90 0 0 la_oenb[30]
port 468 nsew signal input
flabel metal2 s 238106 -800 238218 480 0 FreeSans 1120 90 0 0 la_oenb[31]
port 467 nsew signal input
flabel metal2 s 241652 -800 241764 480 0 FreeSans 1120 90 0 0 la_oenb[32]
port 466 nsew signal input
flabel metal2 s 245198 -800 245310 480 0 FreeSans 1120 90 0 0 la_oenb[33]
port 465 nsew signal input
flabel metal2 s 248744 -800 248856 480 0 FreeSans 1120 90 0 0 la_oenb[34]
port 464 nsew signal input
flabel metal2 s 252290 -800 252402 480 0 FreeSans 1120 90 0 0 la_oenb[35]
port 463 nsew signal input
flabel metal2 s 255836 -800 255948 480 0 FreeSans 1120 90 0 0 la_oenb[36]
port 462 nsew signal input
flabel metal2 s 259382 -800 259494 480 0 FreeSans 1120 90 0 0 la_oenb[37]
port 461 nsew signal input
flabel metal2 s 262928 -800 263040 480 0 FreeSans 1120 90 0 0 la_oenb[38]
port 460 nsew signal input
flabel metal2 s 266474 -800 266586 480 0 FreeSans 1120 90 0 0 la_oenb[39]
port 459 nsew signal input
flabel metal2 s 138818 -800 138930 480 0 FreeSans 1120 90 0 0 la_oenb[3]
port 495 nsew signal input
flabel metal2 s 270020 -800 270132 480 0 FreeSans 1120 90 0 0 la_oenb[40]
port 458 nsew signal input
flabel metal2 s 273566 -800 273678 480 0 FreeSans 1120 90 0 0 la_oenb[41]
port 457 nsew signal input
flabel metal2 s 277112 -800 277224 480 0 FreeSans 1120 90 0 0 la_oenb[42]
port 456 nsew signal input
flabel metal2 s 280658 -800 280770 480 0 FreeSans 1120 90 0 0 la_oenb[43]
port 455 nsew signal input
flabel metal2 s 284204 -800 284316 480 0 FreeSans 1120 90 0 0 la_oenb[44]
port 454 nsew signal input
flabel metal2 s 287750 -800 287862 480 0 FreeSans 1120 90 0 0 la_oenb[45]
port 453 nsew signal input
flabel metal2 s 291296 -800 291408 480 0 FreeSans 1120 90 0 0 la_oenb[46]
port 452 nsew signal input
flabel metal2 s 294842 -800 294954 480 0 FreeSans 1120 90 0 0 la_oenb[47]
port 451 nsew signal input
flabel metal2 s 298388 -800 298500 480 0 FreeSans 1120 90 0 0 la_oenb[48]
port 450 nsew signal input
flabel metal2 s 301934 -800 302046 480 0 FreeSans 1120 90 0 0 la_oenb[49]
port 449 nsew signal input
flabel metal2 s 142364 -800 142476 480 0 FreeSans 1120 90 0 0 la_oenb[4]
port 494 nsew signal input
flabel metal2 s 305480 -800 305592 480 0 FreeSans 1120 90 0 0 la_oenb[50]
port 448 nsew signal input
flabel metal2 s 309026 -800 309138 480 0 FreeSans 1120 90 0 0 la_oenb[51]
port 447 nsew signal input
flabel metal2 s 312572 -800 312684 480 0 FreeSans 1120 90 0 0 la_oenb[52]
port 446 nsew signal input
flabel metal2 s 316118 -800 316230 480 0 FreeSans 1120 90 0 0 la_oenb[53]
port 445 nsew signal input
flabel metal2 s 319664 -800 319776 480 0 FreeSans 1120 90 0 0 la_oenb[54]
port 444 nsew signal input
flabel metal2 s 323210 -800 323322 480 0 FreeSans 1120 90 0 0 la_oenb[55]
port 443 nsew signal input
flabel metal2 s 326756 -800 326868 480 0 FreeSans 1120 90 0 0 la_oenb[56]
port 442 nsew signal input
flabel metal2 s 330302 -800 330414 480 0 FreeSans 1120 90 0 0 la_oenb[57]
port 441 nsew signal input
flabel metal2 s 333848 -800 333960 480 0 FreeSans 1120 90 0 0 la_oenb[58]
port 440 nsew signal input
flabel metal2 s 337394 -800 337506 480 0 FreeSans 1120 90 0 0 la_oenb[59]
port 439 nsew signal input
flabel metal2 s 145910 -800 146022 480 0 FreeSans 1120 90 0 0 la_oenb[5]
port 493 nsew signal input
flabel metal2 s 340940 -800 341052 480 0 FreeSans 1120 90 0 0 la_oenb[60]
port 438 nsew signal input
flabel metal2 s 344486 -800 344598 480 0 FreeSans 1120 90 0 0 la_oenb[61]
port 437 nsew signal input
flabel metal2 s 348032 -800 348144 480 0 FreeSans 1120 90 0 0 la_oenb[62]
port 436 nsew signal input
flabel metal2 s 351578 -800 351690 480 0 FreeSans 1120 90 0 0 la_oenb[63]
port 435 nsew signal input
flabel metal2 s 355124 -800 355236 480 0 FreeSans 1120 90 0 0 la_oenb[64]
port 434 nsew signal input
flabel metal2 s 358670 -800 358782 480 0 FreeSans 1120 90 0 0 la_oenb[65]
port 433 nsew signal input
flabel metal2 s 362216 -800 362328 480 0 FreeSans 1120 90 0 0 la_oenb[66]
port 432 nsew signal input
flabel metal2 s 365762 -800 365874 480 0 FreeSans 1120 90 0 0 la_oenb[67]
port 431 nsew signal input
flabel metal2 s 369308 -800 369420 480 0 FreeSans 1120 90 0 0 la_oenb[68]
port 430 nsew signal input
flabel metal2 s 372854 -800 372966 480 0 FreeSans 1120 90 0 0 la_oenb[69]
port 429 nsew signal input
flabel metal2 s 149456 -800 149568 480 0 FreeSans 1120 90 0 0 la_oenb[6]
port 492 nsew signal input
flabel metal2 s 376400 -800 376512 480 0 FreeSans 1120 90 0 0 la_oenb[70]
port 428 nsew signal input
flabel metal2 s 379946 -800 380058 480 0 FreeSans 1120 90 0 0 la_oenb[71]
port 427 nsew signal input
flabel metal2 s 383492 -800 383604 480 0 FreeSans 1120 90 0 0 la_oenb[72]
port 426 nsew signal input
flabel metal2 s 387038 -800 387150 480 0 FreeSans 1120 90 0 0 la_oenb[73]
port 425 nsew signal input
flabel metal2 s 390584 -800 390696 480 0 FreeSans 1120 90 0 0 la_oenb[74]
port 424 nsew signal input
flabel metal2 s 394130 -800 394242 480 0 FreeSans 1120 90 0 0 la_oenb[75]
port 423 nsew signal input
flabel metal2 s 397676 -800 397788 480 0 FreeSans 1120 90 0 0 la_oenb[76]
port 422 nsew signal input
flabel metal2 s 401222 -800 401334 480 0 FreeSans 1120 90 0 0 la_oenb[77]
port 421 nsew signal input
flabel metal2 s 404768 -800 404880 480 0 FreeSans 1120 90 0 0 la_oenb[78]
port 420 nsew signal input
flabel metal2 s 408314 -800 408426 480 0 FreeSans 1120 90 0 0 la_oenb[79]
port 419 nsew signal input
flabel metal2 s 153002 -800 153114 480 0 FreeSans 1120 90 0 0 la_oenb[7]
port 491 nsew signal input
flabel metal2 s 411860 -800 411972 480 0 FreeSans 1120 90 0 0 la_oenb[80]
port 418 nsew signal input
flabel metal2 s 415406 -800 415518 480 0 FreeSans 1120 90 0 0 la_oenb[81]
port 417 nsew signal input
flabel metal2 s 418952 -800 419064 480 0 FreeSans 1120 90 0 0 la_oenb[82]
port 416 nsew signal input
flabel metal2 s 422498 -800 422610 480 0 FreeSans 1120 90 0 0 la_oenb[83]
port 415 nsew signal input
flabel metal2 s 426044 -800 426156 480 0 FreeSans 1120 90 0 0 la_oenb[84]
port 414 nsew signal input
flabel metal2 s 429590 -800 429702 480 0 FreeSans 1120 90 0 0 la_oenb[85]
port 413 nsew signal input
flabel metal2 s 433136 -800 433248 480 0 FreeSans 1120 90 0 0 la_oenb[86]
port 412 nsew signal input
flabel metal2 s 436682 -800 436794 480 0 FreeSans 1120 90 0 0 la_oenb[87]
port 411 nsew signal input
flabel metal2 s 440228 -800 440340 480 0 FreeSans 1120 90 0 0 la_oenb[88]
port 410 nsew signal input
flabel metal2 s 443774 -800 443886 480 0 FreeSans 1120 90 0 0 la_oenb[89]
port 409 nsew signal input
flabel metal2 s 156548 -800 156660 480 0 FreeSans 1120 90 0 0 la_oenb[8]
port 490 nsew signal input
flabel metal2 s 447320 -800 447432 480 0 FreeSans 1120 90 0 0 la_oenb[90]
port 408 nsew signal input
flabel metal2 s 450866 -800 450978 480 0 FreeSans 1120 90 0 0 la_oenb[91]
port 407 nsew signal input
flabel metal2 s 454412 -800 454524 480 0 FreeSans 1120 90 0 0 la_oenb[92]
port 406 nsew signal input
flabel metal2 s 457958 -800 458070 480 0 FreeSans 1120 90 0 0 la_oenb[93]
port 405 nsew signal input
flabel metal2 s 461504 -800 461616 480 0 FreeSans 1120 90 0 0 la_oenb[94]
port 404 nsew signal input
flabel metal2 s 465050 -800 465162 480 0 FreeSans 1120 90 0 0 la_oenb[95]
port 403 nsew signal input
flabel metal2 s 468596 -800 468708 480 0 FreeSans 1120 90 0 0 la_oenb[96]
port 402 nsew signal input
flabel metal2 s 472142 -800 472254 480 0 FreeSans 1120 90 0 0 la_oenb[97]
port 401 nsew signal input
flabel metal2 s 475688 -800 475800 480 0 FreeSans 1120 90 0 0 la_oenb[98]
port 400 nsew signal input
flabel metal2 s 479234 -800 479346 480 0 FreeSans 1120 90 0 0 la_oenb[99]
port 399 nsew signal input
flabel metal2 s 160094 -800 160206 480 0 FreeSans 1120 90 0 0 la_oenb[9]
port 489 nsew signal input
flabel metal2 s 579704 -800 579816 480 0 FreeSans 1120 90 0 0 user_clock2
port 660 nsew signal input
flabel metal2 s 580886 -800 580998 480 0 FreeSans 1120 90 0 0 user_irq[0]
port 663 nsew signal tristate
flabel metal2 s 582068 -800 582180 480 0 FreeSans 1120 90 0 0 user_irq[1]
port 662 nsew signal tristate
flabel metal2 s 583250 -800 583362 480 0 FreeSans 1120 90 0 0 user_irq[2]
port 661 nsew signal tristate
flabel metal3 s 582340 639784 584800 644584 0 FreeSans 1120 0 0 0 vccd1
port 5 nsew signal bidirectional
flabel metal3 s 582340 629784 584800 634584 0 FreeSans 1120 0 0 0 vccd1
port 5 nsew signal bidirectional
flabel metal3 s 582340 540562 584800 545362 0 FreeSans 1120 0 0 0 vdda1
port 1 nsew signal bidirectional
flabel metal3 s 582340 550562 584800 555362 0 FreeSans 1120 0 0 0 vdda1
port 1 nsew signal bidirectional
flabel metal3 s 582340 235230 584800 240030 0 FreeSans 1120 0 0 0 vdda1
port 1 nsew signal bidirectional
flabel metal3 s 582340 225230 584800 230030 0 FreeSans 1120 0 0 0 vdda1
port 1 nsew signal bidirectional
flabel metal3 s 0 204888 1660 209688 0 FreeSans 1120 0 0 0 vdda2
port 2 nsew signal bidirectional
flabel metal3 s 0 214888 1660 219688 0 FreeSans 1120 0 0 0 vdda2
port 2 nsew signal bidirectional
flabel metal3 s 520594 702340 525394 704800 0 FreeSans 1920 180 0 0 vssa1
port 3 nsew signal bidirectional
flabel metal3 s 510594 702340 515394 704800 0 FreeSans 1920 180 0 0 vssa1
port 3 nsew signal bidirectional
flabel metal3 s 582340 146830 584800 151630 0 FreeSans 1120 0 0 0 vssa1
port 3 nsew signal bidirectional
flabel metal3 s 582340 136830 584800 141630 0 FreeSans 1120 0 0 0 vssa1
port 3 nsew signal bidirectional
flabel metal3 s 582340 191430 584800 196230 0 FreeSans 1120 0 0 0 vssd1
port 7 nsew signal bidirectional
flabel metal3 s 582340 181430 584800 186230 0 FreeSans 1120 0 0 0 vssd1
port 7 nsew signal bidirectional
flabel metal3 s 0 172888 1660 177688 0 FreeSans 1120 0 0 0 vssd2
port 8 nsew signal bidirectional
flabel metal3 s 0 162888 1660 167688 0 FreeSans 1120 0 0 0 vssd2
port 8 nsew signal bidirectional
flabel metal2 s 524 -800 636 480 0 FreeSans 1120 90 0 0 wb_clk_i
port 9 nsew signal input
flabel metal2 s 1706 -800 1818 480 0 FreeSans 1120 90 0 0 wb_rst_i
port 10 nsew signal input
flabel metal2 s 2888 -800 3000 480 0 FreeSans 1120 90 0 0 wbs_ack_o
port 82 nsew signal tristate
flabel metal2 s 7616 -800 7728 480 0 FreeSans 1120 90 0 0 wbs_adr_i[0]
port 81 nsew signal input
flabel metal2 s 47804 -800 47916 480 0 FreeSans 1120 90 0 0 wbs_adr_i[10]
port 71 nsew signal input
flabel metal2 s 51350 -800 51462 480 0 FreeSans 1120 90 0 0 wbs_adr_i[11]
port 70 nsew signal input
flabel metal2 s 54896 -800 55008 480 0 FreeSans 1120 90 0 0 wbs_adr_i[12]
port 69 nsew signal input
flabel metal2 s 58442 -800 58554 480 0 FreeSans 1120 90 0 0 wbs_adr_i[13]
port 68 nsew signal input
flabel metal2 s 61988 -800 62100 480 0 FreeSans 1120 90 0 0 wbs_adr_i[14]
port 67 nsew signal input
flabel metal2 s 65534 -800 65646 480 0 FreeSans 1120 90 0 0 wbs_adr_i[15]
port 66 nsew signal input
flabel metal2 s 69080 -800 69192 480 0 FreeSans 1120 90 0 0 wbs_adr_i[16]
port 65 nsew signal input
flabel metal2 s 72626 -800 72738 480 0 FreeSans 1120 90 0 0 wbs_adr_i[17]
port 64 nsew signal input
flabel metal2 s 76172 -800 76284 480 0 FreeSans 1120 90 0 0 wbs_adr_i[18]
port 63 nsew signal input
flabel metal2 s 79718 -800 79830 480 0 FreeSans 1120 90 0 0 wbs_adr_i[19]
port 62 nsew signal input
flabel metal2 s 12344 -800 12456 480 0 FreeSans 1120 90 0 0 wbs_adr_i[1]
port 80 nsew signal input
flabel metal2 s 83264 -800 83376 480 0 FreeSans 1120 90 0 0 wbs_adr_i[20]
port 61 nsew signal input
flabel metal2 s 86810 -800 86922 480 0 FreeSans 1120 90 0 0 wbs_adr_i[21]
port 60 nsew signal input
flabel metal2 s 90356 -800 90468 480 0 FreeSans 1120 90 0 0 wbs_adr_i[22]
port 59 nsew signal input
flabel metal2 s 93902 -800 94014 480 0 FreeSans 1120 90 0 0 wbs_adr_i[23]
port 58 nsew signal input
flabel metal2 s 97448 -800 97560 480 0 FreeSans 1120 90 0 0 wbs_adr_i[24]
port 57 nsew signal input
flabel metal2 s 100994 -800 101106 480 0 FreeSans 1120 90 0 0 wbs_adr_i[25]
port 56 nsew signal input
flabel metal2 s 104540 -800 104652 480 0 FreeSans 1120 90 0 0 wbs_adr_i[26]
port 55 nsew signal input
flabel metal2 s 108086 -800 108198 480 0 FreeSans 1120 90 0 0 wbs_adr_i[27]
port 54 nsew signal input
flabel metal2 s 111632 -800 111744 480 0 FreeSans 1120 90 0 0 wbs_adr_i[28]
port 53 nsew signal input
flabel metal2 s 115178 -800 115290 480 0 FreeSans 1120 90 0 0 wbs_adr_i[29]
port 52 nsew signal input
flabel metal2 s 17072 -800 17184 480 0 FreeSans 1120 90 0 0 wbs_adr_i[2]
port 79 nsew signal input
flabel metal2 s 118724 -800 118836 480 0 FreeSans 1120 90 0 0 wbs_adr_i[30]
port 51 nsew signal input
flabel metal2 s 122270 -800 122382 480 0 FreeSans 1120 90 0 0 wbs_adr_i[31]
port 50 nsew signal input
flabel metal2 s 21800 -800 21912 480 0 FreeSans 1120 90 0 0 wbs_adr_i[3]
port 78 nsew signal input
flabel metal2 s 26528 -800 26640 480 0 FreeSans 1120 90 0 0 wbs_adr_i[4]
port 77 nsew signal input
flabel metal2 s 30074 -800 30186 480 0 FreeSans 1120 90 0 0 wbs_adr_i[5]
port 76 nsew signal input
flabel metal2 s 33620 -800 33732 480 0 FreeSans 1120 90 0 0 wbs_adr_i[6]
port 75 nsew signal input
flabel metal2 s 37166 -800 37278 480 0 FreeSans 1120 90 0 0 wbs_adr_i[7]
port 74 nsew signal input
flabel metal2 s 40712 -800 40824 480 0 FreeSans 1120 90 0 0 wbs_adr_i[8]
port 73 nsew signal input
flabel metal2 s 44258 -800 44370 480 0 FreeSans 1120 90 0 0 wbs_adr_i[9]
port 72 nsew signal input
flabel metal2 s 4070 -800 4182 480 0 FreeSans 1120 90 0 0 wbs_cyc_i
port 12 nsew signal input
flabel metal2 s 8798 -800 8910 480 0 FreeSans 1120 90 0 0 wbs_dat_i[0]
port 49 nsew signal input
flabel metal2 s 48986 -800 49098 480 0 FreeSans 1120 90 0 0 wbs_dat_i[10]
port 39 nsew signal input
flabel metal2 s 52532 -800 52644 480 0 FreeSans 1120 90 0 0 wbs_dat_i[11]
port 38 nsew signal input
flabel metal2 s 56078 -800 56190 480 0 FreeSans 1120 90 0 0 wbs_dat_i[12]
port 37 nsew signal input
flabel metal2 s 59624 -800 59736 480 0 FreeSans 1120 90 0 0 wbs_dat_i[13]
port 36 nsew signal input
flabel metal2 s 63170 -800 63282 480 0 FreeSans 1120 90 0 0 wbs_dat_i[14]
port 35 nsew signal input
flabel metal2 s 66716 -800 66828 480 0 FreeSans 1120 90 0 0 wbs_dat_i[15]
port 34 nsew signal input
flabel metal2 s 70262 -800 70374 480 0 FreeSans 1120 90 0 0 wbs_dat_i[16]
port 33 nsew signal input
flabel metal2 s 73808 -800 73920 480 0 FreeSans 1120 90 0 0 wbs_dat_i[17]
port 32 nsew signal input
flabel metal2 s 77354 -800 77466 480 0 FreeSans 1120 90 0 0 wbs_dat_i[18]
port 31 nsew signal input
flabel metal2 s 80900 -800 81012 480 0 FreeSans 1120 90 0 0 wbs_dat_i[19]
port 30 nsew signal input
flabel metal2 s 13526 -800 13638 480 0 FreeSans 1120 90 0 0 wbs_dat_i[1]
port 48 nsew signal input
flabel metal2 s 84446 -800 84558 480 0 FreeSans 1120 90 0 0 wbs_dat_i[20]
port 29 nsew signal input
flabel metal2 s 87992 -800 88104 480 0 FreeSans 1120 90 0 0 wbs_dat_i[21]
port 28 nsew signal input
flabel metal2 s 91538 -800 91650 480 0 FreeSans 1120 90 0 0 wbs_dat_i[22]
port 27 nsew signal input
flabel metal2 s 95084 -800 95196 480 0 FreeSans 1120 90 0 0 wbs_dat_i[23]
port 26 nsew signal input
flabel metal2 s 98630 -800 98742 480 0 FreeSans 1120 90 0 0 wbs_dat_i[24]
port 25 nsew signal input
flabel metal2 s 102176 -800 102288 480 0 FreeSans 1120 90 0 0 wbs_dat_i[25]
port 24 nsew signal input
flabel metal2 s 105722 -800 105834 480 0 FreeSans 1120 90 0 0 wbs_dat_i[26]
port 23 nsew signal input
flabel metal2 s 109268 -800 109380 480 0 FreeSans 1120 90 0 0 wbs_dat_i[27]
port 22 nsew signal input
flabel metal2 s 112814 -800 112926 480 0 FreeSans 1120 90 0 0 wbs_dat_i[28]
port 21 nsew signal input
flabel metal2 s 116360 -800 116472 480 0 FreeSans 1120 90 0 0 wbs_dat_i[29]
port 20 nsew signal input
flabel metal2 s 18254 -800 18366 480 0 FreeSans 1120 90 0 0 wbs_dat_i[2]
port 47 nsew signal input
flabel metal2 s 119906 -800 120018 480 0 FreeSans 1120 90 0 0 wbs_dat_i[30]
port 19 nsew signal input
flabel metal2 s 123452 -800 123564 480 0 FreeSans 1120 90 0 0 wbs_dat_i[31]
port 18 nsew signal input
flabel metal2 s 22982 -800 23094 480 0 FreeSans 1120 90 0 0 wbs_dat_i[3]
port 46 nsew signal input
flabel metal2 s 27710 -800 27822 480 0 FreeSans 1120 90 0 0 wbs_dat_i[4]
port 45 nsew signal input
flabel metal2 s 31256 -800 31368 480 0 FreeSans 1120 90 0 0 wbs_dat_i[5]
port 44 nsew signal input
flabel metal2 s 34802 -800 34914 480 0 FreeSans 1120 90 0 0 wbs_dat_i[6]
port 43 nsew signal input
flabel metal2 s 38348 -800 38460 480 0 FreeSans 1120 90 0 0 wbs_dat_i[7]
port 42 nsew signal input
flabel metal2 s 41894 -800 42006 480 0 FreeSans 1120 90 0 0 wbs_dat_i[8]
port 41 nsew signal input
flabel metal2 s 45440 -800 45552 480 0 FreeSans 1120 90 0 0 wbs_dat_i[9]
port 40 nsew signal input
flabel metal2 s 9980 -800 10092 480 0 FreeSans 1120 90 0 0 wbs_dat_o[0]
port 114 nsew signal tristate
flabel metal2 s 50168 -800 50280 480 0 FreeSans 1120 90 0 0 wbs_dat_o[10]
port 104 nsew signal tristate
flabel metal2 s 53714 -800 53826 480 0 FreeSans 1120 90 0 0 wbs_dat_o[11]
port 103 nsew signal tristate
flabel metal2 s 57260 -800 57372 480 0 FreeSans 1120 90 0 0 wbs_dat_o[12]
port 102 nsew signal tristate
flabel metal2 s 60806 -800 60918 480 0 FreeSans 1120 90 0 0 wbs_dat_o[13]
port 101 nsew signal tristate
flabel metal2 s 64352 -800 64464 480 0 FreeSans 1120 90 0 0 wbs_dat_o[14]
port 100 nsew signal tristate
flabel metal2 s 67898 -800 68010 480 0 FreeSans 1120 90 0 0 wbs_dat_o[15]
port 99 nsew signal tristate
flabel metal2 s 71444 -800 71556 480 0 FreeSans 1120 90 0 0 wbs_dat_o[16]
port 98 nsew signal tristate
flabel metal2 s 74990 -800 75102 480 0 FreeSans 1120 90 0 0 wbs_dat_o[17]
port 97 nsew signal tristate
flabel metal2 s 78536 -800 78648 480 0 FreeSans 1120 90 0 0 wbs_dat_o[18]
port 96 nsew signal tristate
flabel metal2 s 82082 -800 82194 480 0 FreeSans 1120 90 0 0 wbs_dat_o[19]
port 95 nsew signal tristate
flabel metal2 s 14708 -800 14820 480 0 FreeSans 1120 90 0 0 wbs_dat_o[1]
port 113 nsew signal tristate
flabel metal2 s 85628 -800 85740 480 0 FreeSans 1120 90 0 0 wbs_dat_o[20]
port 94 nsew signal tristate
flabel metal2 s 89174 -800 89286 480 0 FreeSans 1120 90 0 0 wbs_dat_o[21]
port 93 nsew signal tristate
flabel metal2 s 92720 -800 92832 480 0 FreeSans 1120 90 0 0 wbs_dat_o[22]
port 92 nsew signal tristate
flabel metal2 s 96266 -800 96378 480 0 FreeSans 1120 90 0 0 wbs_dat_o[23]
port 91 nsew signal tristate
flabel metal2 s 99812 -800 99924 480 0 FreeSans 1120 90 0 0 wbs_dat_o[24]
port 90 nsew signal tristate
flabel metal2 s 103358 -800 103470 480 0 FreeSans 1120 90 0 0 wbs_dat_o[25]
port 89 nsew signal tristate
flabel metal2 s 106904 -800 107016 480 0 FreeSans 1120 90 0 0 wbs_dat_o[26]
port 88 nsew signal tristate
flabel metal2 s 110450 -800 110562 480 0 FreeSans 1120 90 0 0 wbs_dat_o[27]
port 87 nsew signal tristate
flabel metal2 s 113996 -800 114108 480 0 FreeSans 1120 90 0 0 wbs_dat_o[28]
port 86 nsew signal tristate
flabel metal2 s 117542 -800 117654 480 0 FreeSans 1120 90 0 0 wbs_dat_o[29]
port 85 nsew signal tristate
flabel metal2 s 19436 -800 19548 480 0 FreeSans 1120 90 0 0 wbs_dat_o[2]
port 112 nsew signal tristate
flabel metal2 s 121088 -800 121200 480 0 FreeSans 1120 90 0 0 wbs_dat_o[30]
port 84 nsew signal tristate
flabel metal2 s 124634 -800 124746 480 0 FreeSans 1120 90 0 0 wbs_dat_o[31]
port 83 nsew signal tristate
flabel metal2 s 24164 -800 24276 480 0 FreeSans 1120 90 0 0 wbs_dat_o[3]
port 111 nsew signal tristate
flabel metal2 s 28892 -800 29004 480 0 FreeSans 1120 90 0 0 wbs_dat_o[4]
port 110 nsew signal tristate
flabel metal2 s 32438 -800 32550 480 0 FreeSans 1120 90 0 0 wbs_dat_o[5]
port 109 nsew signal tristate
flabel metal2 s 35984 -800 36096 480 0 FreeSans 1120 90 0 0 wbs_dat_o[6]
port 108 nsew signal tristate
flabel metal2 s 39530 -800 39642 480 0 FreeSans 1120 90 0 0 wbs_dat_o[7]
port 107 nsew signal tristate
flabel metal2 s 43076 -800 43188 480 0 FreeSans 1120 90 0 0 wbs_dat_o[8]
port 106 nsew signal tristate
flabel metal2 s 46622 -800 46734 480 0 FreeSans 1120 90 0 0 wbs_dat_o[9]
port 105 nsew signal tristate
flabel metal2 s 11162 -800 11274 480 0 FreeSans 1120 90 0 0 wbs_sel_i[0]
port 17 nsew signal input
flabel metal2 s 15890 -800 16002 480 0 FreeSans 1120 90 0 0 wbs_sel_i[1]
port 16 nsew signal input
flabel metal2 s 20618 -800 20730 480 0 FreeSans 1120 90 0 0 wbs_sel_i[2]
port 15 nsew signal input
flabel metal2 s 25346 -800 25458 480 0 FreeSans 1120 90 0 0 wbs_sel_i[3]
port 14 nsew signal input
flabel metal2 s 5252 -800 5364 480 0 FreeSans 1120 90 0 0 wbs_stb_i
port 11 nsew signal input
flabel metal2 s 6434 -800 6546 480 0 FreeSans 1120 90 0 0 wbs_we_i
port 13 nsew signal input
rlabel metal4 41592 695986 41736 696166 1 OTA_GM_0/Vout
rlabel metal1 41376 693876 41602 694036 1 OTA_GM_0/Vmid
flabel metal3 s 0 549442 1660 554242 0 FreeSans 1120 0 0 0 vssa2
port 4 nsew signal bidirectional
flabel metal3 s 0 559442 1660 564242 0 FreeSans 1120 0 0 0 vssa2
port 4 nsew signal bidirectional
flabel metal3 s 0 633842 1660 638642 0 FreeSans 1120 0 0 0 vccd2
port 6 nsew signal bidirectional
flabel metal3 s 0 643842 1660 648642 0 FreeSans 1120 0 0 0 vccd2
port 6 nsew signal bidirectional
flabel metal3 s -800 506802 480 506914 0 FreeSans 1120 0 0 0 io_out[14]
port 565 nsew signal tristate
flabel metal3 s -800 505620 480 505732 0 FreeSans 1120 0 0 0 io_oeb[14]
port 592 nsew signal tristate
flabel metal3 s -800 509166 480 509278 0 FreeSans 1120 0 0 0 io_in_3v3[14]
port 538 nsew signal input
flabel metal3 s -800 507984 480 508096 0 FreeSans 1120 0 0 0 io_in[14]
port 511 nsew signal input
flabel metal3 s 170894 702300 173094 704800 0 FreeSans 1920 180 0 0 io_clamp_low[2]
port 657 nsew signal bidirectional
flabel metal3 s 222594 702300 224794 704800 0 FreeSans 1920 180 0 0 io_clamp_low[1]
port 658 nsew signal bidirectional
flabel metal3 s 324294 702300 326494 704800 0 FreeSans 1920 180 0 0 io_clamp_low[0]
port 659 nsew signal bidirectional
flabel metal3 s 173394 702300 175594 704800 0 FreeSans 1920 180 0 0 io_clamp_high[2]
port 654 nsew signal bidirectional
flabel metal3 s 225094 702300 227294 704800 0 FreeSans 1920 180 0 0 io_clamp_high[1]
port 655 nsew signal bidirectional
flabel metal3 s 326794 702300 328994 704800 0 FreeSans 1920 180 0 0 io_clamp_high[0]
port 656 nsew signal bidirectional
flabel metal4 s 165594 702300 170594 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 647 nsew signal bidirectional
flabel metal3 s 165594 702300 170594 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 647 nsew signal bidirectional
flabel metal4 s 217294 702300 222294 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 648 nsew signal bidirectional
flabel metal3 s 217294 702300 222294 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 648 nsew signal bidirectional
flabel metal4 s 318994 702300 323994 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 649 nsew signal bidirectional
flabel metal3 s 318994 702300 323994 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 649 nsew signal bidirectional
flabel metal3 s 16194 702300 21194 704800 0 FreeSans 1920 180 0 0 io_analog[9]
port 644 nsew signal bidirectional
flabel metal3 s 68194 702300 73194 704800 0 FreeSans 1920 180 0 0 io_analog[8]
port 645 nsew signal bidirectional
flabel metal3 s 120194 702300 125194 704800 0 FreeSans 1920 180 0 0 io_analog[7]
port 646 nsew signal bidirectional
flabel metal4 s 175894 702300 180894 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 647 nsew signal bidirectional
flabel metal3 s 175894 702300 180894 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 647 nsew signal bidirectional
flabel metal4 s 227594 702300 232594 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 648 nsew signal bidirectional
flabel metal3 s 227594 702300 232594 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 648 nsew signal bidirectional
flabel metal4 s 329294 702300 334294 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 649 nsew signal bidirectional
flabel metal3 s 329294 702300 334294 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 649 nsew signal bidirectional
flabel metal3 s 0 680242 1700 685242 0 FreeSans 1120 0 0 0 io_analog[10]
port 643 nsew signal bidirectional
flabel metal3 s -800 510348 480 510460 0 FreeSans 1120 0 0 0 gpio_noesd[7]
port 635 nsew signal bidirectional
flabel metal3 s -800 511530 480 511642 0 FreeSans 1120 0 0 0 gpio_analog[7]
port 617 nsew signal bidirectional
<< end >>
