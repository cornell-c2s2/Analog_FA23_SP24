magic
tech sky130A
magscale 1 2
timestamp 1713626893
<< nwell >>
rect -100 -1800 1790 1140
<< pwell >>
rect -2636 -6210 -2344 -5870
rect 4064 -6210 4356 -5870
rect -2636 -7930 -2344 -7590
rect 4064 -7930 4356 -7590
rect -2636 -9650 -2344 -9310
rect 4064 -9650 4356 -9310
rect -2636 -11130 -2344 -10790
rect 4064 -11130 4356 -10790
rect -2636 -12850 -2344 -12510
rect 4064 -12850 4356 -12510
rect -2636 -14450 -2344 -14110
rect 4064 -14450 4356 -14110
rect -2636 -16170 -2344 -15830
rect 4064 -16170 4356 -15830
rect -2636 -17770 -2344 -17430
rect 4064 -17770 4356 -17430
rect -2636 -19490 -2344 -19150
rect 4064 -19490 4356 -19150
<< psubdiff >>
rect -2610 -5921 -2370 -5896
rect -2610 -6159 -2609 -5921
rect -2371 -6159 -2370 -5921
rect -2610 -6184 -2370 -6159
rect 4090 -5921 4330 -5896
rect 4090 -6159 4091 -5921
rect 4329 -6159 4330 -5921
rect 4090 -6184 4330 -6159
rect -2610 -7641 -2370 -7616
rect -2610 -7879 -2609 -7641
rect -2371 -7879 -2370 -7641
rect -2610 -7904 -2370 -7879
rect 4090 -7641 4330 -7616
rect 4090 -7879 4091 -7641
rect 4329 -7879 4330 -7641
rect 4090 -7904 4330 -7879
rect -2610 -9361 -2370 -9336
rect -2610 -9599 -2609 -9361
rect -2371 -9599 -2370 -9361
rect -2610 -9624 -2370 -9599
rect 4090 -9361 4330 -9336
rect 4090 -9599 4091 -9361
rect 4329 -9599 4330 -9361
rect 4090 -9624 4330 -9599
rect -2610 -10841 -2370 -10816
rect -2610 -11079 -2609 -10841
rect -2371 -11079 -2370 -10841
rect -2610 -11104 -2370 -11079
rect 4090 -10841 4330 -10816
rect 4090 -11079 4091 -10841
rect 4329 -11079 4330 -10841
rect 4090 -11104 4330 -11079
rect -2610 -12561 -2370 -12536
rect -2610 -12799 -2609 -12561
rect -2371 -12799 -2370 -12561
rect -2610 -12824 -2370 -12799
rect 4090 -12561 4330 -12536
rect 4090 -12799 4091 -12561
rect 4329 -12799 4330 -12561
rect 4090 -12824 4330 -12799
rect -2610 -14161 -2370 -14136
rect -2610 -14399 -2609 -14161
rect -2371 -14399 -2370 -14161
rect -2610 -14424 -2370 -14399
rect 4090 -14161 4330 -14136
rect 4090 -14399 4091 -14161
rect 4329 -14399 4330 -14161
rect 4090 -14424 4330 -14399
rect -2610 -15881 -2370 -15856
rect -2610 -16119 -2609 -15881
rect -2371 -16119 -2370 -15881
rect -2610 -16144 -2370 -16119
rect 4090 -15881 4330 -15856
rect 4090 -16119 4091 -15881
rect 4329 -16119 4330 -15881
rect 4090 -16144 4330 -16119
rect -2610 -17481 -2370 -17456
rect -2610 -17719 -2609 -17481
rect -2371 -17719 -2370 -17481
rect -2610 -17744 -2370 -17719
rect 4090 -17481 4330 -17456
rect 4090 -17719 4091 -17481
rect 4329 -17719 4330 -17481
rect 4090 -17744 4330 -17719
rect -2610 -19201 -2370 -19176
rect -2610 -19439 -2609 -19201
rect -2371 -19439 -2370 -19201
rect -2610 -19464 -2370 -19439
rect 4090 -19201 4330 -19176
rect 4090 -19439 4091 -19201
rect 4329 -19439 4330 -19201
rect 4090 -19464 4330 -19439
<< psubdiffcont >>
rect -2609 -6159 -2371 -5921
rect 4091 -6159 4329 -5921
rect -2609 -7879 -2371 -7641
rect 4091 -7879 4329 -7641
rect -2609 -9599 -2371 -9361
rect 4091 -9599 4329 -9361
rect -2609 -11079 -2371 -10841
rect 4091 -11079 4329 -10841
rect -2609 -12799 -2371 -12561
rect 4091 -12799 4329 -12561
rect -2609 -14399 -2371 -14161
rect 4091 -14399 4329 -14161
rect -2609 -16119 -2371 -15881
rect 4091 -16119 4329 -15881
rect -2609 -17719 -2371 -17481
rect 4091 -17719 4329 -17481
rect -2609 -19439 -2371 -19201
rect 4091 -19439 4329 -19201
<< locali >>
rect -70 504 -30 530
rect -70 470 -67 504
rect -33 470 -30 504
rect -70 432 -30 470
rect -70 398 -67 432
rect -33 398 -30 432
rect -70 360 -30 398
rect -70 326 -67 360
rect -33 326 -30 360
rect -70 300 -30 326
rect 1710 504 1750 530
rect 1710 470 1713 504
rect 1747 470 1750 504
rect 1710 432 1750 470
rect 1710 398 1713 432
rect 1747 398 1750 432
rect 1710 360 1750 398
rect 1710 326 1713 360
rect 1747 326 1750 360
rect 1710 300 1750 326
rect -70 -1006 -30 -980
rect -70 -1040 -67 -1006
rect -33 -1040 -30 -1006
rect -70 -1078 -30 -1040
rect -70 -1112 -67 -1078
rect -33 -1112 -30 -1078
rect -70 -1150 -30 -1112
rect -70 -1184 -67 -1150
rect -33 -1184 -30 -1150
rect -70 -1210 -30 -1184
rect 1710 -1006 1750 -980
rect 1710 -1040 1713 -1006
rect 1747 -1040 1750 -1006
rect 1710 -1078 1750 -1040
rect 1710 -1112 1713 -1078
rect 1747 -1112 1750 -1078
rect 1710 -1150 1750 -1112
rect 1710 -1184 1713 -1150
rect 1747 -1184 1750 -1150
rect 1710 -1210 1750 -1184
rect 530 -2346 570 -2320
rect 530 -2380 533 -2346
rect 567 -2380 570 -2346
rect 530 -2418 570 -2380
rect 530 -2452 533 -2418
rect 567 -2452 570 -2418
rect 530 -2490 570 -2452
rect 530 -2524 533 -2490
rect 567 -2524 570 -2490
rect 530 -2550 570 -2524
rect 1080 -2346 1120 -2320
rect 1080 -2380 1083 -2346
rect 1117 -2380 1120 -2346
rect 1080 -2418 1120 -2380
rect 1080 -2452 1083 -2418
rect 1117 -2452 1120 -2418
rect 1080 -2490 1120 -2452
rect 1080 -2524 1083 -2490
rect 1117 -2524 1120 -2490
rect 1080 -2550 1120 -2524
rect 150 -3298 240 -3270
rect 150 -3332 178 -3298
rect 212 -3332 240 -3298
rect 150 -3360 240 -3332
rect 1410 -3293 1490 -3270
rect 1410 -3327 1433 -3293
rect 1467 -3327 1490 -3293
rect 1410 -3350 1490 -3327
rect 690 -3583 930 -3580
rect 690 -3617 721 -3583
rect 755 -3617 793 -3583
rect 827 -3617 865 -3583
rect 899 -3617 930 -3583
rect 690 -3620 930 -3617
rect 690 -3763 930 -3760
rect 690 -3797 721 -3763
rect 755 -3797 793 -3763
rect 827 -3797 865 -3763
rect 899 -3797 930 -3763
rect 690 -3800 930 -3797
rect 690 -5083 930 -5080
rect 690 -5117 721 -5083
rect 755 -5117 793 -5083
rect 827 -5117 865 -5083
rect 899 -5117 930 -5083
rect 690 -5120 930 -5117
rect -2610 -5921 -2370 -5904
rect -2610 -6159 -2609 -5921
rect -2371 -6159 -2370 -5921
rect -2610 -6176 -2370 -6159
rect 4090 -5921 4330 -5904
rect 4090 -6159 4091 -5921
rect 4329 -6159 4330 -5921
rect 4090 -6176 4330 -6159
rect -2610 -7641 -2370 -7624
rect -2610 -7879 -2609 -7641
rect -2371 -7879 -2370 -7641
rect -2610 -7896 -2370 -7879
rect 4090 -7641 4330 -7624
rect 4090 -7879 4091 -7641
rect 4329 -7879 4330 -7641
rect 4090 -7896 4330 -7879
rect -2610 -9361 -2370 -9344
rect -2610 -9599 -2609 -9361
rect -2371 -9599 -2370 -9361
rect -2610 -9616 -2370 -9599
rect 4090 -9361 4330 -9344
rect 4090 -9599 4091 -9361
rect 4329 -9599 4330 -9361
rect 4090 -9616 4330 -9599
rect -2610 -10841 -2370 -10824
rect -2610 -11079 -2609 -10841
rect -2371 -11079 -2370 -10841
rect -2610 -11096 -2370 -11079
rect 4090 -10841 4330 -10824
rect 4090 -11079 4091 -10841
rect 4329 -11079 4330 -10841
rect 4090 -11096 4330 -11079
rect -2610 -12561 -2370 -12544
rect -2610 -12799 -2609 -12561
rect -2371 -12799 -2370 -12561
rect -2610 -12816 -2370 -12799
rect 4090 -12561 4330 -12544
rect 4090 -12799 4091 -12561
rect 4329 -12799 4330 -12561
rect 4090 -12816 4330 -12799
rect -2610 -14161 -2370 -14144
rect -2610 -14399 -2609 -14161
rect -2371 -14399 -2370 -14161
rect -2610 -14416 -2370 -14399
rect 4090 -14161 4330 -14144
rect 4090 -14399 4091 -14161
rect 4329 -14399 4330 -14161
rect 4090 -14416 4330 -14399
rect -2610 -15881 -2370 -15864
rect -2610 -16119 -2609 -15881
rect -2371 -16119 -2370 -15881
rect -2610 -16136 -2370 -16119
rect 4090 -15881 4330 -15864
rect 4090 -16119 4091 -15881
rect 4329 -16119 4330 -15881
rect 4090 -16136 4330 -16119
rect -2610 -17481 -2370 -17464
rect -2610 -17719 -2609 -17481
rect -2371 -17719 -2370 -17481
rect -2610 -17736 -2370 -17719
rect 4090 -17481 4330 -17464
rect 4090 -17719 4091 -17481
rect 4329 -17719 4330 -17481
rect 4090 -17736 4330 -17719
rect -2610 -19201 -2370 -19184
rect -2610 -19439 -2609 -19201
rect -2371 -19439 -2370 -19201
rect -2610 -19456 -2370 -19439
rect 4090 -19201 4330 -19184
rect 4090 -19439 4091 -19201
rect 4329 -19439 4330 -19201
rect 4090 -19456 4330 -19439
<< viali >>
rect -67 470 -33 504
rect -67 398 -33 432
rect -67 326 -33 360
rect 1713 470 1747 504
rect 1713 398 1747 432
rect 1713 326 1747 360
rect -67 -1040 -33 -1006
rect -67 -1112 -33 -1078
rect -67 -1184 -33 -1150
rect 1713 -1040 1747 -1006
rect 1713 -1112 1747 -1078
rect 1713 -1184 1747 -1150
rect 533 -2380 567 -2346
rect 533 -2452 567 -2418
rect 533 -2524 567 -2490
rect 1083 -2380 1117 -2346
rect 1083 -2452 1117 -2418
rect 1083 -2524 1117 -2490
rect 178 -3332 212 -3298
rect 1433 -3327 1467 -3293
rect 721 -3617 755 -3583
rect 793 -3617 827 -3583
rect 865 -3617 899 -3583
rect 721 -3797 755 -3763
rect 793 -3797 827 -3763
rect 865 -3797 899 -3763
rect 721 -5117 755 -5083
rect 793 -5117 827 -5083
rect 865 -5117 899 -5083
rect -2579 -6129 -2401 -5951
rect 4121 -6129 4299 -5951
rect -2579 -7849 -2401 -7671
rect 4121 -7849 4299 -7671
rect -2579 -9569 -2401 -9391
rect 4121 -9569 4299 -9391
rect -2579 -11049 -2401 -10871
rect 4121 -11049 4299 -10871
rect -2579 -12769 -2401 -12591
rect 4121 -12769 4299 -12591
rect -2579 -14369 -2401 -14191
rect 4121 -14369 4299 -14191
rect -2579 -16089 -2401 -15911
rect 4121 -16089 4299 -15911
rect -2579 -17689 -2401 -17511
rect 4121 -17689 4299 -17511
rect -2579 -19409 -2401 -19231
rect 4121 -19409 4299 -19231
<< metal1 >>
rect -210 960 1890 1010
rect -210 -120 -140 960
rect 20 686 120 700
rect 20 634 44 686
rect 96 634 120 686
rect 20 620 120 634
rect 530 686 630 700
rect 530 634 554 686
rect 606 634 630 686
rect 530 620 630 634
rect 1050 686 1150 700
rect 1050 634 1074 686
rect 1126 634 1150 686
rect 1050 620 1150 634
rect 1570 686 1670 700
rect 1570 634 1594 686
rect 1646 634 1670 686
rect 1570 620 1670 634
rect -80 504 90 550
rect -80 470 -67 504
rect -33 470 90 504
rect -80 432 90 470
rect -80 398 -67 432
rect -33 398 90 432
rect -80 360 90 398
rect -80 326 -67 360
rect -33 326 90 360
rect -80 280 90 326
rect 1590 504 1760 550
rect 1590 470 1713 504
rect 1747 470 1760 504
rect 1590 432 1760 470
rect 1590 398 1713 432
rect 1747 398 1760 432
rect 1590 360 1760 398
rect 1590 326 1713 360
rect 1747 326 1760 360
rect 1590 280 1760 326
rect 270 206 370 220
rect 270 154 294 206
rect 346 154 370 206
rect 270 140 370 154
rect 790 206 890 220
rect 790 154 814 206
rect 866 154 890 206
rect 790 140 890 154
rect 1310 206 1410 220
rect 1310 154 1334 206
rect 1386 154 1410 206
rect 1310 140 1410 154
rect 1820 -120 1890 960
rect -210 -139 1890 -120
rect -210 -170 119 -139
rect 100 -191 119 -170
rect 171 -170 819 -139
rect 171 -191 190 -170
rect 100 -200 190 -191
rect 800 -191 819 -170
rect 871 -170 1509 -139
rect 871 -191 890 -170
rect 800 -200 890 -191
rect 1490 -191 1509 -170
rect 1561 -170 1890 -139
rect 1561 -191 1580 -170
rect 1490 -200 1580 -191
rect 100 -469 190 -460
rect 100 -490 119 -469
rect 90 -521 119 -490
rect 171 -490 190 -469
rect 800 -469 890 -460
rect 800 -490 819 -469
rect 171 -521 819 -490
rect 871 -490 890 -469
rect 1490 -469 1580 -460
rect 1490 -490 1509 -469
rect 871 -521 1509 -490
rect 1561 -490 1580 -469
rect 1561 -521 1590 -490
rect 90 -540 1590 -521
rect 300 -700 350 -540
rect 820 -700 870 -540
rect 1330 -700 1380 -540
rect 20 -774 120 -760
rect 20 -826 44 -774
rect 96 -826 120 -774
rect 20 -840 120 -826
rect 530 -774 630 -760
rect 530 -826 554 -774
rect 606 -826 630 -774
rect 530 -840 630 -826
rect 1050 -774 1150 -760
rect 1050 -826 1074 -774
rect 1126 -826 1150 -774
rect 1050 -840 1150 -826
rect 1570 -774 1670 -760
rect 1570 -826 1594 -774
rect 1646 -826 1670 -774
rect 1570 -840 1670 -826
rect -240 -994 -20 -960
rect -240 -1046 -166 -994
rect -114 -1006 -20 -994
rect -114 -1040 -67 -1006
rect -33 -1040 -20 -1006
rect -114 -1046 -20 -1040
rect -240 -1078 -20 -1046
rect -240 -1112 -67 -1078
rect -33 -1112 -20 -1078
rect -240 -1134 -20 -1112
rect -240 -1186 -166 -1134
rect -114 -1150 -20 -1134
rect -114 -1184 -67 -1150
rect -33 -1184 -20 -1150
rect -114 -1186 -20 -1184
rect -240 -1220 -20 -1186
rect 1700 -994 1920 -960
rect 1700 -1006 1794 -994
rect 1700 -1040 1713 -1006
rect 1747 -1040 1794 -1006
rect 1700 -1046 1794 -1040
rect 1846 -1046 1920 -994
rect 1700 -1078 1920 -1046
rect 1700 -1112 1713 -1078
rect 1747 -1112 1920 -1078
rect 1700 -1134 1920 -1112
rect 1700 -1150 1794 -1134
rect 1700 -1184 1713 -1150
rect 1747 -1184 1794 -1150
rect 1700 -1186 1794 -1184
rect 1846 -1186 1920 -1134
rect 1700 -1220 1920 -1186
rect -76 -1222 -24 -1220
rect 1704 -1222 1756 -1220
rect 300 -1620 350 -1460
rect 820 -1620 870 -1450
rect 1330 -1620 1380 -1460
rect -20 -1639 1670 -1620
rect -20 -1654 799 -1639
rect -20 -1706 24 -1654
rect 76 -1670 799 -1654
rect 76 -1706 120 -1670
rect 780 -1691 799 -1670
rect 851 -1654 1670 -1639
rect 851 -1670 1574 -1654
rect 851 -1691 870 -1670
rect 780 -1700 870 -1691
rect -20 -1740 120 -1706
rect 1530 -1706 1574 -1670
rect 1626 -1706 1670 -1654
rect 1530 -1740 1670 -1706
rect 780 -2079 870 -2070
rect 780 -2110 799 -2079
rect 640 -2131 799 -2110
rect 851 -2110 870 -2079
rect 851 -2131 1010 -2110
rect 640 -2160 1010 -2131
rect 524 -2346 576 -2308
rect 524 -2380 533 -2346
rect 567 -2380 576 -2346
rect 640 -2350 690 -2160
rect 960 -2350 1010 -2160
rect 1074 -2346 1126 -2308
rect 1074 -2370 1083 -2346
rect 1070 -2372 1083 -2370
rect 1117 -2370 1126 -2346
rect 1117 -2372 1210 -2370
rect 450 -2382 590 -2380
rect 450 -2498 462 -2382
rect 578 -2498 590 -2382
rect 1070 -2488 1082 -2372
rect 1198 -2488 1210 -2372
rect 1070 -2490 1210 -2488
rect 450 -2500 533 -2498
rect 524 -2524 533 -2500
rect 567 -2500 590 -2498
rect 567 -2524 576 -2500
rect 524 -2562 576 -2524
rect 1074 -2524 1083 -2490
rect 1117 -2524 1126 -2490
rect 780 -2549 870 -2540
rect 780 -2601 799 -2549
rect 851 -2601 870 -2549
rect 1074 -2562 1126 -2524
rect 780 -2610 870 -2601
rect 640 -2720 690 -2680
rect 960 -2720 1010 -2680
rect 640 -2770 1010 -2720
rect 270 -3084 370 -3070
rect 270 -3136 294 -3084
rect 346 -3110 370 -3084
rect 780 -3079 870 -3070
rect 780 -3110 799 -3079
rect 346 -3131 799 -3110
rect 851 -3110 870 -3079
rect 1310 -3084 1410 -3070
rect 1310 -3110 1334 -3084
rect 851 -3131 1334 -3110
rect 346 -3136 1334 -3131
rect 1386 -3136 1410 -3084
rect 270 -3160 1410 -3136
rect 540 -3200 590 -3160
rect 1060 -3190 1110 -3160
rect 130 -3289 360 -3260
rect 1320 -3270 1510 -3260
rect 130 -3298 279 -3289
rect 130 -3332 178 -3298
rect 212 -3332 279 -3298
rect 130 -3341 279 -3332
rect 331 -3341 360 -3289
rect 130 -3370 360 -3341
rect 770 -3289 880 -3270
rect 770 -3341 799 -3289
rect 851 -3341 880 -3289
rect 770 -3360 880 -3341
rect 1280 -3289 1510 -3270
rect 1280 -3341 1309 -3289
rect 1361 -3293 1510 -3289
rect 1361 -3327 1433 -3293
rect 1467 -3327 1510 -3293
rect 1361 -3341 1510 -3327
rect 1280 -3360 1510 -3341
rect 540 -3470 590 -3430
rect 1060 -3470 1110 -3430
rect 330 -3484 1310 -3470
rect 330 -3520 414 -3484
rect 400 -3536 414 -3520
rect 466 -3520 1184 -3484
rect 466 -3536 480 -3520
rect 400 -3540 480 -3536
rect 1170 -3536 1184 -3520
rect 1236 -3520 1310 -3484
rect 1236 -3536 1250 -3520
rect 1170 -3540 1250 -3536
rect 670 -3583 950 -3570
rect 670 -3617 721 -3583
rect 755 -3617 793 -3583
rect 827 -3617 865 -3583
rect 899 -3617 950 -3583
rect 670 -3669 950 -3617
rect 670 -3721 789 -3669
rect 841 -3721 950 -3669
rect 670 -3763 950 -3721
rect 670 -3797 721 -3763
rect 755 -3797 793 -3763
rect 827 -3797 865 -3763
rect 899 -3797 950 -3763
rect 670 -3810 950 -3797
rect 400 -3844 480 -3840
rect 400 -3860 414 -3844
rect -90 -3896 414 -3860
rect 466 -3860 480 -3844
rect 1170 -3844 1250 -3840
rect 1170 -3860 1184 -3844
rect 466 -3896 1184 -3860
rect 1236 -3860 1250 -3844
rect 1236 -3896 1740 -3860
rect -90 -3910 1740 -3896
rect -90 -4970 -30 -3910
rect 10 -4214 90 -4210
rect 10 -4266 24 -4214
rect 76 -4266 90 -4214
rect 10 -4270 90 -4266
rect 530 -4214 610 -4210
rect 530 -4266 544 -4214
rect 596 -4266 610 -4214
rect 530 -4270 610 -4266
rect 1040 -4214 1120 -4210
rect 1040 -4266 1054 -4214
rect 1106 -4266 1120 -4214
rect 1040 -4270 1120 -4266
rect 1560 -4214 1640 -4210
rect 1560 -4266 1574 -4214
rect 1626 -4266 1640 -4214
rect 1560 -4270 1640 -4266
rect 270 -4624 350 -4620
rect 270 -4676 284 -4624
rect 336 -4676 350 -4624
rect 270 -4680 350 -4676
rect 790 -4624 870 -4620
rect 790 -4676 804 -4624
rect 856 -4676 870 -4624
rect 790 -4680 870 -4676
rect 1300 -4624 1380 -4620
rect 1300 -4676 1314 -4624
rect 1366 -4676 1380 -4624
rect 1300 -4680 1380 -4676
rect 1680 -4970 1740 -3910
rect -90 -5020 1740 -4970
rect 670 -5083 950 -5070
rect 670 -5117 721 -5083
rect 755 -5109 793 -5083
rect 827 -5109 865 -5083
rect 755 -5117 789 -5109
rect 841 -5117 865 -5109
rect 899 -5117 950 -5083
rect 670 -5161 789 -5117
rect 841 -5161 950 -5117
rect 670 -5190 950 -5161
rect -1220 -5374 3150 -5350
rect -1220 -5426 284 -5374
rect 336 -5426 1314 -5374
rect 1366 -5426 3150 -5374
rect -1220 -5544 3150 -5426
rect -1220 -5596 284 -5544
rect 336 -5596 1314 -5544
rect 1366 -5596 3150 -5544
rect -1220 -5714 3150 -5596
rect -1220 -5766 284 -5714
rect 336 -5766 1314 -5714
rect 1366 -5766 3150 -5714
rect -1220 -5790 3150 -5766
rect -2622 -5950 -2358 -5914
rect -2622 -6130 -2580 -5950
rect -2400 -6130 -2358 -5950
rect -2622 -6166 -2358 -6130
rect 4078 -5950 4342 -5914
rect 4078 -6130 4120 -5950
rect 4300 -6130 4342 -5950
rect 4078 -6166 4342 -6130
rect -2622 -7670 -2358 -7634
rect -2622 -7850 -2580 -7670
rect -2400 -7850 -2358 -7670
rect -2622 -7886 -2358 -7850
rect 4078 -7670 4342 -7634
rect 4078 -7850 4120 -7670
rect 4300 -7850 4342 -7670
rect 4078 -7886 4342 -7850
rect -2622 -9390 -2358 -9354
rect -2622 -9570 -2580 -9390
rect -2400 -9570 -2358 -9390
rect -2622 -9606 -2358 -9570
rect 4078 -9390 4342 -9354
rect 4078 -9570 4120 -9390
rect 4300 -9570 4342 -9390
rect 4078 -9606 4342 -9570
rect -2622 -10870 -2358 -10834
rect -2622 -11050 -2580 -10870
rect -2400 -11050 -2358 -10870
rect -2622 -11086 -2358 -11050
rect 4078 -10870 4342 -10834
rect 4078 -11050 4120 -10870
rect 4300 -11050 4342 -10870
rect 4078 -11086 4342 -11050
rect -2622 -12590 -2358 -12554
rect -2622 -12770 -2580 -12590
rect -2400 -12770 -2358 -12590
rect -2622 -12806 -2358 -12770
rect 4078 -12590 4342 -12554
rect 4078 -12770 4120 -12590
rect 4300 -12770 4342 -12590
rect 4078 -12806 4342 -12770
rect -2622 -14190 -2358 -14154
rect -2622 -14370 -2580 -14190
rect -2400 -14370 -2358 -14190
rect -2622 -14406 -2358 -14370
rect 4078 -14190 4342 -14154
rect 4078 -14370 4120 -14190
rect 4300 -14370 4342 -14190
rect 4078 -14406 4342 -14370
rect -2622 -15910 -2358 -15874
rect -2622 -16090 -2580 -15910
rect -2400 -16090 -2358 -15910
rect -2622 -16126 -2358 -16090
rect 4078 -15910 4342 -15874
rect 4078 -16090 4120 -15910
rect 4300 -16090 4342 -15910
rect 4078 -16126 4342 -16090
rect -2622 -17510 -2358 -17474
rect -2622 -17690 -2580 -17510
rect -2400 -17690 -2358 -17510
rect -2622 -17726 -2358 -17690
rect 4078 -17510 4342 -17474
rect 4078 -17690 4120 -17510
rect 4300 -17690 4342 -17510
rect 4078 -17726 4342 -17690
rect -2622 -19230 -2358 -19194
rect -2622 -19410 -2580 -19230
rect -2400 -19410 -2358 -19230
rect -2622 -19446 -2358 -19410
rect 4078 -19230 4342 -19194
rect 4078 -19410 4120 -19230
rect 4300 -19410 4342 -19230
rect 4078 -19446 4342 -19410
rect -2630 -19710 4350 -19580
rect -2630 -19890 -2580 -19710
rect -2400 -19890 4120 -19710
rect 4300 -19890 4350 -19710
rect -2630 -20020 4350 -19890
<< via1 >>
rect 44 634 96 686
rect 554 634 606 686
rect 1074 634 1126 686
rect 1594 634 1646 686
rect 294 154 346 206
rect 814 154 866 206
rect 1334 154 1386 206
rect 119 -191 171 -139
rect 819 -191 871 -139
rect 1509 -191 1561 -139
rect 119 -521 171 -469
rect 819 -521 871 -469
rect 1509 -521 1561 -469
rect 44 -826 96 -774
rect 554 -826 606 -774
rect 1074 -826 1126 -774
rect 1594 -826 1646 -774
rect -166 -1046 -114 -994
rect -166 -1186 -114 -1134
rect 1794 -1046 1846 -994
rect 1794 -1186 1846 -1134
rect 24 -1706 76 -1654
rect 799 -1691 851 -1639
rect 1574 -1706 1626 -1654
rect 799 -2131 851 -2079
rect 462 -2418 578 -2382
rect 462 -2452 533 -2418
rect 533 -2452 567 -2418
rect 567 -2452 578 -2418
rect 462 -2490 578 -2452
rect 462 -2498 533 -2490
rect 533 -2498 567 -2490
rect 567 -2498 578 -2490
rect 1082 -2380 1083 -2372
rect 1083 -2380 1117 -2372
rect 1117 -2380 1198 -2372
rect 1082 -2418 1198 -2380
rect 1082 -2452 1083 -2418
rect 1083 -2452 1117 -2418
rect 1117 -2452 1198 -2418
rect 1082 -2488 1198 -2452
rect 799 -2601 851 -2549
rect 294 -3136 346 -3084
rect 799 -3131 851 -3079
rect 1334 -3136 1386 -3084
rect 279 -3341 331 -3289
rect 799 -3341 851 -3289
rect 1309 -3341 1361 -3289
rect 414 -3536 466 -3484
rect 1184 -3536 1236 -3484
rect 789 -3721 841 -3669
rect 414 -3896 466 -3844
rect 1184 -3896 1236 -3844
rect 24 -4266 76 -4214
rect 544 -4266 596 -4214
rect 1054 -4266 1106 -4214
rect 1574 -4266 1626 -4214
rect 284 -4676 336 -4624
rect 804 -4676 856 -4624
rect 1314 -4676 1366 -4624
rect 789 -5117 793 -5109
rect 793 -5117 827 -5109
rect 827 -5117 841 -5109
rect 789 -5161 841 -5117
rect 284 -5426 336 -5374
rect 1314 -5426 1366 -5374
rect 284 -5596 336 -5544
rect 1314 -5596 1366 -5544
rect 284 -5766 336 -5714
rect 1314 -5766 1366 -5714
rect -2580 -5951 -2400 -5950
rect -2580 -6129 -2579 -5951
rect -2579 -6129 -2401 -5951
rect -2401 -6129 -2400 -5951
rect -2580 -6130 -2400 -6129
rect 4120 -5951 4300 -5950
rect 4120 -6129 4121 -5951
rect 4121 -6129 4299 -5951
rect 4299 -6129 4300 -5951
rect 4120 -6130 4300 -6129
rect -2580 -7671 -2400 -7670
rect -2580 -7849 -2579 -7671
rect -2579 -7849 -2401 -7671
rect -2401 -7849 -2400 -7671
rect -2580 -7850 -2400 -7849
rect 4120 -7671 4300 -7670
rect 4120 -7849 4121 -7671
rect 4121 -7849 4299 -7671
rect 4299 -7849 4300 -7671
rect 4120 -7850 4300 -7849
rect -2580 -9391 -2400 -9390
rect -2580 -9569 -2579 -9391
rect -2579 -9569 -2401 -9391
rect -2401 -9569 -2400 -9391
rect -2580 -9570 -2400 -9569
rect 4120 -9391 4300 -9390
rect 4120 -9569 4121 -9391
rect 4121 -9569 4299 -9391
rect 4299 -9569 4300 -9391
rect 4120 -9570 4300 -9569
rect -2580 -10871 -2400 -10870
rect -2580 -11049 -2579 -10871
rect -2579 -11049 -2401 -10871
rect -2401 -11049 -2400 -10871
rect -2580 -11050 -2400 -11049
rect 4120 -10871 4300 -10870
rect 4120 -11049 4121 -10871
rect 4121 -11049 4299 -10871
rect 4299 -11049 4300 -10871
rect 4120 -11050 4300 -11049
rect -2580 -12591 -2400 -12590
rect -2580 -12769 -2579 -12591
rect -2579 -12769 -2401 -12591
rect -2401 -12769 -2400 -12591
rect -2580 -12770 -2400 -12769
rect 4120 -12591 4300 -12590
rect 4120 -12769 4121 -12591
rect 4121 -12769 4299 -12591
rect 4299 -12769 4300 -12591
rect 4120 -12770 4300 -12769
rect -2580 -14191 -2400 -14190
rect -2580 -14369 -2579 -14191
rect -2579 -14369 -2401 -14191
rect -2401 -14369 -2400 -14191
rect -2580 -14370 -2400 -14369
rect 4120 -14191 4300 -14190
rect 4120 -14369 4121 -14191
rect 4121 -14369 4299 -14191
rect 4299 -14369 4300 -14191
rect 4120 -14370 4300 -14369
rect -2580 -15911 -2400 -15910
rect -2580 -16089 -2579 -15911
rect -2579 -16089 -2401 -15911
rect -2401 -16089 -2400 -15911
rect -2580 -16090 -2400 -16089
rect 4120 -15911 4300 -15910
rect 4120 -16089 4121 -15911
rect 4121 -16089 4299 -15911
rect 4299 -16089 4300 -15911
rect 4120 -16090 4300 -16089
rect -2580 -17511 -2400 -17510
rect -2580 -17689 -2579 -17511
rect -2579 -17689 -2401 -17511
rect -2401 -17689 -2400 -17511
rect -2580 -17690 -2400 -17689
rect 4120 -17511 4300 -17510
rect 4120 -17689 4121 -17511
rect 4121 -17689 4299 -17511
rect 4299 -17689 4300 -17511
rect 4120 -17690 4300 -17689
rect -2580 -19231 -2400 -19230
rect -2580 -19409 -2579 -19231
rect -2579 -19409 -2401 -19231
rect -2401 -19409 -2400 -19231
rect -2580 -19410 -2400 -19409
rect 4120 -19231 4300 -19230
rect 4120 -19409 4121 -19231
rect 4121 -19409 4299 -19231
rect 4299 -19409 4300 -19231
rect 4120 -19410 4300 -19409
rect -2580 -19890 -2400 -19710
rect 4120 -19890 4300 -19710
<< metal2 >>
rect 30 688 110 710
rect 30 632 42 688
rect 98 632 110 688
rect 30 610 110 632
rect 540 688 620 710
rect 540 632 552 688
rect 608 632 620 688
rect 540 610 620 632
rect 1060 688 1140 710
rect 1060 632 1072 688
rect 1128 632 1140 688
rect 1060 610 1140 632
rect 1580 688 1660 710
rect 1580 632 1592 688
rect 1648 632 1660 688
rect 1580 610 1660 632
rect 270 208 370 230
rect 270 152 292 208
rect 348 152 370 208
rect 90 -139 200 -120
rect 90 -191 119 -139
rect 171 -191 200 -139
rect 90 -469 200 -191
rect 90 -521 119 -469
rect 171 -521 200 -469
rect 90 -540 200 -521
rect 30 -772 110 -750
rect 30 -828 42 -772
rect 98 -828 110 -772
rect 30 -850 110 -828
rect -180 -992 -100 -970
rect -180 -1048 -168 -992
rect -112 -1048 -100 -992
rect -180 -1070 -100 -1048
rect -180 -1132 -100 -1110
rect -180 -1188 -168 -1132
rect -112 -1188 -100 -1132
rect -180 -1210 -100 -1188
rect -20 -1654 120 -1620
rect -20 -1706 24 -1654
rect 76 -1706 120 -1654
rect -20 -4212 120 -1706
rect 270 -3084 370 152
rect 800 208 880 230
rect 800 152 812 208
rect 868 152 880 208
rect 800 130 880 152
rect 1310 208 1410 230
rect 1310 152 1332 208
rect 1388 152 1410 208
rect 790 -139 900 -120
rect 790 -191 819 -139
rect 871 -191 900 -139
rect 790 -469 900 -191
rect 790 -521 819 -469
rect 871 -521 900 -469
rect 790 -540 900 -521
rect 540 -772 620 -750
rect 540 -828 552 -772
rect 608 -828 620 -772
rect 540 -850 620 -828
rect 1060 -772 1140 -750
rect 1060 -828 1072 -772
rect 1128 -828 1140 -772
rect 1060 -850 1140 -828
rect 780 -1639 870 -1620
rect 780 -1691 799 -1639
rect 851 -1691 870 -1639
rect 780 -2079 870 -1691
rect 780 -2131 799 -2079
rect 851 -2131 870 -2079
rect 780 -2150 870 -2131
rect 460 -2382 580 -2370
rect 460 -2498 462 -2382
rect 578 -2498 580 -2382
rect 460 -2510 580 -2498
rect 1080 -2372 1200 -2360
rect 1080 -2488 1082 -2372
rect 1198 -2488 1200 -2372
rect 1080 -2500 1200 -2488
rect 270 -3136 294 -3084
rect 346 -3136 370 -3084
rect 780 -2549 870 -2530
rect 780 -2601 799 -2549
rect 851 -2601 870 -2549
rect 780 -3079 870 -2601
rect 780 -3110 799 -3079
rect 270 -3160 370 -3136
rect 790 -3131 799 -3110
rect 851 -3110 870 -3079
rect 1310 -3084 1410 152
rect 1480 -139 1590 -120
rect 1480 -191 1509 -139
rect 1561 -191 1590 -139
rect 1480 -469 1590 -191
rect 1480 -521 1509 -469
rect 1561 -521 1590 -469
rect 1480 -540 1590 -521
rect 1580 -772 1660 -750
rect 1580 -828 1592 -772
rect 1648 -828 1660 -772
rect 1580 -850 1660 -828
rect 1780 -992 1860 -970
rect 1780 -1048 1792 -992
rect 1848 -1048 1860 -992
rect 1780 -1070 1860 -1048
rect 1780 -1132 1860 -1110
rect 1780 -1188 1792 -1132
rect 1848 -1188 1860 -1132
rect 1780 -1210 1860 -1188
rect 851 -3131 860 -3110
rect 790 -3150 860 -3131
rect 1310 -3136 1334 -3084
rect 1386 -3136 1410 -3084
rect 1310 -3160 1410 -3136
rect 1530 -1654 1670 -1620
rect 1530 -1706 1574 -1654
rect 1626 -1706 1670 -1654
rect 260 -3287 350 -3260
rect 260 -3343 277 -3287
rect 333 -3343 350 -3287
rect 260 -3370 350 -3343
rect 780 -3287 870 -3260
rect 780 -3343 797 -3287
rect 853 -3343 870 -3287
rect 780 -3370 870 -3343
rect 1290 -3287 1380 -3260
rect 1290 -3343 1307 -3287
rect 1363 -3343 1380 -3287
rect 1290 -3370 1380 -3343
rect 400 -3484 480 -3470
rect 400 -3536 414 -3484
rect 466 -3536 480 -3484
rect 400 -3844 480 -3536
rect 1170 -3484 1250 -3470
rect 1170 -3536 1184 -3484
rect 1236 -3536 1250 -3484
rect 770 -3667 860 -3640
rect 770 -3723 787 -3667
rect 843 -3723 860 -3667
rect 770 -3750 860 -3723
rect 400 -3896 414 -3844
rect 466 -3896 480 -3844
rect 400 -3910 480 -3896
rect 1170 -3844 1250 -3536
rect 1170 -3896 1184 -3844
rect 1236 -3896 1250 -3844
rect 1170 -3910 1250 -3896
rect -20 -4268 22 -4212
rect 78 -4268 120 -4212
rect -20 -4280 120 -4268
rect 540 -4212 600 -4200
rect 540 -4268 542 -4212
rect 598 -4268 600 -4212
rect 540 -4280 600 -4268
rect 1050 -4212 1110 -4200
rect 1050 -4268 1052 -4212
rect 1108 -4268 1110 -4212
rect 1050 -4280 1110 -4268
rect 1530 -4212 1670 -1706
rect 1530 -4268 1572 -4212
rect 1628 -4268 1670 -4212
rect 1530 -4280 1670 -4268
rect 260 -4622 360 -4610
rect 260 -4678 282 -4622
rect 338 -4678 360 -4622
rect 260 -5374 360 -4678
rect 800 -4622 860 -4610
rect 800 -4678 802 -4622
rect 858 -4678 860 -4622
rect 800 -4690 860 -4678
rect 1290 -4622 1390 -4610
rect 1290 -4678 1312 -4622
rect 1368 -4678 1390 -4622
rect 770 -5107 860 -5080
rect 770 -5163 787 -5107
rect 843 -5163 860 -5107
rect 770 -5190 860 -5163
rect 260 -5426 284 -5374
rect 336 -5426 360 -5374
rect 260 -5544 360 -5426
rect 260 -5596 284 -5544
rect 336 -5596 360 -5544
rect 260 -5714 360 -5596
rect 260 -5766 284 -5714
rect 336 -5766 360 -5714
rect 260 -5790 360 -5766
rect 1290 -5374 1390 -4678
rect 1290 -5426 1314 -5374
rect 1366 -5426 1390 -5374
rect 1290 -5544 1390 -5426
rect 1290 -5596 1314 -5544
rect 1366 -5596 1390 -5544
rect 1290 -5714 1390 -5596
rect 1290 -5766 1314 -5714
rect 1366 -5766 1390 -5714
rect 1290 -5790 1390 -5766
rect -2630 -5932 -2350 -5880
rect -2630 -6148 -2598 -5932
rect -2382 -6148 -2350 -5932
rect -2630 -7652 -2350 -6148
rect -2630 -7868 -2598 -7652
rect -2382 -7868 -2350 -7652
rect -2630 -9372 -2350 -7868
rect -2630 -9588 -2598 -9372
rect -2382 -9588 -2350 -9372
rect -2630 -10852 -2350 -9588
rect -2630 -11068 -2598 -10852
rect -2382 -11068 -2350 -10852
rect -2630 -12572 -2350 -11068
rect -2630 -12788 -2598 -12572
rect -2382 -12788 -2350 -12572
rect -2630 -14172 -2350 -12788
rect -2630 -14388 -2598 -14172
rect -2382 -14388 -2350 -14172
rect -2630 -15892 -2350 -14388
rect -2630 -16108 -2598 -15892
rect -2382 -16108 -2350 -15892
rect -2630 -17492 -2350 -16108
rect -2630 -17708 -2598 -17492
rect -2382 -17708 -2350 -17492
rect -2630 -19212 -2350 -17708
rect -2630 -19428 -2598 -19212
rect -2382 -19428 -2350 -19212
rect -2630 -19710 -2350 -19428
rect -2630 -19890 -2580 -19710
rect -2400 -19890 -2350 -19710
rect -2630 -20020 -2350 -19890
rect 4070 -5932 4350 -5880
rect 4070 -6148 4102 -5932
rect 4318 -6148 4350 -5932
rect 4070 -7652 4350 -6148
rect 4070 -7868 4102 -7652
rect 4318 -7868 4350 -7652
rect 4070 -9372 4350 -7868
rect 4070 -9588 4102 -9372
rect 4318 -9588 4350 -9372
rect 4070 -10852 4350 -9588
rect 4070 -11068 4102 -10852
rect 4318 -11068 4350 -10852
rect 4070 -12572 4350 -11068
rect 4070 -12788 4102 -12572
rect 4318 -12788 4350 -12572
rect 4070 -14172 4350 -12788
rect 4070 -14388 4102 -14172
rect 4318 -14388 4350 -14172
rect 4070 -15892 4350 -14388
rect 4070 -16108 4102 -15892
rect 4318 -16108 4350 -15892
rect 4070 -17492 4350 -16108
rect 4070 -17708 4102 -17492
rect 4318 -17708 4350 -17492
rect 4070 -19212 4350 -17708
rect 4070 -19428 4102 -19212
rect 4318 -19428 4350 -19212
rect 4070 -19710 4350 -19428
rect 4070 -19890 4120 -19710
rect 4300 -19890 4350 -19710
rect 4070 -20020 4350 -19890
<< via2 >>
rect 42 686 98 688
rect 42 634 44 686
rect 44 634 96 686
rect 96 634 98 686
rect 42 632 98 634
rect 552 686 608 688
rect 552 634 554 686
rect 554 634 606 686
rect 606 634 608 686
rect 552 632 608 634
rect 1072 686 1128 688
rect 1072 634 1074 686
rect 1074 634 1126 686
rect 1126 634 1128 686
rect 1072 632 1128 634
rect 1592 686 1648 688
rect 1592 634 1594 686
rect 1594 634 1646 686
rect 1646 634 1648 686
rect 1592 632 1648 634
rect 292 206 348 208
rect 292 154 294 206
rect 294 154 346 206
rect 346 154 348 206
rect 292 152 348 154
rect 42 -774 98 -772
rect 42 -826 44 -774
rect 44 -826 96 -774
rect 96 -826 98 -774
rect 42 -828 98 -826
rect -168 -994 -112 -992
rect -168 -1046 -166 -994
rect -166 -1046 -114 -994
rect -114 -1046 -112 -994
rect -168 -1048 -112 -1046
rect -168 -1134 -112 -1132
rect -168 -1186 -166 -1134
rect -166 -1186 -114 -1134
rect -114 -1186 -112 -1134
rect -168 -1188 -112 -1186
rect 812 206 868 208
rect 812 154 814 206
rect 814 154 866 206
rect 866 154 868 206
rect 812 152 868 154
rect 1332 206 1388 208
rect 1332 154 1334 206
rect 1334 154 1386 206
rect 1386 154 1388 206
rect 1332 152 1388 154
rect 552 -774 608 -772
rect 552 -826 554 -774
rect 554 -826 606 -774
rect 606 -826 608 -774
rect 552 -828 608 -826
rect 1072 -774 1128 -772
rect 1072 -826 1074 -774
rect 1074 -826 1126 -774
rect 1126 -826 1128 -774
rect 1072 -828 1128 -826
rect 492 -2468 548 -2412
rect 1112 -2458 1168 -2402
rect 1592 -774 1648 -772
rect 1592 -826 1594 -774
rect 1594 -826 1646 -774
rect 1646 -826 1648 -774
rect 1592 -828 1648 -826
rect 1792 -994 1848 -992
rect 1792 -1046 1794 -994
rect 1794 -1046 1846 -994
rect 1846 -1046 1848 -994
rect 1792 -1048 1848 -1046
rect 1792 -1134 1848 -1132
rect 1792 -1186 1794 -1134
rect 1794 -1186 1846 -1134
rect 1846 -1186 1848 -1134
rect 1792 -1188 1848 -1186
rect 277 -3289 333 -3287
rect 277 -3341 279 -3289
rect 279 -3341 331 -3289
rect 331 -3341 333 -3289
rect 277 -3343 333 -3341
rect 797 -3289 853 -3287
rect 797 -3341 799 -3289
rect 799 -3341 851 -3289
rect 851 -3341 853 -3289
rect 797 -3343 853 -3341
rect 1307 -3289 1363 -3287
rect 1307 -3341 1309 -3289
rect 1309 -3341 1361 -3289
rect 1361 -3341 1363 -3289
rect 1307 -3343 1363 -3341
rect 787 -3669 843 -3667
rect 787 -3721 789 -3669
rect 789 -3721 841 -3669
rect 841 -3721 843 -3669
rect 787 -3723 843 -3721
rect 22 -4214 78 -4212
rect 22 -4266 24 -4214
rect 24 -4266 76 -4214
rect 76 -4266 78 -4214
rect 22 -4268 78 -4266
rect 542 -4214 598 -4212
rect 542 -4266 544 -4214
rect 544 -4266 596 -4214
rect 596 -4266 598 -4214
rect 542 -4268 598 -4266
rect 1052 -4214 1108 -4212
rect 1052 -4266 1054 -4214
rect 1054 -4266 1106 -4214
rect 1106 -4266 1108 -4214
rect 1052 -4268 1108 -4266
rect 1572 -4214 1628 -4212
rect 1572 -4266 1574 -4214
rect 1574 -4266 1626 -4214
rect 1626 -4266 1628 -4214
rect 1572 -4268 1628 -4266
rect 282 -4624 338 -4622
rect 282 -4676 284 -4624
rect 284 -4676 336 -4624
rect 336 -4676 338 -4624
rect 282 -4678 338 -4676
rect 802 -4624 858 -4622
rect 802 -4676 804 -4624
rect 804 -4676 856 -4624
rect 856 -4676 858 -4624
rect 802 -4678 858 -4676
rect 1312 -4624 1368 -4622
rect 1312 -4676 1314 -4624
rect 1314 -4676 1366 -4624
rect 1366 -4676 1368 -4624
rect 1312 -4678 1368 -4676
rect 787 -5109 843 -5107
rect 787 -5161 789 -5109
rect 789 -5161 841 -5109
rect 841 -5161 843 -5109
rect 787 -5163 843 -5161
rect -2598 -5950 -2382 -5932
rect -2598 -6130 -2580 -5950
rect -2580 -6130 -2400 -5950
rect -2400 -6130 -2382 -5950
rect -2598 -6148 -2382 -6130
rect -2598 -7670 -2382 -7652
rect -2598 -7850 -2580 -7670
rect -2580 -7850 -2400 -7670
rect -2400 -7850 -2382 -7670
rect -2598 -7868 -2382 -7850
rect -2598 -9390 -2382 -9372
rect -2598 -9570 -2580 -9390
rect -2580 -9570 -2400 -9390
rect -2400 -9570 -2382 -9390
rect -2598 -9588 -2382 -9570
rect -2598 -10870 -2382 -10852
rect -2598 -11050 -2580 -10870
rect -2580 -11050 -2400 -10870
rect -2400 -11050 -2382 -10870
rect -2598 -11068 -2382 -11050
rect -2598 -12590 -2382 -12572
rect -2598 -12770 -2580 -12590
rect -2580 -12770 -2400 -12590
rect -2400 -12770 -2382 -12590
rect -2598 -12788 -2382 -12770
rect -2598 -14190 -2382 -14172
rect -2598 -14370 -2580 -14190
rect -2580 -14370 -2400 -14190
rect -2400 -14370 -2382 -14190
rect -2598 -14388 -2382 -14370
rect -2598 -15910 -2382 -15892
rect -2598 -16090 -2580 -15910
rect -2580 -16090 -2400 -15910
rect -2400 -16090 -2382 -15910
rect -2598 -16108 -2382 -16090
rect -2598 -17510 -2382 -17492
rect -2598 -17690 -2580 -17510
rect -2580 -17690 -2400 -17510
rect -2400 -17690 -2382 -17510
rect -2598 -17708 -2382 -17690
rect -2598 -19230 -2382 -19212
rect -2598 -19410 -2580 -19230
rect -2580 -19410 -2400 -19230
rect -2400 -19410 -2382 -19230
rect -2598 -19428 -2382 -19410
rect 4102 -5950 4318 -5932
rect 4102 -6130 4120 -5950
rect 4120 -6130 4300 -5950
rect 4300 -6130 4318 -5950
rect 4102 -6148 4318 -6130
rect 4102 -7670 4318 -7652
rect 4102 -7850 4120 -7670
rect 4120 -7850 4300 -7670
rect 4300 -7850 4318 -7670
rect 4102 -7868 4318 -7850
rect 4102 -9390 4318 -9372
rect 4102 -9570 4120 -9390
rect 4120 -9570 4300 -9390
rect 4300 -9570 4318 -9390
rect 4102 -9588 4318 -9570
rect 4102 -10870 4318 -10852
rect 4102 -11050 4120 -10870
rect 4120 -11050 4300 -10870
rect 4300 -11050 4318 -10870
rect 4102 -11068 4318 -11050
rect 4102 -12590 4318 -12572
rect 4102 -12770 4120 -12590
rect 4120 -12770 4300 -12590
rect 4300 -12770 4318 -12590
rect 4102 -12788 4318 -12770
rect 4102 -14190 4318 -14172
rect 4102 -14370 4120 -14190
rect 4120 -14370 4300 -14190
rect 4300 -14370 4318 -14190
rect 4102 -14388 4318 -14370
rect 4102 -15910 4318 -15892
rect 4102 -16090 4120 -15910
rect 4120 -16090 4300 -15910
rect 4300 -16090 4318 -15910
rect 4102 -16108 4318 -16090
rect 4102 -17510 4318 -17492
rect 4102 -17690 4120 -17510
rect 4120 -17690 4300 -17510
rect 4300 -17690 4318 -17510
rect 4102 -17708 4318 -17690
rect 4102 -19230 4318 -19212
rect 4102 -19410 4120 -19230
rect 4120 -19410 4300 -19230
rect 4300 -19410 4318 -19230
rect 4102 -19428 4318 -19410
<< metal3 >>
rect -10 692 1670 720
rect -10 628 28 692
rect 92 688 548 692
rect 98 632 548 688
rect 92 628 548 632
rect 612 628 1068 692
rect 1132 628 1588 692
rect 1652 628 1670 692
rect -10 600 1670 628
rect 40 208 1640 240
rect 40 152 292 208
rect 348 152 812 208
rect 868 152 1332 208
rect 1388 152 1640 208
rect 40 120 1640 152
rect -240 -768 1920 -740
rect -240 -832 -172 -768
rect -108 -772 1788 -768
rect -108 -828 42 -772
rect 98 -828 552 -772
rect 608 -828 1072 -772
rect 1128 -828 1592 -772
rect 1648 -828 1788 -772
rect -108 -832 1788 -828
rect 1852 -832 1920 -768
rect -240 -860 1920 -832
rect -200 -988 -80 -960
rect -200 -1052 -172 -988
rect -108 -1052 -80 -988
rect -200 -1128 -80 -1052
rect -200 -1192 -172 -1128
rect -108 -1192 -80 -1128
rect -200 -1220 -80 -1192
rect 1760 -988 1880 -960
rect 1760 -1052 1788 -988
rect 1852 -1052 1880 -988
rect 1760 -1128 1880 -1052
rect 1760 -1192 1788 -1128
rect 1852 -1192 1880 -1128
rect 1760 -1220 1880 -1192
rect 450 -2408 590 -2375
rect 450 -2472 488 -2408
rect 552 -2472 590 -2408
rect 450 -2505 590 -2472
rect 1070 -2398 1210 -2365
rect 1070 -2462 1108 -2398
rect 1172 -2462 1210 -2398
rect 1070 -2495 1210 -2462
rect 240 -3283 1400 -3250
rect 240 -3287 793 -3283
rect 857 -3287 1400 -3283
rect 240 -3343 277 -3287
rect 333 -3343 793 -3287
rect 857 -3343 1307 -3287
rect 1363 -3343 1400 -3287
rect 240 -3347 793 -3343
rect 857 -3347 1400 -3343
rect 240 -3380 1400 -3347
rect 760 -3663 870 -3645
rect 760 -3727 783 -3663
rect 847 -3727 870 -3663
rect 760 -3745 870 -3727
rect 10 -4212 1640 -4200
rect 10 -4268 22 -4212
rect 78 -4268 542 -4212
rect 598 -4268 1052 -4212
rect 1108 -4268 1572 -4212
rect 1628 -4268 1640 -4212
rect 10 -4280 1640 -4268
rect 30 -4622 1620 -4610
rect 30 -4678 282 -4622
rect 338 -4678 802 -4622
rect 858 -4678 1312 -4622
rect 1368 -4678 1620 -4622
rect 30 -4690 1620 -4678
rect 760 -5103 870 -5085
rect 760 -5167 783 -5103
rect 847 -5167 870 -5103
rect 760 -5185 870 -5167
rect -2620 -5932 -2360 -5915
rect -2620 -6148 -2598 -5932
rect -2382 -6148 -2360 -5932
rect -2620 -6165 -2360 -6148
rect 4080 -5932 4340 -5915
rect 4080 -6148 4102 -5932
rect 4318 -6148 4340 -5932
rect 4080 -6165 4340 -6148
rect -2620 -7652 -2360 -7635
rect -2620 -7868 -2598 -7652
rect -2382 -7868 -2360 -7652
rect -2620 -7885 -2360 -7868
rect 4080 -7652 4340 -7635
rect 4080 -7868 4102 -7652
rect 4318 -7868 4340 -7652
rect 4080 -7885 4340 -7868
rect -2620 -9368 -2360 -9355
rect -2620 -9592 -2602 -9368
rect -2378 -9592 -2360 -9368
rect -2620 -9605 -2360 -9592
rect 4080 -9368 4340 -9355
rect 4080 -9592 4098 -9368
rect 4322 -9592 4340 -9368
rect 4080 -9605 4340 -9592
rect -2620 -10852 -2360 -10835
rect -2620 -11068 -2598 -10852
rect -2382 -11068 -2360 -10852
rect -2620 -11085 -2360 -11068
rect 4080 -10852 4340 -10835
rect 4080 -11068 4102 -10852
rect 4318 -11068 4340 -10852
rect 4080 -11085 4340 -11068
rect -2620 -12568 -2360 -12555
rect -2620 -12792 -2602 -12568
rect -2378 -12792 -2360 -12568
rect -2620 -12805 -2360 -12792
rect 4080 -12568 4340 -12555
rect 4080 -12792 4098 -12568
rect 4322 -12792 4340 -12568
rect 4080 -12805 4340 -12792
rect -2620 -14172 -2360 -14155
rect -2620 -14388 -2598 -14172
rect -2382 -14388 -2360 -14172
rect -2620 -14405 -2360 -14388
rect 4080 -14172 4340 -14155
rect 4080 -14388 4102 -14172
rect 4318 -14388 4340 -14172
rect 4080 -14405 4340 -14388
rect -2620 -15888 -2360 -15875
rect -2620 -16112 -2602 -15888
rect -2378 -16112 -2360 -15888
rect -2620 -16125 -2360 -16112
rect 4080 -15888 4340 -15875
rect 4080 -16112 4098 -15888
rect 4322 -16112 4340 -15888
rect 4080 -16125 4340 -16112
rect -2620 -17492 -2360 -17475
rect -2620 -17708 -2598 -17492
rect -2382 -17708 -2360 -17492
rect -2620 -17725 -2360 -17708
rect 4080 -17492 4340 -17475
rect 4080 -17708 4102 -17492
rect 4318 -17708 4340 -17492
rect 4080 -17725 4340 -17708
rect -2620 -19212 -2360 -19195
rect -2620 -19428 -2598 -19212
rect -2382 -19428 -2360 -19212
rect -2620 -19445 -2360 -19428
rect 4080 -19212 4340 -19195
rect 4080 -19428 4102 -19212
rect 4318 -19428 4340 -19212
rect 4080 -19445 4340 -19428
<< via3 >>
rect 28 688 92 692
rect 548 688 612 692
rect 28 632 42 688
rect 42 632 92 688
rect 548 632 552 688
rect 552 632 608 688
rect 608 632 612 688
rect 28 628 92 632
rect 548 628 612 632
rect 1068 688 1132 692
rect 1068 632 1072 688
rect 1072 632 1128 688
rect 1128 632 1132 688
rect 1068 628 1132 632
rect 1588 688 1652 692
rect 1588 632 1592 688
rect 1592 632 1648 688
rect 1648 632 1652 688
rect 1588 628 1652 632
rect -172 -832 -108 -768
rect 1788 -832 1852 -768
rect -172 -992 -108 -988
rect -172 -1048 -168 -992
rect -168 -1048 -112 -992
rect -112 -1048 -108 -992
rect -172 -1052 -108 -1048
rect -172 -1132 -108 -1128
rect -172 -1188 -168 -1132
rect -168 -1188 -112 -1132
rect -112 -1188 -108 -1132
rect -172 -1192 -108 -1188
rect 1788 -992 1852 -988
rect 1788 -1048 1792 -992
rect 1792 -1048 1848 -992
rect 1848 -1048 1852 -992
rect 1788 -1052 1852 -1048
rect 1788 -1132 1852 -1128
rect 1788 -1188 1792 -1132
rect 1792 -1188 1848 -1132
rect 1848 -1188 1852 -1132
rect 1788 -1192 1852 -1188
rect 488 -2412 552 -2408
rect 488 -2468 492 -2412
rect 492 -2468 548 -2412
rect 548 -2468 552 -2412
rect 488 -2472 552 -2468
rect 1108 -2402 1172 -2398
rect 1108 -2458 1112 -2402
rect 1112 -2458 1168 -2402
rect 1168 -2458 1172 -2402
rect 1108 -2462 1172 -2458
rect 793 -3287 857 -3283
rect 793 -3343 797 -3287
rect 797 -3343 853 -3287
rect 853 -3343 857 -3287
rect 793 -3347 857 -3343
rect 783 -3667 847 -3663
rect 783 -3723 787 -3667
rect 787 -3723 843 -3667
rect 843 -3723 847 -3667
rect 783 -3727 847 -3723
rect 783 -5107 847 -5103
rect 783 -5163 787 -5107
rect 787 -5163 843 -5107
rect 843 -5163 847 -5107
rect 783 -5167 847 -5163
rect -2602 -9372 -2378 -9368
rect -2602 -9588 -2598 -9372
rect -2598 -9588 -2382 -9372
rect -2382 -9588 -2378 -9372
rect -2602 -9592 -2378 -9588
rect 4098 -9372 4322 -9368
rect 4098 -9588 4102 -9372
rect 4102 -9588 4318 -9372
rect 4318 -9588 4322 -9372
rect 4098 -9592 4322 -9588
rect -2602 -12572 -2378 -12568
rect -2602 -12788 -2598 -12572
rect -2598 -12788 -2382 -12572
rect -2382 -12788 -2378 -12572
rect -2602 -12792 -2378 -12788
rect 4098 -12572 4322 -12568
rect 4098 -12788 4102 -12572
rect 4102 -12788 4318 -12572
rect 4318 -12788 4322 -12572
rect 4098 -12792 4322 -12788
rect -2602 -15892 -2378 -15888
rect -2602 -16108 -2598 -15892
rect -2598 -16108 -2382 -15892
rect -2382 -16108 -2378 -15892
rect -2602 -16112 -2378 -16108
rect 4098 -15892 4322 -15888
rect 4098 -16108 4102 -15892
rect 4102 -16108 4318 -15892
rect 4318 -16108 4322 -15892
rect 4098 -16112 4322 -16108
<< metal4 >>
rect -240 778 180 780
rect -240 542 -58 778
rect 178 542 180 778
rect -240 540 180 542
rect 460 778 700 780
rect 460 542 462 778
rect 698 542 700 778
rect 460 540 700 542
rect 980 778 1220 780
rect 980 542 982 778
rect 1218 542 1220 778
rect 980 540 1220 542
rect 1500 778 1920 780
rect 1500 542 1502 778
rect 1738 542 1920 778
rect 1500 540 1920 542
rect -240 -768 -20 540
rect -240 -832 -172 -768
rect -108 -832 -20 -768
rect -240 -988 -20 -832
rect -240 -1052 -172 -988
rect -108 -1052 -20 -988
rect -240 -1128 -20 -1052
rect -240 -1192 -172 -1128
rect -108 -1192 -20 -1128
rect -240 -1220 -20 -1192
rect 1700 -768 1920 540
rect 1700 -832 1788 -768
rect 1852 -832 1920 -768
rect 1700 -988 1920 -832
rect 1700 -1052 1788 -988
rect 1852 -1052 1920 -988
rect 1700 -1128 1920 -1052
rect 1700 -1192 1788 -1128
rect 1852 -1192 1920 -1128
rect 1700 -1220 1920 -1192
rect 320 -2398 1280 -2200
rect 320 -2408 1108 -2398
rect 320 -2472 488 -2408
rect 552 -2462 1108 -2408
rect 1172 -2462 1280 -2398
rect 552 -2472 1280 -2462
rect 320 -3283 1280 -2472
rect 320 -3347 793 -3283
rect 857 -3347 1280 -3283
rect 320 -3663 1280 -3347
rect 320 -3727 783 -3663
rect 847 -3727 1280 -3663
rect 320 -5103 1280 -3727
rect 320 -5167 783 -5103
rect 847 -5167 1280 -5103
rect 320 -8882 1280 -5167
rect 320 -9118 402 -8882
rect 638 -9118 962 -8882
rect 1198 -9118 1280 -8882
rect -2611 -9362 -2369 -9359
rect -2611 -9598 -2608 -9362
rect -2372 -9598 -2369 -9362
rect -2611 -9601 -2369 -9598
rect 320 -9362 1280 -9118
rect 320 -9598 402 -9362
rect 638 -9598 962 -9362
rect 1198 -9598 1280 -9362
rect 320 -9842 1280 -9598
rect 4089 -9362 4331 -9359
rect 4089 -9598 4092 -9362
rect 4328 -9598 4331 -9362
rect 4089 -9601 4331 -9598
rect 320 -10078 402 -9842
rect 638 -10078 962 -9842
rect 1198 -10078 1280 -9842
rect 320 -12082 1280 -10078
rect 320 -12318 402 -12082
rect 638 -12318 962 -12082
rect 1198 -12318 1280 -12082
rect -2611 -12562 -2369 -12559
rect -2611 -12798 -2608 -12562
rect -2372 -12798 -2369 -12562
rect -2611 -12801 -2369 -12798
rect 320 -12562 1280 -12318
rect 320 -12798 402 -12562
rect 638 -12798 962 -12562
rect 1198 -12798 1280 -12562
rect 320 -13042 1280 -12798
rect 4089 -12562 4331 -12559
rect 4089 -12798 4092 -12562
rect 4328 -12798 4331 -12562
rect 4089 -12801 4331 -12798
rect 320 -13278 402 -13042
rect 638 -13278 962 -13042
rect 1198 -13278 1280 -13042
rect 320 -15402 1280 -13278
rect 320 -15638 402 -15402
rect 638 -15638 962 -15402
rect 1198 -15638 1280 -15402
rect -2611 -15882 -2369 -15879
rect -2611 -16118 -2608 -15882
rect -2372 -16118 -2369 -15882
rect -2611 -16121 -2369 -16118
rect 320 -15882 1280 -15638
rect 320 -16118 402 -15882
rect 638 -16118 962 -15882
rect 1198 -16118 1280 -15882
rect 320 -16362 1280 -16118
rect 4089 -15882 4331 -15879
rect 4089 -16118 4092 -15882
rect 4328 -16118 4331 -15882
rect 4089 -16121 4331 -16118
rect 320 -16598 402 -16362
rect 638 -16598 962 -16362
rect 1198 -16598 1280 -16362
rect 320 -16680 1280 -16598
<< via4 >>
rect -58 692 178 778
rect -58 628 28 692
rect 28 628 92 692
rect 92 628 178 692
rect -58 542 178 628
rect 462 692 698 778
rect 462 628 548 692
rect 548 628 612 692
rect 612 628 698 692
rect 462 542 698 628
rect 982 692 1218 778
rect 982 628 1068 692
rect 1068 628 1132 692
rect 1132 628 1218 692
rect 982 542 1218 628
rect 1502 692 1738 778
rect 1502 628 1588 692
rect 1588 628 1652 692
rect 1652 628 1738 692
rect 1502 542 1738 628
rect 402 -9118 638 -8882
rect 962 -9118 1198 -8882
rect -2608 -9368 -2372 -9362
rect -2608 -9592 -2602 -9368
rect -2602 -9592 -2378 -9368
rect -2378 -9592 -2372 -9368
rect -2608 -9598 -2372 -9592
rect 402 -9598 638 -9362
rect 962 -9598 1198 -9362
rect 4092 -9368 4328 -9362
rect 4092 -9592 4098 -9368
rect 4098 -9592 4322 -9368
rect 4322 -9592 4328 -9368
rect 4092 -9598 4328 -9592
rect 402 -10078 638 -9842
rect 962 -10078 1198 -9842
rect 402 -12318 638 -12082
rect 962 -12318 1198 -12082
rect -2608 -12568 -2372 -12562
rect -2608 -12792 -2602 -12568
rect -2602 -12792 -2378 -12568
rect -2378 -12792 -2372 -12568
rect -2608 -12798 -2372 -12792
rect 402 -12798 638 -12562
rect 962 -12798 1198 -12562
rect 4092 -12568 4328 -12562
rect 4092 -12792 4098 -12568
rect 4098 -12792 4322 -12568
rect 4322 -12792 4328 -12568
rect 4092 -12798 4328 -12792
rect 402 -13278 638 -13042
rect 962 -13278 1198 -13042
rect 402 -15638 638 -15402
rect 962 -15638 1198 -15402
rect -2608 -15888 -2372 -15882
rect -2608 -16112 -2602 -15888
rect -2602 -16112 -2378 -15888
rect -2378 -16112 -2372 -15888
rect -2608 -16118 -2372 -16112
rect 402 -16118 638 -15882
rect 962 -16118 1198 -15882
rect 4092 -15888 4328 -15882
rect 4092 -16112 4098 -15888
rect 4098 -16112 4322 -15888
rect 4322 -16112 4328 -15888
rect 4092 -16118 4328 -16112
rect 402 -16598 638 -16362
rect 962 -16598 1198 -16362
<< metal5 >>
rect -320 778 2040 1120
rect -320 542 -58 778
rect 178 542 462 778
rect 698 542 982 778
rect 1218 542 1502 778
rect 1738 542 2040 778
rect -320 480 2040 542
rect -2690 -8882 4420 -8790
rect -2690 -9118 402 -8882
rect 638 -9118 962 -8882
rect 1198 -9118 4420 -8882
rect -2690 -9362 4420 -9118
rect -2690 -9598 -2608 -9362
rect -2372 -9598 402 -9362
rect 638 -9598 962 -9362
rect 1198 -9598 4092 -9362
rect 4328 -9598 4420 -9362
rect -2690 -9842 4420 -9598
rect -2690 -10078 402 -9842
rect 638 -10078 962 -9842
rect 1198 -10078 4420 -9842
rect -2690 -10160 4420 -10078
rect -2700 -12082 4410 -12000
rect -2700 -12318 402 -12082
rect 638 -12318 962 -12082
rect 1198 -12318 4410 -12082
rect -2700 -12562 4410 -12318
rect -2700 -12798 -2608 -12562
rect -2372 -12798 402 -12562
rect 638 -12798 962 -12562
rect 1198 -12798 4092 -12562
rect 4328 -12798 4410 -12562
rect -2700 -13042 4410 -12798
rect -2700 -13278 402 -13042
rect 638 -13278 962 -13042
rect 1198 -13278 4410 -13042
rect -2700 -13370 4410 -13278
rect -2690 -15402 4410 -15320
rect -2690 -15638 402 -15402
rect 638 -15638 962 -15402
rect 1198 -15638 4410 -15402
rect -2690 -15882 4410 -15638
rect -2690 -16118 -2608 -15882
rect -2372 -16118 402 -15882
rect 638 -16118 962 -15882
rect 1198 -16118 4092 -15882
rect 4328 -16118 4410 -15882
rect -2690 -16362 4410 -16118
rect -2690 -16598 402 -16362
rect 638 -16598 962 -16362
rect 1198 -16598 4410 -16362
rect -2690 -16680 4410 -16598
use sky130_fd_pr__nfet_01v8_A5635U  sky130_fd_pr__nfet_01v8_A5635U_0
timestamp 1710000196
transform 1 0 823 0 1 -3315
box -673 -325 673 325
use sky130_fd_pr__nfet_01v8_GLZPWL  sky130_fd_pr__nfet_01v8_GLZPWL_0
timestamp 1710000196
transform 1 0 826 0 1 -4440
box -931 -700 931 700
use sky130_fd_pr__nfet_01v8_H7FLKU  sky130_fd_pr__nfet_01v8_H7FLKU_0
timestamp 1710000196
transform 1 0 825 0 1 -2440
box -315 -450 315 450
use sky130_fd_pr__pfet_01v8_LK874N  sky130_fd_pr__pfet_01v8_LK874N_0
timestamp 1710000196
transform 1 0 841 0 1 419
box -941 -719 941 719
use sky130_fd_pr__pfet_01v8_LK874N  sky130_fd_pr__pfet_01v8_LK874N_1
timestamp 1710000196
transform 1 0 841 0 1 -1081
box -941 -719 941 719
use sky130_fd_pr__res_xhigh_po_5p73_B5N4SD  sky130_fd_pr__res_xhigh_po_5p73_B5N4SD_0
timestamp 1710000196
transform 1 0 1575 0 1 -12688
box -573 -7332 573 7332
use sky130_fd_pr__res_xhigh_po_5p73_B5N4SD  sky130_fd_pr__res_xhigh_po_5p73_B5N4SD_1
timestamp 1710000196
transform 1 0 35 0 1 -12688
box -573 -7332 573 7332
use sky130_fd_pr__res_xhigh_po_5p73_B5N4SD  sky130_fd_pr__res_xhigh_po_5p73_B5N4SD_2
timestamp 1710000196
transform 1 0 -1515 0 1 -12688
box -573 -7332 573 7332
use sky130_fd_pr__res_xhigh_po_5p73_B5N4SD  sky130_fd_pr__res_xhigh_po_5p73_B5N4SD_3
timestamp 1710000196
transform 1 0 3125 0 1 -12688
box -573 -7332 573 7332
<< labels >>
rlabel metal5 s -438 -12860 -438 -12860 4 VSS
rlabel metal3 s 582 184 582 184 4 Vout
rlabel metal5 s 290 1000 290 1000 4 VDD
<< end >>
