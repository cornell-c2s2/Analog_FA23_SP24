magic
tech sky130A
magscale 1 2
timestamp 1710014858
<< pwell >>
rect 3450 -2700 4650 -2600
<< viali >>
rect 1625 50 1675 100
rect 1825 50 1875 100
rect 2050 50 2100 100
rect 2626 92 2666 132
rect 3026 92 3066 132
rect 3426 92 3466 132
rect 3826 92 3866 132
rect 4226 92 4266 132
rect 5026 92 5066 132
rect 5426 92 5466 132
rect 5826 92 5866 132
rect 6226 92 6266 132
rect 6585 90 6625 136
<< metal1 >>
rect 2200 136 6750 150
rect 2200 132 6585 136
rect 1613 100 1687 106
rect 1613 50 1625 100
rect 1675 50 1687 100
rect 1813 100 1887 106
rect 1813 50 1825 100
rect 1875 50 1887 100
rect 2038 100 2112 106
rect 2038 50 2050 100
rect 2100 50 2112 100
rect 2200 100 2626 132
rect 2200 50 2400 100
rect 2614 92 2626 100
rect 2666 100 3026 132
rect 2666 92 2678 100
rect 2614 86 2678 92
rect 3014 92 3026 100
rect 3066 100 3426 132
rect 3066 92 3078 100
rect 3014 86 3078 92
rect 3414 92 3426 100
rect 3466 100 3826 132
rect 3466 92 3478 100
rect 3414 86 3478 92
rect 3814 92 3826 100
rect 3866 100 4226 132
rect 3866 92 3878 100
rect 3814 86 3878 92
rect 4214 92 4226 100
rect 4266 100 5026 132
rect 4266 92 4278 100
rect 4214 86 4278 92
rect 5014 92 5026 100
rect 5066 100 5426 132
rect 5066 92 5078 100
rect 5014 86 5078 92
rect 5414 92 5426 100
rect 5466 100 5826 132
rect 5466 92 5478 100
rect 5414 86 5478 92
rect 5814 92 5826 100
rect 5866 100 6226 132
rect 5866 92 5878 100
rect 5814 86 5878 92
rect 6214 92 6226 100
rect 6266 100 6585 132
rect 6266 92 6278 100
rect 6214 86 6278 92
rect 6569 90 6585 100
rect 6625 100 6750 136
rect 6625 90 6644 100
rect 6569 83 6644 90
rect 1600 -50 2400 50
rect 2500 -50 3450 50
rect 3550 -50 4650 50
rect 4800 -50 5750 50
rect 5850 -50 6800 50
rect 1600 -500 4542 -400
rect 1650 -650 1850 -600
rect 1650 -750 1750 -650
rect 4590 -750 4600 -650
rect 4700 -750 6700 -650
rect 1650 -800 1850 -750
rect 1700 -1250 1950 -1150
rect 2650 -1250 6700 -1150
rect 1850 -1300 1950 -1250
rect 1850 -1400 2300 -1300
rect 2400 -1400 2410 -1300
rect 4550 -1400 4750 -1250
rect 1800 -1500 1950 -1400
rect 3450 -1500 5850 -1400
rect 1700 -1950 1722 -1850
rect 2290 -1900 2300 -1800
rect 2400 -1900 4416 -1800
rect 1686 -2100 1766 -2000
rect 1866 -2100 1940 -2000
rect 4590 -2100 4600 -2000
rect 4700 -2100 5700 -2000
rect 2200 -2600 2400 -2550
rect 5750 -2600 5950 -2550
rect 1700 -2700 2400 -2600
rect 3440 -2700 3450 -2600
rect 3550 -2700 4500 -2600
rect 4700 -2700 5750 -2600
rect 5850 -2700 5950 -2600
rect 2200 -2750 2400 -2700
rect 5750 -2750 5950 -2700
<< via1 >>
rect 3450 -50 3550 50
rect 5750 -50 5850 50
rect 1750 -750 1850 -650
rect 4600 -750 4700 -650
rect 2300 -1400 2400 -1300
rect 2300 -1900 2400 -1800
rect 1766 -2100 1866 -2000
rect 4600 -2100 4700 -2000
rect 3450 -2700 3550 -2600
rect 5750 -2700 5850 -2600
<< metal2 >>
rect 3450 50 3550 60
rect 1750 -650 1850 -640
rect 2300 -650 2400 -628
rect 1850 -750 1866 -652
rect 1750 -760 1866 -750
rect 1766 -2000 1866 -760
rect 2300 -1300 2400 -750
rect 2300 -1800 2400 -1400
rect 2300 -1910 2400 -1900
rect 1766 -2110 1866 -2100
rect 3450 -2600 3550 -50
rect 5750 50 5850 60
rect 4600 -650 4700 -640
rect 4600 -760 4700 -750
rect 4600 -2000 4700 -1990
rect 4600 -2110 4700 -2100
rect 3450 -2710 3550 -2700
rect 5750 -2600 5850 -50
rect 5750 -2710 5850 -2700
<< via2 >>
rect 2300 -750 2400 -650
rect 1766 -2100 1866 -2000
rect 4600 -750 4700 -650
rect 4600 -2100 4700 -2000
<< metal3 >>
rect 2290 -650 2410 -645
rect 4590 -650 4710 -645
rect 2290 -750 2300 -650
rect 2400 -750 4600 -650
rect 4700 -750 4710 -650
rect 2290 -755 2410 -750
rect 4590 -755 4710 -750
rect 1756 -2000 1876 -1995
rect 4590 -2000 4710 -1995
rect 1756 -2100 1766 -2000
rect 1866 -2100 4600 -2000
rect 4700 -2100 4710 -2000
rect 1756 -2105 1876 -2100
rect 4590 -2105 4710 -2100
use sky130_fd_pr__nfet_01v8_6H2JYD  sky130_fd_pr__nfet_01v8_6H2JYD_0
timestamp 1710000826
transform 1 0 1813 0 1 -2040
box -263 -710 263 710
use sky130_fd_pr__pfet_01v8_UJHYGH  sky130_fd_pr__pfet_01v8_UJHYGH_0
timestamp 1709401415
transform 1 0 1859 0 1 -581
box -359 -719 359 719
use sky130_fd_pr__pfet_01v8_BDZ9JN  XM1
timestamp 1709390584
transform 1 0 3579 0 1 -581
box -1079 -719 1079 719
use sky130_fd_pr__nfet_01v8_KBNS5F  XM2
timestamp 1709392794
transform 1 0 4049 0 1 -2040
box -599 -710 599 710
use sky130_fd_pr__pfet_01v8_BDZ9JN  XM3
timestamp 1709390584
transform 1 0 5729 0 1 -581
box -1079 -719 1079 719
use sky130_fd_pr__nfet_01v8_KBNS5F  XM4
timestamp 1709392794
transform 1 0 5249 0 1 -2040
box -599 -710 599 710
<< labels >>
flabel metal1 2200 -2750 2400 -2550 0 FreeSans 256 0 0 0 VSS
port 4 nsew
flabel metal1 4550 -1350 4750 -1150 0 FreeSans 256 0 0 0 OUT
port 2 nsew
flabel metal1 5750 -2750 5950 -2550 0 FreeSans 256 0 0 0 VREF_N
port 5 nsew
flabel metal1 1650 -800 1850 -600 0 FreeSans 256 0 0 0 VIN
port 3 nsew
flabel metal1 2200 -50 2400 150 0 FreeSans 256 0 0 0 VDD
port 1 nsew
flabel metal1 4550 -50 4650 50 0 FreeSans 256 0 0 0 VREF_P
port 6 nsew
<< end >>
