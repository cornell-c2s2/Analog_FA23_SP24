magic
tech sky130A
magscale 1 2
timestamp 1716868724
<< pwell >>
rect -729 1502 729 1588
rect -729 -1502 -643 1502
rect 643 -1502 729 1502
rect -729 -1588 729 -1502
<< psubdiff >>
rect -703 1528 -595 1562
rect -561 1528 -527 1562
rect -493 1528 -459 1562
rect -425 1528 -391 1562
rect -357 1528 -323 1562
rect -289 1528 -255 1562
rect -221 1528 -187 1562
rect -153 1528 -119 1562
rect -85 1528 -51 1562
rect -17 1528 17 1562
rect 51 1528 85 1562
rect 119 1528 153 1562
rect 187 1528 221 1562
rect 255 1528 289 1562
rect 323 1528 357 1562
rect 391 1528 425 1562
rect 459 1528 493 1562
rect 527 1528 561 1562
rect 595 1528 703 1562
rect -703 1445 -669 1528
rect 669 1445 703 1528
rect -703 1377 -669 1411
rect -703 1309 -669 1343
rect -703 1241 -669 1275
rect -703 1173 -669 1207
rect -703 1105 -669 1139
rect -703 1037 -669 1071
rect -703 969 -669 1003
rect -703 901 -669 935
rect -703 833 -669 867
rect -703 765 -669 799
rect -703 697 -669 731
rect -703 629 -669 663
rect -703 561 -669 595
rect -703 493 -669 527
rect -703 425 -669 459
rect -703 357 -669 391
rect -703 289 -669 323
rect -703 221 -669 255
rect -703 153 -669 187
rect -703 85 -669 119
rect -703 17 -669 51
rect -703 -51 -669 -17
rect -703 -119 -669 -85
rect -703 -187 -669 -153
rect -703 -255 -669 -221
rect -703 -323 -669 -289
rect -703 -391 -669 -357
rect -703 -459 -669 -425
rect -703 -527 -669 -493
rect -703 -595 -669 -561
rect -703 -663 -669 -629
rect -703 -731 -669 -697
rect -703 -799 -669 -765
rect -703 -867 -669 -833
rect -703 -935 -669 -901
rect -703 -1003 -669 -969
rect -703 -1071 -669 -1037
rect -703 -1139 -669 -1105
rect -703 -1207 -669 -1173
rect -703 -1275 -669 -1241
rect -703 -1343 -669 -1309
rect -703 -1411 -669 -1377
rect 669 1377 703 1411
rect 669 1309 703 1343
rect 669 1241 703 1275
rect 669 1173 703 1207
rect 669 1105 703 1139
rect 669 1037 703 1071
rect 669 969 703 1003
rect 669 901 703 935
rect 669 833 703 867
rect 669 765 703 799
rect 669 697 703 731
rect 669 629 703 663
rect 669 561 703 595
rect 669 493 703 527
rect 669 425 703 459
rect 669 357 703 391
rect 669 289 703 323
rect 669 221 703 255
rect 669 153 703 187
rect 669 85 703 119
rect 669 17 703 51
rect 669 -51 703 -17
rect 669 -119 703 -85
rect 669 -187 703 -153
rect 669 -255 703 -221
rect 669 -323 703 -289
rect 669 -391 703 -357
rect 669 -459 703 -425
rect 669 -527 703 -493
rect 669 -595 703 -561
rect 669 -663 703 -629
rect 669 -731 703 -697
rect 669 -799 703 -765
rect 669 -867 703 -833
rect 669 -935 703 -901
rect 669 -1003 703 -969
rect 669 -1071 703 -1037
rect 669 -1139 703 -1105
rect 669 -1207 703 -1173
rect 669 -1275 703 -1241
rect 669 -1343 703 -1309
rect 669 -1411 703 -1377
rect -703 -1528 -669 -1445
rect 669 -1528 703 -1445
rect -703 -1562 -595 -1528
rect -561 -1562 -527 -1528
rect -493 -1562 -459 -1528
rect -425 -1562 -391 -1528
rect -357 -1562 -323 -1528
rect -289 -1562 -255 -1528
rect -221 -1562 -187 -1528
rect -153 -1562 -119 -1528
rect -85 -1562 -51 -1528
rect -17 -1562 17 -1528
rect 51 -1562 85 -1528
rect 119 -1562 153 -1528
rect 187 -1562 221 -1528
rect 255 -1562 289 -1528
rect 323 -1562 357 -1528
rect 391 -1562 425 -1528
rect 459 -1562 493 -1528
rect 527 -1562 561 -1528
rect 595 -1562 703 -1528
<< psubdiffcont >>
rect -595 1528 -561 1562
rect -527 1528 -493 1562
rect -459 1528 -425 1562
rect -391 1528 -357 1562
rect -323 1528 -289 1562
rect -255 1528 -221 1562
rect -187 1528 -153 1562
rect -119 1528 -85 1562
rect -51 1528 -17 1562
rect 17 1528 51 1562
rect 85 1528 119 1562
rect 153 1528 187 1562
rect 221 1528 255 1562
rect 289 1528 323 1562
rect 357 1528 391 1562
rect 425 1528 459 1562
rect 493 1528 527 1562
rect 561 1528 595 1562
rect -703 1411 -669 1445
rect -703 1343 -669 1377
rect -703 1275 -669 1309
rect -703 1207 -669 1241
rect -703 1139 -669 1173
rect -703 1071 -669 1105
rect -703 1003 -669 1037
rect -703 935 -669 969
rect -703 867 -669 901
rect -703 799 -669 833
rect -703 731 -669 765
rect -703 663 -669 697
rect -703 595 -669 629
rect -703 527 -669 561
rect -703 459 -669 493
rect -703 391 -669 425
rect -703 323 -669 357
rect -703 255 -669 289
rect -703 187 -669 221
rect -703 119 -669 153
rect -703 51 -669 85
rect -703 -17 -669 17
rect -703 -85 -669 -51
rect -703 -153 -669 -119
rect -703 -221 -669 -187
rect -703 -289 -669 -255
rect -703 -357 -669 -323
rect -703 -425 -669 -391
rect -703 -493 -669 -459
rect -703 -561 -669 -527
rect -703 -629 -669 -595
rect -703 -697 -669 -663
rect -703 -765 -669 -731
rect -703 -833 -669 -799
rect -703 -901 -669 -867
rect -703 -969 -669 -935
rect -703 -1037 -669 -1003
rect -703 -1105 -669 -1071
rect -703 -1173 -669 -1139
rect -703 -1241 -669 -1207
rect -703 -1309 -669 -1275
rect -703 -1377 -669 -1343
rect -703 -1445 -669 -1411
rect 669 1411 703 1445
rect 669 1343 703 1377
rect 669 1275 703 1309
rect 669 1207 703 1241
rect 669 1139 703 1173
rect 669 1071 703 1105
rect 669 1003 703 1037
rect 669 935 703 969
rect 669 867 703 901
rect 669 799 703 833
rect 669 731 703 765
rect 669 663 703 697
rect 669 595 703 629
rect 669 527 703 561
rect 669 459 703 493
rect 669 391 703 425
rect 669 323 703 357
rect 669 255 703 289
rect 669 187 703 221
rect 669 119 703 153
rect 669 51 703 85
rect 669 -17 703 17
rect 669 -85 703 -51
rect 669 -153 703 -119
rect 669 -221 703 -187
rect 669 -289 703 -255
rect 669 -357 703 -323
rect 669 -425 703 -391
rect 669 -493 703 -459
rect 669 -561 703 -527
rect 669 -629 703 -595
rect 669 -697 703 -663
rect 669 -765 703 -731
rect 669 -833 703 -799
rect 669 -901 703 -867
rect 669 -969 703 -935
rect 669 -1037 703 -1003
rect 669 -1105 703 -1071
rect 669 -1173 703 -1139
rect 669 -1241 703 -1207
rect 669 -1309 703 -1275
rect 669 -1377 703 -1343
rect 669 -1445 703 -1411
rect -595 -1562 -561 -1528
rect -527 -1562 -493 -1528
rect -459 -1562 -425 -1528
rect -391 -1562 -357 -1528
rect -323 -1562 -289 -1528
rect -255 -1562 -221 -1528
rect -187 -1562 -153 -1528
rect -119 -1562 -85 -1528
rect -51 -1562 -17 -1528
rect 17 -1562 51 -1528
rect 85 -1562 119 -1528
rect 153 -1562 187 -1528
rect 221 -1562 255 -1528
rect 289 -1562 323 -1528
rect 357 -1562 391 -1528
rect 425 -1562 459 -1528
rect 493 -1562 527 -1528
rect 561 -1562 595 -1528
<< xpolycontact >>
rect -573 1000 573 1432
rect -573 -1432 573 -1000
<< xpolyres >>
rect -573 -1000 573 1000
<< locali >>
rect -703 1528 -595 1562
rect -561 1528 -527 1562
rect -493 1528 -459 1562
rect -425 1528 -391 1562
rect -357 1528 -323 1562
rect -289 1528 -255 1562
rect -221 1528 -187 1562
rect -153 1528 -119 1562
rect -85 1528 -51 1562
rect -17 1528 17 1562
rect 51 1528 85 1562
rect 119 1528 153 1562
rect 187 1528 221 1562
rect 255 1528 289 1562
rect 323 1528 357 1562
rect 391 1528 425 1562
rect 459 1528 493 1562
rect 527 1528 561 1562
rect 595 1528 703 1562
rect -703 1445 -669 1528
rect 669 1445 703 1528
rect -703 1377 -669 1411
rect -703 1309 -669 1343
rect -703 1241 -669 1275
rect -703 1173 -669 1207
rect -703 1105 -669 1139
rect -703 1037 -669 1071
rect -703 969 -669 1003
rect 669 1377 703 1411
rect 669 1309 703 1343
rect 669 1241 703 1275
rect 669 1173 703 1207
rect 669 1105 703 1139
rect 669 1037 703 1071
rect -703 901 -669 935
rect -703 833 -669 867
rect -703 765 -669 799
rect -703 697 -669 731
rect -703 629 -669 663
rect -703 561 -669 595
rect -703 493 -669 527
rect -703 425 -669 459
rect -703 357 -669 391
rect -703 289 -669 323
rect -703 221 -669 255
rect -703 153 -669 187
rect -703 85 -669 119
rect -703 17 -669 51
rect -703 -51 -669 -17
rect -703 -119 -669 -85
rect -703 -187 -669 -153
rect -703 -255 -669 -221
rect -703 -323 -669 -289
rect -703 -391 -669 -357
rect -703 -459 -669 -425
rect -703 -527 -669 -493
rect -703 -595 -669 -561
rect -703 -663 -669 -629
rect -703 -731 -669 -697
rect -703 -799 -669 -765
rect -703 -867 -669 -833
rect -703 -935 -669 -901
rect -703 -1003 -669 -969
rect 669 969 703 1003
rect 669 901 703 935
rect 669 833 703 867
rect 669 765 703 799
rect 669 697 703 731
rect 669 629 703 663
rect 669 561 703 595
rect 669 493 703 527
rect 669 425 703 459
rect 669 357 703 391
rect 669 289 703 323
rect 669 221 703 255
rect 669 153 703 187
rect 669 85 703 119
rect 669 17 703 51
rect 669 -51 703 -17
rect 669 -119 703 -85
rect 669 -187 703 -153
rect 669 -255 703 -221
rect 669 -323 703 -289
rect 669 -391 703 -357
rect 669 -459 703 -425
rect 669 -527 703 -493
rect 669 -595 703 -561
rect 669 -663 703 -629
rect 669 -731 703 -697
rect 669 -799 703 -765
rect 669 -867 703 -833
rect 669 -935 703 -901
rect -703 -1071 -669 -1037
rect -703 -1139 -669 -1105
rect -703 -1207 -669 -1173
rect -703 -1275 -669 -1241
rect -703 -1343 -669 -1309
rect -703 -1411 -669 -1377
rect 669 -1003 703 -969
rect 669 -1071 703 -1037
rect 669 -1139 703 -1105
rect 669 -1207 703 -1173
rect 669 -1275 703 -1241
rect 669 -1343 703 -1309
rect 669 -1411 703 -1377
rect -703 -1528 -669 -1445
rect 669 -1528 703 -1445
rect -703 -1562 -595 -1528
rect -561 -1562 -527 -1528
rect -493 -1562 -459 -1528
rect -425 -1562 -391 -1528
rect -357 -1562 -323 -1528
rect -289 -1562 -255 -1528
rect -221 -1562 -187 -1528
rect -153 -1562 -119 -1528
rect -85 -1562 -51 -1528
rect -17 -1562 17 -1528
rect 51 -1562 85 -1528
rect 119 -1562 153 -1528
rect 187 -1562 221 -1528
rect 255 -1562 289 -1528
rect 323 -1562 357 -1528
rect 391 -1562 425 -1528
rect 459 -1562 493 -1528
rect 527 -1562 561 -1528
rect 595 -1562 703 -1528
<< viali >>
rect -557 1018 557 1412
rect -557 -1413 557 -1019
<< metal1 >>
rect -569 1412 569 1420
rect -569 1018 -557 1412
rect 557 1018 569 1412
rect -569 1011 569 1018
rect -569 -1019 569 -1011
rect -569 -1413 -557 -1019
rect 557 -1413 569 -1019
rect -569 -1420 569 -1413
<< properties >>
string FIXED_BBOX -686 -1545 686 1545
<< end >>
