magic
tech sky130A
magscale 1 2
timestamp 1716868724
<< pwell >>
rect -1963 -700 1963 700
<< nmos >>
rect -1777 -500 -1577 500
rect -1519 -500 -1319 500
rect -1261 -500 -1061 500
rect -1003 -500 -803 500
rect -745 -500 -545 500
rect -487 -500 -287 500
rect -229 -500 -29 500
rect 29 -500 229 500
rect 287 -500 487 500
rect 545 -500 745 500
rect 803 -500 1003 500
rect 1061 -500 1261 500
rect 1319 -500 1519 500
rect 1577 -500 1777 500
<< ndiff >>
rect -1835 459 -1777 500
rect -1835 425 -1823 459
rect -1789 425 -1777 459
rect -1835 391 -1777 425
rect -1835 357 -1823 391
rect -1789 357 -1777 391
rect -1835 323 -1777 357
rect -1835 289 -1823 323
rect -1789 289 -1777 323
rect -1835 255 -1777 289
rect -1835 221 -1823 255
rect -1789 221 -1777 255
rect -1835 187 -1777 221
rect -1835 153 -1823 187
rect -1789 153 -1777 187
rect -1835 119 -1777 153
rect -1835 85 -1823 119
rect -1789 85 -1777 119
rect -1835 51 -1777 85
rect -1835 17 -1823 51
rect -1789 17 -1777 51
rect -1835 -17 -1777 17
rect -1835 -51 -1823 -17
rect -1789 -51 -1777 -17
rect -1835 -85 -1777 -51
rect -1835 -119 -1823 -85
rect -1789 -119 -1777 -85
rect -1835 -153 -1777 -119
rect -1835 -187 -1823 -153
rect -1789 -187 -1777 -153
rect -1835 -221 -1777 -187
rect -1835 -255 -1823 -221
rect -1789 -255 -1777 -221
rect -1835 -289 -1777 -255
rect -1835 -323 -1823 -289
rect -1789 -323 -1777 -289
rect -1835 -357 -1777 -323
rect -1835 -391 -1823 -357
rect -1789 -391 -1777 -357
rect -1835 -425 -1777 -391
rect -1835 -459 -1823 -425
rect -1789 -459 -1777 -425
rect -1835 -500 -1777 -459
rect -1577 459 -1519 500
rect -1577 425 -1565 459
rect -1531 425 -1519 459
rect -1577 391 -1519 425
rect -1577 357 -1565 391
rect -1531 357 -1519 391
rect -1577 323 -1519 357
rect -1577 289 -1565 323
rect -1531 289 -1519 323
rect -1577 255 -1519 289
rect -1577 221 -1565 255
rect -1531 221 -1519 255
rect -1577 187 -1519 221
rect -1577 153 -1565 187
rect -1531 153 -1519 187
rect -1577 119 -1519 153
rect -1577 85 -1565 119
rect -1531 85 -1519 119
rect -1577 51 -1519 85
rect -1577 17 -1565 51
rect -1531 17 -1519 51
rect -1577 -17 -1519 17
rect -1577 -51 -1565 -17
rect -1531 -51 -1519 -17
rect -1577 -85 -1519 -51
rect -1577 -119 -1565 -85
rect -1531 -119 -1519 -85
rect -1577 -153 -1519 -119
rect -1577 -187 -1565 -153
rect -1531 -187 -1519 -153
rect -1577 -221 -1519 -187
rect -1577 -255 -1565 -221
rect -1531 -255 -1519 -221
rect -1577 -289 -1519 -255
rect -1577 -323 -1565 -289
rect -1531 -323 -1519 -289
rect -1577 -357 -1519 -323
rect -1577 -391 -1565 -357
rect -1531 -391 -1519 -357
rect -1577 -425 -1519 -391
rect -1577 -459 -1565 -425
rect -1531 -459 -1519 -425
rect -1577 -500 -1519 -459
rect -1319 459 -1261 500
rect -1319 425 -1307 459
rect -1273 425 -1261 459
rect -1319 391 -1261 425
rect -1319 357 -1307 391
rect -1273 357 -1261 391
rect -1319 323 -1261 357
rect -1319 289 -1307 323
rect -1273 289 -1261 323
rect -1319 255 -1261 289
rect -1319 221 -1307 255
rect -1273 221 -1261 255
rect -1319 187 -1261 221
rect -1319 153 -1307 187
rect -1273 153 -1261 187
rect -1319 119 -1261 153
rect -1319 85 -1307 119
rect -1273 85 -1261 119
rect -1319 51 -1261 85
rect -1319 17 -1307 51
rect -1273 17 -1261 51
rect -1319 -17 -1261 17
rect -1319 -51 -1307 -17
rect -1273 -51 -1261 -17
rect -1319 -85 -1261 -51
rect -1319 -119 -1307 -85
rect -1273 -119 -1261 -85
rect -1319 -153 -1261 -119
rect -1319 -187 -1307 -153
rect -1273 -187 -1261 -153
rect -1319 -221 -1261 -187
rect -1319 -255 -1307 -221
rect -1273 -255 -1261 -221
rect -1319 -289 -1261 -255
rect -1319 -323 -1307 -289
rect -1273 -323 -1261 -289
rect -1319 -357 -1261 -323
rect -1319 -391 -1307 -357
rect -1273 -391 -1261 -357
rect -1319 -425 -1261 -391
rect -1319 -459 -1307 -425
rect -1273 -459 -1261 -425
rect -1319 -500 -1261 -459
rect -1061 459 -1003 500
rect -1061 425 -1049 459
rect -1015 425 -1003 459
rect -1061 391 -1003 425
rect -1061 357 -1049 391
rect -1015 357 -1003 391
rect -1061 323 -1003 357
rect -1061 289 -1049 323
rect -1015 289 -1003 323
rect -1061 255 -1003 289
rect -1061 221 -1049 255
rect -1015 221 -1003 255
rect -1061 187 -1003 221
rect -1061 153 -1049 187
rect -1015 153 -1003 187
rect -1061 119 -1003 153
rect -1061 85 -1049 119
rect -1015 85 -1003 119
rect -1061 51 -1003 85
rect -1061 17 -1049 51
rect -1015 17 -1003 51
rect -1061 -17 -1003 17
rect -1061 -51 -1049 -17
rect -1015 -51 -1003 -17
rect -1061 -85 -1003 -51
rect -1061 -119 -1049 -85
rect -1015 -119 -1003 -85
rect -1061 -153 -1003 -119
rect -1061 -187 -1049 -153
rect -1015 -187 -1003 -153
rect -1061 -221 -1003 -187
rect -1061 -255 -1049 -221
rect -1015 -255 -1003 -221
rect -1061 -289 -1003 -255
rect -1061 -323 -1049 -289
rect -1015 -323 -1003 -289
rect -1061 -357 -1003 -323
rect -1061 -391 -1049 -357
rect -1015 -391 -1003 -357
rect -1061 -425 -1003 -391
rect -1061 -459 -1049 -425
rect -1015 -459 -1003 -425
rect -1061 -500 -1003 -459
rect -803 459 -745 500
rect -803 425 -791 459
rect -757 425 -745 459
rect -803 391 -745 425
rect -803 357 -791 391
rect -757 357 -745 391
rect -803 323 -745 357
rect -803 289 -791 323
rect -757 289 -745 323
rect -803 255 -745 289
rect -803 221 -791 255
rect -757 221 -745 255
rect -803 187 -745 221
rect -803 153 -791 187
rect -757 153 -745 187
rect -803 119 -745 153
rect -803 85 -791 119
rect -757 85 -745 119
rect -803 51 -745 85
rect -803 17 -791 51
rect -757 17 -745 51
rect -803 -17 -745 17
rect -803 -51 -791 -17
rect -757 -51 -745 -17
rect -803 -85 -745 -51
rect -803 -119 -791 -85
rect -757 -119 -745 -85
rect -803 -153 -745 -119
rect -803 -187 -791 -153
rect -757 -187 -745 -153
rect -803 -221 -745 -187
rect -803 -255 -791 -221
rect -757 -255 -745 -221
rect -803 -289 -745 -255
rect -803 -323 -791 -289
rect -757 -323 -745 -289
rect -803 -357 -745 -323
rect -803 -391 -791 -357
rect -757 -391 -745 -357
rect -803 -425 -745 -391
rect -803 -459 -791 -425
rect -757 -459 -745 -425
rect -803 -500 -745 -459
rect -545 459 -487 500
rect -545 425 -533 459
rect -499 425 -487 459
rect -545 391 -487 425
rect -545 357 -533 391
rect -499 357 -487 391
rect -545 323 -487 357
rect -545 289 -533 323
rect -499 289 -487 323
rect -545 255 -487 289
rect -545 221 -533 255
rect -499 221 -487 255
rect -545 187 -487 221
rect -545 153 -533 187
rect -499 153 -487 187
rect -545 119 -487 153
rect -545 85 -533 119
rect -499 85 -487 119
rect -545 51 -487 85
rect -545 17 -533 51
rect -499 17 -487 51
rect -545 -17 -487 17
rect -545 -51 -533 -17
rect -499 -51 -487 -17
rect -545 -85 -487 -51
rect -545 -119 -533 -85
rect -499 -119 -487 -85
rect -545 -153 -487 -119
rect -545 -187 -533 -153
rect -499 -187 -487 -153
rect -545 -221 -487 -187
rect -545 -255 -533 -221
rect -499 -255 -487 -221
rect -545 -289 -487 -255
rect -545 -323 -533 -289
rect -499 -323 -487 -289
rect -545 -357 -487 -323
rect -545 -391 -533 -357
rect -499 -391 -487 -357
rect -545 -425 -487 -391
rect -545 -459 -533 -425
rect -499 -459 -487 -425
rect -545 -500 -487 -459
rect -287 459 -229 500
rect -287 425 -275 459
rect -241 425 -229 459
rect -287 391 -229 425
rect -287 357 -275 391
rect -241 357 -229 391
rect -287 323 -229 357
rect -287 289 -275 323
rect -241 289 -229 323
rect -287 255 -229 289
rect -287 221 -275 255
rect -241 221 -229 255
rect -287 187 -229 221
rect -287 153 -275 187
rect -241 153 -229 187
rect -287 119 -229 153
rect -287 85 -275 119
rect -241 85 -229 119
rect -287 51 -229 85
rect -287 17 -275 51
rect -241 17 -229 51
rect -287 -17 -229 17
rect -287 -51 -275 -17
rect -241 -51 -229 -17
rect -287 -85 -229 -51
rect -287 -119 -275 -85
rect -241 -119 -229 -85
rect -287 -153 -229 -119
rect -287 -187 -275 -153
rect -241 -187 -229 -153
rect -287 -221 -229 -187
rect -287 -255 -275 -221
rect -241 -255 -229 -221
rect -287 -289 -229 -255
rect -287 -323 -275 -289
rect -241 -323 -229 -289
rect -287 -357 -229 -323
rect -287 -391 -275 -357
rect -241 -391 -229 -357
rect -287 -425 -229 -391
rect -287 -459 -275 -425
rect -241 -459 -229 -425
rect -287 -500 -229 -459
rect -29 459 29 500
rect -29 425 -17 459
rect 17 425 29 459
rect -29 391 29 425
rect -29 357 -17 391
rect 17 357 29 391
rect -29 323 29 357
rect -29 289 -17 323
rect 17 289 29 323
rect -29 255 29 289
rect -29 221 -17 255
rect 17 221 29 255
rect -29 187 29 221
rect -29 153 -17 187
rect 17 153 29 187
rect -29 119 29 153
rect -29 85 -17 119
rect 17 85 29 119
rect -29 51 29 85
rect -29 17 -17 51
rect 17 17 29 51
rect -29 -17 29 17
rect -29 -51 -17 -17
rect 17 -51 29 -17
rect -29 -85 29 -51
rect -29 -119 -17 -85
rect 17 -119 29 -85
rect -29 -153 29 -119
rect -29 -187 -17 -153
rect 17 -187 29 -153
rect -29 -221 29 -187
rect -29 -255 -17 -221
rect 17 -255 29 -221
rect -29 -289 29 -255
rect -29 -323 -17 -289
rect 17 -323 29 -289
rect -29 -357 29 -323
rect -29 -391 -17 -357
rect 17 -391 29 -357
rect -29 -425 29 -391
rect -29 -459 -17 -425
rect 17 -459 29 -425
rect -29 -500 29 -459
rect 229 459 287 500
rect 229 425 241 459
rect 275 425 287 459
rect 229 391 287 425
rect 229 357 241 391
rect 275 357 287 391
rect 229 323 287 357
rect 229 289 241 323
rect 275 289 287 323
rect 229 255 287 289
rect 229 221 241 255
rect 275 221 287 255
rect 229 187 287 221
rect 229 153 241 187
rect 275 153 287 187
rect 229 119 287 153
rect 229 85 241 119
rect 275 85 287 119
rect 229 51 287 85
rect 229 17 241 51
rect 275 17 287 51
rect 229 -17 287 17
rect 229 -51 241 -17
rect 275 -51 287 -17
rect 229 -85 287 -51
rect 229 -119 241 -85
rect 275 -119 287 -85
rect 229 -153 287 -119
rect 229 -187 241 -153
rect 275 -187 287 -153
rect 229 -221 287 -187
rect 229 -255 241 -221
rect 275 -255 287 -221
rect 229 -289 287 -255
rect 229 -323 241 -289
rect 275 -323 287 -289
rect 229 -357 287 -323
rect 229 -391 241 -357
rect 275 -391 287 -357
rect 229 -425 287 -391
rect 229 -459 241 -425
rect 275 -459 287 -425
rect 229 -500 287 -459
rect 487 459 545 500
rect 487 425 499 459
rect 533 425 545 459
rect 487 391 545 425
rect 487 357 499 391
rect 533 357 545 391
rect 487 323 545 357
rect 487 289 499 323
rect 533 289 545 323
rect 487 255 545 289
rect 487 221 499 255
rect 533 221 545 255
rect 487 187 545 221
rect 487 153 499 187
rect 533 153 545 187
rect 487 119 545 153
rect 487 85 499 119
rect 533 85 545 119
rect 487 51 545 85
rect 487 17 499 51
rect 533 17 545 51
rect 487 -17 545 17
rect 487 -51 499 -17
rect 533 -51 545 -17
rect 487 -85 545 -51
rect 487 -119 499 -85
rect 533 -119 545 -85
rect 487 -153 545 -119
rect 487 -187 499 -153
rect 533 -187 545 -153
rect 487 -221 545 -187
rect 487 -255 499 -221
rect 533 -255 545 -221
rect 487 -289 545 -255
rect 487 -323 499 -289
rect 533 -323 545 -289
rect 487 -357 545 -323
rect 487 -391 499 -357
rect 533 -391 545 -357
rect 487 -425 545 -391
rect 487 -459 499 -425
rect 533 -459 545 -425
rect 487 -500 545 -459
rect 745 459 803 500
rect 745 425 757 459
rect 791 425 803 459
rect 745 391 803 425
rect 745 357 757 391
rect 791 357 803 391
rect 745 323 803 357
rect 745 289 757 323
rect 791 289 803 323
rect 745 255 803 289
rect 745 221 757 255
rect 791 221 803 255
rect 745 187 803 221
rect 745 153 757 187
rect 791 153 803 187
rect 745 119 803 153
rect 745 85 757 119
rect 791 85 803 119
rect 745 51 803 85
rect 745 17 757 51
rect 791 17 803 51
rect 745 -17 803 17
rect 745 -51 757 -17
rect 791 -51 803 -17
rect 745 -85 803 -51
rect 745 -119 757 -85
rect 791 -119 803 -85
rect 745 -153 803 -119
rect 745 -187 757 -153
rect 791 -187 803 -153
rect 745 -221 803 -187
rect 745 -255 757 -221
rect 791 -255 803 -221
rect 745 -289 803 -255
rect 745 -323 757 -289
rect 791 -323 803 -289
rect 745 -357 803 -323
rect 745 -391 757 -357
rect 791 -391 803 -357
rect 745 -425 803 -391
rect 745 -459 757 -425
rect 791 -459 803 -425
rect 745 -500 803 -459
rect 1003 459 1061 500
rect 1003 425 1015 459
rect 1049 425 1061 459
rect 1003 391 1061 425
rect 1003 357 1015 391
rect 1049 357 1061 391
rect 1003 323 1061 357
rect 1003 289 1015 323
rect 1049 289 1061 323
rect 1003 255 1061 289
rect 1003 221 1015 255
rect 1049 221 1061 255
rect 1003 187 1061 221
rect 1003 153 1015 187
rect 1049 153 1061 187
rect 1003 119 1061 153
rect 1003 85 1015 119
rect 1049 85 1061 119
rect 1003 51 1061 85
rect 1003 17 1015 51
rect 1049 17 1061 51
rect 1003 -17 1061 17
rect 1003 -51 1015 -17
rect 1049 -51 1061 -17
rect 1003 -85 1061 -51
rect 1003 -119 1015 -85
rect 1049 -119 1061 -85
rect 1003 -153 1061 -119
rect 1003 -187 1015 -153
rect 1049 -187 1061 -153
rect 1003 -221 1061 -187
rect 1003 -255 1015 -221
rect 1049 -255 1061 -221
rect 1003 -289 1061 -255
rect 1003 -323 1015 -289
rect 1049 -323 1061 -289
rect 1003 -357 1061 -323
rect 1003 -391 1015 -357
rect 1049 -391 1061 -357
rect 1003 -425 1061 -391
rect 1003 -459 1015 -425
rect 1049 -459 1061 -425
rect 1003 -500 1061 -459
rect 1261 459 1319 500
rect 1261 425 1273 459
rect 1307 425 1319 459
rect 1261 391 1319 425
rect 1261 357 1273 391
rect 1307 357 1319 391
rect 1261 323 1319 357
rect 1261 289 1273 323
rect 1307 289 1319 323
rect 1261 255 1319 289
rect 1261 221 1273 255
rect 1307 221 1319 255
rect 1261 187 1319 221
rect 1261 153 1273 187
rect 1307 153 1319 187
rect 1261 119 1319 153
rect 1261 85 1273 119
rect 1307 85 1319 119
rect 1261 51 1319 85
rect 1261 17 1273 51
rect 1307 17 1319 51
rect 1261 -17 1319 17
rect 1261 -51 1273 -17
rect 1307 -51 1319 -17
rect 1261 -85 1319 -51
rect 1261 -119 1273 -85
rect 1307 -119 1319 -85
rect 1261 -153 1319 -119
rect 1261 -187 1273 -153
rect 1307 -187 1319 -153
rect 1261 -221 1319 -187
rect 1261 -255 1273 -221
rect 1307 -255 1319 -221
rect 1261 -289 1319 -255
rect 1261 -323 1273 -289
rect 1307 -323 1319 -289
rect 1261 -357 1319 -323
rect 1261 -391 1273 -357
rect 1307 -391 1319 -357
rect 1261 -425 1319 -391
rect 1261 -459 1273 -425
rect 1307 -459 1319 -425
rect 1261 -500 1319 -459
rect 1519 459 1577 500
rect 1519 425 1531 459
rect 1565 425 1577 459
rect 1519 391 1577 425
rect 1519 357 1531 391
rect 1565 357 1577 391
rect 1519 323 1577 357
rect 1519 289 1531 323
rect 1565 289 1577 323
rect 1519 255 1577 289
rect 1519 221 1531 255
rect 1565 221 1577 255
rect 1519 187 1577 221
rect 1519 153 1531 187
rect 1565 153 1577 187
rect 1519 119 1577 153
rect 1519 85 1531 119
rect 1565 85 1577 119
rect 1519 51 1577 85
rect 1519 17 1531 51
rect 1565 17 1577 51
rect 1519 -17 1577 17
rect 1519 -51 1531 -17
rect 1565 -51 1577 -17
rect 1519 -85 1577 -51
rect 1519 -119 1531 -85
rect 1565 -119 1577 -85
rect 1519 -153 1577 -119
rect 1519 -187 1531 -153
rect 1565 -187 1577 -153
rect 1519 -221 1577 -187
rect 1519 -255 1531 -221
rect 1565 -255 1577 -221
rect 1519 -289 1577 -255
rect 1519 -323 1531 -289
rect 1565 -323 1577 -289
rect 1519 -357 1577 -323
rect 1519 -391 1531 -357
rect 1565 -391 1577 -357
rect 1519 -425 1577 -391
rect 1519 -459 1531 -425
rect 1565 -459 1577 -425
rect 1519 -500 1577 -459
rect 1777 459 1835 500
rect 1777 425 1789 459
rect 1823 425 1835 459
rect 1777 391 1835 425
rect 1777 357 1789 391
rect 1823 357 1835 391
rect 1777 323 1835 357
rect 1777 289 1789 323
rect 1823 289 1835 323
rect 1777 255 1835 289
rect 1777 221 1789 255
rect 1823 221 1835 255
rect 1777 187 1835 221
rect 1777 153 1789 187
rect 1823 153 1835 187
rect 1777 119 1835 153
rect 1777 85 1789 119
rect 1823 85 1835 119
rect 1777 51 1835 85
rect 1777 17 1789 51
rect 1823 17 1835 51
rect 1777 -17 1835 17
rect 1777 -51 1789 -17
rect 1823 -51 1835 -17
rect 1777 -85 1835 -51
rect 1777 -119 1789 -85
rect 1823 -119 1835 -85
rect 1777 -153 1835 -119
rect 1777 -187 1789 -153
rect 1823 -187 1835 -153
rect 1777 -221 1835 -187
rect 1777 -255 1789 -221
rect 1823 -255 1835 -221
rect 1777 -289 1835 -255
rect 1777 -323 1789 -289
rect 1823 -323 1835 -289
rect 1777 -357 1835 -323
rect 1777 -391 1789 -357
rect 1823 -391 1835 -357
rect 1777 -425 1835 -391
rect 1777 -459 1789 -425
rect 1823 -459 1835 -425
rect 1777 -500 1835 -459
<< ndiffc >>
rect -1823 425 -1789 459
rect -1823 357 -1789 391
rect -1823 289 -1789 323
rect -1823 221 -1789 255
rect -1823 153 -1789 187
rect -1823 85 -1789 119
rect -1823 17 -1789 51
rect -1823 -51 -1789 -17
rect -1823 -119 -1789 -85
rect -1823 -187 -1789 -153
rect -1823 -255 -1789 -221
rect -1823 -323 -1789 -289
rect -1823 -391 -1789 -357
rect -1823 -459 -1789 -425
rect -1565 425 -1531 459
rect -1565 357 -1531 391
rect -1565 289 -1531 323
rect -1565 221 -1531 255
rect -1565 153 -1531 187
rect -1565 85 -1531 119
rect -1565 17 -1531 51
rect -1565 -51 -1531 -17
rect -1565 -119 -1531 -85
rect -1565 -187 -1531 -153
rect -1565 -255 -1531 -221
rect -1565 -323 -1531 -289
rect -1565 -391 -1531 -357
rect -1565 -459 -1531 -425
rect -1307 425 -1273 459
rect -1307 357 -1273 391
rect -1307 289 -1273 323
rect -1307 221 -1273 255
rect -1307 153 -1273 187
rect -1307 85 -1273 119
rect -1307 17 -1273 51
rect -1307 -51 -1273 -17
rect -1307 -119 -1273 -85
rect -1307 -187 -1273 -153
rect -1307 -255 -1273 -221
rect -1307 -323 -1273 -289
rect -1307 -391 -1273 -357
rect -1307 -459 -1273 -425
rect -1049 425 -1015 459
rect -1049 357 -1015 391
rect -1049 289 -1015 323
rect -1049 221 -1015 255
rect -1049 153 -1015 187
rect -1049 85 -1015 119
rect -1049 17 -1015 51
rect -1049 -51 -1015 -17
rect -1049 -119 -1015 -85
rect -1049 -187 -1015 -153
rect -1049 -255 -1015 -221
rect -1049 -323 -1015 -289
rect -1049 -391 -1015 -357
rect -1049 -459 -1015 -425
rect -791 425 -757 459
rect -791 357 -757 391
rect -791 289 -757 323
rect -791 221 -757 255
rect -791 153 -757 187
rect -791 85 -757 119
rect -791 17 -757 51
rect -791 -51 -757 -17
rect -791 -119 -757 -85
rect -791 -187 -757 -153
rect -791 -255 -757 -221
rect -791 -323 -757 -289
rect -791 -391 -757 -357
rect -791 -459 -757 -425
rect -533 425 -499 459
rect -533 357 -499 391
rect -533 289 -499 323
rect -533 221 -499 255
rect -533 153 -499 187
rect -533 85 -499 119
rect -533 17 -499 51
rect -533 -51 -499 -17
rect -533 -119 -499 -85
rect -533 -187 -499 -153
rect -533 -255 -499 -221
rect -533 -323 -499 -289
rect -533 -391 -499 -357
rect -533 -459 -499 -425
rect -275 425 -241 459
rect -275 357 -241 391
rect -275 289 -241 323
rect -275 221 -241 255
rect -275 153 -241 187
rect -275 85 -241 119
rect -275 17 -241 51
rect -275 -51 -241 -17
rect -275 -119 -241 -85
rect -275 -187 -241 -153
rect -275 -255 -241 -221
rect -275 -323 -241 -289
rect -275 -391 -241 -357
rect -275 -459 -241 -425
rect -17 425 17 459
rect -17 357 17 391
rect -17 289 17 323
rect -17 221 17 255
rect -17 153 17 187
rect -17 85 17 119
rect -17 17 17 51
rect -17 -51 17 -17
rect -17 -119 17 -85
rect -17 -187 17 -153
rect -17 -255 17 -221
rect -17 -323 17 -289
rect -17 -391 17 -357
rect -17 -459 17 -425
rect 241 425 275 459
rect 241 357 275 391
rect 241 289 275 323
rect 241 221 275 255
rect 241 153 275 187
rect 241 85 275 119
rect 241 17 275 51
rect 241 -51 275 -17
rect 241 -119 275 -85
rect 241 -187 275 -153
rect 241 -255 275 -221
rect 241 -323 275 -289
rect 241 -391 275 -357
rect 241 -459 275 -425
rect 499 425 533 459
rect 499 357 533 391
rect 499 289 533 323
rect 499 221 533 255
rect 499 153 533 187
rect 499 85 533 119
rect 499 17 533 51
rect 499 -51 533 -17
rect 499 -119 533 -85
rect 499 -187 533 -153
rect 499 -255 533 -221
rect 499 -323 533 -289
rect 499 -391 533 -357
rect 499 -459 533 -425
rect 757 425 791 459
rect 757 357 791 391
rect 757 289 791 323
rect 757 221 791 255
rect 757 153 791 187
rect 757 85 791 119
rect 757 17 791 51
rect 757 -51 791 -17
rect 757 -119 791 -85
rect 757 -187 791 -153
rect 757 -255 791 -221
rect 757 -323 791 -289
rect 757 -391 791 -357
rect 757 -459 791 -425
rect 1015 425 1049 459
rect 1015 357 1049 391
rect 1015 289 1049 323
rect 1015 221 1049 255
rect 1015 153 1049 187
rect 1015 85 1049 119
rect 1015 17 1049 51
rect 1015 -51 1049 -17
rect 1015 -119 1049 -85
rect 1015 -187 1049 -153
rect 1015 -255 1049 -221
rect 1015 -323 1049 -289
rect 1015 -391 1049 -357
rect 1015 -459 1049 -425
rect 1273 425 1307 459
rect 1273 357 1307 391
rect 1273 289 1307 323
rect 1273 221 1307 255
rect 1273 153 1307 187
rect 1273 85 1307 119
rect 1273 17 1307 51
rect 1273 -51 1307 -17
rect 1273 -119 1307 -85
rect 1273 -187 1307 -153
rect 1273 -255 1307 -221
rect 1273 -323 1307 -289
rect 1273 -391 1307 -357
rect 1273 -459 1307 -425
rect 1531 425 1565 459
rect 1531 357 1565 391
rect 1531 289 1565 323
rect 1531 221 1565 255
rect 1531 153 1565 187
rect 1531 85 1565 119
rect 1531 17 1565 51
rect 1531 -51 1565 -17
rect 1531 -119 1565 -85
rect 1531 -187 1565 -153
rect 1531 -255 1565 -221
rect 1531 -323 1565 -289
rect 1531 -391 1565 -357
rect 1531 -459 1565 -425
rect 1789 425 1823 459
rect 1789 357 1823 391
rect 1789 289 1823 323
rect 1789 221 1823 255
rect 1789 153 1823 187
rect 1789 85 1823 119
rect 1789 17 1823 51
rect 1789 -51 1823 -17
rect 1789 -119 1823 -85
rect 1789 -187 1823 -153
rect 1789 -255 1823 -221
rect 1789 -323 1823 -289
rect 1789 -391 1823 -357
rect 1789 -459 1823 -425
<< psubdiff >>
rect -1937 640 -1819 674
rect -1785 640 -1751 674
rect -1717 640 -1683 674
rect -1649 640 -1615 674
rect -1581 640 -1547 674
rect -1513 640 -1479 674
rect -1445 640 -1411 674
rect -1377 640 -1343 674
rect -1309 640 -1275 674
rect -1241 640 -1207 674
rect -1173 640 -1139 674
rect -1105 640 -1071 674
rect -1037 640 -1003 674
rect -969 640 -935 674
rect -901 640 -867 674
rect -833 640 -799 674
rect -765 640 -731 674
rect -697 640 -663 674
rect -629 640 -595 674
rect -561 640 -527 674
rect -493 640 -459 674
rect -425 640 -391 674
rect -357 640 -323 674
rect -289 640 -255 674
rect -221 640 -187 674
rect -153 640 -119 674
rect -85 640 -51 674
rect -17 640 17 674
rect 51 640 85 674
rect 119 640 153 674
rect 187 640 221 674
rect 255 640 289 674
rect 323 640 357 674
rect 391 640 425 674
rect 459 640 493 674
rect 527 640 561 674
rect 595 640 629 674
rect 663 640 697 674
rect 731 640 765 674
rect 799 640 833 674
rect 867 640 901 674
rect 935 640 969 674
rect 1003 640 1037 674
rect 1071 640 1105 674
rect 1139 640 1173 674
rect 1207 640 1241 674
rect 1275 640 1309 674
rect 1343 640 1377 674
rect 1411 640 1445 674
rect 1479 640 1513 674
rect 1547 640 1581 674
rect 1615 640 1649 674
rect 1683 640 1717 674
rect 1751 640 1785 674
rect 1819 640 1937 674
rect -1937 561 -1903 640
rect -1937 493 -1903 527
rect 1903 561 1937 640
rect -1937 425 -1903 459
rect -1937 357 -1903 391
rect -1937 289 -1903 323
rect -1937 221 -1903 255
rect -1937 153 -1903 187
rect -1937 85 -1903 119
rect -1937 17 -1903 51
rect -1937 -51 -1903 -17
rect -1937 -119 -1903 -85
rect -1937 -187 -1903 -153
rect -1937 -255 -1903 -221
rect -1937 -323 -1903 -289
rect -1937 -391 -1903 -357
rect -1937 -459 -1903 -425
rect -1937 -527 -1903 -493
rect 1903 493 1937 527
rect 1903 425 1937 459
rect 1903 357 1937 391
rect 1903 289 1937 323
rect 1903 221 1937 255
rect 1903 153 1937 187
rect 1903 85 1937 119
rect 1903 17 1937 51
rect 1903 -51 1937 -17
rect 1903 -119 1937 -85
rect 1903 -187 1937 -153
rect 1903 -255 1937 -221
rect 1903 -323 1937 -289
rect 1903 -391 1937 -357
rect 1903 -459 1937 -425
rect -1937 -640 -1903 -561
rect 1903 -527 1937 -493
rect 1903 -640 1937 -561
rect -1937 -674 -1819 -640
rect -1785 -674 -1751 -640
rect -1717 -674 -1683 -640
rect -1649 -674 -1615 -640
rect -1581 -674 -1547 -640
rect -1513 -674 -1479 -640
rect -1445 -674 -1411 -640
rect -1377 -674 -1343 -640
rect -1309 -674 -1275 -640
rect -1241 -674 -1207 -640
rect -1173 -674 -1139 -640
rect -1105 -674 -1071 -640
rect -1037 -674 -1003 -640
rect -969 -674 -935 -640
rect -901 -674 -867 -640
rect -833 -674 -799 -640
rect -765 -674 -731 -640
rect -697 -674 -663 -640
rect -629 -674 -595 -640
rect -561 -674 -527 -640
rect -493 -674 -459 -640
rect -425 -674 -391 -640
rect -357 -674 -323 -640
rect -289 -674 -255 -640
rect -221 -674 -187 -640
rect -153 -674 -119 -640
rect -85 -674 -51 -640
rect -17 -674 17 -640
rect 51 -674 85 -640
rect 119 -674 153 -640
rect 187 -674 221 -640
rect 255 -674 289 -640
rect 323 -674 357 -640
rect 391 -674 425 -640
rect 459 -674 493 -640
rect 527 -674 561 -640
rect 595 -674 629 -640
rect 663 -674 697 -640
rect 731 -674 765 -640
rect 799 -674 833 -640
rect 867 -674 901 -640
rect 935 -674 969 -640
rect 1003 -674 1037 -640
rect 1071 -674 1105 -640
rect 1139 -674 1173 -640
rect 1207 -674 1241 -640
rect 1275 -674 1309 -640
rect 1343 -674 1377 -640
rect 1411 -674 1445 -640
rect 1479 -674 1513 -640
rect 1547 -674 1581 -640
rect 1615 -674 1649 -640
rect 1683 -674 1717 -640
rect 1751 -674 1785 -640
rect 1819 -674 1937 -640
<< psubdiffcont >>
rect -1819 640 -1785 674
rect -1751 640 -1717 674
rect -1683 640 -1649 674
rect -1615 640 -1581 674
rect -1547 640 -1513 674
rect -1479 640 -1445 674
rect -1411 640 -1377 674
rect -1343 640 -1309 674
rect -1275 640 -1241 674
rect -1207 640 -1173 674
rect -1139 640 -1105 674
rect -1071 640 -1037 674
rect -1003 640 -969 674
rect -935 640 -901 674
rect -867 640 -833 674
rect -799 640 -765 674
rect -731 640 -697 674
rect -663 640 -629 674
rect -595 640 -561 674
rect -527 640 -493 674
rect -459 640 -425 674
rect -391 640 -357 674
rect -323 640 -289 674
rect -255 640 -221 674
rect -187 640 -153 674
rect -119 640 -85 674
rect -51 640 -17 674
rect 17 640 51 674
rect 85 640 119 674
rect 153 640 187 674
rect 221 640 255 674
rect 289 640 323 674
rect 357 640 391 674
rect 425 640 459 674
rect 493 640 527 674
rect 561 640 595 674
rect 629 640 663 674
rect 697 640 731 674
rect 765 640 799 674
rect 833 640 867 674
rect 901 640 935 674
rect 969 640 1003 674
rect 1037 640 1071 674
rect 1105 640 1139 674
rect 1173 640 1207 674
rect 1241 640 1275 674
rect 1309 640 1343 674
rect 1377 640 1411 674
rect 1445 640 1479 674
rect 1513 640 1547 674
rect 1581 640 1615 674
rect 1649 640 1683 674
rect 1717 640 1751 674
rect 1785 640 1819 674
rect -1937 527 -1903 561
rect 1903 527 1937 561
rect -1937 459 -1903 493
rect -1937 391 -1903 425
rect -1937 323 -1903 357
rect -1937 255 -1903 289
rect -1937 187 -1903 221
rect -1937 119 -1903 153
rect -1937 51 -1903 85
rect -1937 -17 -1903 17
rect -1937 -85 -1903 -51
rect -1937 -153 -1903 -119
rect -1937 -221 -1903 -187
rect -1937 -289 -1903 -255
rect -1937 -357 -1903 -323
rect -1937 -425 -1903 -391
rect -1937 -493 -1903 -459
rect 1903 459 1937 493
rect 1903 391 1937 425
rect 1903 323 1937 357
rect 1903 255 1937 289
rect 1903 187 1937 221
rect 1903 119 1937 153
rect 1903 51 1937 85
rect 1903 -17 1937 17
rect 1903 -85 1937 -51
rect 1903 -153 1937 -119
rect 1903 -221 1937 -187
rect 1903 -289 1937 -255
rect 1903 -357 1937 -323
rect 1903 -425 1937 -391
rect 1903 -493 1937 -459
rect -1937 -561 -1903 -527
rect 1903 -561 1937 -527
rect -1819 -674 -1785 -640
rect -1751 -674 -1717 -640
rect -1683 -674 -1649 -640
rect -1615 -674 -1581 -640
rect -1547 -674 -1513 -640
rect -1479 -674 -1445 -640
rect -1411 -674 -1377 -640
rect -1343 -674 -1309 -640
rect -1275 -674 -1241 -640
rect -1207 -674 -1173 -640
rect -1139 -674 -1105 -640
rect -1071 -674 -1037 -640
rect -1003 -674 -969 -640
rect -935 -674 -901 -640
rect -867 -674 -833 -640
rect -799 -674 -765 -640
rect -731 -674 -697 -640
rect -663 -674 -629 -640
rect -595 -674 -561 -640
rect -527 -674 -493 -640
rect -459 -674 -425 -640
rect -391 -674 -357 -640
rect -323 -674 -289 -640
rect -255 -674 -221 -640
rect -187 -674 -153 -640
rect -119 -674 -85 -640
rect -51 -674 -17 -640
rect 17 -674 51 -640
rect 85 -674 119 -640
rect 153 -674 187 -640
rect 221 -674 255 -640
rect 289 -674 323 -640
rect 357 -674 391 -640
rect 425 -674 459 -640
rect 493 -674 527 -640
rect 561 -674 595 -640
rect 629 -674 663 -640
rect 697 -674 731 -640
rect 765 -674 799 -640
rect 833 -674 867 -640
rect 901 -674 935 -640
rect 969 -674 1003 -640
rect 1037 -674 1071 -640
rect 1105 -674 1139 -640
rect 1173 -674 1207 -640
rect 1241 -674 1275 -640
rect 1309 -674 1343 -640
rect 1377 -674 1411 -640
rect 1445 -674 1479 -640
rect 1513 -674 1547 -640
rect 1581 -674 1615 -640
rect 1649 -674 1683 -640
rect 1717 -674 1751 -640
rect 1785 -674 1819 -640
<< poly >>
rect -1777 572 -1577 588
rect -1777 538 -1728 572
rect -1694 538 -1660 572
rect -1626 538 -1577 572
rect -1777 500 -1577 538
rect -1519 572 -1319 588
rect -1519 538 -1470 572
rect -1436 538 -1402 572
rect -1368 538 -1319 572
rect -1519 500 -1319 538
rect -1261 572 -1061 588
rect -1261 538 -1212 572
rect -1178 538 -1144 572
rect -1110 538 -1061 572
rect -1261 500 -1061 538
rect -1003 572 -803 588
rect -1003 538 -954 572
rect -920 538 -886 572
rect -852 538 -803 572
rect -1003 500 -803 538
rect -745 572 -545 588
rect -745 538 -696 572
rect -662 538 -628 572
rect -594 538 -545 572
rect -745 500 -545 538
rect -487 572 -287 588
rect -487 538 -438 572
rect -404 538 -370 572
rect -336 538 -287 572
rect -487 500 -287 538
rect -229 572 -29 588
rect -229 538 -180 572
rect -146 538 -112 572
rect -78 538 -29 572
rect -229 500 -29 538
rect 29 572 229 588
rect 29 538 78 572
rect 112 538 146 572
rect 180 538 229 572
rect 29 500 229 538
rect 287 572 487 588
rect 287 538 336 572
rect 370 538 404 572
rect 438 538 487 572
rect 287 500 487 538
rect 545 572 745 588
rect 545 538 594 572
rect 628 538 662 572
rect 696 538 745 572
rect 545 500 745 538
rect 803 572 1003 588
rect 803 538 852 572
rect 886 538 920 572
rect 954 538 1003 572
rect 803 500 1003 538
rect 1061 572 1261 588
rect 1061 538 1110 572
rect 1144 538 1178 572
rect 1212 538 1261 572
rect 1061 500 1261 538
rect 1319 572 1519 588
rect 1319 538 1368 572
rect 1402 538 1436 572
rect 1470 538 1519 572
rect 1319 500 1519 538
rect 1577 572 1777 588
rect 1577 538 1626 572
rect 1660 538 1694 572
rect 1728 538 1777 572
rect 1577 500 1777 538
rect -1777 -538 -1577 -500
rect -1777 -572 -1728 -538
rect -1694 -572 -1660 -538
rect -1626 -572 -1577 -538
rect -1777 -588 -1577 -572
rect -1519 -538 -1319 -500
rect -1519 -572 -1470 -538
rect -1436 -572 -1402 -538
rect -1368 -572 -1319 -538
rect -1519 -588 -1319 -572
rect -1261 -538 -1061 -500
rect -1261 -572 -1212 -538
rect -1178 -572 -1144 -538
rect -1110 -572 -1061 -538
rect -1261 -588 -1061 -572
rect -1003 -538 -803 -500
rect -1003 -572 -954 -538
rect -920 -572 -886 -538
rect -852 -572 -803 -538
rect -1003 -588 -803 -572
rect -745 -538 -545 -500
rect -745 -572 -696 -538
rect -662 -572 -628 -538
rect -594 -572 -545 -538
rect -745 -588 -545 -572
rect -487 -538 -287 -500
rect -487 -572 -438 -538
rect -404 -572 -370 -538
rect -336 -572 -287 -538
rect -487 -588 -287 -572
rect -229 -538 -29 -500
rect -229 -572 -180 -538
rect -146 -572 -112 -538
rect -78 -572 -29 -538
rect -229 -588 -29 -572
rect 29 -538 229 -500
rect 29 -572 78 -538
rect 112 -572 146 -538
rect 180 -572 229 -538
rect 29 -588 229 -572
rect 287 -538 487 -500
rect 287 -572 336 -538
rect 370 -572 404 -538
rect 438 -572 487 -538
rect 287 -588 487 -572
rect 545 -538 745 -500
rect 545 -572 594 -538
rect 628 -572 662 -538
rect 696 -572 745 -538
rect 545 -588 745 -572
rect 803 -538 1003 -500
rect 803 -572 852 -538
rect 886 -572 920 -538
rect 954 -572 1003 -538
rect 803 -588 1003 -572
rect 1061 -538 1261 -500
rect 1061 -572 1110 -538
rect 1144 -572 1178 -538
rect 1212 -572 1261 -538
rect 1061 -588 1261 -572
rect 1319 -538 1519 -500
rect 1319 -572 1368 -538
rect 1402 -572 1436 -538
rect 1470 -572 1519 -538
rect 1319 -588 1519 -572
rect 1577 -538 1777 -500
rect 1577 -572 1626 -538
rect 1660 -572 1694 -538
rect 1728 -572 1777 -538
rect 1577 -588 1777 -572
<< polycont >>
rect -1728 538 -1694 572
rect -1660 538 -1626 572
rect -1470 538 -1436 572
rect -1402 538 -1368 572
rect -1212 538 -1178 572
rect -1144 538 -1110 572
rect -954 538 -920 572
rect -886 538 -852 572
rect -696 538 -662 572
rect -628 538 -594 572
rect -438 538 -404 572
rect -370 538 -336 572
rect -180 538 -146 572
rect -112 538 -78 572
rect 78 538 112 572
rect 146 538 180 572
rect 336 538 370 572
rect 404 538 438 572
rect 594 538 628 572
rect 662 538 696 572
rect 852 538 886 572
rect 920 538 954 572
rect 1110 538 1144 572
rect 1178 538 1212 572
rect 1368 538 1402 572
rect 1436 538 1470 572
rect 1626 538 1660 572
rect 1694 538 1728 572
rect -1728 -572 -1694 -538
rect -1660 -572 -1626 -538
rect -1470 -572 -1436 -538
rect -1402 -572 -1368 -538
rect -1212 -572 -1178 -538
rect -1144 -572 -1110 -538
rect -954 -572 -920 -538
rect -886 -572 -852 -538
rect -696 -572 -662 -538
rect -628 -572 -594 -538
rect -438 -572 -404 -538
rect -370 -572 -336 -538
rect -180 -572 -146 -538
rect -112 -572 -78 -538
rect 78 -572 112 -538
rect 146 -572 180 -538
rect 336 -572 370 -538
rect 404 -572 438 -538
rect 594 -572 628 -538
rect 662 -572 696 -538
rect 852 -572 886 -538
rect 920 -572 954 -538
rect 1110 -572 1144 -538
rect 1178 -572 1212 -538
rect 1368 -572 1402 -538
rect 1436 -572 1470 -538
rect 1626 -572 1660 -538
rect 1694 -572 1728 -538
<< locali >>
rect -1937 640 -1819 674
rect -1785 640 -1751 674
rect -1717 640 -1683 674
rect -1649 640 -1615 674
rect -1581 640 -1547 674
rect -1513 640 -1479 674
rect -1445 640 -1411 674
rect -1377 640 -1343 674
rect -1309 640 -1275 674
rect -1241 640 -1207 674
rect -1173 640 -1139 674
rect -1105 640 -1071 674
rect -1037 640 -1003 674
rect -969 640 -935 674
rect -883 640 -867 674
rect -811 640 -799 674
rect -739 640 -731 674
rect -667 640 -663 674
rect -561 640 -557 674
rect -493 640 -485 674
rect -425 640 -413 674
rect -357 640 -341 674
rect -289 640 -269 674
rect -221 640 -197 674
rect -153 640 -125 674
rect -85 640 -53 674
rect -17 640 17 674
rect 53 640 85 674
rect 125 640 153 674
rect 197 640 221 674
rect 269 640 289 674
rect 341 640 357 674
rect 413 640 425 674
rect 485 640 493 674
rect 557 640 561 674
rect 663 640 667 674
rect 731 640 739 674
rect 799 640 811 674
rect 867 640 883 674
rect 935 640 969 674
rect 1003 640 1037 674
rect 1071 640 1105 674
rect 1139 640 1173 674
rect 1207 640 1241 674
rect 1275 640 1309 674
rect 1343 640 1377 674
rect 1411 640 1445 674
rect 1479 640 1513 674
rect 1547 640 1581 674
rect 1615 640 1649 674
rect 1683 640 1717 674
rect 1751 640 1785 674
rect 1819 640 1937 674
rect -1937 561 -1903 640
rect -1777 538 -1730 572
rect -1694 538 -1660 572
rect -1624 538 -1577 572
rect -1519 538 -1472 572
rect -1436 538 -1402 572
rect -1366 538 -1319 572
rect -1261 538 -1214 572
rect -1178 538 -1144 572
rect -1108 538 -1061 572
rect -1003 538 -956 572
rect -920 538 -886 572
rect -850 538 -803 572
rect -745 538 -698 572
rect -662 538 -628 572
rect -592 538 -545 572
rect -487 538 -440 572
rect -404 538 -370 572
rect -334 538 -287 572
rect -229 538 -182 572
rect -146 538 -112 572
rect -76 538 -29 572
rect 29 538 76 572
rect 112 538 146 572
rect 182 538 229 572
rect 287 538 334 572
rect 370 538 404 572
rect 440 538 487 572
rect 545 538 592 572
rect 628 538 662 572
rect 698 538 745 572
rect 803 538 850 572
rect 886 538 920 572
rect 956 538 1003 572
rect 1061 538 1108 572
rect 1144 538 1178 572
rect 1214 538 1261 572
rect 1319 538 1366 572
rect 1402 538 1436 572
rect 1472 538 1519 572
rect 1577 538 1624 572
rect 1660 538 1694 572
rect 1730 538 1777 572
rect 1903 561 1937 640
rect -1937 493 -1903 527
rect -1937 425 -1903 459
rect -1937 357 -1903 391
rect -1937 289 -1903 323
rect -1937 221 -1903 255
rect -1937 153 -1903 187
rect -1937 85 -1903 119
rect -1937 17 -1903 51
rect -1937 -51 -1903 -17
rect -1937 -119 -1903 -85
rect -1937 -187 -1903 -153
rect -1937 -255 -1903 -221
rect -1937 -323 -1903 -289
rect -1937 -391 -1903 -357
rect -1937 -459 -1903 -425
rect -1937 -527 -1903 -493
rect -1823 485 -1789 504
rect -1823 413 -1789 425
rect -1823 341 -1789 357
rect -1823 269 -1789 289
rect -1823 197 -1789 221
rect -1823 125 -1789 153
rect -1823 53 -1789 85
rect -1823 -17 -1789 17
rect -1823 -85 -1789 -53
rect -1823 -153 -1789 -125
rect -1823 -221 -1789 -197
rect -1823 -289 -1789 -269
rect -1823 -357 -1789 -341
rect -1823 -425 -1789 -413
rect -1823 -504 -1789 -485
rect -1565 485 -1531 504
rect -1565 413 -1531 425
rect -1565 341 -1531 357
rect -1565 269 -1531 289
rect -1565 197 -1531 221
rect -1565 125 -1531 153
rect -1565 53 -1531 85
rect -1565 -17 -1531 17
rect -1565 -85 -1531 -53
rect -1565 -153 -1531 -125
rect -1565 -221 -1531 -197
rect -1565 -289 -1531 -269
rect -1565 -357 -1531 -341
rect -1565 -425 -1531 -413
rect -1565 -504 -1531 -485
rect -1307 485 -1273 504
rect -1307 413 -1273 425
rect -1307 341 -1273 357
rect -1307 269 -1273 289
rect -1307 197 -1273 221
rect -1307 125 -1273 153
rect -1307 53 -1273 85
rect -1307 -17 -1273 17
rect -1307 -85 -1273 -53
rect -1307 -153 -1273 -125
rect -1307 -221 -1273 -197
rect -1307 -289 -1273 -269
rect -1307 -357 -1273 -341
rect -1307 -425 -1273 -413
rect -1307 -504 -1273 -485
rect -1049 485 -1015 504
rect -1049 413 -1015 425
rect -1049 341 -1015 357
rect -1049 269 -1015 289
rect -1049 197 -1015 221
rect -1049 125 -1015 153
rect -1049 53 -1015 85
rect -1049 -17 -1015 17
rect -1049 -85 -1015 -53
rect -1049 -153 -1015 -125
rect -1049 -221 -1015 -197
rect -1049 -289 -1015 -269
rect -1049 -357 -1015 -341
rect -1049 -425 -1015 -413
rect -1049 -504 -1015 -485
rect -791 485 -757 504
rect -791 413 -757 425
rect -791 341 -757 357
rect -791 269 -757 289
rect -791 197 -757 221
rect -791 125 -757 153
rect -791 53 -757 85
rect -791 -17 -757 17
rect -791 -85 -757 -53
rect -791 -153 -757 -125
rect -791 -221 -757 -197
rect -791 -289 -757 -269
rect -791 -357 -757 -341
rect -791 -425 -757 -413
rect -791 -504 -757 -485
rect -533 485 -499 504
rect -533 413 -499 425
rect -533 341 -499 357
rect -533 269 -499 289
rect -533 197 -499 221
rect -533 125 -499 153
rect -533 53 -499 85
rect -533 -17 -499 17
rect -533 -85 -499 -53
rect -533 -153 -499 -125
rect -533 -221 -499 -197
rect -533 -289 -499 -269
rect -533 -357 -499 -341
rect -533 -425 -499 -413
rect -533 -504 -499 -485
rect -275 485 -241 504
rect -275 413 -241 425
rect -275 341 -241 357
rect -275 269 -241 289
rect -275 197 -241 221
rect -275 125 -241 153
rect -275 53 -241 85
rect -275 -17 -241 17
rect -275 -85 -241 -53
rect -275 -153 -241 -125
rect -275 -221 -241 -197
rect -275 -289 -241 -269
rect -275 -357 -241 -341
rect -275 -425 -241 -413
rect -275 -504 -241 -485
rect -17 485 17 504
rect -17 413 17 425
rect -17 341 17 357
rect -17 269 17 289
rect -17 197 17 221
rect -17 125 17 153
rect -17 53 17 85
rect -17 -17 17 17
rect -17 -85 17 -53
rect -17 -153 17 -125
rect -17 -221 17 -197
rect -17 -289 17 -269
rect -17 -357 17 -341
rect -17 -425 17 -413
rect -17 -504 17 -485
rect 241 485 275 504
rect 241 413 275 425
rect 241 341 275 357
rect 241 269 275 289
rect 241 197 275 221
rect 241 125 275 153
rect 241 53 275 85
rect 241 -17 275 17
rect 241 -85 275 -53
rect 241 -153 275 -125
rect 241 -221 275 -197
rect 241 -289 275 -269
rect 241 -357 275 -341
rect 241 -425 275 -413
rect 241 -504 275 -485
rect 499 485 533 504
rect 499 413 533 425
rect 499 341 533 357
rect 499 269 533 289
rect 499 197 533 221
rect 499 125 533 153
rect 499 53 533 85
rect 499 -17 533 17
rect 499 -85 533 -53
rect 499 -153 533 -125
rect 499 -221 533 -197
rect 499 -289 533 -269
rect 499 -357 533 -341
rect 499 -425 533 -413
rect 499 -504 533 -485
rect 757 485 791 504
rect 757 413 791 425
rect 757 341 791 357
rect 757 269 791 289
rect 757 197 791 221
rect 757 125 791 153
rect 757 53 791 85
rect 757 -17 791 17
rect 757 -85 791 -53
rect 757 -153 791 -125
rect 757 -221 791 -197
rect 757 -289 791 -269
rect 757 -357 791 -341
rect 757 -425 791 -413
rect 757 -504 791 -485
rect 1015 485 1049 504
rect 1015 413 1049 425
rect 1015 341 1049 357
rect 1015 269 1049 289
rect 1015 197 1049 221
rect 1015 125 1049 153
rect 1015 53 1049 85
rect 1015 -17 1049 17
rect 1015 -85 1049 -53
rect 1015 -153 1049 -125
rect 1015 -221 1049 -197
rect 1015 -289 1049 -269
rect 1015 -357 1049 -341
rect 1015 -425 1049 -413
rect 1015 -504 1049 -485
rect 1273 485 1307 504
rect 1273 413 1307 425
rect 1273 341 1307 357
rect 1273 269 1307 289
rect 1273 197 1307 221
rect 1273 125 1307 153
rect 1273 53 1307 85
rect 1273 -17 1307 17
rect 1273 -85 1307 -53
rect 1273 -153 1307 -125
rect 1273 -221 1307 -197
rect 1273 -289 1307 -269
rect 1273 -357 1307 -341
rect 1273 -425 1307 -413
rect 1273 -504 1307 -485
rect 1531 485 1565 504
rect 1531 413 1565 425
rect 1531 341 1565 357
rect 1531 269 1565 289
rect 1531 197 1565 221
rect 1531 125 1565 153
rect 1531 53 1565 85
rect 1531 -17 1565 17
rect 1531 -85 1565 -53
rect 1531 -153 1565 -125
rect 1531 -221 1565 -197
rect 1531 -289 1565 -269
rect 1531 -357 1565 -341
rect 1531 -425 1565 -413
rect 1531 -504 1565 -485
rect 1789 485 1823 504
rect 1789 413 1823 425
rect 1789 341 1823 357
rect 1789 269 1823 289
rect 1789 197 1823 221
rect 1789 125 1823 153
rect 1789 53 1823 85
rect 1789 -17 1823 17
rect 1789 -85 1823 -53
rect 1789 -153 1823 -125
rect 1789 -221 1823 -197
rect 1789 -289 1823 -269
rect 1789 -357 1823 -341
rect 1789 -425 1823 -413
rect 1789 -504 1823 -485
rect 1903 493 1937 527
rect 1903 425 1937 459
rect 1903 357 1937 391
rect 1903 289 1937 323
rect 1903 221 1937 255
rect 1903 153 1937 187
rect 1903 85 1937 119
rect 1903 17 1937 51
rect 1903 -51 1937 -17
rect 1903 -119 1937 -85
rect 1903 -187 1937 -153
rect 1903 -255 1937 -221
rect 1903 -323 1937 -289
rect 1903 -391 1937 -357
rect 1903 -459 1937 -425
rect 1903 -527 1937 -493
rect -1937 -640 -1903 -561
rect -1777 -572 -1730 -538
rect -1694 -572 -1660 -538
rect -1624 -572 -1577 -538
rect -1519 -572 -1472 -538
rect -1436 -572 -1402 -538
rect -1366 -572 -1319 -538
rect -1261 -572 -1214 -538
rect -1178 -572 -1144 -538
rect -1108 -572 -1061 -538
rect -1003 -572 -956 -538
rect -920 -572 -886 -538
rect -850 -572 -803 -538
rect -745 -572 -698 -538
rect -662 -572 -628 -538
rect -592 -572 -545 -538
rect -487 -572 -440 -538
rect -404 -572 -370 -538
rect -334 -572 -287 -538
rect -229 -572 -182 -538
rect -146 -572 -112 -538
rect -76 -572 -29 -538
rect 29 -572 76 -538
rect 112 -572 146 -538
rect 182 -572 229 -538
rect 287 -572 334 -538
rect 370 -572 404 -538
rect 440 -572 487 -538
rect 545 -572 592 -538
rect 628 -572 662 -538
rect 698 -572 745 -538
rect 803 -572 850 -538
rect 886 -572 920 -538
rect 956 -572 1003 -538
rect 1061 -572 1108 -538
rect 1144 -572 1178 -538
rect 1214 -572 1261 -538
rect 1319 -572 1366 -538
rect 1402 -572 1436 -538
rect 1472 -572 1519 -538
rect 1577 -572 1624 -538
rect 1660 -572 1694 -538
rect 1730 -572 1777 -538
rect 1903 -640 1937 -561
rect -1937 -674 -1819 -640
rect -1785 -674 -1751 -640
rect -1717 -674 -1683 -640
rect -1649 -674 -1615 -640
rect -1581 -674 -1547 -640
rect -1513 -674 -1479 -640
rect -1445 -674 -1411 -640
rect -1377 -674 -1343 -640
rect -1309 -674 -1275 -640
rect -1241 -674 -1207 -640
rect -1173 -674 -1139 -640
rect -1105 -674 -1071 -640
rect -1037 -674 -1003 -640
rect -969 -674 -935 -640
rect -883 -674 -867 -640
rect -811 -674 -799 -640
rect -739 -674 -731 -640
rect -667 -674 -663 -640
rect -561 -674 -557 -640
rect -493 -674 -485 -640
rect -425 -674 -413 -640
rect -357 -674 -341 -640
rect -289 -674 -269 -640
rect -221 -674 -197 -640
rect -153 -674 -125 -640
rect -85 -674 -53 -640
rect -17 -674 17 -640
rect 53 -674 85 -640
rect 125 -674 153 -640
rect 197 -674 221 -640
rect 269 -674 289 -640
rect 341 -674 357 -640
rect 413 -674 425 -640
rect 485 -674 493 -640
rect 557 -674 561 -640
rect 663 -674 667 -640
rect 731 -674 739 -640
rect 799 -674 811 -640
rect 867 -674 883 -640
rect 935 -674 969 -640
rect 1003 -674 1037 -640
rect 1071 -674 1105 -640
rect 1139 -674 1173 -640
rect 1207 -674 1241 -640
rect 1275 -674 1309 -640
rect 1343 -674 1377 -640
rect 1411 -674 1445 -640
rect 1479 -674 1513 -640
rect 1547 -674 1581 -640
rect 1615 -674 1649 -640
rect 1683 -674 1717 -640
rect 1751 -674 1785 -640
rect 1819 -674 1937 -640
<< viali >>
rect -917 640 -901 674
rect -901 640 -883 674
rect -845 640 -833 674
rect -833 640 -811 674
rect -773 640 -765 674
rect -765 640 -739 674
rect -701 640 -697 674
rect -697 640 -667 674
rect -629 640 -595 674
rect -557 640 -527 674
rect -527 640 -523 674
rect -485 640 -459 674
rect -459 640 -451 674
rect -413 640 -391 674
rect -391 640 -379 674
rect -341 640 -323 674
rect -323 640 -307 674
rect -269 640 -255 674
rect -255 640 -235 674
rect -197 640 -187 674
rect -187 640 -163 674
rect -125 640 -119 674
rect -119 640 -91 674
rect -53 640 -51 674
rect -51 640 -19 674
rect 19 640 51 674
rect 51 640 53 674
rect 91 640 119 674
rect 119 640 125 674
rect 163 640 187 674
rect 187 640 197 674
rect 235 640 255 674
rect 255 640 269 674
rect 307 640 323 674
rect 323 640 341 674
rect 379 640 391 674
rect 391 640 413 674
rect 451 640 459 674
rect 459 640 485 674
rect 523 640 527 674
rect 527 640 557 674
rect 595 640 629 674
rect 667 640 697 674
rect 697 640 701 674
rect 739 640 765 674
rect 765 640 773 674
rect 811 640 833 674
rect 833 640 845 674
rect 883 640 901 674
rect 901 640 917 674
rect -1730 538 -1728 572
rect -1728 538 -1696 572
rect -1658 538 -1626 572
rect -1626 538 -1624 572
rect -1472 538 -1470 572
rect -1470 538 -1438 572
rect -1400 538 -1368 572
rect -1368 538 -1366 572
rect -1214 538 -1212 572
rect -1212 538 -1180 572
rect -1142 538 -1110 572
rect -1110 538 -1108 572
rect -956 538 -954 572
rect -954 538 -922 572
rect -884 538 -852 572
rect -852 538 -850 572
rect -698 538 -696 572
rect -696 538 -664 572
rect -626 538 -594 572
rect -594 538 -592 572
rect -440 538 -438 572
rect -438 538 -406 572
rect -368 538 -336 572
rect -336 538 -334 572
rect -182 538 -180 572
rect -180 538 -148 572
rect -110 538 -78 572
rect -78 538 -76 572
rect 76 538 78 572
rect 78 538 110 572
rect 148 538 180 572
rect 180 538 182 572
rect 334 538 336 572
rect 336 538 368 572
rect 406 538 438 572
rect 438 538 440 572
rect 592 538 594 572
rect 594 538 626 572
rect 664 538 696 572
rect 696 538 698 572
rect 850 538 852 572
rect 852 538 884 572
rect 922 538 954 572
rect 954 538 956 572
rect 1108 538 1110 572
rect 1110 538 1142 572
rect 1180 538 1212 572
rect 1212 538 1214 572
rect 1366 538 1368 572
rect 1368 538 1400 572
rect 1438 538 1470 572
rect 1470 538 1472 572
rect 1624 538 1626 572
rect 1626 538 1658 572
rect 1696 538 1728 572
rect 1728 538 1730 572
rect -1823 459 -1789 485
rect -1823 451 -1789 459
rect -1823 391 -1789 413
rect -1823 379 -1789 391
rect -1823 323 -1789 341
rect -1823 307 -1789 323
rect -1823 255 -1789 269
rect -1823 235 -1789 255
rect -1823 187 -1789 197
rect -1823 163 -1789 187
rect -1823 119 -1789 125
rect -1823 91 -1789 119
rect -1823 51 -1789 53
rect -1823 19 -1789 51
rect -1823 -51 -1789 -19
rect -1823 -53 -1789 -51
rect -1823 -119 -1789 -91
rect -1823 -125 -1789 -119
rect -1823 -187 -1789 -163
rect -1823 -197 -1789 -187
rect -1823 -255 -1789 -235
rect -1823 -269 -1789 -255
rect -1823 -323 -1789 -307
rect -1823 -341 -1789 -323
rect -1823 -391 -1789 -379
rect -1823 -413 -1789 -391
rect -1823 -459 -1789 -451
rect -1823 -485 -1789 -459
rect -1565 459 -1531 485
rect -1565 451 -1531 459
rect -1565 391 -1531 413
rect -1565 379 -1531 391
rect -1565 323 -1531 341
rect -1565 307 -1531 323
rect -1565 255 -1531 269
rect -1565 235 -1531 255
rect -1565 187 -1531 197
rect -1565 163 -1531 187
rect -1565 119 -1531 125
rect -1565 91 -1531 119
rect -1565 51 -1531 53
rect -1565 19 -1531 51
rect -1565 -51 -1531 -19
rect -1565 -53 -1531 -51
rect -1565 -119 -1531 -91
rect -1565 -125 -1531 -119
rect -1565 -187 -1531 -163
rect -1565 -197 -1531 -187
rect -1565 -255 -1531 -235
rect -1565 -269 -1531 -255
rect -1565 -323 -1531 -307
rect -1565 -341 -1531 -323
rect -1565 -391 -1531 -379
rect -1565 -413 -1531 -391
rect -1565 -459 -1531 -451
rect -1565 -485 -1531 -459
rect -1307 459 -1273 485
rect -1307 451 -1273 459
rect -1307 391 -1273 413
rect -1307 379 -1273 391
rect -1307 323 -1273 341
rect -1307 307 -1273 323
rect -1307 255 -1273 269
rect -1307 235 -1273 255
rect -1307 187 -1273 197
rect -1307 163 -1273 187
rect -1307 119 -1273 125
rect -1307 91 -1273 119
rect -1307 51 -1273 53
rect -1307 19 -1273 51
rect -1307 -51 -1273 -19
rect -1307 -53 -1273 -51
rect -1307 -119 -1273 -91
rect -1307 -125 -1273 -119
rect -1307 -187 -1273 -163
rect -1307 -197 -1273 -187
rect -1307 -255 -1273 -235
rect -1307 -269 -1273 -255
rect -1307 -323 -1273 -307
rect -1307 -341 -1273 -323
rect -1307 -391 -1273 -379
rect -1307 -413 -1273 -391
rect -1307 -459 -1273 -451
rect -1307 -485 -1273 -459
rect -1049 459 -1015 485
rect -1049 451 -1015 459
rect -1049 391 -1015 413
rect -1049 379 -1015 391
rect -1049 323 -1015 341
rect -1049 307 -1015 323
rect -1049 255 -1015 269
rect -1049 235 -1015 255
rect -1049 187 -1015 197
rect -1049 163 -1015 187
rect -1049 119 -1015 125
rect -1049 91 -1015 119
rect -1049 51 -1015 53
rect -1049 19 -1015 51
rect -1049 -51 -1015 -19
rect -1049 -53 -1015 -51
rect -1049 -119 -1015 -91
rect -1049 -125 -1015 -119
rect -1049 -187 -1015 -163
rect -1049 -197 -1015 -187
rect -1049 -255 -1015 -235
rect -1049 -269 -1015 -255
rect -1049 -323 -1015 -307
rect -1049 -341 -1015 -323
rect -1049 -391 -1015 -379
rect -1049 -413 -1015 -391
rect -1049 -459 -1015 -451
rect -1049 -485 -1015 -459
rect -791 459 -757 485
rect -791 451 -757 459
rect -791 391 -757 413
rect -791 379 -757 391
rect -791 323 -757 341
rect -791 307 -757 323
rect -791 255 -757 269
rect -791 235 -757 255
rect -791 187 -757 197
rect -791 163 -757 187
rect -791 119 -757 125
rect -791 91 -757 119
rect -791 51 -757 53
rect -791 19 -757 51
rect -791 -51 -757 -19
rect -791 -53 -757 -51
rect -791 -119 -757 -91
rect -791 -125 -757 -119
rect -791 -187 -757 -163
rect -791 -197 -757 -187
rect -791 -255 -757 -235
rect -791 -269 -757 -255
rect -791 -323 -757 -307
rect -791 -341 -757 -323
rect -791 -391 -757 -379
rect -791 -413 -757 -391
rect -791 -459 -757 -451
rect -791 -485 -757 -459
rect -533 459 -499 485
rect -533 451 -499 459
rect -533 391 -499 413
rect -533 379 -499 391
rect -533 323 -499 341
rect -533 307 -499 323
rect -533 255 -499 269
rect -533 235 -499 255
rect -533 187 -499 197
rect -533 163 -499 187
rect -533 119 -499 125
rect -533 91 -499 119
rect -533 51 -499 53
rect -533 19 -499 51
rect -533 -51 -499 -19
rect -533 -53 -499 -51
rect -533 -119 -499 -91
rect -533 -125 -499 -119
rect -533 -187 -499 -163
rect -533 -197 -499 -187
rect -533 -255 -499 -235
rect -533 -269 -499 -255
rect -533 -323 -499 -307
rect -533 -341 -499 -323
rect -533 -391 -499 -379
rect -533 -413 -499 -391
rect -533 -459 -499 -451
rect -533 -485 -499 -459
rect -275 459 -241 485
rect -275 451 -241 459
rect -275 391 -241 413
rect -275 379 -241 391
rect -275 323 -241 341
rect -275 307 -241 323
rect -275 255 -241 269
rect -275 235 -241 255
rect -275 187 -241 197
rect -275 163 -241 187
rect -275 119 -241 125
rect -275 91 -241 119
rect -275 51 -241 53
rect -275 19 -241 51
rect -275 -51 -241 -19
rect -275 -53 -241 -51
rect -275 -119 -241 -91
rect -275 -125 -241 -119
rect -275 -187 -241 -163
rect -275 -197 -241 -187
rect -275 -255 -241 -235
rect -275 -269 -241 -255
rect -275 -323 -241 -307
rect -275 -341 -241 -323
rect -275 -391 -241 -379
rect -275 -413 -241 -391
rect -275 -459 -241 -451
rect -275 -485 -241 -459
rect -17 459 17 485
rect -17 451 17 459
rect -17 391 17 413
rect -17 379 17 391
rect -17 323 17 341
rect -17 307 17 323
rect -17 255 17 269
rect -17 235 17 255
rect -17 187 17 197
rect -17 163 17 187
rect -17 119 17 125
rect -17 91 17 119
rect -17 51 17 53
rect -17 19 17 51
rect -17 -51 17 -19
rect -17 -53 17 -51
rect -17 -119 17 -91
rect -17 -125 17 -119
rect -17 -187 17 -163
rect -17 -197 17 -187
rect -17 -255 17 -235
rect -17 -269 17 -255
rect -17 -323 17 -307
rect -17 -341 17 -323
rect -17 -391 17 -379
rect -17 -413 17 -391
rect -17 -459 17 -451
rect -17 -485 17 -459
rect 241 459 275 485
rect 241 451 275 459
rect 241 391 275 413
rect 241 379 275 391
rect 241 323 275 341
rect 241 307 275 323
rect 241 255 275 269
rect 241 235 275 255
rect 241 187 275 197
rect 241 163 275 187
rect 241 119 275 125
rect 241 91 275 119
rect 241 51 275 53
rect 241 19 275 51
rect 241 -51 275 -19
rect 241 -53 275 -51
rect 241 -119 275 -91
rect 241 -125 275 -119
rect 241 -187 275 -163
rect 241 -197 275 -187
rect 241 -255 275 -235
rect 241 -269 275 -255
rect 241 -323 275 -307
rect 241 -341 275 -323
rect 241 -391 275 -379
rect 241 -413 275 -391
rect 241 -459 275 -451
rect 241 -485 275 -459
rect 499 459 533 485
rect 499 451 533 459
rect 499 391 533 413
rect 499 379 533 391
rect 499 323 533 341
rect 499 307 533 323
rect 499 255 533 269
rect 499 235 533 255
rect 499 187 533 197
rect 499 163 533 187
rect 499 119 533 125
rect 499 91 533 119
rect 499 51 533 53
rect 499 19 533 51
rect 499 -51 533 -19
rect 499 -53 533 -51
rect 499 -119 533 -91
rect 499 -125 533 -119
rect 499 -187 533 -163
rect 499 -197 533 -187
rect 499 -255 533 -235
rect 499 -269 533 -255
rect 499 -323 533 -307
rect 499 -341 533 -323
rect 499 -391 533 -379
rect 499 -413 533 -391
rect 499 -459 533 -451
rect 499 -485 533 -459
rect 757 459 791 485
rect 757 451 791 459
rect 757 391 791 413
rect 757 379 791 391
rect 757 323 791 341
rect 757 307 791 323
rect 757 255 791 269
rect 757 235 791 255
rect 757 187 791 197
rect 757 163 791 187
rect 757 119 791 125
rect 757 91 791 119
rect 757 51 791 53
rect 757 19 791 51
rect 757 -51 791 -19
rect 757 -53 791 -51
rect 757 -119 791 -91
rect 757 -125 791 -119
rect 757 -187 791 -163
rect 757 -197 791 -187
rect 757 -255 791 -235
rect 757 -269 791 -255
rect 757 -323 791 -307
rect 757 -341 791 -323
rect 757 -391 791 -379
rect 757 -413 791 -391
rect 757 -459 791 -451
rect 757 -485 791 -459
rect 1015 459 1049 485
rect 1015 451 1049 459
rect 1015 391 1049 413
rect 1015 379 1049 391
rect 1015 323 1049 341
rect 1015 307 1049 323
rect 1015 255 1049 269
rect 1015 235 1049 255
rect 1015 187 1049 197
rect 1015 163 1049 187
rect 1015 119 1049 125
rect 1015 91 1049 119
rect 1015 51 1049 53
rect 1015 19 1049 51
rect 1015 -51 1049 -19
rect 1015 -53 1049 -51
rect 1015 -119 1049 -91
rect 1015 -125 1049 -119
rect 1015 -187 1049 -163
rect 1015 -197 1049 -187
rect 1015 -255 1049 -235
rect 1015 -269 1049 -255
rect 1015 -323 1049 -307
rect 1015 -341 1049 -323
rect 1015 -391 1049 -379
rect 1015 -413 1049 -391
rect 1015 -459 1049 -451
rect 1015 -485 1049 -459
rect 1273 459 1307 485
rect 1273 451 1307 459
rect 1273 391 1307 413
rect 1273 379 1307 391
rect 1273 323 1307 341
rect 1273 307 1307 323
rect 1273 255 1307 269
rect 1273 235 1307 255
rect 1273 187 1307 197
rect 1273 163 1307 187
rect 1273 119 1307 125
rect 1273 91 1307 119
rect 1273 51 1307 53
rect 1273 19 1307 51
rect 1273 -51 1307 -19
rect 1273 -53 1307 -51
rect 1273 -119 1307 -91
rect 1273 -125 1307 -119
rect 1273 -187 1307 -163
rect 1273 -197 1307 -187
rect 1273 -255 1307 -235
rect 1273 -269 1307 -255
rect 1273 -323 1307 -307
rect 1273 -341 1307 -323
rect 1273 -391 1307 -379
rect 1273 -413 1307 -391
rect 1273 -459 1307 -451
rect 1273 -485 1307 -459
rect 1531 459 1565 485
rect 1531 451 1565 459
rect 1531 391 1565 413
rect 1531 379 1565 391
rect 1531 323 1565 341
rect 1531 307 1565 323
rect 1531 255 1565 269
rect 1531 235 1565 255
rect 1531 187 1565 197
rect 1531 163 1565 187
rect 1531 119 1565 125
rect 1531 91 1565 119
rect 1531 51 1565 53
rect 1531 19 1565 51
rect 1531 -51 1565 -19
rect 1531 -53 1565 -51
rect 1531 -119 1565 -91
rect 1531 -125 1565 -119
rect 1531 -187 1565 -163
rect 1531 -197 1565 -187
rect 1531 -255 1565 -235
rect 1531 -269 1565 -255
rect 1531 -323 1565 -307
rect 1531 -341 1565 -323
rect 1531 -391 1565 -379
rect 1531 -413 1565 -391
rect 1531 -459 1565 -451
rect 1531 -485 1565 -459
rect 1789 459 1823 485
rect 1789 451 1823 459
rect 1789 391 1823 413
rect 1789 379 1823 391
rect 1789 323 1823 341
rect 1789 307 1823 323
rect 1789 255 1823 269
rect 1789 235 1823 255
rect 1789 187 1823 197
rect 1789 163 1823 187
rect 1789 119 1823 125
rect 1789 91 1823 119
rect 1789 51 1823 53
rect 1789 19 1823 51
rect 1789 -51 1823 -19
rect 1789 -53 1823 -51
rect 1789 -119 1823 -91
rect 1789 -125 1823 -119
rect 1789 -187 1823 -163
rect 1789 -197 1823 -187
rect 1789 -255 1823 -235
rect 1789 -269 1823 -255
rect 1789 -323 1823 -307
rect 1789 -341 1823 -323
rect 1789 -391 1823 -379
rect 1789 -413 1823 -391
rect 1789 -459 1823 -451
rect 1789 -485 1823 -459
rect -1730 -572 -1728 -538
rect -1728 -572 -1696 -538
rect -1658 -572 -1626 -538
rect -1626 -572 -1624 -538
rect -1472 -572 -1470 -538
rect -1470 -572 -1438 -538
rect -1400 -572 -1368 -538
rect -1368 -572 -1366 -538
rect -1214 -572 -1212 -538
rect -1212 -572 -1180 -538
rect -1142 -572 -1110 -538
rect -1110 -572 -1108 -538
rect -956 -572 -954 -538
rect -954 -572 -922 -538
rect -884 -572 -852 -538
rect -852 -572 -850 -538
rect -698 -572 -696 -538
rect -696 -572 -664 -538
rect -626 -572 -594 -538
rect -594 -572 -592 -538
rect -440 -572 -438 -538
rect -438 -572 -406 -538
rect -368 -572 -336 -538
rect -336 -572 -334 -538
rect -182 -572 -180 -538
rect -180 -572 -148 -538
rect -110 -572 -78 -538
rect -78 -572 -76 -538
rect 76 -572 78 -538
rect 78 -572 110 -538
rect 148 -572 180 -538
rect 180 -572 182 -538
rect 334 -572 336 -538
rect 336 -572 368 -538
rect 406 -572 438 -538
rect 438 -572 440 -538
rect 592 -572 594 -538
rect 594 -572 626 -538
rect 664 -572 696 -538
rect 696 -572 698 -538
rect 850 -572 852 -538
rect 852 -572 884 -538
rect 922 -572 954 -538
rect 954 -572 956 -538
rect 1108 -572 1110 -538
rect 1110 -572 1142 -538
rect 1180 -572 1212 -538
rect 1212 -572 1214 -538
rect 1366 -572 1368 -538
rect 1368 -572 1400 -538
rect 1438 -572 1470 -538
rect 1470 -572 1472 -538
rect 1624 -572 1626 -538
rect 1626 -572 1658 -538
rect 1696 -572 1728 -538
rect 1728 -572 1730 -538
rect -917 -674 -901 -640
rect -901 -674 -883 -640
rect -845 -674 -833 -640
rect -833 -674 -811 -640
rect -773 -674 -765 -640
rect -765 -674 -739 -640
rect -701 -674 -697 -640
rect -697 -674 -667 -640
rect -629 -674 -595 -640
rect -557 -674 -527 -640
rect -527 -674 -523 -640
rect -485 -674 -459 -640
rect -459 -674 -451 -640
rect -413 -674 -391 -640
rect -391 -674 -379 -640
rect -341 -674 -323 -640
rect -323 -674 -307 -640
rect -269 -674 -255 -640
rect -255 -674 -235 -640
rect -197 -674 -187 -640
rect -187 -674 -163 -640
rect -125 -674 -119 -640
rect -119 -674 -91 -640
rect -53 -674 -51 -640
rect -51 -674 -19 -640
rect 19 -674 51 -640
rect 51 -674 53 -640
rect 91 -674 119 -640
rect 119 -674 125 -640
rect 163 -674 187 -640
rect 187 -674 197 -640
rect 235 -674 255 -640
rect 255 -674 269 -640
rect 307 -674 323 -640
rect 323 -674 341 -640
rect 379 -674 391 -640
rect 391 -674 413 -640
rect 451 -674 459 -640
rect 459 -674 485 -640
rect 523 -674 527 -640
rect 527 -674 557 -640
rect 595 -674 629 -640
rect 667 -674 697 -640
rect 697 -674 701 -640
rect 739 -674 765 -640
rect 765 -674 773 -640
rect 811 -674 833 -640
rect 833 -674 845 -640
rect 883 -674 901 -640
rect 901 -674 917 -640
<< metal1 >>
rect -963 674 963 680
rect -963 640 -917 674
rect -883 640 -845 674
rect -811 640 -773 674
rect -739 640 -701 674
rect -667 640 -629 674
rect -595 640 -557 674
rect -523 640 -485 674
rect -451 640 -413 674
rect -379 640 -341 674
rect -307 640 -269 674
rect -235 640 -197 674
rect -163 640 -125 674
rect -91 640 -53 674
rect -19 640 19 674
rect 53 640 91 674
rect 125 640 163 674
rect 197 640 235 674
rect 269 640 307 674
rect 341 640 379 674
rect 413 640 451 674
rect 485 640 523 674
rect 557 640 595 674
rect 629 640 667 674
rect 701 640 739 674
rect 773 640 811 674
rect 845 640 883 674
rect 917 640 963 674
rect -963 634 963 640
rect -1773 572 -1581 578
rect -1773 538 -1730 572
rect -1696 538 -1658 572
rect -1624 538 -1581 572
rect -1773 532 -1581 538
rect -1515 572 -1323 578
rect -1515 538 -1472 572
rect -1438 538 -1400 572
rect -1366 538 -1323 572
rect -1515 532 -1323 538
rect -1257 572 -1065 578
rect -1257 538 -1214 572
rect -1180 538 -1142 572
rect -1108 538 -1065 572
rect -1257 532 -1065 538
rect -999 572 -807 578
rect -999 538 -956 572
rect -922 538 -884 572
rect -850 538 -807 572
rect -999 532 -807 538
rect -741 572 -549 578
rect -741 538 -698 572
rect -664 538 -626 572
rect -592 538 -549 572
rect -741 532 -549 538
rect -483 572 -291 578
rect -483 538 -440 572
rect -406 538 -368 572
rect -334 538 -291 572
rect -483 532 -291 538
rect -225 572 -33 578
rect -225 538 -182 572
rect -148 538 -110 572
rect -76 538 -33 572
rect -225 532 -33 538
rect 33 572 225 578
rect 33 538 76 572
rect 110 538 148 572
rect 182 538 225 572
rect 33 532 225 538
rect 291 572 483 578
rect 291 538 334 572
rect 368 538 406 572
rect 440 538 483 572
rect 291 532 483 538
rect 549 572 741 578
rect 549 538 592 572
rect 626 538 664 572
rect 698 538 741 572
rect 549 532 741 538
rect 807 572 999 578
rect 807 538 850 572
rect 884 538 922 572
rect 956 538 999 572
rect 807 532 999 538
rect 1065 572 1257 578
rect 1065 538 1108 572
rect 1142 538 1180 572
rect 1214 538 1257 572
rect 1065 532 1257 538
rect 1323 572 1515 578
rect 1323 538 1366 572
rect 1400 538 1438 572
rect 1472 538 1515 572
rect 1323 532 1515 538
rect 1581 572 1773 578
rect 1581 538 1624 572
rect 1658 538 1696 572
rect 1730 538 1773 572
rect 1581 532 1773 538
rect -1829 485 -1783 500
rect -1829 451 -1823 485
rect -1789 451 -1783 485
rect -1829 413 -1783 451
rect -1829 379 -1823 413
rect -1789 379 -1783 413
rect -1829 341 -1783 379
rect -1829 307 -1823 341
rect -1789 307 -1783 341
rect -1829 269 -1783 307
rect -1829 235 -1823 269
rect -1789 235 -1783 269
rect -1829 197 -1783 235
rect -1829 163 -1823 197
rect -1789 163 -1783 197
rect -1829 125 -1783 163
rect -1829 91 -1823 125
rect -1789 91 -1783 125
rect -1829 53 -1783 91
rect -1829 19 -1823 53
rect -1789 19 -1783 53
rect -1829 -19 -1783 19
rect -1829 -53 -1823 -19
rect -1789 -53 -1783 -19
rect -1829 -91 -1783 -53
rect -1829 -125 -1823 -91
rect -1789 -125 -1783 -91
rect -1829 -163 -1783 -125
rect -1829 -197 -1823 -163
rect -1789 -197 -1783 -163
rect -1829 -235 -1783 -197
rect -1829 -269 -1823 -235
rect -1789 -269 -1783 -235
rect -1829 -307 -1783 -269
rect -1829 -341 -1823 -307
rect -1789 -341 -1783 -307
rect -1829 -379 -1783 -341
rect -1829 -413 -1823 -379
rect -1789 -413 -1783 -379
rect -1829 -451 -1783 -413
rect -1829 -485 -1823 -451
rect -1789 -485 -1783 -451
rect -1829 -500 -1783 -485
rect -1571 485 -1525 500
rect -1571 451 -1565 485
rect -1531 451 -1525 485
rect -1571 413 -1525 451
rect -1571 379 -1565 413
rect -1531 379 -1525 413
rect -1571 341 -1525 379
rect -1571 307 -1565 341
rect -1531 307 -1525 341
rect -1571 269 -1525 307
rect -1571 235 -1565 269
rect -1531 235 -1525 269
rect -1571 197 -1525 235
rect -1571 163 -1565 197
rect -1531 163 -1525 197
rect -1571 125 -1525 163
rect -1571 91 -1565 125
rect -1531 91 -1525 125
rect -1571 53 -1525 91
rect -1571 19 -1565 53
rect -1531 19 -1525 53
rect -1571 -19 -1525 19
rect -1571 -53 -1565 -19
rect -1531 -53 -1525 -19
rect -1571 -91 -1525 -53
rect -1571 -125 -1565 -91
rect -1531 -125 -1525 -91
rect -1571 -163 -1525 -125
rect -1571 -197 -1565 -163
rect -1531 -197 -1525 -163
rect -1571 -235 -1525 -197
rect -1571 -269 -1565 -235
rect -1531 -269 -1525 -235
rect -1571 -307 -1525 -269
rect -1571 -341 -1565 -307
rect -1531 -341 -1525 -307
rect -1571 -379 -1525 -341
rect -1571 -413 -1565 -379
rect -1531 -413 -1525 -379
rect -1571 -451 -1525 -413
rect -1571 -485 -1565 -451
rect -1531 -485 -1525 -451
rect -1571 -500 -1525 -485
rect -1313 485 -1267 500
rect -1313 451 -1307 485
rect -1273 451 -1267 485
rect -1313 413 -1267 451
rect -1313 379 -1307 413
rect -1273 379 -1267 413
rect -1313 341 -1267 379
rect -1313 307 -1307 341
rect -1273 307 -1267 341
rect -1313 269 -1267 307
rect -1313 235 -1307 269
rect -1273 235 -1267 269
rect -1313 197 -1267 235
rect -1313 163 -1307 197
rect -1273 163 -1267 197
rect -1313 125 -1267 163
rect -1313 91 -1307 125
rect -1273 91 -1267 125
rect -1313 53 -1267 91
rect -1313 19 -1307 53
rect -1273 19 -1267 53
rect -1313 -19 -1267 19
rect -1313 -53 -1307 -19
rect -1273 -53 -1267 -19
rect -1313 -91 -1267 -53
rect -1313 -125 -1307 -91
rect -1273 -125 -1267 -91
rect -1313 -163 -1267 -125
rect -1313 -197 -1307 -163
rect -1273 -197 -1267 -163
rect -1313 -235 -1267 -197
rect -1313 -269 -1307 -235
rect -1273 -269 -1267 -235
rect -1313 -307 -1267 -269
rect -1313 -341 -1307 -307
rect -1273 -341 -1267 -307
rect -1313 -379 -1267 -341
rect -1313 -413 -1307 -379
rect -1273 -413 -1267 -379
rect -1313 -451 -1267 -413
rect -1313 -485 -1307 -451
rect -1273 -485 -1267 -451
rect -1313 -500 -1267 -485
rect -1055 485 -1009 500
rect -1055 451 -1049 485
rect -1015 451 -1009 485
rect -1055 413 -1009 451
rect -1055 379 -1049 413
rect -1015 379 -1009 413
rect -1055 341 -1009 379
rect -1055 307 -1049 341
rect -1015 307 -1009 341
rect -1055 269 -1009 307
rect -1055 235 -1049 269
rect -1015 235 -1009 269
rect -1055 197 -1009 235
rect -1055 163 -1049 197
rect -1015 163 -1009 197
rect -1055 125 -1009 163
rect -1055 91 -1049 125
rect -1015 91 -1009 125
rect -1055 53 -1009 91
rect -1055 19 -1049 53
rect -1015 19 -1009 53
rect -1055 -19 -1009 19
rect -1055 -53 -1049 -19
rect -1015 -53 -1009 -19
rect -1055 -91 -1009 -53
rect -1055 -125 -1049 -91
rect -1015 -125 -1009 -91
rect -1055 -163 -1009 -125
rect -1055 -197 -1049 -163
rect -1015 -197 -1009 -163
rect -1055 -235 -1009 -197
rect -1055 -269 -1049 -235
rect -1015 -269 -1009 -235
rect -1055 -307 -1009 -269
rect -1055 -341 -1049 -307
rect -1015 -341 -1009 -307
rect -1055 -379 -1009 -341
rect -1055 -413 -1049 -379
rect -1015 -413 -1009 -379
rect -1055 -451 -1009 -413
rect -1055 -485 -1049 -451
rect -1015 -485 -1009 -451
rect -1055 -500 -1009 -485
rect -797 485 -751 500
rect -797 451 -791 485
rect -757 451 -751 485
rect -797 413 -751 451
rect -797 379 -791 413
rect -757 379 -751 413
rect -797 341 -751 379
rect -797 307 -791 341
rect -757 307 -751 341
rect -797 269 -751 307
rect -797 235 -791 269
rect -757 235 -751 269
rect -797 197 -751 235
rect -797 163 -791 197
rect -757 163 -751 197
rect -797 125 -751 163
rect -797 91 -791 125
rect -757 91 -751 125
rect -797 53 -751 91
rect -797 19 -791 53
rect -757 19 -751 53
rect -797 -19 -751 19
rect -797 -53 -791 -19
rect -757 -53 -751 -19
rect -797 -91 -751 -53
rect -797 -125 -791 -91
rect -757 -125 -751 -91
rect -797 -163 -751 -125
rect -797 -197 -791 -163
rect -757 -197 -751 -163
rect -797 -235 -751 -197
rect -797 -269 -791 -235
rect -757 -269 -751 -235
rect -797 -307 -751 -269
rect -797 -341 -791 -307
rect -757 -341 -751 -307
rect -797 -379 -751 -341
rect -797 -413 -791 -379
rect -757 -413 -751 -379
rect -797 -451 -751 -413
rect -797 -485 -791 -451
rect -757 -485 -751 -451
rect -797 -500 -751 -485
rect -539 485 -493 500
rect -539 451 -533 485
rect -499 451 -493 485
rect -539 413 -493 451
rect -539 379 -533 413
rect -499 379 -493 413
rect -539 341 -493 379
rect -539 307 -533 341
rect -499 307 -493 341
rect -539 269 -493 307
rect -539 235 -533 269
rect -499 235 -493 269
rect -539 197 -493 235
rect -539 163 -533 197
rect -499 163 -493 197
rect -539 125 -493 163
rect -539 91 -533 125
rect -499 91 -493 125
rect -539 53 -493 91
rect -539 19 -533 53
rect -499 19 -493 53
rect -539 -19 -493 19
rect -539 -53 -533 -19
rect -499 -53 -493 -19
rect -539 -91 -493 -53
rect -539 -125 -533 -91
rect -499 -125 -493 -91
rect -539 -163 -493 -125
rect -539 -197 -533 -163
rect -499 -197 -493 -163
rect -539 -235 -493 -197
rect -539 -269 -533 -235
rect -499 -269 -493 -235
rect -539 -307 -493 -269
rect -539 -341 -533 -307
rect -499 -341 -493 -307
rect -539 -379 -493 -341
rect -539 -413 -533 -379
rect -499 -413 -493 -379
rect -539 -451 -493 -413
rect -539 -485 -533 -451
rect -499 -485 -493 -451
rect -539 -500 -493 -485
rect -281 485 -235 500
rect -281 451 -275 485
rect -241 451 -235 485
rect -281 413 -235 451
rect -281 379 -275 413
rect -241 379 -235 413
rect -281 341 -235 379
rect -281 307 -275 341
rect -241 307 -235 341
rect -281 269 -235 307
rect -281 235 -275 269
rect -241 235 -235 269
rect -281 197 -235 235
rect -281 163 -275 197
rect -241 163 -235 197
rect -281 125 -235 163
rect -281 91 -275 125
rect -241 91 -235 125
rect -281 53 -235 91
rect -281 19 -275 53
rect -241 19 -235 53
rect -281 -19 -235 19
rect -281 -53 -275 -19
rect -241 -53 -235 -19
rect -281 -91 -235 -53
rect -281 -125 -275 -91
rect -241 -125 -235 -91
rect -281 -163 -235 -125
rect -281 -197 -275 -163
rect -241 -197 -235 -163
rect -281 -235 -235 -197
rect -281 -269 -275 -235
rect -241 -269 -235 -235
rect -281 -307 -235 -269
rect -281 -341 -275 -307
rect -241 -341 -235 -307
rect -281 -379 -235 -341
rect -281 -413 -275 -379
rect -241 -413 -235 -379
rect -281 -451 -235 -413
rect -281 -485 -275 -451
rect -241 -485 -235 -451
rect -281 -500 -235 -485
rect -23 485 23 500
rect -23 451 -17 485
rect 17 451 23 485
rect -23 413 23 451
rect -23 379 -17 413
rect 17 379 23 413
rect -23 341 23 379
rect -23 307 -17 341
rect 17 307 23 341
rect -23 269 23 307
rect -23 235 -17 269
rect 17 235 23 269
rect -23 197 23 235
rect -23 163 -17 197
rect 17 163 23 197
rect -23 125 23 163
rect -23 91 -17 125
rect 17 91 23 125
rect -23 53 23 91
rect -23 19 -17 53
rect 17 19 23 53
rect -23 -19 23 19
rect -23 -53 -17 -19
rect 17 -53 23 -19
rect -23 -91 23 -53
rect -23 -125 -17 -91
rect 17 -125 23 -91
rect -23 -163 23 -125
rect -23 -197 -17 -163
rect 17 -197 23 -163
rect -23 -235 23 -197
rect -23 -269 -17 -235
rect 17 -269 23 -235
rect -23 -307 23 -269
rect -23 -341 -17 -307
rect 17 -341 23 -307
rect -23 -379 23 -341
rect -23 -413 -17 -379
rect 17 -413 23 -379
rect -23 -451 23 -413
rect -23 -485 -17 -451
rect 17 -485 23 -451
rect -23 -500 23 -485
rect 235 485 281 500
rect 235 451 241 485
rect 275 451 281 485
rect 235 413 281 451
rect 235 379 241 413
rect 275 379 281 413
rect 235 341 281 379
rect 235 307 241 341
rect 275 307 281 341
rect 235 269 281 307
rect 235 235 241 269
rect 275 235 281 269
rect 235 197 281 235
rect 235 163 241 197
rect 275 163 281 197
rect 235 125 281 163
rect 235 91 241 125
rect 275 91 281 125
rect 235 53 281 91
rect 235 19 241 53
rect 275 19 281 53
rect 235 -19 281 19
rect 235 -53 241 -19
rect 275 -53 281 -19
rect 235 -91 281 -53
rect 235 -125 241 -91
rect 275 -125 281 -91
rect 235 -163 281 -125
rect 235 -197 241 -163
rect 275 -197 281 -163
rect 235 -235 281 -197
rect 235 -269 241 -235
rect 275 -269 281 -235
rect 235 -307 281 -269
rect 235 -341 241 -307
rect 275 -341 281 -307
rect 235 -379 281 -341
rect 235 -413 241 -379
rect 275 -413 281 -379
rect 235 -451 281 -413
rect 235 -485 241 -451
rect 275 -485 281 -451
rect 235 -500 281 -485
rect 493 485 539 500
rect 493 451 499 485
rect 533 451 539 485
rect 493 413 539 451
rect 493 379 499 413
rect 533 379 539 413
rect 493 341 539 379
rect 493 307 499 341
rect 533 307 539 341
rect 493 269 539 307
rect 493 235 499 269
rect 533 235 539 269
rect 493 197 539 235
rect 493 163 499 197
rect 533 163 539 197
rect 493 125 539 163
rect 493 91 499 125
rect 533 91 539 125
rect 493 53 539 91
rect 493 19 499 53
rect 533 19 539 53
rect 493 -19 539 19
rect 493 -53 499 -19
rect 533 -53 539 -19
rect 493 -91 539 -53
rect 493 -125 499 -91
rect 533 -125 539 -91
rect 493 -163 539 -125
rect 493 -197 499 -163
rect 533 -197 539 -163
rect 493 -235 539 -197
rect 493 -269 499 -235
rect 533 -269 539 -235
rect 493 -307 539 -269
rect 493 -341 499 -307
rect 533 -341 539 -307
rect 493 -379 539 -341
rect 493 -413 499 -379
rect 533 -413 539 -379
rect 493 -451 539 -413
rect 493 -485 499 -451
rect 533 -485 539 -451
rect 493 -500 539 -485
rect 751 485 797 500
rect 751 451 757 485
rect 791 451 797 485
rect 751 413 797 451
rect 751 379 757 413
rect 791 379 797 413
rect 751 341 797 379
rect 751 307 757 341
rect 791 307 797 341
rect 751 269 797 307
rect 751 235 757 269
rect 791 235 797 269
rect 751 197 797 235
rect 751 163 757 197
rect 791 163 797 197
rect 751 125 797 163
rect 751 91 757 125
rect 791 91 797 125
rect 751 53 797 91
rect 751 19 757 53
rect 791 19 797 53
rect 751 -19 797 19
rect 751 -53 757 -19
rect 791 -53 797 -19
rect 751 -91 797 -53
rect 751 -125 757 -91
rect 791 -125 797 -91
rect 751 -163 797 -125
rect 751 -197 757 -163
rect 791 -197 797 -163
rect 751 -235 797 -197
rect 751 -269 757 -235
rect 791 -269 797 -235
rect 751 -307 797 -269
rect 751 -341 757 -307
rect 791 -341 797 -307
rect 751 -379 797 -341
rect 751 -413 757 -379
rect 791 -413 797 -379
rect 751 -451 797 -413
rect 751 -485 757 -451
rect 791 -485 797 -451
rect 751 -500 797 -485
rect 1009 485 1055 500
rect 1009 451 1015 485
rect 1049 451 1055 485
rect 1009 413 1055 451
rect 1009 379 1015 413
rect 1049 379 1055 413
rect 1009 341 1055 379
rect 1009 307 1015 341
rect 1049 307 1055 341
rect 1009 269 1055 307
rect 1009 235 1015 269
rect 1049 235 1055 269
rect 1009 197 1055 235
rect 1009 163 1015 197
rect 1049 163 1055 197
rect 1009 125 1055 163
rect 1009 91 1015 125
rect 1049 91 1055 125
rect 1009 53 1055 91
rect 1009 19 1015 53
rect 1049 19 1055 53
rect 1009 -19 1055 19
rect 1009 -53 1015 -19
rect 1049 -53 1055 -19
rect 1009 -91 1055 -53
rect 1009 -125 1015 -91
rect 1049 -125 1055 -91
rect 1009 -163 1055 -125
rect 1009 -197 1015 -163
rect 1049 -197 1055 -163
rect 1009 -235 1055 -197
rect 1009 -269 1015 -235
rect 1049 -269 1055 -235
rect 1009 -307 1055 -269
rect 1009 -341 1015 -307
rect 1049 -341 1055 -307
rect 1009 -379 1055 -341
rect 1009 -413 1015 -379
rect 1049 -413 1055 -379
rect 1009 -451 1055 -413
rect 1009 -485 1015 -451
rect 1049 -485 1055 -451
rect 1009 -500 1055 -485
rect 1267 485 1313 500
rect 1267 451 1273 485
rect 1307 451 1313 485
rect 1267 413 1313 451
rect 1267 379 1273 413
rect 1307 379 1313 413
rect 1267 341 1313 379
rect 1267 307 1273 341
rect 1307 307 1313 341
rect 1267 269 1313 307
rect 1267 235 1273 269
rect 1307 235 1313 269
rect 1267 197 1313 235
rect 1267 163 1273 197
rect 1307 163 1313 197
rect 1267 125 1313 163
rect 1267 91 1273 125
rect 1307 91 1313 125
rect 1267 53 1313 91
rect 1267 19 1273 53
rect 1307 19 1313 53
rect 1267 -19 1313 19
rect 1267 -53 1273 -19
rect 1307 -53 1313 -19
rect 1267 -91 1313 -53
rect 1267 -125 1273 -91
rect 1307 -125 1313 -91
rect 1267 -163 1313 -125
rect 1267 -197 1273 -163
rect 1307 -197 1313 -163
rect 1267 -235 1313 -197
rect 1267 -269 1273 -235
rect 1307 -269 1313 -235
rect 1267 -307 1313 -269
rect 1267 -341 1273 -307
rect 1307 -341 1313 -307
rect 1267 -379 1313 -341
rect 1267 -413 1273 -379
rect 1307 -413 1313 -379
rect 1267 -451 1313 -413
rect 1267 -485 1273 -451
rect 1307 -485 1313 -451
rect 1267 -500 1313 -485
rect 1525 485 1571 500
rect 1525 451 1531 485
rect 1565 451 1571 485
rect 1525 413 1571 451
rect 1525 379 1531 413
rect 1565 379 1571 413
rect 1525 341 1571 379
rect 1525 307 1531 341
rect 1565 307 1571 341
rect 1525 269 1571 307
rect 1525 235 1531 269
rect 1565 235 1571 269
rect 1525 197 1571 235
rect 1525 163 1531 197
rect 1565 163 1571 197
rect 1525 125 1571 163
rect 1525 91 1531 125
rect 1565 91 1571 125
rect 1525 53 1571 91
rect 1525 19 1531 53
rect 1565 19 1571 53
rect 1525 -19 1571 19
rect 1525 -53 1531 -19
rect 1565 -53 1571 -19
rect 1525 -91 1571 -53
rect 1525 -125 1531 -91
rect 1565 -125 1571 -91
rect 1525 -163 1571 -125
rect 1525 -197 1531 -163
rect 1565 -197 1571 -163
rect 1525 -235 1571 -197
rect 1525 -269 1531 -235
rect 1565 -269 1571 -235
rect 1525 -307 1571 -269
rect 1525 -341 1531 -307
rect 1565 -341 1571 -307
rect 1525 -379 1571 -341
rect 1525 -413 1531 -379
rect 1565 -413 1571 -379
rect 1525 -451 1571 -413
rect 1525 -485 1531 -451
rect 1565 -485 1571 -451
rect 1525 -500 1571 -485
rect 1783 485 1829 500
rect 1783 451 1789 485
rect 1823 451 1829 485
rect 1783 413 1829 451
rect 1783 379 1789 413
rect 1823 379 1829 413
rect 1783 341 1829 379
rect 1783 307 1789 341
rect 1823 307 1829 341
rect 1783 269 1829 307
rect 1783 235 1789 269
rect 1823 235 1829 269
rect 1783 197 1829 235
rect 1783 163 1789 197
rect 1823 163 1829 197
rect 1783 125 1829 163
rect 1783 91 1789 125
rect 1823 91 1829 125
rect 1783 53 1829 91
rect 1783 19 1789 53
rect 1823 19 1829 53
rect 1783 -19 1829 19
rect 1783 -53 1789 -19
rect 1823 -53 1829 -19
rect 1783 -91 1829 -53
rect 1783 -125 1789 -91
rect 1823 -125 1829 -91
rect 1783 -163 1829 -125
rect 1783 -197 1789 -163
rect 1823 -197 1829 -163
rect 1783 -235 1829 -197
rect 1783 -269 1789 -235
rect 1823 -269 1829 -235
rect 1783 -307 1829 -269
rect 1783 -341 1789 -307
rect 1823 -341 1829 -307
rect 1783 -379 1829 -341
rect 1783 -413 1789 -379
rect 1823 -413 1829 -379
rect 1783 -451 1829 -413
rect 1783 -485 1789 -451
rect 1823 -485 1829 -451
rect 1783 -500 1829 -485
rect -1773 -538 -1581 -532
rect -1773 -572 -1730 -538
rect -1696 -572 -1658 -538
rect -1624 -572 -1581 -538
rect -1773 -578 -1581 -572
rect -1515 -538 -1323 -532
rect -1515 -572 -1472 -538
rect -1438 -572 -1400 -538
rect -1366 -572 -1323 -538
rect -1515 -578 -1323 -572
rect -1257 -538 -1065 -532
rect -1257 -572 -1214 -538
rect -1180 -572 -1142 -538
rect -1108 -572 -1065 -538
rect -1257 -578 -1065 -572
rect -999 -538 -807 -532
rect -999 -572 -956 -538
rect -922 -572 -884 -538
rect -850 -572 -807 -538
rect -999 -578 -807 -572
rect -741 -538 -549 -532
rect -741 -572 -698 -538
rect -664 -572 -626 -538
rect -592 -572 -549 -538
rect -741 -578 -549 -572
rect -483 -538 -291 -532
rect -483 -572 -440 -538
rect -406 -572 -368 -538
rect -334 -572 -291 -538
rect -483 -578 -291 -572
rect -225 -538 -33 -532
rect -225 -572 -182 -538
rect -148 -572 -110 -538
rect -76 -572 -33 -538
rect -225 -578 -33 -572
rect 33 -538 225 -532
rect 33 -572 76 -538
rect 110 -572 148 -538
rect 182 -572 225 -538
rect 33 -578 225 -572
rect 291 -538 483 -532
rect 291 -572 334 -538
rect 368 -572 406 -538
rect 440 -572 483 -538
rect 291 -578 483 -572
rect 549 -538 741 -532
rect 549 -572 592 -538
rect 626 -572 664 -538
rect 698 -572 741 -538
rect 549 -578 741 -572
rect 807 -538 999 -532
rect 807 -572 850 -538
rect 884 -572 922 -538
rect 956 -572 999 -538
rect 807 -578 999 -572
rect 1065 -538 1257 -532
rect 1065 -572 1108 -538
rect 1142 -572 1180 -538
rect 1214 -572 1257 -538
rect 1065 -578 1257 -572
rect 1323 -538 1515 -532
rect 1323 -572 1366 -538
rect 1400 -572 1438 -538
rect 1472 -572 1515 -538
rect 1323 -578 1515 -572
rect 1581 -538 1773 -532
rect 1581 -572 1624 -538
rect 1658 -572 1696 -538
rect 1730 -572 1773 -538
rect 1581 -578 1773 -572
rect -963 -640 963 -634
rect -963 -674 -917 -640
rect -883 -674 -845 -640
rect -811 -674 -773 -640
rect -739 -674 -701 -640
rect -667 -674 -629 -640
rect -595 -674 -557 -640
rect -523 -674 -485 -640
rect -451 -674 -413 -640
rect -379 -674 -341 -640
rect -307 -674 -269 -640
rect -235 -674 -197 -640
rect -163 -674 -125 -640
rect -91 -674 -53 -640
rect -19 -674 19 -640
rect 53 -674 91 -640
rect 125 -674 163 -640
rect 197 -674 235 -640
rect 269 -674 307 -640
rect 341 -674 379 -640
rect 413 -674 451 -640
rect 485 -674 523 -640
rect 557 -674 595 -640
rect 629 -674 667 -640
rect 701 -674 739 -640
rect 773 -674 811 -640
rect 845 -674 883 -640
rect 917 -674 963 -640
rect -963 -680 963 -674
<< properties >>
string FIXED_BBOX -1920 -657 1920 657
<< end >>
