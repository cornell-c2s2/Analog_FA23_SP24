magic
tech sky130A
magscale 1 2
timestamp 1716868724
<< pwell >>
rect -315 -450 315 450
<< nmos >>
rect -129 -250 -29 250
rect 29 -250 129 250
<< ndiff >>
rect -187 221 -129 250
rect -187 187 -175 221
rect -141 187 -129 221
rect -187 153 -129 187
rect -187 119 -175 153
rect -141 119 -129 153
rect -187 85 -129 119
rect -187 51 -175 85
rect -141 51 -129 85
rect -187 17 -129 51
rect -187 -17 -175 17
rect -141 -17 -129 17
rect -187 -51 -129 -17
rect -187 -85 -175 -51
rect -141 -85 -129 -51
rect -187 -119 -129 -85
rect -187 -153 -175 -119
rect -141 -153 -129 -119
rect -187 -187 -129 -153
rect -187 -221 -175 -187
rect -141 -221 -129 -187
rect -187 -250 -129 -221
rect -29 221 29 250
rect -29 187 -17 221
rect 17 187 29 221
rect -29 153 29 187
rect -29 119 -17 153
rect 17 119 29 153
rect -29 85 29 119
rect -29 51 -17 85
rect 17 51 29 85
rect -29 17 29 51
rect -29 -17 -17 17
rect 17 -17 29 17
rect -29 -51 29 -17
rect -29 -85 -17 -51
rect 17 -85 29 -51
rect -29 -119 29 -85
rect -29 -153 -17 -119
rect 17 -153 29 -119
rect -29 -187 29 -153
rect -29 -221 -17 -187
rect 17 -221 29 -187
rect -29 -250 29 -221
rect 129 221 187 250
rect 129 187 141 221
rect 175 187 187 221
rect 129 153 187 187
rect 129 119 141 153
rect 175 119 187 153
rect 129 85 187 119
rect 129 51 141 85
rect 175 51 187 85
rect 129 17 187 51
rect 129 -17 141 17
rect 175 -17 187 17
rect 129 -51 187 -17
rect 129 -85 141 -51
rect 175 -85 187 -51
rect 129 -119 187 -85
rect 129 -153 141 -119
rect 175 -153 187 -119
rect 129 -187 187 -153
rect 129 -221 141 -187
rect 175 -221 187 -187
rect 129 -250 187 -221
<< ndiffc >>
rect -175 187 -141 221
rect -175 119 -141 153
rect -175 51 -141 85
rect -175 -17 -141 17
rect -175 -85 -141 -51
rect -175 -153 -141 -119
rect -175 -221 -141 -187
rect -17 187 17 221
rect -17 119 17 153
rect -17 51 17 85
rect -17 -17 17 17
rect -17 -85 17 -51
rect -17 -153 17 -119
rect -17 -221 17 -187
rect 141 187 175 221
rect 141 119 175 153
rect 141 51 175 85
rect 141 -17 175 17
rect 141 -85 175 -51
rect 141 -153 175 -119
rect 141 -221 175 -187
<< psubdiff >>
rect -289 390 -187 424
rect -153 390 -119 424
rect -85 390 -51 424
rect -17 390 17 424
rect 51 390 85 424
rect 119 390 153 424
rect 187 390 289 424
rect -289 323 -255 390
rect -289 255 -255 289
rect 255 323 289 390
rect 255 255 289 289
rect -289 187 -255 221
rect -289 119 -255 153
rect -289 51 -255 85
rect -289 -17 -255 17
rect -289 -85 -255 -51
rect -289 -153 -255 -119
rect -289 -221 -255 -187
rect 255 187 289 221
rect 255 119 289 153
rect 255 51 289 85
rect 255 -17 289 17
rect 255 -85 289 -51
rect 255 -153 289 -119
rect 255 -221 289 -187
rect -289 -289 -255 -255
rect -289 -390 -255 -323
rect 255 -289 289 -255
rect 255 -390 289 -323
rect -289 -424 -187 -390
rect -153 -424 -119 -390
rect -85 -424 -51 -390
rect -17 -424 17 -390
rect 51 -424 85 -390
rect 119 -424 153 -390
rect 187 -424 289 -390
<< psubdiffcont >>
rect -187 390 -153 424
rect -119 390 -85 424
rect -51 390 -17 424
rect 17 390 51 424
rect 85 390 119 424
rect 153 390 187 424
rect -289 289 -255 323
rect -289 221 -255 255
rect 255 289 289 323
rect -289 153 -255 187
rect -289 85 -255 119
rect -289 17 -255 51
rect -289 -51 -255 -17
rect -289 -119 -255 -85
rect -289 -187 -255 -153
rect -289 -255 -255 -221
rect 255 221 289 255
rect 255 153 289 187
rect 255 85 289 119
rect 255 17 289 51
rect 255 -51 289 -17
rect 255 -119 289 -85
rect 255 -187 289 -153
rect -289 -323 -255 -289
rect 255 -255 289 -221
rect 255 -323 289 -289
rect -187 -424 -153 -390
rect -119 -424 -85 -390
rect -51 -424 -17 -390
rect 17 -424 51 -390
rect 85 -424 119 -390
rect 153 -424 187 -390
<< poly >>
rect -129 322 -29 338
rect -129 288 -96 322
rect -62 288 -29 322
rect -129 250 -29 288
rect 29 322 129 338
rect 29 288 62 322
rect 96 288 129 322
rect 29 250 129 288
rect -129 -288 -29 -250
rect -129 -322 -96 -288
rect -62 -322 -29 -288
rect -129 -338 -29 -322
rect 29 -288 129 -250
rect 29 -322 62 -288
rect 96 -322 129 -288
rect 29 -338 129 -322
<< polycont >>
rect -96 288 -62 322
rect 62 288 96 322
rect -96 -322 -62 -288
rect 62 -322 96 -288
<< locali >>
rect -289 390 -187 424
rect -153 390 -119 424
rect -85 390 -51 424
rect -17 390 17 424
rect 51 390 85 424
rect 119 390 153 424
rect 187 390 289 424
rect -289 323 -255 390
rect 255 323 289 390
rect -289 255 -255 289
rect -129 288 -96 322
rect -62 288 -29 322
rect 29 288 62 322
rect 96 288 129 322
rect 255 255 289 289
rect -289 187 -255 221
rect -289 119 -255 153
rect -289 51 -255 85
rect -289 -17 -255 17
rect -289 -85 -255 -51
rect -289 -153 -255 -119
rect -289 -221 -255 -187
rect -175 233 -141 254
rect -175 161 -141 187
rect -175 89 -141 119
rect -175 17 -141 51
rect -175 -51 -141 -17
rect -175 -119 -141 -89
rect -175 -187 -141 -161
rect -175 -254 -141 -233
rect -17 233 17 254
rect -17 161 17 187
rect -17 89 17 119
rect -17 17 17 51
rect -17 -51 17 -17
rect -17 -119 17 -89
rect -17 -187 17 -161
rect -17 -254 17 -233
rect 141 233 175 254
rect 141 161 175 187
rect 141 89 175 119
rect 141 17 175 51
rect 141 -51 175 -17
rect 141 -119 175 -89
rect 141 -187 175 -161
rect 141 -254 175 -233
rect 255 187 289 221
rect 255 119 289 153
rect 255 51 289 85
rect 255 -17 289 17
rect 255 -85 289 -51
rect 255 -153 289 -119
rect 255 -221 289 -187
rect -289 -289 -255 -255
rect -129 -322 -96 -288
rect -62 -322 -29 -288
rect 29 -322 62 -288
rect 96 -322 129 -288
rect 255 -289 289 -255
rect -289 -390 -255 -323
rect 255 -390 289 -323
rect -289 -424 -187 -390
rect -153 -424 -119 -390
rect -85 -424 -51 -390
rect -17 -424 17 -390
rect 51 -424 85 -390
rect 119 -424 153 -390
rect 187 -424 289 -390
<< viali >>
rect -96 288 -62 322
rect 62 288 96 322
rect -175 221 -141 233
rect -175 199 -141 221
rect -175 153 -141 161
rect -175 127 -141 153
rect -175 85 -141 89
rect -175 55 -141 85
rect -175 -17 -141 17
rect -175 -85 -141 -55
rect -175 -89 -141 -85
rect -175 -153 -141 -127
rect -175 -161 -141 -153
rect -175 -221 -141 -199
rect -175 -233 -141 -221
rect -17 221 17 233
rect -17 199 17 221
rect -17 153 17 161
rect -17 127 17 153
rect -17 85 17 89
rect -17 55 17 85
rect -17 -17 17 17
rect -17 -85 17 -55
rect -17 -89 17 -85
rect -17 -153 17 -127
rect -17 -161 17 -153
rect -17 -221 17 -199
rect -17 -233 17 -221
rect 141 221 175 233
rect 141 199 175 221
rect 141 153 175 161
rect 141 127 175 153
rect 141 85 175 89
rect 141 55 175 85
rect 141 -17 175 17
rect 141 -85 175 -55
rect 141 -89 175 -85
rect 141 -153 175 -127
rect 141 -161 175 -153
rect 141 -221 175 -199
rect 141 -233 175 -221
rect -96 -322 -62 -288
rect 62 -322 96 -288
<< metal1 >>
rect -125 322 -33 328
rect -125 288 -96 322
rect -62 288 -33 322
rect -125 282 -33 288
rect 33 322 125 328
rect 33 288 62 322
rect 96 288 125 322
rect 33 282 125 288
rect -181 233 -135 250
rect -181 199 -175 233
rect -141 199 -135 233
rect -181 161 -135 199
rect -181 127 -175 161
rect -141 127 -135 161
rect -181 89 -135 127
rect -181 55 -175 89
rect -141 55 -135 89
rect -181 17 -135 55
rect -181 -17 -175 17
rect -141 -17 -135 17
rect -181 -55 -135 -17
rect -181 -89 -175 -55
rect -141 -89 -135 -55
rect -181 -127 -135 -89
rect -181 -161 -175 -127
rect -141 -161 -135 -127
rect -181 -199 -135 -161
rect -181 -233 -175 -199
rect -141 -233 -135 -199
rect -181 -250 -135 -233
rect -23 233 23 250
rect -23 199 -17 233
rect 17 199 23 233
rect -23 161 23 199
rect -23 127 -17 161
rect 17 127 23 161
rect -23 89 23 127
rect -23 55 -17 89
rect 17 55 23 89
rect -23 17 23 55
rect -23 -17 -17 17
rect 17 -17 23 17
rect -23 -55 23 -17
rect -23 -89 -17 -55
rect 17 -89 23 -55
rect -23 -127 23 -89
rect -23 -161 -17 -127
rect 17 -161 23 -127
rect -23 -199 23 -161
rect -23 -233 -17 -199
rect 17 -233 23 -199
rect -23 -250 23 -233
rect 135 233 181 250
rect 135 199 141 233
rect 175 199 181 233
rect 135 161 181 199
rect 135 127 141 161
rect 175 127 181 161
rect 135 89 181 127
rect 135 55 141 89
rect 175 55 181 89
rect 135 17 181 55
rect 135 -17 141 17
rect 175 -17 181 17
rect 135 -55 181 -17
rect 135 -89 141 -55
rect 175 -89 181 -55
rect 135 -127 181 -89
rect 135 -161 141 -127
rect 175 -161 181 -127
rect 135 -199 181 -161
rect 135 -233 141 -199
rect 175 -233 181 -199
rect 135 -250 181 -233
rect -125 -288 -33 -282
rect -125 -322 -96 -288
rect -62 -322 -33 -288
rect -125 -328 -33 -322
rect 33 -288 125 -282
rect 33 -322 62 -288
rect 96 -322 125 -288
rect 33 -328 125 -322
<< properties >>
string FIXED_BBOX -272 -407 272 407
<< end >>
