magic
tech sky130A
magscale 1 2
timestamp 1712340852
<< nwell >>
rect -396 -261 396 261
<< pmos >>
rect -200 -42 200 42
<< pdiff >>
rect -258 30 -200 42
rect -258 -30 -246 30
rect -212 -30 -200 30
rect -258 -42 -200 -30
rect 200 30 258 42
rect 200 -30 212 30
rect 246 -30 258 30
rect 200 -42 258 -30
<< pdiffc >>
rect -246 -30 -212 30
rect 212 -30 246 30
<< nsubdiff >>
rect -360 191 -264 225
rect 264 191 360 225
rect -360 129 -326 191
rect 326 129 360 191
rect -360 -191 -326 -129
rect 326 -191 360 -129
rect -360 -225 360 -191
<< nsubdiffcont >>
rect -264 191 264 225
rect -360 -129 -326 129
rect 326 -129 360 129
<< poly >>
rect -200 123 200 139
rect -200 89 -184 123
rect 184 89 200 123
rect -200 42 200 89
rect -200 -89 200 -42
rect -200 -123 -184 -89
rect 184 -123 200 -89
rect -200 -139 200 -123
<< polycont >>
rect -184 89 184 123
rect -184 -123 184 -89
<< locali >>
rect -360 191 -264 225
rect 264 191 360 225
rect -360 129 -326 191
rect 326 129 360 191
rect -200 89 -184 123
rect 184 89 200 123
rect -246 30 -212 46
rect -246 -46 -212 -30
rect 212 30 246 46
rect 212 -46 246 -30
rect -200 -123 -184 -89
rect 184 -123 200 -89
rect -360 -191 -326 -129
rect 326 -191 360 -129
rect -360 -225 360 -191
<< viali >>
rect -184 89 184 123
rect -246 -30 -212 30
rect 212 -30 246 30
rect -184 -123 184 -89
<< metal1 >>
rect -196 123 196 129
rect -196 89 -184 123
rect 184 89 196 123
rect -196 83 196 89
rect -252 30 -206 42
rect -252 -30 -246 30
rect -212 -30 -206 30
rect -252 -42 -206 -30
rect 206 30 252 42
rect 206 -30 212 30
rect 246 -30 252 30
rect 206 -42 252 -30
rect -196 -89 196 -83
rect -196 -123 -184 -89
rect 184 -123 196 -89
rect -196 -129 196 -123
<< properties >>
string FIXED_BBOX -343 -208 343 208
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 0.42 l 2.0 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
