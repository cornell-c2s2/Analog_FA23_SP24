* NGSPICE file created from PTAT_v0p0p0_mag_ext_flat.ext - technology: sky130A

.subckt PTAT_v0p0p0_mag_ext_flat VDD VOUT VSS
X0 a_n2389_n1015.t16 VSS.t20 VSS.t17 sky130_fd_pr__res_xhigh_po_5p73 l=85.8
X1 a_n2211_n1015.t19 a_n2331_n1103.t4 a_n2389_n1015.t3 VSS.t3 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X2 a_n2211_n1015.t18 a_n2331_n1103.t5 a_n2389_n1015.t6 VSS.t6 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X3 a_n2211_n1015.t17 a_n2331_n1103.t6 a_n2389_n1015.t7 VSS.t7 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X4 a_n2211_n1015.t16 a_n2331_n1103.t7 a_n2389_n1015.t4 VSS.t4 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X5 a_n2211_n1015.t23 a_n2211_n1015.t22 VDD.t5 VDD.t4 sky130_fd_pr__pfet_01v8_lvt ad=5.51 pd=38.6 as=5.51 ps=38.6 w=19 l=1
X6 a_n2211_n1015.t15 a_n2331_n1103.t8 a_n2389_n1015.t8 VSS.t8 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X7 VOUT.t0 a_n2211_n1015.t24 VDD.t3 VDD.t2 sky130_fd_pr__pfet_01v8_lvt ad=5.51 pd=38.6 as=5.51 ps=38.6 w=19 l=1
X8 a_n2211_n1015.t14 a_n2331_n1103.t9 a_n2389_n1015.t10 VSS.t10 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X9 a_n2211_n1015.t13 a_n2331_n1103.t10 a_n2389_n1015.t0 VSS.t0 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X10 VSS.t13 VOUT.t1 VOUT.t2 VSS.t12 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X11 a_n2211_n1015.t12 a_n2331_n1103.t11 a_n2389_n1015.t17 VSS.t21 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X12 a_n2389_n1015.t14 VSS.t18 VSS.t17 sky130_fd_pr__res_xhigh_po_5p73 l=85.8
X13 a_n2331_n1103.t1 a_n2331_n1103.t0 VSS.t26 VSS.t25 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X14 VDD.t1 a_n2211_n1015.t25 a_n2331_n1103.t3 VDD.t0 sky130_fd_pr__pfet_01v8_lvt ad=5.51 pd=38.6 as=5.51 ps=38.6 w=19 l=1
X15 a_n2211_n1015.t11 a_n2331_n1103.t12 a_n2389_n1015.t15 VSS.t19 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X16 a_n2211_n1015.t10 a_n2331_n1103.t13 a_n2389_n1015.t13 VSS.t16 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X17 a_n2211_n1015.t21 a_n2211_n1015.t20 a_n2331_n1103.t2 VSS.t15 sky130_fd_pr__nfet_01v8_lvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X18 a_n2211_n1015.t9 a_n2331_n1103.t14 a_n2389_n1015.t20 VSS.t24 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X19 a_n2211_n1015.t8 a_n2331_n1103.t15 a_n2389_n1015.t18 VSS.t22 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X20 a_n2211_n1015.t7 a_n2331_n1103.t16 a_n2389_n1015.t19 VSS.t23 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X21 a_n2211_n1015.t6 a_n2331_n1103.t17 a_n2389_n1015.t9 VSS.t9 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X22 a_n2211_n1015.t5 a_n2331_n1103.t18 a_n2389_n1015.t11 VSS.t11 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X23 a_n2211_n1015.t4 a_n2331_n1103.t19 a_n2389_n1015.t12 VSS.t14 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X24 a_n2211_n1015.t3 a_n2331_n1103.t20 a_n2389_n1015.t1 VSS.t1 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X25 a_n2211_n1015.t2 a_n2331_n1103.t21 a_n2389_n1015.t21 VSS.t27 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X26 a_n2211_n1015.t1 a_n2331_n1103.t22 a_n2389_n1015.t5 VSS.t5 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X27 a_n2211_n1015.t0 a_n2331_n1103.t23 a_n2389_n1015.t2 VSS.t2 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
R0 a_n2389_n1015.n0 a_n2389_n1015.t1 5.73525
R1 a_n2389_n1015.n18 a_n2389_n1015.t17 5.34571
R2 a_n2389_n1015.n0 a_n2389_n1015.t3 5.18362
R3 a_n2389_n1015.n1 a_n2389_n1015.t20 5.18362
R4 a_n2389_n1015.n2 a_n2389_n1015.t9 5.18362
R5 a_n2389_n1015.n3 a_n2389_n1015.t7 5.18362
R6 a_n2389_n1015.n4 a_n2389_n1015.t19 5.18362
R7 a_n2389_n1015.n5 a_n2389_n1015.t12 5.18362
R8 a_n2389_n1015.n6 a_n2389_n1015.t0 5.18362
R9 a_n2389_n1015.n7 a_n2389_n1015.t13 5.18362
R10 a_n2389_n1015.n8 a_n2389_n1015.t2 5.18362
R11 a_n2389_n1015.n9 a_n2389_n1015.t18 5.18362
R12 a_n2389_n1015.n10 a_n2389_n1015.t4 5.18362
R13 a_n2389_n1015.n11 a_n2389_n1015.t10 5.18362
R14 a_n2389_n1015.n12 a_n2389_n1015.t11 5.18362
R15 a_n2389_n1015.n13 a_n2389_n1015.t6 5.18362
R16 a_n2389_n1015.n14 a_n2389_n1015.t5 5.18362
R17 a_n2389_n1015.n15 a_n2389_n1015.t15 5.18362
R18 a_n2389_n1015.n16 a_n2389_n1015.t8 5.18362
R19 a_n2389_n1015.n17 a_n2389_n1015.t21 5.18362
R20 a_n2389_n1015.n19 a_n2389_n1015.t16 2.79552
R21 a_n2389_n1015.t14 a_n2389_n1015.n19 2.38201
R22 a_n2389_n1015.n9 a_n2389_n1015.n8 1.10376
R23 a_n2389_n1015.n1 a_n2389_n1015.n0 0.55213
R24 a_n2389_n1015.n2 a_n2389_n1015.n1 0.55213
R25 a_n2389_n1015.n3 a_n2389_n1015.n2 0.55213
R26 a_n2389_n1015.n4 a_n2389_n1015.n3 0.55213
R27 a_n2389_n1015.n5 a_n2389_n1015.n4 0.55213
R28 a_n2389_n1015.n6 a_n2389_n1015.n5 0.55213
R29 a_n2389_n1015.n7 a_n2389_n1015.n6 0.55213
R30 a_n2389_n1015.n8 a_n2389_n1015.n7 0.55213
R31 a_n2389_n1015.n10 a_n2389_n1015.n9 0.55213
R32 a_n2389_n1015.n11 a_n2389_n1015.n10 0.55213
R33 a_n2389_n1015.n12 a_n2389_n1015.n11 0.55213
R34 a_n2389_n1015.n13 a_n2389_n1015.n12 0.55213
R35 a_n2389_n1015.n14 a_n2389_n1015.n13 0.55213
R36 a_n2389_n1015.n15 a_n2389_n1015.n14 0.55213
R37 a_n2389_n1015.n16 a_n2389_n1015.n15 0.55213
R38 a_n2389_n1015.n17 a_n2389_n1015.n16 0.512683
R39 a_n2389_n1015.n19 a_n2389_n1015.n18 0.168655
R40 a_n2389_n1015.n18 a_n2389_n1015.n17 0.0581389
R41 VSS.n19 VSS.n3 3876.26
R42 VSS.n58 VSS.n46 3876.26
R43 VSS.n218 VSS.n206 1176.21
R44 VSS.n198 VSS.n190 1176.21
R45 VSS.n183 VSS.n175 1176.21
R46 VSS.n168 VSS.n160 1176.21
R47 VSS.n153 VSS.n145 1176.21
R48 VSS.n133 VSS.n125 1176.21
R49 VSS.n118 VSS.n110 1176.21
R50 VSS.n103 VSS.n95 1176.21
R51 VSS.n88 VSS.n80 1176.21
R52 VSS.n411 VSS.n34 1176.21
R53 VSS.n404 VSS.n403 1176.21
R54 VSS.n389 VSS.n388 1176.21
R55 VSS.n374 VSS.n373 1176.21
R56 VSS.n359 VSS.n358 1176.21
R57 VSS.n344 VSS.n343 1176.21
R58 VSS.n327 VSS.n326 1176.21
R59 VSS.n312 VSS.n311 1176.21
R60 VSS.n296 VSS.n295 1176.21
R61 VSS.n281 VSS.n280 1176.21
R62 VSS.n266 VSS.n265 1176.21
R63 VSS.n245 VSS.n244 1176.21
R64 VSS.n220 VSS.n219 1176.21
R65 VSS.n200 VSS.n199 1176.21
R66 VSS.n185 VSS.n184 1176.21
R67 VSS.n170 VSS.n169 1176.21
R68 VSS.n155 VSS.n154 1176.21
R69 VSS.n135 VSS.n134 1176.21
R70 VSS.n120 VSS.n119 1176.21
R71 VSS.n105 VSS.n104 1176.21
R72 VSS.n90 VSS.n89 1176.21
R73 VSS.n412 VSS.n30 1176.21
R74 VSS.n402 VSS.n397 1176.21
R75 VSS.n387 VSS.n382 1176.21
R76 VSS.n372 VSS.n367 1176.21
R77 VSS.n357 VSS.n352 1176.21
R78 VSS.n342 VSS.n337 1176.21
R79 VSS.n325 VSS.n320 1176.21
R80 VSS.n310 VSS.n305 1176.21
R81 VSS.n294 VSS.n286 1176.21
R82 VSS.n279 VSS.n271 1176.21
R83 VSS.n264 VSS.n254 1176.21
R84 VSS.n243 VSS.n228 1176.21
R85 VSS.n290 VSS.n289 201.412
R86 VSS.n275 VSS.n274 201.412
R87 VSS.n194 VSS.n193 201.412
R88 VSS.n179 VSS.n178 201.412
R89 VSS.n149 VSS.n148 201.412
R90 VSS.n114 VSS.n113 201.412
R91 VSS.n84 VSS.n83 201.412
R92 VSS.n99 VSS.n98 201.412
R93 VSS.n129 VSS.n128 201.412
R94 VSS.n164 VSS.n163 201.412
R95 VSS.n258 VSS.n257 201.412
R96 VSS.n218 VSS.n205 162.236
R97 VSS.t6 VSS.n144 143.446
R98 VSS.n304 VSS.n303 122.082
R99 VSS.n237 VSS.n231 116.329
R100 VSS.t12 VSS.n33 101.605
R101 VSS.t1 VSS.n396 101.605
R102 VSS.t3 VSS.n381 101.605
R103 VSS.t24 VSS.n366 101.605
R104 VSS.t9 VSS.n351 101.605
R105 VSS.t7 VSS.n336 101.605
R106 VSS.t23 VSS.n319 101.605
R107 VSS.n210 VSS.n209 64.093
R108 VSS.n213 VSS.n212 49.3181
R109 VSS.n238 VSS.n237 49.3181
R110 VSS.t14 VSS.n304 41.543
R111 VSS.n426 VSS.t13 26.8697
R112 VSS.n214 VSS.n213 13.4405
R113 VSS.n423 VSS.n422 9.3005
R114 VSS.n333 VSS.n332 9.3005
R115 VSS.n142 VSS.n141 9.3005
R116 VSS.n55 VSS.n54 9.3005
R117 VSS.n457 VSS.n456 9.3005
R118 VSS.n235 VSS.n234 7.12189
R119 VSS.n139 VSS.n138 4.90717
R120 VSS.n227 VSS.t26 4.78444
R121 VSS.n227 VSS.n225 4.5005
R122 VSS.n227 VSS.n226 4.5005
R123 VSS.n428 VSS.n427 4.4805
R124 VSS.n416 VSS.n415 4.4805
R125 VSS.n425 VSS.n424 3.84205
R126 VSS.n67 VSS.n35 3.38533
R127 VSS.n53 VSS.n51 3.20453
R128 VSS.t22 VSS.t15 3.05252
R129 VSS.n59 VSS.n45 3.05252
R130 VSS.n21 VSS.t18 2.36824
R131 VSS.n15 VSS.t20 2.36824
R132 VSS.n53 VSS.n52 1.85757
R133 VSS.n12 VSS.n11 1.70717
R134 VSS.n239 VSS.n238 1.49383
R135 VSS.n66 VSS.n64 1.40675
R136 VSS.n62 VSS.n42 1.40675
R137 VSS.n50 VSS.n48 1.3822
R138 VSS.n56 VSS.n55 1.3822
R139 VSS.n435 VSS.n434 1.2805
R140 VSS.n454 VSS.n442 1.2805
R141 VSS VSS.n27 0.647262
R142 VSS.n37 VSS.n36 0.549071
R143 VSS.n249 VSS.n248 0.427167
R144 VSS.n5 VSS.n4 0.427167
R145 VSS.n414 VSS.n29 0.352931
R146 VSS.n400 VSS.n399 0.352931
R147 VSS.n385 VSS.n384 0.352931
R148 VSS.n370 VSS.n369 0.352931
R149 VSS.n355 VSS.n354 0.352931
R150 VSS.n340 VSS.n339 0.352931
R151 VSS.n323 VSS.n322 0.352931
R152 VSS.n308 VSS.n307 0.352931
R153 VSS.n292 VSS.n291 0.352931
R154 VSS.n277 VSS.n276 0.352931
R155 VSS.n241 VSS.n240 0.352931
R156 VSS.n216 VSS.n215 0.352931
R157 VSS.n196 VSS.n195 0.352931
R158 VSS.n181 VSS.n180 0.352931
R159 VSS.n166 VSS.n165 0.352931
R160 VSS.n151 VSS.n150 0.352931
R161 VSS.n131 VSS.n130 0.352931
R162 VSS.n116 VSS.n115 0.352931
R163 VSS.n101 VSS.n100 0.352931
R164 VSS.n86 VSS.n85 0.352931
R165 VSS.n262 VSS.n261 0.347722
R166 VSS.n438 VSS.n435 0.3205
R167 VSS.n417 VSS.n414 0.302583
R168 VSS.n457 VSS.n455 0.227666
R169 VSS.n409 VSS.n408 0.141472
R170 VSS.n408 VSS.n406 0.141472
R171 VSS.n406 VSS.n393 0.141472
R172 VSS.n393 VSS.n391 0.141472
R173 VSS.n391 VSS.n378 0.141472
R174 VSS.n378 VSS.n376 0.141472
R175 VSS.n376 VSS.n363 0.141472
R176 VSS.n363 VSS.n361 0.141472
R177 VSS.n361 VSS.n348 0.141472
R178 VSS.n348 VSS.n346 0.141472
R179 VSS.n331 VSS.n329 0.141472
R180 VSS.n329 VSS.n316 0.141472
R181 VSS.n316 VSS.n314 0.141472
R182 VSS.n314 VSS.n300 0.141472
R183 VSS.n300 VSS.n298 0.141472
R184 VSS.n298 VSS.n285 0.141472
R185 VSS.n285 VSS.n283 0.141472
R186 VSS.n283 VSS.n270 0.141472
R187 VSS.n270 VSS.n268 0.141472
R188 VSS.n250 VSS.n247 0.141472
R189 VSS.n224 VSS.n222 0.141472
R190 VSS.n222 VSS.n204 0.141472
R191 VSS.n204 VSS.n202 0.141472
R192 VSS.n202 VSS.n189 0.141472
R193 VSS.n189 VSS.n187 0.141472
R194 VSS.n187 VSS.n174 0.141472
R195 VSS.n174 VSS.n172 0.141472
R196 VSS.n172 VSS.n159 0.141472
R197 VSS.n159 VSS.n157 0.141472
R198 VSS.n140 VSS.n137 0.141472
R199 VSS.n137 VSS.n124 0.141472
R200 VSS.n124 VSS.n122 0.141472
R201 VSS.n122 VSS.n109 0.141472
R202 VSS.n109 VSS.n107 0.141472
R203 VSS.n107 VSS.n94 0.141472
R204 VSS.n94 VSS.n92 0.141472
R205 VSS.n92 VSS.n79 0.141472
R206 VSS.n79 VSS.n77 0.141472
R207 VSS.n25 VSS.n23 0.139634
R208 VSS.n21 VSS.n2 0.139634
R209 VSS.n10 VSS.n8 0.137205
R210 VSS.n15 VSS.n14 0.137205
R211 VSS.n268 VSS.n253 0.136611
R212 VSS.n44 VSS.n43 0.134262
R213 VSS.n55 VSS.n53 0.127732
R214 VSS.n157 VSS.n143 0.1255
R215 VSS.n77 VSS.n71 0.117167
R216 VSS.n212 VSS.n211 0.10956
R217 VSS.n211 VSS.n210 0.10956
R218 VSS.n237 VSS.n236 0.10956
R219 VSS.n236 VSS.n235 0.10956
R220 VSS.n231 VSS.n230 0.0944005
R221 VSS.n230 VSS.n229 0.0944005
R222 VSS.n419 VSS.n417 0.0920099
R223 VSS.n42 VSS.n40 0.0853214
R224 VSS.n346 VSS.n333 0.0838333
R225 VSS VSS.n457 0.0771509
R226 VSS.n227 VSS.n224 0.0727222
R227 VSS.n247 VSS.n227 0.06925
R228 VSS.n423 VSS.n421 0.0589677
R229 VSS.n333 VSS.n331 0.0581389
R230 VSS.n67 VSS.n66 0.0540714
R231 VSS.n421 VSS.n419 0.0367903
R232 VSS.n40 VSS.n39 0.0339821
R233 VSS.n27 VSS.n26 0.0321352
R234 VSS.n56 VSS.n50 0.03175
R235 VSS.n441 VSS.n440 0.0179743
R236 VSS.n64 VSS.n62 0.016125
R237 VSS.n148 VSS.n147 0.015169
R238 VSS.n147 VSS.n146 0.015169
R239 VSS.n113 VSS.n112 0.015169
R240 VSS.n112 VSS.n111 0.015169
R241 VSS.n83 VSS.n82 0.015169
R242 VSS.n82 VSS.n81 0.015169
R243 VSS.n98 VSS.n97 0.015169
R244 VSS.n97 VSS.n96 0.015169
R245 VSS.n128 VSS.n127 0.015169
R246 VSS.n127 VSS.n126 0.015169
R247 VSS.n163 VSS.n162 0.015169
R248 VSS.n162 VSS.n161 0.015169
R249 VSS.n178 VSS.n177 0.015169
R250 VSS.n177 VSS.n176 0.015169
R251 VSS.n193 VSS.n192 0.015169
R252 VSS.n192 VSS.n191 0.015169
R253 VSS.n208 VSS.n207 0.015169
R254 VSS.n209 VSS.n208 0.015169
R255 VSS.n233 VSS.n232 0.015169
R256 VSS.n234 VSS.n233 0.015169
R257 VSS.n257 VSS.n256 0.015169
R258 VSS.n256 VSS.n255 0.015169
R259 VSS.n289 VSS.n288 0.015169
R260 VSS.n288 VSS.n287 0.015169
R261 VSS.n274 VSS.n273 0.015169
R262 VSS.n273 VSS.n272 0.015169
R263 VSS.n302 VSS.n301 0.015169
R264 VSS.n303 VSS.n302 0.015169
R265 VSS.n45 VSS.n44 0.015169
R266 VSS.n32 VSS.n31 0.015169
R267 VSS.n33 VSS.n32 0.015169
R268 VSS.n380 VSS.n379 0.015169
R269 VSS.n381 VSS.n380 0.015169
R270 VSS.n350 VSS.n349 0.015169
R271 VSS.n351 VSS.n350 0.015169
R272 VSS.n318 VSS.n317 0.015169
R273 VSS.n319 VSS.n318 0.015169
R274 VSS.n335 VSS.n334 0.015169
R275 VSS.n336 VSS.n335 0.015169
R276 VSS.n365 VSS.n364 0.015169
R277 VSS.n366 VSS.n365 0.015169
R278 VSS.n395 VSS.n394 0.015169
R279 VSS.n396 VSS.n395 0.015169
R280 VSS.n14 VSS.n13 0.0130883
R281 VSS.n2 VSS.n0 0.0122049
R282 VSS.n8 VSS.n6 0.0122049
R283 VSS.n71 VSS.n69 0.0109167
R284 VSS.n143 VSS.n142 0.0102222
R285 VSS.n71 VSS.n70 0.00959091
R286 VSS.n13 VSS.n12 0.00904795
R287 VSS.n431 VSS.n423 0.00856452
R288 VSS.n417 VSS.n416 0.00769258
R289 VSS.n429 VSS.n428 0.00769258
R290 VSS.n450 VSS.n449 0.00744444
R291 VSS.n6 VSS.n5 0.00738379
R292 VSS.n39 VSS.n38 0.00719643
R293 VSS.n142 VSS.n140 0.00675
R294 VSS.n69 VSS.n68 0.0066794
R295 VSS.n38 VSS.n37 0.0066794
R296 VSS.n69 VSS.n67 0.00605556
R297 VSS.n27 VSS.n25 0.00580035
R298 VSS.n261 VSS.n259 0.00570833
R299 VSS.n240 VSS.n239 0.00438796
R300 VSS.n259 VSS.n258 0.00438796
R301 VSS.n165 VSS.n164 0.00438796
R302 VSS.n130 VSS.n129 0.00438796
R303 VSS.n100 VSS.n99 0.00438796
R304 VSS.n85 VSS.n84 0.00438796
R305 VSS.n115 VSS.n114 0.00438796
R306 VSS.n150 VSS.n149 0.00438796
R307 VSS.n180 VSS.n179 0.00438796
R308 VSS.n195 VSS.n194 0.00438796
R309 VSS.n215 VSS.n214 0.00438796
R310 VSS.n399 VSS.n398 0.00438796
R311 VSS.n369 VSS.n368 0.00438796
R312 VSS.n339 VSS.n338 0.00438796
R313 VSS.n307 VSS.n306 0.00438796
R314 VSS.n276 VSS.n275 0.00438796
R315 VSS.n291 VSS.n290 0.00438796
R316 VSS.n322 VSS.n321 0.00438796
R317 VSS.n354 VSS.n353 0.00438796
R318 VSS.n384 VSS.n383 0.00438796
R319 VSS.n29 VSS.n28 0.00438796
R320 VSS.n408 VSS.n407 0.00438796
R321 VSS.n393 VSS.n392 0.00438796
R322 VSS.n378 VSS.n377 0.00438796
R323 VSS.n363 VSS.n362 0.00438796
R324 VSS.n348 VSS.n347 0.00438796
R325 VSS.n331 VSS.n330 0.00438796
R326 VSS.n316 VSS.n315 0.00438796
R327 VSS.n300 VSS.n299 0.00438796
R328 VSS.n285 VSS.n284 0.00438796
R329 VSS.n270 VSS.n269 0.00438796
R330 VSS.n250 VSS.n249 0.00438796
R331 VSS.n224 VSS.n223 0.00438796
R332 VSS.n204 VSS.n203 0.00438796
R333 VSS.n189 VSS.n188 0.00438796
R334 VSS.n174 VSS.n173 0.00438796
R335 VSS.n159 VSS.n158 0.00438796
R336 VSS.n140 VSS.n139 0.00438796
R337 VSS.n124 VSS.n123 0.00438796
R338 VSS.n109 VSS.n108 0.00438796
R339 VSS.n94 VSS.n93 0.00438796
R340 VSS.n79 VSS.n78 0.00438796
R341 VSS.n253 VSS.n251 0.00397222
R342 VSS.n15 VSS.n10 0.00359187
R343 VSS.n73 VSS.n72 0.00299232
R344 VSS.n440 VSS.n439 0.00253688
R345 VSS.n431 VSS.n430 0.00253688
R346 VSS.n87 VSS.n86 0.00250907
R347 VSS.n102 VSS.n101 0.00250907
R348 VSS.n117 VSS.n116 0.00250907
R349 VSS.n132 VSS.n131 0.00250907
R350 VSS.n152 VSS.n151 0.00250907
R351 VSS.n167 VSS.n166 0.00250907
R352 VSS.n182 VSS.n181 0.00250907
R353 VSS.n217 VSS.n216 0.00250907
R354 VSS.n197 VSS.n196 0.00250907
R355 VSS.n263 VSS.n262 0.00250907
R356 VSS.n278 VSS.n277 0.00250907
R357 VSS.n293 VSS.n292 0.00250907
R358 VSS.n242 VSS.n241 0.00250907
R359 VSS.n309 VSS.n308 0.00250907
R360 VSS.n324 VSS.n323 0.00250907
R361 VSS.n341 VSS.n340 0.00250907
R362 VSS.n356 VSS.n355 0.00250907
R363 VSS.n371 VSS.n370 0.00250907
R364 VSS.n386 VSS.n385 0.00250907
R365 VSS.n401 VSS.n400 0.00250907
R366 VSS.n414 VSS.n413 0.00250907
R367 VSS.n410 VSS.n409 0.00250907
R368 VSS.n406 VSS.n405 0.00250907
R369 VSS.n391 VSS.n390 0.00250907
R370 VSS.n376 VSS.n375 0.00250907
R371 VSS.n361 VSS.n360 0.00250907
R372 VSS.n346 VSS.n345 0.00250907
R373 VSS.n329 VSS.n328 0.00250907
R374 VSS.n314 VSS.n313 0.00250907
R375 VSS.n298 VSS.n297 0.00250907
R376 VSS.n283 VSS.n282 0.00250907
R377 VSS.n268 VSS.n267 0.00250907
R378 VSS.n247 VSS.n246 0.00250907
R379 VSS.n222 VSS.n221 0.00250907
R380 VSS.n202 VSS.n201 0.00250907
R381 VSS.n187 VSS.n186 0.00250907
R382 VSS.n172 VSS.n171 0.00250907
R383 VSS.n157 VSS.n156 0.00250907
R384 VSS.n137 VSS.n136 0.00250907
R385 VSS.n122 VSS.n121 0.00250907
R386 VSS.n107 VSS.n106 0.00250907
R387 VSS.n92 VSS.n91 0.00250907
R388 VSS.n77 VSS.n76 0.00250907
R389 VSS.n74 VSS.n73 0.00247763
R390 VSS.t21 VSS.n74 0.00247763
R391 VSS.n88 VSS.n87 0.00247763
R392 VSS.t27 VSS.n88 0.00247763
R393 VSS.n103 VSS.n102 0.00247763
R394 VSS.t8 VSS.n103 0.00247763
R395 VSS.n118 VSS.n117 0.00247763
R396 VSS.t19 VSS.n118 0.00247763
R397 VSS.n133 VSS.n132 0.00247763
R398 VSS.t5 VSS.n133 0.00247763
R399 VSS.n153 VSS.n152 0.00247763
R400 VSS.t6 VSS.n153 0.00247763
R401 VSS.n168 VSS.n167 0.00247763
R402 VSS.t11 VSS.n168 0.00247763
R403 VSS.n183 VSS.n182 0.00247763
R404 VSS.t10 VSS.n183 0.00247763
R405 VSS.n218 VSS.n217 0.00247763
R406 VSS.t22 VSS.n218 0.00247763
R407 VSS.n198 VSS.n197 0.00247763
R408 VSS.t4 VSS.n198 0.00247763
R409 VSS.n264 VSS.n263 0.00247763
R410 VSS.t2 VSS.n264 0.00247763
R411 VSS.n279 VSS.n278 0.00247763
R412 VSS.t16 VSS.n279 0.00247763
R413 VSS.n294 VSS.n293 0.00247763
R414 VSS.t0 VSS.n294 0.00247763
R415 VSS.n296 VSS.t0 0.00247763
R416 VSS.n281 VSS.t16 0.00247763
R417 VSS.n266 VSS.t2 0.00247763
R418 VSS.n245 VSS.t25 0.00247763
R419 VSS.n220 VSS.t22 0.00247763
R420 VSS.n200 VSS.t4 0.00247763
R421 VSS.n185 VSS.t10 0.00247763
R422 VSS.n170 VSS.t11 0.00247763
R423 VSS.n155 VSS.t6 0.00247763
R424 VSS.n135 VSS.t5 0.00247763
R425 VSS.n120 VSS.t19 0.00247763
R426 VSS.n105 VSS.t8 0.00247763
R427 VSS.n90 VSS.t27 0.00247763
R428 VSS.n75 VSS.t21 0.00247763
R429 VSS.n243 VSS.n242 0.00247763
R430 VSS.t25 VSS.n243 0.00247763
R431 VSS.n310 VSS.n309 0.00247763
R432 VSS.t14 VSS.n310 0.00247763
R433 VSS.n325 VSS.n324 0.00247763
R434 VSS.t23 VSS.n325 0.00247763
R435 VSS.n342 VSS.n341 0.00247763
R436 VSS.t7 VSS.n342 0.00247763
R437 VSS.n357 VSS.n356 0.00247763
R438 VSS.t9 VSS.n357 0.00247763
R439 VSS.n372 VSS.n371 0.00247763
R440 VSS.t24 VSS.n372 0.00247763
R441 VSS.n387 VSS.n386 0.00247763
R442 VSS.t3 VSS.n387 0.00247763
R443 VSS.n402 VSS.n401 0.00247763
R444 VSS.t1 VSS.n402 0.00247763
R445 VSS.n413 VSS.n412 0.00247763
R446 VSS.n412 VSS.t12 0.00247763
R447 VSS.t12 VSS.n411 0.00247763
R448 VSS.n404 VSS.t1 0.00247763
R449 VSS.n389 VSS.t3 0.00247763
R450 VSS.n374 VSS.t24 0.00247763
R451 VSS.n359 VSS.t9 0.00247763
R452 VSS.n344 VSS.t7 0.00247763
R453 VSS.n327 VSS.t23 0.00247763
R454 VSS.n312 VSS.t14 0.00247763
R455 VSS.n411 VSS.n410 0.00247763
R456 VSS.n405 VSS.n404 0.00247763
R457 VSS.n390 VSS.n389 0.00247763
R458 VSS.n375 VSS.n374 0.00247763
R459 VSS.n360 VSS.n359 0.00247763
R460 VSS.n345 VSS.n344 0.00247763
R461 VSS.n328 VSS.n327 0.00247763
R462 VSS.n313 VSS.n312 0.00247763
R463 VSS.n297 VSS.n296 0.00247763
R464 VSS.n282 VSS.n281 0.00247763
R465 VSS.n267 VSS.n266 0.00247763
R466 VSS.n246 VSS.n245 0.00247763
R467 VSS.n221 VSS.n220 0.00247763
R468 VSS.n201 VSS.n200 0.00247763
R469 VSS.n186 VSS.n185 0.00247763
R470 VSS.n171 VSS.n170 0.00247763
R471 VSS.n156 VSS.n155 0.00247763
R472 VSS.n136 VSS.n135 0.00247763
R473 VSS.n121 VSS.n120 0.00247763
R474 VSS.n106 VSS.n105 0.00247763
R475 VSS.n91 VSS.n90 0.00247763
R476 VSS.n76 VSS.n75 0.00247763
R477 VSS.n23 VSS.n21 0.00204594
R478 VSS.n251 VSS.n250 0.00188889
R479 VSS.n445 VSS.n444 0.00172549
R480 VSS.n430 VSS.n429 0.00125043
R481 VSS.n455 VSS.n441 0.00114322
R482 VSS.n429 VSS.n426 0.00103602
R483 VSS.n431 VSS.n425 0.00100003
R484 VSS.n439 VSS.n438 0.000966399
R485 VSS.n438 VSS.n437 0.000959101
R486 VSS.n437 VSS.n436 0.000959101
R487 VSS.n57 VSS.n56 0.000864406
R488 VSS.n62 VSS.n61 0.000864406
R489 VSS.n58 VSS.n57 0.000858717
R490 VSS.n59 VSS.n58 0.000858717
R491 VSS.n61 VSS.n60 0.000858717
R492 VSS.n60 VSS.n59 0.000858717
R493 VSS.n20 VSS.n19 0.000858717
R494 VSS.n19 VSS.n18 0.000858717
R495 VSS.n17 VSS.n16 0.000858717
R496 VSS.n18 VSS.n17 0.000858717
R497 VSS.n439 VSS.n433 0.000714408
R498 VSS.n433 VSS.n431 0.000607204
R499 VSS.n419 VSS.n418 0.000567786
R500 VSS.n42 VSS.n41 0.000557678
R501 VSS.n48 VSS.n47 0.000538452
R502 VSS.n2 VSS.n1 0.000537082
R503 VSS.n66 VSS.n65 0.000526656
R504 VSS.n421 VSS.n420 0.000525991
R505 VSS.n8 VSS.n7 0.000524722
R506 VSS.n446 VSS.n445 0.000523819
R507 VSS.n451 VSS.n450 0.000523819
R508 VSS.n455 VSS.n454 0.000523819
R509 VSS.n454 VSS.n453 0.000523446
R510 VSS.n453 VSS.t17 0.000523446
R511 VSS.n447 VSS.n446 0.000523446
R512 VSS.t17 VSS.n447 0.000523446
R513 VSS.n452 VSS.n451 0.000523446
R514 VSS.t17 VSS.n452 0.000523446
R515 VSS.n25 VSS.n24 0.000517138
R516 VSS.n433 VSS.n432 0.00050212
R517 VSS.n21 VSS.n20 0.00050117
R518 VSS.n16 VSS.n15 0.00050117
R519 VSS.n50 VSS.n49 0.000500552
R520 VSS.n64 VSS.n63 0.000500539
R521 VSS.n10 VSS.n9 0.000500355
R522 VSS.n23 VSS.n22 0.000500347
R523 VSS.n253 VSS.n252 0.000500199
R524 VSS.n261 VSS.n260 0.000500107
R525 VSS.n449 VSS.n448 0.000500053
R526 VSS.n444 VSS.n443 0.000500023
R527 a_n2331_n1103.n14 a_n2331_n1103.t21 182.77
R528 a_n2331_n1103.n15 a_n2331_n1103.t8 182.77
R529 a_n2331_n1103.n16 a_n2331_n1103.t12 182.77
R530 a_n2331_n1103.n17 a_n2331_n1103.t22 182.77
R531 a_n2331_n1103.n18 a_n2331_n1103.t5 182.77
R532 a_n2331_n1103.n19 a_n2331_n1103.t18 182.77
R533 a_n2331_n1103.n20 a_n2331_n1103.t9 182.77
R534 a_n2331_n1103.n21 a_n2331_n1103.t7 182.77
R535 a_n2331_n1103.n22 a_n2331_n1103.t15 182.77
R536 a_n2331_n1103.n2 a_n2331_n1103.t0 182.77
R537 a_n2331_n1103.n4 a_n2331_n1103.t4 182.77
R538 a_n2331_n1103.n5 a_n2331_n1103.t14 182.77
R539 a_n2331_n1103.n6 a_n2331_n1103.t17 182.77
R540 a_n2331_n1103.n7 a_n2331_n1103.t6 182.77
R541 a_n2331_n1103.n8 a_n2331_n1103.t16 182.77
R542 a_n2331_n1103.n9 a_n2331_n1103.t19 182.77
R543 a_n2331_n1103.n10 a_n2331_n1103.t10 182.77
R544 a_n2331_n1103.n11 a_n2331_n1103.t13 182.77
R545 a_n2331_n1103.n12 a_n2331_n1103.t23 182.77
R546 a_n2331_n1103.n13 a_n2331_n1103.t11 90.7933
R547 a_n2331_n1103.n3 a_n2331_n1103.t20 90.7875
R548 a_n2331_n1103.n0 a_n2331_n1103.t2 42.4202
R549 a_n2331_n1103.n0 a_n2331_n1103.t1 4.35105
R550 a_n2331_n1103.t3 a_n2331_n1103.n0 2.70045
R551 a_n2331_n1103.n4 a_n2331_n1103.n3 2.03273
R552 a_n2331_n1103.n14 a_n2331_n1103.n13 2.02124
R553 a_n2331_n1103.n0 a_n2331_n1103.n2 1.1178
R554 a_n2331_n1103.n1 a_n2331_n1103.n40 0.835222
R555 a_n2331_n1103.n40 a_n2331_n1103.n39 0.835222
R556 a_n2331_n1103.n39 a_n2331_n1103.n38 0.835222
R557 a_n2331_n1103.n38 a_n2331_n1103.n37 0.835222
R558 a_n2331_n1103.n37 a_n2331_n1103.n36 0.835222
R559 a_n2331_n1103.n36 a_n2331_n1103.n35 0.835222
R560 a_n2331_n1103.n35 a_n2331_n1103.n34 0.835222
R561 a_n2331_n1103.n34 a_n2331_n1103.n33 0.835222
R562 a_n2331_n1103.n33 a_n2331_n1103.n32 0.835222
R563 a_n2331_n1103.n15 a_n2331_n1103.n14 0.835222
R564 a_n2331_n1103.n16 a_n2331_n1103.n15 0.835222
R565 a_n2331_n1103.n17 a_n2331_n1103.n16 0.835222
R566 a_n2331_n1103.n18 a_n2331_n1103.n17 0.835222
R567 a_n2331_n1103.n19 a_n2331_n1103.n18 0.835222
R568 a_n2331_n1103.n20 a_n2331_n1103.n19 0.835222
R569 a_n2331_n1103.n21 a_n2331_n1103.n20 0.835222
R570 a_n2331_n1103.n22 a_n2331_n1103.n21 0.835222
R571 a_n2331_n1103.n2 a_n2331_n1103.n22 0.835222
R572 a_n2331_n1103.n12 a_n2331_n1103.n11 0.835222
R573 a_n2331_n1103.n11 a_n2331_n1103.n10 0.835222
R574 a_n2331_n1103.n10 a_n2331_n1103.n9 0.835222
R575 a_n2331_n1103.n9 a_n2331_n1103.n8 0.835222
R576 a_n2331_n1103.n8 a_n2331_n1103.n7 0.835222
R577 a_n2331_n1103.n7 a_n2331_n1103.n6 0.835222
R578 a_n2331_n1103.n6 a_n2331_n1103.n5 0.835222
R579 a_n2331_n1103.n5 a_n2331_n1103.n4 0.835222
R580 a_n2331_n1103.n24 a_n2331_n1103.n23 0.835222
R581 a_n2331_n1103.n25 a_n2331_n1103.n24 0.835222
R582 a_n2331_n1103.n26 a_n2331_n1103.n25 0.835222
R583 a_n2331_n1103.n27 a_n2331_n1103.n26 0.835222
R584 a_n2331_n1103.n28 a_n2331_n1103.n27 0.835222
R585 a_n2331_n1103.n29 a_n2331_n1103.n28 0.835222
R586 a_n2331_n1103.n30 a_n2331_n1103.n29 0.835222
R587 a_n2331_n1103.n31 a_n2331_n1103.n30 0.835222
R588 a_n2331_n1103.n2 a_n2331_n1103.n12 0.786611
R589 a_n2331_n1103.n1 a_n2331_n1103.n31 0.786611
R590 a_n2331_n1103.n0 a_n2331_n1103.n1 0.750184
R591 a_n2211_n1015.n18 a_n2211_n1015.t24 473.437
R592 a_n2211_n1015.n12 a_n2211_n1015.t25 473.332
R593 a_n2211_n1015.n1 a_n2211_n1015.t22 473.329
R594 a_n2211_n1015.n11 a_n2211_n1015.t20 140.444
R595 a_n2211_n1015.n11 a_n2211_n1015.t21 41.6504
R596 a_n2211_n1015.n2 a_n2211_n1015.t12 5.95597
R597 a_n2211_n1015.n27 a_n2211_n1015.t3 5.95597
R598 a_n2211_n1015.n2 a_n2211_n1015.t2 5.32159
R599 a_n2211_n1015.n3 a_n2211_n1015.t15 5.32159
R600 a_n2211_n1015.n4 a_n2211_n1015.t11 5.32159
R601 a_n2211_n1015.n5 a_n2211_n1015.t1 5.32159
R602 a_n2211_n1015.n6 a_n2211_n1015.t18 5.32159
R603 a_n2211_n1015.n7 a_n2211_n1015.t5 5.32159
R604 a_n2211_n1015.n8 a_n2211_n1015.t14 5.32159
R605 a_n2211_n1015.n9 a_n2211_n1015.t16 5.32159
R606 a_n2211_n1015.n10 a_n2211_n1015.t8 5.32159
R607 a_n2211_n1015.n0 a_n2211_n1015.t0 5.32159
R608 a_n2211_n1015.n1 a_n2211_n1015.t10 5.32159
R609 a_n2211_n1015.n21 a_n2211_n1015.t13 5.32159
R610 a_n2211_n1015.n22 a_n2211_n1015.t4 5.32159
R611 a_n2211_n1015.n23 a_n2211_n1015.t7 5.32159
R612 a_n2211_n1015.n24 a_n2211_n1015.t17 5.32159
R613 a_n2211_n1015.n25 a_n2211_n1015.t6 5.32159
R614 a_n2211_n1015.n26 a_n2211_n1015.t9 5.32159
R615 a_n2211_n1015.t19 a_n2211_n1015.n27 5.32059
R616 a_n2211_n1015.n17 a_n2211_n1015.n16 2.75606
R617 a_n2211_n1015.n20 a_n2211_n1015.n17 2.75328
R618 a_n2211_n1015.n17 a_n2211_n1015.t23 1.50409
R619 a_n2211_n1015.n12 a_n2211_n1015.n11 1.23545
R620 a_n2211_n1015.n0 a_n2211_n1015.n10 1.02772
R621 a_n2211_n1015.n10 a_n2211_n1015.n9 0.634875
R622 a_n2211_n1015.n9 a_n2211_n1015.n8 0.634875
R623 a_n2211_n1015.n8 a_n2211_n1015.n7 0.634875
R624 a_n2211_n1015.n7 a_n2211_n1015.n6 0.634875
R625 a_n2211_n1015.n6 a_n2211_n1015.n5 0.634875
R626 a_n2211_n1015.n5 a_n2211_n1015.n4 0.634875
R627 a_n2211_n1015.n4 a_n2211_n1015.n3 0.634875
R628 a_n2211_n1015.n3 a_n2211_n1015.n2 0.634875
R629 a_n2211_n1015.n27 a_n2211_n1015.n26 0.634875
R630 a_n2211_n1015.n26 a_n2211_n1015.n25 0.634875
R631 a_n2211_n1015.n25 a_n2211_n1015.n24 0.634875
R632 a_n2211_n1015.n24 a_n2211_n1015.n23 0.634875
R633 a_n2211_n1015.n23 a_n2211_n1015.n22 0.634875
R634 a_n2211_n1015.n22 a_n2211_n1015.n21 0.634875
R635 a_n2211_n1015.n1 a_n2211_n1015.n14 0.376529
R636 a_n2211_n1015.n19 a_n2211_n1015.n18 0.271346
R637 a_n2211_n1015.n21 a_n2211_n1015.n1 0.260122
R638 a_n2211_n1015.n14 a_n2211_n1015.n13 0.253053
R639 a_n2211_n1015.n1 a_n2211_n1015.n0 0.12461
R640 a_n2211_n1015.n13 a_n2211_n1015.n12 0.124538
R641 a_n2211_n1015.n20 a_n2211_n1015.n19 0.119076
R642 a_n2211_n1015.n16 a_n2211_n1015.n15 0.113872
R643 a_n2211_n1015.n1 a_n2211_n1015.n20 0.10111
R644 VDD.n37 VDD.n34 437.647
R645 VDD.n52 VDD.n49 430.589
R646 VDD.n4 VDD.n1 430.589
R647 VDD.n17 VDD.n14 420
R648 VDD.n48 VDD.t4 54.472
R649 VDD.n48 VDD.t0 54.472
R650 VDD.n12 VDD.t2 54.2478
R651 VDD.n11 VDD.n8 54.1098
R652 VDD.n45 VDD.n42 54.1091
R653 VDD.n36 VDD.n35 46.6829
R654 VDD.n51 VDD.n50 45.9299
R655 VDD.n3 VDD.n2 45.9299
R656 VDD.n16 VDD.n15 44.8005
R657 VDD.n23 VDD.n22 8.85536
R658 VDD.n24 VDD.n23 4.58799
R659 VDD.n18 VDD.n13 3.5871
R660 VDD.n58 VDD.n26 2.83443
R661 VDD.n58 VDD.n57 2.80943
R662 VDD.n25 VDD.t3 1.50409
R663 VDD.n29 VDD.t5 1.50409
R664 VDD.n29 VDD.t1 1.50409
R665 VDD.n29 VDD.n28 0.800961
R666 VDD.n23 VDD.n21 0.738962
R667 VDD.n18 VDD.n12 0.224662
R668 VDD.n17 VDD.n16 0.107375
R669 VDD.n18 VDD.n17 0.107375
R670 VDD.n53 VDD.n52 0.100461
R671 VDD.n19 VDD.n4 0.100461
R672 VDD.n52 VDD.n51 0.0999624
R673 VDD.n4 VDD.n3 0.0999624
R674 VDD.n40 VDD.n37 0.0960166
R675 VDD.n37 VDD.n36 0.095518
R676 VDD VDD.n58 0.0676185
R677 VDD.n26 VDD.n25 0.0258165
R678 VDD.n25 VDD.n24 0.0183679
R679 VDD.n11 VDD.n10 0.0154506
R680 VDD.n45 VDD.n44 0.015449
R681 VDD.n10 VDD.n9 0.0150463
R682 VDD.n33 VDD.n32 0.0150463
R683 VDD.t4 VDD.n33 0.0150463
R684 VDD.n47 VDD.n46 0.0150463
R685 VDD.t0 VDD.n47 0.0150463
R686 VDD.n44 VDD.n43 0.0150463
R687 VDD.t4 VDD.n31 0.0150463
R688 VDD.n31 VDD.n30 0.0150463
R689 VDD.t2 VDD.n6 0.0150463
R690 VDD.n6 VDD.n5 0.0150463
R691 VDD.n57 VDD.n56 0.0138929
R692 VDD.n26 VDD.n0 0.0108144
R693 VDD.n40 VDD.n39 0.00317113
R694 VDD.n20 VDD.n19 0.00317113
R695 VDD.n39 VDD.n38 0.00267116
R696 VDD.n21 VDD.n20 0.00267116
R697 VDD.n8 VDD.n7 0.00158558
R698 VDD.n42 VDD.n41 0.00158558
R699 VDD.n56 VDD.n29 0.00139286
R700 VDD.t2 VDD.n11 0.00134143
R701 VDD.n54 VDD.n53 0.00111635
R702 VDD.t0 VDD.n45 0.0010973
R703 VDD.n19 VDD.n18 0.00100003
R704 VDD.n48 VDD.n40 0.00100003
R705 VDD.n53 VDD.n48 0.001
R706 VDD.n57 VDD.n27 0.001
R707 VDD.n55 VDD.n54 0.00061635
R708 VDD.n56 VDD.n55 0.000616347
R709 VOUT.n0 VOUT.t1 182.794
R710 VOUT.n6 VOUT.t0 6.11598
R711 VOUT.n2 VOUT.t2 4.35136
R712 VOUT.n3 VOUT.n2 0.807781
R713 VOUT.n6 VOUT.n5 0.749453
R714 VOUT VOUT.n6 0.168769
R715 VOUT.n4 VOUT.n3 0.063
R716 VOUT.n1 VOUT.n0 0.00758218
R717 VOUT.n5 VOUT.n1 0.00620837
R718 VOUT.n5 VOUT.n4 0.00100612
C0 VOUT VDD 2.97f
.ends

