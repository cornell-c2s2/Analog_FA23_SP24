magic
tech sky130A
magscale 1 2
timestamp 1708718597
<< checkpaint >>
rect 38349 752 42183 805
rect 38349 699 43444 752
rect 38349 646 44705 699
rect 38349 -12135 45966 646
rect 39610 -12188 45966 -12135
rect 40871 -12241 45966 -12188
rect 42132 -12294 45966 -12241
<< error_s >>
rect 3822 1897 3857 1931
rect 3823 1878 3857 1897
rect 3842 583 3857 1878
rect 3876 1844 3911 1878
rect 5209 1844 5244 1878
rect 3876 583 3910 1844
rect 5210 1825 5244 1844
rect 6614 1825 6667 1826
rect 3876 549 3891 583
rect 5229 530 5244 1825
rect 5263 1791 5298 1825
rect 6596 1791 6667 1825
rect 5263 530 5297 1791
rect 6597 1790 6667 1791
rect 6614 1756 6685 1790
rect 10195 1756 10230 1790
rect 5263 496 5278 530
rect 6614 477 6684 1756
rect 10196 1737 10230 1756
rect 6614 441 6667 477
rect 10215 424 10230 1737
rect 10249 1703 10284 1737
rect 13794 1703 13829 1737
rect 10249 424 10283 1703
rect 13795 1684 13829 1703
rect 10249 390 10264 424
rect 13814 371 13829 1684
rect 13848 1650 13883 1684
rect 20395 1650 20430 1667
rect 13848 371 13882 1650
rect 20396 1649 20430 1650
rect 20396 1613 20466 1649
rect 20413 1579 20484 1613
rect 13848 337 13863 371
rect 20413 318 20483 1579
rect 20413 282 20466 318
rect 40852 -525 40887 -491
rect 40853 -544 40887 -525
rect 39894 -593 39952 -587
rect 40090 -593 40148 -587
rect 40286 -593 40344 -587
rect 40482 -593 40540 -587
rect 40678 -593 40736 -587
rect 39894 -627 39906 -593
rect 40090 -627 40102 -593
rect 40286 -627 40298 -593
rect 40482 -627 40494 -593
rect 40678 -627 40690 -593
rect 39894 -633 39952 -627
rect 40090 -633 40148 -627
rect 40286 -633 40344 -627
rect 40482 -633 40540 -627
rect 40678 -633 40736 -627
rect 28770 -9119 28804 -9101
rect 28770 -9155 28840 -9119
rect 28787 -9189 28858 -9155
rect 30598 -9189 30633 -9155
rect 28787 -10468 28857 -9189
rect 30599 -9208 30633 -9189
rect 28787 -10504 28840 -10468
rect 30618 -10521 30633 -9208
rect 30652 -9242 30687 -9208
rect 32427 -9242 32462 -9225
rect 30652 -10521 30686 -9242
rect 32428 -9243 32462 -9242
rect 32428 -9279 32498 -9243
rect 32445 -9313 32516 -9279
rect 30652 -10555 30667 -10521
rect 32445 -10574 32515 -9313
rect 34257 -10082 34291 -10028
rect 32445 -10610 32498 -10574
rect 34276 -10627 34291 -10082
rect 34310 -10116 34345 -10082
rect 34310 -10627 34344 -10116
rect 34310 -10661 34325 -10627
rect 35589 -10680 35604 -10082
rect 35623 -10680 35657 -10028
rect 35623 -10714 35638 -10680
rect 36186 -10733 36201 -9885
rect 36220 -10733 36254 -9831
rect 39796 -10703 39854 -10697
rect 39992 -10703 40050 -10697
rect 40188 -10703 40246 -10697
rect 40384 -10703 40442 -10697
rect 40580 -10703 40638 -10697
rect 36220 -10767 36235 -10733
rect 39796 -10737 39808 -10703
rect 39992 -10737 40004 -10703
rect 40188 -10737 40200 -10703
rect 40384 -10737 40396 -10703
rect 40580 -10737 40592 -10703
rect 39796 -10743 39854 -10737
rect 39992 -10743 40050 -10737
rect 40188 -10743 40246 -10737
rect 40384 -10743 40442 -10737
rect 40580 -10743 40638 -10737
rect 40872 -10839 40887 -544
rect 40906 -578 40941 -544
rect 42113 -578 42148 -544
rect 40906 -10839 40940 -578
rect 42114 -597 42148 -578
rect 41155 -646 41213 -640
rect 41351 -646 41409 -640
rect 41547 -646 41605 -640
rect 41743 -646 41801 -640
rect 41939 -646 41997 -640
rect 41155 -680 41167 -646
rect 41351 -680 41363 -646
rect 41547 -680 41559 -646
rect 41743 -680 41755 -646
rect 41939 -680 41951 -646
rect 41155 -686 41213 -680
rect 41351 -686 41409 -680
rect 41547 -686 41605 -680
rect 41743 -686 41801 -680
rect 41939 -686 41997 -680
rect 41057 -10756 41115 -10750
rect 41253 -10756 41311 -10750
rect 41449 -10756 41507 -10750
rect 41645 -10756 41703 -10750
rect 41841 -10756 41899 -10750
rect 41057 -10790 41069 -10756
rect 41253 -10790 41265 -10756
rect 41449 -10790 41461 -10756
rect 41645 -10790 41657 -10756
rect 41841 -10790 41853 -10756
rect 41057 -10796 41115 -10790
rect 41253 -10796 41311 -10790
rect 41449 -10796 41507 -10790
rect 41645 -10796 41703 -10790
rect 41841 -10796 41899 -10790
rect 40906 -10873 40921 -10839
rect 42133 -10892 42148 -597
rect 42167 -631 42202 -597
rect 42167 -10892 42201 -631
rect 42416 -699 42474 -693
rect 42612 -699 42670 -693
rect 42808 -699 42866 -693
rect 43004 -699 43062 -693
rect 43200 -699 43258 -693
rect 42416 -733 42428 -699
rect 42612 -733 42624 -699
rect 42808 -733 42820 -699
rect 43004 -733 43016 -699
rect 43200 -733 43212 -699
rect 42416 -739 42474 -733
rect 42612 -739 42670 -733
rect 42808 -739 42866 -733
rect 43004 -739 43062 -733
rect 43200 -739 43258 -733
rect 42318 -10809 42376 -10803
rect 42514 -10809 42572 -10803
rect 42710 -10809 42768 -10803
rect 42906 -10809 42964 -10803
rect 43102 -10809 43160 -10803
rect 42318 -10843 42330 -10809
rect 42514 -10843 42526 -10809
rect 42710 -10843 42722 -10809
rect 42906 -10843 42918 -10809
rect 43102 -10843 43114 -10809
rect 42318 -10849 42376 -10843
rect 42514 -10849 42572 -10843
rect 42710 -10849 42768 -10843
rect 42906 -10849 42964 -10843
rect 43102 -10849 43160 -10843
rect 42167 -10926 42182 -10892
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
rect 0 -1600 200 -1400
use sky130_fd_pr__res_generic_m3_7P7WHS  R16
timestamp 0
transform 1 0 38662 0 1 -3215
box -1000 -7607 1000 7607
use sky130_fd_pr__cap_mim_m3_1_RJVX7Z  XC2
timestamp 0
transform 1 0 25629 0 1 -3411
box -1786 -7040 1786 7040
use sky130_fd_pr__nfet_01v8_X9T245  XM28
timestamp 0
transform 1 0 1920 0 1 1257
box -1973 -710 1973 710
use sky130_fd_pr__nfet_01v8_F7BW33  XM29
timestamp 0
transform 1 0 4560 0 1 1204
box -720 -710 720 710
use sky130_fd_pr__nfet_01v8_F7BW33  XM30
timestamp 0
transform 1 0 5947 0 1 1151
box -720 -710 720 710
use sky130_fd_pr__pfet_01v8_GCT3F7  XM31
timestamp 0
transform 1 0 8440 0 1 1107
box -1826 -719 1826 719
use sky130_fd_pr__pfet_01v8_GCT3F7  XM32
timestamp 0
transform 1 0 12039 0 1 1054
box -1826 -719 1826 719
use sky130_fd_pr__pfet_01v8_ED7GUS  XM38
timestamp 0
transform 1 0 17139 0 1 1001
box -3327 -719 3327 719
use sky130_fd_pr__nfet_01v8_6JG44H  XM39
timestamp 0
transform 1 0 22128 0 1 939
box -1715 -710 1715 710
use sky130_fd_pr__pfet_01v8_3H5TVM  XM40
timestamp 0
transform 1 0 29728 0 1 -9838
box -941 -719 941 719
use sky130_fd_pr__pfet_01v8_3H5TVM  XM41
timestamp 0
transform 1 0 31557 0 1 -9891
box -941 -719 941 719
use sky130_fd_pr__nfet_01v8_UFMA4B  XM42
timestamp 0
transform 1 0 33386 0 1 -9953
box -941 -710 941 710
use sky130_fd_pr__nfet_01v8_UR5WPG  XM43
timestamp 0
transform 1 0 34957 0 1 -10381
box -683 -335 683 335
use sky130_fd_pr__nfet_01v8_G6BLWB  XM44
timestamp 0
transform 1 0 35912 0 1 -10309
box -325 -460 325 460
use sky130_fd_pr__nfet_01v8_8WJ4K3  XM57
timestamp 0
transform 1 0 40266 0 1 -5665
box -657 -5210 657 5210
use sky130_fd_pr__nfet_01v8_8WJ4K3  XM58
timestamp 0
transform 1 0 41527 0 1 -5718
box -657 -5210 657 5210
use sky130_fd_pr__nfet_01v8_8WJ4K3  XM59
timestamp 0
transform 1 0 42788 0 1 -5771
box -657 -5210 657 5210
use sky130_fd_pr__nfet_01v8_8WJ4K3  XM60
timestamp 0
transform 1 0 44049 0 1 -5824
box -657 -5210 657 5210
use sky130_fd_pr__res_xhigh_po_5p73_ETCMCS  XR6
timestamp 0
transform 1 0 28101 0 1 -8922
box -739 -1582 739 1582
use sky130_fd_pr__res_xhigh_po_5p73_5TXYRS  XR8
timestamp 0
transform 1 0 36923 0 1 -3340
box -739 -7482 739 7482
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 VDD
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 VP
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 VN
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 OUT
port 3 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 256 0 0 0 VSS
port 4 nsew
<< end >>
