magic
tech sky130A
magscale 1 2
timestamp 1711217682
<< nwell >>
rect 450 -220 2250 180
rect 450 -230 2790 -220
rect 450 -540 2250 -230
rect 2780 -540 2790 -230
rect 450 -560 2790 -540
rect 450 -1510 3240 -1180
rect 450 -1870 2590 -1510
rect 450 -2830 3600 -2500
<< metal1 >>
rect -1400 400 -1200 600
rect 480 381 2220 491
rect -1400 0 -1200 200
rect -1400 -400 -1200 -200
rect 480 -209 2210 -59
rect 480 -319 2760 -209
rect 3800 -400 4000 -200
rect -1400 -800 -1200 -600
rect 480 -980 2760 -760
rect 3800 -800 4000 -600
rect -1400 -1200 -1200 -1000
rect 3800 -1200 4000 -1000
rect -1400 -1600 -1200 -1400
rect 480 -1530 3210 -1410
rect 480 -1640 2600 -1530
rect 3800 -1600 4000 -1400
rect -1400 -2000 -1200 -1800
rect 3800 -2000 4000 -1800
rect 480 -2200 2490 -2080
rect -1400 -2400 -1200 -2200
rect 480 -2300 3560 -2200
rect -1400 -2800 -1200 -2600
rect 480 -2850 3570 -2730
use sky130_fd_sc_hd__or4_1  x1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1711211407
transform 1 0 488 0 1 -811
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  x2
timestamp 1711211407
transform 1 0 1118 0 1 -811
box -38 -48 590 592
use sky130_fd_sc_hd__inv_1  x3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 848 0 -1 433
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  x4 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 1748 0 1 -811
box -38 -48 498 592
use sky130_fd_sc_hd__inv_1  x5
timestamp 1701704242
transform 1 0 1568 0 -1 433
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  x6
timestamp 1701704242
transform 1 0 1208 0 -1 433
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  x7
timestamp 1701704242
transform 1 0 1928 0 -1 433
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  x8 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 2288 0 1 -811
box -38 -48 498 592
use sky130_fd_sc_hd__inv_1  x9
timestamp 1701704242
transform 1 0 488 0 -1 433
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  x10
timestamp 1701704242
transform 1 0 488 0 -1 -928
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  x11
timestamp 1701704242
transform 1 0 1028 0 -1 -928
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  x12
timestamp 1701704242
transform 1 0 1568 0 -1 -928
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  x13
timestamp 1701704242
transform 1 0 2108 0 -1 -928
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  x14
timestamp 1711211407
transform 1 0 2648 0 -1 -928
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  x15 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 488 0 1 -2132
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  x16
timestamp 1701704242
transform 1 0 1208 0 1 -2132
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  x17
timestamp 1711211407
transform 1 0 1928 0 1 -2132
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  x18
timestamp 1701704242
transform 1 0 488 0 -1 -2248
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  x19
timestamp 1701704242
transform 1 0 1208 0 -1 -2248
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  x20 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 1928 0 -1 -2248
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  x21
timestamp 1701704242
transform 1 0 2468 0 -1 -2248
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  x22
timestamp 1711211407
transform -1 0 3560 0 -1 -2248
box -38 -48 590 592
<< labels >>
flabel metal1 3800 -2000 4000 -1800 0 FreeSans 256 0 0 0 A0
port 12 nsew
flabel metal1 3800 -1600 4000 -1400 0 FreeSans 256 0 0 0 A1
port 11 nsew
flabel metal1 3800 -1200 4000 -1000 0 FreeSans 256 0 0 0 A2
port 10 nsew
flabel metal1 3800 -400 4000 -200 0 FreeSans 256 0 0 0 EO
port 8 nsew
flabel metal1 3800 -800 4000 -600 0 FreeSans 256 0 0 0 GS
port 9 nsew
flabel metal1 -1400 -2800 -1200 -2600 0 FreeSans 256 0 0 0 I7
port 6 nsew
flabel metal1 -1400 -2400 -1200 -2200 0 FreeSans 256 0 0 0 I6
port 5 nsew
flabel metal1 -1400 -2000 -1200 -1800 0 FreeSans 256 0 0 0 I5
port 1 nsew
flabel metal1 -1400 -1600 -1200 -1400 0 FreeSans 256 0 0 0 I4
port 7 nsew
flabel metal1 -1400 -1200 -1200 -1000 0 FreeSans 256 0 0 0 I3
port 2 nsew
flabel metal1 -1400 -800 -1200 -600 0 FreeSans 256 0 0 0 I2
port 4 nsew
flabel metal1 -1400 -400 -1200 -200 0 FreeSans 256 0 0 0 I1
port 0 nsew
flabel metal1 -1400 0 -1200 200 0 FreeSans 256 0 0 0 I0
port 3 nsew
flabel metal1 -1400 400 -1200 600 0 FreeSans 256 0 0 0 EI
port 13 nsew
<< end >>
