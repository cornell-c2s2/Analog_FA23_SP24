magic
tech sky130A
magscale 1 2
timestamp 1713148681
<< viali >>
rect 1620 100 1660 140
rect 2060 100 2100 140
rect 2626 92 2666 132
rect 3026 92 3066 132
rect 3426 94 3466 133
rect 3826 92 3866 132
rect 4226 92 4266 132
rect 5026 92 5066 132
rect 5426 92 5466 132
rect 5826 92 5866 132
rect 6226 92 6266 132
rect 6585 90 6625 136
rect 1620 -2750 1680 -2700
rect 1940 -2750 2000 -2700
rect 3533 -2744 3583 -2694
rect 3933 -2744 3983 -2694
rect 4333 -2744 4383 -2694
rect 4733 -2744 4783 -2694
rect 5133 -2744 5183 -2694
rect 5533 -2744 5583 -2694
<< metal1 >>
rect 1600 140 1640 200
rect 1600 100 1620 140
rect 1700 100 1830 200
rect 1890 100 2020 200
rect 2080 140 6800 200
rect 2100 136 6800 140
rect 2100 133 6585 136
rect 2100 132 3426 133
rect 2100 100 2626 132
rect 1600 80 1680 100
rect 2040 80 2120 100
rect 2614 92 2626 100
rect 2666 100 3026 132
rect 2666 92 2678 100
rect 2614 86 2678 92
rect 3014 92 3026 100
rect 3066 100 3426 132
rect 3066 92 3078 100
rect 3014 86 3078 92
rect 3409 94 3426 100
rect 3466 132 6585 133
rect 3466 100 3826 132
rect 3466 94 3478 100
rect 3409 89 3478 94
rect 3814 92 3826 100
rect 3866 100 4226 132
rect 3866 92 3878 100
rect 3409 87 3477 89
rect 3814 86 3878 92
rect 4214 92 4226 100
rect 4266 100 5026 132
rect 4266 92 4278 100
rect 4214 86 4278 92
rect 5014 92 5026 100
rect 5066 100 5426 132
rect 5066 92 5078 100
rect 5014 86 5078 92
rect 5414 92 5426 100
rect 5466 100 5826 132
rect 5466 92 5478 100
rect 5414 86 5478 92
rect 5814 92 5826 100
rect 5866 100 6226 132
rect 5866 92 5878 100
rect 5814 86 5878 92
rect 6214 92 6226 100
rect 6266 100 6585 132
rect 6266 92 6278 100
rect 6214 86 6278 92
rect 6569 90 6585 100
rect 6625 100 6800 136
rect 6625 90 6644 100
rect 6569 83 6644 90
rect 1490 -50 1500 50
rect 1600 -50 2116 50
rect 2366 -50 2372 50
rect 2472 -50 4560 50
rect 4660 -50 4670 50
rect 4780 -50 6720 50
rect 6820 -50 6830 50
rect 1630 -400 1640 -300
rect 1700 -400 1710 -300
rect 1820 -400 1830 -300
rect 1890 -400 1900 -300
rect 2010 -400 2020 -300
rect 2080 -400 2090 -300
rect 2720 -394 2730 -294
rect 2790 -394 2800 -294
rect 2920 -394 2930 -294
rect 2990 -394 3000 -294
rect 3110 -394 3120 -294
rect 3180 -394 3190 -294
rect 3300 -394 3310 -294
rect 3370 -394 3380 -294
rect 3490 -394 3500 -294
rect 3560 -394 3570 -294
rect 3680 -394 3690 -294
rect 3750 -394 3760 -294
rect 3880 -394 3890 -294
rect 3950 -394 3960 -294
rect 4070 -394 4080 -294
rect 4140 -394 4150 -294
rect 4260 -394 4270 -294
rect 4330 -394 4340 -294
rect 4450 -394 4460 -294
rect 4520 -394 4530 -294
rect 4870 -400 4880 -300
rect 4940 -400 4950 -300
rect 5070 -400 5080 -300
rect 5140 -400 5150 -300
rect 5260 -400 5270 -300
rect 5330 -400 5340 -300
rect 5450 -400 5460 -300
rect 5520 -400 5530 -300
rect 5640 -400 5650 -300
rect 5710 -400 5720 -300
rect 5830 -400 5840 -300
rect 5900 -400 5910 -300
rect 6030 -400 6040 -300
rect 6100 -400 6110 -300
rect 6220 -400 6230 -300
rect 6290 -400 6300 -300
rect 6410 -400 6420 -300
rect 6480 -400 6490 -300
rect 6600 -400 6610 -300
rect 6670 -400 6680 -300
rect 2630 -900 2640 -800
rect 2700 -900 2710 -800
rect 2820 -900 2830 -800
rect 2890 -900 2900 -800
rect 3010 -900 3020 -800
rect 3080 -900 3090 -800
rect 3200 -900 3210 -800
rect 3270 -900 3280 -800
rect 3400 -900 3410 -800
rect 3470 -900 3480 -800
rect 3590 -900 3600 -800
rect 3660 -900 3670 -800
rect 3780 -900 3790 -800
rect 3850 -900 3860 -800
rect 3970 -900 3980 -800
rect 4040 -900 4050 -800
rect 4160 -900 4170 -800
rect 4230 -900 4240 -800
rect 4350 -900 4360 -800
rect 4420 -900 4430 -800
rect 4780 -900 4790 -800
rect 4850 -900 4860 -800
rect 4970 -900 4980 -800
rect 5040 -900 5050 -800
rect 5160 -900 5170 -800
rect 5230 -900 5240 -800
rect 5350 -900 5360 -800
rect 5420 -900 5430 -800
rect 5550 -900 5560 -800
rect 5620 -900 5630 -800
rect 5740 -900 5750 -800
rect 5810 -900 5820 -800
rect 5930 -900 5940 -800
rect 6000 -900 6010 -800
rect 6120 -900 6130 -800
rect 6190 -900 6200 -800
rect 6310 -900 6320 -800
rect 6380 -900 6390 -800
rect 6500 -900 6510 -800
rect 6570 -900 6580 -800
rect 1720 -1000 1730 -900
rect 1790 -1000 1800 -900
rect 1910 -1000 1920 -900
rect 1980 -1000 1990 -900
rect 1490 -1250 1500 -1150
rect 1600 -1250 2034 -1150
rect 2364 -1250 2370 -1150
rect 2470 -1250 4560 -1150
rect 4660 -1250 4666 -1150
rect 4810 -1250 6720 -1150
rect 6820 -1250 6826 -1150
rect 1494 -1500 1500 -1400
rect 1600 -1500 4540 -1400
rect 4640 -1450 4650 -1400
rect 4640 -1500 4680 -1450
rect 4845 -1500 5765 -1450
rect 5759 -1550 5765 -1500
rect 5865 -1550 5871 -1450
rect 1770 -1800 1780 -1700
rect 1840 -1800 1850 -1700
rect 3670 -1800 3680 -1700
rect 3740 -1800 3750 -1700
rect 3870 -1800 3880 -1700
rect 3940 -1800 3950 -1700
rect 4060 -1800 4070 -1700
rect 4130 -1800 4140 -1700
rect 4250 -1800 4260 -1700
rect 4320 -1800 4330 -1700
rect 4440 -1800 4450 -1700
rect 4510 -1800 4520 -1700
rect 4870 -1800 4880 -1700
rect 4940 -1800 4950 -1700
rect 5070 -1800 5080 -1700
rect 5140 -1800 5150 -1700
rect 5260 -1800 5270 -1700
rect 5330 -1800 5340 -1700
rect 5450 -1800 5460 -1700
rect 5520 -1800 5530 -1700
rect 5640 -1800 5650 -1700
rect 5710 -1800 5720 -1700
rect 1670 -2300 1680 -2200
rect 1740 -2300 1750 -2200
rect 1870 -2300 1880 -2200
rect 1940 -2300 1950 -2200
rect 3570 -2300 3580 -2200
rect 3650 -2300 3660 -2200
rect 3770 -2300 3780 -2200
rect 3840 -2300 3850 -2200
rect 3960 -2300 3970 -2200
rect 4030 -2300 4040 -2200
rect 4150 -2300 4160 -2200
rect 4220 -2300 4230 -2200
rect 4340 -2300 4350 -2200
rect 4420 -2300 4430 -2200
rect 4770 -2300 4780 -2200
rect 4850 -2300 4860 -2200
rect 4970 -2300 4980 -2200
rect 5040 -2300 5050 -2200
rect 5160 -2300 5170 -2200
rect 5230 -2300 5240 -2200
rect 5350 -2300 5360 -2200
rect 5420 -2300 5430 -2200
rect 5540 -2300 5550 -2200
rect 5610 -2300 5620 -2200
rect 1494 -2650 1500 -2550
rect 1600 -2600 1606 -2550
rect 4530 -2600 4540 -2570
rect 1600 -2650 1816 -2600
rect 3600 -2650 4540 -2600
rect 4640 -2650 4650 -2570
rect 5755 -2600 5765 -2570
rect 4860 -2650 5765 -2600
rect 5865 -2650 5875 -2570
rect 1599 -2694 5724 -2680
rect 1599 -2698 3533 -2694
rect 1599 -2700 1680 -2698
rect 1599 -2750 1620 -2700
rect 1740 -2750 1880 -2698
rect 1940 -2700 3533 -2698
rect 2000 -2744 3533 -2700
rect 3583 -2744 3933 -2694
rect 3983 -2744 4333 -2694
rect 4383 -2744 4733 -2694
rect 4783 -2744 5133 -2694
rect 5183 -2744 5533 -2694
rect 5583 -2744 5724 -2694
rect 2000 -2750 5724 -2744
rect 1599 -2780 5724 -2750
<< via1 >>
rect 1640 140 1700 200
rect 1640 100 1660 140
rect 1660 100 1700 140
rect 1830 100 1890 200
rect 2020 140 2080 200
rect 2020 100 2060 140
rect 2060 100 2080 140
rect 1500 -50 1600 50
rect 2372 -50 2472 50
rect 4560 -50 4660 50
rect 6720 -50 6820 50
rect 1640 -400 1700 -300
rect 1830 -400 1890 -300
rect 2020 -400 2080 -300
rect 2730 -394 2790 -294
rect 2930 -394 2990 -294
rect 3120 -394 3180 -294
rect 3310 -394 3370 -294
rect 3500 -394 3560 -294
rect 3690 -394 3750 -294
rect 3890 -394 3950 -294
rect 4080 -394 4140 -294
rect 4270 -394 4330 -294
rect 4460 -394 4520 -294
rect 4880 -400 4940 -300
rect 5080 -400 5140 -300
rect 5270 -400 5330 -300
rect 5460 -400 5520 -300
rect 5650 -400 5710 -300
rect 5840 -400 5900 -300
rect 6040 -400 6100 -300
rect 6230 -400 6290 -300
rect 6420 -400 6480 -300
rect 6610 -400 6670 -300
rect 2640 -900 2700 -800
rect 2830 -900 2890 -800
rect 3020 -900 3080 -800
rect 3210 -900 3270 -800
rect 3410 -900 3470 -800
rect 3600 -900 3660 -800
rect 3790 -900 3850 -800
rect 3980 -900 4040 -800
rect 4170 -900 4230 -800
rect 4360 -900 4420 -800
rect 4790 -900 4850 -800
rect 4980 -900 5040 -800
rect 5170 -900 5230 -800
rect 5360 -900 5420 -800
rect 5560 -900 5620 -800
rect 5750 -900 5810 -800
rect 5940 -900 6000 -800
rect 6130 -900 6190 -800
rect 6320 -900 6380 -800
rect 6510 -900 6570 -800
rect 1730 -1000 1790 -900
rect 1920 -1000 1980 -900
rect 1500 -1250 1600 -1150
rect 2370 -1250 2470 -1150
rect 4560 -1250 4660 -1150
rect 6720 -1250 6820 -1150
rect 1500 -1500 1600 -1400
rect 4540 -1500 4640 -1400
rect 5765 -1550 5865 -1450
rect 1780 -1800 1840 -1700
rect 3680 -1800 3740 -1700
rect 3880 -1800 3940 -1700
rect 4070 -1800 4130 -1700
rect 4260 -1800 4320 -1700
rect 4450 -1800 4510 -1700
rect 4880 -1800 4940 -1700
rect 5080 -1800 5140 -1700
rect 5270 -1800 5330 -1700
rect 5460 -1800 5520 -1700
rect 5650 -1800 5710 -1700
rect 1680 -2300 1740 -2200
rect 1880 -2300 1940 -2200
rect 3580 -2300 3650 -2200
rect 3780 -2300 3840 -2200
rect 3970 -2300 4030 -2200
rect 4160 -2300 4220 -2200
rect 4350 -2300 4420 -2200
rect 4780 -2300 4850 -2200
rect 4980 -2300 5040 -2200
rect 5170 -2300 5230 -2200
rect 5360 -2300 5420 -2200
rect 5550 -2300 5610 -2200
rect 1500 -2650 1600 -2550
rect 4540 -2650 4640 -2570
rect 5765 -2650 5865 -2570
rect 1680 -2750 1740 -2698
rect 1880 -2750 1940 -2698
<< metal2 >>
rect 1640 200 1700 210
rect 1500 50 1600 56
rect 1500 -605 1600 -50
rect 1640 -300 1700 100
rect 1640 -410 1700 -400
rect 1830 200 1890 210
rect 1830 -300 1890 100
rect 1830 -410 1890 -400
rect 2020 200 2080 210
rect 2020 -300 2080 100
rect 2370 50 2472 56
rect 2020 -410 2080 -400
rect 2180 -300 2280 -45
rect 1500 -695 1505 -605
rect 1595 -695 1600 -605
rect 1500 -1150 1600 -695
rect 1500 -1400 1600 -1250
rect 1730 -900 1790 -890
rect 1730 -1290 1790 -1000
rect 1920 -900 1980 -890
rect 1730 -1300 1840 -1290
rect 1730 -1410 1840 -1400
rect 1920 -1300 1980 -1000
rect 1920 -1410 1980 -1400
rect 1500 -2550 1600 -1500
rect 1780 -1700 1840 -1410
rect 1780 -1810 1840 -1800
rect 1500 -2656 1600 -2650
rect 1680 -2200 1740 -2190
rect 1680 -2698 1740 -2300
rect 1680 -2760 1740 -2750
rect 1880 -2200 1940 -2190
rect 1880 -2698 1940 -2300
rect 2180 -2200 2280 -400
rect 2370 -50 2372 50
rect 2370 -56 2472 -50
rect 4560 50 4660 56
rect 2370 -1150 2470 -56
rect 2730 -294 2790 -284
rect 2730 -404 2790 -394
rect 2930 -294 2990 -284
rect 2930 -404 2990 -394
rect 3120 -294 3190 -284
rect 3120 -404 3190 -394
rect 3310 -294 3370 -284
rect 3310 -404 3370 -394
rect 3500 -294 3570 -284
rect 3500 -404 3570 -394
rect 3690 -294 3750 -284
rect 3690 -404 3750 -394
rect 3890 -294 3950 -284
rect 3890 -404 3950 -394
rect 4080 -294 4150 -284
rect 4080 -404 4150 -394
rect 4270 -294 4330 -284
rect 4270 -404 4330 -394
rect 4460 -294 4520 -284
rect 4460 -404 4520 -394
rect 2640 -800 2700 -790
rect 2640 -910 2700 -900
rect 2830 -800 2890 -790
rect 3020 -800 3080 -790
rect 3210 -800 3270 -790
rect 3410 -800 3470 -790
rect 2890 -900 2900 -800
rect 2830 -910 2900 -900
rect 3080 -900 3100 -800
rect 3020 -910 3100 -900
rect 2650 -1240 2700 -910
rect 2850 -1240 2900 -910
rect 3050 -1240 3100 -910
rect 2370 -1300 2470 -1250
rect 2370 -2005 2470 -1400
rect 2640 -1250 2700 -1240
rect 2640 -1410 2700 -1400
rect 2840 -1250 2900 -1240
rect 2840 -1410 2900 -1400
rect 3040 -1250 3100 -1240
rect 3040 -1410 3100 -1400
rect 3200 -900 3210 -800
rect 3200 -910 3270 -900
rect 3400 -900 3410 -800
rect 3400 -910 3470 -900
rect 3600 -800 3660 -790
rect 3600 -910 3660 -900
rect 3790 -800 3850 -790
rect 3790 -910 3850 -900
rect 3980 -800 4040 -790
rect 4170 -800 4230 -790
rect 4360 -800 4420 -790
rect 4040 -900 4050 -800
rect 3980 -910 4050 -900
rect 4230 -900 4250 -800
rect 4170 -910 4250 -900
rect 3200 -1240 3250 -910
rect 3400 -1240 3450 -910
rect 3600 -1240 3650 -910
rect 3800 -1240 3850 -910
rect 4000 -1240 4050 -910
rect 4200 -1240 4250 -910
rect 4350 -900 4360 -800
rect 4350 -910 4420 -900
rect 4350 -1240 4400 -910
rect 3200 -1250 3260 -1240
rect 3200 -1410 3260 -1400
rect 3400 -1250 3460 -1240
rect 3400 -1410 3460 -1400
rect 3600 -1250 3660 -1240
rect 3600 -1410 3660 -1400
rect 3800 -1250 3860 -1240
rect 3800 -1410 3860 -1400
rect 4000 -1250 4060 -1240
rect 4000 -1410 4060 -1400
rect 4200 -1250 4260 -1240
rect 4200 -1410 4260 -1400
rect 4340 -1250 4400 -1240
rect 4560 -1150 4660 -50
rect 6720 50 6820 56
rect 4880 -300 4940 -290
rect 4880 -410 4940 -400
rect 5080 -300 5140 -290
rect 5080 -410 5140 -400
rect 5270 -300 5340 -290
rect 5270 -410 5340 -400
rect 5460 -300 5520 -290
rect 5460 -410 5520 -400
rect 5650 -300 5720 -290
rect 5650 -410 5720 -400
rect 5840 -300 5900 -290
rect 5840 -410 5900 -400
rect 6040 -300 6100 -290
rect 6040 -410 6100 -400
rect 6230 -300 6300 -290
rect 6230 -410 6300 -400
rect 6420 -300 6480 -290
rect 6420 -410 6480 -400
rect 6610 -300 6680 -290
rect 6610 -410 6680 -400
rect 6720 -600 6820 -50
rect 6905 -300 6995 -296
rect 4790 -790 4840 -775
rect 4990 -790 5040 -775
rect 5190 -790 5240 -775
rect 4790 -800 4850 -790
rect 4790 -910 4850 -900
rect 4980 -800 5040 -790
rect 4980 -910 5040 -900
rect 5170 -800 5240 -790
rect 5230 -900 5240 -800
rect 5170 -910 5240 -900
rect 4790 -1240 4840 -910
rect 4990 -1240 5040 -910
rect 5190 -1240 5240 -910
rect 4560 -1256 4660 -1250
rect 4780 -1250 4840 -1240
rect 4340 -1410 4400 -1400
rect 4540 -1400 4640 -1390
rect 3700 -1500 3760 -1490
rect 3700 -1660 3760 -1650
rect 3880 -1500 3940 -1490
rect 3700 -1690 3750 -1660
rect 3680 -1700 3750 -1690
rect 3740 -1750 3750 -1700
rect 3880 -1700 3940 -1650
rect 3680 -1810 3740 -1800
rect 4060 -1500 4120 -1490
rect 4060 -1690 4120 -1650
rect 4260 -1500 4320 -1490
rect 4060 -1700 4130 -1690
rect 4060 -1800 4070 -1700
rect 3880 -1810 3940 -1800
rect 4070 -1810 4130 -1800
rect 4260 -1700 4320 -1650
rect 4440 -1500 4500 -1490
rect 4440 -1690 4500 -1650
rect 4780 -1410 4840 -1400
rect 4980 -1250 5040 -1240
rect 4980 -1410 5040 -1400
rect 5180 -1250 5240 -1240
rect 5180 -1410 5240 -1400
rect 5340 -790 5390 -775
rect 5540 -790 5590 -775
rect 5740 -790 5790 -775
rect 5940 -790 5990 -775
rect 6140 -790 6190 -775
rect 6340 -790 6390 -775
rect 5340 -800 5420 -790
rect 5340 -900 5360 -800
rect 5340 -910 5420 -900
rect 5540 -800 5620 -790
rect 5540 -900 5560 -800
rect 5540 -910 5620 -900
rect 5740 -800 5810 -790
rect 5740 -900 5750 -800
rect 5740 -910 5810 -900
rect 5940 -800 6000 -790
rect 5940 -910 6000 -900
rect 6130 -800 6190 -790
rect 6130 -910 6190 -900
rect 6320 -800 6390 -790
rect 6380 -900 6390 -800
rect 6320 -910 6390 -900
rect 5340 -1240 5390 -910
rect 5540 -1240 5590 -910
rect 5740 -1240 5790 -910
rect 5940 -1240 5990 -910
rect 6140 -1240 6190 -910
rect 6340 -1240 6390 -910
rect 6490 -790 6540 -775
rect 6490 -800 6570 -790
rect 6490 -900 6510 -800
rect 6490 -910 6570 -900
rect 6490 -1240 6540 -910
rect 5340 -1250 5400 -1240
rect 5340 -1410 5400 -1400
rect 5540 -1250 5600 -1240
rect 5540 -1410 5600 -1400
rect 5740 -1250 5800 -1240
rect 5740 -1411 5800 -1400
rect 5940 -1250 6000 -1240
rect 5940 -1410 6000 -1400
rect 6140 -1250 6200 -1240
rect 6140 -1410 6200 -1400
rect 6340 -1250 6400 -1240
rect 6340 -1410 6400 -1400
rect 6480 -1250 6540 -1240
rect 6720 -1150 6820 -700
rect 6720 -1256 6820 -1250
rect 6900 -305 7000 -300
rect 6900 -395 6905 -305
rect 6995 -395 7000 -305
rect 6480 -1410 6540 -1400
rect 5765 -1450 5865 -1444
rect 4440 -1700 4510 -1690
rect 4440 -1800 4450 -1700
rect 4260 -1810 4320 -1800
rect 4450 -1810 4510 -1800
rect 2370 -2095 2375 -2005
rect 2465 -2095 2470 -2005
rect 2370 -2146 2470 -2095
rect 2180 -2600 2280 -2300
rect 3580 -2200 3650 -2190
rect 3580 -2310 3650 -2300
rect 3780 -2200 3840 -2190
rect 3780 -2310 3840 -2300
rect 3970 -2200 4040 -2190
rect 3970 -2310 4040 -2300
rect 4160 -2200 4220 -2190
rect 4160 -2310 4220 -2300
rect 4350 -2200 4420 -2190
rect 4350 -2310 4420 -2300
rect 4540 -2570 4640 -1500
rect 4880 -1500 4940 -1490
rect 4880 -1700 4940 -1650
rect 4880 -1810 4940 -1800
rect 5080 -1500 5140 -1490
rect 5080 -1700 5140 -1650
rect 5280 -1500 5340 -1490
rect 5280 -1690 5340 -1650
rect 5080 -1810 5140 -1800
rect 5270 -1700 5340 -1690
rect 5330 -1800 5340 -1700
rect 5460 -1500 5520 -1490
rect 5460 -1700 5520 -1650
rect 5660 -1500 5720 -1490
rect 5660 -1690 5720 -1650
rect 5270 -1810 5330 -1800
rect 5460 -1810 5520 -1800
rect 5650 -1700 5720 -1690
rect 5710 -1800 5720 -1700
rect 5650 -1810 5710 -1800
rect 5765 -1996 5865 -1550
rect 5755 -2005 5865 -1996
rect 5845 -2095 5865 -2005
rect 5755 -2104 5865 -2095
rect 4780 -2200 4850 -2190
rect 4780 -2310 4850 -2300
rect 4980 -2200 5040 -2190
rect 4980 -2310 5040 -2300
rect 5170 -2200 5240 -2190
rect 5170 -2310 5240 -2300
rect 5360 -2200 5420 -2190
rect 5360 -2310 5420 -2300
rect 5550 -2200 5620 -2190
rect 5550 -2310 5620 -2300
rect 4540 -2660 4640 -2650
rect 5765 -2570 5865 -2104
rect 6900 -2200 7000 -395
rect 6900 -2309 7000 -2300
rect 5765 -2660 5865 -2650
rect 1880 -2760 1940 -2750
<< via2 >>
rect 2180 -400 2280 -300
rect 1505 -695 1595 -605
rect 1730 -1400 1840 -1300
rect 1920 -1400 1980 -1300
rect 2730 -394 2790 -294
rect 2930 -394 2990 -294
rect 3130 -394 3180 -294
rect 3180 -394 3190 -294
rect 3310 -394 3370 -294
rect 3510 -394 3560 -294
rect 3560 -394 3570 -294
rect 3690 -394 3750 -294
rect 3890 -394 3950 -294
rect 4090 -394 4140 -294
rect 4140 -394 4150 -294
rect 4270 -394 4330 -294
rect 4460 -394 4520 -294
rect 2370 -1400 2470 -1300
rect 2640 -1400 2700 -1250
rect 2840 -1400 2900 -1250
rect 3040 -1400 3100 -1250
rect 3200 -1400 3260 -1250
rect 3400 -1400 3460 -1250
rect 3600 -1400 3660 -1250
rect 3800 -1400 3860 -1250
rect 4000 -1400 4060 -1250
rect 4200 -1400 4260 -1250
rect 4340 -1400 4400 -1250
rect 4880 -400 4940 -300
rect 5080 -400 5140 -300
rect 5280 -400 5330 -300
rect 5330 -400 5340 -300
rect 5460 -400 5520 -300
rect 5660 -400 5710 -300
rect 5710 -400 5720 -300
rect 5840 -400 5900 -300
rect 6040 -400 6100 -300
rect 6240 -400 6290 -300
rect 6290 -400 6300 -300
rect 6420 -400 6480 -300
rect 6620 -400 6670 -300
rect 6670 -400 6680 -300
rect 6720 -700 6820 -600
rect 3700 -1650 3760 -1500
rect 3880 -1650 3940 -1500
rect 4060 -1650 4120 -1500
rect 4260 -1650 4320 -1500
rect 4440 -1650 4500 -1500
rect 4780 -1400 4840 -1250
rect 4980 -1400 5040 -1250
rect 5180 -1400 5240 -1250
rect 5340 -1400 5400 -1250
rect 5540 -1400 5600 -1250
rect 5740 -1400 5800 -1250
rect 5940 -1400 6000 -1250
rect 6140 -1400 6200 -1250
rect 6340 -1400 6400 -1250
rect 6480 -1400 6540 -1250
rect 6905 -395 6995 -305
rect 2375 -2095 2465 -2005
rect 2180 -2300 2280 -2200
rect 3580 -2300 3640 -2200
rect 3780 -2300 3840 -2200
rect 3980 -2300 4030 -2200
rect 4030 -2300 4040 -2200
rect 4160 -2300 4220 -2200
rect 4350 -2300 4420 -2200
rect 4880 -1650 4940 -1500
rect 5080 -1650 5140 -1500
rect 5280 -1650 5340 -1500
rect 5460 -1650 5520 -1500
rect 5660 -1650 5720 -1500
rect 5755 -2095 5845 -2005
rect 4780 -2300 4840 -2200
rect 4980 -2300 5040 -2200
rect 5180 -2300 5230 -2200
rect 5230 -2300 5240 -2200
rect 5360 -2300 5420 -2200
rect 5560 -2300 5610 -2200
rect 5610 -2300 5620 -2200
rect 6900 -2300 7000 -2200
<< metal3 >>
rect 2720 -294 2800 -289
rect 2920 -294 3000 -289
rect 3120 -294 3200 -289
rect 3300 -294 3380 -289
rect 3500 -294 3580 -289
rect 3680 -294 3760 -289
rect 3880 -294 3960 -289
rect 4080 -294 4160 -289
rect 4260 -294 4340 -289
rect 4401 -294 4540 -289
rect 2190 -295 2730 -294
rect 2175 -300 2730 -295
rect 2175 -400 2180 -300
rect 2280 -394 2730 -300
rect 2790 -394 2930 -294
rect 2990 -394 3130 -294
rect 3190 -394 3310 -294
rect 3370 -394 3510 -294
rect 3570 -394 3690 -294
rect 3750 -394 3890 -294
rect 3950 -394 4090 -294
rect 4150 -394 4270 -294
rect 4330 -394 4460 -294
rect 4520 -394 4540 -294
rect 4870 -300 4950 -295
rect 5070 -300 5150 -295
rect 5270 -300 5350 -295
rect 5450 -300 5530 -295
rect 5650 -300 5730 -295
rect 5830 -300 5910 -295
rect 6030 -300 6110 -295
rect 6230 -300 6310 -295
rect 6410 -300 6490 -295
rect 6610 -300 6690 -295
rect 2280 -400 2285 -394
rect 2720 -399 2800 -394
rect 2920 -399 3000 -394
rect 3120 -399 3200 -394
rect 3300 -399 3380 -394
rect 3500 -399 3580 -394
rect 3680 -399 3760 -394
rect 3880 -399 3960 -394
rect 4080 -399 4160 -394
rect 4260 -399 4340 -394
rect 4401 -399 4540 -394
rect 4780 -400 4880 -300
rect 4940 -400 5080 -300
rect 5140 -400 5280 -300
rect 5340 -400 5460 -300
rect 5520 -400 5660 -300
rect 5720 -400 5840 -300
rect 5900 -400 6040 -300
rect 6100 -400 6240 -300
rect 6300 -400 6420 -300
rect 6480 -400 6620 -300
rect 6680 -305 7000 -300
rect 6680 -395 6905 -305
rect 6995 -395 7000 -305
rect 6680 -400 7000 -395
rect 2175 -405 2285 -400
rect 4870 -405 4950 -400
rect 5070 -405 5150 -400
rect 5270 -405 5350 -400
rect 5450 -405 5530 -400
rect 5650 -405 5730 -400
rect 5830 -405 5910 -400
rect 6030 -405 6110 -400
rect 6230 -405 6310 -400
rect 6410 -405 6490 -400
rect 6610 -405 6690 -400
rect 6710 -600 6830 -595
rect 1500 -605 6720 -600
rect 1500 -695 1505 -605
rect 1595 -695 6720 -605
rect 1500 -700 6720 -695
rect 6820 -700 6830 -600
rect 6710 -705 6830 -700
rect 2630 -1250 2710 -1245
rect 2830 -1250 2910 -1245
rect 3030 -1250 3110 -1245
rect 3190 -1250 3270 -1245
rect 3390 -1250 3470 -1245
rect 3590 -1250 3670 -1245
rect 3790 -1250 3870 -1245
rect 3990 -1250 4070 -1245
rect 4190 -1250 4270 -1245
rect 4330 -1250 4410 -1245
rect 4770 -1250 4850 -1245
rect 4970 -1250 5050 -1245
rect 5170 -1250 5250 -1245
rect 5330 -1250 5410 -1245
rect 5530 -1250 5610 -1245
rect 5730 -1250 5810 -1245
rect 5930 -1250 6010 -1245
rect 6130 -1250 6210 -1245
rect 6330 -1250 6410 -1245
rect 6470 -1250 6550 -1245
rect 1720 -1300 1850 -1295
rect 1910 -1300 1990 -1295
rect 2365 -1300 2475 -1295
rect 1700 -1400 1730 -1300
rect 1840 -1400 1920 -1300
rect 1980 -1400 2370 -1300
rect 2470 -1400 2475 -1300
rect 1720 -1405 1850 -1400
rect 1910 -1405 1990 -1400
rect 2365 -1405 2475 -1400
rect 2630 -1400 2640 -1250
rect 2700 -1400 2840 -1250
rect 2900 -1400 3040 -1250
rect 3100 -1400 3200 -1250
rect 3260 -1400 3400 -1250
rect 3460 -1400 3600 -1250
rect 3660 -1400 3800 -1250
rect 3860 -1400 4000 -1250
rect 4060 -1400 4200 -1250
rect 4260 -1400 4340 -1250
rect 4400 -1400 4780 -1250
rect 4840 -1400 4980 -1250
rect 5040 -1400 5180 -1250
rect 5240 -1400 5340 -1250
rect 5400 -1400 5540 -1250
rect 5600 -1400 5740 -1250
rect 5800 -1400 5940 -1250
rect 6000 -1400 6140 -1250
rect 6200 -1400 6340 -1250
rect 6400 -1400 6480 -1250
rect 6540 -1400 6640 -1250
rect 2630 -1405 2710 -1400
rect 2830 -1405 2910 -1400
rect 3030 -1405 3110 -1400
rect 3190 -1405 3270 -1400
rect 3390 -1405 3470 -1400
rect 3590 -1405 3670 -1400
rect 3790 -1405 3870 -1400
rect 3990 -1405 4070 -1400
rect 4190 -1405 4270 -1400
rect 4330 -1405 4410 -1400
rect 3690 -1500 3770 -1495
rect 3870 -1500 3950 -1495
rect 4050 -1500 4130 -1495
rect 4250 -1500 4330 -1495
rect 4430 -1500 4510 -1495
rect 4580 -1500 4700 -1400
rect 4770 -1405 4850 -1400
rect 4970 -1405 5050 -1400
rect 5170 -1405 5250 -1400
rect 5330 -1405 5410 -1400
rect 5530 -1405 5610 -1400
rect 5730 -1405 5810 -1400
rect 5930 -1405 6010 -1400
rect 6130 -1405 6210 -1400
rect 6330 -1405 6410 -1400
rect 6470 -1405 6550 -1400
rect 4870 -1500 4950 -1495
rect 5070 -1500 5150 -1495
rect 5270 -1500 5350 -1495
rect 5450 -1500 5530 -1495
rect 5650 -1500 5730 -1495
rect 3500 -1650 3700 -1500
rect 3760 -1650 3880 -1500
rect 3940 -1650 4060 -1500
rect 4120 -1650 4260 -1500
rect 4320 -1650 4440 -1500
rect 4500 -1650 4880 -1500
rect 4940 -1650 5080 -1500
rect 5140 -1650 5280 -1500
rect 5340 -1650 5460 -1500
rect 5520 -1650 5660 -1500
rect 5720 -1650 5740 -1500
rect 3690 -1655 3770 -1650
rect 3870 -1655 3950 -1650
rect 4050 -1655 4130 -1650
rect 4250 -1655 4330 -1650
rect 4430 -1655 4510 -1650
rect 4870 -1655 4950 -1650
rect 5070 -1655 5150 -1650
rect 5270 -1655 5350 -1650
rect 5450 -1655 5530 -1650
rect 5650 -1655 5730 -1650
rect 2356 -2005 5850 -2000
rect 2356 -2095 2375 -2005
rect 2465 -2095 5755 -2005
rect 5845 -2095 5850 -2005
rect 2356 -2100 5850 -2095
rect 2175 -2200 2285 -2195
rect 3570 -2200 3650 -2195
rect 3770 -2200 3850 -2195
rect 3970 -2200 4050 -2195
rect 4150 -2200 4230 -2195
rect 4340 -2200 4430 -2195
rect 4770 -2200 4850 -2195
rect 4970 -2200 5050 -2195
rect 5170 -2200 5250 -2195
rect 5350 -2200 5430 -2195
rect 5550 -2200 5630 -2195
rect 6895 -2200 7005 -2195
rect 2175 -2300 2180 -2200
rect 2280 -2300 3580 -2200
rect 3640 -2300 3780 -2200
rect 3840 -2300 3980 -2200
rect 4040 -2300 4160 -2200
rect 4220 -2300 4350 -2200
rect 4420 -2300 4430 -2200
rect 4680 -2300 4780 -2200
rect 4840 -2300 4980 -2200
rect 5040 -2300 5180 -2200
rect 5240 -2300 5360 -2200
rect 5420 -2300 5560 -2200
rect 5620 -2300 6900 -2200
rect 7000 -2300 7005 -2200
rect 2175 -2305 2285 -2300
rect 3570 -2305 3650 -2300
rect 3770 -2305 3850 -2300
rect 3970 -2305 4050 -2300
rect 4150 -2305 4230 -2300
rect 4340 -2305 4430 -2300
rect 4770 -2305 4850 -2300
rect 4970 -2305 5050 -2300
rect 5170 -2305 5250 -2300
rect 5350 -2305 5430 -2300
rect 5550 -2305 5630 -2300
rect 6895 -2305 7005 -2300
use sky130_fd_pr__nfet_01v8_6H2JYD  sky130_fd_pr__nfet_01v8_6H2JYD_0
timestamp 1710000826
transform 1 0 1813 0 1 -2040
box -263 -710 263 710
use sky130_fd_pr__pfet_01v8_BDZ9JN  sky130_fd_pr__pfet_01v8_BDZ9JN_0
timestamp 1709390584
transform 1 0 3579 0 1 -581
box -1079 -719 1079 719
use sky130_fd_pr__pfet_01v8_UJHYGH  sky130_fd_pr__pfet_01v8_UJHYGH_0
timestamp 1709401415
transform 1 0 1859 0 1 -581
box -359 -719 359 719
use sky130_fd_pr__nfet_01v8_KBNS5F  XM2
timestamp 1709392794
transform 1 0 4049 0 1 -2040
box -599 -710 599 710
use sky130_fd_pr__pfet_01v8_BDZ9JN  XM3
timestamp 1709390584
transform 1 0 5729 0 1 -581
box -1079 -719 1079 719
use sky130_fd_pr__nfet_01v8_KBNS5F  XM4
timestamp 1709392794
transform 1 0 5249 0 1 -2040
box -599 -710 599 710
use sky130_fd_pr__nfet_01v8_J4PS55  XM5
timestamp 1713148681
transform 1 0 6723 0 1 -2146
box 0 0 1 1
use sky130_fd_pr__pfet_01v8_UGNTUG  XM8
timestamp 1713148681
transform 1 0 6154 0 1 -2084
box 0 0 1 1
<< labels >>
rlabel metal2 6900 -2200 7000 -395 1 VREF_N
port 9 n
rlabel metal2 2180 -2600 2280 -45 1 VREF_P
port 10 n
rlabel metal2 1500 -2550 1600 -50 1 VIN
port 13 n
rlabel metal3 4580 -1650 4700 -1250 1 OUT
port 8 n
rlabel metal1 1600 -2780 5720 -2680 1 VSS
port 12 n
rlabel metal1 2180 100 6800 200 1 VDD
port 14 n
<< end >>
