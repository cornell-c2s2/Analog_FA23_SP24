magic
tech sky130A
magscale 1 2
timestamp 1716866472
<< metal4 >>
rect -3349 3039 3349 3080
rect -3349 -3039 3093 3039
rect 3329 -3039 3349 3039
rect -3349 -3080 3349 -3039
<< via4 >>
rect 3093 -3039 3329 3039
<< mimcap2 >>
rect -3269 2960 2731 3000
rect -3269 -2960 -3229 2960
rect 2691 -2960 2731 2960
rect -3269 -3000 2731 -2960
<< mimcap2contact >>
rect -3229 -2960 2691 2960
<< metal5 >>
rect 3051 3039 3371 3081
rect -3253 2960 2715 2984
rect -3253 -2960 -3229 2960
rect 2691 -2960 2715 2960
rect -3253 -2984 2715 -2960
rect 3051 -3039 3093 3039
rect 3329 -3039 3371 3039
rect 3051 -3081 3371 -3039
<< properties >>
string FIXED_BBOX -3349 -3080 2811 3080
string gencell sky130_fd_pr__cap_mim_m3_2
string library sky130
string parameters w 30.0 l 30.0 val 1.822k carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
