magic
tech sky130A
magscale 1 2
timestamp 1709401415
<< error_p >>
rect -77 581 -19 587
rect 115 581 173 587
rect -77 547 -65 581
rect 115 547 127 581
rect -77 541 -19 547
rect 115 541 173 547
rect -173 -547 -115 -541
rect 19 -547 77 -541
rect -173 -581 -161 -547
rect 19 -581 31 -547
rect -173 -587 -115 -581
rect 19 -587 77 -581
<< nwell >>
rect -359 -719 359 719
<< pmos >>
rect -159 -500 -129 500
rect -63 -500 -33 500
rect 33 -500 63 500
rect 129 -500 159 500
<< pdiff >>
rect -221 488 -159 500
rect -221 -488 -209 488
rect -175 -488 -159 488
rect -221 -500 -159 -488
rect -129 488 -63 500
rect -129 -488 -113 488
rect -79 -488 -63 488
rect -129 -500 -63 -488
rect -33 488 33 500
rect -33 -488 -17 488
rect 17 -488 33 488
rect -33 -500 33 -488
rect 63 488 129 500
rect 63 -488 79 488
rect 113 -488 129 488
rect 63 -500 129 -488
rect 159 488 221 500
rect 159 -488 175 488
rect 209 -488 221 488
rect 159 -500 221 -488
<< pdiffc >>
rect -209 -488 -175 488
rect -113 -488 -79 488
rect -17 -488 17 488
rect 79 -488 113 488
rect 175 -488 209 488
<< nsubdiff >>
rect -323 649 -227 683
rect 227 649 323 683
rect -323 587 -289 649
rect 289 587 323 649
rect -323 -649 -289 -587
rect 289 -649 323 -587
rect -323 -683 -227 -649
rect 227 -683 323 -649
<< nsubdiffcont >>
rect -227 649 227 683
rect -323 -587 -289 587
rect 289 -587 323 587
rect -227 -683 227 -649
<< poly >>
rect -81 581 -15 597
rect -81 547 -65 581
rect -31 547 -15 581
rect -81 531 -15 547
rect 111 581 177 597
rect 111 547 127 581
rect 161 547 177 581
rect 111 531 177 547
rect -159 500 -129 526
rect -63 500 -33 531
rect 33 500 63 526
rect 129 500 159 531
rect -159 -531 -129 -500
rect -63 -526 -33 -500
rect 33 -531 63 -500
rect 129 -526 159 -500
rect -177 -547 -111 -531
rect -177 -581 -161 -547
rect -127 -581 -111 -547
rect -177 -597 -111 -581
rect 15 -547 81 -531
rect 15 -581 31 -547
rect 65 -581 81 -547
rect 15 -597 81 -581
<< polycont >>
rect -65 547 -31 581
rect 127 547 161 581
rect -161 -581 -127 -547
rect 31 -581 65 -547
<< locali >>
rect -323 649 -227 683
rect 227 649 323 683
rect -323 587 -289 649
rect 289 587 323 649
rect -81 547 -65 581
rect -31 547 -15 581
rect 111 547 127 581
rect 161 547 177 581
rect -209 488 -175 504
rect -209 -504 -175 -488
rect -113 488 -79 504
rect -113 -504 -79 -488
rect -17 488 17 504
rect -17 -504 17 -488
rect 79 488 113 504
rect 79 -504 113 -488
rect 175 488 209 504
rect 175 -504 209 -488
rect -177 -581 -161 -547
rect -127 -581 -111 -547
rect 15 -581 31 -547
rect 65 -581 81 -547
rect -323 -649 -289 -587
rect 289 -649 323 -587
rect -323 -683 -227 -649
rect 227 -683 323 -649
<< viali >>
rect -65 547 -31 581
rect 127 547 161 581
rect -209 -488 -175 488
rect -113 -488 -79 488
rect -17 -488 17 488
rect 79 -488 113 488
rect 175 -488 209 488
rect -161 -581 -127 -547
rect 31 -581 65 -547
<< metal1 >>
rect -77 581 -19 587
rect -77 547 -65 581
rect -31 547 -19 581
rect -77 541 -19 547
rect 115 581 173 587
rect 115 547 127 581
rect 161 547 173 581
rect 115 541 173 547
rect -215 488 -169 500
rect -215 -488 -209 488
rect -175 -488 -169 488
rect -215 -500 -169 -488
rect -119 488 -73 500
rect -119 -488 -113 488
rect -79 -488 -73 488
rect -119 -500 -73 -488
rect -23 488 23 500
rect -23 -488 -17 488
rect 17 -488 23 488
rect -23 -500 23 -488
rect 73 488 119 500
rect 73 -488 79 488
rect 113 -488 119 488
rect 73 -500 119 -488
rect 169 488 215 500
rect 169 -488 175 488
rect 209 -488 215 488
rect 169 -500 215 -488
rect -173 -547 -115 -541
rect -173 -581 -161 -547
rect -127 -581 -115 -547
rect -173 -587 -115 -581
rect 19 -547 77 -541
rect 19 -581 31 -547
rect 65 -581 77 -547
rect 19 -587 77 -581
<< properties >>
string FIXED_BBOX -306 -666 306 666
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 5 l 0.15 m 1 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
