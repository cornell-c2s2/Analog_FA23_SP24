magic
tech sky130A
magscale 1 2
timestamp 1712465298
<< error_s >>
rect 20 488 130 490
rect 3393 -2385 3451 -2301
rect 3481 -2385 3533 -2301
rect 515 -2745 567 -2661
rect 597 -2745 667 -2661
<< nwell >>
rect -1610 -250 3790 180
rect 450 -320 3790 -250
rect 450 -560 2830 -320
rect 450 -1640 3790 -1180
rect 450 -1880 2480 -1640
rect 450 -2970 3800 -2500
<< pwell >>
rect -1550 494 -247 500
rect -1550 230 170 494
rect 10 -760 2830 -610
rect 10 -1120 3200 -760
rect 10 -2080 2510 -1930
rect 10 -2410 3560 -2080
<< psubdiff >>
rect 20 460 130 490
rect 20 410 50 460
rect 100 410 130 460
rect 20 340 130 410
rect 20 290 50 340
rect 100 290 130 340
rect 20 260 130 290
rect 30 -850 410 -820
rect 30 -900 60 -850
rect 110 -900 200 -850
rect 250 -900 330 -850
rect 380 -900 410 -850
rect 30 -930 410 -900
rect 40 -2170 440 -2140
rect 40 -2220 70 -2170
rect 120 -2220 220 -2170
rect 270 -2220 360 -2170
rect 410 -2220 440 -2170
rect 40 -2250 440 -2220
<< nsubdiff >>
rect -160 0 -50 30
rect -160 -50 -130 0
rect -80 -50 -50 0
rect -160 -130 -50 -50
rect -160 -180 -130 -130
rect -80 -180 -50 -130
rect -160 -210 -50 -180
rect 2860 -170 2970 -140
rect 2860 -220 2890 -170
rect 2940 -220 2970 -170
rect 2860 -250 2970 -220
rect 3080 -170 3190 -140
rect 3080 -220 3110 -170
rect 3160 -220 3190 -170
rect 3080 -250 3190 -220
rect 3310 -170 3420 -140
rect 3310 -220 3340 -170
rect 3390 -220 3420 -170
rect 3310 -250 3420 -220
rect 3530 -170 3640 -140
rect 3530 -220 3560 -170
rect 3610 -220 3640 -170
rect 3530 -250 3640 -220
rect 3260 -1500 3370 -1470
rect 3260 -1550 3290 -1500
rect 3340 -1550 3370 -1500
rect 3260 -1580 3370 -1550
rect 3440 -1500 3550 -1470
rect 3440 -1550 3470 -1500
rect 3520 -1550 3550 -1500
rect 3440 -1580 3550 -1550
rect 3620 -1500 3730 -1470
rect 3620 -1550 3650 -1500
rect 3700 -1550 3730 -1500
rect 3620 -1580 3730 -1550
rect 3620 -2760 3730 -2730
rect 3620 -2810 3650 -2760
rect 3700 -2810 3730 -2760
rect 3620 -2850 3730 -2810
rect 3620 -2900 3650 -2850
rect 3700 -2900 3730 -2850
rect 3620 -2930 3730 -2900
<< psubdiffcont >>
rect 50 410 100 460
rect 50 290 100 340
rect 60 -900 110 -850
rect 200 -900 250 -850
rect 330 -900 380 -850
rect 70 -2220 120 -2170
rect 220 -2220 270 -2170
rect 360 -2220 410 -2170
<< nsubdiffcont >>
rect -130 -50 -80 0
rect -130 -180 -80 -130
rect 2890 -220 2940 -170
rect 3110 -220 3160 -170
rect 3340 -220 3390 -170
rect 3560 -220 3610 -170
rect 3290 -1550 3340 -1500
rect 3470 -1550 3520 -1500
rect 3650 -1550 3700 -1500
rect 3650 -2810 3700 -2760
rect 3650 -2900 3700 -2850
<< locali >>
rect 623 -350 657 -349
rect 745 -350 779 -349
rect 518 -586 552 -552
rect 619 -604 653 -570
rect 698 -601 732 -567
<< viali >>
rect 20 460 130 490
rect 20 410 50 460
rect 50 410 100 460
rect 100 410 130 460
rect 20 340 130 410
rect -1420 279 -1386 313
rect -1148 276 -1114 310
rect -873 277 -839 311
rect -598 277 -564 311
rect -322 275 -288 309
rect 20 290 50 340
rect 50 290 100 340
rect 100 290 130 340
rect 20 260 130 290
rect -1510 180 -1470 220
rect -1420 187 -1386 221
rect -1228 193 -1194 227
rect -1143 187 -1109 221
rect -962 186 -928 220
rect -866 186 -832 220
rect -686 187 -652 221
rect -593 187 -559 221
rect -410 187 -376 221
rect -318 186 -284 220
rect -1420 98 -1386 132
rect -1147 93 -1113 127
rect -875 92 -841 126
rect -598 93 -564 127
rect -322 93 -288 127
rect -872 20 -838 54
rect -160 0 -50 30
rect -160 -50 -130 0
rect -130 -50 -80 0
rect -80 -50 -50 0
rect -160 -130 -50 -50
rect -160 -180 -130 -130
rect -130 -180 -80 -130
rect -80 -180 -50 -130
rect -160 -210 -50 -180
rect 2860 -170 2970 -140
rect 2860 -220 2890 -170
rect 2890 -220 2940 -170
rect 2940 -220 2970 -170
rect 2860 -250 2970 -220
rect 3080 -170 3190 -140
rect 3080 -220 3110 -170
rect 3110 -220 3160 -170
rect 3160 -220 3190 -170
rect 3080 -250 3190 -220
rect 3310 -170 3420 -140
rect 3310 -220 3340 -170
rect 3340 -220 3390 -170
rect 3390 -220 3420 -170
rect 3310 -250 3420 -220
rect 3530 -170 3640 -140
rect 3530 -220 3560 -170
rect 3560 -220 3610 -170
rect 3610 -220 3640 -170
rect 3530 -250 3640 -220
rect 532 -386 567 -351
rect 622 -386 657 -350
rect 745 -386 780 -350
rect 618 -526 652 -492
rect 697 -525 731 -491
rect 806 -598 845 -559
rect 518 -658 552 -624
rect 30 -850 410 -820
rect 30 -900 60 -850
rect 60 -900 110 -850
rect 110 -900 200 -850
rect 200 -900 250 -850
rect 250 -900 330 -850
rect 330 -900 380 -850
rect 380 -900 410 -850
rect 30 -930 410 -900
rect 3260 -1500 3370 -1470
rect 3260 -1550 3290 -1500
rect 3290 -1550 3340 -1500
rect 3340 -1550 3370 -1500
rect 3260 -1580 3370 -1550
rect 3440 -1500 3550 -1470
rect 3440 -1550 3470 -1500
rect 3470 -1550 3520 -1500
rect 3520 -1550 3550 -1500
rect 3440 -1580 3550 -1550
rect 3620 -1500 3730 -1470
rect 3620 -1550 3650 -1500
rect 3650 -1550 3700 -1500
rect 3700 -1550 3730 -1500
rect 3620 -1580 3730 -1550
rect 40 -2170 440 -2140
rect 40 -2220 70 -2170
rect 70 -2220 120 -2170
rect 120 -2220 220 -2170
rect 220 -2220 270 -2170
rect 270 -2220 360 -2170
rect 360 -2220 410 -2170
rect 410 -2220 440 -2170
rect 40 -2250 440 -2220
rect 3620 -2760 3730 -2730
rect 3620 -2810 3650 -2760
rect 3650 -2810 3700 -2760
rect 3700 -2810 3730 -2760
rect 3620 -2850 3730 -2810
rect 3620 -2900 3650 -2850
rect 3650 -2900 3700 -2850
rect 3700 -2900 3730 -2850
rect 3620 -2930 3730 -2900
<< metal1 >>
rect -3910 470 -3710 690
rect -3910 280 -3870 470
rect -3750 280 -3710 470
rect -3910 270 -3710 280
rect -3660 470 -3460 690
rect -3660 280 -3620 470
rect -3500 280 -3460 470
rect -3660 270 -3460 280
rect -3410 470 -3210 690
rect -3410 280 -3370 470
rect -3250 280 -3210 470
rect -3410 270 -3210 280
rect -3160 470 -2960 690
rect -3160 280 -3120 470
rect -3000 280 -2960 470
rect -3160 270 -2960 280
rect -2910 470 -2710 690
rect -2910 280 -2870 470
rect -2750 280 -2710 470
rect -2910 270 -2710 280
rect -2660 470 -2460 690
rect -2660 280 -2620 470
rect -2500 280 -2460 470
rect -2660 270 -2460 280
rect -2410 470 -2210 690
rect -2410 280 -2370 470
rect -2250 280 -2210 470
rect -2410 270 -2210 280
rect -2160 470 -1960 690
rect -2160 280 -2120 470
rect -2000 280 -1960 470
rect -2160 270 -1960 280
rect -1910 470 -1710 690
rect -1677 520 -1664 585
rect -1599 533 741 585
rect -1599 520 -286 533
rect -210 490 170 494
rect -1910 280 -1870 470
rect -1750 280 -1710 470
rect -1590 420 20 490
rect -1590 390 -170 420
rect -1429 330 -1362 336
rect -1910 270 -1710 280
rect -1430 313 -1362 330
rect -1430 279 -1420 313
rect -1386 279 -1362 313
rect -1430 260 -1362 279
rect -1157 310 -1079 338
rect -325 332 -273 338
rect -1157 276 -1148 310
rect -1114 276 -1079 310
rect -1157 260 -1079 276
rect -886 311 -822 327
rect -886 277 -873 311
rect -839 277 -822 311
rect -886 260 -822 277
rect -607 311 -541 324
rect -607 277 -598 311
rect -564 277 -541 311
rect -1430 247 -1326 260
rect -1530 234 -1460 240
rect -3380 182 -3367 234
rect -3250 182 -1677 234
rect -1625 220 -1460 234
rect -1625 182 -1510 220
rect -1530 180 -1510 182
rect -1470 180 -1460 220
rect -1530 160 -1460 180
rect -1430 221 -1417 247
rect -1430 187 -1420 221
rect -1430 169 -1417 187
rect -1339 169 -1326 247
rect -1430 156 -1326 169
rect -1250 248 -1190 249
rect -1250 227 -1188 248
rect -1250 193 -1228 227
rect -1194 193 -1188 227
rect -1250 167 -1188 193
rect -1157 247 -1053 260
rect -1157 169 -1144 247
rect -1066 169 -1053 247
rect -1157 156 -1053 169
rect -988 247 -923 260
rect -886 247 -767 260
rect -607 247 -541 277
rect -331 309 -273 332
rect -331 275 -322 309
rect -288 275 -273 309
rect -331 247 -273 275
rect -208 300 -170 390
rect -30 300 20 420
rect -208 260 20 300
rect 130 260 170 490
rect -208 250 170 260
rect -923 169 -922 234
rect -886 220 -858 247
rect -886 186 -866 220
rect -886 169 -858 186
rect -780 169 -767 247
rect -988 156 -923 169
rect -886 156 -767 169
rect -728 236 -637 247
rect -728 221 -635 236
rect -728 187 -686 221
rect -652 187 -635 221
rect -728 167 -635 187
rect -607 234 -494 247
rect -607 221 -585 234
rect -607 187 -593 221
rect -607 169 -585 187
rect -507 169 -494 234
rect -728 156 -637 167
rect -607 156 -494 169
rect -455 234 -364 247
rect -455 156 -442 234
rect -1430 132 -1362 156
rect -1430 98 -1420 132
rect -1386 98 -1362 132
rect -1430 80 -1362 98
rect -1157 127 -1079 156
rect -1157 93 -1147 127
rect -1113 93 -1079 127
rect -1157 52 -1079 93
rect -2886 0 -2873 52
rect -2756 0 -1079 52
rect -886 126 -822 156
rect -886 92 -875 126
rect -841 92 -822 126
rect -886 54 -822 92
rect -607 127 -541 156
rect -455 143 -364 156
rect -331 234 -247 247
rect -331 220 -299 234
rect -331 186 -318 220
rect -331 156 -299 186
rect -331 143 -247 156
rect -607 93 -598 127
rect -564 93 -541 127
rect -607 76 -541 93
rect -331 127 -273 143
rect -331 93 -322 127
rect -288 93 -273 127
rect -331 74 -273 93
rect -886 20 -872 54
rect -838 20 -822 54
rect -886 7 -822 20
rect -325 0 -273 74
rect -240 40 4220 70
rect -240 30 80 40
rect -240 -50 -160 30
rect -1590 -150 -160 -50
rect -240 -210 -160 -150
rect -50 -210 80 30
rect 340 -90 4220 40
rect 340 -140 3960 -90
rect 340 -210 2860 -140
rect -240 -250 2860 -210
rect 2970 -250 3080 -140
rect 3190 -250 3310 -140
rect 3420 -250 3530 -140
rect 3640 -250 3960 -140
rect 480 -290 3960 -250
rect 4160 -290 4220 -90
rect 5540 -270 5740 -70
rect 480 -312 4220 -290
rect -312 -351 -221 -338
rect -312 -416 -299 -351
rect -234 -416 -221 -351
rect -312 -429 -221 -416
rect 299 -351 403 -338
rect 507 -350 831 -343
rect 507 -351 622 -350
rect 299 -416 312 -351
rect 390 -386 532 -351
rect 567 -386 622 -351
rect 657 -386 745 -350
rect 780 -386 831 -350
rect 390 -403 831 -386
rect 390 -416 559 -403
rect 299 -429 403 -416
rect -299 -455 -234 -429
rect 612 -485 752 -484
rect 604 -488 752 -485
rect 603 -491 754 -488
rect 603 -492 697 -491
rect 603 -526 618 -492
rect 652 -525 697 -492
rect 731 -525 754 -491
rect 652 -526 754 -525
rect 603 -546 754 -526
rect 793 -559 884 -546
rect 506 -624 575 -598
rect 793 -611 806 -559
rect 858 -611 884 -559
rect 793 -624 884 -611
rect 506 -658 518 -624
rect 552 -658 575 -624
rect 506 -663 575 -658
rect 506 -665 573 -663
rect 5540 -670 5740 -470
rect -220 -770 3200 -760
rect -220 -980 -180 -770
rect -20 -820 3200 -770
rect -20 -930 30 -820
rect 410 -930 3200 -820
rect -20 -980 3200 -930
rect -220 -990 10 -980
rect 5540 -1070 5740 -870
rect 480 -1430 4220 -1410
rect 480 -1470 3960 -1430
rect 480 -1580 3260 -1470
rect 3370 -1580 3440 -1470
rect 3550 -1580 3620 -1470
rect 3730 -1580 3960 -1470
rect 480 -1620 3960 -1580
rect 4160 -1620 4220 -1430
rect 5540 -1470 5740 -1270
rect 480 -1640 4220 -1620
rect -220 -2090 3560 -2080
rect -220 -2290 -180 -2090
rect -20 -2140 3560 -2090
rect -20 -2250 40 -2140
rect 440 -2250 3560 -2140
rect -20 -2290 3560 -2250
rect -220 -2300 3560 -2290
rect 480 -2730 4280 -2720
rect 480 -2930 3620 -2730
rect 3730 -2810 4280 -2730
rect 3730 -2880 4020 -2810
rect 4090 -2880 4280 -2810
rect 3730 -2930 4280 -2880
rect 480 -2970 4280 -2930
<< via1 >>
rect -3870 280 -3750 470
rect -3620 280 -3500 470
rect -3370 280 -3250 470
rect -3120 280 -3000 470
rect -2870 280 -2750 470
rect -2620 280 -2500 470
rect -2370 280 -2250 470
rect -2120 280 -2000 470
rect -1664 520 -1599 585
rect -1870 280 -1750 470
rect -3367 182 -3250 234
rect -1677 182 -1625 234
rect -1417 221 -1339 247
rect -1417 187 -1386 221
rect -1386 187 -1339 221
rect -1417 169 -1339 187
rect -1144 221 -1066 247
rect -1144 187 -1143 221
rect -1143 187 -1109 221
rect -1109 187 -1066 221
rect -1144 169 -1066 187
rect -988 220 -923 247
rect -170 300 -30 420
rect -988 186 -962 220
rect -962 186 -928 220
rect -928 186 -923 220
rect -988 169 -923 186
rect -858 220 -780 247
rect -858 186 -832 220
rect -832 186 -780 220
rect -858 169 -780 186
rect -585 221 -507 234
rect -585 187 -559 221
rect -559 187 -507 221
rect -585 169 -507 187
rect -442 221 -364 234
rect -442 187 -410 221
rect -410 187 -376 221
rect -376 187 -364 221
rect -442 156 -364 187
rect -2873 0 -2756 52
rect -299 220 -247 234
rect -299 186 -284 220
rect -284 186 -247 220
rect -299 156 -247 186
rect 80 -210 340 40
rect 3960 -290 4160 -90
rect -299 -416 -234 -351
rect 312 -416 390 -351
rect 806 -598 845 -559
rect 845 -598 858 -559
rect 806 -611 858 -598
rect -180 -980 -20 -770
rect 3960 -1620 4160 -1430
rect -180 -2290 -20 -2090
rect 4020 -2880 4090 -2810
<< metal2 >>
rect -1690 585 -1573 598
rect -1690 520 -1664 585
rect -1599 520 -1573 585
rect -1690 507 -1573 520
rect -3880 470 -3740 480
rect -3880 280 -3870 470
rect -3750 280 -3740 470
rect -3880 -533 -3740 280
rect -3880 -624 -3874 -533
rect -3757 -624 -3740 -533
rect -3880 -650 -3740 -624
rect -3630 470 -3490 480
rect -3630 280 -3620 470
rect -3500 280 -3490 470
rect -3630 -338 -3490 280
rect -3630 -429 -3614 -338
rect -3510 -429 -3490 -338
rect -3630 -3090 -3490 -429
rect -3380 470 -3240 480
rect -3380 280 -3370 470
rect -3250 280 -3240 470
rect -3380 234 -3240 280
rect -3380 182 -3367 234
rect -3250 182 -3240 234
rect -3380 -3090 -3240 182
rect -3130 470 -2990 480
rect -3130 280 -3120 470
rect -3000 280 -2990 470
rect -3130 -3090 -2990 280
rect -2880 470 -2740 480
rect -2880 280 -2870 470
rect -2750 280 -2740 470
rect -2880 52 -2740 280
rect -2880 0 -2873 52
rect -2756 0 -2740 52
rect -2880 -3090 -2740 0
rect -2630 470 -2490 480
rect -2630 280 -2620 470
rect -2500 280 -2490 470
rect -2630 260 -2490 280
rect -2630 156 -2613 260
rect -2496 156 -2490 260
rect -2630 -3090 -2490 156
rect -2380 470 -2240 480
rect -2380 280 -2370 470
rect -2250 280 -2240 470
rect -2380 78 -2240 280
rect -2380 0 -2366 78
rect -2249 0 -2240 78
rect -2380 -3090 -2240 0
rect -2130 470 -1990 480
rect -2130 280 -2120 470
rect -2000 280 -1990 470
rect -2130 -3090 -1990 280
rect -1880 470 -1740 480
rect -1880 280 -1870 470
rect -1750 280 -1740 470
rect -1880 -3090 -1740 280
rect -1690 234 -1612 507
rect -180 420 -20 430
rect -455 390 -351 403
rect -455 325 -442 390
rect -364 325 -351 390
rect -1690 182 -1677 234
rect -1625 182 -1612 234
rect -1690 169 -1612 182
rect -1443 247 -1313 260
rect -1443 169 -1417 247
rect -1339 169 -1313 247
rect -1443 -3094 -1313 169
rect -1157 247 -1027 260
rect -1157 169 -1144 247
rect -1066 169 -1027 247
rect -1157 -3094 -1027 169
rect -988 247 -897 260
rect -910 169 -897 247
rect -988 156 -897 169
rect -858 247 -767 260
rect -780 169 -767 247
rect -858 -52 -767 169
rect -728 104 -637 247
rect -598 234 -494 247
rect -598 169 -585 234
rect -507 169 -494 234
rect -598 156 -494 169
rect -728 26 -715 104
rect -650 26 -637 104
rect -728 13 -637 26
rect -871 -3094 -767 -52
rect -585 -3094 -494 156
rect -455 234 -351 325
rect -180 300 -170 420
rect -30 300 -20 420
rect -180 290 -20 300
rect -455 156 -442 234
rect -364 156 -351 234
rect -455 143 -351 156
rect -312 234 -221 247
rect -312 156 -299 234
rect -247 156 -221 234
rect -312 -351 -221 156
rect 70 40 350 50
rect 70 -210 80 40
rect 340 -210 350 40
rect 70 -220 350 -210
rect 3930 -80 4190 -70
rect 3930 -310 3940 -80
rect 4180 -310 4190 -80
rect 3930 -320 4190 -310
rect -312 -416 -299 -351
rect -234 -416 -221 -351
rect -312 -3094 -221 -416
rect 299 -351 403 -338
rect 299 -416 312 -351
rect 390 -416 403 -351
rect 299 -429 403 -416
rect 780 -546 897 -533
rect 780 -611 793 -546
rect 884 -611 897 -546
rect 780 -624 897 -611
rect -190 -770 -10 -760
rect -190 -980 -180 -770
rect -20 -980 -10 -770
rect -190 -990 -10 -980
rect 3940 -1430 4180 -1420
rect 3940 -1620 3960 -1430
rect 4160 -1620 4180 -1430
rect 3940 -1630 4180 -1620
rect -190 -2090 -10 -2080
rect -190 -2290 -180 -2090
rect -20 -2290 -10 -2090
rect -190 -2300 -10 -2290
rect 4010 -2810 4100 -2800
rect 4010 -2880 4020 -2810
rect 4090 -2880 4100 -2810
rect 4010 -2890 4100 -2880
<< via2 >>
rect -3874 -624 -3757 -533
rect -3614 -429 -3510 -338
rect -2613 156 -2496 260
rect -2366 0 -2249 78
rect -1859 338 -1768 403
rect -442 325 -364 390
rect -988 169 -923 247
rect -923 169 -910 247
rect -715 26 -650 104
rect -170 300 -30 420
rect 80 -210 340 40
rect 3940 -90 4180 -80
rect 3940 -290 3960 -90
rect 3960 -290 4160 -90
rect 4160 -290 4180 -90
rect 3940 -310 4180 -290
rect 312 -416 390 -351
rect 793 -559 884 -546
rect 793 -611 806 -559
rect 806 -611 858 -559
rect 858 -611 884 -559
rect -180 -980 -20 -770
rect 3960 -1620 4160 -1430
rect -180 -2290 -20 -2090
rect 4020 -2880 4090 -2810
<< metal3 >>
rect -190 430 -10 440
rect -1885 403 -1729 416
rect -1885 338 -1859 403
rect -1768 390 -1729 403
rect -455 390 -351 403
rect -1768 338 -442 390
rect -1885 325 -442 338
rect -364 325 -351 390
rect -455 312 -351 325
rect -190 290 -180 430
rect -20 290 -10 430
rect -190 280 -10 290
rect -2639 260 -2470 273
rect -2639 156 -2613 260
rect -2496 247 -897 260
rect -2496 169 -988 247
rect -910 169 -897 247
rect -2496 156 -897 169
rect -2639 143 -2470 156
rect -728 104 -637 117
rect -728 91 -715 104
rect -2379 78 -715 91
rect -2379 0 -2366 78
rect -2249 26 -715 78
rect -650 26 -637 104
rect -2249 13 -637 26
rect 70 40 350 50
rect -2249 0 -2236 13
rect -2379 -13 -2236 0
rect 70 -210 80 40
rect 340 -210 350 40
rect 70 -220 350 -210
rect 3930 -80 4190 -70
rect 3930 -310 3940 -80
rect 4180 -310 4190 -80
rect 3930 -320 4190 -310
rect -3627 -338 -3484 -325
rect -3627 -429 -3614 -338
rect -3510 -351 403 -338
rect -3510 -416 312 -351
rect 390 -416 403 -351
rect -3510 -429 403 -416
rect -3627 -442 -3484 -429
rect -3887 -533 -3744 -520
rect -3887 -624 -3874 -533
rect -3757 -546 897 -533
rect -3757 -611 793 -546
rect 884 -611 897 -546
rect -3757 -624 897 -611
rect -3887 -637 -3744 -624
rect -190 -770 -10 -760
rect -190 -980 -180 -770
rect -20 -980 -10 -770
rect -190 -990 -10 -980
rect 3930 -1420 4190 -1410
rect 3930 -1630 3940 -1420
rect 4180 -1630 4190 -1420
rect 3930 -1640 4190 -1630
rect -190 -2090 -10 -2080
rect -190 -2290 -180 -2090
rect -20 -2290 -10 -2090
rect -190 -2300 -10 -2290
rect 3990 -2790 4120 -2780
rect 3990 -2900 4000 -2790
rect 4110 -2900 4120 -2790
rect 3990 -2910 4120 -2900
<< via3 >>
rect -180 420 -20 430
rect -180 300 -170 420
rect -170 300 -30 420
rect -30 300 -20 420
rect -180 290 -20 300
rect 80 -210 340 40
rect 3940 -310 4180 -80
rect -180 -980 -20 -770
rect 3940 -1430 4180 -1420
rect 3940 -1620 3960 -1430
rect 3960 -1620 4160 -1430
rect 4160 -1620 4180 -1430
rect 3940 -1630 4180 -1620
rect -180 -2290 -20 -2090
rect 4000 -2810 4110 -2790
rect 4000 -2880 4020 -2810
rect 4020 -2880 4090 -2810
rect 4090 -2880 4110 -2810
rect 4000 -2900 4110 -2880
<< metal4 >>
rect -190 430 -10 440
rect -190 290 -180 430
rect -20 290 -10 430
rect -190 -770 -10 290
rect 70 40 350 50
rect 70 -210 80 40
rect 340 -210 350 40
rect 70 -220 350 -210
rect -190 -980 -180 -770
rect -20 -980 -10 -770
rect -190 -2090 -10 -980
rect 3900 -1400 4220 -1390
rect 3900 -1650 3930 -1400
rect 4190 -1650 4220 -1400
rect 3900 -1660 4220 -1650
rect -190 -2290 -180 -2090
rect -20 -2290 -10 -2090
rect -190 -2300 -10 -2290
<< via4 >>
rect 80 -210 340 40
rect 3930 -80 4190 -70
rect 3930 -310 3940 -80
rect 3940 -310 4180 -80
rect 4180 -310 4190 -80
rect 3930 -320 4190 -310
rect 3930 -1420 4190 -1400
rect 3930 -1630 3940 -1420
rect 3940 -1630 4180 -1420
rect 4180 -1630 4190 -1420
rect 3930 -1650 4190 -1630
rect 3930 -2790 4190 -2720
rect 3930 -2900 4000 -2790
rect 4000 -2900 4110 -2790
rect 4110 -2900 4190 -2790
rect 3930 -2970 4190 -2900
<< metal5 >>
rect -1590 40 4220 70
rect -1590 -210 80 40
rect 340 -70 4220 40
rect 340 -210 3930 -70
rect -1590 -250 3930 -210
rect 3900 -320 3930 -250
rect 4190 -320 4220 -70
rect 3900 -1400 4220 -320
rect 3900 -1650 3930 -1400
rect 4190 -1650 4220 -1400
rect 3900 -2720 4220 -1650
rect 3900 -2970 3930 -2720
rect 4190 -2970 4220 -2720
rect 3900 -3000 4220 -2970
use sky130_fd_sc_hd__or4_1  x1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712456748
transform 1 0 488 0 1 -811
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  x2
timestamp 1712456748
transform 1 0 1118 0 1 -811
box -38 -48 590 592
use sky130_fd_sc_hd__inv_1  x3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712456748
transform 1 0 -758 0 -1 442
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  x4 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712456748
transform 1 0 1748 0 1 -811
box -38 -48 498 592
use sky130_fd_sc_hd__inv_1  x5
timestamp 1712456748
transform 1 0 -1034 0 -1 442
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  x6
timestamp 1712456748
transform 1 0 -1308 0 -1 442
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  x7
timestamp 1712456748
transform 1 0 -1584 0 -1 442
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  x8 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712456748
transform 1 0 2288 0 1 -811
box -38 -48 498 592
use sky130_fd_sc_hd__inv_1  x9
timestamp 1712456748
transform 1 0 -482 0 -1 442
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  x10
timestamp 1712456748
transform 1 0 488 0 -1 -928
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  x11
timestamp 1712456748
transform 1 0 1028 0 -1 -928
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  x12
timestamp 1712456748
transform 1 0 1568 0 -1 -928
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  x13
timestamp 1712456748
transform 1 0 2108 0 -1 -928
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  x14
timestamp 1712456748
transform 1 0 2648 0 -1 -928
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  x15 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712456748
transform 1 0 488 0 1 -2132
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  x16
timestamp 1712456748
transform 1 0 1208 0 1 -2132
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  x17
timestamp 1712456748
transform 1 0 1928 0 1 -2132
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  x18
timestamp 1712456748
transform 1 0 488 0 -1 -2248
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  x19
timestamp 1712456748
transform 1 0 1208 0 -1 -2248
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  x20 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712456748
transform 1 0 1928 0 -1 -2248
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  x21
timestamp 1712456748
transform 1 0 2468 0 -1 -2248
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  x22
timestamp 1712456748
transform -1 0 3560 0 -1 -2248
box -38 -48 590 592
<< labels >>
flabel metal1 5540 -1470 5740 -1270 0 FreeSans 256 0 0 0 A1
port 11 nsew
flabel metal1 5540 -1070 5740 -870 0 FreeSans 256 0 0 0 A2
port 10 nsew
flabel metal1 5540 -270 5740 -70 0 FreeSans 256 0 0 0 EO
port 8 nsew
flabel metal1 5540 -670 5740 -470 0 FreeSans 256 0 0 0 GS
port 9 nsew
flabel metal1 -3910 490 -3710 690 0 FreeSans 256 0 0 0 I0
port 3 nsew
flabel metal1 -3660 490 -3460 690 0 FreeSans 256 0 0 0 I1
port 0 nsew
flabel metal1 -3410 490 -3210 690 0 FreeSans 256 0 0 0 I2
port 4 nsew
flabel metal1 -3160 490 -2960 690 0 FreeSans 256 0 0 0 I3
port 2 nsew
flabel metal1 -2910 490 -2710 690 0 FreeSans 256 0 0 0 I4
port 7 nsew
flabel metal1 -2660 490 -2460 690 0 FreeSans 256 0 0 0 I5
port 1 nsew
flabel metal1 -2410 490 -2210 690 0 FreeSans 256 0 0 0 I6
port 5 nsew
flabel metal1 -2160 490 -1960 690 0 FreeSans 256 0 0 0 I7
port 6 nsew
flabel metal1 -1910 490 -1710 690 0 FreeSans 256 0 0 0 EI
port 13 nsew
<< end >>
