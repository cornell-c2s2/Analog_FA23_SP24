magic
tech sky130A
timestamp 1713148681
<< end >>
