magic
tech sky130A
magscale 1 2
timestamp 1710185907
<< locali >>
rect 1250 -331 1450 -325
rect 1250 -369 1256 -331
rect 1294 -369 1406 -331
rect 1444 -369 1450 -331
rect 1250 -375 1450 -369
<< viali >>
rect 1707 -318 1744 -281
rect 1081 -369 1119 -331
rect 1256 -369 1294 -331
rect 1406 -369 1444 -331
rect 1855 -370 1895 -330
rect 2206 -368 2243 -331
rect 2531 -369 2569 -331
rect 2831 -369 2869 -331
rect 3151 -374 3199 -327
rect 3406 -369 3444 -331
rect 3556 -369 3594 -331
rect 3976 -374 4024 -327
rect 4231 -369 4269 -331
rect 4406 -369 4444 -331
rect 1051 -849 1099 -801
rect 1201 -924 1249 -876
rect 1355 -945 1395 -905
rect 1855 -945 1895 -905
rect 2555 -945 2595 -905
rect 2705 -945 2745 -905
rect 3006 -944 3044 -906
rect 3355 -945 3395 -905
rect 3556 -944 3594 -906
rect 3856 -969 3894 -931
rect 4026 -948 4074 -901
rect 4406 -944 4444 -906
rect 4655 -945 4695 -905
rect 4805 -945 4845 -905
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 1700 -250 2250 -200
rect 1700 -281 1750 -250
rect 1700 -318 1707 -281
rect 1744 -318 1750 -281
rect 1075 -331 1125 -319
rect 1700 -325 1750 -318
rect 1075 -369 1081 -331
rect 1119 -369 1125 -331
rect 1075 -425 1125 -369
rect 1244 -331 1456 -325
rect 1701 -330 1750 -325
rect 1244 -369 1256 -331
rect 1294 -369 1406 -331
rect 1444 -369 1456 -331
rect 1244 -375 1456 -369
rect 1843 -376 1849 -324
rect 1901 -376 1907 -324
rect 2200 -325 2250 -250
rect 3400 -275 4450 -225
rect 2693 -325 2699 -324
rect 2200 -331 2249 -325
rect 2200 -368 2206 -331
rect 2243 -368 2249 -331
rect 2200 -380 2249 -368
rect 2519 -331 2699 -325
rect 2519 -369 2531 -331
rect 2569 -369 2699 -331
rect 2519 -375 2699 -369
rect 2693 -376 2699 -375
rect 2751 -376 2757 -324
rect 2825 -331 2875 -319
rect 2825 -369 2831 -331
rect 2869 -369 2875 -331
rect 1343 -425 1349 -424
rect 1075 -475 1349 -425
rect 1343 -476 1349 -475
rect 1401 -476 1407 -424
rect 2543 -476 2549 -424
rect 2601 -425 2607 -424
rect 2825 -425 2875 -369
rect 3139 -380 3145 -320
rect 3205 -380 3211 -320
rect 3400 -331 3450 -275
rect 3400 -369 3406 -331
rect 3444 -369 3450 -331
rect 3400 -381 3450 -369
rect 3550 -331 3600 -319
rect 3550 -369 3556 -331
rect 3594 -369 3600 -331
rect 2601 -475 2875 -425
rect 2601 -476 2607 -475
rect 3343 -476 3349 -424
rect 3401 -425 3407 -424
rect 3550 -425 3600 -369
rect 3964 -380 3970 -320
rect 4030 -380 4036 -320
rect 4225 -331 4275 -319
rect 4225 -369 4231 -331
rect 4269 -369 4275 -331
rect 3401 -475 3600 -425
rect 4225 -425 4275 -369
rect 4400 -331 4450 -275
rect 4400 -369 4406 -331
rect 4444 -369 4450 -331
rect 4400 -381 4450 -369
rect 4799 -424 4851 -418
rect 4225 -475 4799 -425
rect 3401 -476 3407 -475
rect 4799 -482 4851 -476
rect 0 -800 200 -600
rect 1025 -795 1125 -775
rect 1025 -855 1045 -795
rect 1105 -855 1125 -795
rect 1025 -875 1125 -855
rect 3850 -850 4450 -800
rect 1189 -930 1195 -870
rect 1255 -930 1261 -870
rect 1343 -951 1349 -899
rect 1401 -951 1407 -899
rect 1843 -951 1849 -899
rect 1901 -951 1907 -899
rect 2543 -951 2549 -899
rect 2601 -951 2607 -899
rect 2693 -951 2699 -899
rect 2751 -951 2757 -899
rect 3000 -906 3050 -894
rect 3000 -944 3006 -906
rect 3044 -944 3050 -906
rect 2550 -1000 2600 -951
rect 3000 -1000 3050 -944
rect 3343 -951 3349 -899
rect 3401 -951 3407 -899
rect 3550 -906 3600 -894
rect 3550 -944 3556 -906
rect 3594 -944 3600 -906
rect 3550 -1000 3600 -944
rect 3850 -931 3900 -850
rect 3850 -969 3856 -931
rect 3894 -969 3900 -931
rect 4014 -955 4020 -895
rect 4080 -955 4086 -895
rect 4400 -906 4450 -850
rect 4400 -944 4406 -906
rect 4444 -944 4450 -906
rect 4400 -956 4450 -944
rect 4643 -951 4649 -899
rect 4701 -951 4707 -899
rect 4793 -951 4799 -899
rect 4851 -951 4857 -899
rect 3850 -981 3900 -969
rect 0 -1200 200 -1000
rect 2550 -1050 3600 -1000
rect 0 -1600 200 -1400
rect 0 -2000 200 -1800
<< via1 >>
rect 1849 -330 1901 -324
rect 1849 -370 1855 -330
rect 1855 -370 1895 -330
rect 1895 -370 1901 -330
rect 1849 -376 1901 -370
rect 2699 -376 2751 -324
rect 1349 -476 1401 -424
rect 2549 -476 2601 -424
rect 3145 -327 3205 -320
rect 3145 -374 3151 -327
rect 3151 -374 3199 -327
rect 3199 -374 3205 -327
rect 3145 -380 3205 -374
rect 3349 -476 3401 -424
rect 3970 -327 4030 -320
rect 3970 -374 3976 -327
rect 3976 -374 4024 -327
rect 4024 -374 4030 -327
rect 3970 -380 4030 -374
rect 4799 -476 4851 -424
rect 1045 -801 1105 -795
rect 1045 -849 1051 -801
rect 1051 -849 1099 -801
rect 1099 -849 1105 -801
rect 1045 -855 1105 -849
rect 1195 -876 1255 -870
rect 1195 -924 1201 -876
rect 1201 -924 1249 -876
rect 1249 -924 1255 -876
rect 1195 -930 1255 -924
rect 1349 -905 1401 -899
rect 1349 -945 1355 -905
rect 1355 -945 1395 -905
rect 1395 -945 1401 -905
rect 1349 -951 1401 -945
rect 1849 -905 1901 -899
rect 1849 -945 1855 -905
rect 1855 -945 1895 -905
rect 1895 -945 1901 -905
rect 1849 -951 1901 -945
rect 2549 -905 2601 -899
rect 2549 -945 2555 -905
rect 2555 -945 2595 -905
rect 2595 -945 2601 -905
rect 2549 -951 2601 -945
rect 2699 -905 2751 -899
rect 2699 -945 2705 -905
rect 2705 -945 2745 -905
rect 2745 -945 2751 -905
rect 2699 -951 2751 -945
rect 3349 -905 3401 -899
rect 3349 -945 3355 -905
rect 3355 -945 3395 -905
rect 3395 -945 3401 -905
rect 3349 -951 3401 -945
rect 4020 -901 4080 -895
rect 4020 -948 4026 -901
rect 4026 -948 4074 -901
rect 4074 -948 4080 -901
rect 4020 -955 4080 -948
rect 4649 -905 4701 -899
rect 4649 -945 4655 -905
rect 4655 -945 4695 -905
rect 4695 -945 4701 -905
rect 4649 -951 4701 -945
rect 4799 -905 4851 -899
rect 4799 -945 4805 -905
rect 4805 -945 4845 -905
rect 4845 -945 4851 -905
rect 4799 -951 4851 -945
<< metal2 >>
rect 1849 -324 1901 -318
rect 1849 -382 1901 -376
rect 2699 -324 2751 -318
rect 2699 -382 2751 -376
rect 3145 -320 3205 -314
rect 1350 -418 1425 -400
rect 1349 -424 1425 -418
rect 1401 -475 1425 -424
rect 1349 -482 1401 -476
rect 1025 -795 1125 -775
rect 1025 -855 1045 -795
rect 1105 -855 1125 -795
rect 1025 -875 1125 -855
rect 1195 -870 1255 -864
rect 1350 -893 1400 -482
rect 1850 -786 1900 -382
rect 2549 -424 2601 -418
rect 2549 -482 2601 -476
rect 1845 -795 1905 -786
rect 1845 -864 1905 -855
rect 1850 -893 1900 -864
rect 2550 -893 2600 -482
rect 2700 -893 2750 -382
rect 1195 -967 1255 -930
rect 1349 -899 1401 -893
rect 1349 -957 1401 -951
rect 1849 -899 1901 -893
rect 1849 -957 1901 -951
rect 2549 -899 2601 -893
rect 2549 -957 2601 -951
rect 2699 -899 2751 -893
rect 2699 -957 2751 -951
rect 3145 -967 3205 -380
rect 3970 -320 4030 -314
rect 3349 -424 3401 -418
rect 3349 -482 3401 -476
rect 3350 -893 3400 -482
rect 3970 -522 4030 -380
rect 4793 -476 4799 -424
rect 4851 -476 4857 -424
rect 4645 -520 4705 -511
rect 3963 -578 3972 -522
rect 4028 -578 4037 -522
rect 3970 -580 4030 -578
rect 4645 -589 4705 -580
rect 3349 -899 3401 -893
rect 3349 -957 3401 -951
rect 4020 -895 4080 -889
rect 4650 -893 4700 -589
rect 4800 -893 4850 -476
rect 4020 -967 4080 -955
rect 4649 -899 4701 -893
rect 4649 -957 4701 -951
rect 4799 -899 4851 -893
rect 4799 -957 4851 -951
rect 1195 -1023 1197 -967
rect 1253 -1023 1255 -967
rect 3138 -1023 3147 -967
rect 3203 -1023 3212 -967
rect 4020 -1023 4022 -967
rect 4078 -1023 4080 -967
rect 1195 -1025 1255 -1023
rect 3145 -1025 3205 -1023
rect 4020 -1025 4080 -1023
rect 1197 -1032 1253 -1025
rect 4022 -1032 4078 -1025
<< via2 >>
rect 1047 -853 1103 -797
rect 1845 -855 1905 -795
rect 3972 -578 4028 -522
rect 4645 -580 4705 -520
rect 1197 -1023 1253 -967
rect 3147 -1023 3203 -967
rect 4022 -1023 4078 -967
<< metal3 >>
rect 3967 -520 4033 -517
rect 4640 -520 4710 -515
rect 3967 -522 4645 -520
rect 3967 -578 3972 -522
rect 4028 -578 4645 -522
rect 3967 -580 4645 -578
rect 4705 -580 4710 -520
rect 3967 -583 4033 -580
rect 4640 -585 4710 -580
rect 1025 -795 1125 -775
rect 1840 -795 1910 -790
rect 1025 -797 1845 -795
rect 1025 -853 1047 -797
rect 1103 -853 1845 -797
rect 1025 -855 1845 -853
rect 1905 -855 1910 -795
rect 1025 -875 1125 -855
rect 1840 -860 1910 -855
rect 1192 -965 1258 -962
rect 3142 -965 3208 -962
rect 4017 -965 4083 -962
rect 1192 -967 4083 -965
rect 1192 -1023 1197 -967
rect 1253 -1023 3147 -967
rect 3203 -1023 4022 -967
rect 4078 -1023 4083 -967
rect 1192 -1025 4083 -1023
rect 1192 -1028 1258 -1025
rect 3142 -1028 3208 -1025
rect 4017 -1028 4083 -1025
use sky130_fd_sc_hd__nand2_4  x3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform -1 0 2974 0 1 -592
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  x4
timestamp 1701704242
transform 1 0 2142 0 -1 -683
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  x5
timestamp 1701704242
transform -1 0 2146 0 1 -592
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  x6
timestamp 1701704242
transform 1 0 1314 0 -1 -683
box -38 -48 866 592
use sky130_fd_sc_hd__inv_4  x8 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 858 0 1 -592
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_4  x9
timestamp 1701704242
transform 1 0 3802 0 1 -592
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  x10
timestamp 1701704242
transform 1 0 4258 0 -1 -683
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  x11
timestamp 1701704242
transform 1 0 2974 0 1 -592
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  x12
timestamp 1701704242
transform 1 0 3430 0 -1 -683
box -38 -48 866 592
use sky130_fd_sc_hd__inv_4  x13
timestamp 1701704242
transform 1 0 2970 0 -1 -683
box -38 -48 498 592
use sky130_fd_sc_hd__clkinv_1  x14 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 1038 0 -1 -683
box -38 -48 314 592
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 VDD
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 SIG
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 OUT
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 CLK
port 3 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 256 0 0 0 VSS
port 4 nsew
flabel metal1 0 -2000 200 -1800 0 FreeSans 256 0 0 0 VMID
port 5 nsew
<< end >>
