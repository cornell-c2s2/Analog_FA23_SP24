* NGSPICE file created from resistorDivider_v0p0p1.ext - technology: sky130A

.subckt sky130_fd_pr__res_xhigh_po_5p73_QJNTVE a_2532_252# a_n1194_n684# a_n1194_252#
+ a_n5050_n814# a_n4920_n684# a_n2436_252# a_n2436_n684# a_48_252# a_n3678_n684# a_1290_n684#
+ a_3774_252# a_48_n684# a_2532_n684# a_1290_252# a_n3678_252# a_3774_n684# a_n4920_252#
X0 a_n2436_252# a_n2436_n684# a_n5050_n814# sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1 a_1290_252# a_1290_n684# a_n5050_n814# sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X2 a_48_252# a_48_n684# a_n5050_n814# sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X3 a_n4920_252# a_n4920_n684# a_n5050_n814# sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X4 a_3774_252# a_3774_n684# a_n5050_n814# sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X5 a_n1194_252# a_n1194_n684# a_n5050_n814# sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X6 a_2532_252# a_2532_n684# a_n5050_n814# sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X7 a_n3678_252# a_n3678_n684# a_n5050_n814# sky130_fd_pr__res_xhigh_po_5p73 l=2.52
.ends

.subckt sky130_fd_pr__res_xhigh_po_5p73_7KNTDX a_2532_252# a_n1194_n684# a_n1194_252#
+ a_n5050_n814# a_n4920_n684# a_n2436_252# a_n2436_n684# a_48_252# a_n3678_n684# a_1290_n684#
+ a_3774_252# a_48_n684# a_2532_n684# a_1290_252# a_n3678_252# a_3774_n684# a_n4920_252#
X0 a_n2436_252# a_n2436_n684# a_n5050_n814# sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1 a_1290_252# a_1290_n684# a_n5050_n814# sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X2 a_48_252# a_48_n684# a_n5050_n814# sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X3 a_n4920_252# a_n4920_n684# a_n5050_n814# sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X4 a_3774_252# a_3774_n684# a_n5050_n814# sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X5 a_n1194_252# a_n1194_n684# a_n5050_n814# sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X6 a_2532_252# a_2532_n684# a_n5050_n814# sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X7 a_n3678_252# a_n3678_n684# a_n5050_n814# sky130_fd_pr__res_xhigh_po_5p73 l=2.52
.ends

.subckt resistorDivider_v0p0p1 VL VFS V1 V2 V3 V4 V5 V6 V7 V8 V9 V10 V11 V12 V13 V14
+ V15 V16
XXR1 VL V1 VL VL V1 VL V1 VL V1 V1 VL V1 V1 VL VL V1 VL sky130_fd_pr__res_xhigh_po_5p73_QJNTVE
XXR10 V9 V10 V9 VL V10 V9 V10 V9 V10 V10 V9 V10 V10 V9 V9 V10 V9 sky130_fd_pr__res_xhigh_po_5p73_7KNTDX
XXR2 V1 V2 V1 VL V2 V1 V2 V1 V2 V2 V1 V2 V2 V1 V1 V2 V1 sky130_fd_pr__res_xhigh_po_5p73_7KNTDX
XXR11 V10 V11 V10 VL V11 V10 V11 V10 V11 V11 V10 V11 V11 V10 V10 V11 V10 sky130_fd_pr__res_xhigh_po_5p73_7KNTDX
XXR3 V2 V3 V2 VL V3 V2 V3 V2 V3 V3 V2 V3 V3 V2 V2 V3 V2 sky130_fd_pr__res_xhigh_po_5p73_7KNTDX
XXR12 V11 V12 V11 VL V12 V11 V12 V11 V12 V12 V11 V12 V12 V11 V11 V12 V11 sky130_fd_pr__res_xhigh_po_5p73_7KNTDX
XXR5 V4 V5 V4 VL V5 V4 V5 V4 V5 V5 V4 V5 V5 V4 V4 V5 V4 sky130_fd_pr__res_xhigh_po_5p73_7KNTDX
XXR4 V3 V4 V3 VL V4 V3 V4 V3 V4 V4 V3 V4 V4 V3 V3 V4 V3 sky130_fd_pr__res_xhigh_po_5p73_7KNTDX
XXR14 V13 V14 V13 VL V14 V13 V14 V13 V14 V14 V13 V14 V14 V13 V13 V14 V13 sky130_fd_pr__res_xhigh_po_5p73_7KNTDX
XXR13 V12 V13 V12 VL V13 V12 V13 V12 V13 V13 V12 V13 V13 V12 V12 V13 V12 sky130_fd_pr__res_xhigh_po_5p73_7KNTDX
XXR6 V5 V6 V5 VL V6 V5 V6 V5 V6 V6 V5 V6 V6 V5 V5 V6 V5 sky130_fd_pr__res_xhigh_po_5p73_7KNTDX
XXR15 V14 V15 V14 VL V15 V14 V15 V14 V15 V15 V14 V15 V15 V14 V14 V15 V14 sky130_fd_pr__res_xhigh_po_5p73_7KNTDX
XXR7 V6 V7 V6 VL V7 V6 V7 V6 V7 V7 V6 V7 V7 V6 V6 V7 V6 sky130_fd_pr__res_xhigh_po_5p73_7KNTDX
XXR16 V15 V16 V15 VL V16 V15 V16 V15 V16 V16 V15 V16 V16 V15 V15 V16 V15 sky130_fd_pr__res_xhigh_po_5p73_7KNTDX
XXR8 V7 V8 V7 VL V8 V7 V8 V7 V8 V8 V7 V8 V8 V7 V7 V8 V7 sky130_fd_pr__res_xhigh_po_5p73_7KNTDX
XXR17 V16 VFS V16 VL VFS V16 VFS V16 VFS VFS V16 VFS VFS V16 V16 VFS V16 sky130_fd_pr__res_xhigh_po_5p73_7KNTDX
XXR9 V8 V9 V8 VL V9 V8 V9 V8 V9 V9 V8 V9 V9 V8 V8 V9 V8 sky130_fd_pr__res_xhigh_po_5p73_7KNTDX
.ends

