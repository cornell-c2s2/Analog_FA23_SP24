magic
tech sky130A
magscale 1 2
timestamp 1714790421
<< pwell >>
rect -5086 -867 5086 867
<< psubdiff >>
rect -5050 797 -4954 831
rect 4954 797 5050 831
rect -5050 735 -5016 797
rect 5016 735 5050 797
rect -5050 -797 -5016 -735
rect 5016 -797 5050 -735
rect -5050 -831 -4954 -797
rect 4954 -831 5050 -797
<< psubdiffcont >>
rect -4954 797 4954 831
rect -5050 -735 -5016 735
rect 5016 -735 5050 735
rect -4954 -831 4954 -797
<< xpolycontact >>
rect -4920 269 -3774 701
rect -4920 -701 -3774 -269
rect -3678 269 -2532 701
rect -3678 -701 -2532 -269
rect -2436 269 -1290 701
rect -2436 -701 -1290 -269
rect -1194 269 -48 701
rect -1194 -701 -48 -269
rect 48 269 1194 701
rect 48 -701 1194 -269
rect 1290 269 2436 701
rect 1290 -701 2436 -269
rect 2532 269 3678 701
rect 2532 -701 3678 -269
rect 3774 269 4920 701
rect 3774 -701 4920 -269
<< xpolyres >>
rect -4920 -269 -3774 269
rect -3678 -269 -2532 269
rect -2436 -269 -1290 269
rect -1194 -269 -48 269
rect 48 -269 1194 269
rect 1290 -269 2436 269
rect 2532 -269 3678 269
rect 3774 -269 4920 269
<< locali >>
rect -5050 797 -4954 831
rect 4954 797 5050 831
rect -5050 735 -5016 797
rect 5016 735 5050 797
rect -5050 -797 -5016 -735
rect 5016 -797 5050 -735
rect -5050 -831 -4954 -797
rect 4954 -831 5050 -797
<< viali >>
rect -4904 286 -3790 683
rect -3662 286 -2548 683
rect -2420 286 -1306 683
rect -1178 286 -64 683
rect 64 286 1178 683
rect 1306 286 2420 683
rect 2548 286 3662 683
rect 3790 286 4904 683
rect -4904 -683 -3790 -286
rect -3662 -683 -2548 -286
rect -2420 -683 -1306 -286
rect -1178 -683 -64 -286
rect 64 -683 1178 -286
rect 1306 -683 2420 -286
rect 2548 -683 3662 -286
rect 3790 -683 4904 -286
<< metal1 >>
rect -4916 683 -3778 689
rect -4916 286 -4904 683
rect -3790 286 -3778 683
rect -4916 280 -3778 286
rect -3674 683 -2536 689
rect -3674 286 -3662 683
rect -2548 286 -2536 683
rect -3674 280 -2536 286
rect -2432 683 -1294 689
rect -2432 286 -2420 683
rect -1306 286 -1294 683
rect -2432 280 -1294 286
rect -1190 683 -52 689
rect -1190 286 -1178 683
rect -64 286 -52 683
rect -1190 280 -52 286
rect 52 683 1190 689
rect 52 286 64 683
rect 1178 286 1190 683
rect 52 280 1190 286
rect 1294 683 2432 689
rect 1294 286 1306 683
rect 2420 286 2432 683
rect 1294 280 2432 286
rect 2536 683 3674 689
rect 2536 286 2548 683
rect 3662 286 3674 683
rect 2536 280 3674 286
rect 3778 683 4916 689
rect 3778 286 3790 683
rect 4904 286 4916 683
rect 3778 280 4916 286
rect -4916 -286 -3778 -280
rect -4916 -683 -4904 -286
rect -3790 -683 -3778 -286
rect -4916 -689 -3778 -683
rect -3674 -286 -2536 -280
rect -3674 -683 -3662 -286
rect -2548 -683 -2536 -286
rect -3674 -689 -2536 -683
rect -2432 -286 -1294 -280
rect -2432 -683 -2420 -286
rect -1306 -683 -1294 -286
rect -2432 -689 -1294 -683
rect -1190 -286 -52 -280
rect -1190 -683 -1178 -286
rect -64 -683 -52 -286
rect -1190 -689 -52 -683
rect 52 -286 1190 -280
rect 52 -683 64 -286
rect 1178 -683 1190 -286
rect 52 -689 1190 -683
rect 1294 -286 2432 -280
rect 1294 -683 1306 -286
rect 2420 -683 2432 -286
rect 1294 -689 2432 -683
rect 2536 -286 3674 -280
rect 2536 -683 2548 -286
rect 3662 -683 3674 -286
rect 2536 -689 3674 -683
rect 3778 -286 4916 -280
rect 3778 -683 3790 -286
rect 4904 -683 4916 -286
rect 3778 -689 4916 -683
<< properties >>
string FIXED_BBOX -5033 -814 5033 814
string gencell sky130_fd_pr__res_xhigh_po_5p73
string library sky130
string parameters w 5.73 l 2.852 m 1 nx 8 wmin 5.730 lmin 0.50 rho 2000 val 1.061k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 5.730 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
