magic
tech sky130A
magscale 1 2
timestamp 1717179484
<< nwell >>
rect 202 -452 984 -208
rect 380 -870 390 -452
rect 450 -870 470 -850
rect 490 -870 560 -452
rect 860 -560 1260 -470
rect 1740 -550 1990 -480
rect 380 -920 560 -870
rect 380 -930 390 -920
rect 450 -930 470 -920
rect 2290 -930 2390 -900
rect 2400 -920 2460 -860
rect 2480 -930 2490 -860
rect 1600 -1860 1680 -1790
rect 1710 -2030 1870 -1720
rect 1190 -2050 1870 -2030
rect 1721 -2070 1870 -2050
rect 1720 -2280 1870 -2070
rect 1190 -2350 1250 -2340
rect 1721 -2350 1870 -2280
rect 1190 -2370 1870 -2350
<< pwell >>
rect 910 -700 1410 -670
rect 1920 -700 1970 -690
rect 870 -760 1410 -700
rect 870 -1050 940 -760
rect 960 -900 1040 -840
rect 1150 -850 1220 -790
rect 950 -1050 1040 -900
rect 1370 -910 1380 -830
rect 1470 -940 1560 -770
rect 1580 -860 1790 -780
rect 1800 -920 1890 -820
rect 520 -1110 1040 -1050
rect 1910 -1070 1970 -700
rect 520 -1140 530 -1110
rect 540 -1130 610 -1110
rect 540 -1140 890 -1130
rect 930 -1140 940 -1110
rect 1910 -1140 2310 -1070
rect 430 -1260 890 -1140
rect 430 -1290 610 -1260
rect 520 -1870 530 -1290
rect 540 -1850 610 -1290
rect 1050 -1340 1380 -1220
rect 1580 -1340 1790 -1220
rect 1830 -1230 1880 -1220
rect 1670 -1590 1920 -1510
rect 710 -1870 790 -1700
rect 2240 -1850 2310 -1140
rect 1060 -2450 1250 -2420
rect 1060 -2680 1260 -2450
rect 1080 -2690 1260 -2680
rect 1080 -2700 1200 -2690
<< ndiff >>
rect 1150 -850 1220 -790
<< psubdiff >>
rect 1090 -2530 1190 -2500
rect 1090 -2600 1120 -2530
rect 1100 -2650 1120 -2600
rect 1160 -2600 1190 -2530
rect 1160 -2650 1180 -2600
rect 1100 -2680 1180 -2650
<< nsubdiff >>
rect 1730 -1800 1830 -1780
rect 1730 -1840 1760 -1800
rect 1800 -1840 1830 -1800
rect 1730 -1860 1830 -1840
rect 1730 -1940 1830 -1920
rect 1730 -1980 1760 -1940
rect 1800 -1980 1830 -1940
rect 1730 -2000 1830 -1980
rect 1730 -2080 1830 -2060
rect 1730 -2120 1760 -2080
rect 1800 -2120 1830 -2080
rect 1730 -2140 1830 -2120
rect 1730 -2220 1830 -2200
rect 1730 -2260 1760 -2220
rect 1800 -2260 1830 -2220
rect 1730 -2280 1830 -2260
<< psubdiffcont >>
rect 1120 -2650 1160 -2530
<< nsubdiffcont >>
rect 1760 -1840 1800 -1800
rect 1760 -1980 1800 -1940
rect 1760 -2120 1800 -2080
rect 1760 -2260 1800 -2220
<< poly >>
rect 1480 -910 1530 -840
<< locali >>
rect 310 -280 320 -240
rect 620 -280 640 -240
rect 1740 -1800 1820 -1780
rect 1740 -1840 1760 -1800
rect 1800 -1840 1820 -1800
rect 1740 -1860 1820 -1840
rect 1740 -1940 1820 -1920
rect 1740 -1980 1760 -1940
rect 1800 -1980 1820 -1940
rect 1740 -2000 1820 -1980
rect 1740 -2080 1820 -2060
rect 1740 -2120 1760 -2080
rect 1800 -2120 1820 -2080
rect 1740 -2140 1820 -2120
rect 1740 -2220 1820 -2200
rect 1740 -2260 1760 -2220
rect 1800 -2260 1820 -2220
rect 1740 -2280 1820 -2260
rect 1090 -2510 1190 -2500
rect 1090 -2600 1100 -2510
rect 1180 -2600 1190 -2510
<< viali >>
rect 320 -280 620 -240
rect 860 -280 1990 -240
rect 2210 -280 2600 -240
rect 990 -740 1350 -700
rect 1500 -740 1870 -700
rect 890 -970 930 -790
rect 1920 -960 1960 -790
rect 330 -1010 620 -970
rect 2230 -1020 2530 -970
rect 650 -1120 840 -1080
rect 2020 -1120 2200 -1080
rect 560 -1740 600 -1180
rect 1625 -1645 1659 -1611
rect 1260 -1720 1300 -1680
rect 1350 -1720 1390 -1680
rect 1440 -1720 1480 -1680
rect 1520 -1720 1560 -1680
rect 1625 -1719 1659 -1683
rect 2260 -1740 2300 -1180
rect 1625 -1798 1659 -1763
rect 1760 -1840 1800 -1800
rect 1760 -1980 1800 -1940
rect 1760 -2120 1800 -2080
rect 1760 -2260 1800 -2220
rect 1625 -2329 1659 -2294
rect 1260 -2400 1300 -2360
rect 1350 -2400 1390 -2360
rect 1440 -2400 1480 -2360
rect 1520 -2400 1560 -2360
rect 1625 -2402 1659 -2367
rect 1624 -2478 1658 -2443
rect 1100 -2530 1180 -2510
rect 1100 -2650 1120 -2530
rect 1120 -2650 1160 -2530
rect 1160 -2650 1180 -2530
rect 1100 -2680 1180 -2650
<< metal1 >>
rect 1360 110 1560 130
rect 1360 -50 1380 110
rect 1540 -50 1560 110
rect 1360 -70 1560 -50
rect -350 -280 -50 -90
rect 692 -210 786 -208
rect -350 -440 -230 -280
rect -70 -440 -50 -280
rect 250 -220 2620 -210
rect 250 -280 270 -220
rect 330 -240 630 -220
rect 620 -280 630 -240
rect 690 -240 2530 -220
rect 690 -280 860 -240
rect 1990 -280 2160 -240
rect 250 -300 2160 -280
rect 2230 -300 2530 -280
rect 2600 -300 2620 -220
rect 2880 -300 3190 -120
rect 692 -302 786 -300
rect 490 -390 500 -330
rect 560 -390 570 -330
rect 850 -350 2000 -300
rect 730 -390 820 -380
rect 850 -390 1270 -350
rect -350 -620 -50 -440
rect 260 -530 380 -420
rect 260 -590 270 -530
rect 330 -590 380 -530
rect 570 -530 700 -430
rect 730 -480 740 -390
rect 810 -480 820 -390
rect 860 -400 1270 -390
rect 1300 -390 1390 -380
rect 730 -490 820 -480
rect 860 -490 1260 -470
rect 1300 -480 1310 -390
rect 1380 -480 1390 -390
rect 1300 -490 1390 -480
rect 1460 -390 1550 -380
rect 1460 -480 1470 -390
rect 1540 -480 1550 -390
rect 1580 -400 2000 -350
rect 2030 -390 2110 -380
rect 2380 -390 2400 -330
rect 2460 -390 2490 -330
rect 1460 -490 1550 -480
rect 1590 -480 1990 -470
rect 570 -590 620 -530
rect 680 -590 700 -530
rect 860 -550 940 -490
rect 1020 -550 1140 -490
rect 1220 -520 1260 -490
rect 1220 -550 1470 -520
rect 860 -570 1470 -550
rect 1460 -580 1470 -570
rect 1540 -580 1550 -520
rect 1590 -540 1630 -480
rect 1710 -540 1860 -480
rect 1940 -540 1990 -480
rect 2030 -480 2040 -390
rect 2100 -480 2110 -390
rect 2030 -490 2110 -480
rect 2140 -460 2280 -430
rect 1590 -550 1990 -540
rect 2140 -540 2160 -460
rect 2230 -540 2280 -460
rect 260 -640 380 -590
rect 260 -700 270 -640
rect 330 -700 380 -640
rect 420 -600 500 -590
rect 420 -660 430 -600
rect 490 -660 500 -600
rect 420 -670 500 -660
rect 570 -650 700 -590
rect 260 -750 380 -700
rect 260 -810 270 -750
rect 330 -810 380 -750
rect 260 -830 380 -810
rect 570 -710 620 -650
rect 680 -710 700 -650
rect 2140 -590 2280 -540
rect 2480 -460 2620 -430
rect 2480 -540 2530 -460
rect 2600 -540 2620 -460
rect 2140 -670 2160 -590
rect 2230 -670 2280 -590
rect 570 -750 700 -710
rect 570 -810 620 -750
rect 680 -810 700 -750
rect 570 -820 700 -810
rect 600 -830 700 -820
rect 870 -700 1970 -690
rect 870 -740 990 -700
rect 1350 -740 1500 -700
rect 1870 -740 1970 -700
rect 870 -750 1970 -740
rect 870 -790 940 -750
rect 380 -920 390 -860
rect 450 -920 460 -860
rect 380 -930 460 -920
rect 500 -920 510 -860
rect 570 -920 580 -860
rect 500 -930 580 -920
rect 230 -950 340 -940
rect 230 -1010 270 -950
rect 330 -960 340 -950
rect 610 -960 630 -950
rect 330 -970 630 -960
rect 620 -1010 630 -970
rect 690 -1010 710 -950
rect 230 -1020 710 -1010
rect 870 -970 890 -790
rect 930 -970 940 -790
rect 870 -1070 940 -970
rect 970 -890 1040 -840
rect 1070 -850 1150 -790
rect 1220 -850 1270 -790
rect 1070 -860 1270 -850
rect 1030 -950 1040 -890
rect 1070 -950 1090 -890
rect 1260 -950 1270 -890
rect 970 -980 1040 -950
rect 1310 -980 1380 -830
rect 970 -1020 1380 -980
rect 1470 -990 1550 -830
rect 1580 -840 1630 -780
rect 1710 -840 1780 -780
rect 1910 -790 1970 -750
rect 1580 -860 1780 -840
rect 1820 -830 1880 -820
rect 1580 -960 1610 -900
rect 1750 -960 1780 -900
rect 1820 -990 1880 -910
rect 1470 -1020 1880 -990
rect 1910 -960 1920 -790
rect 1960 -960 1970 -790
rect 2140 -710 2280 -670
rect 2330 -570 2400 -560
rect 2390 -680 2400 -570
rect 2480 -590 2620 -540
rect 2480 -600 2530 -590
rect 2500 -670 2530 -600
rect 2600 -670 2620 -590
rect 2880 -440 2920 -300
rect 3060 -440 3190 -300
rect 2880 -670 3190 -440
rect 2330 -690 2400 -680
rect 2140 -790 2160 -710
rect 2230 -790 2280 -710
rect 2140 -820 2280 -790
rect 2480 -710 2620 -670
rect 2480 -790 2530 -710
rect 2600 -790 2620 -710
rect 2480 -820 2620 -790
rect 2510 -830 2620 -820
rect 2290 -920 2300 -860
rect 2360 -920 2370 -860
rect 2290 -930 2370 -920
rect 540 -1080 940 -1070
rect 540 -1120 650 -1080
rect 840 -1120 940 -1080
rect 540 -1140 940 -1120
rect 970 -1090 1390 -1060
rect 540 -1170 610 -1140
rect 430 -1180 610 -1170
rect -300 -1270 -10 -1260
rect -300 -1480 -200 -1270
rect -40 -1480 -10 -1270
rect 430 -1280 440 -1180
rect 530 -1280 560 -1180
rect 430 -1290 560 -1280
rect -300 -1700 -10 -1480
rect 540 -1740 560 -1290
rect 600 -1740 610 -1180
rect 700 -1230 710 -1170
rect 780 -1230 790 -1170
rect 970 -1250 1040 -1090
rect 1070 -1180 1100 -1120
rect 1240 -1180 1270 -1120
rect 1300 -1140 1390 -1090
rect 1070 -1230 1270 -1220
rect 640 -1360 710 -1270
rect 700 -1440 710 -1360
rect 640 -1450 710 -1440
rect 790 -1290 860 -1280
rect 640 -1650 700 -1450
rect 790 -1630 800 -1290
rect 852 -1630 860 -1290
rect 1070 -1320 1080 -1230
rect 1260 -1320 1270 -1230
rect 1300 -1230 1310 -1140
rect 1380 -1230 1390 -1140
rect 1300 -1240 1390 -1230
rect 1460 -1080 1880 -1050
rect 1460 -1140 1550 -1080
rect 1460 -1240 1470 -1140
rect 1540 -1240 1550 -1140
rect 1580 -1170 1590 -1110
rect 1770 -1170 1780 -1110
rect 1460 -1250 1550 -1240
rect 1590 -1230 1780 -1220
rect 1070 -1330 1270 -1320
rect 1820 -1240 1880 -1080
rect 1910 -1070 1970 -960
rect 2140 -1020 2160 -960
rect 2220 -970 2540 -960
rect 2220 -1020 2230 -970
rect 2530 -1020 2540 -970
rect 2600 -1020 2620 -960
rect 2140 -1030 2620 -1020
rect 1910 -1080 2310 -1070
rect 1910 -1120 2020 -1080
rect 2200 -1110 2310 -1080
rect 2200 -1120 2430 -1110
rect 1910 -1140 2310 -1120
rect 2070 -1230 2080 -1170
rect 2140 -1230 2160 -1170
rect 2240 -1180 2310 -1140
rect 2240 -1260 2260 -1180
rect 1590 -1330 1780 -1320
rect 2010 -1280 2090 -1270
rect 1220 -1410 1690 -1390
rect 1220 -1490 1380 -1410
rect 1540 -1490 1690 -1410
rect 1220 -1510 1690 -1490
rect 790 -1640 860 -1630
rect 1040 -1620 1200 -1600
rect 540 -1750 610 -1740
rect 420 -1760 610 -1750
rect 710 -1760 720 -1690
rect 780 -1760 790 -1690
rect 520 -1840 610 -1760
rect 1040 -1770 1050 -1620
rect 1190 -1650 1200 -1620
rect 1600 -1611 1680 -1590
rect 1600 -1645 1625 -1611
rect 1659 -1645 1680 -1611
rect 1190 -1660 1300 -1650
rect 1190 -1680 1570 -1660
rect 1190 -1720 1260 -1680
rect 1300 -1720 1350 -1680
rect 1390 -1720 1440 -1680
rect 1480 -1720 1520 -1680
rect 1560 -1720 1570 -1680
rect 1190 -1740 1570 -1720
rect 1600 -1683 1680 -1645
rect 2010 -1640 2020 -1280
rect 2080 -1640 2090 -1280
rect 2010 -1650 2090 -1640
rect 2150 -1650 2260 -1260
rect 1600 -1719 1625 -1683
rect 1659 -1719 1680 -1683
rect 1190 -1760 1300 -1740
rect 1190 -1770 1200 -1760
rect 1040 -1790 1200 -1770
rect 1600 -1763 1680 -1719
rect 2060 -1750 2080 -1690
rect 2140 -1750 2160 -1690
rect 2240 -1740 2260 -1650
rect 2300 -1230 2310 -1180
rect 2420 -1230 2430 -1120
rect 2300 -1240 2430 -1230
rect 2300 -1740 2310 -1240
rect 2880 -1310 3210 -1160
rect 2880 -1420 2890 -1310
rect 3000 -1420 3210 -1310
rect 2880 -1570 3210 -1420
rect 2240 -1750 2310 -1740
rect 1600 -1790 1625 -1763
rect 1659 -1790 1680 -1763
rect 2240 -1760 2460 -1750
rect 420 -1850 610 -1840
rect 1600 -1850 1610 -1790
rect 1670 -1850 1680 -1790
rect 1600 -1860 1680 -1850
rect 1740 -1790 1820 -1780
rect 1740 -1850 1750 -1790
rect 1810 -1850 1820 -1790
rect 2240 -1840 2330 -1760
rect 2450 -1840 2460 -1760
rect 2240 -1850 2460 -1840
rect 1740 -1860 1820 -1850
rect 1740 -1930 1820 -1920
rect 1740 -1950 1750 -1930
rect 1220 -2050 1750 -1950
rect 1810 -1950 1820 -1930
rect 1810 -2050 1870 -1950
rect 1220 -2070 1870 -2050
rect 1220 -2130 1750 -2070
rect 1810 -2130 1870 -2070
rect 1740 -2140 1820 -2130
rect 1740 -2210 1820 -2200
rect 1740 -2270 1750 -2210
rect 1810 -2270 1820 -2210
rect 1740 -2280 1820 -2270
rect 1610 -2294 1690 -2280
rect 1610 -2329 1625 -2294
rect 1659 -2329 1690 -2294
rect 1110 -2350 1580 -2340
rect 810 -2520 1040 -2350
rect 1110 -2440 1120 -2350
rect 1230 -2360 1580 -2350
rect 1230 -2400 1260 -2360
rect 1300 -2400 1350 -2360
rect 1390 -2400 1440 -2360
rect 1480 -2400 1520 -2360
rect 1560 -2400 1580 -2360
rect 1230 -2440 1580 -2400
rect 1110 -2450 1580 -2440
rect 1610 -2367 1690 -2329
rect 1610 -2402 1625 -2367
rect 1659 -2370 1690 -2367
rect 1659 -2402 2040 -2370
rect 1610 -2440 2040 -2402
rect 2140 -2440 2170 -2370
rect 1610 -2443 2170 -2440
rect 1610 -2478 1624 -2443
rect 1658 -2478 2170 -2443
rect 1610 -2490 2170 -2478
rect 810 -2660 820 -2520
rect 1000 -2660 1040 -2520
rect 810 -2780 1040 -2660
rect 1080 -2510 1200 -2490
rect 1610 -2491 1690 -2490
rect 1080 -2680 1100 -2510
rect 1180 -2570 1200 -2510
rect 1180 -2590 1690 -2570
rect 1180 -2670 1350 -2590
rect 1560 -2670 1690 -2590
rect 1180 -2680 1690 -2670
rect 1080 -2700 1200 -2680
<< via1 >>
rect 1380 -50 1540 110
rect -230 -440 -70 -280
rect 270 -240 330 -220
rect 270 -280 320 -240
rect 320 -280 330 -240
rect 630 -280 690 -220
rect 2530 -240 2600 -220
rect 2160 -280 2210 -240
rect 2210 -280 2230 -240
rect 2530 -280 2600 -240
rect 2160 -300 2230 -280
rect 2530 -300 2600 -280
rect 500 -390 560 -330
rect 270 -590 330 -530
rect 740 -480 810 -390
rect 1310 -480 1380 -390
rect 1470 -480 1540 -390
rect 2400 -390 2460 -330
rect 620 -590 680 -530
rect 940 -550 1020 -490
rect 1140 -550 1220 -490
rect 1470 -580 1540 -520
rect 1630 -540 1710 -480
rect 1860 -540 1940 -480
rect 2040 -480 2100 -390
rect 2160 -540 2230 -460
rect 270 -700 330 -640
rect 430 -660 490 -600
rect 270 -810 330 -750
rect 620 -710 680 -650
rect 2530 -540 2600 -460
rect 2160 -670 2230 -590
rect 620 -810 680 -750
rect 390 -920 450 -860
rect 510 -920 570 -860
rect 270 -1010 330 -950
rect 630 -1010 690 -950
rect 1150 -850 1220 -790
rect 970 -950 1030 -890
rect 1090 -950 1260 -890
rect 1630 -840 1710 -780
rect 1610 -960 1750 -900
rect 1820 -910 1880 -830
rect 2330 -680 2390 -570
rect 2530 -670 2600 -590
rect 2920 -440 3060 -300
rect 2160 -790 2230 -710
rect 2530 -790 2600 -710
rect 2300 -920 2360 -860
rect -200 -1480 -40 -1270
rect 440 -1280 530 -1180
rect 710 -1230 780 -1170
rect 1100 -1180 1240 -1120
rect 640 -1440 700 -1360
rect 800 -1630 852 -1290
rect 1080 -1320 1260 -1230
rect 1310 -1230 1380 -1140
rect 1470 -1240 1540 -1140
rect 1590 -1170 1770 -1110
rect 1590 -1320 1780 -1230
rect 2160 -1020 2220 -960
rect 2540 -1020 2600 -960
rect 2080 -1230 2140 -1170
rect 1380 -1490 1540 -1410
rect 720 -1760 780 -1690
rect 420 -1840 520 -1760
rect 1050 -1770 1190 -1620
rect 2020 -1640 2080 -1280
rect 2080 -1750 2140 -1690
rect 2310 -1230 2420 -1120
rect 2890 -1420 3000 -1310
rect 1610 -1798 1625 -1790
rect 1625 -1798 1659 -1790
rect 1659 -1798 1670 -1790
rect 1610 -1850 1670 -1798
rect 1750 -1800 1810 -1790
rect 1750 -1840 1760 -1800
rect 1760 -1840 1800 -1800
rect 1800 -1840 1810 -1800
rect 1750 -1850 1810 -1840
rect 2330 -1840 2450 -1760
rect 1750 -1940 1810 -1930
rect 1750 -1980 1760 -1940
rect 1760 -1980 1800 -1940
rect 1800 -1980 1810 -1940
rect 1750 -2050 1810 -1980
rect 1750 -2080 1810 -2070
rect 1750 -2120 1760 -2080
rect 1760 -2120 1800 -2080
rect 1800 -2120 1810 -2080
rect 1750 -2130 1810 -2120
rect 1750 -2220 1810 -2210
rect 1750 -2260 1760 -2220
rect 1760 -2260 1800 -2220
rect 1800 -2260 1810 -2220
rect 1750 -2270 1810 -2260
rect 1120 -2440 1230 -2350
rect 2040 -2440 2140 -2370
rect 820 -2660 1000 -2520
rect 1350 -2670 1560 -2590
<< metal2 >>
rect 140 200 700 290
rect 140 -130 230 200
rect 590 -130 700 200
rect 1290 130 1640 170
rect 1290 -70 1360 130
rect 1560 -70 1640 130
rect 1290 -110 1640 -70
rect 140 -210 700 -130
rect 250 -220 340 -210
rect -250 -280 -50 -260
rect -250 -440 -230 -280
rect -70 -440 -50 -280
rect -250 -460 -50 -440
rect 10 -310 160 -270
rect 10 -420 30 -310
rect 140 -420 160 -310
rect -210 -650 -30 -630
rect -210 -730 -190 -650
rect -50 -730 -30 -650
rect -210 -1270 -30 -730
rect -210 -1480 -200 -1270
rect -40 -1480 -30 -1270
rect -210 -1490 -30 -1480
rect 10 -830 160 -420
rect 10 -930 40 -830
rect 140 -930 160 -830
rect 10 -2370 160 -930
rect 250 -280 270 -220
rect 330 -280 340 -220
rect 250 -530 340 -280
rect 610 -220 700 -210
rect 610 -280 630 -220
rect 690 -280 700 -220
rect 490 -320 570 -310
rect 490 -390 500 -320
rect 560 -390 570 -320
rect 500 -400 560 -390
rect 250 -590 270 -530
rect 330 -590 340 -530
rect 250 -640 340 -590
rect 250 -700 270 -640
rect 330 -700 340 -640
rect 420 -600 490 -590
rect 420 -660 430 -600
rect 420 -670 490 -660
rect 250 -750 340 -700
rect 250 -810 270 -750
rect 330 -810 340 -750
rect 250 -950 340 -810
rect 520 -850 560 -400
rect 610 -530 700 -280
rect 2150 -210 2650 290
rect 2150 -240 2240 -210
rect 2150 -300 2160 -240
rect 2230 -300 2240 -240
rect 730 -390 820 -380
rect 730 -480 740 -390
rect 810 -480 820 -390
rect 1300 -390 1390 -380
rect 1300 -480 1310 -390
rect 1380 -480 1390 -390
rect 730 -490 820 -480
rect 920 -490 1030 -480
rect 610 -590 620 -530
rect 680 -590 700 -530
rect 610 -650 700 -590
rect 610 -710 620 -650
rect 680 -710 700 -650
rect 920 -550 940 -490
rect 1020 -550 1030 -490
rect 920 -600 1030 -550
rect 920 -680 930 -600
rect 1020 -680 1030 -600
rect 920 -690 1030 -680
rect 1130 -490 1240 -480
rect 1130 -550 1140 -490
rect 1220 -550 1240 -490
rect 1130 -600 1240 -550
rect 1130 -670 1140 -600
rect 1230 -670 1240 -600
rect 610 -750 700 -710
rect 610 -810 620 -750
rect 680 -810 700 -750
rect 380 -860 470 -850
rect 380 -920 390 -860
rect 450 -920 470 -860
rect 380 -930 470 -920
rect 500 -860 580 -850
rect 500 -920 510 -860
rect 570 -920 580 -860
rect 500 -930 580 -920
rect 250 -960 270 -950
rect 230 -1010 270 -960
rect 330 -960 340 -950
rect 610 -950 700 -810
rect 1130 -790 1240 -670
rect 610 -960 630 -950
rect 330 -1010 630 -960
rect 690 -960 700 -950
rect 950 -890 1060 -840
rect 1130 -850 1150 -790
rect 1220 -850 1240 -790
rect 1300 -630 1390 -480
rect 1300 -690 1330 -630
rect 950 -950 970 -890
rect 1030 -950 1060 -890
rect 950 -960 1060 -950
rect 1090 -890 1270 -880
rect 1260 -950 1270 -890
rect 690 -1010 710 -960
rect 230 -1020 710 -1010
rect 1090 -1120 1260 -950
rect 710 -1170 780 -1160
rect 430 -1180 540 -1170
rect 430 -1280 440 -1180
rect 530 -1280 540 -1180
rect 1080 -1180 1100 -1120
rect 1240 -1180 1260 -1120
rect 1300 -1140 1390 -690
rect 710 -1240 780 -1230
rect 1070 -1230 1270 -1220
rect 430 -1290 540 -1280
rect 610 -1360 700 -1350
rect 610 -1440 620 -1360
rect 610 -1450 700 -1440
rect 730 -1670 760 -1240
rect 790 -1290 860 -1280
rect 790 -1630 800 -1290
rect 1070 -1320 1080 -1230
rect 1260 -1320 1270 -1230
rect 1300 -1230 1310 -1140
rect 1380 -1230 1390 -1140
rect 1300 -1250 1390 -1230
rect 1460 -390 1550 -380
rect 1460 -480 1470 -390
rect 1540 -480 1550 -390
rect 2030 -390 2110 -380
rect 1460 -520 1550 -480
rect 1460 -580 1470 -520
rect 1540 -580 1550 -520
rect 1460 -1140 1550 -580
rect 1610 -480 1730 -470
rect 1610 -540 1630 -480
rect 1710 -540 1730 -480
rect 1610 -580 1730 -540
rect 1610 -680 1620 -580
rect 1710 -680 1730 -580
rect 1610 -780 1730 -680
rect 1840 -480 1960 -470
rect 1840 -540 1860 -480
rect 1940 -540 1960 -480
rect 2030 -480 2040 -390
rect 2100 -480 2110 -390
rect 2030 -490 2110 -480
rect 2150 -460 2240 -300
rect 2520 -220 2610 -210
rect 2520 -300 2530 -220
rect 2600 -300 2610 -220
rect 2380 -330 2490 -320
rect 2380 -390 2400 -330
rect 2460 -390 2490 -330
rect 2410 -400 2470 -390
rect 1840 -580 1960 -540
rect 1840 -680 1860 -580
rect 1950 -680 1960 -580
rect 2150 -540 2160 -460
rect 2230 -540 2240 -460
rect 2150 -590 2240 -540
rect 1840 -690 1960 -680
rect 2000 -630 2090 -620
rect 2000 -690 2020 -630
rect 2080 -690 2090 -630
rect 1610 -840 1630 -780
rect 1710 -840 1730 -780
rect 1610 -850 1730 -840
rect 1800 -830 1890 -820
rect 1580 -960 1610 -900
rect 1750 -960 1770 -900
rect 1800 -910 1810 -830
rect 1880 -910 1890 -830
rect 1800 -920 1890 -910
rect 1580 -970 1770 -960
rect 1590 -1110 1770 -970
rect 1460 -1240 1470 -1140
rect 1540 -1240 1550 -1140
rect 1580 -1170 1590 -1110
rect 1770 -1170 1780 -1110
rect 1580 -1180 1780 -1170
rect 2000 -1130 2090 -690
rect 2150 -670 2160 -590
rect 2230 -670 2240 -590
rect 2150 -710 2240 -670
rect 2330 -570 2390 -560
rect 2330 -690 2390 -680
rect 2150 -790 2160 -710
rect 2230 -790 2240 -710
rect 2150 -960 2240 -790
rect 2420 -850 2470 -400
rect 2520 -460 2610 -300
rect 2890 -280 3090 -270
rect 2520 -540 2530 -460
rect 2600 -540 2610 -460
rect 2520 -590 2610 -540
rect 2520 -670 2530 -590
rect 2600 -670 2610 -590
rect 2520 -710 2610 -670
rect 2520 -790 2530 -710
rect 2600 -790 2610 -710
rect 2290 -860 2370 -850
rect 2360 -920 2370 -860
rect 2290 -930 2370 -920
rect 2400 -860 2490 -850
rect 2400 -920 2410 -860
rect 2470 -920 2490 -860
rect 2400 -930 2490 -920
rect 2520 -960 2610 -790
rect 2690 -330 2840 -320
rect 2690 -390 2740 -330
rect 2810 -390 2840 -330
rect 2690 -860 2840 -390
rect 2890 -460 2900 -280
rect 3080 -460 3090 -280
rect 2890 -470 3090 -460
rect 2690 -920 2740 -860
rect 2810 -920 2840 -860
rect 2140 -1020 2160 -960
rect 2220 -1020 2540 -960
rect 2600 -1020 2620 -960
rect 2140 -1030 2620 -1020
rect 2300 -1120 2430 -1110
rect 1460 -1250 1550 -1240
rect 1580 -1230 1790 -1220
rect 1070 -1330 1270 -1320
rect 1580 -1320 1590 -1230
rect 1780 -1320 1790 -1230
rect 1580 -1330 1790 -1320
rect 2000 -1260 2040 -1130
rect 2070 -1170 2150 -1160
rect 2070 -1230 2080 -1170
rect 2140 -1230 2150 -1170
rect 2300 -1230 2310 -1120
rect 2420 -1230 2430 -1120
rect 2300 -1240 2430 -1230
rect 2000 -1280 2090 -1260
rect 1340 -1410 1580 -1390
rect 1340 -1490 1380 -1410
rect 1540 -1490 1580 -1410
rect 1340 -1510 1580 -1490
rect 790 -1640 860 -1630
rect 1040 -1620 1200 -1600
rect 710 -1690 790 -1670
rect 410 -1760 530 -1750
rect 410 -1840 420 -1760
rect 520 -1840 530 -1760
rect 410 -1850 530 -1840
rect 710 -1760 720 -1690
rect 780 -1760 790 -1690
rect 710 -1860 790 -1760
rect 1040 -1770 1050 -1620
rect 1190 -1770 1200 -1620
rect 2000 -1640 2020 -1280
rect 2080 -1640 2090 -1280
rect 2000 -1650 2090 -1640
rect 2690 -1580 2840 -920
rect 2880 -1310 3010 -1300
rect 2880 -1420 2890 -1310
rect 3000 -1420 3010 -1310
rect 2880 -1430 3010 -1420
rect 1040 -1790 1200 -1770
rect 2030 -1690 2170 -1680
rect 2030 -1750 2080 -1690
rect 2140 -1750 2170 -1690
rect 2690 -1720 2700 -1580
rect 2830 -1720 2840 -1580
rect 2690 -1730 2840 -1720
rect 1740 -1790 1820 -1780
rect 1600 -1850 1610 -1790
rect 1670 -1850 1680 -1790
rect 1600 -1860 1680 -1850
rect 1740 -1850 1750 -1790
rect 1810 -1850 1820 -1790
rect 700 -1870 810 -1860
rect 700 -1940 710 -1870
rect 790 -1940 810 -1870
rect 700 -1950 810 -1940
rect 1740 -1930 1820 -1850
rect 1740 -2050 1750 -1930
rect 1810 -2050 1820 -1930
rect 1740 -2070 1820 -2050
rect 1740 -2130 1750 -2070
rect 1810 -2130 1820 -2070
rect 1740 -2210 1820 -2130
rect 1740 -2270 1750 -2210
rect 1810 -2270 1820 -2210
rect 1740 -2280 1820 -2270
rect 10 -2440 20 -2370
rect 150 -2440 160 -2370
rect 10 -2450 160 -2440
rect 1110 -2350 1240 -2340
rect 1110 -2440 1120 -2350
rect 1230 -2440 1240 -2350
rect 1110 -2450 1240 -2440
rect 810 -2520 1010 -2500
rect 810 -2660 820 -2520
rect 1000 -2660 1010 -2520
rect 810 -2680 1010 -2660
rect 1340 -2590 1570 -2580
rect 1340 -2670 1350 -2590
rect 1560 -2670 1570 -2590
rect 1340 -2680 1570 -2670
rect 1720 -2650 1870 -2280
rect 2030 -2370 2170 -1750
rect 2310 -1760 2460 -1750
rect 2310 -1840 2330 -1760
rect 2450 -1840 2460 -1760
rect 2310 -1850 2460 -1840
rect 2030 -2440 2040 -2370
rect 2140 -2440 2170 -2370
rect 2030 -2460 2170 -2440
rect 1720 -2770 1730 -2650
rect 1860 -2770 1870 -2650
rect 1720 -2800 1870 -2770
<< via2 >>
rect 230 -130 590 200
rect 1360 110 1560 130
rect 1360 -50 1380 110
rect 1380 -50 1540 110
rect 1540 -50 1560 110
rect 1360 -70 1560 -50
rect -230 -440 -70 -280
rect 30 -420 140 -310
rect -190 -730 -50 -650
rect -180 -1440 -60 -1360
rect 40 -930 140 -830
rect 500 -330 560 -320
rect 500 -380 560 -330
rect 430 -660 490 -600
rect 740 -480 810 -390
rect 1310 -480 1380 -390
rect 930 -680 1020 -600
rect 1140 -670 1230 -600
rect 390 -920 450 -860
rect 510 -920 570 -860
rect 1330 -690 1390 -630
rect 970 -950 1030 -890
rect 440 -1280 530 -1180
rect 620 -1440 640 -1360
rect 640 -1440 700 -1360
rect 800 -1630 852 -1290
rect 852 -1630 860 -1290
rect 1080 -1320 1260 -1230
rect 1470 -480 1540 -390
rect 1620 -680 1710 -580
rect 2040 -480 2100 -390
rect 2400 -390 2460 -330
rect 1860 -680 1950 -580
rect 2020 -690 2080 -630
rect 1810 -910 1820 -830
rect 1820 -910 1880 -830
rect 2330 -680 2390 -570
rect 2290 -920 2300 -860
rect 2300 -920 2360 -860
rect 2410 -920 2470 -860
rect 2740 -390 2810 -330
rect 2900 -300 3080 -280
rect 2900 -440 2920 -300
rect 2920 -440 3060 -300
rect 3060 -440 3080 -300
rect 2900 -460 3080 -440
rect 2740 -920 2810 -860
rect 1590 -1320 1780 -1230
rect 2310 -1230 2420 -1120
rect 1380 -1490 1540 -1410
rect 420 -1840 520 -1760
rect 1050 -1770 1190 -1620
rect 2020 -1420 2080 -1310
rect 2890 -1420 3000 -1310
rect 2700 -1720 2830 -1580
rect 1610 -1850 1670 -1790
rect 710 -1940 790 -1870
rect 20 -2440 150 -2370
rect 1120 -2440 1230 -2350
rect 820 -2660 1000 -2520
rect 1350 -2670 1560 -2590
rect 2330 -1840 2450 -1760
rect 1730 -2770 1860 -2650
<< metal3 >>
rect 140 200 700 290
rect 140 -130 230 200
rect 590 -130 700 200
rect 1290 130 1640 170
rect 1290 -70 1360 130
rect 1560 -70 1640 130
rect 1290 -110 1640 -70
rect 140 -210 700 -130
rect 2150 -210 2650 290
rect -250 -270 -50 -260
rect -250 -280 200 -270
rect -250 -440 -230 -280
rect -70 -310 200 -280
rect 2890 -280 3090 -270
rect -70 -420 30 -310
rect 140 -320 570 -310
rect 2890 -320 2900 -280
rect 140 -380 500 -320
rect 560 -380 570 -320
rect 2380 -330 2900 -320
rect 140 -400 570 -380
rect 730 -390 1390 -380
rect 140 -420 200 -400
rect -70 -440 200 -420
rect -250 -450 200 -440
rect -250 -460 -50 -450
rect 730 -480 740 -390
rect 810 -480 1310 -390
rect 1380 -480 1390 -390
rect 730 -490 1390 -480
rect 1460 -390 2110 -380
rect 1460 -480 1470 -390
rect 1540 -480 2040 -390
rect 2100 -480 2110 -390
rect 2380 -390 2400 -330
rect 2460 -390 2740 -330
rect 2810 -390 2900 -330
rect 2380 -400 2900 -390
rect 2650 -440 2900 -400
rect 2890 -460 2900 -440
rect 3080 -460 3090 -280
rect 2890 -470 3090 -460
rect 1460 -490 2110 -480
rect 1590 -570 2400 -550
rect 1590 -580 2330 -570
rect 180 -600 1260 -580
rect 180 -630 430 -600
rect -250 -650 430 -630
rect -250 -730 -190 -650
rect -50 -660 430 -650
rect 490 -660 930 -600
rect -50 -680 930 -660
rect 1020 -670 1140 -600
rect 1230 -670 1260 -600
rect 1590 -620 1620 -580
rect 1020 -680 1260 -670
rect 1320 -630 1620 -620
rect -50 -730 230 -680
rect 920 -690 1030 -680
rect 1320 -690 1330 -630
rect 1390 -680 1620 -630
rect 1710 -680 1860 -580
rect 1950 -630 2330 -580
rect 1950 -680 2020 -630
rect 1390 -690 2020 -680
rect 2080 -680 2330 -630
rect 2390 -680 2400 -570
rect 2080 -690 2400 -680
rect 1320 -700 1730 -690
rect 2000 -700 2400 -690
rect -250 -740 230 -730
rect 0 -830 200 -820
rect 1800 -830 2820 -820
rect 0 -930 40 -830
rect 140 -850 200 -830
rect 140 -860 580 -850
rect 140 -920 390 -860
rect 450 -920 510 -860
rect 570 -920 580 -860
rect 980 -880 1370 -830
rect 140 -930 580 -920
rect 950 -890 1370 -880
rect 0 -1050 200 -930
rect 950 -950 970 -890
rect 1030 -910 1370 -890
rect 1800 -910 1810 -830
rect 1880 -860 2820 -830
rect 1880 -910 2290 -860
rect 1030 -950 1040 -910
rect 1800 -920 1890 -910
rect 2280 -920 2290 -910
rect 2360 -920 2410 -860
rect 2470 -920 2740 -860
rect 2810 -920 2820 -860
rect 2280 -930 2820 -920
rect 950 -1050 1040 -950
rect 0 -1110 1040 -1050
rect 2300 -1120 2430 -1110
rect 430 -1180 540 -1170
rect -300 -1350 -10 -1260
rect 430 -1280 440 -1180
rect 530 -1280 540 -1180
rect 1070 -1230 1270 -1220
rect 430 -1290 540 -1280
rect 790 -1290 880 -1280
rect -300 -1360 710 -1350
rect -300 -1440 -180 -1360
rect -60 -1440 620 -1360
rect 700 -1440 710 -1360
rect -300 -1450 710 -1440
rect -300 -1700 -10 -1450
rect 790 -1630 800 -1290
rect 870 -1630 880 -1290
rect 1070 -1320 1080 -1230
rect 1260 -1320 1270 -1230
rect 1070 -1330 1270 -1320
rect 1580 -1230 1790 -1220
rect 1580 -1320 1590 -1230
rect 1780 -1320 1790 -1230
rect 2300 -1230 2310 -1120
rect 2420 -1230 2430 -1120
rect 2300 -1240 2430 -1230
rect 1580 -1330 1790 -1320
rect 2010 -1310 3010 -1300
rect 1340 -1410 1580 -1390
rect 1340 -1490 1380 -1410
rect 1540 -1490 1580 -1410
rect 2010 -1420 2020 -1310
rect 2080 -1420 2890 -1310
rect 3000 -1420 3010 -1310
rect 2010 -1430 3010 -1420
rect 1340 -1510 1580 -1490
rect 2570 -1580 2850 -1570
rect 2570 -1600 2700 -1580
rect 790 -1640 880 -1630
rect 1040 -1620 2700 -1600
rect 410 -1760 530 -1750
rect 410 -1840 420 -1760
rect 520 -1840 530 -1760
rect 410 -1850 530 -1840
rect 710 -1860 790 -1700
rect 1040 -1770 1050 -1620
rect 1190 -1690 2700 -1620
rect 1190 -1770 1200 -1690
rect 1610 -1720 1670 -1690
rect 2570 -1720 2700 -1690
rect 2830 -1720 2850 -1580
rect 2570 -1730 2850 -1720
rect 1040 -1790 1200 -1770
rect 2310 -1760 2460 -1750
rect 1600 -1790 1680 -1780
rect 1600 -1850 1610 -1790
rect 1670 -1850 1680 -1790
rect 2310 -1840 2330 -1760
rect 2450 -1840 2460 -1760
rect 2310 -1850 2460 -1840
rect 700 -1870 810 -1860
rect 1600 -1870 1680 -1850
rect 700 -1940 710 -1870
rect 790 -1940 1680 -1870
rect 700 -1950 810 -1940
rect 10 -2350 1240 -2340
rect 10 -2370 1120 -2350
rect 10 -2440 20 -2370
rect 150 -2440 1120 -2370
rect 1230 -2440 1240 -2350
rect 10 -2450 1240 -2440
rect 810 -2520 1010 -2510
rect 810 -2660 820 -2520
rect 1000 -2660 1010 -2520
rect 810 -2670 1010 -2660
rect 1340 -2570 1570 -2560
rect 1340 -2590 1360 -2570
rect 1340 -2670 1350 -2590
rect 1560 -2670 1570 -2570
rect 1340 -2680 1570 -2670
rect 1720 -2650 1870 -2640
rect 1720 -2770 1730 -2650
rect 1860 -2770 1870 -2650
rect 1720 -2800 1870 -2770
rect 1640 -2810 1870 -2800
rect 1640 -3010 1670 -2810
rect 1840 -3010 1870 -2810
rect 1640 -3040 1870 -3010
<< via3 >>
rect 230 -130 590 200
rect 1360 -70 1560 130
rect 440 -1280 530 -1180
rect 800 -1630 860 -1290
rect 860 -1630 870 -1290
rect 1080 -1320 1260 -1230
rect 1590 -1320 1780 -1230
rect 2310 -1230 2420 -1120
rect 1380 -1490 1540 -1410
rect 420 -1840 520 -1760
rect 2330 -1840 2450 -1760
rect 820 -2660 1000 -2520
rect 1360 -2590 1560 -2570
rect 1360 -2640 1560 -2590
rect 1670 -3010 1840 -2810
<< metal4 >>
rect 140 200 700 290
rect 140 -130 230 200
rect 590 -130 700 200
rect 2150 200 2650 290
rect 140 -210 700 -130
rect 2150 -130 2230 200
rect 2590 -130 2650 200
rect 2150 -210 2650 -130
rect 940 -980 2070 -970
rect 770 -1090 2070 -980
rect 770 -1140 890 -1090
rect 430 -1180 890 -1140
rect 430 -1280 440 -1180
rect 530 -1260 890 -1180
rect 1340 -1220 1580 -1090
rect 1950 -1110 2070 -1090
rect 1950 -1120 2430 -1110
rect 530 -1280 540 -1260
rect 430 -1290 540 -1280
rect 770 -1290 890 -1260
rect 770 -1630 800 -1290
rect 870 -1630 890 -1290
rect 1050 -1230 1790 -1220
rect 1050 -1320 1080 -1230
rect 1260 -1320 1590 -1230
rect 1780 -1320 1790 -1230
rect 1050 -1340 1790 -1320
rect 1950 -1230 2310 -1120
rect 2420 -1230 2430 -1120
rect 1950 -1240 2430 -1230
rect 770 -1750 890 -1630
rect 410 -1760 890 -1750
rect 410 -1840 420 -1760
rect 520 -1840 890 -1760
rect 410 -1850 890 -1840
rect 1340 -1410 1580 -1340
rect 1340 -1490 1380 -1410
rect 1540 -1490 1580 -1410
rect 1340 -2500 1580 -1490
rect 1950 -1750 2070 -1240
rect 1950 -1760 2460 -1750
rect 1950 -1840 2330 -1760
rect 2450 -1840 2460 -1760
rect 1950 -1850 2460 -1840
rect 810 -2520 1580 -2500
rect 810 -2660 820 -2520
rect 1000 -2570 1580 -2520
rect 1000 -2640 1360 -2570
rect 1560 -2640 1690 -2570
rect 1000 -2660 1690 -2640
rect 810 -2680 1690 -2660
rect 1560 -2760 1870 -2740
rect 1800 -2810 1870 -2760
rect 1560 -3010 1670 -3000
rect 1840 -3010 1870 -2810
rect 1560 -3040 1870 -3010
<< via4 >>
rect 230 -130 590 200
rect 1290 130 1640 170
rect 1290 -70 1360 130
rect 1360 -70 1560 130
rect 1560 -70 1640 130
rect 1290 -110 1640 -70
rect 2230 -130 2590 200
rect 1560 -2810 1800 -2760
rect 1560 -3000 1670 -2810
rect 1670 -3000 1800 -2810
<< metal5 >>
rect 140 200 2650 290
rect 140 -130 230 200
rect 590 170 2230 200
rect 590 -110 1290 170
rect 1640 -110 2230 170
rect 590 -130 2230 -110
rect 2590 -130 2650 200
rect 140 -210 2650 -130
rect 1190 -2760 1880 -210
rect 1190 -3000 1560 -2760
rect 1800 -3000 1880 -2760
rect 1190 -3040 1880 -3000
use sky130_fd_sc_hd__inv_4  x1 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 1228 0 -1 -1458
box -38 -48 498 592
use sky130_fd_sc_hd__inv_4  x2
timestamp 1701704242
transform 1 0 1228 0 1 -2622
box -38 -48 498 592
use sky130_fd_pr__nfet_01v8_8X7CJE  XM1
timestamp 1716869746
transform 0 1 1170 -1 0 -877
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_ENQT6S  XM2
timestamp 1716869746
transform 0 1 1170 -1 0 -1193
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_CBNSG2  XM3
timestamp 1716869746
transform 0 1 1683 -1 0 -876
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_GNLSML  XM4
timestamp 1716869746
transform 0 1 1683 -1 0 -1192
box -211 -310 211 310
use sky130_fd_pr__pfet_01v8_K7FRP5  XM5
timestamp 1716869746
transform 0 1 1059 -1 0 -434
box -226 -419 226 419
use sky130_fd_pr__pfet_01v8_GHY9W9  XM6
timestamp 1716869746
transform 0 1 1789 -1 0 -434
box -226 -419 226 419
use sky130_fd_pr__pfet_01v8_E3L9V7  XM7
timestamp 1716869746
transform 1 0 472 0 1 -627
box -275 -419 275 419
use sky130_fd_pr__pfet_01v8_EDASV7  XM8
timestamp 1716869746
transform 1 0 2379 0 1 -627
box -275 -419 275 419
use sky130_fd_pr__nfet_01v8_4WSMTB  XM9
timestamp 1716869746
transform 1 0 745 0 1 -1460
box -221 -410 221 410
use sky130_fd_pr__nfet_01v8_XJSMYS  XM10
timestamp 1716869746
transform 1 0 2111 0 1 -1460
box -221 -410 221 410
<< labels >>
flabel metal1 1360 -70 1560 130 0 FreeSans 256 0 0 0 VDD
port 0 nsew
flabel metal1 810 -2680 1010 -2480 0 FreeSans 256 0 0 0 GND
port 5 nsew
flabel metal1 2890 -470 3090 -270 0 FreeSans 256 0 0 0 R
port 2 nsew
flabel metal1 -250 -460 -50 -260 0 FreeSans 256 0 0 0 S
port 1 nsew
flabel metal1 3010 -1470 3210 -1270 0 FreeSans 256 0 0 0 Q
port 3 nsew
flabel metal1 -220 -1700 -20 -1500 0 FreeSans 256 0 0 0 QN
port 4 nsew
<< end >>
