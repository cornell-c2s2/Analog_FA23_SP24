magic
tech sky130A
timestamp 1709401280
<< metal1 >>
rect 0 0 100 100
rect 0 -200 100 -100
rect 0 -400 100 -300
rect 0 -600 100 -500
rect 0 -800 100 -700
rect 0 -1000 100 -900
rect 0 -1200 100 -1100
rect 0 -1400 100 -1300
rect 0 -1600 100 -1500
rect 0 -1800 100 -1700
rect 0 -2000 100 -1900
use sky130_fd_sc_hd__or4_4  sky130_fd_sc_hd__or4_4_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 1145 0 1 -1726
box -19 -24 433 296
use sky130_fd_sc_hd__or4_4  sky130_fd_sc_hd__or4_4_1
timestamp 1701704242
transform 1 0 1137 0 1 -2236
box -19 -24 433 296
use sky130_fd_sc_hd__or4_4  x0
timestamp 1701704242
transform 1 0 1142 0 1 28
box -19 -24 433 296
use sky130_fd_sc_hd__or4_4  x1
timestamp 1701704242
transform 1 0 1152 0 1 -572
box -19 -24 433 296
use sky130_fd_sc_hd__or4_4  x2
timestamp 1701704242
transform 1 0 1152 0 1 -1155
box -19 -24 433 296
<< labels >>
flabel metal1 0 0 100 100 0 FreeSans 128 0 0 0 Q0
port 0 nsew
flabel metal1 0 -200 100 -100 0 FreeSans 128 0 0 0 D0
port 1 nsew
flabel metal1 0 -400 100 -300 0 FreeSans 128 0 0 0 D1
port 2 nsew
flabel metal1 0 -600 100 -500 0 FreeSans 128 0 0 0 D2
port 3 nsew
flabel metal1 0 -800 100 -700 0 FreeSans 128 0 0 0 D3
port 4 nsew
flabel metal1 0 -1000 100 -900 0 FreeSans 128 0 0 0 Q1
port 5 nsew
flabel metal1 0 -1200 100 -1100 0 FreeSans 128 0 0 0 D4
port 6 nsew
flabel metal1 0 -1400 100 -1300 0 FreeSans 128 0 0 0 D5
port 7 nsew
flabel metal1 0 -1600 100 -1500 0 FreeSans 128 0 0 0 D6
port 8 nsew
flabel metal1 0 -1800 100 -1700 0 FreeSans 128 0 0 0 D7
port 9 nsew
flabel metal1 0 -2000 100 -1900 0 FreeSans 128 0 0 0 Q2
port 10 nsew
<< end >>
