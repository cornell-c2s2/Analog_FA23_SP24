magic
tech sky130A
magscale 1 2
timestamp 1713486840
<< nwell >>
rect 197 -660 2654 -208
rect 197 -1046 747 -660
rect 2104 -1046 2654 -660
rect 1190 -1720 1726 -1719
rect 1190 -2370 1870 -1720
<< pwell >>
rect 1373 -666 1993 -665
rect 860 -1050 1993 -666
rect 520 -1140 2332 -1050
rect 430 -1290 2332 -1140
rect 520 -1403 2332 -1290
rect 520 -1404 1480 -1403
rect 520 -1870 966 -1404
rect 1257 -1479 1291 -1441
rect 1239 -1510 1677 -1479
rect 1890 -1510 2332 -1403
rect 1239 -1590 2332 -1510
rect 1239 -1661 1677 -1590
rect 1890 -1870 2332 -1590
rect 1239 -2420 1677 -2419
rect 1060 -2601 1677 -2420
rect 1060 -2639 1291 -2601
rect 1060 -2680 1260 -2639
rect 1080 -2690 1260 -2680
rect 1080 -2700 1200 -2690
<< nmos >>
rect 1070 -892 1270 -862
rect 1583 -891 1783 -861
rect 720 -1660 770 -1260
rect 1070 -1208 1270 -1178
rect 1583 -1207 1783 -1177
rect 2086 -1660 2136 -1260
<< scnmos >>
rect 1317 -1635 1347 -1505
rect 1401 -1635 1431 -1505
rect 1485 -1635 1515 -1505
rect 1569 -1635 1599 -1505
rect 1317 -2575 1347 -2445
rect 1401 -2575 1431 -2445
rect 1485 -2575 1515 -2445
rect 1569 -2575 1599 -2445
<< pmos >>
rect 393 -827 443 -427
rect 501 -827 551 -427
rect 859 -464 1259 -404
rect 1589 -464 1989 -404
rect 2300 -827 2350 -427
rect 2408 -827 2458 -427
<< scpmoshvt >>
rect 1317 -1955 1347 -1755
rect 1401 -1955 1431 -1755
rect 1485 -1955 1515 -1755
rect 1569 -1955 1599 -1755
rect 1317 -2325 1347 -2125
rect 1401 -2325 1431 -2125
rect 1485 -2325 1515 -2125
rect 1569 -2325 1599 -2125
<< ndiff >>
rect 1150 -804 1220 -790
rect 1070 -816 1270 -804
rect 1070 -850 1082 -816
rect 1258 -850 1270 -816
rect 1070 -862 1270 -850
rect 1070 -904 1270 -892
rect 1070 -938 1082 -904
rect 1258 -938 1270 -904
rect 1070 -950 1270 -938
rect 1583 -815 1783 -803
rect 1583 -849 1595 -815
rect 1771 -849 1783 -815
rect 1583 -861 1783 -849
rect 1583 -903 1783 -891
rect 1583 -937 1595 -903
rect 1771 -937 1783 -903
rect 1583 -949 1783 -937
rect 662 -1272 720 -1260
rect 662 -1648 674 -1272
rect 708 -1648 720 -1272
rect 662 -1660 720 -1648
rect 770 -1272 828 -1260
rect 770 -1648 782 -1272
rect 816 -1648 828 -1272
rect 770 -1660 828 -1648
rect 1070 -1132 1270 -1120
rect 1070 -1166 1082 -1132
rect 1258 -1166 1270 -1132
rect 1070 -1178 1270 -1166
rect 1070 -1220 1270 -1208
rect 1070 -1254 1082 -1220
rect 1258 -1254 1270 -1220
rect 1070 -1266 1270 -1254
rect 1583 -1131 1783 -1119
rect 1583 -1165 1595 -1131
rect 1771 -1165 1783 -1131
rect 1583 -1177 1783 -1165
rect 1583 -1219 1783 -1207
rect 1583 -1253 1595 -1219
rect 1771 -1253 1783 -1219
rect 1583 -1265 1783 -1253
rect 1265 -1517 1317 -1505
rect 1265 -1551 1273 -1517
rect 1307 -1551 1317 -1517
rect 1265 -1635 1317 -1551
rect 1347 -1525 1401 -1505
rect 1347 -1559 1357 -1525
rect 1391 -1559 1401 -1525
rect 1347 -1635 1401 -1559
rect 1431 -1517 1485 -1505
rect 1431 -1551 1441 -1517
rect 1475 -1551 1485 -1517
rect 1431 -1635 1485 -1551
rect 1515 -1525 1569 -1505
rect 1515 -1559 1525 -1525
rect 1559 -1559 1569 -1525
rect 1515 -1635 1569 -1559
rect 1599 -1518 1651 -1505
rect 1599 -1552 1609 -1518
rect 1643 -1552 1651 -1518
rect 1599 -1635 1651 -1552
rect 2028 -1272 2086 -1260
rect 2028 -1648 2040 -1272
rect 2074 -1648 2086 -1272
rect 2028 -1660 2086 -1648
rect 2136 -1272 2194 -1260
rect 2136 -1648 2148 -1272
rect 2182 -1648 2194 -1272
rect 2136 -1660 2194 -1648
rect 1265 -2529 1317 -2445
rect 1265 -2563 1273 -2529
rect 1307 -2563 1317 -2529
rect 1265 -2575 1317 -2563
rect 1347 -2521 1401 -2445
rect 1347 -2555 1357 -2521
rect 1391 -2555 1401 -2521
rect 1347 -2575 1401 -2555
rect 1431 -2529 1485 -2445
rect 1431 -2563 1441 -2529
rect 1475 -2563 1485 -2529
rect 1431 -2575 1485 -2563
rect 1515 -2521 1569 -2445
rect 1515 -2555 1525 -2521
rect 1559 -2555 1569 -2521
rect 1515 -2575 1569 -2555
rect 1599 -2528 1651 -2445
rect 1599 -2562 1609 -2528
rect 1643 -2562 1651 -2528
rect 1599 -2575 1651 -2562
<< pdiff >>
rect 335 -439 393 -427
rect 335 -815 347 -439
rect 381 -815 393 -439
rect 335 -827 393 -815
rect 443 -439 501 -427
rect 443 -815 455 -439
rect 489 -815 501 -439
rect 443 -827 501 -815
rect 551 -439 609 -427
rect 551 -815 563 -439
rect 597 -815 609 -439
rect 859 -358 1259 -346
rect 859 -392 871 -358
rect 1247 -392 1259 -358
rect 859 -404 1259 -392
rect 859 -476 1259 -464
rect 859 -510 871 -476
rect 1247 -510 1259 -476
rect 859 -522 1259 -510
rect 1589 -358 1989 -346
rect 1589 -392 1601 -358
rect 1977 -392 1989 -358
rect 1589 -404 1989 -392
rect 1589 -476 1989 -464
rect 1589 -510 1601 -476
rect 1977 -510 1989 -476
rect 1589 -522 1989 -510
rect 551 -827 609 -815
rect 2242 -439 2300 -427
rect 2242 -815 2254 -439
rect 2288 -815 2300 -439
rect 2242 -827 2300 -815
rect 2350 -439 2408 -427
rect 2350 -815 2362 -439
rect 2396 -815 2408 -439
rect 2350 -827 2408 -815
rect 2458 -439 2516 -427
rect 2458 -815 2470 -439
rect 2504 -815 2516 -439
rect 2458 -827 2516 -815
rect 1265 -1773 1317 -1755
rect 1265 -1807 1273 -1773
rect 1307 -1807 1317 -1773
rect 1265 -1841 1317 -1807
rect 1265 -1875 1273 -1841
rect 1307 -1875 1317 -1841
rect 1265 -1909 1317 -1875
rect 1265 -1943 1273 -1909
rect 1307 -1943 1317 -1909
rect 1265 -1955 1317 -1943
rect 1347 -1773 1401 -1755
rect 1347 -1807 1357 -1773
rect 1391 -1807 1401 -1773
rect 1347 -1841 1401 -1807
rect 1347 -1875 1357 -1841
rect 1391 -1875 1401 -1841
rect 1347 -1909 1401 -1875
rect 1347 -1943 1357 -1909
rect 1391 -1943 1401 -1909
rect 1347 -1955 1401 -1943
rect 1431 -1841 1485 -1755
rect 1431 -1875 1441 -1841
rect 1475 -1875 1485 -1841
rect 1431 -1909 1485 -1875
rect 1431 -1943 1441 -1909
rect 1475 -1943 1485 -1909
rect 1431 -1955 1485 -1943
rect 1515 -1773 1569 -1755
rect 1515 -1807 1525 -1773
rect 1559 -1807 1569 -1773
rect 1515 -1841 1569 -1807
rect 1515 -1875 1525 -1841
rect 1559 -1875 1569 -1841
rect 1515 -1909 1569 -1875
rect 1515 -1943 1525 -1909
rect 1559 -1943 1569 -1909
rect 1515 -1955 1569 -1943
rect 1599 -1909 1651 -1755
rect 1599 -1943 1609 -1909
rect 1643 -1943 1651 -1909
rect 1599 -1955 1651 -1943
rect 1265 -2137 1317 -2125
rect 1265 -2171 1273 -2137
rect 1307 -2171 1317 -2137
rect 1265 -2205 1317 -2171
rect 1265 -2239 1273 -2205
rect 1307 -2239 1317 -2205
rect 1265 -2273 1317 -2239
rect 1265 -2307 1273 -2273
rect 1307 -2307 1317 -2273
rect 1265 -2325 1317 -2307
rect 1347 -2137 1401 -2125
rect 1347 -2171 1357 -2137
rect 1391 -2171 1401 -2137
rect 1347 -2205 1401 -2171
rect 1347 -2239 1357 -2205
rect 1391 -2239 1401 -2205
rect 1347 -2273 1401 -2239
rect 1347 -2307 1357 -2273
rect 1391 -2307 1401 -2273
rect 1347 -2325 1401 -2307
rect 1431 -2137 1485 -2125
rect 1431 -2171 1441 -2137
rect 1475 -2171 1485 -2137
rect 1431 -2205 1485 -2171
rect 1431 -2239 1441 -2205
rect 1475 -2239 1485 -2205
rect 1431 -2325 1485 -2239
rect 1515 -2137 1569 -2125
rect 1515 -2171 1525 -2137
rect 1559 -2171 1569 -2137
rect 1515 -2205 1569 -2171
rect 1515 -2239 1525 -2205
rect 1559 -2239 1569 -2205
rect 1515 -2273 1569 -2239
rect 1515 -2307 1525 -2273
rect 1559 -2307 1569 -2273
rect 1515 -2325 1569 -2307
rect 1599 -2137 1651 -2125
rect 1599 -2171 1609 -2137
rect 1643 -2171 1651 -2137
rect 1599 -2325 1651 -2171
<< ndiffc >>
rect 1082 -850 1258 -816
rect 1082 -938 1258 -904
rect 1595 -849 1771 -815
rect 1595 -937 1771 -903
rect 674 -1648 708 -1272
rect 782 -1648 816 -1272
rect 1082 -1166 1258 -1132
rect 1082 -1254 1258 -1220
rect 1595 -1165 1771 -1131
rect 1595 -1253 1771 -1219
rect 1273 -1551 1307 -1517
rect 1357 -1559 1391 -1525
rect 1441 -1551 1475 -1517
rect 1525 -1559 1559 -1525
rect 1609 -1552 1643 -1518
rect 2040 -1648 2074 -1272
rect 2148 -1648 2182 -1272
rect 1273 -2563 1307 -2529
rect 1357 -2555 1391 -2521
rect 1441 -2563 1475 -2529
rect 1525 -2555 1559 -2521
rect 1609 -2562 1643 -2528
<< pdiffc >>
rect 347 -815 381 -439
rect 455 -815 489 -439
rect 563 -815 597 -439
rect 871 -392 1247 -358
rect 871 -510 1247 -476
rect 1601 -392 1977 -358
rect 1601 -510 1977 -476
rect 2254 -815 2288 -439
rect 2362 -815 2396 -439
rect 2470 -815 2504 -439
rect 1273 -1807 1307 -1773
rect 1273 -1875 1307 -1841
rect 1273 -1943 1307 -1909
rect 1357 -1807 1391 -1773
rect 1357 -1875 1391 -1841
rect 1357 -1943 1391 -1909
rect 1441 -1875 1475 -1841
rect 1441 -1943 1475 -1909
rect 1525 -1807 1559 -1773
rect 1525 -1875 1559 -1841
rect 1525 -1943 1559 -1909
rect 1609 -1943 1643 -1909
rect 1273 -2171 1307 -2137
rect 1273 -2239 1307 -2205
rect 1273 -2307 1307 -2273
rect 1357 -2171 1391 -2137
rect 1357 -2239 1391 -2205
rect 1357 -2307 1391 -2273
rect 1441 -2171 1475 -2137
rect 1441 -2239 1475 -2205
rect 1525 -2171 1559 -2137
rect 1525 -2239 1559 -2205
rect 1525 -2307 1559 -2273
rect 1609 -2171 1643 -2137
<< psubdiff >>
rect 1409 -702 1505 -701
rect 896 -736 992 -702
rect 1348 -735 1505 -702
rect 1861 -735 1957 -701
rect 1348 -736 1444 -735
rect 896 -798 930 -736
rect 896 -1018 930 -956
rect 1409 -1017 1444 -736
rect 1923 -797 1957 -735
rect 1923 -1017 1957 -955
rect 1409 -1018 1957 -1017
rect 896 -1051 1957 -1018
rect 896 -1052 1444 -1051
rect 896 -1086 930 -1052
rect 560 -1120 656 -1086
rect 834 -1114 930 -1086
rect 834 -1120 896 -1114
rect 560 -1182 594 -1120
rect 896 -1334 930 -1272
rect 1409 -1333 1444 -1052
rect 1923 -1086 1957 -1051
rect 1923 -1113 2022 -1086
rect 1957 -1120 2022 -1113
rect 2200 -1120 2296 -1086
rect 1957 -1271 1960 -1120
rect 2262 -1182 2296 -1120
rect 1923 -1333 1960 -1271
rect 1409 -1334 1505 -1333
rect 896 -1368 992 -1334
rect 1348 -1367 1505 -1334
rect 1861 -1367 1960 -1333
rect 1348 -1368 1444 -1367
rect 560 -1800 594 -1738
rect 896 -1800 930 -1368
rect 560 -1834 656 -1800
rect 834 -1834 930 -1800
rect 1926 -1800 1960 -1367
rect 2262 -1800 2296 -1738
rect 1926 -1834 2022 -1800
rect 2200 -1834 2296 -1800
rect 1090 -2530 1190 -2500
rect 1090 -2600 1120 -2530
rect 1100 -2650 1120 -2600
rect 1160 -2600 1190 -2530
rect 1160 -2650 1180 -2600
rect 1100 -2680 1180 -2650
<< nsubdiff >>
rect 233 -278 329 -244
rect 615 -278 772 -244
rect 1346 -278 1502 -244
rect 2076 -278 2236 -244
rect 2522 -278 2618 -244
rect 233 -340 267 -278
rect 676 -340 711 -278
rect 710 -528 711 -340
rect 676 -590 711 -528
rect 1406 -590 1442 -278
rect 2138 -340 2174 -278
rect 2172 -528 2174 -340
rect 2584 -340 2618 -278
rect 2138 -590 2174 -528
rect 676 -624 772 -590
rect 1346 -624 1502 -590
rect 2076 -624 2174 -590
rect 233 -976 267 -914
rect 677 -976 711 -624
rect 233 -1010 329 -976
rect 615 -1010 711 -976
rect 2140 -976 2174 -624
rect 2584 -976 2618 -914
rect 2140 -1010 2236 -976
rect 2522 -1010 2618 -976
rect 1730 -1800 1830 -1780
rect 1730 -1840 1760 -1800
rect 1800 -1840 1830 -1800
rect 1730 -1860 1830 -1840
rect 1730 -1940 1830 -1920
rect 1730 -1980 1760 -1940
rect 1800 -1980 1830 -1940
rect 1730 -2000 1830 -1980
rect 1730 -2080 1830 -2060
rect 1730 -2120 1760 -2080
rect 1800 -2120 1830 -2080
rect 1730 -2140 1830 -2120
rect 1730 -2220 1830 -2200
rect 1730 -2260 1760 -2220
rect 1800 -2260 1830 -2220
rect 1730 -2280 1830 -2260
<< psubdiffcont >>
rect 992 -736 1348 -702
rect 1505 -735 1861 -701
rect 896 -956 930 -798
rect 1923 -955 1957 -797
rect 656 -1120 834 -1086
rect 560 -1738 594 -1182
rect 896 -1272 930 -1114
rect 1923 -1271 1957 -1113
rect 2022 -1120 2200 -1086
rect 992 -1368 1348 -1334
rect 1505 -1367 1861 -1333
rect 656 -1834 834 -1800
rect 2262 -1738 2296 -1182
rect 2022 -1834 2200 -1800
rect 1120 -2650 1160 -2530
<< nsubdiffcont >>
rect 329 -278 615 -244
rect 772 -278 1346 -244
rect 1502 -278 2076 -244
rect 2236 -278 2522 -244
rect 233 -914 267 -340
rect 676 -528 710 -340
rect 2138 -528 2172 -340
rect 772 -624 1346 -590
rect 1502 -624 2076 -590
rect 329 -1010 615 -976
rect 2584 -914 2618 -340
rect 2236 -1010 2522 -976
rect 1760 -1840 1800 -1800
rect 1760 -1980 1800 -1940
rect 1760 -2120 1800 -2080
rect 1760 -2260 1800 -2220
<< poly >>
rect 493 -346 559 -330
rect 493 -380 509 -346
rect 543 -380 559 -346
rect 493 -396 559 -380
rect 393 -427 443 -401
rect 501 -427 551 -396
rect 762 -404 828 -401
rect 1290 -404 1356 -401
rect 762 -417 859 -404
rect 762 -451 778 -417
rect 812 -451 859 -417
rect 762 -464 859 -451
rect 1259 -417 1356 -404
rect 1259 -451 1306 -417
rect 1340 -451 1356 -417
rect 1259 -464 1356 -451
rect 762 -467 828 -464
rect 1290 -467 1356 -464
rect 1492 -404 1558 -401
rect 2020 -404 2086 -401
rect 1492 -417 1589 -404
rect 1492 -451 1508 -417
rect 1542 -451 1589 -417
rect 1492 -464 1589 -451
rect 1989 -417 2086 -404
rect 1989 -451 2036 -417
rect 2070 -451 2086 -417
rect 1989 -464 2086 -451
rect 1492 -467 1558 -464
rect 2020 -467 2086 -464
rect 2400 -346 2466 -330
rect 2400 -380 2416 -346
rect 2450 -380 2466 -346
rect 2400 -396 2466 -380
rect 2300 -427 2350 -401
rect 2408 -427 2458 -396
rect 393 -858 443 -827
rect 501 -853 551 -827
rect 385 -874 451 -858
rect 385 -908 401 -874
rect 435 -908 451 -874
rect 385 -924 451 -908
rect 982 -860 1048 -844
rect 982 -894 998 -860
rect 1032 -862 1048 -860
rect 1292 -860 1358 -844
rect 1292 -862 1308 -860
rect 1032 -892 1070 -862
rect 1270 -892 1308 -862
rect 1032 -894 1048 -892
rect 982 -910 1048 -894
rect 1292 -894 1308 -892
rect 1342 -894 1358 -860
rect 1292 -910 1358 -894
rect 1480 -843 1530 -840
rect 1480 -859 1561 -843
rect 1480 -893 1511 -859
rect 1545 -861 1561 -859
rect 1805 -859 1871 -843
rect 1805 -861 1821 -859
rect 1545 -891 1583 -861
rect 1783 -891 1821 -861
rect 1545 -893 1561 -891
rect 1480 -909 1561 -893
rect 1480 -910 1530 -909
rect 1805 -893 1821 -891
rect 1855 -893 1871 -859
rect 1805 -909 1871 -893
rect 2300 -858 2350 -827
rect 2408 -853 2458 -827
rect 2292 -874 2358 -858
rect 2292 -908 2308 -874
rect 2342 -908 2358 -874
rect 2292 -924 2358 -908
rect 712 -1188 778 -1172
rect 712 -1222 728 -1188
rect 762 -1222 778 -1188
rect 712 -1238 778 -1222
rect 720 -1260 770 -1238
rect 982 -1176 1048 -1160
rect 982 -1210 998 -1176
rect 1032 -1178 1048 -1176
rect 1292 -1176 1358 -1160
rect 1292 -1178 1308 -1176
rect 1032 -1208 1070 -1178
rect 1270 -1208 1308 -1178
rect 1032 -1210 1048 -1208
rect 982 -1226 1048 -1210
rect 1292 -1210 1308 -1208
rect 1342 -1210 1358 -1176
rect 1292 -1226 1358 -1210
rect 1495 -1175 1561 -1159
rect 1495 -1209 1511 -1175
rect 1545 -1177 1561 -1175
rect 1805 -1175 1871 -1159
rect 1805 -1177 1821 -1175
rect 1545 -1207 1583 -1177
rect 1783 -1207 1821 -1177
rect 1545 -1209 1561 -1207
rect 1495 -1225 1561 -1209
rect 1805 -1209 1821 -1207
rect 1855 -1209 1871 -1175
rect 1805 -1225 1871 -1209
rect 2078 -1188 2144 -1172
rect 2078 -1222 2094 -1188
rect 2128 -1222 2144 -1188
rect 2078 -1238 2144 -1222
rect 2086 -1260 2136 -1238
rect 720 -1682 770 -1660
rect 712 -1698 778 -1682
rect 712 -1732 728 -1698
rect 762 -1732 778 -1698
rect 712 -1748 778 -1732
rect 1317 -1505 1347 -1479
rect 1401 -1505 1431 -1479
rect 1485 -1505 1515 -1479
rect 1569 -1505 1599 -1479
rect 1317 -1657 1347 -1635
rect 1401 -1657 1431 -1635
rect 1485 -1657 1515 -1635
rect 1569 -1657 1599 -1635
rect 1249 -1673 1599 -1657
rect 1249 -1707 1265 -1673
rect 1299 -1707 1357 -1673
rect 1391 -1707 1441 -1673
rect 1475 -1707 1525 -1673
rect 1559 -1707 1599 -1673
rect 1249 -1723 1599 -1707
rect 1317 -1755 1347 -1723
rect 1401 -1755 1431 -1723
rect 1485 -1755 1515 -1723
rect 1569 -1755 1599 -1723
rect 2086 -1682 2136 -1660
rect 2078 -1698 2144 -1682
rect 2078 -1732 2094 -1698
rect 2128 -1732 2144 -1698
rect 2078 -1748 2144 -1732
rect 1317 -1981 1347 -1955
rect 1401 -1981 1431 -1955
rect 1485 -1981 1515 -1955
rect 1569 -1981 1599 -1955
rect 1317 -2125 1347 -2099
rect 1401 -2125 1431 -2099
rect 1485 -2125 1515 -2099
rect 1569 -2125 1599 -2099
rect 1317 -2357 1347 -2325
rect 1401 -2357 1431 -2325
rect 1485 -2357 1515 -2325
rect 1569 -2357 1599 -2325
rect 1249 -2373 1599 -2357
rect 1249 -2407 1265 -2373
rect 1299 -2407 1357 -2373
rect 1391 -2407 1441 -2373
rect 1475 -2407 1525 -2373
rect 1559 -2407 1599 -2373
rect 1249 -2423 1599 -2407
rect 1317 -2445 1347 -2423
rect 1401 -2445 1431 -2423
rect 1485 -2445 1515 -2423
rect 1569 -2445 1599 -2423
rect 1317 -2601 1347 -2575
rect 1401 -2601 1431 -2575
rect 1485 -2601 1515 -2575
rect 1569 -2601 1599 -2575
<< polycont >>
rect 509 -380 543 -346
rect 778 -451 812 -417
rect 1306 -451 1340 -417
rect 1508 -451 1542 -417
rect 2036 -451 2070 -417
rect 2416 -380 2450 -346
rect 401 -908 435 -874
rect 998 -894 1032 -860
rect 1308 -894 1342 -860
rect 1511 -893 1545 -859
rect 1821 -893 1855 -859
rect 2308 -908 2342 -874
rect 728 -1222 762 -1188
rect 998 -1210 1032 -1176
rect 1308 -1210 1342 -1176
rect 1511 -1209 1545 -1175
rect 1821 -1209 1855 -1175
rect 2094 -1222 2128 -1188
rect 728 -1732 762 -1698
rect 1265 -1707 1299 -1673
rect 1357 -1707 1391 -1673
rect 1441 -1707 1475 -1673
rect 1525 -1707 1559 -1673
rect 2094 -1732 2128 -1698
rect 1265 -2407 1299 -2373
rect 1357 -2407 1391 -2373
rect 1441 -2407 1475 -2373
rect 1525 -2407 1559 -2373
<< locali >>
rect 310 -244 320 -240
rect 620 -244 640 -240
rect 233 -278 320 -244
rect 620 -278 772 -244
rect 2076 -278 2210 -244
rect 233 -340 267 -278
rect 310 -280 320 -278
rect 620 -280 640 -278
rect 676 -340 711 -278
rect 493 -380 509 -346
rect 543 -380 559 -346
rect 347 -439 381 -423
rect 347 -831 381 -815
rect 455 -439 489 -423
rect 455 -831 489 -815
rect 563 -439 597 -423
rect 710 -528 711 -340
rect 855 -392 871 -358
rect 1247 -392 1263 -358
rect 778 -417 812 -401
rect 778 -467 812 -451
rect 1306 -417 1340 -401
rect 1306 -467 1340 -451
rect 855 -510 871 -476
rect 1247 -510 1263 -476
rect 676 -590 711 -528
rect 1406 -590 1442 -280
rect 2138 -340 2174 -278
rect 2600 -280 2618 -244
rect 1585 -392 1601 -358
rect 1977 -392 1993 -358
rect 1508 -417 1542 -401
rect 1508 -467 1542 -451
rect 2036 -417 2070 -401
rect 2036 -467 2070 -451
rect 1585 -510 1601 -476
rect 1977 -510 1993 -476
rect 2172 -528 2174 -340
rect 2584 -340 2618 -280
rect 2400 -380 2416 -346
rect 2450 -380 2466 -346
rect 2138 -590 2174 -528
rect 676 -624 772 -590
rect 1346 -624 1502 -590
rect 2076 -624 2174 -590
rect 563 -831 597 -815
rect 385 -908 401 -874
rect 435 -908 451 -874
rect 233 -976 267 -914
rect 677 -976 711 -624
rect 1409 -702 1500 -701
rect 896 -736 990 -702
rect 1350 -735 1500 -702
rect 1870 -735 1957 -701
rect 1350 -736 1444 -735
rect 896 -790 930 -736
rect 998 -860 1032 -844
rect 1066 -850 1082 -816
rect 1258 -850 1274 -816
rect 998 -910 1032 -894
rect 1308 -860 1342 -844
rect 1066 -938 1082 -904
rect 1258 -938 1274 -904
rect 1308 -910 1342 -894
rect 233 -1010 329 -976
rect 620 -1010 711 -976
rect 896 -1018 930 -970
rect 1409 -1017 1444 -736
rect 1923 -790 1957 -735
rect 1511 -859 1545 -843
rect 1579 -849 1595 -815
rect 1771 -849 1787 -815
rect 1511 -909 1545 -893
rect 1821 -859 1855 -843
rect 1579 -937 1595 -903
rect 1771 -937 1787 -903
rect 1821 -909 1855 -893
rect 1923 -1017 1957 -960
rect 2140 -976 2174 -624
rect 2254 -439 2288 -423
rect 2254 -831 2288 -815
rect 2362 -439 2396 -423
rect 2362 -831 2396 -815
rect 2470 -439 2504 -423
rect 2470 -831 2504 -815
rect 2292 -908 2308 -874
rect 2342 -908 2358 -874
rect 2584 -976 2618 -914
rect 2140 -1010 2230 -976
rect 2530 -1010 2618 -976
rect 1409 -1018 1957 -1017
rect 896 -1051 1957 -1018
rect 896 -1052 1444 -1051
rect 896 -1086 930 -1052
rect 560 -1120 650 -1086
rect 840 -1114 930 -1086
rect 840 -1120 896 -1114
rect 560 -1180 594 -1120
rect 712 -1222 728 -1188
rect 762 -1222 778 -1188
rect 674 -1272 708 -1256
rect 674 -1664 708 -1648
rect 782 -1272 816 -1256
rect 782 -1664 816 -1648
rect 998 -1176 1032 -1160
rect 1066 -1166 1082 -1132
rect 1258 -1166 1274 -1132
rect 998 -1226 1032 -1210
rect 1308 -1176 1342 -1160
rect 1066 -1254 1082 -1220
rect 1258 -1254 1274 -1220
rect 1308 -1226 1342 -1210
rect 896 -1334 930 -1272
rect 1409 -1333 1444 -1052
rect 1923 -1086 1957 -1051
rect 1923 -1113 2020 -1086
rect 1511 -1175 1545 -1159
rect 1579 -1165 1595 -1131
rect 1771 -1165 1787 -1131
rect 1511 -1225 1545 -1209
rect 1821 -1175 1855 -1159
rect 1579 -1253 1595 -1219
rect 1771 -1253 1787 -1219
rect 1821 -1225 1855 -1209
rect 1957 -1120 2020 -1113
rect 2200 -1120 2296 -1086
rect 1957 -1271 1960 -1120
rect 2262 -1180 2296 -1120
rect 2078 -1222 2094 -1188
rect 2128 -1222 2144 -1188
rect 1923 -1333 1960 -1271
rect 1409 -1334 1505 -1333
rect 896 -1368 992 -1334
rect 1348 -1367 1505 -1334
rect 1861 -1367 1960 -1333
rect 1348 -1368 1444 -1367
rect 712 -1732 728 -1698
rect 762 -1732 778 -1698
rect 560 -1800 594 -1740
rect 896 -1800 930 -1368
rect 1228 -1475 1257 -1441
rect 1291 -1475 1349 -1441
rect 1383 -1475 1441 -1441
rect 1475 -1475 1533 -1441
rect 1567 -1475 1625 -1441
rect 1659 -1475 1688 -1441
rect 1254 -1517 1307 -1475
rect 1254 -1551 1273 -1517
rect 1254 -1567 1307 -1551
rect 1341 -1525 1407 -1509
rect 1341 -1559 1357 -1525
rect 1391 -1559 1407 -1525
rect 1341 -1603 1407 -1559
rect 1441 -1517 1475 -1475
rect 1441 -1567 1475 -1551
rect 1509 -1525 1575 -1509
rect 1509 -1559 1525 -1525
rect 1559 -1559 1575 -1525
rect 1509 -1603 1575 -1559
rect 1609 -1518 1659 -1475
rect 1643 -1552 1659 -1518
rect 1609 -1568 1659 -1552
rect 1341 -1611 1662 -1603
rect 1341 -1639 1625 -1611
rect 1609 -1645 1625 -1639
rect 1659 -1645 1662 -1611
rect 1249 -1680 1265 -1673
rect 1299 -1680 1357 -1673
rect 1391 -1680 1441 -1673
rect 1475 -1680 1525 -1673
rect 1559 -1680 1575 -1673
rect 1249 -1720 1260 -1680
rect 1300 -1720 1350 -1680
rect 1391 -1707 1440 -1680
rect 1390 -1720 1440 -1707
rect 1480 -1720 1520 -1680
rect 1560 -1720 1575 -1680
rect 1249 -1723 1575 -1720
rect 1609 -1683 1662 -1645
rect 1609 -1719 1625 -1683
rect 1659 -1719 1662 -1683
rect 1609 -1757 1662 -1719
rect 560 -1834 656 -1800
rect 834 -1834 930 -1800
rect 1254 -1773 1307 -1757
rect 1254 -1807 1273 -1773
rect 1254 -1841 1307 -1807
rect 1254 -1875 1273 -1841
rect 1254 -1909 1307 -1875
rect 1254 -1943 1273 -1909
rect 1254 -1985 1307 -1943
rect 1341 -1763 1662 -1757
rect 1341 -1773 1625 -1763
rect 1341 -1807 1357 -1773
rect 1391 -1791 1525 -1773
rect 1391 -1807 1407 -1791
rect 1341 -1841 1407 -1807
rect 1509 -1807 1525 -1791
rect 1559 -1795 1625 -1773
rect 1559 -1807 1575 -1795
rect 1659 -1795 1662 -1763
rect 1341 -1875 1357 -1841
rect 1391 -1875 1407 -1841
rect 1341 -1909 1407 -1875
rect 1341 -1943 1357 -1909
rect 1391 -1943 1407 -1909
rect 1341 -1951 1407 -1943
rect 1441 -1841 1475 -1825
rect 1441 -1909 1475 -1875
rect 1441 -1985 1475 -1943
rect 1509 -1841 1575 -1807
rect 1509 -1875 1525 -1841
rect 1559 -1875 1575 -1841
rect 1740 -1800 1820 -1780
rect 1740 -1840 1760 -1800
rect 1800 -1840 1820 -1800
rect 1926 -1800 1960 -1367
rect 2040 -1272 2074 -1256
rect 2040 -1664 2074 -1648
rect 2148 -1272 2182 -1256
rect 2148 -1664 2182 -1648
rect 2078 -1732 2094 -1698
rect 2128 -1732 2144 -1698
rect 2262 -1800 2296 -1740
rect 1926 -1834 2022 -1800
rect 2200 -1834 2296 -1800
rect 1740 -1860 1820 -1840
rect 1509 -1909 1575 -1875
rect 1509 -1943 1525 -1909
rect 1559 -1943 1575 -1909
rect 1509 -1951 1575 -1943
rect 1609 -1909 1651 -1893
rect 1643 -1943 1651 -1909
rect 1609 -1985 1651 -1943
rect 1740 -1940 1820 -1920
rect 1740 -1980 1760 -1940
rect 1800 -1980 1820 -1940
rect 1228 -2019 1257 -1985
rect 1291 -2019 1349 -1985
rect 1383 -2019 1441 -1985
rect 1475 -2019 1533 -1985
rect 1567 -2019 1625 -1985
rect 1659 -2019 1688 -1985
rect 1740 -2000 1820 -1980
rect 1228 -2095 1257 -2061
rect 1291 -2095 1349 -2061
rect 1383 -2095 1441 -2061
rect 1475 -2095 1533 -2061
rect 1567 -2095 1625 -2061
rect 1659 -2095 1688 -2061
rect 1740 -2080 1820 -2060
rect 1254 -2137 1307 -2095
rect 1254 -2171 1273 -2137
rect 1254 -2205 1307 -2171
rect 1254 -2239 1273 -2205
rect 1254 -2273 1307 -2239
rect 1254 -2307 1273 -2273
rect 1254 -2323 1307 -2307
rect 1341 -2137 1407 -2129
rect 1341 -2171 1357 -2137
rect 1391 -2171 1407 -2137
rect 1341 -2205 1407 -2171
rect 1341 -2239 1357 -2205
rect 1391 -2239 1407 -2205
rect 1341 -2273 1407 -2239
rect 1441 -2137 1475 -2095
rect 1441 -2205 1475 -2171
rect 1441 -2255 1475 -2239
rect 1509 -2137 1575 -2129
rect 1509 -2171 1525 -2137
rect 1559 -2171 1575 -2137
rect 1509 -2205 1575 -2171
rect 1609 -2137 1651 -2095
rect 1643 -2171 1651 -2137
rect 1740 -2120 1760 -2080
rect 1800 -2120 1820 -2080
rect 1740 -2140 1820 -2120
rect 1609 -2187 1651 -2171
rect 1509 -2239 1525 -2205
rect 1559 -2239 1575 -2205
rect 1341 -2307 1357 -2273
rect 1391 -2289 1407 -2273
rect 1509 -2273 1575 -2239
rect 1509 -2289 1525 -2273
rect 1391 -2307 1525 -2289
rect 1559 -2285 1575 -2273
rect 1740 -2220 1820 -2200
rect 1740 -2260 1760 -2220
rect 1800 -2260 1820 -2220
rect 1740 -2280 1820 -2260
rect 1559 -2294 1662 -2285
rect 1559 -2307 1625 -2294
rect 1341 -2323 1625 -2307
rect 1609 -2329 1625 -2323
rect 1659 -2329 1662 -2294
rect 1249 -2360 1575 -2357
rect 1249 -2400 1260 -2360
rect 1300 -2400 1350 -2360
rect 1390 -2373 1440 -2360
rect 1391 -2400 1440 -2373
rect 1480 -2400 1520 -2360
rect 1560 -2400 1575 -2360
rect 1249 -2407 1265 -2400
rect 1299 -2407 1357 -2400
rect 1391 -2407 1441 -2400
rect 1475 -2407 1525 -2400
rect 1559 -2407 1575 -2400
rect 1609 -2367 1662 -2329
rect 1609 -2402 1625 -2367
rect 1659 -2402 1662 -2367
rect 1609 -2441 1662 -2402
rect 1341 -2443 1662 -2441
rect 1341 -2477 1624 -2443
rect 1090 -2510 1190 -2500
rect 1090 -2600 1100 -2510
rect 1180 -2600 1190 -2510
rect 1254 -2529 1307 -2513
rect 1254 -2563 1273 -2529
rect 1254 -2605 1307 -2563
rect 1341 -2521 1407 -2477
rect 1341 -2555 1357 -2521
rect 1391 -2555 1407 -2521
rect 1341 -2571 1407 -2555
rect 1441 -2529 1475 -2513
rect 1441 -2605 1475 -2563
rect 1509 -2521 1575 -2477
rect 1658 -2477 1662 -2443
rect 1509 -2555 1525 -2521
rect 1559 -2555 1575 -2521
rect 1509 -2571 1575 -2555
rect 1609 -2528 1659 -2512
rect 1643 -2562 1659 -2528
rect 1609 -2605 1659 -2562
rect 1228 -2639 1257 -2605
rect 1291 -2639 1349 -2605
rect 1383 -2639 1441 -2605
rect 1475 -2639 1533 -2605
rect 1567 -2639 1625 -2605
rect 1659 -2639 1688 -2605
<< viali >>
rect 320 -244 620 -240
rect 860 -244 1990 -240
rect 2210 -244 2600 -240
rect 320 -278 329 -244
rect 329 -278 615 -244
rect 615 -278 620 -244
rect 860 -278 1346 -244
rect 1346 -278 1502 -244
rect 1502 -278 1990 -244
rect 2210 -278 2236 -244
rect 2236 -278 2522 -244
rect 2522 -278 2600 -244
rect 320 -280 620 -278
rect 860 -280 1990 -278
rect 509 -380 543 -346
rect 347 -815 381 -439
rect 455 -815 489 -439
rect 563 -815 597 -439
rect 871 -392 1247 -358
rect 778 -451 812 -417
rect 1306 -451 1340 -417
rect 871 -510 1247 -476
rect 2210 -280 2600 -278
rect 1601 -392 1977 -358
rect 1508 -451 1542 -417
rect 2036 -451 2070 -417
rect 1601 -510 1977 -476
rect 2416 -380 2450 -346
rect 401 -908 435 -874
rect 330 -976 620 -970
rect 990 -702 1350 -700
rect 1500 -701 1870 -700
rect 990 -736 992 -702
rect 992 -736 1348 -702
rect 1348 -736 1350 -702
rect 1500 -735 1505 -701
rect 1505 -735 1861 -701
rect 1861 -735 1870 -701
rect 990 -740 1350 -736
rect 890 -798 930 -790
rect 890 -956 896 -798
rect 896 -956 930 -798
rect 1082 -850 1258 -816
rect 998 -894 1032 -860
rect 1308 -894 1342 -860
rect 1082 -938 1258 -904
rect 890 -970 930 -956
rect 330 -1010 615 -976
rect 615 -1010 620 -976
rect 1500 -740 1870 -735
rect 1920 -797 1960 -790
rect 1595 -849 1771 -815
rect 1511 -893 1545 -859
rect 1821 -893 1855 -859
rect 1595 -937 1771 -903
rect 1920 -955 1923 -797
rect 1923 -955 1957 -797
rect 1957 -955 1960 -797
rect 1920 -960 1960 -955
rect 2254 -815 2288 -439
rect 2362 -815 2396 -439
rect 2470 -815 2504 -439
rect 2308 -908 2342 -874
rect 2230 -976 2530 -970
rect 2230 -1010 2236 -976
rect 2236 -1010 2522 -976
rect 2522 -1010 2530 -976
rect 2230 -1020 2530 -1010
rect 650 -1086 840 -1080
rect 650 -1120 656 -1086
rect 656 -1120 834 -1086
rect 834 -1120 840 -1086
rect 560 -1182 600 -1180
rect 560 -1738 594 -1182
rect 594 -1738 600 -1182
rect 728 -1222 762 -1188
rect 674 -1648 708 -1272
rect 782 -1648 816 -1272
rect 1082 -1166 1258 -1132
rect 998 -1210 1032 -1176
rect 1308 -1210 1342 -1176
rect 1082 -1254 1258 -1220
rect 2020 -1086 2200 -1080
rect 1595 -1165 1771 -1131
rect 1511 -1209 1545 -1175
rect 1821 -1209 1855 -1175
rect 1595 -1253 1771 -1219
rect 2020 -1120 2022 -1086
rect 2022 -1120 2200 -1086
rect 2260 -1182 2300 -1180
rect 2094 -1222 2128 -1188
rect 728 -1732 762 -1698
rect 560 -1740 600 -1738
rect 1257 -1475 1291 -1441
rect 1349 -1475 1383 -1441
rect 1441 -1475 1475 -1441
rect 1533 -1475 1567 -1441
rect 1625 -1475 1659 -1441
rect 1625 -1645 1659 -1611
rect 1260 -1707 1265 -1680
rect 1265 -1707 1299 -1680
rect 1299 -1707 1300 -1680
rect 1260 -1720 1300 -1707
rect 1350 -1707 1357 -1680
rect 1357 -1707 1390 -1680
rect 1440 -1707 1441 -1680
rect 1441 -1707 1475 -1680
rect 1475 -1707 1480 -1680
rect 1350 -1720 1390 -1707
rect 1440 -1720 1480 -1707
rect 1520 -1707 1525 -1680
rect 1525 -1707 1559 -1680
rect 1559 -1707 1560 -1680
rect 1520 -1720 1560 -1707
rect 1625 -1719 1659 -1683
rect 1625 -1798 1659 -1763
rect 1760 -1840 1800 -1800
rect 2040 -1648 2074 -1272
rect 2148 -1648 2182 -1272
rect 2094 -1732 2128 -1698
rect 2260 -1738 2262 -1182
rect 2262 -1738 2296 -1182
rect 2296 -1738 2300 -1182
rect 2260 -1740 2300 -1738
rect 1760 -1980 1800 -1940
rect 1257 -2019 1291 -1985
rect 1349 -2019 1383 -1985
rect 1441 -2019 1475 -1985
rect 1533 -2019 1567 -1985
rect 1625 -2019 1659 -1985
rect 1257 -2095 1291 -2061
rect 1349 -2095 1383 -2061
rect 1441 -2095 1475 -2061
rect 1533 -2095 1567 -2061
rect 1625 -2095 1659 -2061
rect 1760 -2120 1800 -2080
rect 1760 -2260 1800 -2220
rect 1625 -2329 1659 -2294
rect 1260 -2373 1300 -2360
rect 1260 -2400 1265 -2373
rect 1265 -2400 1299 -2373
rect 1299 -2400 1300 -2373
rect 1350 -2373 1390 -2360
rect 1440 -2373 1480 -2360
rect 1350 -2400 1357 -2373
rect 1357 -2400 1390 -2373
rect 1440 -2400 1441 -2373
rect 1441 -2400 1475 -2373
rect 1475 -2400 1480 -2373
rect 1520 -2373 1560 -2360
rect 1520 -2400 1525 -2373
rect 1525 -2400 1559 -2373
rect 1559 -2400 1560 -2373
rect 1625 -2402 1659 -2367
rect 1100 -2530 1180 -2510
rect 1100 -2650 1120 -2530
rect 1120 -2650 1160 -2530
rect 1160 -2650 1180 -2530
rect 1624 -2478 1658 -2443
rect 1257 -2639 1291 -2605
rect 1349 -2639 1383 -2605
rect 1441 -2639 1475 -2605
rect 1533 -2639 1567 -2605
rect 1625 -2639 1659 -2605
rect 1100 -2680 1180 -2650
<< metal1 >>
rect 1360 110 1560 130
rect 1360 -50 1380 110
rect 1540 -50 1560 110
rect 1360 -70 1560 -50
rect -350 -280 -50 -90
rect 692 -210 786 -208
rect -350 -440 -230 -280
rect -70 -440 -50 -280
rect 250 -220 2620 -210
rect 250 -280 270 -220
rect 330 -240 630 -220
rect 620 -280 630 -240
rect 690 -240 2530 -220
rect 690 -280 860 -240
rect 1990 -280 2160 -240
rect 250 -300 2160 -280
rect 2230 -300 2530 -280
rect 2600 -300 2620 -220
rect 2880 -300 3190 -120
rect 692 -302 786 -300
rect 490 -390 500 -330
rect 560 -390 570 -330
rect 850 -350 2000 -300
rect 850 -358 1270 -350
rect 730 -390 820 -380
rect 850 -390 871 -358
rect -350 -620 -50 -440
rect 260 -427 380 -420
rect 260 -439 387 -427
rect 260 -530 347 -439
rect 260 -590 270 -530
rect 330 -590 347 -530
rect 260 -640 347 -590
rect 260 -700 270 -640
rect 330 -700 347 -640
rect 260 -750 347 -700
rect 260 -810 270 -750
rect 330 -810 347 -750
rect 260 -815 347 -810
rect 381 -815 387 -439
rect 449 -439 495 -427
rect 449 -590 455 -439
rect 420 -600 455 -590
rect 489 -590 495 -439
rect 557 -430 603 -427
rect 557 -439 700 -430
rect 489 -600 500 -590
rect 420 -660 430 -600
rect 490 -660 500 -600
rect 420 -670 455 -660
rect 260 -827 387 -815
rect 449 -815 455 -670
rect 489 -670 500 -660
rect 489 -815 495 -670
rect 449 -827 495 -815
rect 557 -815 563 -439
rect 597 -530 700 -439
rect 730 -480 740 -390
rect 810 -417 820 -390
rect 859 -392 871 -390
rect 1247 -392 1270 -358
rect 1580 -358 2000 -350
rect 859 -398 1270 -392
rect 860 -400 1270 -398
rect 1300 -390 1390 -380
rect 812 -451 820 -417
rect 810 -480 820 -451
rect 1300 -417 1310 -390
rect 1300 -451 1306 -417
rect 730 -490 820 -480
rect 859 -476 1260 -470
rect 859 -510 871 -476
rect 1247 -510 1260 -476
rect 1300 -480 1310 -451
rect 1380 -480 1390 -390
rect 1300 -490 1390 -480
rect 1460 -390 1550 -380
rect 1460 -480 1470 -390
rect 1540 -417 1550 -390
rect 1580 -392 1601 -358
rect 1977 -392 2000 -358
rect 1580 -400 2000 -392
rect 2030 -390 2110 -380
rect 2380 -390 2400 -330
rect 2460 -390 2490 -330
rect 1542 -451 1550 -417
rect 1540 -480 1550 -451
rect 2030 -417 2040 -390
rect 2030 -451 2036 -417
rect 1460 -490 1550 -480
rect 1589 -476 1990 -470
rect 859 -516 940 -510
rect 597 -590 620 -530
rect 680 -590 700 -530
rect 860 -550 940 -516
rect 1020 -550 1140 -510
rect 1220 -520 1260 -510
rect 1589 -510 1601 -476
rect 1977 -510 1990 -476
rect 2030 -480 2040 -451
rect 2100 -480 2110 -390
rect 2248 -430 2294 -427
rect 2030 -490 2110 -480
rect 2140 -439 2294 -430
rect 2140 -460 2254 -439
rect 1589 -516 1630 -510
rect 1220 -550 1470 -520
rect 860 -570 1470 -550
rect 1460 -580 1470 -570
rect 1540 -580 1550 -520
rect 1590 -540 1630 -516
rect 1710 -540 1860 -510
rect 1940 -540 1990 -510
rect 1590 -550 1990 -540
rect 2140 -540 2160 -460
rect 2230 -540 2254 -460
rect 597 -650 700 -590
rect 597 -710 620 -650
rect 680 -710 700 -650
rect 2140 -590 2254 -540
rect 2140 -670 2160 -590
rect 2230 -670 2254 -590
rect 597 -750 700 -710
rect 597 -810 620 -750
rect 680 -810 700 -750
rect 597 -815 700 -810
rect 557 -827 700 -815
rect 260 -830 380 -827
rect 600 -830 700 -827
rect 870 -700 1970 -690
rect 870 -740 990 -700
rect 1350 -740 1500 -700
rect 1870 -740 1970 -700
rect 870 -750 1970 -740
rect 870 -790 940 -750
rect 380 -920 390 -860
rect 450 -920 460 -860
rect 380 -930 460 -920
rect 500 -920 510 -860
rect 570 -920 580 -860
rect 500 -930 580 -920
rect 230 -950 340 -940
rect 230 -1010 270 -950
rect 330 -960 340 -950
rect 610 -960 630 -950
rect 330 -970 630 -960
rect 620 -1010 630 -970
rect 690 -1010 710 -950
rect 230 -1020 710 -1010
rect 870 -970 890 -790
rect 930 -970 940 -790
rect 1070 -816 1150 -790
rect 1220 -816 1270 -790
rect 870 -1070 940 -970
rect 970 -860 1040 -840
rect 1070 -850 1082 -816
rect 1258 -850 1270 -816
rect 1580 -815 1630 -780
rect 1710 -809 1780 -780
rect 1910 -790 1970 -750
rect 1710 -815 1783 -809
rect 1310 -848 1380 -830
rect 1070 -860 1270 -850
rect 1302 -860 1380 -848
rect 970 -890 998 -860
rect 1032 -894 1040 -860
rect 1030 -950 1040 -894
rect 1070 -904 1090 -890
rect 1070 -938 1082 -904
rect 1070 -950 1090 -938
rect 1260 -950 1270 -890
rect 1302 -894 1308 -860
rect 1342 -894 1380 -860
rect 1302 -906 1380 -894
rect 970 -980 1040 -950
rect 1310 -980 1380 -906
rect 970 -1020 1380 -980
rect 1470 -847 1550 -830
rect 1470 -859 1551 -847
rect 1470 -893 1511 -859
rect 1545 -893 1551 -859
rect 1580 -849 1595 -815
rect 1771 -849 1783 -815
rect 1820 -830 1880 -820
rect 1580 -855 1783 -849
rect 1580 -860 1780 -855
rect 1470 -905 1551 -893
rect 1583 -900 1783 -897
rect 1580 -903 1610 -900
rect 1750 -903 1783 -900
rect 1470 -990 1550 -905
rect 1580 -937 1595 -903
rect 1771 -937 1783 -903
rect 1815 -905 1820 -847
rect 1580 -960 1610 -937
rect 1750 -943 1783 -937
rect 1750 -960 1780 -943
rect 1820 -990 1880 -910
rect 1470 -1020 1880 -990
rect 1910 -960 1920 -790
rect 1960 -960 1970 -790
rect 2140 -710 2254 -670
rect 2140 -790 2160 -710
rect 2230 -790 2254 -710
rect 2140 -815 2254 -790
rect 2288 -815 2294 -439
rect 2356 -439 2402 -427
rect 2356 -560 2362 -439
rect 2330 -570 2362 -560
rect 2330 -690 2362 -680
rect 2140 -820 2294 -815
rect 2248 -827 2294 -820
rect 2356 -815 2362 -690
rect 2396 -815 2402 -439
rect 2356 -827 2402 -815
rect 2464 -430 2510 -427
rect 2464 -439 2620 -430
rect 2464 -815 2470 -439
rect 2504 -460 2620 -439
rect 2504 -540 2530 -460
rect 2600 -540 2620 -460
rect 2504 -590 2620 -540
rect 2504 -670 2530 -590
rect 2600 -670 2620 -590
rect 2880 -440 2920 -300
rect 3060 -440 3190 -300
rect 2880 -670 3190 -440
rect 2504 -710 2620 -670
rect 2504 -790 2530 -710
rect 2600 -790 2620 -710
rect 2504 -815 2620 -790
rect 2464 -827 2620 -815
rect 2510 -830 2620 -827
rect 2290 -920 2300 -860
rect 2360 -920 2370 -860
rect 2290 -930 2370 -920
rect 540 -1080 940 -1070
rect 540 -1120 650 -1080
rect 840 -1120 940 -1080
rect 540 -1140 940 -1120
rect 970 -1090 1390 -1060
rect 540 -1170 610 -1140
rect 430 -1180 610 -1170
rect -300 -1270 -10 -1260
rect -300 -1480 -200 -1270
rect -40 -1480 -10 -1270
rect 430 -1280 440 -1180
rect 530 -1280 560 -1180
rect 430 -1290 560 -1280
rect -300 -1700 -10 -1480
rect 540 -1740 560 -1290
rect 600 -1740 610 -1180
rect 700 -1230 710 -1170
rect 780 -1230 790 -1170
rect 970 -1176 1040 -1090
rect 970 -1210 998 -1176
rect 1032 -1210 1040 -1176
rect 1070 -1132 1100 -1120
rect 1240 -1132 1270 -1120
rect 1070 -1166 1082 -1132
rect 1258 -1166 1270 -1132
rect 1070 -1180 1100 -1166
rect 1240 -1180 1270 -1166
rect 1300 -1140 1390 -1090
rect 1300 -1176 1310 -1140
rect 970 -1250 1040 -1210
rect 1300 -1210 1308 -1176
rect 1070 -1220 1270 -1214
rect 1070 -1230 1082 -1220
rect 1258 -1230 1270 -1220
rect 668 -1270 714 -1260
rect 640 -1272 714 -1270
rect 640 -1360 674 -1272
rect 640 -1648 674 -1440
rect 708 -1648 714 -1272
rect 640 -1650 714 -1648
rect 668 -1660 714 -1650
rect 776 -1272 822 -1260
rect 776 -1648 782 -1272
rect 816 -1280 822 -1272
rect 816 -1290 860 -1280
rect 852 -1630 860 -1290
rect 1070 -1320 1080 -1230
rect 1260 -1320 1270 -1230
rect 1300 -1230 1310 -1210
rect 1380 -1230 1390 -1140
rect 1300 -1240 1390 -1230
rect 1460 -1080 1880 -1050
rect 1460 -1140 1550 -1080
rect 1460 -1240 1470 -1140
rect 1540 -1163 1550 -1140
rect 1540 -1175 1551 -1163
rect 1580 -1170 1590 -1110
rect 1770 -1125 1780 -1110
rect 1770 -1131 1783 -1125
rect 1771 -1165 1783 -1131
rect 1820 -1163 1880 -1080
rect 1910 -1070 1970 -960
rect 2140 -1020 2160 -960
rect 2220 -970 2540 -960
rect 2220 -1020 2230 -970
rect 2530 -1020 2540 -970
rect 2600 -1020 2620 -960
rect 2140 -1030 2620 -1020
rect 1910 -1080 2310 -1070
rect 1910 -1120 2020 -1080
rect 2200 -1110 2310 -1080
rect 2200 -1120 2430 -1110
rect 1910 -1140 2310 -1120
rect 1770 -1170 1783 -1165
rect 1583 -1171 1783 -1170
rect 1545 -1209 1551 -1175
rect 1540 -1221 1551 -1209
rect 1815 -1175 1880 -1163
rect 1815 -1209 1821 -1175
rect 1855 -1209 1880 -1175
rect 1583 -1219 1783 -1213
rect 1540 -1240 1550 -1221
rect 1460 -1250 1550 -1240
rect 1583 -1230 1595 -1219
rect 1771 -1230 1783 -1219
rect 1815 -1221 1880 -1209
rect 1583 -1259 1590 -1230
rect 1070 -1330 1270 -1320
rect 1780 -1259 1783 -1230
rect 1820 -1240 1880 -1221
rect 2070 -1230 2080 -1170
rect 2140 -1230 2160 -1170
rect 2240 -1180 2310 -1140
rect 2240 -1260 2260 -1180
rect 2034 -1270 2080 -1260
rect 1590 -1330 1780 -1320
rect 2010 -1272 2090 -1270
rect 2010 -1280 2040 -1272
rect 2074 -1280 2090 -1272
rect 1220 -1410 1690 -1390
rect 1220 -1441 1380 -1410
rect 1540 -1441 1690 -1410
rect 1220 -1475 1257 -1441
rect 1291 -1475 1349 -1441
rect 1567 -1475 1625 -1441
rect 1659 -1475 1690 -1441
rect 1220 -1490 1380 -1475
rect 1540 -1490 1690 -1475
rect 1220 -1510 1690 -1490
rect 816 -1640 860 -1630
rect 1040 -1620 1200 -1600
rect 816 -1648 822 -1640
rect 776 -1660 822 -1648
rect 540 -1750 610 -1740
rect 420 -1760 610 -1750
rect 710 -1760 720 -1690
rect 780 -1760 790 -1690
rect 520 -1840 610 -1760
rect 1040 -1770 1050 -1620
rect 1190 -1650 1200 -1620
rect 1600 -1611 1680 -1590
rect 1600 -1645 1625 -1611
rect 1659 -1645 1680 -1611
rect 1190 -1660 1300 -1650
rect 1190 -1680 1570 -1660
rect 1190 -1720 1260 -1680
rect 1300 -1720 1350 -1680
rect 1390 -1720 1440 -1680
rect 1480 -1720 1520 -1680
rect 1560 -1720 1570 -1680
rect 1190 -1740 1570 -1720
rect 1600 -1683 1680 -1645
rect 2010 -1640 2020 -1280
rect 2080 -1640 2090 -1280
rect 2010 -1648 2040 -1640
rect 2074 -1648 2090 -1640
rect 2010 -1650 2090 -1648
rect 2142 -1272 2260 -1260
rect 2142 -1648 2148 -1272
rect 2182 -1648 2260 -1272
rect 2142 -1650 2260 -1648
rect 2034 -1660 2080 -1650
rect 2142 -1660 2188 -1650
rect 1600 -1719 1625 -1683
rect 1659 -1719 1680 -1683
rect 1190 -1760 1300 -1740
rect 1190 -1770 1200 -1760
rect 1040 -1790 1200 -1770
rect 1600 -1763 1680 -1719
rect 2060 -1750 2080 -1690
rect 2140 -1750 2160 -1690
rect 2240 -1740 2260 -1650
rect 2300 -1230 2310 -1180
rect 2420 -1230 2430 -1120
rect 2300 -1240 2430 -1230
rect 2300 -1740 2310 -1240
rect 2880 -1310 3210 -1160
rect 2880 -1420 2890 -1310
rect 3000 -1420 3210 -1310
rect 2880 -1570 3210 -1420
rect 2240 -1750 2310 -1740
rect 1600 -1790 1625 -1763
rect 1659 -1790 1680 -1763
rect 2240 -1760 2460 -1750
rect 420 -1850 610 -1840
rect 1600 -1850 1610 -1790
rect 1670 -1850 1680 -1790
rect 1600 -1860 1680 -1850
rect 1740 -1790 1820 -1780
rect 1740 -1850 1750 -1790
rect 1810 -1850 1820 -1790
rect 2240 -1840 2330 -1760
rect 2450 -1840 2460 -1760
rect 2240 -1850 2460 -1840
rect 1740 -1860 1820 -1850
rect 1740 -1930 1820 -1920
rect 1740 -1950 1750 -1930
rect 1220 -1985 1750 -1950
rect 1810 -1950 1820 -1930
rect 1220 -2019 1257 -1985
rect 1291 -2019 1349 -1985
rect 1383 -2019 1441 -1985
rect 1475 -2019 1533 -1985
rect 1567 -2019 1625 -1985
rect 1659 -2019 1750 -1985
rect 1220 -2050 1750 -2019
rect 1810 -2050 1870 -1950
rect 1220 -2061 1870 -2050
rect 1220 -2095 1257 -2061
rect 1291 -2095 1349 -2061
rect 1383 -2095 1441 -2061
rect 1475 -2095 1533 -2061
rect 1567 -2095 1625 -2061
rect 1659 -2070 1870 -2061
rect 1659 -2095 1750 -2070
rect 1220 -2130 1750 -2095
rect 1810 -2130 1870 -2070
rect 1740 -2140 1820 -2130
rect 1740 -2210 1820 -2200
rect 1740 -2270 1750 -2210
rect 1810 -2270 1820 -2210
rect 1740 -2280 1820 -2270
rect 1610 -2294 1690 -2280
rect 1610 -2329 1625 -2294
rect 1659 -2329 1690 -2294
rect 1110 -2350 1580 -2340
rect 810 -2520 1040 -2350
rect 1110 -2440 1120 -2350
rect 1230 -2360 1580 -2350
rect 1230 -2400 1260 -2360
rect 1300 -2400 1350 -2360
rect 1390 -2400 1440 -2360
rect 1480 -2400 1520 -2360
rect 1560 -2400 1580 -2360
rect 1230 -2440 1580 -2400
rect 1110 -2450 1580 -2440
rect 1610 -2367 1690 -2329
rect 1610 -2402 1625 -2367
rect 1659 -2370 1690 -2367
rect 1659 -2402 2040 -2370
rect 1610 -2440 2040 -2402
rect 2140 -2440 2170 -2370
rect 1610 -2443 2170 -2440
rect 1610 -2478 1624 -2443
rect 1658 -2478 2170 -2443
rect 1610 -2490 2170 -2478
rect 810 -2660 820 -2520
rect 1000 -2660 1040 -2520
rect 810 -2780 1040 -2660
rect 1080 -2510 1200 -2490
rect 1610 -2491 1690 -2490
rect 1080 -2680 1100 -2510
rect 1180 -2570 1200 -2510
rect 1180 -2590 1690 -2570
rect 1180 -2605 1350 -2590
rect 1560 -2605 1690 -2590
rect 1180 -2639 1257 -2605
rect 1291 -2639 1349 -2605
rect 1567 -2639 1625 -2605
rect 1659 -2639 1690 -2605
rect 1180 -2670 1350 -2639
rect 1560 -2670 1690 -2639
rect 1180 -2680 1690 -2670
rect 1080 -2700 1200 -2680
<< via1 >>
rect 1380 -50 1540 110
rect -230 -440 -70 -280
rect 270 -240 330 -220
rect 270 -280 320 -240
rect 320 -280 330 -240
rect 630 -280 690 -220
rect 2530 -240 2600 -220
rect 2160 -280 2210 -240
rect 2210 -280 2230 -240
rect 2530 -280 2600 -240
rect 2160 -300 2230 -280
rect 2530 -300 2600 -280
rect 500 -346 560 -330
rect 500 -380 509 -346
rect 509 -380 543 -346
rect 543 -380 560 -346
rect 500 -390 560 -380
rect 270 -590 330 -530
rect 270 -700 330 -640
rect 270 -810 330 -750
rect 430 -660 455 -600
rect 455 -660 489 -600
rect 489 -660 490 -600
rect 740 -417 810 -390
rect 740 -451 778 -417
rect 778 -451 810 -417
rect 740 -480 810 -451
rect 1310 -417 1380 -390
rect 1310 -451 1340 -417
rect 1340 -451 1380 -417
rect 940 -510 1020 -490
rect 1140 -510 1220 -490
rect 1310 -480 1380 -451
rect 1470 -417 1540 -390
rect 2400 -346 2460 -330
rect 2400 -380 2416 -346
rect 2416 -380 2450 -346
rect 2450 -380 2460 -346
rect 2400 -390 2460 -380
rect 1470 -451 1508 -417
rect 1508 -451 1540 -417
rect 1470 -480 1540 -451
rect 2040 -417 2100 -390
rect 2040 -451 2070 -417
rect 2070 -451 2100 -417
rect 620 -590 680 -530
rect 940 -550 1020 -510
rect 1140 -550 1220 -510
rect 1630 -510 1710 -480
rect 1860 -510 1940 -480
rect 2040 -480 2100 -451
rect 1470 -580 1540 -520
rect 1630 -540 1710 -510
rect 1860 -540 1940 -510
rect 2160 -540 2230 -460
rect 620 -710 680 -650
rect 2160 -670 2230 -590
rect 620 -810 680 -750
rect 390 -874 450 -860
rect 390 -908 401 -874
rect 401 -908 435 -874
rect 435 -908 450 -874
rect 390 -920 450 -908
rect 510 -920 570 -860
rect 270 -1010 330 -950
rect 630 -1010 690 -950
rect 1150 -816 1220 -790
rect 1150 -850 1220 -816
rect 1630 -815 1710 -780
rect 970 -894 998 -890
rect 998 -894 1030 -890
rect 970 -950 1030 -894
rect 1090 -904 1260 -890
rect 1090 -938 1258 -904
rect 1258 -938 1260 -904
rect 1090 -950 1260 -938
rect 1630 -840 1710 -815
rect 1610 -903 1750 -900
rect 1610 -937 1750 -903
rect 1820 -859 1880 -830
rect 1820 -893 1821 -859
rect 1821 -893 1855 -859
rect 1855 -893 1880 -859
rect 1610 -960 1750 -937
rect 1820 -910 1880 -893
rect 2160 -790 2230 -710
rect 2330 -680 2362 -570
rect 2362 -680 2390 -570
rect 2530 -540 2600 -460
rect 2530 -670 2600 -590
rect 2920 -440 3060 -300
rect 2530 -790 2600 -710
rect 2300 -874 2360 -860
rect 2300 -908 2308 -874
rect 2308 -908 2342 -874
rect 2342 -908 2360 -874
rect 2300 -920 2360 -908
rect -200 -1480 -40 -1270
rect 440 -1280 530 -1180
rect 710 -1188 780 -1170
rect 710 -1222 728 -1188
rect 728 -1222 762 -1188
rect 762 -1222 780 -1188
rect 710 -1230 780 -1222
rect 1100 -1132 1240 -1120
rect 1100 -1166 1240 -1132
rect 1100 -1180 1240 -1166
rect 1310 -1176 1380 -1140
rect 1310 -1210 1342 -1176
rect 1342 -1210 1380 -1176
rect 640 -1440 674 -1360
rect 674 -1440 700 -1360
rect 800 -1630 816 -1290
rect 816 -1630 852 -1290
rect 1080 -1254 1082 -1230
rect 1082 -1254 1258 -1230
rect 1258 -1254 1260 -1230
rect 1080 -1320 1260 -1254
rect 1310 -1230 1380 -1210
rect 1470 -1175 1540 -1140
rect 1590 -1131 1770 -1110
rect 1590 -1165 1595 -1131
rect 1595 -1165 1770 -1131
rect 2160 -1020 2220 -960
rect 2540 -1020 2600 -960
rect 1590 -1170 1770 -1165
rect 1470 -1209 1511 -1175
rect 1511 -1209 1540 -1175
rect 1470 -1240 1540 -1209
rect 1590 -1253 1595 -1230
rect 1595 -1253 1771 -1230
rect 1771 -1253 1780 -1230
rect 1590 -1320 1780 -1253
rect 2080 -1188 2140 -1170
rect 2080 -1222 2094 -1188
rect 2094 -1222 2128 -1188
rect 2128 -1222 2140 -1188
rect 2080 -1230 2140 -1222
rect 1380 -1441 1540 -1410
rect 1380 -1475 1383 -1441
rect 1383 -1475 1441 -1441
rect 1441 -1475 1475 -1441
rect 1475 -1475 1533 -1441
rect 1533 -1475 1540 -1441
rect 1380 -1490 1540 -1475
rect 720 -1698 780 -1690
rect 720 -1732 728 -1698
rect 728 -1732 762 -1698
rect 762 -1732 780 -1698
rect 720 -1760 780 -1732
rect 420 -1840 520 -1760
rect 1050 -1770 1190 -1620
rect 2020 -1640 2040 -1280
rect 2040 -1640 2074 -1280
rect 2074 -1640 2080 -1280
rect 2080 -1698 2140 -1690
rect 2080 -1732 2094 -1698
rect 2094 -1732 2128 -1698
rect 2128 -1732 2140 -1698
rect 2080 -1750 2140 -1732
rect 2310 -1230 2420 -1120
rect 2890 -1420 3000 -1310
rect 1610 -1798 1625 -1790
rect 1625 -1798 1659 -1790
rect 1659 -1798 1670 -1790
rect 1610 -1850 1670 -1798
rect 1750 -1800 1810 -1790
rect 1750 -1840 1760 -1800
rect 1760 -1840 1800 -1800
rect 1800 -1840 1810 -1800
rect 1750 -1850 1810 -1840
rect 2330 -1840 2450 -1760
rect 1750 -1940 1810 -1930
rect 1750 -1980 1760 -1940
rect 1760 -1980 1800 -1940
rect 1800 -1980 1810 -1940
rect 1750 -2050 1810 -1980
rect 1750 -2080 1810 -2070
rect 1750 -2120 1760 -2080
rect 1760 -2120 1800 -2080
rect 1800 -2120 1810 -2080
rect 1750 -2130 1810 -2120
rect 1750 -2220 1810 -2210
rect 1750 -2260 1760 -2220
rect 1760 -2260 1800 -2220
rect 1800 -2260 1810 -2220
rect 1750 -2270 1810 -2260
rect 1120 -2440 1230 -2350
rect 2040 -2440 2140 -2370
rect 820 -2660 1000 -2520
rect 1350 -2605 1560 -2590
rect 1350 -2639 1383 -2605
rect 1383 -2639 1441 -2605
rect 1441 -2639 1475 -2605
rect 1475 -2639 1533 -2605
rect 1533 -2639 1560 -2605
rect 1350 -2670 1560 -2639
<< metal2 >>
rect 140 200 700 290
rect 140 -130 230 200
rect 590 -130 700 200
rect 1290 130 1640 170
rect 1290 -70 1360 130
rect 1560 -70 1640 130
rect 1290 -110 1640 -70
rect 140 -210 700 -130
rect 250 -220 340 -210
rect -250 -280 -50 -260
rect -250 -440 -230 -280
rect -70 -440 -50 -280
rect -250 -460 -50 -440
rect 10 -310 160 -270
rect 10 -420 30 -310
rect 140 -420 160 -310
rect -210 -650 -30 -630
rect -210 -730 -190 -650
rect -50 -730 -30 -650
rect -210 -1270 -30 -730
rect -210 -1480 -200 -1270
rect -40 -1480 -30 -1270
rect -210 -1490 -30 -1480
rect 10 -830 160 -420
rect 10 -930 40 -830
rect 140 -930 160 -830
rect 10 -2370 160 -930
rect 250 -280 270 -220
rect 330 -280 340 -220
rect 250 -530 340 -280
rect 610 -220 700 -210
rect 610 -280 630 -220
rect 690 -280 700 -220
rect 490 -320 570 -310
rect 490 -390 500 -320
rect 560 -390 570 -320
rect 500 -400 560 -390
rect 250 -590 270 -530
rect 330 -590 340 -530
rect 250 -640 340 -590
rect 250 -700 270 -640
rect 330 -700 340 -640
rect 420 -600 490 -590
rect 420 -660 430 -600
rect 420 -670 490 -660
rect 250 -750 340 -700
rect 250 -810 270 -750
rect 330 -810 340 -750
rect 250 -950 340 -810
rect 520 -850 560 -400
rect 610 -530 700 -280
rect 2150 -210 2650 290
rect 2150 -240 2240 -210
rect 2150 -300 2160 -240
rect 2230 -300 2240 -240
rect 730 -390 820 -380
rect 730 -480 740 -390
rect 810 -480 820 -390
rect 1300 -390 1390 -380
rect 1300 -480 1310 -390
rect 1380 -480 1390 -390
rect 730 -490 820 -480
rect 920 -490 1030 -480
rect 610 -590 620 -530
rect 680 -590 700 -530
rect 610 -650 700 -590
rect 610 -710 620 -650
rect 680 -710 700 -650
rect 920 -550 940 -490
rect 1020 -550 1030 -490
rect 920 -600 1030 -550
rect 920 -680 930 -600
rect 1020 -680 1030 -600
rect 920 -690 1030 -680
rect 1130 -490 1240 -480
rect 1130 -550 1140 -490
rect 1220 -550 1240 -490
rect 1130 -600 1240 -550
rect 1130 -670 1140 -600
rect 1230 -670 1240 -600
rect 610 -750 700 -710
rect 610 -810 620 -750
rect 680 -810 700 -750
rect 380 -860 470 -850
rect 380 -920 390 -860
rect 450 -920 470 -860
rect 380 -930 470 -920
rect 500 -860 580 -850
rect 500 -920 510 -860
rect 570 -920 580 -860
rect 500 -930 580 -920
rect 250 -960 270 -950
rect 230 -1010 270 -960
rect 330 -960 340 -950
rect 610 -950 700 -810
rect 1130 -790 1240 -670
rect 610 -960 630 -950
rect 330 -1010 630 -960
rect 690 -960 700 -950
rect 950 -890 1060 -840
rect 1130 -850 1150 -790
rect 1220 -850 1240 -790
rect 1300 -630 1390 -480
rect 1300 -690 1330 -630
rect 950 -950 970 -890
rect 1030 -950 1060 -890
rect 950 -960 1060 -950
rect 1090 -890 1270 -880
rect 1260 -950 1270 -890
rect 690 -1010 710 -960
rect 230 -1020 710 -1010
rect 1090 -1120 1260 -950
rect 710 -1170 780 -1160
rect 430 -1180 540 -1170
rect 430 -1280 440 -1180
rect 530 -1280 540 -1180
rect 1080 -1180 1100 -1120
rect 1240 -1180 1260 -1120
rect 1300 -1140 1390 -690
rect 710 -1240 780 -1230
rect 1070 -1230 1270 -1220
rect 430 -1290 540 -1280
rect 610 -1360 700 -1350
rect 610 -1440 620 -1360
rect 610 -1450 700 -1440
rect 730 -1670 760 -1240
rect 790 -1290 860 -1280
rect 790 -1630 800 -1290
rect 1070 -1320 1080 -1230
rect 1260 -1320 1270 -1230
rect 1300 -1230 1310 -1140
rect 1380 -1230 1390 -1140
rect 1300 -1250 1390 -1230
rect 1460 -390 1550 -380
rect 1460 -480 1470 -390
rect 1540 -480 1550 -390
rect 2030 -390 2110 -380
rect 1460 -520 1550 -480
rect 1460 -580 1470 -520
rect 1540 -580 1550 -520
rect 1460 -1140 1550 -580
rect 1610 -480 1730 -470
rect 1610 -540 1630 -480
rect 1710 -540 1730 -480
rect 1610 -580 1730 -540
rect 1610 -680 1620 -580
rect 1710 -680 1730 -580
rect 1610 -780 1730 -680
rect 1840 -480 1960 -470
rect 1840 -540 1860 -480
rect 1940 -540 1960 -480
rect 2030 -480 2040 -390
rect 2100 -480 2110 -390
rect 2030 -490 2110 -480
rect 2150 -460 2240 -300
rect 2520 -220 2610 -210
rect 2520 -300 2530 -220
rect 2600 -300 2610 -220
rect 2380 -330 2490 -320
rect 2380 -390 2400 -330
rect 2460 -390 2490 -330
rect 2410 -400 2470 -390
rect 1840 -580 1960 -540
rect 1840 -680 1860 -580
rect 1950 -680 1960 -580
rect 2150 -540 2160 -460
rect 2230 -540 2240 -460
rect 2150 -590 2240 -540
rect 1840 -690 1960 -680
rect 2000 -630 2090 -620
rect 2000 -690 2020 -630
rect 2080 -690 2090 -630
rect 1610 -840 1630 -780
rect 1710 -840 1730 -780
rect 1610 -850 1730 -840
rect 1800 -830 1890 -820
rect 1580 -960 1610 -900
rect 1750 -960 1770 -900
rect 1800 -910 1810 -830
rect 1880 -910 1890 -830
rect 1800 -920 1890 -910
rect 1580 -970 1770 -960
rect 1590 -1110 1770 -970
rect 1460 -1240 1470 -1140
rect 1540 -1240 1550 -1140
rect 1580 -1170 1590 -1110
rect 1770 -1170 1780 -1110
rect 1580 -1180 1780 -1170
rect 2000 -1130 2090 -690
rect 2150 -670 2160 -590
rect 2230 -670 2240 -590
rect 2150 -710 2240 -670
rect 2330 -570 2390 -560
rect 2330 -690 2390 -680
rect 2150 -790 2160 -710
rect 2230 -790 2240 -710
rect 2150 -960 2240 -790
rect 2420 -850 2470 -400
rect 2520 -460 2610 -300
rect 2890 -280 3090 -270
rect 2520 -540 2530 -460
rect 2600 -540 2610 -460
rect 2520 -590 2610 -540
rect 2520 -670 2530 -590
rect 2600 -670 2610 -590
rect 2520 -710 2610 -670
rect 2520 -790 2530 -710
rect 2600 -790 2610 -710
rect 2290 -860 2370 -850
rect 2360 -920 2370 -860
rect 2290 -930 2370 -920
rect 2400 -860 2490 -850
rect 2400 -920 2410 -860
rect 2470 -920 2490 -860
rect 2400 -930 2490 -920
rect 2520 -960 2610 -790
rect 2690 -330 2840 -320
rect 2690 -390 2740 -330
rect 2810 -390 2840 -330
rect 2690 -860 2840 -390
rect 2890 -460 2900 -280
rect 3080 -460 3090 -280
rect 2890 -470 3090 -460
rect 2690 -920 2740 -860
rect 2810 -920 2840 -860
rect 2140 -1020 2160 -960
rect 2220 -1020 2540 -960
rect 2600 -1020 2620 -960
rect 2140 -1030 2620 -1020
rect 2300 -1120 2430 -1110
rect 1460 -1250 1550 -1240
rect 1580 -1230 1790 -1220
rect 1070 -1330 1270 -1320
rect 1580 -1320 1590 -1230
rect 1780 -1320 1790 -1230
rect 1580 -1330 1790 -1320
rect 2000 -1260 2040 -1130
rect 2070 -1170 2150 -1160
rect 2070 -1230 2080 -1170
rect 2140 -1230 2150 -1170
rect 2300 -1230 2310 -1120
rect 2420 -1230 2430 -1120
rect 2300 -1240 2430 -1230
rect 2000 -1280 2090 -1260
rect 1340 -1410 1580 -1390
rect 1340 -1490 1380 -1410
rect 1540 -1490 1580 -1410
rect 1340 -1510 1580 -1490
rect 790 -1640 860 -1630
rect 1040 -1620 1200 -1600
rect 710 -1690 790 -1670
rect 410 -1760 530 -1750
rect 410 -1840 420 -1760
rect 520 -1840 530 -1760
rect 410 -1850 530 -1840
rect 710 -1760 720 -1690
rect 780 -1760 790 -1690
rect 710 -1860 790 -1760
rect 1040 -1770 1050 -1620
rect 1190 -1770 1200 -1620
rect 2000 -1640 2020 -1280
rect 2080 -1640 2090 -1280
rect 2000 -1650 2090 -1640
rect 2690 -1580 2840 -920
rect 2880 -1310 3010 -1300
rect 2880 -1420 2890 -1310
rect 3000 -1420 3010 -1310
rect 2880 -1430 3010 -1420
rect 1040 -1790 1200 -1770
rect 2030 -1690 2170 -1680
rect 2030 -1750 2080 -1690
rect 2140 -1750 2170 -1690
rect 2690 -1720 2700 -1580
rect 2830 -1720 2840 -1580
rect 2690 -1730 2840 -1720
rect 1740 -1790 1820 -1780
rect 1600 -1850 1610 -1790
rect 1670 -1850 1680 -1790
rect 1600 -1860 1680 -1850
rect 1740 -1850 1750 -1790
rect 1810 -1850 1820 -1790
rect 700 -1870 810 -1860
rect 700 -1940 710 -1870
rect 790 -1940 810 -1870
rect 700 -1950 810 -1940
rect 1740 -1930 1820 -1850
rect 1740 -2050 1750 -1930
rect 1810 -2050 1820 -1930
rect 1740 -2070 1820 -2050
rect 1740 -2130 1750 -2070
rect 1810 -2130 1820 -2070
rect 1740 -2210 1820 -2130
rect 1740 -2270 1750 -2210
rect 1810 -2270 1820 -2210
rect 1740 -2280 1820 -2270
rect 10 -2440 20 -2370
rect 150 -2440 160 -2370
rect 10 -2450 160 -2440
rect 1110 -2350 1240 -2340
rect 1110 -2440 1120 -2350
rect 1230 -2440 1240 -2350
rect 1110 -2450 1240 -2440
rect 810 -2520 1010 -2500
rect 810 -2660 820 -2520
rect 1000 -2660 1010 -2520
rect 810 -2680 1010 -2660
rect 1340 -2590 1570 -2580
rect 1340 -2670 1350 -2590
rect 1560 -2670 1570 -2590
rect 1340 -2680 1570 -2670
rect 1720 -2650 1870 -2280
rect 2030 -2370 2170 -1750
rect 2310 -1760 2460 -1750
rect 2310 -1840 2330 -1760
rect 2450 -1840 2460 -1760
rect 2310 -1850 2460 -1840
rect 2030 -2440 2040 -2370
rect 2140 -2440 2170 -2370
rect 2030 -2460 2170 -2440
rect 1720 -2770 1730 -2650
rect 1860 -2770 1870 -2650
rect 1720 -2800 1870 -2770
<< via2 >>
rect 230 -130 590 200
rect 1360 110 1560 130
rect 1360 -50 1380 110
rect 1380 -50 1540 110
rect 1540 -50 1560 110
rect 1360 -70 1560 -50
rect -230 -440 -70 -280
rect 30 -420 140 -310
rect -190 -730 -50 -650
rect -180 -1440 -60 -1360
rect 40 -930 140 -830
rect 500 -330 560 -320
rect 500 -380 560 -330
rect 430 -660 490 -600
rect 740 -480 810 -390
rect 1310 -480 1380 -390
rect 930 -680 1020 -600
rect 1140 -670 1230 -600
rect 390 -920 450 -860
rect 510 -920 570 -860
rect 1330 -690 1390 -630
rect 970 -950 1030 -890
rect 440 -1280 530 -1180
rect 620 -1440 640 -1360
rect 640 -1440 700 -1360
rect 800 -1630 852 -1290
rect 852 -1630 860 -1290
rect 1080 -1320 1260 -1230
rect 1470 -480 1540 -390
rect 1620 -680 1710 -580
rect 2040 -480 2100 -390
rect 2400 -390 2460 -330
rect 1860 -680 1950 -580
rect 2020 -690 2080 -630
rect 1810 -910 1820 -830
rect 1820 -910 1880 -830
rect 2330 -680 2390 -570
rect 2290 -920 2300 -860
rect 2300 -920 2360 -860
rect 2410 -920 2470 -860
rect 2740 -390 2810 -330
rect 2900 -300 3080 -280
rect 2900 -440 2920 -300
rect 2920 -440 3060 -300
rect 3060 -440 3080 -300
rect 2900 -460 3080 -440
rect 2740 -920 2810 -860
rect 1590 -1320 1780 -1230
rect 2310 -1230 2420 -1120
rect 1380 -1490 1540 -1410
rect 420 -1840 520 -1760
rect 1050 -1770 1190 -1620
rect 2020 -1420 2080 -1310
rect 2890 -1420 3000 -1310
rect 2700 -1720 2830 -1580
rect 1610 -1850 1670 -1790
rect 710 -1940 790 -1870
rect 20 -2440 150 -2370
rect 1120 -2440 1230 -2350
rect 820 -2660 1000 -2520
rect 1350 -2670 1560 -2590
rect 2330 -1840 2450 -1760
rect 1730 -2770 1860 -2650
<< metal3 >>
rect 140 200 700 290
rect 140 -130 230 200
rect 590 -130 700 200
rect 1290 130 1640 170
rect 1290 -70 1360 130
rect 1560 -70 1640 130
rect 1290 -110 1640 -70
rect 140 -210 700 -130
rect 2150 -210 2650 290
rect -250 -270 -50 -260
rect -250 -280 200 -270
rect -250 -440 -230 -280
rect -70 -310 200 -280
rect 2890 -280 3090 -270
rect -70 -420 30 -310
rect 140 -320 570 -310
rect 2890 -320 2900 -280
rect 140 -380 500 -320
rect 560 -380 570 -320
rect 2380 -330 2900 -320
rect 140 -400 570 -380
rect 730 -390 1390 -380
rect 140 -420 200 -400
rect -70 -440 200 -420
rect -250 -450 200 -440
rect -250 -460 -50 -450
rect 730 -480 740 -390
rect 810 -480 1310 -390
rect 1380 -480 1390 -390
rect 730 -490 1390 -480
rect 1460 -390 2110 -380
rect 1460 -480 1470 -390
rect 1540 -480 2040 -390
rect 2100 -480 2110 -390
rect 2380 -390 2400 -330
rect 2460 -390 2740 -330
rect 2810 -390 2900 -330
rect 2380 -400 2900 -390
rect 2650 -440 2900 -400
rect 2890 -460 2900 -440
rect 3080 -460 3090 -280
rect 2890 -470 3090 -460
rect 1460 -490 2110 -480
rect 1590 -570 2400 -550
rect 1590 -580 2330 -570
rect 180 -600 1260 -580
rect 180 -630 430 -600
rect -250 -650 430 -630
rect -250 -730 -190 -650
rect -50 -660 430 -650
rect 490 -660 930 -600
rect -50 -680 930 -660
rect 1020 -670 1140 -600
rect 1230 -670 1260 -600
rect 1590 -620 1620 -580
rect 1020 -680 1260 -670
rect 1320 -630 1620 -620
rect -50 -730 230 -680
rect 920 -690 1030 -680
rect 1320 -690 1330 -630
rect 1390 -680 1620 -630
rect 1710 -680 1860 -580
rect 1950 -630 2330 -580
rect 1950 -680 2020 -630
rect 1390 -690 2020 -680
rect 2080 -680 2330 -630
rect 2390 -680 2400 -570
rect 2080 -690 2400 -680
rect 1320 -700 1730 -690
rect 2000 -700 2400 -690
rect -250 -740 230 -730
rect 0 -830 200 -820
rect 1800 -830 2820 -820
rect 0 -930 40 -830
rect 140 -850 200 -830
rect 140 -860 580 -850
rect 140 -920 390 -860
rect 450 -920 510 -860
rect 570 -920 580 -860
rect 980 -880 1370 -830
rect 140 -930 580 -920
rect 950 -890 1370 -880
rect 0 -1050 200 -930
rect 950 -950 970 -890
rect 1030 -910 1370 -890
rect 1800 -910 1810 -830
rect 1880 -860 2820 -830
rect 1880 -910 2290 -860
rect 1030 -950 1040 -910
rect 1800 -920 1890 -910
rect 2280 -920 2290 -910
rect 2360 -920 2410 -860
rect 2470 -920 2740 -860
rect 2810 -920 2820 -860
rect 2280 -930 2820 -920
rect 950 -1050 1040 -950
rect 0 -1110 1040 -1050
rect 2300 -1120 2430 -1110
rect 430 -1180 540 -1170
rect -300 -1350 -10 -1260
rect 430 -1280 440 -1180
rect 530 -1280 540 -1180
rect 1070 -1230 1270 -1220
rect 430 -1290 540 -1280
rect 790 -1290 880 -1280
rect -300 -1360 710 -1350
rect -300 -1440 -180 -1360
rect -60 -1440 620 -1360
rect 700 -1440 710 -1360
rect -300 -1450 710 -1440
rect -300 -1700 -10 -1450
rect 790 -1630 800 -1290
rect 870 -1630 880 -1290
rect 1070 -1320 1080 -1230
rect 1260 -1320 1270 -1230
rect 1070 -1330 1270 -1320
rect 1580 -1230 1790 -1220
rect 1580 -1320 1590 -1230
rect 1780 -1320 1790 -1230
rect 2300 -1230 2310 -1120
rect 2420 -1230 2430 -1120
rect 2300 -1240 2430 -1230
rect 1580 -1330 1790 -1320
rect 2010 -1310 3010 -1300
rect 1340 -1410 1580 -1390
rect 1340 -1490 1380 -1410
rect 1540 -1490 1580 -1410
rect 2010 -1420 2020 -1310
rect 2080 -1420 2890 -1310
rect 3000 -1420 3010 -1310
rect 2010 -1430 3010 -1420
rect 1340 -1510 1580 -1490
rect 2570 -1580 2850 -1570
rect 2570 -1600 2700 -1580
rect 790 -1640 880 -1630
rect 1040 -1620 2700 -1600
rect 410 -1760 530 -1750
rect 410 -1840 420 -1760
rect 520 -1840 530 -1760
rect 410 -1850 530 -1840
rect 710 -1860 790 -1700
rect 1040 -1770 1050 -1620
rect 1190 -1690 2700 -1620
rect 1190 -1770 1200 -1690
rect 1610 -1720 1670 -1690
rect 2570 -1720 2700 -1690
rect 2830 -1720 2850 -1580
rect 2570 -1730 2850 -1720
rect 1040 -1790 1200 -1770
rect 2310 -1760 2460 -1750
rect 1600 -1790 1680 -1780
rect 1600 -1850 1610 -1790
rect 1670 -1850 1680 -1790
rect 2310 -1840 2330 -1760
rect 2450 -1840 2460 -1760
rect 2310 -1850 2460 -1840
rect 700 -1870 810 -1860
rect 1600 -1870 1680 -1850
rect 700 -1940 710 -1870
rect 790 -1940 1680 -1870
rect 700 -1950 810 -1940
rect 10 -2350 1240 -2340
rect 10 -2370 1120 -2350
rect 10 -2440 20 -2370
rect 150 -2440 1120 -2370
rect 1230 -2440 1240 -2350
rect 10 -2450 1240 -2440
rect 810 -2520 1010 -2510
rect 810 -2660 820 -2520
rect 1000 -2660 1010 -2520
rect 810 -2670 1010 -2660
rect 1340 -2570 1570 -2560
rect 1340 -2590 1360 -2570
rect 1340 -2670 1350 -2590
rect 1560 -2670 1570 -2570
rect 1340 -2680 1570 -2670
rect 1720 -2650 1870 -2640
rect 1720 -2770 1730 -2650
rect 1860 -2770 1870 -2650
rect 1720 -2800 1870 -2770
rect 1640 -2810 1870 -2800
rect 1640 -3010 1670 -2810
rect 1840 -3010 1870 -2810
rect 1640 -3040 1870 -3010
<< via3 >>
rect 230 -130 590 200
rect 1360 -70 1560 130
rect 440 -1280 530 -1180
rect 800 -1630 860 -1290
rect 860 -1630 870 -1290
rect 1080 -1320 1260 -1230
rect 1590 -1320 1780 -1230
rect 2310 -1230 2420 -1120
rect 1380 -1490 1540 -1410
rect 420 -1840 520 -1760
rect 2330 -1840 2450 -1760
rect 820 -2660 1000 -2520
rect 1360 -2590 1560 -2570
rect 1360 -2640 1560 -2590
rect 1670 -3010 1840 -2810
<< metal4 >>
rect 140 200 700 290
rect 140 -130 230 200
rect 590 -130 700 200
rect 2150 200 2650 290
rect 140 -210 700 -130
rect 2150 -130 2230 200
rect 2590 -130 2650 200
rect 2150 -210 2650 -130
rect 940 -980 2070 -970
rect 770 -1090 2070 -980
rect 770 -1140 890 -1090
rect 430 -1180 890 -1140
rect 430 -1280 440 -1180
rect 530 -1260 890 -1180
rect 1340 -1220 1580 -1090
rect 1950 -1110 2070 -1090
rect 1950 -1120 2430 -1110
rect 530 -1280 540 -1260
rect 430 -1290 540 -1280
rect 770 -1290 890 -1260
rect 770 -1630 800 -1290
rect 870 -1630 890 -1290
rect 1050 -1230 1790 -1220
rect 1050 -1320 1080 -1230
rect 1260 -1320 1590 -1230
rect 1780 -1320 1790 -1230
rect 1050 -1340 1790 -1320
rect 1950 -1230 2310 -1120
rect 2420 -1230 2430 -1120
rect 1950 -1240 2430 -1230
rect 770 -1750 890 -1630
rect 410 -1760 890 -1750
rect 410 -1840 420 -1760
rect 520 -1840 890 -1760
rect 410 -1850 890 -1840
rect 1340 -1410 1580 -1340
rect 1340 -1490 1380 -1410
rect 1540 -1490 1580 -1410
rect 1340 -2500 1580 -1490
rect 1950 -1750 2070 -1240
rect 1950 -1760 2460 -1750
rect 1950 -1840 2330 -1760
rect 2450 -1840 2460 -1760
rect 1950 -1850 2460 -1840
rect 810 -2520 1580 -2500
rect 810 -2660 820 -2520
rect 1000 -2570 1580 -2520
rect 1000 -2640 1360 -2570
rect 1560 -2640 1690 -2570
rect 1000 -2660 1690 -2640
rect 810 -2680 1690 -2660
rect 1560 -2760 1870 -2740
rect 1800 -2810 1870 -2760
rect 1560 -3010 1670 -3000
rect 1840 -3010 1870 -2810
rect 1560 -3040 1870 -3010
<< via4 >>
rect 230 -130 590 200
rect 1290 130 1640 170
rect 1290 -70 1360 130
rect 1360 -70 1560 130
rect 1560 -70 1640 130
rect 1290 -110 1640 -70
rect 2230 -130 2590 200
rect 1560 -2810 1800 -2760
rect 1560 -3000 1670 -2810
rect 1670 -3000 1800 -2810
<< metal5 >>
rect 140 200 2650 290
rect 140 -130 230 200
rect 590 170 2230 200
rect 590 -110 1290 170
rect 1640 -110 2230 170
rect 590 -130 2230 -110
rect 2590 -130 2650 200
rect 140 -210 2650 -130
rect 1190 -2760 1880 -210
rect 1190 -3000 1560 -2760
rect 1800 -3000 1880 -2760
rect 1190 -3040 1880 -3000
<< labels >>
flabel metal1 1360 -70 1560 130 0 FreeSans 256 0 0 0 VDD
port 0 nsew
flabel metal1 810 -2680 1010 -2480 0 FreeSans 256 0 0 0 GND
port 5 nsew
flabel metal1 -220 -1700 -20 -1500 0 FreeSans 256 0 0 0 Q
port 4 nsew
flabel metal1 2890 -470 3090 -270 0 FreeSans 256 0 0 0 R
port 2 nsew
flabel metal1 3010 -1470 3210 -1270 0 FreeSans 256 0 0 0 QN
port 3 nsew
flabel metal1 -250 -460 -50 -260 0 FreeSans 256 0 0 0 S
port 1 nsew
flabel locali 1625 -1645 1659 -1611 0 FreeSans 340 0 0 0 x1.Y
flabel locali 1625 -1713 1659 -1679 0 FreeSans 340 0 0 0 x1.Y
flabel locali 1625 -1781 1659 -1747 0 FreeSans 340 0 0 0 x1.Y
flabel locali 1257 -1713 1291 -1679 0 FreeSans 340 0 0 0 x1.A
flabel locali 1349 -1713 1383 -1679 0 FreeSans 340 0 0 0 x1.A
flabel locali 1441 -1713 1475 -1679 0 FreeSans 340 0 0 0 x1.A
flabel locali 1533 -1713 1567 -1679 0 FreeSans 340 0 0 0 x1.A
flabel nwell 1257 -2019 1291 -1985 0 FreeSans 200 0 0 0 x1.VPB
flabel pwell 1257 -1475 1291 -1441 0 FreeSans 200 0 0 0 x1.VNB
flabel metal1 1257 -2019 1291 -1985 0 FreeSans 200 0 0 0 x1.VPWR
flabel metal1 1257 -1475 1291 -1441 0 FreeSans 200 0 0 0 x1.VGND
rlabel comment 1228 -1458 1228 -1458 2 x1.inv_4
rlabel metal1 1228 -1506 1688 -1410 5 x1.VGND
rlabel metal1 1228 -2050 1688 -1954 5 x1.VPWR
flabel locali 1625 -2469 1659 -2435 0 FreeSans 340 0 0 0 x2.Y
flabel locali 1625 -2401 1659 -2367 0 FreeSans 340 0 0 0 x2.Y
flabel locali 1625 -2333 1659 -2299 0 FreeSans 340 0 0 0 x2.Y
flabel locali 1257 -2401 1291 -2367 0 FreeSans 340 0 0 0 x2.A
flabel locali 1349 -2401 1383 -2367 0 FreeSans 340 0 0 0 x2.A
flabel locali 1441 -2401 1475 -2367 0 FreeSans 340 0 0 0 x2.A
flabel locali 1533 -2401 1567 -2367 0 FreeSans 340 0 0 0 x2.A
flabel nwell 1257 -2095 1291 -2061 0 FreeSans 200 0 0 0 x2.VPB
flabel pwell 1257 -2639 1291 -2605 0 FreeSans 200 0 0 0 x2.VNB
flabel metal1 1257 -2095 1291 -2061 0 FreeSans 200 0 0 0 x2.VPWR
flabel metal1 1257 -2639 1291 -2605 0 FreeSans 200 0 0 0 x2.VGND
rlabel comment 1228 -2622 1228 -2622 4 x2.inv_4
rlabel metal1 1228 -2670 1688 -2574 1 x2.VGND
rlabel metal1 1228 -2126 1688 -2030 1 x2.VPWR
<< end >>
