magic
tech sky130A
timestamp 1710000196
<< metal1 >>
rect 23550 345138 23700 345200
rect 23550 345112 23612 345138
rect 23638 345112 23700 345138
rect 23550 345005 23700 345112
rect 21935 344915 21975 345005
rect 22675 344995 23700 345005
rect 22675 344969 23612 344995
rect 23638 344969 23700 344995
rect 22675 344963 23700 344969
rect 22675 344937 23612 344963
rect 23638 344937 23700 344963
rect 22675 344931 23700 344937
rect 22675 344915 23612 344931
rect 23550 344905 23612 344915
rect 23638 344905 23700 344931
rect 23550 344788 23700 344905
rect 23550 344762 23612 344788
rect 23638 344762 23700 344788
rect 23550 344700 23700 344762
rect 20950 344338 21100 344400
rect 20950 344312 21012 344338
rect 21038 344312 21100 344338
rect 20950 344245 21100 344312
rect 20950 344219 21012 344245
rect 21038 344219 21935 344245
rect 20950 344213 21935 344219
rect 20950 344187 21012 344213
rect 21038 344187 21935 344213
rect 20950 344181 21935 344187
rect 20950 344155 21012 344181
rect 21038 344155 21935 344181
rect 20950 344088 21100 344155
rect 20950 344062 21012 344088
rect 21038 344062 21100 344088
rect 20950 344000 21100 344062
rect 20460 331400 24150 331700
<< via1 >>
rect 23612 345112 23638 345138
rect 23612 344969 23638 344995
rect 23612 344937 23638 344963
rect 23612 344905 23638 344931
rect 23612 344762 23638 344788
rect 21012 344312 21038 344338
rect 21012 344219 21038 344245
rect 21012 344187 21038 344213
rect 21012 344155 21038 344181
rect 21012 344062 21038 344088
<< metal2 >>
rect 23600 345139 23650 345155
rect 23600 345111 23611 345139
rect 23639 345111 23650 345139
rect 23600 345095 23650 345111
rect 23600 344995 23650 345005
rect 23600 344984 23612 344995
rect 23638 344984 23650 344995
rect 23600 344956 23611 344984
rect 23639 344956 23650 344984
rect 23600 344944 23612 344956
rect 23638 344944 23650 344956
rect 23600 344916 23611 344944
rect 23639 344916 23650 344944
rect 23600 344905 23612 344916
rect 23638 344905 23650 344916
rect 23600 344895 23650 344905
rect 23600 344789 23650 344805
rect 23600 344761 23611 344789
rect 23639 344761 23650 344789
rect 23600 344745 23650 344761
rect 21000 344339 21050 344355
rect 21000 344311 21011 344339
rect 21039 344311 21050 344339
rect 21000 344295 21050 344311
rect 21000 344245 21050 344255
rect 21000 344234 21012 344245
rect 21038 344234 21050 344245
rect 21000 344206 21011 344234
rect 21039 344206 21050 344234
rect 21000 344194 21012 344206
rect 21038 344194 21050 344206
rect 21000 344166 21011 344194
rect 21039 344166 21050 344194
rect 21000 344155 21012 344166
rect 21038 344155 21050 344166
rect 21000 344145 21050 344155
rect 21000 344089 21050 344105
rect 21000 344061 21011 344089
rect 21039 344061 21050 344089
rect 21000 344045 21050 344061
rect 21120 341554 21320 342305
rect 21120 341526 21136 341554
rect 21164 341526 21206 341554
rect 21234 341526 21276 341554
rect 21304 341526 21320 341554
rect 21120 341510 21320 341526
rect 23320 341554 23520 342305
rect 23320 341526 23336 341554
rect 23364 341526 23406 341554
rect 23434 341526 23476 341554
rect 23504 341526 23520 341554
rect 23320 341510 23520 341526
<< via2 >>
rect 23611 345138 23639 345139
rect 23611 345112 23612 345138
rect 23612 345112 23638 345138
rect 23638 345112 23639 345138
rect 23611 345111 23639 345112
rect 23611 344969 23612 344984
rect 23612 344969 23638 344984
rect 23638 344969 23639 344984
rect 23611 344963 23639 344969
rect 23611 344956 23612 344963
rect 23612 344956 23638 344963
rect 23638 344956 23639 344963
rect 23611 344937 23612 344944
rect 23612 344937 23638 344944
rect 23638 344937 23639 344944
rect 23611 344931 23639 344937
rect 23611 344916 23612 344931
rect 23612 344916 23638 344931
rect 23638 344916 23639 344931
rect 23611 344788 23639 344789
rect 23611 344762 23612 344788
rect 23612 344762 23638 344788
rect 23638 344762 23639 344788
rect 23611 344761 23639 344762
rect 21011 344338 21039 344339
rect 21011 344312 21012 344338
rect 21012 344312 21038 344338
rect 21038 344312 21039 344338
rect 21011 344311 21039 344312
rect 21011 344219 21012 344234
rect 21012 344219 21038 344234
rect 21038 344219 21039 344234
rect 21011 344213 21039 344219
rect 21011 344206 21012 344213
rect 21012 344206 21038 344213
rect 21038 344206 21039 344213
rect 21011 344187 21012 344194
rect 21012 344187 21038 344194
rect 21038 344187 21039 344194
rect 21011 344181 21039 344187
rect 21011 344166 21012 344181
rect 21012 344166 21038 344181
rect 21038 344166 21039 344181
rect 21011 344088 21039 344089
rect 21011 344062 21012 344088
rect 21012 344062 21038 344088
rect 21038 344062 21039 344088
rect 21011 344061 21039 344062
rect 21136 341526 21164 341554
rect 21206 341526 21234 341554
rect 21276 341526 21304 341554
rect 23336 341526 23364 341554
rect 23406 341526 23434 341554
rect 23476 341526 23504 341554
<< metal3 >>
rect 23160 345780 27603 346020
rect 23550 345139 27603 345200
rect 23550 345111 23611 345139
rect 23639 345111 27603 345139
rect 23550 344984 27603 345111
rect 23550 344956 23611 344984
rect 23639 344956 27603 344984
rect 23550 344944 27603 344956
rect 23550 344916 23611 344944
rect 23639 344916 27603 344944
rect 23550 344789 27603 344916
rect 23550 344761 23611 344789
rect 23639 344761 27603 344789
rect 23550 344700 27603 344761
rect 17085 344339 21100 344400
rect 17085 344311 21011 344339
rect 21039 344311 21100 344339
rect 17085 344234 21100 344311
rect 17085 344206 21011 344234
rect 21039 344206 21100 344234
rect 17085 344194 21100 344206
rect 17085 344166 21011 344194
rect 21039 344166 21100 344194
rect 17085 344089 21100 344166
rect 17085 344061 21011 344089
rect 21039 344061 21100 344089
rect 17085 344000 21100 344061
rect 19222 343500 23900 343700
rect 21120 341554 21955 341570
rect 21120 341526 21136 341554
rect 21164 341526 21206 341554
rect 21234 341526 21276 341554
rect 21304 341526 21955 341554
rect 21120 341510 21955 341526
rect 22680 341554 23520 341570
rect 22680 341526 23336 341554
rect 23364 341526 23406 341554
rect 23434 341526 23476 341554
rect 23504 341526 23520 341554
rect 22680 341510 23520 341526
rect 22720 340930 27603 341160
<< metal4 >>
rect 19335 337683 19665 343025
rect 24960 336984 25290 343050
rect 24960 336866 25066 336984
rect 25184 336866 25290 336984
rect 24960 336784 25290 336866
rect 24960 336666 25066 336784
rect 25184 336666 25290 336784
rect 24960 336584 25290 336666
rect 24960 336466 25066 336584
rect 25184 336466 25290 336584
rect 24960 336350 25290 336466
<< via4 >>
rect 25066 336866 25184 336984
rect 25066 336666 25184 336784
rect 25066 336466 25184 336584
<< metal5 >>
rect 20460 336984 25650 337100
rect 20460 336866 25066 336984
rect 25184 336866 25650 336984
rect 20460 336784 25650 336866
rect 20460 336666 25066 336784
rect 25184 336666 25650 336784
rect 20460 336584 25650 336666
rect 20460 336466 25066 336584
rect 25184 336466 25650 336584
rect 20460 336350 25650 336466
rect 20460 334750 24150 335450
rect 20460 333100 24150 333800
use constant_gm_fingers  constant_gm_fingers_0
timestamp 1710000196
transform 1 0 21905 0 1 341450
box -1350 -10010 2210 570
use OTA_fingers_031123_NON_FLAT  OTA_fingers_031123_NON_FLAT_0
timestamp 1710000196
transform 1 0 21370 0 1 342355
box -2970 -155 4890 8275
<< properties >>
string FIXED_BBOX 0 0 292000 352000
<< end >>
