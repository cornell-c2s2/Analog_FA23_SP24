* NGSPICE file created from flashADC_flat.ext - technology: sky130A

.subckt flashADC_flat VFS OUT3 OUT2 OUT1 OUT0 VL VDD CLK VIN GND VV15 VV14 VV13 VV12 VV11 VV10 VV9 VV8 VV7 VV6 VV5 VV4 VV3 VV2 VV1 VV16 I14 I13 I12
+ I11 I10 I9 I8 I7 I6 I5 I4 I3 I2 I1 I0 I15 S1 R1 S0 R0
X0 GND.t1375 frontAnalog_v0p0p1_7.x65.X frontAnalog_v0p0p1_7.RSfetsym_0.x2.Y GND.t1374 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1 OUT3.t127 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD.t1251 VDD.t1250 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 VDD.t1059 frontAnalog_v0p0p1_15.x63.A.t4 a_57123_n85079# VDD.t1058 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X3 GND.t208 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t63 GND.t207 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X4 VDD.t490 frontAnalog_v0p0p1_10.x63.X I5.t1 VDD.t485 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.25
X5 VDD.t965 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t127 VDD.t964 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 VFS.t3 VV16.t6 GND.t21 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X7 a_78315_n41309# 16to4_PriorityEncoder_v0p0p1_0.x5.x11.X a_78243_n41309# VDD.t290 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X8 a_16719_n13117.t23 a_16599_n13205.t4 a_16541_n13117.t7 GND.t1567 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X9 w_55000_n56928# CLK.t0 frontAnalog_v0p0p1_10.x65.A.t3 VDD.t1084 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X10 VV4.t4 VV3.t5 GND.t244 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X11 frontAnalog_v0p0p1_3.x65.X a_57123_n13359# VDD.t1384 VDD.t1383 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X12 VDD.t1340 frontAnalog_v0p0p1_9.x63.X frontAnalog_v0p0p1_9.RSfetsym_0.x1.Y VDD.t1333 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X13 OUT3.t63 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND.t1312 GND.t1311 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X14 frontAnalog_v0p0p1_14.x65.A.t2 frontAnalog_v0p0p1_14.x63.A.t4 a_55268_n79536# GND.t861 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X15 OUT2.t63 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND.t1012 GND.t1011 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X16 frontAnalog_v0p0p1_5.RSfetsym_0.QN.t0 frontAnalog_v0p0p1_5.RSfetsym_0.x1.Y GND.t11 GND.t10 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.25
X17 16to4_PriorityEncoder_v0p0p1_0.x29.A 16to4_PriorityEncoder_v0p0p1_0.x28.A VDD.t993 VDD.t992 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X18 VV11.t13 VV10.t14 GND.t299 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X19 frontAnalog_v0p0p1_6.x63.X a_57123_n31079# GND.t582 GND.t581 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X20 GND.t1310 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t62 GND.t1309 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X21 GND.t1059 frontAnalog_v0p0p1_8.x63.X frontAnalog_v0p0p1_8.RSfetsym_0.x1.Y GND.t1054 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X22 GND.t1010 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t62 GND.t1009 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X23 OUT3.t126 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD.t1249 VDD.t1248 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X24 VV2.t5 VV1.t2 GND.t12 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X25 a_53630_n84996# VV1.t16 w_55000_n83928# GND.t284 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X26 16to4_PriorityEncoder_v0p0p1_0.x29.Y 16to4_PriorityEncoder_v0p0p1_0.x29.A GND.t241 GND.t240 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X27 GND.t1151 I0.t5 a_77605_n47345# GND.t531 sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X28 VDD.t214 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t127 VDD.t213 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X29 VDD.t1247 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t125 VDD.t1246 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X30 a_55268_n63336# CLK.t1 GND.t1144 GND.t1143 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X31 GND.t486 16to4_PriorityEncoder_v0p0p1_0.x5.x17.A a_78349_n43045# GND.t319 sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X32 frontAnalog_v0p0p1_14.RSfetsym_0.x1.Y R1.t2 VDD.t561 VDD.t560 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X33 a_77605_n51335# I2.t5 VDD.t1065 VDD.t1064 sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.109 ps=1.36 w=0.42 l=0.15
X34 frontAnalog_v0p0p1_5.RSfetsym_0.x1.Y frontAnalog_v0p0p1_5.x63.X GND.t1033 GND.t1029 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X35 VDD.t489 frontAnalog_v0p0p1_10.x63.X frontAnalog_v0p0p1_10.RSfetsym_0.x1.Y VDD.t483 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X36 VDD.t814 VDD.t812 a_77605_n43295# VDD.t813 sky130_fd_pr__pfet_01v8_hvt ad=0.312 pd=1.68 as=0.0588 ps=0.7 w=0.42 l=0.15
X37 VDD.t779 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t127 VDD.t778 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X38 GND.t1308 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t61 GND.t1307 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X39 GND.t1022 frontAnalog_v0p0p1_8.RSfetsym_0.QN.t5 a_59577_n46683# GND.t1021 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X40 GND.t1008 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t61 GND.t1007 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X41 GND.t360 I5.t5 a_59578_n56970# GND.t359 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X42 a_53630_n41796# VV9.t16 w_55000_n40728# GND.t1094 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X43 VDD.t963 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t126 VDD.t962 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X44 VV16.t4 VV15.t3 GND.t80 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X45 OUT1.t63 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND.t846 GND.t845 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X46 GND.t400 frontAnalog_v0p0p1_12.x65.X frontAnalog_v0p0p1_12.RSfetsym_0.x2.Y GND.t399 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X47 OUT2.t125 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD.t961 VDD.t960 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X48 GND.t239 16to4_PriorityEncoder_v0p0p1_0.x29.A 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND.t238 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X49 frontAnalog_v0p0p1_7.RSfetsym_0.x1.Y frontAnalog_v0p0p1_7.x63.X VDD.t587 VDD.t580 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X50 OUT0.t62 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND.t206 GND.t205 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X51 a_77637_n50057# 16to4_PriorityEncoder_v0p0p1_0.x3.EI VDD.t363 VDD.t362 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X52 frontAnalog_v0p0p1_2.x65.A.t3 frontAnalog_v0p0p1_2.x63.A.t4 a_55268_n3936# GND.t503 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X53 VDD.t1 S0.t2 frontAnalog_v0p0p1_15.RSfetsym_0.QN.t4 VDD.t0 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.25
X54 GND.t1306 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t60 GND.t1305 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X55 GND.t204 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t61 GND.t203 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X56 a_82906_n51645# 16to4_PriorityEncoder_v0p0p1_0.x3.A0 GND.t1101 GND.t1100 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X57 OUT3.t124 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD.t1245 VDD.t1244 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X58 frontAnalog_v0p0p1_6.RSfetsym_0.QN.t3 I10.t5 VDD.t641 VDD.t395 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.3
X59 a_77881_n44527# 16to4_PriorityEncoder_v0p0p1_0.x5.x18.C a_77775_n44527# GND.t511 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X60 GND.t1425 I13.t5 a_59578_n13770# GND.t1424 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X61 OUT3.t59 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND.t1304 GND.t1303 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X62 16to4_PriorityEncoder_v0p0p1_0.x36.Y 16to4_PriorityEncoder_v0p0p1_0.x36.A GND.t63 GND.t62 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X63 a_53630_n9396# frontAnalog_v0p0p1_10.IB.t3 GND.t1017 GND.t293 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X64 VDD.t1243 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t123 VDD.t1242 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X65 VDD.t465 frontAnalog_v0p0p1_2.x63.A.t5 a_57123_n4079# VDD.t464 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X66 frontAnalog_v0p0p1_11.x63.X a_57123_n63479# VDD.t1463 VDD.t1462 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X67 a_77723_n41087# VDD.t1502 a_77637_n41087# GND.t691 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X68 VV14.t11 VV13.t12 GND.t299 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X69 GND.t416 frontAnalog_v0p0p1_6.x65.X frontAnalog_v0p0p1_6.RSfetsym_0.x2.Y GND.t415 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X70 GND.t374 16to4_PriorityEncoder_v0p0p1_0.x21.A 16to4_PriorityEncoder_v0p0p1_0.x22.A GND.t373 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X71 w_55000_n79150# VIN.t0 a_53630_n79596# GND.t22 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X72 GND.t1389 R0.t2 frontAnalog_v0p0p1_15.RSfetsym_0.x1.Y GND.t1065 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X73 VIN.t1 w_55000_n51528# error sky130_fd_pr__cap_var_lvt w=2 l=0.18
X74 GND.t844 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t62 GND.t843 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X75 16to4_PriorityEncoder_v0p0p1_0.x5.x19.X a_77605_n44779# VDD.t432 VDD.t431 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.312 ps=1.68 w=1 l=0.15
X76 OUT2.t124 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD.t959 VDD.t958 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X77 VV4.t3 VV3.t3 GND.t401 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X78 16to4_PriorityEncoder_v0p0p1_0.x43.Y 16to4_PriorityEncoder_v0p0p1_0.x43.A VDD.t325 VDD.t324 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X79 VDD.t248 frontAnalog_v0p0p1_4.x65.A.t4 a_57123_n18759# VDD.t247 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X80 VV10.t5 VV9.t5 GND.t12 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X81 OUT0.t126 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD.t212 VDD.t211 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X82 a_78065_n41309# 16to4_PriorityEncoder_v0p0p1_0.x5.x22.A GND.t324 GND.t323 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X83 OUT0.t60 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND.t202 GND.t201 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X84 GND.t200 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t59 GND.t199 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X85 VV3.t7 VV2.t7 GND.t209 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X86 VDD.t361 16to4_PriorityEncoder_v0p0p1_0.x3.EI a_77605_n51335# VDD.t360 sky130_fd_pr__pfet_01v8_hvt ad=0.312 pd=1.68 as=0.0588 ps=0.7 w=0.42 l=0.15
X87 VV13.t0 VV12.t0 GND.t12 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X88 VDD.t210 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t125 VDD.t209 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X89 OUT3.t58 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND.t1302 GND.t1301 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X90 frontAnalog_v0p0p1_9.x65.A.t2 CLK.t2 frontAnalog_v0p0p1_9.x63.A.t2 VDD.t1085 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X91 OUT2.t60 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND.t1006 GND.t1005 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X92 frontAnalog_v0p0p1_12.RSfetsym_0.x2.Y frontAnalog_v0p0p1_12.x65.X VDD.t377 VDD.t372 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X93 VDD.t1241 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t122 VDD.t1240 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X94 frontAnalog_v0p0p1_4.x63.X a_57123_n20279# VDD.t86 VDD.t85 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X95 GND.t842 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t61 GND.t841 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X96 w_55000_n35950# VIN.t2 a_53630_n36396# GND.t281 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X97 GND.t1532 frontAnalog_v0p0p1_1.x63.X frontAnalog_v0p0p1_1.RSfetsym_0.x1.Y GND.t1527 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X98 frontAnalog_v0p0p1_10.RSfetsym_0.x2.Y frontAnalog_v0p0p1_10.x65.X GND.t1181 GND.t1180 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X99 GND.t1300 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t57 GND.t1299 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X100 VDD.t327 I5.t6 a_77637_n49127# VDD.t326 sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X101 GND.t61 16to4_PriorityEncoder_v0p0p1_0.x36.A 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND.t60 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X102 VDD.t344 16to4_PriorityEncoder_v0p0p1_0.x21.A 16to4_PriorityEncoder_v0p0p1_0.x22.A VDD.t343 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X103 frontAnalog_v0p0p1_2.RSfetsym_0.x1.Y frontAnalog_v0p0p1_2.x63.X GND.t480 GND.t475 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X104 VDD.t66 16to4_PriorityEncoder_v0p0p1_0.x36.A 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD.t65 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X105 a_16541_n13117.t1 GND.t1487 GND.t657 sky130_fd_pr__res_xhigh_po_5p73 l=85.8
X106 I1.t3 frontAnalog_v0p0p1_14.RSfetsym_0.x2.Y GND.t602 GND.t594 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.25
X107 GND.t325 frontAnalog_v0p0p1_9.x65.A.t4 a_57123_n51159# GND.t255 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X108 VV3.t1 VV2.t1 GND.t79 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X109 VDD.t1358 I13.t6 a_77605_n45765# VDD.t804 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X110 a_77881_n52567# 16to4_PriorityEncoder_v0p0p1_0.x3.x18.C a_77775_n52567# GND.t67 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X111 16to4_PriorityEncoder_v0p0p1_0.x22.Y 16to4_PriorityEncoder_v0p0p1_0.x22.A GND.t1475 GND.t1474 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X112 frontAnalog_v0p0p1_9.x63.A.t0 frontAnalog_v0p0p1_9.x65.A.t5 a_55268_n52536# GND.t326 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X113 OUT2.t123 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD.t957 VDD.t956 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X114 OUT0.t124 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD.t208 VDD.t207 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X115 VDD.t206 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t123 VDD.t205 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X116 I6.t1 frontAnalog_v0p0p1_9.RSfetsym_0.QN.t5 VDD.t250 VDD.t249 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.3
X117 frontAnalog_v0p0p1_6.RSfetsym_0.x2.Y frontAnalog_v0p0p1_6.x65.X VDD.t390 VDD.t385 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X118 GND.t358 16to4_PriorityEncoder_v0p0p1_0.x43.A 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND.t357 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X119 GND.t840 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t60 GND.t839 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X120 OUT2.t122 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD.t955 VDD.t954 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X121 frontAnalog_v0p0p1_3.RSfetsym_0.x2.Y frontAnalog_v0p0p1_3.x65.X GND.t879 GND.t878 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X122 a_77639_n42341# VDD.t809 VDD.t811 VDD.t810 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X123 frontAnalog_v0p0p1_13.RSfetsym_0.x1.Y frontAnalog_v0p0p1_13.x63.X GND.t1114 GND.t1110 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X124 a_59577_n57483# frontAnalog_v0p0p1_10.x63.X I5.t2 GND.t530 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X125 a_59578_n67770# frontAnalog_v0p0p1_13.x65.X frontAnalog_v0p0p1_13.RSfetsym_0.QN.t2 GND.t1503 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.315 ps=2.72 w=1 l=0.15
X126 a_77687_n45765# I13.t7 a_77605_n45765# GND.t1426 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X127 16to4_PriorityEncoder_v0p0p1_0.x42.A 16to4_PriorityEncoder_v0p0p1_0.x5.GS VDD.t1483 VDD.t1482 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X128 16to4_PriorityEncoder_v0p0p1_0.x3.x19.X a_77605_n52819# VDD.t638 VDD.t637 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.312 ps=1.68 w=1 l=0.15
X129 VV2.t10 VV1.t7 GND.t417 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X130 VDD.t953 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t121 VDD.t952 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X131 OUT1.t59 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND.t838 GND.t837 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X132 frontAnalog_v0p0p1_7.x63.A.t1 frontAnalog_v0p0p1_7.x65.A.t4 VDD.t1378 VDD.t419 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X133 I9.t3 frontAnalog_v0p0p1_7.RSfetsym_0.x2.Y GND.t707 GND.t473 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.25
X134 VV7.t16 w_55000_n52150# error sky130_fd_pr__cap_var_lvt w=2 l=0.18
X135 a_16719_n13117.t22 a_16599_n13205.t5 a_16541_n13117.t6 GND.t1568 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X136 16to4_PriorityEncoder_v0p0p1_0.x5.x11.X a_77637_n41087# GND.t717 GND.t579 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.112 ps=1.04 w=0.65 l=0.15
X137 OUT0.t58 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND.t198 GND.t197 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X138 GND.t1014 16to4_PriorityEncoder_v0p0p1_0.x3.x14.A a_78065_n49349# GND.t1013 sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X139 a_78703_n45515# 16to4_PriorityEncoder_v0p0p1_0.x5.x19.X a_78607_n45515# VDD.t457 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X140 frontAnalog_v0p0p1_2.x65.X a_57123_n2559# GND.t1148 GND.t1147 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X141 16to4_PriorityEncoder_v0p0p1_0.x22.Y 16to4_PriorityEncoder_v0p0p1_0.x22.A VDD.t1416 VDD.t1415 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X142 a_16719_n13117.t3 a_16719_n13117.t2 a_16599_n13205.t0 GND.t1072 sky130_fd_pr__nfet_01v8_lvt ad=0.122 pd=1.42 as=0.122 ps=1.42 w=0.42 l=0.15
X143 VV6.t2 VV5.t4 GND.t21 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X144 VDD.t1263 frontAnalog_v0p0p1_8.x65.X frontAnalog_v0p0p1_8.RSfetsym_0.x2.Y VDD.t1256 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X145 GND.t1298 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t56 GND.t1297 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X146 GND.t1473 16to4_PriorityEncoder_v0p0p1_0.x22.A 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND.t1472 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X147 VDD.t951 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t120 VDD.t950 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X148 VDD.t1068 frontAnalog_v0p0p1_13.x63.A.t4 a_57123_n68879# VDD.t1067 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X149 a_59577_n14283# frontAnalog_v0p0p1_3.x63.X I13.t4 GND.t1513 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X150 a_59578_n24570# frontAnalog_v0p0p1_5.x65.X frontAnalog_v0p0p1_5.RSfetsym_0.QN.t2 GND.t470 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.315 ps=2.72 w=1 l=0.15
X151 16to4_PriorityEncoder_v0p0p1_0.x29.Y 16to4_PriorityEncoder_v0p0p1_0.x29.A GND.t237 GND.t236 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X152 VV7.t5 VV6.t6 GND.t250 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X153 I6.t3 frontAnalog_v0p0p1_9.x63.X VDD.t1339 VDD.t1336 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.25
X154 a_53630_n63396# frontAnalog_v0p0p1_10.IB.t4 GND.t1018 GND.t296 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X155 16to4_PriorityEncoder_v0p0p1_0.x5.x22.A a_77639_n42341# VDD.t566 VDD.t565 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.167 ps=1.39 w=1 l=0.15
X156 frontAnalog_v0p0p1_0.RSfetsym_0.x1.Y frontAnalog_v0p0p1_0.x63.X GND.t75 GND.t71 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X157 16to4_PriorityEncoder_v0p0p1_0.x43.Y 16to4_PriorityEncoder_v0p0p1_0.x43.A GND.t356 GND.t355 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X158 VDD.t267 frontAnalog_v0p0p1_10.x63.A.t4 frontAnalog_v0p0p1_10.x65.A.t0 VDD.t266 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X159 OUT2.t59 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND.t1004 GND.t1003 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X160 frontAnalog_v0p0p1_0.RSfetsym_0.x2.Y frontAnalog_v0p0p1_0.x65.X GND.t1342 GND.t1341 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X161 OUT1.t126 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD.t777 VDD.t776 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X162 w_55000_n8950# VIN.t3 a_53630_n9396# GND.t282 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X163 VDD.t329 I5.t7 a_77605_n53805# VDD.t328 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X164 frontAnalog_v0p0p1_12.x65.X a_57123_n72759# GND.t1534 GND.t1533 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X165 VDD.t775 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t125 VDD.t774 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X166 OUT0.t122 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD.t204 VDD.t203 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X167 frontAnalog_v0p0p1_4.RSfetsym_0.x2.Y frontAnalog_v0p0p1_4.x65.X GND.t1486 GND.t1485 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X168 GND.t1296 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t55 GND.t1295 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X169 VDD.t367 frontAnalog_v0p0p1_5.x63.A.t4 a_57123_n25679# VDD.t366 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X170 GND.t196 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t57 GND.t195 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X171 a_53630_n20196# frontAnalog_v0p0p1_10.IB.t5 GND.t1019 GND.t296 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X172 a_77639_n50381# 16to4_PriorityEncoder_v0p0p1_0.x3.EI VDD.t359 VDD.t358 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X173 VDD.t64 16to4_PriorityEncoder_v0p0p1_0.x36.A 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD.t63 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X174 VDD.t1414 16to4_PriorityEncoder_v0p0p1_0.x22.A 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD.t1413 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X175 VDD.t1016 frontAnalog_v0p0p1_3.x63.A.t4 frontAnalog_v0p0p1_3.x65.A.t0 VDD.t521 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X176 OUT3.t54 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND.t1294 GND.t1293 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X177 VDD.t406 frontAnalog_v0p0p1_15.x65.A.t4 a_57123_n83559# VDD.t405 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X178 GND.t863 frontAnalog_v0p0p1_14.x63.A.t5 a_57123_n79679# GND.t862 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X179 a_55268_n47136# CLK.t3 GND.t1146 GND.t1145 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X180 frontAnalog_v0p0p1_1.RSfetsym_0.x2.Y frontAnalog_v0p0p1_1.x65.X GND.t520 GND.t519 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X181 VDD.t376 frontAnalog_v0p0p1_12.x65.X frontAnalog_v0p0p1_12.RSfetsym_0.x2.Y VDD.t372 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X182 GND.t668 16to4_PriorityEncoder_v0p0p1_0.x3.x15.X a_78349_n51085# GND.t505 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X183 frontAnalog_v0p0p1_4.x65.A.t2 frontAnalog_v0p0p1_4.x63.A.t4 a_55268_n20136# GND.t1390 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X184 frontAnalog_v0p0p1_9.RSfetsym_0.QN.t4 I6.t5 VDD.t1477 VDD.t249 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.3
X185 OUT3.t121 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD.t1239 VDD.t1238 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X186 VV10.t8 VV9.t10 GND.t417 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X187 a_78703_n53555# 16to4_PriorityEncoder_v0p0p1_0.x3.x19.X a_78607_n53555# VDD.t1066 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X188 GND.t194 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t56 GND.t193 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X189 OUT1.t58 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND.t836 GND.t835 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X190 VV12.t5 VV11.t5 GND.t257 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X191 VV3.t6 VV2.t6 GND.t589 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X192 a_77775_n51335# 16to4_PriorityEncoder_v0p0p1_0.x3.x19.C a_77687_n51335# GND.t69 sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
X193 16to4_PriorityEncoder_v0p0p1_0.x43.A 16to4_PriorityEncoder_v0p0p1_0.x42.A VDD.t1279 VDD.t1278 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X194 a_53630_n25596# VV12.t16 w_55000_n24528# GND.t317 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X195 VV13.t7 VV12.t7 GND.t417 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X196 OUT3.t53 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND.t1292 GND.t1291 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X197 16to4_PriorityEncoder_v0p0p1_0.x28.A 16to4_PriorityEncoder_v0p0p1_0.x1.X GND.t403 GND.t402 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X198 VDD.t202 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t121 VDD.t201 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X199 VDD.t949 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t119 VDD.t948 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X200 frontAnalog_v0p0p1_9.RSfetsym_0.x2.Y frontAnalog_v0p0p1_9.x65.X VDD.t1373 VDD.t1368 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X201 VDD.t1354 frontAnalog_v0p0p1_1.x65.A.t4 a_57123_n40359# VDD.t1353 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X202 GND.t1157 frontAnalog_v0p0p1_7.x63.A.t4 a_57123_n36479# GND.t1156 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X203 frontAnalog_v0p0p1_10.RSfetsym_0.QN.t4 frontAnalog_v0p0p1_10.x65.X VDD.t1118 VDD.t1114 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.25
X204 frontAnalog_v0p0p1_9.RSfetsym_0.x1.Y frontAnalog_v0p0p1_9.x63.X GND.t1403 GND.t1398 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X205 VDD.t389 frontAnalog_v0p0p1_6.x65.X frontAnalog_v0p0p1_6.RSfetsym_0.x2.Y VDD.t385 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X206 16to4_PriorityEncoder_v0p0p1_0.x36.Y 16to4_PriorityEncoder_v0p0p1_0.x36.A VDD.t62 VDD.t61 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X207 VDD.t1347 I4.t5 a_77637_n48817# VDD.t1346 sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X208 VDD.t773 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t124 VDD.t772 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X209 VDD.t1440 frontAnalog_v0p0p1_13.x65.X frontAnalog_v0p0p1_13.RSfetsym_0.QN.t4 VDD.t1436 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.25
X210 GND.t192 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t55 GND.t191 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X211 VDD.t200 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t120 VDD.t199 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X212 frontAnalog_v0p0p1_11.RSfetsym_0.x1.Y frontAnalog_v0p0p1_11.x63.X VDD.t12 VDD.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X213 OUT0.t54 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND.t190 GND.t189 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X214 VFS.t1 VV16.t1 GND.t289 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X215 frontAnalog_v0p0p1_3.RSfetsym_0.QN.t4 frontAnalog_v0p0p1_3.x65.X VDD.t835 VDD.t831 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.25
X216 VDD.t1277 16to4_PriorityEncoder_v0p0p1_0.x42.A 16to4_PriorityEncoder_v0p0p1_0.x43.A VDD.t1276 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X217 VDD.t771 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t123 VDD.t770 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X218 VV4.t6 VV3.t9 GND.t80 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X219 VV15.t16 w_55000_n8950# error sky130_fd_pr__cap_var_lvt w=2 l=0.18
X220 16to4_PriorityEncoder_v0p0p1_0.x5.x17.A a_77637_n42017# GND.t1184 GND.t1183 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.112 ps=1.04 w=0.65 l=0.15
X221 VDD.t440 frontAnalog_v0p0p1_5.x65.X frontAnalog_v0p0p1_5.RSfetsym_0.QN.t4 VDD.t436 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.25
X222 VV15.t11 VV14.t12 GND.t244 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X223 GND.t74 frontAnalog_v0p0p1_0.x63.X frontAnalog_v0p0p1_0.RSfetsym_0.x1.Y GND.t71 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X224 VDD.t1237 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t120 VDD.t1236 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X225 16to4_PriorityEncoder_v0p0p1_0.x22.Y 16to4_PriorityEncoder_v0p0p1_0.x22.A GND.t1471 GND.t1470 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X226 VDD.t198 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t119 VDD.t197 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X227 a_16719_n13117.t21 a_16599_n13205.t6 a_16541_n13117.t5 GND.t1569 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X228 frontAnalog_v0p0p1_7.x65.A.t2 CLK.t4 frontAnalog_v0p0p1_7.x63.A.t2 VDD.t1086 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X229 VV7.t14 VV6.t14 GND.t78 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X230 VDD.t562 R1.t3 frontAnalog_v0p0p1_14.RSfetsym_0.x1.Y VDD.t560 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X231 frontAnalog_v0p0p1_6.x63.A.t2 CLK.t5 w_55000_n30550# VDD.t1087 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X232 GND.t1032 frontAnalog_v0p0p1_5.x63.X frontAnalog_v0p0p1_5.RSfetsym_0.x1.Y GND.t1029 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X233 OUT2.t118 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD.t947 VDD.t946 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X234 OUT0.t118 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD.t196 VDD.t195 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X235 a_78607_n45515# 16to4_PriorityEncoder_v0p0p1_0.x5.x20.X a_78525_n45515# VDD.t1443 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X236 VDD.t600 frontAnalog_v0p0p1_2.x65.A.t4 a_57123_n2559# VDD.t599 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X237 frontAnalog_v0p0p1_11.x65.X a_57123_n61959# VDD.t985 VDD.t984 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X238 GND.t1484 frontAnalog_v0p0p1_4.x65.X frontAnalog_v0p0p1_4.RSfetsym_0.x2.Y GND.t1483 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X239 frontAnalog_v0p0p1_10.x63.X a_57123_n58079# GND.t1105 GND.t1104 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X240 OUT1.t122 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD.t769 VDD.t768 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X241 frontAnalog_v0p0p1_9.x63.A.t3 CLK.t6 w_55000_n52150# VDD.t251 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X242 VDD.t1019 CLK.t7 w_55000_n73128# GND.t536 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X243 GND.t1442 frontAnalog_v0p0p1_7.x65.A.t5 a_57123_n34959# GND.t1156 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X244 frontAnalog_v0p0p1_12.RSfetsym_0.QN.t3 frontAnalog_v0p0p1_12.RSfetsym_0.x1.Y GND.t424 GND.t423 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.25
X245 GND.t1002 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t58 GND.t1001 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X246 16to4_PriorityEncoder_v0p0p1_0.x5.x16.X a_77605_n43545# GND.t14 GND.t13 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.196 ps=1.33 w=0.65 l=0.15
X247 GND.t824 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t57 GND.t823 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X248 GND.t518 frontAnalog_v0p0p1_1.x65.X frontAnalog_v0p0p1_1.RSfetsym_0.x2.Y GND.t517 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X249 frontAnalog_v0p0p1_15.RSfetsym_0.x2.Y S0.t3 GND.t1 GND.t0 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X250 frontAnalog_v0p0p1_3.RSfetsym_0.x2.Y frontAnalog_v0p0p1_3.x65.X VDD.t834 VDD.t828 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X251 VDD.t586 frontAnalog_v0p0p1_7.x63.X frontAnalog_v0p0p1_7.RSfetsym_0.x1.Y VDD.t580 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X252 VDD.t11 frontAnalog_v0p0p1_11.x63.X I4.t2 VDD.t5 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.25
X253 VDD.t1020 CLK.t8 w_55000_n73750# GND.t573 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X254 16to4_PriorityEncoder_v0p0p1_0.x22.Y 16to4_PriorityEncoder_v0p0p1_0.x22.A VDD.t1412 VDD.t1411 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X255 VV1.t8 VL.t5 GND.t12 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X256 w_55000_n62328# CLK.t9 frontAnalog_v0p0p1_11.x65.A.t3 VDD.t1021 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X257 a_78243_n41309# 16to4_PriorityEncoder_v0p0p1_0.x5.x17.A a_78147_n41309# VDD.t290 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X258 OUT2.t117 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD.t933 VDD.t932 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X259 VDD.t808 VDD.t806 a_78649_n39527# VDD.t807 sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X260 frontAnalog_v0p0p1_3.x63.X a_57123_n14879# GND.t1358 GND.t1357 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X261 OUT3.t52 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND.t1290 GND.t1289 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X262 VV10.t16 w_55000_n35950# error sky130_fd_pr__cap_var_lvt w=2 l=0.18
X263 frontAnalog_v0p0p1_15.x65.A.t3 frontAnalog_v0p0p1_15.x63.A.t5 a_55268_n84936# GND.t1361 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X264 a_53630_n68796# VV4.t16 w_55000_n67728# GND.t242 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X265 VDD.t945 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t116 VDD.t944 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X266 VV9.t15 VV8.t15 GND.t12 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X267 VDD.t1235 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t119 VDD.t1234 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X268 16to4_PriorityEncoder_v0p0p1_0.x3.x17.A a_77637_n50057# GND.t388 GND.t387 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.112 ps=1.04 w=0.65 l=0.15
X269 OUT0.t53 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND.t188 GND.t187 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X270 GND.t1288 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t51 GND.t1287 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X271 GND.t1402 frontAnalog_v0p0p1_9.x63.X frontAnalog_v0p0p1_9.RSfetsym_0.x1.Y GND.t1398 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X272 OUT3.t118 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD.t1233 VDD.t1232 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X273 16to4_PriorityEncoder_v0p0p1_0.x21.A 16to4_PriorityEncoder_v0p0p1_0.x2.X GND.t848 GND.t847 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X274 VIN.t4 w_55000_n8328# error sky130_fd_pr__cap_var_lvt w=2 l=0.18
X275 GND.t1441 16to4_PriorityEncoder_v0p0p1_0.x5.x21.B a_78183_n45737# GND.t1440 sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X276 VDD.t1022 CLK.t10 w_55000_n30550# GND.t568 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X277 VDD.t574 frontAnalog_v0p0p1_4.x63.X I12.t3 VDD.t567 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.25
X278 w_55000_n19128# CLK.t11 frontAnalog_v0p0p1_4.x65.A.t1 VDD.t1023 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X279 VDD.t323 16to4_PriorityEncoder_v0p0p1_0.x43.A 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD.t322 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X280 GND.t1352 16to4_PriorityEncoder_v0p0p1_0.x42.A 16to4_PriorityEncoder_v0p0p1_0.x43.A GND.t1351 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X281 GND.t1000 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t57 GND.t999 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X282 a_78607_n53555# 16to4_PriorityEncoder_v0p0p1_0.x3.x20.X a_78525_n53555# VDD.t559 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X283 frontAnalog_v0p0p1_1.x65.A.t0 frontAnalog_v0p0p1_1.x63.A.t4 a_55268_n41736# GND.t855 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X284 OUT2.t56 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND.t998 GND.t997 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X285 VDD.t10 frontAnalog_v0p0p1_11.x63.X frontAnalog_v0p0p1_11.RSfetsym_0.x1.Y VDD.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X286 GND.t834 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t56 GND.t833 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X287 VV15.t4 VV14.t3 GND.t401 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X288 16to4_PriorityEncoder_v0p0p1_0.x3.x16.C I5.t8 GND.t362 GND.t361 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X289 OUT0.t117 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD.t194 VDD.t193 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X290 OUT3.t117 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD.t1231 VDD.t1230 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X291 GND.t1179 frontAnalog_v0p0p1_10.x65.X frontAnalog_v0p0p1_10.RSfetsym_0.x2.Y GND.t1178 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X292 VIN.t5 w_55000_n78528# error sky130_fd_pr__cap_var_lvt w=2 l=0.18
X293 OUT1.t55 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND.t832 GND.t831 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X294 frontAnalog_v0p0p1_4.RSfetsym_0.x1.Y frontAnalog_v0p0p1_4.x63.X VDD.t573 VDD.t569 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X295 VDD.t1357 16to4_PriorityEncoder_v0p0p1_0.x1.A a_82988_n47995# VDD.t1356 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X296 GND.t479 frontAnalog_v0p0p1_2.x63.X frontAnalog_v0p0p1_2.RSfetsym_0.x1.Y GND.t475 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X297 16to4_PriorityEncoder_v0p0p1_0.x21.A 16to4_PriorityEncoder_v0p0p1_0.x2.X VDD.t781 VDD.t780 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X298 a_77687_n44779# VDD.t1503 a_77605_n44779# GND.t247 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.109 ps=1.36 w=0.42 l=0.15
X299 a_77723_n42017# VDD.t1504 a_77637_n42017# GND.t692 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X300 VDD.t357 16to4_PriorityEncoder_v0p0p1_0.x3.EI a_78649_n47567# VDD.t356 sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X301 GND.t996 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t55 GND.t995 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X302 OUT2.t54 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND.t994 GND.t993 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X303 frontAnalog_v0p0p1_14.x65.A.t0 CLK.t12 frontAnalog_v0p0p1_14.x63.A.t0 VDD.t1024 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X304 OUT2.t115 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD.t943 VDD.t942 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X305 16to4_PriorityEncoder_v0p0p1_0.x43.Y 16to4_PriorityEncoder_v0p0p1_0.x43.A VDD.t321 VDD.t320 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X306 frontAnalog_v0p0p1_8.x63.X a_57123_n47279# VDD.t454 VDD.t453 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X307 GND.t877 frontAnalog_v0p0p1_3.x65.X frontAnalog_v0p0p1_3.RSfetsym_0.x2.Y GND.t876 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X308 VIN.t6 w_55000_n35328# error sky130_fd_pr__cap_var_lvt w=2 l=0.18
X309 GND.t1113 frontAnalog_v0p0p1_13.x63.X frontAnalog_v0p0p1_13.RSfetsym_0.x1.Y GND.t1110 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X310 16to4_PriorityEncoder_v0p0p1_0.x43.Y 16to4_PriorityEncoder_v0p0p1_0.x43.A GND.t354 GND.t353 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X311 OUT1.t54 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND.t830 GND.t829 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X312 VDD.t941 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t114 VDD.t940 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X313 VDD.t1229 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t116 VDD.t1228 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X314 GND.t601 16to4_PriorityEncoder_v0p0p1_0.x3.x21.B a_78183_n53777# GND.t600 sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X315 a_53630_n74196# frontAnalog_v0p0p1_10.IB.t6 GND.t1020 GND.t296 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X316 w_55000_n84550# VIN.t7 a_53630_n84996# GND.t284 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X317 GND.t1160 frontAnalog_v0p0p1_14.x65.A.t4 a_57123_n78159# GND.t862 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X318 OUT2.t53 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND.t992 GND.t991 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X319 VDD.t619 frontAnalog_v0p0p1_5.x65.A.t4 a_57123_n24159# VDD.t618 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X320 GND.t1392 frontAnalog_v0p0p1_4.x63.A.t5 a_57123_n20279# GND.t1391 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X321 frontAnalog_v0p0p1_14.x63.A.t2 frontAnalog_v0p0p1_14.x65.A.t5 a_55268_n79536# GND.t1161 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X322 GND.t3 S0.t4 frontAnalog_v0p0p1_15.RSfetsym_0.x2.Y GND.t2 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X323 VDD.t767 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t121 VDD.t766 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X324 VDD.t833 frontAnalog_v0p0p1_3.x65.X frontAnalog_v0p0p1_3.RSfetsym_0.x2.Y VDD.t828 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X325 GND.t1286 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t50 GND.t1285 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X326 I1.t4 frontAnalog_v0p0p1_14.RSfetsym_0.QN.t5 VDD.t827 VDD.t279 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.3
X327 frontAnalog_v0p0p1_10.RSfetsym_0.x2.Y frontAnalog_v0p0p1_10.x65.X VDD.t1117 VDD.t1111 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X328 GND.t186 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t52 GND.t185 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X329 GND.t59 16to4_PriorityEncoder_v0p0p1_0.x36.A 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND.t58 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X330 w_55000_n19750# VIN.t8 a_53630_n20196# GND.t446 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X331 VDD.t60 16to4_PriorityEncoder_v0p0p1_0.x36.A 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD.t59 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X332 OUT3.t49 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND.t1284 GND.t1283 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X333 a_77881_n43295# 16to4_PriorityEncoder_v0p0p1_0.x5.x16.C a_77775_n43295# GND.t687 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X334 VV6.t12 VV5.t13 GND.t289 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X335 VDD.t939 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t113 VDD.t938 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X336 VDD.t1227 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t115 VDD.t1226 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X337 VV2.t15 VV1.t15 GND.t299 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X338 GND.t235 16to4_PriorityEncoder_v0p0p1_0.x29.A 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND.t234 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X339 VV2.t16 w_55000_n79150# error sky130_fd_pr__cap_var_lvt w=2 l=0.18
X340 w_55000_n41350# VIN.t9 a_53630_n41796# GND.t1094 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X341 GND.t1340 frontAnalog_v0p0p1_0.x65.X frontAnalog_v0p0p1_0.RSfetsym_0.x2.Y GND.t1339 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X342 frontAnalog_v0p0p1_11.RSfetsym_0.x2.Y frontAnalog_v0p0p1_11.x65.X GND.t31 GND.t30 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X343 a_77723_n50057# 16to4_PriorityEncoder_v0p0p1_0.x3.EI a_77637_n50057# GND.t386 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X344 GND.t1548 16to4_PriorityEncoder_v0p0p1_0.x5.x19.D a_77881_n44779# GND.t247 sky130_fd_pr__nfet_01v8 ad=0.196 pd=1.33 as=0.0693 ps=0.75 w=0.42 l=0.15
X345 frontAnalog_v0p0p1_7.x63.A.t0 frontAnalog_v0p0p1_7.x65.A.t6 a_55268_n36336# GND.t574 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X346 VV1.t4 VL.t2 GND.t417 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X347 VV11.t15 VV10.t15 GND.t244 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X348 I0.t4 frontAnalog_v0p0p1_15.RSfetsym_0.x2.Y GND.t1423 GND.t1422 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.25
X349 OUT1.t53 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND.t828 GND.t827 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X350 a_77775_n44527# I9.t5 a_77687_n44527# GND.t511 sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
X351 I9.t4 frontAnalog_v0p0p1_7.RSfetsym_0.QN.t5 VDD.t640 VDD.t639 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.3
X352 a_59578_n8370# frontAnalog_v0p0p1_0.x65.X frontAnalog_v0p0p1_0.RSfetsym_0.QN.t1 GND.t1338 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.315 ps=2.72 w=1 l=0.15
X353 GND.t990 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t52 GND.t989 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X354 VDD.t937 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t112 VDD.t936 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X355 a_78147_n41309# 16to4_PriorityEncoder_v0p0p1_0.x5.x22.A a_78065_n41309# VDD.t290 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X356 VDD.t192 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t116 VDD.t191 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X357 OUT1.t52 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND.t826 GND.t825 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X358 OUT3.t48 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND.t1282 GND.t1281 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X359 I1.t1 R1.t4 VDD.t564 VDD.t563 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.25
X360 VV9.t8 VV8.t6 GND.t417 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X361 16to4_PriorityEncoder_v0p0p1_0.x36.Y 16to4_PriorityEncoder_v0p0p1_0.x36.A GND.t57 GND.t56 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X362 16to4_PriorityEncoder_v0p0p1_0.x36.Y 16to4_PriorityEncoder_v0p0p1_0.x36.A VDD.t58 VDD.t57 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X363 GND.t822 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t51 GND.t821 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X364 frontAnalog_v0p0p1_12.RSfetsym_0.x1.Y frontAnalog_v0p0p1_12.x63.X GND.t20 GND.t16 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X365 a_59577_n62883# frontAnalog_v0p0p1_11.x63.X I4.t0 GND.t9 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X366 I8.t0 frontAnalog_v0p0p1_1.RSfetsym_0.x2.Y GND.t1323 GND.t1060 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.25
X367 GND.t184 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t51 GND.t183 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X368 16to4_PriorityEncoder_v0p0p1_0.x3.x15.X a_77605_n51335# GND.t1027 GND.t1026 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.196 ps=1.33 w=0.65 l=0.15
X369 16to4_PriorityEncoder_v0p0p1_0.x43.Y 16to4_PriorityEncoder_v0p0p1_0.x43.A GND.t352 GND.t351 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X370 OUT0.t50 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND.t182 GND.t181 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X371 VDD.t1025 CLK.t13 w_55000_n56928# GND.t1071 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X372 GND.t820 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t50 GND.t819 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X373 a_53630_n47196# frontAnalog_v0p0p1_10.IB.t7 GND.t308 GND.t296 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X374 I9.t1 frontAnalog_v0p0p1_7.x63.X VDD.t585 VDD.t582 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.25
X375 OUT1.t120 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD.t765 VDD.t764 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X376 frontAnalog_v0p0p1_15.RSfetsym_0.x1.Y R0.t3 VDD.t1322 VDD.t1006 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X377 VDD.t1372 frontAnalog_v0p0p1_9.x65.X frontAnalog_v0p0p1_9.RSfetsym_0.x2.Y VDD.t1368 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X378 VDD.t783 frontAnalog_v0p0p1_1.x63.A.t5 frontAnalog_v0p0p1_1.x65.A.t1 VDD.t514 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X379 OUT2.t111 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD.t935 VDD.t934 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X380 frontAnalog_v0p0p1_6.RSfetsym_0.x1.Y frontAnalog_v0p0p1_6.x63.X GND.t588 GND.t584 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X381 frontAnalog_v0p0p1_13.RSfetsym_0.x2.Y frontAnalog_v0p0p1_13.x65.X GND.t1502 GND.t1501 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X382 16to4_PriorityEncoder_v0p0p1_0.x5.x14.A a_77637_n40777# VDD.t540 VDD.t539 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.167 ps=1.39 w=1 l=0.15
X383 VDD.t763 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t119 VDD.t762 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X384 16to4_PriorityEncoder_v0p0p1_0.x34.A a_82906_n43855# VDD.t1432 VDD.t1431 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.146 ps=1.34 w=1 l=0.15
X385 frontAnalog_v0p0p1_14.RSfetsym_0.QN.t0 I1.t5 VDD.t280 VDD.t279 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.3
X386 frontAnalog_v0p0p1_10.x65.X a_57123_n56559# GND.t1117 GND.t1104 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X387 GND.t1412 I4.t6 a_59578_n62370# GND.t1411 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X388 GND.t246 frontAnalog_v0p0p1_9.RSfetsym_0.QN.t6 a_59577_n52083# GND.t245 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X389 GND.t1278 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t47 GND.t1277 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X390 16to4_PriorityEncoder_v0p0p1_0.x5.x4.A VDD.t1505 GND.t694 GND.t693 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X391 a_77775_n52567# I1.t6 a_77687_n52567# GND.t67 sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
X392 VV10.t4 VV9.t2 GND.t299 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X393 a_16719_n13117.t20 a_16599_n13205.t7 a_16541_n13117.t4 GND.t1313 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X394 VDD.t190 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t115 VDD.t189 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X395 VDD.t991 16to4_PriorityEncoder_v0p0p1_0.x28.A 16to4_PriorityEncoder_v0p0p1_0.x29.A VDD.t990 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X396 VDD.t1379 CLK.t14 w_55000_n13728# GND.t1128 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X397 OUT3.t46 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND.t1280 GND.t1279 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X398 VV3.t2 VV2.t3 GND.t257 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X399 OUT0.t49 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND.t180 GND.t179 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X400 OUT2.t51 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND.t988 GND.t987 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X401 VV14.t2 VV13.t3 GND.t244 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X402 VV13.t8 VV12.t9 GND.t299 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X403 16to4_PriorityEncoder_v0p0p1_0.x36.A 16to4_PriorityEncoder_v0p0p1_0.x35.A GND.t1142 GND.t1141 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X404 VDD.t1225 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t114 VDD.t1224 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X405 OUT0.t114 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD.t188 VDD.t187 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X406 GND.t233 16to4_PriorityEncoder_v0p0p1_0.x29.A 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND.t232 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X407 OUT2.t110 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD.t931 VDD.t930 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X408 frontAnalog_v0p0p1_1.RSfetsym_0.x1.Y frontAnalog_v0p0p1_1.x63.X VDD.t1473 VDD.t1466 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X409 frontAnalog_v0p0p1_14.RSfetsym_0.x2.Y S1.t2 VDD.t1092 VDD.t420 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X410 GND.t1276 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t45 GND.t1275 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X411 GND.t350 16to4_PriorityEncoder_v0p0p1_0.x43.A 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND.t349 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X412 frontAnalog_v0p0p1_5.RSfetsym_0.x2.Y frontAnalog_v0p0p1_5.x65.X GND.t469 GND.t468 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X413 VDD.t609 frontAnalog_v0p0p1_13.x65.A.t4 a_57123_n67359# VDD.t608 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X414 frontAnalog_v0p0p1_14.RSfetsym_0.x1.Y R1.t5 GND.t866 GND.t606 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X415 VDD.t1380 CLK.t15 w_55000_n14350# GND.t563 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X416 16to4_PriorityEncoder_v0p0p1_0.x5.x16.X a_77605_n43545# VDD.t18 VDD.t17 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.312 ps=1.68 w=1 l=0.15
X417 VDD.t1116 frontAnalog_v0p0p1_10.x65.X frontAnalog_v0p0p1_10.RSfetsym_0.x2.Y VDD.t1111 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X418 OUT1.t118 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD.t761 VDD.t760 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X419 VDD.t759 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t117 VDD.t758 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X420 frontAnalog_v0p0p1_7.RSfetsym_0.QN.t4 I9.t6 VDD.t1425 VDD.t639 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.3
X421 frontAnalog_v0p0p1_3.x65.X a_57123_n13359# GND.t1443 GND.t1357 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X422 GND.t1385 frontAnalog_v0p0p1_15.x63.A.t6 a_57123_n85079# GND.t438 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X423 VV11.t11 VV10.t12 GND.t401 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X424 OUT3.t44 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND.t1274 GND.t1273 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X425 VDD.t281 I1.t7 a_77605_n52567# VDD.t75 sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X426 VV15.t6 VV14.t5 GND.t80 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X427 GND.t1469 16to4_PriorityEncoder_v0p0p1_0.x22.A 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND.t1468 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X428 OUT2.t109 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD.t929 VDD.t928 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X429 frontAnalog_v0p0p1_7.RSfetsym_0.x2.Y frontAnalog_v0p0p1_7.x65.X VDD.t1302 VDD.t1297 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X430 OUT0.t113 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD.t186 VDD.t185 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X431 GND.t818 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t49 GND.t817 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X432 frontAnalog_v0p0p1_7.RSfetsym_0.x1.Y frontAnalog_v0p0p1_7.x63.X GND.t634 GND.t629 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X433 VDD.t927 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t108 VDD.t926 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X434 16to4_PriorityEncoder_v0p0p1_0.x29.Y 16to4_PriorityEncoder_v0p0p1_0.x29.A GND.t231 GND.t230 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X435 OUT0.t48 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND.t178 GND.t177 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X436 16to4_PriorityEncoder_v0p0p1_0.x29.Y 16to4_PriorityEncoder_v0p0p1_0.x29.A VDD.t246 VDD.t245 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X437 GND.t660 frontAnalog_v0p0p1_1.x63.A.t6 a_57123_n41879# GND.t659 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X438 frontAnalog_v0p0p1_11.RSfetsym_0.QN.t1 frontAnalog_v0p0p1_11.x65.X VDD.t34 VDD.t30 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.25
X439 VDD.t1478 I6.t6 a_77637_n50057# VDD.t362 sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X440 a_16719_n13117.t19 a_16599_n13205.t8 a_16541_n13117.t3 GND.t1314 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X441 frontAnalog_v0p0p1_2.RSfetsym_0.x2.Y frontAnalog_v0p0p1_2.x65.X VDD.t1035 VDD.t1028 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X442 a_77723_n40777# VDD.t1506 a_77637_n40777# GND.t691 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X443 OUT0.t47 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND.t176 GND.t175 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X444 16to4_PriorityEncoder_v0p0p1_0.x3.EI 16to4_PriorityEncoder_v0p0p1_0.x5.EO VDD.t537 VDD.t536 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X445 frontAnalog_v0p0p1_8.RSfetsym_0.x1.Y frontAnalog_v0p0p1_8.x63.X VDD.t1002 VDD.t997 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X446 GND.t1272 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t43 GND.t1271 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X447 GND.t174 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t46 GND.t173 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X448 GND.t55 16to4_PriorityEncoder_v0p0p1_0.x36.A 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND.t54 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X449 VDD.t1410 16to4_PriorityEncoder_v0p0p1_0.x22.A 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD.t1409 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X450 GND.t1427 I13.t8 a_77723_n41087# GND.t539 sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X451 VIN.t10 w_55000_n19128# error sky130_fd_pr__cap_var_lvt w=2 l=0.18
X452 frontAnalog_v0p0p1_15.x63.A.t2 frontAnalog_v0p0p1_15.x65.A.t5 VDD.t408 VDD.t407 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X453 VDD.t1271 frontAnalog_v0p0p1_0.x65.X frontAnalog_v0p0p1_0.RSfetsym_0.QN.t3 VDD.t1264 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.25
X454 16to4_PriorityEncoder_v0p0p1_0.x3.x16.X a_77605_n51585# VDD.t554 VDD.t553 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.312 ps=1.68 w=1 l=0.15
X455 VDD.t925 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t107 VDD.t924 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X456 VDD.t319 16to4_PriorityEncoder_v0p0p1_0.x43.A 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD.t318 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X457 a_53630_n57996# frontAnalog_v0p0p1_10.IB.t8 GND.t309 GND.t296 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X458 frontAnalog_v0p0p1_14.x63.A.t1 CLK.t16 w_55000_n79150# VDD.t815 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X459 OUT1.t116 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD.t757 VDD.t756 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X460 OUT0.t112 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD.t184 VDD.t183 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X461 GND.t172 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t45 GND.t171 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X462 VDD.t244 16to4_PriorityEncoder_v0p0p1_0.x29.A 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD.t243 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X463 GND.t1500 frontAnalog_v0p0p1_13.x65.X frontAnalog_v0p0p1_13.RSfetsym_0.x2.Y GND.t1499 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X464 16to4_PriorityEncoder_v0p0p1_0.x3.x19.D I6.t7 GND.t1538 GND.t1537 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X465 frontAnalog_v0p0p1_4.x65.A.t0 CLK.t17 frontAnalog_v0p0p1_4.x63.A.t1 VDD.t1381 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X466 a_59578_n73170# frontAnalog_v0p0p1_12.x65.X frontAnalog_v0p0p1_12.RSfetsym_0.QN.t0 GND.t398 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.315 ps=2.72 w=1 l=0.15
X467 OUT0.t111 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD.t182 VDD.t181 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X468 VV16.t2 VV15.t0 GND.t250 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X469 a_77605_n52567# 16to4_PriorityEncoder_v0p0p1_0.x3.x19.C VDD.t76 VDD.t75 sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.109 ps=1.36 w=0.42 l=0.15
X470 GND.t1270 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t42 GND.t1269 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X471 VV14.t7 VV13.t5 GND.t401 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X472 frontAnalog_v0p0p1_1.x63.A.t1 frontAnalog_v0p0p1_1.x65.A.t5 VDD.t1355 VDD.t1075 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X473 VDD.t180 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t110 VDD.t179 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X474 OUT1.t48 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND.t816 GND.t815 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X475 OUT3.t41 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND.t1268 GND.t1267 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X476 frontAnalog_v0p0p1_8.x65.X a_57123_n45759# VDD.t1306 VDD.t1305 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X477 a_53630_n14796# frontAnalog_v0p0p1_10.IB.t9 GND.t310 GND.t296 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X478 frontAnalog_v0p0p1_7.x63.A.t3 CLK.t18 w_55000_n35950# VDD.t1093 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X479 16to4_PriorityEncoder_v0p0p1_0.x36.Y 16to4_PriorityEncoder_v0p0p1_0.x36.A VDD.t56 VDD.t55 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X480 GND.t1394 frontAnalog_v0p0p1_4.x65.A.t5 a_57123_n18759# GND.t1391 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X481 frontAnalog_v0p0p1_10.RSfetsym_0.QN.t1 frontAnalog_v0p0p1_10.RSfetsym_0.x1.Y GND.t405 GND.t404 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.25
X482 GND.t1526 16to4_PriorityEncoder_v0p0p1_0.x3.x17.A a_78065_n49349# GND.t1525 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X483 GND.t504 frontAnalog_v0p0p1_2.x63.A.t6 a_57123_n4079# GND.t305 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X484 frontAnalog_v0p0p1_0.RSfetsym_0.x2.Y frontAnalog_v0p0p1_0.x65.X VDD.t1270 VDD.t1266 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X485 OUT3.t113 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD.t1223 VDD.t1222 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X486 GND.t467 frontAnalog_v0p0p1_5.x65.X frontAnalog_v0p0p1_5.RSfetsym_0.x2.Y GND.t466 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X487 GND.t867 R1.t6 frontAnalog_v0p0p1_14.RSfetsym_0.x1.Y GND.t606 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X488 VDD.t755 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t115 VDD.t754 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X489 VDD.t1310 frontAnalog_v0p0p1_12.x63.A.t4 a_57123_n74279# VDD.t1309 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X490 I12.t4 frontAnalog_v0p0p1_4.RSfetsym_0.QN.t5 VDD.t1427 VDD.t825 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.3
X491 GND.t1467 16to4_PriorityEncoder_v0p0p1_0.x22.A 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND.t1466 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X492 VDD.t572 frontAnalog_v0p0p1_4.x63.X frontAnalog_v0p0p1_4.RSfetsym_0.x1.Y VDD.t569 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X493 VDD.t178 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t109 VDD.t177 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X494 VDD.t1382 CLK.t19 w_55000_n57550# GND.t269 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X495 VDD.t1001 frontAnalog_v0p0p1_8.x63.X I7.t3 VDD.t995 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.25
X496 VDD.t14 frontAnalog_v0p0p1_11.x63.A.t4 frontAnalog_v0p0p1_11.x65.A.t0 VDD.t13 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X497 w_55000_n46128# CLK.t20 frontAnalog_v0p0p1_8.x65.A.t3 VDD.t393 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X498 16to4_PriorityEncoder_v0p0p1_0.x43.Y 16to4_PriorityEncoder_v0p0p1_0.x43.A GND.t348 GND.t347 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X499 I14.t4 frontAnalog_v0p0p1_0.RSfetsym_0.x2.Y GND.t435 GND.t434 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.25
X500 OUT1.t47 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND.t814 GND.t813 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X501 VDD.t463 I15.t5 a_77639_n42341# VDD.t462 sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X502 VV13.t16 w_55000_n19750# error sky130_fd_pr__cap_var_lvt w=2 l=0.18
X503 a_16719_n13117.t18 a_16599_n13205.t9 a_16541_n13117.t2 GND.t1315 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X504 frontAnalog_v0p0p1_13.x65.A.t3 frontAnalog_v0p0p1_13.x63.A.t5 a_55268_n68736# GND.t1124 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X505 OUT2.t106 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD.t923 VDD.t922 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X506 GND.t812 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t46 GND.t811 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X507 OUT3.t112 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD.t1221 VDD.t1220 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X508 frontAnalog_v0p0p1_3.RSfetsym_0.QN.t1 frontAnalog_v0p0p1_3.RSfetsym_0.x1.Y GND.t628 GND.t434 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.25
X509 VDD.t753 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t114 VDD.t752 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X510 GND.t633 frontAnalog_v0p0p1_7.x63.X frontAnalog_v0p0p1_7.RSfetsym_0.x1.Y GND.t629 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X511 VDD.t448 frontAnalog_v0p0p1_2.x63.X I15.t2 VDD.t441 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.25
X512 VDD.t1460 frontAnalog_v0p0p1_6.x63.A.t4 a_57123_n31079# VDD.t1459 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X513 VDD.t54 16to4_PriorityEncoder_v0p0p1_0.x36.A 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD.t53 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X514 a_53630_n74196# VV3.t16 w_55000_n73128# GND.t471 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X515 VV5.t1 VV4.t0 GND.t12 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X516 VDD.t317 16to4_PriorityEncoder_v0p0p1_0.x43.A 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD.t316 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X517 VV12.t1 VV11.t0 GND.t21 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X518 GND.t170 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t44 GND.t169 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X519 VDD.t1408 16to4_PriorityEncoder_v0p0p1_0.x22.A 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD.t1407 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X520 OUT3.t40 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND.t1266 GND.t1265 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X521 VDD.t1497 16to4_PriorityEncoder_v0p0p1_0.x3.x19.D a_77605_n52567# VDD.t75 sky130_fd_pr__pfet_01v8_hvt ad=0.312 pd=1.68 as=0.0588 ps=0.7 w=0.42 l=0.15
X522 a_55268_n52536# CLK.t21 GND.t301 GND.t300 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X523 16to4_PriorityEncoder_v0p0p1_0.x22.Y 16to4_PriorityEncoder_v0p0p1_0.x22.A GND.t1465 GND.t1464 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X524 frontAnalog_v0p0p1_5.x65.A.t3 frontAnalog_v0p0p1_5.x63.A.t5 a_55268_n25536# GND.t389 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X525 GND.t346 16to4_PriorityEncoder_v0p0p1_0.x43.A 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND.t345 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X526 GND.t986 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t50 GND.t985 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X527 VDD.t1000 frontAnalog_v0p0p1_8.x63.X frontAnalog_v0p0p1_8.RSfetsym_0.x1.Y VDD.t997 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X528 OUT3.t111 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD.t1219 VDD.t1218 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X529 VDD.t751 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t113 VDD.t750 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X530 GND.t260 frontAnalog_v0p0p1_7.RSfetsym_0.QN.t6 a_59577_n35883# GND.t259 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X531 a_53630_n30996# VV11.t16 w_55000_n29928# GND.t286 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X532 16to4_PriorityEncoder_v0p0p1_0.x36.Y 16to4_PriorityEncoder_v0p0p1_0.x36.A GND.t53 GND.t52 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X533 VDD.t1217 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t110 VDD.t1216 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X534 OUT1.t112 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD.t749 VDD.t748 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X535 VDD.t176 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t108 VDD.t175 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X536 a_55268_n9336# CLK.t22 GND.t303 GND.t302 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X537 GND.t29 frontAnalog_v0p0p1_11.x65.X frontAnalog_v0p0p1_11.RSfetsym_0.x2.Y GND.t28 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X538 VIN.t11 w_55000_n83928# error sky130_fd_pr__cap_var_lvt w=2 l=0.18
X539 frontAnalog_v0p0p1_5.RSfetsym_0.x1.Y frontAnalog_v0p0p1_5.x63.X VDD.t983 VDD.t976 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X540 VDD.t456 I7.t5 a_77639_n50381# VDD.t455 sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X541 16to4_PriorityEncoder_v0p0p1_0.x22.Y 16to4_PriorityEncoder_v0p0p1_0.x22.A VDD.t1406 VDD.t1405 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X542 VDD.t467 frontAnalog_v0p0p1_2.x63.A.t7 frontAnalog_v0p0p1_2.x65.A.t2 VDD.t466 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X543 VDD.t375 frontAnalog_v0p0p1_12.x65.X frontAnalog_v0p0p1_12.RSfetsym_0.QN.t2 VDD.t370 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.25
X544 16to4_PriorityEncoder_v0p0p1_0.x5.x21.B a_77605_n44527# GND.t704 GND.t703 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.196 ps=1.33 w=0.65 l=0.15
X545 OUT1.t45 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND.t810 GND.t809 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X546 16to4_PriorityEncoder_v0p0p1_0.x29.Y 16to4_PriorityEncoder_v0p0p1_0.x29.A VDD.t242 VDD.t241 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X547 frontAnalog_v0p0p1_2.x65.A.t1 CLK.t23 frontAnalog_v0p0p1_2.x63.A.t2 VDD.t274 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X548 VV11.t6 VV10.t3 GND.t80 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X549 VDD.t1215 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t109 VDD.t1214 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X550 OUT2.t105 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD.t921 VDD.t920 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X551 GND.t808 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t44 GND.t807 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X552 VV16.t10 VV15.t9 GND.t78 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X553 frontAnalog_v0p0p1_15.x65.A.t1 CLK.t24 frontAnalog_v0p0p1_15.x63.A.t1 VDD.t275 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X554 frontAnalog_v0p0p1_9.x63.X a_57123_n52679# VDD.t1102 VDD.t1101 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X555 OUT0.t43 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND.t168 GND.t167 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X556 w_55000_n68350# VIN.t12 a_53630_n68796# GND.t242 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X557 OUT2.t49 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND.t984 GND.t983 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X558 GND.t708 I10.t6 a_77605_n39305# GND.t267 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X559 GND.t19 frontAnalog_v0p0p1_12.x63.X frontAnalog_v0p0p1_12.RSfetsym_0.x1.Y GND.t16 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X560 VIN.t13 w_55000_n40728# error sky130_fd_pr__cap_var_lvt w=2 l=0.18
X561 VDD.t1269 frontAnalog_v0p0p1_0.x65.X frontAnalog_v0p0p1_0.RSfetsym_0.x2.Y VDD.t1266 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X562 VDD.t1283 16to4_PriorityEncoder_v0p0p1_0.x5.x4.A a_78313_n39305# VDD.t1282 sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X563 VDD.t824 I12.t5 a_77855_n40069# VDD.t823 sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X564 VV1.t9 VL.t6 GND.t299 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X565 GND.t439 frontAnalog_v0p0p1_15.x65.A.t6 a_57123_n83559# GND.t438 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X566 16to4_PriorityEncoder_v0p0p1_0.x3.x18.C I2.t6 GND.t1119 GND.t1118 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X567 a_77723_n49127# 16to4_PriorityEncoder_v0p0p1_0.x3.EI a_77637_n49127# GND.t384 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X568 VDD.t1213 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t108 VDD.t1212 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X569 GND.t229 16to4_PriorityEncoder_v0p0p1_0.x29.A 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND.t228 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X570 frontAnalog_v0p0p1_15.x63.A.t3 frontAnalog_v0p0p1_15.x65.A.t7 a_55268_n84936# GND.t440 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X571 16to4_PriorityEncoder_v0p0p1_0.x3.A2 a_78065_n49349# VDD.t968 VDD.t967 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.148 ps=1.34 w=1 l=0.15
X572 I0.t1 frontAnalog_v0p0p1_15.RSfetsym_0.QN.t5 VDD.t1061 VDD.t1060 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.3
X573 VV9.t9 VV8.t7 GND.t299 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X574 frontAnalog_v0p0p1_1.x65.A.t2 CLK.t25 frontAnalog_v0p0p1_1.x63.A.t2 VDD.t276 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X575 frontAnalog_v0p0p1_11.RSfetsym_0.x2.Y frontAnalog_v0p0p1_11.x65.X VDD.t33 VDD.t27 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X576 VDD.t1007 R0.t4 frontAnalog_v0p0p1_15.RSfetsym_0.x1.Y VDD.t1006 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X577 GND.t806 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t43 GND.t805 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X578 OUT3.t107 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD.t1211 VDD.t1210 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X579 frontAnalog_v0p0p1_2.RSfetsym_0.x1.Y frontAnalog_v0p0p1_2.x63.X VDD.t447 VDD.t443 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X580 w_55000_n25150# VIN.t14 a_53630_n25596# GND.t317 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X581 GND.t587 frontAnalog_v0p0p1_6.x63.X frontAnalog_v0p0p1_6.RSfetsym_0.x1.Y GND.t584 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X582 OUT0.t42 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND.t166 GND.t165 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X583 frontAnalog_v0p0p1_8.RSfetsym_0.x2.Y frontAnalog_v0p0p1_8.x65.X GND.t1333 GND.t1332 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X584 OUT0.t107 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD.t174 VDD.t173 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X585 a_78065_n49349# 16to4_PriorityEncoder_v0p0p1_0.x3.x22.A GND.t510 GND.t509 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X586 frontAnalog_v0p0p1_11.x63.X a_57123_n63479# GND.t1522 GND.t1042 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X587 a_53630_n3996# VV16.t16 w_55000_n2928# GND.t1091 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X588 GND.t164 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t41 GND.t163 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X589 I3.t4 frontAnalog_v0p0p1_13.RSfetsym_0.x2.Y GND.t1551 GND.t423 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.25
X590 VV1.t17 w_55000_n84550# error sky130_fd_pr__cap_var_lvt w=2 l=0.18
X591 a_78065_n41309# 16to4_PriorityEncoder_v0p0p1_0.x5.x11.X GND.t1564 GND.t1563 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X592 OUT1.t111 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD.t747 VDD.t746 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X593 GND.t1418 frontAnalog_v0p0p1_1.x65.A.t6 a_57123_n40359# GND.t659 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X594 16to4_PriorityEncoder_v0p0p1_0.x3.x21.B a_77605_n52567# GND.t502 GND.t501 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.196 ps=1.33 w=0.65 l=0.15
X595 OUT3.t39 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND.t1264 GND.t1263 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X596 OUT2.t48 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND.t982 GND.t981 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X597 a_82988_n43855# 16to4_PriorityEncoder_v0p0p1_0.x3.A2 a_82906_n43855# VDD.t819 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X598 GND.t980 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t47 GND.t979 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X599 16to4_PriorityEncoder_v0p0p1_0.x28.A 16to4_PriorityEncoder_v0p0p1_0.x1.X VDD.t380 VDD.t379 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X600 frontAnalog_v0p0p1_1.x63.A.t0 frontAnalog_v0p0p1_1.x65.A.t7 a_55268_n41736# GND.t1419 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X601 GND.t804 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t42 GND.t803 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X602 I8.t1 frontAnalog_v0p0p1_1.RSfetsym_0.QN.t5 VDD.t1428 VDD.t1307 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.3
X603 GND.t1262 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t38 GND.t1261 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X604 VDD.t1472 frontAnalog_v0p0p1_1.x63.X frontAnalog_v0p0p1_1.RSfetsym_0.x1.Y VDD.t1466 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X605 GND.t978 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t46 GND.t977 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X606 VDD.t421 S1.t3 frontAnalog_v0p0p1_14.RSfetsym_0.x2.Y VDD.t420 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X607 OUT3.t106 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD.t1209 VDD.t1208 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X608 16to4_PriorityEncoder_v0p0p1_0.x29.Y 16to4_PriorityEncoder_v0p0p1_0.x29.A GND.t227 GND.t226 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X609 frontAnalog_v0p0p1_10.RSfetsym_0.x1.Y frontAnalog_v0p0p1_10.x63.X GND.t529 GND.t525 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X610 a_59577_n46683# frontAnalog_v0p0p1_8.x63.X I7.t1 GND.t1058 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X611 VV14.t10 VV13.t11 GND.t80 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X612 a_59578_n56970# frontAnalog_v0p0p1_10.x65.X frontAnalog_v0p0p1_10.RSfetsym_0.QN.t2 GND.t1177 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.315 ps=2.72 w=1 l=0.15
X613 VV5.t11 VV4.t8 GND.t417 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X614 GND.t1120 I2.t7 a_77605_n47345# GND.t531 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X615 16to4_PriorityEncoder_v0p0p1_0.x3.x4.A 16to4_PriorityEncoder_v0p0p1_0.x3.EI VDD.t355 VDD.t354 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X616 OUT0.t106 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD.t172 VDD.t171 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X617 VDD.t1091 16to4_PriorityEncoder_v0p0p1_0.x3.x4.A a_78313_n47345# VDD.t1090 sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X618 VDD.t1207 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t105 VDD.t1206 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X619 I11.t4 frontAnalog_v0p0p1_5.RSfetsym_0.x2.Y GND.t1504 GND.t1154 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.25
X620 VV9.t17 w_55000_n41350# error sky130_fd_pr__cap_var_lvt w=2 l=0.18
X621 GND.t662 frontAnalog_v0p0p1_14.RSfetsym_0.QN.t6 a_59577_n79083# GND.t661 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X622 GND.t718 16to4_PriorityEncoder_v0p0p1_0.x5.x15.X a_78349_n43045# GND.t319 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X623 VDD.t170 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t105 VDD.t169 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X624 16to4_PriorityEncoder_v0p0p1_0.x3.x21.B a_77605_n52567# VDD.t461 VDD.t460 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.312 ps=1.68 w=1 l=0.15
X625 GND.t1260 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t37 GND.t1259 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X626 VDD.t1301 frontAnalog_v0p0p1_7.x65.X frontAnalog_v0p0p1_7.RSfetsym_0.x2.Y VDD.t1297 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X627 frontAnalog_v0p0p1_13.RSfetsym_0.x1.Y frontAnalog_v0p0p1_13.x63.X VDD.t1057 VDD.t1050 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X628 a_77775_n43295# 16to4_PriorityEncoder_v0p0p1_0.x5.x19.C a_77687_n43295# GND.t687 sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
X629 OUT2.t45 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND.t976 GND.t975 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X630 GND.t974 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t44 GND.t973 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X631 frontAnalog_v0p0p1_3.RSfetsym_0.x1.Y frontAnalog_v0p0p1_3.x63.X GND.t1512 GND.t1508 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X632 OUT1.t41 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND.t802 GND.t801 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X633 VDD.t315 16to4_PriorityEncoder_v0p0p1_0.x43.A 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD.t314 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X634 a_59578_n13770# frontAnalog_v0p0p1_3.x65.X frontAnalog_v0p0p1_3.RSfetsym_0.QN.t2 GND.t875 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.315 ps=2.72 w=1 l=0.15
X635 a_53630_n52596# frontAnalog_v0p0p1_10.IB.t10 GND.t311 GND.t296 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X636 I8.t4 frontAnalog_v0p0p1_1.x63.X VDD.t1471 VDD.t1468 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.25
X637 16to4_PriorityEncoder_v0p0p1_0.x1.X a_82906_n47995# GND.t650 GND.t649 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1 ps=0.985 w=0.65 l=0.15
X638 16to4_PriorityEncoder_v0p0p1_0.x5.x17.A a_77637_n42017# VDD.t1120 VDD.t1119 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.167 ps=1.39 w=1 l=0.15
X639 VFS.t7 VV16.t14 GND.t481 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X640 VDD.t642 frontAnalog_v0p0p1_8.x63.A.t4 frontAnalog_v0p0p1_8.x65.A.t1 VDD.t507 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X641 GND.t262 I7.t6 a_59578_n46170# GND.t261 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X642 16to4_PriorityEncoder_v0p0p1_0.x3.EI 16to4_PriorityEncoder_v0p0p1_0.x5.EO GND.t577 GND.t576 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X643 OUT0.t40 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND.t162 GND.t161 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X644 frontAnalog_v0p0p1_2.RSfetsym_0.QN.t1 frontAnalog_v0p0p1_2.RSfetsym_0.x1.Y GND.t611 GND.t610 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.25
X645 VV4.t15 VV3.t15 GND.t250 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X646 VDD.t1034 frontAnalog_v0p0p1_2.x65.X frontAnalog_v0p0p1_2.RSfetsym_0.x2.Y VDD.t1028 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X647 GND.t306 frontAnalog_v0p0p1_2.x65.A.t5 a_57123_n2559# GND.t305 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X648 frontAnalog_v0p0p1_15.RSfetsym_0.QN.t1 I0.t6 VDD.t1095 VDD.t1060 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.3
X649 VV8.t10 VV7.t9 GND.t12 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X650 GND.t1258 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t36 GND.t1257 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X651 frontAnalog_v0p0p1_11.x65.X a_57123_n61959# GND.t1043 GND.t1042 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X652 GND.t160 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t39 GND.t159 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X653 OUT1.t40 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND.t800 GND.t799 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X654 a_77605_n43295# 16to4_PriorityEncoder_v0p0p1_0.x5.x16.C VDD.t1458 VDD.t1457 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X655 VDD.t1018 frontAnalog_v0p0p1_3.x63.A.t5 a_57123_n14879# VDD.t1017 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X656 OUT3.t35 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND.t1256 GND.t1255 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X657 VDD.t1205 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t104 VDD.t1204 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X658 GND.t868 I12.t6 a_77605_n40069# GND.t555 sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X659 frontAnalog_v0p0p1_4.RSfetsym_0.QN.t1 I12.t7 VDD.t826 VDD.t825 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.3
X660 VDD.t400 frontAnalog_v0p0p1_12.x65.A.t4 a_57123_n72759# VDD.t399 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X661 GND.t1125 frontAnalog_v0p0p1_13.x63.A.t6 a_57123_n68879# GND.t1039 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X662 VDD.t919 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t104 VDD.t918 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X663 16to4_PriorityEncoder_v0p0p1_0.x43.Y 16to4_PriorityEncoder_v0p0p1_0.x43.A VDD.t313 VDD.t312 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X664 VDD.t745 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t110 VDD.t744 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X665 VDD.t32 frontAnalog_v0p0p1_11.x65.X frontAnalog_v0p0p1_11.RSfetsym_0.x2.Y VDD.t27 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X666 VDD.t446 frontAnalog_v0p0p1_2.x63.X frontAnalog_v0p0p1_2.RSfetsym_0.x1.Y VDD.t443 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X667 GND.t1463 16to4_PriorityEncoder_v0p0p1_0.x22.A 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND.t1462 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X668 frontAnalog_v0p0p1_1.RSfetsym_0.QN.t0 I8.t5 VDD.t1308 VDD.t1307 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.3
X669 OUT0.t104 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD.t168 VDD.t167 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X670 a_77605_n39305# I11.t5 GND.t709 GND.t267 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X671 GND.t158 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t38 GND.t157 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X672 frontAnalog_v0p0p1_4.RSfetsym_0.x2.Y frontAnalog_v0p0p1_4.x65.X VDD.t1424 VDD.t1419 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X673 VDD.t166 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t103 VDD.t165 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X674 OUT1.t39 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND.t798 GND.t797 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X675 frontAnalog_v0p0p1_4.RSfetsym_0.x1.Y frontAnalog_v0p0p1_4.x63.X GND.t620 GND.t615 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X676 OUT3.t34 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND.t1254 GND.t1253 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X677 a_77855_n40069# I13.t9 a_77783_n40069# VDD.t1359 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X678 VV2.t14 VV1.t13 GND.t244 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X679 OUT2.t43 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND.t972 GND.t971 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X680 VDD.t1203 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t103 VDD.t1202 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X681 a_16719_n13117.t17 a_16599_n13205.t10 a_16541_n13117.t13 GND.t1316 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X682 GND.t796 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t38 GND.t795 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X683 GND.t391 frontAnalog_v0p0p1_5.x63.A.t6 a_57123_n25679# GND.t390 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X684 frontAnalog_v0p0p1_8.RSfetsym_0.QN.t3 frontAnalog_v0p0p1_8.x65.X VDD.t1262 VDD.t1258 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.25
X685 frontAnalog_v0p0p1_1.RSfetsym_0.x1.Y frontAnalog_v0p0p1_1.x63.X GND.t1531 GND.t1527 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X686 OUT3.t102 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD.t1201 VDD.t1200 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X687 GND.t1550 I14.t5 a_77723_n42017# GND.t1549 sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X688 frontAnalog_v0p0p1_2.x63.A.t0 frontAnalog_v0p0p1_2.x65.A.t6 a_55268_n3936# GND.t307 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X689 GND.t156 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t37 GND.t155 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X690 VDD.t1404 16to4_PriorityEncoder_v0p0p1_0.x22.A 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD.t1403 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X691 VDD.t259 I8.t6 a_77855_n39305# VDD.t258 sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X692 OUT3.t33 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND.t1252 GND.t1251 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X693 16to4_PriorityEncoder_v0p0p1_0.x22.Y 16to4_PriorityEncoder_v0p0p1_0.x22.A GND.t1461 GND.t1460 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X694 VDD.t917 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t103 VDD.t916 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X695 VDD.t164 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t102 VDD.t163 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X696 a_77605_n51335# 16to4_PriorityEncoder_v0p0p1_0.x3.x16.C VDD.t1123 VDD.t1122 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X697 frontAnalog_v0p0p1_13.x63.A.t0 frontAnalog_v0p0p1_13.x65.A.t5 VDD.t610 VDD.t531 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X698 a_77881_n52819# 16to4_PriorityEncoder_v0p0p1_0.x3.x19.C a_77775_n52819# GND.t68 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X699 frontAnalog_v0p0p1_2.RSfetsym_0.QN.t4 frontAnalog_v0p0p1_2.x65.X VDD.t1033 VDD.t1031 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.25
X700 GND.t344 16to4_PriorityEncoder_v0p0p1_0.x43.A 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND.t343 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X701 frontAnalog_v0p0p1_9.RSfetsym_0.x1.Y frontAnalog_v0p0p1_9.x63.X VDD.t1338 VDD.t1333 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X702 GND.t794 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t37 GND.t793 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X703 GND.t1413 I4.t7 a_77605_n48109# GND.t263 sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X704 OUT2.t102 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD.t915 VDD.t914 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X705 OUT3.t101 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD.t1199 VDD.t1198 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X706 VDD.t743 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t109 VDD.t742 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X707 OUT1.t108 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD.t741 VDD.t740 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X708 VDD.t832 frontAnalog_v0p0p1_3.x65.X frontAnalog_v0p0p1_3.RSfetsym_0.QN.t3 VDD.t831 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.25
X709 VDD.t162 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t101 VDD.t161 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X710 I0.t0 R0.t5 VDD.t1009 VDD.t1008 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.25
X711 a_77605_n47345# I3.t5 GND.t532 GND.t531 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X712 OUT3.t32 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND.t1250 GND.t1249 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X713 frontAnalog_v0p0p1_5.x63.A.t1 frontAnalog_v0p0p1_5.x65.A.t5 VDD.t620 VDD.t524 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X714 OUT0.t36 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND.t154 GND.t153 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X715 a_59577_n3483# frontAnalog_v0p0p1_2.x63.X I15.t0 GND.t478 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X716 VV12.t8 VV11.t8 GND.t289 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X717 16to4_PriorityEncoder_v0p0p1_0.x2.X a_82906_n51645# GND.t1103 GND.t1102 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1 ps=0.985 w=0.65 l=0.15
X718 16to4_PriorityEncoder_v0p0p1_0.x22.Y 16to4_PriorityEncoder_v0p0p1_0.x22.A VDD.t1402 VDD.t1401 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X719 w_55000_n2928# CLK.t26 frontAnalog_v0p0p1_2.x65.A.t0 VDD.t277 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X720 frontAnalog_v0p0p1_6.x65.X a_57123_n29559# VDD.t1004 VDD.t1003 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X721 GND.t1248 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t31 GND.t1247 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X722 frontAnalog_v0p0p1_4.x63.A.t0 CLK.t27 w_55000_n19750# VDD.t278 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X723 VDD.t913 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t101 VDD.t912 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X724 OUT2.t100 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD.t911 VDD.t910 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X725 16to4_PriorityEncoder_v0p0p1_0.x29.Y 16to4_PriorityEncoder_v0p0p1_0.x29.A GND.t225 GND.t224 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X726 GND.t1540 I6.t8 a_77723_n50057# GND.t1539 sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X727 frontAnalog_v0p0p1_9.x65.X a_57123_n51159# VDD.t1071 VDD.t1070 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X728 VV4.t14 VV3.t14 GND.t78 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X729 frontAnalog_v0p0p1_8.x63.X a_57123_n47279# GND.t488 GND.t487 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X730 VDD.t269 frontAnalog_v0p0p1_10.x63.A.t5 a_57123_n58079# VDD.t268 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X731 OUT1.t107 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD.t739 VDD.t738 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X732 VV10.t0 VV9.t1 GND.t244 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X733 VDD.t260 CLK.t28 w_55000_n62328# GND.t269 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X734 OUT0.t35 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND.t152 GND.t151 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X735 frontAnalog_v0p0p1_11.RSfetsym_0.QN.t3 frontAnalog_v0p0p1_11.RSfetsym_0.x1.Y GND.t1182 GND.t622 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.25
X736 16to4_PriorityEncoder_v0p0p1_0.x5.x16.C I13.t10 GND.t1429 GND.t1428 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X737 a_78349_n51085# 16to4_PriorityEncoder_v0p0p1_0.x3.x16.X GND.t880 GND.t505 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X738 VDD.t1097 I0.t7 a_77855_n47345# VDD.t1096 sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X739 VV3.t0 VV2.t0 GND.t21 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X740 a_77687_n43545# I11.t6 a_77605_n43545# GND.t686 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.109 ps=1.36 w=0.42 l=0.15
X741 VV13.t2 VV12.t3 GND.t244 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X742 a_53630_n9396# frontAnalog_v0p0p1_10.IB.t11 GND.t294 GND.t293 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X743 frontAnalog_v0p0p1_12.RSfetsym_0.x2.Y frontAnalog_v0p0p1_12.x65.X GND.t397 GND.t396 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X744 VDD.t646 I11.t7 a_77605_n44779# VDD.t645 sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X745 VV8.t2 VV7.t2 GND.t417 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X746 OUT2.t99 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD.t909 VDD.t908 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X747 VDD.t982 frontAnalog_v0p0p1_5.x63.X frontAnalog_v0p0p1_5.RSfetsym_0.x1.Y VDD.t976 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X748 VV2.t12 VV1.t11 GND.t401 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X749 OUT0.t100 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD.t160 VDD.t159 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X750 VDD.t452 16to4_PriorityEncoder_v0p0p1_0.x5.x17.A a_78599_n43045# VDD.t451 sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X751 VDD.t1337 frontAnalog_v0p0p1_9.x63.X I6.t2 VDD.t1336 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.25
X752 VDD.t261 CLK.t29 w_55000_n62950# GND.t270 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X753 GND.t1246 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t30 GND.t1245 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X754 16to4_PriorityEncoder_v0p0p1_0.x2.X a_82906_n51645# VDD.t1047 VDD.t1046 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.146 ps=1.34 w=1 l=0.15
X755 w_55000_n51528# CLK.t30 frontAnalog_v0p0p1_9.x65.A.t3 VDD.t262 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X756 OUT1.t36 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND.t792 GND.t791 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X757 VDD.t52 16to4_PriorityEncoder_v0p0p1_0.x36.A 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD.t51 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X758 GND.t619 frontAnalog_v0p0p1_4.x63.X frontAnalog_v0p0p1_4.RSfetsym_0.x1.Y GND.t615 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X759 16to4_PriorityEncoder_v0p0p1_0.x3.x19.C I4.t8 GND.t1407 GND.t1406 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X760 frontAnalog_v0p0p1_12.x65.A.t1 frontAnalog_v0p0p1_12.x63.A.t5 a_55268_n74136# GND.t1379 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X761 a_53630_n57996# VV6.t16 w_55000_n56928# GND.t493 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X762 GND.t223 16to4_PriorityEncoder_v0p0p1_0.x29.A 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND.t222 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X763 VDD.t240 16to4_PriorityEncoder_v0p0p1_0.x29.A 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD.t239 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X764 OUT0.t34 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND.t150 GND.t149 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X765 frontAnalog_v0p0p1_15.RSfetsym_0.x2.Y S0.t5 VDD.t3 VDD.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X766 OUT0.t99 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD.t158 VDD.t157 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X767 GND.t1530 frontAnalog_v0p0p1_1.x63.X frontAnalog_v0p0p1_1.RSfetsym_0.x1.Y GND.t1527 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X768 frontAnalog_v0p0p1_0.x63.X a_57123_n9479# VDD.t626 VDD.t625 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X769 frontAnalog_v0p0p1_6.RSfetsym_0.x2.Y frontAnalog_v0p0p1_6.x65.X GND.t414 GND.t413 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X770 a_55268_n36336# CLK.t31 GND.t272 GND.t271 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X771 frontAnalog_v0p0p1_15.RSfetsym_0.x1.Y R0.t6 GND.t1066 GND.t1065 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X772 GND.t342 16to4_PriorityEncoder_v0p0p1_0.x43.A 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND.t341 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X773 GND.t148 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t33 GND.t147 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X774 VDD.t263 CLK.t32 w_55000_n19750# GND.t273 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X775 VFS.t6 VV16.t13 GND.t537 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X776 VV6.t10 VV5.t10 GND.t481 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X777 OUT1.t106 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD.t737 VDD.t736 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X778 OUT3.t29 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND.t1244 GND.t1243 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X779 VDD.t903 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t98 VDD.t902 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X780 GND.t1088 frontAnalog_v0p0p1_0.RSfetsym_0.QN.t5 a_59577_n8883# GND.t1087 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X781 OUT1.t105 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD.t735 VDD.t734 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X782 a_53630_n14796# VV14.t16 w_55000_n13728# GND.t491 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X783 GND.t870 frontAnalog_v0p0p1_4.RSfetsym_0.QN.t6 a_59577_n19683# GND.t869 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X784 GND.t882 I10.t7 a_59578_n29970# GND.t881 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X785 16to4_PriorityEncoder_v0p0p1_0.x36.Y 16to4_PriorityEncoder_v0p0p1_0.x36.A VDD.t50 VDD.t49 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X786 OUT3.t100 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD.t1197 VDD.t1196 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X787 VDD.t1335 frontAnalog_v0p0p1_9.x63.X frontAnalog_v0p0p1_9.RSfetsym_0.x1.Y VDD.t1333 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X788 VDD.t733 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t104 VDD.t732 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X789 frontAnalog_v0p0p1_1.RSfetsym_0.x2.Y frontAnalog_v0p0p1_1.x65.X VDD.t480 VDD.t473 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X790 R1.t1 a_57123_n79679# VDD.t1289 VDD.t1288 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X791 a_77687_n51585# I3.t6 a_77605_n51585# GND.t66 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.109 ps=1.36 w=0.42 l=0.15
X792 OUT0.t98 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD.t156 VDD.t155 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X793 a_78735_n39527# 16to4_PriorityEncoder_v0p0p1_0.x5.EO a_78649_n39527# GND.t575 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X794 GND.t1331 frontAnalog_v0p0p1_8.x65.X frontAnalog_v0p0p1_8.RSfetsym_0.x2.Y GND.t1330 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X795 16to4_PriorityEncoder_v0p0p1_0.x5.x11.X a_77637_n41087# VDD.t650 VDD.t649 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.167 ps=1.39 w=1 l=0.15
X796 VDD.t1195 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t99 VDD.t1194 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X797 VIN.t15 w_55000_n67728# error sky130_fd_pr__cap_var_lvt w=2 l=0.18
X798 GND.t695 VDD.t1507 a_77881_n43545# GND.t686 sky130_fd_pr__nfet_01v8 ad=0.196 pd=1.33 as=0.0693 ps=0.75 w=0.42 l=0.15
X799 GND.t146 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t32 GND.t145 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X800 VDD.t492 I3.t7 a_77605_n52819# VDD.t491 sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X801 a_77605_n44779# VDD.t803 VDD.t805 VDD.t804 sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.109 ps=1.36 w=0.42 l=0.15
X802 VDD.t1465 16to4_PriorityEncoder_v0p0p1_0.x3.x17.A a_78599_n51085# VDD.t1464 sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X803 GND.t1140 16to4_PriorityEncoder_v0p0p1_0.x35.A 16to4_PriorityEncoder_v0p0p1_0.x36.A GND.t1139 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X804 VDD.t154 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t97 VDD.t153 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X805 VDD.t1115 frontAnalog_v0p0p1_10.x65.X frontAnalog_v0p0p1_10.RSfetsym_0.QN.t3 VDD.t1114 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.25
X806 OUT3.t28 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND.t1242 GND.t1241 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X807 a_77855_n39305# I9.t7 a_77783_n39305# VDD.t1426 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X808 a_78097_n45737# VDD.t800 VDD.t802 VDD.t801 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X809 VDD.t1275 16to4_PriorityEncoder_v0p0p1_0.x42.A 16to4_PriorityEncoder_v0p0p1_0.x43.A VDD.t1274 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X810 VDD.t731 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t103 VDD.t730 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X811 GND.t1240 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t27 GND.t1239 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X812 VV10.t9 VV9.t11 GND.t401 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X813 OUT2.t42 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND.t970 GND.t969 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X814 frontAnalog_v0p0p1_13.x65.A.t1 CLK.t33 frontAnalog_v0p0p1_13.x63.A.t1 VDD.t264 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X815 OUT1.t35 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND.t790 GND.t789 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X816 frontAnalog_v0p0p1_7.x63.X a_57123_n36479# VDD.t1281 VDD.t1280 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X817 GND.t528 frontAnalog_v0p0p1_10.x63.X frontAnalog_v0p0p1_10.RSfetsym_0.x1.Y GND.t525 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X818 VIN.t16 w_55000_n24528# error sky130_fd_pr__cap_var_lvt w=2 l=0.18
X819 VV13.t14 VV12.t14 GND.t401 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X820 a_53630_n3996# frontAnalog_v0p0p1_10.IB.t12 GND.t295 GND.t293 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X821 16to4_PriorityEncoder_v0p0p1_0.x22.Y 16to4_PriorityEncoder_v0p0p1_0.x22.A GND.t1459 GND.t1458 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X822 a_53630_n63396# frontAnalog_v0p0p1_10.IB.t13 GND.t297 GND.t296 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X823 VDD.t152 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t96 VDD.t151 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X824 frontAnalog_v0p0p1_15.x63.A.t0 CLK.t34 w_55000_n84550# VDD.t265 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X825 GND.t1040 frontAnalog_v0p0p1_13.x65.A.t6 a_57123_n67359# GND.t1039 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X826 OUT2.t97 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD.t907 VDD.t906 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X827 frontAnalog_v0p0p1_13.x63.A.t3 frontAnalog_v0p0p1_13.x65.A.t7 a_55268_n68736# GND.t1041 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X828 GND.t395 frontAnalog_v0p0p1_12.x65.X frontAnalog_v0p0p1_12.RSfetsym_0.x2.Y GND.t394 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X829 16to4_PriorityEncoder_v0p0p1_0.x36.A 16to4_PriorityEncoder_v0p0p1_0.x35.A VDD.t1083 VDD.t1082 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X830 VDD.t238 16to4_PriorityEncoder_v0p0p1_0.x29.A 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD.t237 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X831 frontAnalog_v0p0p1_5.x65.A.t1 CLK.t35 frontAnalog_v0p0p1_5.x63.A.t3 VDD.t414 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X832 I3.t3 frontAnalog_v0p0p1_13.RSfetsym_0.QN.t5 VDD.t1109 VDD.t1108 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.3
X833 VDD.t1056 frontAnalog_v0p0p1_13.x63.X frontAnalog_v0p0p1_13.RSfetsym_0.x1.Y VDD.t1050 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X834 frontAnalog_v0p0p1_8.RSfetsym_0.x2.Y frontAnalog_v0p0p1_8.x65.X VDD.t1261 VDD.t1256 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X835 16to4_PriorityEncoder_v0p0p1_0.x5.x15.X a_77605_n43295# GND.t407 GND.t406 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.196 ps=1.33 w=0.65 l=0.15
X836 GND.t1511 frontAnalog_v0p0p1_3.x63.X frontAnalog_v0p0p1_3.RSfetsym_0.x1.Y GND.t1508 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X837 GND.t540 I12.t8 a_77723_n40777# GND.t539 sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X838 a_78735_n47567# 16to4_PriorityEncoder_v0p0p1_0.x3.EO a_78649_n47567# GND.t675 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X839 GND.t385 16to4_PriorityEncoder_v0p0p1_0.x3.EI a_77881_n51585# GND.t66 sky130_fd_pr__nfet_01v8 ad=0.196 pd=1.33 as=0.0693 ps=0.75 w=0.42 l=0.15
X840 a_77605_n52819# 16to4_PriorityEncoder_v0p0p1_0.x3.EI VDD.t353 VDD.t328 sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.109 ps=1.36 w=0.42 l=0.15
X841 VV5.t3 VV4.t2 GND.t299 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X842 16to4_PriorityEncoder_v0p0p1_0.x43.Y 16to4_PriorityEncoder_v0p0p1_0.x43.A VDD.t311 VDD.t310 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X843 VV4.t17 w_55000_n68350# error sky130_fd_pr__cap_var_lvt w=2 l=0.18
X844 OUT0.t31 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND.t144 GND.t143 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X845 VDD.t1490 16to4_PriorityEncoder_v0p0p1_0.x5.x19.D a_77605_n44779# VDD.t1489 sky130_fd_pr__pfet_01v8_hvt ad=0.312 pd=1.68 as=0.0588 ps=0.7 w=0.42 l=0.15
X846 GND.t521 frontAnalog_v0p0p1_5.x65.A.t6 a_57123_n24159# GND.t390 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X847 frontAnalog_v0p0p1_9.RSfetsym_0.x2.Y frontAnalog_v0p0p1_9.x65.X GND.t1439 GND.t1438 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X848 16to4_PriorityEncoder_v0p0p1_0.x22.Y 16to4_PriorityEncoder_v0p0p1_0.x22.A VDD.t1400 VDD.t1399 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X849 frontAnalog_v0p0p1_5.x63.A.t0 frontAnalog_v0p0p1_5.x65.A.t7 a_55268_n25536# GND.t522 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X850 a_78097_n53777# 16to4_PriorityEncoder_v0p0p1_0.x3.EI VDD.t352 VDD.t351 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X851 GND.t1457 16to4_PriorityEncoder_v0p0p1_0.x22.A 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND.t1456 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X852 a_77855_n47345# I1.t8 a_77783_n47345# VDD.t1107 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X853 GND.t412 frontAnalog_v0p0p1_6.x65.X frontAnalog_v0p0p1_6.RSfetsym_0.x2.Y GND.t411 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X854 GND.t1067 R0.t7 frontAnalog_v0p0p1_15.RSfetsym_0.x1.Y GND.t1065 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X855 I11.t0 frontAnalog_v0p0p1_5.RSfetsym_0.QN.t5 VDD.t1476 VDD.t424 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.3
X856 VDD.t729 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t102 VDD.t728 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X857 a_78599_n43045# 16to4_PriorityEncoder_v0p0p1_0.x5.x22.A a_78527_n43045# VDD.t289 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X858 OUT2.t41 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND.t968 GND.t967 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X859 VDD.t1193 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t98 VDD.t1192 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X860 16to4_PriorityEncoder_v0p0p1_0.x29.Y 16to4_PriorityEncoder_v0p0p1_0.x29.A VDD.t236 VDD.t235 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X861 16to4_PriorityEncoder_v0p0p1_0.x5.x15.X a_77605_n43295# VDD.t382 VDD.t381 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.312 ps=1.68 w=1 l=0.15
X862 I3.t2 frontAnalog_v0p0p1_13.x63.X VDD.t1055 VDD.t1052 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.25
X863 a_53630_n79596# frontAnalog_v0p0p1_10.IB.t14 GND.t298 GND.t296 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X864 VV15.t13 VV14.t13 GND.t250 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X865 OUT3.t97 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD.t1191 VDD.t1190 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X866 VV12.t17 w_55000_n25150# error sky130_fd_pr__cap_var_lvt w=2 l=0.18
X867 frontAnalog_v0p0p1_11.RSfetsym_0.x1.Y frontAnalog_v0p0p1_11.x63.X GND.t8 GND.t4 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X868 OUT0.t95 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD.t150 VDD.t149 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X869 I10.t4 frontAnalog_v0p0p1_6.RSfetsym_0.x2.Y GND.t1477 GND.t635 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.25
X870 GND.t1116 frontAnalog_v0p0p1_15.RSfetsym_0.QN.t6 a_59577_n84483# GND.t1115 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X871 VDD.t1398 16to4_PriorityEncoder_v0p0p1_0.x22.A 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD.t1397 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X872 VDD.t48 16to4_PriorityEncoder_v0p0p1_0.x36.A 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD.t47 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X873 VDD.t1423 frontAnalog_v0p0p1_4.x65.X frontAnalog_v0p0p1_4.RSfetsym_0.x2.Y VDD.t1419 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X874 16to4_PriorityEncoder_v0p0p1_0.x3.x14.A a_77637_n48817# GND.t1505 GND.t1023 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.112 ps=1.04 w=0.65 l=0.15
X875 OUT2.t40 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND.t966 GND.t965 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X876 VDD.t286 I9.t8 a_77605_n44527# VDD.t285 sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X877 I11.t3 frontAnalog_v0p0p1_5.x63.X VDD.t981 VDD.t978 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.25
X878 a_53630_n36396# frontAnalog_v0p0p1_10.IB.t15 GND.t710 GND.t296 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X879 16to4_PriorityEncoder_v0p0p1_0.x3.x2.X a_77605_n48109# GND.t674 GND.t673 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.102 ps=0.99 w=0.65 l=0.15
X880 frontAnalog_v0p0p1_12.RSfetsym_0.x1.Y frontAnalog_v0p0p1_12.x63.X VDD.t26 VDD.t19 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X881 VDD.t1461 frontAnalog_v0p0p1_6.x63.A.t5 frontAnalog_v0p0p1_6.x65.A.t1 VDD.t1087 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X882 OUT3.t96 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD.t1189 VDD.t1188 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X883 a_16541_n13117.t0 GND.t658 GND.t657 sky130_fd_pr__res_xhigh_po_5p73 l=85.8
X884 VV2.t13 VV1.t12 GND.t80 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X885 VDD.t1496 16to4_PriorityEncoder_v0p0p1_0.x3.x19.D a_77605_n52819# VDD.t1495 sky130_fd_pr__pfet_01v8_hvt ad=0.312 pd=1.68 as=0.0588 ps=0.7 w=0.42 l=0.15
X886 GND.t322 16to4_PriorityEncoder_v0p0p1_0.x5.x22.A a_78525_n45515# GND.t321 sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X887 frontAnalog_v0p0p1_13.RSfetsym_0.QN.t1 I3.t8 VDD.t1291 VDD.t1108 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.3
X888 GND.t1387 I6.t9 a_59578_n51570# GND.t1386 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X889 frontAnalog_v0p0p1_8.x65.X a_57123_n45759# GND.t1378 GND.t487 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X890 GND.t457 frontAnalog_v0p0p1_1.RSfetsym_0.QN.t6 a_59577_n41283# GND.t456 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X891 OUT0.t30 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND.t142 GND.t141 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X892 16to4_PriorityEncoder_v0p0p1_0.x36.Y 16to4_PriorityEncoder_v0p0p1_0.x36.A GND.t51 GND.t50 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X893 a_78599_n51085# 16to4_PriorityEncoder_v0p0p1_0.x3.x22.A a_78527_n51085# VDD.t471 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X894 OUT1.t101 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD.t727 VDD.t726 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X895 w_55000_n3550# VIN.t17 a_53630_n3996# GND.t1091 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X896 VV6.t3 VV5.t5 GND.t537 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X897 16to4_PriorityEncoder_v0p0p1_0.x3.x15.X a_77605_n51335# VDD.t975 VDD.t974 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.312 ps=1.68 w=1 l=0.15
X898 16to4_PriorityEncoder_v0p0p1_0.x43.Y 16to4_PriorityEncoder_v0p0p1_0.x43.A VDD.t309 VDD.t308 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X899 frontAnalog_v0p0p1_6.RSfetsym_0.x1.Y frontAnalog_v0p0p1_6.x63.X VDD.t550 VDD.t543 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X900 VDD.t1349 frontAnalog_v0p0p1_10.x65.A.t4 a_57123_n56559# VDD.t1348 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X901 VDD.t966 16to4_PriorityEncoder_v0p0p1_0.x3.x14.A a_78315_n49349# VDD.t470 sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X902 frontAnalog_v0p0p1_0.RSfetsym_0.x1.Y frontAnalog_v0p0p1_0.x63.X VDD.t84 VDD.t77 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X903 frontAnalog_v0p0p1_3.RSfetsym_0.x2.Y frontAnalog_v0p0p1_3.x65.X GND.t874 GND.t873 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X904 frontAnalog_v0p0p1_13.RSfetsym_0.x1.Y frontAnalog_v0p0p1_13.x63.X GND.t1112 GND.t1110 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X905 VV7.t6 VV6.t7 GND.t12 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X906 GND.t788 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t34 GND.t787 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X907 VDD.t1260 frontAnalog_v0p0p1_8.x65.X frontAnalog_v0p0p1_8.RSfetsym_0.x2.Y VDD.t1256 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X908 GND.t625 16to4_PriorityEncoder_v0p0p1_0.x5.x2.X a_78159_n39549# GND.t624 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X909 frontAnalog_v0p0p1_5.RSfetsym_0.QN.t1 I11.t8 VDD.t425 VDD.t424 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.3
X910 VV1.t6 VL.t4 GND.t244 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X911 GND.t1380 frontAnalog_v0p0p1_12.x63.A.t6 a_57123_n74279# GND.t665 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X912 OUT2.t39 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND.t964 GND.t963 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X913 VDD.t1187 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t95 VDD.t1186 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X914 16to4_PriorityEncoder_v0p0p1_0.x5.x19.D I14.t6 GND.t1377 GND.t1376 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X915 OUT0.t94 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD.t148 VDD.t147 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X916 OUT1.t100 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD.t725 VDD.t724 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X917 w_55000_n73750# VIN.t18 a_53630_n74196# GND.t471 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X918 VV9.t3 VV8.t3 GND.t244 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X919 a_77605_n44527# 16to4_PriorityEncoder_v0p0p1_0.x5.x19.C VDD.t632 VDD.t285 sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.109 ps=1.36 w=0.42 l=0.15
X920 OUT2.t38 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND.t962 GND.t961 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X921 GND.t960 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t37 GND.t959 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X922 GND.t49 16to4_PriorityEncoder_v0p0p1_0.x36.A 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND.t48 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X923 frontAnalog_v0p0p1_14.RSfetsym_0.x1.Y R1.t7 VDD.t820 VDD.t560 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X924 OUT3.t94 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD.t1185 VDD.t1184 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X925 VDD.t616 frontAnalog_v0p0p1_3.x65.A.t4 a_57123_n13359# VDD.t615 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X926 frontAnalog_v0p0p1_5.RSfetsym_0.x2.Y frontAnalog_v0p0p1_5.x65.X VDD.t439 VDD.t433 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X927 VDD.t723 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t99 VDD.t722 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X928 frontAnalog_v0p0p1_5.RSfetsym_0.x1.Y frontAnalog_v0p0p1_5.x63.X GND.t1031 GND.t1029 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X929 frontAnalog_v0p0p1_6.RSfetsym_0.QN.t1 frontAnalog_v0p0p1_6.x65.X VDD.t388 VDD.t383 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.25
X930 VDD.t1183 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t93 VDD.t1182 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X931 VDD.t307 16to4_PriorityEncoder_v0p0p1_0.x43.A 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD.t306 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X932 GND.t508 16to4_PriorityEncoder_v0p0p1_0.x3.x22.A a_78525_n53555# GND.t507 sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X933 frontAnalog_v0p0p1_0.x65.X a_57123_n7959# VDD.t556 VDD.t555 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X934 GND.t1518 frontAnalog_v0p0p1_6.x63.A.t6 a_57123_n31079# GND.t714 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X935 frontAnalog_v0p0p1_9.RSfetsym_0.QN.t3 frontAnalog_v0p0p1_9.x65.X VDD.t1371 VDD.t1366 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.25
X936 VDD.t479 frontAnalog_v0p0p1_1.x65.X frontAnalog_v0p0p1_1.RSfetsym_0.QN.t4 VDD.t476 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.25
X937 16to4_PriorityEncoder_v0p0p1_0.x5.GS a_78649_n39527# GND.t670 GND.t669 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.112 ps=1.04 w=0.65 l=0.15
X938 GND.t786 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t33 GND.t785 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X939 VV10.t6 VV9.t6 GND.t80 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X940 frontAnalog_v0p0p1_7.RSfetsym_0.x1.Y frontAnalog_v0p0p1_7.x63.X VDD.t584 VDD.t580 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X941 VV15.t15 VV14.t15 GND.t78 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X942 VV3.t8 VV2.t8 GND.t289 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X943 OUT3.t92 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD.t1181 VDD.t1180 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X944 OUT1.t32 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND.t784 GND.t783 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X945 VDD.t905 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t96 VDD.t904 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X946 VV13.t9 VV12.t10 GND.t80 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X947 frontAnalog_v0p0p1_12.x63.A.t0 frontAnalog_v0p0p1_12.x65.A.t5 VDD.t402 VDD.t401 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X948 I2.t4 frontAnalog_v0p0p1_12.RSfetsym_0.x2.Y GND.t1492 GND.t1044 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.25
X949 GND.t958 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t36 GND.t957 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X950 a_77605_n39305# I9.t9 GND.t312 GND.t267 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X951 S1.t1 a_57123_n78159# VDD.t1043 VDD.t1042 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X952 GND.t1410 16to4_PriorityEncoder_v0p0p1_0.x3.x2.X a_78159_n47589# GND.t1409 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X953 16to4_PriorityEncoder_v0p0p1_0.x3.x16.C I5.t9 VDD.t1315 VDD.t1314 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X954 16to4_PriorityEncoder_v0p0p1_0.x36.Y 16to4_PriorityEncoder_v0p0p1_0.x36.A VDD.t46 VDD.t45 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X955 a_77723_n48817# 16to4_PriorityEncoder_v0p0p1_0.x3.EI a_77637_n48817# GND.t384 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X956 frontAnalog_v0p0p1_13.x63.A.t2 CLK.t36 w_55000_n68350# VDD.t415 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X957 a_82988_n51645# 16to4_PriorityEncoder_v0p0p1_0.x3.A0 a_82906_n51645# VDD.t1045 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X958 VDD.t4 S0.t6 frontAnalog_v0p0p1_15.RSfetsym_0.x2.Y VDD.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X959 GND.t956 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t35 GND.t955 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X960 GND.t1382 I5.t10 a_77723_n49127# GND.t1381 sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X961 16to4_PriorityEncoder_v0p0p1_0.x5.GS a_78649_n39527# VDD.t607 VDD.t606 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.167 ps=1.39 w=1 l=0.15
X962 a_59578_n62370# frontAnalog_v0p0p1_11.x65.X frontAnalog_v0p0p1_11.RSfetsym_0.QN.t2 GND.t27 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.315 ps=2.72 w=1 l=0.15
X963 a_59577_n52083# frontAnalog_v0p0p1_9.x63.X I6.t4 GND.t1401 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X964 VV8.t13 VV7.t12 GND.t299 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X965 VDD.t821 R1.t8 I1.t0 VDD.t563 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.25
X966 16to4_PriorityEncoder_v0p0p1_0.x43.Y 16to4_PriorityEncoder_v0p0p1_0.x43.A GND.t340 GND.t339 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X967 frontAnalog_v0p0p1_6.x63.A.t0 frontAnalog_v0p0p1_6.x65.A.t4 VDD.t283 VDD.t282 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X968 GND.t782 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t31 GND.t781 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X969 OUT1.t30 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND.t780 GND.t779 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X970 VDD.t1488 16to4_PriorityEncoder_v0p0p1_0.x5.x19.D a_77605_n44527# VDD.t285 sky130_fd_pr__pfet_01v8_hvt ad=0.312 pd=1.68 as=0.0588 ps=0.7 w=0.42 l=0.15
X971 VDD.t1179 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t91 VDD.t1178 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X972 w_55000_n78528# CLK.t37 frontAnalog_v0p0p1_14.x65.A.t1 VDD.t416 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X973 OUT1.t98 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD.t721 VDD.t720 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X974 16to4_PriorityEncoder_v0p0p1_0.x5.A2 a_78065_n41309# GND.t1363 GND.t1362 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.102 ps=0.99 w=0.65 l=0.15
X975 frontAnalog_v0p0p1_7.x65.X a_57123_n34959# VDD.t398 VDD.t397 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X976 frontAnalog_v0p0p1_5.x63.A.t2 CLK.t38 w_55000_n25150# VDD.t368 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X977 VV1.t3 VL.t1 GND.t401 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X978 VDD.t417 CLK.t39 w_55000_n46128# GND.t447 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X979 VDD.t719 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t97 VDD.t718 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X980 frontAnalog_v0p0p1_8.RSfetsym_0.QN.t1 frontAnalog_v0p0p1_8.RSfetsym_0.x1.Y GND.t1061 GND.t1060 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.25
X981 VDD.t478 frontAnalog_v0p0p1_1.x65.X frontAnalog_v0p0p1_1.RSfetsym_0.x2.Y VDD.t473 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X982 16to4_PriorityEncoder_v0p0p1_0.x3.GS a_78649_n47567# GND.t591 GND.t590 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.112 ps=1.04 w=0.65 l=0.15
X983 OUT2.t95 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD.t901 VDD.t900 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X984 GND.t872 frontAnalog_v0p0p1_3.x65.X frontAnalog_v0p0p1_3.RSfetsym_0.x2.Y GND.t871 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X985 GND.t1238 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t26 GND.t1237 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X986 frontAnalog_v0p0p1_10.RSfetsym_0.x2.Y frontAnalog_v0p0p1_10.x65.X GND.t1176 GND.t1175 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X987 GND.t1111 frontAnalog_v0p0p1_13.x63.X frontAnalog_v0p0p1_13.RSfetsym_0.x1.Y GND.t1110 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X988 VDD.t16 frontAnalog_v0p0p1_11.x63.A.t5 a_57123_n63479# VDD.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X989 VV9.t13 VV8.t9 GND.t401 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X990 VV11.t2 VV10.t1 GND.t250 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X991 OUT1.t29 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND.t778 GND.t777 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X992 VDD.t418 CLK.t40 w_55000_n46750# GND.t448 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X993 frontAnalog_v0p0p1_2.RSfetsym_0.x1.Y frontAnalog_v0p0p1_2.x63.X GND.t477 GND.t475 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X994 VDD.t583 frontAnalog_v0p0p1_7.x63.X I9.t0 VDD.t582 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.25
X995 a_77775_n52819# I3.t9 a_77687_n52819# GND.t68 sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
X996 OUT3.t25 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND.t1236 GND.t1235 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X997 w_55000_n35328# CLK.t41 frontAnalog_v0p0p1_7.x65.A.t1 VDD.t419 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X998 GND.t140 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t29 GND.t139 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X999 VDD.t252 frontAnalog_v0p0p1_9.x63.A.t4 frontAnalog_v0p0p1_9.x65.A.t1 VDD.t251 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1000 VDD.t1177 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t90 VDD.t1176 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1001 frontAnalog_v0p0p1_2.RSfetsym_0.x2.Y frontAnalog_v0p0p1_2.x65.X GND.t1082 GND.t1081 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1002 16to4_PriorityEncoder_v0p0p1_0.x36.A 16to4_PriorityEncoder_v0p0p1_0.x35.A GND.t1138 GND.t1137 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1003 a_55268_n84936# CLK.t42 GND.t644 GND.t643 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1004 GND.t221 16to4_PriorityEncoder_v0p0p1_0.x29.A 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND.t220 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1005 VDD.t234 16to4_PriorityEncoder_v0p0p1_0.x29.A 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD.t233 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1006 a_77605_n47345# I1.t9 GND.t1166 GND.t531 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1007 frontAnalog_v0p0p1_10.x65.A.t1 frontAnalog_v0p0p1_10.x63.A.t6 a_55268_n57936# GND.t274 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1008 OUT3.t89 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD.t1175 VDD.t1174 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1009 VDD.t717 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t96 VDD.t716 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1010 VDD.t822 R1.t9 frontAnalog_v0p0p1_14.RSfetsym_0.x1.Y VDD.t560 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1011 VV7.t7 VV6.t9 GND.t417 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1012 frontAnalog_v0p0p1_13.RSfetsym_0.x2.Y frontAnalog_v0p0p1_13.x65.X VDD.t1439 VDD.t1433 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1013 GND.t1030 frontAnalog_v0p0p1_5.x63.X frontAnalog_v0p0p1_5.RSfetsym_0.x1.Y GND.t1029 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1014 a_78315_n49349# 16to4_PriorityEncoder_v0p0p1_0.x3.x11.X a_78243_n49349# VDD.t470 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X1015 VDD.t1324 frontAnalog_v0p0p1_4.x63.A.t6 a_57123_n20279# VDD.t1323 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1016 a_53630_n63396# VV5.t16 w_55000_n62328# GND.t315 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1017 16to4_PriorityEncoder_v0p0p1_0.x3.GS a_78649_n47567# VDD.t552 VDD.t551 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.167 ps=1.39 w=1 l=0.15
X1018 OUT3.t24 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND.t1234 GND.t1233 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1019 GND.t954 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t34 GND.t953 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1020 a_55268_n41736# CLK.t43 GND.t646 GND.t645 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1021 VIN.t19 w_55000_n2928# error sky130_fd_pr__cap_var_lvt w=2 l=0.18
X1022 OUT2.t94 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD.t899 VDD.t898 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1023 VDD.t146 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t93 VDD.t145 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1024 GND.t776 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t28 GND.t775 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1025 VDD.t897 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t93 VDD.t896 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1026 16to4_PriorityEncoder_v0p0p1_0.x43.Y 16to4_PriorityEncoder_v0p0p1_0.x43.A VDD.t305 VDD.t304 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1027 frontAnalog_v0p0p1_3.x65.A.t1 frontAnalog_v0p0p1_3.x63.A.t6 a_55268_n14736# GND.t1069 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1028 VDD.t715 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t95 VDD.t714 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1029 VDD.t581 frontAnalog_v0p0p1_7.x63.X frontAnalog_v0p0p1_7.RSfetsym_0.x1.Y VDD.t580 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1030 16to4_PriorityEncoder_v0p0p1_0.x29.Y 16to4_PriorityEncoder_v0p0p1_0.x29.A GND.t219 GND.t218 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1031 VDD.t895 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t92 VDD.t894 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1032 16to4_PriorityEncoder_v0p0p1_0.x5.x18.C I10.t8 GND.t884 GND.t883 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1033 16to4_PriorityEncoder_v0p0p1_0.x29.Y 16to4_PriorityEncoder_v0p0p1_0.x29.A VDD.t232 VDD.t231 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1034 GND.t138 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t28 GND.t137 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1035 OUT3.t23 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND.t1232 GND.t1231 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1036 OUT0.t27 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND.t136 GND.t135 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1037 frontAnalog_v0p0p1_0.RSfetsym_0.x2.Y frontAnalog_v0p0p1_0.x65.X GND.t1337 GND.t1336 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1038 GND.t1437 frontAnalog_v0p0p1_9.x65.X frontAnalog_v0p0p1_9.RSfetsym_0.x2.Y GND.t1436 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1039 GND.t1230 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t22 GND.t1229 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1040 VIN.t20 w_55000_n73128# error sky130_fd_pr__cap_var_lvt w=2 l=0.18
X1041 VV14.t8 VV13.t6 GND.t250 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1042 OUT3.t88 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD.t1173 VDD.t1172 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1043 VDD.t31 frontAnalog_v0p0p1_11.x65.X frontAnalog_v0p0p1_11.RSfetsym_0.QN.t0 VDD.t30 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.25
X1044 VDD.t893 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t91 VDD.t892 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1045 OUT2.t90 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD.t891 VDD.t890 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1046 VDD.t303 16to4_PriorityEncoder_v0p0p1_0.x43.A 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD.t302 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1047 OUT1.t94 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD.t713 VDD.t712 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1048 16to4_PriorityEncoder_v0p0p1_0.x1.X a_82906_n47995# VDD.t597 VDD.t596 sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.146 ps=1.34 w=1 l=0.15
X1049 a_16599_n13205.t3 a_16599_n13205.t2 GND.t1566 GND.t1565 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1050 VDD.t144 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t92 VDD.t143 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1051 frontAnalog_v0p0p1_12.x65.A.t3 CLK.t44 frontAnalog_v0p0p1_12.x63.A.t3 VDD.t590 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1052 GND.t134 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t26 GND.t133 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1053 OUT0.t25 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND.t132 GND.t131 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1054 frontAnalog_v0p0p1_1.x63.X a_57123_n41879# VDD.t520 VDD.t519 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1055 a_53630_n47196# frontAnalog_v0p0p1_10.IB.t16 GND.t711 GND.t296 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1056 w_55000_n57550# VIN.t21 a_53630_n57996# GND.t1559 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1057 GND.t7 frontAnalog_v0p0p1_11.x63.X frontAnalog_v0p0p1_11.RSfetsym_0.x1.Y GND.t4 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1058 OUT0.t91 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD.t142 VDD.t141 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1059 16to4_PriorityEncoder_v0p0p1_0.x5.x4.A VDD.t797 VDD.t799 VDD.t798 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1060 frontAnalog_v0p0p1_14.RSfetsym_0.x2.Y S1.t4 GND.t450 GND.t449 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1061 frontAnalog_v0p0p1_0.x63.A.t1 frontAnalog_v0p0p1_0.x65.A.t4 VDD.t1010 VDD.t494 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1062 GND.t1174 frontAnalog_v0p0p1_10.x65.X frontAnalog_v0p0p1_10.RSfetsym_0.x2.Y GND.t1173 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1063 OUT1.t27 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND.t774 GND.t773 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1064 VV16.t17 w_55000_n3550# error sky130_fd_pr__cap_var_lvt w=2 l=0.18
X1065 16to4_PriorityEncoder_v0p0p1_0.x29.A 16to4_PriorityEncoder_v0p0p1_0.x28.A GND.t1053 GND.t1052 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1066 OUT1.t93 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD.t711 VDD.t710 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1067 GND.t476 frontAnalog_v0p0p1_2.x63.X frontAnalog_v0p0p1_2.RSfetsym_0.x1.Y GND.t475 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1068 GND.t666 frontAnalog_v0p0p1_12.x65.A.t6 a_57123_n72759# GND.t665 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X1069 16to4_PriorityEncoder_v0p0p1_0.x5.x21.B a_77605_n44527# VDD.t636 VDD.t635 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.312 ps=1.68 w=1 l=0.15
X1070 OUT0.t24 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND.t130 GND.t129 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1071 a_16719_n13117.t16 a_16599_n13205.t11 a_16541_n13117.t12 GND.t1317 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1072 VV11.t10 VV10.t11 GND.t78 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1073 frontAnalog_v0p0p1_6.x65.A.t2 CLK.t45 frontAnalog_v0p0p1_6.x63.A.t3 VDD.t591 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1074 I2.t3 frontAnalog_v0p0p1_12.RSfetsym_0.QN.t5 VDD.t994 VDD.t332 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.3
X1075 VDD.t25 frontAnalog_v0p0p1_12.x63.X frontAnalog_v0p0p1_12.RSfetsym_0.x1.Y VDD.t19 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1076 frontAnalog_v0p0p1_9.RSfetsym_0.x2.Y frontAnalog_v0p0p1_9.x65.X VDD.t1370 VDD.t1368 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1077 w_55000_n14350# VIN.t22 a_53630_n14796# GND.t491 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1078 frontAnalog_v0p0p1_7.RSfetsym_0.x2.Y frontAnalog_v0p0p1_7.x65.X GND.t1373 GND.t1372 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1079 GND.t1455 16to4_PriorityEncoder_v0p0p1_0.x22.A 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND.t1454 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1080 VDD.t140 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t90 VDD.t139 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1081 OUT0.t89 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD.t138 VDD.t137 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1082 VDD.t1342 I4.t9 a_77855_n48109# VDD.t1341 sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X1083 VDD.t631 16to4_PriorityEncoder_v0p0p1_0.x5.x19.C a_77605_n43545# VDD.t426 sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X1084 frontAnalog_v0p0p1_9.x63.X a_57123_n52679# GND.t1162 GND.t1126 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1085 16to4_PriorityEncoder_v0p0p1_0.x43.Y 16to4_PriorityEncoder_v0p0p1_0.x43.A GND.t338 GND.t337 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1086 I5.t3 frontAnalog_v0p0p1_10.RSfetsym_0.x2.Y GND.t623 GND.t622 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.25
X1087 VV3.t17 w_55000_n73750# error sky130_fd_pr__cap_var_lvt w=2 l=0.18
X1088 OUT1.t92 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD.t709 VDD.t708 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1089 frontAnalog_v0p0p1_6.x63.A.t1 frontAnalog_v0p0p1_6.x65.A.t5 a_55268_n30936# GND.t304 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1090 OUT2.t89 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD.t889 VDD.t888 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1091 a_77687_n51335# I2.t8 a_77605_n51335# GND.t69 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.109 ps=1.36 w=0.42 l=0.15
X1092 VDD.t707 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t91 VDD.t706 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1093 I10.t0 frontAnalog_v0p0p1_6.RSfetsym_0.QN.t5 VDD.t396 VDD.t395 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.3
X1094 VDD.t549 frontAnalog_v0p0p1_6.x63.X frontAnalog_v0p0p1_6.RSfetsym_0.x1.Y VDD.t543 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1095 a_59578_n2970# frontAnalog_v0p0p1_2.x65.X frontAnalog_v0p0p1_2.RSfetsym_0.QN.t2 GND.t1080 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.315 ps=2.72 w=1 l=0.15
X1096 OUT0.t88 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD.t136 VDD.t135 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1097 VDD.t83 frontAnalog_v0p0p1_0.x63.X frontAnalog_v0p0p1_0.RSfetsym_0.x1.Y VDD.t77 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1098 frontAnalog_v0p0p1_8.RSfetsym_0.x1.Y frontAnalog_v0p0p1_8.x63.X GND.t1057 GND.t1054 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1099 GND.t128 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t23 GND.t127 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1100 a_78065_n49349# 16to4_PriorityEncoder_v0p0p1_0.x3.x11.X GND.t857 GND.t856 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1101 a_59577_n35883# frontAnalog_v0p0p1_7.x63.X I9.t2 GND.t632 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1102 a_53630_n84996# frontAnalog_v0p0p1_10.IB.t17 GND.t712 GND.t296 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1103 VDD.t1396 16to4_PriorityEncoder_v0p0p1_0.x22.A 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD.t1395 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1104 a_77637_n42017# VDD.t795 VDD.t796 VDD.t509 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X1105 I13.t0 frontAnalog_v0p0p1_3.RSfetsym_0.x2.Y GND.t548 GND.t547 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.25
X1106 VV11.t17 w_55000_n30550# error sky130_fd_pr__cap_var_lvt w=2 l=0.18
X1107 frontAnalog_v0p0p1_0.x63.A.t3 CLK.t46 w_55000_n8950# VDD.t592 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1108 GND.t1170 frontAnalog_v0p0p1_13.RSfetsym_0.QN.t6 a_59577_n68283# GND.t1169 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1109 16to4_PriorityEncoder_v0p0p1_0.x22.Y 16to4_PriorityEncoder_v0p0p1_0.x22.A GND.t1453 GND.t1452 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1110 GND.t1168 I1.t10 a_59578_n78570# GND.t1167 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1111 GND.t217 16to4_PriorityEncoder_v0p0p1_0.x29.A 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND.t216 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1112 I14.t2 frontAnalog_v0p0p1_0.x63.X VDD.t82 VDD.t80 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.25
X1113 VV1.t14 VL.t7 GND.t80 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1114 GND.t1335 frontAnalog_v0p0p1_0.x65.X frontAnalog_v0p0p1_0.RSfetsym_0.x2.Y GND.t1334 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1115 VDD.t593 CLK.t47 w_55000_n29928# GND.t549 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1116 a_16719_n13117.t15 a_16599_n13205.t12 a_16541_n13117.t11 GND.t1318 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1117 OUT3.t87 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD.t1171 VDD.t1170 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1118 VDD.t705 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t90 VDD.t704 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1119 VDD.t438 frontAnalog_v0p0p1_5.x65.X frontAnalog_v0p0p1_5.RSfetsym_0.x2.Y VDD.t433 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1120 frontAnalog_v0p0p1_10.RSfetsym_0.x1.Y frontAnalog_v0p0p1_10.x63.X VDD.t488 VDD.t483 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1121 OUT2.t33 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND.t952 GND.t951 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1122 VDD.t1169 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t86 VDD.t1168 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1123 VV9.t12 VV8.t8 GND.t80 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1124 a_53630_n41796# frontAnalog_v0p0p1_10.IB.t18 GND.t713 GND.t296 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1125 16to4_PriorityEncoder_v0p0p1_0.x3.x11.X a_77637_n49127# GND.t1024 GND.t1023 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.112 ps=1.04 w=0.65 l=0.15
X1126 I14.t3 frontAnalog_v0p0p1_0.RSfetsym_0.QN.t6 VDD.t624 VDD.t623 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.3
X1127 VDD.t74 16to4_PriorityEncoder_v0p0p1_0.x3.x19.C a_77605_n51585# VDD.t73 sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X1128 a_77605_n43545# I11.t9 VDD.t427 VDD.t426 sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.109 ps=1.36 w=0.42 l=0.15
X1129 VV14.t6 VV13.t4 GND.t78 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1130 VDD.t134 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t87 VDD.t133 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1131 GND.t950 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t32 GND.t949 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1132 GND.t1536 frontAnalog_v0p0p1_5.RSfetsym_0.QN.t6 a_59577_n25083# GND.t1535 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1133 frontAnalog_v0p0p1_6.x65.X a_57123_n29559# GND.t1062 GND.t581 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1134 16to4_PriorityEncoder_v0p0p1_0.x3.x19.D I6.t10 VDD.t1320 VDD.t1319 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1135 GND.t314 I9.t10 a_59578_n35370# GND.t313 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1136 16to4_PriorityEncoder_v0p0p1_0.x5.x2.X a_77605_n40069# VDD.t1492 VDD.t1491 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.148 ps=1.34 w=1 l=0.15
X1137 a_77605_n52567# 16to4_PriorityEncoder_v0p0p1_0.x3.x18.C VDD.t378 VDD.t75 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X1138 16to4_PriorityEncoder_v0p0p1_0.x22.Y 16to4_PriorityEncoder_v0p0p1_0.x22.A VDD.t1394 VDD.t1393 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1139 R0.t1 a_57123_n85079# VDD.t482 VDD.t481 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1140 frontAnalog_v0p0p1_3.RSfetsym_0.x1.Y frontAnalog_v0p0p1_3.x63.X VDD.t1451 VDD.t1444 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1141 VDD.t1167 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t85 VDD.t1166 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1142 16to4_PriorityEncoder_v0p0p1_0.x29.Y 16to4_PriorityEncoder_v0p0p1_0.x29.A VDD.t230 VDD.t229 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1143 GND.t383 16to4_PriorityEncoder_v0p0p1_0.x3.EI a_77881_n51335# GND.t69 sky130_fd_pr__nfet_01v8 ad=0.196 pd=1.33 as=0.0693 ps=0.75 w=0.42 l=0.15
X1144 16to4_PriorityEncoder_v0p0p1_0.x3.x17.A a_77637_n50057# VDD.t365 VDD.t364 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.167 ps=1.39 w=1 l=0.15
X1145 a_77881_n44779# 16to4_PriorityEncoder_v0p0p1_0.x5.x19.C a_77775_n44779# GND.t247 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X1146 16to4_PriorityEncoder_v0p0p1_0.x3.x20.X a_77605_n53805# GND.t1164 GND.t1163 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X1147 VV12.t4 VV11.t4 GND.t481 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1148 OUT0.t22 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND.t126 GND.t125 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1149 VDD.t1364 frontAnalog_v0p0p1_11.x65.A.t4 a_57123_n61959# VDD.t1363 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1150 16to4_PriorityEncoder_v0p0p1_0.x22.A 16to4_PriorityEncoder_v0p0p1_0.x21.A GND.t372 GND.t371 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1151 GND.t276 frontAnalog_v0p0p1_10.x63.A.t7 a_57123_n58079# GND.t275 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X1152 frontAnalog_v0p0p1_14.RSfetsym_0.QN.t1 S1.t5 VDD.t423 VDD.t422 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.25
X1153 VDD.t1369 frontAnalog_v0p0p1_9.x65.X frontAnalog_v0p0p1_9.RSfetsym_0.x2.Y VDD.t1368 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1154 a_77783_n40069# I14.t7 a_77687_n40069# VDD.t1303 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X1155 VDD.t1165 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t84 VDD.t1164 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1156 VDD.t594 CLK.t48 w_55000_n8328# GND.t552 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1157 OUT1.t89 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD.t703 VDD.t702 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1158 VV5.t6 VV4.t5 GND.t244 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1159 GND.t948 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t31 GND.t947 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1160 OUT3.t83 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD.t1163 VDD.t1162 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1161 a_77605_n51585# I3.t10 VDD.t1292 VDD.t73 sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.109 ps=1.36 w=0.42 l=0.15
X1162 VDD.t228 16to4_PriorityEncoder_v0p0p1_0.x29.A 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD.t227 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1163 GND.t1070 frontAnalog_v0p0p1_3.x63.A.t7 a_57123_n14879# GND.t676 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X1164 VDD.t1072 CLK.t49 w_55000_n8950# GND.t1128 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1165 frontAnalog_v0p0p1_7.RSfetsym_0.QN.t3 frontAnalog_v0p0p1_7.x65.X VDD.t1300 VDD.t1295 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.25
X1166 frontAnalog_v0p0p1_12.x63.A.t1 frontAnalog_v0p0p1_12.x65.A.t7 a_55268_n74136# GND.t667 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1167 OUT0.t86 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD.t132 VDD.t131 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1168 VDD.t794 VDD.t793 a_77605_n43545# VDD.t426 sky130_fd_pr__pfet_01v8_hvt ad=0.312 pd=1.68 as=0.0588 ps=0.7 w=0.42 l=0.15
X1169 16to4_PriorityEncoder_v0p0p1_0.x22.A 16to4_PriorityEncoder_v0p0p1_0.x21.A VDD.t342 VDD.t341 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1170 VDD.t1377 16to4_PriorityEncoder_v0p0p1_0.x5.x21.B a_78097_n45737# VDD.t1376 sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X1171 frontAnalog_v0p0p1_4.RSfetsym_0.x1.Y frontAnalog_v0p0p1_4.x63.X VDD.t571 VDD.t569 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1172 a_59577_n79083# R1.t10 I1.t2 GND.t605 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1173 a_77855_n48109# I5.t11 a_77783_n48109# VDD.t1316 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X1174 a_78349_n43045# 16to4_PriorityEncoder_v0p0p1_0.x5.x16.X GND.t578 GND.t319 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X1175 GND.t946 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t30 GND.t945 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1176 a_77605_n45765# 16to4_PriorityEncoder_v0p0p1_0.x5.x19.D VDD.t1487 VDD.t1486 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X1177 GND.t772 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t26 GND.t771 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1178 frontAnalog_v0p0p1_0.RSfetsym_0.QN.t4 I14.t8 VDD.t1304 VDD.t623 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.3
X1179 frontAnalog_v0p0p1_10.x63.A.t1 frontAnalog_v0p0p1_10.x65.A.t5 VDD.t1350 VDD.t1084 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1180 GND.t1079 frontAnalog_v0p0p1_2.x65.X frontAnalog_v0p0p1_2.RSfetsym_0.x2.Y GND.t1078 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1181 a_55268_n3936# CLK.t50 GND.t1130 GND.t1129 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1182 frontAnalog_v0p0p1_1.RSfetsym_0.x1.Y frontAnalog_v0p0p1_1.x63.X VDD.t1470 VDD.t1466 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1183 OUT3.t82 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD.t1161 VDD.t1160 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1184 a_53630_n30996# frontAnalog_v0p0p1_10.IB.t19 GND.t451 GND.t296 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1185 16to4_PriorityEncoder_v0p0p1_0.x29.Y 16to4_PriorityEncoder_v0p0p1_0.x29.A GND.t215 GND.t214 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1186 GND.t1451 16to4_PriorityEncoder_v0p0p1_0.x22.A 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND.t1450 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1187 OUT3.t21 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND.t1228 GND.t1227 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1188 16to4_PriorityEncoder_v0p0p1_0.x5.x19.C I12.t9 GND.t542 GND.t541 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1189 VDD.t1438 frontAnalog_v0p0p1_13.x65.X frontAnalog_v0p0p1_13.RSfetsym_0.x2.Y VDD.t1433 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1190 a_59578_n46170# frontAnalog_v0p0p1_8.x65.X frontAnalog_v0p0p1_8.RSfetsym_0.QN.t4 GND.t1329 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.315 ps=2.72 w=1 l=0.15
X1191 VDD.t1081 16to4_PriorityEncoder_v0p0p1_0.x35.A 16to4_PriorityEncoder_v0p0p1_0.x36.A VDD.t1080 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1192 I2.t2 frontAnalog_v0p0p1_12.x63.X VDD.t24 VDD.t21 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.25
X1193 frontAnalog_v0p0p1_3.x63.A.t0 frontAnalog_v0p0p1_3.x65.A.t5 VDD.t617 VDD.t505 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1194 VDD.t816 frontAnalog_v0p0p1_14.x63.A.t6 frontAnalog_v0p0p1_14.x65.A.t3 VDD.t815 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1195 OUT3.t81 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD.t1159 VDD.t1158 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1196 frontAnalog_v0p0p1_4.x65.X a_57123_n18759# VDD.t576 VDD.t575 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1197 OUT2.t29 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND.t944 GND.t943 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1198 OUT2.t88 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD.t887 VDD.t886 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1199 VDD.t301 16to4_PriorityEncoder_v0p0p1_0.x43.A 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD.t300 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1200 OUT1.t88 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD.t701 VDD.t700 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1201 frontAnalog_v0p0p1_6.RSfetsym_0.QN.t4 frontAnalog_v0p0p1_6.RSfetsym_0.x1.Y GND.t1155 GND.t1154 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.25
X1202 VDD.t350 16to4_PriorityEncoder_v0p0p1_0.x3.EI a_77605_n51585# VDD.t73 sky130_fd_pr__pfet_01v8_hvt ad=0.312 pd=1.68 as=0.0588 ps=0.7 w=0.42 l=0.15
X1203 16to4_PriorityEncoder_v0p0p1_0.x3.A1 a_78349_n51085# GND.t1516 GND.t1026 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.102 ps=0.99 w=0.65 l=0.15
X1204 VV7.t8 VV6.t11 GND.t299 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1205 VDD.t1392 16to4_PriorityEncoder_v0p0p1_0.x22.A 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD.t1391 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1206 OUT1.t25 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND.t770 GND.t769 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1207 VDD.t644 frontAnalog_v0p0p1_8.x63.A.t5 a_57123_n47279# VDD.t643 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1208 VDD.t558 16to4_PriorityEncoder_v0p0p1_0.x3.x21.B a_78097_n53777# VDD.t557 sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X1209 VDD.t1073 CLK.t51 w_55000_n51528# GND.t448 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1210 I10.t3 frontAnalog_v0p0p1_6.x63.X VDD.t548 VDD.t545 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.25
X1211 VDD.t1094 frontAnalog_v0p0p1_7.x63.A.t5 frontAnalog_v0p0p1_7.x65.A.t3 VDD.t1093 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1212 GND.t1226 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t20 GND.t1225 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1213 a_77605_n53805# 16to4_PriorityEncoder_v0p0p1_0.x3.x19.D VDD.t1494 VDD.t1493 sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.0567 ps=0.69 w=0.42 l=0.15
X1214 frontAnalog_v0p0p1_11.RSfetsym_0.x2.Y frontAnalog_v0p0p1_11.x65.X GND.t26 GND.t25 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1215 a_55268_n68736# CLK.t52 GND.t1132 GND.t1131 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1216 OUT3.t80 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD.t1157 VDD.t1156 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1217 VV16.t15 VV15.t14 GND.t12 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1218 VDD.t1074 CLK.t53 w_55000_n52150# GND.t1071 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1219 VV5.t9 VV4.t7 GND.t401 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1220 16to4_PriorityEncoder_v0p0p1_0.x3.x18.C I2.t9 VDD.t331 VDD.t330 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1221 VDD.t1469 frontAnalog_v0p0p1_1.x63.X I8.t3 VDD.t1468 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.25
X1222 OUT3.t19 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND.t1224 GND.t1223 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1223 frontAnalog_v0p0p1_12.RSfetsym_0.QN.t4 I2.t10 VDD.t333 VDD.t332 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.3
X1224 a_77759_n53805# 16to4_PriorityEncoder_v0p0p1_0.x3.x19.D a_77687_n53805# GND.t1557 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X1225 frontAnalog_v0p0p1_9.x65.X a_57123_n51159# GND.t1127 GND.t1126 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1226 w_55000_n40728# CLK.t54 frontAnalog_v0p0p1_1.x65.A.t3 VDD.t1075 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1227 VDD.t1155 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t79 VDD.t1154 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1228 I15.t3 frontAnalog_v0p0p1_2.RSfetsym_0.x2.Y GND.t1073 GND.t688 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.25
X1229 GND.t556 I14.t9 a_77605_n40069# GND.t555 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X1230 GND.t1222 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t18 GND.t1221 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1231 frontAnalog_v0p0p1_11.x65.A.t1 frontAnalog_v0p0p1_11.x63.A.t6 a_55268_n63336# GND.t277 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1232 a_53630_n47196# VV8.t16 w_55000_n46128# GND.t1107 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1233 a_78349_n51085# 16to4_PriorityEncoder_v0p0p1_0.x3.x22.A GND.t506 GND.t505 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1234 GND.t558 I14.t10 a_59578_n8370# GND.t557 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1235 frontAnalog_v0p0p1_12.RSfetsym_0.x2.Y frontAnalog_v0p0p1_12.x65.X VDD.t374 VDD.t372 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1236 a_77637_n41087# VDD.t790 VDD.t792 VDD.t791 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X1237 a_55268_n25536# CLK.t55 GND.t1134 GND.t1133 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1238 frontAnalog_v0p0p1_12.RSfetsym_0.x1.Y frontAnalog_v0p0p1_12.x63.X GND.t18 GND.t16 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1239 a_78243_n49349# 16to4_PriorityEncoder_v0p0p1_0.x3.x17.A a_78147_n49349# VDD.t470 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X1240 GND.t1090 S1.t6 frontAnalog_v0p0p1_14.RSfetsym_0.x2.Y GND.t1089 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1241 OUT1.t24 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND.t768 GND.t767 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1242 a_82988_n47995# 16to4_PriorityEncoder_v0p0p1_0.x3.A1 a_82906_n47995# VDD.t1290 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X1243 GND.t766 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t23 GND.t765 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1244 a_77687_n40069# I15.t6 a_77605_n40069# VDD.t1013 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X1245 VDD.t570 frontAnalog_v0p0p1_4.x63.X frontAnalog_v0p0p1_4.RSfetsym_0.x1.Y VDD.t569 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1246 VDD.t1153 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t78 VDD.t1152 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1247 frontAnalog_v0p0p1_0.x65.A.t0 frontAnalog_v0p0p1_0.x63.A.t4 a_55268_n9336# GND.t258 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1248 GND.t764 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t22 GND.t763 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1249 OUT2.t87 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD.t885 VDD.t884 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1250 a_77687_n44527# 16to4_PriorityEncoder_v0p0p1_0.x5.x19.C a_77605_n44527# GND.t511 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.109 ps=1.36 w=0.42 l=0.15
X1251 GND.t1417 16to4_PriorityEncoder_v0p0p1_0.x5.A2 a_82906_n43855# GND.t1416 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X1252 VDD.t1467 frontAnalog_v0p0p1_1.x63.X frontAnalog_v0p0p1_1.RSfetsym_0.x1.Y VDD.t1466 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1253 frontAnalog_v0p0p1_15.RSfetsym_0.x1.Y R0.t8 VDD.t1326 VDD.t1006 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1254 VDD.t256 frontAnalog_v0p0p1_0.x63.A.t5 a_57123_n9479# VDD.t255 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1255 frontAnalog_v0p0p1_6.RSfetsym_0.x2.Y frontAnalog_v0p0p1_6.x65.X VDD.t387 VDD.t385 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1256 GND.t124 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t21 GND.t123 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1257 frontAnalog_v0p0p1_13.x63.X a_57123_n68879# VDD.t1106 VDD.t1105 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1258 frontAnalog_v0p0p1_6.RSfetsym_0.x1.Y frontAnalog_v0p0p1_6.x63.X GND.t586 GND.t584 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1259 GND.t1371 frontAnalog_v0p0p1_7.x65.X frontAnalog_v0p0p1_7.RSfetsym_0.x2.Y GND.t1370 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1260 VV12.t15 VV11.t14 GND.t537 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1261 a_77783_n39305# I10.t9 a_77687_n39305# VDD.t837 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X1262 VIN.t23 w_55000_n56928# error sky130_fd_pr__cap_var_lvt w=2 l=0.18
X1263 16to4_PriorityEncoder_v0p0p1_0.x22.Y 16to4_PriorityEncoder_v0p0p1_0.x22.A GND.t1449 GND.t1448 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1264 VDD.t299 16to4_PriorityEncoder_v0p0p1_0.x43.A 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD.t298 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1265 frontAnalog_v0p0p1_0.x63.X a_57123_n9479# GND.t681 GND.t598 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1266 VDD.t1259 frontAnalog_v0p0p1_8.x65.X frontAnalog_v0p0p1_8.RSfetsym_0.QN.t2 VDD.t1258 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.25
X1267 GND.t1388 I6.t11 a_77605_n48109# GND.t263 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X1268 OUT1.t21 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND.t762 GND.t761 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1269 GND.t760 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t20 GND.t759 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1270 OUT2.t86 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD.t883 VDD.t882 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1271 OUT3.t77 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD.t1151 VDD.t1150 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1272 frontAnalog_v0p0p1_10.x65.A.t2 CLK.t56 frontAnalog_v0p0p1_10.x63.A.t2 VDD.t526 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1273 frontAnalog_v0p0p1_5.x63.X a_57123_n25679# VDD.t273 VDD.t272 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1274 frontAnalog_v0p0p1_14.RSfetsym_0.x2.Y S1.t7 VDD.t1040 VDD.t420 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1275 GND.t1056 frontAnalog_v0p0p1_8.x63.X frontAnalog_v0p0p1_8.RSfetsym_0.x1.Y GND.t1054 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1276 VV8.t5 VV7.t4 GND.t244 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1277 VIN.t24 w_55000_n13728# error sky130_fd_pr__cap_var_lvt w=2 l=0.18
X1278 frontAnalog_v0p0p1_14.x63.A.t3 frontAnalog_v0p0p1_14.x65.A.t6 VDD.t1098 VDD.t416 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1279 VDD.t130 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t85 VDD.t129 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1280 VDD.t1032 frontAnalog_v0p0p1_2.x65.X frontAnalog_v0p0p1_2.RSfetsym_0.QN.t3 VDD.t1031 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.25
X1281 frontAnalog_v0p0p1_0.RSfetsym_0.x1.Y frontAnalog_v0p0p1_0.x63.X GND.t73 GND.t71 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1282 S0.t1 a_57123_n83559# VDD.t634 VDD.t633 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1283 GND.t942 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t28 GND.t941 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1284 R1.t0 a_57123_n79679# GND.t1364 GND.t1097 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1285 a_53630_n52596# frontAnalog_v0p0p1_10.IB.t20 GND.t452 GND.t296 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1286 16to4_PriorityEncoder_v0p0p1_0.x36.Y 16to4_PriorityEncoder_v0p0p1_0.x36.A VDD.t44 VDD.t43 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1287 frontAnalog_v0p0p1_12.x63.A.t2 CLK.t57 w_55000_n73750# VDD.t527 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1288 16to4_PriorityEncoder_v0p0p1_0.x22.Y 16to4_PriorityEncoder_v0p0p1_0.x22.A VDD.t1390 VDD.t1389 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1289 GND.t1220 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t17 GND.t1219 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1290 VV2.t2 VV1.t0 GND.t250 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1291 GND.t1414 frontAnalog_v0p0p1_10.x65.A.t6 a_57123_n56559# GND.t275 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X1292 OUT0.t20 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND.t122 GND.t121 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1293 a_77687_n52567# 16to4_PriorityEncoder_v0p0p1_0.x3.x19.C a_77605_n52567# GND.t67 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.109 ps=1.36 w=0.42 l=0.15
X1294 OUT3.t76 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD.t1149 VDD.t1148 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1295 frontAnalog_v0p0p1_10.x63.A.t0 frontAnalog_v0p0p1_10.x65.A.t7 a_55268_n57936# GND.t1415 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1296 GND.t24 frontAnalog_v0p0p1_11.x65.X frontAnalog_v0p0p1_11.RSfetsym_0.x2.Y GND.t23 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1297 GND.t1547 16to4_PriorityEncoder_v0p0p1_0.x5.x19.D a_77881_n44527# GND.t511 sky130_fd_pr__nfet_01v8 ad=0.196 pd=1.33 as=0.0693 ps=0.75 w=0.42 l=0.15
X1298 frontAnalog_v0p0p1_3.x65.A.t2 CLK.t58 frontAnalog_v0p0p1_3.x63.A.t2 VDD.t528 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1299 I5.t4 frontAnalog_v0p0p1_10.RSfetsym_0.QN.t5 VDD.t1330 VDD.t1317 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.3
X1300 frontAnalog_v0p0p1_7.RSfetsym_0.x2.Y frontAnalog_v0p0p1_7.x65.X VDD.t1299 VDD.t1297 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1301 VDD.t487 frontAnalog_v0p0p1_10.x63.X frontAnalog_v0p0p1_10.RSfetsym_0.x1.Y VDD.t483 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1302 VDD.t1147 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t75 VDD.t1146 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1303 VDD.t1327 R0.t9 I0.t2 VDD.t1008 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.25
X1304 VDD.t699 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t87 VDD.t698 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1305 frontAnalog_v0p0p1_4.RSfetsym_0.x2.Y frontAnalog_v0p0p1_4.x65.X GND.t1482 GND.t1481 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1306 w_55000_n83928# CLK.t59 frontAnalog_v0p0p1_15.x65.A.t0 VDD.t407 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1307 16to4_PriorityEncoder_v0p0p1_0.x5.x2.X a_77605_n40069# GND.t1553 GND.t1552 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.102 ps=0.99 w=0.65 l=0.15
X1308 a_77783_n47345# I2.t11 a_77687_n47345# VDD.t334 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X1309 frontAnalog_v0p0p1_1.x65.X a_57123_n40359# VDD.t68 VDD.t67 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1310 a_16719_n13117.t14 a_16599_n13205.t13 a_16541_n13117.t10 GND.t428 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1311 frontAnalog_v0p0p1_7.x63.X a_57123_n36479# GND.t1353 GND.t420 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1312 VV6.t17 w_55000_n57550# error sky130_fd_pr__cap_var_lvt w=2 l=0.18
X1313 OUT2.t85 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD.t881 VDD.t880 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1314 GND.t677 frontAnalog_v0p0p1_3.x65.A.t6 a_57123_n13359# GND.t676 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X1315 a_78527_n43045# 16to4_PriorityEncoder_v0p0p1_0.x5.x15.X a_78431_n43045# VDD.t651 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X1316 frontAnalog_v0p0p1_9.RSfetsym_0.QN.t0 frontAnalog_v0p0p1_9.RSfetsym_0.x1.Y GND.t1405 GND.t1404 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.25
X1317 frontAnalog_v0p0p1_2.RSfetsym_0.x2.Y frontAnalog_v0p0p1_2.x65.X VDD.t1030 VDD.t1028 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1318 VV16.t7 VV15.t7 GND.t417 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1319 frontAnalog_v0p0p1_3.x63.A.t1 frontAnalog_v0p0p1_3.x65.A.t7 a_55268_n14736# GND.t678 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1320 GND.t17 frontAnalog_v0p0p1_12.x63.X frontAnalog_v0p0p1_12.RSfetsym_0.x1.Y GND.t16 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1321 OUT1.t19 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND.t758 GND.t757 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1322 OUT2.t84 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD.t879 VDD.t878 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1323 VDD.t877 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t83 VDD.t876 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1324 VDD.t42 16to4_PriorityEncoder_v0p0p1_0.x36.A 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD.t41 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1325 OUT0.t84 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD.t128 VDD.t127 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1326 GND.t1408 I4.t10 a_77723_n48817# GND.t1381 sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X1327 I13.t1 frontAnalog_v0p0p1_3.RSfetsym_0.QN.t5 VDD.t1332 VDD.t1331 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.3
X1328 frontAnalog_v0p0p1_0.x65.X a_57123_n7959# GND.t599 GND.t598 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1329 VDD.t1450 frontAnalog_v0p0p1_3.x63.X frontAnalog_v0p0p1_3.RSfetsym_0.x1.Y VDD.t1444 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1330 a_59577_n19683# frontAnalog_v0p0p1_4.x63.X I12.t1 GND.t618 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1331 OUT0.t19 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND.t120 GND.t119 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1332 a_59578_n29970# frontAnalog_v0p0p1_6.x65.X frontAnalog_v0p0p1_6.RSfetsym_0.QN.t2 GND.t410 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.315 ps=2.72 w=1 l=0.15
X1333 a_53630_n68796# frontAnalog_v0p0p1_10.IB.t21 GND.t453 GND.t296 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1334 GND.t118 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t18 GND.t117 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1335 a_77605_n40069# I15.t7 GND.t1068 GND.t555 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X1336 VV14.t17 w_55000_n14350# error sky130_fd_pr__cap_var_lvt w=2 l=0.18
X1337 GND.t116 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t17 GND.t115 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1338 frontAnalog_v0p0p1_9.RSfetsym_0.x1.Y frontAnalog_v0p0p1_9.x63.X GND.t1400 GND.t1398 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1339 a_16719_n13117.t13 a_16599_n13205.t14 a_16541_n13117.t9 GND.t429 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1340 a_77637_n40777# VDD.t787 VDD.t789 VDD.t788 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X1341 VDD.t1328 R0.t10 frontAnalog_v0p0p1_15.RSfetsym_0.x1.Y VDD.t1006 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1342 VDD.t697 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t86 VDD.t696 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1343 GND.t585 frontAnalog_v0p0p1_6.x63.X frontAnalog_v0p0p1_6.RSfetsym_0.x1.Y GND.t584 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1344 16to4_PriorityEncoder_v0p0p1_0.x43.A 16to4_PriorityEncoder_v0p0p1_0.x42.A GND.t1350 GND.t1349 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1345 GND.t1521 frontAnalog_v0p0p1_12.RSfetsym_0.QN.t6 a_59577_n73683# GND.t1520 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1346 OUT2.t27 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND.t940 GND.t939 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1347 GND.t1153 I0.t8 a_59578_n83970# GND.t1152 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1348 a_78147_n49349# 16to4_PriorityEncoder_v0p0p1_0.x3.x22.A a_78065_n49349# VDD.t470 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X1349 GND.t1556 16to4_PriorityEncoder_v0p0p1_0.x3.x19.D a_77881_n52567# GND.t67 sky130_fd_pr__nfet_01v8 ad=0.196 pd=1.33 as=0.0693 ps=0.75 w=0.42 l=0.15
X1350 OUT1.t85 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD.t695 VDD.t694 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1351 16to4_PriorityEncoder_v0p0p1_0.x5.x19.X a_77605_n44779# GND.t461 GND.t460 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.196 ps=1.33 w=0.65 l=0.15
X1352 GND.t938 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t26 GND.t937 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1353 a_82906_n43855# 16to4_PriorityEncoder_v0p0p1_0.x3.A2 GND.t865 GND.t864 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1354 VDD.t875 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t82 VDD.t874 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1355 a_78313_n39305# 16to4_PriorityEncoder_v0p0p1_0.x5.x1.X a_78241_n39305# VDD.t1005 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X1356 VV8.t14 VV7.t13 GND.t401 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1357 VV10.t13 VV9.t14 GND.t250 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1358 I13.t3 frontAnalog_v0p0p1_3.x63.X VDD.t1449 VDD.t1446 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.25
X1359 a_53630_n25596# frontAnalog_v0p0p1_10.IB.t22 GND.t454 GND.t296 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1360 a_16719_n13117.t12 a_16599_n13205.t15 a_16541_n13117.t8 GND.t430 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1361 VDD.t1325 frontAnalog_v0p0p1_4.x63.A.t7 frontAnalog_v0p0p1_4.x65.A.t3 VDD.t278 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1362 frontAnalog_v0p0p1_11.RSfetsym_0.x1.Y frontAnalog_v0p0p1_11.x63.X VDD.t9 VDD.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1363 OUT0.t83 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD.t126 VDD.t125 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1364 GND.t544 I12.t10 a_59578_n19170# GND.t543 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1365 VV3.t4 VV2.t4 GND.t481 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1366 VDD.t124 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t82 VDD.t123 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1367 VV13.t13 VV12.t13 GND.t250 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1368 OUT0.t16 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND.t114 GND.t113 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1369 GND.t112 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t15 GND.t111 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1370 VV5.t12 VV4.t9 GND.t80 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1371 VDD.t1041 S1.t8 frontAnalog_v0p0p1_14.RSfetsym_0.x2.Y VDD.t420 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1372 a_78527_n51085# 16to4_PriorityEncoder_v0p0p1_0.x3.x15.X a_78431_n51085# VDD.t605 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X1373 GND.t1136 16to4_PriorityEncoder_v0p0p1_0.x35.A 16to4_PriorityEncoder_v0p0p1_0.x36.A GND.t1135 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1374 VDD.t873 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t81 VDD.t872 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1375 VDD.t122 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t81 VDD.t121 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1376 16to4_PriorityEncoder_v0p0p1_0.x3.A0 a_78525_n53555# GND.t444 GND.t443 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.102 ps=0.99 w=0.65 l=0.15
X1377 GND.t419 frontAnalog_v0p0p1_6.RSfetsym_0.QN.t6 a_59577_n30483# GND.t418 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1378 frontAnalog_v0p0p1_10.RSfetsym_0.QN.t0 I5.t12 VDD.t1318 VDD.t1317 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.3
X1379 frontAnalog_v0p0p1_7.x65.X a_57123_n34959# GND.t421 GND.t420 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1380 GND.t266 I8.t7 a_59578_n40770# GND.t265 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1381 frontAnalog_v0p0p1_10.IB.t0 a_16719_n13117.t24 VDD.t1037 VDD.t1036 sky130_fd_pr__pfet_01v8_lvt ad=5.51 pd=38.6 as=5.51 ps=38.6 w=19 l=1
X1382 a_77687_n39305# I11.t10 a_77605_n39305# VDD.t428 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X1383 VDD.t693 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t84 VDD.t692 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1384 OUT1.t83 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD.t691 VDD.t690 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1385 OUT2.t25 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND.t936 GND.t935 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1386 GND.t934 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t24 GND.t933 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1387 16to4_PriorityEncoder_v0p0p1_0.x3.x14.A a_77637_n48817# VDD.t1442 VDD.t1441 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.167 ps=1.39 w=1 l=0.15
X1388 a_77605_n48109# I7.t7 GND.t264 GND.t263 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X1389 VDD.t392 frontAnalog_v0p0p1_8.x65.A.t4 a_57123_n45759# VDD.t391 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1390 VDD.t1298 frontAnalog_v0p0p1_7.x65.X frontAnalog_v0p0p1_7.RSfetsym_0.x2.Y VDD.t1297 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1391 16to4_PriorityEncoder_v0p0p1_0.x5.x16.C I13.t11 VDD.t1361 VDD.t1360 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1392 VV2.t11 VV1.t10 GND.t78 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1393 VFS.t0 VV16.t0 GND.t209 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1394 frontAnalog_v0p0p1_3.RSfetsym_0.QN.t0 I13.t12 VDD.t1362 VDD.t1331 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.3
X1395 OUT0.t80 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD.t120 VDD.t119 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1396 VDD.t118 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t79 VDD.t117 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1397 GND.t697 VDD.t1508 a_78735_n39527# GND.t696 sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X1398 VDD.t1039 a_16719_n13117.t25 a_16599_n13205.t1 VDD.t1038 sky130_fd_pr__pfet_01v8_lvt ad=5.51 pd=38.6 as=5.51 ps=38.6 w=19 l=1
X1399 OUT1.t82 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD.t689 VDD.t688 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1400 VV4.t10 VV3.t11 GND.t12 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1401 16to4_PriorityEncoder_v0p0p1_0.x3.x19.X a_77605_n52819# GND.t706 GND.t705 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.196 ps=1.33 w=0.65 l=0.15
X1402 16to4_PriorityEncoder_v0p0p1_0.x36.A 16to4_PriorityEncoder_v0p0p1_0.x35.A VDD.t1079 VDD.t1078 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1403 VDD.t226 16to4_PriorityEncoder_v0p0p1_0.x29.A 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD.t225 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1404 16to4_PriorityEncoder_v0p0p1_0.x3.x21.X a_78097_n53777# GND.t366 GND.t365 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.112 ps=1.04 w=0.65 l=0.15
X1405 w_55000_n62950# VIN.t25 a_53630_n63396# GND.t315 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1406 frontAnalog_v0p0p1_15.RSfetsym_0.x2.Y S0.t7 GND.t1320 GND.t1319 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1407 a_78313_n47345# 16to4_PriorityEncoder_v0p0p1_0.x3.x1.X a_78241_n47345# VDD.t1110 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X1408 16to4_PriorityEncoder_v0p0p1_0.x36.Y 16to4_PriorityEncoder_v0p0p1_0.x36.A GND.t47 GND.t46 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1409 VDD.t1029 frontAnalog_v0p0p1_2.x65.X frontAnalog_v0p0p1_2.RSfetsym_0.x2.Y VDD.t1028 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1410 frontAnalog_v0p0p1_13.RSfetsym_0.x1.Y frontAnalog_v0p0p1_13.x63.X VDD.t1054 VDD.t1050 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1411 16to4_PriorityEncoder_v0p0p1_0.x3.x19.C I4.t11 VDD.t1344 VDD.t1343 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1412 frontAnalog_v0p0p1_4.RSfetsym_0.QN.t3 frontAnalog_v0p0p1_4.x65.X VDD.t1422 VDD.t1417 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.25
X1413 frontAnalog_v0p0p1_3.RSfetsym_0.x1.Y frontAnalog_v0p0p1_3.x63.X GND.t1510 GND.t1508 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1414 VFS.t5 VV16.t12 GND.t79 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1415 OUT0.t14 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND.t110 GND.t109 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1416 a_77687_n47345# I3.t11 a_77605_n47345# VDD.t782 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X1417 VDD.t871 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t80 VDD.t870 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1418 VDD.t687 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t81 VDD.t686 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1419 frontAnalog_v0p0p1_1.RSfetsym_0.x2.Y frontAnalog_v0p0p1_1.x65.X GND.t516 GND.t515 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1420 frontAnalog_v0p0p1_5.RSfetsym_0.x1.Y frontAnalog_v0p0p1_5.x63.X VDD.t980 VDD.t976 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1421 a_59577_n84483# R0.t11 I0.t3 GND.t1393 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1422 a_77775_n44779# I11.t11 a_77687_n44779# GND.t247 sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
X1423 OUT2.t23 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND.t932 GND.t931 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1424 I4.t4 frontAnalog_v0p0p1_11.RSfetsym_0.x2.Y GND.t1545 GND.t1158 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.25
X1425 16to4_PriorityEncoder_v0p0p1_0.x29.Y 16to4_PriorityEncoder_v0p0p1_0.x29.A VDD.t224 VDD.t223 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1426 frontAnalog_v0p0p1_11.x63.A.t1 frontAnalog_v0p0p1_11.x65.A.t5 VDD.t1365 VDD.t1021 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1427 VDD.t1012 frontAnalog_v0p0p1_0.x65.A.t5 a_57123_n7959# VDD.t1011 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1428 GND.t45 16to4_PriorityEncoder_v0p0p1_0.x36.A 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND.t44 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1429 GND.t382 16to4_PriorityEncoder_v0p0p1_0.x3.EI a_78735_n47567# GND.t381 sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X1430 VDD.t529 CLK.t60 w_55000_n78528# GND.t573 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1431 OUT0.t78 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD.t116 VDD.t115 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1432 I5.t0 frontAnalog_v0p0p1_10.x63.X VDD.t486 VDD.t485 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.25
X1433 GND.t1051 16to4_PriorityEncoder_v0p0p1_0.x28.A 16to4_PriorityEncoder_v0p0p1_0.x29.A GND.t1050 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1434 a_77605_n44779# 16to4_PriorityEncoder_v0p0p1_0.x5.x19.C VDD.t630 VDD.t629 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X1435 VDD.t373 frontAnalog_v0p0p1_12.x65.X frontAnalog_v0p0p1_12.RSfetsym_0.x2.Y VDD.t372 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1436 GND.t380 16to4_PriorityEncoder_v0p0p1_0.x3.EI a_77759_n53805# GND.t379 sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X1437 a_59577_n41283# frontAnalog_v0p0p1_1.x63.X I8.t2 GND.t1529 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1438 VV10.t7 VV9.t7 GND.t78 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1439 a_59578_n51570# frontAnalog_v0p0p1_9.x65.X frontAnalog_v0p0p1_9.RSfetsym_0.QN.t1 GND.t1435 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.315 ps=2.72 w=1 l=0.15
X1440 VDD.t1053 frontAnalog_v0p0p1_13.x63.X I3.t1 VDD.t1052 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.25
X1441 VDD.t530 CLK.t61 w_55000_n79150# GND.t562 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1442 frontAnalog_v0p0p1_4.x63.A.t2 frontAnalog_v0p0p1_4.x65.A.t6 VDD.t1329 VDD.t1023 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1443 I12.t0 frontAnalog_v0p0p1_4.RSfetsym_0.x2.Y GND.t612 GND.t10 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.25
X1444 w_55000_n67728# CLK.t62 frontAnalog_v0p0p1_13.x65.A.t0 VDD.t531 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1445 VDD.t413 frontAnalog_v0p0p1_15.x63.A.t7 frontAnalog_v0p0p1_15.x65.A.t2 VDD.t265 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1446 OUT1.t18 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND.t756 GND.t755 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1447 S1.t0 a_57123_n78159# GND.t1098 GND.t1097 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1448 VV13.t10 VV12.t11 GND.t78 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1449 frontAnalog_v0p0p1_5.x65.X a_57123_n24159# VDD.t1480 VDD.t1479 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1450 frontAnalog_v0p0p1_4.x63.X a_57123_n20279# GND.t77 GND.t76 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1451 GND.t930 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t22 GND.t929 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1452 frontAnalog_v0p0p1_3.x63.A.t3 CLK.t63 w_55000_n14350# VDD.t521 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1453 VDD.t522 CLK.t64 w_55000_n35328# GND.t568 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1454 GND.t490 16to4_PriorityEncoder_v0p0p1_0.x5.x19.X a_78525_n45515# GND.t489 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X1455 frontAnalog_v0p0p1_7.RSfetsym_0.QN.t0 frontAnalog_v0p0p1_7.RSfetsym_0.x1.Y GND.t636 GND.t635 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.25
X1456 VDD.t386 frontAnalog_v0p0p1_6.x65.X frontAnalog_v0p0p1_6.RSfetsym_0.x2.Y VDD.t385 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1457 frontAnalog_v0p0p1_8.RSfetsym_0.x2.Y frontAnalog_v0p0p1_8.x65.X GND.t1328 GND.t1327 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1458 VDD.t254 frontAnalog_v0p0p1_9.x63.A.t5 a_57123_n52679# VDD.t253 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1459 VDD.t979 frontAnalog_v0p0p1_5.x63.X I11.t2 VDD.t978 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.25
X1460 VDD.t523 CLK.t65 w_55000_n35950# GND.t564 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1461 OUT1.t80 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD.t685 VDD.t684 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1462 16to4_PriorityEncoder_v0p0p1_0.x29.A 16to4_PriorityEncoder_v0p0p1_0.x28.A VDD.t989 VDD.t988 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1463 w_55000_n24528# CLK.t66 frontAnalog_v0p0p1_5.x65.A.t0 VDD.t524 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1464 GND.t1218 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t16 GND.t1217 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1465 a_16719_n13117.t1 a_16719_n13117.t0 VDD.t1027 VDD.t1026 sky130_fd_pr__pfet_01v8_lvt ad=5.51 pd=38.6 as=5.51 ps=38.6 w=19 l=1
X1466 a_53630_n3996# frontAnalog_v0p0p1_10.IB.t23 GND.t653 GND.t293 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1467 GND.t928 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t21 GND.t927 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1468 a_55268_n74136# CLK.t67 GND.t570 GND.t569 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1469 16to4_PriorityEncoder_v0p0p1_0.x43.Y 16to4_PriorityEncoder_v0p0p1_0.x43.A VDD.t297 VDD.t296 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1470 frontAnalog_v0p0p1_8.x65.A.t0 frontAnalog_v0p0p1_8.x63.A.t6 a_55268_n47136# GND.t641 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1471 VDD.t510 I14.t11 a_77637_n42017# VDD.t509 sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X1472 16to4_PriorityEncoder_v0p0p1_0.x5.EO a_78159_n39549# GND.t627 GND.t626 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.102 ps=0.99 w=0.65 l=0.15
X1473 VDD.t1051 frontAnalog_v0p0p1_13.x63.X frontAnalog_v0p0p1_13.RSfetsym_0.x1.Y VDD.t1050 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1474 a_77605_n52819# 16to4_PriorityEncoder_v0p0p1_0.x3.x19.C VDD.t72 VDD.t71 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X1475 GND.t1509 frontAnalog_v0p0p1_3.x63.X frontAnalog_v0p0p1_3.RSfetsym_0.x1.Y GND.t1508 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1476 frontAnalog_v0p0p1_10.RSfetsym_0.x2.Y frontAnalog_v0p0p1_10.x65.X VDD.t1113 VDD.t1111 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1477 VFS.t2 VV16.t5 GND.t589 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1478 frontAnalog_v0p0p1_10.RSfetsym_0.x1.Y frontAnalog_v0p0p1_10.x63.X GND.t527 GND.t525 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1479 a_53630_n52596# VV7.t17 w_55000_n51528# GND.t287 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1480 a_16719_n13117.t11 a_16599_n13205.t16 a_16541_n13117.t21 GND.t431 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1481 VV3.t10 VV2.t9 GND.t537 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1482 VDD.t1145 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t74 VDD.t1144 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1483 VV4.t12 VV3.t13 GND.t417 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1484 GND.t72 frontAnalog_v0p0p1_0.x63.X frontAnalog_v0p0p1_0.RSfetsym_0.x1.Y GND.t71 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1485 VV8.t1 VV7.t1 GND.t80 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1486 a_55268_n30936# CLK.t68 GND.t572 GND.t571 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1487 GND.t279 frontAnalog_v0p0p1_11.x63.A.t7 a_57123_n63479# GND.t278 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X1488 frontAnalog_v0p0p1_15.RSfetsym_0.QN.t3 S0.t8 VDD.t1252 VDD.t0 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.25
X1489 GND.t926 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t20 GND.t925 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1490 OUT3.t73 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD.t1143 VDD.t1142 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1491 OUT1.t17 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND.t754 GND.t753 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1492 OUT2.t19 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND.t924 GND.t923 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1493 VDD.t977 frontAnalog_v0p0p1_5.x63.X frontAnalog_v0p0p1_5.RSfetsym_0.x1.Y VDD.t976 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1494 GND.t1123 16to4_PriorityEncoder_v0p0p1_0.x3.x19.X a_78525_n53555# GND.t1122 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X1495 frontAnalog_v0p0p1_3.RSfetsym_0.x2.Y frontAnalog_v0p0p1_3.x65.X VDD.t830 VDD.t828 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1496 16to4_PriorityEncoder_v0p0p1_0.x5.EO a_78159_n39549# VDD.t579 VDD.t578 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.148 ps=1.34 w=1 l=0.15
X1497 GND.t1480 frontAnalog_v0p0p1_4.x65.X frontAnalog_v0p0p1_4.RSfetsym_0.x2.Y GND.t1479 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1498 a_78159_n39549# 16to4_PriorityEncoder_v0p0p1_0.x5.x1.X GND.t1064 GND.t1063 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1499 OUT3.t72 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD.t1141 VDD.t1140 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1500 a_53630_n79596# frontAnalog_v0p0p1_10.IB.t24 GND.t654 GND.t296 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1501 frontAnalog_v0p0p1_1.RSfetsym_0.QN.t3 frontAnalog_v0p0p1_1.x65.X VDD.t477 VDD.t476 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.25
X1502 VDD.t384 frontAnalog_v0p0p1_6.x65.X frontAnalog_v0p0p1_6.RSfetsym_0.QN.t0 VDD.t383 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.25
X1503 VDD.t222 16to4_PriorityEncoder_v0p0p1_0.x29.A 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD.t221 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1504 OUT3.t15 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND.t1216 GND.t1215 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1505 VV6.t5 VV5.t7 GND.t209 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1506 16to4_PriorityEncoder_v0p0p1_0.x36.Y 16to4_PriorityEncoder_v0p0p1_0.x36.A GND.t43 GND.t42 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1507 16to4_PriorityEncoder_v0p0p1_0.x5.x22.A a_77639_n42341# GND.t614 GND.t613 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.112 ps=1.04 w=0.65 l=0.15
X1508 OUT1.t16 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND.t752 GND.t751 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1509 GND.t370 16to4_PriorityEncoder_v0p0p1_0.x21.A 16to4_PriorityEncoder_v0p0p1_0.x22.A GND.t369 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1510 VDD.t1367 frontAnalog_v0p0p1_9.x65.X frontAnalog_v0p0p1_9.RSfetsym_0.QN.t2 VDD.t1366 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.25
X1511 16to4_PriorityEncoder_v0p0p1_0.x3.EO a_78159_n47589# GND.t680 GND.t679 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.102 ps=0.99 w=0.65 l=0.15
X1512 OUT2.t79 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD.t869 VDD.t868 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1513 VV1.t5 VL.t3 GND.t250 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1514 a_77687_n43295# I10.t10 a_77605_n43295# GND.t687 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.109 ps=1.36 w=0.42 l=0.15
X1515 VDD.t867 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t78 VDD.t866 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1516 frontAnalog_v0p0p1_11.x65.A.t2 CLK.t69 frontAnalog_v0p0p1_11.x63.A.t3 VDD.t525 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1517 frontAnalog_v0p0p1_13.x65.X a_57123_n67359# VDD.t459 VDD.t458 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1518 a_53630_n36396# frontAnalog_v0p0p1_10.IB.t25 GND.t655 GND.t296 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1519 OUT0.t13 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND.t108 GND.t107 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1520 OUT3.t71 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD.t1139 VDD.t1138 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1521 frontAnalog_v0p0p1_10.x63.A.t3 CLK.t70 w_55000_n57550# VDD.t266 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1522 GND.t1399 frontAnalog_v0p0p1_9.x63.X frontAnalog_v0p0p1_9.RSfetsym_0.x1.Y GND.t1398 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1523 16to4_PriorityEncoder_v0p0p1_0.x29.Y 16to4_PriorityEncoder_v0p0p1_0.x29.A GND.t213 GND.t212 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1524 VV9.t4 VV8.t4 GND.t250 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1525 frontAnalog_v0p0p1_14.RSfetsym_0.QN.t2 frontAnalog_v0p0p1_14.RSfetsym_0.x1.Y GND.t1045 GND.t1044 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.25
X1526 VV6.t8 VV5.t8 GND.t79 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1527 OUT3.t14 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND.t1214 GND.t1213 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1528 VDD.t1137 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t70 VDD.t1136 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1529 VV16.t8 VV15.t8 GND.t299 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1530 R0.t0 a_57123_n85079# GND.t524 GND.t523 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1531 GND.t1326 frontAnalog_v0p0p1_8.x65.X frontAnalog_v0p0p1_8.RSfetsym_0.x2.Y GND.t1325 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1532 VV7.t3 VV6.t4 GND.t244 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1533 GND.t1212 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t13 GND.t1211 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1534 frontAnalog_v0p0p1_4.RSfetsym_0.x2.Y frontAnalog_v0p0p1_4.x65.X VDD.t1421 VDD.t1419 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1535 GND.t441 frontAnalog_v0p0p1_11.x65.A.t6 a_57123_n61959# GND.t278 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X1536 VDD.t340 16to4_PriorityEncoder_v0p0p1_0.x21.A 16to4_PriorityEncoder_v0p0p1_0.x22.A VDD.t339 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1537 a_16719_n13117.t10 a_16599_n13205.t17 a_16541_n13117.t20 GND.t432 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1538 16to4_PriorityEncoder_v0p0p1_0.x3.EO a_78159_n47589# VDD.t622 VDD.t621 sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.148 ps=1.34 w=1 l=0.15
X1539 a_78159_n47589# 16to4_PriorityEncoder_v0p0p1_0.x3.x1.X GND.t1172 GND.t1171 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1540 VDD.t8 frontAnalog_v0p0p1_11.x63.X frontAnalog_v0p0p1_11.RSfetsym_0.x1.Y VDD.t7 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1541 frontAnalog_v0p0p1_1.RSfetsym_0.x2.Y frontAnalog_v0p0p1_1.x65.X VDD.t475 VDD.t473 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1542 OUT2.t18 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND.t922 GND.t921 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1543 frontAnalog_v0p0p1_5.RSfetsym_0.x2.Y frontAnalog_v0p0p1_5.x65.X GND.t465 GND.t464 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1544 frontAnalog_v0p0p1_14.RSfetsym_0.x1.Y R1.t11 GND.t607 GND.t606 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1545 OUT1.t15 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND.t750 GND.t749 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1546 a_78525_n45515# 16to4_PriorityEncoder_v0p0p1_0.x5.x20.X GND.t1507 GND.t1506 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X1547 OUT0.t77 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD.t114 VDD.t113 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1548 16to4_PriorityEncoder_v0p0p1_0.x5.x19.D I14.t12 VDD.t1312 VDD.t1311 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1549 16to4_PriorityEncoder_v0p0p1_0.x35.A 16to4_PriorityEncoder_v0p0p1_0.x34.A GND.t1544 GND.t1543 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1550 16to4_PriorityEncoder_v0p0p1_0.x3.x22.A a_77639_n50381# GND.t483 GND.t482 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.112 ps=1.04 w=0.65 l=0.15
X1551 frontAnalog_v0p0p1_1.x63.X a_57123_n41879# GND.t567 GND.t64 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1552 GND.t526 frontAnalog_v0p0p1_10.x63.X frontAnalog_v0p0p1_10.RSfetsym_0.x1.Y GND.t525 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1553 VV5.t17 w_55000_n62950# error sky130_fd_pr__cap_var_lvt w=2 l=0.18
X1554 OUT1.t14 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND.t748 GND.t747 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1555 GND.t746 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t13 GND.t745 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1556 GND.t211 16to4_PriorityEncoder_v0p0p1_0.x29.A 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND.t210 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1557 a_77605_n44527# 16to4_PriorityEncoder_v0p0p1_0.x5.x18.C VDD.t472 VDD.t285 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X1558 VDD.t865 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t77 VDD.t864 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1559 a_77881_n43545# 16to4_PriorityEncoder_v0p0p1_0.x5.x16.C a_77775_n43545# GND.t686 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X1560 GND.t698 VDD.t1509 a_77881_n43295# GND.t687 sky130_fd_pr__nfet_01v8 ad=0.196 pd=1.33 as=0.0693 ps=0.75 w=0.42 l=0.15
X1561 a_77725_n42341# VDD.t1510 a_77639_n42341# GND.t699 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X1562 OUT3.t12 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND.t1210 GND.t1209 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1563 frontAnalog_v0p0p1_7.RSfetsym_0.x1.Y frontAnalog_v0p0p1_7.x63.X GND.t631 GND.t629 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1564 OUT0.t12 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND.t106 GND.t105 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1565 16to4_PriorityEncoder_v0p0p1_0.x5.x20.X a_77605_n45765# GND.t1515 GND.t1514 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.132 ps=1.14 w=0.65 l=0.15
X1566 VDD.t288 16to4_PriorityEncoder_v0p0p1_0.x5.x22.A a_78775_n45515# VDD.t287 sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X1567 GND.t1208 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t11 GND.t1207 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1568 GND.t496 frontAnalog_v0p0p1_10.RSfetsym_0.QN.t6 a_59577_n57483# GND.t495 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1569 GND.t854 I3.t12 a_59578_n67770# GND.t853 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1570 VDD.t863 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t76 VDD.t862 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1571 16to4_PriorityEncoder_v0p0p1_0.x43.Y 16to4_PriorityEncoder_v0p0p1_0.x43.A VDD.t295 VDD.t294 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1572 VDD.t683 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t79 VDD.t682 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1573 a_16719_n13117.t9 a_16599_n13205.t18 a_16541_n13117.t19 GND.t433 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1574 16to4_PriorityEncoder_v0p0p1_0.x43.Y 16to4_PriorityEncoder_v0p0p1_0.x43.A GND.t336 GND.t335 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1575 frontAnalog_v0p0p1_2.x63.X a_57123_n4079# VDD.t1499 VDD.t1498 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1576 GND.t744 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t12 GND.t743 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1577 GND.t1322 S0.t9 frontAnalog_v0p0p1_15.RSfetsym_0.x2.Y GND.t1321 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1578 16to4_PriorityEncoder_v0p0p1_0.x29.Y 16to4_PriorityEncoder_v0p0p1_0.x29.A VDD.t220 VDD.t219 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1579 frontAnalog_v0p0p1_8.RSfetsym_0.x1.Y frontAnalog_v0p0p1_8.x63.X VDD.t999 VDD.t997 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1580 VV15.t10 VV14.t9 GND.t12 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1581 a_53630_n30996# frontAnalog_v0p0p1_10.IB.t26 GND.t656 GND.t296 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1582 a_78241_n39305# 16to4_PriorityEncoder_v0p0p1_0.x5.x2.X a_78159_n39549# VDD.t577 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X1583 OUT0.t11 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND.t104 GND.t103 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1584 GND.t638 frontAnalog_v0p0p1_2.RSfetsym_0.QN.t5 a_59577_n3483# GND.t637 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1585 a_78525_n53555# 16to4_PriorityEncoder_v0p0p1_0.x3.x20.X GND.t604 GND.t603 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X1586 OUT0.t76 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD.t112 VDD.t111 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1587 GND.t742 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t11 GND.t741 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1588 16to4_PriorityEncoder_v0p0p1_0.x5.x20.X a_77605_n45765# VDD.t1453 VDD.t1452 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X1589 GND.t1397 frontAnalog_v0p0p1_3.RSfetsym_0.QN.t6 a_59577_n14283# GND.t1396 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1590 frontAnalog_v0p0p1_4.x65.X a_57123_n18759# GND.t621 GND.t76 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1591 GND.t249 I11.t12 a_59578_n24570# GND.t248 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1592 GND.t1206 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t10 GND.t1205 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1593 VV7.t15 VV6.t15 GND.t401 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1594 a_77605_n40069# I13.t13 GND.t1099 GND.t555 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1595 a_16719_n13117.t8 a_16599_n13205.t19 a_16541_n13117.t18 GND.t1034 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1596 frontAnalog_v0p0p1_12.x63.X a_57123_n74279# VDD.t1501 VDD.t1500 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1597 VV6.t13 VV5.t15 GND.t589 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1598 VV1.t1 VL.t0 GND.t78 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1599 a_77881_n51585# 16to4_PriorityEncoder_v0p0p1_0.x3.x16.C a_77775_n51585# GND.t66 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X1600 16to4_PriorityEncoder_v0p0p1_0.x5.A2 a_78065_n41309# VDD.t1287 VDD.t649 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.148 ps=1.34 w=1 l=0.15
X1601 GND.t514 frontAnalog_v0p0p1_1.x65.X frontAnalog_v0p0p1_1.RSfetsym_0.x2.Y GND.t513 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1602 VIN.t26 w_55000_n62328# error sky130_fd_pr__cap_var_lvt w=2 l=0.18
X1603 OUT2.t75 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD.t861 VDD.t860 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1604 GND.t1524 16to4_PriorityEncoder_v0p0p1_0.x3.x17.A a_78349_n51085# GND.t505 sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X1605 VDD.t648 frontAnalog_v0p0p1_6.x65.A.t6 a_57123_n29559# VDD.t647 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1606 16to4_PriorityEncoder_v0p0p1_0.x22.Y 16to4_PriorityEncoder_v0p0p1_0.x22.A GND.t1447 GND.t1446 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1607 16to4_PriorityEncoder_v0p0p1_0.x3.x2.X a_77605_n48109# VDD.t612 VDD.t611 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.148 ps=1.34 w=1 l=0.15
X1608 GND.t920 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t17 GND.t919 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1609 a_77725_n50381# 16to4_PriorityEncoder_v0p0p1_0.x3.EI a_77639_n50381# GND.t378 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X1610 VDD.t1044 I13.t14 a_77637_n41087# VDD.t791 sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X1611 VDD.t1420 frontAnalog_v0p0p1_4.x65.X frontAnalog_v0p0p1_4.RSfetsym_0.x2.Y VDD.t1419 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1612 OUT1.t78 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD.t681 VDD.t680 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1613 VV9.t0 VV8.t0 GND.t78 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1614 VDD.t469 16to4_PriorityEncoder_v0p0p1_0.x3.x22.A a_78775_n53555# VDD.t468 sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X1615 OUT0.t75 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD.t110 VDD.t109 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1616 VDD.t292 frontAnalog_v0p0p1_9.x65.A.t6 a_57123_n51159# VDD.t291 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1617 GND.t642 frontAnalog_v0p0p1_8.x63.A.t7 a_57123_n47279# GND.t425 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X1618 VDD.t474 frontAnalog_v0p0p1_1.x65.X frontAnalog_v0p0p1_1.RSfetsym_0.x2.Y VDD.t473 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1619 frontAnalog_v0p0p1_0.RSfetsym_0.x2.Y frontAnalog_v0p0p1_0.x65.X VDD.t1268 VDD.t1266 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1620 frontAnalog_v0p0p1_6.x63.X a_57123_n31079# VDD.t542 VDD.t541 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1621 frontAnalog_v0p0p1_15.RSfetsym_0.x2.Y S0.t10 VDD.t1253 VDD.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1622 16to4_PriorityEncoder_v0p0p1_0.x42.A 16to4_PriorityEncoder_v0p0p1_0.x5.GS GND.t1542 GND.t1347 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1623 16to4_PriorityEncoder_v0p0p1_0.x29.A 16to4_PriorityEncoder_v0p0p1_0.x28.A GND.t1049 GND.t1048 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1624 w_55000_n46750# VIN.t27 a_53630_n47196# GND.t1107 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1625 frontAnalog_v0p0p1_13.RSfetsym_0.x2.Y frontAnalog_v0p0p1_13.x65.X GND.t1498 GND.t1497 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1626 OUT0.t10 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND.t102 GND.t101 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1627 16to4_PriorityEncoder_v0p0p1_0.x22.Y 16to4_PriorityEncoder_v0p0p1_0.x22.A VDD.t1388 VDD.t1387 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1628 a_78241_n47345# 16to4_PriorityEncoder_v0p0p1_0.x3.x2.X a_78159_n47589# VDD.t1345 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X1629 frontAnalog_v0p0p1_5.RSfetsym_0.QN.t3 frontAnalog_v0p0p1_5.x65.X VDD.t437 VDD.t436 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.25
X1630 frontAnalog_v0p0p1_11.x63.A.t0 frontAnalog_v0p0p1_11.x65.A.t7 a_55268_n63336# GND.t442 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1631 OUT0.t9 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND.t100 GND.t99 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1632 GND.t98 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t8 GND.t97 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1633 GND.t1445 16to4_PriorityEncoder_v0p0p1_0.x22.A 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND.t1444 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1634 16to4_PriorityEncoder_v0p0p1_0.x3.x20.X a_77605_n53805# VDD.t1104 VDD.t1103 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.142 ps=1.34 w=1 l=0.15
X1635 a_77783_n48109# I6.t12 a_77687_n48109# VDD.t1321 sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X1636 16to4_PriorityEncoder_v0p0p1_0.x1.A a_78349_n43045# GND.t538 GND.t406 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.102 ps=0.99 w=0.65 l=0.15
X1637 I4.t3 frontAnalog_v0p0p1_11.RSfetsym_0.QN.t5 VDD.t410 VDD.t409 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.3
X1638 a_77605_n48109# I5.t13 GND.t1383 GND.t263 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1639 GND.t740 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t10 GND.t739 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1640 GND.t1360 16to4_PriorityEncoder_v0p0p1_0.x5.x14.A a_78065_n41309# GND.t1359 sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X1641 VDD.t679 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t77 VDD.t678 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1642 OUT1.t76 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD.t677 VDD.t676 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1643 a_59577_n68283# frontAnalog_v0p0p1_13.x63.X I3.t0 GND.t1109 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1644 a_59578_n78570# S1.t9 frontAnalog_v0p0p1_14.RSfetsym_0.QN.t3 GND.t1489 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.315 ps=2.72 w=1 l=0.15
X1645 GND.t918 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t16 GND.t917 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1646 VDD.t675 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t75 VDD.t674 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1647 I7.t4 frontAnalog_v0p0p1_8.RSfetsym_0.x2.Y GND.t1476 GND.t1404 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.25
X1648 frontAnalog_v0p0p1_8.x63.A.t0 frontAnalog_v0p0p1_8.x65.A.t5 VDD.t394 VDD.t393 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1649 16to4_PriorityEncoder_v0p0p1_0.x5.x18.C I10.t11 VDD.t970 VDD.t969 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1650 OUT0.t74 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD.t108 VDD.t107 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1651 OUT2.t15 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND.t916 GND.t915 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1652 frontAnalog_v0p0p1_4.x63.A.t3 frontAnalog_v0p0p1_4.x65.A.t7 a_55268_n20136# GND.t1395 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1653 a_77759_n45765# 16to4_PriorityEncoder_v0p0p1_0.x5.x19.D a_77687_n45765# GND.t1546 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X1654 VDD.t1352 16to4_PriorityEncoder_v0p0p1_0.x5.A2 a_82988_n43855# VDD.t1351 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X1655 frontAnalog_v0p0p1_1.x63.A.t3 CLK.t71 w_55000_n41350# VDD.t514 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1656 OUT0.t73 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD.t106 VDD.t105 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1657 VDD.t104 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t72 VDD.t103 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1658 VDD.t1386 16to4_PriorityEncoder_v0p0p1_0.x22.A 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD.t1385 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1659 VDD.t1112 frontAnalog_v0p0p1_10.x65.X frontAnalog_v0p0p1_10.RSfetsym_0.x2.Y VDD.t1111 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1660 a_78649_n39527# 16to4_PriorityEncoder_v0p0p1_0.x5.EO VDD.t535 VDD.t534 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X1661 GND.t96 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t7 GND.t95 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1662 16to4_PriorityEncoder_v0p0p1_0.x1.A a_78349_n43045# VDD.t499 VDD.t498 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.148 ps=1.34 w=1 l=0.15
X1663 VDD.t818 frontAnalog_v0p0p1_14.x63.A.t7 a_57123_n79679# VDD.t817 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1664 a_78349_n43045# 16to4_PriorityEncoder_v0p0p1_0.x5.x22.A GND.t320 GND.t319 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1665 a_59577_n25083# frontAnalog_v0p0p1_5.x63.X I11.t1 GND.t1028 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1666 a_59578_n35370# frontAnalog_v0p0p1_7.x65.X frontAnalog_v0p0p1_7.RSfetsym_0.QN.t1 GND.t1369 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.315 ps=2.72 w=1 l=0.15
X1667 VDD.t515 CLK.t72 w_55000_n83928# GND.t562 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1668 I4.t1 frontAnalog_v0p0p1_11.x63.X VDD.t6 VDD.t5 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.25
X1669 a_53630_n74196# frontAnalog_v0p0p1_10.IB.t27 GND.t1083 GND.t296 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1670 a_78775_n45515# 16to4_PriorityEncoder_v0p0p1_0.x5.x21.X a_78703_n45515# VDD.t595 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X1671 VDD.t1069 frontAnalog_v0p0p1_13.x63.A.t7 frontAnalog_v0p0p1_13.x65.A.t2 VDD.t415 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1672 VDD.t673 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t74 VDD.t672 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1673 OUT1.t73 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD.t671 VDD.t670 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1674 GND.t94 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t6 GND.t93 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1675 OUT3.t9 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND.t1204 GND.t1203 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1676 OUT2.t14 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND.t914 GND.t913 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1677 VDD.t516 CLK.t73 w_55000_n19128# GND.t563 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1678 S0.t0 a_57123_n83559# GND.t690 GND.t523 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1679 frontAnalog_v0p0p1_4.RSfetsym_0.QN.t0 frontAnalog_v0p0p1_4.RSfetsym_0.x1.Y GND.t1354 GND.t547 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.25
X1680 16to4_PriorityEncoder_v0p0p1_0.x43.A 16to4_PriorityEncoder_v0p0p1_0.x42.A GND.t1348 GND.t1347 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1681 VDD.t829 frontAnalog_v0p0p1_3.x65.X frontAnalog_v0p0p1_3.RSfetsym_0.x2.Y VDD.t828 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1682 VV15.t1 VV14.t1 GND.t417 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1683 OUT3.t69 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD.t1135 VDD.t1134 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1684 VDD.t81 frontAnalog_v0p0p1_0.x63.X I14.t1 VDD.t80 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.25
X1685 VDD.t1294 frontAnalog_v0p0p1_7.x63.A.t6 a_57123_n36479# VDD.t1293 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1686 a_53630_n79596# VV2.t17 w_55000_n78528# GND.t22 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1687 VDD.t517 CLK.t74 w_55000_n40728# GND.t564 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1688 I12.t2 frontAnalog_v0p0p1_4.x63.X VDD.t568 VDD.t567 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.25
X1689 VFS.t4 VV16.t9 GND.t257 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1690 VDD.t859 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t74 VDD.t858 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1691 VDD.t102 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t71 VDD.t101 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1692 a_77687_n53805# I5.t14 a_77605_n53805# GND.t1384 sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.109 ps=1.36 w=0.42 l=0.15
X1693 VDD.t369 frontAnalog_v0p0p1_5.x63.A.t7 frontAnalog_v0p0p1_5.x65.A.t2 VDD.t368 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1694 VV4.t11 VV3.t12 GND.t299 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1695 frontAnalog_v0p0p1_9.RSfetsym_0.x2.Y frontAnalog_v0p0p1_9.x65.X GND.t1434 GND.t1433 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1696 a_55268_n57936# CLK.t75 GND.t566 GND.t565 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1697 VDD.t1254 S0.t11 frontAnalog_v0p0p1_15.RSfetsym_0.x2.Y VDD.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1698 VDD.t518 CLK.t76 w_55000_n41350# GND.t447 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1699 frontAnalog_v0p0p1_6.x65.A.t0 frontAnalog_v0p0p1_6.x63.A.t7 a_55268_n30936# GND.t1519 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1700 frontAnalog_v0p0p1_11.RSfetsym_0.QN.t4 I4.t12 VDD.t1255 VDD.t409 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.3
X1701 VDD.t100 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t70 VDD.t99 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1702 GND.t41 16to4_PriorityEncoder_v0p0p1_0.x36.A 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND.t40 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1703 frontAnalog_v0p0p1_1.x65.X a_57123_n40359# GND.t65 GND.t64 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1704 VDD.t501 I12.t11 a_77637_n40777# VDD.t500 sky130_fd_pr__pfet_01v8_hvt ad=0.167 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X1705 16to4_PriorityEncoder_v0p0p1_0.x22.A 16to4_PriorityEncoder_v0p0p1_0.x21.A GND.t368 GND.t367 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1706 a_78649_n47567# 16to4_PriorityEncoder_v0p0p1_0.x3.EO VDD.t614 VDD.t613 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X1707 a_53630_n36396# VV10.t17 w_55000_n35328# GND.t281 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1708 16to4_PriorityEncoder_v0p0p1_0.x3.A1 a_78349_n51085# VDD.t1455 VDD.t1454 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.148 ps=1.34 w=1 l=0.15
X1709 GND.t1346 16to4_PriorityEncoder_v0p0p1_0.x42.A 16to4_PriorityEncoder_v0p0p1_0.x43.A GND.t1345 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1710 OUT2.t13 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND.t912 GND.t911 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1711 16to4_PriorityEncoder_v0p0p1_0.x3.x22.A a_77639_n50381# VDD.t450 VDD.t449 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.167 ps=1.39 w=1 l=0.15
X1712 a_78775_n53555# 16to4_PriorityEncoder_v0p0p1_0.x3.x21.X a_78703_n53555# VDD.t598 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X1713 frontAnalog_v0p0p1_11.RSfetsym_0.x2.Y frontAnalog_v0p0p1_11.x65.X VDD.t29 VDD.t27 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1714 frontAnalog_v0p0p1_2.RSfetsym_0.x1.Y frontAnalog_v0p0p1_2.x63.X VDD.t445 VDD.t443 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1715 VV11.t3 VV10.t2 GND.t12 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1716 a_55268_n14736# CLK.t77 GND.t560 GND.t559 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1717 frontAnalog_v0p0p1_11.RSfetsym_0.x1.Y frontAnalog_v0p0p1_11.x63.X GND.t6 GND.t4 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1718 frontAnalog_v0p0p1_13.RSfetsym_0.QN.t3 frontAnalog_v0p0p1_13.x65.X VDD.t1437 VDD.t1436 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.25
X1719 OUT2.t12 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND.t910 GND.t909 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1720 VDD.t1133 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t68 VDD.t1132 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1721 OUT1.t72 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD.t669 VDD.t668 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1722 GND.t1202 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t8 GND.t1201 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1723 GND.t908 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t11 GND.t907 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1724 VDD.t1430 S1.t10 frontAnalog_v0p0p1_14.RSfetsym_0.QN.t4 VDD.t422 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.25
X1725 OUT3.t67 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD.t1131 VDD.t1130 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1726 GND.t92 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t5 GND.t91 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1727 a_77637_n49127# 16to4_PriorityEncoder_v0p0p1_0.x3.EI VDD.t349 VDD.t326 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X1728 frontAnalog_v0p0p1_0.x65.A.t1 CLK.t78 frontAnalog_v0p0p1_0.x63.A.t2 VDD.t511 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1729 VV7.t0 VV6.t0 GND.t80 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1730 VDD.t1129 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t66 VDD.t1128 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1731 16to4_PriorityEncoder_v0p0p1_0.x22.A 16to4_PriorityEncoder_v0p0p1_0.x21.A VDD.t338 VDD.t337 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1732 frontAnalog_v0p0p1_12.RSfetsym_0.x1.Y frontAnalog_v0p0p1_12.x63.X VDD.t23 VDD.t19 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1733 GND.t463 frontAnalog_v0p0p1_5.x65.X frontAnalog_v0p0p1_5.RSfetsym_0.x2.Y GND.t462 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1734 a_77687_n48109# I7.t8 a_77605_n48109# VDD.t257 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X1735 GND.t608 R1.t12 frontAnalog_v0p0p1_14.RSfetsym_0.x1.Y GND.t606 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1736 VIN.t28 w_55000_n46128# error sky130_fd_pr__cap_var_lvt w=2 l=0.18
X1737 GND.t906 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t10 GND.t905 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1738 OUT2.t73 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD.t857 VDD.t856 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1739 frontAnalog_v0p0p1_2.x65.X a_57123_n2559# VDD.t1089 VDD.t1088 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1740 a_16719_n13117.t7 a_16599_n13205.t20 a_16541_n13117.t17 GND.t1035 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1741 a_53630_n84996# frontAnalog_v0p0p1_10.IB.t28 GND.t1084 GND.t296 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1742 VDD.t1296 frontAnalog_v0p0p1_7.x65.X frontAnalog_v0p0p1_7.RSfetsym_0.QN.t2 VDD.t1295 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.25
X1743 a_16719_n13117.t6 a_16599_n13205.t21 a_16541_n13117.t16 GND.t1036 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1744 OUT1.t9 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND.t738 GND.t737 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1745 VDD.t855 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t72 VDD.t854 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1746 VDD.t98 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t69 VDD.t97 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1747 16to4_PriorityEncoder_v0p0p1_0.x3.x11.X a_77637_n49127# VDD.t973 VDD.t967 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.167 ps=1.39 w=1 l=0.15
X1748 frontAnalog_v0p0p1_6.RSfetsym_0.x1.Y frontAnalog_v0p0p1_6.x63.X VDD.t547 VDD.t543 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1749 GND.t736 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t8 GND.t735 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1750 frontAnalog_v0p0p1_8.x65.A.t2 CLK.t79 frontAnalog_v0p0p1_8.x63.A.t2 VDD.t512 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1751 a_77605_n43545# 16to4_PriorityEncoder_v0p0p1_0.x5.x16.C VDD.t1456 VDD.t426 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X1752 frontAnalog_v0p0p1_3.x63.X a_57123_n14879# VDD.t1285 VDD.t1284 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1753 frontAnalog_v0p0p1_13.RSfetsym_0.x2.Y frontAnalog_v0p0p1_13.x65.X VDD.t1435 VDD.t1433 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1754 frontAnalog_v0p0p1_0.RSfetsym_0.x1.Y frontAnalog_v0p0p1_0.x63.X VDD.t79 VDD.t77 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1755 a_53630_n20196# frontAnalog_v0p0p1_10.IB.t29 GND.t1085 GND.t296 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1756 w_55000_n30550# VIN.t29 a_53630_n30996# GND.t286 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1757 GND.t630 frontAnalog_v0p0p1_7.x63.X frontAnalog_v0p0p1_7.RSfetsym_0.x1.Y GND.t629 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1758 VDD.t1077 16to4_PriorityEncoder_v0p0p1_0.x35.A 16to4_PriorityEncoder_v0p0p1_0.x36.A VDD.t1076 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1759 GND.t1200 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t7 GND.t1199 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1760 GND.t1488 frontAnalog_v0p0p1_0.x63.A.t6 a_57123_n9479# GND.t251 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X1761 frontAnalog_v0p0p1_12.x65.X a_57123_n72759# VDD.t1475 VDD.t1474 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1762 frontAnalog_v0p0p1_13.x63.X a_57123_n68879# GND.t1165 GND.t499 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1763 GND.t39 16to4_PriorityEncoder_v0p0p1_0.x36.A 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND.t38 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1764 a_53630_n9396# VV15.t17 w_55000_n8328# GND.t282 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1765 a_53630_n41796# frontAnalog_v0p0p1_10.IB.t30 GND.t1086 GND.t296 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1766 frontAnalog_v0p0p1_11.x63.A.t2 CLK.t80 w_55000_n62950# VDD.t13 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1767 16to4_PriorityEncoder_v0p0p1_0.x5.x1.X a_77605_n39305# GND.t437 GND.t436 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.102 ps=0.99 w=0.65 l=0.15
X1768 VV14.t0 VV13.t1 GND.t12 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1769 GND.t426 frontAnalog_v0p0p1_8.x65.A.t6 a_57123_n45759# GND.t425 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X1770 VV5.t2 VV4.t1 GND.t250 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1771 OUT3.t6 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND.t1198 GND.t1197 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1772 frontAnalog_v0p0p1_15.RSfetsym_0.QN.t0 frontAnalog_v0p0p1_15.RSfetsym_0.x1.Y GND.t595 GND.t594 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.25
X1773 OUT2.t71 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD.t853 VDD.t852 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1774 VDD.t851 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t70 VDD.t850 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1775 GND.t1432 frontAnalog_v0p0p1_9.x65.X frontAnalog_v0p0p1_9.RSfetsym_0.x2.Y GND.t1431 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1776 GND.t334 16to4_PriorityEncoder_v0p0p1_0.x43.A 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND.t333 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1777 I7.t0 frontAnalog_v0p0p1_8.RSfetsym_0.QN.t6 VDD.t271 VDD.t270 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.3
X1778 frontAnalog_v0p0p1_5.RSfetsym_0.x2.Y frontAnalog_v0p0p1_5.x65.X VDD.t435 VDD.t433 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1779 VDD.t513 CLK.t81 w_55000_n84550# GND.t561 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1780 VDD.t998 frontAnalog_v0p0p1_8.x63.X frontAnalog_v0p0p1_8.RSfetsym_0.x1.Y VDD.t997 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1781 VDD.t22 frontAnalog_v0p0p1_12.x63.X I2.t1 VDD.t21 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.25
X1782 w_55000_n73128# CLK.t82 frontAnalog_v0p0p1_12.x65.A.t2 VDD.t401 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1783 frontAnalog_v0p0p1_5.x63.X a_57123_n25679# GND.t291 GND.t290 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1784 GND.t498 frontAnalog_v0p0p1_10.IB.t1 frontAnalog_v0p0p1_10.IB.t2 GND.t497 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1785 VV8.t17 w_55000_n46750# error sky130_fd_pr__cap_var_lvt w=2 l=0.18
X1786 GND.t904 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t9 GND.t903 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1787 frontAnalog_v0p0p1_1.RSfetsym_0.QN.t1 frontAnalog_v0p0p1_1.RSfetsym_0.x1.Y GND.t474 GND.t473 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.25
X1788 16to4_PriorityEncoder_v0p0p1_0.x5.x1.X a_77605_n39305# VDD.t404 VDD.t403 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.148 ps=1.34 w=1 l=0.15
X1789 OUT3.t5 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND.t1196 GND.t1195 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1790 16to4_PriorityEncoder_v0p0p1_0.x2.A a_78525_n45515# GND.t459 GND.t458 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.102 ps=0.99 w=0.65 l=0.15
X1791 16to4_PriorityEncoder_v0p0p1_0.x36.Y 16to4_PriorityEncoder_v0p0p1_0.x36.A GND.t37 GND.t36 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1792 VDD.t1127 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t65 VDD.t1126 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1793 GND.t5 frontAnalog_v0p0p1_11.x63.X frontAnalog_v0p0p1_11.RSfetsym_0.x1.Y GND.t4 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1794 GND.t734 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t7 GND.t733 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1795 16to4_PriorityEncoder_v0p0p1_0.x36.Y 16to4_PriorityEncoder_v0p0p1_0.x36.A VDD.t40 VDD.t39 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1796 VDD.t546 frontAnalog_v0p0p1_6.x63.X I10.t2 VDD.t545 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.25
X1797 a_77605_n51585# 16to4_PriorityEncoder_v0p0p1_0.x3.x16.C VDD.t1121 VDD.t73 sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0777 ps=0.79 w=0.42 l=0.15
X1798 w_55000_n29928# CLK.t83 frontAnalog_v0p0p1_6.x65.A.t3 VDD.t282 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1799 frontAnalog_v0p0p1_4.RSfetsym_0.x1.Y frontAnalog_v0p0p1_4.x63.X GND.t617 GND.t615 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1800 a_53630_n57996# frontAnalog_v0p0p1_10.IB.t31 GND.t849 GND.t296 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1801 a_55268_n79536# CLK.t84 GND.t534 GND.t533 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1802 frontAnalog_v0p0p1_9.x65.A.t0 frontAnalog_v0p0p1_9.x63.A.t6 a_55268_n52536# GND.t254 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1803 16to4_PriorityEncoder_v0p0p1_0.x43.Y 16to4_PriorityEncoder_v0p0p1_0.x43.A GND.t332 GND.t331 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1804 16to4_PriorityEncoder_v0p0p1_0.x3.x1.X a_77605_n47345# GND.t640 GND.t639 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.102 ps=0.99 w=0.65 l=0.15
X1805 VV11.t9 VV10.t10 GND.t417 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1806 VDD.t20 frontAnalog_v0p0p1_12.x63.X frontAnalog_v0p0p1_12.RSfetsym_0.x1.Y VDD.t19 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1807 GND.t732 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t6 GND.t731 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1808 frontAnalog_v0p0p1_0.RSfetsym_0.QN.t0 frontAnalog_v0p0p1_0.RSfetsym_0.x1.Y GND.t689 GND.t688 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.25
X1809 VDD.t1267 frontAnalog_v0p0p1_0.x65.X frontAnalog_v0p0p1_0.RSfetsym_0.x2.Y VDD.t1266 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1810 16to4_PriorityEncoder_v0p0p1_0.x3.x16.X a_77605_n51585# GND.t593 GND.t592 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.196 ps=1.33 w=0.65 l=0.15
X1811 GND.t1194 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t4 GND.t1193 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1812 GND.t252 frontAnalog_v0p0p1_0.x65.A.t6 a_57123_n7959# GND.t251 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X1813 GND.t1344 frontAnalog_v0p0p1_11.RSfetsym_0.QN.t6 a_59577_n62883# GND.t1343 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1814 GND.t1496 frontAnalog_v0p0p1_13.x65.X frontAnalog_v0p0p1_13.RSfetsym_0.x2.Y GND.t1495 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1815 VV6.t1 VV5.t0 GND.t257 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1816 16to4_PriorityEncoder_v0p0p1_0.x2.A a_78525_n45515# VDD.t430 VDD.t429 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.148 ps=1.34 w=1 l=0.15
X1817 OUT2.t69 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD.t849 VDD.t848 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1818 a_78525_n45515# 16to4_PriorityEncoder_v0p0p1_0.x5.x21.X GND.t648 GND.t647 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1819 VDD.t1429 frontAnalog_v0p0p1_0.x63.A.t7 frontAnalog_v0p0p1_0.x65.A.t3 VDD.t592 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1820 16to4_PriorityEncoder_v0p0p1_0.x5.x21.X a_78097_n45737# GND.t546 GND.t545 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.112 ps=1.04 w=0.65 l=0.15
X1821 VDD.t38 16to4_PriorityEncoder_v0p0p1_0.x36.A 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD.t37 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1822 a_53630_n14796# frontAnalog_v0p0p1_10.IB.t32 GND.t850 GND.t296 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1823 a_77637_n48817# 16to4_PriorityEncoder_v0p0p1_0.x3.EI VDD.t348 VDD.t347 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X1824 16to4_PriorityEncoder_v0p0p1_0.x5.x19.C I12.t12 VDD.t1375 VDD.t1374 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1825 frontAnalog_v0p0p1_9.RSfetsym_0.x1.Y frontAnalog_v0p0p1_9.x63.X VDD.t1334 VDD.t1333 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1826 VDD.t1100 frontAnalog_v0p0p1_14.x65.A.t7 a_57123_n78159# VDD.t1099 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1827 VDD.t987 16to4_PriorityEncoder_v0p0p1_0.x28.A 16to4_PriorityEncoder_v0p0p1_0.x29.A VDD.t986 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1828 VDD.t544 frontAnalog_v0p0p1_6.x63.X frontAnalog_v0p0p1_6.RSfetsym_0.x1.Y VDD.t543 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1829 OUT0.t4 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND.t90 GND.t89 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1830 OUT2.t8 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND.t902 GND.t901 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1831 I15.t4 frontAnalog_v0p0p1_2.RSfetsym_0.QN.t6 VDD.t1481 VDD.t1014 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.3
X1832 VDD.t1434 frontAnalog_v0p0p1_13.x65.X frontAnalog_v0p0p1_13.RSfetsym_0.x2.Y VDD.t1433 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1833 VDD.t78 frontAnalog_v0p0p1_0.x63.X frontAnalog_v0p0p1_0.RSfetsym_0.x1.Y VDD.t77 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1834 frontAnalog_v0p0p1_10.x63.X a_57123_n58079# VDD.t1049 VDD.t1048 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1835 16to4_PriorityEncoder_v0p0p1_0.x3.x1.X a_77605_n47345# VDD.t589 VDD.t588 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.148 ps=1.34 w=1 l=0.15
X1836 GND.t1192 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t3 GND.t1191 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1837 GND.t88 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t3 GND.t87 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1838 OUT1.t5 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND.t730 GND.t729 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1839 a_77775_n43545# 16to4_PriorityEncoder_v0p0p1_0.x5.x19.C a_77687_n43545# GND.t686 sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
X1840 16to4_PriorityEncoder_v0p0p1_0.x43.A 16to4_PriorityEncoder_v0p0p1_0.x42.A VDD.t1273 VDD.t1272 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1841 OUT1.t71 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD.t667 VDD.t666 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1842 frontAnalog_v0p0p1_2.RSfetsym_0.x2.Y frontAnalog_v0p0p1_2.x65.X GND.t1077 GND.t1076 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1843 VDD.t847 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t68 VDD.t846 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1844 VDD.t786 VDD.t784 a_77605_n45765# VDD.t785 sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X1845 16to4_PriorityEncoder_v0p0p1_0.x5.x21.X a_78097_n45737# VDD.t503 VDD.t502 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.167 ps=1.39 w=1 l=0.15
X1846 VDD.t533 frontAnalog_v0p0p1_7.x65.A.t7 a_57123_n34959# VDD.t532 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1847 VDD.t434 frontAnalog_v0p0p1_5.x65.X frontAnalog_v0p0p1_5.RSfetsym_0.x2.Y VDD.t433 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1848 VV16.t3 VV15.t2 GND.t244 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1849 VV5.t14 VV4.t13 GND.t78 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1850 OUT2.t7 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND.t900 GND.t899 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1851 OUT0.t68 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD.t96 VDD.t95 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1852 16to4_PriorityEncoder_v0p0p1_0.x3.A0 a_78525_n53555# VDD.t412 VDD.t411 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.148 ps=1.34 w=1 l=0.15
X1853 GND.t898 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t6 GND.t897 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1854 a_78431_n43045# 16to4_PriorityEncoder_v0p0p1_0.x5.x16.X a_78349_n43045# VDD.t538 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X1855 VV14.t14 VV13.t15 GND.t417 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1856 GND.t701 VDD.t1511 a_77759_n45765# GND.t700 sky130_fd_pr__nfet_01v8 ad=0.132 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X1857 VDD.t845 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t67 VDD.t844 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1858 a_78525_n53555# 16to4_PriorityEncoder_v0p0p1_0.x3.x21.X GND.t652 GND.t651 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1859 VDD.t94 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t67 VDD.t93 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1860 a_77687_n52819# 16to4_PriorityEncoder_v0p0p1_0.x3.EI a_77605_n52819# GND.t68 sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.109 ps=1.36 w=0.42 l=0.15
X1861 w_55000_n52150# VIN.t30 a_53630_n52596# GND.t287 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1862 frontAnalog_v0p0p1_12.RSfetsym_0.x2.Y frontAnalog_v0p0p1_12.x65.X GND.t393 GND.t392 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1863 frontAnalog_v0p0p1_0.RSfetsym_0.QN.t2 frontAnalog_v0p0p1_0.x65.X VDD.t1265 VDD.t1264 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.25
X1864 GND.t1356 16to4_PriorityEncoder_v0p0p1_0.x5.x4.A a_78159_n39549# GND.t1355 sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X1865 frontAnalog_v0p0p1_2.x63.A.t1 frontAnalog_v0p0p1_2.x65.A.t7 VDD.t284 VDD.t277 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1866 VDD.t493 CLK.t85 w_55000_n2928# GND.t535 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1867 frontAnalog_v0p0p1_8.x63.A.t1 frontAnalog_v0p0p1_8.x65.A.t7 a_55268_n47136# GND.t427 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1868 VV12.t2 VV11.t1 GND.t209 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1869 GND.t86 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t2 GND.t85 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1870 a_77775_n51585# 16to4_PriorityEncoder_v0p0p1_0.x3.x19.C a_77687_n51585# GND.t66 sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
X1871 16to4_PriorityEncoder_v0p0p1_0.x5.x14.A a_77637_n40777# GND.t580 GND.t579 sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.112 ps=1.04 w=0.65 l=0.15
X1872 VDD.t843 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t66 VDD.t842 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1873 frontAnalog_v0p0p1_6.RSfetsym_0.x2.Y frontAnalog_v0p0p1_6.x65.X GND.t409 GND.t408 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1874 frontAnalog_v0p0p1_15.RSfetsym_0.x1.Y R0.t12 GND.t1430 GND.t1065 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1875 OUT1.t70 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD.t665 VDD.t664 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1876 a_59577_n8883# frontAnalog_v0p0p1_0.x63.X I14.t0 GND.t70 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1877 frontAnalog_v0p0p1_3.RSfetsym_0.x1.Y frontAnalog_v0p0p1_3.x63.X VDD.t1448 VDD.t1444 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1878 w_55000_n8328# CLK.t86 frontAnalog_v0p0p1_0.x65.A.t2 VDD.t494 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1879 a_59577_n73683# frontAnalog_v0p0p1_12.x63.X I2.t0 GND.t15 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1880 a_59578_n83970# S0.t12 frontAnalog_v0p0p1_15.RSfetsym_0.QN.t2 GND.t1324 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.315 ps=2.72 w=1 l=0.15
X1881 VDD.t346 16to4_PriorityEncoder_v0p0p1_0.x3.EI a_77605_n53805# VDD.t345 sky130_fd_pr__pfet_01v8_hvt ad=0.142 pd=1.34 as=0.0662 ps=0.735 w=0.42 l=0.15
X1882 16to4_PriorityEncoder_v0p0p1_0.x3.x21.X a_78097_n53777# VDD.t336 VDD.t335 sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.167 ps=1.39 w=1 l=0.15
X1883 OUT2.t65 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD.t841 VDD.t840 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1884 I6.t0 frontAnalog_v0p0p1_9.RSfetsym_0.x2.Y GND.t609 GND.t404 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.25
X1885 GND.t1421 16to4_PriorityEncoder_v0p0p1_0.x1.A a_82906_n47995# GND.t1420 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X1886 frontAnalog_v0p0p1_2.RSfetsym_0.QN.t0 I15.t8 VDD.t1015 VDD.t1014 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.3
X1887 GND.t84 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t1 GND.t83 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1888 VV12.t12 VV11.t12 GND.t79 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1889 VV8.t12 VV7.t11 GND.t250 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1890 VV15.t5 VV14.t4 GND.t299 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1891 GND.t1190 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t2 GND.t1189 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1892 a_78183_n45737# VDD.t1512 a_78097_n45737# GND.t702 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X1893 VDD.t495 CLK.t87 w_55000_n67728# GND.t270 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1894 a_59578_n19170# frontAnalog_v0p0p1_4.x65.X frontAnalog_v0p0p1_4.RSfetsym_0.QN.t4 GND.t1478 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.315 ps=2.72 w=1 l=0.15
X1895 VDD.t92 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t66 VDD.t91 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1896 a_77881_n51335# 16to4_PriorityEncoder_v0p0p1_0.x3.x16.C a_77775_n51335# GND.t69 sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
X1897 I7.t2 frontAnalog_v0p0p1_8.x63.X VDD.t996 VDD.t995 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.25
X1898 VDD.t28 frontAnalog_v0p0p1_11.x65.X frontAnalog_v0p0p1_11.RSfetsym_0.x2.Y VDD.t27 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1899 a_78431_n51085# 16to4_PriorityEncoder_v0p0p1_0.x3.x16.X a_78349_n51085# VDD.t836 sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.109 ps=1.36 w=0.42 l=0.15
X1900 VDD.t444 frontAnalog_v0p0p1_2.x63.X frontAnalog_v0p0p1_2.RSfetsym_0.x1.Y VDD.t443 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1901 OUT2.t5 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND.t896 GND.t895 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1902 frontAnalog_v0p0p1_1.RSfetsym_0.x1.Y frontAnalog_v0p0p1_1.x63.X GND.t1528 GND.t1527 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1903 frontAnalog_v0p0p1_14.RSfetsym_0.x2.Y S1.t11 GND.t1491 GND.t1490 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1904 OUT1.t69 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD.t663 VDD.t662 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1905 16to4_PriorityEncoder_v0p0p1_0.x36.Y 16to4_PriorityEncoder_v0p0p1_0.x36.A VDD.t36 VDD.t35 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1906 a_59577_n30483# frontAnalog_v0p0p1_6.x63.X I10.t1 GND.t583 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1907 a_59578_n40770# frontAnalog_v0p0p1_1.x65.X frontAnalog_v0p0p1_1.RSfetsym_0.QN.t2 GND.t512 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.315 ps=2.72 w=1 l=0.15
X1908 VDD.t496 CLK.t88 w_55000_n68350# GND.t536 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1909 GND.t1555 16to4_PriorityEncoder_v0p0p1_0.x3.x19.D a_77881_n52819# GND.t68 sky130_fd_pr__nfet_01v8 ad=0.196 pd=1.33 as=0.0693 ps=0.75 w=0.42 l=0.15
X1910 VDD.t1286 16to4_PriorityEncoder_v0p0p1_0.x5.x14.A a_78315_n41309# VDD.t290 sky130_fd_pr__pfet_01v8_hvt ad=0.148 pd=1.34 as=0.0693 ps=0.75 w=0.42 l=0.15
X1911 GND.t1150 16to4_PriorityEncoder_v0p0p1_0.x3.x4.A a_78159_n47589# GND.t1149 sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X1912 GND.t894 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t4 GND.t893 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1913 VDD.t1313 frontAnalog_v0p0p1_12.x63.A.t7 frontAnalog_v0p0p1_12.x65.A.t0 VDD.t527 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1914 frontAnalog_v0p0p1_2.x63.A.t3 CLK.t89 w_55000_n3550# VDD.t466 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1915 frontAnalog_v0p0p1_13.x65.X a_57123_n67359# GND.t500 GND.t499 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1916 GND.t364 I2.t12 a_59578_n73170# GND.t363 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1917 VV16.t11 VV15.t12 GND.t401 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1918 VDD.t90 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0.t65 VDD.t89 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1919 I15.t1 frontAnalog_v0p0p1_2.x63.X VDD.t442 VDD.t441 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.25
X1920 GND.t1075 frontAnalog_v0p0p1_2.x65.X frontAnalog_v0p0p1_2.RSfetsym_0.x2.Y GND.t1074 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1921 VDD.t497 CLK.t90 w_55000_n24528# GND.t273 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1922 OUT0.t0 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND.t82 GND.t81 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1923 GND.t728 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t4 GND.t727 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1924 16to4_PriorityEncoder_v0p0p1_0.x29.Y 16to4_PriorityEncoder_v0p0p1_0.x29.A VDD.t218 VDD.t217 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1925 frontAnalog_v0p0p1_7.RSfetsym_0.x2.Y frontAnalog_v0p0p1_7.x65.X GND.t1368 GND.t1367 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1926 VDD.t602 frontAnalog_v0p0p1_1.x63.A.t7 a_57123_n41879# VDD.t601 sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1927 GND.t35 16to4_PriorityEncoder_v0p0p1_0.x36.A 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND.t34 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1928 VDD.t1447 frontAnalog_v0p0p1_3.x63.X I13.t2 VDD.t1446 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.25
X1929 VDD.t504 CLK.t91 w_55000_n25150# GND.t549 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1930 16to4_PriorityEncoder_v0p0p1_0.x3.A2 a_78065_n49349# GND.t1016 GND.t1015 sky130_fd_pr__nfet_01v8 ad=0.176 pd=1.84 as=0.102 ps=0.99 w=0.65 l=0.15
X1931 w_55000_n13728# CLK.t92 frontAnalog_v0p0p1_3.x65.A.t3 VDD.t505 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1932 frontAnalog_v0p0p1_8.RSfetsym_0.QN.t0 I7.t9 VDD.t508 VDD.t270 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.3
X1933 GND.t892 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t3 GND.t891 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1934 frontAnalog_v0p0p1_5.x65.X a_57123_n24159# GND.t1541 GND.t290 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1935 GND.t683 I15.t9 a_77725_n42341# GND.t682 sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X1936 frontAnalog_v0p0p1_7.x65.A.t0 frontAnalog_v0p0p1_7.x63.A.t7 a_55268_n36336# GND.t292 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1937 a_53630_n20196# VV13.t17 w_55000_n19128# GND.t446 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1938 a_78183_n53777# 16to4_PriorityEncoder_v0p0p1_0.x3.EI a_78097_n53777# GND.t377 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
X1939 OUT2.t64 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD.t839 VDD.t838 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1940 OUT0.t64 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD.t88 VDD.t87 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1941 frontAnalog_v0p0p1_8.RSfetsym_0.x2.Y frontAnalog_v0p0p1_8.x65.X VDD.t1257 VDD.t1256 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1942 OUT1.t68 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD.t661 VDD.t660 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1943 frontAnalog_v0p0p1_8.RSfetsym_0.x1.Y frontAnalog_v0p0p1_8.x63.X GND.t1055 GND.t1054 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1944 16to4_PriorityEncoder_v0p0p1_0.x35.A 16to4_PriorityEncoder_v0p0p1_0.x34.A VDD.t1485 VDD.t1484 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1945 GND.t330 16to4_PriorityEncoder_v0p0p1_0.x43.A 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND.t329 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1946 GND.t890 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2.t2 GND.t889 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1947 VDD.t628 16to4_PriorityEncoder_v0p0p1_0.x5.x19.C a_77605_n43295# VDD.t627 sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X1948 frontAnalog_v0p0p1_0.x63.A.t0 frontAnalog_v0p0p1_0.x65.A.t7 a_55268_n9336# GND.t253 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1949 OUT1.t67 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD.t659 VDD.t658 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1950 VDD.t657 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t66 VDD.t656 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1951 VDD.t216 16to4_PriorityEncoder_v0p0p1_0.x29.A 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD.t215 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1952 GND.t685 I15.t10 a_59578_n2970# GND.t684 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1953 GND.t256 frontAnalog_v0p0p1_9.x63.A.t7 a_57123_n52679# GND.t255 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X1954 a_55268_n20136# CLK.t93 GND.t551 GND.t550 sky130_fd_pr__nfet_01v8_lvt ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.15
X1955 frontAnalog_v0p0p1_12.RSfetsym_0.QN.t1 frontAnalog_v0p0p1_12.x65.X VDD.t371 VDD.t370 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.25
X1956 16to4_PriorityEncoder_v0p0p1_0.x36.Y 16to4_PriorityEncoder_v0p0p1_0.x36.A GND.t33 GND.t32 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1957 a_16719_n13117.t5 a_16599_n13205.t22 a_16541_n13117.t15 GND.t1037 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1958 VDD.t1125 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3.t64 VDD.t1124 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1959 16to4_PriorityEncoder_v0p0p1_0.x3.x4.A 16to4_PriorityEncoder_v0p0p1_0.x3.EI GND.t376 GND.t375 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1960 VDD.t1445 frontAnalog_v0p0p1_3.x63.X frontAnalog_v0p0p1_3.RSfetsym_0.x1.Y VDD.t1444 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1961 frontAnalog_v0p0p1_10.RSfetsym_0.x1.Y frontAnalog_v0p0p1_10.x63.X VDD.t484 VDD.t483 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1962 VV12.t6 VV11.t7 GND.t589 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1963 VIN.t31 w_55000_n29928# error sky130_fd_pr__cap_var_lvt w=2 l=0.18
X1964 GND.t664 16to4_PriorityEncoder_v0p0p1_0.x2.A a_82906_n51645# GND.t663 sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.0567 ps=0.69 w=0.42 l=0.15
X1965 OUT1.t3 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND.t726 GND.t725 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1966 VDD.t506 CLK.t94 w_55000_n3550# GND.t552 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1967 VDD.t1418 frontAnalog_v0p0p1_4.x65.X frontAnalog_v0p0p1_4.RSfetsym_0.QN.t2 VDD.t1417 sky130_fd_pr__pfet_01v8 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.25
X1968 a_53630_n68796# frontAnalog_v0p0p1_10.IB.t33 GND.t851 GND.t296 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1969 OUT3.t1 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND.t1188 GND.t1187 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1970 VV8.t11 VV7.t10 GND.t78 sky130_fd_pr__res_xhigh_po_5p73 l=2.52
X1971 OUT2.t1 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND.t888 GND.t887 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1972 GND.t554 I7.t10 a_77725_n50381# GND.t553 sky130_fd_pr__nfet_01v8 ad=0.112 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X1973 GND.t724 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t2 GND.t723 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1974 a_82906_n47995# 16to4_PriorityEncoder_v0p0p1_0.x3.A1 GND.t1366 GND.t1365 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X1975 VDD.t655 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t65 VDD.t654 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1976 16to4_PriorityEncoder_v0p0p1_0.x34.A a_82906_n43855# GND.t1494 GND.t1493 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1 ps=0.985 w=0.65 l=0.15
X1977 frontAnalog_v0p0p1_2.x63.X a_57123_n4079# GND.t1558 GND.t1147 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1978 GND.t672 S1.t12 frontAnalog_v0p0p1_14.RSfetsym_0.x2.Y GND.t671 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.0878 ps=0.92 w=0.65 l=0.15
X1979 GND.t485 16to4_PriorityEncoder_v0p0p1_0.x5.x17.A a_78065_n41309# GND.t484 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0693 ps=0.75 w=0.42 l=0.15
X1980 GND.t268 I8.t8 a_77605_n39305# GND.t267 sky130_fd_pr__nfet_01v8 ad=0.102 pd=0.99 as=0.0567 ps=0.69 w=0.42 l=0.15
X1981 GND.t616 frontAnalog_v0p0p1_4.x63.X frontAnalog_v0p0p1_4.RSfetsym_0.x1.Y GND.t615 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1982 frontAnalog_v0p0p1_9.x63.A.t1 frontAnalog_v0p0p1_9.x65.A.t7 VDD.t293 VDD.t262 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1983 GND.t1047 16to4_PriorityEncoder_v0p0p1_0.x28.A 16to4_PriorityEncoder_v0p0p1_0.x29.A GND.t1046 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1984 VDD.t653 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t64 VDD.t652 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1985 frontAnalog_v0p0p1_10.x65.X a_57123_n56559# VDD.t1063 VDD.t1062 sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X1986 OUT3.t0 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND.t1186 GND.t1185 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1987 VDD.t70 16to4_PriorityEncoder_v0p0p1_0.x3.x19.C a_77605_n51335# VDD.t69 sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X1988 a_53630_n25596# frontAnalog_v0p0p1_10.IB.t34 GND.t852 GND.t296 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1989 OUT2.t0 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND.t886 GND.t885 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1990 a_77605_n43295# I10.t12 VDD.t972 VDD.t971 sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.109 ps=1.36 w=0.42 l=0.15
X1991 frontAnalog_v0p0p1_8.x63.A.t3 CLK.t95 w_55000_n46750# VDD.t507 sky130_fd_pr__pfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.35
X1992 GND.t715 frontAnalog_v0p0p1_6.x65.A.t7 a_57123_n29559# GND.t714 sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
X1993 VDD.t604 16to4_PriorityEncoder_v0p0p1_0.x2.A a_82988_n51645# VDD.t603 sky130_fd_pr__pfet_01v8_hvt ad=0.146 pd=1.34 as=0.0441 ps=0.63 w=0.42 l=0.15
X1994 a_16719_n13117.t4 a_16599_n13205.t23 a_16541_n13117.t14 GND.t1038 sky130_fd_pr__nfet_01v8_lvt ad=1.16 pd=8.58 as=1.16 ps=8.58 w=4 l=0.6
X1995 frontAnalog_v0p0p1_13.RSfetsym_0.QN.t0 frontAnalog_v0p0p1_13.RSfetsym_0.x1.Y GND.t1159 GND.t1158 sky130_fd_pr__nfet_01v8 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.25
X1996 GND.t328 16to4_PriorityEncoder_v0p0p1_0.x43.A 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND.t327 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1997 frontAnalog_v0p0p1_12.x63.X a_57123_n74279# GND.t1562 GND.t1533 sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1998 OUT1.t1 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND.t722 GND.t721 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
X1999 GND.t720 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1.t0 GND.t719 sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.0878 ps=0.92 w=0.65 l=0.15
R0 GND.n6414 GND.n506 5.63094e+06
R1 GND.n6464 GND 2.276e+06
R2 GND.n6464 GND 2.00869e+06
R3 GND.n6467 GND 334900
R4 GND.n6412 GND 334900
R5 GND.n5652 GND.n994 273240
R6 GND.n7762 GND 271091
R7 GND GND.n5652 271091
R8 GND.n6467 GND.n706 215600
R9 GND.n6413 GND.n6412 215600
R10 GND.n4770 GND.n4769 98120
R11 GND.n4882 GND.n4880 20340.7
R12 GND.n2266 GND.n2264 20340.7
R13 GND.n7661 GND.n7660 20340.7
R14 GND.n1526 GND.n1524 20340.7
R15 GND.n5363 GND.n5361 20340.7
R16 GND.n3932 GND.n3930 20340.7
R17 GND.n5224 GND.n5222 20340.7
R18 GND.n3824 GND.n3822 20340.7
R19 GND.n3501 GND.n3499 20340.7
R20 GND.n1953 GND.n1951 20340.7
R21 GND.n2428 GND.n2426 20340.7
R22 GND.n2737 GND.n2735 20340.7
R23 GND.n2847 GND.n2845 20340.7
R24 GND.n7659 GND.n170 20169.3
R25 GND.n3218 GND.n3217 15044.8
R26 GND.n2845 GND 13209.6
R27 GND.n4880 GND 13209.6
R28 GND GND.n4664 13209.6
R29 GND GND.n170 13209.6
R30 GND.n3217 GND 13209.6
R31 GND.n2264 GND 13209.6
R32 GND GND.n7661 13209.6
R33 GND.n1524 GND 13209.6
R34 GND.n5361 GND 13209.6
R35 GND.n3930 GND 13209.6
R36 GND.n5222 GND 13209.6
R37 GND.n3822 GND 13209.6
R38 GND.n3499 GND 13209.6
R39 GND.n1951 GND 13209.6
R40 GND.n2426 GND 13209.6
R41 GND.n2735 GND 13209.6
R42 GND.n4664 GND.n179 12525.6
R43 GND.t482 GND.n5 10105.3
R44 GND.n6418 GND.t613 10105.3
R45 GND.n2100 GND.n2099 8769.23
R46 GND.t1559 GND.n1659 6847.68
R47 GND.t1015 GND.n6466 5863.39
R48 GND.n6416 GND.t1362 5863.39
R49 GND GND.n7805 4548.57
R50 GND.n1423 GND.n1416 4526.39
R51 GND.n1409 GND.n1407 4526.39
R52 GND.n1412 GND.n1410 4526.07
R53 GND.n1429 GND.n1424 4525.74
R54 GND.n1437 GND.n1436 4525.74
R55 GND.n1398 GND.n1391 4525.74
R56 GND.n1409 GND.n1406 4525.74
R57 GND.n1431 GND.n1365 4525.09
R58 GND.n1352 GND.n1349 4519.41
R59 GND.n4549 GND.n4545 4519.41
R60 GND.n4544 GND.n4541 4519.41
R61 GND.n4544 GND.n4542 4519.41
R62 GND.n4540 GND.n4537 4519.41
R63 GND.n4536 GND.n4532 4519.41
R64 GND.n1354 GND.n1340 4519.41
R65 GND.n1354 GND.n1341 4519.41
R66 GND.n4531 GND.n4527 4519.41
R67 GND.n4526 GND.n4523 4519.41
R68 GND.n4526 GND.n4524 4519.41
R69 GND.n4518 GND.n4516 4519.41
R70 GND.n4515 GND.n4510 4519.41
R71 GND.n4515 GND.n4511 4519.41
R72 GND.n1348 GND.n1346 4519.41
R73 GND.n1348 GND.n1347 4519.41
R74 GND.n4509 GND.n4505 4519.41
R75 GND.n4509 GND.n4506 4519.41
R76 GND.n4504 GND.n4500 4519.41
R77 GND.n1345 GND.n1342 4519.41
R78 GND.n1345 GND.n1343 4519.41
R79 GND.n4499 GND.n4495 4519.41
R80 GND.n4499 GND.n4496 4519.41
R81 GND.n1380 GND.n1376 4377.09
R82 GND.n7659 GND.n180 4215.55
R83 GND.n4569 GND.n4554 3876.26
R84 GND.n4094 GND.n4079 3876.26
R85 GND.n6414 GND.t669 3455.76
R86 GND.t1205 GND.n5657 3428.59
R87 GND.n6412 GND.n6411 3003.29
R88 GND.n6415 GND.n6231 2817.54
R89 GND.n7805 GND.n4 2744.41
R90 GND.n6419 GND.n994 2744.41
R91 GND.n6465 GND.t590 2656.51
R92 GND.n6462 GND.n6461 2243.42
R93 GND.n6463 GND.n6420 1899.15
R94 GND.n3016 GND.n3015 1773
R95 GND.n2585 GND.n2584 1773
R96 GND.n7187 GND.n7186 1773
R97 GND.n7024 GND.n7023 1773
R98 GND.n6870 GND.n6869 1773
R99 GND.n6716 GND.n6715 1773
R100 GND.n6567 GND.n6566 1773
R101 GND.n6592 GND.n6591 1773
R102 GND.n5544 GND.n5543 1773
R103 GND.n1149 GND.n1148 1773
R104 GND.n3675 GND.n3674 1773
R105 GND.n5072 GND.n5071 1773
R106 GND.n467 GND.n466 1773
R107 GND.n329 GND.n328 1773
R108 GND.n227 GND.n226 1773
R109 GND.n7634 GND.n7633 1773
R110 GND.n6464 GND.n6463 1742.45
R111 GND.n6466 GND.n6465 1566.95
R112 GND.n6466 GND.n5 1560.68
R113 GND.n6419 GND.n6418 1548.15
R114 GND.n6420 GND.n6419 1548.15
R115 GND.n7805 GND.n5 1535.61
R116 GND.t1319 GND.n3322 1402.22
R117 GND.n2961 GND.n2958 1390.42
R118 GND.n2537 GND.n2534 1390.42
R119 GND.n7142 GND.n7139 1390.42
R120 GND.n605 GND.n602 1390.42
R121 GND.n615 GND.n612 1390.42
R122 GND.n625 GND.n622 1390.42
R123 GND.n632 GND.n629 1390.42
R124 GND.n5611 GND.n5608 1390.42
R125 GND.n5476 GND.n5473 1390.42
R126 GND.n1133 GND.n1130 1390.42
R127 GND.n3625 GND.n3622 1390.42
R128 GND.n5019 GND.n5016 1390.42
R129 GND.n414 GND.n411 1390.42
R130 GND.n310 GND.n307 1390.42
R131 GND.n208 GND.n205 1390.42
R132 GND.n190 GND.n187 1390.42
R133 GND.n3018 GND.n3016 1384.79
R134 GND.n2587 GND.n2585 1384.79
R135 GND.n7189 GND.n7187 1384.79
R136 GND.n7026 GND.n7024 1384.79
R137 GND.n6872 GND.n6870 1384.79
R138 GND.n6718 GND.n6716 1384.79
R139 GND.n6569 GND.n6567 1384.79
R140 GND.n6594 GND.n6592 1384.79
R141 GND.n5546 GND.n5544 1384.79
R142 GND.n1151 GND.n1149 1384.79
R143 GND.n3677 GND.n3675 1384.79
R144 GND.n5074 GND.n5072 1384.79
R145 GND.n469 GND.n467 1384.79
R146 GND.n331 GND.n329 1384.79
R147 GND.n229 GND.n227 1384.79
R148 GND.n7636 GND.n7634 1384.79
R149 GND.n6417 GND.n6416 1309.97
R150 GND.n6463 GND.t458 1269.38
R151 GND.t1023 GND 1255.01
R152 GND.t579 GND 1255.01
R153 GND.n4259 GND.n4253 1176.21
R154 GND.n4234 GND.n4229 1176.21
R155 GND.n4219 GND.n4214 1176.21
R156 GND.n4204 GND.n4199 1176.21
R157 GND.n4189 GND.n4184 1176.21
R158 GND.n4170 GND.n4165 1176.21
R159 GND.n4155 GND.n4150 1176.21
R160 GND.n4140 GND.n4135 1176.21
R161 GND.n4125 GND.n4120 1176.21
R162 GND.n4444 GND.n4069 1176.21
R163 GND.n4437 GND.n4427 1176.21
R164 GND.n4422 GND.n4421 1176.21
R165 GND.n4407 GND.n4406 1176.21
R166 GND.n4392 GND.n4391 1176.21
R167 GND.n4377 GND.n4376 1176.21
R168 GND.n4360 GND.n4359 1176.21
R169 GND.n4345 GND.n4344 1176.21
R170 GND.n4330 GND.n4329 1176.21
R171 GND.n4315 GND.n4314 1176.21
R172 GND.n4300 GND.n4299 1176.21
R173 GND.n4279 GND.n4278 1176.21
R174 GND.n4261 GND.n4260 1176.21
R175 GND.n4236 GND.n4235 1176.21
R176 GND.n4221 GND.n4220 1176.21
R177 GND.n4206 GND.n4205 1176.21
R178 GND.n4191 GND.n4190 1176.21
R179 GND.n4172 GND.n4171 1176.21
R180 GND.n4157 GND.n4156 1176.21
R181 GND.n4142 GND.n4141 1176.21
R182 GND.n4127 GND.n4126 1176.21
R183 GND.n4445 GND.n4065 1176.21
R184 GND.n4436 GND.n4431 1176.21
R185 GND.n4420 GND.n4415 1176.21
R186 GND.n4405 GND.n4400 1176.21
R187 GND.n4390 GND.n4385 1176.21
R188 GND.n4375 GND.n4370 1176.21
R189 GND.n4358 GND.n4353 1176.21
R190 GND.n4343 GND.n4338 1176.21
R191 GND.n4328 GND.n4323 1176.21
R192 GND.n4313 GND.n4308 1176.21
R193 GND.n4298 GND.n4291 1176.21
R194 GND.n4277 GND.n4271 1176.21
R195 GND.n4940 GND.n4937 1153.03
R196 GND.n4729 GND.n4726 1153.03
R197 GND.n3224 GND.n3194 1153.03
R198 GND.n2885 GND.n2882 1153.03
R199 GND.n2329 GND.n2326 1153.03
R200 GND.n7732 GND.n7729 1153.03
R201 GND.n1588 GND.n1585 1153.03
R202 GND.n5428 GND.n5425 1153.03
R203 GND.n3993 GND.n3990 1153.03
R204 GND.n5293 GND.n5290 1153.03
R205 GND.n3881 GND.n3878 1153.03
R206 GND.n3554 GND.n3551 1153.03
R207 GND.n2013 GND.n2010 1153.03
R208 GND.n2104 GND.n2101 1153.03
R209 GND.n2481 GND.n2478 1153.03
R210 GND.n2775 GND.n2772 1153.03
R211 GND.n7374 GND.t443 1131.09
R212 GND GND.t576 1129.73
R213 GND.n4916 GND.n4909 1077.71
R214 GND.n4914 GND.n4911 1077.71
R215 GND.n4780 GND.n4775 1077.71
R216 GND.n4780 GND.n4776 1077.71
R217 GND.n4774 GND.n4771 1077.71
R218 GND.n4785 GND.n4781 1077.71
R219 GND.n4785 GND.n4782 1077.71
R220 GND.n4790 GND.n4786 1077.71
R221 GND.n4760 GND.n4752 1077.71
R222 GND.n4762 GND.n4750 1077.71
R223 GND.n1610 GND.n1607 1077.71
R224 GND.n3169 GND.n3166 1077.71
R225 GND.n3171 GND.n3164 1077.71
R226 GND.n1606 GND.n1601 1077.71
R227 GND.n1606 GND.n1602 1077.71
R228 GND.n1615 GND.n1611 1077.71
R229 GND.n1615 GND.n1612 1077.71
R230 GND.n1620 GND.n1616 1077.71
R231 GND.n2904 GND.n2901 1077.71
R232 GND.n2906 GND.n2899 1077.71
R233 GND.n1646 GND.n1641 1077.71
R234 GND.n1646 GND.n1642 1077.71
R235 GND.n1650 GND.n1647 1077.71
R236 GND.n2298 GND.n2295 1077.71
R237 GND.n2300 GND.n2293 1077.71
R238 GND.n1670 GND.n1666 1077.71
R239 GND.n1675 GND.n1671 1077.71
R240 GND.n1675 GND.n1672 1077.71
R241 GND.n7702 GND.n7699 1077.71
R242 GND.n7704 GND.n7697 1077.71
R243 GND.n1689 GND.n1686 1077.71
R244 GND.n1695 GND.n1690 1077.71
R245 GND.n1695 GND.n1691 1077.71
R246 GND.n1558 GND.n1555 1077.71
R247 GND.n1560 GND.n1553 1077.71
R248 GND.n1711 GND.n1706 1077.71
R249 GND.n1711 GND.n1707 1077.71
R250 GND.n1715 GND.n1712 1077.71
R251 GND.n5395 GND.n5392 1077.71
R252 GND.n5397 GND.n5390 1077.71
R253 GND.n1740 GND.n1736 1077.71
R254 GND.n1740 GND.n1737 1077.71
R255 GND.n1745 GND.n1741 1077.71
R256 GND.n3970 GND.n3967 1077.71
R257 GND.n3972 GND.n3965 1077.71
R258 GND.n1731 GND.n1726 1077.71
R259 GND.n1731 GND.n1727 1077.71
R260 GND.n1735 GND.n1732 1077.71
R261 GND.n5256 GND.n5253 1077.71
R262 GND.n5258 GND.n5251 1077.71
R263 GND.n1719 GND.n1716 1077.71
R264 GND.n1725 GND.n1720 1077.71
R265 GND.n1725 GND.n1721 1077.71
R266 GND.n3856 GND.n3853 1077.71
R267 GND.n3858 GND.n3851 1077.71
R268 GND.n1700 GND.n1696 1077.71
R269 GND.n1700 GND.n1697 1077.71
R270 GND.n1705 GND.n1701 1077.71
R271 GND.n3533 GND.n3530 1077.71
R272 GND.n3535 GND.n3528 1077.71
R273 GND.n1681 GND.n1676 1077.71
R274 GND.n1681 GND.n1677 1077.71
R275 GND.n1685 GND.n1682 1077.71
R276 GND.n1985 GND.n1982 1077.71
R277 GND.n1987 GND.n1980 1077.71
R278 GND.n1656 GND.n1651 1077.71
R279 GND.n1665 GND.n1657 1077.71
R280 GND.n1665 GND.n1658 1077.71
R281 GND.n2079 GND.n2078 1077.71
R282 GND.n2084 GND.n2083 1077.71
R283 GND.n1634 GND.n1631 1077.71
R284 GND.n1640 GND.n1635 1077.71
R285 GND.n1640 GND.n1636 1077.71
R286 GND.n2460 GND.n2457 1077.71
R287 GND.n2462 GND.n2455 1077.71
R288 GND.n2803 GND.n2796 1077.71
R289 GND.n2801 GND.n2798 1077.71
R290 GND.n1630 GND.n1625 1077.71
R291 GND.n1630 GND.n1626 1077.71
R292 GND.n1624 GND.n1621 1077.71
R293 GND GND.t1065 1058.96
R294 GND GND.t606 1058.96
R295 GND GND.t16 1058.96
R296 GND GND.t1110 1058.96
R297 GND GND.t4 1058.96
R298 GND GND.t525 1058.96
R299 GND GND.t1398 1058.96
R300 GND GND.t1054 1058.96
R301 GND GND.t1527 1058.96
R302 GND GND.t629 1058.96
R303 GND GND.t584 1058.96
R304 GND GND.t1029 1058.96
R305 GND GND.t615 1058.96
R306 GND GND.t1508 1058.96
R307 GND GND.t71 1058.96
R308 GND GND.t475 1058.96
R309 GND.n4916 GND.n4908 1054.53
R310 GND.n4762 GND.n4749 1054.53
R311 GND.n3171 GND.n3163 1054.53
R312 GND.n2906 GND.n2898 1054.53
R313 GND.n2300 GND.n2292 1054.53
R314 GND.n7704 GND.n7696 1054.53
R315 GND.n1560 GND.n1552 1054.53
R316 GND.n5397 GND.n5389 1054.53
R317 GND.n3972 GND.n3964 1054.53
R318 GND.n5258 GND.n5250 1054.53
R319 GND.n3858 GND.n3850 1054.53
R320 GND.n3535 GND.n3527 1054.53
R321 GND.n1987 GND.n1979 1054.53
R322 GND.n2084 GND.n2082 1054.53
R323 GND.n2462 GND.n2454 1054.53
R324 GND.n2803 GND.n2795 1054.53
R325 GND.n5652 GND.n5651 940.789
R326 GND GND.t679 917.571
R327 GND GND.t626 917.571
R328 GND.n3000 GND.n2996 915.471
R329 GND.n3026 GND.n3025 915.471
R330 GND.n3292 GND.n3291 915.471
R331 GND.n2574 GND.n2570 915.471
R332 GND.n2600 GND.n2599 915.471
R333 GND.n2984 GND.n2983 915.471
R334 GND.n7174 GND.n7170 915.471
R335 GND.n7204 GND.n7203 915.471
R336 GND.n2558 GND.n2557 915.471
R337 GND.n7011 GND.n7007 915.471
R338 GND.n7046 GND.n7045 915.471
R339 GND.n7158 GND.n7157 915.471
R340 GND.n6857 GND.n6853 915.471
R341 GND.n6892 GND.n6891 915.471
R342 GND.n6995 GND.n6994 915.471
R343 GND.n6703 GND.n6699 915.471
R344 GND.n6738 GND.n6737 915.471
R345 GND.n6841 GND.n6840 915.471
R346 GND.n6632 GND.n6628 915.471
R347 GND.n6579 GND.n6578 915.471
R348 GND.n6687 GND.n6686 915.471
R349 GND.n5584 GND.n5580 915.471
R350 GND.n5531 GND.n5530 915.471
R351 GND.n6616 GND.n6615 915.471
R352 GND.n1082 GND.n1078 915.471
R353 GND.n1036 GND.n1035 915.471
R354 GND.n5568 GND.n5567 915.471
R355 GND.n1203 GND.n1199 915.471
R356 GND.n1159 GND.n1158 915.471
R357 GND.n1066 GND.n1065 915.471
R358 GND.n3664 GND.n3660 915.471
R359 GND.n3687 GND.n3686 915.471
R360 GND.n1187 GND.n1186 915.471
R361 GND.n5061 GND.n5057 915.471
R362 GND.n5087 GND.n5086 915.471
R363 GND.n3648 GND.n3647 915.471
R364 GND.n456 GND.n452 915.471
R365 GND.n479 GND.n478 915.471
R366 GND.n5045 GND.n5044 915.471
R367 GND.n387 GND.n383 915.471
R368 GND.n341 GND.n340 915.471
R369 GND.n440 GND.n439 915.471
R370 GND.n283 GND.n279 915.471
R371 GND.n237 GND.n236 915.471
R372 GND.n371 GND.n370 915.471
R373 GND.n186 GND.n182 915.471
R374 GND.n7644 GND.n7643 915.471
R375 GND.n267 GND.n266 915.471
R376 GND.n5321 GND.n1845 896.809
R377 GND.n3305 GND.n3302 841.244
R378 GND.n3002 GND.n2994 841.244
R379 GND.n2576 GND.n2568 841.244
R380 GND.n7176 GND.n7168 841.244
R381 GND.n7013 GND.n7005 841.244
R382 GND.n6859 GND.n6851 841.244
R383 GND.n6705 GND.n6697 841.244
R384 GND.n6634 GND.n6626 841.244
R385 GND.n5586 GND.n5578 841.244
R386 GND.n1084 GND.n1076 841.244
R387 GND.n1205 GND.n1197 841.244
R388 GND.n3666 GND.n3658 841.244
R389 GND.n5063 GND.n5055 841.244
R390 GND.n458 GND.n450 841.244
R391 GND.n389 GND.n381 841.244
R392 GND.n285 GND.n277 841.244
R393 GND.t1081 GND.n7571 808.275
R394 GND.t1341 GND.n7509 808.275
R395 GND.t878 GND.n7447 808.275
R396 GND.t1481 GND.n5112 808.275
R397 GND.t464 GND.n3712 808.275
R398 GND.n5458 GND.t408 808.275
R399 GND.n5515 GND.t1372 808.275
R400 GND.t1381 GND.t1023 806.792
R401 GND.t539 GND.t579 806.792
R402 GND.n1373 GND.n1371 806.47
R403 GND GND.t531 784.713
R404 GND GND.t267 784.713
R405 GND.t590 GND.t381 780.297
R406 GND.t669 GND.t696 780.297
R407 GND.n4826 GND.n4821 778.15
R408 GND.n4826 GND.n4822 778.15
R409 GND.n4625 GND.n4620 778.15
R410 GND.n4625 GND.n4621 778.15
R411 GND.n4619 GND.n4614 778.15
R412 GND.n4619 GND.n4615 778.15
R413 GND.n4714 GND.n4710 778.15
R414 GND.n4714 GND.n4713 778.15
R415 GND.n3127 GND.n3122 778.15
R416 GND.n3127 GND.n3123 778.15
R417 GND.n3385 GND.n3380 778.15
R418 GND.n3385 GND.n3381 778.15
R419 GND.n3121 GND.n3116 778.15
R420 GND.n3121 GND.n3117 778.15
R421 GND.n2703 GND.n2698 778.15
R422 GND.n2703 GND.n2699 778.15
R423 GND.n2373 GND.n2368 778.15
R424 GND.n2373 GND.n2369 778.15
R425 GND.n2210 GND.n2205 778.15
R426 GND.n2210 GND.n2206 778.15
R427 GND.n2154 GND.n2149 778.15
R428 GND.n2154 GND.n2150 778.15
R429 GND.n112 GND.n107 778.15
R430 GND.n112 GND.n108 778.15
R431 GND.n1903 GND.n1898 778.15
R432 GND.n1903 GND.n1899 778.15
R433 GND.n1897 GND.n1892 778.15
R434 GND.n1897 GND.n1893 778.15
R435 GND.n1471 GND.n1466 778.15
R436 GND.n1471 GND.n1467 778.15
R437 GND.n3452 GND.n3447 778.15
R438 GND.n3452 GND.n3448 778.15
R439 GND.n3446 GND.n3441 778.15
R440 GND.n3446 GND.n3442 778.15
R441 GND.n1303 GND.n1298 778.15
R442 GND.n1303 GND.n1299 778.15
R443 GND.n3774 GND.n3769 778.15
R444 GND.n3774 GND.n3770 778.15
R445 GND.n3768 GND.n3763 778.15
R446 GND.n3768 GND.n3764 778.15
R447 GND.n4044 GND.n4039 778.15
R448 GND.n4044 GND.n4040 778.15
R449 GND.n4832 GND.n4827 778.15
R450 GND.n4832 GND.n4828 778.15
R451 GND.n5169 GND.n5164 778.15
R452 GND.n5169 GND.n5165 778.15
R453 GND.n4050 GND.n4045 778.15
R454 GND.n4050 GND.n4046 778.15
R455 GND.n5175 GND.n5170 778.15
R456 GND.n5175 GND.n5171 778.15
R457 GND.n1309 GND.n1304 778.15
R458 GND.n1309 GND.n1305 778.15
R459 GND.n1477 GND.n1472 778.15
R460 GND.n1477 GND.n1473 778.15
R461 GND.n2148 GND.n2143 778.15
R462 GND.n2148 GND.n2144 778.15
R463 GND.n126 GND.n113 778.15
R464 GND.n126 GND.n114 778.15
R465 GND.n2216 GND.n2211 778.15
R466 GND.n2216 GND.n2212 778.15
R467 GND.n2697 GND.n2692 778.15
R468 GND.n2697 GND.n2693 778.15
R469 GND.n2379 GND.n2374 778.15
R470 GND.n2379 GND.n2375 778.15
R471 GND.t553 GND.t387 777.333
R472 GND.t1183 GND.t682 777.333
R473 GND GND.t384 754.5
R474 GND GND.t691 754.5
R475 GND.t1013 GND.t1015 732.088
R476 GND.t1359 GND.t1362 732.088
R477 GND.t675 GND 729.721
R478 GND.t575 GND 729.721
R479 GND GND.t386 726
R480 GND.t692 GND 726
R481 GND.t509 GND.t1525 717.149
R482 GND.t323 GND.t484 717.149
R483 GND.t679 GND.t1149 708.047
R484 GND.t626 GND.t1355 708.047
R485 GND.n6826 GND.t1180 706.715
R486 GND.n6980 GND.t30 706.715
R487 GND.t392 GND.n2625 706.715
R488 GND.t449 GND.n3051 706.715
R489 GND GND.t545 654.159
R490 GND.n6231 GND 654.054
R491 GND.t856 GND.t1013 627.505
R492 GND.t1525 GND.t856 627.505
R493 GND.t384 GND.t1381 627.505
R494 GND.t1563 GND.t1359 627.505
R495 GND.t484 GND.t1563 627.505
R496 GND.t691 GND.t539 627.505
R497 GND.t381 GND.t675 606.898
R498 GND.t1149 GND.t1171 606.898
R499 GND.t1171 GND.t1409 606.898
R500 GND.t696 GND.t575 606.898
R501 GND.t1355 GND.t1063 606.898
R502 GND.t1063 GND.t624 606.898
R503 GND.t378 GND.t1539 601.333
R504 GND.t1549 GND.t699 601.333
R505 GND.n7230 GND.t1497 591.866
R506 GND.n5650 GND.t515 550.154
R507 GND GND.t263 546.497
R508 GND GND.t555 546.497
R509 GND.n3000 GND.n2997 521.471
R510 GND.n2574 GND.n2571 521.471
R511 GND.n7174 GND.n7171 521.471
R512 GND.n7011 GND.n7008 521.471
R513 GND.n6857 GND.n6854 521.471
R514 GND.n6703 GND.n6700 521.471
R515 GND.n6632 GND.n6629 521.471
R516 GND.n5584 GND.n5581 521.471
R517 GND.n1082 GND.n1079 521.471
R518 GND.n1203 GND.n1200 521.471
R519 GND.n3664 GND.n3661 521.471
R520 GND.n5061 GND.n5058 521.471
R521 GND.n456 GND.n453 521.471
R522 GND.n387 GND.n384 521.471
R523 GND.n283 GND.n280 521.471
R524 GND.n186 GND.n183 521.471
R525 GND.n3051 GND.n3050 515.509
R526 GND.n2625 GND.n2624 515.509
R527 GND.n7229 GND.n7228 515.509
R528 GND.n6982 GND.n6980 515.509
R529 GND.n6828 GND.n6826 515.509
R530 GND.n5649 GND.n5648 515.509
R531 GND.n5516 GND.n5515 515.509
R532 GND.n5459 GND.n5458 515.509
R533 GND.n3712 GND.n3711 515.509
R534 GND.n5112 GND.n5111 515.509
R535 GND.n7447 GND.n505 515.509
R536 GND.n7509 GND.n7508 515.509
R537 GND.n7571 GND.n7570 515.509
R538 GND.t1345 GND 513.333
R539 GND.t1514 GND.t700 498.408
R540 GND.n2963 GND 484.329
R541 GND.n2539 GND 484.329
R542 GND.n7144 GND 484.329
R543 GND.n607 GND 484.329
R544 GND.n617 GND 484.329
R545 GND.n627 GND 484.329
R546 GND.n634 GND 484.329
R547 GND.n5613 GND 484.329
R548 GND.n5478 GND 484.329
R549 GND.n1135 GND 484.329
R550 GND.n3627 GND 484.329
R551 GND.n5021 GND 484.329
R552 GND.n416 GND 484.329
R553 GND.n312 GND 484.329
R554 GND.n210 GND 484.329
R555 GND.n192 GND 484.329
R556 GND.n4944 GND.n4943 480.913
R557 GND.n4735 GND.n4725 480.913
R558 GND.n3230 GND.n3193 480.913
R559 GND.n2889 GND.n2888 480.913
R560 GND.n2333 GND.n2332 480.913
R561 GND.n7736 GND.n7735 480.913
R562 GND.n1592 GND.n1591 480.913
R563 GND.n5432 GND.n5431 480.913
R564 GND.n3999 GND.n3989 480.913
R565 GND.n5297 GND.n5296 480.913
R566 GND.n3887 GND.n3877 480.913
R567 GND.n3560 GND.n3550 480.913
R568 GND.n2019 GND.n2009 480.913
R569 GND.n2117 GND.n2098 480.913
R570 GND.n2487 GND.n2477 480.913
R571 GND.n2781 GND.n2771 480.913
R572 GND GND.t1514 478.938
R573 GND GND.t509 478.099
R574 GND GND.t323 478.099
R575 GND.n3305 GND.n3303 473.865
R576 GND.n3002 GND.n2995 473.865
R577 GND.n2576 GND.n2569 473.865
R578 GND.n7176 GND.n7169 473.865
R579 GND.n7013 GND.n7006 473.865
R580 GND.n6859 GND.n6852 473.865
R581 GND.n6705 GND.n6698 473.865
R582 GND.n6634 GND.n6627 473.865
R583 GND.n5586 GND.n5579 473.865
R584 GND.n1084 GND.n1077 473.865
R585 GND.n1205 GND.n1198 473.865
R586 GND.n3666 GND.n3659 473.865
R587 GND.n5063 GND.n5056 473.865
R588 GND.n458 GND.n451 473.865
R589 GND.n389 GND.n382 473.865
R590 GND.n285 GND.n278 473.865
R591 GND.n6416 GND.n6415 445.014
R592 GND GND.t1102 426.178
R593 GND.t545 GND.t1440 420.531
R594 GND.n706 GND 420.382
R595 GND.n6413 GND 420.382
R596 GND.t1409 GND.n706 419.048
R597 GND.t624 GND.n6413 419.048
R598 GND.t523 GND.n3153 405.955
R599 GND.t702 GND 393.274
R600 GND.t458 GND.t321 381.594
R601 GND.t489 GND.t1506 373.805
R602 GND.n7445 GND.n506 367.533
R603 GND GND.t69 339.942
R604 GND GND.t687 339.942
R605 GND.n3170 GND.n3165 331.909
R606 GND.n2905 GND.n2900 331.909
R607 GND.n2802 GND.n2797 331.909
R608 GND.n2299 GND.n2294 331.909
R609 GND.n7703 GND.n7698 331.909
R610 GND.n1559 GND.n1554 331.909
R611 GND.n5396 GND.n5391 331.909
R612 GND.n5257 GND.n5252 331.909
R613 GND.n3857 GND.n3852 331.909
R614 GND.n3534 GND.n3529 331.909
R615 GND.n1986 GND.n1981 331.909
R616 GND.n2461 GND.n2456 331.909
R617 GND.n4915 GND.n4910 331.909
R618 GND.n3971 GND.n3966 331.909
R619 GND.n4761 GND.n4751 331.909
R620 GND.n4680 GND.n4679 328.866
R621 GND.n4882 GND.n4881 328.866
R622 GND.n3932 GND.n3931 328.866
R623 GND.n5224 GND.n5223 328.866
R624 GND.n3824 GND.n3823 328.866
R625 GND.n5363 GND.n5362 328.866
R626 GND.n3501 GND.n3500 328.866
R627 GND.n1526 GND.n1525 328.866
R628 GND.n1953 GND.n1952 328.866
R629 GND.n7660 GND.n7659 328.866
R630 GND.n2062 GND.n2061 328.866
R631 GND.n2266 GND.n2265 328.866
R632 GND.n2428 GND.n2427 328.866
R633 GND.n2737 GND.n2736 328.866
R634 GND.n2847 GND.n2846 328.866
R635 GND.t321 GND.t647 327.08
R636 GND.t647 GND.t489 327.08
R637 GND.t1440 GND.t702 327.08
R638 GND.t335 GND.t345 324.212
R639 GND.t357 GND.t347 324.212
R640 GND.t337 GND.t357 324.212
R641 GND.t343 GND.t337 324.212
R642 GND.t353 GND.t343 324.212
R643 GND.t349 GND.t353 324.212
R644 GND.t331 GND.t341 324.212
R645 GND.t339 GND.t327 324.212
R646 GND.t1349 GND.t1345 324.212
R647 GND.t1351 GND.t1349 324.212
R648 GND.t1347 GND.t1351 324.212
R649 GND.t97 GND 308.692
R650 GND GND.t85 308.692
R651 GND.t163 GND 308.692
R652 GND.t1456 GND 308.692
R653 GND GND.t369 306.387
R654 GND.n7806 GND.t847 304.084
R655 GND GND.t339 301.053
R656 GND GND.n6462 299.824
R657 GND.n4498 GND.n4497 293.647
R658 GND.n4503 GND.n4501 293.647
R659 GND.n4503 GND.n4502 293.647
R660 GND.n4508 GND.n4507 293.647
R661 GND.n4514 GND.n4512 293.647
R662 GND.n4514 GND.n4513 293.647
R663 GND.n4521 GND.n4519 293.647
R664 GND.n4521 GND.n4520 293.647
R665 GND.n4530 GND.n4528 293.647
R666 GND.n4530 GND.n4529 293.647
R667 GND.n4535 GND.n4533 293.647
R668 GND.n4535 GND.n4534 293.647
R669 GND.n4539 GND.n4538 293.647
R670 GND.n4548 GND.n4546 293.647
R671 GND.n4548 GND.n4547 293.647
R672 GND.n4493 GND.n4492 293.647
R673 GND.n2112 GND.n2109 290.183
R674 GND.n6229 GND.t351 285.615
R675 GND.n2116 GND.n2100 285.455
R676 GND.t700 GND.t1546 280.354
R677 GND.t1546 GND.t1426 280.354
R678 GND.n3219 GND.n3218 271.185
R679 GND.n6162 GND.t333 270.175
R680 GND.n7804 GND.n7803 267.089
R681 GND GND.t67 266.514
R682 GND GND.t511 266.514
R683 GND.t649 GND 263.26
R684 GND.n5650 GND.n5649 258.123
R685 GND.t1426 GND 253.097
R686 GND.n6418 GND.n6417 250.713
R687 GND.t1506 GND 249.204
R688 GND.t847 GND 244.189
R689 GND GND.t66 230.905
R690 GND GND.t686 230.905
R691 GND GND.t1493 227.501
R692 GND.t1102 GND.t663 223.457
R693 GND.t1100 GND 216.544
R694 GND.t743 GND.n727 214.877
R695 GND.n7803 GND.n7802 213.671
R696 GND.n6465 GND.n6464 213.106
R697 GND.n6230 GND 211.114
R698 GND.n1662 GND.n1661 209.695
R699 GND.n1654 GND.n1653 209.695
R700 GND.n3222 GND.n3221 203.294
R701 GND.n6415 GND.t349 196.843
R702 GND.n4764 GND.n4747 195.531
R703 GND.n3179 GND.n3178 195.531
R704 GND.n2914 GND.n2913 195.531
R705 GND.n2308 GND.n2307 195.531
R706 GND.n7712 GND.n7711 195.531
R707 GND.n1568 GND.n1567 195.531
R708 GND.n5405 GND.n5404 195.531
R709 GND.n3974 GND.n3962 195.531
R710 GND.n5266 GND.n5265 195.531
R711 GND.n3866 GND.n3865 195.531
R712 GND.n3543 GND.n3542 195.531
R713 GND.n1995 GND.n1994 195.531
R714 GND.n2470 GND.n2469 195.531
R715 GND.n2805 GND.n2793 195.531
R716 GND.n4924 GND.n4923 195.531
R717 GND.n1 GND.t368 193.933
R718 GND.n3237 GND.t1067 193.933
R719 GND.n3325 GND.t3 193.933
R720 GND.n7540 GND.t74 193.933
R721 GND.n7512 GND.t1335 193.933
R722 GND.n7602 GND.t476 193.933
R723 GND.n7574 GND.t1075 193.933
R724 GND.n2501 GND.t17 193.933
R725 GND.n2628 GND.t395 193.933
R726 GND.n2918 GND.t867 193.933
R727 GND.n3054 GND.t672 193.933
R728 GND.n6940 GND.t5 193.933
R729 GND.n6925 GND.t24 193.933
R730 GND.n6777 GND.t526 193.933
R731 GND.n6771 GND.t1174 193.933
R732 GND.n66 GND.t1402 193.933
R733 GND.n51 GND.t1432 193.933
R734 GND.n1010 GND.t1530 193.933
R735 GND.n995 GND.t518 193.933
R736 GND.n1239 GND.t585 193.933
R737 GND.n1224 GND.t412 193.933
R738 GND.n7478 GND.t1509 193.933
R739 GND.n7450 GND.t872 193.933
R740 GND.n4977 GND.t619 193.933
R741 GND.n5115 GND.t1484 193.933
R742 GND.n3583 GND.t1030 193.933
R743 GND.n3715 GND.t467 193.933
R744 GND.n1109 GND.t633 193.933
R745 GND.n1103 GND.t1375 193.933
R746 GND.n6531 GND.t1059 193.933
R747 GND.n6503 GND.t1326 193.933
R748 GND.n7109 GND.t1111 193.933
R749 GND.n7081 GND.t1500 193.933
R750 GND.n6201 GND.t1348 193.933
R751 GND.n969 GND.t1049 193.933
R752 GND.n6095 GND.t1138 193.933
R753 GND.t402 GND.n993 193.532
R754 GND.t121 GND.t95 193.508
R755 GND.t207 GND.t121 193.508
R756 GND.t99 GND.t207 193.508
R757 GND.t91 GND.t99 193.508
R758 GND.t113 GND.t91 193.508
R759 GND.t81 GND.t139 193.508
R760 GND.t117 GND.t81 193.508
R761 GND.t187 GND.t117 193.508
R762 GND.t83 GND.t187 193.508
R763 GND.t107 GND.t83 193.508
R764 GND.t171 GND.t107 193.508
R765 GND.t201 GND.t171 193.508
R766 GND.t133 GND.t201 193.508
R767 GND.t177 GND.t133 193.508
R768 GND.t165 GND.t97 193.508
R769 GND.t191 GND.t165 193.508
R770 GND.t89 GND.t191 193.508
R771 GND.t145 GND.t179 193.508
R772 GND.t179 GND.t111 193.508
R773 GND.t111 GND.t149 193.508
R774 GND.t149 GND.t183 193.508
R775 GND.t183 GND.t119 193.508
R776 GND.t119 GND.t199 193.508
R777 GND.t199 GND.t131 193.508
R778 GND.t131 GND.t157 193.508
R779 GND.t157 GND.t205 193.508
R780 GND.t205 GND.t137 193.508
R781 GND.t137 GND.t161 193.508
R782 GND.t85 GND.t143 193.508
R783 GND.t143 GND.t173 193.508
R784 GND.t173 GND.t109 193.508
R785 GND.t109 GND.t195 193.508
R786 GND.t169 GND.t105 193.508
R787 GND.t197 GND.t169 193.508
R788 GND.t127 GND.t197 193.508
R789 GND.t153 GND.t127 193.508
R790 GND.t129 GND.t185 193.508
R791 GND.t155 GND.t129 193.508
R792 GND.t101 GND.t155 193.508
R793 GND.t123 GND.t101 193.508
R794 GND.t141 GND.t123 193.508
R795 GND.t189 GND.t163 193.508
R796 GND.t87 GND.t189 193.508
R797 GND.t167 GND.t87 193.508
R798 GND.t125 GND.t193 193.508
R799 GND.t147 GND.t125 193.508
R800 GND.t181 GND.t147 193.508
R801 GND.t115 GND.t181 193.508
R802 GND.t151 GND.t115 193.508
R803 GND.t93 GND.t151 193.508
R804 GND.t175 GND.t93 193.508
R805 GND.t203 GND.t175 193.508
R806 GND.t135 GND.t203 193.508
R807 GND.t159 GND.t135 193.508
R808 GND.t103 GND.t159 193.508
R809 GND.t1470 GND.t1456 193.508
R810 GND.t1450 GND.t1470 193.508
R811 GND.t1458 GND.t1468 193.508
R812 GND.t1468 GND.t1464 193.508
R813 GND.t1464 GND.t1472 193.508
R814 GND.t1472 GND.t1452 193.508
R815 GND.t1452 GND.t1466 193.508
R816 GND.t1466 GND.t1474 193.508
R817 GND.t1474 GND.t1454 193.508
R818 GND.t1454 GND.t1460 193.508
R819 GND.t1460 GND.t1444 193.508
R820 GND.t1444 GND.t1448 193.508
R821 GND.t1448 GND.t1462 193.508
R822 GND.t1462 GND.t1446 193.508
R823 GND.t369 GND.t371 193.508
R824 GND.t371 GND.t373 193.508
R825 GND.t373 GND.t367 193.508
R826 GND.t663 GND.t1100 193.508
R827 GND.n551 GND.t370 192.982
R828 GND.n3249 GND.t1430 192.982
R829 GND.n3336 GND.t1320 192.982
R830 GND.n7552 GND.t73 192.982
R831 GND.n7523 GND.t1342 192.982
R832 GND.n7614 GND.t480 192.982
R833 GND.n7585 GND.t1082 192.982
R834 GND.n2510 GND.t20 192.982
R835 GND.n2639 GND.t393 192.982
R836 GND.n2927 GND.t607 192.982
R837 GND.n3065 GND.t450 192.982
R838 GND.n6953 GND.t8 192.982
R839 GND.n6931 GND.t31 192.982
R840 GND.n6789 GND.t529 192.982
R841 GND.n6808 GND.t1181 192.982
R842 GND.n79 GND.t1400 192.982
R843 GND.n56 GND.t1439 192.982
R844 GND.n1022 GND.t1528 192.982
R845 GND.n1001 GND.t516 192.982
R846 GND.n1249 GND.t588 192.982
R847 GND.n1230 GND.t409 192.982
R848 GND.n7491 GND.t1512 192.982
R849 GND.n7461 GND.t879 192.982
R850 GND.n4990 GND.t617 192.982
R851 GND.n5126 GND.t1482 192.982
R852 GND.n3592 GND.t1033 192.982
R853 GND.n3726 GND.t465 192.982
R854 GND.n1121 GND.t631 192.982
R855 GND.n5497 GND.t1373 192.982
R856 GND.n6543 GND.t1057 192.982
R857 GND.n6518 GND.t1333 192.982
R858 GND.n7121 GND.t1114 192.982
R859 GND.n7092 GND.t1498 192.982
R860 GND.n6200 GND.t1346 192.982
R861 GND.n959 GND.t1051 192.982
R862 GND.n6085 GND.t1140 192.982
R863 GND GND.t745 190.686
R864 GND.t733 GND 190.686
R865 GND GND.t811 190.686
R866 GND.t222 GND 190.686
R867 GND GND.t1050 189.263
R868 GND.t957 GND.n5861 185.69
R869 GND.t305 GND 185.418
R870 GND GND.t438 185.418
R871 GND GND.t278 185.418
R872 GND.t255 GND 185.418
R873 GND GND.t659 185.418
R874 GND GND.t714 185.418
R875 GND GND.t676 185.418
R876 GND GND.t1391 185.418
R877 GND GND.t390 185.418
R878 GND GND.t1156 185.418
R879 GND GND.t425 185.418
R880 GND GND.t1039 185.418
R881 GND GND.t665 185.418
R882 GND.t275 GND 185.418
R883 GND GND.t251 185.418
R884 GND GND.t862 185.418
R885 GND.n706 GND 182.167
R886 GND.n6413 GND 182.167
R887 GND GND.t68 181.03
R888 GND GND.t247 181.03
R889 GND GND.t177 179.686
R890 GND.t161 GND 179.686
R891 GND GND.t141 179.686
R892 GND.t193 GND.n7375 179.686
R893 GND GND.t103 179.686
R894 GND.t1446 GND 179.686
R895 GND.n4 GND 176.386
R896 GND.n994 GND 176.386
R897 GND.t367 GND 172.775
R898 GND.n2854 GND.n2852 171.047
R899 GND.n3938 GND.n3937 171.047
R900 GND.n5230 GND.n5229 171.047
R901 GND.n3830 GND.n3829 171.047
R902 GND.n5369 GND.n5368 171.047
R903 GND.n3507 GND.n3506 171.047
R904 GND.n1532 GND.n1531 171.047
R905 GND.n1959 GND.n1958 171.047
R906 GND.n7676 GND.n7675 171.047
R907 GND.n2068 GND.n2067 171.047
R908 GND.n2272 GND.n2271 171.047
R909 GND.n2434 GND.n2433 171.047
R910 GND.n2743 GND.n2742 171.047
R911 GND.n4888 GND.n4887 171.047
R912 GND.n4687 GND.n4685 171.047
R913 GND.n3371 GND.n3368 170.613
R914 GND.t959 GND 164.786
R915 GND GND.t947 164.786
R916 GND.t897 GND 164.786
R917 GND GND.t60 164.786
R918 GND GND.t1139 163.555
R919 GND.n6119 GND.t1543 162.326
R920 GND.n4259 GND.n4252 162.236
R921 GND.t105 GND.n7373 161.257
R922 GND.n7797 GND.t1438 159.185
R923 GND.n7826 GND.t1101 154.006
R924 GND.n972 GND.t1366 154.006
R925 GND.n6098 GND.t865 154.006
R926 GND.n4722 GND.n4717 153.601
R927 GND.n4722 GND.n4721 153.601
R928 GND.n3190 GND.n3185 153.601
R929 GND.n3190 GND.n3189 153.601
R930 GND.n2876 GND.n2867 153.601
R931 GND.n2876 GND.n2875 153.601
R932 GND.n2320 GND.n2317 153.601
R933 GND.n2320 GND.n2319 153.601
R934 GND.n7723 GND.n7714 153.601
R935 GND.n7723 GND.n7722 153.601
R936 GND.n1579 GND.n1570 153.601
R937 GND.n1579 GND.n1578 153.601
R938 GND.n5419 GND.n5414 153.601
R939 GND.n5419 GND.n5418 153.601
R940 GND.n3986 GND.n3984 153.601
R941 GND.n3986 GND.n3985 153.601
R942 GND.n5284 GND.n5275 153.601
R943 GND.n5284 GND.n5283 153.601
R944 GND.n3874 GND.n3872 153.601
R945 GND.n3874 GND.n3873 153.601
R946 GND.n3547 GND.n3545 153.601
R947 GND.n3547 GND.n3546 153.601
R948 GND.n2006 GND.n1997 153.601
R949 GND.n2006 GND.n2005 153.601
R950 GND.n2095 GND.n2094 153.601
R951 GND.n2474 GND.n2472 153.601
R952 GND.n2474 GND.n2473 153.601
R953 GND.n2768 GND.n2766 153.601
R954 GND.n2768 GND.n2767 153.601
R955 GND.n4931 GND.n4930 153.601
R956 GND GND.t402 150.841
R957 GND.n28 GND.t604 150.465
R958 GND.n6355 GND.t1507 150.465
R959 GND.n7777 GND.t880 150.465
R960 GND.n653 GND.t510 150.465
R961 GND.n669 GND.t264 150.465
R962 GND.n702 GND.t532 150.465
R963 GND.n6310 GND.t578 150.465
R964 GND.n6281 GND.t324 150.465
R965 GND.n6233 GND.t1068 150.465
R966 GND.n6266 GND.t709 150.465
R967 GND.t1191 GND 149.645
R968 GND.t1221 GND 149.645
R969 GND GND.t1239 149.645
R970 GND GND.t329 149.645
R971 GND.n2852 GND.n2847 148.436
R972 GND.n3937 GND.n3932 148.436
R973 GND.n5229 GND.n5224 148.436
R974 GND.n3829 GND.n3824 148.436
R975 GND.n5368 GND.n5363 148.436
R976 GND.n3506 GND.n3501 148.436
R977 GND.n1531 GND.n1526 148.436
R978 GND.n1958 GND.n1953 148.436
R979 GND.n2067 GND.n2062 148.436
R980 GND.n2271 GND.n2266 148.436
R981 GND.n2433 GND.n2428 148.436
R982 GND.n2742 GND.n2737 148.436
R983 GND.n4887 GND.n4882 148.436
R984 GND.n4685 GND.n4680 148.436
R985 GND.t1332 GND.n6500 140.822
R986 GND.n7805 GND 138.286
R987 GND.n6420 GND 138.286
R988 GND.t1420 GND.t649 138.035
R989 GND.n4758 GND.n4757 137.827
R990 GND.n7763 GND.n7762 137.55
R991 GND GND.t1365 133.766
R992 GND.n4491 GND.n1845 130.844
R993 GND.t1543 GND 130.352
R994 GND.n7376 GND.t1458 129.006
R995 GND.n6415 GND.n6414 128.821
R996 GND.n6417 GND.t335 127.368
R997 GND.n6415 GND.t331 127.368
R998 GND.n7286 GND.t113 124.398
R999 GND.n7287 GND.t145 124.398
R1000 GND.n4698 GND.t1147 123.612
R1001 GND.n3154 GND.t523 123.612
R1002 GND.n2283 GND.t1042 123.612
R1003 GND.n7687 GND.t1126 123.612
R1004 GND.n1543 GND.t64 123.612
R1005 GND.n5380 GND.t581 123.612
R1006 GND.n3949 GND.t1357 123.612
R1007 GND.n5241 GND.t76 123.612
R1008 GND.n3841 GND.t290 123.612
R1009 GND.n3518 GND.t420 123.612
R1010 GND.n1970 GND.t487 123.612
R1011 GND.n2445 GND.t499 123.612
R1012 GND.n2754 GND.t1533 123.612
R1013 GND.n2057 GND.t1104 123.612
R1014 GND.n4899 GND.t598 123.612
R1015 GND.n2822 GND.t1097 123.612
R1016 GND.n4707 GND.n4706 123.472
R1017 GND.n3245 GND.n3244 121.112
R1018 GND.n3346 GND.n3345 121.112
R1019 GND.n7548 GND.n7547 121.112
R1020 GND.n7533 GND.n7532 121.112
R1021 GND.n7610 GND.n7609 121.112
R1022 GND.n7595 GND.n7594 121.112
R1023 GND.n2518 GND.n2517 121.112
R1024 GND.n2649 GND.n2648 121.112
R1025 GND.n2935 GND.n2934 121.112
R1026 GND.n3075 GND.n3074 121.112
R1027 GND.n6948 GND.n6947 121.112
R1028 GND.n6968 GND.n6967 121.112
R1029 GND.n6785 GND.n6784 121.112
R1030 GND.n6805 GND.n6804 121.112
R1031 GND.n74 GND.n73 121.112
R1032 GND.n53 GND.n52 121.112
R1033 GND.n1018 GND.n1017 121.112
R1034 GND.n5630 GND.n5629 121.112
R1035 GND.n1256 GND.n1255 121.112
R1036 GND.n5446 GND.n5445 121.112
R1037 GND.n7486 GND.n7485 121.112
R1038 GND.n7471 GND.n7470 121.112
R1039 GND.n4985 GND.n4984 121.112
R1040 GND.n5136 GND.n5135 121.112
R1041 GND.n3600 GND.n3599 121.112
R1042 GND.n3736 GND.n3735 121.112
R1043 GND.n1117 GND.n1116 121.112
R1044 GND.n5494 GND.n5493 121.112
R1045 GND.n6539 GND.n6538 121.112
R1046 GND.n6515 GND.n6514 121.112
R1047 GND.n7117 GND.n7116 121.112
R1048 GND.n7102 GND.n7101 121.112
R1049 GND.n4665 GND.t305 120.669
R1050 GND.t438 GND.n3216 120.669
R1051 GND.t278 GND.n2263 120.669
R1052 GND.n7662 GND.t255 120.669
R1053 GND.t659 GND.n1523 120.669
R1054 GND.t714 GND.n5360 120.669
R1055 GND.t676 GND.n3929 120.669
R1056 GND.t1391 GND.n5221 120.669
R1057 GND.t390 GND.n3821 120.669
R1058 GND.t1156 GND.n3498 120.669
R1059 GND.t425 GND.n1950 120.669
R1060 GND.t1039 GND.n2425 120.669
R1061 GND.t665 GND.n2734 120.669
R1062 GND.n2046 GND.t275 120.669
R1063 GND.t251 GND.n4879 120.669
R1064 GND.t862 GND.n2844 120.669
R1065 GND.t769 GND.t743 119.534
R1066 GND.t727 GND.t769 119.534
R1067 GND.t747 GND.t727 119.534
R1068 GND.t739 GND.t747 119.534
R1069 GND.t761 GND.t739 119.534
R1070 GND.t787 GND.t729 119.534
R1071 GND.t729 GND.t765 119.534
R1072 GND.t765 GND.t835 119.534
R1073 GND.t835 GND.t731 119.534
R1074 GND.t731 GND.t755 119.534
R1075 GND.t755 GND.t819 119.534
R1076 GND.t819 GND.t721 119.534
R1077 GND.t721 GND.t781 119.534
R1078 GND.t781 GND.t827 119.534
R1079 GND.t745 GND.t813 119.534
R1080 GND.t813 GND.t839 119.534
R1081 GND.t839 GND.t737 119.534
R1082 GND.t829 GND.t793 119.534
R1083 GND.t759 GND.t829 119.534
R1084 GND.t797 GND.t759 119.534
R1085 GND.t833 GND.t797 119.534
R1086 GND.t767 GND.t833 119.534
R1087 GND.t719 GND.t767 119.534
R1088 GND.t779 GND.t719 119.534
R1089 GND.t805 GND.t779 119.534
R1090 GND.t725 GND.t805 119.534
R1091 GND.t785 GND.t725 119.534
R1092 GND.t809 GND.t785 119.534
R1093 GND.t791 GND.t733 119.534
R1094 GND.t821 GND.t791 119.534
R1095 GND.t757 GND.t821 119.534
R1096 GND.t843 GND.t757 119.534
R1097 GND.t753 GND.t817 119.534
R1098 GND.t817 GND.t845 119.534
R1099 GND.t845 GND.t775 119.534
R1100 GND.t775 GND.t801 119.534
R1101 GND.t801 GND.t823 119.534
R1102 GND.t823 GND.t777 119.534
R1103 GND.t777 GND.t803 119.534
R1104 GND.t803 GND.t749 119.534
R1105 GND.t749 GND.t771 119.534
R1106 GND.t771 GND.t789 119.534
R1107 GND.t811 GND.t837 119.534
R1108 GND.t837 GND.t735 119.534
R1109 GND.t735 GND.t815 119.534
R1110 GND.t773 GND.t841 119.534
R1111 GND.t795 GND.t773 119.534
R1112 GND.t831 GND.t795 119.534
R1113 GND.t763 GND.t831 119.534
R1114 GND.t799 GND.t763 119.534
R1115 GND.t741 GND.t799 119.534
R1116 GND.t825 GND.t741 119.534
R1117 GND.t723 GND.t825 119.534
R1118 GND.t783 GND.t723 119.534
R1119 GND.t807 GND.t783 119.534
R1120 GND.t751 GND.t807 119.534
R1121 GND.t236 GND.t222 119.534
R1122 GND.t216 GND.t236 119.534
R1123 GND.t224 GND.t234 119.534
R1124 GND.t234 GND.t230 119.534
R1125 GND.t230 GND.t238 119.534
R1126 GND.t238 GND.t218 119.534
R1127 GND.t218 GND.t232 119.534
R1128 GND.t232 GND.t240 119.534
R1129 GND.t240 GND.t220 119.534
R1130 GND.t220 GND.t226 119.534
R1131 GND.t226 GND.t210 119.534
R1132 GND.t210 GND.t214 119.534
R1133 GND.t214 GND.t228 119.534
R1134 GND.t228 GND.t212 119.534
R1135 GND.t1050 GND.t1052 119.534
R1136 GND.t1052 GND.t1046 119.534
R1137 GND.t1046 GND.t1048 119.534
R1138 GND.t1365 GND.t1420 119.534
R1139 GND.t1493 GND.t1416 119.285
R1140 GND.t531 GND.t639 119.109
R1141 GND.t263 GND.t673 119.109
R1142 GND.t267 GND.t436 119.109
R1143 GND.t555 GND.t1552 119.109
R1144 GND.n7821 GND.n7820 118.1
R1145 GND.n977 GND.n976 118.1
R1146 GND.n6103 GND.n6102 118.1
R1147 GND.n680 GND.n679 117.984
R1148 GND.n6244 GND.n6243 117.984
R1149 GND.n7235 GND.t96 117.626
R1150 GND.n717 GND.t744 117.626
R1151 GND.n5864 GND.t958 117.626
R1152 GND.n5660 GND.t1206 117.007
R1153 GND.t841 GND.n916 116.689
R1154 GND.n4249 GND.n4248 116.329
R1155 GND.n48 GND.n47 116.052
R1156 GND.n6375 GND.n6374 116.052
R1157 GND.t864 GND 115.596
R1158 GND.n3011 GND.n3010 115.201
R1159 GND.n2591 GND.n2590 115.201
R1160 GND.n7195 GND.n7194 115.201
R1161 GND.n7037 GND.n7036 115.201
R1162 GND.n6883 GND.n6882 115.201
R1163 GND.n6729 GND.n6728 115.201
R1164 GND.n6672 GND.n6671 115.201
R1165 GND.n6601 GND.n6600 115.201
R1166 GND.n5553 GND.n5552 115.201
R1167 GND.n1051 GND.n1050 115.201
R1168 GND.n1172 GND.n1171 115.201
R1169 GND.n5078 GND.n5077 115.201
R1170 GND.n5030 GND.n5029 115.201
R1171 GND.n425 GND.n424 115.201
R1172 GND.n356 GND.n355 115.201
R1173 GND.n252 GND.n251 115.201
R1174 GND.n7230 GND.n7229 114.849
R1175 GND.n555 GND.n554 114.713
R1176 GND.n7380 GND.n7379 114.713
R1177 GND.n592 GND.n591 114.713
R1178 GND.n586 GND.n585 114.713
R1179 GND.n582 GND.n581 114.713
R1180 GND.n576 GND.n575 114.713
R1181 GND.n570 GND.n569 114.713
R1182 GND.n564 GND.n563 114.713
R1183 GND.n7427 GND.n7426 114.713
R1184 GND.n7419 GND.n7418 114.713
R1185 GND.n7412 GND.n7411 114.713
R1186 GND.n7408 GND.n7407 114.713
R1187 GND.n7402 GND.n7401 114.713
R1188 GND.n7396 GND.n7395 114.713
R1189 GND.n7390 GND.n7389 114.713
R1190 GND.n7332 GND.n7331 114.713
R1191 GND.n7339 GND.n7338 114.713
R1192 GND.n7365 GND.n7364 114.713
R1193 GND.n7361 GND.n7360 114.713
R1194 GND.n7355 GND.n7354 114.713
R1195 GND.n7349 GND.n7348 114.713
R1196 GND.n7343 GND.n7342 114.713
R1197 GND.n7248 GND.n7247 114.713
R1198 GND.n7291 GND.n7290 114.713
R1199 GND.n7298 GND.n7297 114.713
R1200 GND.n7302 GND.n7301 114.713
R1201 GND.n7308 GND.n7307 114.713
R1202 GND.n7314 GND.n7313 114.713
R1203 GND.n7320 GND.n7319 114.713
R1204 GND.n7234 GND.n7233 114.713
R1205 GND.n7239 GND.n7238 114.713
R1206 GND.n7281 GND.n7280 114.713
R1207 GND.n7276 GND.n7275 114.713
R1208 GND.n7270 GND.n7269 114.713
R1209 GND.n7264 GND.n7263 114.713
R1210 GND.n7258 GND.n7257 114.713
R1211 GND.n6217 GND.n6216 114.713
R1212 GND.n5820 GND.n5819 114.713
R1213 GND.n5814 GND.n5813 114.713
R1214 GND.n5808 GND.n5807 114.713
R1215 GND.n5804 GND.n5803 114.713
R1216 GND.n5798 GND.n5797 114.713
R1217 GND.n5790 GND.n5789 114.713
R1218 GND.n5784 GND.n5783 114.713
R1219 GND.n5774 GND.n5773 114.713
R1220 GND.n5768 GND.n5767 114.713
R1221 GND.n5761 GND.n5760 114.713
R1222 GND.n5692 GND.n5691 114.713
R1223 GND.n5701 GND.n5700 114.713
R1224 GND.n5707 GND.n5706 114.713
R1225 GND.n5713 GND.n5712 114.713
R1226 GND.n5725 GND.n5724 114.713
R1227 GND.n5731 GND.n5730 114.713
R1228 GND.n5751 GND.n5750 114.713
R1229 GND.n5746 GND.n5745 114.713
R1230 GND.n5739 GND.n5738 114.713
R1231 GND.n5654 GND.n5653 114.713
R1232 GND.n6143 GND.n6142 114.713
R1233 GND.n6156 GND.n6155 114.713
R1234 GND.n6166 GND.n6165 114.713
R1235 GND.n6173 GND.n6172 114.713
R1236 GND.n6177 GND.n6176 114.713
R1237 GND.n6183 GND.n6182 114.713
R1238 GND.n6189 GND.n6188 114.713
R1239 GND.n6196 GND.n6195 114.713
R1240 GND.n5663 GND.n5662 114.713
R1241 GND.n5671 GND.n5670 114.713
R1242 GND.n5677 GND.n5676 114.713
R1243 GND.n5681 GND.n5680 114.713
R1244 GND.n5847 GND.n5846 114.713
R1245 GND.n5841 GND.n5840 114.713
R1246 GND.n5835 GND.n5834 114.713
R1247 GND.n964 GND.n963 114.713
R1248 GND.n708 GND.n707 114.713
R1249 GND.n924 GND.n923 114.713
R1250 GND.n930 GND.n929 114.713
R1251 GND.n934 GND.n933 114.713
R1252 GND.n940 GND.n939 114.713
R1253 GND.n946 GND.n945 114.713
R1254 GND.n952 GND.n951 114.713
R1255 GND.n866 GND.n865 114.713
R1256 GND.n911 GND.n910 114.713
R1257 GND.n904 GND.n903 114.713
R1258 GND.n900 GND.n899 114.713
R1259 GND.n894 GND.n893 114.713
R1260 GND.n888 GND.n887 114.713
R1261 GND.n882 GND.n881 114.713
R1262 GND.n779 GND.n778 114.713
R1263 GND.n712 GND.n711 114.713
R1264 GND.n831 GND.n830 114.713
R1265 GND.n835 GND.n834 114.713
R1266 GND.n841 GND.n840 114.713
R1267 GND.n847 GND.n846 114.713
R1268 GND.n853 GND.n852 114.713
R1269 GND.n767 GND.n766 114.713
R1270 GND.n818 GND.n817 114.713
R1271 GND.n811 GND.n810 114.713
R1272 GND.n807 GND.n806 114.713
R1273 GND.n801 GND.n800 114.713
R1274 GND.n795 GND.n794 114.713
R1275 GND.n789 GND.n788 114.713
R1276 GND.n716 GND.n715 114.713
R1277 GND.n721 GND.n720 114.713
R1278 GND.n732 GND.n731 114.713
R1279 GND.n737 GND.n736 114.713
R1280 GND.n743 GND.n742 114.713
R1281 GND.n749 GND.n748 114.713
R1282 GND.n755 GND.n754 114.713
R1283 GND.n6090 GND.n6089 114.713
R1284 GND.n6042 GND.n6041 114.713
R1285 GND.n6050 GND.n6049 114.713
R1286 GND.n6056 GND.n6055 114.713
R1287 GND.n6060 GND.n6059 114.713
R1288 GND.n6066 GND.n6065 114.713
R1289 GND.n6072 GND.n6071 114.713
R1290 GND.n6078 GND.n6077 114.713
R1291 GND.n6128 GND.n6127 114.713
R1292 GND.n5856 GND.n5855 114.713
R1293 GND.n6008 GND.n6007 114.713
R1294 GND.n6012 GND.n6011 114.713
R1295 GND.n6018 GND.n6017 114.713
R1296 GND.n6024 GND.n6023 114.713
R1297 GND.n6030 GND.n6029 114.713
R1298 GND.n5961 GND.n5960 114.713
R1299 GND.n5968 GND.n5967 114.713
R1300 GND.n5994 GND.n5993 114.713
R1301 GND.n5990 GND.n5989 114.713
R1302 GND.n5984 GND.n5983 114.713
R1303 GND.n5978 GND.n5977 114.713
R1304 GND.n5972 GND.n5971 114.713
R1305 GND.n5877 GND.n5876 114.713
R1306 GND.n5920 GND.n5919 114.713
R1307 GND.n5927 GND.n5926 114.713
R1308 GND.n5931 GND.n5930 114.713
R1309 GND.n5937 GND.n5936 114.713
R1310 GND.n5943 GND.n5942 114.713
R1311 GND.n5949 GND.n5948 114.713
R1312 GND.n5863 GND.n5862 114.713
R1313 GND.n5868 GND.n5867 114.713
R1314 GND.n5910 GND.n5909 114.713
R1315 GND.n5905 GND.n5904 114.713
R1316 GND.n5899 GND.n5898 114.713
R1317 GND.n5893 GND.n5892 114.713
R1318 GND.n5887 GND.n5886 114.713
R1319 GND.n549 GND.t1457 113.734
R1320 GND.n546 GND.t164 113.734
R1321 GND.n7327 GND.t86 113.734
R1322 GND.n7245 GND.t98 113.734
R1323 GND.n5826 GND.t1192 113.734
R1324 GND.n5690 GND.t1222 113.734
R1325 GND.n5720 GND.t1240 113.734
R1326 GND.n6151 GND.t330 113.734
R1327 GND.n873 GND.t223 113.734
R1328 GND.n861 GND.t812 113.734
R1329 GND.n774 GND.t734 113.734
R1330 GND.n762 GND.t746 113.734
R1331 GND.n6037 GND.t61 113.734
R1332 GND.n5854 GND.t898 113.734
R1333 GND.n5956 GND.t948 113.734
R1334 GND.n5874 GND.t960 113.734
R1335 GND.n7374 GND.t153 112.88
R1336 GND.n40 GND.n39 111.957
R1337 GND.n6367 GND.n6366 111.957
R1338 GND.n6482 GND.n6481 111.957
R1339 GND.n6484 GND.n6483 111.957
R1340 GND.n655 GND.n654 111.957
R1341 GND.n660 GND.n645 111.957
R1342 GND.n6392 GND.n6391 111.957
R1343 GND.n6394 GND.n6393 111.957
R1344 GND.n6283 GND.n6282 111.957
R1345 GND.n6288 GND.n6273 111.957
R1346 GND.n0 GND.t848 111.924
R1347 GND.n6206 GND.t1542 111.924
R1348 GND.n6203 GND.t577 111.924
R1349 GND.n971 GND.t403 111.924
R1350 GND.n6423 GND.t376 111.924
R1351 GND.n6424 GND.t1538 111.924
R1352 GND.n6425 GND.t362 111.924
R1353 GND.n6426 GND.t1407 111.924
R1354 GND.n6427 GND.t1119 111.924
R1355 GND.n508 GND.t694 111.924
R1356 GND.n509 GND.t1377 111.924
R1357 GND.n510 GND.t1429 111.924
R1358 GND.n511 GND.t542 111.924
R1359 GND.n512 GND.t884 111.924
R1360 GND.n6097 GND.t1544 111.924
R1361 GND.n550 GND.t1447 111.296
R1362 GND.n548 GND.t104 111.296
R1363 GND.n545 GND.t142 111.296
R1364 GND.n7326 GND.t162 111.296
R1365 GND.n7244 GND.t178 111.296
R1366 GND.n5827 GND.t1264 111.296
R1367 GND.n5689 GND.t1188 111.296
R1368 GND.n5719 GND.t1186 111.296
R1369 GND.n6150 GND.t1210 111.296
R1370 GND.n6199 GND.t340 111.296
R1371 GND.n958 GND.t213 111.296
R1372 GND.n872 GND.t752 111.296
R1373 GND.n860 GND.t790 111.296
R1374 GND.n773 GND.t810 111.296
R1375 GND.n761 GND.t828 111.296
R1376 GND.n6084 GND.t51 111.296
R1377 GND.n6036 GND.t966 111.296
R1378 GND.n5853 GND.t1004 111.296
R1379 GND.n5955 GND.t896 111.296
R1380 GND.n5873 GND.t912 111.296
R1381 GND.t827 GND 110.996
R1382 GND GND.t809 110.996
R1383 GND.t789 GND 110.996
R1384 GND GND.t751 110.996
R1385 GND.t212 GND 110.996
R1386 GND.n6468 GND.n6467 110.841
R1387 GND.n4896 GND.n4895 109.394
R1388 GND.n4695 GND.n4694 109.394
R1389 GND.n3150 GND.n3149 109.394
R1390 GND.n2819 GND.n2818 109.394
R1391 GND.n2280 GND.n2279 109.394
R1392 GND.n7684 GND.n7683 109.394
R1393 GND.n1540 GND.n1539 109.394
R1394 GND.n5377 GND.n5376 109.394
R1395 GND.n3946 GND.n3945 109.394
R1396 GND.n5238 GND.n5237 109.394
R1397 GND.n3838 GND.n3837 109.394
R1398 GND.n3515 GND.n3514 109.394
R1399 GND.n1967 GND.n1966 109.394
R1400 GND.n2054 GND.n2053 109.394
R1401 GND.n2442 GND.n2441 109.394
R1402 GND.n2751 GND.n2750 109.394
R1403 GND.n30 GND.n29 109.359
R1404 GND.n6357 GND.n6356 109.359
R1405 GND.n7774 GND.n7773 109.314
R1406 GND.n650 GND.n649 109.314
R1407 GND.n6307 GND.n6306 109.314
R1408 GND.n6278 GND.n6277 109.314
R1409 GND.n12 GND.t1556 108.505
R1410 GND.n9 GND.t1555 108.505
R1411 GND.n7770 GND.t385 108.505
R1412 GND.n7767 GND.t383 108.505
R1413 GND.n6337 GND.t1547 108.505
R1414 GND.n6334 GND.t1548 108.505
R1415 GND.n6303 GND.t695 108.505
R1416 GND.n6300 GND.t698 108.505
R1417 GND.n32 GND.n31 108.016
R1418 GND.n6359 GND.n6358 108.016
R1419 GND.n7775 GND.n7772 108.016
R1420 GND.n648 GND.n647 108.016
R1421 GND.n696 GND.n695 108.016
R1422 GND.n700 GND.n670 108.016
R1423 GND.n676 GND.n675 108.016
R1424 GND.n6308 GND.n6305 108.016
R1425 GND.n6276 GND.n6275 108.016
R1426 GND.n6260 GND.n6259 108.016
R1427 GND.n6264 GND.n6234 108.016
R1428 GND.n6240 GND.n6239 108.016
R1429 GND.n2830 GND.n2829 107.24
R1430 GND.n4865 GND.n4864 107.24
R1431 GND.n4656 GND.n4655 107.24
R1432 GND.n3200 GND.n3199 107.24
R1433 GND.n2249 GND.n2248 107.24
R1434 GND.n157 GND.n156 107.24
R1435 GND.n1509 GND.n1508 107.24
R1436 GND.n5346 GND.n5345 107.24
R1437 GND.n3915 GND.n3914 107.24
R1438 GND.n5207 GND.n5206 107.24
R1439 GND.n3807 GND.n3806 107.24
R1440 GND.n3484 GND.n3483 107.24
R1441 GND.n1936 GND.n1935 107.24
R1442 GND.n2038 GND.n2037 107.24
R1443 GND.n2411 GND.n2410 107.24
R1444 GND.n2720 GND.n2719 107.24
R1445 GND.t1048 GND 106.728
R1446 GND.n693 GND.n692 105.975
R1447 GND.n673 GND.n672 105.975
R1448 GND.n683 GND.n678 105.975
R1449 GND.n6257 GND.n6256 105.975
R1450 GND.n6237 GND.n6236 105.975
R1451 GND.n6247 GND.n6242 105.975
R1452 GND.n824 GND.t753 105.305
R1453 GND.n5651 GND.t375 103.51
R1454 GND.t983 GND.t957 103.299
R1455 GND.t941 GND.t983 103.299
R1456 GND.t961 GND.t941 103.299
R1457 GND.t953 GND.t961 103.299
R1458 GND.t975 GND.t953 103.299
R1459 GND.t943 GND.t1001 103.299
R1460 GND.t979 GND.t943 103.299
R1461 GND.t921 GND.t979 103.299
R1462 GND.t945 GND.t921 103.299
R1463 GND.t969 GND.t945 103.299
R1464 GND.t905 GND.t969 103.299
R1465 GND.t935 GND.t905 103.299
R1466 GND.t995 GND.t935 103.299
R1467 GND.t911 GND.t995 103.299
R1468 GND.t899 GND.t959 103.299
R1469 GND.t925 GND.t899 103.299
R1470 GND.t951 GND.t925 103.299
R1471 GND.t1007 GND.t913 103.299
R1472 GND.t913 GND.t973 103.299
R1473 GND.t973 GND.t1011 103.299
R1474 GND.t1011 GND.t917 103.299
R1475 GND.t917 GND.t981 103.299
R1476 GND.t981 GND.t933 103.299
R1477 GND.t933 GND.t993 103.299
R1478 GND.t993 GND.t891 103.299
R1479 GND.t891 GND.t939 103.299
R1480 GND.t939 GND.t999 103.299
R1481 GND.t999 GND.t895 103.299
R1482 GND.t947 GND.t1005 103.299
R1483 GND.t1005 GND.t907 103.299
R1484 GND.t907 GND.t971 103.299
R1485 GND.t971 GND.t929 103.299
R1486 GND.t903 GND.t967 103.299
R1487 GND.t931 GND.t903 103.299
R1488 GND.t989 GND.t931 103.299
R1489 GND.t887 GND.t989 103.299
R1490 GND.t919 GND.t887 103.299
R1491 GND.t991 GND.t919 103.299
R1492 GND.t889 GND.t991 103.299
R1493 GND.t963 GND.t889 103.299
R1494 GND.t985 GND.t963 103.299
R1495 GND.t1003 GND.t985 103.299
R1496 GND.t923 GND.t897 103.299
R1497 GND.t949 GND.t923 103.299
R1498 GND.t901 GND.t949 103.299
R1499 GND.t927 GND.t987 103.299
R1500 GND.t987 GND.t1009 103.299
R1501 GND.t1009 GND.t915 103.299
R1502 GND.t915 GND.t977 103.299
R1503 GND.t977 GND.t885 103.299
R1504 GND.t885 GND.t955 103.299
R1505 GND.t955 GND.t909 103.299
R1506 GND.t909 GND.t937 103.299
R1507 GND.t937 GND.t997 103.299
R1508 GND.t997 GND.t893 103.299
R1509 GND.t893 GND.t965 103.299
R1510 GND.t60 GND.t42 103.299
R1511 GND.t42 GND.t54 103.299
R1512 GND.t62 GND.t40 103.299
R1513 GND.t40 GND.t36 103.299
R1514 GND.t36 GND.t44 103.299
R1515 GND.t44 GND.t56 103.299
R1516 GND.t56 GND.t38 103.299
R1517 GND.t38 GND.t46 103.299
R1518 GND.t46 GND.t58 103.299
R1519 GND.t58 GND.t32 103.299
R1520 GND.t32 GND.t48 103.299
R1521 GND.t48 GND.t52 103.299
R1522 GND.t52 GND.t34 103.299
R1523 GND.t34 GND.t50 103.299
R1524 GND.t1139 GND.t1141 103.299
R1525 GND.t1141 GND.t1135 103.299
R1526 GND.t1135 GND.t1137 103.299
R1527 GND.t1416 GND.t864 103.299
R1528 GND.n4674 GND.n4673 101.948
R1529 GND.n47 GND.t380 101.43
R1530 GND.n6374 GND.t701 101.43
R1531 GND.n4813 GND.n4804 100.894
R1532 GND.n4606 GND.n4597 100.894
R1533 GND.n2672 GND.n2663 100.894
R1534 GND.n3094 GND.n3085 100.894
R1535 GND.n3362 GND.n3356 100.894
R1536 GND.n2197 GND.n2188 100.894
R1537 GND.n2135 GND.n2126 100.894
R1538 GND.n99 GND.n90 100.894
R1539 GND.n1458 GND.n1449 100.894
R1540 GND.n1290 GND.n1281 100.894
R1541 GND.n4017 GND.n4008 100.894
R1542 GND.n5156 GND.n5147 100.894
R1543 GND.n3755 GND.n3746 100.894
R1544 GND.n3433 GND.n3424 100.894
R1545 GND.n1884 GND.n1875 100.894
R1546 GND.n2360 GND.n2351 100.894
R1547 GND.n7659 GND.n181 100.692
R1548 GND GND.t1537 98.3051
R1549 GND GND.t361 98.3051
R1550 GND GND.t1118 98.3051
R1551 GND GND.t1406 97.1486
R1552 GND GND.t911 95.92
R1553 GND.t895 GND 95.92
R1554 GND GND.t1003 95.92
R1555 GND.n6121 GND.t927 95.92
R1556 GND.t965 GND 95.92
R1557 GND.t50 GND 95.92
R1558 GND.t1223 GND.t1205 93.8076
R1559 GND.t1295 GND.t1195 93.8076
R1560 GND.t1195 GND.t1245 93.8076
R1561 GND.t1245 GND.t1281 93.8076
R1562 GND.t1281 GND.t1199 93.8076
R1563 GND.t1199 GND.t1249 93.8076
R1564 GND.t1249 GND.t1285 93.8076
R1565 GND.t1307 GND.t1273 93.8076
R1566 GND.t1203 GND.t1307 93.8076
R1567 GND.t1277 GND.t1203 93.8076
R1568 GND.t1311 GND.t1277 93.8076
R1569 GND.t1237 GND.t1311 93.8076
R1570 GND.t1241 GND.t1191 93.8076
R1571 GND.t1275 GND.t1241 93.8076
R1572 GND.t1227 GND.t1275 93.8076
R1573 GND.t1189 GND.t1227 93.8076
R1574 GND.t1213 GND.t1189 93.8076
R1575 GND.t1269 GND.t1213 93.8076
R1576 GND.t1301 GND.t1269 93.8076
R1577 GND.t1201 GND.t1301 93.8076
R1578 GND.t1253 GND.t1201 93.8076
R1579 GND.t1305 GND.t1253 93.8076
R1580 GND.t1257 GND.t1231 93.8076
R1581 GND.t1289 GND.t1257 93.8076
R1582 GND.t1225 GND.t1289 93.8076
R1583 GND.t1187 GND.t1225 93.8076
R1584 GND.t1293 GND.t1221 93.8076
R1585 GND.t1207 GND.t1293 93.8076
R1586 GND.t1265 GND.t1207 93.8076
R1587 GND.t1297 GND.t1265 93.8076
R1588 GND.t1197 GND.t1297 93.8076
R1589 GND.t1247 GND.t1197 93.8076
R1590 GND.t1283 GND.t1219 93.8076
R1591 GND.t1219 GND.t1251 93.8076
R1592 GND.t1251 GND.t1217 93.8076
R1593 GND.t1217 GND.t1279 93.8076
R1594 GND.t1279 GND.t1309 93.8076
R1595 GND.t1309 GND.t1235 93.8076
R1596 GND.t1235 GND.t1261 93.8076
R1597 GND.t1261 GND.t1185 93.8076
R1598 GND.t1239 GND.t1291 93.8076
R1599 GND.t1291 GND.t1193 93.8076
R1600 GND.t1193 GND.t1243 93.8076
R1601 GND.t1243 GND.t1211 93.8076
R1602 GND.t1211 GND.t1267 93.8076
R1603 GND.t1299 GND.t1215 93.8076
R1604 GND.t1215 GND.t1271 93.8076
R1605 GND.t1271 GND.t1303 93.8076
R1606 GND.t1303 GND.t1229 93.8076
R1607 GND.t1229 GND.t1255 93.8076
R1608 GND.t1255 GND.t1287 93.8076
R1609 GND.t1287 GND.t1233 93.8076
R1610 GND.t1233 GND.t1259 93.8076
R1611 GND.t1259 GND.t1209 93.8076
R1612 GND.t1137 GND 92.2308
R1613 GND.n4848 GND.n4845 91.8593
R1614 GND.n4641 GND.n4638 91.8593
R1615 GND.n2689 GND.n2686 91.8593
R1616 GND.n3113 GND.n3110 91.8593
R1617 GND.n3377 GND.n3374 91.8593
R1618 GND.n2232 GND.n2229 91.8593
R1619 GND.n2170 GND.n2167 91.8593
R1620 GND.n142 GND.n139 91.8593
R1621 GND.n1493 GND.n1490 91.8593
R1622 GND.n1325 GND.n1322 91.8593
R1623 GND.n4036 GND.n4033 91.8593
R1624 GND.n5191 GND.n5188 91.8593
R1625 GND.n3790 GND.n3787 91.8593
R1626 GND.n3468 GND.n3465 91.8593
R1627 GND.n1919 GND.n1916 91.8593
R1628 GND.n2395 GND.n2392 91.8593
R1629 GND.n3301 GND.n3300 90.3534
R1630 GND.n2993 GND.n2992 90.3534
R1631 GND.n2567 GND.n2566 90.3534
R1632 GND.n7167 GND.n7166 90.3534
R1633 GND.n7004 GND.n7003 90.3534
R1634 GND.n6850 GND.n6849 90.3534
R1635 GND.n6696 GND.n6695 90.3534
R1636 GND.n6625 GND.n6624 90.3534
R1637 GND.n5577 GND.n5576 90.3534
R1638 GND.n1075 GND.n1074 90.3534
R1639 GND.n1196 GND.n1195 90.3534
R1640 GND.n3657 GND.n3656 90.3534
R1641 GND.n5054 GND.n5053 90.3534
R1642 GND.n449 GND.n448 90.3534
R1643 GND.n380 GND.n379 90.3534
R1644 GND.n276 GND.n275 90.3534
R1645 GND.n2960 GND.n2959 90.3427
R1646 GND.n207 GND.n206 90.3427
R1647 GND.n189 GND.n188 90.3427
R1648 GND.n7141 GND.n7140 90.3427
R1649 GND.n2536 GND.n2535 90.3427
R1650 GND.n614 GND.n613 90.3427
R1651 GND.n624 GND.n623 90.3427
R1652 GND.n631 GND.n630 90.3427
R1653 GND.n5475 GND.n5474 90.3427
R1654 GND.n3624 GND.n3623 90.3427
R1655 GND.n309 GND.n308 90.3427
R1656 GND.n413 GND.n412 90.3427
R1657 GND.n5018 GND.n5017 90.3427
R1658 GND.n1132 GND.n1131 90.3427
R1659 GND.n5610 GND.n5609 90.3427
R1660 GND.n604 GND.n603 90.3427
R1661 GND.n7806 GND 87.5398
R1662 GND.n5695 GND.t1237 87.1071
R1663 GND GND.t1263 87.1071
R1664 GND GND.t1187 87.1071
R1665 GND.t1185 GND 87.1071
R1666 GND.t1209 GND 87.1071
R1667 GND.n3268 GND.n3267 86.1558
R1668 GND.n7568 GND.n7567 86.1558
R1669 GND.n199 GND.n198 86.1558
R1670 GND.n7134 GND.n7133 86.1558
R1671 GND.n2948 GND.n2947 86.1558
R1672 GND.n610 GND.n609 86.1558
R1673 GND.n620 GND.n619 86.1558
R1674 GND.n6657 GND.n6656 86.1558
R1675 GND.n5519 GND.n5518 86.1558
R1676 GND.n1267 GND.n1266 86.1558
R1677 GND.n7506 GND.n7505 86.1558
R1678 GND.n5007 GND.n5006 86.1558
R1679 GND.n3613 GND.n3612 86.1558
R1680 GND.n5462 GND.n5461 86.1558
R1681 GND.n5645 GND.n5644 86.1558
R1682 GND.n600 GND.n599 86.1558
R1683 GND.n3320 GND.n3319 86.1558
R1684 GND.n3048 GND.n3047 86.1558
R1685 GND.n2622 GND.n2621 86.1558
R1686 GND.n7226 GND.n7225 86.1558
R1687 GND.n6985 GND.n6984 86.1558
R1688 GND.n6831 GND.n6830 86.1558
R1689 GND.n6667 GND.n6666 86.1558
R1690 GND.n637 GND.n636 86.1558
R1691 GND.n5524 GND.n5523 86.1558
R1692 GND.n5468 GND.n5467 86.1558
R1693 GND.n1139 GND.n1138 86.1558
R1694 GND.n3709 GND.n3708 86.1558
R1695 GND.n5109 GND.n5108 86.1558
R1696 GND.n503 GND.n502 86.1558
R1697 GND.n316 GND.n315 86.1558
R1698 GND.n214 GND.n213 86.1558
R1699 GND.t967 GND.n6002 86.0821
R1700 GND.n917 GND.t224 85.3821
R1701 GND.t643 GND.t440 84.4087
R1702 GND.n3105 GND.n3102 83.5572
R1703 GND.n4028 GND.n4025 83.5572
R1704 GND.n5183 GND.n5180 83.5572
R1705 GND.n3782 GND.n3779 83.5572
R1706 GND.n1317 GND.n1314 83.5572
R1707 GND.n3460 GND.n3457 83.5572
R1708 GND.n1485 GND.n1482 83.5572
R1709 GND.n1911 GND.n1908 83.5572
R1710 GND.n134 GND.n131 83.5572
R1711 GND.n2162 GND.n2159 83.5572
R1712 GND.n2224 GND.n2221 83.5572
R1713 GND.n2387 GND.n2384 83.5572
R1714 GND.n2681 GND.n2678 83.5572
R1715 GND.n4840 GND.n4837 83.5572
R1716 GND.n4633 GND.n4630 83.5572
R1717 GND.t793 GND.n823 82.5361
R1718 GND.n5230 GND.n5201 81.2313
R1719 GND.n5369 GND.n5340 81.2313
R1720 GND.n1532 GND.n1503 81.2313
R1721 GND.n7676 GND.n7670 81.2313
R1722 GND.n2272 GND.n2243 81.2313
R1723 GND.n2743 GND.n2714 81.2313
R1724 GND.n4888 GND.n4859 81.2313
R1725 GND.t185 GND.n7374 80.6288
R1726 GND.t1231 GND.n5696 80.4066
R1727 GND.n7659 GND.n171 79.3342
R1728 GND.n4757 GND.n4756 78.6829
R1729 GND.n4728 GND.n4727 74.9181
R1730 GND.n3223 GND.n3222 74.9181
R1731 GND.n2884 GND.n2883 74.9181
R1732 GND.n2328 GND.n2327 74.9181
R1733 GND.n7731 GND.n7730 74.9181
R1734 GND.n1587 GND.n1586 74.9181
R1735 GND.n5427 GND.n5426 74.9181
R1736 GND.n3992 GND.n3991 74.9181
R1737 GND.n5292 GND.n5291 74.9181
R1738 GND.n3880 GND.n3879 74.9181
R1739 GND.n3553 GND.n3552 74.9181
R1740 GND.n2012 GND.n2011 74.9181
R1741 GND.n2103 GND.n2102 74.9181
R1742 GND.n2480 GND.n2479 74.9181
R1743 GND.n2774 GND.n2773 74.9181
R1744 GND.n4939 GND.n4938 74.9181
R1745 GND.t66 GND.t592 73.7614
R1746 GND.t686 GND.t13 73.7614
R1747 GND.n39 GND.t601 72.8576
R1748 GND.n6366 GND.t1441 72.8576
R1749 GND.n6481 GND.t554 72.8576
R1750 GND.n6483 GND.t1540 72.8576
R1751 GND.n654 GND.t1382 72.8576
R1752 GND.n645 GND.t1408 72.8576
R1753 GND.n679 GND.t382 72.8576
R1754 GND.n6391 GND.t683 72.8576
R1755 GND.n6393 GND.t1550 72.8576
R1756 GND.n6282 GND.t1427 72.8576
R1757 GND.n6273 GND.t540 72.8576
R1758 GND.n6243 GND.t697 72.8576
R1759 GND.t401 GND.t257 72.6261
R1760 GND.t299 GND.t289 72.6261
R1761 GND.t21 GND.t250 72.6261
R1762 GND.t79 GND.t244 72.6261
R1763 GND.t589 GND.t78 72.6261
R1764 GND.n706 GND 72.2501
R1765 GND.n6413 GND 72.2501
R1766 GND.t594 GND.n2964 71.7802
R1767 GND.t1044 GND.n2540 71.7802
R1768 GND.t423 GND.n7145 71.7802
R1769 GND.t1158 GND.n608 71.7802
R1770 GND.t622 GND.n618 71.7802
R1771 GND.t404 GND.n628 71.7802
R1772 GND.t1404 GND.n635 71.7802
R1773 GND.t1060 GND.n5614 71.7802
R1774 GND.t473 GND.n5479 71.7802
R1775 GND.t635 GND.n1136 71.7802
R1776 GND.t1154 GND.n3628 71.7802
R1777 GND.t10 GND.n5022 71.7802
R1778 GND.t547 GND.n417 71.7802
R1779 GND.t434 GND.n313 71.7802
R1780 GND.t688 GND.n211 71.7802
R1781 GND.n728 GND.t761 71.1519
R1782 GND.n4917 GND.n4907 70.024
R1783 GND.n4759 GND.n4758 70.024
R1784 GND.n4784 GND.n4783 70.024
R1785 GND.n4789 GND.n4787 70.024
R1786 GND.n4789 GND.n4788 70.024
R1787 GND.n4763 GND.n4748 70.024
R1788 GND.n1623 GND.n1622 70.024
R1789 GND.n2800 GND.n2799 70.024
R1790 GND.n3172 GND.n3162 70.024
R1791 GND.n3168 GND.n3167 70.024
R1792 GND.n1609 GND.n1608 70.024
R1793 GND.n1605 GND.n1603 70.024
R1794 GND.n1605 GND.n1604 70.024
R1795 GND.n2907 GND.n2897 70.024
R1796 GND.n2903 GND.n2902 70.024
R1797 GND.n1619 GND.n1617 70.024
R1798 GND.n1619 GND.n1618 70.024
R1799 GND.n1614 GND.n1613 70.024
R1800 GND.n2301 GND.n2291 70.024
R1801 GND.n2297 GND.n2296 70.024
R1802 GND.n1649 GND.n1648 70.024
R1803 GND.n1645 GND.n1643 70.024
R1804 GND.n1645 GND.n1644 70.024
R1805 GND.n7705 GND.n7695 70.024
R1806 GND.n7701 GND.n7700 70.024
R1807 GND.n1674 GND.n1673 70.024
R1808 GND.n1669 GND.n1667 70.024
R1809 GND.n1669 GND.n1668 70.024
R1810 GND.n1561 GND.n1551 70.024
R1811 GND.n1557 GND.n1556 70.024
R1812 GND.n1694 GND.n1692 70.024
R1813 GND.n1694 GND.n1693 70.024
R1814 GND.n1688 GND.n1687 70.024
R1815 GND.n5398 GND.n5388 70.024
R1816 GND.n5394 GND.n5393 70.024
R1817 GND.n1714 GND.n1713 70.024
R1818 GND.n1710 GND.n1708 70.024
R1819 GND.n1710 GND.n1709 70.024
R1820 GND.n3969 GND.n3968 70.024
R1821 GND.n1739 GND.n1738 70.024
R1822 GND.n1744 GND.n1742 70.024
R1823 GND.n1744 GND.n1743 70.024
R1824 GND.n3973 GND.n3963 70.024
R1825 GND.n5259 GND.n5249 70.024
R1826 GND.n5255 GND.n5254 70.024
R1827 GND.n1734 GND.n1733 70.024
R1828 GND.n1730 GND.n1728 70.024
R1829 GND.n1730 GND.n1729 70.024
R1830 GND.n3859 GND.n3849 70.024
R1831 GND.n3855 GND.n3854 70.024
R1832 GND.n1724 GND.n1722 70.024
R1833 GND.n1724 GND.n1723 70.024
R1834 GND.n1718 GND.n1717 70.024
R1835 GND.n3536 GND.n3526 70.024
R1836 GND.n3532 GND.n3531 70.024
R1837 GND.n1704 GND.n1702 70.024
R1838 GND.n1704 GND.n1703 70.024
R1839 GND.n1699 GND.n1698 70.024
R1840 GND.n1988 GND.n1978 70.024
R1841 GND.n1984 GND.n1983 70.024
R1842 GND.n1684 GND.n1683 70.024
R1843 GND.n1680 GND.n1678 70.024
R1844 GND.n1680 GND.n1679 70.024
R1845 GND.n1664 GND.n1662 70.024
R1846 GND.n1664 GND.n1663 70.024
R1847 GND.n2080 GND.n2077 70.024
R1848 GND.n2085 GND.n2081 70.024
R1849 GND.n1655 GND.n1654 70.024
R1850 GND.n2463 GND.n2453 70.024
R1851 GND.n2459 GND.n2458 70.024
R1852 GND.n1639 GND.n1637 70.024
R1853 GND.n1639 GND.n1638 70.024
R1854 GND.n1633 GND.n1632 70.024
R1855 GND.n1629 GND.n1627 70.024
R1856 GND.n1629 GND.n1628 70.024
R1857 GND.n2804 GND.n2794 70.024
R1858 GND.n4913 GND.n4912 70.024
R1859 GND.n4779 GND.n4777 70.024
R1860 GND.n4779 GND.n4778 70.024
R1861 GND.n4773 GND.n4772 70.024
R1862 GND.t139 GND.n7286 69.1104
R1863 GND.n7287 GND.t89 69.1104
R1864 GND.n6120 GND.t62 68.8658
R1865 GND.n6500 GND.n6499 68.1084
R1866 GND.n13 GND.n12 67.973
R1867 GND.n10 GND.n9 67.973
R1868 GND.n7781 GND.n7770 67.973
R1869 GND.n7768 GND.n7767 67.973
R1870 GND.n6338 GND.n6337 67.973
R1871 GND.n6335 GND.n6334 67.973
R1872 GND.n6314 GND.n6303 67.973
R1873 GND.n6301 GND.n6300 67.973
R1874 GND.n4717 GND.n4716 67.5205
R1875 GND.n123 GND.n122 67.5205
R1876 GND.n5658 GND.t1223 67.0056
R1877 GND.n5915 GND.t975 66.4063
R1878 GND.n5916 GND.t1007 66.4063
R1879 GND.t1267 GND.n5756 64.7721
R1880 GND.n7376 GND.t1450 64.5031
R1881 GND.n7659 GND.n179 64.3169
R1882 GND.t375 GND 61.2963
R1883 GND.t1537 GND 61.2963
R1884 GND.t361 GND 61.2963
R1885 GND.t1406 GND 61.2963
R1886 GND.t1118 GND 61.2963
R1887 GND.n2999 GND.n2998 59.4829
R1888 GND.n282 GND.n281 59.4829
R1889 GND.n185 GND.n184 59.4829
R1890 GND.n7173 GND.n7172 59.4829
R1891 GND.n2573 GND.n2572 59.4829
R1892 GND.n6856 GND.n6855 59.4829
R1893 GND.n6702 GND.n6701 59.4829
R1894 GND.n6631 GND.n6630 59.4829
R1895 GND.n1081 GND.n1080 59.4829
R1896 GND.n3663 GND.n3662 59.4829
R1897 GND.n386 GND.n385 59.4829
R1898 GND.n455 GND.n454 59.4829
R1899 GND.n5060 GND.n5059 59.4829
R1900 GND.n1202 GND.n1201 59.4829
R1901 GND.n5583 GND.n5582 59.4829
R1902 GND.n7010 GND.n7009 59.4829
R1903 GND.n2086 GND.n2080 57.977
R1904 GND.t67 GND.t501 57.8291
R1905 GND.t68 GND.t705 57.8291
R1906 GND.t511 GND.t703 57.8291
R1907 GND.t247 GND.t460 57.8291
R1908 GND.n4924 GND.n4917 57.224
R1909 GND.n4764 GND.n4763 57.224
R1910 GND.n3179 GND.n3172 57.224
R1911 GND.n2914 GND.n2907 57.224
R1912 GND.n2308 GND.n2301 57.224
R1913 GND.n7712 GND.n7705 57.224
R1914 GND.n1568 GND.n1561 57.224
R1915 GND.n5405 GND.n5398 57.224
R1916 GND.n3974 GND.n3973 57.224
R1917 GND.n5266 GND.n5259 57.224
R1918 GND.n3866 GND.n3859 57.224
R1919 GND.n3543 GND.n3536 57.224
R1920 GND.n1995 GND.n1988 57.224
R1921 GND.n2086 GND.n2085 57.224
R1922 GND.n2470 GND.n2463 57.224
R1923 GND.n2805 GND.n2804 57.224
R1924 GND.n6417 GND.t329 56.9548
R1925 GND.n7820 GND.t664 55.7148
R1926 GND.n976 GND.t1421 55.7148
R1927 GND.n6102 GND.t1417 55.7148
R1928 GND.n4754 GND.n4753 54.813
R1929 GND.n3306 GND.n3301 54.66
R1930 GND.n3003 GND.n2993 54.66
R1931 GND.n2577 GND.n2567 54.66
R1932 GND.n7177 GND.n7167 54.66
R1933 GND.n7014 GND.n7004 54.66
R1934 GND.n6860 GND.n6850 54.66
R1935 GND.n6706 GND.n6696 54.66
R1936 GND.n6635 GND.n6625 54.66
R1937 GND.n5587 GND.n5577 54.66
R1938 GND.n1085 GND.n1075 54.66
R1939 GND.n1206 GND.n1196 54.66
R1940 GND.n3667 GND.n3657 54.66
R1941 GND.n5064 GND.n5054 54.66
R1942 GND.n459 GND.n449 54.66
R1943 GND.n390 GND.n380 54.66
R1944 GND.n286 GND.n276 54.66
R1945 GND.t505 GND.t1026 54.5194
R1946 GND.n4 GND 54.5194
R1947 GND.t319 GND.t406 54.5194
R1948 GND.n994 GND 54.5194
R1949 GND.n6162 GND.t355 54.0356
R1950 GND.n5757 GND.t1283 53.6046
R1951 GND.t293 GND.n4791 52.9309
R1952 GND.n4964 GND.t293 52.9309
R1953 GND.n29 GND.t508 52.8576
R1954 GND.n6356 GND.t322 52.8576
R1955 GND.n7773 GND.t1524 52.8576
R1956 GND.n649 GND.t1014 52.8576
R1957 GND.n692 GND.t1413 52.8576
R1958 GND.n672 GND.t1151 52.8576
R1959 GND.n678 GND.t1150 52.8576
R1960 GND.n6306 GND.t486 52.8576
R1961 GND.n6277 GND.t1360 52.8576
R1962 GND.n6256 GND.t868 52.8576
R1963 GND.n6236 GND.t268 52.8576
R1964 GND.n6242 GND.t1356 52.8576
R1965 GND.n7659 GND.n169 51.4154
R1966 GND.n7659 GND.n173 51.4154
R1967 GND.n7659 GND.n175 51.4154
R1968 GND.n7659 GND.n178 51.4154
R1969 GND.n7659 GND.n177 51.4154
R1970 GND.n7659 GND.n176 51.4154
R1971 GND.n7659 GND.n174 51.4154
R1972 GND.n7659 GND.n172 51.4154
R1973 GND.n7659 GND.n167 51.4154
R1974 GND.n7659 GND.n168 51.4154
R1975 GND.n7659 GND.n165 51.4154
R1976 GND.n7659 GND.n166 51.4154
R1977 GND.n4825 GND.n4823 50.5605
R1978 GND.n4825 GND.n4824 50.5605
R1979 GND.n4618 GND.n4616 50.5605
R1980 GND.n4618 GND.n4617 50.5605
R1981 GND.n4716 GND.n4715 50.5605
R1982 GND.n3384 GND.n3382 50.5605
R1983 GND.n3384 GND.n3383 50.5605
R1984 GND.n3126 GND.n3124 50.5605
R1985 GND.n3126 GND.n3125 50.5605
R1986 GND.n3120 GND.n3118 50.5605
R1987 GND.n3120 GND.n3119 50.5605
R1988 GND.n2702 GND.n2700 50.5605
R1989 GND.n2702 GND.n2701 50.5605
R1990 GND.n2209 GND.n2207 50.5605
R1991 GND.n2209 GND.n2208 50.5605
R1992 GND.n2153 GND.n2151 50.5605
R1993 GND.n2153 GND.n2152 50.5605
R1994 GND.n111 GND.n109 50.5605
R1995 GND.n111 GND.n110 50.5605
R1996 GND.n1902 GND.n1900 50.5605
R1997 GND.n1902 GND.n1901 50.5605
R1998 GND.n1470 GND.n1468 50.5605
R1999 GND.n1470 GND.n1469 50.5605
R2000 GND.n3451 GND.n3449 50.5605
R2001 GND.n3451 GND.n3450 50.5605
R2002 GND.n1302 GND.n1300 50.5605
R2003 GND.n1302 GND.n1301 50.5605
R2004 GND.n3773 GND.n3771 50.5605
R2005 GND.n3773 GND.n3772 50.5605
R2006 GND.n4043 GND.n4041 50.5605
R2007 GND.n4043 GND.n4042 50.5605
R2008 GND.n4831 GND.n4829 50.5605
R2009 GND.n4831 GND.n4830 50.5605
R2010 GND.n5168 GND.n5166 50.5605
R2011 GND.n5168 GND.n5167 50.5605
R2012 GND.n4049 GND.n4047 50.5605
R2013 GND.n4049 GND.n4048 50.5605
R2014 GND.n3767 GND.n3765 50.5605
R2015 GND.n3767 GND.n3766 50.5605
R2016 GND.n5174 GND.n5172 50.5605
R2017 GND.n5174 GND.n5173 50.5605
R2018 GND.n3445 GND.n3443 50.5605
R2019 GND.n3445 GND.n3444 50.5605
R2020 GND.n1308 GND.n1306 50.5605
R2021 GND.n1308 GND.n1307 50.5605
R2022 GND.n1896 GND.n1894 50.5605
R2023 GND.n1896 GND.n1895 50.5605
R2024 GND.n1476 GND.n1474 50.5605
R2025 GND.n1476 GND.n1475 50.5605
R2026 GND.n2147 GND.n2145 50.5605
R2027 GND.n2147 GND.n2146 50.5605
R2028 GND.n125 GND.n123 50.5605
R2029 GND.n125 GND.n124 50.5605
R2030 GND.n2372 GND.n2370 50.5605
R2031 GND.n2372 GND.n2371 50.5605
R2032 GND.n2215 GND.n2213 50.5605
R2033 GND.n2215 GND.n2214 50.5605
R2034 GND.n2696 GND.n2694 50.5605
R2035 GND.n2696 GND.n2695 50.5605
R2036 GND.n2378 GND.n2376 50.5605
R2037 GND.n2378 GND.n2377 50.5605
R2038 GND.n4624 GND.n4622 50.5605
R2039 GND.n4624 GND.n4623 50.5605
R2040 GND.n7658 GND.t684 50.1906
R2041 GND.n728 GND.t787 48.3834
R2042 GND.n993 GND 48.3834
R2043 GND.n7805 GND 47.7719
R2044 GND.n6420 GND 47.7719
R2045 GND.n4570 GND.t537 47.2072
R2046 GND.n4096 GND.n4095 47.1486
R2047 GND GND.n6119 46.7305
R2048 GND.n4902 GND.n4894 46.2978
R2049 GND.n3157 GND.n3148 46.2978
R2050 GND.n2286 GND.n2278 46.2978
R2051 GND.n7690 GND.n7682 46.2978
R2052 GND.n1546 GND.n1538 46.2978
R2053 GND.n5383 GND.n5375 46.2978
R2054 GND.n3952 GND.n3944 46.2978
R2055 GND.n5244 GND.n5236 46.2978
R2056 GND.n3844 GND.n3836 46.2978
R2057 GND.n3521 GND.n3513 46.2978
R2058 GND.n1973 GND.n1965 46.2978
R2059 GND.n2448 GND.n2440 46.2978
R2060 GND.n4701 GND.n4693 46.2978
R2061 GND.n2757 GND.n2749 46.2978
R2062 GND.n2861 GND.n2860 46.2978
R2063 GND.n2075 GND.n2074 46.2978
R2064 GND.n7572 GND 46.1266
R2065 GND.n7510 GND 46.1266
R2066 GND.n7448 GND 46.1266
R2067 GND.n5113 GND 46.1266
R2068 GND.n3713 GND 46.1266
R2069 GND GND.n5457 46.1266
R2070 GND GND.n5514 46.1266
R2071 GND GND.n5641 46.1266
R2072 GND.n6501 GND 46.1266
R2073 GND.t610 GND.n192 43.4986
R2074 GND GND.n5650 43.3696
R2075 GND.n4678 GND.n4677 42.8187
R2076 GND.n2052 GND.n2031 42.8187
R2077 GND.n3206 GND.n3205 42.8174
R2078 GND.n2817 GND.n2816 42.8174
R2079 GND.n2242 GND.n2241 42.8174
R2080 GND.n7669 GND.n7668 42.8174
R2081 GND.n1502 GND.n1501 42.8174
R2082 GND.n5339 GND.n5338 42.8174
R2083 GND.n3908 GND.n3907 42.8174
R2084 GND.n5200 GND.n5199 42.8174
R2085 GND.n3800 GND.n3799 42.8174
R2086 GND.n3477 GND.n3476 42.8174
R2087 GND.n1929 GND.n1928 42.8174
R2088 GND.n2404 GND.n2403 42.8174
R2089 GND.n2713 GND.n2712 42.8174
R2090 GND.n4858 GND.n4857 42.8174
R2091 GND.t693 GND.n7445 42.5398
R2092 GND.t561 GND.n3145 40.7031
R2093 GND GND.n6825 40.3307
R2094 GND GND.n6979 40.3307
R2095 GND.n7079 GND 40.3307
R2096 GND.n2626 GND 40.3307
R2097 GND.n3052 GND 40.3307
R2098 GND.n3323 GND 40.3307
R2099 GND.n5757 GND.t1247 40.2035
R2100 GND.t209 GND.n4550 40.0617
R2101 GND.n1353 GND.t417 40.0617
R2102 GND.n4765 GND.n4741 39.6805
R2103 GND.n3180 GND.n3161 39.6805
R2104 GND.n2915 GND.n2896 39.6805
R2105 GND.n2309 GND.n2290 39.6805
R2106 GND.n7713 GND.n7694 39.6805
R2107 GND.n1569 GND.n1550 39.6805
R2108 GND.n5406 GND.n5387 39.6805
R2109 GND.n3975 GND.n3956 39.6805
R2110 GND.n5267 GND.n5248 39.6805
R2111 GND.n3867 GND.n3848 39.6805
R2112 GND.n3544 GND.n3525 39.6805
R2113 GND.n1996 GND.n1977 39.6805
R2114 GND.n2471 GND.n2452 39.6805
R2115 GND.n2806 GND.n2787 39.6805
R2116 GND.n4925 GND.n4906 39.6805
R2117 GND.n6212 GND.n6202 39.2858
R2118 GND.n23 GND.n22 39.2858
R2119 GND.n7791 GND.n7790 39.2858
R2120 GND.n6488 GND.n6478 39.2858
R2121 GND.n6492 GND.n6491 39.2858
R2122 GND.n665 GND.n664 39.2858
R2123 GND.n6348 GND.n6347 39.2858
R2124 GND.n6324 GND.n6323 39.2858
R2125 GND.n6398 GND.n6388 39.2858
R2126 GND.n6402 GND.n6401 39.2858
R2127 GND.n6293 GND.n6292 39.2858
R2128 GND.n19 GND.n6 38.7881
R2129 GND.n7787 GND.n7764 38.7881
R2130 GND.n661 GND.n642 38.7881
R2131 GND.n6344 GND.n6331 38.7881
R2132 GND.n6320 GND.n6297 38.7881
R2133 GND.n6289 GND.n6270 38.7881
R2134 GND.n12 GND.t502 38.7697
R2135 GND.n9 GND.t706 38.7697
R2136 GND.n7770 GND.t593 38.7697
R2137 GND.n7767 GND.t1027 38.7697
R2138 GND.n6337 GND.t704 38.7697
R2139 GND.n6334 GND.t461 38.7697
R2140 GND.n6303 GND.t14 38.7697
R2141 GND.n6300 GND.t407 38.7697
R2142 GND.n682 GND.n680 38.7523
R2143 GND.n6246 GND.n6244 38.7523
R2144 GND.t327 GND.n6229 38.597
R2145 GND.n31 GND.t652 38.5719
R2146 GND.n31 GND.t1123 38.5719
R2147 GND.n6358 GND.t648 38.5719
R2148 GND.n6358 GND.t490 38.5719
R2149 GND.n7772 GND.t506 38.5719
R2150 GND.n7772 GND.t668 38.5719
R2151 GND.n647 GND.t857 38.5719
R2152 GND.n647 GND.t1526 38.5719
R2153 GND.n695 GND.t1383 38.5719
R2154 GND.n695 GND.t1388 38.5719
R2155 GND.n670 GND.t1166 38.5719
R2156 GND.n670 GND.t1120 38.5719
R2157 GND.n675 GND.t1172 38.5719
R2158 GND.n675 GND.t1410 38.5719
R2159 GND.n6305 GND.t320 38.5719
R2160 GND.n6305 GND.t718 38.5719
R2161 GND.n6275 GND.t1564 38.5719
R2162 GND.n6275 GND.t485 38.5719
R2163 GND.n6259 GND.t1099 38.5719
R2164 GND.n6259 GND.t556 38.5719
R2165 GND.n6234 GND.t312 38.5719
R2166 GND.n6234 GND.t708 38.5719
R2167 GND.n6239 GND.t1064 38.5719
R2168 GND.n6239 GND.t625 38.5719
R2169 GND.n823 GND.t737 36.9992
R2170 GND.t1001 GND.n5915 36.8926
R2171 GND.n5916 GND.t951 36.8926
R2172 GND.t533 GND.t1361 36.3723
R2173 GND.t559 GND.t1390 36.3723
R2174 GND.t550 GND.t389 36.3723
R2175 GND.t1133 GND.t1519 36.3723
R2176 GND.t571 GND.t292 36.3723
R2177 GND.t271 GND.t855 36.3723
R2178 GND.t645 GND.t641 36.3723
R2179 GND.t1145 GND.t254 36.3723
R2180 GND.t300 GND.t274 36.3723
R2181 GND.t565 GND.t277 36.3723
R2182 GND.t1143 GND.t1124 36.3723
R2183 GND.t1131 GND.t1379 36.3723
R2184 GND.t569 GND.t861 36.3723
R2185 GND.t302 GND.t1069 36.3723
R2186 GND.t1129 GND.t258 36.3723
R2187 GND.t80 GND.n4553 36.3719
R2188 GND.n2854 GND.n2853 35.6515
R2189 GND.n2434 GND.n2405 35.6515
R2190 GND.n2068 GND.n2060 35.6515
R2191 GND.n1959 GND.n1930 35.6515
R2192 GND.n3507 GND.n3478 35.6515
R2193 GND.n3830 GND.n3801 35.6515
R2194 GND.n3938 GND.n3909 35.6515
R2195 GND.n4687 GND.n4686 35.6515
R2196 GND.n7816 GND.n7815 34.6358
R2197 GND.n38 GND.n37 34.6358
R2198 GND.n41 GND.n26 34.6358
R2199 GND.n45 GND.n26 34.6358
R2200 GND.n46 GND.n45 34.6358
R2201 GND.n6365 GND.n6364 34.6358
R2202 GND.n6368 GND.n6353 34.6358
R2203 GND.n6372 GND.n6353 34.6358
R2204 GND.n6373 GND.n6372 34.6358
R2205 GND.n984 GND.n983 34.6358
R2206 GND.n15 GND.n14 34.6358
R2207 GND.n14 GND.n7 34.6358
R2208 GND.n22 GND.n7 34.6358
R2209 GND.n18 GND.n17 34.6358
R2210 GND.n19 GND.n18 34.6358
R2211 GND.n7783 GND.n7782 34.6358
R2212 GND.n7782 GND.n7765 34.6358
R2213 GND.n7790 GND.n7765 34.6358
R2214 GND.n7786 GND.n7785 34.6358
R2215 GND.n7787 GND.n7786 34.6358
R2216 GND.n6488 GND.n6487 34.6358
R2217 GND.n6491 GND.n6479 34.6358
R2218 GND.n664 GND.n643 34.6358
R2219 GND.n657 GND.n656 34.6358
R2220 GND.n689 GND.n688 34.6358
R2221 GND.n6451 GND.n6450 34.6358
R2222 GND.n6445 GND.n6444 34.6358
R2223 GND.n6433 GND.n6432 34.6358
R2224 GND.n6340 GND.n6339 34.6358
R2225 GND.n6339 GND.n6332 34.6358
R2226 GND.n6347 GND.n6332 34.6358
R2227 GND.n6343 GND.n6342 34.6358
R2228 GND.n6344 GND.n6343 34.6358
R2229 GND.n6316 GND.n6315 34.6358
R2230 GND.n6315 GND.n6298 34.6358
R2231 GND.n6323 GND.n6298 34.6358
R2232 GND.n6319 GND.n6318 34.6358
R2233 GND.n6320 GND.n6319 34.6358
R2234 GND.n6398 GND.n6397 34.6358
R2235 GND.n6401 GND.n6389 34.6358
R2236 GND.n6292 GND.n6271 34.6358
R2237 GND.n6285 GND.n6284 34.6358
R2238 GND.n6253 GND.n6252 34.6358
R2239 GND.n536 GND.n535 34.6358
R2240 GND.n530 GND.n529 34.6358
R2241 GND.n518 GND.n517 34.6358
R2242 GND.n6110 GND.n6109 34.6358
R2243 GND.t54 GND.n6120 34.4331
R2244 GND.n917 GND.t216 34.1532
R2245 GND.n3360 GND.n3359 34.1229
R2246 GND.n6439 GND.n6438 33.8829
R2247 GND.n524 GND.n523 33.8829
R2248 GND.n2829 GND.t1098 33.462
R2249 GND.n2829 GND.t1160 33.462
R2250 GND.n4864 GND.t599 33.462
R2251 GND.n4864 GND.t252 33.462
R2252 GND.n4895 GND.t681 33.462
R2253 GND.n4895 GND.t1488 33.462
R2254 GND.n4655 GND.t1148 33.462
R2255 GND.n4655 GND.t306 33.462
R2256 GND.n4694 GND.t1558 33.462
R2257 GND.n4694 GND.t504 33.462
R2258 GND.n3199 GND.t690 33.462
R2259 GND.n3199 GND.t439 33.462
R2260 GND.n3149 GND.t524 33.462
R2261 GND.n3149 GND.t1385 33.462
R2262 GND.n2818 GND.t1364 33.462
R2263 GND.n2818 GND.t863 33.462
R2264 GND.n2248 GND.t1043 33.462
R2265 GND.n2248 GND.t441 33.462
R2266 GND.n2279 GND.t1522 33.462
R2267 GND.n2279 GND.t279 33.462
R2268 GND.n156 GND.t1127 33.462
R2269 GND.n156 GND.t325 33.462
R2270 GND.n7683 GND.t1162 33.462
R2271 GND.n7683 GND.t256 33.462
R2272 GND.n1508 GND.t65 33.462
R2273 GND.n1508 GND.t1418 33.462
R2274 GND.n1539 GND.t567 33.462
R2275 GND.n1539 GND.t660 33.462
R2276 GND.n5345 GND.t1062 33.462
R2277 GND.n5345 GND.t715 33.462
R2278 GND.n5376 GND.t582 33.462
R2279 GND.n5376 GND.t1518 33.462
R2280 GND.n3914 GND.t1443 33.462
R2281 GND.n3914 GND.t677 33.462
R2282 GND.n3945 GND.t1358 33.462
R2283 GND.n3945 GND.t1070 33.462
R2284 GND.n5206 GND.t621 33.462
R2285 GND.n5206 GND.t1394 33.462
R2286 GND.n5237 GND.t77 33.462
R2287 GND.n5237 GND.t1392 33.462
R2288 GND.n3806 GND.t1541 33.462
R2289 GND.n3806 GND.t521 33.462
R2290 GND.n3837 GND.t291 33.462
R2291 GND.n3837 GND.t391 33.462
R2292 GND.n3483 GND.t421 33.462
R2293 GND.n3483 GND.t1442 33.462
R2294 GND.n3514 GND.t1353 33.462
R2295 GND.n3514 GND.t1157 33.462
R2296 GND.n1935 GND.t1378 33.462
R2297 GND.n1935 GND.t426 33.462
R2298 GND.n1966 GND.t488 33.462
R2299 GND.n1966 GND.t642 33.462
R2300 GND.n2053 GND.t1105 33.462
R2301 GND.n2053 GND.t276 33.462
R2302 GND.n2037 GND.t1117 33.462
R2303 GND.n2037 GND.t1414 33.462
R2304 GND.n2410 GND.t500 33.462
R2305 GND.n2410 GND.t1040 33.462
R2306 GND.n2441 GND.t1165 33.462
R2307 GND.n2441 GND.t1125 33.462
R2308 GND.n2719 GND.t1534 33.462
R2309 GND.n2719 GND.t666 33.462
R2310 GND.n2750 GND.t1562 33.462
R2311 GND.n2750 GND.t1380 33.462
R2312 GND.n7373 GND.t195 32.2518
R2313 GND.n7781 GND.n7780 32.1329
R2314 GND.n6314 GND.n6313 32.1329
R2315 GND.n7659 GND.n7658 31.7876
R2316 GND.n3307 GND.n3306 30.7897
R2317 GND.n3004 GND.n3003 30.7897
R2318 GND.n2578 GND.n2577 30.7897
R2319 GND.n7178 GND.n7177 30.7897
R2320 GND.n7015 GND.n7014 30.7897
R2321 GND.n6861 GND.n6860 30.7897
R2322 GND.n6707 GND.n6706 30.7897
R2323 GND.n6636 GND.n6635 30.7897
R2324 GND.n5588 GND.n5587 30.7897
R2325 GND.n1086 GND.n1085 30.7897
R2326 GND.n1207 GND.n1206 30.7897
R2327 GND.n3668 GND.n3667 30.7897
R2328 GND.n5065 GND.n5064 30.7897
R2329 GND.n460 GND.n459 30.7897
R2330 GND.n391 GND.n390 30.7897
R2331 GND.n287 GND.n286 30.7897
R2332 GND.n2963 GND.n2957 30.5561
R2333 GND.n5756 GND.t1299 29.036
R2334 GND.n7447 GND.n7446 29.0202
R2335 GND.n4818 GND.n4813 28.9511
R2336 GND.n4611 GND.n4606 28.9511
R2337 GND.n2677 GND.n2672 28.9511
R2338 GND.n3099 GND.n3094 28.9511
R2339 GND.n3367 GND.n3362 28.9511
R2340 GND.n2202 GND.n2197 28.9511
R2341 GND.n2140 GND.n2135 28.9511
R2342 GND.n104 GND.n99 28.9511
R2343 GND.n1463 GND.n1458 28.9511
R2344 GND.n1295 GND.n1290 28.9511
R2345 GND.n4022 GND.n4017 28.9511
R2346 GND.n5161 GND.n5156 28.9511
R2347 GND.n3760 GND.n3755 28.9511
R2348 GND.n3438 GND.n3433 28.9511
R2349 GND.n1889 GND.n1884 28.9511
R2350 GND.n2365 GND.n2360 28.9511
R2351 GND.n2963 GND.n2962 28.8988
R2352 GND.n2539 GND.n2538 28.8988
R2353 GND.n7144 GND.n7143 28.8988
R2354 GND.n607 GND.n606 28.8988
R2355 GND.n617 GND.n616 28.8988
R2356 GND.n627 GND.n626 28.8988
R2357 GND.n634 GND.n633 28.8988
R2358 GND.n5613 GND.n5612 28.8988
R2359 GND.n5478 GND.n5477 28.8988
R2360 GND.n1135 GND.n1134 28.8988
R2361 GND.n3627 GND.n3626 28.8988
R2362 GND.n5021 GND.n5020 28.8988
R2363 GND.n416 GND.n415 28.8988
R2364 GND.n312 GND.n311 28.8988
R2365 GND.n210 GND.n209 28.8988
R2366 GND.n3296 GND.n3295 28.8193
R2367 GND.n2988 GND.n2987 28.8193
R2368 GND.n2562 GND.n2561 28.8193
R2369 GND.n7162 GND.n7161 28.8193
R2370 GND.n6999 GND.n6998 28.8193
R2371 GND.n6845 GND.n6844 28.8193
R2372 GND.n6691 GND.n6690 28.8193
R2373 GND.n6620 GND.n6619 28.8193
R2374 GND.n5572 GND.n5571 28.8193
R2375 GND.n1070 GND.n1069 28.8193
R2376 GND.n1191 GND.n1190 28.8193
R2377 GND.n3652 GND.n3651 28.8193
R2378 GND.n5049 GND.n5048 28.8193
R2379 GND.n444 GND.n443 28.8193
R2380 GND.n375 GND.n374 28.8193
R2381 GND.n271 GND.n270 28.8193
R2382 GND.n549 GND.n548 27.8593
R2383 GND.n546 GND.n545 27.8593
R2384 GND.n7327 GND.n7326 27.8593
R2385 GND.n7245 GND.n7244 27.8593
R2386 GND.n5827 GND.n5826 27.8593
R2387 GND.n5720 GND.n5719 27.8593
R2388 GND.n6151 GND.n6150 27.8593
R2389 GND.n873 GND.n872 27.8593
R2390 GND.n861 GND.n860 27.8593
R2391 GND.n774 GND.n773 27.8593
R2392 GND.n762 GND.n761 27.8593
R2393 GND.n6037 GND.n6036 27.8593
R2394 GND.n5854 GND.n5853 27.8593
R2395 GND.n5956 GND.n5955 27.8593
R2396 GND.n5874 GND.n5873 27.8593
R2397 GND.n29 GND.t444 27.5691
R2398 GND.n6356 GND.t459 27.5691
R2399 GND.n7773 GND.t1516 27.5691
R2400 GND.n649 GND.t1016 27.5691
R2401 GND.n692 GND.t674 27.5691
R2402 GND.n672 GND.t640 27.5691
R2403 GND.n678 GND.t680 27.5691
R2404 GND.n6306 GND.t538 27.5691
R2405 GND.n6277 GND.t1363 27.5691
R2406 GND.n6256 GND.t1553 27.5691
R2407 GND.n6236 GND.t437 27.5691
R2408 GND.n6242 GND.t627 27.5691
R2409 GND.n6210 GND.n6201 27.1064
R2410 GND GND.n7796 26.9763
R2411 GND.n4459 GND.t498 26.8697
R2412 GND.n7820 GND.t1103 26.8576
R2413 GND.n976 GND.t650 26.8576
R2414 GND.n6102 GND.t1494 26.8576
R2415 GND.n5658 GND.t1295 26.8025
R2416 GND.n3032 GND.n3031 26.7111
R2417 GND.n243 GND.n242 26.7111
R2418 GND.n7650 GND.n7649 26.7111
R2419 GND.n7210 GND.n7209 26.7111
R2420 GND.n2606 GND.n2605 26.7111
R2421 GND.n6898 GND.n6897 26.7111
R2422 GND.n6744 GND.n6743 26.7111
R2423 GND.n6585 GND.n6584 26.7111
R2424 GND.n1042 GND.n1041 26.7111
R2425 GND.n3693 GND.n3692 26.7111
R2426 GND.n347 GND.n346 26.7111
R2427 GND.n485 GND.n484 26.7111
R2428 GND.n5093 GND.n5092 26.7111
R2429 GND.n1165 GND.n1164 26.7111
R2430 GND.n5537 GND.n5536 26.7111
R2431 GND.n7052 GND.n7051 26.7111
R2432 GND.n6230 GND.t1347 26.1036
R2433 GND.n47 GND.t1164 25.9346
R2434 GND.n6374 GND.t1515 25.9346
R2435 GND.t1074 GND.t1076 25.66
R2436 GND.t1076 GND.t1078 25.66
R2437 GND.t1078 GND.t1081 25.66
R2438 GND.t1334 GND.t1336 25.66
R2439 GND.t1336 GND.t1339 25.66
R2440 GND.t1339 GND.t1341 25.66
R2441 GND.t871 GND.t873 25.66
R2442 GND.t873 GND.t876 25.66
R2443 GND.t876 GND.t878 25.66
R2444 GND.t1483 GND.t1485 25.66
R2445 GND.t1485 GND.t1479 25.66
R2446 GND.t1479 GND.t1481 25.66
R2447 GND.t466 GND.t468 25.66
R2448 GND.t468 GND.t462 25.66
R2449 GND.t462 GND.t464 25.66
R2450 GND.t413 GND.t411 25.66
R2451 GND.t415 GND.t413 25.66
R2452 GND.t408 GND.t415 25.66
R2453 GND.t1367 GND.t1374 25.66
R2454 GND.t1370 GND.t1367 25.66
R2455 GND.t1372 GND.t1370 25.66
R2456 GND.t519 GND.t517 25.66
R2457 GND.t513 GND.t519 25.66
R2458 GND.t515 GND.t513 25.66
R2459 GND.t1325 GND.t1327 25.66
R2460 GND.t1327 GND.t1330 25.66
R2461 GND.t1330 GND.t1332 25.66
R2462 GND.n4570 GND.t12 25.4195
R2463 GND.n4849 GND.n4848 25.0358
R2464 GND.n4642 GND.n4641 25.0358
R2465 GND.n2708 GND.n2689 25.0358
R2466 GND.n3132 GND.n3113 25.0358
R2467 GND.n3388 GND.n3377 25.0358
R2468 GND.n2233 GND.n2232 25.0358
R2469 GND.n2171 GND.n2170 25.0358
R2470 GND.n143 GND.n142 25.0358
R2471 GND.n1494 GND.n1493 25.0358
R2472 GND.n1326 GND.n1325 25.0358
R2473 GND.n4055 GND.n4036 25.0358
R2474 GND.n5192 GND.n5191 25.0358
R2475 GND.n3791 GND.n3790 25.0358
R2476 GND.n3469 GND.n3468 25.0358
R2477 GND.n1920 GND.n1919 25.0358
R2478 GND.n2396 GND.n2395 25.0358
R2479 GND.n554 GND.t372 24.9236
R2480 GND.n554 GND.t374 24.9236
R2481 GND.n7379 GND.t1471 24.9236
R2482 GND.n7379 GND.t1451 24.9236
R2483 GND.n591 GND.t1459 24.9236
R2484 GND.n591 GND.t1469 24.9236
R2485 GND.n585 GND.t1465 24.9236
R2486 GND.n585 GND.t1473 24.9236
R2487 GND.n581 GND.t1453 24.9236
R2488 GND.n581 GND.t1467 24.9236
R2489 GND.n575 GND.t1475 24.9236
R2490 GND.n575 GND.t1455 24.9236
R2491 GND.n569 GND.t1461 24.9236
R2492 GND.n569 GND.t1445 24.9236
R2493 GND.n563 GND.t1449 24.9236
R2494 GND.n563 GND.t1463 24.9236
R2495 GND.n7426 GND.t190 24.9236
R2496 GND.n7426 GND.t88 24.9236
R2497 GND.n7418 GND.t168 24.9236
R2498 GND.n7418 GND.t194 24.9236
R2499 GND.n7411 GND.t126 24.9236
R2500 GND.n7411 GND.t148 24.9236
R2501 GND.n7407 GND.t182 24.9236
R2502 GND.n7407 GND.t116 24.9236
R2503 GND.n7401 GND.t152 24.9236
R2504 GND.n7401 GND.t94 24.9236
R2505 GND.n7395 GND.t176 24.9236
R2506 GND.n7395 GND.t204 24.9236
R2507 GND.n7389 GND.t136 24.9236
R2508 GND.n7389 GND.t160 24.9236
R2509 GND.n7331 GND.t144 24.9236
R2510 GND.n7331 GND.t174 24.9236
R2511 GND.n7338 GND.t110 24.9236
R2512 GND.n7338 GND.t196 24.9236
R2513 GND.n7364 GND.t106 24.9236
R2514 GND.n7364 GND.t170 24.9236
R2515 GND.n7360 GND.t198 24.9236
R2516 GND.n7360 GND.t128 24.9236
R2517 GND.n7354 GND.t154 24.9236
R2518 GND.n7354 GND.t186 24.9236
R2519 GND.n7348 GND.t130 24.9236
R2520 GND.n7348 GND.t156 24.9236
R2521 GND.n7342 GND.t102 24.9236
R2522 GND.n7342 GND.t124 24.9236
R2523 GND.n7247 GND.t166 24.9236
R2524 GND.n7247 GND.t192 24.9236
R2525 GND.n7290 GND.t90 24.9236
R2526 GND.n7290 GND.t146 24.9236
R2527 GND.n7297 GND.t180 24.9236
R2528 GND.n7297 GND.t112 24.9236
R2529 GND.n7301 GND.t150 24.9236
R2530 GND.n7301 GND.t184 24.9236
R2531 GND.n7307 GND.t120 24.9236
R2532 GND.n7307 GND.t200 24.9236
R2533 GND.n7313 GND.t132 24.9236
R2534 GND.n7313 GND.t158 24.9236
R2535 GND.n7319 GND.t206 24.9236
R2536 GND.n7319 GND.t138 24.9236
R2537 GND.n7233 GND.t122 24.9236
R2538 GND.n7233 GND.t208 24.9236
R2539 GND.n7238 GND.t100 24.9236
R2540 GND.n7238 GND.t92 24.9236
R2541 GND.n7280 GND.t114 24.9236
R2542 GND.n7280 GND.t140 24.9236
R2543 GND.n7275 GND.t82 24.9236
R2544 GND.n7275 GND.t118 24.9236
R2545 GND.n7269 GND.t188 24.9236
R2546 GND.n7269 GND.t84 24.9236
R2547 GND.n7263 GND.t108 24.9236
R2548 GND.n7263 GND.t172 24.9236
R2549 GND.n7257 GND.t202 24.9236
R2550 GND.n7257 GND.t134 24.9236
R2551 GND.n3244 GND.t1066 24.9236
R2552 GND.n3244 GND.t1389 24.9236
R2553 GND.n3345 GND.t1 24.9236
R2554 GND.n3345 GND.t1322 24.9236
R2555 GND.n7547 GND.t75 24.9236
R2556 GND.n7547 GND.t72 24.9236
R2557 GND.n7532 GND.t1337 24.9236
R2558 GND.n7532 GND.t1340 24.9236
R2559 GND.n7609 GND.t477 24.9236
R2560 GND.n7609 GND.t479 24.9236
R2561 GND.n7594 GND.t1077 24.9236
R2562 GND.n7594 GND.t1079 24.9236
R2563 GND.n2517 GND.t18 24.9236
R2564 GND.n2517 GND.t19 24.9236
R2565 GND.n2648 GND.t397 24.9236
R2566 GND.n2648 GND.t400 24.9236
R2567 GND.n2934 GND.t866 24.9236
R2568 GND.n2934 GND.t608 24.9236
R2569 GND.n3074 GND.t1491 24.9236
R2570 GND.n3074 GND.t1090 24.9236
R2571 GND.n6947 GND.t6 24.9236
R2572 GND.n6947 GND.t7 24.9236
R2573 GND.n6967 GND.t26 24.9236
R2574 GND.n6967 GND.t29 24.9236
R2575 GND.n6784 GND.t527 24.9236
R2576 GND.n6784 GND.t528 24.9236
R2577 GND.n6804 GND.t1176 24.9236
R2578 GND.n6804 GND.t1179 24.9236
R2579 GND.n73 GND.t1403 24.9236
R2580 GND.n73 GND.t1399 24.9236
R2581 GND.n52 GND.t1434 24.9236
R2582 GND.n52 GND.t1437 24.9236
R2583 GND.n1017 GND.t1531 24.9236
R2584 GND.n1017 GND.t1532 24.9236
R2585 GND.n5629 GND.t520 24.9236
R2586 GND.n5629 GND.t514 24.9236
R2587 GND.n1255 GND.t586 24.9236
R2588 GND.n1255 GND.t587 24.9236
R2589 GND.n5445 GND.t414 24.9236
R2590 GND.n5445 GND.t416 24.9236
R2591 GND.n7485 GND.t1510 24.9236
R2592 GND.n7485 GND.t1511 24.9236
R2593 GND.n7470 GND.t874 24.9236
R2594 GND.n7470 GND.t877 24.9236
R2595 GND.n4984 GND.t620 24.9236
R2596 GND.n4984 GND.t616 24.9236
R2597 GND.n5135 GND.t1486 24.9236
R2598 GND.n5135 GND.t1480 24.9236
R2599 GND.n3599 GND.t1031 24.9236
R2600 GND.n3599 GND.t1032 24.9236
R2601 GND.n3735 GND.t469 24.9236
R2602 GND.n3735 GND.t463 24.9236
R2603 GND.n1116 GND.t634 24.9236
R2604 GND.n1116 GND.t630 24.9236
R2605 GND.n5493 GND.t1368 24.9236
R2606 GND.n5493 GND.t1371 24.9236
R2607 GND.n6538 GND.t1055 24.9236
R2608 GND.n6538 GND.t1056 24.9236
R2609 GND.n6514 GND.t1328 24.9236
R2610 GND.n6514 GND.t1331 24.9236
R2611 GND.n7116 GND.t1112 24.9236
R2612 GND.n7116 GND.t1113 24.9236
R2613 GND.n7101 GND.t1502 24.9236
R2614 GND.n7101 GND.t1496 24.9236
R2615 GND.n6216 GND.t1350 24.9236
R2616 GND.n6216 GND.t1352 24.9236
R2617 GND.n5819 GND.t1242 24.9236
R2618 GND.n5819 GND.t1276 24.9236
R2619 GND.n5813 GND.t1228 24.9236
R2620 GND.n5813 GND.t1190 24.9236
R2621 GND.n5807 GND.t1214 24.9236
R2622 GND.n5807 GND.t1270 24.9236
R2623 GND.n5803 GND.t1302 24.9236
R2624 GND.n5803 GND.t1202 24.9236
R2625 GND.n5797 GND.t1254 24.9236
R2626 GND.n5797 GND.t1306 24.9236
R2627 GND.n5789 GND.t1232 24.9236
R2628 GND.n5789 GND.t1258 24.9236
R2629 GND.n5783 GND.t1290 24.9236
R2630 GND.n5783 GND.t1226 24.9236
R2631 GND.n5773 GND.t1294 24.9236
R2632 GND.n5773 GND.t1208 24.9236
R2633 GND.n5767 GND.t1266 24.9236
R2634 GND.n5767 GND.t1298 24.9236
R2635 GND.n5760 GND.t1198 24.9236
R2636 GND.n5760 GND.t1248 24.9236
R2637 GND.n5691 GND.t1284 24.9236
R2638 GND.n5691 GND.t1220 24.9236
R2639 GND.n5700 GND.t1252 24.9236
R2640 GND.n5700 GND.t1218 24.9236
R2641 GND.n5706 GND.t1280 24.9236
R2642 GND.n5706 GND.t1310 24.9236
R2643 GND.n5712 GND.t1236 24.9236
R2644 GND.n5712 GND.t1262 24.9236
R2645 GND.n5724 GND.t1292 24.9236
R2646 GND.n5724 GND.t1194 24.9236
R2647 GND.n5730 GND.t1244 24.9236
R2648 GND.n5730 GND.t1212 24.9236
R2649 GND.n5750 GND.t1268 24.9236
R2650 GND.n5750 GND.t1300 24.9236
R2651 GND.n5745 GND.t1216 24.9236
R2652 GND.n5745 GND.t1272 24.9236
R2653 GND.n5738 GND.t1304 24.9236
R2654 GND.n5738 GND.t1230 24.9236
R2655 GND.n5653 GND.t1256 24.9236
R2656 GND.n5653 GND.t1288 24.9236
R2657 GND.n6142 GND.t1234 24.9236
R2658 GND.n6142 GND.t1260 24.9236
R2659 GND.n6155 GND.t336 24.9236
R2660 GND.n6155 GND.t346 24.9236
R2661 GND.n6165 GND.t356 24.9236
R2662 GND.n6165 GND.t334 24.9236
R2663 GND.n6172 GND.t348 24.9236
R2664 GND.n6172 GND.t358 24.9236
R2665 GND.n6176 GND.t338 24.9236
R2666 GND.n6176 GND.t344 24.9236
R2667 GND.n6182 GND.t354 24.9236
R2668 GND.n6182 GND.t350 24.9236
R2669 GND.n6188 GND.t332 24.9236
R2670 GND.n6188 GND.t342 24.9236
R2671 GND.n6195 GND.t352 24.9236
R2672 GND.n6195 GND.t328 24.9236
R2673 GND.n5662 GND.t1224 24.9236
R2674 GND.n5662 GND.t1296 24.9236
R2675 GND.n5670 GND.t1196 24.9236
R2676 GND.n5670 GND.t1246 24.9236
R2677 GND.n5676 GND.t1282 24.9236
R2678 GND.n5676 GND.t1200 24.9236
R2679 GND.n5680 GND.t1250 24.9236
R2680 GND.n5680 GND.t1286 24.9236
R2681 GND.n5846 GND.t1274 24.9236
R2682 GND.n5846 GND.t1308 24.9236
R2683 GND.n5840 GND.t1204 24.9236
R2684 GND.n5840 GND.t1278 24.9236
R2685 GND.n5834 GND.t1312 24.9236
R2686 GND.n5834 GND.t1238 24.9236
R2687 GND.n963 GND.t1053 24.9236
R2688 GND.n963 GND.t1047 24.9236
R2689 GND.n707 GND.t237 24.9236
R2690 GND.n707 GND.t217 24.9236
R2691 GND.n923 GND.t225 24.9236
R2692 GND.n923 GND.t235 24.9236
R2693 GND.n929 GND.t231 24.9236
R2694 GND.n929 GND.t239 24.9236
R2695 GND.n933 GND.t219 24.9236
R2696 GND.n933 GND.t233 24.9236
R2697 GND.n939 GND.t241 24.9236
R2698 GND.n939 GND.t221 24.9236
R2699 GND.n945 GND.t227 24.9236
R2700 GND.n945 GND.t211 24.9236
R2701 GND.n951 GND.t215 24.9236
R2702 GND.n951 GND.t229 24.9236
R2703 GND.n865 GND.t838 24.9236
R2704 GND.n865 GND.t736 24.9236
R2705 GND.n910 GND.t816 24.9236
R2706 GND.n910 GND.t842 24.9236
R2707 GND.n903 GND.t774 24.9236
R2708 GND.n903 GND.t796 24.9236
R2709 GND.n899 GND.t832 24.9236
R2710 GND.n899 GND.t764 24.9236
R2711 GND.n893 GND.t800 24.9236
R2712 GND.n893 GND.t742 24.9236
R2713 GND.n887 GND.t826 24.9236
R2714 GND.n887 GND.t724 24.9236
R2715 GND.n881 GND.t784 24.9236
R2716 GND.n881 GND.t808 24.9236
R2717 GND.n778 GND.t792 24.9236
R2718 GND.n778 GND.t822 24.9236
R2719 GND.n711 GND.t758 24.9236
R2720 GND.n711 GND.t844 24.9236
R2721 GND.n830 GND.t754 24.9236
R2722 GND.n830 GND.t818 24.9236
R2723 GND.n834 GND.t846 24.9236
R2724 GND.n834 GND.t776 24.9236
R2725 GND.n840 GND.t802 24.9236
R2726 GND.n840 GND.t824 24.9236
R2727 GND.n846 GND.t778 24.9236
R2728 GND.n846 GND.t804 24.9236
R2729 GND.n852 GND.t750 24.9236
R2730 GND.n852 GND.t772 24.9236
R2731 GND.n766 GND.t814 24.9236
R2732 GND.n766 GND.t840 24.9236
R2733 GND.n817 GND.t738 24.9236
R2734 GND.n817 GND.t794 24.9236
R2735 GND.n810 GND.t830 24.9236
R2736 GND.n810 GND.t760 24.9236
R2737 GND.n806 GND.t798 24.9236
R2738 GND.n806 GND.t834 24.9236
R2739 GND.n800 GND.t768 24.9236
R2740 GND.n800 GND.t720 24.9236
R2741 GND.n794 GND.t780 24.9236
R2742 GND.n794 GND.t806 24.9236
R2743 GND.n788 GND.t726 24.9236
R2744 GND.n788 GND.t786 24.9236
R2745 GND.n715 GND.t770 24.9236
R2746 GND.n715 GND.t728 24.9236
R2747 GND.n720 GND.t748 24.9236
R2748 GND.n720 GND.t740 24.9236
R2749 GND.n731 GND.t762 24.9236
R2750 GND.n731 GND.t788 24.9236
R2751 GND.n736 GND.t730 24.9236
R2752 GND.n736 GND.t766 24.9236
R2753 GND.n742 GND.t836 24.9236
R2754 GND.n742 GND.t732 24.9236
R2755 GND.n748 GND.t756 24.9236
R2756 GND.n748 GND.t820 24.9236
R2757 GND.n754 GND.t722 24.9236
R2758 GND.n754 GND.t782 24.9236
R2759 GND.n6089 GND.t1142 24.9236
R2760 GND.n6089 GND.t1136 24.9236
R2761 GND.n6041 GND.t43 24.9236
R2762 GND.n6041 GND.t55 24.9236
R2763 GND.n6049 GND.t63 24.9236
R2764 GND.n6049 GND.t41 24.9236
R2765 GND.n6055 GND.t37 24.9236
R2766 GND.n6055 GND.t45 24.9236
R2767 GND.n6059 GND.t57 24.9236
R2768 GND.n6059 GND.t39 24.9236
R2769 GND.n6065 GND.t47 24.9236
R2770 GND.n6065 GND.t59 24.9236
R2771 GND.n6071 GND.t33 24.9236
R2772 GND.n6071 GND.t49 24.9236
R2773 GND.n6077 GND.t53 24.9236
R2774 GND.n6077 GND.t35 24.9236
R2775 GND.n6127 GND.t924 24.9236
R2776 GND.n6127 GND.t950 24.9236
R2777 GND.n5855 GND.t902 24.9236
R2778 GND.n5855 GND.t928 24.9236
R2779 GND.n6007 GND.t988 24.9236
R2780 GND.n6007 GND.t1010 24.9236
R2781 GND.n6011 GND.t916 24.9236
R2782 GND.n6011 GND.t978 24.9236
R2783 GND.n6017 GND.t886 24.9236
R2784 GND.n6017 GND.t956 24.9236
R2785 GND.n6023 GND.t910 24.9236
R2786 GND.n6023 GND.t938 24.9236
R2787 GND.n6029 GND.t998 24.9236
R2788 GND.n6029 GND.t894 24.9236
R2789 GND.n5960 GND.t1006 24.9236
R2790 GND.n5960 GND.t908 24.9236
R2791 GND.n5967 GND.t972 24.9236
R2792 GND.n5967 GND.t930 24.9236
R2793 GND.n5993 GND.t968 24.9236
R2794 GND.n5993 GND.t904 24.9236
R2795 GND.n5989 GND.t932 24.9236
R2796 GND.n5989 GND.t990 24.9236
R2797 GND.n5983 GND.t888 24.9236
R2798 GND.n5983 GND.t920 24.9236
R2799 GND.n5977 GND.t992 24.9236
R2800 GND.n5977 GND.t890 24.9236
R2801 GND.n5971 GND.t964 24.9236
R2802 GND.n5971 GND.t986 24.9236
R2803 GND.n5876 GND.t900 24.9236
R2804 GND.n5876 GND.t926 24.9236
R2805 GND.n5919 GND.t952 24.9236
R2806 GND.n5919 GND.t1008 24.9236
R2807 GND.n5926 GND.t914 24.9236
R2808 GND.n5926 GND.t974 24.9236
R2809 GND.n5930 GND.t1012 24.9236
R2810 GND.n5930 GND.t918 24.9236
R2811 GND.n5936 GND.t982 24.9236
R2812 GND.n5936 GND.t934 24.9236
R2813 GND.n5942 GND.t994 24.9236
R2814 GND.n5942 GND.t892 24.9236
R2815 GND.n5948 GND.t940 24.9236
R2816 GND.n5948 GND.t1000 24.9236
R2817 GND.n5862 GND.t984 24.9236
R2818 GND.n5862 GND.t942 24.9236
R2819 GND.n5867 GND.t962 24.9236
R2820 GND.n5867 GND.t954 24.9236
R2821 GND.n5909 GND.t976 24.9236
R2822 GND.n5909 GND.t1002 24.9236
R2823 GND.n5904 GND.t944 24.9236
R2824 GND.n5904 GND.t980 24.9236
R2825 GND.n5898 GND.t922 24.9236
R2826 GND.n5898 GND.t946 24.9236
R2827 GND.n5892 GND.t970 24.9236
R2828 GND.n5892 GND.t906 24.9236
R2829 GND.n5886 GND.t936 24.9236
R2830 GND.n5886 GND.t996 24.9236
R2831 GND.n551 GND.n550 24.4711
R2832 GND.n37 GND.n28 24.4711
R2833 GND.n6364 GND.n6355 24.4711
R2834 GND.n6200 GND.n6199 24.4711
R2835 GND.n959 GND.n958 24.4711
R2836 GND.n657 GND.n653 24.4711
R2837 GND.n683 GND.n682 24.4711
R2838 GND.n6285 GND.n6281 24.4711
R2839 GND.n6247 GND.n6246 24.4711
R2840 GND.n6085 GND.n6084 24.4711
R2841 GND.t562 GND.n2855 23.9028
R2842 GND.t563 GND.n3939 23.9028
R2843 GND.t549 GND.n3831 23.9028
R2844 GND.t564 GND.n3508 23.9028
R2845 GND.t448 GND.n1960 23.9028
R2846 GND.t269 GND.n2069 23.9028
R2847 GND.t536 GND.n2435 23.9028
R2848 GND.t552 GND.n4688 23.9028
R2849 GND.n689 GND.n673 23.7181
R2850 GND.n6253 GND.n6237 23.7181
R2851 GND.n4765 GND.n4764 23.4245
R2852 GND.n3180 GND.n3179 23.4245
R2853 GND.n2915 GND.n2914 23.4245
R2854 GND.n2309 GND.n2308 23.4245
R2855 GND.n7713 GND.n7712 23.4245
R2856 GND.n1569 GND.n1568 23.4245
R2857 GND.n5406 GND.n5405 23.4245
R2858 GND.n3975 GND.n3974 23.4245
R2859 GND.n5267 GND.n5266 23.4245
R2860 GND.n3867 GND.n3866 23.4245
R2861 GND.n3544 GND.n3543 23.4245
R2862 GND.n1996 GND.n1995 23.4245
R2863 GND.n2087 GND.n2086 23.4245
R2864 GND.n2471 GND.n2470 23.4245
R2865 GND.n2806 GND.n2805 23.4245
R2866 GND.n4925 GND.n4924 23.4245
R2867 GND.n33 GND.n32 22.9652
R2868 GND.n6360 GND.n6359 22.9652
R2869 GND.n7776 GND.n7775 22.9652
R2870 GND.n652 GND.n648 22.9652
R2871 GND.n696 GND.n694 22.9652
R2872 GND.n701 GND.n700 22.9652
R2873 GND.n6309 GND.n6308 22.9652
R2874 GND.n6280 GND.n6276 22.9652
R2875 GND.n6260 GND.n6258 22.9652
R2876 GND.n6265 GND.n6264 22.9652
R2877 GND.n3308 GND.n3307 22.9087
R2878 GND.n3005 GND.n3004 22.9087
R2879 GND.n2579 GND.n2578 22.9087
R2880 GND.n7179 GND.n7178 22.9087
R2881 GND.n7016 GND.n7015 22.9087
R2882 GND.n6862 GND.n6861 22.9087
R2883 GND.n6708 GND.n6707 22.9087
R2884 GND.n6637 GND.n6636 22.9087
R2885 GND.n5589 GND.n5588 22.9087
R2886 GND.n1087 GND.n1086 22.9087
R2887 GND.n1208 GND.n1207 22.9087
R2888 GND.n3669 GND.n3668 22.9087
R2889 GND.n5066 GND.n5065 22.9087
R2890 GND.n461 GND.n460 22.9087
R2891 GND.n392 GND.n391 22.9087
R2892 GND.n288 GND.n287 22.9087
R2893 GND.t273 GND.n5231 22.765
R2894 GND.t568 GND.n5370 22.765
R2895 GND.t447 GND.n1533 22.765
R2896 GND.t1071 GND.n7677 22.765
R2897 GND.t270 GND.n2273 22.765
R2898 GND.t573 GND.n2744 22.765
R2899 GND.t1128 GND.n4889 22.765
R2900 GND.n3012 GND.n3011 22.5323
R2901 GND.n7196 GND.n7195 22.5323
R2902 GND.n2592 GND.n2591 22.5323
R2903 GND.n6884 GND.n6883 22.5323
R2904 GND.n6730 GND.n6729 22.5323
R2905 GND.n5079 GND.n5078 22.5323
R2906 GND.n7038 GND.n7037 22.5323
R2907 GND.t1433 GND.t1431 22.4359
R2908 GND.t1436 GND.t1433 22.4359
R2909 GND.t1438 GND.t1436 22.4359
R2910 GND.t1175 GND.t1173 22.4359
R2911 GND.t1178 GND.t1175 22.4359
R2912 GND.t1180 GND.t1178 22.4359
R2913 GND.t25 GND.t23 22.4359
R2914 GND.t28 GND.t25 22.4359
R2915 GND.t30 GND.t28 22.4359
R2916 GND.t1499 GND.t1501 22.4359
R2917 GND.t1501 GND.t1495 22.4359
R2918 GND.t1495 GND.t1497 22.4359
R2919 GND.t394 GND.t396 22.4359
R2920 GND.t396 GND.t399 22.4359
R2921 GND.t399 GND.t392 22.4359
R2922 GND.t671 GND.t1490 22.4359
R2923 GND.t1490 GND.t1089 22.4359
R2924 GND.t1089 GND.t449 22.4359
R2925 GND.t2 GND.t0 22.4359
R2926 GND.t0 GND.t1321 22.4359
R2927 GND.t1321 GND.t1319 22.4359
R2928 GND.n253 GND.n252 22.4086
R2929 GND.n357 GND.n356 22.4086
R2930 GND.n426 GND.n425 22.4086
R2931 GND.n5031 GND.n5030 22.4086
R2932 GND.n1173 GND.n1172 22.4086
R2933 GND.n1052 GND.n1051 22.4086
R2934 GND.n5554 GND.n5553 22.4086
R2935 GND.n6602 GND.n6601 22.4086
R2936 GND.n6673 GND.n6672 22.4086
R2937 GND.n39 GND.t366 22.3257
R2938 GND.n6366 GND.t546 22.3257
R2939 GND.n6481 GND.t483 22.3257
R2940 GND.n6483 GND.t388 22.3257
R2941 GND.n654 GND.t1024 22.3257
R2942 GND.n645 GND.t1505 22.3257
R2943 GND.n679 GND.t591 22.3257
R2944 GND.n6391 GND.t614 22.3257
R2945 GND.n6393 GND.t1184 22.3257
R2946 GND.n6282 GND.t717 22.3257
R2947 GND.n6273 GND.t580 22.3257
R2948 GND.n6243 GND.t670 22.3257
R2949 GND.n688 GND.n676 22.2123
R2950 GND.n684 GND.n676 22.2123
R2951 GND.n6252 GND.n6240 22.2123
R2952 GND.n6248 GND.n6240 22.2123
R2953 GND GND.t365 22.1322
R2954 GND.n3035 GND.n3034 22.0429
R2955 GND.n246 GND.n245 22.0429
R2956 GND.n7653 GND.n7652 22.0429
R2957 GND.n7213 GND.n7212 22.0429
R2958 GND.n2609 GND.n2608 22.0429
R2959 GND.n6901 GND.n6900 22.0429
R2960 GND.n6747 GND.n6746 22.0429
R2961 GND.n6588 GND.n6587 22.0429
R2962 GND.n1045 GND.n1044 22.0429
R2963 GND.n3696 GND.n3695 22.0429
R2964 GND.n350 GND.n349 22.0429
R2965 GND.n488 GND.n487 22.0429
R2966 GND.n5096 GND.n5095 22.0429
R2967 GND.n1168 GND.n1167 22.0429
R2968 GND.n5540 GND.n5539 22.0429
R2969 GND.n7055 GND.n7054 22.0429
R2970 GND.n3238 GND.n3237 21.8358
R2971 GND.n7541 GND.n7540 21.8358
R2972 GND.n7603 GND.n7602 21.8358
R2973 GND.n2502 GND.n2501 21.8358
R2974 GND.n2919 GND.n2918 21.8358
R2975 GND.n6941 GND.n6940 21.8358
R2976 GND.n6778 GND.n6777 21.8358
R2977 GND.n67 GND.n66 21.8358
R2978 GND.n1011 GND.n1010 21.8358
R2979 GND.n1240 GND.n1239 21.8358
R2980 GND.n7479 GND.n7478 21.8358
R2981 GND.n4978 GND.n4977 21.8358
R2982 GND.n3584 GND.n3583 21.8358
R2983 GND.n1110 GND.n1109 21.8358
R2984 GND.n6532 GND.n6531 21.8358
R2985 GND.n7110 GND.n7109 21.8358
R2986 GND.n48 GND.n46 21.4593
R2987 GND.n6375 GND.n6373 21.4593
R2988 GND.n15 GND.n13 21.4593
R2989 GND.n17 GND.n10 21.4593
R2990 GND.n7783 GND.n7781 21.4593
R2991 GND.n7785 GND.n7768 21.4593
R2992 GND.n697 GND.n696 21.4593
R2993 GND.n700 GND.n699 21.4593
R2994 GND.n6340 GND.n6338 21.4593
R2995 GND.n6342 GND.n6335 21.4593
R2996 GND.n6316 GND.n6314 21.4593
R2997 GND.n6318 GND.n6301 21.4593
R2998 GND.n6261 GND.n6260 21.4593
R2999 GND.n6264 GND.n6263 21.4593
R3000 GND.n7805 GND.n7804 21.3675
R3001 GND.n3229 GND.n3228 20.6255
R3002 GND.n2886 GND.n2881 20.6255
R3003 GND.n2486 GND.n2485 20.6255
R3004 GND.n2018 GND.n2017 20.6255
R3005 GND.n3559 GND.n3558 20.6255
R3006 GND.n3886 GND.n3885 20.6255
R3007 GND.n3998 GND.n3997 20.6255
R3008 GND.n5294 GND.n5289 20.6255
R3009 GND.n5429 GND.n5424 20.6255
R3010 GND.n1589 GND.n1584 20.6255
R3011 GND.n7733 GND.n7728 20.6255
R3012 GND.n2330 GND.n2325 20.6255
R3013 GND.n2780 GND.n2779 20.6255
R3014 GND.n4941 GND.n4936 20.6255
R3015 GND.n4734 GND.n4733 20.6255
R3016 GND.n4791 GND.n4770 20.0775
R3017 GND.n33 GND.n28 19.9534
R3018 GND.n6360 GND.n6355 19.9534
R3019 GND.n7777 GND.n7776 19.9534
R3020 GND.n653 GND.n652 19.9534
R3021 GND.n694 GND.n669 19.9534
R3022 GND.n702 GND.n701 19.9534
R3023 GND.n6310 GND.n6309 19.9534
R3024 GND.n6281 GND.n6280 19.9534
R3025 GND.n6258 GND.n6233 19.9534
R3026 GND.n6266 GND.n6265 19.9534
R3027 GND.t69 GND.t505 19.2425
R3028 GND.t687 GND.t319 19.2425
R3029 GND.n4677 GND.n4676 19.2005
R3030 GND.n3372 GND.n3371 17.9597
R3031 GND.n7562 GND.t558 17.475
R3032 GND.n7624 GND.t685 17.475
R3033 GND.n2529 GND.t364 17.475
R3034 GND.n2952 GND.t1168 17.475
R3035 GND.n6961 GND.t1412 17.475
R3036 GND.n6798 GND.t360 17.475
R3037 GND.n6661 GND.t1387 17.475
R3038 GND.n5623 GND.t266 17.475
R3039 GND.n1276 GND.t882 17.475
R3040 GND.n7500 GND.t1425 17.475
R3041 GND.n5011 GND.t544 17.475
R3042 GND.n3617 GND.t249 17.475
R3043 GND.n5488 GND.t314 17.475
R3044 GND.n6553 GND.t262 17.475
R3045 GND.n7131 GND.t854 17.475
R3046 GND.n3260 GND.t1153 17.475
R3047 GND.n4850 GND.t303 17.4601
R3048 GND.n4643 GND.t1130 17.4601
R3049 GND.n2657 GND.t570 17.4601
R3050 GND.n3100 GND.t534 17.4601
R3051 GND.n3389 GND.t644 17.4601
R3052 GND.n2234 GND.t1144 17.4601
R3053 GND.n2172 GND.t566 17.4601
R3054 GND.n144 GND.t301 17.4601
R3055 GND.n1495 GND.t646 17.4601
R3056 GND.n1327 GND.t572 17.4601
R3057 GND.n4023 GND.t560 17.4601
R3058 GND.n5193 GND.t551 17.4601
R3059 GND.n3792 GND.t1134 17.4601
R3060 GND.n3470 GND.t272 17.4601
R3061 GND.n1921 GND.t1146 17.4601
R3062 GND.n2397 GND.t1132 17.4601
R3063 GND.n7562 GND.t1088 17.4528
R3064 GND.n7624 GND.t638 17.4528
R3065 GND.n2529 GND.t1521 17.4528
R3066 GND.n2952 GND.t662 17.4528
R3067 GND.n6961 GND.t1344 17.4528
R3068 GND.n6798 GND.t496 17.4528
R3069 GND.n6661 GND.t246 17.4528
R3070 GND.n5623 GND.t457 17.4528
R3071 GND.n1276 GND.t419 17.4528
R3072 GND.n7500 GND.t1397 17.4528
R3073 GND.n5011 GND.t870 17.4528
R3074 GND.n3617 GND.t1536 17.4528
R3075 GND.n5488 GND.t260 17.4528
R3076 GND.n6553 GND.t1022 17.4528
R3077 GND.n7131 GND.t1170 17.4528
R3078 GND.n3260 GND.t1116 17.4528
R3079 GND.n192 GND.n191 17.2882
R3080 GND.n6002 GND.t929 17.2168
R3081 GND.t1376 GND 17.1372
R3082 GND.t1428 GND 17.1372
R3083 GND.t883 GND 17.1372
R3084 GND.n583 GND.n582 16.9417
R3085 GND.n7409 GND.n7408 16.9417
R3086 GND.n7362 GND.n7361 16.9417
R3087 GND.n7303 GND.n7302 16.9417
R3088 GND.n7277 GND.n7276 16.9417
R3089 GND.n5805 GND.n5804 16.9417
R3090 GND.n5693 GND.n5692 16.9417
R3091 GND.n5747 GND.n5746 16.9417
R3092 GND.n6178 GND.n6177 16.9417
R3093 GND.n5682 GND.n5681 16.9417
R3094 GND.n935 GND.n934 16.9417
R3095 GND.n901 GND.n900 16.9417
R3096 GND.n836 GND.n835 16.9417
R3097 GND.n808 GND.n807 16.9417
R3098 GND.n738 GND.n737 16.9417
R3099 GND.n697 GND.n693 16.9417
R3100 GND.n699 GND.n673 16.9417
R3101 GND.n6261 GND.n6257 16.9417
R3102 GND.n6263 GND.n6237 16.9417
R3103 GND.n6061 GND.n6060 16.9417
R3104 GND.n6013 GND.n6012 16.9417
R3105 GND.n5991 GND.n5990 16.9417
R3106 GND.n5932 GND.n5931 16.9417
R3107 GND.n5906 GND.n5905 16.9417
R3108 GND.t541 GND 16.9356
R3109 GND.t1163 GND.t379 16.8628
R3110 GND GND.t1163 16.2041
R3111 GND.n3326 GND.n3325 16.1887
R3112 GND.n7513 GND.n7512 16.1887
R3113 GND.n7575 GND.n7574 16.1887
R3114 GND.n2629 GND.n2628 16.1887
R3115 GND.n3055 GND.n3054 16.1887
R3116 GND.n6976 GND.n6925 16.1887
R3117 GND.n6822 GND.n6771 16.1887
R3118 GND.n7758 GND.n51 16.1887
R3119 GND.n5638 GND.n995 16.1887
R3120 GND.n5454 GND.n1224 16.1887
R3121 GND.n7451 GND.n7450 16.1887
R3122 GND.n5116 GND.n5115 16.1887
R3123 GND.n3716 GND.n3715 16.1887
R3124 GND.n5511 GND.n1103 16.1887
R3125 GND.n6504 GND.n6503 16.1887
R3126 GND.n7082 GND.n7081 16.1887
R3127 GND.n684 GND.n683 16.1887
R3128 GND.n6248 GND.n6247 16.1887
R3129 GND.n3979 GND.n3978 14.7755
R3130 GND.n4928 GND.n4926 14.7755
R3131 GND.n4719 GND.n4718 14.7755
R3132 GND.n4708 GND.n4703 14.7755
R3133 GND.n3187 GND.n3186 14.7755
R3134 GND.n3183 GND.n3181 14.7755
R3135 GND.n2865 GND.n2863 14.7755
R3136 GND.n2873 GND.n2868 14.7755
R3137 GND.n2762 GND.n2760 14.7755
R3138 GND.n2315 GND.n2310 14.7755
R3139 GND.n2090 GND.n2089 14.7755
R3140 GND.n118 GND.n116 14.7755
R3141 GND.n7720 GND.n7715 14.7755
R3142 GND.n7718 GND.n7716 14.7755
R3143 GND.n2001 GND.n1999 14.7755
R3144 GND.n1576 GND.n1571 14.7755
R3145 GND.n1574 GND.n1572 14.7755
R3146 GND.n5412 GND.n5407 14.7755
R3147 GND.n5416 GND.n5415 14.7755
R3148 GND.n3870 GND.n3868 14.7755
R3149 GND.n5279 GND.n5277 14.7755
R3150 GND.n3982 GND.n3981 14.7755
R3151 GND.n5273 GND.n5268 14.7755
R3152 GND.n5281 GND.n5276 14.7755
R3153 GND.n5271 GND.n5269 14.7755
R3154 GND.n5410 GND.n5408 14.7755
R3155 GND.n2003 GND.n1998 14.7755
R3156 GND.n2092 GND.n2088 14.7755
R3157 GND.n120 GND.n115 14.7755
R3158 GND.n2313 GND.n2311 14.7755
R3159 GND.n2871 GND.n2869 14.7755
R3160 GND.n2764 GND.n2759 14.7755
R3161 GND.t387 GND.t482 14.6672
R3162 GND.t1539 GND.t553 14.6672
R3163 GND.t386 GND.t378 14.6672
R3164 GND.t613 GND.t1183 14.6672
R3165 GND.t682 GND.t1549 14.6672
R3166 GND.t699 GND.t692 14.6672
R3167 GND.n7807 GND.n3 14.5711
R3168 GND.n992 GND.n968 14.5711
R3169 GND.n6118 GND.n6094 14.5711
R3170 GND.t535 GND.n4674 14.4569
R3171 GND.n824 GND.t843 14.2308
R3172 GND.t365 GND.t600 14.228
R3173 GND.n7375 GND.t167 13.8225
R3174 GND.n6485 GND.n6482 13.5727
R3175 GND.n6395 GND.n6392 13.5727
R3176 GND.n6485 GND.n6484 13.5705
R3177 GND.n6395 GND.n6394 13.5705
R3178 GND.n660 GND.n659 13.5646
R3179 GND.n6288 GND.n6287 13.5646
R3180 GND.n4255 GND.n4254 13.4405
R3181 GND.n5696 GND.t1305 13.4015
R3182 GND.n7796 GND.n7761 13.3549
R3183 GND.t377 GND 13.3059
R3184 GND.t443 GND.t507 12.9107
R3185 GND.t1122 GND.t603 12.6472
R3186 GND.n3386 GND.t643 12.5719
R3187 GND GND.t1074 12.5248
R3188 GND GND.t1334 12.5248
R3189 GND GND.t871 12.5248
R3190 GND GND.t1483 12.5248
R3191 GND GND.t466 12.5248
R3192 GND.t411 GND 12.5248
R3193 GND.t1374 GND 12.5248
R3194 GND.t517 GND 12.5248
R3195 GND GND.t1325 12.5248
R3196 GND.t296 GND.n1746 11.89
R3197 GND.n5321 GND.t296 11.89
R3198 GND.t497 GND.n4068 11.89
R3199 GND.t430 GND.n4430 11.89
R3200 GND.t1314 GND.n4414 11.89
R3201 GND.t1038 GND.n4399 11.89
R3202 GND.t1318 GND.n4384 11.89
R3203 GND.t1035 GND.n4369 11.89
R3204 GND.t428 GND.n4352 11.89
R3205 GND.t1313 GND.n4337 11.89
R3206 GND.t1037 GND.n4322 11.89
R3207 GND.t1317 GND.n4307 11.89
R3208 GND.t431 GND.n4290 11.89
R3209 GND.t1565 GND.n4270 11.89
R3210 GND.t1315 GND.n4228 11.89
R3211 GND.t1034 GND.n4213 11.89
R3212 GND.t1567 GND.n4198 11.89
R3213 GND.t433 GND.n4183 11.89
R3214 GND.t1316 GND.n4164 11.89
R3215 GND.t1569 GND.n4149 11.89
R3216 GND.t429 GND.n4134 11.89
R3217 GND.t1036 GND.n4119 11.89
R3218 GND.n587 GND.n586 11.6711
R3219 GND.n7413 GND.n7412 11.6711
R3220 GND.n7366 GND.n7365 11.6711
R3221 GND.n7299 GND.n7298 11.6711
R3222 GND.n7282 GND.n7281 11.6711
R3223 GND.n5809 GND.n5808 11.6711
R3224 GND.n5762 GND.n5761 11.6711
R3225 GND.n5752 GND.n5751 11.6711
R3226 GND.n6174 GND.n6173 11.6711
R3227 GND.n5678 GND.n5677 11.6711
R3228 GND.n931 GND.n930 11.6711
R3229 GND.n905 GND.n904 11.6711
R3230 GND.n832 GND.n831 11.6711
R3231 GND.n812 GND.n811 11.6711
R3232 GND.n733 GND.n732 11.6711
R3233 GND.n6057 GND.n6056 11.6711
R3234 GND.n6009 GND.n6008 11.6711
R3235 GND.n5995 GND.n5994 11.6711
R3236 GND.n5928 GND.n5927 11.6711
R3237 GND.n5911 GND.n5910 11.6711
R3238 GND.t1568 GND.n4243 11.48
R3239 GND.n6206 GND.n6205 11.427
R3240 GND.n6204 GND.n6203 11.427
R3241 GND.n6428 GND.n6427 11.427
R3242 GND.n513 GND.n512 11.427
R3243 GND.t507 GND.t651 11.0664
R3244 GND.t651 GND.t1122 11.0664
R3245 GND.t600 GND.t377 11.0664
R3246 GND.t1431 GND 10.9511
R3247 GND.t1173 GND 10.9511
R3248 GND.t23 GND 10.9511
R3249 GND GND.t1499 10.9511
R3250 GND GND.t394 10.9511
R3251 GND GND.t671 10.9511
R3252 GND GND.t2 10.9511
R3253 GND.n577 GND.n576 10.9181
R3254 GND.n7403 GND.n7402 10.9181
R3255 GND.n7356 GND.n7355 10.9181
R3256 GND.n7309 GND.n7308 10.9181
R3257 GND.n7271 GND.n7270 10.9181
R3258 GND.n5799 GND.n5798 10.9181
R3259 GND.n5702 GND.n5701 10.9181
R3260 GND.n5740 GND.n5739 10.9181
R3261 GND.n6184 GND.n6183 10.9181
R3262 GND.n5848 GND.n5847 10.9181
R3263 GND.n941 GND.n940 10.9181
R3264 GND.n895 GND.n894 10.9181
R3265 GND.n842 GND.n841 10.9181
R3266 GND.n802 GND.n801 10.9181
R3267 GND.n744 GND.n743 10.9181
R3268 GND.n6067 GND.n6066 10.9181
R3269 GND.n6019 GND.n6018 10.9181
R3270 GND.n5985 GND.n5984 10.9181
R3271 GND.n5938 GND.n5937 10.9181
R3272 GND.n5900 GND.n5899 10.9181
R3273 GND.n4581 GND.n4578 10.7897
R3274 GND GND.t693 10.6857
R3275 GND GND.t1376 10.6857
R3276 GND GND.t1428 10.6857
R3277 GND GND.t541 10.6857
R3278 GND GND.t883 10.6857
R3279 GND.n6207 GND.n6206 10.5417
R3280 GND GND.n7230 10.1442
R3281 GND.n3091 GND.n3088 9.8307
R3282 GND.t1361 GND.t1161 9.8307
R3283 GND.n3108 GND.n3105 9.8307
R3284 GND.n4014 GND.n4011 9.8307
R3285 GND.t1390 GND.t678 9.8307
R3286 GND.n4031 GND.n4028 9.8307
R3287 GND.n5153 GND.n5150 9.8307
R3288 GND.t389 GND.t1395 9.8307
R3289 GND.n5186 GND.n5183 9.8307
R3290 GND.n3752 GND.n3749 9.8307
R3291 GND.t1519 GND.t522 9.8307
R3292 GND.n3785 GND.n3782 9.8307
R3293 GND.n1287 GND.n1284 9.8307
R3294 GND.t292 GND.t304 9.8307
R3295 GND.n1320 GND.n1317 9.8307
R3296 GND.n3430 GND.n3427 9.8307
R3297 GND.t855 GND.t574 9.8307
R3298 GND.n3463 GND.n3460 9.8307
R3299 GND.n1455 GND.n1452 9.8307
R3300 GND.t641 GND.t1419 9.8307
R3301 GND.n1488 GND.n1485 9.8307
R3302 GND.n1881 GND.n1878 9.8307
R3303 GND.t254 GND.t427 9.8307
R3304 GND.n1914 GND.n1911 9.8307
R3305 GND.n96 GND.n95 9.8307
R3306 GND.t274 GND.t326 9.8307
R3307 GND.n137 GND.n134 9.8307
R3308 GND.n2132 GND.n2129 9.8307
R3309 GND.t277 GND.t1415 9.8307
R3310 GND.n2165 GND.n2162 9.8307
R3311 GND.n2194 GND.n2191 9.8307
R3312 GND.t1124 GND.t442 9.8307
R3313 GND.n2227 GND.n2224 9.8307
R3314 GND.n2357 GND.n2356 9.8307
R3315 GND.t1379 GND.t1041 9.8307
R3316 GND.n2390 GND.n2387 9.8307
R3317 GND.n2669 GND.n2666 9.8307
R3318 GND.t861 GND.t667 9.8307
R3319 GND.n2684 GND.n2681 9.8307
R3320 GND.n4810 GND.n4807 9.8307
R3321 GND.t1069 GND.t253 9.8307
R3322 GND.n4843 GND.n4840 9.8307
R3323 GND.n4603 GND.n4600 9.8307
R3324 GND.t258 GND.t307 9.8307
R3325 GND.n4636 GND.n4633 9.8307
R3326 GND.t379 GND.t1557 9.48553
R3327 GND.t1557 GND.t1384 9.48553
R3328 GND.n40 GND.n38 9.41227
R3329 GND.n6367 GND.n6365 9.41227
R3330 GND.n656 GND.n655 9.41227
R3331 GND.n6284 GND.n6283 9.41227
R3332 GND.n3252 GND.n3251 9.3005
R3333 GND.n3239 GND.n3238 9.3005
R3334 GND.n3241 GND.n3240 9.3005
R3335 GND.n3254 GND.n3253 9.3005
R3336 GND.n3339 GND.n3338 9.3005
R3337 GND.n3327 GND.n3326 9.3005
R3338 GND.n7555 GND.n7554 9.3005
R3339 GND.n7542 GND.n7541 9.3005
R3340 GND.n7544 GND.n7543 9.3005
R3341 GND.n7557 GND.n7556 9.3005
R3342 GND.n7526 GND.n7525 9.3005
R3343 GND.n7514 GND.n7513 9.3005
R3344 GND.n233 GND.n232 9.3005
R3345 GND.n353 GND.n352 9.3005
R3346 GND.n244 GND.n243 9.3005
R3347 GND.n235 GND.n234 9.3005
R3348 GND.n247 GND.n246 9.3005
R3349 GND.n300 GND.n299 9.3005
R3350 GND.n7567 GND.n7566 9.3005
R3351 GND.n302 GND.n301 9.3005
R3352 GND.n7617 GND.n7616 9.3005
R3353 GND.n7604 GND.n7603 9.3005
R3354 GND.n7606 GND.n7605 9.3005
R3355 GND.n7619 GND.n7618 9.3005
R3356 GND.n7588 GND.n7587 9.3005
R3357 GND.n7576 GND.n7575 9.3005
R3358 GND.n7640 GND.n7639 9.3005
R3359 GND.n249 GND.n248 9.3005
R3360 GND.n7651 GND.n7650 9.3005
R3361 GND.n7642 GND.n7641 9.3005
R3362 GND.n7654 GND.n7653 9.3005
R3363 GND.n7631 GND.n7630 9.3005
R3364 GND.n200 GND.n199 9.3005
R3365 GND.n7629 GND.n7628 9.3005
R3366 GND.n2513 GND.n2512 9.3005
R3367 GND.n2503 GND.n2502 9.3005
R3368 GND.n2505 GND.n2504 9.3005
R3369 GND.n2515 GND.n2514 9.3005
R3370 GND.n2642 GND.n2641 9.3005
R3371 GND.n2630 GND.n2629 9.3005
R3372 GND.n7200 GND.n7199 9.3005
R3373 GND.n7197 GND.n7196 9.3005
R3374 GND.n7211 GND.n7210 9.3005
R3375 GND.n7202 GND.n7201 9.3005
R3376 GND.n7214 GND.n7213 9.3005
R3377 GND.n7184 GND.n7183 9.3005
R3378 GND.n7135 GND.n7134 9.3005
R3379 GND.n2525 GND.n2524 9.3005
R3380 GND.n2930 GND.n2929 9.3005
R3381 GND.n2920 GND.n2919 9.3005
R3382 GND.n2922 GND.n2921 9.3005
R3383 GND.n2932 GND.n2931 9.3005
R3384 GND.n3068 GND.n3067 9.3005
R3385 GND.n3056 GND.n3055 9.3005
R3386 GND.n2596 GND.n2595 9.3005
R3387 GND.n2593 GND.n2592 9.3005
R3388 GND.n2607 GND.n2606 9.3005
R3389 GND.n2598 GND.n2597 9.3005
R3390 GND.n2610 GND.n2609 9.3005
R3391 GND.n2942 GND.n2941 9.3005
R3392 GND.n2949 GND.n2948 9.3005
R3393 GND.n2944 GND.n2943 9.3005
R3394 GND.n3231 GND.n3230 9.3005
R3395 GND.n3230 GND.n3229 9.3005
R3396 GND.n2890 GND.n2889 9.3005
R3397 GND.n6956 GND.n6955 9.3005
R3398 GND.n6942 GND.n6941 9.3005
R3399 GND.n6944 GND.n6943 9.3005
R3400 GND.n6934 GND.n6933 9.3005
R3401 GND.n6977 GND.n6976 9.3005
R3402 GND.n6888 GND.n6887 9.3005
R3403 GND.n6885 GND.n6884 9.3005
R3404 GND.n6899 GND.n6898 9.3005
R3405 GND.n6890 GND.n6889 9.3005
R3406 GND.n6902 GND.n6901 9.3005
R3407 GND.n6867 GND.n6866 9.3005
R3408 GND.n611 GND.n610 9.3005
R3409 GND.n6920 GND.n6919 9.3005
R3410 GND.n6792 GND.n6791 9.3005
R3411 GND.n6779 GND.n6778 9.3005
R3412 GND.n6781 GND.n6780 9.3005
R3413 GND.n6794 GND.n6793 9.3005
R3414 GND.n6811 GND.n6810 9.3005
R3415 GND.n6823 GND.n6822 9.3005
R3416 GND.n6734 GND.n6733 9.3005
R3417 GND.n6731 GND.n6730 9.3005
R3418 GND.n6745 GND.n6744 9.3005
R3419 GND.n6736 GND.n6735 9.3005
R3420 GND.n6748 GND.n6747 9.3005
R3421 GND.n6713 GND.n6712 9.3005
R3422 GND.n621 GND.n620 9.3005
R3423 GND.n6766 GND.n6765 9.3005
R3424 GND.n82 GND.n81 9.3005
R3425 GND.n68 GND.n67 9.3005
R3426 GND.n70 GND.n69 9.3005
R3427 GND.n59 GND.n58 9.3005
R3428 GND.n7759 GND.n7758 9.3005
R3429 GND.n6575 GND.n6574 9.3005
R3430 GND.n6572 GND.n6571 9.3005
R3431 GND.n6586 GND.n6585 9.3005
R3432 GND.n6577 GND.n6576 9.3005
R3433 GND.n6589 GND.n6588 9.3005
R3434 GND.n6649 GND.n6648 9.3005
R3435 GND.n6658 GND.n6657 9.3005
R3436 GND.n6651 GND.n6650 9.3005
R3437 GND.n1025 GND.n1024 9.3005
R3438 GND.n1012 GND.n1011 9.3005
R3439 GND.n1014 GND.n1013 9.3005
R3440 GND.n1027 GND.n1026 9.3005
R3441 GND.n1004 GND.n1003 9.3005
R3442 GND.n5639 GND.n5638 9.3005
R3443 GND.n1032 GND.n1031 9.3005
R3444 GND.n5550 GND.n5549 9.3005
R3445 GND.n1043 GND.n1042 9.3005
R3446 GND.n1034 GND.n1033 9.3005
R3447 GND.n1046 GND.n1045 9.3005
R3448 GND.n1099 GND.n1098 9.3005
R3449 GND.n5520 GND.n5519 9.3005
R3450 GND.n1101 GND.n1100 9.3005
R3451 GND.n1252 GND.n1251 9.3005
R3452 GND.n1241 GND.n1240 9.3005
R3453 GND.n1243 GND.n1242 9.3005
R3454 GND.n1233 GND.n1232 9.3005
R3455 GND.n5455 GND.n5454 9.3005
R3456 GND.n3683 GND.n3682 9.3005
R3457 GND.n3680 GND.n3679 9.3005
R3458 GND.n3694 GND.n3693 9.3005
R3459 GND.n3685 GND.n3684 9.3005
R3460 GND.n3697 GND.n3696 9.3005
R3461 GND.n1261 GND.n1260 9.3005
R3462 GND.n1268 GND.n1267 9.3005
R3463 GND.n1263 GND.n1262 9.3005
R3464 GND.n4000 GND.n3999 9.3005
R3465 GND.n3999 GND.n3998 9.3005
R3466 GND.n7494 GND.n7493 9.3005
R3467 GND.n7480 GND.n7479 9.3005
R3468 GND.n7482 GND.n7481 9.3005
R3469 GND.n7464 GND.n7463 9.3005
R3470 GND.n7452 GND.n7451 9.3005
R3471 GND.n337 GND.n336 9.3005
R3472 GND.n334 GND.n333 9.3005
R3473 GND.n348 GND.n347 9.3005
R3474 GND.n339 GND.n338 9.3005
R3475 GND.n351 GND.n350 9.3005
R3476 GND.n404 GND.n403 9.3005
R3477 GND.n7505 GND.n7504 9.3005
R3478 GND.n406 GND.n405 9.3005
R3479 GND.n4993 GND.n4992 9.3005
R3480 GND.n4979 GND.n4978 9.3005
R3481 GND.n4981 GND.n4980 9.3005
R3482 GND.n5129 GND.n5128 9.3005
R3483 GND.n5117 GND.n5116 9.3005
R3484 GND.n475 GND.n474 9.3005
R3485 GND.n472 GND.n471 9.3005
R3486 GND.n486 GND.n485 9.3005
R3487 GND.n477 GND.n476 9.3005
R3488 GND.n489 GND.n488 9.3005
R3489 GND.n5001 GND.n5000 9.3005
R3490 GND.n5008 GND.n5007 9.3005
R3491 GND.n5003 GND.n5002 9.3005
R3492 GND.n5298 GND.n5297 9.3005
R3493 GND.n3595 GND.n3594 9.3005
R3494 GND.n3585 GND.n3584 9.3005
R3495 GND.n3587 GND.n3586 9.3005
R3496 GND.n3597 GND.n3596 9.3005
R3497 GND.n3729 GND.n3728 9.3005
R3498 GND.n3717 GND.n3716 9.3005
R3499 GND.n5083 GND.n5082 9.3005
R3500 GND.n5080 GND.n5079 9.3005
R3501 GND.n5094 GND.n5093 9.3005
R3502 GND.n5085 GND.n5084 9.3005
R3503 GND.n5097 GND.n5096 9.3005
R3504 GND.n3607 GND.n3606 9.3005
R3505 GND.n3614 GND.n3613 9.3005
R3506 GND.n3609 GND.n3608 9.3005
R3507 GND.n3888 GND.n3887 9.3005
R3508 GND.n3887 GND.n3886 9.3005
R3509 GND.n5433 GND.n5432 9.3005
R3510 GND.n1124 GND.n1123 9.3005
R3511 GND.n1111 GND.n1110 9.3005
R3512 GND.n1113 GND.n1112 9.3005
R3513 GND.n1126 GND.n1125 9.3005
R3514 GND.n5500 GND.n5499 9.3005
R3515 GND.n5512 GND.n5511 9.3005
R3516 GND.n1155 GND.n1154 9.3005
R3517 GND.n1048 GND.n1047 9.3005
R3518 GND.n1166 GND.n1165 9.3005
R3519 GND.n1157 GND.n1156 9.3005
R3520 GND.n1169 GND.n1168 9.3005
R3521 GND.n1220 GND.n1219 9.3005
R3522 GND.n5463 GND.n5462 9.3005
R3523 GND.n1222 GND.n1221 9.3005
R3524 GND.n3561 GND.n3560 9.3005
R3525 GND.n3560 GND.n3559 9.3005
R3526 GND.n1593 GND.n1592 9.3005
R3527 GND.n6546 GND.n6545 9.3005
R3528 GND.n6533 GND.n6532 9.3005
R3529 GND.n6535 GND.n6534 9.3005
R3530 GND.n6548 GND.n6547 9.3005
R3531 GND.n6521 GND.n6520 9.3005
R3532 GND.n6505 GND.n6504 9.3005
R3533 GND.n5527 GND.n5526 9.3005
R3534 GND.n6598 GND.n6597 9.3005
R3535 GND.n5538 GND.n5537 9.3005
R3536 GND.n5529 GND.n5528 9.3005
R3537 GND.n5541 GND.n5540 9.3005
R3538 GND.n5601 GND.n5600 9.3005
R3539 GND.n5644 GND.n5643 9.3005
R3540 GND.n5603 GND.n5602 9.3005
R3541 GND.n2020 GND.n2019 9.3005
R3542 GND.n2019 GND.n2018 9.3005
R3543 GND.n7737 GND.n7736 9.3005
R3544 GND.n2118 GND.n2117 9.3005
R3545 GND.n2117 GND.n2116 9.3005
R3546 GND.n2334 GND.n2333 9.3005
R3547 GND.n7124 GND.n7123 9.3005
R3548 GND.n7111 GND.n7110 9.3005
R3549 GND.n7113 GND.n7112 9.3005
R3550 GND.n7126 GND.n7125 9.3005
R3551 GND.n7095 GND.n7094 9.3005
R3552 GND.n7083 GND.n7082 9.3005
R3553 GND.n7042 GND.n7041 9.3005
R3554 GND.n7039 GND.n7038 9.3005
R3555 GND.n7053 GND.n7052 9.3005
R3556 GND.n7044 GND.n7043 9.3005
R3557 GND.n7056 GND.n7055 9.3005
R3558 GND.n7021 GND.n7020 9.3005
R3559 GND.n601 GND.n600 9.3005
R3560 GND.n7074 GND.n7073 9.3005
R3561 GND.n2488 GND.n2487 9.3005
R3562 GND.n2487 GND.n2486 9.3005
R3563 GND.n2782 GND.n2781 9.3005
R3564 GND.n2781 GND.n2780 9.3005
R3565 GND.n4945 GND.n4944 9.3005
R3566 GND.n4179 GND.n4178 9.3005
R3567 GND.n4091 GND.n4090 9.3005
R3568 GND.n4593 GND.n4592 9.3005
R3569 GND.n4366 GND.n4365 9.3005
R3570 GND.n4456 GND.n4455 9.3005
R3571 GND.n4736 GND.n4735 9.3005
R3572 GND.n4735 GND.n4734 9.3005
R3573 GND.n3269 GND.n3268 9.3005
R3574 GND.n3264 GND.n3263 9.3005
R3575 GND.n3036 GND.n3035 9.3005
R3576 GND.n3262 GND.n3261 9.3005
R3577 GND.n3033 GND.n3032 9.3005
R3578 GND.n3024 GND.n3023 9.3005
R3579 GND.n3022 GND.n3021 9.3005
R3580 GND.n3013 GND.n3012 9.3005
R3581 GND.n3277 GND.n3276 9.3005
R3582 GND.n3319 GND.n3318 9.3005
R3583 GND.n3309 GND.n3308 9.3005
R3584 GND.n3288 GND.n3287 9.3005
R3585 GND.n3297 GND.n3296 9.3005
R3586 GND.n3279 GND.n3278 9.3005
R3587 GND.n3286 GND.n3285 9.3005
R3588 GND.n2969 GND.n2968 9.3005
R3589 GND.n3047 GND.n3046 9.3005
R3590 GND.n3006 GND.n3005 9.3005
R3591 GND.n2980 GND.n2979 9.3005
R3592 GND.n2989 GND.n2988 9.3005
R3593 GND.n2971 GND.n2970 9.3005
R3594 GND.n2978 GND.n2977 9.3005
R3595 GND.n2545 GND.n2544 9.3005
R3596 GND.n2621 GND.n2620 9.3005
R3597 GND.n2580 GND.n2579 9.3005
R3598 GND.n2554 GND.n2553 9.3005
R3599 GND.n2563 GND.n2562 9.3005
R3600 GND.n7192 GND.n7191 9.3005
R3601 GND.n2552 GND.n2551 9.3005
R3602 GND.n7150 GND.n7149 9.3005
R3603 GND.n7225 GND.n7224 9.3005
R3604 GND.n7180 GND.n7179 9.3005
R3605 GND.n7154 GND.n7153 9.3005
R3606 GND.n7163 GND.n7162 9.3005
R3607 GND.n7034 GND.n7033 9.3005
R3608 GND.n7152 GND.n7151 9.3005
R3609 GND.n7066 GND.n7065 9.3005
R3610 GND.n6986 GND.n6985 9.3005
R3611 GND.n7017 GND.n7016 9.3005
R3612 GND.n6991 GND.n6990 9.3005
R3613 GND.n7000 GND.n6999 9.3005
R3614 GND.n6880 GND.n6879 9.3005
R3615 GND.n6989 GND.n6988 9.3005
R3616 GND.n6912 GND.n6911 9.3005
R3617 GND.n6832 GND.n6831 9.3005
R3618 GND.n6863 GND.n6862 9.3005
R3619 GND.n6837 GND.n6836 9.3005
R3620 GND.n6846 GND.n6845 9.3005
R3621 GND.n6726 GND.n6725 9.3005
R3622 GND.n6835 GND.n6834 9.3005
R3623 GND.n6758 GND.n6757 9.3005
R3624 GND.n6668 GND.n6667 9.3005
R3625 GND.n6709 GND.n6708 9.3005
R3626 GND.n6683 GND.n6682 9.3005
R3627 GND.n6692 GND.n6691 9.3005
R3628 GND.n6674 GND.n6673 9.3005
R3629 GND.n6681 GND.n6680 9.3005
R3630 GND.n6558 GND.n6557 9.3005
R3631 GND.n638 GND.n637 9.3005
R3632 GND.n6638 GND.n6637 9.3005
R3633 GND.n6612 GND.n6611 9.3005
R3634 GND.n6621 GND.n6620 9.3005
R3635 GND.n6603 GND.n6602 9.3005
R3636 GND.n6610 GND.n6609 9.3005
R3637 GND.n5619 GND.n5618 9.3005
R3638 GND.n5525 GND.n5524 9.3005
R3639 GND.n5590 GND.n5589 9.3005
R3640 GND.n5564 GND.n5563 9.3005
R3641 GND.n5573 GND.n5572 9.3005
R3642 GND.n5555 GND.n5554 9.3005
R3643 GND.n5562 GND.n5561 9.3005
R3644 GND.n5484 GND.n5483 9.3005
R3645 GND.n5469 GND.n5468 9.3005
R3646 GND.n1088 GND.n1087 9.3005
R3647 GND.n1062 GND.n1061 9.3005
R3648 GND.n1071 GND.n1070 9.3005
R3649 GND.n1053 GND.n1052 9.3005
R3650 GND.n1060 GND.n1059 9.3005
R3651 GND.n1272 GND.n1271 9.3005
R3652 GND.n1140 GND.n1139 9.3005
R3653 GND.n1209 GND.n1208 9.3005
R3654 GND.n1183 GND.n1182 9.3005
R3655 GND.n1192 GND.n1191 9.3005
R3656 GND.n1174 GND.n1173 9.3005
R3657 GND.n1181 GND.n1180 9.3005
R3658 GND.n3633 GND.n3632 9.3005
R3659 GND.n3708 GND.n3707 9.3005
R3660 GND.n3670 GND.n3669 9.3005
R3661 GND.n3644 GND.n3643 9.3005
R3662 GND.n3653 GND.n3652 9.3005
R3663 GND.n3635 GND.n3634 9.3005
R3664 GND.n3642 GND.n3641 9.3005
R3665 GND.n5027 GND.n5026 9.3005
R3666 GND.n5108 GND.n5107 9.3005
R3667 GND.n5067 GND.n5066 9.3005
R3668 GND.n5041 GND.n5040 9.3005
R3669 GND.n5050 GND.n5049 9.3005
R3670 GND.n5032 GND.n5031 9.3005
R3671 GND.n5039 GND.n5038 9.3005
R3672 GND.n422 GND.n421 9.3005
R3673 GND.n502 GND.n501 9.3005
R3674 GND.n462 GND.n461 9.3005
R3675 GND.n436 GND.n435 9.3005
R3676 GND.n445 GND.n444 9.3005
R3677 GND.n427 GND.n426 9.3005
R3678 GND.n434 GND.n433 9.3005
R3679 GND.n320 GND.n319 9.3005
R3680 GND.n317 GND.n316 9.3005
R3681 GND.n393 GND.n392 9.3005
R3682 GND.n367 GND.n366 9.3005
R3683 GND.n376 GND.n375 9.3005
R3684 GND.n358 GND.n357 9.3005
R3685 GND.n365 GND.n364 9.3005
R3686 GND.n218 GND.n217 9.3005
R3687 GND.n215 GND.n214 9.3005
R3688 GND.n289 GND.n288 9.3005
R3689 GND.n263 GND.n262 9.3005
R3690 GND.n272 GND.n271 9.3005
R3691 GND.n254 GND.n253 9.3005
R3692 GND.n261 GND.n260 9.3005
R3693 GND.n4944 GND.n4942 9.1766
R3694 GND.n2889 GND.n2887 9.1766
R3695 GND.n2333 GND.n2331 9.1766
R3696 GND.n7736 GND.n7734 9.1766
R3697 GND.n1592 GND.n1590 9.1766
R3698 GND.n5432 GND.n5430 9.1766
R3699 GND.n5297 GND.n5295 9.1766
R3700 GND.n3092 GND.n3091 8.84768
R3701 GND.n4015 GND.n4014 8.84768
R3702 GND.n5154 GND.n5153 8.84768
R3703 GND.n3753 GND.n3752 8.84768
R3704 GND.n1288 GND.n1287 8.84768
R3705 GND.n3431 GND.n3430 8.84768
R3706 GND.n1456 GND.n1455 8.84768
R3707 GND.n1882 GND.n1881 8.84768
R3708 GND.n97 GND.n96 8.84768
R3709 GND.n2133 GND.n2132 8.84768
R3710 GND.n2195 GND.n2194 8.84768
R3711 GND.n2358 GND.n2357 8.84768
R3712 GND.n2670 GND.n2669 8.84768
R3713 GND.n4811 GND.n4810 8.84768
R3714 GND.n4604 GND.n4603 8.84768
R3715 GND.n3270 GND.t595 8.70904
R3716 GND.n7565 GND.t689 8.70904
R3717 GND.n201 GND.t611 8.70904
R3718 GND.n2527 GND.t424 8.70904
R3719 GND.n2950 GND.t1045 8.70904
R3720 GND.n6922 GND.t1182 8.70904
R3721 GND.n6768 GND.t405 8.70904
R3722 GND.n6659 GND.t1405 8.70904
R3723 GND.n5521 GND.t474 8.70904
R3724 GND.n1269 GND.t1155 8.70904
R3725 GND.n7503 GND.t628 8.70904
R3726 GND.n5009 GND.t1354 8.70904
R3727 GND.n3615 GND.t11 8.70904
R3728 GND.n5464 GND.t636 8.70904
R3729 GND.n5642 GND.t1061 8.70904
R3730 GND.n7076 GND.t1159 8.70904
R3731 GND.n3275 GND.t1423 8.70236
R3732 GND.n321 GND.t435 8.70236
R3733 GND.n219 GND.t1073 8.70236
R3734 GND.n2543 GND.t1492 8.70236
R3735 GND.n2967 GND.t602 8.70236
R3736 GND.n7067 GND.t1545 8.70236
R3737 GND.n6913 GND.t623 8.70236
R3738 GND.n6759 GND.t609 8.70236
R3739 GND.n5617 GND.t1323 8.70236
R3740 GND.n1141 GND.t1477 8.70236
R3741 GND.n420 GND.t548 8.70236
R3742 GND.n5025 GND.t612 8.70236
R3743 GND.n3631 GND.t1504 8.70236
R3744 GND.n5482 GND.t707 8.70236
R3745 GND.n6559 GND.t1476 8.70236
R3746 GND.n7148 GND.t1551 8.70236
R3747 GND.t1384 GND 8.56337
R3748 GND.t603 GND 8.43164
R3749 GND.t1152 GND.t1115 8.20945
R3750 GND.t1167 GND.t661 8.20945
R3751 GND.t363 GND.t1520 8.20945
R3752 GND.t853 GND.t1169 8.20945
R3753 GND.t1411 GND.t1343 8.20945
R3754 GND.t359 GND.t495 8.20945
R3755 GND.t1386 GND.t245 8.20945
R3756 GND.t261 GND.t1021 8.20945
R3757 GND.t265 GND.t456 8.20945
R3758 GND.t313 GND.t259 8.20945
R3759 GND.t881 GND.t418 8.20945
R3760 GND.t248 GND.t1535 8.20945
R3761 GND.t543 GND.t869 8.20945
R3762 GND.t1424 GND.t1396 8.20945
R3763 GND.t557 GND.t1087 8.20945
R3764 GND.t684 GND.t637 8.20945
R3765 GND.n4896 GND 8.05791
R3766 GND.n4695 GND 8.05791
R3767 GND.n3150 GND 8.05791
R3768 GND.n2819 GND 8.05791
R3769 GND.n2280 GND 8.05791
R3770 GND.n7684 GND 8.05791
R3771 GND.n1540 GND 8.05791
R3772 GND.n5377 GND 8.05791
R3773 GND.n3946 GND 8.05791
R3774 GND.n5238 GND 8.05791
R3775 GND.n3838 GND 8.05791
R3776 GND.n3515 GND 8.05791
R3777 GND.n1967 GND 8.05791
R3778 GND.n2054 GND 8.05791
R3779 GND.n2442 GND 8.05791
R3780 GND.n2751 GND 8.05791
R3781 GND.t1072 GND.n4251 8.02446
R3782 GND.n4894 GND.n4893 7.90638
R3783 GND.n4693 GND.n4692 7.90638
R3784 GND.n3148 GND.n3147 7.90638
R3785 GND.n2860 GND.n2859 7.90638
R3786 GND.n2278 GND.n2277 7.90638
R3787 GND.n7682 GND.n7681 7.90638
R3788 GND.n1538 GND.n1537 7.90638
R3789 GND.n5375 GND.n5374 7.90638
R3790 GND.n3944 GND.n3943 7.90638
R3791 GND.n5236 GND.n5235 7.90638
R3792 GND.n3836 GND.n3835 7.90638
R3793 GND.n3513 GND.n3512 7.90638
R3794 GND.n1965 GND.n1964 7.90638
R3795 GND.n2074 GND.n2073 7.90638
R3796 GND.n2440 GND.n2439 7.90638
R3797 GND.n2749 GND.n2748 7.90638
R3798 GND.n7446 GND 7.56079
R3799 GND.n6121 GND.t901 7.37892
R3800 GND.n3130 GND.t533 6.88164
R3801 GND.n4053 GND.t559 6.88164
R3802 GND.n5178 GND.t550 6.88164
R3803 GND.n3777 GND.t1133 6.88164
R3804 GND.n1312 GND.t571 6.88164
R3805 GND.n3455 GND.t271 6.88164
R3806 GND.n1480 GND.t645 6.88164
R3807 GND.n1906 GND.t1145 6.88164
R3808 GND.n129 GND.t300 6.88164
R3809 GND.n2157 GND.t565 6.88164
R3810 GND.n2219 GND.t1143 6.88164
R3811 GND.n2382 GND.t1131 6.88164
R3812 GND.n2706 GND.t569 6.88164
R3813 GND.n4835 GND.t302 6.88164
R3814 GND.n4628 GND.t1129 6.88164
R3815 GND.n7815 GND.n0 6.77697
R3816 GND.n984 GND.n971 6.77697
R3817 GND.n6451 GND.n6423 6.77697
R3818 GND.n6445 GND.n6424 6.77697
R3819 GND.n6439 GND.n6425 6.77697
R3820 GND.n6433 GND.n6426 6.77697
R3821 GND.n536 GND.n508 6.77697
R3822 GND.n530 GND.n509 6.77697
R3823 GND.n524 GND.n510 6.77697
R3824 GND.n518 GND.n511 6.77697
R3825 GND.n6110 GND.n6097 6.77697
R3826 GND.t1263 GND.n5695 6.70101
R3827 GND.n2769 GND.n2768 6.52989
R3828 GND.n4723 GND.n4722 6.5285
R3829 GND.n3191 GND.n3190 6.5285
R3830 GND.n2877 GND.n2876 6.5285
R3831 GND.n2321 GND.n2320 6.5285
R3832 GND.n7724 GND.n7723 6.5285
R3833 GND.n1580 GND.n1579 6.5285
R3834 GND.n5420 GND.n5419 6.5285
R3835 GND.n3987 GND.n3986 6.5285
R3836 GND.n5285 GND.n5284 6.5285
R3837 GND.n3875 GND.n3874 6.5285
R3838 GND.n3548 GND.n3547 6.5285
R3839 GND.n2007 GND.n2006 6.5285
R3840 GND.n2096 GND.n2095 6.5285
R3841 GND.n2475 GND.n2474 6.5285
R3842 GND.n4932 GND.n4931 6.5285
R3843 GND.n41 GND.n40 6.4005
R3844 GND.n6368 GND.n6367 6.4005
R3845 GND.n6487 GND.n6482 6.4005
R3846 GND.n6484 GND.n6479 6.4005
R3847 GND.n655 GND.n643 6.4005
R3848 GND.n661 GND.n660 6.4005
R3849 GND.n6397 GND.n6392 6.4005
R3850 GND.n6394 GND.n6389 6.4005
R3851 GND.n6283 GND.n6271 6.4005
R3852 GND.n6289 GND.n6288 6.4005
R3853 GND.n7827 GND.n7826 6.15638
R3854 GND.n973 GND.n972 6.15638
R3855 GND.n6099 GND.n6098 6.15638
R3856 GND.n7758 GND.n7757 6.02403
R3857 GND.n593 GND.n592 5.64756
R3858 GND.n7420 GND.n7419 5.64756
R3859 GND.n7340 GND.n7339 5.64756
R3860 GND.n7292 GND.n7291 5.64756
R3861 GND.n7240 GND.n7239 5.64756
R3862 GND.n2839 GND 5.64756
R3863 GND.n4874 GND 5.64756
R3864 GND.n4660 GND 5.64756
R3865 GND.n3211 GND 5.64756
R3866 GND.n2258 GND 5.64756
R3867 GND.n161 GND 5.64756
R3868 GND.n1518 GND 5.64756
R3869 GND.n5355 GND 5.64756
R3870 GND.n3924 GND 5.64756
R3871 GND.n5216 GND 5.64756
R3872 GND.n3816 GND 5.64756
R3873 GND.n3493 GND 5.64756
R3874 GND.n1945 GND 5.64756
R3875 GND.n2042 GND 5.64756
R3876 GND.n2420 GND 5.64756
R3877 GND.n2729 GND 5.64756
R3878 GND.n5815 GND.n5814 5.64756
R3879 GND.n5769 GND.n5768 5.64756
R3880 GND.n5732 GND.n5731 5.64756
R3881 GND.n6167 GND.n6166 5.64756
R3882 GND.n5672 GND.n5671 5.64756
R3883 GND.n925 GND.n924 5.64756
R3884 GND.n912 GND.n911 5.64756
R3885 GND.n713 GND.n712 5.64756
R3886 GND.n819 GND.n818 5.64756
R3887 GND.n722 GND.n721 5.64756
R3888 GND.n6051 GND.n6050 5.64756
R3889 GND.n5857 GND.n5856 5.64756
R3890 GND.n5969 GND.n5968 5.64756
R3891 GND.n5921 GND.n5920 5.64756
R3892 GND.n5869 GND.n5868 5.64756
R3893 GND.n3015 GND.n3014 5.62907
R3894 GND.n2584 GND.n2583 5.62907
R3895 GND.n7186 GND.n7185 5.62907
R3896 GND.n7023 GND.n7022 5.62907
R3897 GND.n6869 GND.n6868 5.62907
R3898 GND.n6715 GND.n6714 5.62907
R3899 GND.n6566 GND.n6565 5.62907
R3900 GND.n6591 GND.n6590 5.62907
R3901 GND.n5543 GND.n5542 5.62907
R3902 GND.n1148 GND.n1147 5.62907
R3903 GND.n3674 GND.n3673 5.62907
R3904 GND.n5071 GND.n5070 5.62907
R3905 GND.n466 GND.n465 5.62907
R3906 GND.n328 GND.n327 5.62907
R3907 GND.n226 GND.n225 5.62907
R3908 GND.n7633 GND.n7632 5.62907
R3909 GND.n4849 GND.n4818 5.1205
R3910 GND.n4642 GND.n4611 5.1205
R3911 GND.n2708 GND.n2677 5.1205
R3912 GND.n3132 GND.n3099 5.1205
R3913 GND.n3388 GND.n3367 5.1205
R3914 GND.n2233 GND.n2202 5.1205
R3915 GND.n2171 GND.n2140 5.1205
R3916 GND.n143 GND.n104 5.1205
R3917 GND.n1494 GND.n1463 5.1205
R3918 GND.n1326 GND.n1295 5.1205
R3919 GND.n4055 GND.n4022 5.1205
R3920 GND.n5192 GND.n5161 5.1205
R3921 GND.n3791 GND.n3760 5.1205
R3922 GND.n3469 GND.n3438 5.1205
R3923 GND.n1920 GND.n1889 5.1205
R3924 GND.n2396 GND.n2365 5.1205
R3925 GND.n4176 GND.n4175 4.90717
R3926 GND.n571 GND.n570 4.89462
R3927 GND.n7397 GND.n7396 4.89462
R3928 GND.n7350 GND.n7349 4.89462
R3929 GND.n7315 GND.n7314 4.89462
R3930 GND.n7265 GND.n7264 4.89462
R3931 GND.n6952 GND.n6951 4.89462
R3932 GND.n78 GND.n77 4.89462
R3933 GND.n1248 GND.n1247 4.89462
R3934 GND.n7490 GND.n7489 4.89462
R3935 GND.n4989 GND.n4988 4.89462
R3936 GND.n5791 GND.n5790 4.89462
R3937 GND.n5708 GND.n5707 4.89462
R3938 GND.n5655 GND.n5654 4.89462
R3939 GND.n6190 GND.n6189 4.89462
R3940 GND.n5842 GND.n5841 4.89462
R3941 GND.n947 GND.n946 4.89462
R3942 GND.n889 GND.n888 4.89462
R3943 GND.n848 GND.n847 4.89462
R3944 GND.n796 GND.n795 4.89462
R3945 GND.n750 GND.n749 4.89462
R3946 GND.n6073 GND.n6072 4.89462
R3947 GND.n6025 GND.n6024 4.89462
R3948 GND.n5979 GND.n5978 4.89462
R3949 GND.n5944 GND.n5943 4.89462
R3950 GND.n5894 GND.n5893 4.89462
R3951 GND.n4267 GND.t1566 4.78444
R3952 GND.n3237 GND 4.66821
R3953 GND.n7540 GND 4.66821
R3954 GND.n7602 GND 4.66821
R3955 GND.n2501 GND 4.66821
R3956 GND.n2918 GND 4.66821
R3957 GND.n6940 GND 4.66821
R3958 GND.n6777 GND 4.66821
R3959 GND.n66 GND 4.66821
R3960 GND.n1010 GND 4.66821
R3961 GND.n1239 GND 4.66821
R3962 GND.n7478 GND 4.66821
R3963 GND.n4977 GND 4.66821
R3964 GND.n3583 GND 4.66821
R3965 GND.n1109 GND 4.66821
R3966 GND.n6531 GND 4.66821
R3967 GND.n7109 GND 4.66821
R3968 GND.n35 GND.n28 4.6505
R3969 GND.n46 GND.n25 4.6505
R3970 GND.n45 GND.n44 4.6505
R3971 GND.n43 GND.n26 4.6505
R3972 GND.n42 GND.n41 4.6505
R3973 GND.n38 GND.n27 4.6505
R3974 GND.n37 GND.n36 4.6505
R3975 GND.n34 GND.n33 4.6505
R3976 GND.n3250 GND.n3249 4.6505
R3977 GND.n3325 GND.n3324 4.6505
R3978 GND.n3337 GND.n3336 4.6505
R3979 GND.n7553 GND.n7552 4.6505
R3980 GND.n7512 GND.n7511 4.6505
R3981 GND.n7524 GND.n7523 4.6505
R3982 GND.n7615 GND.n7614 4.6505
R3983 GND.n7574 GND.n7573 4.6505
R3984 GND.n7586 GND.n7585 4.6505
R3985 GND.n2511 GND.n2510 4.6505
R3986 GND.n2628 GND.n2627 4.6505
R3987 GND.n2640 GND.n2639 4.6505
R3988 GND.n2928 GND.n2927 4.6505
R3989 GND.n3054 GND.n3053 4.6505
R3990 GND.n3066 GND.n3065 4.6505
R3991 GND.n6954 GND.n6953 4.6505
R3992 GND.n6978 GND.n6925 4.6505
R3993 GND.n6932 GND.n6931 4.6505
R3994 GND.n6790 GND.n6789 4.6505
R3995 GND.n6824 GND.n6771 4.6505
R3996 GND.n6809 GND.n6808 4.6505
R3997 GND.n80 GND.n79 4.6505
R3998 GND.n7760 GND.n51 4.6505
R3999 GND.n57 GND.n56 4.6505
R4000 GND.n1023 GND.n1022 4.6505
R4001 GND.n5640 GND.n995 4.6505
R4002 GND.n1002 GND.n1001 4.6505
R4003 GND.n1250 GND.n1249 4.6505
R4004 GND.n5456 GND.n1224 4.6505
R4005 GND.n1231 GND.n1230 4.6505
R4006 GND.n7492 GND.n7491 4.6505
R4007 GND.n7450 GND.n7449 4.6505
R4008 GND.n7462 GND.n7461 4.6505
R4009 GND.n4991 GND.n4990 4.6505
R4010 GND.n5115 GND.n5114 4.6505
R4011 GND.n5127 GND.n5126 4.6505
R4012 GND.n3593 GND.n3592 4.6505
R4013 GND.n3715 GND.n3714 4.6505
R4014 GND.n3727 GND.n3726 4.6505
R4015 GND.n1122 GND.n1121 4.6505
R4016 GND.n5513 GND.n1103 4.6505
R4017 GND.n5498 GND.n5497 4.6505
R4018 GND.n6544 GND.n6543 4.6505
R4019 GND.n6503 GND.n6502 4.6505
R4020 GND.n6519 GND.n6518 4.6505
R4021 GND.n7122 GND.n7121 4.6505
R4022 GND.n7081 GND.n7080 4.6505
R4023 GND.n7093 GND.n7092 4.6505
R4024 GND.n6362 GND.n6355 4.6505
R4025 GND.n6373 GND.n6352 4.6505
R4026 GND.n6372 GND.n6371 4.6505
R4027 GND.n6370 GND.n6353 4.6505
R4028 GND.n6369 GND.n6368 4.6505
R4029 GND.n6365 GND.n6354 4.6505
R4030 GND.n6364 GND.n6363 4.6505
R4031 GND.n6361 GND.n6360 4.6505
R4032 GND.n6209 GND.n6202 4.6505
R4033 GND.n6221 GND.n6200 4.6505
R4034 GND.n6213 GND.n6201 4.6505
R4035 GND.n6220 GND.n6219 4.6505
R4036 GND.n6218 GND.n6217 4.6505
R4037 GND.n6215 GND.n6214 4.6505
R4038 GND.n6211 GND.n6210 4.6505
R4039 GND.n6208 GND.n6207 4.6505
R4040 GND.n6150 GND.n6149 4.6505
R4041 GND.n6152 GND.n6151 4.6505
R4042 GND.n6223 GND.n6199 4.6505
R4043 GND.n6154 GND.n6153 4.6505
R4044 GND.n6158 GND.n6157 4.6505
R4045 GND.n6161 GND.n6160 4.6505
R4046 GND.n6168 GND.n6167 4.6505
R4047 GND.n6171 GND.n6170 4.6505
R4048 GND.n6175 GND.n6174 4.6505
R4049 GND.n6179 GND.n6178 4.6505
R4050 GND.n6181 GND.n6180 4.6505
R4051 GND.n6185 GND.n6184 4.6505
R4052 GND.n6187 GND.n6186 4.6505
R4053 GND.n6191 GND.n6190 4.6505
R4054 GND.n6193 GND.n6192 4.6505
R4055 GND.n6198 GND.n6197 4.6505
R4056 GND.n6226 GND.n6225 4.6505
R4057 GND.n5743 GND.n5742 4.6505
R4058 GND.n5741 GND.n5740 4.6505
R4059 GND.n5737 GND.n5736 4.6505
R4060 GND.n5656 GND.n5655 4.6505
R4061 GND.n6141 GND.n6140 4.6505
R4062 GND.n6145 GND.n6144 4.6505
R4063 GND.n6147 GND.n6146 4.6505
R4064 GND.n5826 GND.n5825 4.6505
R4065 GND.n5780 GND.n5689 4.6505
R4066 GND.n5779 GND.n5690 4.6505
R4067 GND.n5719 GND.n5718 4.6505
R4068 GND.n5721 GND.n5720 4.6505
R4069 GND.n5824 GND.n5823 4.6505
R4070 GND.n5822 GND.n5821 4.6505
R4071 GND.n5818 GND.n5817 4.6505
R4072 GND.n5816 GND.n5815 4.6505
R4073 GND.n5812 GND.n5811 4.6505
R4074 GND.n5810 GND.n5809 4.6505
R4075 GND.n5806 GND.n5805 4.6505
R4076 GND.n5802 GND.n5801 4.6505
R4077 GND.n5800 GND.n5799 4.6505
R4078 GND.n5795 GND.n5794 4.6505
R4079 GND.n5792 GND.n5791 4.6505
R4080 GND.n5788 GND.n5787 4.6505
R4081 GND.n5786 GND.n5785 4.6505
R4082 GND.n5782 GND.n5781 4.6505
R4083 GND.n5778 GND.n5777 4.6505
R4084 GND.n5776 GND.n5775 4.6505
R4085 GND.n5772 GND.n5771 4.6505
R4086 GND.n5770 GND.n5769 4.6505
R4087 GND.n5766 GND.n5765 4.6505
R4088 GND.n5763 GND.n5762 4.6505
R4089 GND.n5694 GND.n5693 4.6505
R4090 GND.n5699 GND.n5698 4.6505
R4091 GND.n5703 GND.n5702 4.6505
R4092 GND.n5705 GND.n5704 4.6505
R4093 GND.n5709 GND.n5708 4.6505
R4094 GND.n5711 GND.n5710 4.6505
R4095 GND.n5715 GND.n5714 4.6505
R4096 GND.n5717 GND.n5716 4.6505
R4097 GND.n5723 GND.n5722 4.6505
R4098 GND.n5727 GND.n5726 4.6505
R4099 GND.n5729 GND.n5728 4.6505
R4100 GND.n5733 GND.n5732 4.6505
R4101 GND.n5735 GND.n5734 4.6505
R4102 GND.n5753 GND.n5752 4.6505
R4103 GND.n5748 GND.n5747 4.6505
R4104 GND.n5828 GND.n5827 4.6505
R4105 GND.n5831 GND.n5830 4.6505
R4106 GND.n5665 GND.n5664 4.6505
R4107 GND.n5668 GND.n5667 4.6505
R4108 GND.n5673 GND.n5672 4.6505
R4109 GND.n5675 GND.n5674 4.6505
R4110 GND.n5679 GND.n5678 4.6505
R4111 GND.n5683 GND.n5682 4.6505
R4112 GND.n5685 GND.n5684 4.6505
R4113 GND.n5849 GND.n5848 4.6505
R4114 GND.n5845 GND.n5844 4.6505
R4115 GND.n5843 GND.n5842 4.6505
R4116 GND.n5839 GND.n5838 4.6505
R4117 GND.n5837 GND.n5836 4.6505
R4118 GND.n761 GND.n760 4.6505
R4119 GND.n763 GND.n762 4.6505
R4120 GND.n785 GND.n773 4.6505
R4121 GND.n784 GND.n774 4.6505
R4122 GND.n860 GND.n859 4.6505
R4123 GND.n862 GND.n861 4.6505
R4124 GND.n878 GND.n872 4.6505
R4125 GND.n877 GND.n873 4.6505
R4126 GND.n958 GND.n957 4.6505
R4127 GND.n960 GND.n959 4.6505
R4128 GND.n970 GND.n969 4.6505
R4129 GND.n719 GND.n718 4.6505
R4130 GND.n723 GND.n722 4.6505
R4131 GND.n726 GND.n725 4.6505
R4132 GND.n734 GND.n733 4.6505
R4133 GND.n739 GND.n738 4.6505
R4134 GND.n741 GND.n740 4.6505
R4135 GND.n745 GND.n744 4.6505
R4136 GND.n747 GND.n746 4.6505
R4137 GND.n751 GND.n750 4.6505
R4138 GND.n753 GND.n752 4.6505
R4139 GND.n757 GND.n756 4.6505
R4140 GND.n759 GND.n758 4.6505
R4141 GND.n765 GND.n764 4.6505
R4142 GND.n769 GND.n768 4.6505
R4143 GND.n772 GND.n771 4.6505
R4144 GND.n820 GND.n819 4.6505
R4145 GND.n815 GND.n814 4.6505
R4146 GND.n813 GND.n812 4.6505
R4147 GND.n809 GND.n808 4.6505
R4148 GND.n805 GND.n804 4.6505
R4149 GND.n803 GND.n802 4.6505
R4150 GND.n799 GND.n798 4.6505
R4151 GND.n797 GND.n796 4.6505
R4152 GND.n793 GND.n792 4.6505
R4153 GND.n791 GND.n790 4.6505
R4154 GND.n787 GND.n786 4.6505
R4155 GND.n783 GND.n782 4.6505
R4156 GND.n781 GND.n780 4.6505
R4157 GND.n777 GND.n776 4.6505
R4158 GND.n714 GND.n713 4.6505
R4159 GND.n828 GND.n827 4.6505
R4160 GND.n833 GND.n832 4.6505
R4161 GND.n837 GND.n836 4.6505
R4162 GND.n839 GND.n838 4.6505
R4163 GND.n843 GND.n842 4.6505
R4164 GND.n845 GND.n844 4.6505
R4165 GND.n849 GND.n848 4.6505
R4166 GND.n851 GND.n850 4.6505
R4167 GND.n855 GND.n854 4.6505
R4168 GND.n858 GND.n857 4.6505
R4169 GND.n864 GND.n863 4.6505
R4170 GND.n868 GND.n867 4.6505
R4171 GND.n871 GND.n870 4.6505
R4172 GND.n913 GND.n912 4.6505
R4173 GND.n908 GND.n907 4.6505
R4174 GND.n906 GND.n905 4.6505
R4175 GND.n902 GND.n901 4.6505
R4176 GND.n898 GND.n897 4.6505
R4177 GND.n896 GND.n895 4.6505
R4178 GND.n892 GND.n891 4.6505
R4179 GND.n890 GND.n889 4.6505
R4180 GND.n886 GND.n885 4.6505
R4181 GND.n884 GND.n883 4.6505
R4182 GND.n880 GND.n879 4.6505
R4183 GND.n876 GND.n875 4.6505
R4184 GND.n710 GND.n709 4.6505
R4185 GND.n921 GND.n920 4.6505
R4186 GND.n926 GND.n925 4.6505
R4187 GND.n928 GND.n927 4.6505
R4188 GND.n932 GND.n931 4.6505
R4189 GND.n936 GND.n935 4.6505
R4190 GND.n938 GND.n937 4.6505
R4191 GND.n942 GND.n941 4.6505
R4192 GND.n944 GND.n943 4.6505
R4193 GND.n948 GND.n947 4.6505
R4194 GND.n950 GND.n949 4.6505
R4195 GND.n954 GND.n953 4.6505
R4196 GND.n956 GND.n955 4.6505
R4197 GND.n962 GND.n961 4.6505
R4198 GND.n965 GND.n964 4.6505
R4199 GND.n967 GND.n966 4.6505
R4200 GND.n990 GND.n989 4.6505
R4201 GND.n987 GND.n986 4.6505
R4202 GND.n985 GND.n984 4.6505
R4203 GND.n983 GND.n982 4.6505
R4204 GND.n981 GND.n980 4.6505
R4205 GND.n979 GND.n978 4.6505
R4206 GND.n975 GND.n974 4.6505
R4207 GND.n20 GND.n19 4.6505
R4208 GND.n18 GND.n8 4.6505
R4209 GND.n17 GND.n16 4.6505
R4210 GND.n16 GND.n15 4.6505
R4211 GND.n14 GND.n8 4.6505
R4212 GND.n20 GND.n7 4.6505
R4213 GND.n22 GND.n21 4.6505
R4214 GND.n7776 GND.n7771 4.6505
R4215 GND.n7778 GND.n7777 4.6505
R4216 GND.n7785 GND.n7784 4.6505
R4217 GND.n7786 GND.n7766 4.6505
R4218 GND.n7788 GND.n7787 4.6505
R4219 GND.n7781 GND.n7769 4.6505
R4220 GND.n7784 GND.n7783 4.6505
R4221 GND.n7782 GND.n7766 4.6505
R4222 GND.n7788 GND.n7765 4.6505
R4223 GND.n7790 GND.n7789 4.6505
R4224 GND.n6480 GND.n6479 4.6505
R4225 GND.n6491 GND.n6490 4.6505
R4226 GND.n6487 GND.n6486 4.6505
R4227 GND.n6489 GND.n6488 4.6505
R4228 GND.n662 GND.n661 4.6505
R4229 GND.n653 GND.n646 4.6505
R4230 GND.n652 GND.n651 4.6505
R4231 GND.n658 GND.n657 4.6505
R4232 GND.n656 GND.n644 4.6505
R4233 GND.n662 GND.n643 4.6505
R4234 GND.n664 GND.n663 4.6505
R4235 GND.n683 GND.n677 4.6505
R4236 GND.n686 GND.n676 4.6505
R4237 GND.n674 GND.n673 4.6505
R4238 GND.n700 GND.n671 4.6505
R4239 GND.n682 GND.n681 4.6505
R4240 GND.n685 GND.n684 4.6505
R4241 GND.n688 GND.n687 4.6505
R4242 GND.n690 GND.n689 4.6505
R4243 GND.n699 GND.n698 4.6505
R4244 GND.n701 GND.n668 4.6505
R4245 GND.n703 GND.n702 4.6505
R4246 GND.n696 GND.n671 4.6505
R4247 GND.n698 GND.n697 4.6505
R4248 GND.n694 GND.n668 4.6505
R4249 GND.n703 GND.n669 4.6505
R4250 GND.n6430 GND.n6429 4.6505
R4251 GND.n6432 GND.n6431 4.6505
R4252 GND.n6434 GND.n6433 4.6505
R4253 GND.n6436 GND.n6435 4.6505
R4254 GND.n6438 GND.n6437 4.6505
R4255 GND.n6440 GND.n6439 4.6505
R4256 GND.n6442 GND.n6441 4.6505
R4257 GND.n6444 GND.n6443 4.6505
R4258 GND.n6446 GND.n6445 4.6505
R4259 GND.n6448 GND.n6447 4.6505
R4260 GND.n6450 GND.n6449 4.6505
R4261 GND.n6452 GND.n6451 4.6505
R4262 GND.n6345 GND.n6344 4.6505
R4263 GND.n6343 GND.n6333 4.6505
R4264 GND.n6342 GND.n6341 4.6505
R4265 GND.n6341 GND.n6340 4.6505
R4266 GND.n6339 GND.n6333 4.6505
R4267 GND.n6345 GND.n6332 4.6505
R4268 GND.n6347 GND.n6346 4.6505
R4269 GND.n6309 GND.n6304 4.6505
R4270 GND.n6311 GND.n6310 4.6505
R4271 GND.n6318 GND.n6317 4.6505
R4272 GND.n6319 GND.n6299 4.6505
R4273 GND.n6321 GND.n6320 4.6505
R4274 GND.n6314 GND.n6302 4.6505
R4275 GND.n6317 GND.n6316 4.6505
R4276 GND.n6315 GND.n6299 4.6505
R4277 GND.n6321 GND.n6298 4.6505
R4278 GND.n6323 GND.n6322 4.6505
R4279 GND.n6390 GND.n6389 4.6505
R4280 GND.n6401 GND.n6400 4.6505
R4281 GND.n6397 GND.n6396 4.6505
R4282 GND.n6399 GND.n6398 4.6505
R4283 GND.n6290 GND.n6289 4.6505
R4284 GND.n6281 GND.n6274 4.6505
R4285 GND.n6280 GND.n6279 4.6505
R4286 GND.n6286 GND.n6285 4.6505
R4287 GND.n6284 GND.n6272 4.6505
R4288 GND.n6290 GND.n6271 4.6505
R4289 GND.n6292 GND.n6291 4.6505
R4290 GND.n6247 GND.n6241 4.6505
R4291 GND.n6250 GND.n6240 4.6505
R4292 GND.n6238 GND.n6237 4.6505
R4293 GND.n6264 GND.n6235 4.6505
R4294 GND.n6246 GND.n6245 4.6505
R4295 GND.n6249 GND.n6248 4.6505
R4296 GND.n6252 GND.n6251 4.6505
R4297 GND.n6254 GND.n6253 4.6505
R4298 GND.n6263 GND.n6262 4.6505
R4299 GND.n6265 GND.n6232 4.6505
R4300 GND.n6267 GND.n6266 4.6505
R4301 GND.n6260 GND.n6235 4.6505
R4302 GND.n6262 GND.n6261 4.6505
R4303 GND.n6258 GND.n6232 4.6505
R4304 GND.n6267 GND.n6233 4.6505
R4305 GND.n515 GND.n514 4.6505
R4306 GND.n517 GND.n516 4.6505
R4307 GND.n519 GND.n518 4.6505
R4308 GND.n521 GND.n520 4.6505
R4309 GND.n523 GND.n522 4.6505
R4310 GND.n525 GND.n524 4.6505
R4311 GND.n527 GND.n526 4.6505
R4312 GND.n529 GND.n528 4.6505
R4313 GND.n531 GND.n530 4.6505
R4314 GND.n533 GND.n532 4.6505
R4315 GND.n535 GND.n534 4.6505
R4316 GND.n537 GND.n536 4.6505
R4317 GND.n5883 GND.n5873 4.6505
R4318 GND.n5882 GND.n5874 4.6505
R4319 GND.n5955 GND.n5954 4.6505
R4320 GND.n5957 GND.n5956 4.6505
R4321 GND.n6134 GND.n5853 4.6505
R4322 GND.n6133 GND.n5854 4.6505
R4323 GND.n6036 GND.n6035 4.6505
R4324 GND.n6038 GND.n6037 4.6505
R4325 GND.n6084 GND.n6083 4.6505
R4326 GND.n6086 GND.n6085 4.6505
R4327 GND.n6096 GND.n6095 4.6505
R4328 GND.n5866 GND.n5865 4.6505
R4329 GND.n5870 GND.n5869 4.6505
R4330 GND.n5872 GND.n5871 4.6505
R4331 GND.n5912 GND.n5911 4.6505
R4332 GND.n5907 GND.n5906 4.6505
R4333 GND.n5903 GND.n5902 4.6505
R4334 GND.n5901 GND.n5900 4.6505
R4335 GND.n5897 GND.n5896 4.6505
R4336 GND.n5895 GND.n5894 4.6505
R4337 GND.n5891 GND.n5890 4.6505
R4338 GND.n5889 GND.n5888 4.6505
R4339 GND.n5885 GND.n5884 4.6505
R4340 GND.n5881 GND.n5880 4.6505
R4341 GND.n5879 GND.n5878 4.6505
R4342 GND.n5860 GND.n5859 4.6505
R4343 GND.n5922 GND.n5921 4.6505
R4344 GND.n5925 GND.n5924 4.6505
R4345 GND.n5929 GND.n5928 4.6505
R4346 GND.n5933 GND.n5932 4.6505
R4347 GND.n5935 GND.n5934 4.6505
R4348 GND.n5939 GND.n5938 4.6505
R4349 GND.n5941 GND.n5940 4.6505
R4350 GND.n5945 GND.n5944 4.6505
R4351 GND.n5947 GND.n5946 4.6505
R4352 GND.n5951 GND.n5950 4.6505
R4353 GND.n5953 GND.n5952 4.6505
R4354 GND.n5959 GND.n5958 4.6505
R4355 GND.n5963 GND.n5962 4.6505
R4356 GND.n5965 GND.n5964 4.6505
R4357 GND.n5970 GND.n5969 4.6505
R4358 GND.n5999 GND.n5998 4.6505
R4359 GND.n5996 GND.n5995 4.6505
R4360 GND.n5992 GND.n5991 4.6505
R4361 GND.n5988 GND.n5987 4.6505
R4362 GND.n5986 GND.n5985 4.6505
R4363 GND.n5982 GND.n5981 4.6505
R4364 GND.n5980 GND.n5979 4.6505
R4365 GND.n5976 GND.n5975 4.6505
R4366 GND.n5974 GND.n5973 4.6505
R4367 GND.n5852 GND.n5851 4.6505
R4368 GND.n6132 GND.n6131 4.6505
R4369 GND.n6130 GND.n6129 4.6505
R4370 GND.n6125 GND.n6124 4.6505
R4371 GND.n5858 GND.n5857 4.6505
R4372 GND.n6006 GND.n6005 4.6505
R4373 GND.n6010 GND.n6009 4.6505
R4374 GND.n6014 GND.n6013 4.6505
R4375 GND.n6016 GND.n6015 4.6505
R4376 GND.n6020 GND.n6019 4.6505
R4377 GND.n6022 GND.n6021 4.6505
R4378 GND.n6026 GND.n6025 4.6505
R4379 GND.n6028 GND.n6027 4.6505
R4380 GND.n6032 GND.n6031 4.6505
R4381 GND.n6034 GND.n6033 4.6505
R4382 GND.n6040 GND.n6039 4.6505
R4383 GND.n6044 GND.n6043 4.6505
R4384 GND.n6047 GND.n6046 4.6505
R4385 GND.n6052 GND.n6051 4.6505
R4386 GND.n6054 GND.n6053 4.6505
R4387 GND.n6058 GND.n6057 4.6505
R4388 GND.n6062 GND.n6061 4.6505
R4389 GND.n6064 GND.n6063 4.6505
R4390 GND.n6068 GND.n6067 4.6505
R4391 GND.n6070 GND.n6069 4.6505
R4392 GND.n6074 GND.n6073 4.6505
R4393 GND.n6076 GND.n6075 4.6505
R4394 GND.n6080 GND.n6079 4.6505
R4395 GND.n6082 GND.n6081 4.6505
R4396 GND.n6088 GND.n6087 4.6505
R4397 GND.n6091 GND.n6090 4.6505
R4398 GND.n6093 GND.n6092 4.6505
R4399 GND.n6116 GND.n6115 4.6505
R4400 GND.n6113 GND.n6112 4.6505
R4401 GND.n6111 GND.n6110 4.6505
R4402 GND.n6109 GND.n6108 4.6505
R4403 GND.n6107 GND.n6106 4.6505
R4404 GND.n6105 GND.n6104 4.6505
R4405 GND.n6101 GND.n6100 4.6505
R4406 GND.n7254 GND.n7244 4.6505
R4407 GND.n7253 GND.n7245 4.6505
R4408 GND.n7326 GND.n7325 4.6505
R4409 GND.n7328 GND.n7327 4.6505
R4410 GND.n7433 GND.n545 4.6505
R4411 GND.n7432 GND.n546 4.6505
R4412 GND.n7386 GND.n548 4.6505
R4413 GND.n7385 GND.n549 4.6505
R4414 GND.n560 GND.n550 4.6505
R4415 GND.n559 GND.n551 4.6505
R4416 GND.n2 GND.n1 4.6505
R4417 GND.n7237 GND.n7236 4.6505
R4418 GND.n7241 GND.n7240 4.6505
R4419 GND.n7243 GND.n7242 4.6505
R4420 GND.n7283 GND.n7282 4.6505
R4421 GND.n7278 GND.n7277 4.6505
R4422 GND.n7274 GND.n7273 4.6505
R4423 GND.n7272 GND.n7271 4.6505
R4424 GND.n7268 GND.n7267 4.6505
R4425 GND.n7266 GND.n7265 4.6505
R4426 GND.n7262 GND.n7261 4.6505
R4427 GND.n7260 GND.n7259 4.6505
R4428 GND.n7256 GND.n7255 4.6505
R4429 GND.n7252 GND.n7251 4.6505
R4430 GND.n7250 GND.n7249 4.6505
R4431 GND.n7232 GND.n7231 4.6505
R4432 GND.n7293 GND.n7292 4.6505
R4433 GND.n7296 GND.n7295 4.6505
R4434 GND.n7300 GND.n7299 4.6505
R4435 GND.n7304 GND.n7303 4.6505
R4436 GND.n7306 GND.n7305 4.6505
R4437 GND.n7310 GND.n7309 4.6505
R4438 GND.n7312 GND.n7311 4.6505
R4439 GND.n7316 GND.n7315 4.6505
R4440 GND.n7318 GND.n7317 4.6505
R4441 GND.n7322 GND.n7321 4.6505
R4442 GND.n7324 GND.n7323 4.6505
R4443 GND.n7330 GND.n7329 4.6505
R4444 GND.n7334 GND.n7333 4.6505
R4445 GND.n7336 GND.n7335 4.6505
R4446 GND.n7341 GND.n7340 4.6505
R4447 GND.n7370 GND.n7369 4.6505
R4448 GND.n7367 GND.n7366 4.6505
R4449 GND.n7363 GND.n7362 4.6505
R4450 GND.n7359 GND.n7358 4.6505
R4451 GND.n7357 GND.n7356 4.6505
R4452 GND.n7353 GND.n7352 4.6505
R4453 GND.n7351 GND.n7350 4.6505
R4454 GND.n7347 GND.n7346 4.6505
R4455 GND.n7345 GND.n7344 4.6505
R4456 GND.n544 GND.n543 4.6505
R4457 GND.n7431 GND.n7430 4.6505
R4458 GND.n7429 GND.n7428 4.6505
R4459 GND.n7424 GND.n7423 4.6505
R4460 GND.n7421 GND.n7420 4.6505
R4461 GND.n7416 GND.n7415 4.6505
R4462 GND.n7414 GND.n7413 4.6505
R4463 GND.n7410 GND.n7409 4.6505
R4464 GND.n7406 GND.n7405 4.6505
R4465 GND.n7404 GND.n7403 4.6505
R4466 GND.n7400 GND.n7399 4.6505
R4467 GND.n7398 GND.n7397 4.6505
R4468 GND.n7394 GND.n7393 4.6505
R4469 GND.n7392 GND.n7391 4.6505
R4470 GND.n7388 GND.n7387 4.6505
R4471 GND.n7384 GND.n7383 4.6505
R4472 GND.n7382 GND.n7381 4.6505
R4473 GND.n597 GND.n596 4.6505
R4474 GND.n594 GND.n593 4.6505
R4475 GND.n590 GND.n589 4.6505
R4476 GND.n588 GND.n587 4.6505
R4477 GND.n584 GND.n583 4.6505
R4478 GND.n580 GND.n579 4.6505
R4479 GND.n578 GND.n577 4.6505
R4480 GND.n574 GND.n573 4.6505
R4481 GND.n572 GND.n571 4.6505
R4482 GND.n568 GND.n567 4.6505
R4483 GND.n566 GND.n565 4.6505
R4484 GND.n562 GND.n561 4.6505
R4485 GND.n558 GND.n557 4.6505
R4486 GND.n556 GND.n555 4.6505
R4487 GND.n553 GND.n552 4.6505
R4488 GND.n7810 GND.n7809 4.6505
R4489 GND.n7813 GND.n7812 4.6505
R4490 GND.n7815 GND.n7814 4.6505
R4491 GND.n7817 GND.n7816 4.6505
R4492 GND.n7819 GND.n7818 4.6505
R4493 GND.n7823 GND.n7822 4.6505
R4494 GND.n7825 GND.n7824 4.6505
R4495 GND.n1376 GND.n1375 4.52281
R4496 GND.n1746 GND.n1600 4.51032
R4497 GND.n3243 GND.n3242 4.5005
R4498 GND.n3255 GND.n3248 4.5005
R4499 GND.n3331 GND.n3330 4.5005
R4500 GND.n3341 GND.n3335 4.5005
R4501 GND.n7546 GND.n7545 4.5005
R4502 GND.n7558 GND.n7551 4.5005
R4503 GND.n7518 GND.n7517 4.5005
R4504 GND.n7528 GND.n7522 4.5005
R4505 GND.n7608 GND.n7607 4.5005
R4506 GND.n7620 GND.n7613 4.5005
R4507 GND.n7580 GND.n7579 4.5005
R4508 GND.n7590 GND.n7584 4.5005
R4509 GND.n2507 GND.n2506 4.5005
R4510 GND.n2516 GND.n2509 4.5005
R4511 GND.n2634 GND.n2633 4.5005
R4512 GND.n2644 GND.n2638 4.5005
R4513 GND.n2924 GND.n2923 4.5005
R4514 GND.n2933 GND.n2926 4.5005
R4515 GND.n3060 GND.n3059 4.5005
R4516 GND.n3070 GND.n3064 4.5005
R4517 GND.n6946 GND.n6945 4.5005
R4518 GND.n6958 GND.n6952 4.5005
R4519 GND.n6974 GND.n6927 4.5005
R4520 GND.n6936 GND.n6930 4.5005
R4521 GND.n6783 GND.n6782 4.5005
R4522 GND.n6795 GND.n6788 4.5005
R4523 GND.n6820 GND.n6773 4.5005
R4524 GND.n6813 GND.n6807 4.5005
R4525 GND.n72 GND.n71 4.5005
R4526 GND.n84 GND.n78 4.5005
R4527 GND.n61 GND.n55 4.5005
R4528 GND.n1016 GND.n1015 4.5005
R4529 GND.n1028 GND.n1021 4.5005
R4530 GND.n5636 GND.n997 4.5005
R4531 GND.n1006 GND.n1000 4.5005
R4532 GND.n1245 GND.n1244 4.5005
R4533 GND.n1254 GND.n1248 4.5005
R4534 GND.n5452 GND.n1226 4.5005
R4535 GND.n1235 GND.n1229 4.5005
R4536 GND.n7484 GND.n7483 4.5005
R4537 GND.n7496 GND.n7490 4.5005
R4538 GND.n7456 GND.n7455 4.5005
R4539 GND.n7466 GND.n7460 4.5005
R4540 GND.n4983 GND.n4982 4.5005
R4541 GND.n4995 GND.n4989 4.5005
R4542 GND.n5121 GND.n5120 4.5005
R4543 GND.n5131 GND.n5125 4.5005
R4544 GND.n3589 GND.n3588 4.5005
R4545 GND.n3598 GND.n3591 4.5005
R4546 GND.n3721 GND.n3720 4.5005
R4547 GND.n3731 GND.n3725 4.5005
R4548 GND.n1115 GND.n1114 4.5005
R4549 GND.n1127 GND.n1120 4.5005
R4550 GND.n5509 GND.n1105 4.5005
R4551 GND.n5502 GND.n5496 4.5005
R4552 GND.n6537 GND.n6536 4.5005
R4553 GND.n6549 GND.n6542 4.5005
R4554 GND.n6509 GND.n6508 4.5005
R4555 GND.n6523 GND.n6517 4.5005
R4556 GND.n7115 GND.n7114 4.5005
R4557 GND.n7127 GND.n7120 4.5005
R4558 GND.n7087 GND.n7086 4.5005
R4559 GND.n7097 GND.n7091 4.5005
R4560 GND.n4267 GND.n4070 4.5005
R4561 GND.n4267 GND.n4266 4.5005
R4562 GND.n4461 GND.n4460 4.4805
R4563 GND.n4449 GND.n4448 4.4805
R4564 GND.n7235 GND.n7234 4.45136
R4565 GND.n717 GND.n716 4.45136
R4566 GND.n5864 GND.n5863 4.45136
R4567 GND.n4954 GND.t294 4.41708
R4568 GND.n4970 GND.t653 4.41708
R4569 GND.n2812 GND.t1020 4.41708
R4570 GND.n3399 GND.t1084 4.41708
R4571 GND.n3141 GND.t654 4.41708
R4572 GND.n2343 GND.t297 4.41708
R4573 GND.n2182 GND.t309 4.41708
R4574 GND.n1866 GND.t452 4.41708
R4575 GND.n5327 GND.t1086 4.41708
R4576 GND.n3576 GND.t451 4.41708
R4577 GND.n5315 GND.t310 4.41708
R4578 GND.n5307 GND.t1085 4.41708
R4579 GND.n3897 GND.t852 4.41708
R4580 GND.n3570 GND.t655 4.41708
R4581 GND.n3413 GND.t711 4.41708
R4582 GND.n2497 GND.t851 4.41708
R4583 GND.n4801 GND.t1017 4.35136
R4584 GND.n4971 GND.t295 4.35136
R4585 GND.n3400 GND.t712 4.35136
R4586 GND.n3142 GND.t298 4.35136
R4587 GND.n2344 GND.t1018 4.35136
R4588 GND.n1864 GND.t311 4.35136
R4589 GND.n5328 GND.t713 4.35136
R4590 GND.n1332 GND.t656 4.35136
R4591 GND.n3906 GND.t850 4.35136
R4592 GND.n5308 GND.t1019 4.35136
R4593 GND.n3582 GND.t454 4.35136
R4594 GND.n3419 GND.t710 4.35136
R4595 GND.n1872 GND.t308 4.35136
R4596 GND.n2183 GND.t849 4.35136
R4597 GND.n2498 GND.t453 4.35136
R4598 GND.n2813 GND.t1083 4.35136
R4599 GND.n6231 GND.n6230 4.25025
R4600 GND.n49 GND.n48 4.06709
R4601 GND.n6376 GND.n6375 4.06709
R4602 GND.n11 GND.n10 4.06409
R4603 GND.n6336 GND.n6335 4.06409
R4604 GND.n13 GND.n11 4.0631
R4605 GND.n6338 GND.n6336 4.0631
R4606 GND.n7779 GND.n7768 4.05611
R4607 GND.n6312 GND.n6301 4.05611
R4608 GND.n693 GND.n691 3.98881
R4609 GND.n6257 GND.n6255 3.98881
R4610 GND.n4737 GND.n4736 3.9685
R4611 GND.n2783 GND.n2782 3.9685
R4612 GND.n4458 GND.n4457 3.84205
R4613 GND.n7775 GND.n7774 3.80559
R4614 GND.n650 GND.n648 3.80559
R4615 GND.n6308 GND.n6307 3.80559
R4616 GND.n6278 GND.n6276 3.80559
R4617 GND.n32 GND.n30 3.80083
R4618 GND.n6359 GND.n6357 3.80083
R4619 GND.n4251 GND.n4246 3.69035
R4620 GND.n2116 GND.n2115 3.63686
R4621 GND.n4104 GND.n4071 3.38533
R4622 GND.n4089 GND.n4087 3.20453
R4623 GND.n3246 GND.n3245 3.03311
R4624 GND.n3347 GND.n3346 3.03311
R4625 GND.n7549 GND.n7548 3.03311
R4626 GND.n7534 GND.n7533 3.03311
R4627 GND.n7611 GND.n7610 3.03311
R4628 GND.n7596 GND.n7595 3.03311
R4629 GND.n4657 GND.n4656 3.03311
R4630 GND.n4661 GND.n4660 3.03311
R4631 GND.n2519 GND.n2518 3.03311
R4632 GND.n2650 GND.n2649 3.03311
R4633 GND.n2936 GND.n2935 3.03311
R4634 GND.n3076 GND.n3075 3.03311
R4635 GND.n3201 GND.n3200 3.03311
R4636 GND.n3212 GND.n3211 3.03311
R4637 GND.n6949 GND.n6948 3.03311
R4638 GND.n6969 GND.n6968 3.03311
R4639 GND.n2250 GND.n2249 3.03311
R4640 GND.n2259 GND.n2258 3.03311
R4641 GND.n6786 GND.n6785 3.03311
R4642 GND.n6815 GND.n6805 3.03311
R4643 GND.n75 GND.n74 3.03311
R4644 GND.n64 GND.n53 3.03311
R4645 GND.n158 GND.n157 3.03311
R4646 GND.n162 GND.n161 3.03311
R4647 GND.n1019 GND.n1018 3.03311
R4648 GND.n5631 GND.n5630 3.03311
R4649 GND.n1510 GND.n1509 3.03311
R4650 GND.n1519 GND.n1518 3.03311
R4651 GND.n1257 GND.n1256 3.03311
R4652 GND.n5447 GND.n5446 3.03311
R4653 GND.n5347 GND.n5346 3.03311
R4654 GND.n5356 GND.n5355 3.03311
R4655 GND.n3916 GND.n3915 3.03311
R4656 GND.n3925 GND.n3924 3.03311
R4657 GND.n7487 GND.n7486 3.03311
R4658 GND.n7472 GND.n7471 3.03311
R4659 GND.n4986 GND.n4985 3.03311
R4660 GND.n5137 GND.n5136 3.03311
R4661 GND.n5208 GND.n5207 3.03311
R4662 GND.n5217 GND.n5216 3.03311
R4663 GND.n3601 GND.n3600 3.03311
R4664 GND.n3737 GND.n3736 3.03311
R4665 GND.n3808 GND.n3807 3.03311
R4666 GND.n3817 GND.n3816 3.03311
R4667 GND.n1118 GND.n1117 3.03311
R4668 GND.n5504 GND.n5494 3.03311
R4669 GND.n3485 GND.n3484 3.03311
R4670 GND.n3494 GND.n3493 3.03311
R4671 GND.n6540 GND.n6539 3.03311
R4672 GND.n6525 GND.n6515 3.03311
R4673 GND.n1937 GND.n1936 3.03311
R4674 GND.n1946 GND.n1945 3.03311
R4675 GND.n2039 GND.n2038 3.03311
R4676 GND.n2043 GND.n2042 3.03311
R4677 GND.n7118 GND.n7117 3.03311
R4678 GND.n7103 GND.n7102 3.03311
R4679 GND.n2412 GND.n2411 3.03311
R4680 GND.n2421 GND.n2420 3.03311
R4681 GND.n2721 GND.n2720 3.03311
R4682 GND.n2730 GND.n2729 3.03311
R4683 GND.n4866 GND.n4865 3.03311
R4684 GND.n4875 GND.n4874 3.03311
R4685 GND.n2831 GND.n2830 3.03311
R4686 GND.n2840 GND.n2839 3.03311
R4687 GND.n4898 GND 3.0005
R4688 GND.n4697 GND 3.0005
R4689 GND.n3152 GND 3.0005
R4690 GND.n2821 GND 3.0005
R4691 GND.n2282 GND 3.0005
R4692 GND.n7686 GND 3.0005
R4693 GND.n1542 GND 3.0005
R4694 GND.n5379 GND 3.0005
R4695 GND.n3948 GND 3.0005
R4696 GND.n5240 GND 3.0005
R4697 GND.n3840 GND 3.0005
R4698 GND.n3517 GND 3.0005
R4699 GND.n1969 GND 3.0005
R4700 GND.n2056 GND 3.0005
R4701 GND.n2444 GND 3.0005
R4702 GND.n2753 GND 3.0005
R4703 GND.n916 GND.t815 2.84655
R4704 GND.n5231 GND.n5230 2.5872
R4705 GND.n5370 GND.n5369 2.5872
R4706 GND.n1533 GND.n1532 2.5872
R4707 GND.n7677 GND.n7676 2.5872
R4708 GND.n2273 GND.n2272 2.5872
R4709 GND.n2744 GND.n2743 2.5872
R4710 GND.n4889 GND.n4888 2.5872
R4711 GND.n2855 GND.n2854 2.56838
R4712 GND.n3939 GND.n3938 2.56838
R4713 GND.n3831 GND.n3830 2.56838
R4714 GND.n3508 GND.n3507 2.56838
R4715 GND.n1960 GND.n1959 2.56838
R4716 GND.n2069 GND.n2068 2.56838
R4717 GND.n2435 GND.n2434 2.56838
R4718 GND.n4688 GND.n4687 2.56838
R4719 GND.n4561 GND.t1487 2.36824
R4720 GND.n4562 GND.t658 2.36824
R4721 GND.n7822 GND.n7821 2.25932
R4722 GND.n978 GND.n977 2.25932
R4723 GND.n6104 GND.n6103 2.25932
R4724 GND.n3377 GND.n3376 1.93119
R4725 GND.n3376 GND.n3375 1.93119
R4726 GND.n3113 GND.n3112 1.93119
R4727 GND.n3112 GND.n3111 1.93119
R4728 GND.n4036 GND.n4035 1.93119
R4729 GND.n4035 GND.n4034 1.93119
R4730 GND.n5191 GND.n5190 1.93119
R4731 GND.n5190 GND.n5189 1.93119
R4732 GND.n3790 GND.n3789 1.93119
R4733 GND.n3789 GND.n3788 1.93119
R4734 GND.n1325 GND.n1324 1.93119
R4735 GND.n1324 GND.n1323 1.93119
R4736 GND.n3468 GND.n3467 1.93119
R4737 GND.n3467 GND.n3466 1.93119
R4738 GND.n1493 GND.n1492 1.93119
R4739 GND.n1492 GND.n1491 1.93119
R4740 GND.n1919 GND.n1918 1.93119
R4741 GND.n1918 GND.n1917 1.93119
R4742 GND.n142 GND.n141 1.93119
R4743 GND.n141 GND.n140 1.93119
R4744 GND.n2170 GND.n2169 1.93119
R4745 GND.n2169 GND.n2168 1.93119
R4746 GND.n2232 GND.n2231 1.93119
R4747 GND.n2231 GND.n2230 1.93119
R4748 GND.n2395 GND.n2394 1.93119
R4749 GND.n2394 GND.n2393 1.93119
R4750 GND.n2689 GND.n2688 1.93119
R4751 GND.n2688 GND.n2687 1.93119
R4752 GND.n4848 GND.n4847 1.93119
R4753 GND.n4847 GND.n4846 1.93119
R4754 GND.n4641 GND.n4640 1.93119
R4755 GND.n4640 GND.n4639 1.93119
R4756 GND.n4089 GND.n4088 1.85757
R4757 GND.n2115 GND.n2112 1.81868
R4758 GND.n4856 GND.n305 1.71871
R4759 GND.n2711 GND.n2656 1.71871
R4760 GND.n3137 GND.n3082 1.71871
R4761 GND.n7745 GND.n7744 1.71871
R4762 GND.n5441 GND.n5440 1.71871
R4763 GND.n4060 GND.n499 1.71871
R4764 GND.n5198 GND.n5143 1.71871
R4765 GND.n3798 GND.n3743 1.71871
R4766 GND.n3475 GND.n3420 1.71871
R4767 GND.n2402 GND.n2347 1.71871
R4768 GND.n3395 GND.n3353 1.71871
R4769 GND.n4576 GND.n4575 1.70717
R4770 GND.n3233 GND.n3232 1.64041
R4771 GND.n2892 GND.n2891 1.64041
R4772 GND.n2336 GND.n2335 1.64041
R4773 GND.n7739 GND.n7738 1.64041
R4774 GND.n1595 GND.n1594 1.64041
R4775 GND.n5435 GND.n5434 1.64041
R4776 GND.n4002 GND.n4001 1.64041
R4777 GND.n5300 GND.n5299 1.64041
R4778 GND.n3890 GND.n3889 1.64041
R4779 GND.n3563 GND.n3562 1.64041
R4780 GND.n2022 GND.n2021 1.64041
R4781 GND.n2120 GND.n2119 1.64041
R4782 GND.n2490 GND.n2489 1.64041
R4783 GND.n4947 GND.n4946 1.64041
R4784 GND.n3232 GND.n3231 1.63319
R4785 GND.n2891 GND.n2890 1.63319
R4786 GND.n4001 GND.n4000 1.63319
R4787 GND.n5299 GND.n5298 1.63319
R4788 GND.n3889 GND.n3888 1.63319
R4789 GND.n5434 GND.n5433 1.63319
R4790 GND.n3562 GND.n3561 1.63319
R4791 GND.n1594 GND.n1593 1.63319
R4792 GND.n2021 GND.n2020 1.63319
R4793 GND.n7738 GND.n7737 1.63319
R4794 GND.n2119 GND.n2118 1.63319
R4795 GND.n2335 GND.n2334 1.63319
R4796 GND.n2489 GND.n2488 1.63319
R4797 GND.n4946 GND.n4945 1.63319
R4798 GND.n4273 GND.n4272 1.49383
R4799 GND.n7436 GND 1.48176
R4800 GND.n4103 GND.n4101 1.40675
R4801 GND.n4099 GND.n4075 1.40675
R4802 GND.n4086 GND.n4084 1.3822
R4803 GND.n4092 GND.n4091 1.3822
R4804 GND.n4590 GND.n4475 1.2805
R4805 GND.n4468 GND.n4467 1.2805
R4806 GND.n565 GND.n564 1.12991
R4807 GND.n7391 GND.n7390 1.12991
R4808 GND.n7344 GND.n7343 1.12991
R4809 GND.n7321 GND.n7320 1.12991
R4810 GND.n7259 GND.n7258 1.12991
R4811 GND.n3335 GND.n3334 1.12991
R4812 GND.n7522 GND.n7521 1.12991
R4813 GND.n7584 GND.n7583 1.12991
R4814 GND.n2638 GND.n2637 1.12991
R4815 GND.n3064 GND.n3063 1.12991
R4816 GND.n6930 GND.n6929 1.12991
R4817 GND.n6807 GND.n6806 1.12991
R4818 GND.n55 GND.n54 1.12991
R4819 GND.n1000 GND.n999 1.12991
R4820 GND.n1229 GND.n1228 1.12991
R4821 GND.n7460 GND.n7459 1.12991
R4822 GND.n5125 GND.n5124 1.12991
R4823 GND.n3725 GND.n3724 1.12991
R4824 GND.n5496 GND.n5495 1.12991
R4825 GND.n6517 GND.n6516 1.12991
R4826 GND.n7091 GND.n7090 1.12991
R4827 GND.n5785 GND.n5784 1.12991
R4828 GND.n5714 GND.n5713 1.12991
R4829 GND.n6144 GND.n6143 1.12991
R4830 GND.n6197 GND.n6196 1.12991
R4831 GND.n5836 GND.n5835 1.12991
R4832 GND.n953 GND.n952 1.12991
R4833 GND.n883 GND.n882 1.12991
R4834 GND.n854 GND.n853 1.12991
R4835 GND.n790 GND.n789 1.12991
R4836 GND.n756 GND.n755 1.12991
R4837 GND.n6079 GND.n6078 1.12991
R4838 GND.n6031 GND.n6030 1.12991
R4839 GND.n5973 GND.n5972 1.12991
R4840 GND.n5950 GND.n5949 1.12991
R4841 GND.n5888 GND.n5887 1.12991
R4842 GND.n2916 GND.n2893 1.10214
R4843 GND.n4766 GND.n4738 1.10164
R4844 GND.n4949 GND.n4948 1.10116
R4845 GND.n3235 GND.n3234 1.10116
R4846 GND.n2338 GND.n2337 1.10116
R4847 GND.n2122 GND.n2121 1.10116
R4848 GND.n7741 GND.n7740 1.10116
R4849 GND.n1597 GND.n1596 1.10116
R4850 GND.n5437 GND.n5436 1.10116
R4851 GND.n4004 GND.n4003 1.10116
R4852 GND.n5302 GND.n5301 1.10116
R4853 GND.n3892 GND.n3891 1.10116
R4854 GND.n3565 GND.n3564 1.10116
R4855 GND.n2024 GND.n2023 1.10116
R4856 GND.n2492 GND.n2491 1.10116
R4857 GND.n2807 GND.n2784 1.10114
R4858 GND.n3977 GND.n3976 0.9605
R4859 GND.n4721 GND.n4720 0.9605
R4860 GND.n4717 GND.n4709 0.9605
R4861 GND.n3185 GND.n3184 0.9605
R4862 GND.n3189 GND.n3188 0.9605
R4863 GND.n2867 GND.n2866 0.9605
R4864 GND.n2875 GND.n2874 0.9605
R4865 GND.n2317 GND.n2316 0.9605
R4866 GND.n2319 GND.n2318 0.9605
R4867 GND.n7722 GND.n7721 0.9605
R4868 GND.n1578 GND.n1577 0.9605
R4869 GND.n5414 GND.n5413 0.9605
R4870 GND.n5418 GND.n5417 0.9605
R4871 GND.n3984 GND.n3983 0.9605
R4872 GND.n5275 GND.n5274 0.9605
R4873 GND.n5283 GND.n5282 0.9605
R4874 GND.n3872 GND.n3871 0.9605
R4875 GND.n2005 GND.n2004 0.9605
R4876 GND.n2094 GND.n2093 0.9605
R4877 GND.n122 GND.n121 0.9605
R4878 GND.n2766 GND.n2765 0.9605
R4879 GND.n4930 GND.n4929 0.9605
R4880 GND.n2964 GND.n2963 0.932703
R4881 GND.n3001 GND.t1152 0.932703
R4882 GND.n2540 GND.n2539 0.932703
R4883 GND.n2575 GND.t1167 0.932703
R4884 GND.n7145 GND.n7144 0.932703
R4885 GND.n7175 GND.t363 0.932703
R4886 GND.n608 GND.n607 0.932703
R4887 GND.n7012 GND.t853 0.932703
R4888 GND.n618 GND.n617 0.932703
R4889 GND.n6858 GND.t1411 0.932703
R4890 GND.n628 GND.n627 0.932703
R4891 GND.n6704 GND.t359 0.932703
R4892 GND.n635 GND.n634 0.932703
R4893 GND.n6633 GND.t1386 0.932703
R4894 GND.n5614 GND.n5613 0.932703
R4895 GND.n5585 GND.t261 0.932703
R4896 GND.n5479 GND.n5478 0.932703
R4897 GND.n1083 GND.t265 0.932703
R4898 GND.n1136 GND.n1135 0.932703
R4899 GND.n1204 GND.t313 0.932703
R4900 GND.n3628 GND.n3627 0.932703
R4901 GND.n3665 GND.t881 0.932703
R4902 GND.n5022 GND.n5021 0.932703
R4903 GND.n5062 GND.t248 0.932703
R4904 GND.n417 GND.n416 0.932703
R4905 GND.n457 GND.t543 0.932703
R4906 GND.n313 GND.n312 0.932703
R4907 GND.n388 GND.t1424 0.932703
R4908 GND.n211 GND.n210 0.932703
R4909 GND.n284 GND.t557 0.932703
R4910 GND.n4967 GND.n4966 0.795683
R4911 GND.n1854 GND.n1853 0.795683
R4912 GND.n1848 GND.n1847 0.795683
R4913 GND.n1851 GND.n1850 0.795683
R4914 GND.n1860 GND.n1859 0.795683
R4915 GND.n1871 GND.n1870 0.795683
R4916 GND.n5324 GND.n5323 0.795683
R4917 GND.n3581 GND.n3580 0.795683
R4918 GND.n5320 GND.n5319 0.795683
R4919 GND.n3905 GND.n3904 0.795683
R4920 GND.n3902 GND.n3901 0.795683
R4921 GND.n3575 GND.n3574 0.795683
R4922 GND.n3418 GND.n3417 0.795683
R4923 GND.n1863 GND.n1862 0.795683
R4924 GND.n1857 GND.n1856 0.795683
R4925 GND.n1847 GND.n1846 0.795337
R4926 GND.n1850 GND.n1849 0.795337
R4927 GND.n1853 GND.n1852 0.795337
R4928 GND.n1856 GND.n1855 0.795337
R4929 GND.n1859 GND.n1858 0.795337
R4930 GND.n1862 GND.n1861 0.795337
R4931 GND.n1870 GND.n1869 0.795337
R4932 GND.n3417 GND.n3416 0.795337
R4933 GND.n5323 GND.n5322 0.795337
R4934 GND.n3574 GND.n3573 0.795337
R4935 GND.n3580 GND.n3579 0.795337
R4936 GND.n3901 GND.n3900 0.795337
R4937 GND.n3904 GND.n3903 0.795337
R4938 GND.n5319 GND.n5318 0.795337
R4939 GND.n4966 GND.n4965 0.795337
R4940 GND.n4963 GND.n4962 0.795337
R4941 GND.n4964 GND.n4963 0.795337
R4942 GND.n5661 GND.n5660 0.705542
R4943 GND.n7436 GND.n7435 0.701583
R4944 GND.n4560 GND.n4558 0.6255
R4945 GND.n4567 GND.n4566 0.6255
R4946 GND.n4482 GND.n4480 0.614587
R4947 GND.n4574 GND.n4573 0.614587
R4948 GND.n4081 GND.n4080 0.549071
R4949 GND.n2620 GND.n2619 0.533636
R4950 GND.n3046 GND.n3045 0.533636
R4951 GND.n6987 GND.n6986 0.533636
R4952 GND.n6833 GND.n6832 0.533636
R4953 GND.n6669 GND.n6668 0.533636
R4954 GND.n501 GND.n498 0.533636
R4955 GND.n5107 GND.n5106 0.533636
R4956 GND.n3707 GND.n3706 0.533636
R4957 GND.n7224 GND.n7223 0.533636
R4958 GND.n3318 GND.n3317 0.533636
R4959 GND.n6138 GND.n5850 0.53211
R4960 GND.n4951 GND.n4950 0.520438
R4961 GND.n4768 GND.n4767 0.520438
R4962 GND.n3396 GND.n3236 0.520438
R4963 GND.n2340 GND.n2339 0.520438
R4964 GND.n7743 GND.n7742 0.520438
R4965 GND.n1599 GND.n1598 0.520438
R4966 GND.n5439 GND.n5438 0.520438
R4967 GND.n4061 GND.n4005 0.520438
R4968 GND.n5304 GND.n5303 0.520438
R4969 GND.n3894 GND.n3893 0.520438
R4970 GND.n3567 GND.n3566 0.520438
R4971 GND.n2026 GND.n2025 0.520438
R4972 GND.n2179 GND.n2123 0.520438
R4973 GND.n2494 GND.n2493 0.520438
R4974 GND.n2809 GND.n2808 0.520438
R4975 GND.n3138 GND.n2917 0.520438
R4976 GND.n7136 GND.n7135 0.498714
R4977 GND.n6918 GND.n611 0.498714
R4978 GND.n6764 GND.n621 0.498714
R4979 GND.n7072 GND.n601 0.498714
R4980 GND.n6136 GND.n6135 0.48654
R4981 GND.n856 GND.n542 0.479239
R4982 GND.n3362 GND.n3361 0.436742
R4983 GND.n3361 GND.n3360 0.436742
R4984 GND.n3094 GND.n3093 0.436742
R4985 GND.n3093 GND.n3092 0.436742
R4986 GND.n4017 GND.n4016 0.436742
R4987 GND.n4016 GND.n4015 0.436742
R4988 GND.n5156 GND.n5155 0.436742
R4989 GND.n5155 GND.n5154 0.436742
R4990 GND.n3755 GND.n3754 0.436742
R4991 GND.n3754 GND.n3753 0.436742
R4992 GND.n1290 GND.n1289 0.436742
R4993 GND.n1289 GND.n1288 0.436742
R4994 GND.n3433 GND.n3432 0.436742
R4995 GND.n3432 GND.n3431 0.436742
R4996 GND.n1458 GND.n1457 0.436742
R4997 GND.n1457 GND.n1456 0.436742
R4998 GND.n1884 GND.n1883 0.436742
R4999 GND.n1883 GND.n1882 0.436742
R5000 GND.n99 GND.n98 0.436742
R5001 GND.n98 GND.n97 0.436742
R5002 GND.n2135 GND.n2134 0.436742
R5003 GND.n2134 GND.n2133 0.436742
R5004 GND.n2197 GND.n2196 0.436742
R5005 GND.n2196 GND.n2195 0.436742
R5006 GND.n2360 GND.n2359 0.436742
R5007 GND.n2359 GND.n2358 0.436742
R5008 GND.n2672 GND.n2671 0.436742
R5009 GND.n2671 GND.n2670 0.436742
R5010 GND.n4813 GND.n4812 0.436742
R5011 GND.n4812 GND.n4811 0.436742
R5012 GND.n4606 GND.n4605 0.436742
R5013 GND.n4605 GND.n4604 0.436742
R5014 GND.n4477 GND.n4476 0.427167
R5015 GND.n4283 GND.n4282 0.427167
R5016 GND.n3270 GND.n3269 0.425574
R5017 GND.n7566 GND.n7565 0.425574
R5018 GND.n201 GND.n200 0.425574
R5019 GND.n2950 GND.n2949 0.425574
R5020 GND.n6659 GND.n6658 0.425574
R5021 GND.n5521 GND.n5520 0.425574
R5022 GND.n1269 GND.n1268 0.425574
R5023 GND.n7504 GND.n7503 0.425574
R5024 GND.n5009 GND.n5008 0.425574
R5025 GND.n3615 GND.n3614 0.425574
R5026 GND.n5464 GND.n5463 0.425574
R5027 GND.n5643 GND.n5642 0.425574
R5028 GND.n7801 GND.n7800 0.414845
R5029 GND.n6379 GND.n6378 0.414845
R5030 GND.n393 GND.n376 0.38056
R5031 GND.n289 GND.n272 0.38056
R5032 GND.n2580 GND.n2563 0.38056
R5033 GND.n3006 GND.n2989 0.38056
R5034 GND.n7017 GND.n7000 0.38056
R5035 GND.n6863 GND.n6846 0.38056
R5036 GND.n6709 GND.n6692 0.38056
R5037 GND.n5590 GND.n5573 0.38056
R5038 GND.n1209 GND.n1192 0.38056
R5039 GND.n462 GND.n445 0.38056
R5040 GND.n5067 GND.n5050 0.38056
R5041 GND.n3670 GND.n3653 0.38056
R5042 GND.n1088 GND.n1071 0.38056
R5043 GND.n6638 GND.n6621 0.38056
R5044 GND.n7180 GND.n7163 0.38056
R5045 GND.n3309 GND.n3297 0.38056
R5046 GND.n4951 GND.n4856 0.378813
R5047 GND.n4768 GND.n4649 0.378813
R5048 GND.n2809 GND.n2711 0.378813
R5049 GND.n3138 GND.n3137 0.378813
R5050 GND.n2340 GND.n2240 0.378813
R5051 GND.n2179 GND.n2178 0.378813
R5052 GND.n7744 GND.n7743 0.378813
R5053 GND.n1599 GND.n1500 0.378813
R5054 GND.n5440 GND.n5439 0.378813
R5055 GND.n4061 GND.n4060 0.378813
R5056 GND.n5304 GND.n5198 0.378813
R5057 GND.n3894 GND.n3798 0.378813
R5058 GND.n3567 GND.n3475 0.378813
R5059 GND.n2026 GND.n1927 0.378813
R5060 GND.n2494 GND.n2402 0.378813
R5061 GND.n3396 GND.n3395 0.378813
R5062 GND.n365 GND.n363 0.377583
R5063 GND.n261 GND.n259 0.377583
R5064 GND.n2552 GND.n2550 0.377583
R5065 GND.n2978 GND.n2976 0.377583
R5066 GND.n6681 GND.n6679 0.377583
R5067 GND.n5562 GND.n5560 0.377583
R5068 GND.n1181 GND.n1179 0.377583
R5069 GND.n434 GND.n432 0.377583
R5070 GND.n5039 GND.n5037 0.377583
R5071 GND.n3642 GND.n3640 0.377583
R5072 GND.n1060 GND.n1058 0.377583
R5073 GND.n6610 GND.n6608 0.377583
R5074 GND.n3286 GND.n3284 0.377583
R5075 GND.n7381 GND.n7380 0.376971
R5076 GND.n7428 GND.n7427 0.376971
R5077 GND.n7333 GND.n7332 0.376971
R5078 GND.n7249 GND.n7248 0.376971
R5079 GND.n3330 GND.n3329 0.376971
R5080 GND.n7517 GND.n7516 0.376971
R5081 GND.n7579 GND.n7578 0.376971
R5082 GND.n2633 GND.n2632 0.376971
R5083 GND.n3059 GND.n3058 0.376971
R5084 GND.n6927 GND.n6926 0.376971
R5085 GND.n6773 GND.n6772 0.376971
R5086 GND.n7757 GND.n7756 0.376971
R5087 GND.n997 GND.n996 0.376971
R5088 GND.n1226 GND.n1225 0.376971
R5089 GND.n7455 GND.n7454 0.376971
R5090 GND.n5120 GND.n5119 0.376971
R5091 GND.n3720 GND.n3719 0.376971
R5092 GND.n1105 GND.n1104 0.376971
R5093 GND.n6508 GND.n6507 0.376971
R5094 GND.n7086 GND.n7085 0.376971
R5095 GND.n5821 GND.n5820 0.376971
R5096 GND.n5775 GND.n5774 0.376971
R5097 GND.n5726 GND.n5725 0.376971
R5098 GND.n6157 GND.n6156 0.376971
R5099 GND.n5664 GND.n5663 0.376971
R5100 GND.n709 GND.n708 0.376971
R5101 GND.n867 GND.n866 0.376971
R5102 GND.n780 GND.n779 0.376971
R5103 GND.n768 GND.n767 0.376971
R5104 GND.n6043 GND.n6042 0.376971
R5105 GND.n6129 GND.n6128 0.376971
R5106 GND.n5962 GND.n5961 0.376971
R5107 GND.n5878 GND.n5877 0.376971
R5108 GND.n7799 GND.n7798 0.375505
R5109 GND.n6380 GND.n6351 0.375505
R5110 GND.n361 GND.n358 0.3755
R5111 GND.n257 GND.n254 0.3755
R5112 GND.n2974 GND.n2971 0.3755
R5113 GND.n6880 GND.n6878 0.3755
R5114 GND.n6726 GND.n6724 0.3755
R5115 GND.n6677 GND.n6674 0.3755
R5116 GND.n5558 GND.n5555 0.3755
R5117 GND.n1177 GND.n1174 0.3755
R5118 GND.n430 GND.n427 0.3755
R5119 GND.n5035 GND.n5032 0.3755
R5120 GND.n3638 GND.n3635 0.3755
R5121 GND.n1056 GND.n1053 0.3755
R5122 GND.n6606 GND.n6603 0.3755
R5123 GND.n7034 GND.n7032 0.3755
R5124 GND.n3282 GND.n3279 0.3755
R5125 GND.n233 GND.n231 0.373417
R5126 GND.n7640 GND.n7638 0.373417
R5127 GND.n7200 GND.n7198 0.373417
R5128 GND.n7198 GND.n7197 0.373417
R5129 GND.n2596 GND.n2594 0.373417
R5130 GND.n2594 GND.n2593 0.373417
R5131 GND.n6888 GND.n6886 0.373417
R5132 GND.n6886 GND.n6885 0.373417
R5133 GND.n6734 GND.n6732 0.373417
R5134 GND.n6732 GND.n6731 0.373417
R5135 GND.n6575 GND.n6573 0.373417
R5136 GND.n6573 GND.n6572 0.373417
R5137 GND.n5550 GND.n5548 0.373417
R5138 GND.n3683 GND.n3681 0.373417
R5139 GND.n3681 GND.n3680 0.373417
R5140 GND.n337 GND.n335 0.373417
R5141 GND.n335 GND.n334 0.373417
R5142 GND.n475 GND.n473 0.373417
R5143 GND.n473 GND.n472 0.373417
R5144 GND.n5083 GND.n5081 0.373417
R5145 GND.n5081 GND.n5080 0.373417
R5146 GND.n1155 GND.n1153 0.373417
R5147 GND.n6598 GND.n6596 0.373417
R5148 GND.n7042 GND.n7040 0.373417
R5149 GND.n7040 GND.n7039 0.373417
R5150 GND.n3022 GND.n3020 0.373417
R5151 GND.n3020 GND.n3013 0.373417
R5152 GND.n3010 GND.n3009 0.366214
R5153 GND.n2590 GND.n2589 0.366214
R5154 GND.n7194 GND.n7193 0.366214
R5155 GND.n7036 GND.n7035 0.366214
R5156 GND.n6882 GND.n6881 0.366214
R5157 GND.n6728 GND.n6727 0.366214
R5158 GND.n6671 GND.n6670 0.366214
R5159 GND.n6600 GND.n6599 0.366214
R5160 GND.n5552 GND.n5551 0.366214
R5161 GND.n1050 GND.n1049 0.366214
R5162 GND.n1171 GND.n1170 0.366214
R5163 GND.n5077 GND.n5076 0.366214
R5164 GND.n5029 GND.n5028 0.366214
R5165 GND.n424 GND.n423 0.366214
R5166 GND.n355 GND.n354 0.366214
R5167 GND.n251 GND.n250 0.366214
R5168 GND.n2618 GND.n2617 0.355857
R5169 GND.n3044 GND.n3043 0.355857
R5170 GND.n7064 GND.n7063 0.355857
R5171 GND.n6910 GND.n6909 0.355857
R5172 GND.n6756 GND.n6755 0.355857
R5173 GND.n497 GND.n496 0.355857
R5174 GND.n5105 GND.n5104 0.355857
R5175 GND.n3705 GND.n3704 0.355857
R5176 GND.n7222 GND.n7221 0.355857
R5177 GND.n3316 GND.n3315 0.355857
R5178 GND.n4898 GND 0.354667
R5179 GND.n4697 GND 0.354667
R5180 GND.n3152 GND 0.354667
R5181 GND.n2821 GND 0.354667
R5182 GND.n2282 GND 0.354667
R5183 GND.n7686 GND 0.354667
R5184 GND.n1542 GND 0.354667
R5185 GND.n5379 GND 0.354667
R5186 GND.n3948 GND 0.354667
R5187 GND.n5240 GND 0.354667
R5188 GND.n3840 GND 0.354667
R5189 GND.n3517 GND 0.354667
R5190 GND.n1969 GND 0.354667
R5191 GND.n2056 GND 0.354667
R5192 GND.n2444 GND 0.354667
R5193 GND.n2753 GND 0.354667
R5194 GND.n4447 GND.n4064 0.352931
R5195 GND.n4434 GND.n4433 0.352931
R5196 GND.n4418 GND.n4417 0.352931
R5197 GND.n4403 GND.n4402 0.352931
R5198 GND.n4388 GND.n4387 0.352931
R5199 GND.n4373 GND.n4372 0.352931
R5200 GND.n4356 GND.n4355 0.352931
R5201 GND.n4341 GND.n4340 0.352931
R5202 GND.n4326 GND.n4325 0.352931
R5203 GND.n4311 GND.n4310 0.352931
R5204 GND.n4275 GND.n4274 0.352931
R5205 GND.n4257 GND.n4256 0.352931
R5206 GND.n4232 GND.n4231 0.352931
R5207 GND.n4217 GND.n4216 0.352931
R5208 GND.n4202 GND.n4201 0.352931
R5209 GND.n4187 GND.n4186 0.352931
R5210 GND.n4168 GND.n4167 0.352931
R5211 GND.n4153 GND.n4152 0.352931
R5212 GND.n4138 GND.n4137 0.352931
R5213 GND.n4123 GND.n4122 0.352931
R5214 GND.n4296 GND.n4295 0.347722
R5215 GND.n303 GND.n224 0.345738
R5216 GND.n7627 GND.n195 0.345738
R5217 GND.n6921 GND.n6918 0.345738
R5218 GND.n6767 GND.n6764 0.345738
R5219 GND.n6652 GND.n6564 0.345738
R5220 GND.n5470 GND.n1102 0.345738
R5221 GND.n407 GND.n326 0.345738
R5222 GND.n1223 GND.n1146 0.345738
R5223 GND.n5605 GND.n5604 0.345738
R5224 GND.n7075 GND.n7072 0.345738
R5225 GND.n7794 GND.n50 0.33677
R5226 GND.n6381 GND.n6329 0.33677
R5227 GND.n6137 GND.n6136 0.336652
R5228 GND.n6454 GND 0.327423
R5229 GND.n539 GND 0.327423
R5230 GND.n6498 GND.n6497 0.326891
R5231 GND.n6407 GND.n6295 0.326891
R5232 GND.n6471 GND.n6470 0.325812
R5233 GND.n6409 GND.n6408 0.325812
R5234 GND.n4902 GND.n4901 0.321569
R5235 GND.n4678 GND.n4670 0.321569
R5236 GND.n4701 GND.n4700 0.321569
R5237 GND.n3157 GND.n3156 0.321569
R5238 GND.n3207 GND.n3206 0.321569
R5239 GND.n2861 GND.n2824 0.321569
R5240 GND.n2286 GND.n2285 0.321569
R5241 GND.n2254 GND.n2242 0.321569
R5242 GND.n7690 GND.n7689 0.321569
R5243 GND.n7669 GND.n7667 0.321569
R5244 GND.n1546 GND.n1545 0.321569
R5245 GND.n1514 GND.n1502 0.321569
R5246 GND.n5383 GND.n5382 0.321569
R5247 GND.n5351 GND.n5339 0.321569
R5248 GND.n3952 GND.n3951 0.321569
R5249 GND.n3920 GND.n3908 0.321569
R5250 GND.n5244 GND.n5243 0.321569
R5251 GND.n5212 GND.n5200 0.321569
R5252 GND.n3844 GND.n3843 0.321569
R5253 GND.n3812 GND.n3800 0.321569
R5254 GND.n3521 GND.n3520 0.321569
R5255 GND.n3489 GND.n3477 0.321569
R5256 GND.n1973 GND.n1972 0.321569
R5257 GND.n1941 GND.n1929 0.321569
R5258 GND.n2075 GND.n2059 0.321569
R5259 GND.n2052 GND.n2051 0.321569
R5260 GND.n2448 GND.n2447 0.321569
R5261 GND.n2416 GND.n2404 0.321569
R5262 GND.n2725 GND.n2713 0.321569
R5263 GND.n2757 GND.n2756 0.321569
R5264 GND.n4870 GND.n4858 0.321569
R5265 GND.n2835 GND.n2817 0.321569
R5266 GND.n358 GND.n353 0.321333
R5267 GND.n254 GND.n249 0.321333
R5268 GND.n7197 GND.n7192 0.321333
R5269 GND.n6885 GND.n6880 0.321333
R5270 GND.n6731 GND.n6726 0.321333
R5271 GND.n5555 GND.n5550 0.321333
R5272 GND.n1053 GND.n1048 0.321333
R5273 GND.n6603 GND.n6598 0.321333
R5274 GND.n7039 GND.n7034 0.321333
R5275 GND.n4471 GND.n4468 0.3205
R5276 GND.n6138 GND.n6137 0.31982
R5277 GND.n4950 GND.n4903 0.314812
R5278 GND.n4767 GND.n4702 0.314812
R5279 GND.n3236 GND.n3158 0.314812
R5280 GND.n2339 GND.n2287 0.314812
R5281 GND.n7742 GND.n7691 0.314812
R5282 GND.n1598 GND.n1547 0.314812
R5283 GND.n5438 GND.n5384 0.314812
R5284 GND.n4005 GND.n3953 0.314812
R5285 GND.n5303 GND.n5245 0.314812
R5286 GND.n3893 GND.n3845 0.314812
R5287 GND.n3566 GND.n3522 0.314812
R5288 GND.n2025 GND.n1974 0.314812
R5289 GND.n2123 GND.n2076 0.314812
R5290 GND.n2493 GND.n2449 0.314812
R5291 GND.n2808 GND.n2758 0.314812
R5292 GND.n2917 GND.n2862 0.314812
R5293 GND.n247 GND.n244 0.313
R5294 GND.n7654 GND.n7651 0.313
R5295 GND.n7214 GND.n7211 0.313
R5296 GND.n2610 GND.n2607 0.313
R5297 GND.n6902 GND.n6899 0.313
R5298 GND.n6748 GND.n6745 0.313
R5299 GND.n6589 GND.n6586 0.313
R5300 GND.n1046 GND.n1043 0.313
R5301 GND.n3697 GND.n3694 0.313
R5302 GND.n351 GND.n348 0.313
R5303 GND.n489 GND.n486 0.313
R5304 GND.n5097 GND.n5094 0.313
R5305 GND.n1169 GND.n1166 0.313
R5306 GND.n5541 GND.n5538 0.313
R5307 GND.n7056 GND.n7053 0.313
R5308 GND.n3036 GND.n3033 0.313
R5309 GND.n7435 GND.n542 0.309146
R5310 GND.n4450 GND.n4447 0.302583
R5311 GND.n321 GND.n317 0.300798
R5312 GND.n219 GND.n215 0.300798
R5313 GND.n5617 GND.n5525 0.300798
R5314 GND.n1141 GND.n1140 0.300798
R5315 GND.n5482 GND.n5469 0.300798
R5316 GND.n6559 GND.n638 0.300798
R5317 GND GND.n49 0.295209
R5318 GND GND.n6376 0.295209
R5319 GND.n4898 GND.n4896 0.295052
R5320 GND.n4697 GND.n4695 0.295052
R5321 GND.n3152 GND.n3150 0.295052
R5322 GND.n2821 GND.n2819 0.295052
R5323 GND.n2282 GND.n2280 0.295052
R5324 GND.n7686 GND.n7684 0.295052
R5325 GND.n1542 GND.n1540 0.295052
R5326 GND.n5379 GND.n5377 0.295052
R5327 GND.n3948 GND.n3946 0.295052
R5328 GND.n5240 GND.n5238 0.295052
R5329 GND.n3840 GND.n3838 0.295052
R5330 GND.n3517 GND.n3515 0.295052
R5331 GND.n1969 GND.n1967 0.295052
R5332 GND.n2056 GND.n2054 0.295052
R5333 GND.n2444 GND.n2442 0.295052
R5334 GND.n2753 GND.n2751 0.295052
R5335 GND.n3277 GND.n3275 0.290381
R5336 GND.n321 GND.n320 0.290381
R5337 GND.n219 GND.n218 0.290381
R5338 GND.n2545 GND.n2543 0.290381
R5339 GND.n2969 GND.n2967 0.290381
R5340 GND.n7067 GND.n7066 0.290381
R5341 GND.n6913 GND.n6912 0.290381
R5342 GND.n6759 GND.n6758 0.290381
R5343 GND.n5619 GND.n5617 0.290381
R5344 GND.n422 GND.n420 0.290381
R5345 GND.n5027 GND.n5025 0.290381
R5346 GND.n3633 GND.n3631 0.290381
R5347 GND.n5484 GND.n5482 0.290381
R5348 GND.n6559 GND.n6558 0.290381
R5349 GND.n7150 GND.n7148 0.290381
R5350 GND.n7437 GND.n7436 0.283189
R5351 GND.n6136 GND.n542 0.282159
R5352 GND.n6496 GND.n6495 0.280127
R5353 GND.n6406 GND.n6405 0.280127
R5354 GND.n4578 GND.n4577 0.270108
R5355 GND.n1374 GND.n1373 0.260982
R5356 GND.n1373 GND.n1372 0.2605
R5357 GND.n3403 GND 0.246986
R5358 GND.n367 GND.n365 0.24425
R5359 GND.n263 GND.n261 0.24425
R5360 GND.n2554 GND.n2552 0.24425
R5361 GND.n2980 GND.n2978 0.24425
R5362 GND.n6991 GND.n6989 0.24425
R5363 GND.n6837 GND.n6835 0.24425
R5364 GND.n6683 GND.n6681 0.24425
R5365 GND.n5564 GND.n5562 0.24425
R5366 GND.n1183 GND.n1181 0.24425
R5367 GND.n436 GND.n434 0.24425
R5368 GND.n5041 GND.n5039 0.24425
R5369 GND.n3644 GND.n3642 0.24425
R5370 GND.n1062 GND.n1060 0.24425
R5371 GND.n6612 GND.n6610 0.24425
R5372 GND.n7154 GND.n7152 0.24425
R5373 GND.n3288 GND.n3286 0.24425
R5374 GND.n7564 GND.n7563 0.243155
R5375 GND.n7626 GND.n7625 0.243155
R5376 GND.n2530 GND.n2528 0.243155
R5377 GND.n2953 GND.n2951 0.243155
R5378 GND.n6924 GND.n6923 0.243155
R5379 GND.n6770 GND.n6769 0.243155
R5380 GND.n6662 GND.n6660 0.243155
R5381 GND.n5622 GND.n5522 0.243155
R5382 GND.n1275 GND.n1270 0.243155
R5383 GND.n7502 GND.n7501 0.243155
R5384 GND.n5012 GND.n5010 0.243155
R5385 GND.n3618 GND.n3616 0.243155
R5386 GND.n5487 GND.n5465 0.243155
R5387 GND.n6554 GND.n639 0.243155
R5388 GND.n7132 GND.n7077 0.243155
R5389 GND.n3272 GND.n3271 0.243155
R5390 GND.n235 GND.n233 0.238893
R5391 GND.n7642 GND.n7640 0.238893
R5392 GND.n7202 GND.n7200 0.238893
R5393 GND.n2598 GND.n2596 0.238893
R5394 GND.n6890 GND.n6888 0.238893
R5395 GND.n6736 GND.n6734 0.238893
R5396 GND.n6577 GND.n6575 0.238893
R5397 GND.n1034 GND.n1032 0.238893
R5398 GND.n3685 GND.n3683 0.238893
R5399 GND.n339 GND.n337 0.238893
R5400 GND.n477 GND.n475 0.238893
R5401 GND.n5085 GND.n5083 0.238893
R5402 GND.n1157 GND.n1155 0.238893
R5403 GND.n5529 GND.n5527 0.238893
R5404 GND.n7044 GND.n7042 0.238893
R5405 GND.n3024 GND.n3022 0.238893
R5406 GND.n5744 GND 0.228789
R5407 GND.n34 GND.n30 0.226583
R5408 GND.n6361 GND.n6357 0.226583
R5409 GND.n7561 GND.n7539 0.224247
R5410 GND.n7623 GND.n7601 0.224247
R5411 GND.n2655 GND.n2522 0.224247
R5412 GND.n3081 GND.n2939 0.224247
R5413 GND.n6964 GND.n6962 0.224247
R5414 GND.n6801 GND.n6799 0.224247
R5415 GND.n7746 GND.n87 0.224247
R5416 GND.n5626 GND.n5624 0.224247
R5417 GND.n5442 GND.n1277 0.224247
R5418 GND.n7499 GND.n7477 0.224247
R5419 GND.n5142 GND.n4998 0.224247
R5420 GND.n3742 GND.n3604 0.224247
R5421 GND.n5490 GND.n5489 0.224247
R5422 GND.n6552 GND.n6530 0.224247
R5423 GND.n7130 GND.n7108 0.224247
R5424 GND.n3352 GND.n3258 0.224247
R5425 GND.n5669 GND 0.209082
R5426 GND.n302 GND.n300 0.200996
R5427 GND.n7631 GND.n7629 0.200996
R5428 GND.n2944 GND.n2942 0.200996
R5429 GND.n6651 GND.n6649 0.200996
R5430 GND.n1101 GND.n1099 0.200996
R5431 GND.n1263 GND.n1261 0.200996
R5432 GND.n406 GND.n404 0.200996
R5433 GND.n5003 GND.n5001 0.200996
R5434 GND.n3609 GND.n3607 0.200996
R5435 GND.n1222 GND.n1220 0.200996
R5436 GND.n5603 GND.n5601 0.200996
R5437 GND.n3264 GND.n3262 0.200996
R5438 GND.n4666 GND.n4663 0.197423
R5439 GND.n3215 GND.n3195 0.197423
R5440 GND.n2262 GND.n2244 0.197423
R5441 GND.n7663 GND.n164 0.197423
R5442 GND.n1522 GND.n1504 0.197423
R5443 GND.n5359 GND.n5341 0.197423
R5444 GND.n3928 GND.n3910 0.197423
R5445 GND.n5220 GND.n5202 0.197423
R5446 GND.n3820 GND.n3802 0.197423
R5447 GND.n3497 GND.n3479 0.197423
R5448 GND.n1949 GND.n1931 0.197423
R5449 GND.n2047 GND.n2045 0.197423
R5450 GND.n2424 GND.n2406 0.197423
R5451 GND.n2733 GND.n2715 0.197423
R5452 GND.n4878 GND.n4860 0.197423
R5453 GND.n2843 GND.n2825 0.197423
R5454 GND.n4563 GND.n4562 0.196239
R5455 GND.n4564 GND.n4561 0.190273
R5456 GND.n7774 GND.n7771 0.189094
R5457 GND.n651 GND.n650 0.189094
R5458 GND.n6307 GND.n6304 0.189094
R5459 GND.n6279 GND.n6278 0.189094
R5460 GND.n4561 GND.n4062 0.188284
R5461 GND.n4593 GND.n4591 0.181849
R5462 GND.n3317 GND.n3316 0.181736
R5463 GND.n318 GND.n304 0.181736
R5464 GND.n216 GND.n202 0.181736
R5465 GND.n2619 GND.n2618 0.181736
R5466 GND.n3045 GND.n3044 0.181736
R5467 GND.n7064 GND.n6987 0.181736
R5468 GND.n6910 GND.n6833 0.181736
R5469 GND.n6756 GND.n6669 0.181736
R5470 GND.n5621 GND.n5620 0.181736
R5471 GND.n1274 GND.n1273 0.181736
R5472 GND.n498 GND.n497 0.181736
R5473 GND.n5106 GND.n5105 0.181736
R5474 GND.n3706 GND.n3705 0.181736
R5475 GND.n5486 GND.n5485 0.181736
R5476 GND.n6556 GND.n6555 0.181736
R5477 GND.n7223 GND.n7222 0.181736
R5478 GND.n4975 GND 0.180197
R5479 GND.n4974 GND 0.180197
R5480 GND.n3406 GND 0.180197
R5481 GND.n3408 GND 0.180197
R5482 GND.n5332 GND 0.180197
R5483 GND GND.n5336 0.180197
R5484 GND GND.n5312 0.180197
R5485 GND.n5311 GND 0.180197
R5486 GND GND.n1334 0.180197
R5487 GND.n5335 GND 0.180197
R5488 GND GND.n3410 0.180197
R5489 GND.n3407 GND 0.180197
R5490 GND.n3405 GND 0.180197
R5491 GND.n3404 GND 0.180197
R5492 GND.n3403 GND 0.180197
R5493 GND.n3317 GND.n3272 0.17675
R5494 GND.n7563 GND.n304 0.17675
R5495 GND.n7625 GND.n202 0.17675
R5496 GND.n2619 GND.n2530 0.17675
R5497 GND.n3045 GND.n2953 0.17675
R5498 GND.n6987 GND.n6924 0.17675
R5499 GND.n6833 GND.n6770 0.17675
R5500 GND.n6669 GND.n6662 0.17675
R5501 GND.n5622 GND.n5621 0.17675
R5502 GND.n1275 GND.n1274 0.17675
R5503 GND.n7501 GND.n498 0.17675
R5504 GND.n5106 GND.n5012 0.17675
R5505 GND.n3706 GND.n3618 0.17675
R5506 GND.n5487 GND.n5486 0.17675
R5507 GND.n6555 GND.n6554 0.17675
R5508 GND.n7223 GND.n7132 0.17675
R5509 GND.t1568 GND.t1072 0.176207
R5510 GND.n4096 GND.n4078 0.176207
R5511 GND.n369 GND.n367 0.171333
R5512 GND.n265 GND.n263 0.171333
R5513 GND.n2556 GND.n2554 0.171333
R5514 GND.n2982 GND.n2980 0.171333
R5515 GND.n6993 GND.n6991 0.171333
R5516 GND.n6839 GND.n6837 0.171333
R5517 GND.n6685 GND.n6683 0.171333
R5518 GND.n5566 GND.n5564 0.171333
R5519 GND.n1185 GND.n1183 0.171333
R5520 GND.n438 GND.n436 0.171333
R5521 GND.n5043 GND.n5041 0.171333
R5522 GND.n3646 GND.n3644 0.171333
R5523 GND.n1064 GND.n1062 0.171333
R5524 GND.n6614 GND.n6612 0.171333
R5525 GND.n7156 GND.n7154 0.171333
R5526 GND.n3290 GND.n3288 0.171333
R5527 GND.n376 GND.n373 0.16925
R5528 GND.n272 GND.n269 0.16925
R5529 GND.n2563 GND.n2560 0.16925
R5530 GND.n2989 GND.n2986 0.16925
R5531 GND.n7000 GND.n6997 0.16925
R5532 GND.n6846 GND.n6843 0.16925
R5533 GND.n6692 GND.n6689 0.16925
R5534 GND.n5573 GND.n5570 0.16925
R5535 GND.n1192 GND.n1189 0.16925
R5536 GND.n445 GND.n442 0.16925
R5537 GND.n5050 GND.n5047 0.16925
R5538 GND.n3653 GND.n3650 0.16925
R5539 GND.n1071 GND.n1068 0.16925
R5540 GND.n6621 GND.n6618 0.16925
R5541 GND.n7163 GND.n7160 0.16925
R5542 GND.n3297 GND.n3294 0.16925
R5543 GND.n541 GND 0.165163
R5544 GND.n300 GND.n298 0.164786
R5545 GND.n298 GND.n247 0.164786
R5546 GND.n7655 GND.n7631 0.164786
R5547 GND.n7655 GND.n7654 0.164786
R5548 GND.n7215 GND.n7184 0.164786
R5549 GND.n7215 GND.n7214 0.164786
R5550 GND.n2611 GND.n2610 0.164786
R5551 GND.n6903 GND.n6867 0.164786
R5552 GND.n6903 GND.n6902 0.164786
R5553 GND.n6749 GND.n6713 0.164786
R5554 GND.n6749 GND.n6748 0.164786
R5555 GND.n6649 GND.n6647 0.164786
R5556 GND.n6647 GND.n6589 0.164786
R5557 GND.n1099 GND.n1097 0.164786
R5558 GND.n1097 GND.n1046 0.164786
R5559 GND.n3698 GND.n3697 0.164786
R5560 GND.n404 GND.n402 0.164786
R5561 GND.n402 GND.n351 0.164786
R5562 GND.n490 GND.n489 0.164786
R5563 GND.n5098 GND.n5097 0.164786
R5564 GND.n1220 GND.n1218 0.164786
R5565 GND.n1218 GND.n1169 0.164786
R5566 GND.n5601 GND.n5599 0.164786
R5567 GND.n5599 GND.n5541 0.164786
R5568 GND.n7057 GND.n7021 0.164786
R5569 GND.n7057 GND.n7056 0.164786
R5570 GND.n3037 GND.n3036 0.164786
R5571 GND.n395 GND.n393 0.159429
R5572 GND.n291 GND.n289 0.159429
R5573 GND.n2582 GND.n2580 0.159429
R5574 GND.n3008 GND.n3006 0.159429
R5575 GND.n7019 GND.n7017 0.159429
R5576 GND.n6865 GND.n6863 0.159429
R5577 GND.n6711 GND.n6709 0.159429
R5578 GND.n5592 GND.n5590 0.159429
R5579 GND.n1211 GND.n1209 0.159429
R5580 GND.n464 GND.n462 0.159429
R5581 GND.n5069 GND.n5067 0.159429
R5582 GND.n3672 GND.n3670 0.159429
R5583 GND.n1090 GND.n1088 0.159429
R5584 GND.n6640 GND.n6638 0.159429
R5585 GND.n7182 GND.n7180 0.159429
R5586 GND.n3311 GND.n3309 0.159429
R5587 GND.n6454 GND.n6453 0.15606
R5588 GND.n539 GND.n538 0.15606
R5589 GND.n244 GND.n241 0.148714
R5590 GND.n239 GND.n235 0.148714
R5591 GND.n7651 GND.n7648 0.148714
R5592 GND.n7646 GND.n7642 0.148714
R5593 GND.n7211 GND.n7208 0.148714
R5594 GND.n7206 GND.n7202 0.148714
R5595 GND.n2607 GND.n2604 0.148714
R5596 GND.n2602 GND.n2598 0.148714
R5597 GND.n6899 GND.n6896 0.148714
R5598 GND.n6894 GND.n6890 0.148714
R5599 GND.n6745 GND.n6742 0.148714
R5600 GND.n6740 GND.n6736 0.148714
R5601 GND.n6586 GND.n6583 0.148714
R5602 GND.n6581 GND.n6577 0.148714
R5603 GND.n1043 GND.n1040 0.148714
R5604 GND.n1038 GND.n1034 0.148714
R5605 GND.n3694 GND.n3691 0.148714
R5606 GND.n3689 GND.n3685 0.148714
R5607 GND.n348 GND.n345 0.148714
R5608 GND.n343 GND.n339 0.148714
R5609 GND.n486 GND.n483 0.148714
R5610 GND.n481 GND.n477 0.148714
R5611 GND.n5094 GND.n5091 0.148714
R5612 GND.n5089 GND.n5085 0.148714
R5613 GND.n1166 GND.n1163 0.148714
R5614 GND.n1161 GND.n1157 0.148714
R5615 GND.n5538 GND.n5535 0.148714
R5616 GND.n5533 GND.n5529 0.148714
R5617 GND.n7053 GND.n7050 0.148714
R5618 GND.n7048 GND.n7044 0.148714
R5619 GND.n3033 GND.n3030 0.148714
R5620 GND.n3028 GND.n3024 0.148714
R5621 GND.n4594 GND.n4062 0.148287
R5622 GND.n4953 GND.n4801 0.142154
R5623 GND.n4972 GND.n4971 0.142154
R5624 GND.n3401 GND.n3400 0.142154
R5625 GND.n3143 GND.n3142 0.142154
R5626 GND.n2345 GND.n2344 0.142154
R5627 GND.n1865 GND.n1864 0.142154
R5628 GND.n5329 GND.n5328 0.142154
R5629 GND.n1333 GND.n1332 0.142154
R5630 GND.n5314 GND.n3906 0.142154
R5631 GND.n5309 GND.n5308 0.142154
R5632 GND.n3896 GND.n3582 0.142154
R5633 GND.n3569 GND.n3419 0.142154
R5634 GND.n3412 GND.n1872 0.142154
R5635 GND.n2184 GND.n2183 0.142154
R5636 GND.n2499 GND.n2498 0.142154
R5637 GND.n2814 GND.n2813 0.142154
R5638 GND.n4442 GND.n4441 0.141472
R5639 GND.n4441 GND.n4439 0.141472
R5640 GND.n4439 GND.n4426 0.141472
R5641 GND.n4426 GND.n4424 0.141472
R5642 GND.n4424 GND.n4411 0.141472
R5643 GND.n4411 GND.n4409 0.141472
R5644 GND.n4409 GND.n4396 0.141472
R5645 GND.n4396 GND.n4394 0.141472
R5646 GND.n4394 GND.n4381 0.141472
R5647 GND.n4381 GND.n4379 0.141472
R5648 GND.n4364 GND.n4362 0.141472
R5649 GND.n4362 GND.n4349 0.141472
R5650 GND.n4349 GND.n4347 0.141472
R5651 GND.n4347 GND.n4334 0.141472
R5652 GND.n4334 GND.n4332 0.141472
R5653 GND.n4332 GND.n4319 0.141472
R5654 GND.n4319 GND.n4317 0.141472
R5655 GND.n4317 GND.n4304 0.141472
R5656 GND.n4304 GND.n4302 0.141472
R5657 GND.n4284 GND.n4281 0.141472
R5658 GND.n4265 GND.n4263 0.141472
R5659 GND.n4263 GND.n4240 0.141472
R5660 GND.n4240 GND.n4238 0.141472
R5661 GND.n4238 GND.n4225 0.141472
R5662 GND.n4225 GND.n4223 0.141472
R5663 GND.n4223 GND.n4210 0.141472
R5664 GND.n4210 GND.n4208 0.141472
R5665 GND.n4208 GND.n4195 0.141472
R5666 GND.n4195 GND.n4193 0.141472
R5667 GND.n4177 GND.n4174 0.141472
R5668 GND.n4174 GND.n4161 0.141472
R5669 GND.n4161 GND.n4159 0.141472
R5670 GND.n4159 GND.n4146 0.141472
R5671 GND.n4146 GND.n4144 0.141472
R5672 GND.n4144 GND.n4131 0.141472
R5673 GND.n4131 GND.n4129 0.141472
R5674 GND.n4129 GND.n4116 0.141472
R5675 GND.n4116 GND.n4114 0.141472
R5676 GND.n2109 GND.n2108 0.140882
R5677 GND.n6455 GND 0.140869
R5678 GND.n540 GND 0.140869
R5679 GND.n4302 GND.n4287 0.136611
R5680 GND.n7801 GND 0.134348
R5681 GND.n6378 GND 0.134348
R5682 GND.n4077 GND.n4076 0.134262
R5683 GND.n3224 GND.n3223 0.131784
R5684 GND.n2885 GND.n2884 0.131784
R5685 GND.n2886 GND.n2885 0.131784
R5686 GND.n3993 GND.n3992 0.131784
R5687 GND.n5293 GND.n5292 0.131784
R5688 GND.n5294 GND.n5293 0.131784
R5689 GND.n3881 GND.n3880 0.131784
R5690 GND.n5428 GND.n5427 0.131784
R5691 GND.n5429 GND.n5428 0.131784
R5692 GND.n3554 GND.n3553 0.131784
R5693 GND.n1588 GND.n1587 0.131784
R5694 GND.n1589 GND.n1588 0.131784
R5695 GND.n2013 GND.n2012 0.131784
R5696 GND.n7732 GND.n7731 0.131784
R5697 GND.n7733 GND.n7732 0.131784
R5698 GND.n2104 GND.n2103 0.131784
R5699 GND.n2329 GND.n2328 0.131784
R5700 GND.n2330 GND.n2329 0.131784
R5701 GND.n2481 GND.n2480 0.131784
R5702 GND.n2775 GND.n2774 0.131784
R5703 GND.n4940 GND.n4939 0.131784
R5704 GND.n4941 GND.n4940 0.131784
R5705 GND.n4729 GND.n4728 0.131784
R5706 GND.n3227 GND.n3224 0.13084
R5707 GND.n3996 GND.n3993 0.13084
R5708 GND.n3884 GND.n3881 0.13084
R5709 GND.n3557 GND.n3554 0.13084
R5710 GND.n2016 GND.n2013 0.13084
R5711 GND.n2107 GND.n2104 0.13084
R5712 GND.n2484 GND.n2481 0.13084
R5713 GND.n2778 GND.n2775 0.13084
R5714 GND.n4732 GND.n4729 0.13084
R5715 GND.n6453 GND.n6452 0.12814
R5716 GND.n538 GND.n537 0.12814
R5717 GND.n4091 GND.n4089 0.127732
R5718 GND.n3226 GND.n3225 0.126877
R5719 GND.n2880 GND.n2879 0.126877
R5720 GND.n3995 GND.n3994 0.126877
R5721 GND.n5288 GND.n5287 0.126877
R5722 GND.n3883 GND.n3882 0.126877
R5723 GND.n5423 GND.n5422 0.126877
R5724 GND.n3556 GND.n3555 0.126877
R5725 GND.n1583 GND.n1582 0.126877
R5726 GND.n2015 GND.n2014 0.126877
R5727 GND.n7727 GND.n7726 0.126877
R5728 GND.n2106 GND.n2105 0.126877
R5729 GND.n2324 GND.n2323 0.126877
R5730 GND.n2483 GND.n2482 0.126877
R5731 GND.n2777 GND.n2776 0.126877
R5732 GND.n4935 GND.n4934 0.126877
R5733 GND.n4731 GND.n4730 0.126877
R5734 GND.n4732 GND.n4731 0.125988
R5735 GND.n3227 GND.n3226 0.125988
R5736 GND.n3996 GND.n3995 0.125988
R5737 GND.n3884 GND.n3883 0.125988
R5738 GND.n3557 GND.n3556 0.125988
R5739 GND.n2016 GND.n2015 0.125988
R5740 GND.n2107 GND.n2106 0.125988
R5741 GND.n2484 GND.n2483 0.125988
R5742 GND.n2778 GND.n2777 0.125988
R5743 GND.n2887 GND.n2880 0.125687
R5744 GND.n5295 GND.n5288 0.125687
R5745 GND.n5430 GND.n5423 0.125687
R5746 GND.n1590 GND.n1583 0.125687
R5747 GND.n7734 GND.n7727 0.125687
R5748 GND.n2331 GND.n2324 0.125687
R5749 GND.n4942 GND.n4935 0.125687
R5750 GND.n4193 GND.n4180 0.1255
R5751 GND.n7573 GND.n7572 0.122064
R5752 GND.n7511 GND.n7510 0.122064
R5753 GND.n7449 GND.n7448 0.122064
R5754 GND.n5114 GND.n5113 0.122064
R5755 GND.n3714 GND.n3713 0.122064
R5756 GND.n5457 GND.n5456 0.122064
R5757 GND.n5514 GND.n5513 0.122064
R5758 GND.n5641 GND.n5640 0.122064
R5759 GND.n6502 GND.n6501 0.122064
R5760 GND.n7761 GND.n7760 0.122064
R5761 GND.n6825 GND.n6824 0.122064
R5762 GND.n6979 GND.n6978 0.122064
R5763 GND.n7080 GND.n7079 0.122064
R5764 GND.n2627 GND.n2626 0.122064
R5765 GND.n3053 GND.n3052 0.122064
R5766 GND.n3324 GND.n3323 0.122064
R5767 GND.n4084 GND.n4082 0.118804
R5768 GND.n4976 GND.n4594 0.118
R5769 GND.n4550 GND.n4491 0.117638
R5770 GND.t12 GND.t209 0.117638
R5771 GND.t537 GND.t401 0.117638
R5772 GND.t257 GND.t299 0.117638
R5773 GND.t289 GND.t80 0.117638
R5774 GND.t250 GND.t481 0.117638
R5775 GND.t244 GND.t21 0.117638
R5776 GND.t78 GND.t79 0.117638
R5777 GND.t417 GND.t589 0.117638
R5778 GND.n4114 GND.n4108 0.117167
R5779 GND.n6449 GND.n6448 0.1155
R5780 GND.n6448 GND.n6446 0.1155
R5781 GND.n6443 GND.n6442 0.1155
R5782 GND.n6442 GND.n6440 0.1155
R5783 GND.n6437 GND.n6436 0.1155
R5784 GND.n6436 GND.n6434 0.1155
R5785 GND.n6431 GND.n6430 0.1155
R5786 GND.n6430 GND.n6428 0.1155
R5787 GND.n534 GND.n533 0.1155
R5788 GND.n533 GND.n531 0.1155
R5789 GND.n528 GND.n527 0.1155
R5790 GND.n527 GND.n525 0.1155
R5791 GND.n522 GND.n521 0.1155
R5792 GND.n521 GND.n519 0.1155
R5793 GND.n516 GND.n515 0.1155
R5794 GND.n515 GND.n513 0.1155
R5795 GND.n7564 GND.n303 0.112135
R5796 GND.n7627 GND.n7626 0.112135
R5797 GND.n2528 GND.n2526 0.112135
R5798 GND.n2951 GND.n2945 0.112135
R5799 GND.n6923 GND.n6921 0.112135
R5800 GND.n6769 GND.n6767 0.112135
R5801 GND.n6660 GND.n6652 0.112135
R5802 GND.n5522 GND.n1102 0.112135
R5803 GND.n1270 GND.n1264 0.112135
R5804 GND.n7502 GND.n407 0.112135
R5805 GND.n5010 GND.n5004 0.112135
R5806 GND.n3616 GND.n3610 0.112135
R5807 GND.n5465 GND.n1223 0.112135
R5808 GND.n5604 GND.n639 0.112135
R5809 GND.n7077 GND.n7075 0.112135
R5810 GND.n3271 GND.n3265 0.112135
R5811 GND.n49 GND.n25 0.110055
R5812 GND.n6376 GND.n6352 0.110055
R5813 GND.n3374 GND.n3373 0.10956
R5814 GND.n3373 GND.n3372 0.10956
R5815 GND.n3356 GND.n3355 0.10956
R5816 GND.n3355 GND.n3354 0.10956
R5817 GND.n3379 GND.n3378 0.10956
R5818 GND.t440 GND.n3379 0.10956
R5819 GND.n3385 GND.n3384 0.10956
R5820 GND.t440 GND.n3385 0.10956
R5821 GND.n3110 GND.n3109 0.10956
R5822 GND.n3109 GND.n3108 0.10956
R5823 GND.n3085 GND.n3084 0.10956
R5824 GND.n3084 GND.n3083 0.10956
R5825 GND.n3129 GND.n3128 0.10956
R5826 GND.t1361 GND.n3129 0.10956
R5827 GND.t1361 GND.n3127 0.10956
R5828 GND.n3127 GND.n3126 0.10956
R5829 GND.n3115 GND.n3114 0.10956
R5830 GND.t1161 GND.n3115 0.10956
R5831 GND.n3121 GND.n3120 0.10956
R5832 GND.t1161 GND.n3121 0.10956
R5833 GND.n4033 GND.n4032 0.10956
R5834 GND.n4032 GND.n4031 0.10956
R5835 GND.n4008 GND.n4007 0.10956
R5836 GND.n4007 GND.n4006 0.10956
R5837 GND.n4052 GND.n4051 0.10956
R5838 GND.t1390 GND.n4052 0.10956
R5839 GND.t1390 GND.n4050 0.10956
R5840 GND.n4050 GND.n4049 0.10956
R5841 GND.n4038 GND.n4037 0.10956
R5842 GND.t678 GND.n4038 0.10956
R5843 GND.n4044 GND.n4043 0.10956
R5844 GND.t678 GND.n4044 0.10956
R5845 GND.n5188 GND.n5187 0.10956
R5846 GND.n5187 GND.n5186 0.10956
R5847 GND.n5147 GND.n5146 0.10956
R5848 GND.n5146 GND.n5145 0.10956
R5849 GND.n5163 GND.n5162 0.10956
R5850 GND.t1395 GND.n5163 0.10956
R5851 GND.n5169 GND.n5168 0.10956
R5852 GND.t1395 GND.n5169 0.10956
R5853 GND.n5177 GND.n5176 0.10956
R5854 GND.t389 GND.n5177 0.10956
R5855 GND.t389 GND.n5175 0.10956
R5856 GND.n5175 GND.n5174 0.10956
R5857 GND.n3787 GND.n3786 0.10956
R5858 GND.n3786 GND.n3785 0.10956
R5859 GND.n3746 GND.n3745 0.10956
R5860 GND.n3745 GND.n3744 0.10956
R5861 GND.n3776 GND.n3775 0.10956
R5862 GND.t1519 GND.n3776 0.10956
R5863 GND.t1519 GND.n3774 0.10956
R5864 GND.n3774 GND.n3773 0.10956
R5865 GND.n3762 GND.n3761 0.10956
R5866 GND.t522 GND.n3762 0.10956
R5867 GND.n3768 GND.n3767 0.10956
R5868 GND.t522 GND.n3768 0.10956
R5869 GND.n1322 GND.n1321 0.10956
R5870 GND.n1321 GND.n1320 0.10956
R5871 GND.n1281 GND.n1280 0.10956
R5872 GND.n1280 GND.n1279 0.10956
R5873 GND.n1297 GND.n1296 0.10956
R5874 GND.t304 GND.n1297 0.10956
R5875 GND.n1303 GND.n1302 0.10956
R5876 GND.t304 GND.n1303 0.10956
R5877 GND.n1311 GND.n1310 0.10956
R5878 GND.t292 GND.n1311 0.10956
R5879 GND.t292 GND.n1309 0.10956
R5880 GND.n1309 GND.n1308 0.10956
R5881 GND.n3465 GND.n3464 0.10956
R5882 GND.n3464 GND.n3463 0.10956
R5883 GND.n3424 GND.n3423 0.10956
R5884 GND.n3423 GND.n3422 0.10956
R5885 GND.n3454 GND.n3453 0.10956
R5886 GND.t855 GND.n3454 0.10956
R5887 GND.t855 GND.n3452 0.10956
R5888 GND.n3452 GND.n3451 0.10956
R5889 GND.n3440 GND.n3439 0.10956
R5890 GND.t574 GND.n3440 0.10956
R5891 GND.n3446 GND.n3445 0.10956
R5892 GND.t574 GND.n3446 0.10956
R5893 GND.n1490 GND.n1489 0.10956
R5894 GND.n1489 GND.n1488 0.10956
R5895 GND.n1449 GND.n1448 0.10956
R5896 GND.n1448 GND.n1447 0.10956
R5897 GND.n1465 GND.n1464 0.10956
R5898 GND.t1419 GND.n1465 0.10956
R5899 GND.n1471 GND.n1470 0.10956
R5900 GND.t1419 GND.n1471 0.10956
R5901 GND.n1479 GND.n1478 0.10956
R5902 GND.t641 GND.n1479 0.10956
R5903 GND.t641 GND.n1477 0.10956
R5904 GND.n1477 GND.n1476 0.10956
R5905 GND.n1916 GND.n1915 0.10956
R5906 GND.n1915 GND.n1914 0.10956
R5907 GND.n1875 GND.n1874 0.10956
R5908 GND.n1874 GND.n1873 0.10956
R5909 GND.n1905 GND.n1904 0.10956
R5910 GND.t254 GND.n1905 0.10956
R5911 GND.t254 GND.n1903 0.10956
R5912 GND.n1903 GND.n1902 0.10956
R5913 GND.n1891 GND.n1890 0.10956
R5914 GND.t427 GND.n1891 0.10956
R5915 GND.n1897 GND.n1896 0.10956
R5916 GND.t427 GND.n1897 0.10956
R5917 GND.n139 GND.n138 0.10956
R5918 GND.n138 GND.n137 0.10956
R5919 GND.n90 GND.n89 0.10956
R5920 GND.n89 GND.n88 0.10956
R5921 GND.n106 GND.n105 0.10956
R5922 GND.t326 GND.n106 0.10956
R5923 GND.n112 GND.n111 0.10956
R5924 GND.t326 GND.n112 0.10956
R5925 GND.n128 GND.n127 0.10956
R5926 GND.t274 GND.n128 0.10956
R5927 GND.t274 GND.n126 0.10956
R5928 GND.n126 GND.n125 0.10956
R5929 GND.n2167 GND.n2166 0.10956
R5930 GND.n2166 GND.n2165 0.10956
R5931 GND.n2126 GND.n2125 0.10956
R5932 GND.n2125 GND.n2124 0.10956
R5933 GND.n2156 GND.n2155 0.10956
R5934 GND.t277 GND.n2156 0.10956
R5935 GND.t277 GND.n2154 0.10956
R5936 GND.n2154 GND.n2153 0.10956
R5937 GND.n2142 GND.n2141 0.10956
R5938 GND.t1415 GND.n2142 0.10956
R5939 GND.n2148 GND.n2147 0.10956
R5940 GND.t1415 GND.n2148 0.10956
R5941 GND.n2229 GND.n2228 0.10956
R5942 GND.n2228 GND.n2227 0.10956
R5943 GND.n2188 GND.n2187 0.10956
R5944 GND.n2187 GND.n2186 0.10956
R5945 GND.n2204 GND.n2203 0.10956
R5946 GND.t442 GND.n2204 0.10956
R5947 GND.n2210 GND.n2209 0.10956
R5948 GND.t442 GND.n2210 0.10956
R5949 GND.n2218 GND.n2217 0.10956
R5950 GND.t1124 GND.n2218 0.10956
R5951 GND.t1124 GND.n2216 0.10956
R5952 GND.n2216 GND.n2215 0.10956
R5953 GND.n2392 GND.n2391 0.10956
R5954 GND.n2391 GND.n2390 0.10956
R5955 GND.n2351 GND.n2350 0.10956
R5956 GND.n2350 GND.n2349 0.10956
R5957 GND.n2381 GND.n2380 0.10956
R5958 GND.t1379 GND.n2381 0.10956
R5959 GND.n2367 GND.n2366 0.10956
R5960 GND.t1041 GND.n2367 0.10956
R5961 GND.n2373 GND.n2372 0.10956
R5962 GND.t1041 GND.n2373 0.10956
R5963 GND.n2686 GND.n2685 0.10956
R5964 GND.n2685 GND.n2684 0.10956
R5965 GND.n2663 GND.n2662 0.10956
R5966 GND.n2662 GND.n2661 0.10956
R5967 GND.n2705 GND.n2704 0.10956
R5968 GND.t861 GND.n2705 0.10956
R5969 GND.t861 GND.n2703 0.10956
R5970 GND.n2703 GND.n2702 0.10956
R5971 GND.n2691 GND.n2690 0.10956
R5972 GND.t667 GND.n2691 0.10956
R5973 GND.n2697 GND.n2696 0.10956
R5974 GND.t667 GND.n2697 0.10956
R5975 GND.t1379 GND.n2379 0.10956
R5976 GND.n2379 GND.n2378 0.10956
R5977 GND.n4845 GND.n4844 0.10956
R5978 GND.n4844 GND.n4843 0.10956
R5979 GND.n4804 GND.n4803 0.10956
R5980 GND.n4803 GND.n4802 0.10956
R5981 GND.n4834 GND.n4833 0.10956
R5982 GND.t1069 GND.n4834 0.10956
R5983 GND.t1069 GND.n4832 0.10956
R5984 GND.n4832 GND.n4831 0.10956
R5985 GND.n4820 GND.n4819 0.10956
R5986 GND.t253 GND.n4820 0.10956
R5987 GND.n4826 GND.n4825 0.10956
R5988 GND.t253 GND.n4826 0.10956
R5989 GND.n4242 GND.n4241 0.10956
R5990 GND.n4243 GND.n4242 0.10956
R5991 GND.n4250 GND.n4249 0.10956
R5992 GND.n4251 GND.n4250 0.10956
R5993 GND.n4613 GND.n4612 0.10956
R5994 GND.t307 GND.n4613 0.10956
R5995 GND.n4619 GND.n4618 0.10956
R5996 GND.t307 GND.n4619 0.10956
R5997 GND.n4638 GND.n4637 0.10956
R5998 GND.n4637 GND.n4636 0.10956
R5999 GND.n4597 GND.n4596 0.10956
R6000 GND.n4596 GND.n4595 0.10956
R6001 GND.n4627 GND.n4626 0.10956
R6002 GND.t258 GND.n4627 0.10956
R6003 GND.t258 GND.n4625 0.10956
R6004 GND.n4625 GND.n4624 0.10956
R6005 GND.n4714 GND.t503 0.10956
R6006 GND.n4712 GND.n4711 0.10956
R6007 GND.t503 GND.n4712 0.10956
R6008 GND.n4715 GND.n4714 0.10956
R6009 GND.n3306 GND.n3305 0.10956
R6010 GND.n3305 GND.n3304 0.10956
R6011 GND.n3000 GND.n2999 0.10956
R6012 GND.t1152 GND.n3000 0.10956
R6013 GND.n3003 GND.n3002 0.10956
R6014 GND.n3002 GND.n3001 0.10956
R6015 GND.n2574 GND.n2573 0.10956
R6016 GND.t1167 GND.n2574 0.10956
R6017 GND.n2577 GND.n2576 0.10956
R6018 GND.n2576 GND.n2575 0.10956
R6019 GND.n7174 GND.n7173 0.10956
R6020 GND.t363 GND.n7174 0.10956
R6021 GND.n7177 GND.n7176 0.10956
R6022 GND.n7176 GND.n7175 0.10956
R6023 GND.n7011 GND.n7010 0.10956
R6024 GND.t853 GND.n7011 0.10956
R6025 GND.n7014 GND.n7013 0.10956
R6026 GND.n7013 GND.n7012 0.10956
R6027 GND.n6857 GND.n6856 0.10956
R6028 GND.t1411 GND.n6857 0.10956
R6029 GND.n6860 GND.n6859 0.10956
R6030 GND.n6859 GND.n6858 0.10956
R6031 GND.n6703 GND.n6702 0.10956
R6032 GND.t359 GND.n6703 0.10956
R6033 GND.n6706 GND.n6705 0.10956
R6034 GND.n6705 GND.n6704 0.10956
R6035 GND.n6632 GND.n6631 0.10956
R6036 GND.t1386 GND.n6632 0.10956
R6037 GND.n6635 GND.n6634 0.10956
R6038 GND.n6634 GND.n6633 0.10956
R6039 GND.n5584 GND.n5583 0.10956
R6040 GND.t261 GND.n5584 0.10956
R6041 GND.n5587 GND.n5586 0.10956
R6042 GND.n5586 GND.n5585 0.10956
R6043 GND.n1082 GND.n1081 0.10956
R6044 GND.t265 GND.n1082 0.10956
R6045 GND.n1085 GND.n1084 0.10956
R6046 GND.n1084 GND.n1083 0.10956
R6047 GND.n1203 GND.n1202 0.10956
R6048 GND.t313 GND.n1203 0.10956
R6049 GND.n1206 GND.n1205 0.10956
R6050 GND.n1205 GND.n1204 0.10956
R6051 GND.n3664 GND.n3663 0.10956
R6052 GND.t881 GND.n3664 0.10956
R6053 GND.n3667 GND.n3666 0.10956
R6054 GND.n3666 GND.n3665 0.10956
R6055 GND.n5061 GND.n5060 0.10956
R6056 GND.t248 GND.n5061 0.10956
R6057 GND.n5064 GND.n5063 0.10956
R6058 GND.n5063 GND.n5062 0.10956
R6059 GND.n456 GND.n455 0.10956
R6060 GND.t543 GND.n456 0.10956
R6061 GND.n459 GND.n458 0.10956
R6062 GND.n458 GND.n457 0.10956
R6063 GND.n387 GND.n386 0.10956
R6064 GND.t1424 GND.n387 0.10956
R6065 GND.n390 GND.n389 0.10956
R6066 GND.n389 GND.n388 0.10956
R6067 GND.n283 GND.n282 0.10956
R6068 GND.t557 GND.n283 0.10956
R6069 GND.n286 GND.n285 0.10956
R6070 GND.n285 GND.n284 0.10956
R6071 GND.n186 GND.n185 0.10956
R6072 GND.t684 GND.n186 0.10956
R6073 GND.n4974 GND 0.104579
R6074 GND.n3367 GND.n3366 0.104537
R6075 GND.n3366 GND.n3365 0.104537
R6076 GND.n3099 GND.n3098 0.104537
R6077 GND.n3098 GND.n3097 0.104537
R6078 GND.n4022 GND.n4021 0.104537
R6079 GND.n4021 GND.n4020 0.104537
R6080 GND.n5161 GND.n5160 0.104537
R6081 GND.n5160 GND.n5159 0.104537
R6082 GND.n3760 GND.n3759 0.104537
R6083 GND.n3759 GND.n3758 0.104537
R6084 GND.n1295 GND.n1294 0.104537
R6085 GND.n1294 GND.n1293 0.104537
R6086 GND.n3438 GND.n3437 0.104537
R6087 GND.n3437 GND.n3436 0.104537
R6088 GND.n1463 GND.n1462 0.104537
R6089 GND.n1462 GND.n1461 0.104537
R6090 GND.n1889 GND.n1888 0.104537
R6091 GND.n1888 GND.n1887 0.104537
R6092 GND.n104 GND.n103 0.104537
R6093 GND.n103 GND.n102 0.104537
R6094 GND.n2140 GND.n2139 0.104537
R6095 GND.n2139 GND.n2138 0.104537
R6096 GND.n2202 GND.n2201 0.104537
R6097 GND.n2201 GND.n2200 0.104537
R6098 GND.n2365 GND.n2364 0.104537
R6099 GND.n2364 GND.n2363 0.104537
R6100 GND.n2677 GND.n2676 0.104537
R6101 GND.n2676 GND.n2675 0.104537
R6102 GND.n4818 GND.n4817 0.104537
R6103 GND.n4817 GND.n4816 0.104537
R6104 GND.n4611 GND.n4610 0.104537
R6105 GND.n4610 GND.n4609 0.104537
R6106 GND.n6351 GND.n6330 0.102336
R6107 GND.n7798 GND.n7797 0.102336
R6108 GND.n7565 GND.n7564 0.102333
R6109 GND.n7626 GND.n201 0.102333
R6110 GND.n2528 GND.n2527 0.102333
R6111 GND.n2951 GND.n2950 0.102333
R6112 GND.n6923 GND.n6922 0.102333
R6113 GND.n6769 GND.n6768 0.102333
R6114 GND.n6660 GND.n6659 0.102333
R6115 GND.n5522 GND.n5521 0.102333
R6116 GND.n1270 GND.n1269 0.102333
R6117 GND.n7503 GND.n7502 0.102333
R6118 GND.n5010 GND.n5009 0.102333
R6119 GND.n3616 GND.n3615 0.102333
R6120 GND.n5465 GND.n5464 0.102333
R6121 GND.n5642 GND.n639 0.102333
R6122 GND.n7077 GND.n7076 0.102333
R6123 GND.n3271 GND.n3270 0.102333
R6124 GND.n7780 GND 0.101889
R6125 GND.n6313 GND 0.101889
R6126 GND.n4594 GND 0.0991625
R6127 GND.n35 GND.n34 0.0963333
R6128 GND.n36 GND.n27 0.0963333
R6129 GND.n42 GND.n27 0.0963333
R6130 GND.n43 GND.n42 0.0963333
R6131 GND.n44 GND.n43 0.0963333
R6132 GND.n6362 GND.n6361 0.0963333
R6133 GND.n6363 GND.n6354 0.0963333
R6134 GND.n6369 GND.n6354 0.0963333
R6135 GND.n6370 GND.n6369 0.0963333
R6136 GND.n6371 GND.n6370 0.0963333
R6137 GND.n4248 GND.n4247 0.0944005
R6138 GND.n3321 GND.n3320 0.0944005
R6139 GND.n3322 GND.n3321 0.0944005
R6140 GND.n3267 GND.n3266 0.0944005
R6141 GND.n3049 GND.n3048 0.0944005
R6142 GND.n3050 GND.n3049 0.0944005
R6143 GND.n2947 GND.n2946 0.0944005
R6144 GND.n2623 GND.n2622 0.0944005
R6145 GND.n2624 GND.n2623 0.0944005
R6146 GND.n7228 GND.n598 0.0944005
R6147 GND.n7227 GND.n7226 0.0944005
R6148 GND.n7228 GND.n7227 0.0944005
R6149 GND.n6982 GND.n6981 0.0944005
R6150 GND.n6984 GND.n6983 0.0944005
R6151 GND.n6983 GND.n6982 0.0944005
R6152 GND.n6828 GND.n6827 0.0944005
R6153 GND.n6830 GND.n6829 0.0944005
R6154 GND.n6829 GND.n6828 0.0944005
R6155 GND.n6664 GND.n6663 0.0944005
R6156 GND.n6666 GND.n6665 0.0944005
R6157 GND.n6665 GND.n6664 0.0944005
R6158 GND.n6656 GND.n6655 0.0944005
R6159 GND.n6655 GND.n6654 0.0944005
R6160 GND.n6654 GND.n6653 0.0944005
R6161 GND.n5646 GND.n5645 0.0944005
R6162 GND.n5648 GND.n5646 0.0944005
R6163 GND.n5648 GND.n5647 0.0944005
R6164 GND.n5518 GND.n5517 0.0944005
R6165 GND.n5517 GND.n5516 0.0944005
R6166 GND.n5467 GND.n5466 0.0944005
R6167 GND.n5461 GND.n5460 0.0944005
R6168 GND.n5460 GND.n5459 0.0944005
R6169 GND.n1138 GND.n1137 0.0944005
R6170 GND.n1266 GND.n1265 0.0944005
R6171 GND.n3710 GND.n3709 0.0944005
R6172 GND.n3711 GND.n3710 0.0944005
R6173 GND.n3612 GND.n3611 0.0944005
R6174 GND.n5110 GND.n5109 0.0944005
R6175 GND.n5111 GND.n5110 0.0944005
R6176 GND.n5006 GND.n5005 0.0944005
R6177 GND.n504 GND.n503 0.0944005
R6178 GND.n505 GND.n504 0.0944005
R6179 GND.n7507 GND.n7506 0.0944005
R6180 GND.n7508 GND.n7507 0.0944005
R6181 GND.n315 GND.n314 0.0944005
R6182 GND.n7569 GND.n7568 0.0944005
R6183 GND.n7570 GND.n7569 0.0944005
R6184 GND.n213 GND.n212 0.0944005
R6185 GND.n198 GND.n197 0.0944005
R6186 GND.n197 GND.n196 0.0944005
R6187 GND.n3252 GND.n3250 0.0921667
R6188 GND.n7555 GND.n7553 0.0921667
R6189 GND.n7617 GND.n7615 0.0921667
R6190 GND.n2513 GND.n2511 0.0921667
R6191 GND.n2930 GND.n2928 0.0921667
R6192 GND.n6956 GND.n6954 0.0921667
R6193 GND.n6792 GND.n6790 0.0921667
R6194 GND.n82 GND.n80 0.0921667
R6195 GND.n1025 GND.n1023 0.0921667
R6196 GND.n1252 GND.n1250 0.0921667
R6197 GND.n7494 GND.n7492 0.0921667
R6198 GND.n4993 GND.n4991 0.0921667
R6199 GND.n3595 GND.n3593 0.0921667
R6200 GND.n1124 GND.n1122 0.0921667
R6201 GND.n6546 GND.n6544 0.0921667
R6202 GND.n7124 GND.n7122 0.0921667
R6203 GND.n4452 GND.n4450 0.0920099
R6204 GND.n719 GND.n717 0.0894537
R6205 GND.n5866 GND.n5864 0.0894537
R6206 GND.n7237 GND.n7235 0.0894537
R6207 GND.n3339 GND.n3337 0.0891364
R6208 GND.n7526 GND.n7524 0.0891364
R6209 GND.n7588 GND.n7586 0.0891364
R6210 GND.n2642 GND.n2640 0.0891364
R6211 GND.n3068 GND.n3066 0.0891364
R6212 GND.n6934 GND.n6932 0.0891364
R6213 GND.n6811 GND.n6809 0.0891364
R6214 GND.n59 GND.n57 0.0891364
R6215 GND.n1004 GND.n1002 0.0891364
R6216 GND.n1233 GND.n1231 0.0891364
R6217 GND.n7464 GND.n7462 0.0891364
R6218 GND.n5129 GND.n5127 0.0891364
R6219 GND.n3729 GND.n3727 0.0891364
R6220 GND.n5500 GND.n5498 0.0891364
R6221 GND.n6521 GND.n6519 0.0891364
R6222 GND.n7095 GND.n7093 0.0891364
R6223 GND.n4903 GND.n4902 0.08745
R6224 GND.n4702 GND.n4701 0.08745
R6225 GND.n3158 GND.n3157 0.08745
R6226 GND.n2287 GND.n2286 0.08745
R6227 GND.n7691 GND.n7690 0.08745
R6228 GND.n1547 GND.n1546 0.08745
R6229 GND.n5384 GND.n5383 0.08745
R6230 GND.n3953 GND.n3952 0.08745
R6231 GND.n5245 GND.n5244 0.08745
R6232 GND.n3845 GND.n3844 0.08745
R6233 GND.n3522 GND.n3521 0.08745
R6234 GND.n1974 GND.n1973 0.08745
R6235 GND.n2076 GND.n2075 0.08745
R6236 GND.n2449 GND.n2448 0.08745
R6237 GND.n2758 GND.n2757 0.08745
R6238 GND.n2862 GND.n2861 0.08745
R6239 GND.n4903 GND.n4858 0.0868625
R6240 GND.n4702 GND.n4678 0.0868625
R6241 GND.n3206 GND.n3158 0.0868625
R6242 GND.n2287 GND.n2242 0.0868625
R6243 GND.n7691 GND.n7669 0.0868625
R6244 GND.n1547 GND.n1502 0.0868625
R6245 GND.n5384 GND.n5339 0.0868625
R6246 GND.n3953 GND.n3908 0.0868625
R6247 GND.n5245 GND.n5200 0.0868625
R6248 GND.n3845 GND.n3800 0.0868625
R6249 GND.n3522 GND.n3477 0.0868625
R6250 GND.n1974 GND.n1929 0.0868625
R6251 GND.n2076 GND.n2052 0.0868625
R6252 GND.n2449 GND.n2404 0.0868625
R6253 GND.n2758 GND.n2713 0.0868625
R6254 GND.n2862 GND.n2817 0.0868625
R6255 GND.n4075 GND.n4073 0.0853214
R6256 GND.n7539 GND.n305 0.0845572
R6257 GND.n7601 GND.n203 0.0845572
R6258 GND.n2656 GND.n2655 0.0845572
R6259 GND.n3082 GND.n3081 0.0845572
R6260 GND.n6964 GND.n6963 0.0845572
R6261 GND.n6801 GND.n6800 0.0845572
R6262 GND.n7746 GND.n7745 0.0845572
R6263 GND.n5626 GND.n5625 0.0845572
R6264 GND.n5442 GND.n5441 0.0845572
R6265 GND.n7477 GND.n499 0.0845572
R6266 GND.n5143 GND.n5142 0.0845572
R6267 GND.n3743 GND.n3742 0.0845572
R6268 GND.n6530 GND.n640 0.0845572
R6269 GND.n3353 GND.n3352 0.0845572
R6270 GND.n4379 GND.n4366 0.0838333
R6271 GND.n6498 GND 0.0824444
R6272 GND.n6295 GND 0.0824444
R6273 GND.n3239 GND 0.0775833
R6274 GND.n7542 GND 0.0775833
R6275 GND.n7604 GND 0.0775833
R6276 GND.n2503 GND 0.0775833
R6277 GND.n2920 GND 0.0775833
R6278 GND.n6942 GND 0.0775833
R6279 GND.n6779 GND 0.0775833
R6280 GND.n68 GND 0.0775833
R6281 GND.n1012 GND 0.0775833
R6282 GND.n1241 GND 0.0775833
R6283 GND.n7480 GND 0.0775833
R6284 GND.n4979 GND 0.0775833
R6285 GND.n3585 GND 0.0775833
R6286 GND.n1111 GND 0.0775833
R6287 GND.n6533 GND 0.0775833
R6288 GND.n7111 GND 0.0775833
R6289 GND.n6406 GND.n6381 0.0740087
R6290 GND.n6496 GND.n50 0.0740087
R6291 GND.n6407 GND.n6406 0.0732412
R6292 GND.n6497 GND.n6496 0.0732412
R6293 GND.n6408 GND.n6407 0.0727407
R6294 GND.n6497 GND.n6471 0.0727407
R6295 GND.n4267 GND.n4265 0.0727222
R6296 GND.n6471 GND.n666 0.0714246
R6297 GND.n7435 GND.n7434 0.0711855
R6298 GND.n6457 GND.n6456 0.0696598
R6299 GND.n7439 GND.n7438 0.0696598
R6300 GND.n6381 GND.n6380 0.0692593
R6301 GND.n7799 GND.n50 0.0692593
R6302 GND.n4281 GND.n4267 0.06925
R6303 GND.n3327 GND 0.0675455
R6304 GND.n7514 GND 0.0675455
R6305 GND.n7576 GND 0.0675455
R6306 GND.n2630 GND 0.0675455
R6307 GND.n3056 GND 0.0675455
R6308 GND GND.n6977 0.0675455
R6309 GND GND.n6823 0.0675455
R6310 GND GND.n7759 0.0675455
R6311 GND GND.n5639 0.0675455
R6312 GND GND.n5455 0.0675455
R6313 GND.n7452 GND 0.0675455
R6314 GND.n5117 GND 0.0675455
R6315 GND.n3717 GND 0.0675455
R6316 GND GND.n5512 0.0675455
R6317 GND.n6505 GND 0.0675455
R6318 GND.n7083 GND 0.0675455
R6319 GND.n4975 GND.n4974 0.0672895
R6320 GND.n5312 GND.n5311 0.0672895
R6321 GND.n5311 GND.n1334 0.0672895
R6322 GND.n5336 GND.n1334 0.0672895
R6323 GND.n5336 GND.n5335 0.0672895
R6324 GND.n3408 GND.n3407 0.0672895
R6325 GND.n3407 GND.n3406 0.0672895
R6326 GND.n3406 GND.n3405 0.0672895
R6327 GND.n3405 GND.n3404 0.0672895
R6328 GND.n3404 GND.n3403 0.0672895
R6329 GND.n16 GND.n11 0.0659695
R6330 GND.n6341 GND.n6336 0.0659695
R6331 GND.n1379 GND.n1378 0.0653227
R6332 GND.n6221 GND.n6220 0.0643889
R6333 GND.n6220 GND.n6218 0.0643889
R6334 GND.n6218 GND.n6215 0.0643889
R6335 GND.n6215 GND.n6213 0.0643889
R6336 GND.n16 GND.n8 0.0643889
R6337 GND.n20 GND.n8 0.0643889
R6338 GND.n21 GND.n20 0.0643889
R6339 GND.n7778 GND.n7771 0.0643889
R6340 GND.n7784 GND.n7769 0.0643889
R6341 GND.n7784 GND.n7766 0.0643889
R6342 GND.n7788 GND.n7766 0.0643889
R6343 GND.n7789 GND.n7788 0.0643889
R6344 GND.n651 GND.n646 0.0643889
R6345 GND.n662 GND.n644 0.0643889
R6346 GND.n663 GND.n662 0.0643889
R6347 GND.n6341 GND.n6333 0.0643889
R6348 GND.n6345 GND.n6333 0.0643889
R6349 GND.n6346 GND.n6345 0.0643889
R6350 GND.n6311 GND.n6304 0.0643889
R6351 GND.n6317 GND.n6302 0.0643889
R6352 GND.n6317 GND.n6299 0.0643889
R6353 GND.n6321 GND.n6299 0.0643889
R6354 GND.n6322 GND.n6321 0.0643889
R6355 GND.n6279 GND.n6274 0.0643889
R6356 GND.n6290 GND.n6272 0.0643889
R6357 GND.n6291 GND.n6290 0.0643889
R6358 GND.n3146 GND.t561 0.0636886
R6359 GND.n3147 GND.n3146 0.0636886
R6360 GND.n3169 GND.n3168 0.0636886
R6361 GND.n3170 GND.n3169 0.0636886
R6362 GND.n3172 GND.n3171 0.0636886
R6363 GND.n3171 GND.n3170 0.0636886
R6364 GND.n2904 GND.n2903 0.0636886
R6365 GND.n2905 GND.n2904 0.0636886
R6366 GND.n2907 GND.n2906 0.0636886
R6367 GND.n2906 GND.n2905 0.0636886
R6368 GND.t562 GND.n2857 0.0636886
R6369 GND.n2857 GND.n2856 0.0636886
R6370 GND.n2858 GND.t562 0.0636886
R6371 GND.n2859 GND.n2858 0.0636886
R6372 GND.n2298 GND.n2297 0.0636886
R6373 GND.n2299 GND.n2298 0.0636886
R6374 GND.n2301 GND.n2300 0.0636886
R6375 GND.n2300 GND.n2299 0.0636886
R6376 GND.n7702 GND.n7701 0.0636886
R6377 GND.n7703 GND.n7702 0.0636886
R6378 GND.n7705 GND.n7704 0.0636886
R6379 GND.n7704 GND.n7703 0.0636886
R6380 GND.n1558 GND.n1557 0.0636886
R6381 GND.n1559 GND.n1558 0.0636886
R6382 GND.n1561 GND.n1560 0.0636886
R6383 GND.n1560 GND.n1559 0.0636886
R6384 GND.n5395 GND.n5394 0.0636886
R6385 GND.n5396 GND.n5395 0.0636886
R6386 GND.n5398 GND.n5397 0.0636886
R6387 GND.n5397 GND.n5396 0.0636886
R6388 GND.n5256 GND.n5255 0.0636886
R6389 GND.n5257 GND.n5256 0.0636886
R6390 GND.n5259 GND.n5258 0.0636886
R6391 GND.n5258 GND.n5257 0.0636886
R6392 GND.t563 GND.n3941 0.0636886
R6393 GND.n3941 GND.n3940 0.0636886
R6394 GND.n3942 GND.t563 0.0636886
R6395 GND.n3943 GND.n3942 0.0636886
R6396 GND.n5235 GND.n5234 0.0636886
R6397 GND.n5234 GND.t273 0.0636886
R6398 GND.n5233 GND.n5232 0.0636886
R6399 GND.t273 GND.n5233 0.0636886
R6400 GND.n3856 GND.n3855 0.0636886
R6401 GND.n3857 GND.n3856 0.0636886
R6402 GND.n3859 GND.n3858 0.0636886
R6403 GND.n3858 GND.n3857 0.0636886
R6404 GND.n3833 GND.n3832 0.0636886
R6405 GND.t549 GND.n3833 0.0636886
R6406 GND.n3834 GND.t549 0.0636886
R6407 GND.n3835 GND.n3834 0.0636886
R6408 GND.n5374 GND.n5373 0.0636886
R6409 GND.n5373 GND.t568 0.0636886
R6410 GND.n5372 GND.n5371 0.0636886
R6411 GND.t568 GND.n5372 0.0636886
R6412 GND.n3533 GND.n3532 0.0636886
R6413 GND.n3534 GND.n3533 0.0636886
R6414 GND.n3536 GND.n3535 0.0636886
R6415 GND.n3535 GND.n3534 0.0636886
R6416 GND.n3510 GND.n3509 0.0636886
R6417 GND.t564 GND.n3510 0.0636886
R6418 GND.n3511 GND.t564 0.0636886
R6419 GND.n3512 GND.n3511 0.0636886
R6420 GND.n1537 GND.n1536 0.0636886
R6421 GND.n1536 GND.t447 0.0636886
R6422 GND.n1535 GND.n1534 0.0636886
R6423 GND.t447 GND.n1535 0.0636886
R6424 GND.n1985 GND.n1984 0.0636886
R6425 GND.n1986 GND.n1985 0.0636886
R6426 GND.n1988 GND.n1987 0.0636886
R6427 GND.n1987 GND.n1986 0.0636886
R6428 GND.n1962 GND.n1961 0.0636886
R6429 GND.t448 GND.n1962 0.0636886
R6430 GND.n1963 GND.t448 0.0636886
R6431 GND.n1964 GND.n1963 0.0636886
R6432 GND.n7681 GND.n7680 0.0636886
R6433 GND.n7680 GND.t1071 0.0636886
R6434 GND.t1071 GND.n7679 0.0636886
R6435 GND.n7679 GND.n7678 0.0636886
R6436 GND.n2080 GND.n2079 0.0636886
R6437 GND.n2085 GND.n2084 0.0636886
R6438 GND.n2071 GND.n2070 0.0636886
R6439 GND.t269 GND.n2071 0.0636886
R6440 GND.n2072 GND.t269 0.0636886
R6441 GND.n2073 GND.n2072 0.0636886
R6442 GND.n2277 GND.n2276 0.0636886
R6443 GND.n2276 GND.t270 0.0636886
R6444 GND.n2275 GND.n2274 0.0636886
R6445 GND.t270 GND.n2275 0.0636886
R6446 GND.n2460 GND.n2459 0.0636886
R6447 GND.n2461 GND.n2460 0.0636886
R6448 GND.n2463 GND.n2462 0.0636886
R6449 GND.n2462 GND.n2461 0.0636886
R6450 GND.n2439 GND.n2438 0.0636886
R6451 GND.n2438 GND.t536 0.0636886
R6452 GND.n2746 GND.n2745 0.0636886
R6453 GND.t573 GND.n2746 0.0636886
R6454 GND.n2748 GND.n2747 0.0636886
R6455 GND.n2747 GND.t573 0.0636886
R6456 GND.n2437 GND.n2436 0.0636886
R6457 GND.t536 GND.n2437 0.0636886
R6458 GND.n2801 GND.n2800 0.0636886
R6459 GND.n2802 GND.n2801 0.0636886
R6460 GND.n2804 GND.n2803 0.0636886
R6461 GND.n2803 GND.n2802 0.0636886
R6462 GND.n4914 GND.n4913 0.0636886
R6463 GND.n4915 GND.n4914 0.0636886
R6464 GND.n4917 GND.n4916 0.0636886
R6465 GND.n4916 GND.n4915 0.0636886
R6466 GND.n4891 GND.n4890 0.0636886
R6467 GND.t1128 GND.n4891 0.0636886
R6468 GND.n4892 GND.t1128 0.0636886
R6469 GND.n4893 GND.n4892 0.0636886
R6470 GND.n3970 GND.n3969 0.0636886
R6471 GND.n3971 GND.n3970 0.0636886
R6472 GND.n3973 GND.n3972 0.0636886
R6473 GND.n3972 GND.n3971 0.0636886
R6474 GND.n1610 GND.n1609 0.0636886
R6475 GND.n1746 GND.n1610 0.0636886
R6476 GND.n1606 GND.n1605 0.0636886
R6477 GND.n1746 GND.n1606 0.0636886
R6478 GND.n1748 GND.n1747 0.0636886
R6479 GND.t296 GND.n1748 0.0636886
R6480 GND.n1620 GND.n1619 0.0636886
R6481 GND.n1746 GND.n1620 0.0636886
R6482 GND.n1615 GND.n1614 0.0636886
R6483 GND.n1746 GND.n1615 0.0636886
R6484 GND.n1750 GND.n1749 0.0636886
R6485 GND.t296 GND.n1750 0.0636886
R6486 GND.n1630 GND.n1629 0.0636886
R6487 GND.n1746 GND.n1630 0.0636886
R6488 GND.n1624 GND.n1623 0.0636886
R6489 GND.n1746 GND.n1624 0.0636886
R6490 GND.n1752 GND.n1751 0.0636886
R6491 GND.t296 GND.n1752 0.0636886
R6492 GND.n1640 GND.n1639 0.0636886
R6493 GND.n1746 GND.n1640 0.0636886
R6494 GND.n1634 GND.n1633 0.0636886
R6495 GND.n1746 GND.n1634 0.0636886
R6496 GND.n1754 GND.n1753 0.0636886
R6497 GND.t296 GND.n1754 0.0636886
R6498 GND.n1650 GND.n1649 0.0636886
R6499 GND.n1746 GND.n1650 0.0636886
R6500 GND.n1646 GND.n1645 0.0636886
R6501 GND.n1746 GND.n1646 0.0636886
R6502 GND.n1756 GND.n1755 0.0636886
R6503 GND.t296 GND.n1756 0.0636886
R6504 GND.n1665 GND.n1664 0.0636886
R6505 GND.n1746 GND.n1665 0.0636886
R6506 GND.n1656 GND.n1655 0.0636886
R6507 GND.n1746 GND.n1656 0.0636886
R6508 GND.n1758 GND.n1757 0.0636886
R6509 GND.t296 GND.n1758 0.0636886
R6510 GND.n1675 GND.n1674 0.0636886
R6511 GND.n1746 GND.n1675 0.0636886
R6512 GND.n1670 GND.n1669 0.0636886
R6513 GND.n1746 GND.n1670 0.0636886
R6514 GND.n1760 GND.n1759 0.0636886
R6515 GND.t296 GND.n1760 0.0636886
R6516 GND.n1685 GND.n1684 0.0636886
R6517 GND.n1746 GND.n1685 0.0636886
R6518 GND.n1681 GND.n1680 0.0636886
R6519 GND.n1746 GND.n1681 0.0636886
R6520 GND.n1762 GND.n1761 0.0636886
R6521 GND.t296 GND.n1762 0.0636886
R6522 GND.n1695 GND.n1694 0.0636886
R6523 GND.n1746 GND.n1695 0.0636886
R6524 GND.n1689 GND.n1688 0.0636886
R6525 GND.n1746 GND.n1689 0.0636886
R6526 GND.n1764 GND.n1763 0.0636886
R6527 GND.t296 GND.n1764 0.0636886
R6528 GND.n1705 GND.n1704 0.0636886
R6529 GND.n1746 GND.n1705 0.0636886
R6530 GND.n1700 GND.n1699 0.0636886
R6531 GND.n1746 GND.n1700 0.0636886
R6532 GND.n1766 GND.n1765 0.0636886
R6533 GND.t296 GND.n1766 0.0636886
R6534 GND.n1715 GND.n1714 0.0636886
R6535 GND.n1746 GND.n1715 0.0636886
R6536 GND.n1711 GND.n1710 0.0636886
R6537 GND.n1746 GND.n1711 0.0636886
R6538 GND.n1768 GND.n1767 0.0636886
R6539 GND.t296 GND.n1768 0.0636886
R6540 GND.n1725 GND.n1724 0.0636886
R6541 GND.n1746 GND.n1725 0.0636886
R6542 GND.n1719 GND.n1718 0.0636886
R6543 GND.n1746 GND.n1719 0.0636886
R6544 GND.n1770 GND.n1769 0.0636886
R6545 GND.t296 GND.n1770 0.0636886
R6546 GND.n1735 GND.n1734 0.0636886
R6547 GND.n1746 GND.n1735 0.0636886
R6548 GND.n1731 GND.n1730 0.0636886
R6549 GND.n1746 GND.n1731 0.0636886
R6550 GND.n1772 GND.n1771 0.0636886
R6551 GND.t296 GND.n1772 0.0636886
R6552 GND.n1745 GND.n1744 0.0636886
R6553 GND.n1746 GND.n1745 0.0636886
R6554 GND.n1740 GND.n1739 0.0636886
R6555 GND.n1746 GND.n1740 0.0636886
R6556 GND.n1774 GND.n1773 0.0636886
R6557 GND.t296 GND.n1774 0.0636886
R6558 GND.n4790 GND.n4789 0.0636886
R6559 GND.n4791 GND.n4790 0.0636886
R6560 GND.n4785 GND.n4784 0.0636886
R6561 GND.n4791 GND.n4785 0.0636886
R6562 GND.n4795 GND.n4794 0.0636886
R6563 GND.t293 GND.n4795 0.0636886
R6564 GND.n4780 GND.n4779 0.0636886
R6565 GND.n4791 GND.n4780 0.0636886
R6566 GND.n4774 GND.n4773 0.0636886
R6567 GND.n4791 GND.n4774 0.0636886
R6568 GND.n4793 GND.n4792 0.0636886
R6569 GND.t293 GND.n4793 0.0636886
R6570 GND.n4760 GND.n4759 0.0636886
R6571 GND.n4761 GND.n4760 0.0636886
R6572 GND.n4763 GND.n4762 0.0636886
R6573 GND.n4762 GND.n4761 0.0636886
R6574 GND.n4692 GND.n4691 0.0636886
R6575 GND.n4691 GND.t552 0.0636886
R6576 GND.t552 GND.n4690 0.0636886
R6577 GND.n4690 GND.n4689 0.0636886
R6578 GND.n4676 GND.n4675 0.0636886
R6579 GND.n4675 GND.t535 0.0636886
R6580 GND.n6350 GND.n6349 0.0636834
R6581 GND.n7804 GND.n24 0.0636834
R6582 GND.n6380 GND 0.0628765
R6583 GND GND.n7799 0.0628765
R6584 GND.n1445 GND.n1444 0.0612287
R6585 GND.n681 GND.n677 0.0610263
R6586 GND.n685 GND.n677 0.0610263
R6587 GND.n686 GND.n685 0.0610263
R6588 GND.n687 GND.n686 0.0610263
R6589 GND.n698 GND.n674 0.0610263
R6590 GND.n698 GND.n671 0.0610263
R6591 GND.n671 GND.n668 0.0610263
R6592 GND.n703 GND.n668 0.0610263
R6593 GND.n6245 GND.n6241 0.0610263
R6594 GND.n6249 GND.n6241 0.0610263
R6595 GND.n6250 GND.n6249 0.0610263
R6596 GND.n6251 GND.n6250 0.0610263
R6597 GND.n6262 GND.n6238 0.0610263
R6598 GND.n6262 GND.n6235 0.0610263
R6599 GND.n6235 GND.n6232 0.0610263
R6600 GND.n6267 GND.n6232 0.0610263
R6601 GND.n3353 GND 0.060284
R6602 GND.n305 GND 0.060284
R6603 GND.n203 GND 0.060284
R6604 GND.n2656 GND 0.060284
R6605 GND.n3082 GND 0.060284
R6606 GND.n6963 GND 0.060284
R6607 GND.n6800 GND 0.060284
R6608 GND.n7745 GND 0.060284
R6609 GND.n5625 GND 0.060284
R6610 GND.n5441 GND 0.060284
R6611 GND.n499 GND 0.060284
R6612 GND.n5143 GND 0.060284
R6613 GND.n3743 GND 0.060284
R6614 GND.n3420 GND 0.060284
R6615 GND.n640 GND 0.060284
R6616 GND.n2347 GND 0.060284
R6617 GND.n6408 GND.n541 0.0593951
R6618 GND.n4456 GND.n4454 0.0589677
R6619 GND.n2058 GND.n2057 0.0588369
R6620 GND.n2823 GND.n2822 0.0588369
R6621 GND.n4900 GND.n4899 0.0588344
R6622 GND.n4699 GND.n4698 0.0588344
R6623 GND.n3155 GND.n3154 0.0588344
R6624 GND.n2284 GND.n2283 0.0588344
R6625 GND.n7688 GND.n7687 0.0588344
R6626 GND.n1544 GND.n1543 0.0588344
R6627 GND.n5381 GND.n5380 0.0588344
R6628 GND.n3950 GND.n3949 0.0588344
R6629 GND.n5242 GND.n5241 0.0588344
R6630 GND.n3842 GND.n3841 0.0588344
R6631 GND.n3519 GND.n3518 0.0588344
R6632 GND.n1971 GND.n1970 0.0588344
R6633 GND.n2446 GND.n2445 0.0588344
R6634 GND.n2755 GND.n2754 0.0588344
R6635 GND.n3256 GND.n3255 0.0582982
R6636 GND.n7559 GND.n7558 0.0582982
R6637 GND.n7621 GND.n7620 0.0582982
R6638 GND.n2520 GND.n2516 0.0582982
R6639 GND.n2937 GND.n2933 0.0582982
R6640 GND.n6959 GND.n6958 0.0582982
R6641 GND.n6796 GND.n6795 0.0582982
R6642 GND.n85 GND.n84 0.0582982
R6643 GND.n1029 GND.n1028 0.0582982
R6644 GND.n1258 GND.n1254 0.0582982
R6645 GND.n7497 GND.n7496 0.0582982
R6646 GND.n4996 GND.n4995 0.0582982
R6647 GND.n3602 GND.n3598 0.0582982
R6648 GND.n1128 GND.n1127 0.0582982
R6649 GND.n6550 GND.n6549 0.0582982
R6650 GND.n7128 GND.n7127 0.0582982
R6651 GND.n4366 GND.n4364 0.0581389
R6652 GND.n6486 GND.n6485 0.0580634
R6653 GND.n6396 GND.n6395 0.0580634
R6654 GND.n23 GND.n6 0.0580441
R6655 GND.n7791 GND.n7764 0.0580441
R6656 GND.n659 GND.n658 0.0580441
R6657 GND.n665 GND.n642 0.0580441
R6658 GND.n6348 GND.n6331 0.0580441
R6659 GND.n6324 GND.n6297 0.0580441
R6660 GND.n6287 GND.n6286 0.0580441
R6661 GND.n6293 GND.n6270 0.0580441
R6662 GND.n6449 GND 0.058
R6663 GND.n6443 GND 0.058
R6664 GND.n6431 GND 0.058
R6665 GND.n534 GND 0.058
R6666 GND.n528 GND 0.058
R6667 GND.n516 GND 0.058
R6668 GND.n4577 GND.n4574 0.0570476
R6669 GND.n3333 GND.n3259 0.05675
R6670 GND.n7520 GND.n306 0.05675
R6671 GND.n7582 GND.n204 0.05675
R6672 GND.n2636 GND.n2523 0.05675
R6673 GND.n3062 GND.n2940 0.05675
R6674 GND.n6972 GND.n6928 0.05675
R6675 GND.n6818 GND.n6774 0.05675
R6676 GND.n7752 GND.n7751 0.05675
R6677 GND.n5634 GND.n998 0.05675
R6678 GND.n5450 GND.n1227 0.05675
R6679 GND.n7458 GND.n500 0.05675
R6680 GND.n5123 GND.n4999 0.05675
R6681 GND.n3723 GND.n3605 0.05675
R6682 GND.n5507 GND.n1106 0.05675
R6683 GND.n6511 GND.n641 0.05675
R6684 GND.n7089 GND.n7078 0.05675
R6685 GND.n6489 GND.n6480 0.05675
R6686 GND.n6490 GND.n6478 0.05675
R6687 GND.n6399 GND.n6390 0.05675
R6688 GND.n6400 GND.n6388 0.05675
R6689 GND.n7780 GND.n7779 0.0567153
R6690 GND.n6313 GND.n6312 0.0567153
R6691 GND.n3343 GND.n3342 0.0560434
R6692 GND.n7530 GND.n7529 0.0560434
R6693 GND.n7592 GND.n7591 0.0560434
R6694 GND.n2646 GND.n2645 0.0560434
R6695 GND.n3072 GND.n3071 0.0560434
R6696 GND.n6938 GND.n6937 0.0560434
R6697 GND.n63 GND.n62 0.0560434
R6698 GND.n1008 GND.n1007 0.0560434
R6699 GND.n1237 GND.n1236 0.0560434
R6700 GND.n7468 GND.n7467 0.0560434
R6701 GND.n5133 GND.n5132 0.0560434
R6702 GND.n3733 GND.n3732 0.0560434
R6703 GND.n7099 GND.n7098 0.0560434
R6704 GND.n6456 GND.n6455 0.0558279
R6705 GND.n7438 GND.n540 0.0558279
R6706 GND.n6437 GND 0.0555
R6707 GND.n522 GND 0.0555
R6708 GND.n3349 GND.n3333 0.05425
R6709 GND.n7536 GND.n7520 0.05425
R6710 GND.n7598 GND.n7582 0.05425
R6711 GND.n2652 GND.n2636 0.05425
R6712 GND.n3078 GND.n3062 0.05425
R6713 GND.n6972 GND.n6971 0.05425
R6714 GND.n6818 GND.n6817 0.05425
R6715 GND.n5634 GND.n5633 0.05425
R6716 GND.n5450 GND.n5449 0.05425
R6717 GND.n7474 GND.n7458 0.05425
R6718 GND.n5139 GND.n5123 0.05425
R6719 GND.n3739 GND.n3723 0.05425
R6720 GND.n5507 GND.n5506 0.05425
R6721 GND.n6527 GND.n6511 0.05425
R6722 GND.n7105 GND.n7089 0.05425
R6723 GND.n4104 GND.n4103 0.0540714
R6724 GND.n6815 GND.n6814 0.0532741
R6725 GND.n64 GND.n63 0.0532741
R6726 GND.n5504 GND.n5503 0.0532741
R6727 GND.n6525 GND.n6524 0.0532741
R6728 GND.n4480 GND.n4478 0.0530794
R6729 GND.n691 GND.n690 0.052907
R6730 GND.n6255 GND.n6254 0.052907
R6731 GND.n4800 GND.n4797 0.0528195
R6732 GND.n1834 GND.n1833 0.0528195
R6733 GND.n1844 GND.n1843 0.0528195
R6734 GND.n1839 GND.n1838 0.0528195
R6735 GND.n1824 GND.n1823 0.0528195
R6736 GND.n1814 GND.n1813 0.0528195
R6737 GND.n1804 GND.n1803 0.0528195
R6738 GND.n1794 GND.n1793 0.0528195
R6739 GND.n1779 GND.n1776 0.0528195
R6740 GND.n1784 GND.n1783 0.0528195
R6741 GND.n1789 GND.n1788 0.0528195
R6742 GND.n1799 GND.n1798 0.0528195
R6743 GND.n1809 GND.n1808 0.0528195
R6744 GND.n1819 GND.n1818 0.0528195
R6745 GND.n1829 GND.n1828 0.0528195
R6746 GND.n3337 GND 0.0527727
R6747 GND.n7524 GND 0.0527727
R6748 GND.n7586 GND 0.0527727
R6749 GND.n2640 GND 0.0527727
R6750 GND.n3066 GND 0.0527727
R6751 GND.n6932 GND 0.0527727
R6752 GND.n6809 GND 0.0527727
R6753 GND.n57 GND 0.0527727
R6754 GND.n1002 GND 0.0527727
R6755 GND.n1231 GND 0.0527727
R6756 GND.n7462 GND 0.0527727
R6757 GND.n5127 GND 0.0527727
R6758 GND.n3727 GND 0.0527727
R6759 GND.n5498 GND 0.0527727
R6760 GND.n6519 GND 0.0527727
R6761 GND.n7093 GND 0.0527727
R6762 GND.n3364 GND.n3363 0.0525185
R6763 GND.n3365 GND.n3364 0.0525185
R6764 GND.n3370 GND.n3369 0.0525185
R6765 GND.n3371 GND.n3370 0.0525185
R6766 GND.n3358 GND.n3357 0.0525185
R6767 GND.n3359 GND.n3358 0.0525185
R6768 GND.n3096 GND.n3095 0.0525185
R6769 GND.n3097 GND.n3096 0.0525185
R6770 GND.n3090 GND.n3089 0.0525185
R6771 GND.n3091 GND.n3090 0.0525185
R6772 GND.n3107 GND.n3106 0.0525185
R6773 GND.n3108 GND.n3107 0.0525185
R6774 GND.n3087 GND.n3086 0.0525185
R6775 GND.n3088 GND.n3087 0.0525185
R6776 GND.n3104 GND.n3103 0.0525185
R6777 GND.n3105 GND.n3104 0.0525185
R6778 GND.n4019 GND.n4018 0.0525185
R6779 GND.n4020 GND.n4019 0.0525185
R6780 GND.n4013 GND.n4012 0.0525185
R6781 GND.n4014 GND.n4013 0.0525185
R6782 GND.n4030 GND.n4029 0.0525185
R6783 GND.n4031 GND.n4030 0.0525185
R6784 GND.n4010 GND.n4009 0.0525185
R6785 GND.n4011 GND.n4010 0.0525185
R6786 GND.n4027 GND.n4026 0.0525185
R6787 GND.n4028 GND.n4027 0.0525185
R6788 GND.n5158 GND.n5157 0.0525185
R6789 GND.n5159 GND.n5158 0.0525185
R6790 GND.n5149 GND.n5148 0.0525185
R6791 GND.n5150 GND.n5149 0.0525185
R6792 GND.n5182 GND.n5181 0.0525185
R6793 GND.n5183 GND.n5182 0.0525185
R6794 GND.n5152 GND.n5151 0.0525185
R6795 GND.n5153 GND.n5152 0.0525185
R6796 GND.n5185 GND.n5184 0.0525185
R6797 GND.n5186 GND.n5185 0.0525185
R6798 GND.n3757 GND.n3756 0.0525185
R6799 GND.n3758 GND.n3757 0.0525185
R6800 GND.n3751 GND.n3750 0.0525185
R6801 GND.n3752 GND.n3751 0.0525185
R6802 GND.n3784 GND.n3783 0.0525185
R6803 GND.n3785 GND.n3784 0.0525185
R6804 GND.n3748 GND.n3747 0.0525185
R6805 GND.n3749 GND.n3748 0.0525185
R6806 GND.n3781 GND.n3780 0.0525185
R6807 GND.n3782 GND.n3781 0.0525185
R6808 GND.n1292 GND.n1291 0.0525185
R6809 GND.n1293 GND.n1292 0.0525185
R6810 GND.n1283 GND.n1282 0.0525185
R6811 GND.n1284 GND.n1283 0.0525185
R6812 GND.n1316 GND.n1315 0.0525185
R6813 GND.n1317 GND.n1316 0.0525185
R6814 GND.n1286 GND.n1285 0.0525185
R6815 GND.n1287 GND.n1286 0.0525185
R6816 GND.n1319 GND.n1318 0.0525185
R6817 GND.n1320 GND.n1319 0.0525185
R6818 GND.n3435 GND.n3434 0.0525185
R6819 GND.n3436 GND.n3435 0.0525185
R6820 GND.n3429 GND.n3428 0.0525185
R6821 GND.n3430 GND.n3429 0.0525185
R6822 GND.n3462 GND.n3461 0.0525185
R6823 GND.n3463 GND.n3462 0.0525185
R6824 GND.n3426 GND.n3425 0.0525185
R6825 GND.n3427 GND.n3426 0.0525185
R6826 GND.n3459 GND.n3458 0.0525185
R6827 GND.n3460 GND.n3459 0.0525185
R6828 GND.n1460 GND.n1459 0.0525185
R6829 GND.n1461 GND.n1460 0.0525185
R6830 GND.n1451 GND.n1450 0.0525185
R6831 GND.n1452 GND.n1451 0.0525185
R6832 GND.n1484 GND.n1483 0.0525185
R6833 GND.n1485 GND.n1484 0.0525185
R6834 GND.n1454 GND.n1453 0.0525185
R6835 GND.n1455 GND.n1454 0.0525185
R6836 GND.n1487 GND.n1486 0.0525185
R6837 GND.n1488 GND.n1487 0.0525185
R6838 GND.n1886 GND.n1885 0.0525185
R6839 GND.n1887 GND.n1886 0.0525185
R6840 GND.n1880 GND.n1879 0.0525185
R6841 GND.n1881 GND.n1880 0.0525185
R6842 GND.n1913 GND.n1912 0.0525185
R6843 GND.n1914 GND.n1913 0.0525185
R6844 GND.n1877 GND.n1876 0.0525185
R6845 GND.n1878 GND.n1877 0.0525185
R6846 GND.n1910 GND.n1909 0.0525185
R6847 GND.n1911 GND.n1910 0.0525185
R6848 GND.n101 GND.n100 0.0525185
R6849 GND.n102 GND.n101 0.0525185
R6850 GND.n94 GND.n93 0.0525185
R6851 GND.n95 GND.n94 0.0525185
R6852 GND.n133 GND.n132 0.0525185
R6853 GND.n134 GND.n133 0.0525185
R6854 GND.n92 GND.n91 0.0525185
R6855 GND.n96 GND.n92 0.0525185
R6856 GND.n136 GND.n135 0.0525185
R6857 GND.n137 GND.n136 0.0525185
R6858 GND.n2137 GND.n2136 0.0525185
R6859 GND.n2138 GND.n2137 0.0525185
R6860 GND.n2131 GND.n2130 0.0525185
R6861 GND.n2132 GND.n2131 0.0525185
R6862 GND.n2164 GND.n2163 0.0525185
R6863 GND.n2165 GND.n2164 0.0525185
R6864 GND.n2128 GND.n2127 0.0525185
R6865 GND.n2129 GND.n2128 0.0525185
R6866 GND.n2161 GND.n2160 0.0525185
R6867 GND.n2162 GND.n2161 0.0525185
R6868 GND.n2199 GND.n2198 0.0525185
R6869 GND.n2200 GND.n2199 0.0525185
R6870 GND.n2190 GND.n2189 0.0525185
R6871 GND.n2191 GND.n2190 0.0525185
R6872 GND.n2223 GND.n2222 0.0525185
R6873 GND.n2224 GND.n2223 0.0525185
R6874 GND.n2193 GND.n2192 0.0525185
R6875 GND.n2194 GND.n2193 0.0525185
R6876 GND.n2226 GND.n2225 0.0525185
R6877 GND.n2227 GND.n2226 0.0525185
R6878 GND.n2362 GND.n2361 0.0525185
R6879 GND.n2363 GND.n2362 0.0525185
R6880 GND.n2353 GND.n2352 0.0525185
R6881 GND.n2357 GND.n2353 0.0525185
R6882 GND.n2389 GND.n2388 0.0525185
R6883 GND.n2390 GND.n2389 0.0525185
R6884 GND.n2355 GND.n2354 0.0525185
R6885 GND.n2356 GND.n2355 0.0525185
R6886 GND.n2386 GND.n2385 0.0525185
R6887 GND.n2387 GND.n2386 0.0525185
R6888 GND.n2674 GND.n2673 0.0525185
R6889 GND.n2675 GND.n2674 0.0525185
R6890 GND.n2668 GND.n2667 0.0525185
R6891 GND.n2669 GND.n2668 0.0525185
R6892 GND.n2683 GND.n2682 0.0525185
R6893 GND.n2684 GND.n2683 0.0525185
R6894 GND.n2680 GND.n2679 0.0525185
R6895 GND.n2681 GND.n2680 0.0525185
R6896 GND.n2665 GND.n2664 0.0525185
R6897 GND.n2666 GND.n2665 0.0525185
R6898 GND.n4815 GND.n4814 0.0525185
R6899 GND.n4816 GND.n4815 0.0525185
R6900 GND.n4809 GND.n4808 0.0525185
R6901 GND.n4810 GND.n4809 0.0525185
R6902 GND.n4842 GND.n4841 0.0525185
R6903 GND.n4843 GND.n4842 0.0525185
R6904 GND.n4806 GND.n4805 0.0525185
R6905 GND.n4807 GND.n4806 0.0525185
R6906 GND.n4839 GND.n4838 0.0525185
R6907 GND.n4840 GND.n4839 0.0525185
R6908 GND.n4599 GND.n4598 0.0525185
R6909 GND.n4600 GND.n4599 0.0525185
R6910 GND.n4632 GND.n4631 0.0525185
R6911 GND.n4633 GND.n4632 0.0525185
R6912 GND.n4608 GND.n4607 0.0525185
R6913 GND.n4609 GND.n4608 0.0525185
R6914 GND.n4602 GND.n4601 0.0525185
R6915 GND.n4603 GND.n4602 0.0525185
R6916 GND.n4635 GND.n4634 0.0525185
R6917 GND.n4636 GND.n4635 0.0525185
R6918 GND.n4705 GND.n4704 0.0525185
R6919 GND.n4706 GND.n4705 0.0525185
R6920 GND.n4756 GND.n4755 0.0525185
R6921 GND.n4755 GND.n4754 0.0525185
R6922 GND.n1843 GND.n1842 0.0523204
R6923 GND.n1838 GND.n1837 0.0523204
R6924 GND.n1833 GND.n1832 0.0523204
R6925 GND.n1828 GND.n1827 0.0523204
R6926 GND.n1823 GND.n1822 0.0523204
R6927 GND.n1818 GND.n1817 0.0523204
R6928 GND.n1813 GND.n1812 0.0523204
R6929 GND.n1808 GND.n1807 0.0523204
R6930 GND.n1803 GND.n1802 0.0523204
R6931 GND.n1798 GND.n1797 0.0523204
R6932 GND.n1793 GND.n1792 0.0523204
R6933 GND.n1788 GND.n1787 0.0523204
R6934 GND.n1783 GND.n1782 0.0523204
R6935 GND.n1776 GND.n1775 0.0523204
R6936 GND.n4797 GND.n4796 0.0523204
R6937 GND.n4961 GND.n4960 0.0523204
R6938 GND.n4964 GND.n4961 0.0523204
R6939 GND.n3332 GND.n3331 0.0516364
R6940 GND.n7519 GND.n7518 0.0516364
R6941 GND.n7581 GND.n7580 0.0516364
R6942 GND.n2635 GND.n2634 0.0516364
R6943 GND.n3061 GND.n3060 0.0516364
R6944 GND.n6974 GND.n6973 0.0516364
R6945 GND.n6820 GND.n6819 0.0516364
R6946 GND.n7754 GND.n7753 0.0516364
R6947 GND.n5636 GND.n5635 0.0516364
R6948 GND.n5452 GND.n5451 0.0516364
R6949 GND.n7457 GND.n7456 0.0516364
R6950 GND.n5122 GND.n5121 0.0516364
R6951 GND.n3722 GND.n3721 0.0516364
R6952 GND.n5509 GND.n5508 0.0516364
R6953 GND.n6510 GND.n6509 0.0516364
R6954 GND.n7088 GND.n7087 0.0516364
R6955 GND.n6379 GND.n666 0.0500734
R6956 GND.n7563 GND.n7562 0.0494583
R6957 GND.n7625 GND.n7624 0.0494583
R6958 GND.n2530 GND.n2529 0.0494583
R6959 GND.n2953 GND.n2952 0.0494583
R6960 GND.n6961 GND.n6924 0.0494583
R6961 GND.n6798 GND.n6770 0.0494583
R6962 GND.n6662 GND.n6661 0.0494583
R6963 GND.n5623 GND.n5622 0.0494583
R6964 GND.n1276 GND.n1275 0.0494583
R6965 GND.n7501 GND.n7500 0.0494583
R6966 GND.n5012 GND.n5011 0.0494583
R6967 GND.n3618 GND.n3617 0.0494583
R6968 GND.n5488 GND.n5487 0.0494583
R6969 GND.n6554 GND.n6553 0.0494583
R6970 GND.n7132 GND.n7131 0.0494583
R6971 GND.n3272 GND.n3260 0.0494583
R6972 GND.n7753 GND.n7750 0.0493636
R6973 GND GND.n680 0.0490201
R6974 GND GND.n6244 0.0490201
R6975 GND.n3257 GND.n3247 0.0486039
R6976 GND.n7560 GND.n7550 0.0486039
R6977 GND.n7622 GND.n7612 0.0486039
R6978 GND.n2521 GND.n2508 0.0486039
R6979 GND.n2938 GND.n2925 0.0486039
R6980 GND.n6960 GND.n6950 0.0486039
R6981 GND.n6797 GND.n6787 0.0486039
R6982 GND.n86 GND.n76 0.0486039
R6983 GND.n1030 GND.n1020 0.0486039
R6984 GND.n1259 GND.n1246 0.0486039
R6985 GND.n7498 GND.n7488 0.0486039
R6986 GND.n4997 GND.n4987 0.0486039
R6987 GND.n3603 GND.n3590 0.0486039
R6988 GND.n1129 GND.n1119 0.0486039
R6989 GND.n6551 GND.n6541 0.0486039
R6990 GND.n7129 GND.n7119 0.0486039
R6991 GND.n36 GND 0.0484167
R6992 GND GND.n25 0.0484167
R6993 GND.n3250 GND 0.0484167
R6994 GND.n7553 GND 0.0484167
R6995 GND.n7615 GND 0.0484167
R6996 GND.n2511 GND 0.0484167
R6997 GND.n2928 GND 0.0484167
R6998 GND.n6954 GND 0.0484167
R6999 GND.n6790 GND 0.0484167
R7000 GND.n80 GND 0.0484167
R7001 GND.n1023 GND 0.0484167
R7002 GND.n1250 GND 0.0484167
R7003 GND.n7492 GND 0.0484167
R7004 GND.n4991 GND 0.0484167
R7005 GND.n3593 GND 0.0484167
R7006 GND.n1122 GND 0.0484167
R7007 GND.n6544 GND 0.0484167
R7008 GND.n7122 GND 0.0484167
R7009 GND.n6363 GND 0.0484167
R7010 GND GND.n6352 0.0484167
R7011 GND.n3342 GND.n3341 0.0483725
R7012 GND.n7529 GND.n7528 0.0483725
R7013 GND.n7591 GND.n7590 0.0483725
R7014 GND.n2645 GND.n2644 0.0483725
R7015 GND.n3071 GND.n3070 0.0483725
R7016 GND.n6937 GND.n6936 0.0483725
R7017 GND.n6814 GND.n6813 0.0483725
R7018 GND.n63 GND.n61 0.0483725
R7019 GND.n1007 GND.n1006 0.0483725
R7020 GND.n1236 GND.n1235 0.0483725
R7021 GND.n7467 GND.n7466 0.0483725
R7022 GND.n5132 GND.n5131 0.0483725
R7023 GND.n3732 GND.n3731 0.0483725
R7024 GND.n5503 GND.n5502 0.0483725
R7025 GND.n6524 GND.n6523 0.0483725
R7026 GND.n7098 GND.n7097 0.0483725
R7027 GND.n4558 GND.n4556 0.048348
R7028 GND.n4954 GND.n4953 0.0483051
R7029 GND.n4972 GND.n4970 0.0483051
R7030 GND.n3401 GND.n3399 0.0483051
R7031 GND.n3143 GND.n3141 0.0483051
R7032 GND.n2345 GND.n2343 0.0483051
R7033 GND.n1866 GND.n1865 0.0483051
R7034 GND.n5329 GND.n5327 0.0483051
R7035 GND.n3576 GND.n1333 0.0483051
R7036 GND.n5315 GND.n5314 0.0483051
R7037 GND.n5309 GND.n5307 0.0483051
R7038 GND.n3897 GND.n3896 0.0483051
R7039 GND.n3570 GND.n3569 0.0483051
R7040 GND.n3413 GND.n3412 0.0483051
R7041 GND.n2184 GND.n2182 0.0483051
R7042 GND.n2499 GND.n2497 0.0483051
R7043 GND.n2814 GND.n2812 0.0483051
R7044 GND.n3247 GND.n3246 0.0464802
R7045 GND.n7550 GND.n7549 0.0464802
R7046 GND.n7612 GND.n7611 0.0464802
R7047 GND.n6950 GND.n6949 0.0464802
R7048 GND.n6787 GND.n6786 0.0464802
R7049 GND.n76 GND.n75 0.0464802
R7050 GND.n1020 GND.n1019 0.0464802
R7051 GND.n7488 GND.n7487 0.0464802
R7052 GND.n4987 GND.n4986 0.0464802
R7053 GND.n1119 GND.n1118 0.0464802
R7054 GND.n6541 GND.n6540 0.0464802
R7055 GND.n7119 GND.n7118 0.0464802
R7056 GND.n7792 GND 0.04425
R7057 GND.n6325 GND 0.04425
R7058 GND.n3409 GND.n3408 0.0436389
R7059 GND.n3300 GND.n3299 0.0425017
R7060 GND.n3299 GND.n3298 0.0425017
R7061 GND.n2961 GND.n2960 0.0425017
R7062 GND.n2962 GND.n2961 0.0425017
R7063 GND.n2992 GND.n2991 0.0425017
R7064 GND.n2991 GND.n2990 0.0425017
R7065 GND.n2537 GND.n2536 0.0425017
R7066 GND.n2538 GND.n2537 0.0425017
R7067 GND.n2566 GND.n2565 0.0425017
R7068 GND.n2565 GND.n2564 0.0425017
R7069 GND.n7142 GND.n7141 0.0425017
R7070 GND.n7143 GND.n7142 0.0425017
R7071 GND.n7166 GND.n7165 0.0425017
R7072 GND.n7165 GND.n7164 0.0425017
R7073 GND.n605 GND.n604 0.0425017
R7074 GND.n606 GND.n605 0.0425017
R7075 GND.n7003 GND.n7002 0.0425017
R7076 GND.n7002 GND.n7001 0.0425017
R7077 GND.n615 GND.n614 0.0425017
R7078 GND.n616 GND.n615 0.0425017
R7079 GND.n6849 GND.n6848 0.0425017
R7080 GND.n6848 GND.n6847 0.0425017
R7081 GND.n625 GND.n624 0.0425017
R7082 GND.n626 GND.n625 0.0425017
R7083 GND.n6695 GND.n6694 0.0425017
R7084 GND.n6694 GND.n6693 0.0425017
R7085 GND.n632 GND.n631 0.0425017
R7086 GND.n633 GND.n632 0.0425017
R7087 GND.n6624 GND.n6623 0.0425017
R7088 GND.n6623 GND.n6622 0.0425017
R7089 GND.n5611 GND.n5610 0.0425017
R7090 GND.n5612 GND.n5611 0.0425017
R7091 GND.n5576 GND.n5575 0.0425017
R7092 GND.n5575 GND.n5574 0.0425017
R7093 GND.n5476 GND.n5475 0.0425017
R7094 GND.n5477 GND.n5476 0.0425017
R7095 GND.n1074 GND.n1073 0.0425017
R7096 GND.n1073 GND.n1072 0.0425017
R7097 GND.n1133 GND.n1132 0.0425017
R7098 GND.n1134 GND.n1133 0.0425017
R7099 GND.n1195 GND.n1194 0.0425017
R7100 GND.n1194 GND.n1193 0.0425017
R7101 GND.n3625 GND.n3624 0.0425017
R7102 GND.n3626 GND.n3625 0.0425017
R7103 GND.n3656 GND.n3655 0.0425017
R7104 GND.n3655 GND.n3654 0.0425017
R7105 GND.n5019 GND.n5018 0.0425017
R7106 GND.n5020 GND.n5019 0.0425017
R7107 GND.n5053 GND.n5052 0.0425017
R7108 GND.n5052 GND.n5051 0.0425017
R7109 GND.n414 GND.n413 0.0425017
R7110 GND.n415 GND.n414 0.0425017
R7111 GND.n448 GND.n447 0.0425017
R7112 GND.n447 GND.n446 0.0425017
R7113 GND.n310 GND.n309 0.0425017
R7114 GND.n311 GND.n310 0.0425017
R7115 GND.n379 GND.n378 0.0425017
R7116 GND.n378 GND.n377 0.0425017
R7117 GND.n208 GND.n207 0.0425017
R7118 GND.n209 GND.n208 0.0425017
R7119 GND.n275 GND.n274 0.0425017
R7120 GND.n274 GND.n273 0.0425017
R7121 GND.n190 GND.n189 0.0425017
R7122 GND.n191 GND.n190 0.0425017
R7123 GND.n4651 GND.n4650 0.0415714
R7124 GND.n3203 GND.n3202 0.0415714
R7125 GND.n2252 GND.n2251 0.0415714
R7126 GND.n152 GND.n151 0.0415714
R7127 GND.n1512 GND.n1511 0.0415714
R7128 GND.n5349 GND.n5348 0.0415714
R7129 GND.n3918 GND.n3917 0.0415714
R7130 GND.n5210 GND.n5209 0.0415714
R7131 GND.n3810 GND.n3809 0.0415714
R7132 GND.n3487 GND.n3486 0.0415714
R7133 GND.n1939 GND.n1938 0.0415714
R7134 GND.n2033 GND.n2032 0.0415714
R7135 GND.n2414 GND.n2413 0.0415714
R7136 GND.n2723 GND.n2722 0.0415714
R7137 GND.n4868 GND.n4867 0.0415714
R7138 GND.n2833 GND.n2832 0.0415714
R7139 GND.n4670 GND.n4669 0.0406786
R7140 GND.n3207 GND.n3204 0.0406786
R7141 GND.n2254 GND.n2253 0.0406786
R7142 GND.n7667 GND.n7666 0.0406786
R7143 GND.n1514 GND.n1513 0.0406786
R7144 GND.n5351 GND.n5350 0.0406786
R7145 GND.n3920 GND.n3919 0.0406786
R7146 GND.n5212 GND.n5211 0.0406786
R7147 GND.n3812 GND.n3811 0.0406786
R7148 GND.n3489 GND.n3488 0.0406786
R7149 GND.n1941 GND.n1940 0.0406786
R7150 GND.n2051 GND.n2050 0.0406786
R7151 GND.n2416 GND.n2415 0.0406786
R7152 GND.n2725 GND.n2724 0.0406786
R7153 GND.n4870 GND.n4869 0.0406786
R7154 GND.n2835 GND.n2834 0.0406786
R7155 GND.n1427 GND.n1426 0.0390862
R7156 GND.n4801 GND 0.0386944
R7157 GND.n4971 GND 0.0386944
R7158 GND.n3400 GND 0.0386944
R7159 GND.n3142 GND 0.0386944
R7160 GND.n2344 GND 0.0386944
R7161 GND.n1864 GND 0.0386944
R7162 GND.n5328 GND 0.0386944
R7163 GND.n1332 GND 0.0386944
R7164 GND.n3906 GND 0.0386944
R7165 GND.n5308 GND 0.0386944
R7166 GND.n3582 GND 0.0386944
R7167 GND.n3419 GND 0.0386944
R7168 GND.n1872 GND 0.0386944
R7169 GND.n2183 GND 0.0386944
R7170 GND.n2498 GND 0.0386944
R7171 GND.n2813 GND 0.0386944
R7172 GND.n4566 GND.n4564 0.0381984
R7173 GND.n4454 GND.n4452 0.0367903
R7174 GND.n4976 GND.n4975 0.0363684
R7175 GND.n7798 GND.n24 0.0356562
R7176 GND.n6351 GND.n6350 0.0356562
R7177 GND.n704 GND 0.0353684
R7178 GND.n6268 GND 0.0353684
R7179 GND.n6209 GND.n6208 0.0352222
R7180 GND.n5335 GND.n5334 0.0351316
R7181 GND.n303 GND.n302 0.0345278
R7182 GND.n7629 GND.n7627 0.0345278
R7183 GND.n2526 GND.n2525 0.0345278
R7184 GND.n2945 GND.n2944 0.0345278
R7185 GND.n6921 GND.n6920 0.0345278
R7186 GND.n6767 GND.n6766 0.0345278
R7187 GND.n6652 GND.n6651 0.0345278
R7188 GND.n1102 GND.n1101 0.0345278
R7189 GND.n1264 GND.n1263 0.0345278
R7190 GND.n407 GND.n406 0.0345278
R7191 GND.n5004 GND.n5003 0.0345278
R7192 GND.n3610 GND.n3609 0.0345278
R7193 GND.n1223 GND.n1222 0.0345278
R7194 GND.n5604 GND.n5603 0.0345278
R7195 GND.n7075 GND.n7074 0.0345278
R7196 GND.n3265 GND.n3264 0.0345278
R7197 GND.n4073 GND.n4072 0.0339821
R7198 GND.n7562 GND.n7561 0.0337917
R7199 GND.n7624 GND.n7623 0.0337917
R7200 GND.n2529 GND.n2522 0.0337917
R7201 GND.n2952 GND.n2939 0.0337917
R7202 GND.n6962 GND.n6961 0.0337917
R7203 GND.n6799 GND.n6798 0.0337917
R7204 GND.n6661 GND.n87 0.0337917
R7205 GND.n5624 GND.n5623 0.0337917
R7206 GND.n1277 GND.n1276 0.0337917
R7207 GND.n7500 GND.n7499 0.0337917
R7208 GND.n5011 GND.n4998 0.0337917
R7209 GND.n3617 GND.n3604 0.0337917
R7210 GND.n5489 GND.n5488 0.0337917
R7211 GND.n6553 GND.n6552 0.0337917
R7212 GND.n7131 GND.n7130 0.0337917
R7213 GND.n3260 GND.n3258 0.0337917
R7214 GND.n6493 GND 0.033625
R7215 GND.n6403 GND 0.033625
R7216 GND.n3247 GND.n3243 0.0335935
R7217 GND.n7550 GND.n7546 0.0335935
R7218 GND.n7612 GND.n7608 0.0335935
R7219 GND.n2508 GND.n2507 0.0335935
R7220 GND.n2925 GND.n2924 0.0335935
R7221 GND.n6950 GND.n6946 0.0335935
R7222 GND.n6787 GND.n6783 0.0335935
R7223 GND.n76 GND.n72 0.0335935
R7224 GND.n1020 GND.n1016 0.0335935
R7225 GND.n1246 GND.n1245 0.0335935
R7226 GND.n7488 GND.n7484 0.0335935
R7227 GND.n4987 GND.n4983 0.0335935
R7228 GND.n3590 GND.n3589 0.0335935
R7229 GND.n1119 GND.n1115 0.0335935
R7230 GND.n6541 GND.n6537 0.0335935
R7231 GND.n7119 GND.n7115 0.0335935
R7232 GND GND.n6221 0.0324444
R7233 GND GND.n6211 0.0324444
R7234 GND.n658 GND 0.0324444
R7235 GND.n6286 GND 0.0324444
R7236 GND.n4092 GND.n4086 0.03175
R7237 GND.n7793 GND.n7792 0.03175
R7238 GND.n6326 GND.n6325 0.03175
R7239 GND.n5312 GND.n4976 0.0314211
R7240 GND.n6154 GND.n6152 0.0307632
R7241 GND.n6158 GND.n6154 0.0307632
R7242 GND.n6175 GND.n6171 0.0307632
R7243 GND.n6179 GND.n6175 0.0307632
R7244 GND.n6181 GND.n6179 0.0307632
R7245 GND.n6185 GND.n6181 0.0307632
R7246 GND.n6187 GND.n6185 0.0307632
R7247 GND.n6191 GND.n6187 0.0307632
R7248 GND.n6193 GND.n6191 0.0307632
R7249 GND.n5825 GND.n5824 0.0307632
R7250 GND.n5824 GND.n5822 0.0307632
R7251 GND.n5822 GND.n5818 0.0307632
R7252 GND.n5818 GND.n5816 0.0307632
R7253 GND.n5816 GND.n5812 0.0307632
R7254 GND.n5812 GND.n5810 0.0307632
R7255 GND.n5810 GND.n5806 0.0307632
R7256 GND.n5806 GND.n5802 0.0307632
R7257 GND.n5802 GND.n5800 0.0307632
R7258 GND.n5792 GND.n5788 0.0307632
R7259 GND.n5788 GND.n5786 0.0307632
R7260 GND.n5786 GND.n5782 0.0307632
R7261 GND.n5782 GND.n5780 0.0307632
R7262 GND.n5779 GND.n5778 0.0307632
R7263 GND.n5778 GND.n5776 0.0307632
R7264 GND.n5776 GND.n5772 0.0307632
R7265 GND.n5772 GND.n5770 0.0307632
R7266 GND.n5770 GND.n5766 0.0307632
R7267 GND.n5703 GND.n5699 0.0307632
R7268 GND.n5705 GND.n5703 0.0307632
R7269 GND.n5709 GND.n5705 0.0307632
R7270 GND.n5711 GND.n5709 0.0307632
R7271 GND.n5715 GND.n5711 0.0307632
R7272 GND.n5717 GND.n5715 0.0307632
R7273 GND.n5718 GND.n5717 0.0307632
R7274 GND.n5723 GND.n5721 0.0307632
R7275 GND.n5727 GND.n5723 0.0307632
R7276 GND.n5729 GND.n5727 0.0307632
R7277 GND.n5733 GND.n5729 0.0307632
R7278 GND.n5735 GND.n5733 0.0307632
R7279 GND.n681 GND 0.0307632
R7280 GND.n690 GND 0.0307632
R7281 GND.n6245 GND 0.0307632
R7282 GND.n6254 GND 0.0307632
R7283 GND.n4851 GND.n4850 0.0307537
R7284 GND.n4644 GND.n4643 0.0307537
R7285 GND.n2235 GND.n2234 0.0307537
R7286 GND.n2173 GND.n2172 0.0307537
R7287 GND.n145 GND.n144 0.0307537
R7288 GND.n1496 GND.n1495 0.0307537
R7289 GND.n1328 GND.n1327 0.0307537
R7290 GND.n5194 GND.n5193 0.0307537
R7291 GND.n3793 GND.n3792 0.0307537
R7292 GND.n3471 GND.n3470 0.0307537
R7293 GND.n1922 GND.n1921 0.0307537
R7294 GND.n2398 GND.n2397 0.0307537
R7295 GND.n705 GND.n704 0.0301053
R7296 GND.n6269 GND.n6268 0.0301053
R7297 GND GND.n4593 0.0300162
R7298 GND.n6211 GND.n6209 0.0296667
R7299 GND.n6208 GND.n6204 0.0296667
R7300 GND.n2658 GND.n2657 0.0296391
R7301 GND.n3101 GND.n3100 0.0296391
R7302 GND.n3390 GND.n3389 0.0296391
R7303 GND.n4024 GND.n4023 0.0296391
R7304 GND.n5748 GND.n5744 0.0294474
R7305 GND.n6494 GND.n6493 0.028625
R7306 GND.n6495 GND.n6494 0.028625
R7307 GND.n6404 GND.n6403 0.028625
R7308 GND.n6405 GND.n6404 0.028625
R7309 GND.n6224 GND.n6223 0.0284605
R7310 GND.n5800 GND.n5796 0.0282663
R7311 GND.n24 GND 0.0268889
R7312 GND.n6350 GND 0.0268889
R7313 GND.n5754 GND.n5735 0.0262926
R7314 GND.n5334 GND.n5333 0.0246184
R7315 GND.n6159 GND.n6158 0.0238553
R7316 GND.n5766 GND.n5764 0.0231974
R7317 GND.n5829 GND.n5828 0.0225395
R7318 GND.n5699 GND.n5697 0.0225395
R7319 GND.n6171 GND.n6169 0.0218816
R7320 GND.n6452 GND 0.02175
R7321 GND.n6446 GND 0.02175
R7322 GND.n6440 GND 0.02175
R7323 GND.n6434 GND 0.02175
R7324 GND.n6428 GND 0.02175
R7325 GND.n537 GND 0.02175
R7326 GND.n531 GND 0.02175
R7327 GND.n525 GND 0.02175
R7328 GND.n519 GND 0.02175
R7329 GND.n513 GND 0.02175
R7330 GND.n6227 GND.n6226 0.0212237
R7331 GND.n6458 GND.n6457 0.0209918
R7332 GND.n7440 GND.n7439 0.0209918
R7333 GND.n4654 GND.n4653 0.0208901
R7334 GND.n4657 GND.n4654 0.0208901
R7335 GND.n4662 GND.n4661 0.0208901
R7336 GND.n3198 GND.n3197 0.0208901
R7337 GND.n3201 GND.n3198 0.0208901
R7338 GND.n3213 GND.n3212 0.0208901
R7339 GND.n2247 GND.n2246 0.0208901
R7340 GND.n2250 GND.n2247 0.0208901
R7341 GND.n2260 GND.n2259 0.0208901
R7342 GND.n155 GND.n154 0.0208901
R7343 GND.n158 GND.n155 0.0208901
R7344 GND.n163 GND.n162 0.0208901
R7345 GND.n1507 GND.n1506 0.0208901
R7346 GND.n1510 GND.n1507 0.0208901
R7347 GND.n1520 GND.n1519 0.0208901
R7348 GND.n5344 GND.n5343 0.0208901
R7349 GND.n5347 GND.n5344 0.0208901
R7350 GND.n5357 GND.n5356 0.0208901
R7351 GND.n3913 GND.n3912 0.0208901
R7352 GND.n3916 GND.n3913 0.0208901
R7353 GND.n3926 GND.n3925 0.0208901
R7354 GND.n5205 GND.n5204 0.0208901
R7355 GND.n5208 GND.n5205 0.0208901
R7356 GND.n5218 GND.n5217 0.0208901
R7357 GND.n3805 GND.n3804 0.0208901
R7358 GND.n3808 GND.n3805 0.0208901
R7359 GND.n3818 GND.n3817 0.0208901
R7360 GND.n3482 GND.n3481 0.0208901
R7361 GND.n3485 GND.n3482 0.0208901
R7362 GND.n3495 GND.n3494 0.0208901
R7363 GND.n1934 GND.n1933 0.0208901
R7364 GND.n1937 GND.n1934 0.0208901
R7365 GND.n1947 GND.n1946 0.0208901
R7366 GND.n2036 GND.n2035 0.0208901
R7367 GND.n2039 GND.n2036 0.0208901
R7368 GND.n2044 GND.n2043 0.0208901
R7369 GND.n2409 GND.n2408 0.0208901
R7370 GND.n2412 GND.n2409 0.0208901
R7371 GND.n2422 GND.n2421 0.0208901
R7372 GND.n2718 GND.n2717 0.0208901
R7373 GND.n2721 GND.n2718 0.0208901
R7374 GND.n2731 GND.n2730 0.0208901
R7375 GND.n4863 GND.n4862 0.0208901
R7376 GND.n4866 GND.n4863 0.0208901
R7377 GND.n4876 GND.n4875 0.0208901
R7378 GND.n2828 GND.n2827 0.0208901
R7379 GND.n2831 GND.n2828 0.0208901
R7380 GND.n2841 GND.n2840 0.0208901
R7381 GND.n5795 GND.n5793 0.0205658
R7382 GND.n1374 GND.n1370 0.0202922
R7383 GND.n4900 GND.n4898 0.0200011
R7384 GND.n4699 GND.n4697 0.0200011
R7385 GND.n3155 GND.n3152 0.0200011
R7386 GND.n2823 GND.n2821 0.0200011
R7387 GND.n2284 GND.n2282 0.0200011
R7388 GND.n7688 GND.n7686 0.0200011
R7389 GND.n1544 GND.n1542 0.0200011
R7390 GND.n5381 GND.n5379 0.0200011
R7391 GND.n3950 GND.n3948 0.0200011
R7392 GND.n5242 GND.n5240 0.0200011
R7393 GND.n3842 GND.n3840 0.0200011
R7394 GND.n3519 GND.n3517 0.0200011
R7395 GND.n1971 GND.n1969 0.0200011
R7396 GND.n2058 GND.n2056 0.0200011
R7397 GND.n2446 GND.n2444 0.0200011
R7398 GND.n2755 GND.n2753 0.0200011
R7399 GND.n3410 GND.n3409 0.0198933
R7400 GND.n3324 GND 0.0198182
R7401 GND.n7511 GND 0.0198182
R7402 GND.n7573 GND 0.0198182
R7403 GND.n2627 GND 0.0198182
R7404 GND.n3053 GND 0.0198182
R7405 GND.n6978 GND 0.0198182
R7406 GND.n6824 GND 0.0198182
R7407 GND.n7760 GND 0.0198182
R7408 GND.n5640 GND 0.0198182
R7409 GND.n5456 GND 0.0198182
R7410 GND.n7449 GND 0.0198182
R7411 GND.n5114 GND 0.0198182
R7412 GND.n3714 GND 0.0198182
R7413 GND.n5513 GND 0.0198182
R7414 GND.n6502 GND 0.0198182
R7415 GND.n7080 GND 0.0198182
R7416 GND.n1370 GND.n1369 0.0197936
R7417 GND.n2030 GND.n2029 0.0197605
R7418 GND.n4667 GND.n4662 0.0195603
R7419 GND.n3214 GND.n3213 0.0195603
R7420 GND.n2261 GND.n2260 0.0195603
R7421 GND.n7664 GND.n163 0.0195603
R7422 GND.n1521 GND.n1520 0.0195603
R7423 GND.n5358 GND.n5357 0.0195603
R7424 GND.n3927 GND.n3926 0.0195603
R7425 GND.n5219 GND.n5218 0.0195603
R7426 GND.n3819 GND.n3818 0.0195603
R7427 GND.n3496 GND.n3495 0.0195603
R7428 GND.n1948 GND.n1947 0.0195603
R7429 GND.n2048 GND.n2044 0.0195603
R7430 GND.n2423 GND.n2422 0.0195603
R7431 GND.n2732 GND.n2731 0.0195603
R7432 GND.n4877 GND.n4876 0.0195603
R7433 GND.n2842 GND.n2841 0.0195603
R7434 GND.n3328 GND.n3327 0.0186818
R7435 GND.n7515 GND.n7514 0.0186818
R7436 GND.n7577 GND.n7576 0.0186818
R7437 GND.n2631 GND.n2630 0.0186818
R7438 GND.n3057 GND.n3056 0.0186818
R7439 GND.n6977 GND.n6975 0.0186818
R7440 GND.n6823 GND.n6821 0.0186818
R7441 GND.n7759 GND.n7755 0.0186818
R7442 GND.n5639 GND.n5637 0.0186818
R7443 GND.n5455 GND.n5453 0.0186818
R7444 GND.n7453 GND.n7452 0.0186818
R7445 GND.n5118 GND.n5117 0.0186818
R7446 GND.n3718 GND.n3717 0.0186818
R7447 GND.n5512 GND.n5510 0.0186818
R7448 GND.n6506 GND.n6505 0.0186818
R7449 GND.n7084 GND.n7083 0.0186818
R7450 GND.n5753 GND.n5749 0.0185921
R7451 GND.n44 GND 0.0182083
R7452 GND.n6371 GND 0.0182083
R7453 GND.n4474 GND.n4473 0.0179743
R7454 GND GND.n6212 0.0178611
R7455 GND.n4724 GND.n4723 0.0176904
R7456 GND.n3192 GND.n3191 0.0176904
R7457 GND.n2878 GND.n2877 0.0176904
R7458 GND.n2322 GND.n2321 0.0176904
R7459 GND.n7725 GND.n7724 0.0176904
R7460 GND.n1581 GND.n1580 0.0176904
R7461 GND.n5421 GND.n5420 0.0176904
R7462 GND.n3988 GND.n3987 0.0176904
R7463 GND.n5286 GND.n5285 0.0176904
R7464 GND.n3876 GND.n3875 0.0176904
R7465 GND.n3549 GND.n3548 0.0176904
R7466 GND.n2008 GND.n2007 0.0176904
R7467 GND.n2097 GND.n2096 0.0176904
R7468 GND.n2476 GND.n2475 0.0176904
R7469 GND.n4933 GND.n4932 0.0176904
R7470 GND.n5334 GND.n1445 0.0175762
R7471 GND.n6194 GND.n6193 0.0172763
R7472 GND.n2770 GND.n2769 0.0172687
R7473 GND GND.n35 0.0171667
R7474 GND.n3243 GND.n3241 0.0171667
R7475 GND.n7546 GND.n7544 0.0171667
R7476 GND.n7608 GND.n7606 0.0171667
R7477 GND.n2507 GND.n2505 0.0171667
R7478 GND.n2924 GND.n2922 0.0171667
R7479 GND.n6946 GND.n6944 0.0171667
R7480 GND.n6783 GND.n6781 0.0171667
R7481 GND.n72 GND.n70 0.0171667
R7482 GND.n1016 GND.n1014 0.0171667
R7483 GND.n1245 GND.n1243 0.0171667
R7484 GND.n7484 GND.n7482 0.0171667
R7485 GND.n4983 GND.n4981 0.0171667
R7486 GND.n3589 GND.n3587 0.0171667
R7487 GND.n1115 GND.n1113 0.0171667
R7488 GND.n6537 GND.n6535 0.0171667
R7489 GND.n7115 GND.n7113 0.0171667
R7490 GND GND.n6362 0.0171667
R7491 GND.n5743 GND.n5741 0.0171667
R7492 GND.n5741 GND.n5737 0.0171667
R7493 GND.n5737 GND.n5656 0.0171667
R7494 GND.n6145 GND.n6141 0.0171667
R7495 GND.n6147 GND.n6145 0.0171667
R7496 GND.n4577 GND.n4576 0.0167601
R7497 GND.n2710 GND.n2709 0.0166817
R7498 GND.n3136 GND.n3135 0.0166817
R7499 GND.n4059 GND.n4058 0.0166817
R7500 GND.n6164 GND.n6161 0.0166184
R7501 GND.n3340 GND.n3339 0.0164091
R7502 GND.n7527 GND.n7526 0.0164091
R7503 GND.n7589 GND.n7588 0.0164091
R7504 GND.n2643 GND.n2642 0.0164091
R7505 GND.n3069 GND.n3068 0.0164091
R7506 GND.n6935 GND.n6934 0.0164091
R7507 GND.n6812 GND.n6811 0.0164091
R7508 GND.n60 GND.n59 0.0164091
R7509 GND.n1005 GND.n1004 0.0164091
R7510 GND.n1234 GND.n1233 0.0164091
R7511 GND.n7465 GND.n7464 0.0164091
R7512 GND.n5130 GND.n5129 0.0164091
R7513 GND.n3730 GND.n3729 0.0164091
R7514 GND.n5501 GND.n5500 0.0164091
R7515 GND.n6522 GND.n6521 0.0164091
R7516 GND.n7096 GND.n7095 0.0164091
R7517 GND.n4101 GND.n4099 0.016125
R7518 GND.n5763 GND.n5759 0.0159605
R7519 GND.n5832 GND 0.0158101
R7520 GND.n5332 GND.n5331 0.0157734
R7521 GND.n6148 GND.n6147 0.0157174
R7522 GND.n1498 GND.n1497 0.0157059
R7523 GND.n1329 GND.n1278 0.0157059
R7524 GND.n5196 GND.n5195 0.0157059
R7525 GND.n3472 GND.n3421 0.0157059
R7526 GND.n2399 GND.n2348 0.0157059
R7527 GND.n6152 GND 0.0156316
R7528 GND.n5825 GND 0.0156316
R7529 GND GND.n5779 0.0156316
R7530 GND.n5721 GND 0.0156316
R7531 GND.n5759 GND.n5694 0.0153026
R7532 GND.n4855 GND.n4853 0.0152059
R7533 GND.n4648 GND.n4646 0.0152059
R7534 GND.n2710 GND.n2660 0.0152059
R7535 GND.n3394 GND.n3393 0.0152059
R7536 GND.n2239 GND.n2237 0.0152059
R7537 GND.n2177 GND.n2175 0.0152059
R7538 GND.n149 GND.n147 0.0152059
R7539 GND.n1499 GND.n1446 0.0152059
R7540 GND.n1331 GND.n1330 0.0152059
R7541 GND.n5197 GND.n5144 0.0152059
R7542 GND.n3797 GND.n3795 0.0152059
R7543 GND.n3474 GND.n3473 0.0152059
R7544 GND.n1926 GND.n1924 0.0152059
R7545 GND.n2401 GND.n2400 0.0152059
R7546 GND.n3184 GND.n3183 0.015169
R7547 GND.n3183 GND.n3182 0.015169
R7548 GND.n3221 GND.n3220 0.015169
R7549 GND.n3220 GND.n3219 0.015169
R7550 GND.n3178 GND.n3177 0.015169
R7551 GND.n3177 GND.t284 0.015169
R7552 GND.n3176 GND.n3175 0.015169
R7553 GND.t284 GND.n3176 0.015169
R7554 GND.n3174 GND.n3173 0.015169
R7555 GND.t284 GND.n3174 0.015169
R7556 GND.n2913 GND.n2912 0.015169
R7557 GND.n2912 GND.t22 0.015169
R7558 GND.n2911 GND.n2910 0.015169
R7559 GND.t22 GND.n2911 0.015169
R7560 GND.n2909 GND.n2908 0.015169
R7561 GND.t22 GND.n2909 0.015169
R7562 GND.n3188 GND.n3187 0.015169
R7563 GND.n2849 GND.n2848 0.015169
R7564 GND.n2852 GND.n2849 0.015169
R7565 GND.n2851 GND.n2850 0.015169
R7566 GND.n2852 GND.n2851 0.015169
R7567 GND.n2866 GND.n2865 0.015169
R7568 GND.n2865 GND.n2864 0.015169
R7569 GND.n2307 GND.n2306 0.015169
R7570 GND.n2306 GND.t315 0.015169
R7571 GND.n2305 GND.n2304 0.015169
R7572 GND.t315 GND.n2305 0.015169
R7573 GND.n2303 GND.n2302 0.015169
R7574 GND.t315 GND.n2303 0.015169
R7575 GND.n7711 GND.n7710 0.015169
R7576 GND.n7710 GND.t287 0.015169
R7577 GND.n7709 GND.n7708 0.015169
R7578 GND.t287 GND.n7709 0.015169
R7579 GND.n7707 GND.n7706 0.015169
R7580 GND.t287 GND.n7707 0.015169
R7581 GND.n1567 GND.n1566 0.015169
R7582 GND.n1566 GND.t1094 0.015169
R7583 GND.n1565 GND.n1564 0.015169
R7584 GND.t1094 GND.n1565 0.015169
R7585 GND.n1563 GND.n1562 0.015169
R7586 GND.t1094 GND.n1563 0.015169
R7587 GND.n5404 GND.n5403 0.015169
R7588 GND.n5403 GND.t286 0.015169
R7589 GND.n5402 GND.n5401 0.015169
R7590 GND.t286 GND.n5402 0.015169
R7591 GND.n5400 GND.n5399 0.015169
R7592 GND.t286 GND.n5400 0.015169
R7593 GND.n5265 GND.n5264 0.015169
R7594 GND.n5264 GND.t446 0.015169
R7595 GND.n5263 GND.n5262 0.015169
R7596 GND.t446 GND.n5263 0.015169
R7597 GND.n5261 GND.n5260 0.015169
R7598 GND.t446 GND.n5261 0.015169
R7599 GND.n5282 GND.n5281 0.015169
R7600 GND.n5281 GND.n5280 0.015169
R7601 GND.n3934 GND.n3933 0.015169
R7602 GND.n3937 GND.n3934 0.015169
R7603 GND.n3936 GND.n3935 0.015169
R7604 GND.n3937 GND.n3936 0.015169
R7605 GND.n5279 GND.n5278 0.015169
R7606 GND.n5280 GND.n5279 0.015169
R7607 GND.n5228 GND.n5227 0.015169
R7608 GND.n5229 GND.n5228 0.015169
R7609 GND.n5274 GND.n5273 0.015169
R7610 GND.n5273 GND.n5272 0.015169
R7611 GND.n5226 GND.n5225 0.015169
R7612 GND.n5229 GND.n5226 0.015169
R7613 GND.n5271 GND.n5270 0.015169
R7614 GND.n5272 GND.n5271 0.015169
R7615 GND.n3865 GND.n3864 0.015169
R7616 GND.n3864 GND.t317 0.015169
R7617 GND.n3863 GND.n3862 0.015169
R7618 GND.t317 GND.n3863 0.015169
R7619 GND.n3861 GND.n3860 0.015169
R7620 GND.t317 GND.n3861 0.015169
R7621 GND.n5417 GND.n5416 0.015169
R7622 GND.n3826 GND.n3825 0.015169
R7623 GND.n3829 GND.n3826 0.015169
R7624 GND.n3828 GND.n3827 0.015169
R7625 GND.n3829 GND.n3828 0.015169
R7626 GND.n3871 GND.n3870 0.015169
R7627 GND.n3870 GND.n3869 0.015169
R7628 GND.n5367 GND.n5366 0.015169
R7629 GND.n5368 GND.n5367 0.015169
R7630 GND.n5413 GND.n5412 0.015169
R7631 GND.n5412 GND.n5411 0.015169
R7632 GND.n5365 GND.n5364 0.015169
R7633 GND.n5368 GND.n5365 0.015169
R7634 GND.n5410 GND.n5409 0.015169
R7635 GND.n5411 GND.n5410 0.015169
R7636 GND.n3542 GND.n3541 0.015169
R7637 GND.n3541 GND.t281 0.015169
R7638 GND.n3540 GND.n3539 0.015169
R7639 GND.t281 GND.n3540 0.015169
R7640 GND.n3538 GND.n3537 0.015169
R7641 GND.t281 GND.n3538 0.015169
R7642 GND.n1577 GND.n1576 0.015169
R7643 GND.n1576 GND.n1575 0.015169
R7644 GND.n3503 GND.n3502 0.015169
R7645 GND.n3506 GND.n3503 0.015169
R7646 GND.n3505 GND.n3504 0.015169
R7647 GND.n3506 GND.n3505 0.015169
R7648 GND.n1574 GND.n1573 0.015169
R7649 GND.n1575 GND.n1574 0.015169
R7650 GND.n1530 GND.n1529 0.015169
R7651 GND.n1531 GND.n1530 0.015169
R7652 GND.n2001 GND.n2000 0.015169
R7653 GND.n2002 GND.n2001 0.015169
R7654 GND.n1528 GND.n1527 0.015169
R7655 GND.n1531 GND.n1528 0.015169
R7656 GND.n2004 GND.n2003 0.015169
R7657 GND.n2003 GND.n2002 0.015169
R7658 GND.n1994 GND.n1993 0.015169
R7659 GND.n1993 GND.t1107 0.015169
R7660 GND.n1992 GND.n1991 0.015169
R7661 GND.t1107 GND.n1992 0.015169
R7662 GND.n1990 GND.n1989 0.015169
R7663 GND.t1107 GND.n1990 0.015169
R7664 GND.n7721 GND.n7720 0.015169
R7665 GND.n7720 GND.n7719 0.015169
R7666 GND.n1955 GND.n1954 0.015169
R7667 GND.n1958 GND.n1955 0.015169
R7668 GND.n1957 GND.n1956 0.015169
R7669 GND.n1958 GND.n1957 0.015169
R7670 GND.n7718 GND.n7717 0.015169
R7671 GND.n7719 GND.n7718 0.015169
R7672 GND.n7672 GND.n7671 0.015169
R7673 GND.n7675 GND.n7672 0.015169
R7674 GND.n118 GND.n117 0.015169
R7675 GND.n119 GND.n118 0.015169
R7676 GND.n7674 GND.n7673 0.015169
R7677 GND.n7675 GND.n7674 0.015169
R7678 GND.n121 GND.n120 0.015169
R7679 GND.n120 GND.n119 0.015169
R7680 GND.n1661 GND.n1660 0.015169
R7681 GND.n1660 GND.t1559 0.015169
R7682 GND.n2114 GND.n2113 0.015169
R7683 GND.n2115 GND.n2114 0.015169
R7684 GND.n1653 GND.n1652 0.015169
R7685 GND.n1652 GND.t493 0.015169
R7686 GND.n2091 GND.n2090 0.015169
R7687 GND.n2064 GND.n2063 0.015169
R7688 GND.n2067 GND.n2064 0.015169
R7689 GND.n2066 GND.n2065 0.015169
R7690 GND.n2067 GND.n2066 0.015169
R7691 GND.n2093 GND.n2092 0.015169
R7692 GND.n2092 GND.n2091 0.015169
R7693 GND.n2270 GND.n2269 0.015169
R7694 GND.n2271 GND.n2270 0.015169
R7695 GND.n2316 GND.n2315 0.015169
R7696 GND.n2315 GND.n2314 0.015169
R7697 GND.n2268 GND.n2267 0.015169
R7698 GND.n2271 GND.n2268 0.015169
R7699 GND.n2313 GND.n2312 0.015169
R7700 GND.n2314 GND.n2313 0.015169
R7701 GND.n2469 GND.n2468 0.015169
R7702 GND.n2468 GND.t242 0.015169
R7703 GND.n2467 GND.n2466 0.015169
R7704 GND.t242 GND.n2467 0.015169
R7705 GND.n2465 GND.n2464 0.015169
R7706 GND.t242 GND.n2465 0.015169
R7707 GND.n2432 GND.n2431 0.015169
R7708 GND.n2433 GND.n2432 0.015169
R7709 GND.n2762 GND.n2761 0.015169
R7710 GND.n2763 GND.n2762 0.015169
R7711 GND.n2874 GND.n2873 0.015169
R7712 GND.n2873 GND.n2872 0.015169
R7713 GND.n2739 GND.n2738 0.015169
R7714 GND.n2742 GND.n2739 0.015169
R7715 GND.n2871 GND.n2870 0.015169
R7716 GND.n2872 GND.n2871 0.015169
R7717 GND.n2430 GND.n2429 0.015169
R7718 GND.n2433 GND.n2430 0.015169
R7719 GND.n2741 GND.n2740 0.015169
R7720 GND.n2742 GND.n2741 0.015169
R7721 GND.n2793 GND.n2792 0.015169
R7722 GND.n2792 GND.t471 0.015169
R7723 GND.n2791 GND.n2790 0.015169
R7724 GND.t471 GND.n2791 0.015169
R7725 GND.n2765 GND.n2764 0.015169
R7726 GND.n2764 GND.n2763 0.015169
R7727 GND.n2789 GND.n2788 0.015169
R7728 GND.t471 GND.n2789 0.015169
R7729 GND.n4923 GND.n4922 0.015169
R7730 GND.n4922 GND.t282 0.015169
R7731 GND.n4921 GND.n4920 0.015169
R7732 GND.t282 GND.n4921 0.015169
R7733 GND.n4919 GND.n4918 0.015169
R7734 GND.t282 GND.n4919 0.015169
R7735 GND.n3983 GND.n3982 0.015169
R7736 GND.n3982 GND.n3980 0.015169
R7737 GND.n4884 GND.n4883 0.015169
R7738 GND.n4887 GND.n4884 0.015169
R7739 GND.n4886 GND.n4885 0.015169
R7740 GND.n4887 GND.n4886 0.015169
R7741 GND.n3979 GND.n3977 0.015169
R7742 GND.n3980 GND.n3979 0.015169
R7743 GND.n3962 GND.n3961 0.015169
R7744 GND.n3961 GND.t491 0.015169
R7745 GND.n3960 GND.n3959 0.015169
R7746 GND.t491 GND.n3960 0.015169
R7747 GND.n3958 GND.n3957 0.015169
R7748 GND.t491 GND.n3958 0.015169
R7749 GND.n4118 GND.n4117 0.015169
R7750 GND.n4119 GND.n4118 0.015169
R7751 GND.n4133 GND.n4132 0.015169
R7752 GND.n4134 GND.n4133 0.015169
R7753 GND.n4148 GND.n4147 0.015169
R7754 GND.n4149 GND.n4148 0.015169
R7755 GND.n4163 GND.n4162 0.015169
R7756 GND.n4164 GND.n4163 0.015169
R7757 GND.n4182 GND.n4181 0.015169
R7758 GND.n4183 GND.n4182 0.015169
R7759 GND.n4197 GND.n4196 0.015169
R7760 GND.n4198 GND.n4197 0.015169
R7761 GND.n4212 GND.n4211 0.015169
R7762 GND.n4213 GND.n4212 0.015169
R7763 GND.n4227 GND.n4226 0.015169
R7764 GND.n4228 GND.n4227 0.015169
R7765 GND.n4245 GND.n4244 0.015169
R7766 GND.n4246 GND.n4245 0.015169
R7767 GND.n4269 GND.n4268 0.015169
R7768 GND.n4270 GND.n4269 0.015169
R7769 GND.n4289 GND.n4288 0.015169
R7770 GND.n4290 GND.n4289 0.015169
R7771 GND.n4306 GND.n4305 0.015169
R7772 GND.n4307 GND.n4306 0.015169
R7773 GND.n4321 GND.n4320 0.015169
R7774 GND.n4322 GND.n4321 0.015169
R7775 GND.n4336 GND.n4335 0.015169
R7776 GND.n4337 GND.n4336 0.015169
R7777 GND.n4351 GND.n4350 0.015169
R7778 GND.n4352 GND.n4351 0.015169
R7779 GND.n4368 GND.n4367 0.015169
R7780 GND.n4369 GND.n4368 0.015169
R7781 GND.n4383 GND.n4382 0.015169
R7782 GND.n4384 GND.n4383 0.015169
R7783 GND.n4398 GND.n4397 0.015169
R7784 GND.n4399 GND.n4398 0.015169
R7785 GND.n4413 GND.n4412 0.015169
R7786 GND.n4414 GND.n4413 0.015169
R7787 GND.n4078 GND.n4077 0.015169
R7788 GND.n4429 GND.n4428 0.015169
R7789 GND.n4430 GND.n4429 0.015169
R7790 GND.n4067 GND.n4066 0.015169
R7791 GND.n4068 GND.n4067 0.015169
R7792 GND.n4745 GND.n4744 0.015169
R7793 GND.t1091 GND.n4745 0.015169
R7794 GND.n4746 GND.t1091 0.015169
R7795 GND.n4747 GND.n4746 0.015169
R7796 GND.n4743 GND.n4742 0.015169
R7797 GND.t1091 GND.n4743 0.015169
R7798 GND.n4720 GND.n4719 0.015169
R7799 GND.n4929 GND.n4928 0.015169
R7800 GND.n4928 GND.n4927 0.015169
R7801 GND.n4682 GND.n4681 0.015169
R7802 GND.n4685 GND.n4682 0.015169
R7803 GND.n4684 GND.n4683 0.015169
R7804 GND.n4685 GND.n4684 0.015169
R7805 GND.n4709 GND.n4708 0.015169
R7806 GND.n4708 GND.n4707 0.015169
R7807 GND.n4672 GND.n4671 0.015169
R7808 GND.n4673 GND.n4672 0.015169
R7809 GND.n4959 GND.n4958 0.014943
R7810 GND.n1844 GND.n1841 0.014943
R7811 GND.n1839 GND.n1836 0.014943
R7812 GND.n1834 GND.n1831 0.014943
R7813 GND.n1829 GND.n1826 0.014943
R7814 GND.n1824 GND.n1821 0.014943
R7815 GND.n1819 GND.n1816 0.014943
R7816 GND.n1814 GND.n1811 0.014943
R7817 GND.n1809 GND.n1806 0.014943
R7818 GND.n1804 GND.n1801 0.014943
R7819 GND.n1799 GND.n1796 0.014943
R7820 GND.n1794 GND.n1791 0.014943
R7821 GND.n1789 GND.n1786 0.014943
R7822 GND.n1784 GND.n1781 0.014943
R7823 GND.n1779 GND.n1778 0.014943
R7824 GND.n4800 GND.n4799 0.014943
R7825 GND.n6168 GND.n6164 0.0146447
R7826 GND.n5668 GND.n5666 0.0146077
R7827 GND.n1841 GND.n1840 0.0144432
R7828 GND.n1836 GND.n1835 0.0144432
R7829 GND.n1831 GND.n1830 0.0144432
R7830 GND.n1826 GND.n1825 0.0144432
R7831 GND.n1821 GND.n1820 0.0144432
R7832 GND.n1816 GND.n1815 0.0144432
R7833 GND.n1811 GND.n1810 0.0144432
R7834 GND.n1806 GND.n1805 0.0144432
R7835 GND.n1801 GND.n1800 0.0144432
R7836 GND.n1796 GND.n1795 0.0144432
R7837 GND.n1791 GND.n1790 0.0144432
R7838 GND.n1786 GND.n1785 0.0144432
R7839 GND.n1781 GND.n1780 0.0144432
R7840 GND.n1778 GND.n1777 0.0144432
R7841 GND.n4799 GND.n4798 0.0144432
R7842 GND.n4958 GND.n4957 0.0144432
R7843 GND.n4573 GND.n4482 0.0143889
R7844 GND.n3255 GND.n3254 0.0140417
R7845 GND.n7558 GND.n7557 0.0140417
R7846 GND.n7620 GND.n7619 0.0140417
R7847 GND.n2516 GND.n2515 0.0140417
R7848 GND.n2933 GND.n2932 0.0140417
R7849 GND.n6958 GND.n6957 0.0140417
R7850 GND.n6795 GND.n6794 0.0140417
R7851 GND.n84 GND.n83 0.0140417
R7852 GND.n1028 GND.n1027 0.0140417
R7853 GND.n1254 GND.n1253 0.0140417
R7854 GND.n7496 GND.n7495 0.0140417
R7855 GND.n4995 GND.n4994 0.0140417
R7856 GND.n3598 GND.n3597 0.0140417
R7857 GND.n1127 GND.n1126 0.0140417
R7858 GND.n6549 GND.n6548 0.0140417
R7859 GND.n7127 GND.n7126 0.0140417
R7860 GND.n6198 GND.n6194 0.0139868
R7861 GND.n4659 GND.n4658 0.0138596
R7862 GND.n3210 GND.n3209 0.0138596
R7863 GND.n2257 GND.n2256 0.0138596
R7864 GND.n160 GND.n159 0.0138596
R7865 GND.n1517 GND.n1516 0.0138596
R7866 GND.n5354 GND.n5353 0.0138596
R7867 GND.n3923 GND.n3922 0.0138596
R7868 GND.n5215 GND.n5214 0.0138596
R7869 GND.n3815 GND.n3814 0.0138596
R7870 GND.n3492 GND.n3491 0.0138596
R7871 GND.n1944 GND.n1943 0.0138596
R7872 GND.n2041 GND.n2040 0.0138596
R7873 GND.n2419 GND.n2418 0.0138596
R7874 GND.n2728 GND.n2727 0.0138596
R7875 GND.n4873 GND.n4872 0.0138596
R7876 GND.n2838 GND.n2837 0.0138596
R7877 GND.n723 GND.n719 0.012734
R7878 GND.n741 GND.n739 0.012734
R7879 GND.n745 GND.n741 0.012734
R7880 GND.n747 GND.n745 0.012734
R7881 GND.n751 GND.n747 0.012734
R7882 GND.n753 GND.n751 0.012734
R7883 GND.n757 GND.n753 0.012734
R7884 GND.n759 GND.n757 0.012734
R7885 GND.n760 GND.n759 0.012734
R7886 GND.n765 GND.n763 0.012734
R7887 GND.n769 GND.n765 0.012734
R7888 GND.n815 GND.n813 0.012734
R7889 GND.n813 GND.n809 0.012734
R7890 GND.n809 GND.n805 0.012734
R7891 GND.n805 GND.n803 0.012734
R7892 GND.n803 GND.n799 0.012734
R7893 GND.n799 GND.n797 0.012734
R7894 GND.n797 GND.n793 0.012734
R7895 GND.n793 GND.n791 0.012734
R7896 GND.n791 GND.n787 0.012734
R7897 GND.n787 GND.n785 0.012734
R7898 GND.n784 GND.n783 0.012734
R7899 GND.n783 GND.n781 0.012734
R7900 GND.n781 GND.n777 0.012734
R7901 GND.n837 GND.n833 0.012734
R7902 GND.n839 GND.n837 0.012734
R7903 GND.n843 GND.n839 0.012734
R7904 GND.n845 GND.n843 0.012734
R7905 GND.n849 GND.n845 0.012734
R7906 GND.n851 GND.n849 0.012734
R7907 GND.n855 GND.n851 0.012734
R7908 GND.n859 GND.n858 0.012734
R7909 GND.n864 GND.n862 0.012734
R7910 GND.n868 GND.n864 0.012734
R7911 GND.n908 GND.n906 0.012734
R7912 GND.n906 GND.n902 0.012734
R7913 GND.n902 GND.n898 0.012734
R7914 GND.n898 GND.n896 0.012734
R7915 GND.n896 GND.n892 0.012734
R7916 GND.n892 GND.n890 0.012734
R7917 GND.n890 GND.n886 0.012734
R7918 GND.n886 GND.n884 0.012734
R7919 GND.n884 GND.n880 0.012734
R7920 GND.n880 GND.n878 0.012734
R7921 GND.n877 GND.n876 0.012734
R7922 GND.n928 GND.n926 0.012734
R7923 GND.n932 GND.n928 0.012734
R7924 GND.n936 GND.n932 0.012734
R7925 GND.n938 GND.n936 0.012734
R7926 GND.n942 GND.n938 0.012734
R7927 GND.n944 GND.n942 0.012734
R7928 GND.n948 GND.n944 0.012734
R7929 GND.n950 GND.n948 0.012734
R7930 GND.n954 GND.n950 0.012734
R7931 GND.n956 GND.n954 0.012734
R7932 GND.n957 GND.n956 0.012734
R7933 GND.n962 GND.n960 0.012734
R7934 GND.n965 GND.n962 0.012734
R7935 GND.n967 GND.n965 0.012734
R7936 GND.n987 GND.n985 0.012734
R7937 GND.n982 GND.n981 0.012734
R7938 GND.n981 GND.n979 0.012734
R7939 GND.n979 GND.n975 0.012734
R7940 GND.n975 GND.n973 0.012734
R7941 GND.n5870 GND.n5866 0.012734
R7942 GND.n5872 GND.n5870 0.012734
R7943 GND.n5907 GND.n5903 0.012734
R7944 GND.n5903 GND.n5901 0.012734
R7945 GND.n5901 GND.n5897 0.012734
R7946 GND.n5897 GND.n5895 0.012734
R7947 GND.n5895 GND.n5891 0.012734
R7948 GND.n5891 GND.n5889 0.012734
R7949 GND.n5889 GND.n5885 0.012734
R7950 GND.n5885 GND.n5883 0.012734
R7951 GND.n5882 GND.n5881 0.012734
R7952 GND.n5881 GND.n5879 0.012734
R7953 GND.n5929 GND.n5925 0.012734
R7954 GND.n5933 GND.n5929 0.012734
R7955 GND.n5935 GND.n5933 0.012734
R7956 GND.n5939 GND.n5935 0.012734
R7957 GND.n5941 GND.n5939 0.012734
R7958 GND.n5945 GND.n5941 0.012734
R7959 GND.n5947 GND.n5945 0.012734
R7960 GND.n5951 GND.n5947 0.012734
R7961 GND.n5953 GND.n5951 0.012734
R7962 GND.n5954 GND.n5953 0.012734
R7963 GND.n5959 GND.n5957 0.012734
R7964 GND.n5963 GND.n5959 0.012734
R7965 GND.n5965 GND.n5963 0.012734
R7966 GND.n5996 GND.n5992 0.012734
R7967 GND.n5992 GND.n5988 0.012734
R7968 GND.n5988 GND.n5986 0.012734
R7969 GND.n5986 GND.n5982 0.012734
R7970 GND.n5982 GND.n5980 0.012734
R7971 GND.n5980 GND.n5976 0.012734
R7972 GND.n5976 GND.n5974 0.012734
R7973 GND.n5974 GND.n5852 0.012734
R7974 GND.n6133 GND.n6132 0.012734
R7975 GND.n6132 GND.n6130 0.012734
R7976 GND.n6010 GND.n6006 0.012734
R7977 GND.n6014 GND.n6010 0.012734
R7978 GND.n6016 GND.n6014 0.012734
R7979 GND.n6020 GND.n6016 0.012734
R7980 GND.n6022 GND.n6020 0.012734
R7981 GND.n6026 GND.n6022 0.012734
R7982 GND.n6028 GND.n6026 0.012734
R7983 GND.n6032 GND.n6028 0.012734
R7984 GND.n6034 GND.n6032 0.012734
R7985 GND.n6035 GND.n6034 0.012734
R7986 GND.n6040 GND.n6038 0.012734
R7987 GND.n6044 GND.n6040 0.012734
R7988 GND.n6054 GND.n6052 0.012734
R7989 GND.n6058 GND.n6054 0.012734
R7990 GND.n6062 GND.n6058 0.012734
R7991 GND.n6064 GND.n6062 0.012734
R7992 GND.n6068 GND.n6064 0.012734
R7993 GND.n6070 GND.n6068 0.012734
R7994 GND.n6074 GND.n6070 0.012734
R7995 GND.n6076 GND.n6074 0.012734
R7996 GND.n6080 GND.n6076 0.012734
R7997 GND.n6082 GND.n6080 0.012734
R7998 GND.n6083 GND.n6082 0.012734
R7999 GND.n6088 GND.n6086 0.012734
R8000 GND.n6091 GND.n6088 0.012734
R8001 GND.n6093 GND.n6091 0.012734
R8002 GND.n6113 GND.n6111 0.012734
R8003 GND.n6108 GND.n6107 0.012734
R8004 GND.n6107 GND.n6105 0.012734
R8005 GND.n6105 GND.n6101 0.012734
R8006 GND.n6101 GND.n6099 0.012734
R8007 GND.n7241 GND.n7237 0.012734
R8008 GND.n7243 GND.n7241 0.012734
R8009 GND.n7278 GND.n7274 0.012734
R8010 GND.n7274 GND.n7272 0.012734
R8011 GND.n7272 GND.n7268 0.012734
R8012 GND.n7268 GND.n7266 0.012734
R8013 GND.n7266 GND.n7262 0.012734
R8014 GND.n7262 GND.n7260 0.012734
R8015 GND.n7260 GND.n7256 0.012734
R8016 GND.n7256 GND.n7254 0.012734
R8017 GND.n7253 GND.n7252 0.012734
R8018 GND.n7252 GND.n7250 0.012734
R8019 GND.n7300 GND.n7296 0.012734
R8020 GND.n7304 GND.n7300 0.012734
R8021 GND.n7306 GND.n7304 0.012734
R8022 GND.n7310 GND.n7306 0.012734
R8023 GND.n7312 GND.n7310 0.012734
R8024 GND.n7316 GND.n7312 0.012734
R8025 GND.n7318 GND.n7316 0.012734
R8026 GND.n7322 GND.n7318 0.012734
R8027 GND.n7324 GND.n7322 0.012734
R8028 GND.n7325 GND.n7324 0.012734
R8029 GND.n7330 GND.n7328 0.012734
R8030 GND.n7334 GND.n7330 0.012734
R8031 GND.n7336 GND.n7334 0.012734
R8032 GND.n7367 GND.n7363 0.012734
R8033 GND.n7363 GND.n7359 0.012734
R8034 GND.n7359 GND.n7357 0.012734
R8035 GND.n7357 GND.n7353 0.012734
R8036 GND.n7353 GND.n7351 0.012734
R8037 GND.n7351 GND.n7347 0.012734
R8038 GND.n7347 GND.n7345 0.012734
R8039 GND.n7345 GND.n544 0.012734
R8040 GND.n7432 GND.n7431 0.012734
R8041 GND.n7431 GND.n7429 0.012734
R8042 GND.n7416 GND.n7414 0.012734
R8043 GND.n7414 GND.n7410 0.012734
R8044 GND.n7410 GND.n7406 0.012734
R8045 GND.n7406 GND.n7404 0.012734
R8046 GND.n7404 GND.n7400 0.012734
R8047 GND.n7400 GND.n7398 0.012734
R8048 GND.n7398 GND.n7394 0.012734
R8049 GND.n7394 GND.n7392 0.012734
R8050 GND.n7392 GND.n7388 0.012734
R8051 GND.n7388 GND.n7386 0.012734
R8052 GND.n7385 GND.n7384 0.012734
R8053 GND.n7384 GND.n7382 0.012734
R8054 GND.n594 GND.n590 0.012734
R8055 GND.n590 GND.n588 0.012734
R8056 GND.n588 GND.n584 0.012734
R8057 GND.n584 GND.n580 0.012734
R8058 GND.n580 GND.n578 0.012734
R8059 GND.n578 GND.n574 0.012734
R8060 GND.n574 GND.n572 0.012734
R8061 GND.n572 GND.n568 0.012734
R8062 GND.n568 GND.n566 0.012734
R8063 GND.n566 GND.n562 0.012734
R8064 GND.n562 GND.n560 0.012734
R8065 GND.n559 GND.n558 0.012734
R8066 GND.n558 GND.n556 0.012734
R8067 GND.n556 GND.n553 0.012734
R8068 GND.n7814 GND.n7813 0.012734
R8069 GND.n7819 GND.n7817 0.012734
R8070 GND.n7823 GND.n7819 0.012734
R8071 GND.n7825 GND.n7823 0.012734
R8072 GND.n7827 GND.n7825 0.012734
R8073 GND.n5749 GND.n5748 0.0126711
R8074 GND.n724 GND.n723 0.0126011
R8075 GND.n6135 GND.n6134 0.0126011
R8076 GND.n7434 GND.n7433 0.0126011
R8077 GND.n687 GND 0.0123421
R8078 GND.n6251 GND 0.0123421
R8079 GND.n856 GND.n855 0.0123351
R8080 GND.n876 GND.n874 0.0123351
R8081 GND.n6213 GND 0.0123056
R8082 GND GND.n6204 0.0123056
R8083 GND.n6205 GND 0.0123056
R8084 GND GND.n23 0.0123056
R8085 GND GND.n7791 0.0123056
R8086 GND GND.n665 0.0123056
R8087 GND GND.n6348 0.0123056
R8088 GND GND.n6324 0.0123056
R8089 GND GND.n6293 0.0123056
R8090 GND.n4898 GND.n4897 0.0120741
R8091 GND.n4697 GND.n4696 0.0120741
R8092 GND.n3152 GND.n3151 0.0120741
R8093 GND.n2821 GND.n2820 0.0120741
R8094 GND.n2282 GND.n2281 0.0120741
R8095 GND.n7686 GND.n7685 0.0120741
R8096 GND.n1542 GND.n1541 0.0120741
R8097 GND.n5379 GND.n5378 0.0120741
R8098 GND.n3948 GND.n3947 0.0120741
R8099 GND.n5240 GND.n5239 0.0120741
R8100 GND.n3840 GND.n3839 0.0120741
R8101 GND.n3517 GND.n3516 0.0120741
R8102 GND.n1969 GND.n1968 0.0120741
R8103 GND.n2056 GND.n2055 0.0120741
R8104 GND.n2444 GND.n2443 0.0120741
R8105 GND.n2753 GND.n2752 0.0120741
R8106 GND.n5879 GND.n5875 0.0120691
R8107 GND.n7250 GND.n7246 0.0120691
R8108 GND.n6141 GND.n6139 0.0117319
R8109 GND GND.n7778 0.0116111
R8110 GND.n646 GND 0.0116111
R8111 GND GND.n6311 0.0116111
R8112 GND.n6274 GND 0.0116111
R8113 GND.n770 GND.n769 0.0115372
R8114 GND.n320 GND.n318 0.0112143
R8115 GND.n218 GND.n216 0.0112143
R8116 GND.n2618 GND.n2545 0.0112143
R8117 GND.n3044 GND.n2969 0.0112143
R8118 GND.n7066 GND.n7064 0.0112143
R8119 GND.n6912 GND.n6910 0.0112143
R8120 GND.n6758 GND.n6756 0.0112143
R8121 GND.n5620 GND.n5619 0.0112143
R8122 GND.n1273 GND.n1272 0.0112143
R8123 GND.n497 GND.n422 0.0112143
R8124 GND.n5105 GND.n5027 0.0112143
R8125 GND.n3705 GND.n3633 0.0112143
R8126 GND.n5485 GND.n5484 0.0112143
R8127 GND.n6558 GND.n6556 0.0112143
R8128 GND.n7222 GND.n7150 0.0112143
R8129 GND.n3316 GND.n3277 0.0112143
R8130 GND.n4897 GND 0.0111481
R8131 GND.n4696 GND 0.0111481
R8132 GND.n3151 GND 0.0111481
R8133 GND.n2820 GND 0.0111481
R8134 GND.n2281 GND 0.0111481
R8135 GND.n7685 GND 0.0111481
R8136 GND.n1541 GND 0.0111481
R8137 GND.n5378 GND 0.0111481
R8138 GND.n3947 GND 0.0111481
R8139 GND.n5239 GND 0.0111481
R8140 GND.n3839 GND 0.0111481
R8141 GND.n3516 GND 0.0111481
R8142 GND.n1968 GND 0.0111481
R8143 GND.n2055 GND 0.0111481
R8144 GND.n2443 GND 0.0111481
R8145 GND.n2752 GND 0.0111481
R8146 GND GND.n703 0.0110263
R8147 GND GND.n6267 0.0110263
R8148 GND.n4108 GND.n4106 0.0109167
R8149 GND.n833 GND.n829 0.0107394
R8150 GND.n909 GND.n908 0.0107394
R8151 GND.n6094 GND.n6093 0.0107394
R8152 GND.n553 GND.n3 0.0107394
R8153 GND.n5913 GND.n5872 0.0107015
R8154 GND.n7284 GND.n7243 0.0107015
R8155 GND.n5793 GND.n5792 0.0106974
R8156 GND.n6045 GND.n6044 0.0104355
R8157 GND.n7382 GND.n7378 0.0104355
R8158 GND.n4180 GND.n4179 0.0102222
R8159 GND.n968 GND.n967 0.0102074
R8160 GND.n5997 GND.n5996 0.0102074
R8161 GND.n6006 GND.n6004 0.0102074
R8162 GND.n7368 GND.n7367 0.0102074
R8163 GND.n7417 GND.n7416 0.0102074
R8164 GND.n4490 GND.n4489 0.0101468
R8165 GND.n4491 GND.n4490 0.0101468
R8166 GND.n4549 GND.n4548 0.0101468
R8167 GND.n4550 GND.n4549 0.0101468
R8168 GND.n4544 GND.n4543 0.0101468
R8169 GND.n4550 GND.n4544 0.0101468
R8170 GND.n4540 GND.n4539 0.0101468
R8171 GND.n4550 GND.n4540 0.0101468
R8172 GND.n4536 GND.n4535 0.0101468
R8173 GND.n4550 GND.n4536 0.0101468
R8174 GND.n4488 GND.n4487 0.0101468
R8175 GND.n4491 GND.n4488 0.0101468
R8176 GND.n4531 GND.n4530 0.0101468
R8177 GND.n4550 GND.n4531 0.0101468
R8178 GND.n4526 GND.n4525 0.0101468
R8179 GND.n4550 GND.n4526 0.0101468
R8180 GND.n4522 GND.n4521 0.0101468
R8181 GND.n4550 GND.n4522 0.0101468
R8182 GND.n4518 GND.n4517 0.0101468
R8183 GND.n4550 GND.n4518 0.0101468
R8184 GND.n4515 GND.n4514 0.0101468
R8185 GND.n4550 GND.n4515 0.0101468
R8186 GND.n4486 GND.n4485 0.0101468
R8187 GND.n4491 GND.n4486 0.0101468
R8188 GND.n4509 GND.n4508 0.0101468
R8189 GND.n4550 GND.n4509 0.0101468
R8190 GND.n4504 GND.n4503 0.0101468
R8191 GND.n4550 GND.n4504 0.0101468
R8192 GND.n4484 GND.n4483 0.0101468
R8193 GND.n4491 GND.n4484 0.0101468
R8194 GND.n4499 GND.n4498 0.0101468
R8195 GND.n4550 GND.n4499 0.0101468
R8196 GND.n4494 GND.n4493 0.0101468
R8197 GND.n4550 GND.n4494 0.0101468
R8198 GND.n6227 GND.n6198 0.0100395
R8199 GND.n5665 GND.n5661 0.0100149
R8200 GND GND.n6492 0.009875
R8201 GND GND.n6402 0.009875
R8202 GND.n730 GND.n726 0.00967553
R8203 GND.n4108 GND.n4107 0.00959091
R8204 GND.n691 GND.n674 0.00950855
R8205 GND.n6255 GND.n6238 0.00950855
R8206 GND.n5675 GND.n5673 0.00941473
R8207 GND.n5679 GND.n5675 0.00941473
R8208 GND.n5683 GND.n5679 0.00941473
R8209 GND.n5685 GND.n5683 0.00941473
R8210 GND.n5849 GND.n5845 0.00941473
R8211 GND.n5845 GND.n5843 0.00941473
R8212 GND.n5843 GND.n5839 0.00941473
R8213 GND.n5839 GND.n5837 0.00941473
R8214 GND.n919 GND.n710 0.00940957
R8215 GND.n6169 GND.n6168 0.00938158
R8216 GND.n5918 GND.n5860 0.00914362
R8217 GND.n7289 GND.n7232 0.00914362
R8218 GND.n7779 GND.n7769 0.00906279
R8219 GND.n6312 GND.n6302 0.00906279
R8220 GND.n1385 GND.n1384 0.00904142
R8221 GND.n1421 GND.n1420 0.00898517
R8222 GND.n1339 GND.n1337 0.00898517
R8223 GND.n1356 GND.n1339 0.00898517
R8224 GND.n1403 GND.n1402 0.00898517
R8225 GND.n1388 GND.n1387 0.00898517
R8226 GND.n1387 GND.n1385 0.00898517
R8227 GND.n1337 GND.n1336 0.00897458
R8228 GND.n1421 GND.n1418 0.00896398
R8229 GND.n1358 GND.n1356 0.00896398
R8230 GND.n1361 GND.n1358 0.00896398
R8231 GND.n1363 GND.n1361 0.00896398
R8232 GND.n1364 GND.n1363 0.00896398
R8233 GND.n1435 GND.n1433 0.00896398
R8234 GND.n1395 GND.n1393 0.00896398
R8235 GND.n1396 GND.n1395 0.00896398
R8236 GND.n1388 GND.n1382 0.00896398
R8237 GND.n1403 GND.n1400 0.0089428
R8238 GND.n988 GND.n987 0.00887766
R8239 GND.n5966 GND.n5965 0.00887766
R8240 GND.n6130 GND.n6126 0.00887766
R8241 GND.n7337 GND.n7336 0.00887766
R8242 GND.n7429 GND.n7425 0.00887766
R8243 GND.n5831 GND.n5829 0.00872368
R8244 GND.n5697 GND.n5694 0.00872368
R8245 GND.n821 GND.n772 0.0086117
R8246 GND.n4464 GND.n4456 0.00856452
R8247 GND.n5333 GND.n5332 0.00853947
R8248 GND.n3409 GND.n2030 0.00853768
R8249 GND.n777 GND.n775 0.00834574
R8250 GND.n869 GND.n868 0.00834574
R8251 GND.n6114 GND.n6113 0.00834574
R8252 GND.n7813 GND.n7811 0.00834574
R8253 GND GND.n1435 0.00822246
R8254 GND GND.n6222 0.00806579
R8255 GND.n5764 GND.n5763 0.00806579
R8256 GND.n4661 GND.n4659 0.00783909
R8257 GND.n3212 GND.n3210 0.00783909
R8258 GND.n2259 GND.n2257 0.00783909
R8259 GND.n162 GND.n160 0.00783909
R8260 GND.n1519 GND.n1517 0.00783909
R8261 GND.n5356 GND.n5354 0.00783909
R8262 GND.n3925 GND.n3923 0.00783909
R8263 GND.n5217 GND.n5215 0.00783909
R8264 GND.n3817 GND.n3815 0.00783909
R8265 GND.n3494 GND.n3492 0.00783909
R8266 GND.n1946 GND.n1944 0.00783909
R8267 GND.n2043 GND.n2041 0.00783909
R8268 GND.n2421 GND.n2419 0.00783909
R8269 GND.n2730 GND.n2728 0.00783909
R8270 GND.n4875 GND.n4873 0.00783909
R8271 GND.n2840 GND.n2838 0.00783909
R8272 GND.n1443 GND.n1441 0.00781992
R8273 GND.n828 GND.n826 0.00781383
R8274 GND.n914 GND.n913 0.00781383
R8275 GND.n4556 GND.n4555 0.00779984
R8276 GND.n21 GND.n6 0.00775202
R8277 GND.n7789 GND.n7764 0.00775202
R8278 GND.n659 GND.n644 0.00775202
R8279 GND.n663 GND.n642 0.00775202
R8280 GND.n6346 GND.n6331 0.00775202
R8281 GND.n6322 GND.n6297 0.00775202
R8282 GND.n6287 GND.n6272 0.00775202
R8283 GND.n6291 GND.n6270 0.00775202
R8284 GND.n4462 GND.n4461 0.00769258
R8285 GND.n4450 GND.n4449 0.00769258
R8286 GND.n816 GND.n815 0.00754787
R8287 GND.n4586 GND.n4585 0.00744444
R8288 GND.n4567 GND.n4560 0.00744444
R8289 GND.n6161 GND.n6159 0.00740789
R8290 GND.n4653 GND.n4652 0.00739975
R8291 GND.n3197 GND.n3196 0.00739975
R8292 GND.n2246 GND.n2245 0.00739975
R8293 GND.n154 GND.n153 0.00739975
R8294 GND.n1506 GND.n1505 0.00739975
R8295 GND.n5343 GND.n5342 0.00739975
R8296 GND.n3912 GND.n3911 0.00739975
R8297 GND.n5204 GND.n5203 0.00739975
R8298 GND.n3804 GND.n3803 0.00739975
R8299 GND.n3481 GND.n3480 0.00739975
R8300 GND.n1933 GND.n1932 0.00739975
R8301 GND.n2035 GND.n2034 0.00739975
R8302 GND.n2408 GND.n2407 0.00739975
R8303 GND.n2717 GND.n2716 0.00739975
R8304 GND.n4862 GND.n4861 0.00739975
R8305 GND.n2827 GND.n2826 0.00739975
R8306 GND.n4478 GND.n4477 0.00738379
R8307 GND.n5912 GND.n5908 0.00728191
R8308 GND.n6000 GND.n5999 0.00728191
R8309 GND.n6123 GND.n5858 0.00728191
R8310 GND.n7283 GND.n7279 0.00728191
R8311 GND.n7371 GND.n7370 0.00728191
R8312 GND.n7422 GND.n7421 0.00728191
R8313 GND.n2028 GND.n1445 0.00720761
R8314 GND.n5832 GND.n5831 0.00707895
R8315 GND.n5925 GND.n5923 0.00701596
R8316 GND.n6048 GND.n6047 0.00701596
R8317 GND.n7296 GND.n7294 0.00701596
R8318 GND.n597 GND.n595 0.00701596
R8319 GND.n4179 GND.n4177 0.00675
R8320 GND.n735 GND.n734 0.00675
R8321 GND.n926 GND.n922 0.00675
R8322 GND.n4106 GND.n4105 0.0066794
R8323 GND.n4082 GND.n4081 0.0066794
R8324 GND.n763 GND 0.00661702
R8325 GND GND.n784 0.00661702
R8326 GND.n862 GND 0.00661702
R8327 GND GND.n877 0.00661702
R8328 GND.n960 GND 0.00661702
R8329 GND.n982 GND 0.00661702
R8330 GND GND.n5882 0.00661702
R8331 GND.n5957 GND 0.00661702
R8332 GND GND.n6133 0.00661702
R8333 GND.n6038 GND 0.00661702
R8334 GND.n6086 GND 0.00661702
R8335 GND.n6108 GND 0.00661702
R8336 GND GND.n7253 0.00661702
R8337 GND.n7328 GND 0.00661702
R8338 GND GND.n7432 0.00661702
R8339 GND GND.n7385 0.00661702
R8340 GND GND.n559 0.00661702
R8341 GND.n7817 GND 0.00661702
R8342 GND.n739 GND.n735 0.00648404
R8343 GND.n922 GND.n921 0.00648404
R8344 GND.n5669 GND.n5668 0.00647015
R8345 GND.n5673 GND.n5669 0.00631395
R8346 GND.n5923 GND.n5922 0.00621809
R8347 GND.n6052 GND.n6048 0.00621809
R8348 GND.n7294 GND.n7293 0.00621809
R8349 GND.n595 GND.n594 0.00621809
R8350 GND.n6149 GND 0.00609211
R8351 GND.n6223 GND 0.00609211
R8352 GND.n5780 GND 0.00609211
R8353 GND.n5718 GND 0.00609211
R8354 GND.n4106 GND.n4104 0.00605556
R8355 GND.n991 GND.n990 0.00595213
R8356 GND.n5908 GND.n5907 0.00595213
R8357 GND.n6000 GND.n5970 0.00595213
R8358 GND.n6125 GND.n6123 0.00595213
R8359 GND.n7279 GND.n7278 0.00595213
R8360 GND.n7371 GND.n7341 0.00595213
R8361 GND.n7424 GND.n7422 0.00595213
R8362 GND.n6139 GND.n5656 0.00593478
R8363 GND.n5754 GND.n5753 0.00593421
R8364 GND.n241 GND.n239 0.00585714
R8365 GND.n7648 GND.n7646 0.00585714
R8366 GND.n7208 GND.n7206 0.00585714
R8367 GND.n2604 GND.n2602 0.00585714
R8368 GND.n6896 GND.n6894 0.00585714
R8369 GND.n6742 GND.n6740 0.00585714
R8370 GND.n6583 GND.n6581 0.00585714
R8371 GND.n1040 GND.n1038 0.00585714
R8372 GND.n3691 GND.n3689 0.00585714
R8373 GND.n345 GND.n343 0.00585714
R8374 GND.n483 GND.n481 0.00585714
R8375 GND.n5091 GND.n5089 0.00585714
R8376 GND.n1163 GND.n1161 0.00585714
R8377 GND.n5535 GND.n5533 0.00585714
R8378 GND.n7050 GND.n7048 0.00585714
R8379 GND.n3030 GND.n3028 0.00585714
R8380 GND.n1444 GND.n1364 0.00571186
R8381 GND.n4295 GND.n4293 0.00570833
R8382 GND.n820 GND.n816 0.00568617
R8383 GND.n4738 GND.n4724 0.00557093
R8384 GND.n826 GND.n714 0.00542021
R8385 GND.n914 GND.n871 0.00542021
R8386 GND.n6117 GND.n6116 0.00542021
R8387 GND.n7810 GND.n7808 0.00542021
R8388 GND.n5850 GND.n5849 0.00534496
R8389 GND GND.n5687 0.00510526
R8390 GND.n4948 GND.n4933 0.00507317
R8391 GND.n2784 GND.n2770 0.00507317
R8392 GND.n3234 GND.n3192 0.00507317
R8393 GND.n2893 GND.n2878 0.00507317
R8394 GND.n2337 GND.n2322 0.00507317
R8395 GND.n2121 GND.n2097 0.00507317
R8396 GND.n7740 GND.n7725 0.00507317
R8397 GND.n1596 GND.n1581 0.00507317
R8398 GND.n5436 GND.n5421 0.00507317
R8399 GND.n4003 GND.n3988 0.00507317
R8400 GND.n5301 GND.n5286 0.00507317
R8401 GND.n3891 GND.n3876 0.00507317
R8402 GND.n3564 GND.n3549 0.00507317
R8403 GND.n2023 GND.n2008 0.00507317
R8404 GND.n2491 GND.n2476 0.00507317
R8405 GND.n5837 GND.n5833 0.00505426
R8406 GND.n6148 GND 0.00502899
R8407 GND.n7437 GND.n541 0.00498679
R8408 GND.n775 GND.n714 0.0048883
R8409 GND.n871 GND.n869 0.0048883
R8410 GND.n6116 GND.n6114 0.0048883
R8411 GND.n7811 GND.n7810 0.0048883
R8412 GND.n4564 GND.n4563 0.00476136
R8413 GND.n3132 GND.n3101 0.00469846
R8414 GND.n3390 GND.n3388 0.00469846
R8415 GND.n4055 GND.n4024 0.00469846
R8416 GND.n3254 GND.n3252 0.00466667
R8417 GND.n7557 GND.n7555 0.00466667
R8418 GND.n363 GND.n361 0.00466667
R8419 GND.n7619 GND.n7617 0.00466667
R8420 GND.n259 GND.n257 0.00466667
R8421 GND.n2515 GND.n2513 0.00466667
R8422 GND.n2550 GND.n2548 0.00466667
R8423 GND.n2932 GND.n2930 0.00466667
R8424 GND.n2976 GND.n2974 0.00466667
R8425 GND.n6957 GND.n6956 0.00466667
R8426 GND.n6878 GND.n6875 0.00466667
R8427 GND.n6794 GND.n6792 0.00466667
R8428 GND.n6724 GND.n6721 0.00466667
R8429 GND.n83 GND.n82 0.00466667
R8430 GND.n6679 GND.n6677 0.00466667
R8431 GND.n1027 GND.n1025 0.00466667
R8432 GND.n5560 GND.n5558 0.00466667
R8433 GND.n1253 GND.n1252 0.00466667
R8434 GND.n1179 GND.n1177 0.00466667
R8435 GND.n7495 GND.n7494 0.00466667
R8436 GND.n432 GND.n430 0.00466667
R8437 GND.n4994 GND.n4993 0.00466667
R8438 GND.n5037 GND.n5035 0.00466667
R8439 GND.n3597 GND.n3595 0.00466667
R8440 GND.n3640 GND.n3638 0.00466667
R8441 GND.n1126 GND.n1124 0.00466667
R8442 GND.n1058 GND.n1056 0.00466667
R8443 GND.n6548 GND.n6546 0.00466667
R8444 GND.n6608 GND.n6606 0.00466667
R8445 GND.n7126 GND.n7124 0.00466667
R8446 GND.n7032 GND.n7029 0.00466667
R8447 GND.n3284 GND.n3282 0.00466667
R8448 GND.n6222 GND 0.00466667
R8449 GND.n821 GND.n820 0.00462234
R8450 GND.n5850 GND.n5685 0.00456977
R8451 GND.n7800 GND 0.00456173
R8452 GND.n5666 GND.n5665 0.00454478
R8453 GND.n4116 GND.n4115 0.00438796
R8454 GND.n4131 GND.n4130 0.00438796
R8455 GND.n4146 GND.n4145 0.00438796
R8456 GND.n4161 GND.n4160 0.00438796
R8457 GND.n4177 GND.n4176 0.00438796
R8458 GND.n4195 GND.n4194 0.00438796
R8459 GND.n4210 GND.n4209 0.00438796
R8460 GND.n4225 GND.n4224 0.00438796
R8461 GND.n4240 GND.n4239 0.00438796
R8462 GND.n4265 GND.n4264 0.00438796
R8463 GND.n4284 GND.n4283 0.00438796
R8464 GND.n4304 GND.n4303 0.00438796
R8465 GND.n4319 GND.n4318 0.00438796
R8466 GND.n4334 GND.n4333 0.00438796
R8467 GND.n4349 GND.n4348 0.00438796
R8468 GND.n4364 GND.n4363 0.00438796
R8469 GND.n4381 GND.n4380 0.00438796
R8470 GND.n4396 GND.n4395 0.00438796
R8471 GND.n4411 GND.n4410 0.00438796
R8472 GND.n4426 GND.n4425 0.00438796
R8473 GND.n4441 GND.n4440 0.00438796
R8474 GND.n4064 GND.n4063 0.00438796
R8475 GND.n4433 GND.n4432 0.00438796
R8476 GND.n4417 GND.n4416 0.00438796
R8477 GND.n4402 GND.n4401 0.00438796
R8478 GND.n4387 GND.n4386 0.00438796
R8479 GND.n4372 GND.n4371 0.00438796
R8480 GND.n4355 GND.n4354 0.00438796
R8481 GND.n4340 GND.n4339 0.00438796
R8482 GND.n4325 GND.n4324 0.00438796
R8483 GND.n4310 GND.n4309 0.00438796
R8484 GND.n4293 GND.n4292 0.00438796
R8485 GND.n4274 GND.n4273 0.00438796
R8486 GND.n4256 GND.n4255 0.00438796
R8487 GND.n4231 GND.n4230 0.00438796
R8488 GND.n4216 GND.n4215 0.00438796
R8489 GND.n4201 GND.n4200 0.00438796
R8490 GND.n4186 GND.n4185 0.00438796
R8491 GND.n4167 GND.n4166 0.00438796
R8492 GND.n4152 GND.n4151 0.00438796
R8493 GND.n4137 GND.n4136 0.00438796
R8494 GND.n4122 GND.n4121 0.00438796
R8495 GND.n990 GND.n988 0.00435638
R8496 GND.n5970 GND.n5966 0.00435638
R8497 GND.n6126 GND.n6125 0.00435638
R8498 GND.n7341 GND.n7337 0.00435638
R8499 GND.n7425 GND.n7424 0.00435638
R8500 GND.n3349 GND.n3344 0.00425
R8501 GND.n7536 GND.n7531 0.00425
R8502 GND.n7598 GND.n7593 0.00425
R8503 GND.n2652 GND.n2647 0.00425
R8504 GND.n3078 GND.n3073 0.00425
R8505 GND.n6971 GND.n6939 0.00425
R8506 GND.n6817 GND.n6776 0.00425
R8507 GND.n7749 GND.n65 0.00425
R8508 GND.n5633 GND.n1009 0.00425
R8509 GND.n5449 GND.n1238 0.00425
R8510 GND.n7474 GND.n7469 0.00425
R8511 GND.n5139 GND.n5134 0.00425
R8512 GND.n3739 GND.n3734 0.00425
R8513 GND.n5506 GND.n1108 0.00425
R8514 GND.n6527 GND.n6513 0.00425
R8515 GND.n7105 GND.n7100 0.00425
R8516 GND.n3388 GND.n3387 0.00420666
R8517 GND.n3387 GND.n3386 0.00420666
R8518 GND.n3132 GND.n3131 0.00420666
R8519 GND.n3131 GND.n3130 0.00420666
R8520 GND.n4055 GND.n4054 0.00420666
R8521 GND.n4054 GND.n4053 0.00420666
R8522 GND.n5192 GND.n5179 0.00420666
R8523 GND.n5179 GND.n5178 0.00420666
R8524 GND.n3791 GND.n3778 0.00420666
R8525 GND.n3778 GND.n3777 0.00420666
R8526 GND.n1326 GND.n1313 0.00420666
R8527 GND.n1313 GND.n1312 0.00420666
R8528 GND.n3469 GND.n3456 0.00420666
R8529 GND.n3456 GND.n3455 0.00420666
R8530 GND.n1494 GND.n1481 0.00420666
R8531 GND.n1481 GND.n1480 0.00420666
R8532 GND.n1920 GND.n1907 0.00420666
R8533 GND.n1907 GND.n1906 0.00420666
R8534 GND.n143 GND.n130 0.00420666
R8535 GND.n130 GND.n129 0.00420666
R8536 GND.n2171 GND.n2158 0.00420666
R8537 GND.n2158 GND.n2157 0.00420666
R8538 GND.n2233 GND.n2220 0.00420666
R8539 GND.n2220 GND.n2219 0.00420666
R8540 GND.n2396 GND.n2383 0.00420666
R8541 GND.n2383 GND.n2382 0.00420666
R8542 GND.n2708 GND.n2707 0.00420666
R8543 GND.n2707 GND.n2706 0.00420666
R8544 GND.n4849 GND.n4836 0.00420666
R8545 GND.n4836 GND.n4835 0.00420666
R8546 GND.n4642 GND.n4629 0.00420666
R8547 GND.n4629 GND.n4628 0.00420666
R8548 GND.n5922 GND.n5918 0.00409043
R8549 GND.n7293 GND.n7289 0.00409043
R8550 GND.n4287 GND.n4285 0.00397222
R8551 GND.n3028 GND.n3027 0.00396756
R8552 GND.n3294 GND.n3293 0.00396756
R8553 GND.n2602 GND.n2601 0.00396756
R8554 GND.n2986 GND.n2985 0.00396756
R8555 GND.n7206 GND.n7205 0.00396756
R8556 GND.n2560 GND.n2559 0.00396756
R8557 GND.n7048 GND.n7047 0.00396756
R8558 GND.n7160 GND.n7159 0.00396756
R8559 GND.n6894 GND.n6893 0.00396756
R8560 GND.n6997 GND.n6996 0.00396756
R8561 GND.n6740 GND.n6739 0.00396756
R8562 GND.n6843 GND.n6842 0.00396756
R8563 GND.n6581 GND.n6580 0.00396756
R8564 GND.n6689 GND.n6688 0.00396756
R8565 GND.n5533 GND.n5532 0.00396756
R8566 GND.n6618 GND.n6617 0.00396756
R8567 GND.n1038 GND.n1037 0.00396756
R8568 GND.n5570 GND.n5569 0.00396756
R8569 GND.n1161 GND.n1160 0.00396756
R8570 GND.n1068 GND.n1067 0.00396756
R8571 GND.n3689 GND.n3688 0.00396756
R8572 GND.n1189 GND.n1188 0.00396756
R8573 GND.n5089 GND.n5088 0.00396756
R8574 GND.n3650 GND.n3649 0.00396756
R8575 GND.n481 GND.n480 0.00396756
R8576 GND.n5047 GND.n5046 0.00396756
R8577 GND.n343 GND.n342 0.00396756
R8578 GND.n442 GND.n441 0.00396756
R8579 GND.n239 GND.n238 0.00396756
R8580 GND.n373 GND.n372 0.00396756
R8581 GND.n7646 GND.n7645 0.00396756
R8582 GND.n269 GND.n268 0.00396756
R8583 GND.n5796 GND.n5795 0.00396053
R8584 GND.n7539 GND.n7538 0.00395031
R8585 GND.n7601 GND.n7600 0.00395031
R8586 GND.n2655 GND.n2654 0.00395031
R8587 GND.n3081 GND.n3080 0.00395031
R8588 GND.n6965 GND.n6964 0.00395031
R8589 GND.n6802 GND.n6801 0.00395031
R8590 GND.n7747 GND.n7746 0.00395031
R8591 GND.n5627 GND.n5626 0.00395031
R8592 GND.n5443 GND.n5442 0.00395031
R8593 GND.n7477 GND.n7476 0.00395031
R8594 GND.n5142 GND.n5141 0.00395031
R8595 GND.n3742 GND.n3741 0.00395031
R8596 GND.n5491 GND.n5490 0.00395031
R8597 GND.n6530 GND.n6529 0.00395031
R8598 GND.n7108 GND.n7107 0.00395031
R8599 GND.n3352 GND.n3351 0.00395031
R8600 GND.n3027 GND.n3026 0.0039133
R8601 GND.n3026 GND.t1324 0.0039133
R8602 GND.n3293 GND.n3292 0.0039133
R8603 GND.n3292 GND.t1393 0.0039133
R8604 GND.n2601 GND.n2600 0.0039133
R8605 GND.n2600 GND.t1489 0.0039133
R8606 GND.n2985 GND.n2984 0.0039133
R8607 GND.n2984 GND.t605 0.0039133
R8608 GND.n7205 GND.n7204 0.0039133
R8609 GND.n7204 GND.t398 0.0039133
R8610 GND.n2559 GND.n2558 0.0039133
R8611 GND.n2558 GND.t15 0.0039133
R8612 GND.n7047 GND.n7046 0.0039133
R8613 GND.n7046 GND.t1503 0.0039133
R8614 GND.n7159 GND.n7158 0.0039133
R8615 GND.n7158 GND.t1109 0.0039133
R8616 GND.n6893 GND.n6892 0.0039133
R8617 GND.n6892 GND.t27 0.0039133
R8618 GND.n6996 GND.n6995 0.0039133
R8619 GND.n6995 GND.t9 0.0039133
R8620 GND.n6739 GND.n6738 0.0039133
R8621 GND.n6738 GND.t1177 0.0039133
R8622 GND.n6842 GND.n6841 0.0039133
R8623 GND.n6841 GND.t530 0.0039133
R8624 GND.n6580 GND.n6579 0.0039133
R8625 GND.n6579 GND.t1435 0.0039133
R8626 GND.n6688 GND.n6687 0.0039133
R8627 GND.n6687 GND.t1401 0.0039133
R8628 GND.n5532 GND.n5531 0.0039133
R8629 GND.n5531 GND.t1329 0.0039133
R8630 GND.n6617 GND.n6616 0.0039133
R8631 GND.n6616 GND.t1058 0.0039133
R8632 GND.n1037 GND.n1036 0.0039133
R8633 GND.n1036 GND.t512 0.0039133
R8634 GND.n5569 GND.n5568 0.0039133
R8635 GND.n5568 GND.t1529 0.0039133
R8636 GND.n1160 GND.n1159 0.0039133
R8637 GND.n1159 GND.t1369 0.0039133
R8638 GND.n1067 GND.n1066 0.0039133
R8639 GND.n1066 GND.t632 0.0039133
R8640 GND.n3688 GND.n3687 0.0039133
R8641 GND.n3687 GND.t410 0.0039133
R8642 GND.n1188 GND.n1187 0.0039133
R8643 GND.n1187 GND.t583 0.0039133
R8644 GND.n5088 GND.n5087 0.0039133
R8645 GND.n5087 GND.t470 0.0039133
R8646 GND.n3649 GND.n3648 0.0039133
R8647 GND.n3648 GND.t1028 0.0039133
R8648 GND.n480 GND.n479 0.0039133
R8649 GND.n479 GND.t1478 0.0039133
R8650 GND.n5046 GND.n5045 0.0039133
R8651 GND.n5045 GND.t618 0.0039133
R8652 GND.n342 GND.n341 0.0039133
R8653 GND.n341 GND.t875 0.0039133
R8654 GND.n441 GND.n440 0.0039133
R8655 GND.n440 GND.t1513 0.0039133
R8656 GND.n238 GND.n237 0.0039133
R8657 GND.n237 GND.t1338 0.0039133
R8658 GND.n372 GND.n371 0.0039133
R8659 GND.n371 GND.t70 0.0039133
R8660 GND.n7645 GND.n7644 0.0039133
R8661 GND.n7644 GND.t1080 0.0039133
R8662 GND.n268 GND.n267 0.0039133
R8663 GND.n267 GND.t478 0.0039133
R8664 GND.n3348 GND.n3347 0.00390909
R8665 GND.n3341 GND.n3340 0.00390909
R8666 GND.n7535 GND.n7534 0.00390909
R8667 GND.n7528 GND.n7527 0.00390909
R8668 GND.n7597 GND.n7596 0.00390909
R8669 GND.n7590 GND.n7589 0.00390909
R8670 GND.n2651 GND.n2650 0.00390909
R8671 GND.n2644 GND.n2643 0.00390909
R8672 GND.n3077 GND.n3076 0.00390909
R8673 GND.n3070 GND.n3069 0.00390909
R8674 GND.n6970 GND.n6969 0.00390909
R8675 GND.n6936 GND.n6935 0.00390909
R8676 GND.n6816 GND.n6815 0.00390909
R8677 GND.n6813 GND.n6812 0.00390909
R8678 GND.n7750 GND.n64 0.00390909
R8679 GND.n61 GND.n60 0.00390909
R8680 GND.n5632 GND.n5631 0.00390909
R8681 GND.n1006 GND.n1005 0.00390909
R8682 GND.n5448 GND.n5447 0.00390909
R8683 GND.n1235 GND.n1234 0.00390909
R8684 GND.n7473 GND.n7472 0.00390909
R8685 GND.n7466 GND.n7465 0.00390909
R8686 GND.n5138 GND.n5137 0.00390909
R8687 GND.n5131 GND.n5130 0.00390909
R8688 GND.n3738 GND.n3737 0.00390909
R8689 GND.n3731 GND.n3730 0.00390909
R8690 GND.n5505 GND.n5504 0.00390909
R8691 GND.n5502 GND.n5501 0.00390909
R8692 GND.n6526 GND.n6525 0.00390909
R8693 GND.n6523 GND.n6522 0.00390909
R8694 GND.n7104 GND.n7103 0.00390909
R8695 GND.n7097 GND.n7096 0.00390909
R8696 GND.n921 GND.n919 0.00382447
R8697 GND.n6047 GND.n6045 0.00379255
R8698 GND.n7378 GND.n597 0.00379255
R8699 GND.n1444 GND.n1443 0.00377331
R8700 GND.n734 GND.n730 0.00355851
R8701 GND.n5913 GND.n5912 0.0035266
R8702 GND.n7284 GND.n7283 0.0035266
R8703 GND.n3315 GND.n3314 0.0034846
R8704 GND.n3043 GND.n3042 0.0034846
R8705 GND.n2617 GND.n2616 0.0034846
R8706 GND.n7221 GND.n7220 0.0034846
R8707 GND.n7063 GND.n7062 0.0034846
R8708 GND.n6909 GND.n6908 0.0034846
R8709 GND.n6755 GND.n6754 0.0034846
R8710 GND.n6642 GND.n6641 0.0034846
R8711 GND.n5594 GND.n5593 0.0034846
R8712 GND.n1092 GND.n1091 0.0034846
R8713 GND.n1213 GND.n1212 0.0034846
R8714 GND.n3704 GND.n3703 0.0034846
R8715 GND.n5104 GND.n5103 0.0034846
R8716 GND.n496 GND.n495 0.0034846
R8717 GND.n397 GND.n396 0.0034846
R8718 GND.n293 GND.n292 0.0034846
R8719 GND.n3314 GND.n3313 0.00343883
R8720 GND.n3313 GND.n3312 0.00343883
R8721 GND.n3039 GND.n3038 0.00343883
R8722 GND.n3040 GND.n3039 0.00343883
R8723 GND.n3042 GND.n3041 0.00343883
R8724 GND.n3041 GND.n3040 0.00343883
R8725 GND.n2613 GND.n2612 0.00343883
R8726 GND.n2614 GND.n2613 0.00343883
R8727 GND.n2616 GND.n2615 0.00343883
R8728 GND.n2615 GND.n2614 0.00343883
R8729 GND.n7217 GND.n7216 0.00343883
R8730 GND.n7218 GND.n7217 0.00343883
R8731 GND.n7220 GND.n7219 0.00343883
R8732 GND.n7219 GND.n7218 0.00343883
R8733 GND.n7059 GND.n7058 0.00343883
R8734 GND.n7060 GND.n7059 0.00343883
R8735 GND.n7062 GND.n7061 0.00343883
R8736 GND.n7061 GND.n7060 0.00343883
R8737 GND.n6905 GND.n6904 0.00343883
R8738 GND.n6906 GND.n6905 0.00343883
R8739 GND.n6908 GND.n6907 0.00343883
R8740 GND.n6907 GND.n6906 0.00343883
R8741 GND.n6751 GND.n6750 0.00343883
R8742 GND.n6752 GND.n6751 0.00343883
R8743 GND.n6754 GND.n6753 0.00343883
R8744 GND.n6753 GND.n6752 0.00343883
R8745 GND.n6646 GND.n6645 0.00343883
R8746 GND.n6645 GND.n6644 0.00343883
R8747 GND.n6643 GND.n6642 0.00343883
R8748 GND.n6644 GND.n6643 0.00343883
R8749 GND.n5598 GND.n5597 0.00343883
R8750 GND.n5597 GND.n5596 0.00343883
R8751 GND.n5595 GND.n5594 0.00343883
R8752 GND.n5596 GND.n5595 0.00343883
R8753 GND.n1096 GND.n1095 0.00343883
R8754 GND.n1095 GND.n1094 0.00343883
R8755 GND.n1093 GND.n1092 0.00343883
R8756 GND.n1094 GND.n1093 0.00343883
R8757 GND.n1217 GND.n1216 0.00343883
R8758 GND.n1216 GND.n1215 0.00343883
R8759 GND.n1214 GND.n1213 0.00343883
R8760 GND.n1215 GND.n1214 0.00343883
R8761 GND.n3700 GND.n3699 0.00343883
R8762 GND.n3701 GND.n3700 0.00343883
R8763 GND.n3703 GND.n3702 0.00343883
R8764 GND.n3702 GND.n3701 0.00343883
R8765 GND.n5100 GND.n5099 0.00343883
R8766 GND.n5101 GND.n5100 0.00343883
R8767 GND.n5103 GND.n5102 0.00343883
R8768 GND.n5102 GND.n5101 0.00343883
R8769 GND.n492 GND.n491 0.00343883
R8770 GND.n493 GND.n492 0.00343883
R8771 GND.n495 GND.n494 0.00343883
R8772 GND.n494 GND.n493 0.00343883
R8773 GND.n401 GND.n400 0.00343883
R8774 GND.n400 GND.n399 0.00343883
R8775 GND.n398 GND.n397 0.00343883
R8776 GND.n399 GND.n398 0.00343883
R8777 GND.n297 GND.n296 0.00343883
R8778 GND.n296 GND.n295 0.00343883
R8779 GND.n294 GND.n293 0.00343883
R8780 GND.n295 GND.n294 0.00343883
R8781 GND.n7657 GND.n7656 0.00343883
R8782 GND.n7658 GND.n7657 0.00343883
R8783 GND GND.n6379 0.00340123
R8784 GND.n7800 GND 0.00340123
R8785 GND.n6212 GND 0.00327778
R8786 GND.n6205 GND 0.00327778
R8787 GND.n6149 GND.n6148 0.00313158
R8788 GND.n2520 GND.n2519 0.00308428
R8789 GND.n2937 GND.n2936 0.00308428
R8790 GND.n1258 GND.n1257 0.00308428
R8791 GND.n3602 GND.n3601 0.00308428
R8792 GND.n6422 GND.n6421 0.00307458
R8793 GND.n970 GND.n968 0.0030266
R8794 GND.n5999 GND.n5997 0.0030266
R8795 GND.n6004 GND.n5858 0.0030266
R8796 GND.n7370 GND.n7368 0.0030266
R8797 GND.n7421 GND.n7417 0.0030266
R8798 GND.n3344 GND.n3343 0.003
R8799 GND.n7531 GND.n7530 0.003
R8800 GND.n7593 GND.n7592 0.003
R8801 GND.n2647 GND.n2646 0.003
R8802 GND.n3073 GND.n3072 0.003
R8803 GND.n6939 GND.n6938 0.003
R8804 GND.n6776 GND.n6775 0.003
R8805 GND.n1009 GND.n1008 0.003
R8806 GND.n1238 GND.n1237 0.003
R8807 GND.n7469 GND.n7468 0.003
R8808 GND.n5134 GND.n5133 0.003
R8809 GND.n3734 GND.n3733 0.003
R8810 GND.n1108 GND.n1107 0.003
R8811 GND.n6513 GND.n6512 0.003
R8812 GND.n7100 GND.n7099 0.003
R8813 GND.n4110 GND.n4109 0.00299232
R8814 GND.n5833 GND.n5832 0.00292248
R8815 GND.n6455 GND.n6454 0.00290385
R8816 GND.n540 GND.n539 0.00290385
R8817 GND.n4952 GND.n4951 0.00285
R8818 GND.n4973 GND.n4768 0.00285
R8819 GND.n2346 GND.n2340 0.00285
R8820 GND.n7743 GND.n150 0.00285
R8821 GND.n5330 GND.n1599 0.00285
R8822 GND.n5439 GND.n5337 0.00285
R8823 GND.n5313 GND.n4061 0.00285
R8824 GND.n5310 GND.n5304 0.00285
R8825 GND.n3895 GND.n3894 0.00285
R8826 GND.n3568 GND.n3567 0.00285
R8827 GND.n3411 GND.n2026 0.00285
R8828 GND.n2185 GND.n2179 0.00285
R8829 GND.n2500 GND.n2494 0.00285
R8830 GND.n2815 GND.n2809 0.00285
R8831 GND.n3144 GND.n3138 0.00285
R8832 GND.n3402 GND.n3396 0.00285
R8833 GND.n6226 GND.n6224 0.00280263
R8834 GND.n6477 GND.n6474 0.00277946
R8835 GND.n6387 GND.n6384 0.00277946
R8836 GND.n760 GND 0.00276064
R8837 GND.n785 GND 0.00276064
R8838 GND.n859 GND 0.00276064
R8839 GND.n878 GND 0.00276064
R8840 GND.n957 GND 0.00276064
R8841 GND GND.n970 0.00276064
R8842 GND.n985 GND 0.00276064
R8843 GND.n973 GND 0.00276064
R8844 GND.n5883 GND 0.00276064
R8845 GND.n5954 GND 0.00276064
R8846 GND.n6134 GND 0.00276064
R8847 GND.n6035 GND 0.00276064
R8848 GND.n6083 GND 0.00276064
R8849 GND GND.n6096 0.00276064
R8850 GND.n6111 GND 0.00276064
R8851 GND.n6099 GND 0.00276064
R8852 GND.n7254 GND 0.00276064
R8853 GND.n7325 GND 0.00276064
R8854 GND.n7433 GND 0.00276064
R8855 GND.n7386 GND 0.00276064
R8856 GND.n560 GND 0.00276064
R8857 GND.n2 GND 0.00276064
R8858 GND.n7814 GND 0.00276064
R8859 GND GND.n7827 0.00276064
R8860 GND.n2887 GND.n2886 0.00266776
R8861 GND.n5295 GND.n5294 0.00266776
R8862 GND.n5430 GND.n5429 0.00266776
R8863 GND.n1590 GND.n1589 0.00266776
R8864 GND.n7734 GND.n7733 0.00266776
R8865 GND.n2331 GND.n2330 0.00266776
R8866 GND.n4942 GND.n4941 0.00266776
R8867 GND.n373 GND.n369 0.00258333
R8868 GND.n269 GND.n265 0.00258333
R8869 GND.n2560 GND.n2556 0.00258333
R8870 GND.n2986 GND.n2982 0.00258333
R8871 GND.n6997 GND.n6993 0.00258333
R8872 GND.n6843 GND.n6839 0.00258333
R8873 GND.n6689 GND.n6685 0.00258333
R8874 GND.n5570 GND.n5566 0.00258333
R8875 GND.n1189 GND.n1185 0.00258333
R8876 GND.n442 GND.n438 0.00258333
R8877 GND.n5047 GND.n5043 0.00258333
R8878 GND.n3650 GND.n3646 0.00258333
R8879 GND.n1068 GND.n1064 0.00258333
R8880 GND.n6618 GND.n6614 0.00258333
R8881 GND.n7160 GND.n7156 0.00258333
R8882 GND.n3294 GND.n3290 0.00258333
R8883 GND.n4473 GND.n4472 0.00253688
R8884 GND.n4464 GND.n4463 0.00253688
R8885 GND.n4447 GND.n4446 0.00250907
R8886 GND.n4435 GND.n4434 0.00250907
R8887 GND.n4419 GND.n4418 0.00250907
R8888 GND.n4404 GND.n4403 0.00250907
R8889 GND.n4389 GND.n4388 0.00250907
R8890 GND.n4374 GND.n4373 0.00250907
R8891 GND.n4357 GND.n4356 0.00250907
R8892 GND.n4342 GND.n4341 0.00250907
R8893 GND.n4327 GND.n4326 0.00250907
R8894 GND.n4312 GND.n4311 0.00250907
R8895 GND.n4297 GND.n4296 0.00250907
R8896 GND.n4276 GND.n4275 0.00250907
R8897 GND.n4258 GND.n4257 0.00250907
R8898 GND.n4233 GND.n4232 0.00250907
R8899 GND.n4218 GND.n4217 0.00250907
R8900 GND.n4203 GND.n4202 0.00250907
R8901 GND.n4188 GND.n4187 0.00250907
R8902 GND.n4169 GND.n4168 0.00250907
R8903 GND.n4154 GND.n4153 0.00250907
R8904 GND.n4139 GND.n4138 0.00250907
R8905 GND.n4124 GND.n4123 0.00250907
R8906 GND.n4114 GND.n4113 0.00250907
R8907 GND.n4129 GND.n4128 0.00250907
R8908 GND.n4144 GND.n4143 0.00250907
R8909 GND.n4159 GND.n4158 0.00250907
R8910 GND.n4174 GND.n4173 0.00250907
R8911 GND.n4193 GND.n4192 0.00250907
R8912 GND.n4208 GND.n4207 0.00250907
R8913 GND.n4223 GND.n4222 0.00250907
R8914 GND.n4238 GND.n4237 0.00250907
R8915 GND.n4263 GND.n4262 0.00250907
R8916 GND.n4281 GND.n4280 0.00250907
R8917 GND.n4302 GND.n4301 0.00250907
R8918 GND.n4317 GND.n4316 0.00250907
R8919 GND.n4332 GND.n4331 0.00250907
R8920 GND.n4347 GND.n4346 0.00250907
R8921 GND.n4362 GND.n4361 0.00250907
R8922 GND.n4379 GND.n4378 0.00250907
R8923 GND.n4394 GND.n4393 0.00250907
R8924 GND.n4409 GND.n4408 0.00250907
R8925 GND.n4424 GND.n4423 0.00250907
R8926 GND.n4439 GND.n4438 0.00250907
R8927 GND.n4443 GND.n4442 0.00250907
R8928 GND.n829 GND.n828 0.00249468
R8929 GND.n913 GND.n909 0.00249468
R8930 GND.n6096 GND.n6094 0.00249468
R8931 GND.n3 GND.n2 0.00249468
R8932 GND.n4112 GND.t432 0.00247763
R8933 GND.n4127 GND.t1036 0.00247763
R8934 GND.n4142 GND.t429 0.00247763
R8935 GND.n4157 GND.t1569 0.00247763
R8936 GND.n4172 GND.t1316 0.00247763
R8937 GND.n4191 GND.t433 0.00247763
R8938 GND.n4206 GND.t1567 0.00247763
R8939 GND.n4221 GND.t1034 0.00247763
R8940 GND.n4236 GND.t1315 0.00247763
R8941 GND.n4261 GND.t1568 0.00247763
R8942 GND.n4279 GND.t1565 0.00247763
R8943 GND.n4300 GND.t431 0.00247763
R8944 GND.n4315 GND.t1317 0.00247763
R8945 GND.n4330 GND.t1037 0.00247763
R8946 GND.n4345 GND.t1313 0.00247763
R8947 GND.n4360 GND.t428 0.00247763
R8948 GND.n4377 GND.t1035 0.00247763
R8949 GND.n4392 GND.t1318 0.00247763
R8950 GND.n4407 GND.t1038 0.00247763
R8951 GND.n4422 GND.t1314 0.00247763
R8952 GND.n4420 GND.n4419 0.00247763
R8953 GND.t1314 GND.n4420 0.00247763
R8954 GND.n4405 GND.n4404 0.00247763
R8955 GND.t1038 GND.n4405 0.00247763
R8956 GND.n4390 GND.n4389 0.00247763
R8957 GND.t1318 GND.n4390 0.00247763
R8958 GND.n4375 GND.n4374 0.00247763
R8959 GND.t1035 GND.n4375 0.00247763
R8960 GND.n4358 GND.n4357 0.00247763
R8961 GND.t428 GND.n4358 0.00247763
R8962 GND.n4343 GND.n4342 0.00247763
R8963 GND.t1313 GND.n4343 0.00247763
R8964 GND.n4328 GND.n4327 0.00247763
R8965 GND.t1037 GND.n4328 0.00247763
R8966 GND.n4313 GND.n4312 0.00247763
R8967 GND.t1317 GND.n4313 0.00247763
R8968 GND.n4298 GND.n4297 0.00247763
R8969 GND.t431 GND.n4298 0.00247763
R8970 GND.n4277 GND.n4276 0.00247763
R8971 GND.t1565 GND.n4277 0.00247763
R8972 GND.n4259 GND.n4258 0.00247763
R8973 GND.t1568 GND.n4259 0.00247763
R8974 GND.n4234 GND.n4233 0.00247763
R8975 GND.t1315 GND.n4234 0.00247763
R8976 GND.n4219 GND.n4218 0.00247763
R8977 GND.t1034 GND.n4219 0.00247763
R8978 GND.n4204 GND.n4203 0.00247763
R8979 GND.t1567 GND.n4204 0.00247763
R8980 GND.n4189 GND.n4188 0.00247763
R8981 GND.t433 GND.n4189 0.00247763
R8982 GND.n4170 GND.n4169 0.00247763
R8983 GND.t1316 GND.n4170 0.00247763
R8984 GND.n4155 GND.n4154 0.00247763
R8985 GND.t1569 GND.n4155 0.00247763
R8986 GND.n4140 GND.n4139 0.00247763
R8987 GND.t429 GND.n4140 0.00247763
R8988 GND.n4125 GND.n4124 0.00247763
R8989 GND.t1036 GND.n4125 0.00247763
R8990 GND.n4111 GND.n4110 0.00247763
R8991 GND.t432 GND.n4111 0.00247763
R8992 GND.n4113 GND.n4112 0.00247763
R8993 GND.n4128 GND.n4127 0.00247763
R8994 GND.n4143 GND.n4142 0.00247763
R8995 GND.n4158 GND.n4157 0.00247763
R8996 GND.n4173 GND.n4172 0.00247763
R8997 GND.n4192 GND.n4191 0.00247763
R8998 GND.n4207 GND.n4206 0.00247763
R8999 GND.n4222 GND.n4221 0.00247763
R9000 GND.n4237 GND.n4236 0.00247763
R9001 GND.n4262 GND.n4261 0.00247763
R9002 GND.n4280 GND.n4279 0.00247763
R9003 GND.n4301 GND.n4300 0.00247763
R9004 GND.n4316 GND.n4315 0.00247763
R9005 GND.n4331 GND.n4330 0.00247763
R9006 GND.n4346 GND.n4345 0.00247763
R9007 GND.n4361 GND.n4360 0.00247763
R9008 GND.n4378 GND.n4377 0.00247763
R9009 GND.n4393 GND.n4392 0.00247763
R9010 GND.n4408 GND.n4407 0.00247763
R9011 GND.n4423 GND.n4422 0.00247763
R9012 GND.n4438 GND.n4437 0.00247763
R9013 GND.n4437 GND.t430 0.00247763
R9014 GND.n4436 GND.n4435 0.00247763
R9015 GND.t430 GND.n4436 0.00247763
R9016 GND.n4446 GND.n4445 0.00247763
R9017 GND.n4445 GND.t497 0.00247763
R9018 GND.t497 GND.n4444 0.00247763
R9019 GND.n4444 GND.n4443 0.00247763
R9020 GND.n6222 GND 0.00247368
R9021 GND.n3351 GND.n3350 0.00245833
R9022 GND.n7538 GND.n7537 0.00245833
R9023 GND.n7600 GND.n7599 0.00245833
R9024 GND.n2654 GND.n2653 0.00245833
R9025 GND.n3080 GND.n3079 0.00245833
R9026 GND.n6966 GND.n6965 0.00245833
R9027 GND.n6803 GND.n6802 0.00245833
R9028 GND.n7748 GND.n7747 0.00245833
R9029 GND.n5628 GND.n5627 0.00245833
R9030 GND.n5444 GND.n5443 0.00245833
R9031 GND.n7476 GND.n7475 0.00245833
R9032 GND.n5141 GND.n5140 0.00245833
R9033 GND.n3741 GND.n3740 0.00245833
R9034 GND.n5492 GND.n5491 0.00245833
R9035 GND.n6529 GND.n6528 0.00245833
R9036 GND.n7107 GND.n7106 0.00245833
R9037 GND.n396 GND.n395 0.00228571
R9038 GND.n292 GND.n291 0.00228571
R9039 GND.n2617 GND.n2582 0.00228571
R9040 GND.n3043 GND.n3008 0.00228571
R9041 GND.n7063 GND.n7019 0.00228571
R9042 GND.n6909 GND.n6865 0.00228571
R9043 GND.n6755 GND.n6711 0.00228571
R9044 GND.n5593 GND.n5592 0.00228571
R9045 GND.n1212 GND.n1211 0.00228571
R9046 GND.n496 GND.n464 0.00228571
R9047 GND.n5104 GND.n5069 0.00228571
R9048 GND.n3704 GND.n3672 0.00228571
R9049 GND.n1091 GND.n1090 0.00228571
R9050 GND.n6641 GND.n6640 0.00228571
R9051 GND.n7221 GND.n7182 0.00228571
R9052 GND.n3315 GND.n3311 0.00228571
R9053 GND.n4658 GND 0.00217027
R9054 GND.n3209 GND 0.00217027
R9055 GND.n2256 GND 0.00217027
R9056 GND.n159 GND 0.00217027
R9057 GND.n1516 GND 0.00217027
R9058 GND.n5353 GND 0.00217027
R9059 GND.n3922 GND 0.00217027
R9060 GND.n5214 GND 0.00217027
R9061 GND.n3814 GND 0.00217027
R9062 GND.n3491 GND 0.00217027
R9063 GND.n1943 GND 0.00217027
R9064 GND.n2040 GND 0.00217027
R9065 GND.n2418 GND 0.00217027
R9066 GND.n2727 GND 0.00217027
R9067 GND.n4872 GND 0.00217027
R9068 GND.n2837 GND 0.00217027
R9069 GND.n2030 GND.n2028 0.00200519
R9070 GND.n4767 GND.n4766 0.00199276
R9071 GND.n2808 GND.n2807 0.00199276
R9072 GND.n2028 GND.n2027 0.00195117
R9073 GND.n6387 GND.n6386 0.00193331
R9074 GND.n6477 GND.n6476 0.00193331
R9075 GND.n4285 GND.n4284 0.00188889
R9076 GND.n4552 GND.n4551 0.00186977
R9077 GND.n4553 GND.n4552 0.00186977
R9078 GND.n3282 GND.n3281 0.00183506
R9079 GND.n2974 GND.n2973 0.00183506
R9080 GND.n2548 GND.n2547 0.00183506
R9081 GND.n7032 GND.n7031 0.00183506
R9082 GND.n6878 GND.n6877 0.00183506
R9083 GND.n6724 GND.n6723 0.00183506
R9084 GND.n6677 GND.n6676 0.00183506
R9085 GND.n6606 GND.n6605 0.00183506
R9086 GND.n5558 GND.n5557 0.00183506
R9087 GND.n1056 GND.n1055 0.00183506
R9088 GND.n1177 GND.n1176 0.00183506
R9089 GND.n3638 GND.n3637 0.00183506
R9090 GND.n5035 GND.n5034 0.00183506
R9091 GND.n430 GND.n429 0.00183506
R9092 GND.n361 GND.n360 0.00183506
R9093 GND.n257 GND.n256 0.00183506
R9094 GND.n3281 GND.n3280 0.00181454
R9095 GND.n3019 GND.n3018 0.00181454
R9096 GND.n3018 GND.n3017 0.00181454
R9097 GND.n2973 GND.n2972 0.00181454
R9098 GND.n2588 GND.n2587 0.00181454
R9099 GND.n2587 GND.n2586 0.00181454
R9100 GND.n2547 GND.n2546 0.00181454
R9101 GND.n7190 GND.n7189 0.00181454
R9102 GND.n7189 GND.n7188 0.00181454
R9103 GND.n7031 GND.n7030 0.00181454
R9104 GND.n7027 GND.n7026 0.00181454
R9105 GND.n7026 GND.n7025 0.00181454
R9106 GND.n6877 GND.n6876 0.00181454
R9107 GND.n6873 GND.n6872 0.00181454
R9108 GND.n6872 GND.n6871 0.00181454
R9109 GND.n6723 GND.n6722 0.00181454
R9110 GND.n6719 GND.n6718 0.00181454
R9111 GND.n6718 GND.n6717 0.00181454
R9112 GND.n6676 GND.n6675 0.00181454
R9113 GND.n6570 GND.n6569 0.00181454
R9114 GND.n6569 GND.n6568 0.00181454
R9115 GND.n6605 GND.n6604 0.00181454
R9116 GND.n6595 GND.n6594 0.00181454
R9117 GND.n6594 GND.n6593 0.00181454
R9118 GND.n5557 GND.n5556 0.00181454
R9119 GND.n5547 GND.n5546 0.00181454
R9120 GND.n5546 GND.n5545 0.00181454
R9121 GND.n1055 GND.n1054 0.00181454
R9122 GND.n1152 GND.n1151 0.00181454
R9123 GND.n1151 GND.n1150 0.00181454
R9124 GND.n1176 GND.n1175 0.00181454
R9125 GND.n3678 GND.n3677 0.00181454
R9126 GND.n3677 GND.n3676 0.00181454
R9127 GND.n3637 GND.n3636 0.00181454
R9128 GND.n5075 GND.n5074 0.00181454
R9129 GND.n5074 GND.n5073 0.00181454
R9130 GND.n5034 GND.n5033 0.00181454
R9131 GND.n470 GND.n469 0.00181454
R9132 GND.n469 GND.n468 0.00181454
R9133 GND.n429 GND.n428 0.00181454
R9134 GND.n332 GND.n331 0.00181454
R9135 GND.n331 GND.n330 0.00181454
R9136 GND.n360 GND.n359 0.00181454
R9137 GND.n230 GND.n229 0.00181454
R9138 GND.n229 GND.n228 0.00181454
R9139 GND.n256 GND.n255 0.00181454
R9140 GND.n7637 GND.n7636 0.00181454
R9141 GND.n7636 GND.n7635 0.00181454
R9142 GND.n4952 GND 0.00175333
R9143 GND GND.n4973 0.00175333
R9144 GND GND.n2346 0.00175333
R9145 GND GND.n150 0.00175333
R9146 GND GND.n5330 0.00175333
R9147 GND.n5337 GND 0.00175333
R9148 GND.n5313 GND 0.00175333
R9149 GND GND.n5310 0.00175333
R9150 GND.n3895 GND 0.00175333
R9151 GND.n3568 GND 0.00175333
R9152 GND.n3411 GND 0.00175333
R9153 GND GND.n2185 0.00175333
R9154 GND GND.n2500 0.00175333
R9155 GND GND.n2815 0.00175333
R9156 GND GND.n3144 0.00175333
R9157 GND GND.n3402 0.00175333
R9158 GND.n6486 GND.n6480 0.00175
R9159 GND.n6490 GND.n6489 0.00175
R9160 GND.n6492 GND.n6478 0.00175
R9161 GND.n6396 GND.n6390 0.00175
R9162 GND.n6400 GND.n6399 0.00175
R9163 GND.n6402 GND.n6388 0.00175
R9164 GND.n2659 GND.n2658 0.00174202
R9165 GND.n3392 GND.n3390 0.00174202
R9166 GND.n4581 GND.n4580 0.00172549
R9167 GND.n3229 GND.n3227 0.001708
R9168 GND.n3998 GND.n3996 0.001708
R9169 GND.n3886 GND.n3884 0.001708
R9170 GND.n3559 GND.n3557 0.001708
R9171 GND.n2018 GND.n2016 0.001708
R9172 GND.n2116 GND.n2107 0.001708
R9173 GND.n2486 GND.n2484 0.001708
R9174 GND.n2780 GND.n2778 0.001708
R9175 GND.n4734 GND.n4732 0.001708
R9176 GND.n772 GND.n770 0.00169681
R9177 GND.n6117 GND 0.00169681
R9178 GND.n7808 GND 0.00169681
R9179 GND.n1441 GND.n1439 0.00166525
R9180 GND.n3331 GND.n3328 0.00163636
R9181 GND.n7518 GND.n7515 0.00163636
R9182 GND.n7580 GND.n7577 0.00163636
R9183 GND.n2634 GND.n2631 0.00163636
R9184 GND.n3060 GND.n3057 0.00163636
R9185 GND.n6975 GND.n6974 0.00163636
R9186 GND.n6821 GND.n6820 0.00163636
R9187 GND.n7755 GND.n7754 0.00163636
R9188 GND.n5637 GND.n5636 0.00163636
R9189 GND.n5453 GND.n5452 0.00163636
R9190 GND.n7456 GND.n7453 0.00163636
R9191 GND.n5121 GND.n5118 0.00163636
R9192 GND.n3721 GND.n3718 0.00163636
R9193 GND.n5510 GND.n5509 0.00163636
R9194 GND.n6509 GND.n6506 0.00163636
R9195 GND.n7087 GND.n7084 0.00163636
R9196 GND.n3241 GND.n3239 0.00154167
R9197 GND.n7544 GND.n7542 0.00154167
R9198 GND.n7606 GND.n7604 0.00154167
R9199 GND.n2505 GND.n2503 0.00154167
R9200 GND.n2922 GND.n2920 0.00154167
R9201 GND.n6944 GND.n6942 0.00154167
R9202 GND.n6781 GND.n6779 0.00154167
R9203 GND.n70 GND.n68 0.00154167
R9204 GND.n1014 GND.n1012 0.00154167
R9205 GND.n1243 GND.n1241 0.00154167
R9206 GND.n7482 GND.n7480 0.00154167
R9207 GND.n4981 GND.n4979 0.00154167
R9208 GND.n3587 GND.n3585 0.00154167
R9209 GND.n1113 GND.n1111 0.00154167
R9210 GND.n6535 GND.n6533 0.00154167
R9211 GND.n7113 GND.n7111 0.00154167
R9212 GND.n3234 GND.n3233 0.00150729
R9213 GND.n2893 GND.n2892 0.00150729
R9214 GND.n2337 GND.n2336 0.00150729
R9215 GND.n7740 GND.n7739 0.00150729
R9216 GND.n1596 GND.n1595 0.00150729
R9217 GND.n5436 GND.n5435 0.00150729
R9218 GND.n4003 GND.n4002 0.00150729
R9219 GND.n5301 GND.n5300 0.00150729
R9220 GND.n3891 GND.n3890 0.00150729
R9221 GND.n3564 GND.n3563 0.00150729
R9222 GND.n2023 GND.n2022 0.00150729
R9223 GND.n2121 GND.n2120 0.00150729
R9224 GND.n2491 GND.n2490 0.00150729
R9225 GND.n4948 GND.n4947 0.00150729
R9226 GND.n4851 GND.n4849 0.00150234
R9227 GND.n4644 GND.n4642 0.00150234
R9228 GND.n2235 GND.n2233 0.00150234
R9229 GND.n2173 GND.n2171 0.00150234
R9230 GND.n145 GND.n143 0.00150234
R9231 GND.n1496 GND.n1494 0.00150234
R9232 GND.n1328 GND.n1326 0.00150234
R9233 GND.n5194 GND.n5192 0.00150234
R9234 GND.n3793 GND.n3791 0.00150234
R9235 GND.n3471 GND.n3469 0.00150234
R9236 GND.n1922 GND.n1920 0.00150234
R9237 GND.n2398 GND.n2396 0.00150234
R9238 GND.n7438 GND.n7437 0.00150166
R9239 GND.n4852 GND.n4851 0.00150164
R9240 GND.n4645 GND.n4644 0.00150164
R9241 GND.n2236 GND.n2235 0.00150164
R9242 GND.n2174 GND.n2173 0.00150164
R9243 GND.n146 GND.n145 0.00150164
R9244 GND.n1497 GND.n1496 0.00150164
R9245 GND.n1329 GND.n1328 0.00150164
R9246 GND.n5195 GND.n5194 0.00150164
R9247 GND.n3794 GND.n3793 0.00150164
R9248 GND.n3472 GND.n3471 0.00150164
R9249 GND.n1923 GND.n1922 0.00150164
R9250 GND.n2399 GND.n2398 0.00150164
R9251 GND.n6456 GND.n666 0.00150121
R9252 GND.n5828 GND.n5687 0.00148684
R9253 GND.n4670 GND.n4651 0.00139286
R9254 GND.n3207 GND.n3203 0.00139286
R9255 GND.n2254 GND.n2252 0.00139286
R9256 GND.n7667 GND.n152 0.00139286
R9257 GND.n1514 GND.n1512 0.00139286
R9258 GND.n5351 GND.n5349 0.00139286
R9259 GND.n3920 GND.n3918 0.00139286
R9260 GND.n5212 GND.n5210 0.00139286
R9261 GND.n3812 GND.n3810 0.00139286
R9262 GND.n3489 GND.n3487 0.00139286
R9263 GND.n1941 GND.n1939 0.00139286
R9264 GND.n2051 GND.n2033 0.00139286
R9265 GND.n2416 GND.n2414 0.00139286
R9266 GND.n2725 GND.n2723 0.00139286
R9267 GND.n4870 GND.n4868 0.00139286
R9268 GND.n2835 GND.n2833 0.00139286
R9269 GND.n4668 GND.n4667 0.00138653
R9270 GND.n3214 GND.n3208 0.00138653
R9271 GND.n2261 GND.n2255 0.00138653
R9272 GND.n7665 GND.n7664 0.00138653
R9273 GND.n1521 GND.n1515 0.00138653
R9274 GND.n5358 GND.n5352 0.00138653
R9275 GND.n3927 GND.n3921 0.00138653
R9276 GND.n5219 GND.n5213 0.00138653
R9277 GND.n3819 GND.n3813 0.00138653
R9278 GND.n3496 GND.n3490 0.00138653
R9279 GND.n1948 GND.n1942 0.00138653
R9280 GND.n2049 GND.n2048 0.00138653
R9281 GND.n2423 GND.n2417 0.00138653
R9282 GND.n2732 GND.n2726 0.00138653
R9283 GND.n4877 GND.n4871 0.00138653
R9284 GND.n2842 GND.n2836 0.00138653
R9285 GND.n4959 GND.n4956 0.00132676
R9286 GND.n3397 GND.n1848 0.0013267
R9287 GND.n3139 GND.n1851 0.0013267
R9288 GND.n2810 GND.n1854 0.0013267
R9289 GND.n2495 GND.n1857 0.0013267
R9290 GND.n2341 GND.n1860 0.0013267
R9291 GND.n2180 GND.n1863 0.0013267
R9292 GND.n1871 GND.n1868 0.0013267
R9293 GND.n3418 GND.n3415 0.0013267
R9294 GND.n5325 GND.n5324 0.0013267
R9295 GND.n3575 GND.n3572 0.0013267
R9296 GND.n3581 GND.n3578 0.0013267
R9297 GND.n3902 GND.n3899 0.0013267
R9298 GND.n5305 GND.n3905 0.0013267
R9299 GND.n5320 GND.n5317 0.0013267
R9300 GND.n4968 GND.n4967 0.0013267
R9301 GND.n3273 GND.t1422 0.00131092
R9302 GND.n3274 GND.n3273 0.00131092
R9303 GND.n2956 GND.n2955 0.00131092
R9304 GND.t594 GND.n2956 0.00131092
R9305 GND.n2965 GND.t594 0.00131092
R9306 GND.n2966 GND.n2965 0.00131092
R9307 GND.n2533 GND.n2532 0.00131092
R9308 GND.t1044 GND.n2533 0.00131092
R9309 GND.n2541 GND.t1044 0.00131092
R9310 GND.n2542 GND.n2541 0.00131092
R9311 GND.n7138 GND.n7137 0.00131092
R9312 GND.t423 GND.n7138 0.00131092
R9313 GND.n7146 GND.t423 0.00131092
R9314 GND.n7147 GND.n7146 0.00131092
R9315 GND.n7071 GND.n7070 0.00131092
R9316 GND.n7070 GND.t1158 0.00131092
R9317 GND.t1158 GND.n7069 0.00131092
R9318 GND.n7069 GND.n7068 0.00131092
R9319 GND.n6917 GND.n6916 0.00131092
R9320 GND.n6916 GND.t622 0.00131092
R9321 GND.t622 GND.n6915 0.00131092
R9322 GND.n6915 GND.n6914 0.00131092
R9323 GND.n6763 GND.n6762 0.00131092
R9324 GND.n6762 GND.t404 0.00131092
R9325 GND.t404 GND.n6761 0.00131092
R9326 GND.n6761 GND.n6760 0.00131092
R9327 GND.n6563 GND.n6562 0.00131092
R9328 GND.n6562 GND.t1404 0.00131092
R9329 GND.t1404 GND.n6561 0.00131092
R9330 GND.n6561 GND.n6560 0.00131092
R9331 GND.n5607 GND.n5606 0.00131092
R9332 GND.t1060 GND.n5607 0.00131092
R9333 GND.n5615 GND.t1060 0.00131092
R9334 GND.n5616 GND.n5615 0.00131092
R9335 GND.n5472 GND.n5471 0.00131092
R9336 GND.t473 GND.n5472 0.00131092
R9337 GND.n5480 GND.t473 0.00131092
R9338 GND.n5481 GND.n5480 0.00131092
R9339 GND.n1145 GND.n1144 0.00131092
R9340 GND.n1144 GND.t635 0.00131092
R9341 GND.t635 GND.n1143 0.00131092
R9342 GND.n1143 GND.n1142 0.00131092
R9343 GND.n3621 GND.n3620 0.00131092
R9344 GND.t1154 GND.n3621 0.00131092
R9345 GND.n3629 GND.t1154 0.00131092
R9346 GND.n3630 GND.n3629 0.00131092
R9347 GND.n5015 GND.n5014 0.00131092
R9348 GND.t10 GND.n5015 0.00131092
R9349 GND.n5023 GND.t10 0.00131092
R9350 GND.n5024 GND.n5023 0.00131092
R9351 GND.n410 GND.n409 0.00131092
R9352 GND.t547 GND.n410 0.00131092
R9353 GND.n418 GND.t547 0.00131092
R9354 GND.n419 GND.n418 0.00131092
R9355 GND.n325 GND.n324 0.00131092
R9356 GND.n324 GND.t434 0.00131092
R9357 GND.t434 GND.n323 0.00131092
R9358 GND.n323 GND.n322 0.00131092
R9359 GND.n223 GND.n222 0.00131092
R9360 GND.n222 GND.t688 0.00131092
R9361 GND.t688 GND.n221 0.00131092
R9362 GND.n221 GND.n220 0.00131092
R9363 GND.n194 GND.n193 0.00131092
R9364 GND.n193 GND.t610 0.00131092
R9365 GND.n4463 GND.n4462 0.00125043
R9366 GND.n1439 GND 0.00124153
R9367 GND.n5744 GND.n5743 0.00122464
R9368 GND.n991 GND 0.00116489
R9369 GND.n5875 GND.n5860 0.00116489
R9370 GND.n7246 GND.n7232 0.00116489
R9371 GND.n7444 GND.n7442 0.00115206
R9372 GND.n7444 GND.n7443 0.00115206
R9373 GND.n4591 GND.n4474 0.00114322
R9374 GND.n6461 GND.n6460 0.00109111
R9375 GND.n6494 GND.n6477 0.00108327
R9376 GND.n6404 GND.n6387 0.00108327
R9377 GND.n6460 GND.n6459 0.00107707
R9378 GND.n7442 GND.n7441 0.00107707
R9379 GND.n6378 GND.n6377 0.00107231
R9380 GND.n7803 GND.n7801 0.00107231
R9381 GND.n4901 GND.n4900 0.00103916
R9382 GND.n4700 GND.n4699 0.00103916
R9383 GND.n3156 GND.n3155 0.00103916
R9384 GND.n2824 GND.n2823 0.00103916
R9385 GND.n2285 GND.n2284 0.00103916
R9386 GND.n7689 GND.n7688 0.00103916
R9387 GND.n1545 GND.n1544 0.00103916
R9388 GND.n5382 GND.n5381 0.00103916
R9389 GND.n3951 GND.n3950 0.00103916
R9390 GND.n5243 GND.n5242 0.00103916
R9391 GND.n3843 GND.n3842 0.00103916
R9392 GND.n3520 GND.n3519 0.00103916
R9393 GND.n1972 GND.n1971 0.00103916
R9394 GND.n2059 GND.n2058 0.00103916
R9395 GND.n2447 GND.n2446 0.00103916
R9396 GND.n2756 GND.n2755 0.00103916
R9397 GND.n4462 GND.n4459 0.00103602
R9398 GND.n4766 GND.n4765 0.00102722
R9399 GND.n2807 GND.n2806 0.00102722
R9400 GND.n4950 GND.n4949 0.00101312
R9401 GND.n3236 GND.n3235 0.00101312
R9402 GND.n2339 GND.n2338 0.00101312
R9403 GND.n2123 GND.n2122 0.00101312
R9404 GND.n7742 GND.n7741 0.00101312
R9405 GND.n1598 GND.n1597 0.00101312
R9406 GND.n5438 GND.n5437 0.00101312
R9407 GND.n4005 GND.n4004 0.00101312
R9408 GND.n5303 GND.n5302 0.00101312
R9409 GND.n3893 GND.n3892 0.00101312
R9410 GND.n3566 GND.n3565 0.00101312
R9411 GND.n2025 GND.n2024 0.00101312
R9412 GND.n2493 GND.n2492 0.00101312
R9413 GND.n2917 GND.n2916 0.00101312
R9414 GND.n4738 GND.n4737 0.00100729
R9415 GND.n2916 GND.n2915 0.00100714
R9416 GND.n4949 GND.n4925 0.00100714
R9417 GND.n3235 GND.n3180 0.00100714
R9418 GND.n2338 GND.n2309 0.00100714
R9419 GND.n2122 GND.n2087 0.00100714
R9420 GND.n7741 GND.n7713 0.00100714
R9421 GND.n1597 GND.n1569 0.00100714
R9422 GND.n5437 GND.n5406 0.00100714
R9423 GND.n4004 GND.n3975 0.00100714
R9424 GND.n5302 GND.n5267 0.00100714
R9425 GND.n3892 GND.n3867 0.00100714
R9426 GND.n3565 GND.n3544 0.00100714
R9427 GND.n2024 GND.n1996 0.00100714
R9428 GND.n2492 GND.n2471 0.00100714
R9429 GND.n1378 GND.n1377 0.00100417
R9430 GND.n2709 GND.n2708 0.001004
R9431 GND.n3135 GND.n3132 0.001004
R9432 GND.n4058 GND.n4055 0.001004
R9433 GND.n1351 GND.n1350 0.00100271
R9434 GND.n7795 GND.n7794 0.00100171
R9435 GND.n6470 GND.n6469 0.00100171
R9436 GND.n6329 GND.n6328 0.00100171
R9437 GND.n6410 GND.n6409 0.00100171
R9438 GND.n7794 GND.n7793 0.00100166
R9439 GND.n6470 GND.n705 0.00100166
R9440 GND.n6329 GND.n6326 0.00100166
R9441 GND.n6409 GND.n6269 0.00100166
R9442 GND.n1430 GND.n1374 0.00100126
R9443 GND.n7378 GND.n7377 0.00100097
R9444 GND.n5914 GND.n5913 0.00100097
R9445 GND.n6045 GND.n6003 0.00100097
R9446 GND.n7285 GND.n7284 0.00100097
R9447 GND.n5666 GND.n5659 0.00100097
R9448 GND.n5796 GND.n5688 0.00100097
R9449 GND.n5755 GND.n5754 0.00100097
R9450 GND.n3257 GND.n3256 0.00100095
R9451 GND.n7560 GND.n7559 0.00100095
R9452 GND.n7622 GND.n7621 0.00100095
R9453 GND.n2521 GND.n2520 0.00100095
R9454 GND.n2938 GND.n2937 0.00100095
R9455 GND.n6960 GND.n6959 0.00100095
R9456 GND.n6797 GND.n6796 0.00100095
R9457 GND.n86 GND.n85 0.00100095
R9458 GND.n1030 GND.n1029 0.00100095
R9459 GND.n1259 GND.n1258 0.00100095
R9460 GND.n7498 GND.n7497 0.00100095
R9461 GND.n4997 GND.n4996 0.00100095
R9462 GND.n3603 GND.n3602 0.00100095
R9463 GND.n1129 GND.n1128 0.00100095
R9464 GND.n6551 GND.n6550 0.00100095
R9465 GND.n7129 GND.n7128 0.00100095
R9466 GND.n6458 GND.n6422 0.00100086
R9467 GND.n7440 GND.n507 0.00100086
R9468 GND.n4855 GND.n4854 0.00100064
R9469 GND.n4648 GND.n4647 0.00100064
R9470 GND.n2239 GND.n2238 0.00100064
R9471 GND.n2177 GND.n2176 0.00100064
R9472 GND.n149 GND.n148 0.00100064
R9473 GND.n1499 GND.n1498 0.00100064
R9474 GND.n5197 GND.n5196 0.00100064
R9475 GND.n3797 GND.n3796 0.00100064
R9476 GND.n1926 GND.n1925 0.00100064
R9477 GND.n5321 GND.n1844 0.00100018
R9478 GND.n5321 GND.n1839 0.00100018
R9479 GND.n5321 GND.n1834 0.00100018
R9480 GND.n5321 GND.n1829 0.00100018
R9481 GND.n5321 GND.n1824 0.00100018
R9482 GND.n5321 GND.n1819 0.00100018
R9483 GND.n5321 GND.n1814 0.00100018
R9484 GND.n5321 GND.n1809 0.00100018
R9485 GND.n5321 GND.n1804 0.00100018
R9486 GND.n5321 GND.n1799 0.00100018
R9487 GND.n5321 GND.n1794 0.00100018
R9488 GND.n5321 GND.n1789 0.00100018
R9489 GND.n5321 GND.n1784 0.00100018
R9490 GND.n5321 GND.n1779 0.00100018
R9491 GND.n4964 GND.n4800 0.00100018
R9492 GND.n7441 GND.n7440 0.00100017
R9493 GND.n6459 GND.n6458 0.00100017
R9494 GND.n5321 GND.n1848 0.00100006
R9495 GND.n5321 GND.n1851 0.00100006
R9496 GND.n5321 GND.n1854 0.00100006
R9497 GND.n5321 GND.n1857 0.00100006
R9498 GND.n5321 GND.n1860 0.00100006
R9499 GND.n5321 GND.n1863 0.00100006
R9500 GND.n5321 GND.n1871 0.00100006
R9501 GND.n5321 GND.n3418 0.00100006
R9502 GND.n5324 GND.n5321 0.00100006
R9503 GND.n5321 GND.n3575 0.00100006
R9504 GND.n5321 GND.n3581 0.00100006
R9505 GND.n5321 GND.n3902 0.00100006
R9506 GND.n5321 GND.n3905 0.00100006
R9507 GND.n5321 GND.n5320 0.00100006
R9508 GND.n4967 GND.n4964 0.00100006
R9509 GND.n4464 GND.n4458 0.00100003
R9510 GND.n3135 GND.n3134 0.00100001
R9511 GND.n3392 GND.n3391 0.00100001
R9512 GND.n4058 GND.n4057 0.00100001
R9513 GND.n4964 GND.n4959 0.001
R9514 GND.n6499 GND.n6498 0.001
R9515 GND.n7445 GND.n7444 0.001
R9516 GND.n6295 GND.n6294 0.001
R9517 GND.n4472 GND.n4471 0.000966399
R9518 GND.n4471 GND.n4470 0.000959101
R9519 GND.n4470 GND.n4469 0.000959101
R9520 GND.n4668 GND.n4657 0.000943262
R9521 GND.n3208 GND.n3201 0.000943262
R9522 GND.n2255 GND.n2250 0.000943262
R9523 GND.n7665 GND.n158 0.000943262
R9524 GND.n1515 GND.n1510 0.000943262
R9525 GND.n5352 GND.n5347 0.000943262
R9526 GND.n3921 GND.n3916 0.000943262
R9527 GND.n5213 GND.n5208 0.000943262
R9528 GND.n3813 GND.n3808 0.000943262
R9529 GND.n3490 GND.n3485 0.000943262
R9530 GND.n1942 GND.n1937 0.000943262
R9531 GND.n2049 GND.n2039 0.000943262
R9532 GND.n2417 GND.n2412 0.000943262
R9533 GND.n2726 GND.n2721 0.000943262
R9534 GND.n4871 GND.n4866 0.000943262
R9535 GND.n2836 GND.n2831 0.000943262
R9536 GND.n858 GND.n856 0.000898936
R9537 GND.n874 GND.n710 0.000898936
R9538 GND.n4093 GND.n4092 0.000864406
R9539 GND.n4099 GND.n4098 0.000864406
R9540 GND.n4094 GND.n4093 0.000858717
R9541 GND.n4096 GND.n4094 0.000858717
R9542 GND.n4098 GND.n4097 0.000858717
R9543 GND.n4097 GND.n4096 0.000858717
R9544 GND.n4569 GND.n4568 0.000858717
R9545 GND.n4570 GND.n4569 0.000858717
R9546 GND.n4572 GND.n4571 0.000858717
R9547 GND.n4571 GND.n4570 0.000858717
R9548 GND.n1380 GND.n1379 0.000840211
R9549 GND.n1430 GND.n1380 0.000840211
R9550 GND.n3398 GND.n3397 0.000826763
R9551 GND.n3140 GND.n3139 0.000826763
R9552 GND.n2811 GND.n2810 0.000826763
R9553 GND.n2496 GND.n2495 0.000826763
R9554 GND.n2342 GND.n2341 0.000826763
R9555 GND.n2181 GND.n2180 0.000826763
R9556 GND.n1868 GND.n1867 0.000826763
R9557 GND.n3415 GND.n3414 0.000826763
R9558 GND.n5326 GND.n5325 0.000826763
R9559 GND.n3572 GND.n3571 0.000826763
R9560 GND.n3578 GND.n3577 0.000826763
R9561 GND.n3899 GND.n3898 0.000826763
R9562 GND.n5306 GND.n5305 0.000826763
R9563 GND.n5317 GND.n5316 0.000826763
R9564 GND.n4969 GND.n4968 0.000826763
R9565 GND.n4956 GND.n4955 0.000826763
R9566 GND.n1352 GND.n1351 0.000801918
R9567 GND.n1353 GND.n1352 0.000801918
R9568 GND.n1429 GND.n1428 0.000801918
R9569 GND.n1430 GND.n1429 0.000801918
R9570 GND.n1423 GND.n1422 0.000801918
R9571 GND.n1430 GND.n1423 0.000801918
R9572 GND.n1415 GND.n1414 0.000801918
R9573 GND.n1430 GND.n1415 0.000801918
R9574 GND.n1412 GND.n1411 0.000801918
R9575 GND.n1430 GND.n1412 0.000801918
R9576 GND.n1355 GND.n1354 0.000801918
R9577 GND.n1354 GND.n1353 0.000801918
R9578 GND.n1360 GND.n1359 0.000801918
R9579 GND.n1409 GND.n1408 0.000801918
R9580 GND.n1430 GND.n1409 0.000801918
R9581 GND.n1438 GND.n1437 0.000801918
R9582 GND.n1432 GND.n1431 0.000801918
R9583 GND.n1431 GND.n1430 0.000801918
R9584 GND.n1405 GND.n1404 0.000801918
R9585 GND.n1430 GND.n1405 0.000801918
R9586 GND.n1353 GND.n1348 0.000801918
R9587 GND.n1398 GND.n1397 0.000801918
R9588 GND.n1430 GND.n1398 0.000801918
R9589 GND.n1390 GND.n1389 0.000801918
R9590 GND.n1430 GND.n1390 0.000801918
R9591 GND.n1345 GND.n1344 0.000801918
R9592 GND.n1353 GND.n1345 0.000801918
R9593 GND.n1368 GND.n1367 0.000801918
R9594 GND.n1430 GND.n1368 0.000801918
R9595 GND.n4741 GND.n4740 0.000756235
R9596 GND.n4740 GND.n4739 0.000756235
R9597 GND.n3161 GND.n3160 0.000756235
R9598 GND.n3160 GND.n3159 0.000756235
R9599 GND.n2896 GND.n2895 0.000756235
R9600 GND.n2895 GND.n2894 0.000756235
R9601 GND.n2290 GND.n2289 0.000756235
R9602 GND.n2289 GND.n2288 0.000756235
R9603 GND.n7694 GND.n7693 0.000756235
R9604 GND.n7693 GND.n7692 0.000756235
R9605 GND.n1550 GND.n1549 0.000756235
R9606 GND.n1549 GND.n1548 0.000756235
R9607 GND.n5387 GND.n5386 0.000756235
R9608 GND.n5386 GND.n5385 0.000756235
R9609 GND.n5248 GND.n5247 0.000756235
R9610 GND.n5247 GND.n5246 0.000756235
R9611 GND.n3848 GND.n3847 0.000756235
R9612 GND.n3847 GND.n3846 0.000756235
R9613 GND.n3525 GND.n3524 0.000756235
R9614 GND.n3524 GND.n3523 0.000756235
R9615 GND.n1977 GND.n1976 0.000756235
R9616 GND.n1976 GND.n1975 0.000756235
R9617 GND.n2111 GND.n2110 0.000756235
R9618 GND.n2112 GND.n2111 0.000756235
R9619 GND.n2452 GND.n2451 0.000756235
R9620 GND.n2451 GND.n2450 0.000756235
R9621 GND.n2787 GND.n2786 0.000756235
R9622 GND.n2786 GND.n2785 0.000756235
R9623 GND.n4906 GND.n4905 0.000756235
R9624 GND.n4905 GND.n4904 0.000756235
R9625 GND.n3956 GND.n3955 0.000756235
R9626 GND.n3955 GND.n3954 0.000756235
R9627 GND.n4472 GND.n4466 0.000714408
R9628 GND.n726 GND.n724 0.000632979
R9629 GND.n6135 GND.n5852 0.000632979
R9630 GND.n7434 GND.n544 0.000632979
R9631 GND.n4466 GND.n4464 0.000607204
R9632 GND.n4452 GND.n4451 0.000567786
R9633 GND.n6326 GND.n6296 0.000560793
R9634 GND.n705 GND.n667 0.000560793
R9635 GND.n7793 GND.n7763 0.000560793
R9636 GND.n6411 GND.n6410 0.000557763
R9637 GND.n6328 GND.n6327 0.000557763
R9638 GND.n6469 GND.n6468 0.000557763
R9639 GND.n7796 GND.n7795 0.000557763
R9640 GND.n4075 GND.n4074 0.000557678
R9641 GND.n3333 GND.n3332 0.000544755
R9642 GND.n7520 GND.n7519 0.000544755
R9643 GND.n7582 GND.n7581 0.000544755
R9644 GND.n2636 GND.n2635 0.000544755
R9645 GND.n3062 GND.n3061 0.000544755
R9646 GND.n6973 GND.n6972 0.000544755
R9647 GND.n6819 GND.n6818 0.000544755
R9648 GND.n7753 GND.n7752 0.000544755
R9649 GND.n5635 GND.n5634 0.000544755
R9650 GND.n5451 GND.n5450 0.000544755
R9651 GND.n7458 GND.n7457 0.000544755
R9652 GND.n5123 GND.n5122 0.000544755
R9653 GND.n3723 GND.n3722 0.000544755
R9654 GND.n5508 GND.n5507 0.000544755
R9655 GND.n6511 GND.n6510 0.000544755
R9656 GND.n7089 GND.n7088 0.000544755
R9657 GND.n4084 GND.n4083 0.000538452
R9658 GND.n4566 GND.n4565 0.000537082
R9659 GND.n3290 GND.n3289 0.000530553
R9660 GND.n2982 GND.n2981 0.000530553
R9661 GND.n2556 GND.n2555 0.000530553
R9662 GND.n7156 GND.n7155 0.000530553
R9663 GND.n6993 GND.n6992 0.000530553
R9664 GND.n6839 GND.n6838 0.000530553
R9665 GND.n6685 GND.n6684 0.000530553
R9666 GND.n6614 GND.n6613 0.000530553
R9667 GND.n5566 GND.n5565 0.000530553
R9668 GND.n1064 GND.n1063 0.000530553
R9669 GND.n1185 GND.n1184 0.000530553
R9670 GND.n3646 GND.n3645 0.000530553
R9671 GND.n5043 GND.n5042 0.000530553
R9672 GND.n438 GND.n437 0.000530553
R9673 GND.n369 GND.n368 0.000530553
R9674 GND.n265 GND.n264 0.000530553
R9675 GND.n6384 GND.n6383 0.000528881
R9676 GND.n6383 GND.n6382 0.000528881
R9677 GND.n6386 GND.n6385 0.000528881
R9678 GND.n6474 GND.n6473 0.000528881
R9679 GND.n6473 GND.n6472 0.000528881
R9680 GND.n6476 GND.n6475 0.000528881
R9681 GND.n3311 GND.n3310 0.00052846
R9682 GND.n3008 GND.n3007 0.00052846
R9683 GND.n2582 GND.n2581 0.00052846
R9684 GND.n7182 GND.n7181 0.00052846
R9685 GND.n7019 GND.n7018 0.00052846
R9686 GND.n6865 GND.n6864 0.00052846
R9687 GND.n6711 GND.n6710 0.00052846
R9688 GND.n6640 GND.n6639 0.00052846
R9689 GND.n5592 GND.n5591 0.00052846
R9690 GND.n1090 GND.n1089 0.00052846
R9691 GND.n1211 GND.n1210 0.00052846
R9692 GND.n3672 GND.n3671 0.00052846
R9693 GND.n5069 GND.n5068 0.00052846
R9694 GND.n464 GND.n463 0.00052846
R9695 GND.n395 GND.n394 0.00052846
R9696 GND.n291 GND.n290 0.00052846
R9697 GND.n241 GND.n240 0.00052846
R9698 GND.n7648 GND.n7647 0.00052846
R9699 GND.n7208 GND.n7207 0.00052846
R9700 GND.n2604 GND.n2603 0.00052846
R9701 GND.n6896 GND.n6895 0.00052846
R9702 GND.n6742 GND.n6741 0.00052846
R9703 GND.n6583 GND.n6582 0.00052846
R9704 GND.n1040 GND.n1039 0.00052846
R9705 GND.n3691 GND.n3690 0.00052846
R9706 GND.n345 GND.n344 0.00052846
R9707 GND.n483 GND.n482 0.00052846
R9708 GND.n5091 GND.n5090 0.00052846
R9709 GND.n1163 GND.n1162 0.00052846
R9710 GND.n5535 GND.n5534 0.00052846
R9711 GND.n7050 GND.n7049 0.00052846
R9712 GND.n3030 GND.n3029 0.00052846
R9713 GND.n4103 GND.n4102 0.000526656
R9714 GND.n3038 GND.n3037 0.0005264
R9715 GND.n298 GND.n297 0.0005264
R9716 GND.n7656 GND.n7655 0.0005264
R9717 GND.n7216 GND.n7215 0.0005264
R9718 GND.n2612 GND.n2611 0.0005264
R9719 GND.n6904 GND.n6903 0.0005264
R9720 GND.n6750 GND.n6749 0.0005264
R9721 GND.n6647 GND.n6646 0.0005264
R9722 GND.n1097 GND.n1096 0.0005264
R9723 GND.n3699 GND.n3698 0.0005264
R9724 GND.n402 GND.n401 0.0005264
R9725 GND.n491 GND.n490 0.0005264
R9726 GND.n5099 GND.n5098 0.0005264
R9727 GND.n1218 GND.n1217 0.0005264
R9728 GND.n5599 GND.n5598 0.0005264
R9729 GND.n7058 GND.n7057 0.0005264
R9730 GND.n4454 GND.n4453 0.000525991
R9731 GND.n4480 GND.n4479 0.000524722
R9732 GND.n4587 GND.n4586 0.000523819
R9733 GND.n4591 GND.n4590 0.000523819
R9734 GND.n4582 GND.n4581 0.000523819
R9735 GND.t657 GND.n4588 0.000523446
R9736 GND.n4590 GND.n4589 0.000523446
R9737 GND.n4589 GND.t657 0.000523446
R9738 GND.n4588 GND.n4587 0.000523446
R9739 GND.n4583 GND.n4582 0.000523446
R9740 GND.t657 GND.n4583 0.000523446
R9741 GND.n4558 GND.n4557 0.000517138
R9742 GND.n231 GND.n230 0.000512627
R9743 GND.n7638 GND.n7637 0.000512627
R9744 GND.n7198 GND.n7190 0.000512627
R9745 GND.n2594 GND.n2588 0.000512627
R9746 GND.n6886 GND.n6873 0.000512627
R9747 GND.n6732 GND.n6719 0.000512627
R9748 GND.n6573 GND.n6570 0.000512627
R9749 GND.n5548 GND.n5547 0.000512627
R9750 GND.n3681 GND.n3678 0.000512627
R9751 GND.n335 GND.n332 0.000512627
R9752 GND.n473 GND.n470 0.000512627
R9753 GND.n5081 GND.n5075 0.000512627
R9754 GND.n1153 GND.n1152 0.000512627
R9755 GND.n6596 GND.n6595 0.000512627
R9756 GND.n7040 GND.n7027 0.000512627
R9757 GND.n3020 GND.n3019 0.000512627
R9758 GND.n3284 GND.n3283 0.000512369
R9759 GND.n2976 GND.n2975 0.000512369
R9760 GND.n2550 GND.n2549 0.000512369
R9761 GND.n7029 GND.n7028 0.000512369
R9762 GND.n6875 GND.n6874 0.000512369
R9763 GND.n6721 GND.n6720 0.000512369
R9764 GND.n6679 GND.n6678 0.000512369
R9765 GND.n6608 GND.n6607 0.000512369
R9766 GND.n5560 GND.n5559 0.000512369
R9767 GND.n1058 GND.n1057 0.000512369
R9768 GND.n1179 GND.n1178 0.000512369
R9769 GND.n3640 GND.n3639 0.000512369
R9770 GND.n5037 GND.n5036 0.000512369
R9771 GND.n432 GND.n431 0.000512369
R9772 GND.n363 GND.n362 0.000512369
R9773 GND.n259 GND.n258 0.000512369
R9774 GND.n1389 GND.n1388 0.000508571
R9775 GND.n1397 GND.n1396 0.000508571
R9776 GND.n1404 GND.n1403 0.000508571
R9777 GND.n1433 GND.n1432 0.000508571
R9778 GND.n1439 GND.n1438 0.000508571
R9779 GND.n1408 GND.n1364 0.000508571
R9780 GND.n1361 GND.n1360 0.000508571
R9781 GND.n1414 GND.n1413 0.000508571
R9782 GND.n1422 GND.n1421 0.000508571
R9783 GND.n1428 GND.n1427 0.000508571
R9784 GND.n1367 GND.n1366 0.000508571
R9785 GND.n2955 GND.n2954 0.000507826
R9786 GND.n2532 GND.n2531 0.000507826
R9787 GND.n7137 GND.n7136 0.000507826
R9788 GND.n7072 GND.n7071 0.000507826
R9789 GND.n6918 GND.n6917 0.000507826
R9790 GND.n6764 GND.n6763 0.000507826
R9791 GND.n6564 GND.n6563 0.000507826
R9792 GND.n5606 GND.n5605 0.000507826
R9793 GND.n5471 GND.n5470 0.000507826
R9794 GND.n1146 GND.n1145 0.000507826
R9795 GND.n3620 GND.n3619 0.000507826
R9796 GND.n5014 GND.n5013 0.000507826
R9797 GND.n409 GND.n408 0.000507826
R9798 GND.n326 GND.n325 0.000507826
R9799 GND.n224 GND.n223 0.000507826
R9800 GND.n195 GND.n194 0.000507826
R9801 GND.n3275 GND.n3274 0.000507826
R9802 GND.n2967 GND.n2966 0.000507826
R9803 GND.n2543 GND.n2542 0.000507826
R9804 GND.n7148 GND.n7147 0.000507826
R9805 GND.n7068 GND.n7067 0.000507826
R9806 GND.n6914 GND.n6913 0.000507826
R9807 GND.n6760 GND.n6759 0.000507826
R9808 GND.n6560 GND.n6559 0.000507826
R9809 GND.n5617 GND.n5616 0.000507826
R9810 GND.n5482 GND.n5481 0.000507826
R9811 GND.n1142 GND.n1141 0.000507826
R9812 GND.n3631 GND.n3630 0.000507826
R9813 GND.n5025 GND.n5024 0.000507826
R9814 GND.n420 GND.n419 0.000507826
R9815 GND.n322 GND.n321 0.000507826
R9816 GND.n220 GND.n219 0.000507826
R9817 GND.n2784 GND.n2783 0.000507291
R9818 GND.n5915 GND.n5914 0.000506774
R9819 GND.n5917 GND.n5916 0.000506774
R9820 GND.n6120 GND.n6003 0.000506774
R9821 GND.n6119 GND.n6118 0.000506774
R9822 GND.n6122 GND.n6121 0.000506774
R9823 GND.n6002 GND.n6001 0.000506774
R9824 GND.n729 GND.n728 0.000506774
R9825 GND.n823 GND.n822 0.000506774
R9826 GND.n918 GND.n917 0.000506774
R9827 GND.n993 GND.n992 0.000506774
R9828 GND.n916 GND.n915 0.000506774
R9829 GND.n825 GND.n824 0.000506774
R9830 GND.n5696 GND.n5688 0.000506774
R9831 GND.n5756 GND.n5755 0.000506774
R9832 GND.n5659 GND.n5658 0.000506774
R9833 GND.n5695 GND.n5686 0.000506774
R9834 GND.n5758 GND.n5757 0.000506774
R9835 GND.n6229 GND.n6228 0.000506774
R9836 GND.n6163 GND.n6162 0.000506774
R9837 GND.n7288 GND.n7287 0.000506774
R9838 GND.n7377 GND.n7376 0.000506774
R9839 GND.n7807 GND.n7806 0.000506774
R9840 GND.n7375 GND.n547 0.000506774
R9841 GND.n7373 GND.n7372 0.000506774
R9842 GND.n7286 GND.n7285 0.000506774
R9843 GND.n4666 GND.n4665 0.000505544
R9844 GND.n3216 GND.n3215 0.000505544
R9845 GND.n2263 GND.n2262 0.000505544
R9846 GND.n7663 GND.n7662 0.000505544
R9847 GND.n1523 GND.n1522 0.000505544
R9848 GND.n5360 GND.n5359 0.000505544
R9849 GND.n3929 GND.n3928 0.000505544
R9850 GND.n5221 GND.n5220 0.000505544
R9851 GND.n3821 GND.n3820 0.000505544
R9852 GND.n3498 GND.n3497 0.000505544
R9853 GND.n1950 GND.n1949 0.000505544
R9854 GND.n2425 GND.n2424 0.000505544
R9855 GND.n2734 GND.n2733 0.000505544
R9856 GND.n2047 GND.n2046 0.000505544
R9857 GND.n4879 GND.n4878 0.000505544
R9858 GND.n2844 GND.n2843 0.000505544
R9859 GND.n3258 GND.n3257 0.000504863
R9860 GND.n7561 GND.n7560 0.000504863
R9861 GND.n7623 GND.n7622 0.000504863
R9862 GND.n2522 GND.n2521 0.000504863
R9863 GND.n2939 GND.n2938 0.000504863
R9864 GND.n6962 GND.n6960 0.000504863
R9865 GND.n6799 GND.n6797 0.000504863
R9866 GND.n87 GND.n86 0.000504863
R9867 GND.n5624 GND.n1030 0.000504863
R9868 GND.n1277 GND.n1259 0.000504863
R9869 GND.n7499 GND.n7498 0.000504863
R9870 GND.n4998 GND.n4997 0.000504863
R9871 GND.n3604 GND.n3603 0.000504863
R9872 GND.n5489 GND.n1129 0.000504863
R9873 GND.n6552 GND.n6551 0.000504863
R9874 GND.n7130 GND.n7129 0.000504863
R9875 GND.n1400 GND.n1399 0.000504378
R9876 GND.n1393 GND.n1392 0.000504346
R9877 GND.n1356 GND.n1355 0.000504346
R9878 GND.n1426 GND.n1425 0.00050424
R9879 GND.n1418 GND.n1417 0.00050424
R9880 GND.n1358 GND.n1357 0.00050424
R9881 GND.n1363 GND.n1362 0.00050424
R9882 GND.n1435 GND.n1434 0.00050424
R9883 GND.n1395 GND.n1394 0.00050424
R9884 GND.n1382 GND.n1381 0.00050424
R9885 GND.n1384 GND.n1383 0.00050424
R9886 GND.n1336 GND.n1335 0.000504176
R9887 GND.n1420 GND.n1419 0.000504112
R9888 GND.n1339 GND.n1338 0.000504112
R9889 GND.n1443 GND.n1442 0.000504112
R9890 GND.n1402 GND.n1401 0.000504112
R9891 GND.n1387 GND.n1386 0.000504112
R9892 GND.n4853 GND.n4852 0.000504005
R9893 GND.n4646 GND.n4645 0.000504005
R9894 GND.n2660 GND.n2659 0.000504005
R9895 GND.n3134 GND.n3133 0.000504005
R9896 GND.n3393 GND.n3392 0.000504005
R9897 GND.n2237 GND.n2236 0.000504005
R9898 GND.n2175 GND.n2174 0.000504005
R9899 GND.n147 GND.n146 0.000504005
R9900 GND.n1330 GND.n1329 0.000504005
R9901 GND.n4057 GND.n4056 0.000504005
R9902 GND.n3795 GND.n3794 0.000504005
R9903 GND.n3473 GND.n3472 0.000504005
R9904 GND.n1924 GND.n1923 0.000504005
R9905 GND.n2400 GND.n2399 0.000504005
R9906 GND.n4466 GND.n4465 0.00050212
R9907 GND.n4856 GND.n4855 0.000501449
R9908 GND.n4649 GND.n4648 0.000501449
R9909 GND.n2711 GND.n2710 0.000501449
R9910 GND.n3137 GND.n3136 0.000501449
R9911 GND.n2240 GND.n2239 0.000501449
R9912 GND.n2178 GND.n2177 0.000501449
R9913 GND.n7744 GND.n149 0.000501449
R9914 GND.n1500 GND.n1499 0.000501449
R9915 GND.n5440 GND.n1331 0.000501449
R9916 GND.n4060 GND.n4059 0.000501449
R9917 GND.n5198 GND.n5197 0.000501449
R9918 GND.n3798 GND.n3797 0.000501449
R9919 GND.n3475 GND.n3474 0.000501449
R9920 GND.n1927 GND.n1926 0.000501449
R9921 GND.n2402 GND.n2401 0.000501449
R9922 GND.n3395 GND.n3394 0.000501449
R9923 GND.n3350 GND.n3349 0.000501292
R9924 GND.n3349 GND.n3348 0.000501292
R9925 GND.n7537 GND.n7536 0.000501292
R9926 GND.n7536 GND.n7535 0.000501292
R9927 GND.n7599 GND.n7598 0.000501292
R9928 GND.n7598 GND.n7597 0.000501292
R9929 GND.n2653 GND.n2652 0.000501292
R9930 GND.n2652 GND.n2651 0.000501292
R9931 GND.n3079 GND.n3078 0.000501292
R9932 GND.n3078 GND.n3077 0.000501292
R9933 GND.n6971 GND.n6966 0.000501292
R9934 GND.n6971 GND.n6970 0.000501292
R9935 GND.n6817 GND.n6803 0.000501292
R9936 GND.n6817 GND.n6816 0.000501292
R9937 GND.n7749 GND.n7748 0.000501292
R9938 GND.n7750 GND.n7749 0.000501292
R9939 GND.n5633 GND.n5628 0.000501292
R9940 GND.n5633 GND.n5632 0.000501292
R9941 GND.n5449 GND.n5444 0.000501292
R9942 GND.n5449 GND.n5448 0.000501292
R9943 GND.n7475 GND.n7474 0.000501292
R9944 GND.n7474 GND.n7473 0.000501292
R9945 GND.n5140 GND.n5139 0.000501292
R9946 GND.n5139 GND.n5138 0.000501292
R9947 GND.n3740 GND.n3739 0.000501292
R9948 GND.n3739 GND.n3738 0.000501292
R9949 GND.n5506 GND.n5492 0.000501292
R9950 GND.n5506 GND.n5505 0.000501292
R9951 GND.n6528 GND.n6527 0.000501292
R9952 GND.n6527 GND.n6526 0.000501292
R9953 GND.n7106 GND.n7105 0.000501292
R9954 GND.n7105 GND.n7104 0.000501292
R9955 GND.n4568 GND.n4567 0.00050117
R9956 GND.n4573 GND.n4572 0.00050117
R9957 GND.n5918 GND.n5917 0.00050097
R9958 GND.n6118 GND.n6117 0.00050097
R9959 GND.n6123 GND.n6122 0.00050097
R9960 GND.n6001 GND.n6000 0.00050097
R9961 GND.n730 GND.n729 0.00050097
R9962 GND.n822 GND.n821 0.00050097
R9963 GND.n919 GND.n918 0.00050097
R9964 GND.n992 GND.n991 0.00050097
R9965 GND.n915 GND.n914 0.00050097
R9966 GND.n826 GND.n825 0.00050097
R9967 GND.n5759 GND.n5758 0.00050097
R9968 GND.n6228 GND.n6227 0.00050097
R9969 GND.n6164 GND.n6163 0.00050097
R9970 GND.n7289 GND.n7288 0.00050097
R9971 GND.n7808 GND.n7807 0.00050097
R9972 GND.n7422 GND.n547 0.00050097
R9973 GND.n7372 GND.n7371 0.00050097
R9974 GND.n5829 GND.n5686 0.00050097
R9975 GND.n4667 GND.n4666 0.000500915
R9976 GND.n3215 GND.n3214 0.000500915
R9977 GND.n2262 GND.n2261 0.000500915
R9978 GND.n7664 GND.n7663 0.000500915
R9979 GND.n1522 GND.n1521 0.000500915
R9980 GND.n5359 GND.n5358 0.000500915
R9981 GND.n3928 GND.n3927 0.000500915
R9982 GND.n5220 GND.n5219 0.000500915
R9983 GND.n3820 GND.n3819 0.000500915
R9984 GND.n3497 GND.n3496 0.000500915
R9985 GND.n1949 GND.n1948 0.000500915
R9986 GND.n2424 GND.n2423 0.000500915
R9987 GND.n2733 GND.n2732 0.000500915
R9988 GND.n2048 GND.n2047 0.000500915
R9989 GND.n4878 GND.n4877 0.000500915
R9990 GND.n2843 GND.n2842 0.000500915
R9991 GND.n4086 GND.n4085 0.000500552
R9992 GND.n4101 GND.n4100 0.000500539
R9993 GND.n4955 GND.n4954 0.000500526
R9994 GND.n4970 GND.n4969 0.000500526
R9995 GND.n3399 GND.n3398 0.000500526
R9996 GND.n3141 GND.n3140 0.000500526
R9997 GND.n2343 GND.n2342 0.000500526
R9998 GND.n1867 GND.n1866 0.000500526
R9999 GND.n5327 GND.n5326 0.000500526
R10000 GND.n3577 GND.n3576 0.000500526
R10001 GND.n5316 GND.n5315 0.000500526
R10002 GND.n5307 GND.n5306 0.000500526
R10003 GND.n3898 GND.n3897 0.000500526
R10004 GND.n3571 GND.n3570 0.000500526
R10005 GND.n3414 GND.n3413 0.000500526
R10006 GND.n2182 GND.n2181 0.000500526
R10007 GND.n2497 GND.n2496 0.000500526
R10008 GND.n2812 GND.n2811 0.000500526
R10009 GND.n4482 GND.n4481 0.000500355
R10010 GND.n4560 GND.n4559 0.000500347
R10011 GND.n4670 GND.n4668 0.000500286
R10012 GND.n3208 GND.n3207 0.000500286
R10013 GND.n2255 GND.n2254 0.000500286
R10014 GND.n7667 GND.n7665 0.000500286
R10015 GND.n1515 GND.n1514 0.000500286
R10016 GND.n5352 GND.n5351 0.000500286
R10017 GND.n3921 GND.n3920 0.000500286
R10018 GND.n5213 GND.n5212 0.000500286
R10019 GND.n3813 GND.n3812 0.000500286
R10020 GND.n3490 GND.n3489 0.000500286
R10021 GND.n1942 GND.n1941 0.000500286
R10022 GND.n2051 GND.n2049 0.000500286
R10023 GND.n2417 GND.n2416 0.000500286
R10024 GND.n2726 GND.n2725 0.000500286
R10025 GND.n4871 GND.n4870 0.000500286
R10026 GND.n2836 GND.n2835 0.000500286
R10027 GND.n4287 GND.n4286 0.000500199
R10028 GND.n6139 GND.n6138 0.00050016
R10029 GND.n4295 GND.n4294 0.000500107
R10030 GND.n4953 GND.n4952 0.000500059
R10031 GND.n4973 GND.n4972 0.000500059
R10032 GND.n2346 GND.n2345 0.000500059
R10033 GND.n1865 GND.n150 0.000500059
R10034 GND.n5330 GND.n5329 0.000500059
R10035 GND.n5337 GND.n1333 0.000500059
R10036 GND.n5314 GND.n5313 0.000500059
R10037 GND.n5310 GND.n5309 0.000500059
R10038 GND.n3896 GND.n3895 0.000500059
R10039 GND.n3569 GND.n3568 0.000500059
R10040 GND.n3412 GND.n3411 0.000500059
R10041 GND.n2185 GND.n2184 0.000500059
R10042 GND.n2500 GND.n2499 0.000500059
R10043 GND.n2815 GND.n2814 0.000500059
R10044 GND.n3144 GND.n3143 0.000500059
R10045 GND.n3402 GND.n3401 0.000500059
R10046 GND.n4585 GND.n4584 0.000500053
R10047 GND.n4580 GND.n4579 0.000500023
R10048 GND.n1441 GND.n1440 0.00050002
R10049 VDD.n1970 VDD.n1931 8089.41
R10050 VDD.n1951 VDD.n1949 8089.41
R10051 VDD.n1954 VDD.n1948 6801.18
R10052 VDD.n1913 VDD.n1895 2565.88
R10053 VDD.n1913 VDD.n1896 2565.88
R10054 VDD.n1878 VDD.n1823 2565.88
R10055 VDD.n1859 VDD.n1848 2565.88
R10056 VDD.n1864 VDD.n1848 2565.88
R10057 VDD.n2180 VDD.n2169 2565.88
R10058 VDD.n2185 VDD.n2169 2565.88
R10059 VDD.n2199 VDD.n2144 2565.88
R10060 VDD.n2234 VDD.n2216 2565.88
R10061 VDD.n2234 VDD.n2217 2565.88
R10062 VDD.n2438 VDD.n2427 2565.88
R10063 VDD.n2443 VDD.n2427 2565.88
R10064 VDD.n2457 VDD.n2402 2565.88
R10065 VDD.n2492 VDD.n2474 2565.88
R10066 VDD.n2492 VDD.n2475 2565.88
R10067 VDD.n2696 VDD.n2685 2565.88
R10068 VDD.n2701 VDD.n2685 2565.88
R10069 VDD.n2715 VDD.n2660 2565.88
R10070 VDD.n2750 VDD.n2732 2565.88
R10071 VDD.n2750 VDD.n2733 2565.88
R10072 VDD.n2954 VDD.n2943 2565.88
R10073 VDD.n2959 VDD.n2943 2565.88
R10074 VDD.n2973 VDD.n2918 2565.88
R10075 VDD.n3008 VDD.n2990 2565.88
R10076 VDD.n3008 VDD.n2991 2565.88
R10077 VDD.n3212 VDD.n3201 2565.88
R10078 VDD.n3217 VDD.n3201 2565.88
R10079 VDD.n3231 VDD.n3176 2565.88
R10080 VDD.n3266 VDD.n3248 2565.88
R10081 VDD.n3266 VDD.n3249 2565.88
R10082 VDD.n3470 VDD.n3459 2565.88
R10083 VDD.n3475 VDD.n3459 2565.88
R10084 VDD.n3489 VDD.n3434 2565.88
R10085 VDD.n3524 VDD.n3506 2565.88
R10086 VDD.n3524 VDD.n3507 2565.88
R10087 VDD.n5790 VDD.n5779 2565.88
R10088 VDD.n5795 VDD.n5779 2565.88
R10089 VDD.n5809 VDD.n5754 2565.88
R10090 VDD.n5844 VDD.n5826 2565.88
R10091 VDD.n5844 VDD.n5827 2565.88
R10092 VDD.n5536 VDD.n5525 2565.88
R10093 VDD.n5541 VDD.n5525 2565.88
R10094 VDD.n5555 VDD.n5500 2565.88
R10095 VDD.n5590 VDD.n5572 2565.88
R10096 VDD.n5590 VDD.n5573 2565.88
R10097 VDD.n3728 VDD.n3717 2565.88
R10098 VDD.n3733 VDD.n3717 2565.88
R10099 VDD.n3747 VDD.n3692 2565.88
R10100 VDD.n3782 VDD.n3764 2565.88
R10101 VDD.n3782 VDD.n3765 2565.88
R10102 VDD.n3986 VDD.n3975 2565.88
R10103 VDD.n3991 VDD.n3975 2565.88
R10104 VDD.n4005 VDD.n3950 2565.88
R10105 VDD.n4040 VDD.n4022 2565.88
R10106 VDD.n4040 VDD.n4023 2565.88
R10107 VDD.n4244 VDD.n4233 2565.88
R10108 VDD.n4249 VDD.n4233 2565.88
R10109 VDD.n4263 VDD.n4208 2565.88
R10110 VDD.n4298 VDD.n4280 2565.88
R10111 VDD.n4298 VDD.n4281 2565.88
R10112 VDD.n4502 VDD.n4491 2565.88
R10113 VDD.n4507 VDD.n4491 2565.88
R10114 VDD.n4521 VDD.n4466 2565.88
R10115 VDD.n4556 VDD.n4538 2565.88
R10116 VDD.n4556 VDD.n4539 2565.88
R10117 VDD.n4760 VDD.n4749 2565.88
R10118 VDD.n4765 VDD.n4749 2565.88
R10119 VDD.n4779 VDD.n4724 2565.88
R10120 VDD.n4814 VDD.n4796 2565.88
R10121 VDD.n4814 VDD.n4797 2565.88
R10122 VDD.n5018 VDD.n5007 2565.88
R10123 VDD.n5023 VDD.n5007 2565.88
R10124 VDD.n5037 VDD.n4982 2565.88
R10125 VDD.n5072 VDD.n5054 2565.88
R10126 VDD.n5072 VDD.n5055 2565.88
R10127 VDD.n5276 VDD.n5265 2565.88
R10128 VDD.n5281 VDD.n5265 2565.88
R10129 VDD.n5295 VDD.n5240 2565.88
R10130 VDD.n5330 VDD.n5312 2565.88
R10131 VDD.n5330 VDD.n5313 2565.88
R10132 VDD.n1744 VDD.n1713 2082.55
R10133 VDD.n2093 VDD.n2062 2082.55
R10134 VDD.n2323 VDD.n2292 2082.55
R10135 VDD.n2581 VDD.n2550 2082.55
R10136 VDD.n2839 VDD.n2808 2082.55
R10137 VDD.n3097 VDD.n3066 2082.55
R10138 VDD.n3355 VDD.n3324 2082.55
R10139 VDD.n5678 VDD.n5647 2082.55
R10140 VDD.n5424 VDD.n5393 2082.55
R10141 VDD.n3613 VDD.n3582 2082.55
R10142 VDD.n3871 VDD.n3840 2082.55
R10143 VDD.n4129 VDD.n4098 2082.55
R10144 VDD.n4387 VDD.n4356 2082.55
R10145 VDD.n4645 VDD.n4614 2082.55
R10146 VDD.n4903 VDD.n4872 2082.55
R10147 VDD.n5161 VDD.n5130 2082.55
R10148 VDD.n1694 VDD.n1674 2080.64
R10149 VDD.n2043 VDD.n2023 2080.64
R10150 VDD.n2273 VDD.n2253 2080.64
R10151 VDD.n2531 VDD.n2511 2080.64
R10152 VDD.n2789 VDD.n2769 2080.64
R10153 VDD.n3047 VDD.n3027 2080.64
R10154 VDD.n3305 VDD.n3285 2080.64
R10155 VDD.n5628 VDD.n5608 2080.64
R10156 VDD.n5374 VDD.n5354 2080.64
R10157 VDD.n3563 VDD.n3543 2080.64
R10158 VDD.n3821 VDD.n3801 2080.64
R10159 VDD.n4079 VDD.n4059 2080.64
R10160 VDD.n4337 VDD.n4317 2080.64
R10161 VDD.n4595 VDD.n4575 2080.64
R10162 VDD.n4853 VDD.n4833 2080.64
R10163 VDD.n5111 VDD.n5091 2080.64
R10164 VDD.n1742 VDD.n1712 2015.29
R10165 VDD.n1698 VDD.n1678 2015.29
R10166 VDD.n2091 VDD.n2061 2015.29
R10167 VDD.n2047 VDD.n2027 2015.29
R10168 VDD.n2321 VDD.n2291 2015.29
R10169 VDD.n2277 VDD.n2257 2015.29
R10170 VDD.n2579 VDD.n2549 2015.29
R10171 VDD.n2535 VDD.n2515 2015.29
R10172 VDD.n2837 VDD.n2807 2015.29
R10173 VDD.n2793 VDD.n2773 2015.29
R10174 VDD.n3095 VDD.n3065 2015.29
R10175 VDD.n3051 VDD.n3031 2015.29
R10176 VDD.n3353 VDD.n3323 2015.29
R10177 VDD.n3309 VDD.n3289 2015.29
R10178 VDD.n5676 VDD.n5646 2015.29
R10179 VDD.n5632 VDD.n5612 2015.29
R10180 VDD.n5422 VDD.n5392 2015.29
R10181 VDD.n5378 VDD.n5358 2015.29
R10182 VDD.n3611 VDD.n3581 2015.29
R10183 VDD.n3567 VDD.n3547 2015.29
R10184 VDD.n3869 VDD.n3839 2015.29
R10185 VDD.n3825 VDD.n3805 2015.29
R10186 VDD.n4127 VDD.n4097 2015.29
R10187 VDD.n4083 VDD.n4063 2015.29
R10188 VDD.n4385 VDD.n4355 2015.29
R10189 VDD.n4341 VDD.n4321 2015.29
R10190 VDD.n4643 VDD.n4613 2015.29
R10191 VDD.n4599 VDD.n4579 2015.29
R10192 VDD.n4901 VDD.n4871 2015.29
R10193 VDD.n4857 VDD.n4837 2015.29
R10194 VDD.n5159 VDD.n5129 2015.29
R10195 VDD.n5115 VDD.n5095 2015.29
R10196 VDD.n1904 VDD.n1894 1997.65
R10197 VDD.n1899 VDD.n1894 1997.65
R10198 VDD.n1868 VDD.n1850 1997.65
R10199 VDD.n1868 VDD.n1851 1997.65
R10200 VDD.n2189 VDD.n2171 1997.65
R10201 VDD.n2189 VDD.n2172 1997.65
R10202 VDD.n2225 VDD.n2215 1997.65
R10203 VDD.n2220 VDD.n2215 1997.65
R10204 VDD.n2447 VDD.n2429 1997.65
R10205 VDD.n2447 VDD.n2430 1997.65
R10206 VDD.n2483 VDD.n2473 1997.65
R10207 VDD.n2478 VDD.n2473 1997.65
R10208 VDD.n2705 VDD.n2687 1997.65
R10209 VDD.n2705 VDD.n2688 1997.65
R10210 VDD.n2741 VDD.n2731 1997.65
R10211 VDD.n2736 VDD.n2731 1997.65
R10212 VDD.n2963 VDD.n2945 1997.65
R10213 VDD.n2963 VDD.n2946 1997.65
R10214 VDD.n2999 VDD.n2989 1997.65
R10215 VDD.n2994 VDD.n2989 1997.65
R10216 VDD.n3221 VDD.n3203 1997.65
R10217 VDD.n3221 VDD.n3204 1997.65
R10218 VDD.n3257 VDD.n3247 1997.65
R10219 VDD.n3252 VDD.n3247 1997.65
R10220 VDD.n3479 VDD.n3461 1997.65
R10221 VDD.n3479 VDD.n3462 1997.65
R10222 VDD.n3515 VDD.n3505 1997.65
R10223 VDD.n3510 VDD.n3505 1997.65
R10224 VDD.n5799 VDD.n5781 1997.65
R10225 VDD.n5799 VDD.n5782 1997.65
R10226 VDD.n5835 VDD.n5825 1997.65
R10227 VDD.n5830 VDD.n5825 1997.65
R10228 VDD.n5545 VDD.n5527 1997.65
R10229 VDD.n5545 VDD.n5528 1997.65
R10230 VDD.n5581 VDD.n5571 1997.65
R10231 VDD.n5576 VDD.n5571 1997.65
R10232 VDD.n3737 VDD.n3719 1997.65
R10233 VDD.n3737 VDD.n3720 1997.65
R10234 VDD.n3773 VDD.n3763 1997.65
R10235 VDD.n3768 VDD.n3763 1997.65
R10236 VDD.n3995 VDD.n3977 1997.65
R10237 VDD.n3995 VDD.n3978 1997.65
R10238 VDD.n4031 VDD.n4021 1997.65
R10239 VDD.n4026 VDD.n4021 1997.65
R10240 VDD.n4253 VDD.n4235 1997.65
R10241 VDD.n4253 VDD.n4236 1997.65
R10242 VDD.n4289 VDD.n4279 1997.65
R10243 VDD.n4284 VDD.n4279 1997.65
R10244 VDD.n4511 VDD.n4493 1997.65
R10245 VDD.n4511 VDD.n4494 1997.65
R10246 VDD.n4547 VDD.n4537 1997.65
R10247 VDD.n4542 VDD.n4537 1997.65
R10248 VDD.n4769 VDD.n4751 1997.65
R10249 VDD.n4769 VDD.n4752 1997.65
R10250 VDD.n4805 VDD.n4795 1997.65
R10251 VDD.n4800 VDD.n4795 1997.65
R10252 VDD.n5027 VDD.n5009 1997.65
R10253 VDD.n5027 VDD.n5010 1997.65
R10254 VDD.n5063 VDD.n5053 1997.65
R10255 VDD.n5058 VDD.n5053 1997.65
R10256 VDD.n5285 VDD.n5267 1997.65
R10257 VDD.n5285 VDD.n5268 1997.65
R10258 VDD.n5321 VDD.n5311 1997.65
R10259 VDD.n5316 VDD.n5311 1997.65
R10260 VDD.n1878 VDD.n1819 1814.12
R10261 VDD.n2199 VDD.n2140 1814.12
R10262 VDD.n2457 VDD.n2398 1814.12
R10263 VDD.n2715 VDD.n2656 1814.12
R10264 VDD.n2973 VDD.n2914 1814.12
R10265 VDD.n3231 VDD.n3172 1814.12
R10266 VDD.n3489 VDD.n3430 1814.12
R10267 VDD.n5809 VDD.n5750 1814.12
R10268 VDD.n5555 VDD.n5496 1814.12
R10269 VDD.n3747 VDD.n3688 1814.12
R10270 VDD.n4005 VDD.n3946 1814.12
R10271 VDD.n4263 VDD.n4204 1814.12
R10272 VDD.n4521 VDD.n4462 1814.12
R10273 VDD.n4779 VDD.n4720 1814.12
R10274 VDD.n5037 VDD.n4978 1814.12
R10275 VDD.n5295 VDD.n5236 1814.12
R10276 VDD.n1881 VDD.n1880 1598.82
R10277 VDD.n2202 VDD.n2201 1598.82
R10278 VDD.n2460 VDD.n2459 1598.82
R10279 VDD.n2718 VDD.n2717 1598.82
R10280 VDD.n2976 VDD.n2975 1598.82
R10281 VDD.n3234 VDD.n3233 1598.82
R10282 VDD.n3492 VDD.n3491 1598.82
R10283 VDD.n5812 VDD.n5811 1598.82
R10284 VDD.n5558 VDD.n5557 1598.82
R10285 VDD.n3750 VDD.n3749 1598.82
R10286 VDD.n4008 VDD.n4007 1598.82
R10287 VDD.n4266 VDD.n4265 1598.82
R10288 VDD.n4524 VDD.n4523 1598.82
R10289 VDD.n4782 VDD.n4781 1598.82
R10290 VDD.n5040 VDD.n5039 1598.82
R10291 VDD.n5298 VDD.n5297 1598.82
R10292 VDD.n1698 VDD.n1697 1514.12
R10293 VDD.n2047 VDD.n2046 1514.12
R10294 VDD.n2277 VDD.n2276 1514.12
R10295 VDD.n2535 VDD.n2534 1514.12
R10296 VDD.n2793 VDD.n2792 1514.12
R10297 VDD.n3051 VDD.n3050 1514.12
R10298 VDD.n3309 VDD.n3308 1514.12
R10299 VDD.n5632 VDD.n5631 1514.12
R10300 VDD.n5378 VDD.n5377 1514.12
R10301 VDD.n3567 VDD.n3566 1514.12
R10302 VDD.n3825 VDD.n3824 1514.12
R10303 VDD.n4083 VDD.n4082 1514.12
R10304 VDD.n4341 VDD.n4340 1514.12
R10305 VDD.n4599 VDD.n4598 1514.12
R10306 VDD.n4857 VDD.n4856 1514.12
R10307 VDD.n5115 VDD.n5114 1514.12
R10308 VDD.n1856 VDD.n1844 1440
R10309 VDD.n1869 VDD.n1846 1440
R10310 VDD.n2177 VDD.n2165 1440
R10311 VDD.n2190 VDD.n2167 1440
R10312 VDD.n2435 VDD.n2423 1440
R10313 VDD.n2448 VDD.n2425 1440
R10314 VDD.n2693 VDD.n2681 1440
R10315 VDD.n2706 VDD.n2683 1440
R10316 VDD.n2951 VDD.n2939 1440
R10317 VDD.n2964 VDD.n2941 1440
R10318 VDD.n3209 VDD.n3197 1440
R10319 VDD.n3222 VDD.n3199 1440
R10320 VDD.n3467 VDD.n3455 1440
R10321 VDD.n3480 VDD.n3457 1440
R10322 VDD.n5787 VDD.n5775 1440
R10323 VDD.n5800 VDD.n5777 1440
R10324 VDD.n5533 VDD.n5521 1440
R10325 VDD.n5546 VDD.n5523 1440
R10326 VDD.n3725 VDD.n3713 1440
R10327 VDD.n3738 VDD.n3715 1440
R10328 VDD.n3983 VDD.n3971 1440
R10329 VDD.n3996 VDD.n3973 1440
R10330 VDD.n4241 VDD.n4229 1440
R10331 VDD.n4254 VDD.n4231 1440
R10332 VDD.n4499 VDD.n4487 1440
R10333 VDD.n4512 VDD.n4489 1440
R10334 VDD.n4757 VDD.n4745 1440
R10335 VDD.n4770 VDD.n4747 1440
R10336 VDD.n5015 VDD.n5003 1440
R10337 VDD.n5028 VDD.n5005 1440
R10338 VDD.n5273 VDD.n5261 1440
R10339 VDD.n5286 VDD.n5263 1440
R10340 VDD.n1915 VDD.n1890 1422.35
R10341 VDD.n1900 VDD.n1891 1422.35
R10342 VDD.n2236 VDD.n2211 1422.35
R10343 VDD.n2221 VDD.n2212 1422.35
R10344 VDD.n2494 VDD.n2469 1422.35
R10345 VDD.n2479 VDD.n2470 1422.35
R10346 VDD.n2752 VDD.n2727 1422.35
R10347 VDD.n2737 VDD.n2728 1422.35
R10348 VDD.n3010 VDD.n2985 1422.35
R10349 VDD.n2995 VDD.n2986 1422.35
R10350 VDD.n3268 VDD.n3243 1422.35
R10351 VDD.n3253 VDD.n3244 1422.35
R10352 VDD.n3526 VDD.n3501 1422.35
R10353 VDD.n3511 VDD.n3502 1422.35
R10354 VDD.n5846 VDD.n5821 1422.35
R10355 VDD.n5831 VDD.n5822 1422.35
R10356 VDD.n5592 VDD.n5567 1422.35
R10357 VDD.n5577 VDD.n5568 1422.35
R10358 VDD.n3784 VDD.n3759 1422.35
R10359 VDD.n3769 VDD.n3760 1422.35
R10360 VDD.n4042 VDD.n4017 1422.35
R10361 VDD.n4027 VDD.n4018 1422.35
R10362 VDD.n4300 VDD.n4275 1422.35
R10363 VDD.n4285 VDD.n4276 1422.35
R10364 VDD.n4558 VDD.n4533 1422.35
R10365 VDD.n4543 VDD.n4534 1422.35
R10366 VDD.n4816 VDD.n4791 1422.35
R10367 VDD.n4801 VDD.n4792 1422.35
R10368 VDD.n5074 VDD.n5049 1422.35
R10369 VDD.n5059 VDD.n5050 1422.35
R10370 VDD.n5332 VDD.n5307 1422.35
R10371 VDD.n5317 VDD.n5308 1422.35
R10372 VDD.n857 VDD 1319.65
R10373 VDD.n1240 VDD 1319.65
R10374 VDD.n1713 VDD.n1676 1231.76
R10375 VDD.n2062 VDD.n2025 1231.76
R10376 VDD.n2292 VDD.n2255 1231.76
R10377 VDD.n2550 VDD.n2513 1231.76
R10378 VDD.n2808 VDD.n2771 1231.76
R10379 VDD.n3066 VDD.n3029 1231.76
R10380 VDD.n3324 VDD.n3287 1231.76
R10381 VDD.n5647 VDD.n5610 1231.76
R10382 VDD.n5393 VDD.n5356 1231.76
R10383 VDD.n3582 VDD.n3545 1231.76
R10384 VDD.n3840 VDD.n3803 1231.76
R10385 VDD.n4098 VDD.n4061 1231.76
R10386 VDD.n4356 VDD.n4319 1231.76
R10387 VDD.n4614 VDD.n4577 1231.76
R10388 VDD.n4872 VDD.n4835 1231.76
R10389 VDD.n5130 VDD.n5093 1231.76
R10390 VDD.n1765 VDD.n1674 1228.24
R10391 VDD.n2114 VDD.n2023 1228.24
R10392 VDD.n2344 VDD.n2253 1228.24
R10393 VDD.n2602 VDD.n2511 1228.24
R10394 VDD.n2860 VDD.n2769 1228.24
R10395 VDD.n3118 VDD.n3027 1228.24
R10396 VDD.n3376 VDD.n3285 1228.24
R10397 VDD.n5699 VDD.n5608 1228.24
R10398 VDD.n5445 VDD.n5354 1228.24
R10399 VDD.n3634 VDD.n3543 1228.24
R10400 VDD.n3892 VDD.n3801 1228.24
R10401 VDD.n4150 VDD.n4059 1228.24
R10402 VDD.n4408 VDD.n4317 1228.24
R10403 VDD.n4666 VDD.n4575 1228.24
R10404 VDD.n4924 VDD.n4833 1228.24
R10405 VDD.n5182 VDD.n5091 1228.24
R10406 VDD.n1765 VDD.n1675 1224.71
R10407 VDD.n1676 VDD.n1675 1224.71
R10408 VDD.n2114 VDD.n2024 1224.71
R10409 VDD.n2025 VDD.n2024 1224.71
R10410 VDD.n2344 VDD.n2254 1224.71
R10411 VDD.n2255 VDD.n2254 1224.71
R10412 VDD.n2602 VDD.n2512 1224.71
R10413 VDD.n2513 VDD.n2512 1224.71
R10414 VDD.n2860 VDD.n2770 1224.71
R10415 VDD.n2771 VDD.n2770 1224.71
R10416 VDD.n3118 VDD.n3028 1224.71
R10417 VDD.n3029 VDD.n3028 1224.71
R10418 VDD.n3376 VDD.n3286 1224.71
R10419 VDD.n3287 VDD.n3286 1224.71
R10420 VDD.n5699 VDD.n5609 1224.71
R10421 VDD.n5610 VDD.n5609 1224.71
R10422 VDD.n5445 VDD.n5355 1224.71
R10423 VDD.n5356 VDD.n5355 1224.71
R10424 VDD.n3634 VDD.n3544 1224.71
R10425 VDD.n3545 VDD.n3544 1224.71
R10426 VDD.n3892 VDD.n3802 1224.71
R10427 VDD.n3803 VDD.n3802 1224.71
R10428 VDD.n4150 VDD.n4060 1224.71
R10429 VDD.n4061 VDD.n4060 1224.71
R10430 VDD.n4408 VDD.n4318 1224.71
R10431 VDD.n4319 VDD.n4318 1224.71
R10432 VDD.n4666 VDD.n4576 1224.71
R10433 VDD.n4577 VDD.n4576 1224.71
R10434 VDD.n4924 VDD.n4834 1224.71
R10435 VDD.n4835 VDD.n4834 1224.71
R10436 VDD.n5182 VDD.n5092 1224.71
R10437 VDD.n5093 VDD.n5092 1224.71
R10438 VDD.n1718 VDD.n1675 1153.33
R10439 VDD.n2067 VDD.n2024 1153.33
R10440 VDD.n2297 VDD.n2254 1153.33
R10441 VDD.n2555 VDD.n2512 1153.33
R10442 VDD.n2813 VDD.n2770 1153.33
R10443 VDD.n3071 VDD.n3028 1153.33
R10444 VDD.n3329 VDD.n3286 1153.33
R10445 VDD.n5652 VDD.n5609 1153.33
R10446 VDD.n5398 VDD.n5355 1153.33
R10447 VDD.n3587 VDD.n3544 1153.33
R10448 VDD.n3845 VDD.n3802 1153.33
R10449 VDD.n4103 VDD.n4060 1153.33
R10450 VDD.n4361 VDD.n4318 1153.33
R10451 VDD.n4619 VDD.n4576 1153.33
R10452 VDD.n4877 VDD.n4834 1153.33
R10453 VDD.n5135 VDD.n5092 1153.33
R10454 VDD.n1902 VDD.n1900 1143.53
R10455 VDD.n2223 VDD.n2221 1143.53
R10456 VDD.n2481 VDD.n2479 1143.53
R10457 VDD.n2739 VDD.n2737 1143.53
R10458 VDD.n2997 VDD.n2995 1143.53
R10459 VDD.n3255 VDD.n3253 1143.53
R10460 VDD.n3513 VDD.n3511 1143.53
R10461 VDD.n5833 VDD.n5831 1143.53
R10462 VDD.n5579 VDD.n5577 1143.53
R10463 VDD.n3771 VDD.n3769 1143.53
R10464 VDD.n4029 VDD.n4027 1143.53
R10465 VDD.n4287 VDD.n4285 1143.53
R10466 VDD.n4545 VDD.n4543 1143.53
R10467 VDD.n4803 VDD.n4801 1143.53
R10468 VDD.n5061 VDD.n5059 1143.53
R10469 VDD.n5319 VDD.n5317 1143.53
R10470 VDD.n1862 VDD.n1846 1125.88
R10471 VDD.n2183 VDD.n2167 1125.88
R10472 VDD.n2441 VDD.n2425 1125.88
R10473 VDD.n2699 VDD.n2683 1125.88
R10474 VDD.n2957 VDD.n2941 1125.88
R10475 VDD.n3215 VDD.n3199 1125.88
R10476 VDD.n3473 VDD.n3457 1125.88
R10477 VDD.n5793 VDD.n5777 1125.88
R10478 VDD.n5539 VDD.n5523 1125.88
R10479 VDD.n3731 VDD.n3715 1125.88
R10480 VDD.n3989 VDD.n3973 1125.88
R10481 VDD.n4247 VDD.n4231 1125.88
R10482 VDD.n4505 VDD.n4489 1125.88
R10483 VDD.n4763 VDD.n4747 1125.88
R10484 VDD.n5021 VDD.n5005 1125.88
R10485 VDD.n5279 VDD.n5263 1125.88
R10486 VDD.n1756 VDD.n1718 1072.94
R10487 VDD.n2105 VDD.n2067 1072.94
R10488 VDD.n2335 VDD.n2297 1072.94
R10489 VDD.n2593 VDD.n2555 1072.94
R10490 VDD.n2851 VDD.n2813 1072.94
R10491 VDD.n3109 VDD.n3071 1072.94
R10492 VDD.n3367 VDD.n3329 1072.94
R10493 VDD.n5690 VDD.n5652 1072.94
R10494 VDD.n5436 VDD.n5398 1072.94
R10495 VDD.n3625 VDD.n3587 1072.94
R10496 VDD.n3883 VDD.n3845 1072.94
R10497 VDD.n4141 VDD.n4103 1072.94
R10498 VDD.n4399 VDD.n4361 1072.94
R10499 VDD.n4657 VDD.n4619 1072.94
R10500 VDD.n4915 VDD.n4877 1072.94
R10501 VDD.n5173 VDD.n5135 1072.94
R10502 VDD.n1718 VDD.n1670 1069.41
R10503 VDD.n2067 VDD.n2019 1069.41
R10504 VDD.n2297 VDD.n2249 1069.41
R10505 VDD.n2555 VDD.n2507 1069.41
R10506 VDD.n2813 VDD.n2765 1069.41
R10507 VDD.n3071 VDD.n3023 1069.41
R10508 VDD.n3329 VDD.n3281 1069.41
R10509 VDD.n5652 VDD.n5604 1069.41
R10510 VDD.n5398 VDD.n5350 1069.41
R10511 VDD.n3587 VDD.n3539 1069.41
R10512 VDD.n3845 VDD.n3797 1069.41
R10513 VDD.n4103 VDD.n4055 1069.41
R10514 VDD.n4361 VDD.n4313 1069.41
R10515 VDD.n4619 VDD.n4571 1069.41
R10516 VDD.n4877 VDD.n4829 1069.41
R10517 VDD.n5135 VDD.n5087 1069.41
R10518 VDD.n1906 VDD.n1890 1051.76
R10519 VDD.n1856 VDD.n1855 1051.76
R10520 VDD.n2177 VDD.n2176 1051.76
R10521 VDD.n2227 VDD.n2211 1051.76
R10522 VDD.n2435 VDD.n2434 1051.76
R10523 VDD.n2485 VDD.n2469 1051.76
R10524 VDD.n2693 VDD.n2692 1051.76
R10525 VDD.n2743 VDD.n2727 1051.76
R10526 VDD.n2951 VDD.n2950 1051.76
R10527 VDD.n3001 VDD.n2985 1051.76
R10528 VDD.n3209 VDD.n3208 1051.76
R10529 VDD.n3259 VDD.n3243 1051.76
R10530 VDD.n3467 VDD.n3466 1051.76
R10531 VDD.n3517 VDD.n3501 1051.76
R10532 VDD.n5787 VDD.n5786 1051.76
R10533 VDD.n5837 VDD.n5821 1051.76
R10534 VDD.n5533 VDD.n5532 1051.76
R10535 VDD.n5583 VDD.n5567 1051.76
R10536 VDD.n3725 VDD.n3724 1051.76
R10537 VDD.n3775 VDD.n3759 1051.76
R10538 VDD.n3983 VDD.n3982 1051.76
R10539 VDD.n4033 VDD.n4017 1051.76
R10540 VDD.n4241 VDD.n4240 1051.76
R10541 VDD.n4291 VDD.n4275 1051.76
R10542 VDD.n4499 VDD.n4498 1051.76
R10543 VDD.n4549 VDD.n4533 1051.76
R10544 VDD.n4757 VDD.n4756 1051.76
R10545 VDD.n4807 VDD.n4791 1051.76
R10546 VDD.n5015 VDD.n5014 1051.76
R10547 VDD.n5065 VDD.n5049 1051.76
R10548 VDD.n5273 VDD.n5272 1051.76
R10549 VDD.n5323 VDD.n5307 1051.76
R10550 VDD.n1960 VDD.n1942 862.871
R10551 VDD.n1950 VDD.n1942 862.871
R10552 VDD.n1971 VDD.n1930 862.871
R10553 VDD.n1967 VDD.n1930 862.871
R10554 VDD.n1759 VDD.n1758 861.178
R10555 VDD.n2108 VDD.n2107 861.178
R10556 VDD.n2338 VDD.n2337 861.178
R10557 VDD.n2596 VDD.n2595 861.178
R10558 VDD.n2854 VDD.n2853 861.178
R10559 VDD.n3112 VDD.n3111 861.178
R10560 VDD.n3370 VDD.n3369 861.178
R10561 VDD.n5693 VDD.n5692 861.178
R10562 VDD.n5439 VDD.n5438 861.178
R10563 VDD.n3628 VDD.n3627 861.178
R10564 VDD.n3886 VDD.n3885 861.178
R10565 VDD.n4144 VDD.n4143 861.178
R10566 VDD.n4402 VDD.n4401 861.178
R10567 VDD.n4660 VDD.n4659 861.178
R10568 VDD.n4918 VDD.n4917 861.178
R10569 VDD.n5176 VDD.n5175 861.178
R10570 VDD.n1962 VDD.n1961 857.648
R10571 VDD.n1963 VDD.n1962 857.648
R10572 VDD.n1963 VDD.n1928 857.648
R10573 VDD.n1970 VDD.n1928 857.648
R10574 VDD.n1951 VDD.n1938 857.648
R10575 VDD.n1964 VDD.n1938 857.648
R10576 VDD.n1964 VDD.n1932 857.648
R10577 VDD.n1968 VDD.n1932 857.648
R10578 VDD.n1883 VDD.n1819 751.765
R10579 VDD.n2204 VDD.n2140 751.765
R10580 VDD.n2462 VDD.n2398 751.765
R10581 VDD.n2720 VDD.n2656 751.765
R10582 VDD.n2978 VDD.n2914 751.765
R10583 VDD.n3236 VDD.n3172 751.765
R10584 VDD.n3494 VDD.n3430 751.765
R10585 VDD.n5814 VDD.n5750 751.765
R10586 VDD.n5560 VDD.n5496 751.765
R10587 VDD.n3752 VDD.n3688 751.765
R10588 VDD.n4010 VDD.n3946 751.765
R10589 VDD.n4268 VDD.n4204 751.765
R10590 VDD.n4526 VDD.n4462 751.765
R10591 VDD.n4784 VDD.n4720 751.765
R10592 VDD.n5042 VDD.n4978 751.765
R10593 VDD.n5300 VDD.n5236 751.765
R10594 VDD.n1714 VDD.n1712 723.529
R10595 VDD.n2063 VDD.n2061 723.529
R10596 VDD.n2293 VDD.n2291 723.529
R10597 VDD.n2551 VDD.n2549 723.529
R10598 VDD.n2809 VDD.n2807 723.529
R10599 VDD.n3067 VDD.n3065 723.529
R10600 VDD.n3325 VDD.n3323 723.529
R10601 VDD.n5648 VDD.n5646 723.529
R10602 VDD.n5394 VDD.n5392 723.529
R10603 VDD.n3583 VDD.n3581 723.529
R10604 VDD.n3841 VDD.n3839 723.529
R10605 VDD.n4099 VDD.n4097 723.529
R10606 VDD.n4357 VDD.n4355 723.529
R10607 VDD.n4615 VDD.n4613 723.529
R10608 VDD.n4873 VDD.n4871 723.529
R10609 VDD.n5131 VDD.n5129 723.529
R10610 VDD.n1680 VDD.n1678 720
R10611 VDD.n2029 VDD.n2027 720
R10612 VDD.n2259 VDD.n2257 720
R10613 VDD.n2517 VDD.n2515 720
R10614 VDD.n2775 VDD.n2773 720
R10615 VDD.n3033 VDD.n3031 720
R10616 VDD.n3291 VDD.n3289 720
R10617 VDD.n5614 VDD.n5612 720
R10618 VDD.n5360 VDD.n5358 720
R10619 VDD.n3549 VDD.n3547 720
R10620 VDD.n3807 VDD.n3805 720
R10621 VDD.n4065 VDD.n4063 720
R10622 VDD.n4323 VDD.n4321 720
R10623 VDD.n4581 VDD.n4579 720
R10624 VDD.n4839 VDD.n4837 720
R10625 VDD.n5097 VDD.n5095 720
R10626 VDD.n1695 VDD.t1031 632.183
R10627 VDD.n2044 VDD.t1264 632.183
R10628 VDD.n2274 VDD.t831 632.183
R10629 VDD.n2532 VDD.t1417 632.183
R10630 VDD.n2790 VDD.t436 632.183
R10631 VDD.n3048 VDD.t383 632.183
R10632 VDD.n3306 VDD.t1295 632.183
R10633 VDD.n5629 VDD.t476 632.183
R10634 VDD.n5375 VDD.t1258 632.183
R10635 VDD.n3564 VDD.t1366 632.183
R10636 VDD.n3822 VDD.t1114 632.183
R10637 VDD.n4080 VDD.t30 632.183
R10638 VDD.n4338 VDD.t1436 632.183
R10639 VDD.n4596 VDD.t370 632.183
R10640 VDD.n4854 VDD.t422 632.183
R10641 VDD.n5112 VDD.t0 632.183
R10642 VDD.n1677 VDD.n1674 593.144
R10643 VDD.n1680 VDD.n1677 593.144
R10644 VDD.n2026 VDD.n2023 593.144
R10645 VDD.n2029 VDD.n2026 593.144
R10646 VDD.n2256 VDD.n2253 593.144
R10647 VDD.n2259 VDD.n2256 593.144
R10648 VDD.n2514 VDD.n2511 593.144
R10649 VDD.n2517 VDD.n2514 593.144
R10650 VDD.n2772 VDD.n2769 593.144
R10651 VDD.n2775 VDD.n2772 593.144
R10652 VDD.n3030 VDD.n3027 593.144
R10653 VDD.n3033 VDD.n3030 593.144
R10654 VDD.n3288 VDD.n3285 593.144
R10655 VDD.n3291 VDD.n3288 593.144
R10656 VDD.n5611 VDD.n5608 593.144
R10657 VDD.n5614 VDD.n5611 593.144
R10658 VDD.n5357 VDD.n5354 593.144
R10659 VDD.n5360 VDD.n5357 593.144
R10660 VDD.n3546 VDD.n3543 593.144
R10661 VDD.n3549 VDD.n3546 593.144
R10662 VDD.n3804 VDD.n3801 593.144
R10663 VDD.n3807 VDD.n3804 593.144
R10664 VDD.n4062 VDD.n4059 593.144
R10665 VDD.n4065 VDD.n4062 593.144
R10666 VDD.n4320 VDD.n4317 593.144
R10667 VDD.n4323 VDD.n4320 593.144
R10668 VDD.n4578 VDD.n4575 593.144
R10669 VDD.n4581 VDD.n4578 593.144
R10670 VDD.n4836 VDD.n4833 593.144
R10671 VDD.n4839 VDD.n4836 593.144
R10672 VDD.n5094 VDD.n5091 593.144
R10673 VDD.n5097 VDD.n5094 593.144
R10674 VDD.n1795 VDD.t445 584.644
R10675 VDD.n1781 VDD.t1035 584.644
R10676 VDD.n2003 VDD.t84 584.644
R10677 VDD.n1989 VDD.t1268 584.644
R10678 VDD.n2374 VDD.t1451 584.644
R10679 VDD.n2360 VDD.t830 584.644
R10680 VDD.n2632 VDD.t573 584.644
R10681 VDD.n2618 VDD.t1424 584.644
R10682 VDD.n2890 VDD.t983 584.644
R10683 VDD.n2876 VDD.t439 584.644
R10684 VDD.n3148 VDD.t550 584.644
R10685 VDD.n3134 VDD.t387 584.644
R10686 VDD.n3406 VDD.t587 584.644
R10687 VDD.n3392 VDD.t1302 584.644
R10688 VDD.n5729 VDD.t1473 584.644
R10689 VDD.n5715 VDD.t480 584.644
R10690 VDD.n5475 VDD.t999 584.644
R10691 VDD.n5461 VDD.t1257 584.644
R10692 VDD.n3664 VDD.t1334 584.644
R10693 VDD.n3650 VDD.t1373 584.644
R10694 VDD.n3922 VDD.t488 584.644
R10695 VDD.n3908 VDD.t1113 584.644
R10696 VDD.n4180 VDD.t9 584.644
R10697 VDD.n4166 VDD.t29 584.644
R10698 VDD.n4438 VDD.t1057 584.644
R10699 VDD.n4424 VDD.t1439 584.644
R10700 VDD.n4696 VDD.t26 584.644
R10701 VDD.n4682 VDD.t374 584.644
R10702 VDD.n4954 VDD.t561 584.644
R10703 VDD.n4940 VDD.t1092 584.644
R10704 VDD.n5212 VDD.t1322 584.644
R10705 VDD.n5198 VDD.t3 584.644
R10706 VDD.n523 VDD.t340 584.644
R10707 VDD.n873 VDD.t1081 584.644
R10708 VDD.n122 VDD.t987 584.644
R10709 VDD.n1348 VDD.t1277 584.644
R10710 VDD.n1763 VDD.n1713 576.668
R10711 VDD.n1763 VDD.n1714 576.668
R10712 VDD.n2112 VDD.n2062 576.668
R10713 VDD.n2112 VDD.n2063 576.668
R10714 VDD.n2342 VDD.n2292 576.668
R10715 VDD.n2342 VDD.n2293 576.668
R10716 VDD.n2600 VDD.n2550 576.668
R10717 VDD.n2600 VDD.n2551 576.668
R10718 VDD.n2858 VDD.n2808 576.668
R10719 VDD.n2858 VDD.n2809 576.668
R10720 VDD.n3116 VDD.n3066 576.668
R10721 VDD.n3116 VDD.n3067 576.668
R10722 VDD.n3374 VDD.n3324 576.668
R10723 VDD.n3374 VDD.n3325 576.668
R10724 VDD.n5697 VDD.n5647 576.668
R10725 VDD.n5697 VDD.n5648 576.668
R10726 VDD.n5443 VDD.n5393 576.668
R10727 VDD.n5443 VDD.n5394 576.668
R10728 VDD.n3632 VDD.n3582 576.668
R10729 VDD.n3632 VDD.n3583 576.668
R10730 VDD.n3890 VDD.n3840 576.668
R10731 VDD.n3890 VDD.n3841 576.668
R10732 VDD.n4148 VDD.n4098 576.668
R10733 VDD.n4148 VDD.n4099 576.668
R10734 VDD.n4406 VDD.n4356 576.668
R10735 VDD.n4406 VDD.n4357 576.668
R10736 VDD.n4664 VDD.n4614 576.668
R10737 VDD.n4664 VDD.n4615 576.668
R10738 VDD.n4922 VDD.n4872 576.668
R10739 VDD.n4922 VDD.n4873 576.668
R10740 VDD.n5180 VDD.n5130 576.668
R10741 VDD.n5180 VDD.n5131 576.668
R10742 VDD.n1906 VDD.n1904 568.236
R10743 VDD.n1899 VDD.n1896 568.236
R10744 VDD.n1902 VDD.n1899 568.236
R10745 VDD.n1904 VDD.n1895 568.236
R10746 VDD.n1859 VDD.n1850 568.236
R10747 VDD.n1862 VDD.n1851 568.236
R10748 VDD.n1864 VDD.n1851 568.236
R10749 VDD.n1855 VDD.n1850 568.236
R10750 VDD.n2180 VDD.n2171 568.236
R10751 VDD.n2183 VDD.n2172 568.236
R10752 VDD.n2185 VDD.n2172 568.236
R10753 VDD.n2176 VDD.n2171 568.236
R10754 VDD.n2227 VDD.n2225 568.236
R10755 VDD.n2220 VDD.n2217 568.236
R10756 VDD.n2223 VDD.n2220 568.236
R10757 VDD.n2225 VDD.n2216 568.236
R10758 VDD.n2438 VDD.n2429 568.236
R10759 VDD.n2441 VDD.n2430 568.236
R10760 VDD.n2443 VDD.n2430 568.236
R10761 VDD.n2434 VDD.n2429 568.236
R10762 VDD.n2485 VDD.n2483 568.236
R10763 VDD.n2478 VDD.n2475 568.236
R10764 VDD.n2481 VDD.n2478 568.236
R10765 VDD.n2483 VDD.n2474 568.236
R10766 VDD.n2696 VDD.n2687 568.236
R10767 VDD.n2699 VDD.n2688 568.236
R10768 VDD.n2701 VDD.n2688 568.236
R10769 VDD.n2692 VDD.n2687 568.236
R10770 VDD.n2743 VDD.n2741 568.236
R10771 VDD.n2736 VDD.n2733 568.236
R10772 VDD.n2739 VDD.n2736 568.236
R10773 VDD.n2741 VDD.n2732 568.236
R10774 VDD.n2954 VDD.n2945 568.236
R10775 VDD.n2957 VDD.n2946 568.236
R10776 VDD.n2959 VDD.n2946 568.236
R10777 VDD.n2950 VDD.n2945 568.236
R10778 VDD.n3001 VDD.n2999 568.236
R10779 VDD.n2994 VDD.n2991 568.236
R10780 VDD.n2997 VDD.n2994 568.236
R10781 VDD.n2999 VDD.n2990 568.236
R10782 VDD.n3212 VDD.n3203 568.236
R10783 VDD.n3215 VDD.n3204 568.236
R10784 VDD.n3217 VDD.n3204 568.236
R10785 VDD.n3208 VDD.n3203 568.236
R10786 VDD.n3259 VDD.n3257 568.236
R10787 VDD.n3252 VDD.n3249 568.236
R10788 VDD.n3255 VDD.n3252 568.236
R10789 VDD.n3257 VDD.n3248 568.236
R10790 VDD.n3470 VDD.n3461 568.236
R10791 VDD.n3473 VDD.n3462 568.236
R10792 VDD.n3475 VDD.n3462 568.236
R10793 VDD.n3466 VDD.n3461 568.236
R10794 VDD.n3517 VDD.n3515 568.236
R10795 VDD.n3510 VDD.n3507 568.236
R10796 VDD.n3513 VDD.n3510 568.236
R10797 VDD.n3515 VDD.n3506 568.236
R10798 VDD.n5790 VDD.n5781 568.236
R10799 VDD.n5793 VDD.n5782 568.236
R10800 VDD.n5795 VDD.n5782 568.236
R10801 VDD.n5786 VDD.n5781 568.236
R10802 VDD.n5837 VDD.n5835 568.236
R10803 VDD.n5830 VDD.n5827 568.236
R10804 VDD.n5833 VDD.n5830 568.236
R10805 VDD.n5835 VDD.n5826 568.236
R10806 VDD.n5536 VDD.n5527 568.236
R10807 VDD.n5539 VDD.n5528 568.236
R10808 VDD.n5541 VDD.n5528 568.236
R10809 VDD.n5532 VDD.n5527 568.236
R10810 VDD.n5583 VDD.n5581 568.236
R10811 VDD.n5576 VDD.n5573 568.236
R10812 VDD.n5579 VDD.n5576 568.236
R10813 VDD.n5581 VDD.n5572 568.236
R10814 VDD.n3728 VDD.n3719 568.236
R10815 VDD.n3731 VDD.n3720 568.236
R10816 VDD.n3733 VDD.n3720 568.236
R10817 VDD.n3724 VDD.n3719 568.236
R10818 VDD.n3775 VDD.n3773 568.236
R10819 VDD.n3768 VDD.n3765 568.236
R10820 VDD.n3771 VDD.n3768 568.236
R10821 VDD.n3773 VDD.n3764 568.236
R10822 VDD.n3986 VDD.n3977 568.236
R10823 VDD.n3989 VDD.n3978 568.236
R10824 VDD.n3991 VDD.n3978 568.236
R10825 VDD.n3982 VDD.n3977 568.236
R10826 VDD.n4033 VDD.n4031 568.236
R10827 VDD.n4026 VDD.n4023 568.236
R10828 VDD.n4029 VDD.n4026 568.236
R10829 VDD.n4031 VDD.n4022 568.236
R10830 VDD.n4244 VDD.n4235 568.236
R10831 VDD.n4247 VDD.n4236 568.236
R10832 VDD.n4249 VDD.n4236 568.236
R10833 VDD.n4240 VDD.n4235 568.236
R10834 VDD.n4291 VDD.n4289 568.236
R10835 VDD.n4284 VDD.n4281 568.236
R10836 VDD.n4287 VDD.n4284 568.236
R10837 VDD.n4289 VDD.n4280 568.236
R10838 VDD.n4502 VDD.n4493 568.236
R10839 VDD.n4505 VDD.n4494 568.236
R10840 VDD.n4507 VDD.n4494 568.236
R10841 VDD.n4498 VDD.n4493 568.236
R10842 VDD.n4549 VDD.n4547 568.236
R10843 VDD.n4542 VDD.n4539 568.236
R10844 VDD.n4545 VDD.n4542 568.236
R10845 VDD.n4547 VDD.n4538 568.236
R10846 VDD.n4760 VDD.n4751 568.236
R10847 VDD.n4763 VDD.n4752 568.236
R10848 VDD.n4765 VDD.n4752 568.236
R10849 VDD.n4756 VDD.n4751 568.236
R10850 VDD.n4807 VDD.n4805 568.236
R10851 VDD.n4800 VDD.n4797 568.236
R10852 VDD.n4803 VDD.n4800 568.236
R10853 VDD.n4805 VDD.n4796 568.236
R10854 VDD.n5018 VDD.n5009 568.236
R10855 VDD.n5021 VDD.n5010 568.236
R10856 VDD.n5023 VDD.n5010 568.236
R10857 VDD.n5014 VDD.n5009 568.236
R10858 VDD.n5065 VDD.n5063 568.236
R10859 VDD.n5058 VDD.n5055 568.236
R10860 VDD.n5061 VDD.n5058 568.236
R10861 VDD.n5063 VDD.n5054 568.236
R10862 VDD.n5276 VDD.n5267 568.236
R10863 VDD.n5279 VDD.n5268 568.236
R10864 VDD.n5281 VDD.n5268 568.236
R10865 VDD.n5272 VDD.n5267 568.236
R10866 VDD.n5323 VDD.n5321 568.236
R10867 VDD.n5316 VDD.n5313 568.236
R10868 VDD.n5319 VDD.n5316 568.236
R10869 VDD.n5321 VDD.n5312 568.236
R10870 VDD.n857 VDD.t354 533.735
R10871 VDD.n1240 VDD.t798 533.735
R10872 VDD.n1744 VDD.n1743 481.226
R10873 VDD.n2093 VDD.n2092 481.226
R10874 VDD.n2323 VDD.n2322 481.226
R10875 VDD.n2581 VDD.n2580 481.226
R10876 VDD.n2839 VDD.n2838 481.226
R10877 VDD.n3097 VDD.n3096 481.226
R10878 VDD.n3355 VDD.n3354 481.226
R10879 VDD.n5678 VDD.n5677 481.226
R10880 VDD.n5424 VDD.n5423 481.226
R10881 VDD.n3613 VDD.n3612 481.226
R10882 VDD.n3871 VDD.n3870 481.226
R10883 VDD.n4129 VDD.n4128 481.226
R10884 VDD.n4387 VDD.n4386 481.226
R10885 VDD.n4645 VDD.n4644 481.226
R10886 VDD.n4903 VDD.n4902 481.226
R10887 VDD.n5161 VDD.n5160 481.226
R10888 VDD.n1857 VDD.n1847 473.839
R10889 VDD.t466 VDD.n1849 473.839
R10890 VDD.n2178 VDD.n2168 473.839
R10891 VDD.t592 VDD.n2170 473.839
R10892 VDD.n2436 VDD.n2426 473.839
R10893 VDD.t521 VDD.n2428 473.839
R10894 VDD.n2694 VDD.n2684 473.839
R10895 VDD.t278 VDD.n2686 473.839
R10896 VDD.n2952 VDD.n2942 473.839
R10897 VDD.t368 VDD.n2944 473.839
R10898 VDD.n3210 VDD.n3200 473.839
R10899 VDD.t1087 VDD.n3202 473.839
R10900 VDD.n3468 VDD.n3458 473.839
R10901 VDD.t1093 VDD.n3460 473.839
R10902 VDD.n5788 VDD.n5778 473.839
R10903 VDD.t514 VDD.n5780 473.839
R10904 VDD.n5534 VDD.n5524 473.839
R10905 VDD.t507 VDD.n5526 473.839
R10906 VDD.n3726 VDD.n3716 473.839
R10907 VDD.t251 VDD.n3718 473.839
R10908 VDD.n3984 VDD.n3974 473.839
R10909 VDD.t266 VDD.n3976 473.839
R10910 VDD.n4242 VDD.n4232 473.839
R10911 VDD.t13 VDD.n4234 473.839
R10912 VDD.n4500 VDD.n4490 473.839
R10913 VDD.t415 VDD.n4492 473.839
R10914 VDD.n4758 VDD.n4748 473.839
R10915 VDD.t527 VDD.n4750 473.839
R10916 VDD.n5016 VDD.n5006 473.839
R10917 VDD.t815 VDD.n5008 473.839
R10918 VDD.n5274 VDD.n5264 473.839
R10919 VDD.t265 VDD.n5266 473.839
R10920 VDD.n1914 VDD.n1892 468.033
R10921 VDD.t277 VDD.n1893 468.033
R10922 VDD.n2235 VDD.n2213 468.033
R10923 VDD.t494 VDD.n2214 468.033
R10924 VDD.n2493 VDD.n2471 468.033
R10925 VDD.t505 VDD.n2472 468.033
R10926 VDD.n2751 VDD.n2729 468.033
R10927 VDD.t1023 VDD.n2730 468.033
R10928 VDD.n3009 VDD.n2987 468.033
R10929 VDD.t524 VDD.n2988 468.033
R10930 VDD.n3267 VDD.n3245 468.033
R10931 VDD.t282 VDD.n3246 468.033
R10932 VDD.n3525 VDD.n3503 468.033
R10933 VDD.t419 VDD.n3504 468.033
R10934 VDD.n5845 VDD.n5823 468.033
R10935 VDD.t1075 VDD.n5824 468.033
R10936 VDD.n5591 VDD.n5569 468.033
R10937 VDD.t393 VDD.n5570 468.033
R10938 VDD.n3783 VDD.n3761 468.033
R10939 VDD.t262 VDD.n3762 468.033
R10940 VDD.n4041 VDD.n4019 468.033
R10941 VDD.t1084 VDD.n4020 468.033
R10942 VDD.n4299 VDD.n4277 468.033
R10943 VDD.t1021 VDD.n4278 468.033
R10944 VDD.n4557 VDD.n4535 468.033
R10945 VDD.t531 VDD.n4536 468.033
R10946 VDD.n4815 VDD.n4793 468.033
R10947 VDD.t401 VDD.n4794 468.033
R10948 VDD.n5073 VDD.n5051 468.033
R10949 VDD.t416 VDD.n5052 468.033
R10950 VDD.n5331 VDD.n5309 468.033
R10951 VDD.t407 VDD.n5310 468.033
R10952 VDD.n1933 VDD.n1925 459.009
R10953 VDD.n1935 VDD.n1932 437.647
R10954 VDD.n1974 VDD.n1928 430.589
R10955 VDD.n1962 VDD.n1940 430.589
R10956 VDD.n483 VDD.n482 425.228
R10957 VDD.n81 VDD.n80 425.228
R10958 VDD VDD.t536 421.082
R10959 VDD.n1948 VDD.n1938 420
R10960 VDD.n407 VDD.t611 396.079
R10961 VDD.n1565 VDD.t1491 396.079
R10962 VDD.n9 VDD.t359 382.793
R10963 VDD.n465 VDD.t352 382.793
R10964 VDD.n412 VDD.t363 382.793
R10965 VDD.n411 VDD.t349 382.793
R10966 VDD.n393 VDD.t348 382.793
R10967 VDD.n63 VDD.t802 382.793
R10968 VDD.n1153 VDD.t811 382.793
R10969 VDD.n1570 VDD.t796 382.793
R10970 VDD.n1569 VDD.t792 382.793
R10971 VDD.n1551 VDD.t789 382.793
R10972 VDD.n805 VDD.t614 382.793
R10973 VDD.n1188 VDD.t535 382.793
R10974 VDD VDD.t1319 374.711
R10975 VDD VDD.t1314 374.711
R10976 VDD VDD.t330 374.711
R10977 VDD VDD.t1311 374.711
R10978 VDD VDD.t1360 374.711
R10979 VDD VDD.t969 374.711
R10980 VDD.n1709 VDD.n1680 370.589
R10981 VDD.n1759 VDD.n1714 370.589
R10982 VDD.n2058 VDD.n2029 370.589
R10983 VDD.n2108 VDD.n2063 370.589
R10984 VDD.n2288 VDD.n2259 370.589
R10985 VDD.n2338 VDD.n2293 370.589
R10986 VDD.n2546 VDD.n2517 370.589
R10987 VDD.n2596 VDD.n2551 370.589
R10988 VDD.n2804 VDD.n2775 370.589
R10989 VDD.n2854 VDD.n2809 370.589
R10990 VDD.n3062 VDD.n3033 370.589
R10991 VDD.n3112 VDD.n3067 370.589
R10992 VDD.n3320 VDD.n3291 370.589
R10993 VDD.n3370 VDD.n3325 370.589
R10994 VDD.n5643 VDD.n5614 370.589
R10995 VDD.n5693 VDD.n5648 370.589
R10996 VDD.n5389 VDD.n5360 370.589
R10997 VDD.n5439 VDD.n5394 370.589
R10998 VDD.n3578 VDD.n3549 370.589
R10999 VDD.n3628 VDD.n3583 370.589
R11000 VDD.n3836 VDD.n3807 370.589
R11001 VDD.n3886 VDD.n3841 370.589
R11002 VDD.n4094 VDD.n4065 370.589
R11003 VDD.n4144 VDD.n4099 370.589
R11004 VDD.n4352 VDD.n4323 370.589
R11005 VDD.n4402 VDD.n4357 370.589
R11006 VDD.n4610 VDD.n4581 370.589
R11007 VDD.n4660 VDD.n4615 370.589
R11008 VDD.n4868 VDD.n4839 370.589
R11009 VDD.n4918 VDD.n4873 370.589
R11010 VDD.n5126 VDD.n5097 370.589
R11011 VDD.n5176 VDD.n5131 370.589
R11012 VDD.n12 VDD.t1065 370.341
R11013 VDD.n473 VDD.t353 370.341
R11014 VDD.n445 VDD.t1292 370.341
R11015 VDD.n446 VDD.t76 370.341
R11016 VDD.n71 VDD.t805 370.341
R11017 VDD.n42 VDD.t427 370.341
R11018 VDD.n43 VDD.t632 370.341
R11019 VDD.n1156 VDD.t972 370.341
R11020 VDD VDD.t1343 370.303
R11021 VDD VDD.t1374 370.303
R11022 VDD.t1014 VDD.t1031 333.365
R11023 VDD.t1014 VDD.t441 333.365
R11024 VDD.t623 VDD.t1264 333.365
R11025 VDD.t623 VDD.t80 333.365
R11026 VDD.t1331 VDD.t831 333.365
R11027 VDD.t1331 VDD.t1446 333.365
R11028 VDD.t825 VDD.t1417 333.365
R11029 VDD.t825 VDD.t567 333.365
R11030 VDD.t424 VDD.t436 333.365
R11031 VDD.t424 VDD.t978 333.365
R11032 VDD.t395 VDD.t383 333.365
R11033 VDD.t395 VDD.t545 333.365
R11034 VDD.t639 VDD.t1295 333.365
R11035 VDD.t639 VDD.t582 333.365
R11036 VDD.t1307 VDD.t476 333.365
R11037 VDD.t1307 VDD.t1468 333.365
R11038 VDD.t270 VDD.t1258 333.365
R11039 VDD.t270 VDD.t995 333.365
R11040 VDD.t249 VDD.t1366 333.365
R11041 VDD.t249 VDD.t1336 333.365
R11042 VDD.t1317 VDD.t1114 333.365
R11043 VDD.t1317 VDD.t485 333.365
R11044 VDD.t409 VDD.t30 333.365
R11045 VDD.t409 VDD.t5 333.365
R11046 VDD.t1108 VDD.t1436 333.365
R11047 VDD.t1108 VDD.t1052 333.365
R11048 VDD.t332 VDD.t370 333.365
R11049 VDD.t332 VDD.t21 333.365
R11050 VDD.t279 VDD.t422 333.365
R11051 VDD.t279 VDD.t563 333.365
R11052 VDD.t1060 VDD.t0 333.365
R11053 VDD.t1060 VDD.t1008 333.365
R11054 VDD VDD.t974 331.981
R11055 VDD VDD.t381 331.981
R11056 VDD.n1634 VDD.t812 330.12
R11057 VDD.n1635 VDD.t793 330.002
R11058 VDD.n1541 VDD 323.514
R11059 VDD.n1643 VDD.t803 323.342
R11060 VDD.n34 VDD.t1454 321.801
R11061 VDD.n1178 VDD.t498 321.801
R11062 VDD.n476 VDD.n475 318.678
R11063 VDD.n74 VDD.n73 318.678
R11064 VDD.n511 VDD.t411 318.108
R11065 VDD.n109 VDD.t429 318.108
R11066 VDD VDD.t1046 313.839
R11067 VDD VDD.t1431 313.839
R11068 VDD VDD.t596 313.839
R11069 VDD.n8 VDD.n7 307.24
R11070 VDD.n472 VDD.n471 307.24
R11071 VDD.n442 VDD.n441 307.24
R11072 VDD.n444 VDD.n443 307.24
R11073 VDD.n70 VDD.n69 307.24
R11074 VDD.n39 VDD.n38 307.24
R11075 VDD.n41 VDD.n40 307.24
R11076 VDD.n1152 VDD.n1151 307.24
R11077 VDD.t1014 VDD.n1678 298.82
R11078 VDD.t1014 VDD.n1712 298.82
R11079 VDD.t623 VDD.n2027 298.82
R11080 VDD.t623 VDD.n2061 298.82
R11081 VDD.t1331 VDD.n2257 298.82
R11082 VDD.t1331 VDD.n2291 298.82
R11083 VDD.t825 VDD.n2515 298.82
R11084 VDD.t825 VDD.n2549 298.82
R11085 VDD.t424 VDD.n2773 298.82
R11086 VDD.t424 VDD.n2807 298.82
R11087 VDD.t395 VDD.n3031 298.82
R11088 VDD.t395 VDD.n3065 298.82
R11089 VDD.t639 VDD.n3289 298.82
R11090 VDD.t639 VDD.n3323 298.82
R11091 VDD.t1307 VDD.n5612 298.82
R11092 VDD.t1307 VDD.n5646 298.82
R11093 VDD.t270 VDD.n5358 298.82
R11094 VDD.t270 VDD.n5392 298.82
R11095 VDD.t249 VDD.n3547 298.82
R11096 VDD.t249 VDD.n3581 298.82
R11097 VDD.t1317 VDD.n3805 298.82
R11098 VDD.t1317 VDD.n3839 298.82
R11099 VDD.t409 VDD.n4063 298.82
R11100 VDD.t409 VDD.n4097 298.82
R11101 VDD.t1108 VDD.n4321 298.82
R11102 VDD.t1108 VDD.n4355 298.82
R11103 VDD.t332 VDD.n4579 298.82
R11104 VDD.t332 VDD.n4613 298.82
R11105 VDD.t279 VDD.n4837 298.82
R11106 VDD.t279 VDD.n4871 298.82
R11107 VDD.t1060 VDD.n5095 298.82
R11108 VDD.t1060 VDD.n5129 298.82
R11109 VDD.n1912 VDD.n1897 273.695
R11110 VDD.n1912 VDD.n1911 273.695
R11111 VDD.n1877 VDD.n1824 273.695
R11112 VDD.n1824 VDD.n1822 273.695
R11113 VDD.n1861 VDD.n1860 273.695
R11114 VDD.n1865 VDD.n1861 273.695
R11115 VDD.n2182 VDD.n2181 273.695
R11116 VDD.n2186 VDD.n2182 273.695
R11117 VDD.n2198 VDD.n2145 273.695
R11118 VDD.n2145 VDD.n2143 273.695
R11119 VDD.n2233 VDD.n2218 273.695
R11120 VDD.n2233 VDD.n2232 273.695
R11121 VDD.n2440 VDD.n2439 273.695
R11122 VDD.n2444 VDD.n2440 273.695
R11123 VDD.n2456 VDD.n2403 273.695
R11124 VDD.n2403 VDD.n2401 273.695
R11125 VDD.n2491 VDD.n2476 273.695
R11126 VDD.n2491 VDD.n2490 273.695
R11127 VDD.n2698 VDD.n2697 273.695
R11128 VDD.n2702 VDD.n2698 273.695
R11129 VDD.n2714 VDD.n2661 273.695
R11130 VDD.n2661 VDD.n2659 273.695
R11131 VDD.n2749 VDD.n2734 273.695
R11132 VDD.n2749 VDD.n2748 273.695
R11133 VDD.n2956 VDD.n2955 273.695
R11134 VDD.n2960 VDD.n2956 273.695
R11135 VDD.n2972 VDD.n2919 273.695
R11136 VDD.n2919 VDD.n2917 273.695
R11137 VDD.n3007 VDD.n2992 273.695
R11138 VDD.n3007 VDD.n3006 273.695
R11139 VDD.n3214 VDD.n3213 273.695
R11140 VDD.n3218 VDD.n3214 273.695
R11141 VDD.n3230 VDD.n3177 273.695
R11142 VDD.n3177 VDD.n3175 273.695
R11143 VDD.n3265 VDD.n3250 273.695
R11144 VDD.n3265 VDD.n3264 273.695
R11145 VDD.n3472 VDD.n3471 273.695
R11146 VDD.n3476 VDD.n3472 273.695
R11147 VDD.n3488 VDD.n3435 273.695
R11148 VDD.n3435 VDD.n3433 273.695
R11149 VDD.n3523 VDD.n3508 273.695
R11150 VDD.n3523 VDD.n3522 273.695
R11151 VDD.n5792 VDD.n5791 273.695
R11152 VDD.n5796 VDD.n5792 273.695
R11153 VDD.n5808 VDD.n5755 273.695
R11154 VDD.n5755 VDD.n5753 273.695
R11155 VDD.n5843 VDD.n5828 273.695
R11156 VDD.n5843 VDD.n5842 273.695
R11157 VDD.n5538 VDD.n5537 273.695
R11158 VDD.n5542 VDD.n5538 273.695
R11159 VDD.n5554 VDD.n5501 273.695
R11160 VDD.n5501 VDD.n5499 273.695
R11161 VDD.n5589 VDD.n5574 273.695
R11162 VDD.n5589 VDD.n5588 273.695
R11163 VDD.n3730 VDD.n3729 273.695
R11164 VDD.n3734 VDD.n3730 273.695
R11165 VDD.n3746 VDD.n3693 273.695
R11166 VDD.n3693 VDD.n3691 273.695
R11167 VDD.n3781 VDD.n3766 273.695
R11168 VDD.n3781 VDD.n3780 273.695
R11169 VDD.n3988 VDD.n3987 273.695
R11170 VDD.n3992 VDD.n3988 273.695
R11171 VDD.n4004 VDD.n3951 273.695
R11172 VDD.n3951 VDD.n3949 273.695
R11173 VDD.n4039 VDD.n4024 273.695
R11174 VDD.n4039 VDD.n4038 273.695
R11175 VDD.n4246 VDD.n4245 273.695
R11176 VDD.n4250 VDD.n4246 273.695
R11177 VDD.n4262 VDD.n4209 273.695
R11178 VDD.n4209 VDD.n4207 273.695
R11179 VDD.n4297 VDD.n4282 273.695
R11180 VDD.n4297 VDD.n4296 273.695
R11181 VDD.n4504 VDD.n4503 273.695
R11182 VDD.n4508 VDD.n4504 273.695
R11183 VDD.n4520 VDD.n4467 273.695
R11184 VDD.n4467 VDD.n4465 273.695
R11185 VDD.n4555 VDD.n4540 273.695
R11186 VDD.n4555 VDD.n4554 273.695
R11187 VDD.n4762 VDD.n4761 273.695
R11188 VDD.n4766 VDD.n4762 273.695
R11189 VDD.n4778 VDD.n4725 273.695
R11190 VDD.n4725 VDD.n4723 273.695
R11191 VDD.n4813 VDD.n4798 273.695
R11192 VDD.n4813 VDD.n4812 273.695
R11193 VDD.n5020 VDD.n5019 273.695
R11194 VDD.n5024 VDD.n5020 273.695
R11195 VDD.n5036 VDD.n4983 273.695
R11196 VDD.n4983 VDD.n4981 273.695
R11197 VDD.n5071 VDD.n5056 273.695
R11198 VDD.n5071 VDD.n5070 273.695
R11199 VDD.n5278 VDD.n5277 273.695
R11200 VDD.n5282 VDD.n5278 273.695
R11201 VDD.n5294 VDD.n5241 273.695
R11202 VDD.n5241 VDD.n5239 273.695
R11203 VDD.n5329 VDD.n5314 273.695
R11204 VDD.n5329 VDD.n5328 273.695
R11205 VDD.n1616 VDD.t806 260.435
R11206 VDD.n1624 VDD.t787 256.07
R11207 VDD.n1627 VDD.t790 256.07
R11208 VDD.n1629 VDD.t795 256.07
R11209 VDD.n1632 VDD.t809 256.07
R11210 VDD.n1649 VDD.t800 251.637
R11211 VDD.t974 VDD.t360 246.023
R11212 VDD.t381 VDD.t813 246.023
R11213 VDD VDD.t335 241.819
R11214 VDD VDD.t502 241.819
R11215 VDD.t354 VDD 233.643
R11216 VDD.t1319 VDD 233.643
R11217 VDD.t1314 VDD 233.643
R11218 VDD.t1343 VDD 233.643
R11219 VDD.t330 VDD 233.643
R11220 VDD.t798 VDD 233.643
R11221 VDD.t1311 VDD 233.643
R11222 VDD.t1360 VDD 233.643
R11223 VDD.t1374 VDD 233.643
R11224 VDD.t969 VDD 233.643
R11225 VDD.n1605 VDD.t797 229.433
R11226 VDD.t103 VDD 227.321
R11227 VDD VDD.t91 227.321
R11228 VDD.t169 VDD 227.321
R11229 VDD.t1397 VDD 227.321
R11230 VDD.t876 VDD 227.321
R11231 VDD VDD.t864 227.321
R11232 VDD.t944 VDD 227.321
R11233 VDD.t53 VDD 227.321
R11234 VDD.t656 VDD 227.321
R11235 VDD VDD.t772 227.321
R11236 VDD.t722 VDD 227.321
R11237 VDD.t227 VDD 227.321
R11238 VDD.t339 VDD 225.625
R11239 VDD.t1080 VDD 225.625
R11240 VDD.t986 VDD 225.625
R11241 VDD.n1909 VDD.n1908 213.083
R11242 VDD.n1910 VDD.n1909 213.083
R11243 VDD.n1867 VDD.n1852 213.083
R11244 VDD.n1867 VDD.n1866 213.083
R11245 VDD.n2188 VDD.n2173 213.083
R11246 VDD.n2188 VDD.n2187 213.083
R11247 VDD.n2230 VDD.n2229 213.083
R11248 VDD.n2231 VDD.n2230 213.083
R11249 VDD.n2446 VDD.n2431 213.083
R11250 VDD.n2446 VDD.n2445 213.083
R11251 VDD.n2488 VDD.n2487 213.083
R11252 VDD.n2489 VDD.n2488 213.083
R11253 VDD.n2704 VDD.n2689 213.083
R11254 VDD.n2704 VDD.n2703 213.083
R11255 VDD.n2746 VDD.n2745 213.083
R11256 VDD.n2747 VDD.n2746 213.083
R11257 VDD.n2962 VDD.n2947 213.083
R11258 VDD.n2962 VDD.n2961 213.083
R11259 VDD.n3004 VDD.n3003 213.083
R11260 VDD.n3005 VDD.n3004 213.083
R11261 VDD.n3220 VDD.n3205 213.083
R11262 VDD.n3220 VDD.n3219 213.083
R11263 VDD.n3262 VDD.n3261 213.083
R11264 VDD.n3263 VDD.n3262 213.083
R11265 VDD.n3478 VDD.n3463 213.083
R11266 VDD.n3478 VDD.n3477 213.083
R11267 VDD.n3520 VDD.n3519 213.083
R11268 VDD.n3521 VDD.n3520 213.083
R11269 VDD.n5798 VDD.n5783 213.083
R11270 VDD.n5798 VDD.n5797 213.083
R11271 VDD.n5840 VDD.n5839 213.083
R11272 VDD.n5841 VDD.n5840 213.083
R11273 VDD.n5544 VDD.n5529 213.083
R11274 VDD.n5544 VDD.n5543 213.083
R11275 VDD.n5586 VDD.n5585 213.083
R11276 VDD.n5587 VDD.n5586 213.083
R11277 VDD.n3736 VDD.n3721 213.083
R11278 VDD.n3736 VDD.n3735 213.083
R11279 VDD.n3778 VDD.n3777 213.083
R11280 VDD.n3779 VDD.n3778 213.083
R11281 VDD.n3994 VDD.n3979 213.083
R11282 VDD.n3994 VDD.n3993 213.083
R11283 VDD.n4036 VDD.n4035 213.083
R11284 VDD.n4037 VDD.n4036 213.083
R11285 VDD.n4252 VDD.n4237 213.083
R11286 VDD.n4252 VDD.n4251 213.083
R11287 VDD.n4294 VDD.n4293 213.083
R11288 VDD.n4295 VDD.n4294 213.083
R11289 VDD.n4510 VDD.n4495 213.083
R11290 VDD.n4510 VDD.n4509 213.083
R11291 VDD.n4552 VDD.n4551 213.083
R11292 VDD.n4553 VDD.n4552 213.083
R11293 VDD.n4768 VDD.n4753 213.083
R11294 VDD.n4768 VDD.n4767 213.083
R11295 VDD.n4810 VDD.n4809 213.083
R11296 VDD.n4811 VDD.n4810 213.083
R11297 VDD.n5026 VDD.n5011 213.083
R11298 VDD.n5026 VDD.n5025 213.083
R11299 VDD.n5068 VDD.n5067 213.083
R11300 VDD.n5069 VDD.n5068 213.083
R11301 VDD.n5284 VDD.n5269 213.083
R11302 VDD.n5284 VDD.n5283 213.083
R11303 VDD.n5326 VDD.n5325 213.083
R11304 VDD.n5327 VDD.n5326 213.083
R11305 VDD.n531 VDD.t102 204.903
R11306 VDD.n881 VDD.t875 204.903
R11307 VDD.n130 VDD.t655 204.903
R11308 VDD.n1249 VDD.t1241 204.9
R11309 VDD.n1634 VDD.t1509 201.587
R11310 VDD.n542 VDD.t104 201.012
R11311 VDD.n621 VDD.t92 201.012
R11312 VDD.n517 VDD.t170 201.012
R11313 VDD.n520 VDD.t1398 201.012
R11314 VDD.n892 VDD.t877 201.012
R11315 VDD.n971 VDD.t865 201.012
R11316 VDD.n867 VDD.t945 201.012
R11317 VDD.n870 VDD.t54 201.012
R11318 VDD.n141 VDD.t657 201.012
R11319 VDD.n220 VDD.t773 201.012
R11320 VDD.n116 VDD.t723 201.012
R11321 VDD.n119 VDD.t228 201.012
R11322 VDD.n1313 VDD.t1147 201.012
R11323 VDD.n1342 VDD.t319 201.012
R11324 VDD.n1263 VDD.t1129 201.012
R11325 VDD.n1260 VDD.t1227 201.012
R11326 VDD.n1635 VDD.t1507 200.782
R11327 VDD.n1643 VDD.t1503 194.809
R11328 VDD.n1901 VDD.n1893 189.304
R11329 VDD.n2222 VDD.n2214 189.304
R11330 VDD.n2480 VDD.n2472 189.304
R11331 VDD.n2738 VDD.n2730 189.304
R11332 VDD.n2996 VDD.n2988 189.304
R11333 VDD.n3254 VDD.n3246 189.304
R11334 VDD.n3512 VDD.n3504 189.304
R11335 VDD.n5832 VDD.n5824 189.304
R11336 VDD.n5578 VDD.n5570 189.304
R11337 VDD.n3770 VDD.n3762 189.304
R11338 VDD.n4028 VDD.n4020 189.304
R11339 VDD.n4286 VDD.n4278 189.304
R11340 VDD.n4544 VDD.n4536 189.304
R11341 VDD.n4802 VDD.n4794 189.304
R11342 VDD.n5060 VDD.n5052 189.304
R11343 VDD.n5318 VDD.n5310 189.304
R11344 VDD.n1954 VDD.n1939 185
R11345 VDD.n1900 VDD.n1898 185
R11346 VDD.n1900 VDD.n1893 185
R11347 VDD.n1890 VDD.n1888 185
R11348 VDD.n1892 VDD.n1890 185
R11349 VDD.n1697 VDD.n1682 185
R11350 VDD.n2046 VDD.n2031 185
R11351 VDD.n2221 VDD.n2219 185
R11352 VDD.n2221 VDD.n2214 185
R11353 VDD.n2211 VDD.n2209 185
R11354 VDD.n2213 VDD.n2211 185
R11355 VDD.n2276 VDD.n2261 185
R11356 VDD.n2479 VDD.n2477 185
R11357 VDD.n2479 VDD.n2472 185
R11358 VDD.n2469 VDD.n2467 185
R11359 VDD.n2471 VDD.n2469 185
R11360 VDD.n2534 VDD.n2519 185
R11361 VDD.n2737 VDD.n2735 185
R11362 VDD.n2737 VDD.n2730 185
R11363 VDD.n2727 VDD.n2725 185
R11364 VDD.n2729 VDD.n2727 185
R11365 VDD.n2792 VDD.n2777 185
R11366 VDD.n2995 VDD.n2993 185
R11367 VDD.n2995 VDD.n2988 185
R11368 VDD.n2985 VDD.n2983 185
R11369 VDD.n2987 VDD.n2985 185
R11370 VDD.n3050 VDD.n3035 185
R11371 VDD.n3253 VDD.n3251 185
R11372 VDD.n3253 VDD.n3246 185
R11373 VDD.n3243 VDD.n3241 185
R11374 VDD.n3245 VDD.n3243 185
R11375 VDD.n3308 VDD.n3293 185
R11376 VDD.n3511 VDD.n3509 185
R11377 VDD.n3511 VDD.n3504 185
R11378 VDD.n3501 VDD.n3499 185
R11379 VDD.n3503 VDD.n3501 185
R11380 VDD.n5631 VDD.n5616 185
R11381 VDD.n5831 VDD.n5829 185
R11382 VDD.n5831 VDD.n5824 185
R11383 VDD.n5821 VDD.n5819 185
R11384 VDD.n5823 VDD.n5821 185
R11385 VDD.n5377 VDD.n5362 185
R11386 VDD.n5577 VDD.n5575 185
R11387 VDD.n5577 VDD.n5570 185
R11388 VDD.n5567 VDD.n5565 185
R11389 VDD.n5569 VDD.n5567 185
R11390 VDD.n3566 VDD.n3551 185
R11391 VDD.n3769 VDD.n3767 185
R11392 VDD.n3769 VDD.n3762 185
R11393 VDD.n3759 VDD.n3757 185
R11394 VDD.n3761 VDD.n3759 185
R11395 VDD.n3824 VDD.n3809 185
R11396 VDD.n4027 VDD.n4025 185
R11397 VDD.n4027 VDD.n4020 185
R11398 VDD.n4017 VDD.n4015 185
R11399 VDD.n4019 VDD.n4017 185
R11400 VDD.n4082 VDD.n4067 185
R11401 VDD.n4285 VDD.n4283 185
R11402 VDD.n4285 VDD.n4278 185
R11403 VDD.n4275 VDD.n4273 185
R11404 VDD.n4277 VDD.n4275 185
R11405 VDD.n4340 VDD.n4325 185
R11406 VDD.n4543 VDD.n4541 185
R11407 VDD.n4543 VDD.n4536 185
R11408 VDD.n4533 VDD.n4531 185
R11409 VDD.n4535 VDD.n4533 185
R11410 VDD.n4598 VDD.n4583 185
R11411 VDD.n4801 VDD.n4799 185
R11412 VDD.n4801 VDD.n4794 185
R11413 VDD.n4791 VDD.n4789 185
R11414 VDD.n4793 VDD.n4791 185
R11415 VDD.n4856 VDD.n4841 185
R11416 VDD.n5059 VDD.n5057 185
R11417 VDD.n5059 VDD.n5052 185
R11418 VDD.n5049 VDD.n5047 185
R11419 VDD.n5051 VDD.n5049 185
R11420 VDD.n5114 VDD.n5099 185
R11421 VDD.n5317 VDD.n5315 185
R11422 VDD.n5317 VDD.n5310 185
R11423 VDD.n5307 VDD.n5305 185
R11424 VDD.n5309 VDD.n5307 185
R11425 VDD.n1863 VDD.n1849 183.496
R11426 VDD.n2184 VDD.n2170 183.496
R11427 VDD.n2442 VDD.n2428 183.496
R11428 VDD.n2700 VDD.n2686 183.496
R11429 VDD.n2958 VDD.n2944 183.496
R11430 VDD.n3216 VDD.n3202 183.496
R11431 VDD.n3474 VDD.n3460 183.496
R11432 VDD.n5794 VDD.n5780 183.496
R11433 VDD.n5540 VDD.n5526 183.496
R11434 VDD.n3732 VDD.n3718 183.496
R11435 VDD.n3990 VDD.n3976 183.496
R11436 VDD.n4248 VDD.n4234 183.496
R11437 VDD.n4506 VDD.n4492 183.496
R11438 VDD.n4764 VDD.n4750 183.496
R11439 VDD.n5022 VDD.n5008 183.496
R11440 VDD.n5280 VDD.n5266 183.496
R11441 VDD.n807 VDD.n806 183.363
R11442 VDD.n1190 VDD.n1189 183.363
R11443 VDD.n1793 VDD.n1792 180.994
R11444 VDD.n1790 VDD.n1788 180.994
R11445 VDD.n2001 VDD.n2000 180.994
R11446 VDD.n1998 VDD.n1996 180.994
R11447 VDD.n2372 VDD.n2371 180.994
R11448 VDD.n2369 VDD.n2367 180.994
R11449 VDD.n2630 VDD.n2629 180.994
R11450 VDD.n2627 VDD.n2625 180.994
R11451 VDD.n2888 VDD.n2887 180.994
R11452 VDD.n2885 VDD.n2883 180.994
R11453 VDD.n3146 VDD.n3145 180.994
R11454 VDD.n3143 VDD.n3141 180.994
R11455 VDD.n3404 VDD.n3403 180.994
R11456 VDD.n3401 VDD.n3399 180.994
R11457 VDD.n5727 VDD.n5726 180.994
R11458 VDD.n5724 VDD.n5722 180.994
R11459 VDD.n5473 VDD.n5472 180.994
R11460 VDD.n5470 VDD.n5468 180.994
R11461 VDD.n3662 VDD.n3661 180.994
R11462 VDD.n3659 VDD.n3657 180.994
R11463 VDD.n3920 VDD.n3919 180.994
R11464 VDD.n3917 VDD.n3915 180.994
R11465 VDD.n4178 VDD.n4177 180.994
R11466 VDD.n4175 VDD.n4173 180.994
R11467 VDD.n4436 VDD.n4435 180.994
R11468 VDD.n4433 VDD.n4431 180.994
R11469 VDD.n4694 VDD.n4693 180.994
R11470 VDD.n4691 VDD.n4689 180.994
R11471 VDD.n4952 VDD.n4951 180.994
R11472 VDD.n4949 VDD.n4947 180.994
R11473 VDD.n5210 VDD.n5209 180.994
R11474 VDD.n5207 VDD.n5205 180.994
R11475 VDD.t780 VDD 179.821
R11476 VDD.t1045 VDD 179.821
R11477 VDD.t1484 VDD 179.821
R11478 VDD.t819 VDD 179.821
R11479 VDD.n265 VDD.t379 179.821
R11480 VDD.t379 VDD 179.821
R11481 VDD.t1290 VDD 179.821
R11482 VDD.n19 VDD.n5 179.131
R11483 VDD.n495 VDD.n494 179.131
R11484 VDD.n423 VDD.n422 179.131
R11485 VDD.n419 VDD.n418 179.131
R11486 VDD.n402 VDD.n401 179.131
R11487 VDD.n93 VDD.n92 179.131
R11488 VDD.n1163 VDD.n1149 179.131
R11489 VDD.n1581 VDD.n1580 179.131
R11490 VDD.n1577 VDD.n1576 179.131
R11491 VDD.n1560 VDD.n1559 179.131
R11492 VDD.t1028 VDD.n1803 174.632
R11493 VDD.t1266 VDD.n2011 174.632
R11494 VDD.t828 VDD.n2382 174.632
R11495 VDD.t1419 VDD.n2640 174.632
R11496 VDD.t433 VDD.n2898 174.632
R11497 VDD.t385 VDD.n3156 174.632
R11498 VDD.t1297 VDD.n3414 174.632
R11499 VDD.t473 VDD.n5737 174.632
R11500 VDD.t1256 VDD.n5483 174.632
R11501 VDD.t1368 VDD.n3672 174.632
R11502 VDD.t1111 VDD.n3930 174.632
R11503 VDD.t27 VDD.n4188 174.632
R11504 VDD.t1433 VDD.n4446 174.632
R11505 VDD.t372 VDD.n4704 174.632
R11506 VDD.t420 VDD.n4962 174.632
R11507 VDD.t2 VDD.n5220 174.632
R11508 VDD.t621 VDD 174.602
R11509 VDD.t578 VDD 174.602
R11510 VDD.n693 VDD.n692 174.595
R11511 VDD.n556 VDD.n555 174.595
R11512 VDD.n562 VDD.n561 174.595
R11513 VDD.n568 VDD.n567 174.595
R11514 VDD.n574 VDD.n573 174.595
R11515 VDD.n579 VDD.n578 174.595
R11516 VDD.n535 VDD.n534 174.595
R11517 VDD.n530 VDD.n529 174.595
R11518 VDD.n614 VDD.n613 174.595
R11519 VDD.n608 VDD.n607 174.595
R11520 VDD.n602 VDD.n601 174.595
R11521 VDD.n596 VDD.n595 174.595
R11522 VDD.n592 VDD.n591 174.595
R11523 VDD.n526 VDD.n525 174.595
R11524 VDD.n546 VDD.n545 174.595
R11525 VDD.n639 VDD.n638 174.595
R11526 VDD.n645 VDD.n644 174.595
R11527 VDD.n651 VDD.n650 174.595
R11528 VDD.n657 VDD.n656 174.595
R11529 VDD.n662 VDD.n661 174.595
R11530 VDD.n632 VDD.n631 174.595
R11531 VDD.n626 VDD.n625 174.595
R11532 VDD.n749 VDD.n748 174.595
R11533 VDD.n755 VDD.n754 174.595
R11534 VDD.n761 VDD.n760 174.595
R11535 VDD.n767 VDD.n766 174.595
R11536 VDD.n771 VDD.n770 174.595
R11537 VDD.n778 VDD.n777 174.595
R11538 VDD.n786 VDD.n785 174.595
R11539 VDD.n702 VDD.n701 174.595
R11540 VDD.n708 VDD.n707 174.595
R11541 VDD.n714 VDD.n713 174.595
R11542 VDD.n720 VDD.n719 174.595
R11543 VDD.n724 VDD.n723 174.595
R11544 VDD.n730 VDD.n729 174.595
R11545 VDD.n738 VDD.n737 174.595
R11546 VDD.n1043 VDD.n1042 174.595
R11547 VDD.n906 VDD.n905 174.595
R11548 VDD.n912 VDD.n911 174.595
R11549 VDD.n918 VDD.n917 174.595
R11550 VDD.n924 VDD.n923 174.595
R11551 VDD.n929 VDD.n928 174.595
R11552 VDD.n885 VDD.n884 174.595
R11553 VDD.n880 VDD.n879 174.595
R11554 VDD.n964 VDD.n963 174.595
R11555 VDD.n958 VDD.n957 174.595
R11556 VDD.n952 VDD.n951 174.595
R11557 VDD.n946 VDD.n945 174.595
R11558 VDD.n942 VDD.n941 174.595
R11559 VDD.n876 VDD.n875 174.595
R11560 VDD.n896 VDD.n895 174.595
R11561 VDD.n989 VDD.n988 174.595
R11562 VDD.n995 VDD.n994 174.595
R11563 VDD.n1001 VDD.n1000 174.595
R11564 VDD.n1007 VDD.n1006 174.595
R11565 VDD.n1012 VDD.n1011 174.595
R11566 VDD.n982 VDD.n981 174.595
R11567 VDD.n976 VDD.n975 174.595
R11568 VDD.n1099 VDD.n1098 174.595
R11569 VDD.n1105 VDD.n1104 174.595
R11570 VDD.n1111 VDD.n1110 174.595
R11571 VDD.n1117 VDD.n1116 174.595
R11572 VDD.n1121 VDD.n1120 174.595
R11573 VDD.n1128 VDD.n1127 174.595
R11574 VDD.n1136 VDD.n1135 174.595
R11575 VDD.n1052 VDD.n1051 174.595
R11576 VDD.n1058 VDD.n1057 174.595
R11577 VDD.n1064 VDD.n1063 174.595
R11578 VDD.n1070 VDD.n1069 174.595
R11579 VDD.n1074 VDD.n1073 174.595
R11580 VDD.n1080 VDD.n1079 174.595
R11581 VDD.n1088 VDD.n1087 174.595
R11582 VDD.n288 VDD.n287 174.595
R11583 VDD.n155 VDD.n154 174.595
R11584 VDD.n161 VDD.n160 174.595
R11585 VDD.n167 VDD.n166 174.595
R11586 VDD.n173 VDD.n172 174.595
R11587 VDD.n178 VDD.n177 174.595
R11588 VDD.n134 VDD.n133 174.595
R11589 VDD.n129 VDD.n128 174.595
R11590 VDD.n213 VDD.n212 174.595
R11591 VDD.n207 VDD.n206 174.595
R11592 VDD.n201 VDD.n200 174.595
R11593 VDD.n195 VDD.n194 174.595
R11594 VDD.n191 VDD.n190 174.595
R11595 VDD.n125 VDD.n124 174.595
R11596 VDD.n145 VDD.n144 174.595
R11597 VDD.n112 VDD.n111 174.595
R11598 VDD.n240 VDD.n239 174.595
R11599 VDD.n246 VDD.n245 174.595
R11600 VDD.n252 VDD.n251 174.595
R11601 VDD.n257 VDD.n256 174.595
R11602 VDD.n231 VDD.n230 174.595
R11603 VDD.n225 VDD.n224 174.595
R11604 VDD.n344 VDD.n343 174.595
R11605 VDD.n350 VDD.n349 174.595
R11606 VDD.n356 VDD.n355 174.595
R11607 VDD.n362 VDD.n361 174.595
R11608 VDD.n366 VDD.n365 174.595
R11609 VDD.n373 VDD.n372 174.595
R11610 VDD.n381 VDD.n380 174.595
R11611 VDD.n297 VDD.n296 174.595
R11612 VDD.n303 VDD.n302 174.595
R11613 VDD.n309 VDD.n308 174.595
R11614 VDD.n315 VDD.n314 174.595
R11615 VDD.n319 VDD.n318 174.595
R11616 VDD.n325 VDD.n324 174.595
R11617 VDD.n333 VDD.n332 174.595
R11618 VDD.n1353 VDD.n1352 174.595
R11619 VDD.n1335 VDD.n1334 174.595
R11620 VDD.n1329 VDD.n1328 174.595
R11621 VDD.n1322 VDD.n1321 174.595
R11622 VDD.n1435 VDD.n1434 174.595
R11623 VDD.n1439 VDD.n1438 174.595
R11624 VDD.n1445 VDD.n1444 174.595
R11625 VDD.n1451 VDD.n1450 174.595
R11626 VDD.n1379 VDD.n1378 174.595
R11627 VDD.n1385 VDD.n1384 174.595
R11628 VDD.n1391 VDD.n1390 174.595
R11629 VDD.n1403 VDD.n1402 174.595
R11630 VDD.n1408 VDD.n1407 174.595
R11631 VDD.n1414 VDD.n1413 174.595
R11632 VDD.n1420 VDD.n1419 174.595
R11633 VDD.n1306 VDD.n1305 174.595
R11634 VDD.n1299 VDD.n1298 174.595
R11635 VDD.n1293 VDD.n1292 174.595
R11636 VDD.n1268 VDD.n1267 174.595
R11637 VDD.n1272 VDD.n1271 174.595
R11638 VDD.n1278 VDD.n1277 174.595
R11639 VDD.n1265 VDD.n1264 174.595
R11640 VDD.n1465 VDD.n1464 174.595
R11641 VDD.n1471 VDD.n1470 174.595
R11642 VDD.n1477 VDD.n1476 174.595
R11643 VDD.n1483 VDD.n1482 174.595
R11644 VDD.n1487 VDD.n1486 174.595
R11645 VDD.n1493 VDD.n1492 174.595
R11646 VDD.n1499 VDD.n1498 174.595
R11647 VDD.n1515 VDD.n1514 174.595
R11648 VDD.n1521 VDD.n1520 174.595
R11649 VDD.n1257 VDD.n1256 174.595
R11650 VDD.n1531 VDD.n1530 174.595
R11651 VDD.n1535 VDD.n1534 174.595
R11652 VDD.n1253 VDD.n1252 174.595
R11653 VDD.n1248 VDD.n1247 174.595
R11654 VDD VDD.t1128 174.385
R11655 VDD VDD.t1146 174.385
R11656 VDD VDD.t1276 173.083
R11657 VDD.n670 VDD.t780 173.036
R11658 VDD.n1020 VDD.t1484 173.036
R11659 VDD.n1822 VDD.n1820 170.542
R11660 VDD.n2143 VDD.n2141 170.542
R11661 VDD.n2401 VDD.n2399 170.542
R11662 VDD.n2659 VDD.n2657 170.542
R11663 VDD.n2917 VDD.n2915 170.542
R11664 VDD.n3175 VDD.n3173 170.542
R11665 VDD.n3433 VDD.n3431 170.542
R11666 VDD.n5753 VDD.n5751 170.542
R11667 VDD.n5499 VDD.n5497 170.542
R11668 VDD.n3691 VDD.n3689 170.542
R11669 VDD.n3949 VDD.n3947 170.542
R11670 VDD.n4207 VDD.n4205 170.542
R11671 VDD.n4465 VDD.n4463 170.542
R11672 VDD.n4723 VDD.n4721 170.542
R11673 VDD.n4981 VDD.n4979 170.542
R11674 VDD.n5239 VDD.n5237 170.542
R11675 VDD.t588 VDD 170.478
R11676 VDD.t403 VDD 170.478
R11677 VDD VDD.n1428 169.179
R11678 VDD.n32 VDD.n31 169.107
R11679 VDD.n509 VDD.n508 169.107
R11680 VDD.n436 VDD.n435 169.107
R11681 VDD.n405 VDD.n404 169.107
R11682 VDD.n107 VDD.n106 169.107
R11683 VDD.n1176 VDD.n1175 169.107
R11684 VDD.n1594 VDD.n1593 169.107
R11685 VDD.n1563 VDD.n1562 169.107
R11686 VDD.n819 VDD.n800 169.107
R11687 VDD.n812 VDD.n803 169.107
R11688 VDD.n1202 VDD.n1183 169.107
R11689 VDD.n1195 VDD.n1186 169.107
R11690 VDD.n673 VDD.n672 169.017
R11691 VDD.n1023 VDD.n1022 169.017
R11692 VDD.n268 VDD.n267 169.017
R11693 VDD.n1645 VDD.t784 168.561
R11694 VDD.n1689 VDD.n1673 167.234
R11695 VDD.n2038 VDD.n2022 167.234
R11696 VDD.n2268 VDD.n2252 167.234
R11697 VDD.n2526 VDD.n2510 167.234
R11698 VDD.n2784 VDD.n2768 167.234
R11699 VDD.n3042 VDD.n3026 167.234
R11700 VDD.n3300 VDD.n3284 167.234
R11701 VDD.n5623 VDD.n5607 167.234
R11702 VDD.n5369 VDD.n5353 167.234
R11703 VDD.n3558 VDD.n3542 167.234
R11704 VDD.n3816 VDD.n3800 167.234
R11705 VDD.n4074 VDD.n4058 167.234
R11706 VDD.n4332 VDD.n4316 167.234
R11707 VDD.n4590 VDD.n4574 167.234
R11708 VDD.n4848 VDD.n4832 167.234
R11709 VDD.n5106 VDD.n5090 167.234
R11710 VDD.n1746 VDD.n1715 166.812
R11711 VDD.n2095 VDD.n2064 166.812
R11712 VDD.n2325 VDD.n2294 166.812
R11713 VDD.n2583 VDD.n2552 166.812
R11714 VDD.n2841 VDD.n2810 166.812
R11715 VDD.n3099 VDD.n3068 166.812
R11716 VDD.n3357 VDD.n3326 166.812
R11717 VDD.n5680 VDD.n5649 166.812
R11718 VDD.n5426 VDD.n5395 166.812
R11719 VDD.n3615 VDD.n3584 166.812
R11720 VDD.n3873 VDD.n3842 166.812
R11721 VDD.n4131 VDD.n4100 166.812
R11722 VDD.n4389 VDD.n4358 166.812
R11723 VDD.n4647 VDD.n4616 166.812
R11724 VDD.n4905 VDD.n4874 166.812
R11725 VDD.n5163 VDD.n5132 166.812
R11726 VDD.n1645 VDD.t1511 166.328
R11727 VDD.n1834 VDD.n1830 165.767
R11728 VDD.n1814 VDD.n1813 165.767
R11729 VDD.n2135 VDD.n2134 165.767
R11730 VDD.n2155 VDD.n2151 165.767
R11731 VDD.n2393 VDD.n2392 165.767
R11732 VDD.n2413 VDD.n2409 165.767
R11733 VDD.n2651 VDD.n2650 165.767
R11734 VDD.n2671 VDD.n2667 165.767
R11735 VDD.n2909 VDD.n2908 165.767
R11736 VDD.n2929 VDD.n2925 165.767
R11737 VDD.n3167 VDD.n3166 165.767
R11738 VDD.n3187 VDD.n3183 165.767
R11739 VDD.n3425 VDD.n3424 165.767
R11740 VDD.n3445 VDD.n3441 165.767
R11741 VDD.n5745 VDD.n5744 165.767
R11742 VDD.n5765 VDD.n5761 165.767
R11743 VDD.n5491 VDD.n5490 165.767
R11744 VDD.n5511 VDD.n5507 165.767
R11745 VDD.n3683 VDD.n3682 165.767
R11746 VDD.n3703 VDD.n3699 165.767
R11747 VDD.n3941 VDD.n3940 165.767
R11748 VDD.n3961 VDD.n3957 165.767
R11749 VDD.n4199 VDD.n4198 165.767
R11750 VDD.n4219 VDD.n4215 165.767
R11751 VDD.n4457 VDD.n4456 165.767
R11752 VDD.n4477 VDD.n4473 165.767
R11753 VDD.n4715 VDD.n4714 165.767
R11754 VDD.n4735 VDD.n4731 165.767
R11755 VDD.n4973 VDD.n4972 165.767
R11756 VDD.n4993 VDD.n4989 165.767
R11757 VDD.n5231 VDD.n5230 165.767
R11758 VDD.n5251 VDD.n5247 165.767
R11759 VDD.t1046 VDD.t603 164.554
R11760 VDD.t1431 VDD.t1351 164.554
R11761 VDD.t596 VDD.t1356 164.554
R11762 VDD.n24 VDD.n1 164.215
R11763 VDD.n488 VDD.n468 164.215
R11764 VDD.n440 VDD.n439 164.215
R11765 VDD.n460 VDD.n459 164.215
R11766 VDD.n86 VDD.n66 164.215
R11767 VDD.n37 VDD.n36 164.215
R11768 VDD.n57 VDD.n56 164.215
R11769 VDD.n1168 VDD.n1145 164.215
R11770 VDD.n1699 VDD.n1682 161.506
R11771 VDD.n2048 VDD.n2031 161.506
R11772 VDD.n2278 VDD.n2261 161.506
R11773 VDD.n2536 VDD.n2519 161.506
R11774 VDD.n2794 VDD.n2777 161.506
R11775 VDD.n3052 VDD.n3035 161.506
R11776 VDD.n3310 VDD.n3293 161.506
R11777 VDD.n5633 VDD.n5616 161.506
R11778 VDD.n5379 VDD.n5362 161.506
R11779 VDD.n3568 VDD.n3551 161.506
R11780 VDD.n3826 VDD.n3809 161.506
R11781 VDD.n4084 VDD.n4067 161.506
R11782 VDD.n4342 VDD.n4325 161.506
R11783 VDD.n4600 VDD.n4583 161.506
R11784 VDD.n4858 VDD.n4841 161.506
R11785 VDD.n5116 VDD.n5099 161.506
R11786 VDD.n1741 VDD.n1728 159.143
R11787 VDD.n2090 VDD.n2077 159.143
R11788 VDD.n2320 VDD.n2307 159.143
R11789 VDD.n2578 VDD.n2565 159.143
R11790 VDD.n2836 VDD.n2823 159.143
R11791 VDD.n3094 VDD.n3081 159.143
R11792 VDD.n3352 VDD.n3339 159.143
R11793 VDD.n5675 VDD.n5662 159.143
R11794 VDD.n5421 VDD.n5408 159.143
R11795 VDD.n3610 VDD.n3597 159.143
R11796 VDD.n3868 VDD.n3855 159.143
R11797 VDD.n4126 VDD.n4113 159.143
R11798 VDD.n4384 VDD.n4371 159.143
R11799 VDD.n4642 VDD.n4629 159.143
R11800 VDD.n4900 VDD.n4887 159.143
R11801 VDD.n5158 VDD.n5145 159.143
R11802 VDD.n1905 VDD.n1892 159.108
R11803 VDD.n1858 VDD.n1857 159.108
R11804 VDD.n2179 VDD.n2178 159.108
R11805 VDD.n2226 VDD.n2213 159.108
R11806 VDD.n2437 VDD.n2436 159.108
R11807 VDD.n2484 VDD.n2471 159.108
R11808 VDD.n2695 VDD.n2694 159.108
R11809 VDD.n2742 VDD.n2729 159.108
R11810 VDD.n2953 VDD.n2952 159.108
R11811 VDD.n3000 VDD.n2987 159.108
R11812 VDD.n3211 VDD.n3210 159.108
R11813 VDD.n3258 VDD.n3245 159.108
R11814 VDD.n3469 VDD.n3468 159.108
R11815 VDD.n3516 VDD.n3503 159.108
R11816 VDD.n5789 VDD.n5788 159.108
R11817 VDD.n5836 VDD.n5823 159.108
R11818 VDD.n5535 VDD.n5534 159.108
R11819 VDD.n5582 VDD.n5569 159.108
R11820 VDD.n3727 VDD.n3726 159.108
R11821 VDD.n3774 VDD.n3761 159.108
R11822 VDD.n3985 VDD.n3984 159.108
R11823 VDD.n4032 VDD.n4019 159.108
R11824 VDD.n4243 VDD.n4242 159.108
R11825 VDD.n4290 VDD.n4277 159.108
R11826 VDD.n4501 VDD.n4500 159.108
R11827 VDD.n4548 VDD.n4535 159.108
R11828 VDD.n4759 VDD.n4758 159.108
R11829 VDD.n4806 VDD.n4793 159.108
R11830 VDD.n5017 VDD.n5016 159.108
R11831 VDD.n5064 VDD.n5051 159.108
R11832 VDD.n5275 VDD.n5274 159.108
R11833 VDD.n5322 VDD.n5309 159.108
R11834 VDD.n1605 VDD.t1505 158.886
R11835 VDD.n1700 VDD.n1699 158.776
R11836 VDD.n2049 VDD.n2048 158.776
R11837 VDD.n2279 VDD.n2278 158.776
R11838 VDD.n2537 VDD.n2536 158.776
R11839 VDD.n2795 VDD.n2794 158.776
R11840 VDD.n3053 VDD.n3052 158.776
R11841 VDD.n3311 VDD.n3310 158.776
R11842 VDD.n5634 VDD.n5633 158.776
R11843 VDD.n5380 VDD.n5379 158.776
R11844 VDD.n3569 VDD.n3568 158.776
R11845 VDD.n3827 VDD.n3826 158.776
R11846 VDD.n4085 VDD.n4084 158.776
R11847 VDD.n4343 VDD.n4342 158.776
R11848 VDD.n4601 VDD.n4600 158.776
R11849 VDD.n4859 VDD.n4858 158.776
R11850 VDD.n5117 VDD.n5116 158.776
R11851 VDD.n541 VDD.t184 158.117
R11852 VDD.n620 VDD.t168 158.117
R11853 VDD.n516 VDD.t148 158.117
R11854 VDD.n519 VDD.t110 158.117
R11855 VDD.n522 VDD.t1388 158.117
R11856 VDD.n891 VDD.t957 158.117
R11857 VDD.n970 VDD.t943 158.117
R11858 VDD.n866 VDD.t921 158.117
R11859 VDD.n869 VDD.t883 158.117
R11860 VDD.n872 VDD.t44 158.117
R11861 VDD.n140 VDD.t737 158.117
R11862 VDD.n219 VDD.t721 158.117
R11863 VDD.n115 VDD.t701 158.117
R11864 VDD.n118 VDD.t663 158.117
R11865 VDD.n121 VDD.t218 158.117
R11866 VDD.n1341 VDD.t1245 158.117
R11867 VDD.n1347 VDD.t297 158.117
R11868 VDD.n1312 VDD.t1221 158.117
R11869 VDD.n1262 VDD.t1223 158.117
R11870 VDD.n1259 VDD.t1171 158.117
R11871 VDD.n671 VDD.t781 158.06
R11872 VDD.n1021 VDD.t1485 158.06
R11873 VDD.n266 VDD.t380 158.06
R11874 VDD.n1362 VDD.t1483 158.06
R11875 VDD.n826 VDD.t331 158.06
R11876 VDD.n825 VDD.t1344 158.06
R11877 VDD.n824 VDD.t1315 158.06
R11878 VDD.n823 VDD.t1320 158.06
R11879 VDD.n822 VDD.t355 158.06
R11880 VDD.n1542 VDD.t537 158.06
R11881 VDD.n1209 VDD.t970 158.06
R11882 VDD.n1208 VDD.t1375 158.06
R11883 VDD.n1207 VDD.t1361 158.06
R11884 VDD.n1206 VDD.t1312 158.06
R11885 VDD.n1205 VDD.t799 158.06
R11886 VDD.n1616 VDD.t1508 156.403
R11887 VDD.t335 VDD.t557 155.456
R11888 VDD.t502 VDD.t1376 155.456
R11889 VDD.n1679 VDD.n1670 155.294
R11890 VDD.n2028 VDD.n2019 155.294
R11891 VDD.n2258 VDD.n2249 155.294
R11892 VDD.n2516 VDD.n2507 155.294
R11893 VDD.n2774 VDD.n2765 155.294
R11894 VDD.n3032 VDD.n3023 155.294
R11895 VDD.n3290 VDD.n3281 155.294
R11896 VDD.n5613 VDD.n5604 155.294
R11897 VDD.n5359 VDD.n5350 155.294
R11898 VDD.n3548 VDD.n3539 155.294
R11899 VDD.n3806 VDD.n3797 155.294
R11900 VDD.n4064 VDD.n4055 155.294
R11901 VDD.n4322 VDD.n4313 155.294
R11902 VDD.n4580 VDD.n4571 155.294
R11903 VDD.n4838 VDD.n4829 155.294
R11904 VDD.n5096 VDD.n5087 155.294
R11905 VDD.n1507 VDD.t1226 153.562
R11906 VDD VDD.t1495 151.137
R11907 VDD VDD.t1489 151.137
R11908 VDD.n1784 VDD.t446 151.123
R11909 VDD.n1786 VDD.t1029 151.123
R11910 VDD.n1992 VDD.t78 151.123
R11911 VDD.n1994 VDD.t1269 151.123
R11912 VDD.n2363 VDD.t1445 151.123
R11913 VDD.n2365 VDD.t833 151.123
R11914 VDD.n2621 VDD.t570 151.123
R11915 VDD.n2623 VDD.t1420 151.123
R11916 VDD.n2879 VDD.t977 151.123
R11917 VDD.n2881 VDD.t434 151.123
R11918 VDD.n3137 VDD.t544 151.123
R11919 VDD.n3139 VDD.t389 151.123
R11920 VDD.n3395 VDD.t581 151.123
R11921 VDD.n3397 VDD.t1298 151.123
R11922 VDD.n5718 VDD.t1467 151.123
R11923 VDD.n5720 VDD.t474 151.123
R11924 VDD.n5464 VDD.t1000 151.123
R11925 VDD.n5466 VDD.t1260 151.123
R11926 VDD.n3653 VDD.t1335 151.123
R11927 VDD.n3655 VDD.t1369 151.123
R11928 VDD.n3911 VDD.t489 151.123
R11929 VDD.n3913 VDD.t1116 151.123
R11930 VDD.n4169 VDD.t10 151.123
R11931 VDD.n4171 VDD.t32 151.123
R11932 VDD.n4427 VDD.t1051 151.123
R11933 VDD.n4429 VDD.t1434 151.123
R11934 VDD.n4685 VDD.t20 151.123
R11935 VDD.n4687 VDD.t376 151.123
R11936 VDD.n4943 VDD.t822 151.123
R11937 VDD.n4945 VDD.t1041 151.123
R11938 VDD.n5201 VDD.t1328 151.123
R11939 VDD.n5203 VDD.t1254 151.123
R11940 VDD.n524 VDD.t338 151.123
R11941 VDD.n874 VDD.t1079 151.123
R11942 VDD.n123 VDD.t993 151.123
R11943 VDD.n1357 VDD.t1279 151.123
R11944 VDD.n1624 VDD.t1506 150.03
R11945 VDD.n1627 VDD.t1502 150.03
R11946 VDD.n1629 VDD.t1504 150.03
R11947 VDD.n1632 VDD.t1510 150.03
R11948 VDD.t356 VDD.t551 148.481
R11949 VDD.t807 VDD.t606 148.481
R11950 VDD.n1802 VDD.t443 146.691
R11951 VDD.n2010 VDD.t77 146.691
R11952 VDD.n2381 VDD.t1444 146.691
R11953 VDD.n2639 VDD.t569 146.691
R11954 VDD.n2897 VDD.t976 146.691
R11955 VDD.n3155 VDD.t543 146.691
R11956 VDD.n3413 VDD.t580 146.691
R11957 VDD.n5736 VDD.t1466 146.691
R11958 VDD.n5482 VDD.t997 146.691
R11959 VDD.n3671 VDD.t1333 146.691
R11960 VDD.n3929 VDD.t483 146.691
R11961 VDD.n4187 VDD.t7 146.691
R11962 VDD.n4445 VDD.t1050 146.691
R11963 VDD.n4703 VDD.t19 146.691
R11964 VDD.n4961 VDD.t560 146.691
R11965 VDD.n5219 VDD.t1006 146.691
R11966 VDD.t1454 VDD.t1464 145.243
R11967 VDD.t498 VDD.t451 145.243
R11968 VDD.n1647 VDD.t1512 145.043
R11969 VDD.n1741 VDD.n1740 143.435
R11970 VDD.n2090 VDD.n2089 143.435
R11971 VDD.n2320 VDD.n2319 143.435
R11972 VDD.n2578 VDD.n2577 143.435
R11973 VDD.n2836 VDD.n2835 143.435
R11974 VDD.n3094 VDD.n3093 143.435
R11975 VDD.n3352 VDD.n3351 143.435
R11976 VDD.n5675 VDD.n5674 143.435
R11977 VDD.n5421 VDD.n5420 143.435
R11978 VDD.n3610 VDD.n3609 143.435
R11979 VDD.n3868 VDD.n3867 143.435
R11980 VDD.n4126 VDD.n4125 143.435
R11981 VDD.n4384 VDD.n4383 143.435
R11982 VDD.n4642 VDD.n4641 143.435
R11983 VDD.n4900 VDD.n4899 143.435
R11984 VDD.n5158 VDD.n5157 143.435
R11985 VDD.t611 VDD.t1341 143.232
R11986 VDD.t1491 VDD.t823 143.232
R11987 VDD.t127 VDD.t101 142.5
R11988 VDD.t213 VDD.t127 142.5
R11989 VDD.t105 VDD.t213 142.5
R11990 VDD.t97 VDD.t105 142.5
R11991 VDD.t119 VDD.t97 142.5
R11992 VDD.t87 VDD.t145 142.5
R11993 VDD.t123 VDD.t87 142.5
R11994 VDD.t193 VDD.t123 142.5
R11995 VDD.t89 VDD.t193 142.5
R11996 VDD.t113 VDD.t89 142.5
R11997 VDD.t177 VDD.t113 142.5
R11998 VDD.t207 VDD.t177 142.5
R11999 VDD.t139 VDD.t207 142.5
R12000 VDD.t183 VDD.t139 142.5
R12001 VDD.t171 VDD.t103 142.5
R12002 VDD.t197 VDD.t171 142.5
R12003 VDD.t95 VDD.t197 142.5
R12004 VDD.t151 VDD.t95 142.5
R12005 VDD.t185 VDD.t117 142.5
R12006 VDD.t117 VDD.t155 142.5
R12007 VDD.t155 VDD.t189 142.5
R12008 VDD.t189 VDD.t125 142.5
R12009 VDD.t125 VDD.t205 142.5
R12010 VDD.t205 VDD.t137 142.5
R12011 VDD.t137 VDD.t163 142.5
R12012 VDD.t163 VDD.t211 142.5
R12013 VDD.t211 VDD.t143 142.5
R12014 VDD.t143 VDD.t167 142.5
R12015 VDD.t91 VDD.t149 142.5
R12016 VDD.t149 VDD.t179 142.5
R12017 VDD.t179 VDD.t115 142.5
R12018 VDD.t115 VDD.t201 142.5
R12019 VDD.t201 VDD.t111 142.5
R12020 VDD.t203 VDD.t175 142.5
R12021 VDD.t133 VDD.t203 142.5
R12022 VDD.t159 VDD.t133 142.5
R12023 VDD.t191 VDD.t159 142.5
R12024 VDD.t135 VDD.t191 142.5
R12025 VDD.t161 VDD.t135 142.5
R12026 VDD.t107 VDD.t161 142.5
R12027 VDD.t129 VDD.t107 142.5
R12028 VDD.t147 VDD.t129 142.5
R12029 VDD.t195 VDD.t169 142.5
R12030 VDD.t93 VDD.t195 142.5
R12031 VDD.t173 VDD.t93 142.5
R12032 VDD.t131 VDD.t199 142.5
R12033 VDD.t153 VDD.t131 142.5
R12034 VDD.t187 VDD.t153 142.5
R12035 VDD.t121 VDD.t187 142.5
R12036 VDD.t157 VDD.t121 142.5
R12037 VDD.t99 VDD.t157 142.5
R12038 VDD.t181 VDD.t99 142.5
R12039 VDD.t209 VDD.t181 142.5
R12040 VDD.t141 VDD.t209 142.5
R12041 VDD.t165 VDD.t141 142.5
R12042 VDD.t109 VDD.t165 142.5
R12043 VDD.t1411 VDD.t1397 142.5
R12044 VDD.t1399 VDD.t1391 142.5
R12045 VDD.t1409 VDD.t1399 142.5
R12046 VDD.t1405 VDD.t1409 142.5
R12047 VDD.t1413 VDD.t1405 142.5
R12048 VDD.t1393 VDD.t1413 142.5
R12049 VDD.t1407 VDD.t1393 142.5
R12050 VDD.t1415 VDD.t1407 142.5
R12051 VDD.t1395 VDD.t1415 142.5
R12052 VDD.t1401 VDD.t1395 142.5
R12053 VDD.t1385 VDD.t1401 142.5
R12054 VDD.t1389 VDD.t1385 142.5
R12055 VDD.t1403 VDD.t1389 142.5
R12056 VDD.t1387 VDD.t1403 142.5
R12057 VDD.t341 VDD.t339 142.5
R12058 VDD.t343 VDD.t341 142.5
R12059 VDD.t337 VDD.t343 142.5
R12060 VDD.t900 VDD.t874 142.5
R12061 VDD.t858 VDD.t900 142.5
R12062 VDD.t878 VDD.t858 142.5
R12063 VDD.t870 VDD.t878 142.5
R12064 VDD.t890 VDD.t870 142.5
R12065 VDD.t860 VDD.t918 142.5
R12066 VDD.t896 VDD.t860 142.5
R12067 VDD.t838 VDD.t896 142.5
R12068 VDD.t862 VDD.t838 142.5
R12069 VDD.t886 VDD.t862 142.5
R12070 VDD.t950 VDD.t886 142.5
R12071 VDD.t852 VDD.t950 142.5
R12072 VDD.t912 VDD.t852 142.5
R12073 VDD.t956 VDD.t912 142.5
R12074 VDD.t932 VDD.t876 142.5
R12075 VDD.t842 VDD.t932 142.5
R12076 VDD.t868 VDD.t842 142.5
R12077 VDD.t924 VDD.t868 142.5
R12078 VDD.t958 VDD.t892 142.5
R12079 VDD.t892 VDD.t928 142.5
R12080 VDD.t928 VDD.t962 142.5
R12081 VDD.t962 VDD.t898 142.5
R12082 VDD.t898 VDD.t850 142.5
R12083 VDD.t850 VDD.t910 142.5
R12084 VDD.t910 VDD.t938 142.5
R12085 VDD.t938 VDD.t856 142.5
R12086 VDD.t856 VDD.t916 142.5
R12087 VDD.t916 VDD.t942 142.5
R12088 VDD.t864 VDD.t922 142.5
R12089 VDD.t922 VDD.t952 142.5
R12090 VDD.t952 VDD.t888 142.5
R12091 VDD.t888 VDD.t846 142.5
R12092 VDD.t846 VDD.t884 142.5
R12093 VDD.t848 VDD.t948 142.5
R12094 VDD.t902 VDD.t848 142.5
R12095 VDD.t934 VDD.t902 142.5
R12096 VDD.t964 VDD.t934 142.5
R12097 VDD.t908 VDD.t964 142.5
R12098 VDD.t936 VDD.t908 142.5
R12099 VDD.t880 VDD.t936 142.5
R12100 VDD.t904 VDD.t880 142.5
R12101 VDD.t920 VDD.t904 142.5
R12102 VDD.t840 VDD.t944 142.5
R12103 VDD.t866 VDD.t840 142.5
R12104 VDD.t946 VDD.t866 142.5
R12105 VDD.t906 VDD.t844 142.5
R12106 VDD.t926 VDD.t906 142.5
R12107 VDD.t960 VDD.t926 142.5
R12108 VDD.t894 VDD.t960 142.5
R12109 VDD.t930 VDD.t894 142.5
R12110 VDD.t872 VDD.t930 142.5
R12111 VDD.t954 VDD.t872 142.5
R12112 VDD.t854 VDD.t954 142.5
R12113 VDD.t914 VDD.t854 142.5
R12114 VDD.t940 VDD.t914 142.5
R12115 VDD.t882 VDD.t940 142.5
R12116 VDD.t35 VDD.t53 142.5
R12117 VDD.t55 VDD.t47 142.5
R12118 VDD.t65 VDD.t55 142.5
R12119 VDD.t61 VDD.t65 142.5
R12120 VDD.t37 VDD.t61 142.5
R12121 VDD.t49 VDD.t37 142.5
R12122 VDD.t63 VDD.t49 142.5
R12123 VDD.t39 VDD.t63 142.5
R12124 VDD.t51 VDD.t39 142.5
R12125 VDD.t57 VDD.t51 142.5
R12126 VDD.t41 VDD.t57 142.5
R12127 VDD.t45 VDD.t41 142.5
R12128 VDD.t59 VDD.t45 142.5
R12129 VDD.t43 VDD.t59 142.5
R12130 VDD.t1082 VDD.t1080 142.5
R12131 VDD.t1076 VDD.t1082 142.5
R12132 VDD.t1078 VDD.t1076 142.5
R12133 VDD.t680 VDD.t654 142.5
R12134 VDD.t766 VDD.t680 142.5
R12135 VDD.t658 VDD.t766 142.5
R12136 VDD.t778 VDD.t658 142.5
R12137 VDD.t670 VDD.t778 142.5
R12138 VDD.t768 VDD.t698 142.5
R12139 VDD.t678 VDD.t768 142.5
R12140 VDD.t746 VDD.t678 142.5
R12141 VDD.t770 VDD.t746 142.5
R12142 VDD.t666 VDD.t770 142.5
R12143 VDD.t730 VDD.t666 142.5
R12144 VDD.t760 VDD.t730 142.5
R12145 VDD.t692 VDD.t760 142.5
R12146 VDD.t736 VDD.t692 142.5
R12147 VDD.t724 VDD.t656 142.5
R12148 VDD.t750 VDD.t724 142.5
R12149 VDD.t776 VDD.t750 142.5
R12150 VDD.t704 VDD.t776 142.5
R12151 VDD.t738 VDD.t672 142.5
R12152 VDD.t672 VDD.t708 142.5
R12153 VDD.t708 VDD.t742 142.5
R12154 VDD.t742 VDD.t676 142.5
R12155 VDD.t676 VDD.t758 142.5
R12156 VDD.t758 VDD.t690 142.5
R12157 VDD.t690 VDD.t716 142.5
R12158 VDD.t716 VDD.t764 142.5
R12159 VDD.t764 VDD.t696 142.5
R12160 VDD.t696 VDD.t720 142.5
R12161 VDD.t772 VDD.t702 142.5
R12162 VDD.t702 VDD.t732 142.5
R12163 VDD.t732 VDD.t668 142.5
R12164 VDD.t668 VDD.t754 142.5
R12165 VDD.t754 VDD.t664 142.5
R12166 VDD.t756 VDD.t728 142.5
R12167 VDD.t686 VDD.t756 142.5
R12168 VDD.t712 VDD.t686 142.5
R12169 VDD.t744 VDD.t712 142.5
R12170 VDD.t688 VDD.t744 142.5
R12171 VDD.t714 VDD.t688 142.5
R12172 VDD.t660 VDD.t714 142.5
R12173 VDD.t682 VDD.t660 142.5
R12174 VDD.t700 VDD.t682 142.5
R12175 VDD.t748 VDD.t722 142.5
R12176 VDD.t774 VDD.t748 142.5
R12177 VDD.t726 VDD.t774 142.5
R12178 VDD.t684 VDD.t752 142.5
R12179 VDD.t706 VDD.t684 142.5
R12180 VDD.t740 VDD.t706 142.5
R12181 VDD.t674 VDD.t740 142.5
R12182 VDD.t710 VDD.t674 142.5
R12183 VDD.t652 VDD.t710 142.5
R12184 VDD.t734 VDD.t652 142.5
R12185 VDD.t762 VDD.t734 142.5
R12186 VDD.t694 VDD.t762 142.5
R12187 VDD.t718 VDD.t694 142.5
R12188 VDD.t662 VDD.t718 142.5
R12189 VDD.t241 VDD.t227 142.5
R12190 VDD.t229 VDD.t221 142.5
R12191 VDD.t239 VDD.t229 142.5
R12192 VDD.t235 VDD.t239 142.5
R12193 VDD.t243 VDD.t235 142.5
R12194 VDD.t223 VDD.t243 142.5
R12195 VDD.t237 VDD.t223 142.5
R12196 VDD.t245 VDD.t237 142.5
R12197 VDD.t225 VDD.t245 142.5
R12198 VDD.t231 VDD.t225 142.5
R12199 VDD.t215 VDD.t231 142.5
R12200 VDD.t219 VDD.t215 142.5
R12201 VDD.t233 VDD.t219 142.5
R12202 VDD.t217 VDD.t233 142.5
R12203 VDD.t988 VDD.t986 142.5
R12204 VDD.t990 VDD.t988 142.5
R12205 VDD.t992 VDD.t990 142.5
R12206 VDD.t1464 VDD.t471 142.279
R12207 VDD.t605 VDD.t836 142.279
R12208 VDD.t451 VDD.t289 142.279
R12209 VDD.t651 VDD.t538 142.279
R12210 VDD.t411 VDD.t468 141.061
R12211 VDD.t429 VDD.t287 141.061
R12212 VDD.n669 VDD.t1411 139.107
R12213 VDD.n1019 VDD.t35 139.107
R12214 VDD.t752 VDD.n263 139.107
R12215 VDD VDD.t613 138.857
R12216 VDD VDD.t534 138.857
R12217 VDD.t468 VDD.t598 138.183
R12218 VDD.t1066 VDD.t559 138.183
R12219 VDD.t287 VDD.t595 138.183
R12220 VDD.t457 VDD.t1443 138.183
R12221 VDD.t1482 VDD 137.946
R12222 VDD.t274 VDD.n1821 136.591
R12223 VDD.t511 VDD.n2142 136.591
R12224 VDD.t528 VDD.n2400 136.591
R12225 VDD.t1381 VDD.n2658 136.591
R12226 VDD.t414 VDD.n2916 136.591
R12227 VDD.t591 VDD.n3174 136.591
R12228 VDD.t1086 VDD.n3432 136.591
R12229 VDD.t276 VDD.n5752 136.591
R12230 VDD.t512 VDD.n5498 136.591
R12231 VDD.t1085 VDD.n3690 136.591
R12232 VDD.t526 VDD.n3948 136.591
R12233 VDD.t525 VDD.n4206 136.591
R12234 VDD.t264 VDD.n4464 136.591
R12235 VDD.t590 VDD.n4722 136.591
R12236 VDD.t1024 VDD.n4980 136.591
R12237 VDD.t275 VDD.n5238 136.591
R12238 VDD.n1697 VDD.n1696 135.117
R12239 VDD.n2046 VDD.n2045 135.117
R12240 VDD.n2276 VDD.n2275 135.117
R12241 VDD.n2534 VDD.n2533 135.117
R12242 VDD.n2792 VDD.n2791 135.117
R12243 VDD.n3050 VDD.n3049 135.117
R12244 VDD.n3308 VDD.n3307 135.117
R12245 VDD.n5631 VDD.n5630 135.117
R12246 VDD.n5377 VDD.n5376 135.117
R12247 VDD.n3566 VDD.n3565 135.117
R12248 VDD.n3824 VDD.n3823 135.117
R12249 VDD.n4082 VDD.n4081 135.117
R12250 VDD.n4340 VDD.n4339 135.117
R12251 VDD.n4598 VDD.n4597 135.117
R12252 VDD.n4856 VDD.n4855 135.117
R12253 VDD.n5114 VDD.n5113 135.117
R12254 VDD.t1090 VDD.t621 134.732
R12255 VDD.t1096 VDD.t588 134.732
R12256 VDD.t1282 VDD.t578 134.732
R12257 VDD.t258 VDD.t403 134.732
R12258 VDD.n1371 VDD.t1482 132.74
R12259 VDD VDD.t183 132.321
R12260 VDD.t167 VDD 132.321
R12261 VDD VDD.t147 132.321
R12262 VDD.t199 VDD.n668 132.321
R12263 VDD VDD.t109 132.321
R12264 VDD VDD.t1387 132.321
R12265 VDD VDD.t956 132.321
R12266 VDD.t942 VDD 132.321
R12267 VDD VDD.t920 132.321
R12268 VDD.t844 VDD.n1018 132.321
R12269 VDD VDD.t882 132.321
R12270 VDD VDD.t43 132.321
R12271 VDD VDD.t736 132.321
R12272 VDD.t720 VDD 132.321
R12273 VDD VDD.t700 132.321
R12274 VDD VDD.t662 132.321
R12275 VDD.n264 VDD.t241 132.321
R12276 VDD VDD.t217 132.321
R12277 VDD.t1110 VDD.t1090 131.983
R12278 VDD.t1107 VDD.t1096 131.983
R12279 VDD.t782 VDD.t334 131.983
R12280 VDD.t1005 VDD.t1282 131.983
R12281 VDD.t1426 VDD.t258 131.983
R12282 VDD.t428 VDD.t837 131.983
R12283 VDD.n1715 VDD.n1672 131.388
R12284 VDD.n2064 VDD.n2021 131.388
R12285 VDD.n2294 VDD.n2251 131.388
R12286 VDD.n2552 VDD.n2509 131.388
R12287 VDD.n2810 VDD.n2767 131.388
R12288 VDD.n3068 VDD.n3025 131.388
R12289 VDD.n3326 VDD.n3283 131.388
R12290 VDD.n5649 VDD.n5606 131.388
R12291 VDD.n5395 VDD.n5352 131.388
R12292 VDD.n3584 VDD.n3541 131.388
R12293 VDD.n3842 VDD.n3799 131.388
R12294 VDD.n4100 VDD.n4057 131.388
R12295 VDD.n4358 VDD.n4315 131.388
R12296 VDD.n4616 VDD.n4573 131.388
R12297 VDD.n4874 VDD.n4831 131.388
R12298 VDD.n5132 VDD.n5089 131.388
R12299 VDD.n1766 VDD.n1673 131.012
R12300 VDD.n2115 VDD.n2022 131.012
R12301 VDD.n2345 VDD.n2252 131.012
R12302 VDD.n2603 VDD.n2510 131.012
R12303 VDD.n2861 VDD.n2768 131.012
R12304 VDD.n3119 VDD.n3026 131.012
R12305 VDD.n3377 VDD.n3284 131.012
R12306 VDD.n5700 VDD.n5607 131.012
R12307 VDD.n5446 VDD.n5353 131.012
R12308 VDD.n3635 VDD.n3542 131.012
R12309 VDD.n3893 VDD.n3800 131.012
R12310 VDD.n4151 VDD.n4058 131.012
R12311 VDD.n4409 VDD.n4316 131.012
R12312 VDD.n4667 VDD.n4574 131.012
R12313 VDD.n4925 VDD.n4832 131.012
R12314 VDD.n5183 VDD.n5090 131.012
R12315 VDD.n1767 VDD.n1672 130.636
R12316 VDD.n1767 VDD.n1766 130.636
R12317 VDD.n2116 VDD.n2021 130.636
R12318 VDD.n2116 VDD.n2115 130.636
R12319 VDD.n2346 VDD.n2251 130.636
R12320 VDD.n2346 VDD.n2345 130.636
R12321 VDD.n2604 VDD.n2509 130.636
R12322 VDD.n2604 VDD.n2603 130.636
R12323 VDD.n2862 VDD.n2767 130.636
R12324 VDD.n2862 VDD.n2861 130.636
R12325 VDD.n3120 VDD.n3025 130.636
R12326 VDD.n3120 VDD.n3119 130.636
R12327 VDD.n3378 VDD.n3283 130.636
R12328 VDD.n3378 VDD.n3377 130.636
R12329 VDD.n5701 VDD.n5606 130.636
R12330 VDD.n5701 VDD.n5700 130.636
R12331 VDD.n5447 VDD.n5352 130.636
R12332 VDD.n5447 VDD.n5446 130.636
R12333 VDD.n3636 VDD.n3541 130.636
R12334 VDD.n3636 VDD.n3635 130.636
R12335 VDD.n3894 VDD.n3799 130.636
R12336 VDD.n3894 VDD.n3893 130.636
R12337 VDD.n4152 VDD.n4057 130.636
R12338 VDD.n4152 VDD.n4151 130.636
R12339 VDD.n4410 VDD.n4315 130.636
R12340 VDD.n4410 VDD.n4409 130.636
R12341 VDD.n4668 VDD.n4573 130.636
R12342 VDD.n4668 VDD.n4667 130.636
R12343 VDD.n4926 VDD.n4831 130.636
R12344 VDD.n4926 VDD.n4925 130.636
R12345 VDD.n5184 VDD.n5089 130.636
R12346 VDD.n5184 VDD.n5183 130.636
R12347 VDD.n1879 VDD.n1823 129.691
R12348 VDD.n2200 VDD.n2144 129.691
R12349 VDD.n2458 VDD.n2402 129.691
R12350 VDD.n2716 VDD.n2660 129.691
R12351 VDD.n2974 VDD.n2918 129.691
R12352 VDD.n3232 VDD.n3176 129.691
R12353 VDD.n3490 VDD.n3434 129.691
R12354 VDD.n5810 VDD.n5754 129.691
R12355 VDD.n5556 VDD.n5500 129.691
R12356 VDD.n3748 VDD.n3692 129.691
R12357 VDD.n4006 VDD.n3950 129.691
R12358 VDD.n4264 VDD.n4208 129.691
R12359 VDD.n4522 VDD.n4466 129.691
R12360 VDD.n4780 VDD.n4724 129.691
R12361 VDD.n5038 VDD.n4982 129.691
R12362 VDD.n5296 VDD.n5240 129.691
R12363 VDD VDD.t326 129.228
R12364 VDD VDD.t791 129.228
R12365 VDD VDD.t337 127.233
R12366 VDD VDD.t1078 127.233
R12367 VDD VDD.t992 127.233
R12368 VDD.t599 VDD 126.02
R12369 VDD.t1011 VDD 126.02
R12370 VDD.t615 VDD 126.02
R12371 VDD.t247 VDD 126.02
R12372 VDD.t618 VDD 126.02
R12373 VDD.t647 VDD 126.02
R12374 VDD.t532 VDD 126.02
R12375 VDD.t1353 VDD 126.02
R12376 VDD.t391 VDD 126.02
R12377 VDD.t291 VDD 126.02
R12378 VDD.t1348 VDD 126.02
R12379 VDD.t1363 VDD 126.02
R12380 VDD.t608 VDD 126.02
R12381 VDD.t399 VDD 126.02
R12382 VDD.t1099 VDD 126.02
R12383 VDD.t405 VDD 126.02
R12384 VDD.t603 VDD.t1045 122.144
R12385 VDD.t1351 VDD.t819 122.144
R12386 VDD.t1356 VDD.t1290 122.144
R12387 VDD.n1903 VDD.n1898 121.977
R12388 VDD.n2224 VDD.n2219 121.977
R12389 VDD.n2482 VDD.n2477 121.977
R12390 VDD.n2740 VDD.n2735 121.977
R12391 VDD.n2998 VDD.n2993 121.977
R12392 VDD.n3256 VDD.n3251 121.977
R12393 VDD.n3514 VDD.n3509 121.977
R12394 VDD.n5834 VDD.n5829 121.977
R12395 VDD.n5580 VDD.n5575 121.977
R12396 VDD.n3772 VDD.n3767 121.977
R12397 VDD.n4030 VDD.n4025 121.977
R12398 VDD.n4288 VDD.n4283 121.977
R12399 VDD.n4546 VDD.n4541 121.977
R12400 VDD.n4804 VDD.n4799 121.977
R12401 VDD.n5062 VDD.n5057 121.977
R12402 VDD.n5320 VDD.n5315 121.977
R12403 VDD.t1122 VDD.t455 121.529
R12404 VDD.t1457 VDD.t462 121.529
R12405 VDD.n1764 VDD.t1014 121.114
R12406 VDD.t1014 VDD.n1711 121.114
R12407 VDD.n2113 VDD.t623 121.114
R12408 VDD.t623 VDD.n2060 121.114
R12409 VDD.n2343 VDD.t1331 121.114
R12410 VDD.t1331 VDD.n2290 121.114
R12411 VDD.n2601 VDD.t825 121.114
R12412 VDD.t825 VDD.n2548 121.114
R12413 VDD.n2859 VDD.t424 121.114
R12414 VDD.t424 VDD.n2806 121.114
R12415 VDD.n3117 VDD.t395 121.114
R12416 VDD.t395 VDD.n3064 121.114
R12417 VDD.n3375 VDD.t639 121.114
R12418 VDD.t639 VDD.n3322 121.114
R12419 VDD.n5698 VDD.t1307 121.114
R12420 VDD.t1307 VDD.n5645 121.114
R12421 VDD.n5444 VDD.t270 121.114
R12422 VDD.t270 VDD.n5391 121.114
R12423 VDD.n3633 VDD.t249 121.114
R12424 VDD.t249 VDD.n3580 121.114
R12425 VDD.n3891 VDD.t1317 121.114
R12426 VDD.t1317 VDD.n3838 121.114
R12427 VDD.n4149 VDD.t409 121.114
R12428 VDD.t409 VDD.n4096 121.114
R12429 VDD.n4407 VDD.t1108 121.114
R12430 VDD.t1108 VDD.n4354 121.114
R12431 VDD.n4665 VDD.t332 121.114
R12432 VDD.t332 VDD.n4612 121.114
R12433 VDD.n4923 VDD.t279 121.114
R12434 VDD.t279 VDD.n4870 121.114
R12435 VDD.n5181 VDD.t1060 121.114
R12436 VDD.t1060 VDD.n5128 121.114
R12437 VDD.t557 VDD.t351 120.909
R12438 VDD.t1493 VDD.t328 120.909
R12439 VDD.t1376 VDD.t801 120.909
R12440 VDD.t1486 VDD.t804 120.909
R12441 VDD.n1853 VDD.n1845 120.094
R12442 VDD.n2174 VDD.n2166 120.094
R12443 VDD.n2432 VDD.n2424 120.094
R12444 VDD.n2690 VDD.n2682 120.094
R12445 VDD.n2948 VDD.n2940 120.094
R12446 VDD.n3206 VDD.n3198 120.094
R12447 VDD.n3464 VDD.n3456 120.094
R12448 VDD.n5784 VDD.n5776 120.094
R12449 VDD.n5530 VDD.n5522 120.094
R12450 VDD.n3722 VDD.n3714 120.094
R12451 VDD.n3980 VDD.n3972 120.094
R12452 VDD.n4238 VDD.n4230 120.094
R12453 VDD.n4496 VDD.n4488 120.094
R12454 VDD.n4754 VDD.n4746 120.094
R12455 VDD.n5012 VDD.n5004 120.094
R12456 VDD.n5270 VDD.n5262 120.094
R12457 VDD.n1 VDD.t361 117.451
R12458 VDD.n468 VDD.t1496 117.451
R12459 VDD.n439 VDD.t350 117.451
R12460 VDD.n459 VDD.t1497 117.451
R12461 VDD.n66 VDD.t1490 117.451
R12462 VDD.n36 VDD.t794 117.451
R12463 VDD.n56 VDD.t1488 117.451
R12464 VDD.n1145 VDD.t814 117.451
R12465 VDD.n5 VDD.t456 116.322
R12466 VDD.n494 VDD.t558 116.322
R12467 VDD.n422 VDD.t1478 116.322
R12468 VDD.n418 VDD.t327 116.322
R12469 VDD.n401 VDD.t1347 116.322
R12470 VDD.n92 VDD.t1377 116.322
R12471 VDD.n1149 VDD.t463 116.322
R12472 VDD.n1580 VDD.t510 116.322
R12473 VDD.n1576 VDD.t1044 116.322
R12474 VDD.n1559 VDD.t501 116.322
R12475 VDD.n806 VDD.t357 116.322
R12476 VDD.n1189 VDD.t808 116.322
R12477 VDD.n1768 VDD.n1767 116.267
R12478 VDD.n2117 VDD.n2116 116.267
R12479 VDD.n2347 VDD.n2346 116.267
R12480 VDD.n2605 VDD.n2604 116.267
R12481 VDD.n2863 VDD.n2862 116.267
R12482 VDD.n3121 VDD.n3120 116.267
R12483 VDD.n3379 VDD.n3378 116.267
R12484 VDD.n5702 VDD.n5701 116.267
R12485 VDD.n5448 VDD.n5447 116.267
R12486 VDD.n3637 VDD.n3636 116.267
R12487 VDD.n3895 VDD.n3894 116.267
R12488 VDD.n4153 VDD.n4152 116.267
R12489 VDD.n4411 VDD.n4410 116.267
R12490 VDD.n4669 VDD.n4668 116.267
R12491 VDD.n4927 VDD.n4926 116.267
R12492 VDD.n5185 VDD.n5184 116.267
R12493 VDD.t613 VDD.t356 115.486
R12494 VDD.t534 VDD.t807 115.486
R12495 VDD.n670 VDD 115.358
R12496 VDD.n1020 VDD 115.358
R12497 VDD.t728 VDD.n262 115.358
R12498 VDD.n1907 VDD.n1888 112.189
R12499 VDD.n1854 VDD.n1843 112.189
R12500 VDD.n2175 VDD.n2164 112.189
R12501 VDD.n2228 VDD.n2209 112.189
R12502 VDD.n2433 VDD.n2422 112.189
R12503 VDD.n2486 VDD.n2467 112.189
R12504 VDD.n2691 VDD.n2680 112.189
R12505 VDD.n2744 VDD.n2725 112.189
R12506 VDD.n2949 VDD.n2938 112.189
R12507 VDD.n3002 VDD.n2983 112.189
R12508 VDD.n3207 VDD.n3196 112.189
R12509 VDD.n3260 VDD.n3241 112.189
R12510 VDD.n3465 VDD.n3454 112.189
R12511 VDD.n3518 VDD.n3499 112.189
R12512 VDD.n5785 VDD.n5774 112.189
R12513 VDD.n5838 VDD.n5819 112.189
R12514 VDD.n5531 VDD.n5520 112.189
R12515 VDD.n5584 VDD.n5565 112.189
R12516 VDD.n3723 VDD.n3712 112.189
R12517 VDD.n3776 VDD.n3757 112.189
R12518 VDD.n3981 VDD.n3970 112.189
R12519 VDD.n4034 VDD.n4015 112.189
R12520 VDD.n4239 VDD.n4228 112.189
R12521 VDD.n4292 VDD.n4273 112.189
R12522 VDD.n4497 VDD.n4486 112.189
R12523 VDD.n4550 VDD.n4531 112.189
R12524 VDD.n4755 VDD.n4744 112.189
R12525 VDD.n4808 VDD.n4789 112.189
R12526 VDD.n5013 VDD.n5002 112.189
R12527 VDD.n5066 VDD.n5047 112.189
R12528 VDD.n5271 VDD.n5260 112.189
R12529 VDD.n5324 VDD.n5305 112.189
R12530 VDD.t345 VDD.t491 110.834
R12531 VDD.t785 VDD.t645 110.834
R12532 VDD.t1130 VDD.t1240 109.316
R12533 VDD.t1202 VDD.t1130 109.316
R12534 VDD.t1230 VDD.t1202 109.316
R12535 VDD.t1152 VDD.t1230 109.316
R12536 VDD.t1188 VDD.t1152 109.316
R12537 VDD.t1234 VDD.t1188 109.316
R12538 VDD.t1156 VDD.t1234 109.316
R12539 VDD.t1192 VDD.t1156 109.316
R12540 VDD.t1180 VDD.t1192 109.316
R12541 VDD.t1214 VDD.t1180 109.316
R12542 VDD.t1238 VDD.t1214 109.316
R12543 VDD.t1186 VDD.t1238 109.316
R12544 VDD.t1218 VDD.t1186 109.316
R12545 VDD.t1144 VDD.t1218 109.316
R12546 VDD.t1170 VDD.t1144 109.316
R12547 VDD.t1226 VDD.t1148 109.316
R12548 VDD.t1148 VDD.t1182 109.316
R12549 VDD.t1182 VDD.t1134 109.316
R12550 VDD.t1134 VDD.t1224 109.316
R12551 VDD.t1224 VDD.t1248 109.316
R12552 VDD.t1248 VDD.t1176 109.316
R12553 VDD.t1176 VDD.t1208 109.316
R12554 VDD.t1160 VDD.t1236 109.316
R12555 VDD.t1212 VDD.t1160 109.316
R12556 VDD.t1138 VDD.t1212 109.316
R12557 VDD.t1164 VDD.t1138 109.316
R12558 VDD.t1196 VDD.t1164 109.316
R12559 VDD.t1132 VDD.t1196 109.316
R12560 VDD.t1222 VDD.t1132 109.316
R12561 VDD.t1128 VDD.t1200 109.316
R12562 VDD.t1142 VDD.t1168 109.316
R12563 VDD.t1168 VDD.t1220 109.316
R12564 VDD.t1198 VDD.t1228 109.316
R12565 VDD.t1228 VDD.t1150 109.316
R12566 VDD.t1150 VDD.t1246 109.316
R12567 VDD.t1206 VDD.t1174 109.316
R12568 VDD.t1250 VDD.t1206 109.316
R12569 VDD.t1178 VDD.t1250 109.316
R12570 VDD.t1210 VDD.t1136 109.316
R12571 VDD.t1136 VDD.t1162 109.316
R12572 VDD.t1162 VDD.t1194 109.316
R12573 VDD.t1194 VDD.t1140 109.316
R12574 VDD.t1140 VDD.t1166 109.316
R12575 VDD.t1166 VDD.t1244 109.316
R12576 VDD.t318 VDD.t324 109.316
R12577 VDD.t324 VDD.t302 109.316
R12578 VDD.t302 VDD.t312 109.316
R12579 VDD.t304 VDD.t322 109.316
R12580 VDD.t314 VDD.t304 109.316
R12581 VDD.t294 VDD.t314 109.316
R12582 VDD.t300 VDD.t310 109.316
R12583 VDD.t310 VDD.t306 109.316
R12584 VDD.t306 VDD.t320 109.316
R12585 VDD.t308 VDD.t298 109.316
R12586 VDD.t316 VDD.t308 109.316
R12587 VDD.t1276 VDD.t1272 109.316
R12588 VDD.t1272 VDD.t1274 109.316
R12589 VDD.t1274 VDD.t1278 109.316
R12590 VDD.t175 VDD.n667 108.572
R12591 VDD.t948 VDD.n1017 108.572
R12592 VDD.n265 VDD 108.572
R12593 VDD.t471 VDD.t605 106.709
R12594 VDD.t289 VDD.t651 106.709
R12595 VDD.t598 VDD.t1066 103.636
R12596 VDD.t595 VDD.t457 103.636
R12597 VDD.n1769 VDD.n1768 102.721
R12598 VDD.n1755 VDD.n1671 102.721
R12599 VDD.n2118 VDD.n2117 102.721
R12600 VDD.n2104 VDD.n2020 102.721
R12601 VDD.n2348 VDD.n2347 102.721
R12602 VDD.n2334 VDD.n2250 102.721
R12603 VDD.n2606 VDD.n2605 102.721
R12604 VDD.n2592 VDD.n2508 102.721
R12605 VDD.n2864 VDD.n2863 102.721
R12606 VDD.n2850 VDD.n2766 102.721
R12607 VDD.n3122 VDD.n3121 102.721
R12608 VDD.n3108 VDD.n3024 102.721
R12609 VDD.n3380 VDD.n3379 102.721
R12610 VDD.n3366 VDD.n3282 102.721
R12611 VDD.n5703 VDD.n5702 102.721
R12612 VDD.n5689 VDD.n5605 102.721
R12613 VDD.n5449 VDD.n5448 102.721
R12614 VDD.n5435 VDD.n5351 102.721
R12615 VDD.n3638 VDD.n3637 102.721
R12616 VDD.n3624 VDD.n3540 102.721
R12617 VDD.n3896 VDD.n3895 102.721
R12618 VDD.n3882 VDD.n3798 102.721
R12619 VDD.n4154 VDD.n4153 102.721
R12620 VDD.n4140 VDD.n4056 102.721
R12621 VDD.n4412 VDD.n4411 102.721
R12622 VDD.n4398 VDD.n4314 102.721
R12623 VDD.n4670 VDD.n4669 102.721
R12624 VDD.n4656 VDD.n4572 102.721
R12625 VDD.n4928 VDD.n4927 102.721
R12626 VDD.n4914 VDD.n4830 102.721
R12627 VDD.n5186 VDD.n5185 102.721
R12628 VDD.n5172 VDD.n5088 102.721
R12629 VDD VDD.t1170 101.507
R12630 VDD.t1220 VDD 101.507
R12631 VDD.t1244 VDD 101.507
R12632 VDD.t296 VDD 101.507
R12633 VDD.t464 VDD 99.5973
R12634 VDD.t255 VDD 99.5973
R12635 VDD.t1017 VDD 99.5973
R12636 VDD.t1323 VDD 99.5973
R12637 VDD.t366 VDD 99.5973
R12638 VDD.t1459 VDD 99.5973
R12639 VDD.t1293 VDD 99.5973
R12640 VDD.t601 VDD 99.5973
R12641 VDD.t643 VDD 99.5973
R12642 VDD.t253 VDD 99.5973
R12643 VDD.t268 VDD 99.5973
R12644 VDD.t15 VDD 99.5973
R12645 VDD.t1067 VDD 99.5973
R12646 VDD.t1309 VDD 99.5973
R12647 VDD.t817 VDD 99.5973
R12648 VDD.t1058 VDD 99.5973
R12649 VDD VDD.t362 99.5409
R12650 VDD VDD.t509 99.5409
R12651 VDD.t1345 VDD.t1110 98.9875
R12652 VDD.t334 VDD.t1107 98.9875
R12653 VDD.t577 VDD.t1005 98.9875
R12654 VDD.t837 VDD.t1426 98.9875
R12655 VDD.n1429 VDD.t1178 98.9046
R12656 VDD.t1103 VDD.t71 97.8793
R12657 VDD.t1452 VDD.t629 97.8793
R12658 VDD.t1278 VDD 97.6032
R12659 VDD.n31 VDD.t1465 96.1553
R12660 VDD.n672 VDD.t604 96.1553
R12661 VDD.n508 VDD.t469 96.1553
R12662 VDD.n435 VDD.t966 96.1553
R12663 VDD.n404 VDD.t1342 96.1553
R12664 VDD.n106 VDD.t288 96.1553
R12665 VDD.n1175 VDD.t452 96.1553
R12666 VDD.n1593 VDD.t1286 96.1553
R12667 VDD.n1562 VDD.t824 96.1553
R12668 VDD.n800 VDD.t1097 96.1553
R12669 VDD.n803 VDD.t1091 96.1553
R12670 VDD.n1022 VDD.t1352 96.1553
R12671 VDD.n267 VDD.t1357 96.1553
R12672 VDD.n1183 VDD.t259 96.1553
R12673 VDD.n1186 VDD.t1283 96.1553
R12674 VDD.n585 VDD.t151 95.0005
R12675 VDD.n935 VDD.t924 95.0005
R12676 VDD.t836 VDD 94.8523
R12677 VDD.t538 VDD 94.8523
R12678 VDD.n482 VDD.t346 93.81
R12679 VDD.n80 VDD.t786 93.81
R12680 VDD.t328 VDD 93.5611
R12681 VDD.t804 VDD 93.5611
R12682 VDD.t257 VDD 93.539
R12683 VDD.t1013 VDD 93.539
R12684 VDD VDD.t1345 93.4882
R12685 VDD VDD.t577 93.4882
R12686 VDD.t1064 VDD 93.3702
R12687 VDD.t971 VDD 93.3702
R12688 VDD.n1733 VDD.n1730 92.5005
R12689 VDD.n2082 VDD.n2079 92.5005
R12690 VDD.n2312 VDD.n2309 92.5005
R12691 VDD.n2570 VDD.n2567 92.5005
R12692 VDD.n2828 VDD.n2825 92.5005
R12693 VDD.n3086 VDD.n3083 92.5005
R12694 VDD.n3344 VDD.n3341 92.5005
R12695 VDD.n5667 VDD.n5664 92.5005
R12696 VDD.n5413 VDD.n5410 92.5005
R12697 VDD.n3602 VDD.n3599 92.5005
R12698 VDD.n3860 VDD.n3857 92.5005
R12699 VDD.n4118 VDD.n4115 92.5005
R12700 VDD.n4376 VDD.n4373 92.5005
R12701 VDD.n4634 VDD.n4631 92.5005
R12702 VDD.n4892 VDD.n4889 92.5005
R12703 VDD.n5150 VDD.n5147 92.5005
R12704 VDD.t559 VDD 92.1217
R12705 VDD.t1443 VDD 92.1217
R12706 VDD.t69 VDD.t358 91.8882
R12707 VDD.t627 VDD.t810 91.8882
R12708 VDD.n1915 VDD.n1891 91.7652
R12709 VDD.n2236 VDD.n2212 91.7652
R12710 VDD.n2494 VDD.n2470 91.7652
R12711 VDD.n2752 VDD.n2728 91.7652
R12712 VDD.n3010 VDD.n2986 91.7652
R12713 VDD.n3268 VDD.n3244 91.7652
R12714 VDD.n3526 VDD.n3502 91.7652
R12715 VDD.n5846 VDD.n5822 91.7652
R12716 VDD.n5592 VDD.n5568 91.7652
R12717 VDD.n3784 VDD.n3760 91.7652
R12718 VDD.n4042 VDD.n4018 91.7652
R12719 VDD.n4300 VDD.n4276 91.7652
R12720 VDD.n4558 VDD.n4534 91.7652
R12721 VDD.n4816 VDD.n4792 91.7652
R12722 VDD.n5074 VDD.n5050 91.7652
R12723 VDD.n5332 VDD.n5308 91.7652
R12724 VDD.t698 VDD.n183 91.6076
R12725 VDD.n1960 VDD.n1959 91.4829
R12726 VDD.n1959 VDD.n1929 91.4829
R12727 VDD.n1972 VDD.n1929 91.4829
R12728 VDD.n1972 VDD.n1971 91.4829
R12729 VDD.n1950 VDD.n1937 91.4829
R12730 VDD.n1965 VDD.n1937 91.4829
R12731 VDD.n1966 VDD.n1965 91.4829
R12732 VDD.n1967 VDD.n1966 91.4829
R12733 VDD.n1884 VDD.n1820 91.343
R12734 VDD.n2205 VDD.n2141 91.343
R12735 VDD.n2463 VDD.n2399 91.343
R12736 VDD.n2721 VDD.n2657 91.343
R12737 VDD.n2979 VDD.n2915 91.343
R12738 VDD.n3237 VDD.n3173 91.343
R12739 VDD.n3495 VDD.n3431 91.343
R12740 VDD.n5815 VDD.n5751 91.343
R12741 VDD.n5561 VDD.n5497 91.343
R12742 VDD.n3753 VDD.n3689 91.343
R12743 VDD.n4011 VDD.n3947 91.343
R12744 VDD.n4269 VDD.n4205 91.343
R12745 VDD.n4527 VDD.n4463 91.343
R12746 VDD.n4785 VDD.n4721 91.343
R12747 VDD.n5043 VDD.n4979 91.343
R12748 VDD.n5301 VDD.n5237 91.343
R12749 VDD.n1372 VDD.t316 91.0964
R12750 VDD.n1827 VDD.t599 89.1694
R12751 VDD.n2148 VDD.t1011 89.1694
R12752 VDD.n2406 VDD.t615 89.1694
R12753 VDD.n2664 VDD.t247 89.1694
R12754 VDD.n2922 VDD.t618 89.1694
R12755 VDD.n3180 VDD.t647 89.1694
R12756 VDD.n3438 VDD.t532 89.1694
R12757 VDD.n5758 VDD.t1353 89.1694
R12758 VDD.n5504 VDD.t391 89.1694
R12759 VDD.n3696 VDD.t291 89.1694
R12760 VDD.n3954 VDD.t1348 89.1694
R12761 VDD.n4212 VDD.t1363 89.1694
R12762 VDD.n4470 VDD.t608 89.1694
R12763 VDD.n4728 VDD.t399 89.1694
R12764 VDD.n4986 VDD.t1099 89.1694
R12765 VDD.n5244 VDD.t405 89.1694
R12766 VDD.t360 VDD.t449 88.9241
R12767 VDD.t813 VDD.t565 88.9241
R12768 VDD VDD.n1371 88.4936
R12769 VDD.n184 VDD.t704 88.2148
R12770 VDD VDD.t782 87.9889
R12771 VDD VDD.t428 87.9889
R12772 VDD.t637 VDD 87.8035
R12773 VDD.t431 VDD 87.8035
R12774 VDD.t1441 VDD.t1316 87.6928
R12775 VDD.t1321 VDD.t347 87.6928
R12776 VDD.t539 VDD.t1359 87.6928
R12777 VDD.t1303 VDD.t788 87.6928
R12778 VDD.n7 VDD.t1123 86.7743
R12779 VDD.n7 VDD.t70 86.7743
R12780 VDD.n471 VDD.t72 86.7743
R12781 VDD.n471 VDD.t492 86.7743
R12782 VDD.n441 VDD.t1121 86.7743
R12783 VDD.n441 VDD.t74 86.7743
R12784 VDD.n443 VDD.t378 86.7743
R12785 VDD.n443 VDD.t281 86.7743
R12786 VDD.n69 VDD.t630 86.7743
R12787 VDD.n69 VDD.t646 86.7743
R12788 VDD.n38 VDD.t1456 86.7743
R12789 VDD.n38 VDD.t631 86.7743
R12790 VDD.n40 VDD.t472 86.7743
R12791 VDD.n40 VDD.t286 86.7743
R12792 VDD.n1151 VDD.t1458 86.7743
R12793 VDD.n1151 VDD.t628 86.7743
R12794 VDD.t145 VDD.n584 84.8219
R12795 VDD.t918 VDD.n934 84.8219
R12796 VDD.n438 VDD.n408 83.3098
R12797 VDD.n1596 VDD.n1566 83.3098
R12798 VDD.n1827 VDD.t1088 81.2688
R12799 VDD.n2148 VDD.t555 81.2688
R12800 VDD.n2406 VDD.t1383 81.2688
R12801 VDD.n2664 VDD.t575 81.2688
R12802 VDD.n2922 VDD.t1479 81.2688
R12803 VDD.n3180 VDD.t1003 81.2688
R12804 VDD.n3438 VDD.t397 81.2688
R12805 VDD.n5758 VDD.t67 81.2688
R12806 VDD.n5504 VDD.t1305 81.2688
R12807 VDD.n3696 VDD.t1070 81.2688
R12808 VDD.n3954 VDD.t1062 81.2688
R12809 VDD.n4212 VDD.t984 81.2688
R12810 VDD.n4470 VDD.t458 81.2688
R12811 VDD.n4728 VDD.t1474 81.2688
R12812 VDD.n4986 VDD.t1042 81.2688
R12813 VDD.n5244 VDD.t633 81.2688
R12814 VDD.n1457 VDD.t1222 80.6854
R12815 VDD.n1760 VDD.n1717 80.5087
R12816 VDD.n2109 VDD.n2066 80.5087
R12817 VDD.n2339 VDD.n2296 80.5087
R12818 VDD.n2597 VDD.n2554 80.5087
R12819 VDD.n2855 VDD.n2812 80.5087
R12820 VDD.n3113 VDD.n3070 80.5087
R12821 VDD.n3371 VDD.n3328 80.5087
R12822 VDD.n5694 VDD.n5651 80.5087
R12823 VDD.n5440 VDD.n5397 80.5087
R12824 VDD.n3629 VDD.n3586 80.5087
R12825 VDD.n3887 VDD.n3844 80.5087
R12826 VDD.n4145 VDD.n4102 80.5087
R12827 VDD.n4403 VDD.n4360 80.5087
R12828 VDD.n4661 VDD.n4618 80.5087
R12829 VDD.n4919 VDD.n4876 80.5087
R12830 VDD.n5177 VDD.n5134 80.5087
R12831 VDD.n1708 VDD.n1669 80.2452
R12832 VDD.n2057 VDD.n2018 80.2452
R12833 VDD.n2287 VDD.n2248 80.2452
R12834 VDD.n2545 VDD.n2506 80.2452
R12835 VDD.n2803 VDD.n2764 80.2452
R12836 VDD.n3061 VDD.n3022 80.2452
R12837 VDD.n3319 VDD.n3280 80.2452
R12838 VDD.n5642 VDD.n5603 80.2452
R12839 VDD.n5388 VDD.n5349 80.2452
R12840 VDD.n3577 VDD.n3538 80.2452
R12841 VDD.n3835 VDD.n3796 80.2452
R12842 VDD.n4093 VDD.n4054 80.2452
R12843 VDD.n4351 VDD.n4312 80.2452
R12844 VDD.n4609 VDD.n4570 80.2452
R12845 VDD.n4867 VDD.n4828 80.2452
R12846 VDD.n5125 VDD.n5086 80.2452
R12847 VDD VDD.n1643 79.5475
R12848 VDD.t1200 VDD.t1242 78.5727
R12849 VDD VDD.n1634 78.5148
R12850 VDD.n1633 VDD.n1632 77.1383
R12851 VDD.n1870 VDD.n1845 76.5328
R12852 VDD.n2191 VDD.n2166 76.5328
R12853 VDD.n2449 VDD.n2424 76.5328
R12854 VDD.n2707 VDD.n2682 76.5328
R12855 VDD.n2965 VDD.n2940 76.5328
R12856 VDD.n3223 VDD.n3198 76.5328
R12857 VDD.n3481 VDD.n3456 76.5328
R12858 VDD.n5801 VDD.n5776 76.5328
R12859 VDD.n5547 VDD.n5522 76.5328
R12860 VDD.n3739 VDD.n3714 76.5328
R12861 VDD.n3997 VDD.n3972 76.5328
R12862 VDD.n4255 VDD.n4230 76.5328
R12863 VDD.n4513 VDD.n4488 76.5328
R12864 VDD.n4771 VDD.n4746 76.5328
R12865 VDD.n5029 VDD.n5004 76.5328
R12866 VDD.n5287 VDD.n5262 76.5328
R12867 VDD.n1625 VDD.n1624 76.0005
R12868 VDD.n1628 VDD.n1627 76.0005
R12869 VDD.n1630 VDD.n1629 76.0005
R12870 VDD.n1397 VDD.t294 75.48
R12871 VDD.n1869 VDD.n1844 74.1181
R12872 VDD.n2190 VDD.n2165 74.1181
R12873 VDD.n2448 VDD.n2423 74.1181
R12874 VDD.n2706 VDD.n2681 74.1181
R12875 VDD.n2964 VDD.n2939 74.1181
R12876 VDD.n3222 VDD.n3197 74.1181
R12877 VDD.n3480 VDD.n3455 74.1181
R12878 VDD.n5800 VDD.n5775 74.1181
R12879 VDD.n5546 VDD.n5521 74.1181
R12880 VDD.n3738 VDD.n3713 74.1181
R12881 VDD.n3996 VDD.n3971 74.1181
R12882 VDD.n4254 VDD.n4229 74.1181
R12883 VDD.n4512 VDD.n4487 74.1181
R12884 VDD.n4770 VDD.n4745 74.1181
R12885 VDD.n5028 VDD.n5003 74.1181
R12886 VDD.n5286 VDD.n5261 74.1181
R12887 VDD.n1871 VDD.n1843 71.6136
R12888 VDD.n2192 VDD.n2164 71.6136
R12889 VDD.n2450 VDD.n2422 71.6136
R12890 VDD.n2708 VDD.n2680 71.6136
R12891 VDD.n2966 VDD.n2938 71.6136
R12892 VDD.n3224 VDD.n3196 71.6136
R12893 VDD.n3482 VDD.n3454 71.6136
R12894 VDD.n5802 VDD.n5774 71.6136
R12895 VDD.n5548 VDD.n5520 71.6136
R12896 VDD.n3740 VDD.n3712 71.6136
R12897 VDD.n3998 VDD.n3970 71.6136
R12898 VDD.n4256 VDD.n4228 71.6136
R12899 VDD.n4514 VDD.n4486 71.6136
R12900 VDD.n4772 VDD.n4744 71.6136
R12901 VDD.n5030 VDD.n5002 71.6136
R12902 VDD.n5288 VDD.n5260 71.6136
R12903 VDD.n1809 VDD.t464 70.4844
R12904 VDD.n2130 VDD.t255 70.4844
R12905 VDD.n2388 VDD.t1017 70.4844
R12906 VDD.n2646 VDD.t1323 70.4844
R12907 VDD.n2904 VDD.t366 70.4844
R12908 VDD.n3162 VDD.t1459 70.4844
R12909 VDD.n3420 VDD.t1293 70.4844
R12910 VDD.n5740 VDD.t601 70.4844
R12911 VDD.n5486 VDD.t643 70.4844
R12912 VDD.n3678 VDD.t253 70.4844
R12913 VDD.n3936 VDD.t268 70.4844
R12914 VDD.n4194 VDD.t15 70.4844
R12915 VDD.n4452 VDD.t1067 70.4844
R12916 VDD.n4710 VDD.t1309 70.4844
R12917 VDD.n4968 VDD.t817 70.4844
R12918 VDD.n5226 VDD.t1058 70.4844
R12919 VDD.t1316 VDD.t1346 70.1543
R12920 VDD.t1359 VDD.t500 70.1543
R12921 VDD.n1877 VDD.n1876 66.2808
R12922 VDD.n2198 VDD.n2197 66.2808
R12923 VDD.n2456 VDD.n2455 66.2808
R12924 VDD.n2714 VDD.n2713 66.2808
R12925 VDD.n2972 VDD.n2971 66.2808
R12926 VDD.n3230 VDD.n3229 66.2808
R12927 VDD.n3488 VDD.n3487 66.2808
R12928 VDD.n5808 VDD.n5807 66.2808
R12929 VDD.n5554 VDD.n5553 66.2808
R12930 VDD.n3746 VDD.n3745 66.2808
R12931 VDD.n4004 VDD.n4003 66.2808
R12932 VDD.n4262 VDD.n4261 66.2808
R12933 VDD.n4520 VDD.n4519 66.2808
R12934 VDD.n4778 VDD.n4777 66.2808
R12935 VDD.n5036 VDD.n5035 66.2808
R12936 VDD.n5294 VDD.n5293 66.2808
R12937 VDD.n1898 VDD.n1889 65.0929
R12938 VDD.n2219 VDD.n2210 65.0929
R12939 VDD.n2477 VDD.n2468 65.0929
R12940 VDD.n2735 VDD.n2726 65.0929
R12941 VDD.n2993 VDD.n2984 65.0929
R12942 VDD.n3251 VDD.n3242 65.0929
R12943 VDD.n3509 VDD.n3500 65.0929
R12944 VDD.n5829 VDD.n5820 65.0929
R12945 VDD.n5575 VDD.n5566 65.0929
R12946 VDD.n3767 VDD.n3758 65.0929
R12947 VDD.n4025 VDD.n4016 65.0929
R12948 VDD.n4283 VDD.n4274 65.0929
R12949 VDD.n4541 VDD.n4532 65.0929
R12950 VDD.n4799 VDD.n4790 65.0929
R12951 VDD.n5057 VDD.n5048 65.0929
R12952 VDD.n5315 VDD.n5306 65.0929
R12953 VDD.n1809 VDD.t1498 64.3553
R12954 VDD.n2130 VDD.t625 64.3553
R12955 VDD.n2388 VDD.t1284 64.3553
R12956 VDD.n2646 VDD.t85 64.3553
R12957 VDD.n2904 VDD.t272 64.3553
R12958 VDD.n3162 VDD.t541 64.3553
R12959 VDD.n3420 VDD.t1280 64.3553
R12960 VDD.n5740 VDD.t519 64.3553
R12961 VDD.n5486 VDD.t453 64.3553
R12962 VDD.n3678 VDD.t1101 64.3553
R12963 VDD.n3936 VDD.t1048 64.3553
R12964 VDD.n4194 VDD.t1462 64.3553
R12965 VDD.n4452 VDD.t1105 64.3553
R12966 VDD.n4710 VDD.t1500 64.3553
R12967 VDD.n4968 VDD.t1288 64.3553
R12968 VDD.n5226 VDD.t481 64.3553
R12969 VDD.n475 VDD.t1494 63.3219
R12970 VDD.n475 VDD.t329 63.3219
R12971 VDD.n73 VDD.t1487 63.3219
R12972 VDD.n73 VDD.t1358 63.3219
R12973 VDD.n1706 VDD.n1673 63.2691
R12974 VDD.n1707 VDD.n1706 63.2691
R12975 VDD.n2055 VDD.n2022 63.2691
R12976 VDD.n2056 VDD.n2055 63.2691
R12977 VDD.n2285 VDD.n2252 63.2691
R12978 VDD.n2286 VDD.n2285 63.2691
R12979 VDD.n2543 VDD.n2510 63.2691
R12980 VDD.n2544 VDD.n2543 63.2691
R12981 VDD.n2801 VDD.n2768 63.2691
R12982 VDD.n2802 VDD.n2801 63.2691
R12983 VDD.n3059 VDD.n3026 63.2691
R12984 VDD.n3060 VDD.n3059 63.2691
R12985 VDD.n3317 VDD.n3284 63.2691
R12986 VDD.n3318 VDD.n3317 63.2691
R12987 VDD.n5640 VDD.n5607 63.2691
R12988 VDD.n5641 VDD.n5640 63.2691
R12989 VDD.n5386 VDD.n5353 63.2691
R12990 VDD.n5387 VDD.n5386 63.2691
R12991 VDD.n3575 VDD.n3542 63.2691
R12992 VDD.n3576 VDD.n3575 63.2691
R12993 VDD.n3833 VDD.n3800 63.2691
R12994 VDD.n3834 VDD.n3833 63.2691
R12995 VDD.n4091 VDD.n4058 63.2691
R12996 VDD.n4092 VDD.n4091 63.2691
R12997 VDD.n4349 VDD.n4316 63.2691
R12998 VDD.n4350 VDD.n4349 63.2691
R12999 VDD.n4607 VDD.n4574 63.2691
R13000 VDD.n4608 VDD.n4607 63.2691
R13001 VDD.n4865 VDD.n4832 63.2691
R13002 VDD.n4866 VDD.n4865 63.2691
R13003 VDD.n5123 VDD.n5090 63.2691
R13004 VDD.n5124 VDD.n5123 63.2691
R13005 VDD.n1762 VDD.n1715 61.5116
R13006 VDD.n1762 VDD.n1761 61.5116
R13007 VDD.n2111 VDD.n2064 61.5116
R13008 VDD.n2111 VDD.n2110 61.5116
R13009 VDD.n2341 VDD.n2294 61.5116
R13010 VDD.n2341 VDD.n2340 61.5116
R13011 VDD.n2599 VDD.n2552 61.5116
R13012 VDD.n2599 VDD.n2598 61.5116
R13013 VDD.n2857 VDD.n2810 61.5116
R13014 VDD.n2857 VDD.n2856 61.5116
R13015 VDD.n3115 VDD.n3068 61.5116
R13016 VDD.n3115 VDD.n3114 61.5116
R13017 VDD.n3373 VDD.n3326 61.5116
R13018 VDD.n3373 VDD.n3372 61.5116
R13019 VDD.n5696 VDD.n5649 61.5116
R13020 VDD.n5696 VDD.n5695 61.5116
R13021 VDD.n5442 VDD.n5395 61.5116
R13022 VDD.n5442 VDD.n5441 61.5116
R13023 VDD.n3631 VDD.n3584 61.5116
R13024 VDD.n3631 VDD.n3630 61.5116
R13025 VDD.n3889 VDD.n3842 61.5116
R13026 VDD.n3889 VDD.n3888 61.5116
R13027 VDD.n4147 VDD.n4100 61.5116
R13028 VDD.n4147 VDD.n4146 61.5116
R13029 VDD.n4405 VDD.n4358 61.5116
R13030 VDD.n4405 VDD.n4404 61.5116
R13031 VDD.n4663 VDD.n4616 61.5116
R13032 VDD.n4663 VDD.n4662 61.5116
R13033 VDD.n4921 VDD.n4874 61.5116
R13034 VDD.n4921 VDD.n4920 61.5116
R13035 VDD.n5179 VDD.n5132 61.5116
R13036 VDD.n5179 VDD.n5178 61.5116
R13037 VDD.n1908 VDD.n1897 60.6123
R13038 VDD.n1911 VDD.n1910 60.6123
R13039 VDD.n1910 VDD.n1903 60.6123
R13040 VDD.n1908 VDD.n1907 60.6123
R13041 VDD.n1860 VDD.n1852 60.6123
R13042 VDD.n1866 VDD.n1853 60.6123
R13043 VDD.n1866 VDD.n1865 60.6123
R13044 VDD.n1854 VDD.n1852 60.6123
R13045 VDD.n2181 VDD.n2173 60.6123
R13046 VDD.n2187 VDD.n2174 60.6123
R13047 VDD.n2187 VDD.n2186 60.6123
R13048 VDD.n2175 VDD.n2173 60.6123
R13049 VDD.n2229 VDD.n2218 60.6123
R13050 VDD.n2232 VDD.n2231 60.6123
R13051 VDD.n2231 VDD.n2224 60.6123
R13052 VDD.n2229 VDD.n2228 60.6123
R13053 VDD.n2439 VDD.n2431 60.6123
R13054 VDD.n2445 VDD.n2432 60.6123
R13055 VDD.n2445 VDD.n2444 60.6123
R13056 VDD.n2433 VDD.n2431 60.6123
R13057 VDD.n2487 VDD.n2476 60.6123
R13058 VDD.n2490 VDD.n2489 60.6123
R13059 VDD.n2489 VDD.n2482 60.6123
R13060 VDD.n2487 VDD.n2486 60.6123
R13061 VDD.n2697 VDD.n2689 60.6123
R13062 VDD.n2703 VDD.n2690 60.6123
R13063 VDD.n2703 VDD.n2702 60.6123
R13064 VDD.n2691 VDD.n2689 60.6123
R13065 VDD.n2745 VDD.n2734 60.6123
R13066 VDD.n2748 VDD.n2747 60.6123
R13067 VDD.n2747 VDD.n2740 60.6123
R13068 VDD.n2745 VDD.n2744 60.6123
R13069 VDD.n2955 VDD.n2947 60.6123
R13070 VDD.n2961 VDD.n2948 60.6123
R13071 VDD.n2961 VDD.n2960 60.6123
R13072 VDD.n2949 VDD.n2947 60.6123
R13073 VDD.n3003 VDD.n2992 60.6123
R13074 VDD.n3006 VDD.n3005 60.6123
R13075 VDD.n3005 VDD.n2998 60.6123
R13076 VDD.n3003 VDD.n3002 60.6123
R13077 VDD.n3213 VDD.n3205 60.6123
R13078 VDD.n3219 VDD.n3206 60.6123
R13079 VDD.n3219 VDD.n3218 60.6123
R13080 VDD.n3207 VDD.n3205 60.6123
R13081 VDD.n3261 VDD.n3250 60.6123
R13082 VDD.n3264 VDD.n3263 60.6123
R13083 VDD.n3263 VDD.n3256 60.6123
R13084 VDD.n3261 VDD.n3260 60.6123
R13085 VDD.n3471 VDD.n3463 60.6123
R13086 VDD.n3477 VDD.n3464 60.6123
R13087 VDD.n3477 VDD.n3476 60.6123
R13088 VDD.n3465 VDD.n3463 60.6123
R13089 VDD.n3519 VDD.n3508 60.6123
R13090 VDD.n3522 VDD.n3521 60.6123
R13091 VDD.n3521 VDD.n3514 60.6123
R13092 VDD.n3519 VDD.n3518 60.6123
R13093 VDD.n5791 VDD.n5783 60.6123
R13094 VDD.n5797 VDD.n5784 60.6123
R13095 VDD.n5797 VDD.n5796 60.6123
R13096 VDD.n5785 VDD.n5783 60.6123
R13097 VDD.n5839 VDD.n5828 60.6123
R13098 VDD.n5842 VDD.n5841 60.6123
R13099 VDD.n5841 VDD.n5834 60.6123
R13100 VDD.n5839 VDD.n5838 60.6123
R13101 VDD.n5537 VDD.n5529 60.6123
R13102 VDD.n5543 VDD.n5530 60.6123
R13103 VDD.n5543 VDD.n5542 60.6123
R13104 VDD.n5531 VDD.n5529 60.6123
R13105 VDD.n5585 VDD.n5574 60.6123
R13106 VDD.n5588 VDD.n5587 60.6123
R13107 VDD.n5587 VDD.n5580 60.6123
R13108 VDD.n5585 VDD.n5584 60.6123
R13109 VDD.n3729 VDD.n3721 60.6123
R13110 VDD.n3735 VDD.n3722 60.6123
R13111 VDD.n3735 VDD.n3734 60.6123
R13112 VDD.n3723 VDD.n3721 60.6123
R13113 VDD.n3777 VDD.n3766 60.6123
R13114 VDD.n3780 VDD.n3779 60.6123
R13115 VDD.n3779 VDD.n3772 60.6123
R13116 VDD.n3777 VDD.n3776 60.6123
R13117 VDD.n3987 VDD.n3979 60.6123
R13118 VDD.n3993 VDD.n3980 60.6123
R13119 VDD.n3993 VDD.n3992 60.6123
R13120 VDD.n3981 VDD.n3979 60.6123
R13121 VDD.n4035 VDD.n4024 60.6123
R13122 VDD.n4038 VDD.n4037 60.6123
R13123 VDD.n4037 VDD.n4030 60.6123
R13124 VDD.n4035 VDD.n4034 60.6123
R13125 VDD.n4245 VDD.n4237 60.6123
R13126 VDD.n4251 VDD.n4238 60.6123
R13127 VDD.n4251 VDD.n4250 60.6123
R13128 VDD.n4239 VDD.n4237 60.6123
R13129 VDD.n4293 VDD.n4282 60.6123
R13130 VDD.n4296 VDD.n4295 60.6123
R13131 VDD.n4295 VDD.n4288 60.6123
R13132 VDD.n4293 VDD.n4292 60.6123
R13133 VDD.n4503 VDD.n4495 60.6123
R13134 VDD.n4509 VDD.n4496 60.6123
R13135 VDD.n4509 VDD.n4508 60.6123
R13136 VDD.n4497 VDD.n4495 60.6123
R13137 VDD.n4551 VDD.n4540 60.6123
R13138 VDD.n4554 VDD.n4553 60.6123
R13139 VDD.n4553 VDD.n4546 60.6123
R13140 VDD.n4551 VDD.n4550 60.6123
R13141 VDD.n4761 VDD.n4753 60.6123
R13142 VDD.n4767 VDD.n4754 60.6123
R13143 VDD.n4767 VDD.n4766 60.6123
R13144 VDD.n4755 VDD.n4753 60.6123
R13145 VDD.n4809 VDD.n4798 60.6123
R13146 VDD.n4812 VDD.n4811 60.6123
R13147 VDD.n4811 VDD.n4804 60.6123
R13148 VDD.n4809 VDD.n4808 60.6123
R13149 VDD.n5019 VDD.n5011 60.6123
R13150 VDD.n5025 VDD.n5012 60.6123
R13151 VDD.n5025 VDD.n5024 60.6123
R13152 VDD.n5013 VDD.n5011 60.6123
R13153 VDD.n5067 VDD.n5056 60.6123
R13154 VDD.n5070 VDD.n5069 60.6123
R13155 VDD.n5069 VDD.n5062 60.6123
R13156 VDD.n5067 VDD.n5066 60.6123
R13157 VDD.n5277 VDD.n5269 60.6123
R13158 VDD.n5283 VDD.n5270 60.6123
R13159 VDD.n5283 VDD.n5282 60.6123
R13160 VDD.n5271 VDD.n5269 60.6123
R13161 VDD.n5325 VDD.n5314 60.6123
R13162 VDD.n5328 VDD.n5327 60.6123
R13163 VDD.n5327 VDD.n5320 60.6123
R13164 VDD.n5325 VDD.n5324 60.6123
R13165 VDD.n1456 VDD.t1198 59.8635
R13166 VDD.n1916 VDD.n1888 58.0325
R13167 VDD.n2237 VDD.n2209 58.0325
R13168 VDD.n2495 VDD.n2467 58.0325
R13169 VDD.n2753 VDD.n2725 58.0325
R13170 VDD.n3011 VDD.n2983 58.0325
R13171 VDD.n3269 VDD.n3241 58.0325
R13172 VDD.n3527 VDD.n3499 58.0325
R13173 VDD.n5847 VDD.n5819 58.0325
R13174 VDD.n5593 VDD.n5565 58.0325
R13175 VDD.n3785 VDD.n3757 58.0325
R13176 VDD.n4043 VDD.n4015 58.0325
R13177 VDD.n4301 VDD.n4273 58.0325
R13178 VDD.n4559 VDD.n4531 58.0325
R13179 VDD.n4817 VDD.n4789 58.0325
R13180 VDD.n5075 VDD.n5047 58.0325
R13181 VDD.n5333 VDD.n5305 58.0325
R13182 VDD.n584 VDD.t119 57.6791
R13183 VDD.n934 VDD.t890 57.6791
R13184 VDD.t351 VDD.t637 57.5763
R13185 VDD.t801 VDD.t431 57.5763
R13186 VDD VDD.t73 57.5434
R13187 VDD VDD.t426 57.5434
R13188 VDD.t358 VDD.t1064 56.3188
R13189 VDD.t810 VDD.t971 56.3188
R13190 VDD.n1732 VDD.n1731 55.4672
R13191 VDD.n1733 VDD.n1729 55.4672
R13192 VDD.n2081 VDD.n2080 55.4672
R13193 VDD.n2082 VDD.n2078 55.4672
R13194 VDD.n2311 VDD.n2310 55.4672
R13195 VDD.n2312 VDD.n2308 55.4672
R13196 VDD.n2569 VDD.n2568 55.4672
R13197 VDD.n2570 VDD.n2566 55.4672
R13198 VDD.n2827 VDD.n2826 55.4672
R13199 VDD.n2828 VDD.n2824 55.4672
R13200 VDD.n3085 VDD.n3084 55.4672
R13201 VDD.n3086 VDD.n3082 55.4672
R13202 VDD.n3343 VDD.n3342 55.4672
R13203 VDD.n3344 VDD.n3340 55.4672
R13204 VDD.n5666 VDD.n5665 55.4672
R13205 VDD.n5667 VDD.n5663 55.4672
R13206 VDD.n5412 VDD.n5411 55.4672
R13207 VDD.n5413 VDD.n5409 55.4672
R13208 VDD.n3601 VDD.n3600 55.4672
R13209 VDD.n3602 VDD.n3598 55.4672
R13210 VDD.n3859 VDD.n3858 55.4672
R13211 VDD.n3860 VDD.n3856 55.4672
R13212 VDD.n4117 VDD.n4116 55.4672
R13213 VDD.n4118 VDD.n4114 55.4672
R13214 VDD.n4375 VDD.n4374 55.4672
R13215 VDD.n4376 VDD.n4372 55.4672
R13216 VDD.n4633 VDD.n4632 55.4672
R13217 VDD.n4634 VDD.n4630 55.4672
R13218 VDD.n4891 VDD.n4890 55.4672
R13219 VDD.n4892 VDD.n4888 55.4672
R13220 VDD.n5149 VDD.n5148 55.4672
R13221 VDD.n5150 VDD.n5146 55.4672
R13222 VDD.n1803 VDD 54.4858
R13223 VDD.n2011 VDD 54.4858
R13224 VDD.n2382 VDD 54.4858
R13225 VDD.n2640 VDD 54.4858
R13226 VDD.n2898 VDD 54.4858
R13227 VDD.n3156 VDD 54.4858
R13228 VDD.n3414 VDD 54.4858
R13229 VDD.n5737 VDD 54.4858
R13230 VDD.n5483 VDD 54.4858
R13231 VDD.n3672 VDD 54.4858
R13232 VDD.n3930 VDD 54.4858
R13233 VDD.n4188 VDD 54.4858
R13234 VDD.n4446 VDD 54.4858
R13235 VDD.n4704 VDD 54.4858
R13236 VDD.n4962 VDD 54.4858
R13237 VDD.n5220 VDD 54.4858
R13238 VDD.t1026 VDD.n1927 54.472
R13239 VDD.t1038 VDD.n1927 54.472
R13240 VDD.n184 VDD.t738 54.2862
R13241 VDD.n1953 VDD.t1036 54.2478
R13242 VDD.n1949 VDD.n1941 54.1098
R13243 VDD.n1969 VDD.n1931 54.1091
R13244 VDD.t1341 VDD.t1441 52.6159
R13245 VDD.t347 VDD.t257 52.6159
R13246 VDD.t823 VDD.t539 52.6159
R13247 VDD.t788 VDD.t1013 52.6159
R13248 VDD.n183 VDD.t670 50.8934
R13249 VDD.t1026 VDD.n1939 50.8854
R13250 VDD.t967 VDD.t470 50.6439
R13251 VDD.t649 VDD.t290 50.6439
R13252 VDD.n1876 VDD.n1818 50.1034
R13253 VDD.n2197 VDD.n2139 50.1034
R13254 VDD.n2455 VDD.n2397 50.1034
R13255 VDD.n2713 VDD.n2655 50.1034
R13256 VDD.n2971 VDD.n2913 50.1034
R13257 VDD.n3229 VDD.n3171 50.1034
R13258 VDD.n3487 VDD.n3429 50.1034
R13259 VDD.n5807 VDD.n5749 50.1034
R13260 VDD.n5553 VDD.n5495 50.1034
R13261 VDD.n3745 VDD.n3687 50.1034
R13262 VDD.n4003 VDD.n3945 50.1034
R13263 VDD.n4261 VDD.n4203 50.1034
R13264 VDD.n4519 VDD.n4461 50.1034
R13265 VDD.n4777 VDD.n4719 50.1034
R13266 VDD.n5035 VDD.n4977 50.1034
R13267 VDD.n5293 VDD.n5235 50.1034
R13268 VDD.t1146 VDD.n1456 49.4526
R13269 VDD.t1242 VDD.t1172 49.2598
R13270 VDD.t1172 VDD.t1204 49.2598
R13271 VDD.t1204 VDD.t1232 49.2598
R13272 VDD.t1232 VDD.t1154 49.2598
R13273 VDD.t1154 VDD.t1190 49.2598
R13274 VDD.t1190 VDD.t1126 49.2598
R13275 VDD.t1126 VDD.t1158 49.2598
R13276 VDD.t1158 VDD.t1124 49.2598
R13277 VDD.t1124 VDD.t1184 49.2598
R13278 VDD.t1184 VDD.t1216 49.2598
R13279 VDD.t443 VDD.n1801 49.1183
R13280 VDD.t77 VDD.n2009 49.1183
R13281 VDD.t1444 VDD.n2380 49.1183
R13282 VDD.t569 VDD.n2638 49.1183
R13283 VDD.t976 VDD.n2896 49.1183
R13284 VDD.t543 VDD.n3154 49.1183
R13285 VDD.t580 VDD.n3412 49.1183
R13286 VDD.t1466 VDD.n5735 49.1183
R13287 VDD.t997 VDD.n5481 49.1183
R13288 VDD.t1333 VDD.n3670 49.1183
R13289 VDD.t483 VDD.n3928 49.1183
R13290 VDD.t7 VDD.n4186 49.1183
R13291 VDD.t1050 VDD.n4444 49.1183
R13292 VDD.t19 VDD.n4702 49.1183
R13293 VDD.t560 VDD.n4960 49.1183
R13294 VDD.t1006 VDD.n5218 49.1183
R13295 VDD.t1216 VDD.t1142 47.9846
R13296 VDD.n585 VDD.t185 47.5005
R13297 VDD.n935 VDD.t958 47.5005
R13298 VDD.n1700 VDD.n1681 47.0405
R13299 VDD.n2049 VDD.n2030 47.0405
R13300 VDD.n2279 VDD.n2260 47.0405
R13301 VDD.n2537 VDD.n2518 47.0405
R13302 VDD.n2795 VDD.n2776 47.0405
R13303 VDD.n3053 VDD.n3034 47.0405
R13304 VDD.n3311 VDD.n3292 47.0405
R13305 VDD.n5634 VDD.n5615 47.0405
R13306 VDD.n5380 VDD.n5361 47.0405
R13307 VDD.n3569 VDD.n3550 47.0405
R13308 VDD.n3827 VDD.n3808 47.0405
R13309 VDD.n4085 VDD.n4066 47.0405
R13310 VDD.n4343 VDD.n4324 47.0405
R13311 VDD.n4601 VDD.n4582 47.0405
R13312 VDD.n4859 VDD.n4840 47.0405
R13313 VDD.n5117 VDD.n5098 47.0405
R13314 VDD.n1966 VDD.n1936 46.6829
R13315 VDD.n1973 VDD.n1972 45.9299
R13316 VDD.n1959 VDD.n1958 45.9299
R13317 VDD.n1705 VDD.n1704 45.7605
R13318 VDD.n1689 VDD.n1685 45.7605
R13319 VDD.n2054 VDD.n2053 45.7605
R13320 VDD.n2038 VDD.n2034 45.7605
R13321 VDD.n2284 VDD.n2283 45.7605
R13322 VDD.n2268 VDD.n2264 45.7605
R13323 VDD.n2542 VDD.n2541 45.7605
R13324 VDD.n2526 VDD.n2522 45.7605
R13325 VDD.n2800 VDD.n2799 45.7605
R13326 VDD.n2784 VDD.n2780 45.7605
R13327 VDD.n3058 VDD.n3057 45.7605
R13328 VDD.n3042 VDD.n3038 45.7605
R13329 VDD.n3316 VDD.n3315 45.7605
R13330 VDD.n3300 VDD.n3296 45.7605
R13331 VDD.n5639 VDD.n5638 45.7605
R13332 VDD.n5623 VDD.n5619 45.7605
R13333 VDD.n5385 VDD.n5384 45.7605
R13334 VDD.n5369 VDD.n5365 45.7605
R13335 VDD.n3574 VDD.n3573 45.7605
R13336 VDD.n3558 VDD.n3554 45.7605
R13337 VDD.n3832 VDD.n3831 45.7605
R13338 VDD.n3816 VDD.n3812 45.7605
R13339 VDD.n4090 VDD.n4089 45.7605
R13340 VDD.n4074 VDD.n4070 45.7605
R13341 VDD.n4348 VDD.n4347 45.7605
R13342 VDD.n4332 VDD.n4328 45.7605
R13343 VDD.n4606 VDD.n4605 45.7605
R13344 VDD.n4590 VDD.n4586 45.7605
R13345 VDD.n4864 VDD.n4863 45.7605
R13346 VDD.n4848 VDD.n4844 45.7605
R13347 VDD.n5122 VDD.n5121 45.7605
R13348 VDD.n5106 VDD.n5102 45.7605
R13349 VDD.n1684 VDD.n1682 45.4405
R13350 VDD.n2033 VDD.n2031 45.4405
R13351 VDD.n2263 VDD.n2261 45.4405
R13352 VDD.n2521 VDD.n2519 45.4405
R13353 VDD.n2779 VDD.n2777 45.4405
R13354 VDD.n3037 VDD.n3035 45.4405
R13355 VDD.n3295 VDD.n3293 45.4405
R13356 VDD.n5618 VDD.n5616 45.4405
R13357 VDD.n5364 VDD.n5362 45.4405
R13358 VDD.n3553 VDD.n3551 45.4405
R13359 VDD.n3811 VDD.n3809 45.4405
R13360 VDD.n4069 VDD.n4067 45.4405
R13361 VDD.n4327 VDD.n4325 45.4405
R13362 VDD.n4585 VDD.n4583 45.4405
R13363 VDD.n4843 VDD.n4841 45.4405
R13364 VDD.n5101 VDD.n5099 45.4405
R13365 VDD.n1947 VDD.n1937 44.8005
R13366 VDD.n408 VDD 43.6586
R13367 VDD.n1566 VDD 43.6586
R13368 VDD.n1 VDD.t975 42.3555
R13369 VDD.n468 VDD.t638 42.3555
R13370 VDD.n439 VDD.t554 42.3555
R13371 VDD.n459 VDD.t461 42.3555
R13372 VDD.n66 VDD.t432 42.3555
R13373 VDD.n36 VDD.t18 42.3555
R13374 VDD.n56 VDD.t636 42.3555
R13375 VDD.n1145 VDD.t382 42.3555
R13376 VDD.n1947 VDD.n1946 41.323
R13377 VDD.n1936 VDD.n1933 41.2617
R13378 VDD.n1708 VDD.n1707 39.5299
R13379 VDD.n1761 VDD.n1760 39.5299
R13380 VDD.n2057 VDD.n2056 39.5299
R13381 VDD.n2110 VDD.n2109 39.5299
R13382 VDD.n2287 VDD.n2286 39.5299
R13383 VDD.n2340 VDD.n2339 39.5299
R13384 VDD.n2545 VDD.n2544 39.5299
R13385 VDD.n2598 VDD.n2597 39.5299
R13386 VDD.n2803 VDD.n2802 39.5299
R13387 VDD.n2856 VDD.n2855 39.5299
R13388 VDD.n3061 VDD.n3060 39.5299
R13389 VDD.n3114 VDD.n3113 39.5299
R13390 VDD.n3319 VDD.n3318 39.5299
R13391 VDD.n3372 VDD.n3371 39.5299
R13392 VDD.n5642 VDD.n5641 39.5299
R13393 VDD.n5695 VDD.n5694 39.5299
R13394 VDD.n5388 VDD.n5387 39.5299
R13395 VDD.n5441 VDD.n5440 39.5299
R13396 VDD.n3577 VDD.n3576 39.5299
R13397 VDD.n3630 VDD.n3629 39.5299
R13398 VDD.n3835 VDD.n3834 39.5299
R13399 VDD.n3888 VDD.n3887 39.5299
R13400 VDD.n4093 VDD.n4092 39.5299
R13401 VDD.n4146 VDD.n4145 39.5299
R13402 VDD.n4351 VDD.n4350 39.5299
R13403 VDD.n4404 VDD.n4403 39.5299
R13404 VDD.n4609 VDD.n4608 39.5299
R13405 VDD.n4662 VDD.n4661 39.5299
R13406 VDD.n4867 VDD.n4866 39.5299
R13407 VDD.n4920 VDD.n4919 39.5299
R13408 VDD.n5125 VDD.n5124 39.5299
R13409 VDD.n5178 VDD.n5177 39.5299
R13410 VDD.n20 VDD.n3 39.2858
R13411 VDD.n1164 VDD.n1147 39.2858
R13412 VDD VDD.t75 39.0862
R13413 VDD VDD.t285 39.0862
R13414 VDD.n1885 VDD.n1884 38.9491
R13415 VDD.n2206 VDD.n2205 38.9491
R13416 VDD.n2464 VDD.n2463 38.9491
R13417 VDD.n2722 VDD.n2721 38.9491
R13418 VDD.n2980 VDD.n2979 38.9491
R13419 VDD.n3238 VDD.n3237 38.9491
R13420 VDD.n3496 VDD.n3495 38.9491
R13421 VDD.n5816 VDD.n5815 38.9491
R13422 VDD.n5562 VDD.n5561 38.9491
R13423 VDD.n3754 VDD.n3753 38.9491
R13424 VDD.n4012 VDD.n4011 38.9491
R13425 VDD.n4270 VDD.n4269 38.9491
R13426 VDD.n4528 VDD.n4527 38.9491
R13427 VDD.n4786 VDD.n4785 38.9491
R13428 VDD.n5044 VDD.n5043 38.9491
R13429 VDD.n5302 VDD.n5301 38.9491
R13430 VDD.t71 VDD.t345 38.8641
R13431 VDD.t629 VDD.t785 38.8641
R13432 VDD.t449 VDD.t1122 38.534
R13433 VDD.t565 VDD.t1457 38.534
R13434 VDD.n1746 VDD.n1745 37.3765
R13435 VDD.n1728 VDD.n1725 37.3765
R13436 VDD.n2095 VDD.n2094 37.3765
R13437 VDD.n2077 VDD.n2074 37.3765
R13438 VDD.n2325 VDD.n2324 37.3765
R13439 VDD.n2307 VDD.n2304 37.3765
R13440 VDD.n2583 VDD.n2582 37.3765
R13441 VDD.n2565 VDD.n2562 37.3765
R13442 VDD.n2841 VDD.n2840 37.3765
R13443 VDD.n2823 VDD.n2820 37.3765
R13444 VDD.n3099 VDD.n3098 37.3765
R13445 VDD.n3081 VDD.n3078 37.3765
R13446 VDD.n3357 VDD.n3356 37.3765
R13447 VDD.n3339 VDD.n3336 37.3765
R13448 VDD.n5680 VDD.n5679 37.3765
R13449 VDD.n5662 VDD.n5659 37.3765
R13450 VDD.n5426 VDD.n5425 37.3765
R13451 VDD.n5408 VDD.n5405 37.3765
R13452 VDD.n3615 VDD.n3614 37.3765
R13453 VDD.n3597 VDD.n3594 37.3765
R13454 VDD.n3873 VDD.n3872 37.3765
R13455 VDD.n3855 VDD.n3852 37.3765
R13456 VDD.n4131 VDD.n4130 37.3765
R13457 VDD.n4113 VDD.n4110 37.3765
R13458 VDD.n4389 VDD.n4388 37.3765
R13459 VDD.n4371 VDD.n4368 37.3765
R13460 VDD.n4647 VDD.n4646 37.3765
R13461 VDD.n4629 VDD.n4626 37.3765
R13462 VDD.n4905 VDD.n4904 37.3765
R13463 VDD.n4887 VDD.n4884 37.3765
R13464 VDD.n5163 VDD.n5162 37.3765
R13465 VDD.n5145 VDD.n5142 37.3765
R13466 VDD.n1830 VDD.t1089 36.1587
R13467 VDD.n1830 VDD.t600 36.1587
R13468 VDD.n1813 VDD.t1499 36.1587
R13469 VDD.n1813 VDD.t465 36.1587
R13470 VDD.n2134 VDD.t626 36.1587
R13471 VDD.n2134 VDD.t256 36.1587
R13472 VDD.n2151 VDD.t556 36.1587
R13473 VDD.n2151 VDD.t1012 36.1587
R13474 VDD.n2392 VDD.t1285 36.1587
R13475 VDD.n2392 VDD.t1018 36.1587
R13476 VDD.n2409 VDD.t1384 36.1587
R13477 VDD.n2409 VDD.t616 36.1587
R13478 VDD.n2650 VDD.t86 36.1587
R13479 VDD.n2650 VDD.t1324 36.1587
R13480 VDD.n2667 VDD.t576 36.1587
R13481 VDD.n2667 VDD.t248 36.1587
R13482 VDD.n2908 VDD.t273 36.1587
R13483 VDD.n2908 VDD.t367 36.1587
R13484 VDD.n2925 VDD.t1480 36.1587
R13485 VDD.n2925 VDD.t619 36.1587
R13486 VDD.n3166 VDD.t542 36.1587
R13487 VDD.n3166 VDD.t1460 36.1587
R13488 VDD.n3183 VDD.t1004 36.1587
R13489 VDD.n3183 VDD.t648 36.1587
R13490 VDD.n3424 VDD.t1281 36.1587
R13491 VDD.n3424 VDD.t1294 36.1587
R13492 VDD.n3441 VDD.t398 36.1587
R13493 VDD.n3441 VDD.t533 36.1587
R13494 VDD.n5744 VDD.t520 36.1587
R13495 VDD.n5744 VDD.t602 36.1587
R13496 VDD.n5761 VDD.t68 36.1587
R13497 VDD.n5761 VDD.t1354 36.1587
R13498 VDD.n5490 VDD.t454 36.1587
R13499 VDD.n5490 VDD.t644 36.1587
R13500 VDD.n5507 VDD.t1306 36.1587
R13501 VDD.n5507 VDD.t392 36.1587
R13502 VDD.n3682 VDD.t1102 36.1587
R13503 VDD.n3682 VDD.t254 36.1587
R13504 VDD.n3699 VDD.t1071 36.1587
R13505 VDD.n3699 VDD.t292 36.1587
R13506 VDD.n3940 VDD.t1049 36.1587
R13507 VDD.n3940 VDD.t269 36.1587
R13508 VDD.n3957 VDD.t1063 36.1587
R13509 VDD.n3957 VDD.t1349 36.1587
R13510 VDD.n4198 VDD.t1463 36.1587
R13511 VDD.n4198 VDD.t16 36.1587
R13512 VDD.n4215 VDD.t985 36.1587
R13513 VDD.n4215 VDD.t1364 36.1587
R13514 VDD.n4456 VDD.t1106 36.1587
R13515 VDD.n4456 VDD.t1068 36.1587
R13516 VDD.n4473 VDD.t459 36.1587
R13517 VDD.n4473 VDD.t609 36.1587
R13518 VDD.n4714 VDD.t1501 36.1587
R13519 VDD.n4714 VDD.t1310 36.1587
R13520 VDD.n4731 VDD.t1475 36.1587
R13521 VDD.n4731 VDD.t400 36.1587
R13522 VDD.n4972 VDD.t1289 36.1587
R13523 VDD.n4972 VDD.t818 36.1587
R13524 VDD.n4989 VDD.t1043 36.1587
R13525 VDD.n4989 VDD.t1100 36.1587
R13526 VDD.n5230 VDD.t482 36.1587
R13527 VDD.n5230 VDD.t1059 36.1587
R13528 VDD.n5247 VDD.t634 36.1587
R13529 VDD.n5247 VDD.t406 36.1587
R13530 VDD.t1346 VDD.t1321 35.0774
R13531 VDD.t500 VDD.t1303 35.0774
R13532 VDD VDD.n1802 34.927
R13533 VDD VDD.n2010 34.927
R13534 VDD VDD.n2381 34.927
R13535 VDD VDD.n2639 34.927
R13536 VDD VDD.n2897 34.927
R13537 VDD VDD.n3155 34.927
R13538 VDD VDD.n3413 34.927
R13539 VDD VDD.n5736 34.927
R13540 VDD VDD.n5482 34.927
R13541 VDD VDD.n3671 34.927
R13542 VDD VDD.n3929 34.927
R13543 VDD VDD.n4187 34.927
R13544 VDD VDD.n4445 34.927
R13545 VDD VDD.n4703 34.927
R13546 VDD VDD.n4961 34.927
R13547 VDD VDD.n5219 34.927
R13548 VDD.n23 VDD.n2 34.6358
R13549 VDD.n18 VDD.n6 34.6358
R13550 VDD.n679 VDD.n678 34.6358
R13551 VDD.n500 VDD.n499 34.6358
R13552 VDD.n427 VDD.n426 34.6358
R13553 VDD.n98 VDD.n97 34.6358
R13554 VDD.n1167 VDD.n1146 34.6358
R13555 VDD.n1162 VDD.n1150 34.6358
R13556 VDD.n1585 VDD.n1584 34.6358
R13557 VDD.n832 VDD.n831 34.6358
R13558 VDD.n844 VDD.n843 34.6358
R13559 VDD.n850 VDD.n849 34.6358
R13560 VDD.n813 VDD.n801 34.6358
R13561 VDD.n817 VDD.n801 34.6358
R13562 VDD.n818 VDD.n817 34.6358
R13563 VDD.n811 VDD.n804 34.6358
R13564 VDD.n1029 VDD.n1028 34.6358
R13565 VDD.n274 VDD.n273 34.6358
R13566 VDD.n1215 VDD.n1214 34.6358
R13567 VDD.n1227 VDD.n1226 34.6358
R13568 VDD.n1233 VDD.n1232 34.6358
R13569 VDD.n1196 VDD.n1184 34.6358
R13570 VDD.n1200 VDD.n1184 34.6358
R13571 VDD.n1201 VDD.n1200 34.6358
R13572 VDD.n1194 VDD.n1187 34.6358
R13573 VDD.n667 VDD.t111 33.9291
R13574 VDD.n1017 VDD.t884 33.9291
R13575 VDD.n838 VDD.n837 33.8829
R13576 VDD.n1221 VDD.n1220 33.8829
R13577 VDD.n1958 VDD.n1957 33.8422
R13578 VDD.n1397 VDD.t300 33.8361
R13579 VDD.n1973 VDD.n1923 33.6292
R13580 VDD.t455 VDD.t69 32.6058
R13581 VDD.t462 VDD.t627 32.6058
R13582 VDD.t73 VDD.t553 31.4862
R13583 VDD.t75 VDD.t460 31.4862
R13584 VDD.t426 VDD.t17 31.4862
R13585 VDD.t285 VDD.t635 31.4862
R13586 VDD.n1914 VDD.t277 30.1961
R13587 VDD.n2235 VDD.t494 30.1961
R13588 VDD.n2493 VDD.t505 30.1961
R13589 VDD.n2751 VDD.t1023 30.1961
R13590 VDD.n3009 VDD.t524 30.1961
R13591 VDD.n3267 VDD.t282 30.1961
R13592 VDD.n3525 VDD.t419 30.1961
R13593 VDD.n5845 VDD.t1075 30.1961
R13594 VDD.n5591 VDD.t393 30.1961
R13595 VDD.n3783 VDD.t262 30.1961
R13596 VDD.n4041 VDD.t1084 30.1961
R13597 VDD.n4299 VDD.t1021 30.1961
R13598 VDD.n4557 VDD.t531 30.1961
R13599 VDD.n4815 VDD.t401 30.1961
R13600 VDD.n5073 VDD.t416 30.1961
R13601 VDD.n5331 VDD.t407 30.1961
R13602 VDD.n542 VDD.n541 29.3652
R13603 VDD.n621 VDD.n620 29.3652
R13604 VDD.n517 VDD.n516 29.3652
R13605 VDD.n520 VDD.n519 29.3652
R13606 VDD.n892 VDD.n891 29.3652
R13607 VDD.n971 VDD.n970 29.3652
R13608 VDD.n867 VDD.n866 29.3652
R13609 VDD.n870 VDD.n869 29.3652
R13610 VDD.n141 VDD.n140 29.3652
R13611 VDD.n220 VDD.n219 29.3652
R13612 VDD.n116 VDD.n115 29.3652
R13613 VDD.n119 VDD.n118 29.3652
R13614 VDD.n1313 VDD.n1312 29.3652
R13615 VDD.n1342 VDD.n1341 29.3652
R13616 VDD.n523 VDD.n522 28.9887
R13617 VDD.n873 VDD.n872 28.9887
R13618 VDD.n122 VDD.n121 28.9887
R13619 VDD.n1348 VDD.n1347 28.9887
R13620 VDD.n5 VDD.t450 28.4628
R13621 VDD.n494 VDD.t336 28.4628
R13622 VDD.n422 VDD.t365 28.4628
R13623 VDD.n418 VDD.t973 28.4628
R13624 VDD.n401 VDD.t1442 28.4628
R13625 VDD.n92 VDD.t503 28.4628
R13626 VDD.n1149 VDD.t566 28.4628
R13627 VDD.n1580 VDD.t1120 28.4628
R13628 VDD.n1576 VDD.t650 28.4628
R13629 VDD.n1559 VDD.t540 28.4628
R13630 VDD.n806 VDD.t552 28.4628
R13631 VDD.n1189 VDD.t607 28.4628
R13632 VDD.n1793 VDD.n1782 28.2358
R13633 VDD.n1794 VDD.n1793 28.2358
R13634 VDD.n1790 VDD.n1787 28.2358
R13635 VDD.n1790 VDD.n1789 28.2358
R13636 VDD.n2001 VDD.n1990 28.2358
R13637 VDD.n2002 VDD.n2001 28.2358
R13638 VDD.n1998 VDD.n1995 28.2358
R13639 VDD.n1998 VDD.n1997 28.2358
R13640 VDD.n2372 VDD.n2361 28.2358
R13641 VDD.n2373 VDD.n2372 28.2358
R13642 VDD.n2369 VDD.n2366 28.2358
R13643 VDD.n2369 VDD.n2368 28.2358
R13644 VDD.n2630 VDD.n2619 28.2358
R13645 VDD.n2631 VDD.n2630 28.2358
R13646 VDD.n2627 VDD.n2624 28.2358
R13647 VDD.n2627 VDD.n2626 28.2358
R13648 VDD.n2888 VDD.n2877 28.2358
R13649 VDD.n2889 VDD.n2888 28.2358
R13650 VDD.n2885 VDD.n2882 28.2358
R13651 VDD.n2885 VDD.n2884 28.2358
R13652 VDD.n3146 VDD.n3135 28.2358
R13653 VDD.n3147 VDD.n3146 28.2358
R13654 VDD.n3143 VDD.n3140 28.2358
R13655 VDD.n3143 VDD.n3142 28.2358
R13656 VDD.n3404 VDD.n3393 28.2358
R13657 VDD.n3405 VDD.n3404 28.2358
R13658 VDD.n3401 VDD.n3398 28.2358
R13659 VDD.n3401 VDD.n3400 28.2358
R13660 VDD.n5727 VDD.n5716 28.2358
R13661 VDD.n5728 VDD.n5727 28.2358
R13662 VDD.n5724 VDD.n5721 28.2358
R13663 VDD.n5724 VDD.n5723 28.2358
R13664 VDD.n5473 VDD.n5462 28.2358
R13665 VDD.n5474 VDD.n5473 28.2358
R13666 VDD.n5470 VDD.n5467 28.2358
R13667 VDD.n5470 VDD.n5469 28.2358
R13668 VDD.n3662 VDD.n3651 28.2358
R13669 VDD.n3663 VDD.n3662 28.2358
R13670 VDD.n3659 VDD.n3656 28.2358
R13671 VDD.n3659 VDD.n3658 28.2358
R13672 VDD.n3920 VDD.n3909 28.2358
R13673 VDD.n3921 VDD.n3920 28.2358
R13674 VDD.n3917 VDD.n3914 28.2358
R13675 VDD.n3917 VDD.n3916 28.2358
R13676 VDD.n4178 VDD.n4167 28.2358
R13677 VDD.n4179 VDD.n4178 28.2358
R13678 VDD.n4175 VDD.n4172 28.2358
R13679 VDD.n4175 VDD.n4174 28.2358
R13680 VDD.n4436 VDD.n4425 28.2358
R13681 VDD.n4437 VDD.n4436 28.2358
R13682 VDD.n4433 VDD.n4430 28.2358
R13683 VDD.n4433 VDD.n4432 28.2358
R13684 VDD.n4694 VDD.n4683 28.2358
R13685 VDD.n4695 VDD.n4694 28.2358
R13686 VDD.n4691 VDD.n4688 28.2358
R13687 VDD.n4691 VDD.n4690 28.2358
R13688 VDD.n4952 VDD.n4941 28.2358
R13689 VDD.n4953 VDD.n4952 28.2358
R13690 VDD.n4949 VDD.n4946 28.2358
R13691 VDD.n4949 VDD.n4948 28.2358
R13692 VDD.n5210 VDD.n5199 28.2358
R13693 VDD.n5211 VDD.n5210 28.2358
R13694 VDD.n5207 VDD.n5204 28.2358
R13695 VDD.n5207 VDD.n5206 28.2358
R13696 VDD.n13 VDD.n8 28.2358
R13697 VDD.n1157 VDD.n1152 28.2358
R13698 VDD.n463 VDD 28.2291
R13699 VDD.n60 VDD 28.2291
R13700 VDD.n262 VDD.t664 27.1434
R13701 VDD.n482 VDD.t1104 26.9729
R13702 VDD.n80 VDD.t1453 26.9729
R13703 VDD.n1835 VDD.n1834 26.8623
R13704 VDD.n2156 VDD.n2155 26.8623
R13705 VDD.n2414 VDD.n2413 26.8623
R13706 VDD.n2672 VDD.n2671 26.8623
R13707 VDD.n2930 VDD.n2929 26.8623
R13708 VDD.n3188 VDD.n3187 26.8623
R13709 VDD.n3446 VDD.n3445 26.8623
R13710 VDD.n5766 VDD.n5765 26.8623
R13711 VDD.n5512 VDD.n5511 26.8623
R13712 VDD.n3704 VDD.n3703 26.8623
R13713 VDD.n3962 VDD.n3961 26.8623
R13714 VDD.n4220 VDD.n4219 26.8623
R13715 VDD.n4478 VDD.n4477 26.8623
R13716 VDD.n4736 VDD.n4735 26.8623
R13717 VDD.n4994 VDD.n4993 26.8623
R13718 VDD.n5252 VDD.n5251 26.8623
R13719 VDD.n1656 VDD 26.615
R13720 VDD.n31 VDD.t1455 26.5955
R13721 VDD.n508 VDD.t412 26.5955
R13722 VDD.n435 VDD.t968 26.5955
R13723 VDD.n404 VDD.t612 26.5955
R13724 VDD.n106 VDD.t430 26.5955
R13725 VDD.n1175 VDD.t499 26.5955
R13726 VDD.n1593 VDD.t1287 26.5955
R13727 VDD.n1562 VDD.t1492 26.5955
R13728 VDD.n800 VDD.t589 26.5955
R13729 VDD.n803 VDD.t622 26.5955
R13730 VDD.n1183 VDD.t404 26.5955
R13731 VDD.n1186 VDD.t579 26.5955
R13732 VDD.n1792 VDD.t447 26.5955
R13733 VDD.n1792 VDD.t444 26.5955
R13734 VDD.n1788 VDD.t1030 26.5955
R13735 VDD.n1788 VDD.t1034 26.5955
R13736 VDD.n2000 VDD.t79 26.5955
R13737 VDD.n2000 VDD.t83 26.5955
R13738 VDD.n1996 VDD.t1270 26.5955
R13739 VDD.n1996 VDD.t1267 26.5955
R13740 VDD.n2371 VDD.t1448 26.5955
R13741 VDD.n2371 VDD.t1450 26.5955
R13742 VDD.n2367 VDD.t834 26.5955
R13743 VDD.n2367 VDD.t829 26.5955
R13744 VDD.n2629 VDD.t571 26.5955
R13745 VDD.n2629 VDD.t572 26.5955
R13746 VDD.n2625 VDD.t1421 26.5955
R13747 VDD.n2625 VDD.t1423 26.5955
R13748 VDD.n2887 VDD.t980 26.5955
R13749 VDD.n2887 VDD.t982 26.5955
R13750 VDD.n2883 VDD.t435 26.5955
R13751 VDD.n2883 VDD.t438 26.5955
R13752 VDD.n3145 VDD.t547 26.5955
R13753 VDD.n3145 VDD.t549 26.5955
R13754 VDD.n3141 VDD.t390 26.5955
R13755 VDD.n3141 VDD.t386 26.5955
R13756 VDD.n3403 VDD.t584 26.5955
R13757 VDD.n3403 VDD.t586 26.5955
R13758 VDD.n3399 VDD.t1299 26.5955
R13759 VDD.n3399 VDD.t1301 26.5955
R13760 VDD.n5726 VDD.t1470 26.5955
R13761 VDD.n5726 VDD.t1472 26.5955
R13762 VDD.n5722 VDD.t475 26.5955
R13763 VDD.n5722 VDD.t478 26.5955
R13764 VDD.n5472 VDD.t1002 26.5955
R13765 VDD.n5472 VDD.t998 26.5955
R13766 VDD.n5468 VDD.t1261 26.5955
R13767 VDD.n5468 VDD.t1263 26.5955
R13768 VDD.n3661 VDD.t1338 26.5955
R13769 VDD.n3661 VDD.t1340 26.5955
R13770 VDD.n3657 VDD.t1370 26.5955
R13771 VDD.n3657 VDD.t1372 26.5955
R13772 VDD.n3919 VDD.t484 26.5955
R13773 VDD.n3919 VDD.t487 26.5955
R13774 VDD.n3915 VDD.t1117 26.5955
R13775 VDD.n3915 VDD.t1112 26.5955
R13776 VDD.n4177 VDD.t12 26.5955
R13777 VDD.n4177 VDD.t8 26.5955
R13778 VDD.n4173 VDD.t33 26.5955
R13779 VDD.n4173 VDD.t28 26.5955
R13780 VDD.n4435 VDD.t1054 26.5955
R13781 VDD.n4435 VDD.t1056 26.5955
R13782 VDD.n4431 VDD.t1435 26.5955
R13783 VDD.n4431 VDD.t1438 26.5955
R13784 VDD.n4693 VDD.t23 26.5955
R13785 VDD.n4693 VDD.t25 26.5955
R13786 VDD.n4689 VDD.t377 26.5955
R13787 VDD.n4689 VDD.t373 26.5955
R13788 VDD.n4951 VDD.t820 26.5955
R13789 VDD.n4951 VDD.t562 26.5955
R13790 VDD.n4947 VDD.t1040 26.5955
R13791 VDD.n4947 VDD.t421 26.5955
R13792 VDD.n5209 VDD.t1326 26.5955
R13793 VDD.n5209 VDD.t1007 26.5955
R13794 VDD.n5205 VDD.t1253 26.5955
R13795 VDD.n5205 VDD.t4 26.5955
R13796 VDD.n692 VDD.t342 26.5955
R13797 VDD.n692 VDD.t344 26.5955
R13798 VDD.n555 VDD.t208 26.5955
R13799 VDD.n555 VDD.t140 26.5955
R13800 VDD.n561 VDD.t114 26.5955
R13801 VDD.n561 VDD.t178 26.5955
R13802 VDD.n567 VDD.t194 26.5955
R13803 VDD.n567 VDD.t90 26.5955
R13804 VDD.n573 VDD.t88 26.5955
R13805 VDD.n573 VDD.t124 26.5955
R13806 VDD.n578 VDD.t120 26.5955
R13807 VDD.n578 VDD.t146 26.5955
R13808 VDD.n534 VDD.t106 26.5955
R13809 VDD.n534 VDD.t98 26.5955
R13810 VDD.n529 VDD.t128 26.5955
R13811 VDD.n529 VDD.t214 26.5955
R13812 VDD.n613 VDD.t212 26.5955
R13813 VDD.n613 VDD.t144 26.5955
R13814 VDD.n607 VDD.t138 26.5955
R13815 VDD.n607 VDD.t164 26.5955
R13816 VDD.n601 VDD.t126 26.5955
R13817 VDD.n601 VDD.t206 26.5955
R13818 VDD.n595 VDD.t156 26.5955
R13819 VDD.n595 VDD.t190 26.5955
R13820 VDD.n591 VDD.t186 26.5955
R13821 VDD.n591 VDD.t118 26.5955
R13822 VDD.n525 VDD.t96 26.5955
R13823 VDD.n525 VDD.t152 26.5955
R13824 VDD.n545 VDD.t172 26.5955
R13825 VDD.n545 VDD.t198 26.5955
R13826 VDD.n638 VDD.t108 26.5955
R13827 VDD.n638 VDD.t130 26.5955
R13828 VDD.n644 VDD.t136 26.5955
R13829 VDD.n644 VDD.t162 26.5955
R13830 VDD.n650 VDD.t160 26.5955
R13831 VDD.n650 VDD.t192 26.5955
R13832 VDD.n656 VDD.t204 26.5955
R13833 VDD.n656 VDD.t134 26.5955
R13834 VDD.n661 VDD.t112 26.5955
R13835 VDD.n661 VDD.t176 26.5955
R13836 VDD.n631 VDD.t116 26.5955
R13837 VDD.n631 VDD.t202 26.5955
R13838 VDD.n625 VDD.t150 26.5955
R13839 VDD.n625 VDD.t180 26.5955
R13840 VDD.n748 VDD.t142 26.5955
R13841 VDD.n748 VDD.t166 26.5955
R13842 VDD.n754 VDD.t182 26.5955
R13843 VDD.n754 VDD.t210 26.5955
R13844 VDD.n760 VDD.t158 26.5955
R13845 VDD.n760 VDD.t100 26.5955
R13846 VDD.n766 VDD.t188 26.5955
R13847 VDD.n766 VDD.t122 26.5955
R13848 VDD.n770 VDD.t132 26.5955
R13849 VDD.n770 VDD.t154 26.5955
R13850 VDD.n777 VDD.t174 26.5955
R13851 VDD.n777 VDD.t200 26.5955
R13852 VDD.n785 VDD.t196 26.5955
R13853 VDD.n785 VDD.t94 26.5955
R13854 VDD.n701 VDD.t1390 26.5955
R13855 VDD.n701 VDD.t1404 26.5955
R13856 VDD.n707 VDD.t1402 26.5955
R13857 VDD.n707 VDD.t1386 26.5955
R13858 VDD.n713 VDD.t1416 26.5955
R13859 VDD.n713 VDD.t1396 26.5955
R13860 VDD.n719 VDD.t1394 26.5955
R13861 VDD.n719 VDD.t1408 26.5955
R13862 VDD.n723 VDD.t1406 26.5955
R13863 VDD.n723 VDD.t1414 26.5955
R13864 VDD.n729 VDD.t1400 26.5955
R13865 VDD.n729 VDD.t1410 26.5955
R13866 VDD.n737 VDD.t1412 26.5955
R13867 VDD.n737 VDD.t1392 26.5955
R13868 VDD.n1042 VDD.t1083 26.5955
R13869 VDD.n1042 VDD.t1077 26.5955
R13870 VDD.n905 VDD.t853 26.5955
R13871 VDD.n905 VDD.t913 26.5955
R13872 VDD.n911 VDD.t887 26.5955
R13873 VDD.n911 VDD.t951 26.5955
R13874 VDD.n917 VDD.t839 26.5955
R13875 VDD.n917 VDD.t863 26.5955
R13876 VDD.n923 VDD.t861 26.5955
R13877 VDD.n923 VDD.t897 26.5955
R13878 VDD.n928 VDD.t891 26.5955
R13879 VDD.n928 VDD.t919 26.5955
R13880 VDD.n884 VDD.t879 26.5955
R13881 VDD.n884 VDD.t871 26.5955
R13882 VDD.n879 VDD.t901 26.5955
R13883 VDD.n879 VDD.t859 26.5955
R13884 VDD.n963 VDD.t857 26.5955
R13885 VDD.n963 VDD.t917 26.5955
R13886 VDD.n957 VDD.t911 26.5955
R13887 VDD.n957 VDD.t939 26.5955
R13888 VDD.n951 VDD.t899 26.5955
R13889 VDD.n951 VDD.t851 26.5955
R13890 VDD.n945 VDD.t929 26.5955
R13891 VDD.n945 VDD.t963 26.5955
R13892 VDD.n941 VDD.t959 26.5955
R13893 VDD.n941 VDD.t893 26.5955
R13894 VDD.n875 VDD.t869 26.5955
R13895 VDD.n875 VDD.t925 26.5955
R13896 VDD.n895 VDD.t933 26.5955
R13897 VDD.n895 VDD.t843 26.5955
R13898 VDD.n988 VDD.t881 26.5955
R13899 VDD.n988 VDD.t905 26.5955
R13900 VDD.n994 VDD.t909 26.5955
R13901 VDD.n994 VDD.t937 26.5955
R13902 VDD.n1000 VDD.t935 26.5955
R13903 VDD.n1000 VDD.t965 26.5955
R13904 VDD.n1006 VDD.t849 26.5955
R13905 VDD.n1006 VDD.t903 26.5955
R13906 VDD.n1011 VDD.t885 26.5955
R13907 VDD.n1011 VDD.t949 26.5955
R13908 VDD.n981 VDD.t889 26.5955
R13909 VDD.n981 VDD.t847 26.5955
R13910 VDD.n975 VDD.t923 26.5955
R13911 VDD.n975 VDD.t953 26.5955
R13912 VDD.n1098 VDD.t915 26.5955
R13913 VDD.n1098 VDD.t941 26.5955
R13914 VDD.n1104 VDD.t955 26.5955
R13915 VDD.n1104 VDD.t855 26.5955
R13916 VDD.n1110 VDD.t931 26.5955
R13917 VDD.n1110 VDD.t873 26.5955
R13918 VDD.n1116 VDD.t961 26.5955
R13919 VDD.n1116 VDD.t895 26.5955
R13920 VDD.n1120 VDD.t907 26.5955
R13921 VDD.n1120 VDD.t927 26.5955
R13922 VDD.n1127 VDD.t947 26.5955
R13923 VDD.n1127 VDD.t845 26.5955
R13924 VDD.n1135 VDD.t841 26.5955
R13925 VDD.n1135 VDD.t867 26.5955
R13926 VDD.n1051 VDD.t46 26.5955
R13927 VDD.n1051 VDD.t60 26.5955
R13928 VDD.n1057 VDD.t58 26.5955
R13929 VDD.n1057 VDD.t42 26.5955
R13930 VDD.n1063 VDD.t40 26.5955
R13931 VDD.n1063 VDD.t52 26.5955
R13932 VDD.n1069 VDD.t50 26.5955
R13933 VDD.n1069 VDD.t64 26.5955
R13934 VDD.n1073 VDD.t62 26.5955
R13935 VDD.n1073 VDD.t38 26.5955
R13936 VDD.n1079 VDD.t56 26.5955
R13937 VDD.n1079 VDD.t66 26.5955
R13938 VDD.n1087 VDD.t36 26.5955
R13939 VDD.n1087 VDD.t48 26.5955
R13940 VDD.n287 VDD.t989 26.5955
R13941 VDD.n287 VDD.t991 26.5955
R13942 VDD.n154 VDD.t761 26.5955
R13943 VDD.n154 VDD.t693 26.5955
R13944 VDD.n160 VDD.t667 26.5955
R13945 VDD.n160 VDD.t731 26.5955
R13946 VDD.n166 VDD.t747 26.5955
R13947 VDD.n166 VDD.t771 26.5955
R13948 VDD.n172 VDD.t769 26.5955
R13949 VDD.n172 VDD.t679 26.5955
R13950 VDD.n177 VDD.t671 26.5955
R13951 VDD.n177 VDD.t699 26.5955
R13952 VDD.n133 VDD.t659 26.5955
R13953 VDD.n133 VDD.t779 26.5955
R13954 VDD.n128 VDD.t681 26.5955
R13955 VDD.n128 VDD.t767 26.5955
R13956 VDD.n212 VDD.t765 26.5955
R13957 VDD.n212 VDD.t697 26.5955
R13958 VDD.n206 VDD.t691 26.5955
R13959 VDD.n206 VDD.t717 26.5955
R13960 VDD.n200 VDD.t677 26.5955
R13961 VDD.n200 VDD.t759 26.5955
R13962 VDD.n194 VDD.t709 26.5955
R13963 VDD.n194 VDD.t743 26.5955
R13964 VDD.n190 VDD.t739 26.5955
R13965 VDD.n190 VDD.t673 26.5955
R13966 VDD.n124 VDD.t777 26.5955
R13967 VDD.n124 VDD.t705 26.5955
R13968 VDD.n144 VDD.t725 26.5955
R13969 VDD.n144 VDD.t751 26.5955
R13970 VDD.n111 VDD.t661 26.5955
R13971 VDD.n111 VDD.t683 26.5955
R13972 VDD.n239 VDD.t689 26.5955
R13973 VDD.n239 VDD.t715 26.5955
R13974 VDD.n245 VDD.t713 26.5955
R13975 VDD.n245 VDD.t745 26.5955
R13976 VDD.n251 VDD.t757 26.5955
R13977 VDD.n251 VDD.t687 26.5955
R13978 VDD.n256 VDD.t665 26.5955
R13979 VDD.n256 VDD.t729 26.5955
R13980 VDD.n230 VDD.t669 26.5955
R13981 VDD.n230 VDD.t755 26.5955
R13982 VDD.n224 VDD.t703 26.5955
R13983 VDD.n224 VDD.t733 26.5955
R13984 VDD.n343 VDD.t695 26.5955
R13985 VDD.n343 VDD.t719 26.5955
R13986 VDD.n349 VDD.t735 26.5955
R13987 VDD.n349 VDD.t763 26.5955
R13988 VDD.n355 VDD.t711 26.5955
R13989 VDD.n355 VDD.t653 26.5955
R13990 VDD.n361 VDD.t741 26.5955
R13991 VDD.n361 VDD.t675 26.5955
R13992 VDD.n365 VDD.t685 26.5955
R13993 VDD.n365 VDD.t707 26.5955
R13994 VDD.n372 VDD.t727 26.5955
R13995 VDD.n372 VDD.t753 26.5955
R13996 VDD.n380 VDD.t749 26.5955
R13997 VDD.n380 VDD.t775 26.5955
R13998 VDD.n296 VDD.t220 26.5955
R13999 VDD.n296 VDD.t234 26.5955
R14000 VDD.n302 VDD.t232 26.5955
R14001 VDD.n302 VDD.t216 26.5955
R14002 VDD.n308 VDD.t246 26.5955
R14003 VDD.n308 VDD.t226 26.5955
R14004 VDD.n314 VDD.t224 26.5955
R14005 VDD.n314 VDD.t238 26.5955
R14006 VDD.n318 VDD.t236 26.5955
R14007 VDD.n318 VDD.t244 26.5955
R14008 VDD.n324 VDD.t230 26.5955
R14009 VDD.n324 VDD.t240 26.5955
R14010 VDD.n332 VDD.t242 26.5955
R14011 VDD.n332 VDD.t222 26.5955
R14012 VDD.n1352 VDD.t1273 26.5955
R14013 VDD.n1352 VDD.t1275 26.5955
R14014 VDD.n1334 VDD.t1141 26.5955
R14015 VDD.n1334 VDD.t1167 26.5955
R14016 VDD.n1328 VDD.t1163 26.5955
R14017 VDD.n1328 VDD.t1195 26.5955
R14018 VDD.n1321 VDD.t1211 26.5955
R14019 VDD.n1321 VDD.t1137 26.5955
R14020 VDD.n1434 VDD.t1251 26.5955
R14021 VDD.n1434 VDD.t1179 26.5955
R14022 VDD.n1438 VDD.t1175 26.5955
R14023 VDD.n1438 VDD.t1207 26.5955
R14024 VDD.n1444 VDD.t1151 26.5955
R14025 VDD.n1444 VDD.t1247 26.5955
R14026 VDD.n1450 VDD.t1199 26.5955
R14027 VDD.n1450 VDD.t1229 26.5955
R14028 VDD.n1378 VDD.t309 26.5955
R14029 VDD.n1378 VDD.t317 26.5955
R14030 VDD.n1384 VDD.t321 26.5955
R14031 VDD.n1384 VDD.t299 26.5955
R14032 VDD.n1390 VDD.t311 26.5955
R14033 VDD.n1390 VDD.t307 26.5955
R14034 VDD.n1402 VDD.t295 26.5955
R14035 VDD.n1402 VDD.t301 26.5955
R14036 VDD.n1407 VDD.t305 26.5955
R14037 VDD.n1407 VDD.t315 26.5955
R14038 VDD.n1413 VDD.t313 26.5955
R14039 VDD.n1413 VDD.t323 26.5955
R14040 VDD.n1419 VDD.t325 26.5955
R14041 VDD.n1419 VDD.t303 26.5955
R14042 VDD.n1305 VDD.t1143 26.5955
R14043 VDD.n1305 VDD.t1169 26.5955
R14044 VDD.n1298 VDD.t1185 26.5955
R14045 VDD.n1298 VDD.t1217 26.5955
R14046 VDD.n1292 VDD.t1159 26.5955
R14047 VDD.n1292 VDD.t1125 26.5955
R14048 VDD.n1267 VDD.t1191 26.5955
R14049 VDD.n1267 VDD.t1127 26.5955
R14050 VDD.n1271 VDD.t1233 26.5955
R14051 VDD.n1271 VDD.t1155 26.5955
R14052 VDD.n1277 VDD.t1173 26.5955
R14053 VDD.n1277 VDD.t1205 26.5955
R14054 VDD.n1264 VDD.t1201 26.5955
R14055 VDD.n1264 VDD.t1243 26.5955
R14056 VDD.n1464 VDD.t1197 26.5955
R14057 VDD.n1464 VDD.t1133 26.5955
R14058 VDD.n1470 VDD.t1139 26.5955
R14059 VDD.n1470 VDD.t1165 26.5955
R14060 VDD.n1476 VDD.t1161 26.5955
R14061 VDD.n1476 VDD.t1213 26.5955
R14062 VDD.n1482 VDD.t1209 26.5955
R14063 VDD.n1482 VDD.t1237 26.5955
R14064 VDD.n1486 VDD.t1249 26.5955
R14065 VDD.n1486 VDD.t1177 26.5955
R14066 VDD.n1492 VDD.t1135 26.5955
R14067 VDD.n1492 VDD.t1225 26.5955
R14068 VDD.n1498 VDD.t1149 26.5955
R14069 VDD.n1498 VDD.t1183 26.5955
R14070 VDD.n1514 VDD.t1219 26.5955
R14071 VDD.n1514 VDD.t1145 26.5955
R14072 VDD.n1520 VDD.t1239 26.5955
R14073 VDD.n1520 VDD.t1187 26.5955
R14074 VDD.n1256 VDD.t1181 26.5955
R14075 VDD.n1256 VDD.t1215 26.5955
R14076 VDD.n1530 VDD.t1157 26.5955
R14077 VDD.n1530 VDD.t1193 26.5955
R14078 VDD.n1534 VDD.t1189 26.5955
R14079 VDD.n1534 VDD.t1235 26.5955
R14080 VDD.n1252 VDD.t1231 26.5955
R14081 VDD.n1252 VDD.t1153 26.5955
R14082 VDD.n1247 VDD.t1131 26.5955
R14083 VDD.n1247 VDD.t1203 26.5955
R14084 VDD.n812 VDD.n811 25.977
R14085 VDD.n1195 VDD.n1194 25.977
R14086 VDD.t1495 VDD.t1103 25.9096
R14087 VDD.t1489 VDD.t1452 25.9096
R14088 VDD.n672 VDD.t1047 25.6105
R14089 VDD.n1022 VDD.t1432 25.6105
R14090 VDD.n267 VDD.t597 25.6105
R14091 VDD.n819 VDD.n818 25.224
R14092 VDD.n1202 VDD.n1201 25.224
R14093 VDD.t466 VDD.n1847 24.3893
R14094 VDD.t592 VDD.n2168 24.3893
R14095 VDD.t521 VDD.n2426 24.3893
R14096 VDD.t278 VDD.n2684 24.3893
R14097 VDD.t368 VDD.n2942 24.3893
R14098 VDD.t1087 VDD.n3200 24.3893
R14099 VDD.t1093 VDD.n3458 24.3893
R14100 VDD.t514 VDD.n5778 24.3893
R14101 VDD.t507 VDD.n5524 24.3893
R14102 VDD.t251 VDD.n3716 24.3893
R14103 VDD.t266 VDD.n3974 24.3893
R14104 VDD.t13 VDD.n4232 24.3893
R14105 VDD.t415 VDD.n4490 24.3893
R14106 VDD.t527 VDD.n4748 24.3893
R14107 VDD.t815 VDD.n5006 24.3893
R14108 VDD.t265 VDD.n5264 24.3893
R14109 VDD.t491 VDD.t1493 23.0308
R14110 VDD.t645 VDD.t1486 23.0308
R14111 VDD.n408 VDD 22.7027
R14112 VDD.n1566 VDD 22.7027
R14113 VDD.n1660 VDD.n1626 22.5125
R14114 VDD.n1834 VDD.n1833 22.2123
R14115 VDD.n1814 VDD.n1812 22.2123
R14116 VDD.n1784 VDD.n1782 22.2123
R14117 VDD.n1795 VDD.n1794 22.2123
R14118 VDD.n1787 VDD.n1786 22.2123
R14119 VDD.n1789 VDD.n1781 22.2123
R14120 VDD.n2135 VDD.n2133 22.2123
R14121 VDD.n2155 VDD.n2154 22.2123
R14122 VDD.n1992 VDD.n1990 22.2123
R14123 VDD.n2003 VDD.n2002 22.2123
R14124 VDD.n1995 VDD.n1994 22.2123
R14125 VDD.n1997 VDD.n1989 22.2123
R14126 VDD.n2393 VDD.n2391 22.2123
R14127 VDD.n2413 VDD.n2412 22.2123
R14128 VDD.n2363 VDD.n2361 22.2123
R14129 VDD.n2374 VDD.n2373 22.2123
R14130 VDD.n2366 VDD.n2365 22.2123
R14131 VDD.n2368 VDD.n2360 22.2123
R14132 VDD.n2651 VDD.n2649 22.2123
R14133 VDD.n2671 VDD.n2670 22.2123
R14134 VDD.n2621 VDD.n2619 22.2123
R14135 VDD.n2632 VDD.n2631 22.2123
R14136 VDD.n2624 VDD.n2623 22.2123
R14137 VDD.n2626 VDD.n2618 22.2123
R14138 VDD.n2909 VDD.n2907 22.2123
R14139 VDD.n2929 VDD.n2928 22.2123
R14140 VDD.n2879 VDD.n2877 22.2123
R14141 VDD.n2890 VDD.n2889 22.2123
R14142 VDD.n2882 VDD.n2881 22.2123
R14143 VDD.n2884 VDD.n2876 22.2123
R14144 VDD.n3167 VDD.n3165 22.2123
R14145 VDD.n3187 VDD.n3186 22.2123
R14146 VDD.n3137 VDD.n3135 22.2123
R14147 VDD.n3148 VDD.n3147 22.2123
R14148 VDD.n3140 VDD.n3139 22.2123
R14149 VDD.n3142 VDD.n3134 22.2123
R14150 VDD.n3425 VDD.n3423 22.2123
R14151 VDD.n3445 VDD.n3444 22.2123
R14152 VDD.n3395 VDD.n3393 22.2123
R14153 VDD.n3406 VDD.n3405 22.2123
R14154 VDD.n3398 VDD.n3397 22.2123
R14155 VDD.n3400 VDD.n3392 22.2123
R14156 VDD.n5745 VDD.n5743 22.2123
R14157 VDD.n5765 VDD.n5764 22.2123
R14158 VDD.n5718 VDD.n5716 22.2123
R14159 VDD.n5729 VDD.n5728 22.2123
R14160 VDD.n5721 VDD.n5720 22.2123
R14161 VDD.n5723 VDD.n5715 22.2123
R14162 VDD.n5491 VDD.n5489 22.2123
R14163 VDD.n5511 VDD.n5510 22.2123
R14164 VDD.n5464 VDD.n5462 22.2123
R14165 VDD.n5475 VDD.n5474 22.2123
R14166 VDD.n5467 VDD.n5466 22.2123
R14167 VDD.n5469 VDD.n5461 22.2123
R14168 VDD.n3683 VDD.n3681 22.2123
R14169 VDD.n3703 VDD.n3702 22.2123
R14170 VDD.n3653 VDD.n3651 22.2123
R14171 VDD.n3664 VDD.n3663 22.2123
R14172 VDD.n3656 VDD.n3655 22.2123
R14173 VDD.n3658 VDD.n3650 22.2123
R14174 VDD.n3941 VDD.n3939 22.2123
R14175 VDD.n3961 VDD.n3960 22.2123
R14176 VDD.n3911 VDD.n3909 22.2123
R14177 VDD.n3922 VDD.n3921 22.2123
R14178 VDD.n3914 VDD.n3913 22.2123
R14179 VDD.n3916 VDD.n3908 22.2123
R14180 VDD.n4199 VDD.n4197 22.2123
R14181 VDD.n4219 VDD.n4218 22.2123
R14182 VDD.n4169 VDD.n4167 22.2123
R14183 VDD.n4180 VDD.n4179 22.2123
R14184 VDD.n4172 VDD.n4171 22.2123
R14185 VDD.n4174 VDD.n4166 22.2123
R14186 VDD.n4457 VDD.n4455 22.2123
R14187 VDD.n4477 VDD.n4476 22.2123
R14188 VDD.n4427 VDD.n4425 22.2123
R14189 VDD.n4438 VDD.n4437 22.2123
R14190 VDD.n4430 VDD.n4429 22.2123
R14191 VDD.n4432 VDD.n4424 22.2123
R14192 VDD.n4715 VDD.n4713 22.2123
R14193 VDD.n4735 VDD.n4734 22.2123
R14194 VDD.n4685 VDD.n4683 22.2123
R14195 VDD.n4696 VDD.n4695 22.2123
R14196 VDD.n4688 VDD.n4687 22.2123
R14197 VDD.n4690 VDD.n4682 22.2123
R14198 VDD.n4973 VDD.n4971 22.2123
R14199 VDD.n4993 VDD.n4992 22.2123
R14200 VDD.n4943 VDD.n4941 22.2123
R14201 VDD.n4954 VDD.n4953 22.2123
R14202 VDD.n4946 VDD.n4945 22.2123
R14203 VDD.n4948 VDD.n4940 22.2123
R14204 VDD.n5231 VDD.n5229 22.2123
R14205 VDD.n5251 VDD.n5250 22.2123
R14206 VDD.n5201 VDD.n5199 22.2123
R14207 VDD.n5212 VDD.n5211 22.2123
R14208 VDD.n5204 VDD.n5203 22.2123
R14209 VDD.n5206 VDD.n5198 22.2123
R14210 VDD.n813 VDD.n812 22.2123
R14211 VDD.n1196 VDD.n1195 22.2123
R14212 VDD.n1804 VDD.t1028 20.9587
R14213 VDD.n2012 VDD.t1266 20.9587
R14214 VDD.n2383 VDD.t828 20.9587
R14215 VDD.n2641 VDD.t1419 20.9587
R14216 VDD.n2899 VDD.t433 20.9587
R14217 VDD.n3157 VDD.t385 20.9587
R14218 VDD.n3415 VDD.t1297 20.9587
R14219 VDD.n5738 VDD.t473 20.9587
R14220 VDD.n5484 VDD.t1256 20.9587
R14221 VDD.n3673 VDD.t1368 20.9587
R14222 VDD.n3931 VDD.t1111 20.9587
R14223 VDD.n4189 VDD.t27 20.9587
R14224 VDD.n4447 VDD.t1433 20.9587
R14225 VDD.n4705 VDD.t372 20.9587
R14226 VDD.n4963 VDD.t420 20.9587
R14227 VDD.n5221 VDD.t2 20.9587
R14228 VDD.n1507 VDD 20.8224
R14229 VDD.n1457 VDD 20.8224
R14230 VDD.n1707 VDD.n1705 20.5934
R14231 VDD.n2056 VDD.n2054 20.5934
R14232 VDD.n2286 VDD.n2284 20.5934
R14233 VDD.n2544 VDD.n2542 20.5934
R14234 VDD.n2802 VDD.n2800 20.5934
R14235 VDD.n3060 VDD.n3058 20.5934
R14236 VDD.n3318 VDD.n3316 20.5934
R14237 VDD.n5641 VDD.n5639 20.5934
R14238 VDD.n5387 VDD.n5385 20.5934
R14239 VDD.n3576 VDD.n3574 20.5934
R14240 VDD.n3834 VDD.n3832 20.5934
R14241 VDD.n4092 VDD.n4090 20.5934
R14242 VDD.n4350 VDD.n4348 20.5934
R14243 VDD.n4608 VDD.n4606 20.5934
R14244 VDD.n4866 VDD.n4864 20.5934
R14245 VDD.n5124 VDD.n5122 20.5934
R14246 VDD.n13 VDD.n12 19.9534
R14247 VDD.n1157 VDD.n1156 19.9534
R14248 VDD.n1840 VDD.n1839 18.6543
R14249 VDD.n2161 VDD.n2160 18.6543
R14250 VDD.n2419 VDD.n2418 18.6543
R14251 VDD.n2677 VDD.n2676 18.6543
R14252 VDD.n2935 VDD.n2934 18.6543
R14253 VDD.n3193 VDD.n3192 18.6543
R14254 VDD.n3451 VDD.n3450 18.6543
R14255 VDD.n5771 VDD.n5770 18.6543
R14256 VDD.n5517 VDD.n5516 18.6543
R14257 VDD.n3709 VDD.n3708 18.6543
R14258 VDD.n3967 VDD.n3966 18.6543
R14259 VDD.n4225 VDD.n4224 18.6543
R14260 VDD.n4483 VDD.n4482 18.6543
R14261 VDD.n4741 VDD.n4740 18.6543
R14262 VDD.n4999 VDD.n4998 18.6543
R14263 VDD.n5257 VDD.n5256 18.6543
R14264 VDD.n1372 VDD.t296 18.2197
R14265 VDD.n1654 VDD 17.4176
R14266 VDD.n1761 VDD.n1716 17.109
R14267 VDD.n2110 VDD.n2065 17.109
R14268 VDD.n2340 VDD.n2295 17.109
R14269 VDD.n2598 VDD.n2553 17.109
R14270 VDD.n2856 VDD.n2811 17.109
R14271 VDD.n3114 VDD.n3069 17.109
R14272 VDD.n3372 VDD.n3327 17.109
R14273 VDD.n5695 VDD.n5650 17.109
R14274 VDD.n5441 VDD.n5396 17.109
R14275 VDD.n3630 VDD.n3585 17.109
R14276 VDD.n3888 VDD.n3843 17.109
R14277 VDD.n4146 VDD.n4101 17.109
R14278 VDD.n4404 VDD.n4359 17.109
R14279 VDD.n4662 VDD.n4617 17.109
R14280 VDD.n4920 VDD.n4875 17.109
R14281 VDD.n5178 VDD.n5133 17.109
R14282 VDD.n24 VDD.n23 16.9417
R14283 VDD.n575 VDD.n574 16.9417
R14284 VDD.n597 VDD.n596 16.9417
R14285 VDD.n658 VDD.n657 16.9417
R14286 VDD.n768 VDD.n767 16.9417
R14287 VDD.n721 VDD.n720 16.9417
R14288 VDD.n488 VDD.n487 16.9417
R14289 VDD.n86 VDD.n85 16.9417
R14290 VDD.n1168 VDD.n1167 16.9417
R14291 VDD.n925 VDD.n924 16.9417
R14292 VDD.n947 VDD.n946 16.9417
R14293 VDD.n1008 VDD.n1007 16.9417
R14294 VDD.n1118 VDD.n1117 16.9417
R14295 VDD.n1071 VDD.n1070 16.9417
R14296 VDD.n174 VDD.n173 16.9417
R14297 VDD.n196 VDD.n195 16.9417
R14298 VDD.n253 VDD.n252 16.9417
R14299 VDD.n363 VDD.n362 16.9417
R14300 VDD.n316 VDD.n315 16.9417
R14301 VDD.n1436 VDD.n1435 16.9417
R14302 VDD.n1404 VDD.n1403 16.9417
R14303 VDD.n1269 VDD.n1268 16.9417
R14304 VDD.n1484 VDD.n1483 16.9417
R14305 VDD.n1532 VDD.n1531 16.9417
R14306 VDD.n8 VDD.n2 16.1887
R14307 VDD.n1152 VDD.n1146 16.1887
R14308 VDD.n688 VDD.n687 14.5711
R14309 VDD.n1038 VDD.n1037 14.5711
R14310 VDD.n283 VDD.n282 14.5711
R14311 VDD.n1659 VDD 14.551
R14312 VDD.n1686 VDD.t1032 14.2962
R14313 VDD.n2035 VDD.t1271 14.2962
R14314 VDD.n2265 VDD.t832 14.2962
R14315 VDD.n2523 VDD.t1418 14.2962
R14316 VDD.n2781 VDD.t440 14.2962
R14317 VDD.n3039 VDD.t384 14.2962
R14318 VDD.n3297 VDD.t1296 14.2962
R14319 VDD.n5620 VDD.t479 14.2962
R14320 VDD.n5366 VDD.t1259 14.2962
R14321 VDD.n3555 VDD.t1367 14.2962
R14322 VDD.n3813 VDD.t1115 14.2962
R14323 VDD.n4071 VDD.t31 14.2962
R14324 VDD.n4329 VDD.t1440 14.2962
R14325 VDD.n4587 VDD.t375 14.2962
R14326 VDD.n4845 VDD.t1430 14.2962
R14327 VDD.n5103 VDD.t1 14.2962
R14328 VDD.n1666 VDD.t1033 14.2955
R14329 VDD.n2015 VDD.t1265 14.2955
R14330 VDD.n2245 VDD.t835 14.2955
R14331 VDD.n2503 VDD.t1422 14.2955
R14332 VDD.n2761 VDD.t437 14.2955
R14333 VDD.n3019 VDD.t388 14.2955
R14334 VDD.n3277 VDD.t1300 14.2955
R14335 VDD.n5600 VDD.t477 14.2955
R14336 VDD.n5346 VDD.t1262 14.2955
R14337 VDD.n3535 VDD.t1371 14.2955
R14338 VDD.n3793 VDD.t1118 14.2955
R14339 VDD.n4051 VDD.t34 14.2955
R14340 VDD.n4309 VDD.t1437 14.2955
R14341 VDD.n4567 VDD.t371 14.2955
R14342 VDD.n4825 VDD.t423 14.2955
R14343 VDD.n5083 VDD.t1252 14.2955
R14344 VDD.n1749 VDD.t448 14.2865
R14345 VDD.n2098 VDD.t81 14.2865
R14346 VDD.n2328 VDD.t1447 14.2865
R14347 VDD.n2586 VDD.t574 14.2865
R14348 VDD.n2844 VDD.t979 14.2865
R14349 VDD.n3102 VDD.t546 14.2865
R14350 VDD.n3360 VDD.t583 14.2865
R14351 VDD.n5683 VDD.t1469 14.2865
R14352 VDD.n5429 VDD.t1001 14.2865
R14353 VDD.n3618 VDD.t1337 14.2865
R14354 VDD.n3876 VDD.t490 14.2865
R14355 VDD.n4134 VDD.t11 14.2865
R14356 VDD.n4392 VDD.t1053 14.2865
R14357 VDD.n4650 VDD.t22 14.2865
R14358 VDD.n4908 VDD.t821 14.2865
R14359 VDD.n5166 VDD.t1327 14.2865
R14360 VDD.n1737 VDD.t442 14.2864
R14361 VDD.n2086 VDD.t82 14.2864
R14362 VDD.n2316 VDD.t1449 14.2864
R14363 VDD.n2574 VDD.t568 14.2864
R14364 VDD.n2832 VDD.t981 14.2864
R14365 VDD.n3090 VDD.t548 14.2864
R14366 VDD.n3348 VDD.t585 14.2864
R14367 VDD.n5671 VDD.t1471 14.2864
R14368 VDD.n5417 VDD.t996 14.2864
R14369 VDD.n3606 VDD.t1339 14.2864
R14370 VDD.n3864 VDD.t486 14.2864
R14371 VDD.n4122 VDD.t6 14.2864
R14372 VDD.n4380 VDD.t1055 14.2864
R14373 VDD.n4638 VDD.t24 14.2864
R14374 VDD.n4896 VDD.t564 14.2864
R14375 VDD.n5154 VDD.t1009 14.2864
R14376 VDD.n1771 VDD.t1015 14.2849
R14377 VDD.n1753 VDD.t1481 14.2849
R14378 VDD.n2120 VDD.t1304 14.2849
R14379 VDD.n2102 VDD.t624 14.2849
R14380 VDD.n2350 VDD.t1362 14.2849
R14381 VDD.n2332 VDD.t1332 14.2849
R14382 VDD.n2608 VDD.t826 14.2849
R14383 VDD.n2590 VDD.t1427 14.2849
R14384 VDD.n2866 VDD.t425 14.2849
R14385 VDD.n2848 VDD.t1476 14.2849
R14386 VDD.n3124 VDD.t641 14.2849
R14387 VDD.n3106 VDD.t396 14.2849
R14388 VDD.n3382 VDD.t1425 14.2849
R14389 VDD.n3364 VDD.t640 14.2849
R14390 VDD.n5705 VDD.t1308 14.2849
R14391 VDD.n5687 VDD.t1428 14.2849
R14392 VDD.n5451 VDD.t508 14.2849
R14393 VDD.n5433 VDD.t271 14.2849
R14394 VDD.n3640 VDD.t1477 14.2849
R14395 VDD.n3622 VDD.t250 14.2849
R14396 VDD.n3898 VDD.t1318 14.2849
R14397 VDD.n3880 VDD.t1330 14.2849
R14398 VDD.n4156 VDD.t1255 14.2849
R14399 VDD.n4138 VDD.t410 14.2849
R14400 VDD.n4414 VDD.t1291 14.2849
R14401 VDD.n4396 VDD.t1109 14.2849
R14402 VDD.n4672 VDD.t333 14.2849
R14403 VDD.n4654 VDD.t994 14.2849
R14404 VDD.n4930 VDD.t280 14.2849
R14405 VDD.n4912 VDD.t827 14.2849
R14406 VDD.n5188 VDD.t1095 14.2849
R14407 VDD.n5170 VDD.t1061 14.2849
R14408 VDD.n1620 VDD.n1619 14.1868
R14409 VDD.n1769 VDD.n1669 14.0805
R14410 VDD.n2118 VDD.n2018 14.0805
R14411 VDD.n2348 VDD.n2248 14.0805
R14412 VDD.n2606 VDD.n2506 14.0805
R14413 VDD.n2864 VDD.n2764 14.0805
R14414 VDD.n3122 VDD.n3022 14.0805
R14415 VDD.n3380 VDD.n3280 14.0805
R14416 VDD.n5703 VDD.n5603 14.0805
R14417 VDD.n5449 VDD.n5349 14.0805
R14418 VDD.n3638 VDD.n3538 14.0805
R14419 VDD.n3896 VDD.n3796 14.0805
R14420 VDD.n4154 VDD.n4054 14.0805
R14421 VDD.n4412 VDD.n4312 14.0805
R14422 VDD.n4670 VDD.n4570 14.0805
R14423 VDD.n4928 VDD.n4828 14.0805
R14424 VDD.n5186 VDD.n5086 14.0805
R14425 VDD.t326 VDD.t967 13.9711
R14426 VDD.t362 VDD.t364 13.9711
R14427 VDD.t791 VDD.t649 13.9711
R14428 VDD.t509 VDD.t1119 13.9711
R14429 VDD.n1755 VDD.n1717 13.7605
R14430 VDD.n2104 VDD.n2066 13.7605
R14431 VDD.n2334 VDD.n2296 13.7605
R14432 VDD.n2592 VDD.n2554 13.7605
R14433 VDD.n2850 VDD.n2812 13.7605
R14434 VDD.n3108 VDD.n3070 13.7605
R14435 VDD.n3366 VDD.n3328 13.7605
R14436 VDD.n5689 VDD.n5651 13.7605
R14437 VDD.n5435 VDD.n5397 13.7605
R14438 VDD.n3624 VDD.n3586 13.7605
R14439 VDD.n3882 VDD.n3844 13.7605
R14440 VDD.n4140 VDD.n4102 13.7605
R14441 VDD.n4398 VDD.n4360 13.7605
R14442 VDD.n4656 VDD.n4618 13.7605
R14443 VDD.n4914 VDD.n4876 13.7605
R14444 VDD.n5172 VDD.n5134 13.7605
R14445 VDD.n1658 VDD.n1631 13.4428
R14446 VDD.n1657 VDD 13.4235
R14447 VDD.n807 VDD.n805 13.3488
R14448 VDD.n1190 VDD.n1188 13.3488
R14449 VDD.n827 VDD.n826 12.9329
R14450 VDD.n1543 VDD.n1542 12.9329
R14451 VDD.n1363 VDD.n1362 12.9329
R14452 VDD.n1210 VDD.n1209 12.9329
R14453 VDD.n580 VDD.n579 11.6711
R14454 VDD.n593 VDD.n592 11.6711
R14455 VDD.n663 VDD.n662 11.6711
R14456 VDD.n772 VDD.n771 11.6711
R14457 VDD.n725 VDD.n724 11.6711
R14458 VDD.n930 VDD.n929 11.6711
R14459 VDD.n943 VDD.n942 11.6711
R14460 VDD.n1013 VDD.n1012 11.6711
R14461 VDD.n1122 VDD.n1121 11.6711
R14462 VDD.n1075 VDD.n1074 11.6711
R14463 VDD.n179 VDD.n178 11.6711
R14464 VDD.n192 VDD.n191 11.6711
R14465 VDD.n258 VDD.n257 11.6711
R14466 VDD.n367 VDD.n366 11.6711
R14467 VDD.n320 VDD.n319 11.6711
R14468 VDD.n1440 VDD.n1439 11.6711
R14469 VDD.n1409 VDD.n1408 11.6711
R14470 VDD.n1273 VDD.n1272 11.6711
R14471 VDD.n1488 VDD.n1487 11.6711
R14472 VDD.n1536 VDD.n1535 11.6711
R14473 VDD.n569 VDD.n568 10.9181
R14474 VDD.n603 VDD.n602 10.9181
R14475 VDD.n652 VDD.n651 10.9181
R14476 VDD.n762 VDD.n761 10.9181
R14477 VDD.n715 VDD.n714 10.9181
R14478 VDD.n919 VDD.n918 10.9181
R14479 VDD.n953 VDD.n952 10.9181
R14480 VDD.n1002 VDD.n1001 10.9181
R14481 VDD.n1112 VDD.n1111 10.9181
R14482 VDD.n1065 VDD.n1064 10.9181
R14483 VDD.n168 VDD.n167 10.9181
R14484 VDD.n202 VDD.n201 10.9181
R14485 VDD.n247 VDD.n246 10.9181
R14486 VDD.n357 VDD.n356 10.9181
R14487 VDD.n310 VDD.n309 10.9181
R14488 VDD.n1323 VDD.n1322 10.9181
R14489 VDD.n1392 VDD.n1391 10.9181
R14490 VDD.n1294 VDD.n1293 10.9181
R14491 VDD.n1478 VDD.n1477 10.9181
R14492 VDD.n1258 VDD.n1257 10.9181
R14493 VDD.n1957 VDD.n1956 10.8802
R14494 VDD.n463 VDD 10.8576
R14495 VDD.n60 VDD 10.8576
R14496 VDD.n1955 VDD.n1954 10.5887
R14497 VDD.n1429 VDD.t1210 10.4115
R14498 VDD.n668 VDD.t173 10.1791
R14499 VDD.n1018 VDD.t946 10.1791
R14500 VDD.t221 VDD.n264 10.1791
R14501 VDD.n1617 VDD 9.58775
R14502 VDD.n9 VDD.n6 9.41227
R14503 VDD.n1153 VDD.n1150 9.41227
R14504 VDD.n1954 VDD.n1953 9.3005
R14505 VDD.n1916 VDD.n1915 9.3005
R14506 VDD.n1915 VDD.n1914 9.3005
R14507 VDD.n1828 VDD.n1826 9.3005
R14508 VDD.n1747 VDD.n1746 9.3005
R14509 VDD.n1728 VDD.n1727 9.3005
R14510 VDD.n1731 VDD.n1722 9.3005
R14511 VDD.n1705 VDD.n1667 9.3005
R14512 VDD.n1690 VDD.n1689 9.3005
R14513 VDD.n2096 VDD.n2095 9.3005
R14514 VDD.n2077 VDD.n2076 9.3005
R14515 VDD.n2080 VDD.n2071 9.3005
R14516 VDD.n2054 VDD.n2016 9.3005
R14517 VDD.n2039 VDD.n2038 9.3005
R14518 VDD.n2237 VDD.n2236 9.3005
R14519 VDD.n2236 VDD.n2235 9.3005
R14520 VDD.n2149 VDD.n2147 9.3005
R14521 VDD.n2326 VDD.n2325 9.3005
R14522 VDD.n2307 VDD.n2306 9.3005
R14523 VDD.n2310 VDD.n2301 9.3005
R14524 VDD.n2284 VDD.n2246 9.3005
R14525 VDD.n2269 VDD.n2268 9.3005
R14526 VDD.n2495 VDD.n2494 9.3005
R14527 VDD.n2494 VDD.n2493 9.3005
R14528 VDD.n2407 VDD.n2405 9.3005
R14529 VDD.n2584 VDD.n2583 9.3005
R14530 VDD.n2565 VDD.n2564 9.3005
R14531 VDD.n2568 VDD.n2559 9.3005
R14532 VDD.n2542 VDD.n2504 9.3005
R14533 VDD.n2527 VDD.n2526 9.3005
R14534 VDD.n2753 VDD.n2752 9.3005
R14535 VDD.n2752 VDD.n2751 9.3005
R14536 VDD.n2665 VDD.n2663 9.3005
R14537 VDD.n2842 VDD.n2841 9.3005
R14538 VDD.n2823 VDD.n2822 9.3005
R14539 VDD.n2826 VDD.n2817 9.3005
R14540 VDD.n2800 VDD.n2762 9.3005
R14541 VDD.n2785 VDD.n2784 9.3005
R14542 VDD.n3011 VDD.n3010 9.3005
R14543 VDD.n3010 VDD.n3009 9.3005
R14544 VDD.n2923 VDD.n2921 9.3005
R14545 VDD.n3100 VDD.n3099 9.3005
R14546 VDD.n3081 VDD.n3080 9.3005
R14547 VDD.n3084 VDD.n3075 9.3005
R14548 VDD.n3058 VDD.n3020 9.3005
R14549 VDD.n3043 VDD.n3042 9.3005
R14550 VDD.n3269 VDD.n3268 9.3005
R14551 VDD.n3268 VDD.n3267 9.3005
R14552 VDD.n3181 VDD.n3179 9.3005
R14553 VDD.n3358 VDD.n3357 9.3005
R14554 VDD.n3339 VDD.n3338 9.3005
R14555 VDD.n3342 VDD.n3333 9.3005
R14556 VDD.n3316 VDD.n3278 9.3005
R14557 VDD.n3301 VDD.n3300 9.3005
R14558 VDD.n3527 VDD.n3526 9.3005
R14559 VDD.n3526 VDD.n3525 9.3005
R14560 VDD.n3439 VDD.n3437 9.3005
R14561 VDD.n5681 VDD.n5680 9.3005
R14562 VDD.n5662 VDD.n5661 9.3005
R14563 VDD.n5665 VDD.n5656 9.3005
R14564 VDD.n5639 VDD.n5601 9.3005
R14565 VDD.n5624 VDD.n5623 9.3005
R14566 VDD.n5847 VDD.n5846 9.3005
R14567 VDD.n5846 VDD.n5845 9.3005
R14568 VDD.n5759 VDD.n5757 9.3005
R14569 VDD.n5427 VDD.n5426 9.3005
R14570 VDD.n5408 VDD.n5407 9.3005
R14571 VDD.n5411 VDD.n5402 9.3005
R14572 VDD.n5385 VDD.n5347 9.3005
R14573 VDD.n5370 VDD.n5369 9.3005
R14574 VDD.n5593 VDD.n5592 9.3005
R14575 VDD.n5592 VDD.n5591 9.3005
R14576 VDD.n5505 VDD.n5503 9.3005
R14577 VDD.n3616 VDD.n3615 9.3005
R14578 VDD.n3597 VDD.n3596 9.3005
R14579 VDD.n3600 VDD.n3591 9.3005
R14580 VDD.n3574 VDD.n3536 9.3005
R14581 VDD.n3559 VDD.n3558 9.3005
R14582 VDD.n3785 VDD.n3784 9.3005
R14583 VDD.n3784 VDD.n3783 9.3005
R14584 VDD.n3697 VDD.n3695 9.3005
R14585 VDD.n3874 VDD.n3873 9.3005
R14586 VDD.n3855 VDD.n3854 9.3005
R14587 VDD.n3858 VDD.n3849 9.3005
R14588 VDD.n3832 VDD.n3794 9.3005
R14589 VDD.n3817 VDD.n3816 9.3005
R14590 VDD.n4043 VDD.n4042 9.3005
R14591 VDD.n4042 VDD.n4041 9.3005
R14592 VDD.n3955 VDD.n3953 9.3005
R14593 VDD.n4132 VDD.n4131 9.3005
R14594 VDD.n4113 VDD.n4112 9.3005
R14595 VDD.n4116 VDD.n4107 9.3005
R14596 VDD.n4090 VDD.n4052 9.3005
R14597 VDD.n4075 VDD.n4074 9.3005
R14598 VDD.n4301 VDD.n4300 9.3005
R14599 VDD.n4300 VDD.n4299 9.3005
R14600 VDD.n4213 VDD.n4211 9.3005
R14601 VDD.n4390 VDD.n4389 9.3005
R14602 VDD.n4371 VDD.n4370 9.3005
R14603 VDD.n4374 VDD.n4365 9.3005
R14604 VDD.n4348 VDD.n4310 9.3005
R14605 VDD.n4333 VDD.n4332 9.3005
R14606 VDD.n4559 VDD.n4558 9.3005
R14607 VDD.n4558 VDD.n4557 9.3005
R14608 VDD.n4471 VDD.n4469 9.3005
R14609 VDD.n4648 VDD.n4647 9.3005
R14610 VDD.n4629 VDD.n4628 9.3005
R14611 VDD.n4632 VDD.n4623 9.3005
R14612 VDD.n4606 VDD.n4568 9.3005
R14613 VDD.n4591 VDD.n4590 9.3005
R14614 VDD.n4817 VDD.n4816 9.3005
R14615 VDD.n4816 VDD.n4815 9.3005
R14616 VDD.n4729 VDD.n4727 9.3005
R14617 VDD.n4906 VDD.n4905 9.3005
R14618 VDD.n4887 VDD.n4886 9.3005
R14619 VDD.n4890 VDD.n4881 9.3005
R14620 VDD.n4864 VDD.n4826 9.3005
R14621 VDD.n4849 VDD.n4848 9.3005
R14622 VDD.n5075 VDD.n5074 9.3005
R14623 VDD.n5074 VDD.n5073 9.3005
R14624 VDD.n4987 VDD.n4985 9.3005
R14625 VDD.n5164 VDD.n5163 9.3005
R14626 VDD.n5145 VDD.n5144 9.3005
R14627 VDD.n5148 VDD.n5139 9.3005
R14628 VDD.n5122 VDD.n5084 9.3005
R14629 VDD.n5107 VDD.n5106 9.3005
R14630 VDD.n5333 VDD.n5332 9.3005
R14631 VDD.n5332 VDD.n5331 9.3005
R14632 VDD.n5245 VDD.n5243 9.3005
R14633 VDD.n1618 VDD.n1617 9.3005
R14634 VDD VDD.n1628 9.22489
R14635 VDD.n1646 VDD.n1645 9.0245
R14636 VDD.n1734 VDD.n1733 8.88939
R14637 VDD.n2083 VDD.n2082 8.88939
R14638 VDD.n2313 VDD.n2312 8.88939
R14639 VDD.n2571 VDD.n2570 8.88939
R14640 VDD.n2829 VDD.n2828 8.88939
R14641 VDD.n3087 VDD.n3086 8.88939
R14642 VDD.n3345 VDD.n3344 8.88939
R14643 VDD.n5668 VDD.n5667 8.88939
R14644 VDD.n5414 VDD.n5413 8.88939
R14645 VDD.n3603 VDD.n3602 8.88939
R14646 VDD.n3861 VDD.n3860 8.88939
R14647 VDD.n4119 VDD.n4118 8.88939
R14648 VDD.n4377 VDD.n4376 8.88939
R14649 VDD.n4635 VDD.n4634 8.88939
R14650 VDD.n4893 VDD.n4892 8.88939
R14651 VDD.n5151 VDD.n5150 8.88939
R14652 VDD.n1954 VDD.n1943 8.85536
R14653 VDD.n10 VDD.n9 8.79168
R14654 VDD.n413 VDD.n412 8.79168
R14655 VDD.n413 VDD.n411 8.79168
R14656 VDD.n394 VDD.n393 8.79168
R14657 VDD.n1154 VDD.n1153 8.79168
R14658 VDD.n1571 VDD.n1570 8.79168
R14659 VDD.n1571 VDD.n1569 8.79168
R14660 VDD.n1552 VDD.n1551 8.79168
R14661 VDD.n1652 VDD.n1649 8.76429
R14662 VDD.n679 VDD.n671 8.28285
R14663 VDD.n832 VDD.n825 8.28285
R14664 VDD.n838 VDD.n824 8.28285
R14665 VDD.n844 VDD.n823 8.28285
R14666 VDD.n850 VDD.n822 8.28285
R14667 VDD.n1029 VDD.n1021 8.28285
R14668 VDD.n274 VDD.n266 8.28285
R14669 VDD.n1215 VDD.n1208 8.28285
R14670 VDD.n1221 VDD.n1207 8.28285
R14671 VDD.n1227 VDD.n1206 8.28285
R14672 VDD.n1233 VDD.n1205 8.28285
R14673 VDD.n1977 VDD.n1923 7.681
R14674 VDD.n1628 VDD 7.6805
R14675 VDD.n1618 VDD.n1616 7.60183
R14676 VDD.n424 VDD.n423 7.54105
R14677 VDD.n403 VDD.n402 7.54105
R14678 VDD.n1582 VDD.n1581 7.54105
R14679 VDD.n1561 VDD.n1560 7.54105
R14680 VDD.n1885 VDD.n1818 7.49764
R14681 VDD.n2206 VDD.n2139 7.49764
R14682 VDD.n2464 VDD.n2397 7.49764
R14683 VDD.n2722 VDD.n2655 7.49764
R14684 VDD.n2980 VDD.n2913 7.49764
R14685 VDD.n3238 VDD.n3171 7.49764
R14686 VDD.n3496 VDD.n3429 7.49764
R14687 VDD.n5816 VDD.n5749 7.49764
R14688 VDD.n5562 VDD.n5495 7.49764
R14689 VDD.n3754 VDD.n3687 7.49764
R14690 VDD.n4012 VDD.n3945 7.49764
R14691 VDD.n4270 VDD.n4203 7.49764
R14692 VDD.n4528 VDD.n4461 7.49764
R14693 VDD.n4786 VDD.n4719 7.49764
R14694 VDD.n5044 VDD.n4977 7.49764
R14695 VDD.n5302 VDD.n5235 7.49764
R14696 VDD.n1606 VDD.n1605 7.39078
R14697 VDD.n1636 VDD.n1635 7.27155
R14698 VDD.n1917 VDD.t284 7.15136
R14699 VDD.n2238 VDD.t1010 7.15136
R14700 VDD.n2496 VDD.t617 7.15136
R14701 VDD.n2754 VDD.t1329 7.15136
R14702 VDD.n3012 VDD.t620 7.15136
R14703 VDD.n3270 VDD.t283 7.15136
R14704 VDD.n3528 VDD.t1378 7.15136
R14705 VDD.n5848 VDD.t1355 7.15136
R14706 VDD.n5594 VDD.t394 7.15136
R14707 VDD.n3786 VDD.t293 7.15136
R14708 VDD.n4044 VDD.t1350 7.15136
R14709 VDD.n4302 VDD.t1365 7.15136
R14710 VDD.n4560 VDD.t610 7.15136
R14711 VDD.n4818 VDD.t402 7.15136
R14712 VDD.n5076 VDD.t1098 7.15136
R14713 VDD.n5334 VDD.t408 7.15136
R14714 VDD.n1872 VDD.t467 7.14897
R14715 VDD.n2193 VDD.t1429 7.14897
R14716 VDD.n2451 VDD.t1016 7.14897
R14717 VDD.n2709 VDD.t1325 7.14897
R14718 VDD.n2967 VDD.t369 7.14897
R14719 VDD.n3225 VDD.t1461 7.14897
R14720 VDD.n3483 VDD.t1094 7.14897
R14721 VDD.n5803 VDD.t783 7.14897
R14722 VDD.n5549 VDD.t642 7.14897
R14723 VDD.n3741 VDD.t252 7.14897
R14724 VDD.n3999 VDD.t267 7.14897
R14725 VDD.n4257 VDD.t14 7.14897
R14726 VDD.n4515 VDD.t1069 7.14897
R14727 VDD.n4773 VDD.t1313 7.14897
R14728 VDD.n5031 VDD.t816 7.14897
R14729 VDD.n5289 VDD.t413 7.14897
R14730 VDD.n1976 VDD.n1926 7.05932
R14731 VDD.n1625 VDD 6.73734
R14732 VDD.n1833 VDD 6.4005
R14733 VDD.n1812 VDD 6.4005
R14734 VDD.n2133 VDD 6.4005
R14735 VDD.n2154 VDD 6.4005
R14736 VDD.n2391 VDD 6.4005
R14737 VDD.n2412 VDD 6.4005
R14738 VDD.n2649 VDD 6.4005
R14739 VDD.n2670 VDD 6.4005
R14740 VDD.n2907 VDD 6.4005
R14741 VDD.n2928 VDD 6.4005
R14742 VDD.n3165 VDD 6.4005
R14743 VDD.n3186 VDD 6.4005
R14744 VDD.n3423 VDD 6.4005
R14745 VDD.n3444 VDD 6.4005
R14746 VDD.n5743 VDD 6.4005
R14747 VDD.n5764 VDD 6.4005
R14748 VDD.n5489 VDD 6.4005
R14749 VDD.n5510 VDD 6.4005
R14750 VDD.n3681 VDD 6.4005
R14751 VDD.n3702 VDD 6.4005
R14752 VDD.n3939 VDD 6.4005
R14753 VDD.n3960 VDD 6.4005
R14754 VDD.n4197 VDD 6.4005
R14755 VDD.n4218 VDD 6.4005
R14756 VDD.n4455 VDD 6.4005
R14757 VDD.n4476 VDD 6.4005
R14758 VDD.n4713 VDD 6.4005
R14759 VDD.n4734 VDD 6.4005
R14760 VDD.n4971 VDD 6.4005
R14761 VDD.n4992 VDD 6.4005
R14762 VDD.n5229 VDD 6.4005
R14763 VDD.n5250 VDD 6.4005
R14764 VDD.n19 VDD.n18 6.4005
R14765 VDD.n1163 VDD.n1162 6.4005
R14766 VDD.n1646 VDD.n1644 6.23487
R14767 VDD.n1652 VDD 5.65631
R14768 VDD.n1631 VDD 5.65631
R14769 VDD.n536 VDD.n535 5.64756
R14770 VDD.n527 VDD.n526 5.64756
R14771 VDD.n633 VDD.n632 5.64756
R14772 VDD.n779 VDD.n778 5.64756
R14773 VDD.n731 VDD.n730 5.64756
R14774 VDD.n886 VDD.n885 5.64756
R14775 VDD.n877 VDD.n876 5.64756
R14776 VDD.n983 VDD.n982 5.64756
R14777 VDD.n1129 VDD.n1128 5.64756
R14778 VDD.n1081 VDD.n1080 5.64756
R14779 VDD.n135 VDD.n134 5.64756
R14780 VDD.n126 VDD.n125 5.64756
R14781 VDD.n232 VDD.n231 5.64756
R14782 VDD.n374 VDD.n373 5.64756
R14783 VDD.n326 VDD.n325 5.64756
R14784 VDD.n1446 VDD.n1445 5.64756
R14785 VDD.n1415 VDD.n1414 5.64756
R14786 VDD.n1279 VDD.n1278 5.64756
R14787 VDD.n1494 VDD.n1493 5.64756
R14788 VDD.n1254 VDD.n1253 5.64756
R14789 VDD.n2128 VDD.n2013 5.34133
R14790 VDD.n1626 VDD 5.31371
R14791 VDD.n1360 VDD.n1359 5.27114
R14792 VDD.n1505 VDD.n1504 5.27114
R14793 VDD.n1288 VDD.n1287 5.27114
R14794 VDD.n1428 VDD.t318 5.20598
R14795 VDD.n1653 VDD.n1652 4.99699
R14796 VDD.n1648 VDD.n1647 4.98671
R14797 VDD.n563 VDD.n562 4.89462
R14798 VDD.n609 VDD.n608 4.89462
R14799 VDD.n646 VDD.n645 4.89462
R14800 VDD.n756 VDD.n755 4.89462
R14801 VDD.n709 VDD.n708 4.89462
R14802 VDD.n913 VDD.n912 4.89462
R14803 VDD.n959 VDD.n958 4.89462
R14804 VDD.n996 VDD.n995 4.89462
R14805 VDD.n1106 VDD.n1105 4.89462
R14806 VDD.n1059 VDD.n1058 4.89462
R14807 VDD.n162 VDD.n161 4.89462
R14808 VDD.n208 VDD.n207 4.89462
R14809 VDD.n241 VDD.n240 4.89462
R14810 VDD.n351 VDD.n350 4.89462
R14811 VDD.n304 VDD.n303 4.89462
R14812 VDD.n1330 VDD.n1329 4.89462
R14813 VDD.n1386 VDD.n1385 4.89462
R14814 VDD.n1300 VDD.n1299 4.89462
R14815 VDD.n1472 VDD.n1471 4.89462
R14816 VDD.n1522 VDD.n1521 4.89462
R14817 VDD.n1618 VDD 4.8645
R14818 VDD.n1833 VDD.n1832 4.6505
R14819 VDD.n1834 VDD.n1829 4.6505
R14820 VDD.n1812 VDD.n1811 4.6505
R14821 VDD.n1796 VDD.n1781 4.6505
R14822 VDD.n1796 VDD.n1795 4.6505
R14823 VDD.n1791 VDD.n1790 4.6505
R14824 VDD.n1793 VDD.n1791 4.6505
R14825 VDD.n1789 VDD.n1780 4.6505
R14826 VDD.n1787 VDD.n1783 4.6505
R14827 VDD.n1786 VDD.n1785 4.6505
R14828 VDD.n1794 VDD.n1780 4.6505
R14829 VDD.n1783 VDD.n1782 4.6505
R14830 VDD.n1785 VDD.n1784 4.6505
R14831 VDD.n2133 VDD.n2132 4.6505
R14832 VDD.n2154 VDD.n2153 4.6505
R14833 VDD.n2155 VDD.n2150 4.6505
R14834 VDD.n2004 VDD.n1989 4.6505
R14835 VDD.n2004 VDD.n2003 4.6505
R14836 VDD.n1999 VDD.n1998 4.6505
R14837 VDD.n2001 VDD.n1999 4.6505
R14838 VDD.n1997 VDD.n1988 4.6505
R14839 VDD.n1995 VDD.n1991 4.6505
R14840 VDD.n1994 VDD.n1993 4.6505
R14841 VDD.n2002 VDD.n1988 4.6505
R14842 VDD.n1991 VDD.n1990 4.6505
R14843 VDD.n1993 VDD.n1992 4.6505
R14844 VDD.n2391 VDD.n2390 4.6505
R14845 VDD.n2412 VDD.n2411 4.6505
R14846 VDD.n2413 VDD.n2408 4.6505
R14847 VDD.n2375 VDD.n2360 4.6505
R14848 VDD.n2375 VDD.n2374 4.6505
R14849 VDD.n2370 VDD.n2369 4.6505
R14850 VDD.n2372 VDD.n2370 4.6505
R14851 VDD.n2368 VDD.n2359 4.6505
R14852 VDD.n2366 VDD.n2362 4.6505
R14853 VDD.n2365 VDD.n2364 4.6505
R14854 VDD.n2373 VDD.n2359 4.6505
R14855 VDD.n2362 VDD.n2361 4.6505
R14856 VDD.n2364 VDD.n2363 4.6505
R14857 VDD.n2649 VDD.n2648 4.6505
R14858 VDD.n2670 VDD.n2669 4.6505
R14859 VDD.n2671 VDD.n2666 4.6505
R14860 VDD.n2633 VDD.n2618 4.6505
R14861 VDD.n2633 VDD.n2632 4.6505
R14862 VDD.n2628 VDD.n2627 4.6505
R14863 VDD.n2630 VDD.n2628 4.6505
R14864 VDD.n2626 VDD.n2617 4.6505
R14865 VDD.n2624 VDD.n2620 4.6505
R14866 VDD.n2623 VDD.n2622 4.6505
R14867 VDD.n2631 VDD.n2617 4.6505
R14868 VDD.n2620 VDD.n2619 4.6505
R14869 VDD.n2622 VDD.n2621 4.6505
R14870 VDD.n2907 VDD.n2906 4.6505
R14871 VDD.n2928 VDD.n2927 4.6505
R14872 VDD.n2929 VDD.n2924 4.6505
R14873 VDD.n2891 VDD.n2876 4.6505
R14874 VDD.n2891 VDD.n2890 4.6505
R14875 VDD.n2886 VDD.n2885 4.6505
R14876 VDD.n2888 VDD.n2886 4.6505
R14877 VDD.n2884 VDD.n2875 4.6505
R14878 VDD.n2882 VDD.n2878 4.6505
R14879 VDD.n2881 VDD.n2880 4.6505
R14880 VDD.n2889 VDD.n2875 4.6505
R14881 VDD.n2878 VDD.n2877 4.6505
R14882 VDD.n2880 VDD.n2879 4.6505
R14883 VDD.n3165 VDD.n3164 4.6505
R14884 VDD.n3186 VDD.n3185 4.6505
R14885 VDD.n3187 VDD.n3182 4.6505
R14886 VDD.n3149 VDD.n3134 4.6505
R14887 VDD.n3149 VDD.n3148 4.6505
R14888 VDD.n3144 VDD.n3143 4.6505
R14889 VDD.n3146 VDD.n3144 4.6505
R14890 VDD.n3142 VDD.n3133 4.6505
R14891 VDD.n3140 VDD.n3136 4.6505
R14892 VDD.n3139 VDD.n3138 4.6505
R14893 VDD.n3147 VDD.n3133 4.6505
R14894 VDD.n3136 VDD.n3135 4.6505
R14895 VDD.n3138 VDD.n3137 4.6505
R14896 VDD.n3423 VDD.n3422 4.6505
R14897 VDD.n3444 VDD.n3443 4.6505
R14898 VDD.n3445 VDD.n3440 4.6505
R14899 VDD.n3407 VDD.n3392 4.6505
R14900 VDD.n3407 VDD.n3406 4.6505
R14901 VDD.n3402 VDD.n3401 4.6505
R14902 VDD.n3404 VDD.n3402 4.6505
R14903 VDD.n3400 VDD.n3391 4.6505
R14904 VDD.n3398 VDD.n3394 4.6505
R14905 VDD.n3397 VDD.n3396 4.6505
R14906 VDD.n3405 VDD.n3391 4.6505
R14907 VDD.n3394 VDD.n3393 4.6505
R14908 VDD.n3396 VDD.n3395 4.6505
R14909 VDD.n5743 VDD.n5742 4.6505
R14910 VDD.n5764 VDD.n5763 4.6505
R14911 VDD.n5765 VDD.n5760 4.6505
R14912 VDD.n5730 VDD.n5715 4.6505
R14913 VDD.n5730 VDD.n5729 4.6505
R14914 VDD.n5725 VDD.n5724 4.6505
R14915 VDD.n5727 VDD.n5725 4.6505
R14916 VDD.n5723 VDD.n5714 4.6505
R14917 VDD.n5721 VDD.n5717 4.6505
R14918 VDD.n5720 VDD.n5719 4.6505
R14919 VDD.n5728 VDD.n5714 4.6505
R14920 VDD.n5717 VDD.n5716 4.6505
R14921 VDD.n5719 VDD.n5718 4.6505
R14922 VDD.n5489 VDD.n5488 4.6505
R14923 VDD.n5510 VDD.n5509 4.6505
R14924 VDD.n5511 VDD.n5506 4.6505
R14925 VDD.n5476 VDD.n5461 4.6505
R14926 VDD.n5476 VDD.n5475 4.6505
R14927 VDD.n5471 VDD.n5470 4.6505
R14928 VDD.n5473 VDD.n5471 4.6505
R14929 VDD.n5469 VDD.n5460 4.6505
R14930 VDD.n5467 VDD.n5463 4.6505
R14931 VDD.n5466 VDD.n5465 4.6505
R14932 VDD.n5474 VDD.n5460 4.6505
R14933 VDD.n5463 VDD.n5462 4.6505
R14934 VDD.n5465 VDD.n5464 4.6505
R14935 VDD.n3681 VDD.n3680 4.6505
R14936 VDD.n3702 VDD.n3701 4.6505
R14937 VDD.n3703 VDD.n3698 4.6505
R14938 VDD.n3665 VDD.n3650 4.6505
R14939 VDD.n3665 VDD.n3664 4.6505
R14940 VDD.n3660 VDD.n3659 4.6505
R14941 VDD.n3662 VDD.n3660 4.6505
R14942 VDD.n3658 VDD.n3649 4.6505
R14943 VDD.n3656 VDD.n3652 4.6505
R14944 VDD.n3655 VDD.n3654 4.6505
R14945 VDD.n3663 VDD.n3649 4.6505
R14946 VDD.n3652 VDD.n3651 4.6505
R14947 VDD.n3654 VDD.n3653 4.6505
R14948 VDD.n3939 VDD.n3938 4.6505
R14949 VDD.n3960 VDD.n3959 4.6505
R14950 VDD.n3961 VDD.n3956 4.6505
R14951 VDD.n3923 VDD.n3908 4.6505
R14952 VDD.n3923 VDD.n3922 4.6505
R14953 VDD.n3918 VDD.n3917 4.6505
R14954 VDD.n3920 VDD.n3918 4.6505
R14955 VDD.n3916 VDD.n3907 4.6505
R14956 VDD.n3914 VDD.n3910 4.6505
R14957 VDD.n3913 VDD.n3912 4.6505
R14958 VDD.n3921 VDD.n3907 4.6505
R14959 VDD.n3910 VDD.n3909 4.6505
R14960 VDD.n3912 VDD.n3911 4.6505
R14961 VDD.n4197 VDD.n4196 4.6505
R14962 VDD.n4218 VDD.n4217 4.6505
R14963 VDD.n4219 VDD.n4214 4.6505
R14964 VDD.n4181 VDD.n4166 4.6505
R14965 VDD.n4181 VDD.n4180 4.6505
R14966 VDD.n4176 VDD.n4175 4.6505
R14967 VDD.n4178 VDD.n4176 4.6505
R14968 VDD.n4174 VDD.n4165 4.6505
R14969 VDD.n4172 VDD.n4168 4.6505
R14970 VDD.n4171 VDD.n4170 4.6505
R14971 VDD.n4179 VDD.n4165 4.6505
R14972 VDD.n4168 VDD.n4167 4.6505
R14973 VDD.n4170 VDD.n4169 4.6505
R14974 VDD.n4455 VDD.n4454 4.6505
R14975 VDD.n4476 VDD.n4475 4.6505
R14976 VDD.n4477 VDD.n4472 4.6505
R14977 VDD.n4439 VDD.n4424 4.6505
R14978 VDD.n4439 VDD.n4438 4.6505
R14979 VDD.n4434 VDD.n4433 4.6505
R14980 VDD.n4436 VDD.n4434 4.6505
R14981 VDD.n4432 VDD.n4423 4.6505
R14982 VDD.n4430 VDD.n4426 4.6505
R14983 VDD.n4429 VDD.n4428 4.6505
R14984 VDD.n4437 VDD.n4423 4.6505
R14985 VDD.n4426 VDD.n4425 4.6505
R14986 VDD.n4428 VDD.n4427 4.6505
R14987 VDD.n4713 VDD.n4712 4.6505
R14988 VDD.n4734 VDD.n4733 4.6505
R14989 VDD.n4735 VDD.n4730 4.6505
R14990 VDD.n4697 VDD.n4682 4.6505
R14991 VDD.n4697 VDD.n4696 4.6505
R14992 VDD.n4692 VDD.n4691 4.6505
R14993 VDD.n4694 VDD.n4692 4.6505
R14994 VDD.n4690 VDD.n4681 4.6505
R14995 VDD.n4688 VDD.n4684 4.6505
R14996 VDD.n4687 VDD.n4686 4.6505
R14997 VDD.n4695 VDD.n4681 4.6505
R14998 VDD.n4684 VDD.n4683 4.6505
R14999 VDD.n4686 VDD.n4685 4.6505
R15000 VDD.n4971 VDD.n4970 4.6505
R15001 VDD.n4992 VDD.n4991 4.6505
R15002 VDD.n4993 VDD.n4988 4.6505
R15003 VDD.n4955 VDD.n4940 4.6505
R15004 VDD.n4955 VDD.n4954 4.6505
R15005 VDD.n4950 VDD.n4949 4.6505
R15006 VDD.n4952 VDD.n4950 4.6505
R15007 VDD.n4948 VDD.n4939 4.6505
R15008 VDD.n4946 VDD.n4942 4.6505
R15009 VDD.n4945 VDD.n4944 4.6505
R15010 VDD.n4953 VDD.n4939 4.6505
R15011 VDD.n4942 VDD.n4941 4.6505
R15012 VDD.n4944 VDD.n4943 4.6505
R15013 VDD.n5229 VDD.n5228 4.6505
R15014 VDD.n5250 VDD.n5249 4.6505
R15015 VDD.n5251 VDD.n5246 4.6505
R15016 VDD.n5213 VDD.n5198 4.6505
R15017 VDD.n5213 VDD.n5212 4.6505
R15018 VDD.n5208 VDD.n5207 4.6505
R15019 VDD.n5210 VDD.n5208 4.6505
R15020 VDD.n5206 VDD.n5197 4.6505
R15021 VDD.n5204 VDD.n5200 4.6505
R15022 VDD.n5203 VDD.n5202 4.6505
R15023 VDD.n5211 VDD.n5197 4.6505
R15024 VDD.n5200 VDD.n5199 4.6505
R15025 VDD.n5202 VDD.n5201 4.6505
R15026 VDD.n12 VDD.n11 4.6505
R15027 VDD.n14 VDD.n13 4.6505
R15028 VDD.n16 VDD.n8 4.6505
R15029 VDD.n4 VDD.n2 4.6505
R15030 VDD.n23 VDD.n22 4.6505
R15031 VDD.n15 VDD.n6 4.6505
R15032 VDD.n18 VDD.n17 4.6505
R15033 VDD.n21 VDD.n20 4.6505
R15034 VDD.n30 VDD.n29 4.6505
R15035 VDD.n689 VDD.n524 4.6505
R15036 VDD.n697 VDD.n523 4.6505
R15037 VDD.n698 VDD.n522 4.6505
R15038 VDD.n744 VDD.n520 4.6505
R15039 VDD.n745 VDD.n519 4.6505
R15040 VDD.n791 VDD.n517 4.6505
R15041 VDD.n792 VDD.n516 4.6505
R15042 VDD.n622 VDD.n621 4.6505
R15043 VDD.n620 VDD.n619 4.6505
R15044 VDD.n551 VDD.n542 4.6505
R15045 VDD.n552 VDD.n541 4.6505
R15046 VDD.n676 VDD.n675 4.6505
R15047 VDD.n678 VDD.n677 4.6505
R15048 VDD.n680 VDD.n679 4.6505
R15049 VDD.n682 VDD.n681 4.6505
R15050 VDD.n685 VDD.n684 4.6505
R15051 VDD.n691 VDD.n690 4.6505
R15052 VDD.n694 VDD.n693 4.6505
R15053 VDD.n696 VDD.n695 4.6505
R15054 VDD.n700 VDD.n699 4.6505
R15055 VDD.n704 VDD.n703 4.6505
R15056 VDD.n706 VDD.n705 4.6505
R15057 VDD.n710 VDD.n709 4.6505
R15058 VDD.n712 VDD.n711 4.6505
R15059 VDD.n716 VDD.n715 4.6505
R15060 VDD.n718 VDD.n717 4.6505
R15061 VDD.n722 VDD.n721 4.6505
R15062 VDD.n726 VDD.n725 4.6505
R15063 VDD.n728 VDD.n727 4.6505
R15064 VDD.n732 VDD.n731 4.6505
R15065 VDD.n735 VDD.n734 4.6505
R15066 VDD.n740 VDD.n739 4.6505
R15067 VDD.n743 VDD.n742 4.6505
R15068 VDD.n747 VDD.n746 4.6505
R15069 VDD.n751 VDD.n750 4.6505
R15070 VDD.n753 VDD.n752 4.6505
R15071 VDD.n757 VDD.n756 4.6505
R15072 VDD.n759 VDD.n758 4.6505
R15073 VDD.n763 VDD.n762 4.6505
R15074 VDD.n765 VDD.n764 4.6505
R15075 VDD.n769 VDD.n768 4.6505
R15076 VDD.n773 VDD.n772 4.6505
R15077 VDD.n775 VDD.n774 4.6505
R15078 VDD.n780 VDD.n779 4.6505
R15079 VDD.n783 VDD.n782 4.6505
R15080 VDD.n788 VDD.n787 4.6505
R15081 VDD.n790 VDD.n789 4.6505
R15082 VDD.n515 VDD.n514 4.6505
R15083 VDD.n641 VDD.n640 4.6505
R15084 VDD.n643 VDD.n642 4.6505
R15085 VDD.n647 VDD.n646 4.6505
R15086 VDD.n649 VDD.n648 4.6505
R15087 VDD.n653 VDD.n652 4.6505
R15088 VDD.n655 VDD.n654 4.6505
R15089 VDD.n659 VDD.n658 4.6505
R15090 VDD.n664 VDD.n663 4.6505
R15091 VDD.n637 VDD.n636 4.6505
R15092 VDD.n634 VDD.n633 4.6505
R15093 VDD.n630 VDD.n629 4.6505
R15094 VDD.n628 VDD.n627 4.6505
R15095 VDD.n624 VDD.n623 4.6505
R15096 VDD.n618 VDD.n617 4.6505
R15097 VDD.n616 VDD.n615 4.6505
R15098 VDD.n612 VDD.n611 4.6505
R15099 VDD.n610 VDD.n609 4.6505
R15100 VDD.n606 VDD.n605 4.6505
R15101 VDD.n604 VDD.n603 4.6505
R15102 VDD.n600 VDD.n599 4.6505
R15103 VDD.n598 VDD.n597 4.6505
R15104 VDD.n594 VDD.n593 4.6505
R15105 VDD.n589 VDD.n588 4.6505
R15106 VDD.n528 VDD.n527 4.6505
R15107 VDD.n544 VDD.n543 4.6505
R15108 VDD.n548 VDD.n547 4.6505
R15109 VDD.n550 VDD.n549 4.6505
R15110 VDD.n554 VDD.n553 4.6505
R15111 VDD.n558 VDD.n557 4.6505
R15112 VDD.n560 VDD.n559 4.6505
R15113 VDD.n564 VDD.n563 4.6505
R15114 VDD.n566 VDD.n565 4.6505
R15115 VDD.n570 VDD.n569 4.6505
R15116 VDD.n572 VDD.n571 4.6505
R15117 VDD.n576 VDD.n575 4.6505
R15118 VDD.n581 VDD.n580 4.6505
R15119 VDD.n540 VDD.n539 4.6505
R15120 VDD.n537 VDD.n536 4.6505
R15121 VDD.n533 VDD.n532 4.6505
R15122 VDD.n474 VDD.n473 4.6505
R15123 VDD.n480 VDD.n472 4.6505
R15124 VDD.n480 VDD.n470 4.6505
R15125 VDD.n479 VDD.n478 4.6505
R15126 VDD.n485 VDD.n483 4.6505
R15127 VDD.n486 VDD.n469 4.6505
R15128 VDD.n467 VDD.n466 4.6505
R15129 VDD.n491 VDD.n490 4.6505
R15130 VDD.n493 VDD.n492 4.6505
R15131 VDD.n497 VDD.n496 4.6505
R15132 VDD.n499 VDD.n498 4.6505
R15133 VDD.n501 VDD.n500 4.6505
R15134 VDD.n503 VDD.n502 4.6505
R15135 VDD.n505 VDD.n504 4.6505
R15136 VDD.n507 VDD.n506 4.6505
R15137 VDD.n485 VDD.n484 4.6505
R15138 VDD.n487 VDD.n486 4.6505
R15139 VDD.n447 VDD.n446 4.6505
R15140 VDD.n451 VDD.n444 4.6505
R15141 VDD.n450 VDD.n448 4.6505
R15142 VDD.n454 VDD.n452 4.6505
R15143 VDD.n457 VDD.n455 4.6505
R15144 VDD.n447 VDD.n445 4.6505
R15145 VDD.n450 VDD.n449 4.6505
R15146 VDD.n451 VDD.n442 4.6505
R15147 VDD.n454 VDD.n453 4.6505
R15148 VDD.n457 VDD.n456 4.6505
R15149 VDD.n458 VDD.n440 4.6505
R15150 VDD.n415 VDD.n410 4.6505
R15151 VDD.n417 VDD.n409 4.6505
R15152 VDD.n415 VDD.n414 4.6505
R15153 VDD.n417 VDD.n416 4.6505
R15154 VDD.n421 VDD.n420 4.6505
R15155 VDD.n426 VDD.n425 4.6505
R15156 VDD.n428 VDD.n427 4.6505
R15157 VDD.n430 VDD.n429 4.6505
R15158 VDD.n432 VDD.n431 4.6505
R15159 VDD.n434 VDD.n433 4.6505
R15160 VDD.n396 VDD.n392 4.6505
R15161 VDD.n398 VDD.n391 4.6505
R15162 VDD.n398 VDD.n397 4.6505
R15163 VDD.n400 VDD.n399 4.6505
R15164 VDD.n72 VDD.n71 4.6505
R15165 VDD.n78 VDD.n70 4.6505
R15166 VDD.n78 VDD.n68 4.6505
R15167 VDD.n77 VDD.n76 4.6505
R15168 VDD.n83 VDD.n81 4.6505
R15169 VDD.n84 VDD.n67 4.6505
R15170 VDD.n65 VDD.n64 4.6505
R15171 VDD.n89 VDD.n88 4.6505
R15172 VDD.n91 VDD.n90 4.6505
R15173 VDD.n95 VDD.n94 4.6505
R15174 VDD.n97 VDD.n96 4.6505
R15175 VDD.n99 VDD.n98 4.6505
R15176 VDD.n101 VDD.n100 4.6505
R15177 VDD.n103 VDD.n102 4.6505
R15178 VDD.n105 VDD.n104 4.6505
R15179 VDD.n83 VDD.n82 4.6505
R15180 VDD.n85 VDD.n84 4.6505
R15181 VDD.n44 VDD.n43 4.6505
R15182 VDD.n48 VDD.n41 4.6505
R15183 VDD.n47 VDD.n45 4.6505
R15184 VDD.n51 VDD.n49 4.6505
R15185 VDD.n54 VDD.n52 4.6505
R15186 VDD.n44 VDD.n42 4.6505
R15187 VDD.n47 VDD.n46 4.6505
R15188 VDD.n48 VDD.n39 4.6505
R15189 VDD.n51 VDD.n50 4.6505
R15190 VDD.n54 VDD.n53 4.6505
R15191 VDD.n55 VDD.n37 4.6505
R15192 VDD.n1156 VDD.n1155 4.6505
R15193 VDD.n1158 VDD.n1157 4.6505
R15194 VDD.n1160 VDD.n1152 4.6505
R15195 VDD.n1148 VDD.n1146 4.6505
R15196 VDD.n1167 VDD.n1166 4.6505
R15197 VDD.n1159 VDD.n1150 4.6505
R15198 VDD.n1162 VDD.n1161 4.6505
R15199 VDD.n1165 VDD.n1164 4.6505
R15200 VDD.n1174 VDD.n1173 4.6505
R15201 VDD.n1573 VDD.n1568 4.6505
R15202 VDD.n1575 VDD.n1567 4.6505
R15203 VDD.n1573 VDD.n1572 4.6505
R15204 VDD.n1575 VDD.n1574 4.6505
R15205 VDD.n1579 VDD.n1578 4.6505
R15206 VDD.n1584 VDD.n1583 4.6505
R15207 VDD.n1586 VDD.n1585 4.6505
R15208 VDD.n1588 VDD.n1587 4.6505
R15209 VDD.n1590 VDD.n1589 4.6505
R15210 VDD.n1592 VDD.n1591 4.6505
R15211 VDD.n1554 VDD.n1550 4.6505
R15212 VDD.n1556 VDD.n1549 4.6505
R15213 VDD.n1556 VDD.n1555 4.6505
R15214 VDD.n1558 VDD.n1557 4.6505
R15215 VDD.n851 VDD.n850 4.6505
R15216 VDD.n849 VDD.n848 4.6505
R15217 VDD.n847 VDD.n846 4.6505
R15218 VDD.n845 VDD.n844 4.6505
R15219 VDD.n843 VDD.n842 4.6505
R15220 VDD.n841 VDD.n840 4.6505
R15221 VDD.n839 VDD.n838 4.6505
R15222 VDD.n837 VDD.n836 4.6505
R15223 VDD.n835 VDD.n834 4.6505
R15224 VDD.n833 VDD.n832 4.6505
R15225 VDD.n831 VDD.n830 4.6505
R15226 VDD.n829 VDD.n828 4.6505
R15227 VDD.n808 VDD.n804 4.6505
R15228 VDD.n812 VDD.n802 4.6505
R15229 VDD.n818 VDD.n799 4.6505
R15230 VDD.n817 VDD.n816 4.6505
R15231 VDD.n815 VDD.n801 4.6505
R15232 VDD.n814 VDD.n813 4.6505
R15233 VDD.n811 VDD.n810 4.6505
R15234 VDD.n1546 VDD.n1545 4.6505
R15235 VDD.n1039 VDD.n874 4.6505
R15236 VDD.n1047 VDD.n873 4.6505
R15237 VDD.n1048 VDD.n872 4.6505
R15238 VDD.n1094 VDD.n870 4.6505
R15239 VDD.n1095 VDD.n869 4.6505
R15240 VDD.n1141 VDD.n867 4.6505
R15241 VDD.n1142 VDD.n866 4.6505
R15242 VDD.n972 VDD.n971 4.6505
R15243 VDD.n970 VDD.n969 4.6505
R15244 VDD.n901 VDD.n892 4.6505
R15245 VDD.n902 VDD.n891 4.6505
R15246 VDD.n1026 VDD.n1025 4.6505
R15247 VDD.n1028 VDD.n1027 4.6505
R15248 VDD.n1030 VDD.n1029 4.6505
R15249 VDD.n1032 VDD.n1031 4.6505
R15250 VDD.n1035 VDD.n1034 4.6505
R15251 VDD.n1041 VDD.n1040 4.6505
R15252 VDD.n1044 VDD.n1043 4.6505
R15253 VDD.n1046 VDD.n1045 4.6505
R15254 VDD.n1050 VDD.n1049 4.6505
R15255 VDD.n1054 VDD.n1053 4.6505
R15256 VDD.n1056 VDD.n1055 4.6505
R15257 VDD.n1060 VDD.n1059 4.6505
R15258 VDD.n1062 VDD.n1061 4.6505
R15259 VDD.n1066 VDD.n1065 4.6505
R15260 VDD.n1068 VDD.n1067 4.6505
R15261 VDD.n1072 VDD.n1071 4.6505
R15262 VDD.n1076 VDD.n1075 4.6505
R15263 VDD.n1078 VDD.n1077 4.6505
R15264 VDD.n1082 VDD.n1081 4.6505
R15265 VDD.n1085 VDD.n1084 4.6505
R15266 VDD.n1090 VDD.n1089 4.6505
R15267 VDD.n1093 VDD.n1092 4.6505
R15268 VDD.n1097 VDD.n1096 4.6505
R15269 VDD.n1101 VDD.n1100 4.6505
R15270 VDD.n1103 VDD.n1102 4.6505
R15271 VDD.n1107 VDD.n1106 4.6505
R15272 VDD.n1109 VDD.n1108 4.6505
R15273 VDD.n1113 VDD.n1112 4.6505
R15274 VDD.n1115 VDD.n1114 4.6505
R15275 VDD.n1119 VDD.n1118 4.6505
R15276 VDD.n1123 VDD.n1122 4.6505
R15277 VDD.n1125 VDD.n1124 4.6505
R15278 VDD.n1130 VDD.n1129 4.6505
R15279 VDD.n1133 VDD.n1132 4.6505
R15280 VDD.n1138 VDD.n1137 4.6505
R15281 VDD.n1140 VDD.n1139 4.6505
R15282 VDD.n865 VDD.n864 4.6505
R15283 VDD.n991 VDD.n990 4.6505
R15284 VDD.n993 VDD.n992 4.6505
R15285 VDD.n997 VDD.n996 4.6505
R15286 VDD.n999 VDD.n998 4.6505
R15287 VDD.n1003 VDD.n1002 4.6505
R15288 VDD.n1005 VDD.n1004 4.6505
R15289 VDD.n1009 VDD.n1008 4.6505
R15290 VDD.n1014 VDD.n1013 4.6505
R15291 VDD.n987 VDD.n986 4.6505
R15292 VDD.n984 VDD.n983 4.6505
R15293 VDD.n980 VDD.n979 4.6505
R15294 VDD.n978 VDD.n977 4.6505
R15295 VDD.n974 VDD.n973 4.6505
R15296 VDD.n968 VDD.n967 4.6505
R15297 VDD.n966 VDD.n965 4.6505
R15298 VDD.n962 VDD.n961 4.6505
R15299 VDD.n960 VDD.n959 4.6505
R15300 VDD.n956 VDD.n955 4.6505
R15301 VDD.n954 VDD.n953 4.6505
R15302 VDD.n950 VDD.n949 4.6505
R15303 VDD.n948 VDD.n947 4.6505
R15304 VDD.n944 VDD.n943 4.6505
R15305 VDD.n939 VDD.n938 4.6505
R15306 VDD.n878 VDD.n877 4.6505
R15307 VDD.n894 VDD.n893 4.6505
R15308 VDD.n898 VDD.n897 4.6505
R15309 VDD.n900 VDD.n899 4.6505
R15310 VDD.n904 VDD.n903 4.6505
R15311 VDD.n908 VDD.n907 4.6505
R15312 VDD.n910 VDD.n909 4.6505
R15313 VDD.n914 VDD.n913 4.6505
R15314 VDD.n916 VDD.n915 4.6505
R15315 VDD.n920 VDD.n919 4.6505
R15316 VDD.n922 VDD.n921 4.6505
R15317 VDD.n926 VDD.n925 4.6505
R15318 VDD.n931 VDD.n930 4.6505
R15319 VDD.n890 VDD.n889 4.6505
R15320 VDD.n887 VDD.n886 4.6505
R15321 VDD.n883 VDD.n882 4.6505
R15322 VDD.n284 VDD.n123 4.6505
R15323 VDD.n292 VDD.n122 4.6505
R15324 VDD.n293 VDD.n121 4.6505
R15325 VDD.n339 VDD.n119 4.6505
R15326 VDD.n340 VDD.n118 4.6505
R15327 VDD.n386 VDD.n116 4.6505
R15328 VDD.n387 VDD.n115 4.6505
R15329 VDD.n221 VDD.n220 4.6505
R15330 VDD.n219 VDD.n218 4.6505
R15331 VDD.n150 VDD.n141 4.6505
R15332 VDD.n151 VDD.n140 4.6505
R15333 VDD.n271 VDD.n270 4.6505
R15334 VDD.n273 VDD.n272 4.6505
R15335 VDD.n275 VDD.n274 4.6505
R15336 VDD.n277 VDD.n276 4.6505
R15337 VDD.n280 VDD.n279 4.6505
R15338 VDD.n286 VDD.n285 4.6505
R15339 VDD.n289 VDD.n288 4.6505
R15340 VDD.n291 VDD.n290 4.6505
R15341 VDD.n295 VDD.n294 4.6505
R15342 VDD.n299 VDD.n298 4.6505
R15343 VDD.n301 VDD.n300 4.6505
R15344 VDD.n305 VDD.n304 4.6505
R15345 VDD.n307 VDD.n306 4.6505
R15346 VDD.n311 VDD.n310 4.6505
R15347 VDD.n313 VDD.n312 4.6505
R15348 VDD.n317 VDD.n316 4.6505
R15349 VDD.n321 VDD.n320 4.6505
R15350 VDD.n323 VDD.n322 4.6505
R15351 VDD.n327 VDD.n326 4.6505
R15352 VDD.n330 VDD.n329 4.6505
R15353 VDD.n335 VDD.n334 4.6505
R15354 VDD.n338 VDD.n337 4.6505
R15355 VDD.n342 VDD.n341 4.6505
R15356 VDD.n346 VDD.n345 4.6505
R15357 VDD.n348 VDD.n347 4.6505
R15358 VDD.n352 VDD.n351 4.6505
R15359 VDD.n354 VDD.n353 4.6505
R15360 VDD.n358 VDD.n357 4.6505
R15361 VDD.n360 VDD.n359 4.6505
R15362 VDD.n364 VDD.n363 4.6505
R15363 VDD.n368 VDD.n367 4.6505
R15364 VDD.n370 VDD.n369 4.6505
R15365 VDD.n375 VDD.n374 4.6505
R15366 VDD.n378 VDD.n377 4.6505
R15367 VDD.n383 VDD.n382 4.6505
R15368 VDD.n385 VDD.n384 4.6505
R15369 VDD.n389 VDD.n388 4.6505
R15370 VDD.n114 VDD.n113 4.6505
R15371 VDD.n238 VDD.n237 4.6505
R15372 VDD.n242 VDD.n241 4.6505
R15373 VDD.n244 VDD.n243 4.6505
R15374 VDD.n248 VDD.n247 4.6505
R15375 VDD.n250 VDD.n249 4.6505
R15376 VDD.n254 VDD.n253 4.6505
R15377 VDD.n259 VDD.n258 4.6505
R15378 VDD.n236 VDD.n235 4.6505
R15379 VDD.n233 VDD.n232 4.6505
R15380 VDD.n229 VDD.n228 4.6505
R15381 VDD.n227 VDD.n226 4.6505
R15382 VDD.n223 VDD.n222 4.6505
R15383 VDD.n217 VDD.n216 4.6505
R15384 VDD.n215 VDD.n214 4.6505
R15385 VDD.n211 VDD.n210 4.6505
R15386 VDD.n209 VDD.n208 4.6505
R15387 VDD.n205 VDD.n204 4.6505
R15388 VDD.n203 VDD.n202 4.6505
R15389 VDD.n199 VDD.n198 4.6505
R15390 VDD.n197 VDD.n196 4.6505
R15391 VDD.n193 VDD.n192 4.6505
R15392 VDD.n188 VDD.n187 4.6505
R15393 VDD.n127 VDD.n126 4.6505
R15394 VDD.n143 VDD.n142 4.6505
R15395 VDD.n147 VDD.n146 4.6505
R15396 VDD.n149 VDD.n148 4.6505
R15397 VDD.n153 VDD.n152 4.6505
R15398 VDD.n157 VDD.n156 4.6505
R15399 VDD.n159 VDD.n158 4.6505
R15400 VDD.n163 VDD.n162 4.6505
R15401 VDD.n165 VDD.n164 4.6505
R15402 VDD.n169 VDD.n168 4.6505
R15403 VDD.n171 VDD.n170 4.6505
R15404 VDD.n175 VDD.n174 4.6505
R15405 VDD.n180 VDD.n179 4.6505
R15406 VDD.n139 VDD.n138 4.6505
R15407 VDD.n136 VDD.n135 4.6505
R15408 VDD.n132 VDD.n131 4.6505
R15409 VDD.n1358 VDD.n1357 4.6505
R15410 VDD.n1349 VDD.n1348 4.6505
R15411 VDD.n1347 VDD.n1346 4.6505
R15412 VDD.n1343 VDD.n1342 4.6505
R15413 VDD.n1341 VDD.n1340 4.6505
R15414 VDD.n1314 VDD.n1313 4.6505
R15415 VDD.n1365 VDD.n1364 4.6505
R15416 VDD.n1368 VDD.n1367 4.6505
R15417 VDD.n1356 VDD.n1355 4.6505
R15418 VDD.n1354 VDD.n1353 4.6505
R15419 VDD.n1351 VDD.n1350 4.6505
R15420 VDD.n1376 VDD.n1375 4.6505
R15421 VDD.n1381 VDD.n1380 4.6505
R15422 VDD.n1383 VDD.n1382 4.6505
R15423 VDD.n1387 VDD.n1386 4.6505
R15424 VDD.n1389 VDD.n1388 4.6505
R15425 VDD.n1393 VDD.n1392 4.6505
R15426 VDD.n1396 VDD.n1395 4.6505
R15427 VDD.n1405 VDD.n1404 4.6505
R15428 VDD.n1410 VDD.n1409 4.6505
R15429 VDD.n1412 VDD.n1411 4.6505
R15430 VDD.n1416 VDD.n1415 4.6505
R15431 VDD.n1418 VDD.n1417 4.6505
R15432 VDD.n1422 VDD.n1421 4.6505
R15433 VDD.n1425 VDD.n1424 4.6505
R15434 VDD.n1339 VDD.n1338 4.6505
R15435 VDD.n1337 VDD.n1336 4.6505
R15436 VDD.n1333 VDD.n1332 4.6505
R15437 VDD.n1331 VDD.n1330 4.6505
R15438 VDD.n1327 VDD.n1326 4.6505
R15439 VDD.n1324 VDD.n1323 4.6505
R15440 VDD.n1433 VDD.n1432 4.6505
R15441 VDD.n1437 VDD.n1436 4.6505
R15442 VDD.n1441 VDD.n1440 4.6505
R15443 VDD.n1443 VDD.n1442 4.6505
R15444 VDD.n1447 VDD.n1446 4.6505
R15445 VDD.n1449 VDD.n1448 4.6505
R15446 VDD.n1453 VDD.n1452 4.6505
R15447 VDD.n1317 VDD.n1316 4.6505
R15448 VDD.n1312 VDD.n1311 4.6505
R15449 VDD.n1310 VDD.n1309 4.6505
R15450 VDD.n1308 VDD.n1307 4.6505
R15451 VDD.n1527 VDD.n1258 4.6505
R15452 VDD.n1529 VDD.n1528 4.6505
R15453 VDD.n1533 VDD.n1532 4.6505
R15454 VDD.n1537 VDD.n1536 4.6505
R15455 VDD.n1539 VDD.n1538 4.6505
R15456 VDD.n1255 VDD.n1254 4.6505
R15457 VDD.n1251 VDD.n1250 4.6505
R15458 VDD.n1286 VDD.n1263 4.6505
R15459 VDD.n1460 VDD.n1262 4.6505
R15460 VDD.n1261 VDD.n1260 4.6505
R15461 VDD.n1510 VDD.n1259 4.6505
R15462 VDD.n1283 VDD.n1266 4.6505
R15463 VDD.n1285 VDD.n1284 4.6505
R15464 VDD.n1463 VDD.n1462 4.6505
R15465 VDD.n1467 VDD.n1466 4.6505
R15466 VDD.n1469 VDD.n1468 4.6505
R15467 VDD.n1473 VDD.n1472 4.6505
R15468 VDD.n1475 VDD.n1474 4.6505
R15469 VDD.n1479 VDD.n1478 4.6505
R15470 VDD.n1481 VDD.n1480 4.6505
R15471 VDD.n1485 VDD.n1484 4.6505
R15472 VDD.n1489 VDD.n1488 4.6505
R15473 VDD.n1491 VDD.n1490 4.6505
R15474 VDD.n1495 VDD.n1494 4.6505
R15475 VDD.n1497 VDD.n1496 4.6505
R15476 VDD.n1501 VDD.n1500 4.6505
R15477 VDD.n1503 VDD.n1502 4.6505
R15478 VDD.n1513 VDD.n1512 4.6505
R15479 VDD.n1517 VDD.n1516 4.6505
R15480 VDD.n1519 VDD.n1518 4.6505
R15481 VDD.n1523 VDD.n1522 4.6505
R15482 VDD.n1525 VDD.n1524 4.6505
R15483 VDD.n1303 VDD.n1302 4.6505
R15484 VDD.n1301 VDD.n1300 4.6505
R15485 VDD.n1297 VDD.n1296 4.6505
R15486 VDD.n1295 VDD.n1294 4.6505
R15487 VDD.n1291 VDD.n1290 4.6505
R15488 VDD.n1270 VDD.n1269 4.6505
R15489 VDD.n1274 VDD.n1273 4.6505
R15490 VDD.n1276 VDD.n1275 4.6505
R15491 VDD.n1280 VDD.n1279 4.6505
R15492 VDD.n1282 VDD.n1281 4.6505
R15493 VDD.n1234 VDD.n1233 4.6505
R15494 VDD.n1232 VDD.n1231 4.6505
R15495 VDD.n1230 VDD.n1229 4.6505
R15496 VDD.n1228 VDD.n1227 4.6505
R15497 VDD.n1226 VDD.n1225 4.6505
R15498 VDD.n1224 VDD.n1223 4.6505
R15499 VDD.n1222 VDD.n1221 4.6505
R15500 VDD.n1220 VDD.n1219 4.6505
R15501 VDD.n1218 VDD.n1217 4.6505
R15502 VDD.n1216 VDD.n1215 4.6505
R15503 VDD.n1214 VDD.n1213 4.6505
R15504 VDD.n1212 VDD.n1211 4.6505
R15505 VDD.n1191 VDD.n1187 4.6505
R15506 VDD.n1195 VDD.n1185 4.6505
R15507 VDD.n1201 VDD.n1182 4.6505
R15508 VDD.n1200 VDD.n1199 4.6505
R15509 VDD.n1198 VDD.n1184 4.6505
R15510 VDD.n1197 VDD.n1196 4.6505
R15511 VDD.n1194 VDD.n1193 4.6505
R15512 VDD.n1653 VDD.n1646 4.61128
R15513 VDD.n1946 VDD.n1943 4.58799
R15514 VDD.n1751 VDD.n1721 4.5005
R15515 VDD.n1751 VDD.n1716 4.5005
R15516 VDD.n1751 VDD.n1750 4.5005
R15517 VDD.n1777 VDD.n1776 4.5005
R15518 VDD.n1800 VDD.n1779 4.5005
R15519 VDD.n1800 VDD.n1799 4.5005
R15520 VDD.n1797 VDD.n1779 4.5005
R15521 VDD.n2100 VDD.n2070 4.5005
R15522 VDD.n2100 VDD.n2065 4.5005
R15523 VDD.n2100 VDD.n2099 4.5005
R15524 VDD.n1985 VDD.n1984 4.5005
R15525 VDD.n2008 VDD.n1987 4.5005
R15526 VDD.n2008 VDD.n2007 4.5005
R15527 VDD.n2005 VDD.n1987 4.5005
R15528 VDD.n2330 VDD.n2300 4.5005
R15529 VDD.n2330 VDD.n2295 4.5005
R15530 VDD.n2330 VDD.n2329 4.5005
R15531 VDD.n2356 VDD.n2355 4.5005
R15532 VDD.n2379 VDD.n2358 4.5005
R15533 VDD.n2379 VDD.n2378 4.5005
R15534 VDD.n2376 VDD.n2358 4.5005
R15535 VDD.n2588 VDD.n2558 4.5005
R15536 VDD.n2588 VDD.n2553 4.5005
R15537 VDD.n2588 VDD.n2587 4.5005
R15538 VDD.n2614 VDD.n2613 4.5005
R15539 VDD.n2637 VDD.n2616 4.5005
R15540 VDD.n2637 VDD.n2636 4.5005
R15541 VDD.n2634 VDD.n2616 4.5005
R15542 VDD.n2846 VDD.n2816 4.5005
R15543 VDD.n2846 VDD.n2811 4.5005
R15544 VDD.n2846 VDD.n2845 4.5005
R15545 VDD.n2872 VDD.n2871 4.5005
R15546 VDD.n2895 VDD.n2874 4.5005
R15547 VDD.n2895 VDD.n2894 4.5005
R15548 VDD.n2892 VDD.n2874 4.5005
R15549 VDD.n3104 VDD.n3074 4.5005
R15550 VDD.n3104 VDD.n3069 4.5005
R15551 VDD.n3104 VDD.n3103 4.5005
R15552 VDD.n3130 VDD.n3129 4.5005
R15553 VDD.n3153 VDD.n3132 4.5005
R15554 VDD.n3153 VDD.n3152 4.5005
R15555 VDD.n3150 VDD.n3132 4.5005
R15556 VDD.n3362 VDD.n3332 4.5005
R15557 VDD.n3362 VDD.n3327 4.5005
R15558 VDD.n3362 VDD.n3361 4.5005
R15559 VDD.n3388 VDD.n3387 4.5005
R15560 VDD.n3411 VDD.n3390 4.5005
R15561 VDD.n3411 VDD.n3410 4.5005
R15562 VDD.n3408 VDD.n3390 4.5005
R15563 VDD.n5685 VDD.n5655 4.5005
R15564 VDD.n5685 VDD.n5650 4.5005
R15565 VDD.n5685 VDD.n5684 4.5005
R15566 VDD.n5711 VDD.n5710 4.5005
R15567 VDD.n5734 VDD.n5713 4.5005
R15568 VDD.n5734 VDD.n5733 4.5005
R15569 VDD.n5731 VDD.n5713 4.5005
R15570 VDD.n5431 VDD.n5401 4.5005
R15571 VDD.n5431 VDD.n5396 4.5005
R15572 VDD.n5431 VDD.n5430 4.5005
R15573 VDD.n5457 VDD.n5456 4.5005
R15574 VDD.n5480 VDD.n5459 4.5005
R15575 VDD.n5480 VDD.n5479 4.5005
R15576 VDD.n5477 VDD.n5459 4.5005
R15577 VDD.n3620 VDD.n3590 4.5005
R15578 VDD.n3620 VDD.n3585 4.5005
R15579 VDD.n3620 VDD.n3619 4.5005
R15580 VDD.n3646 VDD.n3645 4.5005
R15581 VDD.n3669 VDD.n3648 4.5005
R15582 VDD.n3669 VDD.n3668 4.5005
R15583 VDD.n3666 VDD.n3648 4.5005
R15584 VDD.n3878 VDD.n3848 4.5005
R15585 VDD.n3878 VDD.n3843 4.5005
R15586 VDD.n3878 VDD.n3877 4.5005
R15587 VDD.n3904 VDD.n3903 4.5005
R15588 VDD.n3927 VDD.n3906 4.5005
R15589 VDD.n3927 VDD.n3926 4.5005
R15590 VDD.n3924 VDD.n3906 4.5005
R15591 VDD.n4136 VDD.n4106 4.5005
R15592 VDD.n4136 VDD.n4101 4.5005
R15593 VDD.n4136 VDD.n4135 4.5005
R15594 VDD.n4162 VDD.n4161 4.5005
R15595 VDD.n4185 VDD.n4164 4.5005
R15596 VDD.n4185 VDD.n4184 4.5005
R15597 VDD.n4182 VDD.n4164 4.5005
R15598 VDD.n4394 VDD.n4364 4.5005
R15599 VDD.n4394 VDD.n4359 4.5005
R15600 VDD.n4394 VDD.n4393 4.5005
R15601 VDD.n4420 VDD.n4419 4.5005
R15602 VDD.n4443 VDD.n4422 4.5005
R15603 VDD.n4443 VDD.n4442 4.5005
R15604 VDD.n4440 VDD.n4422 4.5005
R15605 VDD.n4652 VDD.n4622 4.5005
R15606 VDD.n4652 VDD.n4617 4.5005
R15607 VDD.n4652 VDD.n4651 4.5005
R15608 VDD.n4678 VDD.n4677 4.5005
R15609 VDD.n4701 VDD.n4680 4.5005
R15610 VDD.n4701 VDD.n4700 4.5005
R15611 VDD.n4698 VDD.n4680 4.5005
R15612 VDD.n4910 VDD.n4880 4.5005
R15613 VDD.n4910 VDD.n4875 4.5005
R15614 VDD.n4910 VDD.n4909 4.5005
R15615 VDD.n4936 VDD.n4935 4.5005
R15616 VDD.n4959 VDD.n4938 4.5005
R15617 VDD.n4959 VDD.n4958 4.5005
R15618 VDD.n4956 VDD.n4938 4.5005
R15619 VDD.n5168 VDD.n5138 4.5005
R15620 VDD.n5168 VDD.n5133 4.5005
R15621 VDD.n5168 VDD.n5167 4.5005
R15622 VDD.n5194 VDD.n5193 4.5005
R15623 VDD.n5217 VDD.n5196 4.5005
R15624 VDD.n5217 VDD.n5216 4.5005
R15625 VDD.n5214 VDD.n5196 4.5005
R15626 VDD.n1249 VDD.n1248 4.45149
R15627 VDD.n531 VDD.n530 4.4514
R15628 VDD.n881 VDD.n880 4.4514
R15629 VDD.n130 VDD.n129 4.4514
R15630 VDD.n1649 VDD.n1648 4.43268
R15631 VDD.n1887 VDD.t506 4.35136
R15632 VDD.n1874 VDD.t493 4.35136
R15633 VDD.n2195 VDD.t594 4.35136
R15634 VDD.n2208 VDD.t1072 4.35136
R15635 VDD.n2453 VDD.t1379 4.35136
R15636 VDD.n2466 VDD.t1380 4.35136
R15637 VDD.n2711 VDD.t516 4.35136
R15638 VDD.n2724 VDD.t263 4.35136
R15639 VDD.n2969 VDD.t497 4.35136
R15640 VDD.n2982 VDD.t504 4.35136
R15641 VDD.n3227 VDD.t593 4.35136
R15642 VDD.n3240 VDD.t1022 4.35136
R15643 VDD.n3485 VDD.t522 4.35136
R15644 VDD.n3498 VDD.t523 4.35136
R15645 VDD.n5805 VDD.t517 4.35136
R15646 VDD.n5818 VDD.t518 4.35136
R15647 VDD.n5551 VDD.t417 4.35136
R15648 VDD.n5564 VDD.t418 4.35136
R15649 VDD.n3743 VDD.t1073 4.35136
R15650 VDD.n3756 VDD.t1074 4.35136
R15651 VDD.n4001 VDD.t1025 4.35136
R15652 VDD.n4014 VDD.t1382 4.35136
R15653 VDD.n4259 VDD.t260 4.35136
R15654 VDD.n4272 VDD.t261 4.35136
R15655 VDD.n4517 VDD.t495 4.35136
R15656 VDD.n4530 VDD.t496 4.35136
R15657 VDD.n4775 VDD.t1019 4.35136
R15658 VDD.n4788 VDD.t1020 4.35136
R15659 VDD.n5033 VDD.t529 4.35136
R15660 VDD.n5046 VDD.t530 4.35136
R15661 VDD.n5291 VDD.t515 4.35136
R15662 VDD.n5304 VDD.t513 4.35136
R15663 VDD.n1633 VDD 4.26717
R15664 VDD.n674 VDD.n673 4.14756
R15665 VDD.n1024 VDD.n1023 4.14756
R15666 VDD.n269 VDD.n268 4.14756
R15667 VDD.n466 VDD.n465 4.14168
R15668 VDD.n64 VDD.n63 4.14168
R15669 VDD.n805 VDD.n804 4.14168
R15670 VDD.n1188 VDD.n1187 4.14168
R15671 VDD.n489 VDD.n488 4.05611
R15672 VDD.n87 VDD.n86 4.05611
R15673 VDD.n25 VDD.n24 4.05569
R15674 VDD.n461 VDD.n460 4.05569
R15675 VDD.n58 VDD.n57 4.05569
R15676 VDD.n1169 VDD.n1168 4.05569
R15677 VDD.n1626 VDD.n1625 4.04261
R15678 VDD.n510 VDD.n509 4.01726
R15679 VDD.n437 VDD.n436 4.01726
R15680 VDD.n406 VDD.n405 4.01726
R15681 VDD.n108 VDD.n107 4.01726
R15682 VDD.n1595 VDD.n1594 4.01726
R15683 VDD.n1564 VDD.n1563 4.01726
R15684 VDD.n33 VDD.n32 4.01682
R15685 VDD.n1177 VDD.n1176 4.01682
R15686 VDD.n1815 VDD.n1814 3.96837
R15687 VDD.n2136 VDD.n2135 3.96837
R15688 VDD.n2394 VDD.n2393 3.96837
R15689 VDD.n2652 VDD.n2651 3.96837
R15690 VDD.n2910 VDD.n2909 3.96837
R15691 VDD.n3168 VDD.n3167 3.96837
R15692 VDD.n3426 VDD.n3425 3.96837
R15693 VDD.n5746 VDD.n5745 3.96837
R15694 VDD.n5492 VDD.n5491 3.96837
R15695 VDD.n3684 VDD.n3683 3.96837
R15696 VDD.n3942 VDD.n3941 3.96837
R15697 VDD.n4200 VDD.n4199 3.96837
R15698 VDD.n4458 VDD.n4457 3.96837
R15699 VDD.n4716 VDD.n4715 3.96837
R15700 VDD.n4974 VDD.n4973 3.96837
R15701 VDD.n5232 VDD.n5231 3.96837
R15702 VDD.n820 VDD.n819 3.96556
R15703 VDD.n1203 VDD.n1202 3.96556
R15704 VDD.n1638 VDD.n1637 3.88621
R15705 VDD.n1952 VDD.n1939 3.5871
R15706 VDD.n1694 VDD.n1683 3.52991
R15707 VDD.n2043 VDD.n2032 3.52991
R15708 VDD.n2273 VDD.n2262 3.52991
R15709 VDD.n2531 VDD.n2520 3.52991
R15710 VDD.n2789 VDD.n2778 3.52991
R15711 VDD.n3047 VDD.n3036 3.52991
R15712 VDD.n3305 VDD.n3294 3.52991
R15713 VDD.n5628 VDD.n5617 3.52991
R15714 VDD.n5374 VDD.n5363 3.52991
R15715 VDD.n3563 VDD.n3552 3.52991
R15716 VDD.n3821 VDD.n3810 3.52991
R15717 VDD.n4079 VDD.n4068 3.52991
R15718 VDD.n4337 VDD.n4326 3.52991
R15719 VDD.n4595 VDD.n4584 3.52991
R15720 VDD.n4853 VDD.n4842 3.52991
R15721 VDD.n5111 VDD.n5100 3.52991
R15722 VDD.n1608 VDD.n1607 3.46717
R15723 VDD.t1391 VDD.n669 3.39336
R15724 VDD.t47 VDD.n1019 3.39336
R15725 VDD.n263 VDD.t726 3.39336
R15726 VDD.n20 VDD.n19 3.38874
R15727 VDD.n496 VDD.n495 3.38874
R15728 VDD.n420 VDD.n419 3.38874
R15729 VDD.n94 VDD.n93 3.38874
R15730 VDD.n1164 VDD.n1163 3.38874
R15731 VDD.n1578 VDD.n1577 3.38874
R15732 VDD.n1980 VDD.n1922 3.1102
R15733 VDD.n1980 VDD.n1979 3.08146
R15734 VDD.n1701 VDD.n1700 3.03311
R15735 VDD.n2050 VDD.n2049 3.03311
R15736 VDD.n2280 VDD.n2279 3.03311
R15737 VDD.n2538 VDD.n2537 3.03311
R15738 VDD.n2796 VDD.n2795 3.03311
R15739 VDD.n3054 VDD.n3053 3.03311
R15740 VDD.n3312 VDD.n3311 3.03311
R15741 VDD.n5635 VDD.n5634 3.03311
R15742 VDD.n5381 VDD.n5380 3.03311
R15743 VDD.n3570 VDD.n3569 3.03311
R15744 VDD.n3828 VDD.n3827 3.03311
R15745 VDD.n4086 VDD.n4085 3.03311
R15746 VDD.n4344 VDD.n4343 3.03311
R15747 VDD.n4602 VDD.n4601 3.03311
R15748 VDD.n4860 VDD.n4859 3.03311
R15749 VDD.n5118 VDD.n5117 3.03311
R15750 VDD.n1609 VDD.n1608 3.03311
R15751 VDD VDD.n1622 3.02091
R15752 VDD.n1831 VDD 3.0005
R15753 VDD.n2152 VDD 3.0005
R15754 VDD.n2410 VDD 3.0005
R15755 VDD.n2668 VDD 3.0005
R15756 VDD.n2926 VDD 3.0005
R15757 VDD.n3184 VDD 3.0005
R15758 VDD.n3442 VDD 3.0005
R15759 VDD.n5762 VDD 3.0005
R15760 VDD.n5508 VDD 3.0005
R15761 VDD.n3700 VDD 3.0005
R15762 VDD.n3958 VDD 3.0005
R15763 VDD.n4216 VDD 3.0005
R15764 VDD.n4474 VDD 3.0005
R15765 VDD.n4732 VDD 3.0005
R15766 VDD.n4990 VDD 3.0005
R15767 VDD.n5248 VDD 3.0005
R15768 VDD.n1871 VDD.n1870 2.98717
R15769 VDD.n2192 VDD.n2191 2.98717
R15770 VDD.n2450 VDD.n2449 2.98717
R15771 VDD.n2708 VDD.n2707 2.98717
R15772 VDD.n2966 VDD.n2965 2.98717
R15773 VDD.n3224 VDD.n3223 2.98717
R15774 VDD.n3482 VDD.n3481 2.98717
R15775 VDD.n5802 VDD.n5801 2.98717
R15776 VDD.n5548 VDD.n5547 2.98717
R15777 VDD.n3740 VDD.n3739 2.98717
R15778 VDD.n3998 VDD.n3997 2.98717
R15779 VDD.n4256 VDD.n4255 2.98717
R15780 VDD.n4514 VDD.n4513 2.98717
R15781 VDD.n4772 VDD.n4771 2.98717
R15782 VDD.n5030 VDD.n5029 2.98717
R15783 VDD.n5288 VDD.n5287 2.98717
R15784 VDD.n1916 VDD.n1889 2.72837
R15785 VDD.n2237 VDD.n2210 2.72837
R15786 VDD.n2495 VDD.n2468 2.72837
R15787 VDD.n2753 VDD.n2726 2.72837
R15788 VDD.n3011 VDD.n2984 2.72837
R15789 VDD.n3269 VDD.n3242 2.72837
R15790 VDD.n3527 VDD.n3500 2.72837
R15791 VDD.n5847 VDD.n5820 2.72837
R15792 VDD.n5593 VDD.n5566 2.72837
R15793 VDD.n3785 VDD.n3758 2.72837
R15794 VDD.n4043 VDD.n4016 2.72837
R15795 VDD.n4301 VDD.n4274 2.72837
R15796 VDD.n4559 VDD.n4532 2.72837
R15797 VDD.n4817 VDD.n4790 2.72837
R15798 VDD.n5075 VDD.n5048 2.72837
R15799 VDD.n5333 VDD.n5306 2.72837
R15800 VDD.n477 VDD.n476 2.30978
R15801 VDD.n75 VDD.n74 2.30978
R15802 VDD.n1622 VDD.n1614 2.251
R15803 VDD.n1778 VDD.n1777 2.2278
R15804 VDD.n1986 VDD.n1985 2.2278
R15805 VDD.n2357 VDD.n2356 2.2278
R15806 VDD.n2615 VDD.n2614 2.2278
R15807 VDD.n2873 VDD.n2872 2.2278
R15808 VDD.n3131 VDD.n3130 2.2278
R15809 VDD.n3389 VDD.n3388 2.2278
R15810 VDD.n5712 VDD.n5711 2.2278
R15811 VDD.n5458 VDD.n5457 2.2278
R15812 VDD.n3647 VDD.n3646 2.2278
R15813 VDD.n3905 VDD.n3904 2.2278
R15814 VDD.n4163 VDD.n4162 2.2278
R15815 VDD.n4421 VDD.n4420 2.2278
R15816 VDD.n4679 VDD.n4678 2.2278
R15817 VDD.n4937 VDD.n4936 2.2278
R15818 VDD.n5195 VDD.n5194 2.2278
R15819 VDD VDD.n1633 2.13383
R15820 VDD.n1644 VDD 2.11184
R15821 VDD.n1655 VDD.n1642 1.59861
R15822 VDD.n1630 VDD 1.53093
R15823 VDD.n1981 VDD 1.52828
R15824 VDD.n1772 VDD.n1771 1.51475
R15825 VDD.n2121 VDD.n2120 1.51475
R15826 VDD.n2351 VDD.n2350 1.51475
R15827 VDD.n2609 VDD.n2608 1.51475
R15828 VDD.n2867 VDD.n2866 1.51475
R15829 VDD.n3125 VDD.n3124 1.51475
R15830 VDD.n3383 VDD.n3382 1.51475
R15831 VDD.n5706 VDD.n5705 1.51475
R15832 VDD.n5452 VDD.n5451 1.51475
R15833 VDD.n3641 VDD.n3640 1.51475
R15834 VDD.n3899 VDD.n3898 1.51475
R15835 VDD.n4157 VDD.n4156 1.51475
R15836 VDD.n4415 VDD.n4414 1.51475
R15837 VDD.n4673 VDD.n4672 1.51475
R15838 VDD.n4931 VDD.n4930 1.51475
R15839 VDD.n5189 VDD.n5188 1.51475
R15840 VDD.n1945 VDD.t1037 1.50409
R15841 VDD.n1924 VDD.t1027 1.50409
R15842 VDD.n1924 VDD.t1039 1.50409
R15843 VDD.n1918 VDD.n1917 1.49778
R15844 VDD.n2239 VDD.n2238 1.49778
R15845 VDD.n2497 VDD.n2496 1.49778
R15846 VDD.n2755 VDD.n2754 1.49778
R15847 VDD.n3013 VDD.n3012 1.49778
R15848 VDD.n3271 VDD.n3270 1.49778
R15849 VDD.n3529 VDD.n3528 1.49778
R15850 VDD.n5849 VDD.n5848 1.49778
R15851 VDD.n5595 VDD.n5594 1.49778
R15852 VDD.n3787 VDD.n3786 1.49778
R15853 VDD.n4045 VDD.n4044 1.49778
R15854 VDD.n4303 VDD.n4302 1.49778
R15855 VDD.n4561 VDD.n4560 1.49778
R15856 VDD.n4819 VDD.n4818 1.49778
R15857 VDD.n5077 VDD.n5076 1.49778
R15858 VDD.n5335 VDD.n5334 1.49778
R15859 VDD.n2013 VDD.n2012 1.47642
R15860 VDD.n1661 VDD.n1660 1.43354
R15861 VDD.n1740 VDD.n1729 1.42272
R15862 VDD.n2089 VDD.n2078 1.42272
R15863 VDD.n2319 VDD.n2308 1.42272
R15864 VDD.n2577 VDD.n2566 1.42272
R15865 VDD.n2835 VDD.n2824 1.42272
R15866 VDD.n3093 VDD.n3082 1.42272
R15867 VDD.n3351 VDD.n3340 1.42272
R15868 VDD.n5674 VDD.n5663 1.42272
R15869 VDD.n5420 VDD.n5409 1.42272
R15870 VDD.n3609 VDD.n3598 1.42272
R15871 VDD.n3867 VDD.n3856 1.42272
R15872 VDD.n4125 VDD.n4114 1.42272
R15873 VDD.n4383 VDD.n4372 1.42272
R15874 VDD.n4641 VDD.n4630 1.42272
R15875 VDD.n4899 VDD.n4888 1.42272
R15876 VDD.n5157 VDD.n5146 1.42272
R15877 VDD.n1663 VDD.n1662 1.39179
R15878 VDD.n1887 VDD.n1886 1.25748
R15879 VDD.n2208 VDD.n2207 1.25748
R15880 VDD.n2466 VDD.n2465 1.25748
R15881 VDD.n2724 VDD.n2723 1.25748
R15882 VDD.n2982 VDD.n2981 1.25748
R15883 VDD.n3240 VDD.n3239 1.25748
R15884 VDD.n3498 VDD.n3497 1.25748
R15885 VDD.n5818 VDD.n5817 1.25748
R15886 VDD.n5564 VDD.n5563 1.25748
R15887 VDD.n3756 VDD.n3755 1.25748
R15888 VDD.n4014 VDD.n4013 1.25748
R15889 VDD.n4272 VDD.n4271 1.25748
R15890 VDD.n4530 VDD.n4529 1.25748
R15891 VDD.n4788 VDD.n4787 1.25748
R15892 VDD.n5046 VDD.n5045 1.25748
R15893 VDD.n5304 VDD.n5303 1.25748
R15894 VDD.n1651 VDD.n1650 1.25267
R15895 VDD.n1655 VDD.n1654 1.21925
R15896 VDD.n557 VDD.n556 1.12991
R15897 VDD.n615 VDD.n614 1.12991
R15898 VDD.n640 VDD.n639 1.12991
R15899 VDD.n750 VDD.n749 1.12991
R15900 VDD.n703 VDD.n702 1.12991
R15901 VDD.n907 VDD.n906 1.12991
R15902 VDD.n965 VDD.n964 1.12991
R15903 VDD.n990 VDD.n989 1.12991
R15904 VDD.n1100 VDD.n1099 1.12991
R15905 VDD.n1053 VDD.n1052 1.12991
R15906 VDD.n156 VDD.n155 1.12991
R15907 VDD.n214 VDD.n213 1.12991
R15908 VDD.n113 VDD.n112 1.12991
R15909 VDD.n345 VDD.n344 1.12991
R15910 VDD.n298 VDD.n297 1.12991
R15911 VDD.n1336 VDD.n1335 1.12991
R15912 VDD.n1380 VDD.n1379 1.12991
R15913 VDD.n1307 VDD.n1306 1.12991
R15914 VDD.n1466 VDD.n1465 1.12991
R15915 VDD.n1516 VDD.n1515 1.12991
R15916 VDD.n1652 VDD.n1651 1.11354
R15917 VDD.n1631 VDD.n1630 1.11354
R15918 VDD.n1623 VDD.n1613 1.10388
R15919 VDD.n1731 VDD.n1716 1.06717
R15920 VDD.n2080 VDD.n2065 1.06717
R15921 VDD.n2310 VDD.n2295 1.06717
R15922 VDD.n2568 VDD.n2553 1.06717
R15923 VDD.n2826 VDD.n2811 1.06717
R15924 VDD.n3084 VDD.n3069 1.06717
R15925 VDD.n3342 VDD.n3327 1.06717
R15926 VDD.n5665 VDD.n5650 1.06717
R15927 VDD.n5411 VDD.n5396 1.06717
R15928 VDD.n3600 VDD.n3585 1.06717
R15929 VDD.n3858 VDD.n3843 1.06717
R15930 VDD.n4116 VDD.n4101 1.06717
R15931 VDD.n4374 VDD.n4359 1.06717
R15932 VDD.n4632 VDD.n4617 1.06717
R15933 VDD.n4890 VDD.n4875 1.06717
R15934 VDD.n5148 VDD.n5133 1.06717
R15935 VDD.n1608 VDD.n1606 1.06717
R15936 VDD.n1607 VDD 1.06717
R15937 VDD.n1873 VDD.n1872 1.00783
R15938 VDD.n2194 VDD.n2193 1.00687
R15939 VDD.n2452 VDD.n2451 1.00687
R15940 VDD.n2710 VDD.n2709 1.00687
R15941 VDD.n2968 VDD.n2967 1.00687
R15942 VDD.n3226 VDD.n3225 1.00687
R15943 VDD.n3484 VDD.n3483 1.00687
R15944 VDD.n5804 VDD.n5803 1.00687
R15945 VDD.n5550 VDD.n5549 1.00687
R15946 VDD.n3742 VDD.n3741 1.00687
R15947 VDD.n4000 VDD.n3999 1.00687
R15948 VDD.n4258 VDD.n4257 1.00687
R15949 VDD.n4516 VDD.n4515 1.00687
R15950 VDD.n4774 VDD.n4773 1.00687
R15951 VDD.n5032 VDD.n5031 1.00687
R15952 VDD.n5290 VDD.n5289 1.00687
R15953 VDD.n1644 VDD 0.970197
R15954 VDD.n1704 VDD.n1681 0.9605
R15955 VDD.n2053 VDD.n2030 0.9605
R15956 VDD.n2283 VDD.n2260 0.9605
R15957 VDD.n2541 VDD.n2518 0.9605
R15958 VDD.n2799 VDD.n2776 0.9605
R15959 VDD.n3057 VDD.n3034 0.9605
R15960 VDD.n3315 VDD.n3292 0.9605
R15961 VDD.n5638 VDD.n5615 0.9605
R15962 VDD.n5384 VDD.n5361 0.9605
R15963 VDD.n3573 VDD.n3550 0.9605
R15964 VDD.n3831 VDD.n3808 0.9605
R15965 VDD.n4089 VDD.n4066 0.9605
R15966 VDD.n4347 VDD.n4324 0.9605
R15967 VDD.n4605 VDD.n4582 0.9605
R15968 VDD.n4863 VDD.n4840 0.9605
R15969 VDD.n5121 VDD.n5098 0.9605
R15970 VDD.n1603 VDD.n1245 0.939577
R15971 VDD.n5859 VDD.n1982 0.885753
R15972 VDD.n1662 VDD.n1661 0.87764
R15973 VDD.n796 VDD.n407 0.826983
R15974 VDD.n1598 VDD.n1565 0.826983
R15975 VDD.n1933 VDD.n1924 0.800961
R15976 VDD.n5861 VDD 0.78236
R15977 VDD.n1619 VDD.n1618 0.7685
R15978 VDD.n1956 VDD.n1943 0.738962
R15979 VDD.n1638 VDD.n1636 0.686214
R15980 VDD.n1657 VDD.n1656 0.683536
R15981 VDD.n1663 VDD.n1603 0.673542
R15982 VDD.n1693 VDD.n1685 0.6405
R15983 VDD.n2042 VDD.n2034 0.6405
R15984 VDD.n2272 VDD.n2264 0.6405
R15985 VDD.n2530 VDD.n2522 0.6405
R15986 VDD.n2788 VDD.n2780 0.6405
R15987 VDD.n3046 VDD.n3038 0.6405
R15988 VDD.n3304 VDD.n3296 0.6405
R15989 VDD.n5627 VDD.n5619 0.6405
R15990 VDD.n5373 VDD.n5365 0.6405
R15991 VDD.n3562 VDD.n3554 0.6405
R15992 VDD.n3820 VDD.n3812 0.6405
R15993 VDD.n4078 VDD.n4070 0.6405
R15994 VDD.n4336 VDD.n4328 0.6405
R15995 VDD.n4594 VDD.n4586 0.6405
R15996 VDD.n4852 VDD.n4844 0.6405
R15997 VDD.n5110 VDD.n5102 0.6405
R15998 VDD.n1688 VDD.n1687 0.590778
R15999 VDD.n2037 VDD.n2036 0.590778
R16000 VDD.n2267 VDD.n2266 0.590778
R16001 VDD.n2525 VDD.n2524 0.590778
R16002 VDD.n2783 VDD.n2782 0.590778
R16003 VDD.n3041 VDD.n3040 0.590778
R16004 VDD.n3299 VDD.n3298 0.590778
R16005 VDD.n5622 VDD.n5621 0.590778
R16006 VDD.n5368 VDD.n5367 0.590778
R16007 VDD.n3557 VDD.n3556 0.590778
R16008 VDD.n3815 VDD.n3814 0.590778
R16009 VDD.n4073 VDD.n4072 0.590778
R16010 VDD.n4331 VDD.n4330 0.590778
R16011 VDD.n4589 VDD.n4588 0.590778
R16012 VDD.n4847 VDD.n4846 0.590778
R16013 VDD.n5105 VDD.n5104 0.590778
R16014 VDD.n5739 VDD.n5738 0.588569
R16015 VDD.n5485 VDD.n5484 0.588569
R16016 VDD.n1805 VDD.n1804 0.580785
R16017 VDD.n2384 VDD.n2383 0.580785
R16018 VDD.n2642 VDD.n2641 0.580785
R16019 VDD.n2900 VDD.n2899 0.580785
R16020 VDD.n3158 VDD.n3157 0.580785
R16021 VDD.n3416 VDD.n3415 0.580785
R16022 VDD.n3674 VDD.n3673 0.580785
R16023 VDD.n3932 VDD.n3931 0.580785
R16024 VDD.n4190 VDD.n4189 0.580785
R16025 VDD.n4448 VDD.n4447 0.580785
R16026 VDD.n4706 VDD.n4705 0.580785
R16027 VDD.n4964 VDD.n4963 0.580785
R16028 VDD.n5222 VDD.n5221 0.580785
R16029 VDD.n1658 VDD.n1657 0.571929
R16030 VDD.n1660 VDD.n1659 0.558536
R16031 VDD.n795 VDD.n438 0.557954
R16032 VDD.n1597 VDD.n1596 0.557954
R16033 VDD.n1659 VDD.n1658 0.549607
R16034 VDD.n1748 VDD.n1723 0.514389
R16035 VDD.n2097 VDD.n2072 0.514389
R16036 VDD.n2327 VDD.n2302 0.514389
R16037 VDD.n2585 VDD.n2560 0.514389
R16038 VDD.n2843 VDD.n2818 0.514389
R16039 VDD.n3101 VDD.n3076 0.514389
R16040 VDD.n3359 VDD.n3334 0.514389
R16041 VDD.n5682 VDD.n5657 0.514389
R16042 VDD.n5428 VDD.n5403 0.514389
R16043 VDD.n3617 VDD.n3592 0.514389
R16044 VDD.n3875 VDD.n3850 0.514389
R16045 VDD.n4133 VDD.n4108 0.514389
R16046 VDD.n4391 VDD.n4366 0.514389
R16047 VDD.n4649 VDD.n4624 0.514389
R16048 VDD.n4907 VDD.n4882 0.514389
R16049 VDD.n5165 VDD.n5140 0.514389
R16050 VDD.n1977 VDD.n1925 0.5125
R16051 VDD.n1839 VDD.n1826 0.492808
R16052 VDD.n2160 VDD.n2147 0.492808
R16053 VDD.n2418 VDD.n2405 0.492808
R16054 VDD.n2676 VDD.n2663 0.492808
R16055 VDD.n2934 VDD.n2921 0.492808
R16056 VDD.n3192 VDD.n3179 0.492808
R16057 VDD.n3450 VDD.n3437 0.492808
R16058 VDD.n5770 VDD.n5757 0.492808
R16059 VDD.n5516 VDD.n5503 0.492808
R16060 VDD.n3708 VDD.n3695 0.492808
R16061 VDD.n3966 VDD.n3953 0.492808
R16062 VDD.n4224 VDD.n4211 0.492808
R16063 VDD.n4482 VDD.n4469 0.492808
R16064 VDD.n4740 VDD.n4727 0.492808
R16065 VDD.n4998 VDD.n4985 0.492808
R16066 VDD.n5256 VDD.n5243 0.492808
R16067 VDD.n26 VDD 0.476404
R16068 VDD.n1170 VDD 0.476404
R16069 VDD.n1686 VDD.n1665 0.471224
R16070 VDD.n2035 VDD.n2014 0.471224
R16071 VDD.n2265 VDD.n2244 0.471224
R16072 VDD.n2523 VDD.n2502 0.471224
R16073 VDD.n2781 VDD.n2760 0.471224
R16074 VDD.n3039 VDD.n3018 0.471224
R16075 VDD.n3297 VDD.n3276 0.471224
R16076 VDD.n5620 VDD.n5599 0.471224
R16077 VDD.n5366 VDD.n5345 0.471224
R16078 VDD.n3555 VDD.n3534 0.471224
R16079 VDD.n3813 VDD.n3792 0.471224
R16080 VDD.n4071 VDD.n4050 0.471224
R16081 VDD.n4329 VDD.n4308 0.471224
R16082 VDD.n4587 VDD.n4566 0.471224
R16083 VDD.n4845 VDD.n4824 0.471224
R16084 VDD.n5103 VDD.n5082 0.471224
R16085 VDD.n1773 VDD.n1666 0.467504
R16086 VDD.n2122 VDD.n2015 0.467504
R16087 VDD.n2352 VDD.n2245 0.467504
R16088 VDD.n2610 VDD.n2503 0.467504
R16089 VDD.n2868 VDD.n2761 0.467504
R16090 VDD.n3126 VDD.n3019 0.467504
R16091 VDD.n3384 VDD.n3277 0.467504
R16092 VDD.n5707 VDD.n5600 0.467504
R16093 VDD.n5453 VDD.n5346 0.467504
R16094 VDD.n3642 VDD.n3535 0.467504
R16095 VDD.n3900 VDD.n3793 0.467504
R16096 VDD.n4158 VDD.n4051 0.467504
R16097 VDD.n4416 VDD.n4309 0.467504
R16098 VDD.n4674 VDD.n4567 0.467504
R16099 VDD.n4932 VDD.n4825 0.467504
R16100 VDD.n5190 VDD.n5083 0.467504
R16101 VDD.n1654 VDD.n1653 0.464786
R16102 VDD.n1637 VDD 0.457643
R16103 VDD.n1661 VDD.n1623 0.424377
R16104 VDD.n1810 VDD 0.411214
R16105 VDD.n2131 VDD 0.411214
R16106 VDD.n2389 VDD 0.411214
R16107 VDD.n2647 VDD 0.411214
R16108 VDD.n2905 VDD 0.411214
R16109 VDD.n3163 VDD 0.411214
R16110 VDD.n3421 VDD 0.411214
R16111 VDD.n5741 VDD 0.411214
R16112 VDD.n5487 VDD 0.411214
R16113 VDD.n3679 VDD 0.411214
R16114 VDD.n3937 VDD 0.411214
R16115 VDD.n4195 VDD 0.411214
R16116 VDD.n4453 VDD 0.411214
R16117 VDD.n4711 VDD 0.411214
R16118 VDD.n4969 VDD 0.411214
R16119 VDD.n5227 VDD 0.411214
R16120 VDD.n1753 VDD.n1752 0.410606
R16121 VDD.n2102 VDD.n2101 0.410606
R16122 VDD.n2332 VDD.n2331 0.410606
R16123 VDD.n2590 VDD.n2589 0.410606
R16124 VDD.n2848 VDD.n2847 0.410606
R16125 VDD.n3106 VDD.n3105 0.410606
R16126 VDD.n3364 VDD.n3363 0.410606
R16127 VDD.n5687 VDD.n5686 0.410606
R16128 VDD.n5433 VDD.n5432 0.410606
R16129 VDD.n3622 VDD.n3621 0.410606
R16130 VDD.n3880 VDD.n3879 0.410606
R16131 VDD.n4138 VDD.n4137 0.410606
R16132 VDD.n4396 VDD.n4395 0.410606
R16133 VDD.n4654 VDD.n4653 0.410606
R16134 VDD.n4912 VDD.n4911 0.410606
R16135 VDD.n5170 VDD.n5169 0.410606
R16136 VDD.n1921 VDD.n1920 0.409102
R16137 VDD.n2242 VDD.n2241 0.409102
R16138 VDD.n2500 VDD.n2499 0.409102
R16139 VDD.n2758 VDD.n2757 0.409102
R16140 VDD.n3016 VDD.n3015 0.409102
R16141 VDD.n3274 VDD.n3273 0.409102
R16142 VDD.n3532 VDD.n3531 0.409102
R16143 VDD.n3790 VDD.n3789 0.409102
R16144 VDD.n4048 VDD.n4047 0.409102
R16145 VDD.n4306 VDD.n4305 0.409102
R16146 VDD.n4564 VDD.n4563 0.409102
R16147 VDD.n4822 VDD.n4821 0.409102
R16148 VDD.n5080 VDD.n5079 0.409102
R16149 VDD.n5338 VDD.n5337 0.409102
R16150 VDD VDD.n26 0.403703
R16151 VDD VDD.n1170 0.403703
R16152 VDD.n1738 VDD.n1737 0.399706
R16153 VDD.n2087 VDD.n2086 0.399706
R16154 VDD.n2317 VDD.n2316 0.399706
R16155 VDD.n2575 VDD.n2574 0.399706
R16156 VDD.n2833 VDD.n2832 0.399706
R16157 VDD.n3091 VDD.n3090 0.399706
R16158 VDD.n3349 VDD.n3348 0.399706
R16159 VDD.n5672 VDD.n5671 0.399706
R16160 VDD.n5418 VDD.n5417 0.399706
R16161 VDD.n3607 VDD.n3606 0.399706
R16162 VDD.n3865 VDD.n3864 0.399706
R16163 VDD.n4123 VDD.n4122 0.399706
R16164 VDD.n4381 VDD.n4380 0.399706
R16165 VDD.n4639 VDD.n4638 0.399706
R16166 VDD.n4897 VDD.n4896 0.399706
R16167 VDD.n5155 VDD.n5154 0.399706
R16168 VDD.n513 VDD.n464 0.399037
R16169 VDD.n62 VDD.n61 0.399037
R16170 VDD.n1749 VDD.n1748 0.398914
R16171 VDD.n2098 VDD.n2097 0.398914
R16172 VDD.n2328 VDD.n2327 0.398914
R16173 VDD.n2586 VDD.n2585 0.398914
R16174 VDD.n2844 VDD.n2843 0.398914
R16175 VDD.n3102 VDD.n3101 0.398914
R16176 VDD.n3360 VDD.n3359 0.398914
R16177 VDD.n5683 VDD.n5682 0.398914
R16178 VDD.n5429 VDD.n5428 0.398914
R16179 VDD.n3618 VDD.n3617 0.398914
R16180 VDD.n3876 VDD.n3875 0.398914
R16181 VDD.n4134 VDD.n4133 0.398914
R16182 VDD.n4392 VDD.n4391 0.398914
R16183 VDD.n4650 VDD.n4649 0.398914
R16184 VDD.n4908 VDD.n4907 0.398914
R16185 VDD.n5166 VDD.n5165 0.398914
R16186 VDD.n1737 VDD.n1723 0.398403
R16187 VDD.n2086 VDD.n2072 0.398403
R16188 VDD.n2316 VDD.n2302 0.398403
R16189 VDD.n2574 VDD.n2560 0.398403
R16190 VDD.n2832 VDD.n2818 0.398403
R16191 VDD.n3090 VDD.n3076 0.398403
R16192 VDD.n3348 VDD.n3334 0.398403
R16193 VDD.n5671 VDD.n5657 0.398403
R16194 VDD.n5417 VDD.n5403 0.398403
R16195 VDD.n3606 VDD.n3592 0.398403
R16196 VDD.n3864 VDD.n3850 0.398403
R16197 VDD.n4122 VDD.n4108 0.398403
R16198 VDD.n4380 VDD.n4366 0.398403
R16199 VDD.n4638 VDD.n4624 0.398403
R16200 VDD.n4896 VDD.n4882 0.398403
R16201 VDD.n5154 VDD.n5140 0.398403
R16202 VDD.n1656 VDD.n1655 0.384429
R16203 VDD.n1807 VDD.n1806 0.3805
R16204 VDD.n2127 VDD.n2126 0.3805
R16205 VDD.n2386 VDD.n2385 0.3805
R16206 VDD.n2644 VDD.n2643 0.3805
R16207 VDD.n2902 VDD.n2901 0.3805
R16208 VDD.n3160 VDD.n3159 0.3805
R16209 VDD.n3418 VDD.n3417 0.3805
R16210 VDD.n3676 VDD.n3675 0.3805
R16211 VDD.n3934 VDD.n3933 0.3805
R16212 VDD.n4192 VDD.n4191 0.3805
R16213 VDD.n4450 VDD.n4449 0.3805
R16214 VDD.n4708 VDD.n4707 0.3805
R16215 VDD.n4966 VDD.n4965 0.3805
R16216 VDD.n5224 VDD.n5223 0.3805
R16217 VDD.n547 VDD.n546 0.376971
R16218 VDD.n627 VDD.n626 0.376971
R16219 VDD.n787 VDD.n786 0.376971
R16220 VDD.n739 VDD.n738 0.376971
R16221 VDD.n897 VDD.n896 0.376971
R16222 VDD.n977 VDD.n976 0.376971
R16223 VDD.n1137 VDD.n1136 0.376971
R16224 VDD.n1089 VDD.n1088 0.376971
R16225 VDD.n146 VDD.n145 0.376971
R16226 VDD.n226 VDD.n225 0.376971
R16227 VDD.n382 VDD.n381 0.376971
R16228 VDD.n334 VDD.n333 0.376971
R16229 VDD.n1452 VDD.n1451 0.376971
R16230 VDD.n1421 VDD.n1420 0.376971
R16231 VDD.n1266 VDD.n1265 0.376971
R16232 VDD.n1500 VDD.n1499 0.376971
R16233 VDD.n1687 VDD.n1686 0.368458
R16234 VDD.n2036 VDD.n2035 0.368458
R16235 VDD.n2266 VDD.n2265 0.368458
R16236 VDD.n2524 VDD.n2523 0.368458
R16237 VDD.n2782 VDD.n2781 0.368458
R16238 VDD.n3040 VDD.n3039 0.368458
R16239 VDD.n3298 VDD.n3297 0.368458
R16240 VDD.n5621 VDD.n5620 0.368458
R16241 VDD.n5367 VDD.n5366 0.368458
R16242 VDD.n3556 VDD.n3555 0.368458
R16243 VDD.n3814 VDD.n3813 0.368458
R16244 VDD.n4072 VDD.n4071 0.368458
R16245 VDD.n4330 VDD.n4329 0.368458
R16246 VDD.n4588 VDD.n4587 0.368458
R16247 VDD.n4846 VDD.n4845 0.368458
R16248 VDD.n5104 VDD.n5103 0.368458
R16249 VDD.n1688 VDD.n1666 0.361663
R16250 VDD.n2037 VDD.n2015 0.361663
R16251 VDD.n2267 VDD.n2245 0.361663
R16252 VDD.n2525 VDD.n2503 0.361663
R16253 VDD.n2783 VDD.n2761 0.361663
R16254 VDD.n3041 VDD.n3019 0.361663
R16255 VDD.n3299 VDD.n3277 0.361663
R16256 VDD.n5622 VDD.n5600 0.361663
R16257 VDD.n5368 VDD.n5346 0.361663
R16258 VDD.n3557 VDD.n3535 0.361663
R16259 VDD.n3815 VDD.n3793 0.361663
R16260 VDD.n4073 VDD.n4051 0.361663
R16261 VDD.n4331 VDD.n4309 0.361663
R16262 VDD.n4589 VDD.n4567 0.361663
R16263 VDD.n4847 VDD.n4825 0.361663
R16264 VDD.n5105 VDD.n5083 0.361663
R16265 VDD.n1750 VDD.n1749 0.357683
R16266 VDD.n2099 VDD.n2098 0.357683
R16267 VDD.n2329 VDD.n2328 0.357683
R16268 VDD.n2587 VDD.n2586 0.357683
R16269 VDD.n2845 VDD.n2844 0.357683
R16270 VDD.n3103 VDD.n3102 0.357683
R16271 VDD.n3361 VDD.n3360 0.357683
R16272 VDD.n5684 VDD.n5683 0.357683
R16273 VDD.n5430 VDD.n5429 0.357683
R16274 VDD.n3619 VDD.n3618 0.357683
R16275 VDD.n3877 VDD.n3876 0.357683
R16276 VDD.n4135 VDD.n4134 0.357683
R16277 VDD.n4393 VDD.n4392 0.357683
R16278 VDD.n4651 VDD.n4650 0.357683
R16279 VDD.n4909 VDD.n4908 0.357683
R16280 VDD.n5167 VDD.n5166 0.357683
R16281 VDD.n1734 VDD.n1732 0.356056
R16282 VDD.n2083 VDD.n2081 0.356056
R16283 VDD.n2313 VDD.n2311 0.356056
R16284 VDD.n2571 VDD.n2569 0.356056
R16285 VDD.n2829 VDD.n2827 0.356056
R16286 VDD.n3087 VDD.n3085 0.356056
R16287 VDD.n3345 VDD.n3343 0.356056
R16288 VDD.n5668 VDD.n5666 0.356056
R16289 VDD.n5414 VDD.n5412 0.356056
R16290 VDD.n3603 VDD.n3601 0.356056
R16291 VDD.n3861 VDD.n3859 0.356056
R16292 VDD.n4119 VDD.n4117 0.356056
R16293 VDD.n4377 VDD.n4375 0.356056
R16294 VDD.n4635 VDD.n4633 0.356056
R16295 VDD.n4893 VDD.n4891 0.356056
R16296 VDD.n5151 VDD.n5149 0.356056
R16297 VDD.n35 VDD.n34 0.35558
R16298 VDD.n1179 VDD.n1178 0.35558
R16299 VDD.n1836 VDD 0.355332
R16300 VDD.n2157 VDD 0.355332
R16301 VDD.n2415 VDD 0.355332
R16302 VDD.n2673 VDD 0.355332
R16303 VDD.n2931 VDD 0.355332
R16304 VDD.n3189 VDD 0.355332
R16305 VDD.n3447 VDD 0.355332
R16306 VDD.n5767 VDD 0.355332
R16307 VDD.n5513 VDD 0.355332
R16308 VDD.n3705 VDD 0.355332
R16309 VDD.n3963 VDD 0.355332
R16310 VDD.n4221 VDD 0.355332
R16311 VDD.n4479 VDD 0.355332
R16312 VDD.n4737 VDD 0.355332
R16313 VDD.n4995 VDD 0.355332
R16314 VDD.n5253 VDD 0.355332
R16315 VDD.n1918 VDD.n1887 0.349136
R16316 VDD.n2239 VDD.n2208 0.349136
R16317 VDD.n2497 VDD.n2466 0.349136
R16318 VDD.n2755 VDD.n2724 0.349136
R16319 VDD.n3013 VDD.n2982 0.349136
R16320 VDD.n3271 VDD.n3240 0.349136
R16321 VDD.n3529 VDD.n3498 0.349136
R16322 VDD.n5849 VDD.n5818 0.349136
R16323 VDD.n5595 VDD.n5564 0.349136
R16324 VDD.n3787 VDD.n3756 0.349136
R16325 VDD.n4045 VDD.n4014 0.349136
R16326 VDD.n4303 VDD.n4272 0.349136
R16327 VDD.n4561 VDD.n4530 0.349136
R16328 VDD.n4819 VDD.n4788 0.349136
R16329 VDD.n5077 VDD.n5046 0.349136
R16330 VDD.n5335 VDD.n5304 0.349136
R16331 VDD.n0 VDD 0.340206
R16332 VDD.n1144 VDD 0.340206
R16333 VDD.n1692 VDD.n1687 0.340142
R16334 VDD.n2041 VDD.n2036 0.340142
R16335 VDD.n2271 VDD.n2266 0.340142
R16336 VDD.n2529 VDD.n2524 0.340142
R16337 VDD.n2787 VDD.n2782 0.340142
R16338 VDD.n3045 VDD.n3040 0.340142
R16339 VDD.n3303 VDD.n3298 0.340142
R16340 VDD.n5626 VDD.n5621 0.340142
R16341 VDD.n5372 VDD.n5367 0.340142
R16342 VDD.n3561 VDD.n3556 0.340142
R16343 VDD.n3819 VDD.n3814 0.340142
R16344 VDD.n4077 VDD.n4072 0.340142
R16345 VDD.n4335 VDD.n4330 0.340142
R16346 VDD.n4593 VDD.n4588 0.340142
R16347 VDD.n4851 VDD.n4846 0.340142
R16348 VDD.n5109 VDD.n5104 0.340142
R16349 VDD.n1283 VDD 0.330819
R16350 VDD.n1768 VDD.n1671 0.3205
R16351 VDD.n1693 VDD.n1684 0.3205
R16352 VDD.n2117 VDD.n2020 0.3205
R16353 VDD.n2042 VDD.n2033 0.3205
R16354 VDD.n2347 VDD.n2250 0.3205
R16355 VDD.n2272 VDD.n2263 0.3205
R16356 VDD.n2605 VDD.n2508 0.3205
R16357 VDD.n2530 VDD.n2521 0.3205
R16358 VDD.n2863 VDD.n2766 0.3205
R16359 VDD.n2788 VDD.n2779 0.3205
R16360 VDD.n3121 VDD.n3024 0.3205
R16361 VDD.n3046 VDD.n3037 0.3205
R16362 VDD.n3379 VDD.n3282 0.3205
R16363 VDD.n3304 VDD.n3295 0.3205
R16364 VDD.n5702 VDD.n5605 0.3205
R16365 VDD.n5627 VDD.n5618 0.3205
R16366 VDD.n5448 VDD.n5351 0.3205
R16367 VDD.n5373 VDD.n5364 0.3205
R16368 VDD.n3637 VDD.n3540 0.3205
R16369 VDD.n3562 VDD.n3553 0.3205
R16370 VDD.n3895 VDD.n3798 0.3205
R16371 VDD.n3820 VDD.n3811 0.3205
R16372 VDD.n4153 VDD.n4056 0.3205
R16373 VDD.n4078 VDD.n4069 0.3205
R16374 VDD.n4411 VDD.n4314 0.3205
R16375 VDD.n4336 VDD.n4327 0.3205
R16376 VDD.n4669 VDD.n4572 0.3205
R16377 VDD.n4594 VDD.n4585 0.3205
R16378 VDD.n4927 VDD.n4830 0.3205
R16379 VDD.n4852 VDD.n4843 0.3205
R16380 VDD.n5185 VDD.n5088 0.3205
R16381 VDD.n5110 VDD.n5101 0.3205
R16382 VDD.n1919 VDD.n1918 0.314572
R16383 VDD.n2240 VDD.n2239 0.314572
R16384 VDD.n2498 VDD.n2497 0.314572
R16385 VDD.n2756 VDD.n2755 0.314572
R16386 VDD.n3014 VDD.n3013 0.314572
R16387 VDD.n3272 VDD.n3271 0.314572
R16388 VDD.n3530 VDD.n3529 0.314572
R16389 VDD.n5850 VDD.n5849 0.314572
R16390 VDD.n5596 VDD.n5595 0.314572
R16391 VDD.n3788 VDD.n3787 0.314572
R16392 VDD.n4046 VDD.n4045 0.314572
R16393 VDD.n4304 VDD.n4303 0.314572
R16394 VDD.n4562 VDD.n4561 0.314572
R16395 VDD.n4820 VDD.n4819 0.314572
R16396 VDD.n5078 VDD.n5077 0.314572
R16397 VDD.n5336 VDD.n5335 0.314572
R16398 VDD.n1874 VDD.n1873 0.311403
R16399 VDD.n2195 VDD.n2194 0.311403
R16400 VDD.n2453 VDD.n2452 0.311403
R16401 VDD.n2711 VDD.n2710 0.311403
R16402 VDD.n2969 VDD.n2968 0.311403
R16403 VDD.n3227 VDD.n3226 0.311403
R16404 VDD.n3485 VDD.n3484 0.311403
R16405 VDD.n5805 VDD.n5804 0.311403
R16406 VDD.n5551 VDD.n5550 0.311403
R16407 VDD.n3743 VDD.n3742 0.311403
R16408 VDD.n4001 VDD.n4000 0.311403
R16409 VDD.n4259 VDD.n4258 0.311403
R16410 VDD.n4517 VDD.n4516 0.311403
R16411 VDD.n4775 VDD.n4774 0.311403
R16412 VDD.n5033 VDD.n5032 0.311403
R16413 VDD.n5291 VDD.n5290 0.311403
R16414 VDD.n1691 VDD.n1690 0.296036
R16415 VDD.n2040 VDD.n2039 0.296036
R16416 VDD.n2270 VDD.n2269 0.296036
R16417 VDD.n2528 VDD.n2527 0.296036
R16418 VDD.n2786 VDD.n2785 0.296036
R16419 VDD.n3044 VDD.n3043 0.296036
R16420 VDD.n3302 VDD.n3301 0.296036
R16421 VDD.n5625 VDD.n5624 0.296036
R16422 VDD.n5371 VDD.n5370 0.296036
R16423 VDD.n3560 VDD.n3559 0.296036
R16424 VDD.n3818 VDD.n3817 0.296036
R16425 VDD.n4076 VDD.n4075 0.296036
R16426 VDD.n4334 VDD.n4333 0.296036
R16427 VDD.n4592 VDD.n4591 0.296036
R16428 VDD.n4850 VDD.n4849 0.296036
R16429 VDD.n5108 VDD.n5107 0.296036
R16430 VDD.n1650 VDD 0.278761
R16431 VDD VDD.n5863 0.273495
R16432 VDD.n1747 VDD.n1724 0.261214
R16433 VDD.n1727 VDD.n1726 0.261214
R16434 VDD.n2096 VDD.n2073 0.261214
R16435 VDD.n2076 VDD.n2075 0.261214
R16436 VDD.n2326 VDD.n2303 0.261214
R16437 VDD.n2306 VDD.n2305 0.261214
R16438 VDD.n2584 VDD.n2561 0.261214
R16439 VDD.n2564 VDD.n2563 0.261214
R16440 VDD.n2842 VDD.n2819 0.261214
R16441 VDD.n2822 VDD.n2821 0.261214
R16442 VDD.n3100 VDD.n3077 0.261214
R16443 VDD.n3080 VDD.n3079 0.261214
R16444 VDD.n3358 VDD.n3335 0.261214
R16445 VDD.n3338 VDD.n3337 0.261214
R16446 VDD.n5681 VDD.n5658 0.261214
R16447 VDD.n5661 VDD.n5660 0.261214
R16448 VDD.n5427 VDD.n5404 0.261214
R16449 VDD.n5407 VDD.n5406 0.261214
R16450 VDD.n3616 VDD.n3593 0.261214
R16451 VDD.n3596 VDD.n3595 0.261214
R16452 VDD.n3874 VDD.n3851 0.261214
R16453 VDD.n3854 VDD.n3853 0.261214
R16454 VDD.n4132 VDD.n4109 0.261214
R16455 VDD.n4112 VDD.n4111 0.261214
R16456 VDD.n4390 VDD.n4367 0.261214
R16457 VDD.n4370 VDD.n4369 0.261214
R16458 VDD.n4648 VDD.n4625 0.261214
R16459 VDD.n4628 VDD.n4627 0.261214
R16460 VDD.n4906 VDD.n4883 0.261214
R16461 VDD.n4886 VDD.n4885 0.261214
R16462 VDD.n5164 VDD.n5141 0.261214
R16463 VDD.n5144 VDD.n5143 0.261214
R16464 VDD.n1745 VDD.n1725 0.2565
R16465 VDD.n2094 VDD.n2074 0.2565
R16466 VDD.n2324 VDD.n2304 0.2565
R16467 VDD.n2582 VDD.n2562 0.2565
R16468 VDD.n2840 VDD.n2820 0.2565
R16469 VDD.n3098 VDD.n3078 0.2565
R16470 VDD.n3356 VDD.n3336 0.2565
R16471 VDD.n5679 VDD.n5659 0.2565
R16472 VDD.n5425 VDD.n5405 0.2565
R16473 VDD.n3614 VDD.n3594 0.2565
R16474 VDD.n3872 VDD.n3852 0.2565
R16475 VDD.n4130 VDD.n4110 0.2565
R16476 VDD.n4388 VDD.n4368 0.2565
R16477 VDD.n4646 VDD.n4626 0.2565
R16478 VDD.n4904 VDD.n4884 0.2565
R16479 VDD.n5162 VDD.n5142 0.2565
R16480 VDD.n1736 VDD.n1735 0.251889
R16481 VDD.n2085 VDD.n2084 0.251889
R16482 VDD.n2315 VDD.n2314 0.251889
R16483 VDD.n2573 VDD.n2572 0.251889
R16484 VDD.n2831 VDD.n2830 0.251889
R16485 VDD.n3089 VDD.n3088 0.251889
R16486 VDD.n3347 VDD.n3346 0.251889
R16487 VDD.n5670 VDD.n5669 0.251889
R16488 VDD.n5416 VDD.n5415 0.251889
R16489 VDD.n3605 VDD.n3604 0.251889
R16490 VDD.n3863 VDD.n3862 0.251889
R16491 VDD.n4121 VDD.n4120 0.251889
R16492 VDD.n4379 VDD.n4378 0.251889
R16493 VDD.n4637 VDD.n4636 0.251889
R16494 VDD.n4895 VDD.n4894 0.251889
R16495 VDD.n5153 VDD.n5152 0.251889
R16496 VDD.n5851 VDD.n5739 0.25042
R16497 VDD.n5597 VDD.n5485 0.25042
R16498 VDD.n1754 VDD.n1719 0.248103
R16499 VDD.n2103 VDD.n2068 0.248103
R16500 VDD.n2333 VDD.n2298 0.248103
R16501 VDD.n2591 VDD.n2556 0.248103
R16502 VDD.n2849 VDD.n2814 0.248103
R16503 VDD.n3107 VDD.n3072 0.248103
R16504 VDD.n3365 VDD.n3330 0.248103
R16505 VDD.n5688 VDD.n5653 0.248103
R16506 VDD.n5434 VDD.n5399 0.248103
R16507 VDD.n3623 VDD.n3588 0.248103
R16508 VDD.n3881 VDD.n3846 0.248103
R16509 VDD.n4139 VDD.n4104 0.248103
R16510 VDD.n4397 VDD.n4362 0.248103
R16511 VDD.n4655 VDD.n4620 0.248103
R16512 VDD.n4913 VDD.n4878 0.248103
R16513 VDD.n5171 VDD.n5136 0.248103
R16514 VDD.n1770 VDD.n1668 0.247868
R16515 VDD.n2119 VDD.n2017 0.247868
R16516 VDD.n2349 VDD.n2247 0.247868
R16517 VDD.n2607 VDD.n2505 0.247868
R16518 VDD.n2865 VDD.n2763 0.247868
R16519 VDD.n3123 VDD.n3021 0.247868
R16520 VDD.n3381 VDD.n3279 0.247868
R16521 VDD.n5704 VDD.n5602 0.247868
R16522 VDD.n5450 VDD.n5348 0.247868
R16523 VDD.n3639 VDD.n3537 0.247868
R16524 VDD.n3897 VDD.n3795 0.247868
R16525 VDD.n4155 VDD.n4053 0.247868
R16526 VDD.n4413 VDD.n4311 0.247868
R16527 VDD.n4671 VDD.n4569 0.247868
R16528 VDD.n4929 VDD.n4827 0.247868
R16529 VDD.n5187 VDD.n5085 0.247868
R16530 VDD.n808 VDD.n807 0.240091
R16531 VDD.n1191 VDD.n1190 0.240091
R16532 VDD.n1738 VDD.n1721 0.232755
R16533 VDD.n2087 VDD.n2070 0.232755
R16534 VDD.n2317 VDD.n2300 0.232755
R16535 VDD.n2575 VDD.n2558 0.232755
R16536 VDD.n2833 VDD.n2816 0.232755
R16537 VDD.n3091 VDD.n3074 0.232755
R16538 VDD.n3349 VDD.n3332 0.232755
R16539 VDD.n5672 VDD.n5655 0.232755
R16540 VDD.n5418 VDD.n5401 0.232755
R16541 VDD.n3607 VDD.n3590 0.232755
R16542 VDD.n3865 VDD.n3848 0.232755
R16543 VDD.n4123 VDD.n4106 0.232755
R16544 VDD.n4381 VDD.n4364 0.232755
R16545 VDD.n4639 VDD.n4622 0.232755
R16546 VDD.n4897 VDD.n4880 0.232755
R16547 VDD.n5155 VDD.n5138 0.232755
R16548 VDD.n5862 VDD.n1181 0.231188
R16549 VDD.n1953 VDD.n1952 0.224662
R16550 VDD.n1730 VDD.n1722 0.217167
R16551 VDD.n2079 VDD.n2071 0.217167
R16552 VDD.n2309 VDD.n2301 0.217167
R16553 VDD.n2567 VDD.n2559 0.217167
R16554 VDD.n2825 VDD.n2817 0.217167
R16555 VDD.n3083 VDD.n3075 0.217167
R16556 VDD.n3341 VDD.n3333 0.217167
R16557 VDD.n5664 VDD.n5656 0.217167
R16558 VDD.n5410 VDD.n5402 0.217167
R16559 VDD.n3599 VDD.n3591 0.217167
R16560 VDD.n3857 VDD.n3849 0.217167
R16561 VDD.n4115 VDD.n4107 0.217167
R16562 VDD.n4373 VDD.n4365 0.217167
R16563 VDD.n4631 VDD.n4623 0.217167
R16564 VDD.n4889 VDD.n4881 0.217167
R16565 VDD.n5147 VDD.n5139 0.217167
R16566 VDD.n512 VDD.n511 0.212557
R16567 VDD.n110 VDD.n109 0.212557
R16568 VDD.n407 VDD.n406 0.211096
R16569 VDD.n1565 VDD.n1564 0.211096
R16570 VDD.n481 VDD 0.210222
R16571 VDD.n79 VDD 0.210222
R16572 VDD.n1702 VDD.n1701 0.204667
R16573 VDD.n2051 VDD.n2050 0.204667
R16574 VDD.n2281 VDD.n2280 0.204667
R16575 VDD.n2539 VDD.n2538 0.204667
R16576 VDD.n2797 VDD.n2796 0.204667
R16577 VDD.n3055 VDD.n3054 0.204667
R16578 VDD.n3313 VDD.n3312 0.204667
R16579 VDD.n5636 VDD.n5635 0.204667
R16580 VDD.n5382 VDD.n5381 0.204667
R16581 VDD.n3571 VDD.n3570 0.204667
R16582 VDD.n3829 VDD.n3828 0.204667
R16583 VDD.n4087 VDD.n4086 0.204667
R16584 VDD.n4345 VDD.n4344 0.204667
R16585 VDD.n4603 VDD.n4602 0.204667
R16586 VDD.n4861 VDD.n4860 0.204667
R16587 VDD.n5119 VDD.n5118 0.204667
R16588 VDD.n1662 VDD 0.2005
R16589 VDD.n1703 VDD.n1667 0.199111
R16590 VDD.n2052 VDD.n2016 0.199111
R16591 VDD.n2282 VDD.n2246 0.199111
R16592 VDD.n2540 VDD.n2504 0.199111
R16593 VDD.n2798 VDD.n2762 0.199111
R16594 VDD.n3056 VDD.n3020 0.199111
R16595 VDD.n3314 VDD.n3278 0.199111
R16596 VDD.n5637 VDD.n5601 0.199111
R16597 VDD.n5383 VDD.n5347 0.199111
R16598 VDD.n3572 VDD.n3536 0.199111
R16599 VDD.n3830 VDD.n3794 0.199111
R16600 VDD.n4088 VDD.n4052 0.199111
R16601 VDD.n4346 VDD.n4310 0.199111
R16602 VDD.n4604 VDD.n4568 0.199111
R16603 VDD.n4862 VDD.n4826 0.199111
R16604 VDD.n5120 VDD.n5084 0.199111
R16605 VDD.n28 VDD 0.196824
R16606 VDD.n1172 VDD 0.196824
R16607 VDD.n1816 VDD.n1815 0.192557
R16608 VDD.n2137 VDD.n2136 0.192557
R16609 VDD.n2395 VDD.n2394 0.192557
R16610 VDD.n2653 VDD.n2652 0.192557
R16611 VDD.n2911 VDD.n2910 0.192557
R16612 VDD.n3169 VDD.n3168 0.192557
R16613 VDD.n3427 VDD.n3426 0.192557
R16614 VDD.n5747 VDD.n5746 0.192557
R16615 VDD.n5493 VDD.n5492 0.192557
R16616 VDD.n3685 VDD.n3684 0.192557
R16617 VDD.n3943 VDD.n3942 0.192557
R16618 VDD.n4201 VDD.n4200 0.192557
R16619 VDD.n4459 VDD.n4458 0.192557
R16620 VDD.n4717 VDD.n4716 0.192557
R16621 VDD.n4975 VDD.n4974 0.192557
R16622 VDD.n5233 VDD.n5232 0.192557
R16623 VDD.n1811 VDD.n1810 0.192167
R16624 VDD.n2132 VDD.n2131 0.192167
R16625 VDD.n2390 VDD.n2389 0.192167
R16626 VDD.n2648 VDD.n2647 0.192167
R16627 VDD.n2906 VDD.n2905 0.192167
R16628 VDD.n3164 VDD.n3163 0.192167
R16629 VDD.n3422 VDD.n3421 0.192167
R16630 VDD.n5742 VDD.n5741 0.192167
R16631 VDD.n5488 VDD.n5487 0.192167
R16632 VDD.n3680 VDD.n3679 0.192167
R16633 VDD.n3938 VDD.n3937 0.192167
R16634 VDD.n4196 VDD.n4195 0.192167
R16635 VDD.n4454 VDD.n4453 0.192167
R16636 VDD.n4712 VDD.n4711 0.192167
R16637 VDD.n4970 VDD.n4969 0.192167
R16638 VDD.n5228 VDD.n5227 0.192167
R16639 VDD.n5863 VDD.n863 0.189
R16640 VDD.n34 VDD.n33 0.183651
R16641 VDD.n1178 VDD.n1177 0.183651
R16642 VDD.n1804 VDD.n1776 0.180841
R16643 VDD.n2012 VDD.n1984 0.180841
R16644 VDD.n2383 VDD.n2355 0.180841
R16645 VDD.n2641 VDD.n2613 0.180841
R16646 VDD.n2899 VDD.n2871 0.180841
R16647 VDD.n3157 VDD.n3129 0.180841
R16648 VDD.n3415 VDD.n3387 0.180841
R16649 VDD.n5738 VDD.n5710 0.180841
R16650 VDD.n5484 VDD.n5456 0.180841
R16651 VDD.n3673 VDD.n3645 0.180841
R16652 VDD.n3931 VDD.n3903 0.180841
R16653 VDD.n4189 VDD.n4161 0.180841
R16654 VDD.n4447 VDD.n4419 0.180841
R16655 VDD.n4705 VDD.n4677 0.180841
R16656 VDD.n4963 VDD.n4935 0.180841
R16657 VDD.n5221 VDD.n5193 0.180841
R16658 VDD.n511 VDD.n510 0.175873
R16659 VDD.n109 VDD.n108 0.175873
R16660 VDD.n1599 VDD.n1548 0.168948
R16661 VDD.n1760 VDD.n1759 0.164944
R16662 VDD.n1759 VDD.n1711 0.164944
R16663 VDD.n2109 VDD.n2108 0.164944
R16664 VDD.n2108 VDD.n2060 0.164944
R16665 VDD.n2339 VDD.n2338 0.164944
R16666 VDD.n2338 VDD.n2290 0.164944
R16667 VDD.n2597 VDD.n2596 0.164944
R16668 VDD.n2596 VDD.n2548 0.164944
R16669 VDD.n2855 VDD.n2854 0.164944
R16670 VDD.n2854 VDD.n2806 0.164944
R16671 VDD.n3113 VDD.n3112 0.164944
R16672 VDD.n3112 VDD.n3064 0.164944
R16673 VDD.n3371 VDD.n3370 0.164944
R16674 VDD.n3370 VDD.n3322 0.164944
R16675 VDD.n5694 VDD.n5693 0.164944
R16676 VDD.n5693 VDD.n5645 0.164944
R16677 VDD.n5440 VDD.n5439 0.164944
R16678 VDD.n5439 VDD.n5391 0.164944
R16679 VDD.n3629 VDD.n3628 0.164944
R16680 VDD.n3628 VDD.n3580 0.164944
R16681 VDD.n3887 VDD.n3886 0.164944
R16682 VDD.n3886 VDD.n3838 0.164944
R16683 VDD.n4145 VDD.n4144 0.164944
R16684 VDD.n4144 VDD.n4096 0.164944
R16685 VDD.n4403 VDD.n4402 0.164944
R16686 VDD.n4402 VDD.n4354 0.164944
R16687 VDD.n4661 VDD.n4660 0.164944
R16688 VDD.n4660 VDD.n4612 0.164944
R16689 VDD.n4919 VDD.n4918 0.164944
R16690 VDD.n4918 VDD.n4870 0.164944
R16691 VDD.n5177 VDD.n5176 0.164944
R16692 VDD.n5176 VDD.n5128 0.164944
R16693 VDD.n1710 VDD.n1709 0.159358
R16694 VDD.n2059 VDD.n2058 0.159358
R16695 VDD.n2289 VDD.n2288 0.159358
R16696 VDD.n2547 VDD.n2546 0.159358
R16697 VDD.n2805 VDD.n2804 0.159358
R16698 VDD.n3063 VDD.n3062 0.159358
R16699 VDD.n3321 VDD.n3320 0.159358
R16700 VDD.n5644 VDD.n5643 0.159358
R16701 VDD.n5390 VDD.n5389 0.159358
R16702 VDD.n3579 VDD.n3578 0.159358
R16703 VDD.n3837 VDD.n3836 0.159358
R16704 VDD.n4095 VDD.n4094 0.159358
R16705 VDD.n4353 VDD.n4352 0.159358
R16706 VDD.n4611 VDD.n4610 0.159358
R16707 VDD.n4869 VDD.n4868 0.159358
R16708 VDD.n5127 VDD.n5126 0.159358
R16709 VDD.n1709 VDD.n1708 0.15889
R16710 VDD.n2058 VDD.n2057 0.15889
R16711 VDD.n2288 VDD.n2287 0.15889
R16712 VDD.n2546 VDD.n2545 0.15889
R16713 VDD.n2804 VDD.n2803 0.15889
R16714 VDD.n3062 VDD.n3061 0.15889
R16715 VDD.n3320 VDD.n3319 0.15889
R16716 VDD.n5643 VDD.n5642 0.15889
R16717 VDD.n5389 VDD.n5388 0.15889
R16718 VDD.n3578 VDD.n3577 0.15889
R16719 VDD.n3836 VDD.n3835 0.15889
R16720 VDD.n4094 VDD.n4093 0.15889
R16721 VDD.n4352 VDD.n4351 0.15889
R16722 VDD.n4610 VDD.n4609 0.15889
R16723 VDD.n4868 VDD.n4867 0.15889
R16724 VDD.n5126 VDD.n5125 0.15889
R16725 VDD.n438 VDD.n437 0.155541
R16726 VDD.n1596 VDD.n1595 0.155541
R16727 VDD.n27 VDD 0.145087
R16728 VDD.n1171 VDD 0.145087
R16729 VDD VDD.n820 0.137071
R16730 VDD VDD.n1203 0.137071
R16731 VDD.n5339 VDD.n5338 0.135642
R16732 VDD.n5861 VDD.n1663 0.134625
R16733 VDD.n852 VDD.n851 0.128415
R16734 VDD.n1235 VDD.n1234 0.128415
R16735 VDD.n464 VDD.n462 0.120987
R16736 VDD.n61 VDD.n59 0.120987
R16737 VDD.n853 VDD.n852 0.119283
R16738 VDD.n1236 VDD.n1235 0.119283
R16739 VDD.n5851 VDD.n5850 0.118114
R16740 VDD.n5597 VDD.n5596 0.118114
R16741 VDD.n1774 VDD.n1773 0.117306
R16742 VDD.n2123 VDD.n2122 0.117306
R16743 VDD.n2353 VDD.n2352 0.117306
R16744 VDD.n2611 VDD.n2610 0.117306
R16745 VDD.n2869 VDD.n2868 0.117306
R16746 VDD.n3127 VDD.n3126 0.117306
R16747 VDD.n3385 VDD.n3384 0.117306
R16748 VDD.n5708 VDD.n5707 0.117306
R16749 VDD.n5454 VDD.n5453 0.117306
R16750 VDD.n3643 VDD.n3642 0.117306
R16751 VDD.n3901 VDD.n3900 0.117306
R16752 VDD.n4159 VDD.n4158 0.117306
R16753 VDD.n4417 VDD.n4416 0.117306
R16754 VDD.n4675 VDD.n4674 0.117306
R16755 VDD.n4933 VDD.n4932 0.117306
R16756 VDD.n5191 VDD.n5190 0.117306
R16757 VDD.n794 VDD.n793 0.116581
R16758 VDD.n848 VDD.n847 0.1155
R16759 VDD.n847 VDD.n845 0.1155
R16760 VDD.n842 VDD.n841 0.1155
R16761 VDD.n841 VDD.n839 0.1155
R16762 VDD.n836 VDD.n835 0.1155
R16763 VDD.n835 VDD.n833 0.1155
R16764 VDD.n830 VDD.n829 0.1155
R16765 VDD.n829 VDD.n827 0.1155
R16766 VDD.n1231 VDD.n1230 0.1155
R16767 VDD.n1230 VDD.n1228 0.1155
R16768 VDD.n1225 VDD.n1224 0.1155
R16769 VDD.n1224 VDD.n1222 0.1155
R16770 VDD.n1219 VDD.n1218 0.1155
R16771 VDD.n1218 VDD.n1216 0.1155
R16772 VDD.n1213 VDD.n1212 0.1155
R16773 VDD.n1212 VDD.n1210 0.1155
R16774 VDD.n862 VDD 0.109094
R16775 VDD.n1245 VDD 0.109094
R16776 VDD.n862 VDD.n861 0.107922
R16777 VDD.n1245 VDD.n1244 0.107922
R16778 VDD.n1948 VDD.n1947 0.107375
R16779 VDD.n1952 VDD.n1948 0.107375
R16780 VDD.n1856 VDD.n1843 0.104784
R16781 VDD.n1857 VDD.n1856 0.104784
R16782 VDD.n2177 VDD.n2164 0.104784
R16783 VDD.n2178 VDD.n2177 0.104784
R16784 VDD.n2435 VDD.n2422 0.104784
R16785 VDD.n2436 VDD.n2435 0.104784
R16786 VDD.n2693 VDD.n2680 0.104784
R16787 VDD.n2694 VDD.n2693 0.104784
R16788 VDD.n2951 VDD.n2938 0.104784
R16789 VDD.n2952 VDD.n2951 0.104784
R16790 VDD.n3209 VDD.n3196 0.104784
R16791 VDD.n3210 VDD.n3209 0.104784
R16792 VDD.n3467 VDD.n3454 0.104784
R16793 VDD.n3468 VDD.n3467 0.104784
R16794 VDD.n5787 VDD.n5774 0.104784
R16795 VDD.n5788 VDD.n5787 0.104784
R16796 VDD.n5533 VDD.n5520 0.104784
R16797 VDD.n5534 VDD.n5533 0.104784
R16798 VDD.n3725 VDD.n3712 0.104784
R16799 VDD.n3726 VDD.n3725 0.104784
R16800 VDD.n3983 VDD.n3970 0.104784
R16801 VDD.n3984 VDD.n3983 0.104784
R16802 VDD.n4241 VDD.n4228 0.104784
R16803 VDD.n4242 VDD.n4241 0.104784
R16804 VDD.n4499 VDD.n4486 0.104784
R16805 VDD.n4500 VDD.n4499 0.104784
R16806 VDD.n4757 VDD.n4744 0.104784
R16807 VDD.n4758 VDD.n4757 0.104784
R16808 VDD.n5015 VDD.n5002 0.104784
R16809 VDD.n5016 VDD.n5015 0.104784
R16810 VDD.n5273 VDD.n5260 0.104784
R16811 VDD.n5274 VDD.n5273 0.104784
R16812 VDD.n797 VDD.n390 0.102139
R16813 VDD.n1975 VDD.n1974 0.100461
R16814 VDD.n1944 VDD.n1940 0.100461
R16815 VDD.n1974 VDD.n1973 0.0999624
R16816 VDD.n1958 VDD.n1940 0.0999624
R16817 VDD.n1873 VDD.n1842 0.0972991
R16818 VDD.n2194 VDD.n2163 0.0972991
R16819 VDD.n2452 VDD.n2421 0.0972991
R16820 VDD.n2710 VDD.n2679 0.0972991
R16821 VDD.n2968 VDD.n2937 0.0972991
R16822 VDD.n3226 VDD.n3195 0.0972991
R16823 VDD.n3484 VDD.n3453 0.0972991
R16824 VDD.n5804 VDD.n5773 0.0972991
R16825 VDD.n5550 VDD.n5519 0.0972991
R16826 VDD.n3742 VDD.n3711 0.0972991
R16827 VDD.n4000 VDD.n3969 0.0972991
R16828 VDD.n4258 VDD.n4227 0.0972991
R16829 VDD.n4516 VDD.n4485 0.0972991
R16830 VDD.n4774 VDD.n4743 0.0972991
R16831 VDD.n5032 VDD.n5001 0.0972991
R16832 VDD.n5290 VDD.n5259 0.0972991
R16833 VDD.n1811 VDD 0.0963333
R16834 VDD.n2132 VDD 0.0963333
R16835 VDD.n2390 VDD 0.0963333
R16836 VDD.n2648 VDD 0.0963333
R16837 VDD.n2906 VDD 0.0963333
R16838 VDD.n3164 VDD 0.0963333
R16839 VDD.n3422 VDD 0.0963333
R16840 VDD.n5742 VDD 0.0963333
R16841 VDD.n5488 VDD 0.0963333
R16842 VDD.n3680 VDD 0.0963333
R16843 VDD.n3938 VDD 0.0963333
R16844 VDD.n4196 VDD 0.0963333
R16845 VDD.n4454 VDD 0.0963333
R16846 VDD.n4712 VDD 0.0963333
R16847 VDD.n4970 VDD 0.0963333
R16848 VDD.n5228 VDD 0.0963333
R16849 VDD.n1935 VDD.n1934 0.0960166
R16850 VDD.n1936 VDD.n1935 0.095518
R16851 VDD.n853 VDD 0.0950313
R16852 VDD.n1236 VDD 0.0950313
R16853 VDD.n1841 VDD 0.0948131
R16854 VDD.n2162 VDD 0.0948131
R16855 VDD.n2420 VDD 0.0948131
R16856 VDD.n2678 VDD 0.0948131
R16857 VDD.n2936 VDD 0.0948131
R16858 VDD.n3194 VDD 0.0948131
R16859 VDD.n3452 VDD 0.0948131
R16860 VDD.n5772 VDD 0.0948131
R16861 VDD.n5518 VDD 0.0948131
R16862 VDD.n3710 VDD 0.0948131
R16863 VDD.n3968 VDD 0.0948131
R16864 VDD.n4226 VDD 0.0948131
R16865 VDD.n4484 VDD 0.0948131
R16866 VDD.n4742 VDD 0.0948131
R16867 VDD.n5000 VDD 0.0948131
R16868 VDD.n5258 VDD 0.0948131
R16869 VDD.n1875 VDD.n1817 0.0945934
R16870 VDD.n2196 VDD.n2138 0.0945934
R16871 VDD.n2454 VDD.n2396 0.0945934
R16872 VDD.n2712 VDD.n2654 0.0945934
R16873 VDD.n2970 VDD.n2912 0.0945934
R16874 VDD.n3228 VDD.n3170 0.0945934
R16875 VDD.n3486 VDD.n3428 0.0945934
R16876 VDD.n5806 VDD.n5748 0.0945934
R16877 VDD.n5552 VDD.n5494 0.0945934
R16878 VDD.n3744 VDD.n3686 0.0945934
R16879 VDD.n4002 VDD.n3944 0.0945934
R16880 VDD.n4260 VDD.n4202 0.0945934
R16881 VDD.n4518 VDD.n4460 0.0945934
R16882 VDD.n4776 VDD.n4718 0.0945934
R16883 VDD.n5034 VDD.n4976 0.0945934
R16884 VDD.n5292 VDD.n5234 0.0945934
R16885 VDD.n5860 VDD.n1921 0.0944319
R16886 VDD.n5858 VDD.n2242 0.0944319
R16887 VDD.n5857 VDD.n2500 0.0944319
R16888 VDD.n5856 VDD.n2758 0.0944319
R16889 VDD.n5855 VDD.n3016 0.0944319
R16890 VDD.n5854 VDD.n3274 0.0944319
R16891 VDD.n5853 VDD.n3532 0.0944319
R16892 VDD.n5344 VDD.n3790 0.0944319
R16893 VDD.n5343 VDD.n4048 0.0944319
R16894 VDD.n5342 VDD.n4306 0.0944319
R16895 VDD.n5341 VDD.n4564 0.0944319
R16896 VDD.n5340 VDD.n4822 0.0944319
R16897 VDD.n5339 VDD.n5080 0.0944319
R16898 VDD.n1836 VDD 0.0902606
R16899 VDD.n2157 VDD 0.0902606
R16900 VDD.n2415 VDD 0.0902606
R16901 VDD.n2673 VDD 0.0902606
R16902 VDD.n2931 VDD 0.0902606
R16903 VDD.n3189 VDD 0.0902606
R16904 VDD.n3447 VDD 0.0902606
R16905 VDD.n5767 VDD 0.0902606
R16906 VDD.n5513 VDD 0.0902606
R16907 VDD.n3705 VDD 0.0902606
R16908 VDD.n3963 VDD 0.0902606
R16909 VDD.n4221 VDD 0.0902606
R16910 VDD.n4479 VDD 0.0902606
R16911 VDD.n4737 VDD 0.0902606
R16912 VDD.n4995 VDD 0.0902606
R16913 VDD.n5253 VDD 0.0902606
R16914 VDD.n794 VDD 0.0900726
R16915 VDD.n533 VDD.n531 0.0892839
R16916 VDD.n883 VDD.n881 0.0892839
R16917 VDD.n132 VDD.n130 0.0892839
R16918 VDD.n1251 VDD.n1249 0.088354
R16919 VDD.n1797 VDD.n1778 0.0864543
R16920 VDD.n1800 VDD.n1778 0.0864543
R16921 VDD.n2005 VDD.n1986 0.0864543
R16922 VDD.n2008 VDD.n1986 0.0864543
R16923 VDD.n2376 VDD.n2357 0.0864543
R16924 VDD.n2379 VDD.n2357 0.0864543
R16925 VDD.n2634 VDD.n2615 0.0864543
R16926 VDD.n2637 VDD.n2615 0.0864543
R16927 VDD.n2892 VDD.n2873 0.0864543
R16928 VDD.n2895 VDD.n2873 0.0864543
R16929 VDD.n3150 VDD.n3131 0.0864543
R16930 VDD.n3153 VDD.n3131 0.0864543
R16931 VDD.n3408 VDD.n3389 0.0864543
R16932 VDD.n3411 VDD.n3389 0.0864543
R16933 VDD.n5731 VDD.n5712 0.0864543
R16934 VDD.n5734 VDD.n5712 0.0864543
R16935 VDD.n5477 VDD.n5458 0.0864543
R16936 VDD.n5480 VDD.n5458 0.0864543
R16937 VDD.n3666 VDD.n3647 0.0864543
R16938 VDD.n3669 VDD.n3647 0.0864543
R16939 VDD.n3924 VDD.n3905 0.0864543
R16940 VDD.n3927 VDD.n3905 0.0864543
R16941 VDD.n4182 VDD.n4163 0.0864543
R16942 VDD.n4185 VDD.n4163 0.0864543
R16943 VDD.n4440 VDD.n4421 0.0864543
R16944 VDD.n4443 VDD.n4421 0.0864543
R16945 VDD.n4698 VDD.n4679 0.0864543
R16946 VDD.n4701 VDD.n4679 0.0864543
R16947 VDD.n4956 VDD.n4937 0.0864543
R16948 VDD.n4959 VDD.n4937 0.0864543
R16949 VDD.n5214 VDD.n5195 0.0864543
R16950 VDD.n5217 VDD.n5195 0.0864543
R16951 VDD.n5862 VDD.n5861 0.0862917
R16952 VDD.n1774 VDD.n1665 0.0855148
R16953 VDD.n2123 VDD.n2014 0.0855148
R16954 VDD.n2353 VDD.n2244 0.0855148
R16955 VDD.n2611 VDD.n2502 0.0855148
R16956 VDD.n2869 VDD.n2760 0.0855148
R16957 VDD.n3127 VDD.n3018 0.0855148
R16958 VDD.n3385 VDD.n3276 0.0855148
R16959 VDD.n5708 VDD.n5599 0.0855148
R16960 VDD.n5454 VDD.n5345 0.0855148
R16961 VDD.n3643 VDD.n3534 0.0855148
R16962 VDD.n3901 VDD.n3792 0.0855148
R16963 VDD.n4159 VDD.n4050 0.0855148
R16964 VDD.n4417 VDD.n4308 0.0855148
R16965 VDD.n4675 VDD.n4566 0.0855148
R16966 VDD.n4933 VDD.n4824 0.0855148
R16967 VDD.n5191 VDD.n5082 0.0855148
R16968 VDD.n26 VDD.n25 0.0849867
R16969 VDD.n1170 VDD.n1169 0.0849867
R16970 VDD.n5851 VDD.n5709 0.0841827
R16971 VDD.n5597 VDD.n5455 0.0841827
R16972 VDD.n1832 VDD.n1825 0.0832206
R16973 VDD.n2153 VDD.n2146 0.0832206
R16974 VDD.n2411 VDD.n2404 0.0832206
R16975 VDD.n2669 VDD.n2662 0.0832206
R16976 VDD.n2927 VDD.n2920 0.0832206
R16977 VDD.n3185 VDD.n3178 0.0832206
R16978 VDD.n3443 VDD.n3436 0.0832206
R16979 VDD.n5763 VDD.n5756 0.0832206
R16980 VDD.n5509 VDD.n5502 0.0832206
R16981 VDD.n3701 VDD.n3694 0.0832206
R16982 VDD.n3959 VDD.n3952 0.0832206
R16983 VDD.n4217 VDD.n4210 0.0832206
R16984 VDD.n4475 VDD.n4468 0.0832206
R16985 VDD.n4733 VDD.n4726 0.0832206
R16986 VDD.n4991 VDD.n4984 0.0832206
R16987 VDD.n5249 VDD.n5242 0.0832206
R16988 VDD.n1180 VDD.n1143 0.082109
R16989 VDD.n1727 VDD.n1723 0.07913
R16990 VDD.n2076 VDD.n2072 0.07913
R16991 VDD.n2306 VDD.n2302 0.07913
R16992 VDD.n2564 VDD.n2560 0.07913
R16993 VDD.n2822 VDD.n2818 0.07913
R16994 VDD.n3080 VDD.n3076 0.07913
R16995 VDD.n3338 VDD.n3334 0.07913
R16996 VDD.n5661 VDD.n5657 0.07913
R16997 VDD.n5407 VDD.n5403 0.07913
R16998 VDD.n3596 VDD.n3592 0.07913
R16999 VDD.n3854 VDD.n3850 0.07913
R17000 VDD.n4112 VDD.n4108 0.07913
R17001 VDD.n4370 VDD.n4366 0.07913
R17002 VDD.n4628 VDD.n4624 0.07913
R17003 VDD.n4886 VDD.n4882 0.07913
R17004 VDD.n5144 VDD.n5140 0.07913
R17005 VDD.n1835 VDD.n1828 0.078625
R17006 VDD.n2156 VDD.n2149 0.078625
R17007 VDD.n2414 VDD.n2407 0.078625
R17008 VDD.n2672 VDD.n2665 0.078625
R17009 VDD.n2930 VDD.n2923 0.078625
R17010 VDD.n3188 VDD.n3181 0.078625
R17011 VDD.n3446 VDD.n3439 0.078625
R17012 VDD.n5766 VDD.n5759 0.078625
R17013 VDD.n5512 VDD.n5505 0.078625
R17014 VDD.n3704 VDD.n3697 0.078625
R17015 VDD.n3962 VDD.n3955 0.078625
R17016 VDD.n4220 VDD.n4213 0.078625
R17017 VDD.n4478 VDD.n4471 0.078625
R17018 VDD.n4736 VDD.n4729 0.078625
R17019 VDD.n4994 VDD.n4987 0.078625
R17020 VDD.n5252 VDD.n5245 0.078625
R17021 VDD.n33 VDD.n30 0.0777407
R17022 VDD.n1177 VDD.n1174 0.0777407
R17023 VDD.n1748 VDD.n1747 0.0773443
R17024 VDD.n2097 VDD.n2096 0.0773443
R17025 VDD.n2327 VDD.n2326 0.0773443
R17026 VDD.n2585 VDD.n2584 0.0773443
R17027 VDD.n2843 VDD.n2842 0.0773443
R17028 VDD.n3101 VDD.n3100 0.0773443
R17029 VDD.n3359 VDD.n3358 0.0773443
R17030 VDD.n5682 VDD.n5681 0.0773443
R17031 VDD.n5428 VDD.n5427 0.0773443
R17032 VDD.n3617 VDD.n3616 0.0773443
R17033 VDD.n3875 VDD.n3874 0.0773443
R17034 VDD.n4133 VDD.n4132 0.0773443
R17035 VDD.n4391 VDD.n4390 0.0773443
R17036 VDD.n4649 VDD.n4648 0.0773443
R17037 VDD.n4907 VDD.n4906 0.0773443
R17038 VDD.n5165 VDD.n5164 0.0773443
R17039 VDD.n1690 VDD.n1688 0.0755586
R17040 VDD.n2039 VDD.n2037 0.0755586
R17041 VDD.n2269 VDD.n2267 0.0755586
R17042 VDD.n2527 VDD.n2525 0.0755586
R17043 VDD.n2785 VDD.n2783 0.0755586
R17044 VDD.n3043 VDD.n3041 0.0755586
R17045 VDD.n3301 VDD.n3299 0.0755586
R17046 VDD.n5624 VDD.n5622 0.0755586
R17047 VDD.n5370 VDD.n5368 0.0755586
R17048 VDD.n3559 VDD.n3557 0.0755586
R17049 VDD.n3817 VDD.n3815 0.0755586
R17050 VDD.n4075 VDD.n4073 0.0755586
R17051 VDD.n4333 VDD.n4331 0.0755586
R17052 VDD.n4591 VDD.n4589 0.0755586
R17053 VDD.n4849 VDD.n4847 0.0755586
R17054 VDD.n5107 VDD.n5105 0.0755586
R17055 VDD.n510 VDD.n507 0.0734782
R17056 VDD.n437 VDD.n434 0.0734782
R17057 VDD.n108 VDD.n105 0.0734782
R17058 VDD.n1595 VDD.n1592 0.0734782
R17059 VDD.n1842 VDD.n1841 0.0710611
R17060 VDD.n2163 VDD.n2162 0.0710611
R17061 VDD.n2421 VDD.n2420 0.0710611
R17062 VDD.n2679 VDD.n2678 0.0710611
R17063 VDD.n2937 VDD.n2936 0.0710611
R17064 VDD.n3195 VDD.n3194 0.0710611
R17065 VDD.n3453 VDD.n3452 0.0710611
R17066 VDD.n5773 VDD.n5772 0.0710611
R17067 VDD.n5519 VDD.n5518 0.0710611
R17068 VDD.n3711 VDD.n3710 0.0710611
R17069 VDD.n3969 VDD.n3968 0.0710611
R17070 VDD.n4227 VDD.n4226 0.0710611
R17071 VDD.n4485 VDD.n4484 0.0710611
R17072 VDD.n4743 VDD.n4742 0.0710611
R17073 VDD.n5001 VDD.n5000 0.0710611
R17074 VDD.n5259 VDD.n5258 0.0710611
R17075 VDD.n1919 VDD.n1816 0.0705353
R17076 VDD.n2240 VDD.n2137 0.0705353
R17077 VDD.n2498 VDD.n2395 0.0705353
R17078 VDD.n2756 VDD.n2653 0.0705353
R17079 VDD.n3014 VDD.n2911 0.0705353
R17080 VDD.n3272 VDD.n3169 0.0705353
R17081 VDD.n3530 VDD.n3427 0.0705353
R17082 VDD.n5850 VDD.n5747 0.0705353
R17083 VDD.n5596 VDD.n5493 0.0705353
R17084 VDD.n3788 VDD.n3685 0.0705353
R17085 VDD.n4046 VDD.n3943 0.0705353
R17086 VDD.n4304 VDD.n4201 0.0705353
R17087 VDD.n4562 VDD.n4459 0.0705353
R17088 VDD.n4820 VDD.n4717 0.0705353
R17089 VDD.n5078 VDD.n4975 0.0705353
R17090 VDD.n5336 VDD.n5233 0.0705353
R17091 VDD.n1846 VDD.n1845 0.0694784
R17092 VDD.n1849 VDD.n1846 0.0694784
R17093 VDD.n2167 VDD.n2166 0.0694784
R17094 VDD.n2170 VDD.n2167 0.0694784
R17095 VDD.n2425 VDD.n2424 0.0694784
R17096 VDD.n2428 VDD.n2425 0.0694784
R17097 VDD.n2683 VDD.n2682 0.0694784
R17098 VDD.n2686 VDD.n2683 0.0694784
R17099 VDD.n2941 VDD.n2940 0.0694784
R17100 VDD.n2944 VDD.n2941 0.0694784
R17101 VDD.n3199 VDD.n3198 0.0694784
R17102 VDD.n3202 VDD.n3199 0.0694784
R17103 VDD.n3457 VDD.n3456 0.0694784
R17104 VDD.n3460 VDD.n3457 0.0694784
R17105 VDD.n5777 VDD.n5776 0.0694784
R17106 VDD.n5780 VDD.n5777 0.0694784
R17107 VDD.n5523 VDD.n5522 0.0694784
R17108 VDD.n5526 VDD.n5523 0.0694784
R17109 VDD.n3715 VDD.n3714 0.0694784
R17110 VDD.n3718 VDD.n3715 0.0694784
R17111 VDD.n3973 VDD.n3972 0.0694784
R17112 VDD.n3976 VDD.n3973 0.0694784
R17113 VDD.n4231 VDD.n4230 0.0694784
R17114 VDD.n4234 VDD.n4231 0.0694784
R17115 VDD.n4489 VDD.n4488 0.0694784
R17116 VDD.n4492 VDD.n4489 0.0694784
R17117 VDD.n4747 VDD.n4746 0.0694784
R17118 VDD.n4750 VDD.n4747 0.0694784
R17119 VDD.n5005 VDD.n5004 0.0694784
R17120 VDD.n5008 VDD.n5005 0.0694784
R17121 VDD.n5263 VDD.n5262 0.0694784
R17122 VDD.n5266 VDD.n5263 0.0694784
R17123 VDD.n458 VDD.n457 0.0681471
R17124 VDD.n457 VDD.n454 0.0681471
R17125 VDD.n454 VDD.n451 0.0681471
R17126 VDD.n451 VDD.n450 0.0681471
R17127 VDD.n450 VDD.n447 0.0681471
R17128 VDD.n55 VDD.n54 0.0681471
R17129 VDD.n54 VDD.n51 0.0681471
R17130 VDD.n51 VDD.n48 0.0681471
R17131 VDD.n48 VDD.n47 0.0681471
R17132 VDD.n47 VDD.n44 0.0681471
R17133 VDD.n406 VDD.n403 0.0671334
R17134 VDD.n1564 VDD.n1561 0.0671334
R17135 VDD.n22 VDD.n21 0.065907
R17136 VDD.n17 VDD.n4 0.065907
R17137 VDD.n16 VDD.n15 0.065907
R17138 VDD.n14 VDD.n10 0.065907
R17139 VDD.n1166 VDD.n1165 0.065907
R17140 VDD.n1161 VDD.n1148 0.065907
R17141 VDD.n1160 VDD.n1159 0.065907
R17142 VDD.n1158 VDD.n1154 0.065907
R17143 VDD.n480 VDD.n479 0.0658409
R17144 VDD.n78 VDD.n77 0.0658409
R17145 VDD.n5739 VDD 0.0644514
R17146 VDD.n5485 VDD 0.0644514
R17147 VDD.n1791 VDD.n1783 0.0643889
R17148 VDD.n1791 VDD.n1780 0.0643889
R17149 VDD.n1796 VDD.n1780 0.0643889
R17150 VDD.n1999 VDD.n1991 0.0643889
R17151 VDD.n1999 VDD.n1988 0.0643889
R17152 VDD.n2004 VDD.n1988 0.0643889
R17153 VDD.n2370 VDD.n2362 0.0643889
R17154 VDD.n2370 VDD.n2359 0.0643889
R17155 VDD.n2375 VDD.n2359 0.0643889
R17156 VDD.n2628 VDD.n2620 0.0643889
R17157 VDD.n2628 VDD.n2617 0.0643889
R17158 VDD.n2633 VDD.n2617 0.0643889
R17159 VDD.n2886 VDD.n2878 0.0643889
R17160 VDD.n2886 VDD.n2875 0.0643889
R17161 VDD.n2891 VDD.n2875 0.0643889
R17162 VDD.n3144 VDD.n3136 0.0643889
R17163 VDD.n3144 VDD.n3133 0.0643889
R17164 VDD.n3149 VDD.n3133 0.0643889
R17165 VDD.n3402 VDD.n3394 0.0643889
R17166 VDD.n3402 VDD.n3391 0.0643889
R17167 VDD.n3407 VDD.n3391 0.0643889
R17168 VDD.n5725 VDD.n5717 0.0643889
R17169 VDD.n5725 VDD.n5714 0.0643889
R17170 VDD.n5730 VDD.n5714 0.0643889
R17171 VDD.n5471 VDD.n5463 0.0643889
R17172 VDD.n5471 VDD.n5460 0.0643889
R17173 VDD.n5476 VDD.n5460 0.0643889
R17174 VDD.n3660 VDD.n3652 0.0643889
R17175 VDD.n3660 VDD.n3649 0.0643889
R17176 VDD.n3665 VDD.n3649 0.0643889
R17177 VDD.n3918 VDD.n3910 0.0643889
R17178 VDD.n3918 VDD.n3907 0.0643889
R17179 VDD.n3923 VDD.n3907 0.0643889
R17180 VDD.n4176 VDD.n4168 0.0643889
R17181 VDD.n4176 VDD.n4165 0.0643889
R17182 VDD.n4181 VDD.n4165 0.0643889
R17183 VDD.n4434 VDD.n4426 0.0643889
R17184 VDD.n4434 VDD.n4423 0.0643889
R17185 VDD.n4439 VDD.n4423 0.0643889
R17186 VDD.n4692 VDD.n4684 0.0643889
R17187 VDD.n4692 VDD.n4681 0.0643889
R17188 VDD.n4697 VDD.n4681 0.0643889
R17189 VDD.n4950 VDD.n4942 0.0643889
R17190 VDD.n4950 VDD.n4939 0.0643889
R17191 VDD.n4955 VDD.n4939 0.0643889
R17192 VDD.n5208 VDD.n5200 0.0643889
R17193 VDD.n5208 VDD.n5197 0.0643889
R17194 VDD.n5213 VDD.n5197 0.0643889
R17195 VDD.n507 VDD.n505 0.0643889
R17196 VDD.n505 VDD.n503 0.0643889
R17197 VDD.n503 VDD.n501 0.0643889
R17198 VDD.n498 VDD.n497 0.0643889
R17199 VDD.n497 VDD.n493 0.0643889
R17200 VDD.n493 VDD.n491 0.0643889
R17201 VDD.n486 VDD.n485 0.0643889
R17202 VDD.n434 VDD.n432 0.0643889
R17203 VDD.n432 VDD.n430 0.0643889
R17204 VDD.n430 VDD.n428 0.0643889
R17205 VDD.n421 VDD.n417 0.0643889
R17206 VDD.n417 VDD.n415 0.0643889
R17207 VDD.n415 VDD.n413 0.0643889
R17208 VDD.n400 VDD.n398 0.0643889
R17209 VDD.n398 VDD.n396 0.0643889
R17210 VDD.n105 VDD.n103 0.0643889
R17211 VDD.n103 VDD.n101 0.0643889
R17212 VDD.n101 VDD.n99 0.0643889
R17213 VDD.n96 VDD.n95 0.0643889
R17214 VDD.n95 VDD.n91 0.0643889
R17215 VDD.n91 VDD.n89 0.0643889
R17216 VDD.n84 VDD.n83 0.0643889
R17217 VDD.n1592 VDD.n1590 0.0643889
R17218 VDD.n1590 VDD.n1588 0.0643889
R17219 VDD.n1588 VDD.n1586 0.0643889
R17220 VDD.n1579 VDD.n1575 0.0643889
R17221 VDD.n1575 VDD.n1573 0.0643889
R17222 VDD.n1573 VDD.n1571 0.0643889
R17223 VDD.n1558 VDD.n1556 0.0643889
R17224 VDD.n1556 VDD.n1554 0.0643889
R17225 VDD.n1526 VDD 0.0639804
R17226 VDD.n1806 VDD 0.0630006
R17227 VDD.n2126 VDD 0.0630006
R17228 VDD.n2385 VDD 0.0630006
R17229 VDD.n2643 VDD 0.0630006
R17230 VDD.n2901 VDD 0.0630006
R17231 VDD.n3159 VDD 0.0630006
R17232 VDD.n3417 VDD 0.0630006
R17233 VDD.n3675 VDD 0.0630006
R17234 VDD.n3933 VDD 0.0630006
R17235 VDD.n4191 VDD 0.0630006
R17236 VDD.n4449 VDD 0.0630006
R17237 VDD.n4707 VDD 0.0630006
R17238 VDD.n4965 VDD 0.0630006
R17239 VDD.n5223 VDD 0.0630006
R17240 VDD.n1623 VDD 0.0604792
R17241 VDD.n462 VDD.n461 0.0599867
R17242 VDD.n59 VDD.n58 0.0599867
R17243 VDD.n1772 VDD.n1667 0.0588333
R17244 VDD.n2121 VDD.n2016 0.0588333
R17245 VDD.n2351 VDD.n2246 0.0588333
R17246 VDD.n2609 VDD.n2504 0.0588333
R17247 VDD.n2867 VDD.n2762 0.0588333
R17248 VDD.n3125 VDD.n3020 0.0588333
R17249 VDD.n3383 VDD.n3278 0.0588333
R17250 VDD.n5706 VDD.n5601 0.0588333
R17251 VDD.n5452 VDD.n5347 0.0588333
R17252 VDD.n3641 VDD.n3536 0.0588333
R17253 VDD.n3899 VDD.n3794 0.0588333
R17254 VDD.n4157 VDD.n4052 0.0588333
R17255 VDD.n4415 VDD.n4310 0.0588333
R17256 VDD.n4673 VDD.n4568 0.0588333
R17257 VDD.n4931 VDD.n4826 0.0588333
R17258 VDD.n5189 VDD.n5084 0.0588333
R17259 VDD.n395 VDD.n394 0.0587674
R17260 VDD.n1553 VDD.n1552 0.0587674
R17261 VDD.n425 VDD.n424 0.0580441
R17262 VDD.n1583 VDD.n1582 0.0580441
R17263 VDD.n848 VDD 0.058
R17264 VDD.n842 VDD 0.058
R17265 VDD.n830 VDD 0.058
R17266 VDD.n1231 VDD 0.058
R17267 VDD.n1225 VDD 0.058
R17268 VDD.n1213 VDD 0.058
R17269 VDD.n491 VDD.n489 0.0567153
R17270 VDD.n89 VDD.n87 0.0567153
R17271 VDD.n5863 VDD.n5862 0.0560833
R17272 VDD.n836 VDD 0.0555
R17273 VDD.n1219 VDD 0.0555
R17274 VDD.n5852 VDD.n5851 0.0554144
R17275 VDD.n5598 VDD.n5597 0.0554144
R17276 VDD VDD.n5860 0.0546184
R17277 VDD VDD.n1783 0.0525833
R17278 VDD VDD.n1991 0.0525833
R17279 VDD VDD.n2362 0.0525833
R17280 VDD VDD.n2620 0.0525833
R17281 VDD VDD.n2878 0.0525833
R17282 VDD VDD.n3136 0.0525833
R17283 VDD VDD.n3394 0.0525833
R17284 VDD VDD.n5717 0.0525833
R17285 VDD VDD.n5463 0.0525833
R17286 VDD VDD.n3652 0.0525833
R17287 VDD VDD.n3910 0.0525833
R17288 VDD VDD.n4168 0.0525833
R17289 VDD VDD.n4426 0.0525833
R17290 VDD VDD.n4684 0.0525833
R17291 VDD VDD.n4942 0.0525833
R17292 VDD VDD.n5200 0.0525833
R17293 VDD.n481 VDD.n480 0.0516364
R17294 VDD.n79 VDD.n78 0.0516364
R17295 VDD.n1799 VDD 0.0470278
R17296 VDD.n2007 VDD 0.0470278
R17297 VDD.n2378 VDD 0.0470278
R17298 VDD.n2636 VDD 0.0470278
R17299 VDD.n2894 VDD 0.0470278
R17300 VDD.n3152 VDD 0.0470278
R17301 VDD.n3410 VDD 0.0470278
R17302 VDD.n5733 VDD 0.0470278
R17303 VDD.n5479 VDD 0.0470278
R17304 VDD.n3668 VDD 0.0470278
R17305 VDD.n3926 VDD 0.0470278
R17306 VDD.n4184 VDD 0.0470278
R17307 VDD.n4442 VDD 0.0470278
R17308 VDD.n4700 VDD 0.0470278
R17309 VDD.n4958 VDD 0.0470278
R17310 VDD.n5216 VDD 0.0470278
R17311 VDD.n5852 VDD.n5598 0.0430009
R17312 VDD.n5853 VDD.n5852 0.0425691
R17313 VDD.n5598 VDD.n5344 0.0421424
R17314 VDD.n25 VDD.n0 0.0418891
R17315 VDD.n1169 VDD.n1144 0.0418891
R17316 VDD.n5858 VDD.n5857 0.0417105
R17317 VDD.n5857 VDD.n5856 0.0417105
R17318 VDD.n5856 VDD.n5855 0.0417105
R17319 VDD.n5855 VDD.n5854 0.0417105
R17320 VDD.n5854 VDD.n5853 0.0417105
R17321 VDD.n5344 VDD.n5343 0.0417105
R17322 VDD.n5343 VDD.n5342 0.0417105
R17323 VDD.n5342 VDD.n5341 0.0417105
R17324 VDD.n5341 VDD.n5340 0.0417105
R17325 VDD.n5340 VDD.n5339 0.0417105
R17326 VDD.n1832 VDD.n1831 0.0409412
R17327 VDD.n2153 VDD.n2152 0.0409412
R17328 VDD.n2411 VDD.n2410 0.0409412
R17329 VDD.n2669 VDD.n2668 0.0409412
R17330 VDD.n2927 VDD.n2926 0.0409412
R17331 VDD.n3185 VDD.n3184 0.0409412
R17332 VDD.n3443 VDD.n3442 0.0409412
R17333 VDD.n5763 VDD.n5762 0.0409412
R17334 VDD.n5509 VDD.n5508 0.0409412
R17335 VDD.n3701 VDD.n3700 0.0409412
R17336 VDD.n3959 VDD.n3958 0.0409412
R17337 VDD.n4217 VDD.n4216 0.0409412
R17338 VDD.n4475 VDD.n4474 0.0409412
R17339 VDD.n4733 VDD.n4732 0.0409412
R17340 VDD.n4991 VDD.n4990 0.0409412
R17341 VDD.n5249 VDD.n5248 0.0409412
R17342 VDD.n30 VDD.n28 0.0409412
R17343 VDD.n1174 VDD.n1172 0.0409412
R17344 VDD.n5709 VDD.n5708 0.0399318
R17345 VDD.n5455 VDD.n5454 0.0399318
R17346 VDD.n5860 VDD.n5859 0.0398026
R17347 VDD.n820 VDD.n799 0.03976
R17348 VDD.n1203 VDD.n1182 0.03976
R17349 VDD.n1797 VDD.n1776 0.0395625
R17350 VDD.n2005 VDD.n1984 0.0395625
R17351 VDD.n2376 VDD.n2355 0.0395625
R17352 VDD.n2634 VDD.n2613 0.0395625
R17353 VDD.n2892 VDD.n2871 0.0395625
R17354 VDD.n3150 VDD.n3129 0.0395625
R17355 VDD.n3408 VDD.n3387 0.0395625
R17356 VDD.n5731 VDD.n5710 0.0395625
R17357 VDD.n5477 VDD.n5456 0.0395625
R17358 VDD.n3666 VDD.n3645 0.0395625
R17359 VDD.n3924 VDD.n3903 0.0395625
R17360 VDD.n4182 VDD.n4161 0.0395625
R17361 VDD.n4440 VDD.n4419 0.0395625
R17362 VDD.n4698 VDD.n4677 0.0395625
R17363 VDD.n4956 VDD.n4935 0.0395625
R17364 VDD.n5214 VDD.n5193 0.0395625
R17365 VDD.n797 VDD 0.0390887
R17366 VDD.n854 VDD.n853 0.0376094
R17367 VDD.n1237 VDD.n1236 0.0376094
R17368 VDD.n1836 VDD.n1835 0.0372647
R17369 VDD.n2157 VDD.n2156 0.0372647
R17370 VDD.n2415 VDD.n2414 0.0372647
R17371 VDD.n2673 VDD.n2672 0.0372647
R17372 VDD.n2931 VDD.n2930 0.0372647
R17373 VDD.n3189 VDD.n3188 0.0372647
R17374 VDD.n3447 VDD.n3446 0.0372647
R17375 VDD.n5767 VDD.n5766 0.0372647
R17376 VDD.n5513 VDD.n5512 0.0372647
R17377 VDD.n3705 VDD.n3704 0.0372647
R17378 VDD.n3963 VDD.n3962 0.0372647
R17379 VDD.n4221 VDD.n4220 0.0372647
R17380 VDD.n4479 VDD.n4478 0.0372647
R17381 VDD.n4737 VDD.n4736 0.0372647
R17382 VDD.n4995 VDD.n4994 0.0372647
R17383 VDD.n5253 VDD.n5252 0.0372647
R17384 VDD.n28 VDD.n27 0.0371297
R17385 VDD.n1172 VDD.n1171 0.0371297
R17386 VDD.n1701 VDD.n1665 0.0364409
R17387 VDD.n2050 VDD.n2014 0.0364409
R17388 VDD.n2280 VDD.n2244 0.0364409
R17389 VDD.n2538 VDD.n2502 0.0364409
R17390 VDD.n2796 VDD.n2760 0.0364409
R17391 VDD.n3054 VDD.n3018 0.0364409
R17392 VDD.n3312 VDD.n3276 0.0364409
R17393 VDD.n5635 VDD.n5599 0.0364409
R17394 VDD.n5381 VDD.n5345 0.0364409
R17395 VDD.n3570 VDD.n3534 0.0364409
R17396 VDD.n3828 VDD.n3792 0.0364409
R17397 VDD.n4086 VDD.n4050 0.0364409
R17398 VDD.n4344 VDD.n4308 0.0364409
R17399 VDD.n4602 VDD.n4566 0.0364409
R17400 VDD.n4860 VDD.n4824 0.0364409
R17401 VDD.n5118 VDD.n5082 0.0364409
R17402 VDD.n1837 VDD.n1836 0.0361152
R17403 VDD.n2158 VDD.n2157 0.0361152
R17404 VDD.n2416 VDD.n2415 0.0361152
R17405 VDD.n2674 VDD.n2673 0.0361152
R17406 VDD.n2932 VDD.n2931 0.0361152
R17407 VDD.n3190 VDD.n3189 0.0361152
R17408 VDD.n3448 VDD.n3447 0.0361152
R17409 VDD.n5768 VDD.n5767 0.0361152
R17410 VDD.n5514 VDD.n5513 0.0361152
R17411 VDD.n3706 VDD.n3705 0.0361152
R17412 VDD.n3964 VDD.n3963 0.0361152
R17413 VDD.n4222 VDD.n4221 0.0361152
R17414 VDD.n4480 VDD.n4479 0.0361152
R17415 VDD.n4738 VDD.n4737 0.0361152
R17416 VDD.n4996 VDD.n4995 0.0361152
R17417 VDD.n5254 VDD.n5253 0.0361152
R17418 VDD.n1752 VDD.n1751 0.0357224
R17419 VDD.n2101 VDD.n2100 0.0357224
R17420 VDD.n2331 VDD.n2330 0.0357224
R17421 VDD.n2589 VDD.n2588 0.0357224
R17422 VDD.n2847 VDD.n2846 0.0357224
R17423 VDD.n3105 VDD.n3104 0.0357224
R17424 VDD.n3363 VDD.n3362 0.0357224
R17425 VDD.n5686 VDD.n5685 0.0357224
R17426 VDD.n5432 VDD.n5431 0.0357224
R17427 VDD.n3621 VDD.n3620 0.0357224
R17428 VDD.n3879 VDD.n3878 0.0357224
R17429 VDD.n4137 VDD.n4136 0.0357224
R17430 VDD.n4395 VDD.n4394 0.0357224
R17431 VDD.n4653 VDD.n4652 0.0357224
R17432 VDD.n4911 VDD.n4910 0.0357224
R17433 VDD.n5169 VDD.n5168 0.0357224
R17434 VDD.n1684 VDD.n1683 0.034445
R17435 VDD.n2033 VDD.n2032 0.034445
R17436 VDD.n2263 VDD.n2262 0.034445
R17437 VDD.n2521 VDD.n2520 0.034445
R17438 VDD.n2779 VDD.n2778 0.034445
R17439 VDD.n3037 VDD.n3036 0.034445
R17440 VDD.n3295 VDD.n3294 0.034445
R17441 VDD.n5618 VDD.n5617 0.034445
R17442 VDD.n5364 VDD.n5363 0.034445
R17443 VDD.n3553 VDD.n3552 0.034445
R17444 VDD.n3811 VDD.n3810 0.034445
R17445 VDD.n4069 VDD.n4068 0.034445
R17446 VDD.n4327 VDD.n4326 0.034445
R17447 VDD.n4585 VDD.n4584 0.034445
R17448 VDD.n4843 VDD.n4842 0.034445
R17449 VDD.n5101 VDD.n5100 0.034445
R17450 VDD.n3 VDD.n0 0.0339302
R17451 VDD.n1147 VDD.n1144 0.0339302
R17452 VDD.n810 VDD.n802 0.033737
R17453 VDD.n814 VDD.n802 0.033737
R17454 VDD.n815 VDD.n814 0.033737
R17455 VDD.n816 VDD.n815 0.033737
R17456 VDD.n1193 VDD.n1185 0.033737
R17457 VDD.n1197 VDD.n1185 0.033737
R17458 VDD.n1198 VDD.n1197 0.033737
R17459 VDD.n1199 VDD.n1198 0.033737
R17460 VDD.n479 VDD.n477 0.0334425
R17461 VDD.n477 VDD.n474 0.0334425
R17462 VDD.n77 VDD.n75 0.0334425
R17463 VDD.n75 VDD.n72 0.0334425
R17464 VDD.n1548 VDD.n1547 0.0333707
R17465 VDD.n863 VDD.n798 0.0325611
R17466 VDD VDD.n1796 0.0324444
R17467 VDD VDD.n2004 0.0324444
R17468 VDD VDD.n2375 0.0324444
R17469 VDD VDD.n2633 0.0324444
R17470 VDD VDD.n2891 0.0324444
R17471 VDD VDD.n3149 0.0324444
R17472 VDD VDD.n3407 0.0324444
R17473 VDD VDD.n5730 0.0324444
R17474 VDD VDD.n5476 0.0324444
R17475 VDD VDD.n3665 0.0324444
R17476 VDD VDD.n3923 0.0324444
R17477 VDD VDD.n4181 0.0324444
R17478 VDD VDD.n4439 0.0324444
R17479 VDD VDD.n4697 0.0324444
R17480 VDD VDD.n4955 0.0324444
R17481 VDD VDD.n5213 0.0324444
R17482 VDD.n498 VDD 0.0324444
R17483 VDD.n486 VDD 0.0324444
R17484 VDD.n425 VDD 0.0324444
R17485 VDD.n96 VDD 0.0324444
R17486 VDD.n84 VDD 0.0324444
R17487 VDD.n1583 VDD 0.0324444
R17488 VDD.n1640 VDD.n1639 0.0308571
R17489 VDD.n110 VDD.n62 0.0299677
R17490 VDD.n798 VDD.n110 0.0299677
R17491 VDD.n513 VDD.n512 0.0299677
R17492 VDD.n1771 VDD.n1770 0.0294474
R17493 VDD.n2120 VDD.n2119 0.0294474
R17494 VDD.n2350 VDD.n2349 0.0294474
R17495 VDD.n2608 VDD.n2607 0.0294474
R17496 VDD.n2866 VDD.n2865 0.0294474
R17497 VDD.n3124 VDD.n3123 0.0294474
R17498 VDD.n3382 VDD.n3381 0.0294474
R17499 VDD.n5705 VDD.n5704 0.0294474
R17500 VDD.n5451 VDD.n5450 0.0294474
R17501 VDD.n3640 VDD.n3639 0.0294474
R17502 VDD.n3898 VDD.n3897 0.0294474
R17503 VDD.n4156 VDD.n4155 0.0294474
R17504 VDD.n4414 VDD.n4413 0.0294474
R17505 VDD.n4672 VDD.n4671 0.0294474
R17506 VDD.n4930 VDD.n4929 0.0294474
R17507 VDD.n5188 VDD.n5187 0.0294474
R17508 VDD.n1598 VDD.n1597 0.0292661
R17509 VDD.n796 VDD.n795 0.0292661
R17510 VDD.n1754 VDD.n1753 0.0287895
R17511 VDD.n2103 VDD.n2102 0.0287895
R17512 VDD.n2333 VDD.n2332 0.0287895
R17513 VDD.n2591 VDD.n2590 0.0287895
R17514 VDD.n2849 VDD.n2848 0.0287895
R17515 VDD.n3107 VDD.n3106 0.0287895
R17516 VDD.n3365 VDD.n3364 0.0287895
R17517 VDD.n5688 VDD.n5687 0.0287895
R17518 VDD.n5434 VDD.n5433 0.0287895
R17519 VDD.n3623 VDD.n3622 0.0287895
R17520 VDD.n3881 VDD.n3880 0.0287895
R17521 VDD.n4139 VDD.n4138 0.0287895
R17522 VDD.n4397 VDD.n4396 0.0287895
R17523 VDD.n4655 VDD.n4654 0.0287895
R17524 VDD.n4913 VDD.n4912 0.0287895
R17525 VDD.n5171 VDD.n5170 0.0287895
R17526 VDD.n1750 VDD.n1720 0.0282778
R17527 VDD.n2099 VDD.n2069 0.0282778
R17528 VDD.n2329 VDD.n2299 0.0282778
R17529 VDD.n2587 VDD.n2557 0.0282778
R17530 VDD.n2845 VDD.n2815 0.0282778
R17531 VDD.n3103 VDD.n3073 0.0282778
R17532 VDD.n3361 VDD.n3331 0.0282778
R17533 VDD.n5684 VDD.n5654 0.0282778
R17534 VDD.n5430 VDD.n5400 0.0282778
R17535 VDD.n3619 VDD.n3589 0.0282778
R17536 VDD.n3877 VDD.n3847 0.0282778
R17537 VDD.n4135 VDD.n4105 0.0282778
R17538 VDD.n4393 VDD.n4363 0.0282778
R17539 VDD.n4651 VDD.n4621 0.0282778
R17540 VDD.n4909 VDD.n4879 0.0282778
R17541 VDD.n5167 VDD.n5137 0.0282778
R17542 VDD.t1014 VDD.n1763 0.0282694
R17543 VDD.n1763 VDD.n1762 0.0282694
R17544 VDD.t1014 VDD.n1677 0.0282694
R17545 VDD.n1706 VDD.n1677 0.0282694
R17546 VDD.t623 VDD.n2112 0.0282694
R17547 VDD.n2112 VDD.n2111 0.0282694
R17548 VDD.t623 VDD.n2026 0.0282694
R17549 VDD.n2055 VDD.n2026 0.0282694
R17550 VDD.t1331 VDD.n2342 0.0282694
R17551 VDD.n2342 VDD.n2341 0.0282694
R17552 VDD.t1331 VDD.n2256 0.0282694
R17553 VDD.n2285 VDD.n2256 0.0282694
R17554 VDD.t825 VDD.n2600 0.0282694
R17555 VDD.n2600 VDD.n2599 0.0282694
R17556 VDD.t825 VDD.n2514 0.0282694
R17557 VDD.n2543 VDD.n2514 0.0282694
R17558 VDD.t424 VDD.n2858 0.0282694
R17559 VDD.n2858 VDD.n2857 0.0282694
R17560 VDD.t424 VDD.n2772 0.0282694
R17561 VDD.n2801 VDD.n2772 0.0282694
R17562 VDD.t395 VDD.n3116 0.0282694
R17563 VDD.n3116 VDD.n3115 0.0282694
R17564 VDD.t395 VDD.n3030 0.0282694
R17565 VDD.n3059 VDD.n3030 0.0282694
R17566 VDD.t639 VDD.n3374 0.0282694
R17567 VDD.n3374 VDD.n3373 0.0282694
R17568 VDD.t639 VDD.n3288 0.0282694
R17569 VDD.n3317 VDD.n3288 0.0282694
R17570 VDD.t1307 VDD.n5697 0.0282694
R17571 VDD.n5697 VDD.n5696 0.0282694
R17572 VDD.t1307 VDD.n5611 0.0282694
R17573 VDD.n5640 VDD.n5611 0.0282694
R17574 VDD.t270 VDD.n5443 0.0282694
R17575 VDD.n5443 VDD.n5442 0.0282694
R17576 VDD.t270 VDD.n5357 0.0282694
R17577 VDD.n5386 VDD.n5357 0.0282694
R17578 VDD.t249 VDD.n3632 0.0282694
R17579 VDD.n3632 VDD.n3631 0.0282694
R17580 VDD.t249 VDD.n3546 0.0282694
R17581 VDD.n3575 VDD.n3546 0.0282694
R17582 VDD.t1317 VDD.n3890 0.0282694
R17583 VDD.n3890 VDD.n3889 0.0282694
R17584 VDD.t1317 VDD.n3804 0.0282694
R17585 VDD.n3833 VDD.n3804 0.0282694
R17586 VDD.t409 VDD.n4148 0.0282694
R17587 VDD.n4148 VDD.n4147 0.0282694
R17588 VDD.t409 VDD.n4062 0.0282694
R17589 VDD.n4091 VDD.n4062 0.0282694
R17590 VDD.t1108 VDD.n4406 0.0282694
R17591 VDD.n4406 VDD.n4405 0.0282694
R17592 VDD.t1108 VDD.n4320 0.0282694
R17593 VDD.n4349 VDD.n4320 0.0282694
R17594 VDD.t332 VDD.n4664 0.0282694
R17595 VDD.n4664 VDD.n4663 0.0282694
R17596 VDD.t332 VDD.n4578 0.0282694
R17597 VDD.n4607 VDD.n4578 0.0282694
R17598 VDD.t279 VDD.n4922 0.0282694
R17599 VDD.n4922 VDD.n4921 0.0282694
R17600 VDD.t279 VDD.n4836 0.0282694
R17601 VDD.n4865 VDD.n4836 0.0282694
R17602 VDD.t1060 VDD.n5180 0.0282694
R17603 VDD.n5180 VDD.n5179 0.0282694
R17604 VDD.t1060 VDD.n5094 0.0282694
R17605 VDD.n5123 VDD.n5094 0.0282694
R17606 VDD.n674 VDD 0.0279106
R17607 VDD.n1024 VDD 0.0279106
R17608 VDD.n269 VDD 0.0279106
R17609 VDD.n1897 VDD.n1895 0.0265784
R17610 VDD.n1905 VDD.n1895 0.0265784
R17611 VDD.n1911 VDD.n1896 0.0265784
R17612 VDD.n1901 VDD.n1896 0.0265784
R17613 VDD.n1903 VDD.n1902 0.0265784
R17614 VDD.n1902 VDD.n1901 0.0265784
R17615 VDD.n1907 VDD.n1906 0.0265784
R17616 VDD.n1906 VDD.n1905 0.0265784
R17617 VDD.n1878 VDD.n1877 0.0265784
R17618 VDD.t274 VDD.n1878 0.0265784
R17619 VDD.n1880 VDD.n1822 0.0265784
R17620 VDD.n1860 VDD.n1859 0.0265784
R17621 VDD.n1859 VDD.n1858 0.0265784
R17622 VDD.n1862 VDD.n1853 0.0265784
R17623 VDD.n1863 VDD.n1862 0.0265784
R17624 VDD.n1865 VDD.n1864 0.0265784
R17625 VDD.n1864 VDD.n1863 0.0265784
R17626 VDD.n1858 VDD.n1855 0.0265784
R17627 VDD.n1855 VDD.n1854 0.0265784
R17628 VDD.n2181 VDD.n2180 0.0265784
R17629 VDD.n2180 VDD.n2179 0.0265784
R17630 VDD.n2183 VDD.n2174 0.0265784
R17631 VDD.n2184 VDD.n2183 0.0265784
R17632 VDD.n2186 VDD.n2185 0.0265784
R17633 VDD.n2185 VDD.n2184 0.0265784
R17634 VDD.n2179 VDD.n2176 0.0265784
R17635 VDD.n2176 VDD.n2175 0.0265784
R17636 VDD.n2199 VDD.n2198 0.0265784
R17637 VDD.t511 VDD.n2199 0.0265784
R17638 VDD.n2201 VDD.n2143 0.0265784
R17639 VDD.n2218 VDD.n2216 0.0265784
R17640 VDD.n2226 VDD.n2216 0.0265784
R17641 VDD.n2232 VDD.n2217 0.0265784
R17642 VDD.n2222 VDD.n2217 0.0265784
R17643 VDD.n2224 VDD.n2223 0.0265784
R17644 VDD.n2223 VDD.n2222 0.0265784
R17645 VDD.n2228 VDD.n2227 0.0265784
R17646 VDD.n2227 VDD.n2226 0.0265784
R17647 VDD.n2439 VDD.n2438 0.0265784
R17648 VDD.n2438 VDD.n2437 0.0265784
R17649 VDD.n2441 VDD.n2432 0.0265784
R17650 VDD.n2442 VDD.n2441 0.0265784
R17651 VDD.n2444 VDD.n2443 0.0265784
R17652 VDD.n2443 VDD.n2442 0.0265784
R17653 VDD.n2437 VDD.n2434 0.0265784
R17654 VDD.n2434 VDD.n2433 0.0265784
R17655 VDD.n2457 VDD.n2456 0.0265784
R17656 VDD.t528 VDD.n2457 0.0265784
R17657 VDD.n2459 VDD.n2401 0.0265784
R17658 VDD.n2476 VDD.n2474 0.0265784
R17659 VDD.n2484 VDD.n2474 0.0265784
R17660 VDD.n2490 VDD.n2475 0.0265784
R17661 VDD.n2480 VDD.n2475 0.0265784
R17662 VDD.n2482 VDD.n2481 0.0265784
R17663 VDD.n2481 VDD.n2480 0.0265784
R17664 VDD.n2486 VDD.n2485 0.0265784
R17665 VDD.n2485 VDD.n2484 0.0265784
R17666 VDD.n2697 VDD.n2696 0.0265784
R17667 VDD.n2696 VDD.n2695 0.0265784
R17668 VDD.n2699 VDD.n2690 0.0265784
R17669 VDD.n2700 VDD.n2699 0.0265784
R17670 VDD.n2702 VDD.n2701 0.0265784
R17671 VDD.n2701 VDD.n2700 0.0265784
R17672 VDD.n2695 VDD.n2692 0.0265784
R17673 VDD.n2692 VDD.n2691 0.0265784
R17674 VDD.n2715 VDD.n2714 0.0265784
R17675 VDD.t1381 VDD.n2715 0.0265784
R17676 VDD.n2717 VDD.n2659 0.0265784
R17677 VDD.n2734 VDD.n2732 0.0265784
R17678 VDD.n2742 VDD.n2732 0.0265784
R17679 VDD.n2748 VDD.n2733 0.0265784
R17680 VDD.n2738 VDD.n2733 0.0265784
R17681 VDD.n2740 VDD.n2739 0.0265784
R17682 VDD.n2739 VDD.n2738 0.0265784
R17683 VDD.n2744 VDD.n2743 0.0265784
R17684 VDD.n2743 VDD.n2742 0.0265784
R17685 VDD.n2955 VDD.n2954 0.0265784
R17686 VDD.n2954 VDD.n2953 0.0265784
R17687 VDD.n2957 VDD.n2948 0.0265784
R17688 VDD.n2958 VDD.n2957 0.0265784
R17689 VDD.n2960 VDD.n2959 0.0265784
R17690 VDD.n2959 VDD.n2958 0.0265784
R17691 VDD.n2953 VDD.n2950 0.0265784
R17692 VDD.n2950 VDD.n2949 0.0265784
R17693 VDD.n2973 VDD.n2972 0.0265784
R17694 VDD.t414 VDD.n2973 0.0265784
R17695 VDD.n2975 VDD.n2917 0.0265784
R17696 VDD.n2992 VDD.n2990 0.0265784
R17697 VDD.n3000 VDD.n2990 0.0265784
R17698 VDD.n3006 VDD.n2991 0.0265784
R17699 VDD.n2996 VDD.n2991 0.0265784
R17700 VDD.n2998 VDD.n2997 0.0265784
R17701 VDD.n2997 VDD.n2996 0.0265784
R17702 VDD.n3002 VDD.n3001 0.0265784
R17703 VDD.n3001 VDD.n3000 0.0265784
R17704 VDD.n3213 VDD.n3212 0.0265784
R17705 VDD.n3212 VDD.n3211 0.0265784
R17706 VDD.n3215 VDD.n3206 0.0265784
R17707 VDD.n3216 VDD.n3215 0.0265784
R17708 VDD.n3218 VDD.n3217 0.0265784
R17709 VDD.n3217 VDD.n3216 0.0265784
R17710 VDD.n3211 VDD.n3208 0.0265784
R17711 VDD.n3208 VDD.n3207 0.0265784
R17712 VDD.n3231 VDD.n3230 0.0265784
R17713 VDD.t591 VDD.n3231 0.0265784
R17714 VDD.n3233 VDD.n3175 0.0265784
R17715 VDD.n3250 VDD.n3248 0.0265784
R17716 VDD.n3258 VDD.n3248 0.0265784
R17717 VDD.n3264 VDD.n3249 0.0265784
R17718 VDD.n3254 VDD.n3249 0.0265784
R17719 VDD.n3256 VDD.n3255 0.0265784
R17720 VDD.n3255 VDD.n3254 0.0265784
R17721 VDD.n3260 VDD.n3259 0.0265784
R17722 VDD.n3259 VDD.n3258 0.0265784
R17723 VDD.n3471 VDD.n3470 0.0265784
R17724 VDD.n3470 VDD.n3469 0.0265784
R17725 VDD.n3473 VDD.n3464 0.0265784
R17726 VDD.n3474 VDD.n3473 0.0265784
R17727 VDD.n3476 VDD.n3475 0.0265784
R17728 VDD.n3475 VDD.n3474 0.0265784
R17729 VDD.n3469 VDD.n3466 0.0265784
R17730 VDD.n3466 VDD.n3465 0.0265784
R17731 VDD.n3489 VDD.n3488 0.0265784
R17732 VDD.t1086 VDD.n3489 0.0265784
R17733 VDD.n3491 VDD.n3433 0.0265784
R17734 VDD.n3508 VDD.n3506 0.0265784
R17735 VDD.n3516 VDD.n3506 0.0265784
R17736 VDD.n3522 VDD.n3507 0.0265784
R17737 VDD.n3512 VDD.n3507 0.0265784
R17738 VDD.n3514 VDD.n3513 0.0265784
R17739 VDD.n3513 VDD.n3512 0.0265784
R17740 VDD.n3518 VDD.n3517 0.0265784
R17741 VDD.n3517 VDD.n3516 0.0265784
R17742 VDD.n5791 VDD.n5790 0.0265784
R17743 VDD.n5790 VDD.n5789 0.0265784
R17744 VDD.n5793 VDD.n5784 0.0265784
R17745 VDD.n5794 VDD.n5793 0.0265784
R17746 VDD.n5796 VDD.n5795 0.0265784
R17747 VDD.n5795 VDD.n5794 0.0265784
R17748 VDD.n5789 VDD.n5786 0.0265784
R17749 VDD.n5786 VDD.n5785 0.0265784
R17750 VDD.n5809 VDD.n5808 0.0265784
R17751 VDD.t276 VDD.n5809 0.0265784
R17752 VDD.n5811 VDD.n5753 0.0265784
R17753 VDD.n5828 VDD.n5826 0.0265784
R17754 VDD.n5836 VDD.n5826 0.0265784
R17755 VDD.n5842 VDD.n5827 0.0265784
R17756 VDD.n5832 VDD.n5827 0.0265784
R17757 VDD.n5834 VDD.n5833 0.0265784
R17758 VDD.n5833 VDD.n5832 0.0265784
R17759 VDD.n5838 VDD.n5837 0.0265784
R17760 VDD.n5837 VDD.n5836 0.0265784
R17761 VDD.n5537 VDD.n5536 0.0265784
R17762 VDD.n5536 VDD.n5535 0.0265784
R17763 VDD.n5539 VDD.n5530 0.0265784
R17764 VDD.n5540 VDD.n5539 0.0265784
R17765 VDD.n5542 VDD.n5541 0.0265784
R17766 VDD.n5541 VDD.n5540 0.0265784
R17767 VDD.n5535 VDD.n5532 0.0265784
R17768 VDD.n5532 VDD.n5531 0.0265784
R17769 VDD.n5555 VDD.n5554 0.0265784
R17770 VDD.t512 VDD.n5555 0.0265784
R17771 VDD.n5557 VDD.n5499 0.0265784
R17772 VDD.n5574 VDD.n5572 0.0265784
R17773 VDD.n5582 VDD.n5572 0.0265784
R17774 VDD.n5588 VDD.n5573 0.0265784
R17775 VDD.n5578 VDD.n5573 0.0265784
R17776 VDD.n5580 VDD.n5579 0.0265784
R17777 VDD.n5579 VDD.n5578 0.0265784
R17778 VDD.n5584 VDD.n5583 0.0265784
R17779 VDD.n5583 VDD.n5582 0.0265784
R17780 VDD.n3729 VDD.n3728 0.0265784
R17781 VDD.n3728 VDD.n3727 0.0265784
R17782 VDD.n3731 VDD.n3722 0.0265784
R17783 VDD.n3732 VDD.n3731 0.0265784
R17784 VDD.n3734 VDD.n3733 0.0265784
R17785 VDD.n3733 VDD.n3732 0.0265784
R17786 VDD.n3727 VDD.n3724 0.0265784
R17787 VDD.n3724 VDD.n3723 0.0265784
R17788 VDD.n3747 VDD.n3746 0.0265784
R17789 VDD.t1085 VDD.n3747 0.0265784
R17790 VDD.n3749 VDD.n3691 0.0265784
R17791 VDD.n3766 VDD.n3764 0.0265784
R17792 VDD.n3774 VDD.n3764 0.0265784
R17793 VDD.n3780 VDD.n3765 0.0265784
R17794 VDD.n3770 VDD.n3765 0.0265784
R17795 VDD.n3772 VDD.n3771 0.0265784
R17796 VDD.n3771 VDD.n3770 0.0265784
R17797 VDD.n3776 VDD.n3775 0.0265784
R17798 VDD.n3775 VDD.n3774 0.0265784
R17799 VDD.n3987 VDD.n3986 0.0265784
R17800 VDD.n3986 VDD.n3985 0.0265784
R17801 VDD.n3989 VDD.n3980 0.0265784
R17802 VDD.n3990 VDD.n3989 0.0265784
R17803 VDD.n3992 VDD.n3991 0.0265784
R17804 VDD.n3991 VDD.n3990 0.0265784
R17805 VDD.n3985 VDD.n3982 0.0265784
R17806 VDD.n3982 VDD.n3981 0.0265784
R17807 VDD.n4005 VDD.n4004 0.0265784
R17808 VDD.t526 VDD.n4005 0.0265784
R17809 VDD.n4007 VDD.n3949 0.0265784
R17810 VDD.n4024 VDD.n4022 0.0265784
R17811 VDD.n4032 VDD.n4022 0.0265784
R17812 VDD.n4038 VDD.n4023 0.0265784
R17813 VDD.n4028 VDD.n4023 0.0265784
R17814 VDD.n4030 VDD.n4029 0.0265784
R17815 VDD.n4029 VDD.n4028 0.0265784
R17816 VDD.n4034 VDD.n4033 0.0265784
R17817 VDD.n4033 VDD.n4032 0.0265784
R17818 VDD.n4245 VDD.n4244 0.0265784
R17819 VDD.n4244 VDD.n4243 0.0265784
R17820 VDD.n4247 VDD.n4238 0.0265784
R17821 VDD.n4248 VDD.n4247 0.0265784
R17822 VDD.n4250 VDD.n4249 0.0265784
R17823 VDD.n4249 VDD.n4248 0.0265784
R17824 VDD.n4243 VDD.n4240 0.0265784
R17825 VDD.n4240 VDD.n4239 0.0265784
R17826 VDD.n4263 VDD.n4262 0.0265784
R17827 VDD.t525 VDD.n4263 0.0265784
R17828 VDD.n4265 VDD.n4207 0.0265784
R17829 VDD.n4282 VDD.n4280 0.0265784
R17830 VDD.n4290 VDD.n4280 0.0265784
R17831 VDD.n4296 VDD.n4281 0.0265784
R17832 VDD.n4286 VDD.n4281 0.0265784
R17833 VDD.n4288 VDD.n4287 0.0265784
R17834 VDD.n4287 VDD.n4286 0.0265784
R17835 VDD.n4292 VDD.n4291 0.0265784
R17836 VDD.n4291 VDD.n4290 0.0265784
R17837 VDD.n4503 VDD.n4502 0.0265784
R17838 VDD.n4502 VDD.n4501 0.0265784
R17839 VDD.n4505 VDD.n4496 0.0265784
R17840 VDD.n4506 VDD.n4505 0.0265784
R17841 VDD.n4508 VDD.n4507 0.0265784
R17842 VDD.n4507 VDD.n4506 0.0265784
R17843 VDD.n4501 VDD.n4498 0.0265784
R17844 VDD.n4498 VDD.n4497 0.0265784
R17845 VDD.n4521 VDD.n4520 0.0265784
R17846 VDD.t264 VDD.n4521 0.0265784
R17847 VDD.n4523 VDD.n4465 0.0265784
R17848 VDD.n4540 VDD.n4538 0.0265784
R17849 VDD.n4548 VDD.n4538 0.0265784
R17850 VDD.n4554 VDD.n4539 0.0265784
R17851 VDD.n4544 VDD.n4539 0.0265784
R17852 VDD.n4546 VDD.n4545 0.0265784
R17853 VDD.n4545 VDD.n4544 0.0265784
R17854 VDD.n4550 VDD.n4549 0.0265784
R17855 VDD.n4549 VDD.n4548 0.0265784
R17856 VDD.n4761 VDD.n4760 0.0265784
R17857 VDD.n4760 VDD.n4759 0.0265784
R17858 VDD.n4763 VDD.n4754 0.0265784
R17859 VDD.n4764 VDD.n4763 0.0265784
R17860 VDD.n4766 VDD.n4765 0.0265784
R17861 VDD.n4765 VDD.n4764 0.0265784
R17862 VDD.n4759 VDD.n4756 0.0265784
R17863 VDD.n4756 VDD.n4755 0.0265784
R17864 VDD.n4779 VDD.n4778 0.0265784
R17865 VDD.t590 VDD.n4779 0.0265784
R17866 VDD.n4781 VDD.n4723 0.0265784
R17867 VDD.n4798 VDD.n4796 0.0265784
R17868 VDD.n4806 VDD.n4796 0.0265784
R17869 VDD.n4812 VDD.n4797 0.0265784
R17870 VDD.n4802 VDD.n4797 0.0265784
R17871 VDD.n4804 VDD.n4803 0.0265784
R17872 VDD.n4803 VDD.n4802 0.0265784
R17873 VDD.n4808 VDD.n4807 0.0265784
R17874 VDD.n4807 VDD.n4806 0.0265784
R17875 VDD.n5019 VDD.n5018 0.0265784
R17876 VDD.n5018 VDD.n5017 0.0265784
R17877 VDD.n5021 VDD.n5012 0.0265784
R17878 VDD.n5022 VDD.n5021 0.0265784
R17879 VDD.n5024 VDD.n5023 0.0265784
R17880 VDD.n5023 VDD.n5022 0.0265784
R17881 VDD.n5017 VDD.n5014 0.0265784
R17882 VDD.n5014 VDD.n5013 0.0265784
R17883 VDD.n5037 VDD.n5036 0.0265784
R17884 VDD.t1024 VDD.n5037 0.0265784
R17885 VDD.n5039 VDD.n4981 0.0265784
R17886 VDD.n5056 VDD.n5054 0.0265784
R17887 VDD.n5064 VDD.n5054 0.0265784
R17888 VDD.n5070 VDD.n5055 0.0265784
R17889 VDD.n5060 VDD.n5055 0.0265784
R17890 VDD.n5062 VDD.n5061 0.0265784
R17891 VDD.n5061 VDD.n5060 0.0265784
R17892 VDD.n5066 VDD.n5065 0.0265784
R17893 VDD.n5065 VDD.n5064 0.0265784
R17894 VDD.n5277 VDD.n5276 0.0265784
R17895 VDD.n5276 VDD.n5275 0.0265784
R17896 VDD.n5279 VDD.n5270 0.0265784
R17897 VDD.n5280 VDD.n5279 0.0265784
R17898 VDD.n5282 VDD.n5281 0.0265784
R17899 VDD.n5281 VDD.n5280 0.0265784
R17900 VDD.n5275 VDD.n5272 0.0265784
R17901 VDD.n5272 VDD.n5271 0.0265784
R17902 VDD.n5295 VDD.n5294 0.0265784
R17903 VDD.t275 VDD.n5295 0.0265784
R17904 VDD.n5297 VDD.n5239 0.0265784
R17905 VDD.n5314 VDD.n5312 0.0265784
R17906 VDD.n5322 VDD.n5312 0.0265784
R17907 VDD.n5328 VDD.n5313 0.0265784
R17908 VDD.n5318 VDD.n5313 0.0265784
R17909 VDD.n5320 VDD.n5319 0.0265784
R17910 VDD.n5319 VDD.n5318 0.0265784
R17911 VDD.n5324 VDD.n5323 0.0265784
R17912 VDD.n5323 VDD.n5322 0.0265784
R17913 VDD.n1840 VDD.n1825 0.0261194
R17914 VDD.n2161 VDD.n2146 0.0261194
R17915 VDD.n2419 VDD.n2404 0.0261194
R17916 VDD.n2677 VDD.n2662 0.0261194
R17917 VDD.n2935 VDD.n2920 0.0261194
R17918 VDD.n3193 VDD.n3178 0.0261194
R17919 VDD.n3451 VDD.n3436 0.0261194
R17920 VDD.n5771 VDD.n5756 0.0261194
R17921 VDD.n5517 VDD.n5502 0.0261194
R17922 VDD.n3709 VDD.n3694 0.0261194
R17923 VDD.n3967 VDD.n3952 0.0261194
R17924 VDD.n4225 VDD.n4210 0.0261194
R17925 VDD.n4483 VDD.n4468 0.0261194
R17926 VDD.n4741 VDD.n4726 0.0261194
R17927 VDD.n4999 VDD.n4984 0.0261194
R17928 VDD.n5257 VDD.n5242 0.0261194
R17929 VDD.n1304 VDD 0.0260435
R17930 VDD.n1945 VDD.n1922 0.0258165
R17931 VDD.n1696 VDD.n1683 0.0257918
R17932 VDD.n2045 VDD.n2032 0.0257918
R17933 VDD.n2275 VDD.n2262 0.0257918
R17934 VDD.n2533 VDD.n2520 0.0257918
R17935 VDD.n2791 VDD.n2778 0.0257918
R17936 VDD.n3049 VDD.n3036 0.0257918
R17937 VDD.n3307 VDD.n3294 0.0257918
R17938 VDD.n5630 VDD.n5617 0.0257918
R17939 VDD.n5376 VDD.n5363 0.0257918
R17940 VDD.n3565 VDD.n3552 0.0257918
R17941 VDD.n3823 VDD.n3810 0.0257918
R17942 VDD.n4081 VDD.n4068 0.0257918
R17943 VDD.n4339 VDD.n4326 0.0257918
R17944 VDD.n4597 VDD.n4584 0.0257918
R17945 VDD.n4855 VDD.n4842 0.0257918
R17946 VDD.n5113 VDD.n5100 0.0257918
R17947 VDD.n1880 VDD.n1879 0.02576
R17948 VDD.n2201 VDD.n2200 0.02576
R17949 VDD.n2459 VDD.n2458 0.02576
R17950 VDD.n2717 VDD.n2716 0.02576
R17951 VDD.n2975 VDD.n2974 0.02576
R17952 VDD.n3233 VDD.n3232 0.02576
R17953 VDD.n3491 VDD.n3490 0.02576
R17954 VDD.n5811 VDD.n5810 0.02576
R17955 VDD.n5557 VDD.n5556 0.02576
R17956 VDD.n3749 VDD.n3748 0.02576
R17957 VDD.n4007 VDD.n4006 0.02576
R17958 VDD.n4265 VDD.n4264 0.02576
R17959 VDD.n4523 VDD.n4522 0.02576
R17960 VDD.n4781 VDD.n4780 0.02576
R17961 VDD.n5039 VDD.n5038 0.02576
R17962 VDD.n5297 VDD.n5296 0.02576
R17963 VDD.n1315 VDD.n1314 0.0254026
R17964 VDD.n1310 VDD.n1308 0.0249681
R17965 VDD.n1311 VDD.n1310 0.0249681
R17966 VDD.n1453 VDD.n1449 0.0249681
R17967 VDD.n1449 VDD.n1447 0.0249681
R17968 VDD.n1447 VDD.n1443 0.0249681
R17969 VDD.n1443 VDD.n1441 0.0249681
R17970 VDD.n1441 VDD.n1437 0.0249681
R17971 VDD.n1437 VDD.n1433 0.0249681
R17972 VDD.n1331 VDD.n1327 0.0249681
R17973 VDD.n1333 VDD.n1331 0.0249681
R17974 VDD.n1337 VDD.n1333 0.0249681
R17975 VDD.n1339 VDD.n1337 0.0249681
R17976 VDD.n1340 VDD.n1339 0.0249681
R17977 VDD.n1422 VDD.n1418 0.0249681
R17978 VDD.n1418 VDD.n1416 0.0249681
R17979 VDD.n1416 VDD.n1412 0.0249681
R17980 VDD.n1412 VDD.n1410 0.0249681
R17981 VDD.n1393 VDD.n1389 0.0249681
R17982 VDD.n1389 VDD.n1387 0.0249681
R17983 VDD.n1387 VDD.n1383 0.0249681
R17984 VDD.n1383 VDD.n1381 0.0249681
R17985 VDD.n1351 VDD.n1349 0.0249681
R17986 VDD.n1354 VDD.n1351 0.0249681
R17987 VDD.n1356 VDD.n1354 0.0249681
R17988 VDD.n1358 VDD.n1356 0.0249681
R17989 VDD.n1365 VDD.n1363 0.0249681
R17990 VDD.n1525 VDD.n1523 0.0249681
R17991 VDD.n1523 VDD.n1519 0.0249681
R17992 VDD.n1519 VDD.n1517 0.0249681
R17993 VDD.n1517 VDD.n1513 0.0249681
R17994 VDD.n1503 VDD.n1501 0.0249681
R17995 VDD.n1501 VDD.n1497 0.0249681
R17996 VDD.n1497 VDD.n1495 0.0249681
R17997 VDD.n1495 VDD.n1491 0.0249681
R17998 VDD.n1491 VDD.n1489 0.0249681
R17999 VDD.n1489 VDD.n1485 0.0249681
R18000 VDD.n1485 VDD.n1481 0.0249681
R18001 VDD.n1481 VDD.n1479 0.0249681
R18002 VDD.n1479 VDD.n1475 0.0249681
R18003 VDD.n1475 VDD.n1473 0.0249681
R18004 VDD.n1473 VDD.n1469 0.0249681
R18005 VDD.n1469 VDD.n1467 0.0249681
R18006 VDD.n1467 VDD.n1463 0.0249681
R18007 VDD.n1286 VDD.n1285 0.0249681
R18008 VDD.n1285 VDD.n1283 0.0249681
R18009 VDD.n1546 VDD.n1544 0.0243281
R18010 VDD.n1454 VDD.n1453 0.0241145
R18011 VDD.n1882 VDD.n1881 0.0228205
R18012 VDD.n2203 VDD.n2202 0.0228205
R18013 VDD.n2461 VDD.n2460 0.0228205
R18014 VDD.n2719 VDD.n2718 0.0228205
R18015 VDD.n2977 VDD.n2976 0.0228205
R18016 VDD.n3235 VDD.n3234 0.0228205
R18017 VDD.n3493 VDD.n3492 0.0228205
R18018 VDD.n5813 VDD.n5812 0.0228205
R18019 VDD.n5559 VDD.n5558 0.0228205
R18020 VDD.n3751 VDD.n3750 0.0228205
R18021 VDD.n4009 VDD.n4008 0.0228205
R18022 VDD.n4267 VDD.n4266 0.0228205
R18023 VDD.n4525 VDD.n4524 0.0228205
R18024 VDD.n4783 VDD.n4782 0.0228205
R18025 VDD.n5041 VDD.n5040 0.0228205
R18026 VDD.n5299 VDD.n5298 0.0228205
R18027 VDD.n1881 VDD.n1820 0.0223212
R18028 VDD.n2202 VDD.n2141 0.0223212
R18029 VDD.n2460 VDD.n2399 0.0223212
R18030 VDD.n2718 VDD.n2657 0.0223212
R18031 VDD.n2976 VDD.n2915 0.0223212
R18032 VDD.n3234 VDD.n3173 0.0223212
R18033 VDD.n3492 VDD.n3431 0.0223212
R18034 VDD.n5812 VDD.n5751 0.0223212
R18035 VDD.n5558 VDD.n5497 0.0223212
R18036 VDD.n3750 VDD.n3689 0.0223212
R18037 VDD.n4008 VDD.n3947 0.0223212
R18038 VDD.n4266 VDD.n4205 0.0223212
R18039 VDD.n4524 VDD.n4463 0.0223212
R18040 VDD.n4782 VDD.n4721 0.0223212
R18041 VDD.n5040 VDD.n4979 0.0223212
R18042 VDD.n5298 VDD.n5237 0.0223212
R18043 VDD.n1374 VDD.n1346 0.0218724
R18044 VDD.n851 VDD 0.02175
R18045 VDD.n845 VDD 0.02175
R18046 VDD.n839 VDD 0.02175
R18047 VDD.n833 VDD 0.02175
R18048 VDD.n827 VDD 0.02175
R18049 VDD.n1234 VDD 0.02175
R18050 VDD.n1228 VDD 0.02175
R18051 VDD.n1222 VDD 0.02175
R18052 VDD.n1216 VDD 0.02175
R18053 VDD.n1210 VDD 0.02175
R18054 VDD.n1600 VDD 0.0213145
R18055 VDD.n1410 VDD.n1406 0.0212447
R18056 VDD.n1504 VDD.n1503 0.0207128
R18057 VDD.n1622 VDD.n1621 0.0205312
R18058 VDD.n1433 VDD.n1431 0.0198592
R18059 VDD.n1461 VDD.n1460 0.0188511
R18060 VDD.n1946 VDD.n1945 0.0183679
R18061 VDD.n1799 VDD.n1798 0.0182941
R18062 VDD.n2007 VDD.n2006 0.0182941
R18063 VDD.n2378 VDD.n2377 0.0182941
R18064 VDD.n2636 VDD.n2635 0.0182941
R18065 VDD.n2894 VDD.n2893 0.0182941
R18066 VDD.n3152 VDD.n3151 0.0182941
R18067 VDD.n3410 VDD.n3409 0.0182941
R18068 VDD.n5733 VDD.n5732 0.0182941
R18069 VDD.n5479 VDD.n5478 0.0182941
R18070 VDD.n3668 VDD.n3667 0.0182941
R18071 VDD.n3926 VDD.n3925 0.0182941
R18072 VDD.n4184 VDD.n4183 0.0182941
R18073 VDD.n4442 VDD.n4441 0.0182941
R18074 VDD.n4700 VDD.n4699 0.0182941
R18075 VDD.n4958 VDD.n4957 0.0182941
R18076 VDD.n5216 VDD.n5215 0.0182941
R18077 VDD.n1779 VDD.n1777 0.0178611
R18078 VDD.n1987 VDD.n1985 0.0178611
R18079 VDD.n2358 VDD.n2356 0.0178611
R18080 VDD.n2616 VDD.n2614 0.0178611
R18081 VDD.n2874 VDD.n2872 0.0178611
R18082 VDD.n3132 VDD.n3130 0.0178611
R18083 VDD.n3390 VDD.n3388 0.0178611
R18084 VDD.n5713 VDD.n5711 0.0178611
R18085 VDD.n5459 VDD.n5457 0.0178611
R18086 VDD.n3648 VDD.n3646 0.0178611
R18087 VDD.n3906 VDD.n3904 0.0178611
R18088 VDD.n4164 VDD.n4162 0.0178611
R18089 VDD.n4422 VDD.n4420 0.0178611
R18090 VDD.n4680 VDD.n4678 0.0178611
R18091 VDD.n4938 VDD.n4936 0.0178611
R18092 VDD.n5196 VDD.n5194 0.0178611
R18093 VDD.n1808 VDD.n1807 0.0177731
R18094 VDD.n2387 VDD.n2386 0.0177731
R18095 VDD.n2645 VDD.n2644 0.0177731
R18096 VDD.n2903 VDD.n2902 0.0177731
R18097 VDD.n3161 VDD.n3160 0.0177731
R18098 VDD.n3419 VDD.n3418 0.0177731
R18099 VDD.n3677 VDD.n3676 0.0177731
R18100 VDD.n3935 VDD.n3934 0.0177731
R18101 VDD.n4193 VDD.n4192 0.0177731
R18102 VDD.n4451 VDD.n4450 0.0177731
R18103 VDD.n4709 VDD.n4708 0.0177731
R18104 VDD.n4967 VDD.n4966 0.0177731
R18105 VDD.n5225 VDD.n5224 0.0177731
R18106 VDD.n1368 VDD.n1366 0.0172553
R18107 VDD.n810 VDD 0.0171185
R18108 VDD VDD.n799 0.0171185
R18109 VDD.n1193 VDD 0.0171185
R18110 VDD VDD.n1182 0.0171185
R18111 VDD.n1758 VDD.n1757 0.0168386
R18112 VDD.n2107 VDD.n2106 0.0168386
R18113 VDD.n2337 VDD.n2336 0.0168386
R18114 VDD.n2595 VDD.n2594 0.0168386
R18115 VDD.n2853 VDD.n2852 0.0168386
R18116 VDD.n3111 VDD.n3110 0.0168386
R18117 VDD.n3369 VDD.n3368 0.0168386
R18118 VDD.n5692 VDD.n5691 0.0168386
R18119 VDD.n5438 VDD.n5437 0.0168386
R18120 VDD.n3627 VDD.n3626 0.0168386
R18121 VDD.n3885 VDD.n3884 0.0168386
R18122 VDD.n4143 VDD.n4142 0.0168386
R18123 VDD.n4401 VDD.n4400 0.0168386
R18124 VDD.n4659 VDD.n4658 0.0168386
R18125 VDD.n4917 VDD.n4916 0.0168386
R18126 VDD.n5175 VDD.n5174 0.0168386
R18127 VDD.n1710 VDD.n1679 0.0168372
R18128 VDD.n2059 VDD.n2028 0.0168372
R18129 VDD.n2289 VDD.n2258 0.0168372
R18130 VDD.n2547 VDD.n2516 0.0168372
R18131 VDD.n2805 VDD.n2774 0.0168372
R18132 VDD.n3063 VDD.n3032 0.0168372
R18133 VDD.n3321 VDD.n3290 0.0168372
R18134 VDD.n5644 VDD.n5613 0.0168372
R18135 VDD.n5390 VDD.n5359 0.0168372
R18136 VDD.n3579 VDD.n3548 0.0168372
R18137 VDD.n3837 VDD.n3806 0.0168372
R18138 VDD.n4095 VDD.n4064 0.0168372
R18139 VDD.n4353 VDD.n4322 0.0168372
R18140 VDD.n4611 VDD.n4580 0.0168372
R18141 VDD.n4869 VDD.n4838 0.0168372
R18142 VDD.n5127 VDD.n5096 0.0168372
R18143 VDD.n861 VDD.n860 0.0165987
R18144 VDD.n1244 VDD.n1243 0.0165987
R18145 VDD.n1679 VDD.n1669 0.0163404
R18146 VDD.n1758 VDD.n1717 0.0163404
R18147 VDD.n2028 VDD.n2018 0.0163404
R18148 VDD.n2107 VDD.n2066 0.0163404
R18149 VDD.n2258 VDD.n2248 0.0163404
R18150 VDD.n2337 VDD.n2296 0.0163404
R18151 VDD.n2516 VDD.n2506 0.0163404
R18152 VDD.n2595 VDD.n2554 0.0163404
R18153 VDD.n2774 VDD.n2764 0.0163404
R18154 VDD.n2853 VDD.n2812 0.0163404
R18155 VDD.n3032 VDD.n3022 0.0163404
R18156 VDD.n3111 VDD.n3070 0.0163404
R18157 VDD.n3290 VDD.n3280 0.0163404
R18158 VDD.n3369 VDD.n3328 0.0163404
R18159 VDD.n5613 VDD.n5603 0.0163404
R18160 VDD.n5692 VDD.n5651 0.0163404
R18161 VDD.n5359 VDD.n5349 0.0163404
R18162 VDD.n5438 VDD.n5397 0.0163404
R18163 VDD.n3548 VDD.n3538 0.0163404
R18164 VDD.n3627 VDD.n3586 0.0163404
R18165 VDD.n3806 VDD.n3796 0.0163404
R18166 VDD.n3885 VDD.n3844 0.0163404
R18167 VDD.n4064 VDD.n4054 0.0163404
R18168 VDD.n4143 VDD.n4102 0.0163404
R18169 VDD.n4322 VDD.n4312 0.0163404
R18170 VDD.n4401 VDD.n4360 0.0163404
R18171 VDD.n4580 VDD.n4570 0.0163404
R18172 VDD.n4659 VDD.n4618 0.0163404
R18173 VDD.n4838 VDD.n4828 0.0163404
R18174 VDD.n4917 VDD.n4876 0.0163404
R18175 VDD.n5096 VDD.n5086 0.0163404
R18176 VDD.n5175 VDD.n5134 0.0163404
R18177 VDD.n1423 VDD.n1422 0.0161915
R18178 VDD.n855 VDD.n854 0.016125
R18179 VDD.n1238 VDD.n1237 0.016125
R18180 VDD.n1961 VDD.n1941 0.0154506
R18181 VDD.n1969 VDD.n1968 0.015449
R18182 VDD.n1405 VDD.n1401 0.0153936
R18183 VDD.n1513 VDD.n1511 0.0151277
R18184 VDD.n1971 VDD.n1970 0.0150463
R18185 VDD.n1970 VDD.t1038 0.0150463
R18186 VDD.n1963 VDD.n1929 0.0150463
R18187 VDD.t1026 VDD.n1963 0.0150463
R18188 VDD.n1961 VDD.n1960 0.0150463
R18189 VDD.n1964 VDD.t1026 0.0150463
R18190 VDD.n1968 VDD.n1967 0.0150463
R18191 VDD.n1965 VDD.n1964 0.0150463
R18192 VDD.t1036 VDD.n1951 0.0150463
R18193 VDD.n1951 VDD.n1950 0.0150463
R18194 VDD.n794 VDD.n513 0.015
R18195 VDD.n1839 VDD.n1827 0.0149834
R18196 VDD.n2160 VDD.n2148 0.0149834
R18197 VDD.n2418 VDD.n2406 0.0149834
R18198 VDD.n2676 VDD.n2664 0.0149834
R18199 VDD.n2934 VDD.n2922 0.0149834
R18200 VDD.n3192 VDD.n3180 0.0149834
R18201 VDD.n3450 VDD.n3438 0.0149834
R18202 VDD.n5770 VDD.n5758 0.0149834
R18203 VDD.n5516 VDD.n5504 0.0149834
R18204 VDD.n3708 VDD.n3696 0.0149834
R18205 VDD.n3966 VDD.n3954 0.0149834
R18206 VDD.n4224 VDD.n4212 0.0149834
R18207 VDD.n4482 VDD.n4470 0.0149834
R18208 VDD.n4740 VDD.n4728 0.0149834
R18209 VDD.n4998 VDD.n4986 0.0149834
R18210 VDD.n5256 VDD.n5244 0.0149834
R18211 VDD.n1325 VDD.n1324 0.0148617
R18212 VDD.n676 VDD.n674 0.0146339
R18213 VDD.n1026 VDD.n1024 0.0146339
R18214 VDD.n271 VDD.n269 0.0146339
R18215 VDD.n1394 VDD.n1393 0.0145957
R18216 VDD.n1377 VDD.n1376 0.0145957
R18217 VDD.n1886 VDD.n1817 0.0145797
R18218 VDD.n2207 VDD.n2138 0.0145797
R18219 VDD.n2465 VDD.n2396 0.0145797
R18220 VDD.n2723 VDD.n2654 0.0145797
R18221 VDD.n2981 VDD.n2912 0.0145797
R18222 VDD.n3239 VDD.n3170 0.0145797
R18223 VDD.n3497 VDD.n3428 0.0145797
R18224 VDD.n5817 VDD.n5748 0.0145797
R18225 VDD.n5563 VDD.n5494 0.0145797
R18226 VDD.n3755 VDD.n3686 0.0145797
R18227 VDD.n4013 VDD.n3944 0.0145797
R18228 VDD.n4271 VDD.n4202 0.0145797
R18229 VDD.n4529 VDD.n4460 0.0145797
R18230 VDD.n4787 VDD.n4718 0.0145797
R18231 VDD.n5045 VDD.n4976 0.0145797
R18232 VDD.n5303 VDD.n5234 0.0145797
R18233 VDD.n1721 VDD.n1720 0.0143889
R18234 VDD.n2070 VDD.n2069 0.0143889
R18235 VDD.n2300 VDD.n2299 0.0143889
R18236 VDD.n2558 VDD.n2557 0.0143889
R18237 VDD.n2816 VDD.n2815 0.0143889
R18238 VDD.n3074 VDD.n3073 0.0143889
R18239 VDD.n3332 VDD.n3331 0.0143889
R18240 VDD.n5655 VDD.n5654 0.0143889
R18241 VDD.n5401 VDD.n5400 0.0143889
R18242 VDD.n3590 VDD.n3589 0.0143889
R18243 VDD.n3848 VDD.n3847 0.0143889
R18244 VDD.n4106 VDD.n4105 0.0143889
R18245 VDD.n4364 VDD.n4363 0.0143889
R18246 VDD.n4622 VDD.n4621 0.0143889
R18247 VDD.n4880 VDD.n4879 0.0143889
R18248 VDD.n5138 VDD.n5137 0.0143889
R18249 VDD.n485 VDD.n481 0.0143889
R18250 VDD.n83 VDD.n79 0.0143889
R18251 VDD.n1308 VDD.n1304 0.0143298
R18252 VDD.n1180 VDD.n1179 0.0142984
R18253 VDD.n1979 VDD.n1978 0.0138929
R18254 VDD.n1345 VDD.n1343 0.0137979
R18255 VDD VDD.n1840 0.0131689
R18256 VDD VDD.n2161 0.0131689
R18257 VDD VDD.n2419 0.0131689
R18258 VDD VDD.n2677 0.0131689
R18259 VDD VDD.n2935 0.0131689
R18260 VDD VDD.n3193 0.0131689
R18261 VDD VDD.n3451 0.0131689
R18262 VDD VDD.n5771 0.0131689
R18263 VDD VDD.n5517 0.0131689
R18264 VDD VDD.n3709 0.0131689
R18265 VDD VDD.n3967 0.0131689
R18266 VDD VDD.n4225 0.0131689
R18267 VDD VDD.n4483 0.0131689
R18268 VDD VDD.n4741 0.0131689
R18269 VDD VDD.n4999 0.0131689
R18270 VDD VDD.n5257 0.0131689
R18271 VDD.n447 VDD 0.013
R18272 VDD.n44 VDD 0.013
R18273 VDD.n1314 VDD 0.012734
R18274 VDD.n1349 VDD 0.012734
R18275 VDD.n1261 VDD 0.012734
R18276 VDD.n1544 VDD.n1543 0.0126094
R18277 VDD.n537 VDD.n533 0.0126053
R18278 VDD.n576 VDD.n572 0.0126053
R18279 VDD.n572 VDD.n570 0.0126053
R18280 VDD.n570 VDD.n566 0.0126053
R18281 VDD.n566 VDD.n564 0.0126053
R18282 VDD.n564 VDD.n560 0.0126053
R18283 VDD.n560 VDD.n558 0.0126053
R18284 VDD.n558 VDD.n554 0.0126053
R18285 VDD.n554 VDD.n552 0.0126053
R18286 VDD.n551 VDD.n550 0.0126053
R18287 VDD.n550 VDD.n548 0.0126053
R18288 VDD.n548 VDD.n544 0.0126053
R18289 VDD.n544 VDD.n528 0.0126053
R18290 VDD.n598 VDD.n594 0.0126053
R18291 VDD.n600 VDD.n598 0.0126053
R18292 VDD.n604 VDD.n600 0.0126053
R18293 VDD.n606 VDD.n604 0.0126053
R18294 VDD.n610 VDD.n606 0.0126053
R18295 VDD.n612 VDD.n610 0.0126053
R18296 VDD.n616 VDD.n612 0.0126053
R18297 VDD.n618 VDD.n616 0.0126053
R18298 VDD.n619 VDD.n618 0.0126053
R18299 VDD.n624 VDD.n622 0.0126053
R18300 VDD.n628 VDD.n624 0.0126053
R18301 VDD.n630 VDD.n628 0.0126053
R18302 VDD.n634 VDD.n630 0.0126053
R18303 VDD.n659 VDD.n655 0.0126053
R18304 VDD.n655 VDD.n653 0.0126053
R18305 VDD.n653 VDD.n649 0.0126053
R18306 VDD.n649 VDD.n647 0.0126053
R18307 VDD.n647 VDD.n643 0.0126053
R18308 VDD.n643 VDD.n641 0.0126053
R18309 VDD.n641 VDD.n515 0.0126053
R18310 VDD.n791 VDD.n790 0.0126053
R18311 VDD.n790 VDD.n788 0.0126053
R18312 VDD.n775 VDD.n773 0.0126053
R18313 VDD.n773 VDD.n769 0.0126053
R18314 VDD.n769 VDD.n765 0.0126053
R18315 VDD.n765 VDD.n763 0.0126053
R18316 VDD.n763 VDD.n759 0.0126053
R18317 VDD.n759 VDD.n757 0.0126053
R18318 VDD.n757 VDD.n753 0.0126053
R18319 VDD.n753 VDD.n751 0.0126053
R18320 VDD.n751 VDD.n747 0.0126053
R18321 VDD.n747 VDD.n745 0.0126053
R18322 VDD.n744 VDD.n743 0.0126053
R18323 VDD.n732 VDD.n728 0.0126053
R18324 VDD.n728 VDD.n726 0.0126053
R18325 VDD.n726 VDD.n722 0.0126053
R18326 VDD.n722 VDD.n718 0.0126053
R18327 VDD.n718 VDD.n716 0.0126053
R18328 VDD.n716 VDD.n712 0.0126053
R18329 VDD.n712 VDD.n710 0.0126053
R18330 VDD.n710 VDD.n706 0.0126053
R18331 VDD.n706 VDD.n704 0.0126053
R18332 VDD.n704 VDD.n700 0.0126053
R18333 VDD.n700 VDD.n698 0.0126053
R18334 VDD.n697 VDD.n696 0.0126053
R18335 VDD.n696 VDD.n694 0.0126053
R18336 VDD.n694 VDD.n691 0.0126053
R18337 VDD.n691 VDD.n689 0.0126053
R18338 VDD.n682 VDD.n680 0.0126053
R18339 VDD.n677 VDD.n676 0.0126053
R18340 VDD.n887 VDD.n883 0.0126053
R18341 VDD.n926 VDD.n922 0.0126053
R18342 VDD.n922 VDD.n920 0.0126053
R18343 VDD.n920 VDD.n916 0.0126053
R18344 VDD.n916 VDD.n914 0.0126053
R18345 VDD.n914 VDD.n910 0.0126053
R18346 VDD.n910 VDD.n908 0.0126053
R18347 VDD.n908 VDD.n904 0.0126053
R18348 VDD.n904 VDD.n902 0.0126053
R18349 VDD.n901 VDD.n900 0.0126053
R18350 VDD.n900 VDD.n898 0.0126053
R18351 VDD.n898 VDD.n894 0.0126053
R18352 VDD.n894 VDD.n878 0.0126053
R18353 VDD.n948 VDD.n944 0.0126053
R18354 VDD.n950 VDD.n948 0.0126053
R18355 VDD.n954 VDD.n950 0.0126053
R18356 VDD.n956 VDD.n954 0.0126053
R18357 VDD.n960 VDD.n956 0.0126053
R18358 VDD.n962 VDD.n960 0.0126053
R18359 VDD.n966 VDD.n962 0.0126053
R18360 VDD.n968 VDD.n966 0.0126053
R18361 VDD.n969 VDD.n968 0.0126053
R18362 VDD.n974 VDD.n972 0.0126053
R18363 VDD.n978 VDD.n974 0.0126053
R18364 VDD.n980 VDD.n978 0.0126053
R18365 VDD.n984 VDD.n980 0.0126053
R18366 VDD.n1009 VDD.n1005 0.0126053
R18367 VDD.n1005 VDD.n1003 0.0126053
R18368 VDD.n1003 VDD.n999 0.0126053
R18369 VDD.n999 VDD.n997 0.0126053
R18370 VDD.n997 VDD.n993 0.0126053
R18371 VDD.n993 VDD.n991 0.0126053
R18372 VDD.n991 VDD.n865 0.0126053
R18373 VDD.n1141 VDD.n1140 0.0126053
R18374 VDD.n1140 VDD.n1138 0.0126053
R18375 VDD.n1125 VDD.n1123 0.0126053
R18376 VDD.n1123 VDD.n1119 0.0126053
R18377 VDD.n1119 VDD.n1115 0.0126053
R18378 VDD.n1115 VDD.n1113 0.0126053
R18379 VDD.n1113 VDD.n1109 0.0126053
R18380 VDD.n1109 VDD.n1107 0.0126053
R18381 VDD.n1107 VDD.n1103 0.0126053
R18382 VDD.n1103 VDD.n1101 0.0126053
R18383 VDD.n1101 VDD.n1097 0.0126053
R18384 VDD.n1097 VDD.n1095 0.0126053
R18385 VDD.n1094 VDD.n1093 0.0126053
R18386 VDD.n1082 VDD.n1078 0.0126053
R18387 VDD.n1078 VDD.n1076 0.0126053
R18388 VDD.n1076 VDD.n1072 0.0126053
R18389 VDD.n1072 VDD.n1068 0.0126053
R18390 VDD.n1068 VDD.n1066 0.0126053
R18391 VDD.n1066 VDD.n1062 0.0126053
R18392 VDD.n1062 VDD.n1060 0.0126053
R18393 VDD.n1060 VDD.n1056 0.0126053
R18394 VDD.n1056 VDD.n1054 0.0126053
R18395 VDD.n1054 VDD.n1050 0.0126053
R18396 VDD.n1050 VDD.n1048 0.0126053
R18397 VDD.n1047 VDD.n1046 0.0126053
R18398 VDD.n1046 VDD.n1044 0.0126053
R18399 VDD.n1044 VDD.n1041 0.0126053
R18400 VDD.n1041 VDD.n1039 0.0126053
R18401 VDD.n1032 VDD.n1030 0.0126053
R18402 VDD.n1027 VDD.n1026 0.0126053
R18403 VDD.n136 VDD.n132 0.0126053
R18404 VDD.n175 VDD.n171 0.0126053
R18405 VDD.n171 VDD.n169 0.0126053
R18406 VDD.n169 VDD.n165 0.0126053
R18407 VDD.n165 VDD.n163 0.0126053
R18408 VDD.n163 VDD.n159 0.0126053
R18409 VDD.n159 VDD.n157 0.0126053
R18410 VDD.n157 VDD.n153 0.0126053
R18411 VDD.n153 VDD.n151 0.0126053
R18412 VDD.n150 VDD.n149 0.0126053
R18413 VDD.n149 VDD.n147 0.0126053
R18414 VDD.n147 VDD.n143 0.0126053
R18415 VDD.n143 VDD.n127 0.0126053
R18416 VDD.n197 VDD.n193 0.0126053
R18417 VDD.n199 VDD.n197 0.0126053
R18418 VDD.n203 VDD.n199 0.0126053
R18419 VDD.n205 VDD.n203 0.0126053
R18420 VDD.n209 VDD.n205 0.0126053
R18421 VDD.n211 VDD.n209 0.0126053
R18422 VDD.n215 VDD.n211 0.0126053
R18423 VDD.n217 VDD.n215 0.0126053
R18424 VDD.n218 VDD.n217 0.0126053
R18425 VDD.n223 VDD.n221 0.0126053
R18426 VDD.n227 VDD.n223 0.0126053
R18427 VDD.n229 VDD.n227 0.0126053
R18428 VDD.n233 VDD.n229 0.0126053
R18429 VDD.n254 VDD.n250 0.0126053
R18430 VDD.n250 VDD.n248 0.0126053
R18431 VDD.n248 VDD.n244 0.0126053
R18432 VDD.n244 VDD.n242 0.0126053
R18433 VDD.n242 VDD.n238 0.0126053
R18434 VDD.n238 VDD.n114 0.0126053
R18435 VDD.n389 VDD.n387 0.0126053
R18436 VDD.n386 VDD.n385 0.0126053
R18437 VDD.n385 VDD.n383 0.0126053
R18438 VDD.n370 VDD.n368 0.0126053
R18439 VDD.n368 VDD.n364 0.0126053
R18440 VDD.n364 VDD.n360 0.0126053
R18441 VDD.n360 VDD.n358 0.0126053
R18442 VDD.n358 VDD.n354 0.0126053
R18443 VDD.n354 VDD.n352 0.0126053
R18444 VDD.n352 VDD.n348 0.0126053
R18445 VDD.n348 VDD.n346 0.0126053
R18446 VDD.n346 VDD.n342 0.0126053
R18447 VDD.n342 VDD.n340 0.0126053
R18448 VDD.n339 VDD.n338 0.0126053
R18449 VDD.n327 VDD.n323 0.0126053
R18450 VDD.n323 VDD.n321 0.0126053
R18451 VDD.n321 VDD.n317 0.0126053
R18452 VDD.n317 VDD.n313 0.0126053
R18453 VDD.n313 VDD.n311 0.0126053
R18454 VDD.n311 VDD.n307 0.0126053
R18455 VDD.n307 VDD.n305 0.0126053
R18456 VDD.n305 VDD.n301 0.0126053
R18457 VDD.n301 VDD.n299 0.0126053
R18458 VDD.n299 VDD.n295 0.0126053
R18459 VDD.n295 VDD.n293 0.0126053
R18460 VDD.n292 VDD.n291 0.0126053
R18461 VDD.n291 VDD.n289 0.0126053
R18462 VDD.n289 VDD.n286 0.0126053
R18463 VDD.n286 VDD.n284 0.0126053
R18464 VDD.n277 VDD.n275 0.0126053
R18465 VDD.n272 VDD.n271 0.0126053
R18466 VDD.n474 VDD 0.0125739
R18467 VDD.n72 VDD 0.0125739
R18468 VDD.n1611 VDD.n1609 0.0125192
R18469 VDD.n793 VDD.n792 0.0124737
R18470 VDD.n1143 VDD.n1142 0.0124737
R18471 VDD.n1785 VDD 0.0123056
R18472 VDD.n1993 VDD 0.0123056
R18473 VDD.n2364 VDD 0.0123056
R18474 VDD.n2622 VDD 0.0123056
R18475 VDD.n2880 VDD 0.0123056
R18476 VDD.n3138 VDD 0.0123056
R18477 VDD.n3396 VDD 0.0123056
R18478 VDD.n5719 VDD 0.0123056
R18479 VDD.n5465 VDD 0.0123056
R18480 VDD.n3654 VDD 0.0123056
R18481 VDD.n3912 VDD 0.0123056
R18482 VDD.n4170 VDD 0.0123056
R18483 VDD.n4428 VDD 0.0123056
R18484 VDD.n4686 VDD 0.0123056
R18485 VDD.n4944 VDD 0.0123056
R18486 VDD.n5202 VDD 0.0123056
R18487 VDD VDD.n467 0.0123056
R18488 VDD.n413 VDD 0.0123056
R18489 VDD VDD.n65 0.0123056
R18490 VDD.n1571 VDD 0.0123056
R18491 VDD.n390 VDD.n114 0.0122105
R18492 VDD.n587 VDD.n528 0.0119152
R18493 VDD.n937 VDD.n878 0.0119152
R18494 VDD.n1842 VDD 0.0118881
R18495 VDD.n2163 VDD 0.0118881
R18496 VDD.n2421 VDD 0.0118881
R18497 VDD.n2679 VDD 0.0118881
R18498 VDD.n2937 VDD 0.0118881
R18499 VDD.n3195 VDD 0.0118881
R18500 VDD.n3453 VDD 0.0118881
R18501 VDD.n5773 VDD 0.0118881
R18502 VDD.n5519 VDD 0.0118881
R18503 VDD.n3711 VDD 0.0118881
R18504 VDD.n3969 VDD 0.0118881
R18505 VDD.n4227 VDD 0.0118881
R18506 VDD.n4485 VDD 0.0118881
R18507 VDD.n4743 VDD 0.0118881
R18508 VDD.n5001 VDD 0.0118881
R18509 VDD.n5259 VDD 0.0118881
R18510 VDD.n1255 VDD.n1251 0.0117745
R18511 VDD.n1539 VDD.n1537 0.0117745
R18512 VDD.n1537 VDD.n1533 0.0117745
R18513 VDD.n1533 VDD.n1529 0.0117745
R18514 VDD.n1529 VDD.n1527 0.0117745
R18515 VDD.n1613 VDD.n1611 0.0117367
R18516 VDD.n501 VDD 0.0116111
R18517 VDD.n428 VDD 0.0116111
R18518 VDD.n394 VDD 0.0116111
R18519 VDD.n99 VDD 0.0116111
R18520 VDD.n1586 VDD 0.0116111
R18521 VDD.n1552 VDD 0.0116111
R18522 VDD.n11 VDD 0.0114012
R18523 VDD.n1155 VDD 0.0114012
R18524 VDD.n186 VDD.n127 0.0113889
R18525 VDD.n1875 VDD.n1874 0.0111456
R18526 VDD.n2196 VDD.n2195 0.0111456
R18527 VDD.n2454 VDD.n2453 0.0111456
R18528 VDD.n2712 VDD.n2711 0.0111456
R18529 VDD.n2970 VDD.n2969 0.0111456
R18530 VDD.n3228 VDD.n3227 0.0111456
R18531 VDD.n3486 VDD.n3485 0.0111456
R18532 VDD.n5806 VDD.n5805 0.0111456
R18533 VDD.n5552 VDD.n5551 0.0111456
R18534 VDD.n3744 VDD.n3743 0.0111456
R18535 VDD.n4002 VDD.n4001 0.0111456
R18536 VDD.n4260 VDD.n4259 0.0111456
R18537 VDD.n4518 VDD.n4517 0.0111456
R18538 VDD.n4776 VDD.n4775 0.0111456
R18539 VDD.n5034 VDD.n5033 0.0111456
R18540 VDD.n5292 VDD.n5291 0.0111456
R18541 VDD.n255 VDD.n254 0.0108947
R18542 VDD.n1396 VDD.n1394 0.0108723
R18543 VDD.n1381 VDD.n1377 0.0108723
R18544 VDD.n1957 VDD.n1922 0.0108144
R18545 VDD.n371 VDD.n370 0.0106316
R18546 VDD.n328 VDD.n327 0.0106316
R18547 VDD.n1327 VDD.n1325 0.0106064
R18548 VDD.n538 VDD.n537 0.0103684
R18549 VDD.n660 VDD.n659 0.0103684
R18550 VDD.n888 VDD.n887 0.0103684
R18551 VDD.n1010 VDD.n1009 0.0103684
R18552 VDD.n1426 VDD.n1425 0.0103404
R18553 VDD.n1511 VDD.n1510 0.0103404
R18554 VDD.n1527 VDD.n1526 0.0103039
R18555 VDD.n1696 VDD.n1695 0.0101514
R18556 VDD.n2045 VDD.n2044 0.0101514
R18557 VDD.n2275 VDD.n2274 0.0101514
R18558 VDD.n2533 VDD.n2532 0.0101514
R18559 VDD.n2791 VDD.n2790 0.0101514
R18560 VDD.n3049 VDD.n3048 0.0101514
R18561 VDD.n3307 VDD.n3306 0.0101514
R18562 VDD.n5630 VDD.n5629 0.0101514
R18563 VDD.n5376 VDD.n5375 0.0101514
R18564 VDD.n3565 VDD.n3564 0.0101514
R18565 VDD.n3823 VDD.n3822 0.0101514
R18566 VDD.n4081 VDD.n4080 0.0101514
R18567 VDD.n4339 VDD.n4338 0.0101514
R18568 VDD.n4597 VDD.n4596 0.0101514
R18569 VDD.n4855 VDD.n4854 0.0101514
R18570 VDD.n5113 VDD.n5112 0.0101514
R18571 VDD.n776 VDD.n775 0.0101053
R18572 VDD.n733 VDD.n732 0.0101053
R18573 VDD.n1126 VDD.n1125 0.0101053
R18574 VDD.n1083 VDD.n1082 0.0101053
R18575 VDD.n1883 VDD.n1882 0.0101
R18576 VDD.n2204 VDD.n2203 0.0101
R18577 VDD.n2462 VDD.n2461 0.0101
R18578 VDD.n2720 VDD.n2719 0.0101
R18579 VDD.n2978 VDD.n2977 0.0101
R18580 VDD.n3236 VDD.n3235 0.0101
R18581 VDD.n3494 VDD.n3493 0.0101
R18582 VDD.n5814 VDD.n5813 0.0101
R18583 VDD.n5560 VDD.n5559 0.0101
R18584 VDD.n3752 VDD.n3751 0.0101
R18585 VDD.n4010 VDD.n4009 0.0101
R18586 VDD.n4268 VDD.n4267 0.0101
R18587 VDD.n4526 VDD.n4525 0.0101
R18588 VDD.n4784 VDD.n4783 0.0101
R18589 VDD.n5042 VDD.n5041 0.0101
R18590 VDD.n5300 VDD.n5299 0.0101
R18591 VDD.n1597 VDD.n1181 0.00985484
R18592 VDD.n137 VDD.n136 0.00984211
R18593 VDD.n2129 VDD.n2128 0.00977468
R18594 VDD.n1884 VDD.n1883 0.0096003
R18595 VDD.n1870 VDD.n1869 0.0096003
R18596 VDD.n1869 VDD.t466 0.0096003
R18597 VDD.n2191 VDD.n2190 0.0096003
R18598 VDD.n2190 VDD.t592 0.0096003
R18599 VDD.n2205 VDD.n2204 0.0096003
R18600 VDD.n2449 VDD.n2448 0.0096003
R18601 VDD.n2448 VDD.t521 0.0096003
R18602 VDD.n2463 VDD.n2462 0.0096003
R18603 VDD.n2707 VDD.n2706 0.0096003
R18604 VDD.n2706 VDD.t278 0.0096003
R18605 VDD.n2721 VDD.n2720 0.0096003
R18606 VDD.n2965 VDD.n2964 0.0096003
R18607 VDD.n2964 VDD.t368 0.0096003
R18608 VDD.n2979 VDD.n2978 0.0096003
R18609 VDD.n3223 VDD.n3222 0.0096003
R18610 VDD.n3222 VDD.t1087 0.0096003
R18611 VDD.n3237 VDD.n3236 0.0096003
R18612 VDD.n3481 VDD.n3480 0.0096003
R18613 VDD.n3480 VDD.t1093 0.0096003
R18614 VDD.n3495 VDD.n3494 0.0096003
R18615 VDD.n5801 VDD.n5800 0.0096003
R18616 VDD.n5800 VDD.t514 0.0096003
R18617 VDD.n5815 VDD.n5814 0.0096003
R18618 VDD.n5547 VDD.n5546 0.0096003
R18619 VDD.n5546 VDD.t507 0.0096003
R18620 VDD.n5561 VDD.n5560 0.0096003
R18621 VDD.n3739 VDD.n3738 0.0096003
R18622 VDD.n3738 VDD.t251 0.0096003
R18623 VDD.n3753 VDD.n3752 0.0096003
R18624 VDD.n3997 VDD.n3996 0.0096003
R18625 VDD.n3996 VDD.t266 0.0096003
R18626 VDD.n4011 VDD.n4010 0.0096003
R18627 VDD.n4255 VDD.n4254 0.0096003
R18628 VDD.n4254 VDD.t13 0.0096003
R18629 VDD.n4269 VDD.n4268 0.0096003
R18630 VDD.n4513 VDD.n4512 0.0096003
R18631 VDD.n4512 VDD.t415 0.0096003
R18632 VDD.n4527 VDD.n4526 0.0096003
R18633 VDD.n4771 VDD.n4770 0.0096003
R18634 VDD.n4770 VDD.t527 0.0096003
R18635 VDD.n4785 VDD.n4784 0.0096003
R18636 VDD.n5029 VDD.n5028 0.0096003
R18637 VDD.n5028 VDD.t815 0.0096003
R18638 VDD.n5043 VDD.n5042 0.0096003
R18639 VDD.n5287 VDD.n5286 0.0096003
R18640 VDD.n5286 VDD.t265 0.0096003
R18641 VDD.n5301 VDD.n5300 0.0096003
R18642 VDD.t277 VDD.n1891 0.00959985
R18643 VDD.n1891 VDD.n1889 0.00959985
R18644 VDD.t494 VDD.n2212 0.00959985
R18645 VDD.n2212 VDD.n2210 0.00959985
R18646 VDD.t505 VDD.n2470 0.00959985
R18647 VDD.n2470 VDD.n2468 0.00959985
R18648 VDD.t1023 VDD.n2728 0.00959985
R18649 VDD.n2728 VDD.n2726 0.00959985
R18650 VDD.t524 VDD.n2986 0.00959985
R18651 VDD.n2986 VDD.n2984 0.00959985
R18652 VDD.t282 VDD.n3244 0.00959985
R18653 VDD.n3244 VDD.n3242 0.00959985
R18654 VDD.t419 VDD.n3502 0.00959985
R18655 VDD.n3502 VDD.n3500 0.00959985
R18656 VDD.t1075 VDD.n5822 0.00959985
R18657 VDD.n5822 VDD.n5820 0.00959985
R18658 VDD.t393 VDD.n5568 0.00959985
R18659 VDD.n5568 VDD.n5566 0.00959985
R18660 VDD.t262 VDD.n3760 0.00959985
R18661 VDD.n3760 VDD.n3758 0.00959985
R18662 VDD.t1084 VDD.n4018 0.00959985
R18663 VDD.n4018 VDD.n4016 0.00959985
R18664 VDD.t1021 VDD.n4276 0.00959985
R18665 VDD.n4276 VDD.n4274 0.00959985
R18666 VDD.t531 VDD.n4534 0.00959985
R18667 VDD.n4534 VDD.n4532 0.00959985
R18668 VDD.t401 VDD.n4792 0.00959985
R18669 VDD.n4792 VDD.n4790 0.00959985
R18670 VDD.t416 VDD.n5050 0.00959985
R18671 VDD.n5050 VDD.n5048 0.00959985
R18672 VDD.t407 VDD.n5308 0.00959985
R18673 VDD.n5308 VDD.n5306 0.00959985
R18674 VDD.n1361 VDD 0.00954255
R18675 VDD.n461 VDD.n458 0.0095362
R18676 VDD.n58 VDD.n55 0.0095362
R18677 VDD.n1425 VDD.n1423 0.0092766
R18678 VDD.n489 VDD.n467 0.00906279
R18679 VDD.n87 VDD.n65 0.00906279
R18680 VDD.n176 VDD.n175 0.00905263
R18681 VDD.n1283 VDD.n1282 0.00883333
R18682 VDD.n1282 VDD.n1280 0.00883333
R18683 VDD.n1280 VDD.n1276 0.00883333
R18684 VDD.n1276 VDD.n1274 0.00883333
R18685 VDD.n1274 VDD.n1270 0.00883333
R18686 VDD.n1295 VDD.n1291 0.00883333
R18687 VDD.n1297 VDD.n1295 0.00883333
R18688 VDD.n1301 VDD.n1297 0.00883333
R18689 VDD.n1303 VDD.n1301 0.00883333
R18690 VDD.n788 VDD.n784 0.00878947
R18691 VDD.n743 VDD.n741 0.00878947
R18692 VDD.n685 VDD.n683 0.00878947
R18693 VDD.n1138 VDD.n1134 0.00878947
R18694 VDD.n1093 VDD.n1091 0.00878947
R18695 VDD.n1035 VDD.n1033 0.00878947
R18696 VDD.n1399 VDD.n1396 0.00874468
R18697 VDD.n577 VDD.n576 0.00852632
R18698 VDD.n590 VDD.n589 0.00852632
R18699 VDD.n635 VDD.n634 0.00852632
R18700 VDD.n927 VDD.n926 0.00852632
R18701 VDD.n940 VDD.n939 0.00852632
R18702 VDD.n985 VDD.n984 0.00852632
R18703 VDD.n2128 VDD.n2127 0.00849839
R18704 VDD.n1287 VDD 0.00847872
R18705 VDD.n1742 VDD.n1741 0.0084202
R18706 VDD.n1699 VDD.n1698 0.0084202
R18707 VDD.n1698 VDD.t1031 0.0084202
R18708 VDD.n1676 VDD.n1672 0.0084202
R18709 VDD.n1764 VDD.n1676 0.0084202
R18710 VDD.n1766 VDD.n1765 0.0084202
R18711 VDD.n1765 VDD.n1764 0.0084202
R18712 VDD.n2091 VDD.n2090 0.0084202
R18713 VDD.n2048 VDD.n2047 0.0084202
R18714 VDD.n2047 VDD.t1264 0.0084202
R18715 VDD.n2025 VDD.n2021 0.0084202
R18716 VDD.n2113 VDD.n2025 0.0084202
R18717 VDD.n2115 VDD.n2114 0.0084202
R18718 VDD.n2114 VDD.n2113 0.0084202
R18719 VDD.n2321 VDD.n2320 0.0084202
R18720 VDD.n2278 VDD.n2277 0.0084202
R18721 VDD.n2277 VDD.t831 0.0084202
R18722 VDD.n2255 VDD.n2251 0.0084202
R18723 VDD.n2343 VDD.n2255 0.0084202
R18724 VDD.n2345 VDD.n2344 0.0084202
R18725 VDD.n2344 VDD.n2343 0.0084202
R18726 VDD.n2579 VDD.n2578 0.0084202
R18727 VDD.n2536 VDD.n2535 0.0084202
R18728 VDD.n2535 VDD.t1417 0.0084202
R18729 VDD.n2513 VDD.n2509 0.0084202
R18730 VDD.n2601 VDD.n2513 0.0084202
R18731 VDD.n2603 VDD.n2602 0.0084202
R18732 VDD.n2602 VDD.n2601 0.0084202
R18733 VDD.n2837 VDD.n2836 0.0084202
R18734 VDD.n2794 VDD.n2793 0.0084202
R18735 VDD.n2793 VDD.t436 0.0084202
R18736 VDD.n2771 VDD.n2767 0.0084202
R18737 VDD.n2859 VDD.n2771 0.0084202
R18738 VDD.n2861 VDD.n2860 0.0084202
R18739 VDD.n2860 VDD.n2859 0.0084202
R18740 VDD.n3095 VDD.n3094 0.0084202
R18741 VDD.n3052 VDD.n3051 0.0084202
R18742 VDD.n3051 VDD.t383 0.0084202
R18743 VDD.n3029 VDD.n3025 0.0084202
R18744 VDD.n3117 VDD.n3029 0.0084202
R18745 VDD.n3119 VDD.n3118 0.0084202
R18746 VDD.n3118 VDD.n3117 0.0084202
R18747 VDD.n3353 VDD.n3352 0.0084202
R18748 VDD.n3310 VDD.n3309 0.0084202
R18749 VDD.n3309 VDD.t1295 0.0084202
R18750 VDD.n3287 VDD.n3283 0.0084202
R18751 VDD.n3375 VDD.n3287 0.0084202
R18752 VDD.n3377 VDD.n3376 0.0084202
R18753 VDD.n3376 VDD.n3375 0.0084202
R18754 VDD.n5676 VDD.n5675 0.0084202
R18755 VDD.n5633 VDD.n5632 0.0084202
R18756 VDD.n5632 VDD.t476 0.0084202
R18757 VDD.n5610 VDD.n5606 0.0084202
R18758 VDD.n5698 VDD.n5610 0.0084202
R18759 VDD.n5700 VDD.n5699 0.0084202
R18760 VDD.n5699 VDD.n5698 0.0084202
R18761 VDD.n5422 VDD.n5421 0.0084202
R18762 VDD.n5379 VDD.n5378 0.0084202
R18763 VDD.n5378 VDD.t1258 0.0084202
R18764 VDD.n5356 VDD.n5352 0.0084202
R18765 VDD.n5444 VDD.n5356 0.0084202
R18766 VDD.n5446 VDD.n5445 0.0084202
R18767 VDD.n5445 VDD.n5444 0.0084202
R18768 VDD.n3611 VDD.n3610 0.0084202
R18769 VDD.n3568 VDD.n3567 0.0084202
R18770 VDD.n3567 VDD.t1366 0.0084202
R18771 VDD.n3545 VDD.n3541 0.0084202
R18772 VDD.n3633 VDD.n3545 0.0084202
R18773 VDD.n3635 VDD.n3634 0.0084202
R18774 VDD.n3634 VDD.n3633 0.0084202
R18775 VDD.n3869 VDD.n3868 0.0084202
R18776 VDD.n3826 VDD.n3825 0.0084202
R18777 VDD.n3825 VDD.t1114 0.0084202
R18778 VDD.n3803 VDD.n3799 0.0084202
R18779 VDD.n3891 VDD.n3803 0.0084202
R18780 VDD.n3893 VDD.n3892 0.0084202
R18781 VDD.n3892 VDD.n3891 0.0084202
R18782 VDD.n4127 VDD.n4126 0.0084202
R18783 VDD.n4084 VDD.n4083 0.0084202
R18784 VDD.n4083 VDD.t30 0.0084202
R18785 VDD.n4061 VDD.n4057 0.0084202
R18786 VDD.n4149 VDD.n4061 0.0084202
R18787 VDD.n4151 VDD.n4150 0.0084202
R18788 VDD.n4150 VDD.n4149 0.0084202
R18789 VDD.n4385 VDD.n4384 0.0084202
R18790 VDD.n4342 VDD.n4341 0.0084202
R18791 VDD.n4341 VDD.t1436 0.0084202
R18792 VDD.n4319 VDD.n4315 0.0084202
R18793 VDD.n4407 VDD.n4319 0.0084202
R18794 VDD.n4409 VDD.n4408 0.0084202
R18795 VDD.n4408 VDD.n4407 0.0084202
R18796 VDD.n4643 VDD.n4642 0.0084202
R18797 VDD.n4600 VDD.n4599 0.0084202
R18798 VDD.n4599 VDD.t370 0.0084202
R18799 VDD.n4577 VDD.n4573 0.0084202
R18800 VDD.n4665 VDD.n4577 0.0084202
R18801 VDD.n4667 VDD.n4666 0.0084202
R18802 VDD.n4666 VDD.n4665 0.0084202
R18803 VDD.n4901 VDD.n4900 0.0084202
R18804 VDD.n4858 VDD.n4857 0.0084202
R18805 VDD.n4857 VDD.t422 0.0084202
R18806 VDD.n4835 VDD.n4831 0.0084202
R18807 VDD.n4923 VDD.n4835 0.0084202
R18808 VDD.n4925 VDD.n4924 0.0084202
R18809 VDD.n4924 VDD.n4923 0.0084202
R18810 VDD.n5159 VDD.n5158 0.0084202
R18811 VDD.n5116 VDD.n5115 0.0084202
R18812 VDD.n5115 VDD.t0 0.0084202
R18813 VDD.n5093 VDD.n5089 0.0084202
R18814 VDD.n5181 VDD.n5093 0.0084202
R18815 VDD.n5183 VDD.n5182 0.0084202
R18816 VDD.n5182 VDD.n5181 0.0084202
R18817 VDD.n1615 VDD.n1614 0.0083125
R18818 VDD.n383 VDD.n379 0.00826316
R18819 VDD.n338 VDD.n336 0.00826316
R18820 VDD.n280 VDD.n278 0.00826316
R18821 VDD.n1366 VDD.n1365 0.00821277
R18822 VDD.n396 VDD.n395 0.00802802
R18823 VDD.n1554 VDD.n1553 0.00802802
R18824 VDD.n189 VDD.n188 0.008
R18825 VDD.n234 VDD.n233 0.008
R18826 VDD.n260 VDD.n259 0.008
R18827 VDD.n424 VDD.n421 0.00775202
R18828 VDD.n403 VDD.n400 0.00775202
R18829 VDD.n1582 VDD.n1579 0.00775202
R18830 VDD.n1561 VDD.n1558 0.00775202
R18831 VDD.n376 VDD.n375 0.00773684
R18832 VDD.n331 VDD.n330 0.00773684
R18833 VDD.n582 VDD.n540 0.00747368
R18834 VDD.n665 VDD.n664 0.00747368
R18835 VDD.n932 VDD.n890 0.00747368
R18836 VDD.n1015 VDD.n1014 0.00747368
R18837 VDD VDD.n1320 0.00741489
R18838 VDD.n781 VDD.n780 0.00721053
R18839 VDD.n736 VDD.n735 0.00721053
R18840 VDD.n1131 VDD.n1130 0.00721053
R18841 VDD.n1086 VDD.n1085 0.00721053
R18842 VDD.n1543 VDD 0.00714063
R18843 VDD.n1743 VDD.n1742 0.00702894
R18844 VDD.n2092 VDD.n2091 0.00702894
R18845 VDD.n2322 VDD.n2321 0.00702894
R18846 VDD.n2580 VDD.n2579 0.00702894
R18847 VDD.n2838 VDD.n2837 0.00702894
R18848 VDD.n3096 VDD.n3095 0.00702894
R18849 VDD.n3354 VDD.n3353 0.00702894
R18850 VDD.n5677 VDD.n5676 0.00702894
R18851 VDD.n5423 VDD.n5422 0.00702894
R18852 VDD.n3612 VDD.n3611 0.00702894
R18853 VDD.n3870 VDD.n3869 0.00702894
R18854 VDD.n4128 VDD.n4127 0.00702894
R18855 VDD.n4386 VDD.n4385 0.00702894
R18856 VDD.n4644 VDD.n4643 0.00702894
R18857 VDD.n4902 VDD.n4901 0.00702894
R18858 VDD.n5160 VDD.n5159 0.00702894
R18859 VDD.n1291 VDD.n1246 0.00702174
R18860 VDD.n816 VDD 0.00700289
R18861 VDD.n1199 VDD 0.00700289
R18862 VDD.n181 VDD.n139 0.00694737
R18863 VDD.n1829 VDD.n1828 0.00693382
R18864 VDD.n2150 VDD.n2149 0.00693382
R18865 VDD.n2408 VDD.n2407 0.00693382
R18866 VDD.n2666 VDD.n2665 0.00693382
R18867 VDD.n2924 VDD.n2923 0.00693382
R18868 VDD.n3182 VDD.n3181 0.00693382
R18869 VDD.n3440 VDD.n3439 0.00693382
R18870 VDD.n5760 VDD.n5759 0.00693382
R18871 VDD.n5506 VDD.n5505 0.00693382
R18872 VDD.n3698 VDD.n3697 0.00693382
R18873 VDD.n3956 VDD.n3955 0.00693382
R18874 VDD.n4214 VDD.n4213 0.00693382
R18875 VDD.n4472 VDD.n4471 0.00693382
R18876 VDD.n4730 VDD.n4729 0.00693382
R18877 VDD.n4988 VDD.n4987 0.00693382
R18878 VDD.n5246 VDD.n5245 0.00693382
R18879 VDD.n1181 VDD.n1180 0.00681452
R18880 VDD.n809 VDD 0.00675
R18881 VDD.n1192 VDD 0.00675
R18882 VDD.n1540 VDD.n1255 0.00662745
R18883 VDD.n1463 VDD.n1461 0.00661702
R18884 VDD VDD.n551 0.00655263
R18885 VDD.n622 VDD 0.00655263
R18886 VDD VDD.n791 0.00655263
R18887 VDD VDD.n744 0.00655263
R18888 VDD VDD.n697 0.00655263
R18889 VDD.n677 VDD 0.00655263
R18890 VDD VDD.n901 0.00655263
R18891 VDD.n972 VDD 0.00655263
R18892 VDD VDD.n1141 0.00655263
R18893 VDD VDD.n1094 0.00655263
R18894 VDD VDD.n1047 0.00655263
R18895 VDD.n1027 VDD 0.00655263
R18896 VDD VDD.n150 0.00655263
R18897 VDD.n221 VDD 0.00655263
R18898 VDD VDD.n386 0.00655263
R18899 VDD VDD.n339 0.00655263
R18900 VDD VDD.n292 0.00655263
R18901 VDD.n272 VDD 0.00655263
R18902 VDD.n794 VDD.n35 0.00638056
R18903 VDD.n181 VDD.n180 0.00615789
R18904 VDD VDD.n808 0.00609211
R18905 VDD VDD.n1191 0.00609211
R18906 VDD.n1739 VDD.n1736 0.00605556
R18907 VDD.n2088 VDD.n2085 0.00605556
R18908 VDD.n2318 VDD.n2315 0.00605556
R18909 VDD.n2576 VDD.n2573 0.00605556
R18910 VDD.n2834 VDD.n2831 0.00605556
R18911 VDD.n3092 VDD.n3089 0.00605556
R18912 VDD.n3350 VDD.n3347 0.00605556
R18913 VDD.n5673 VDD.n5670 0.00605556
R18914 VDD.n5419 VDD.n5416 0.00605556
R18915 VDD.n3608 VDD.n3605 0.00605556
R18916 VDD.n3866 VDD.n3863 0.00605556
R18917 VDD.n4124 VDD.n4121 0.00605556
R18918 VDD.n4382 VDD.n4379 0.00605556
R18919 VDD.n4640 VDD.n4637 0.00605556
R18920 VDD.n4898 VDD.n4895 0.00605556
R18921 VDD.n5156 VDD.n5153 0.00605556
R18922 VDD.n783 VDD.n781 0.00589474
R18923 VDD.n740 VDD.n736 0.00589474
R18924 VDD.n1133 VDD.n1131 0.00589474
R18925 VDD.n1090 VDD.n1086 0.00589474
R18926 VDD.n1343 VDD.n1320 0.00581915
R18927 VDD.n1982 VDD.n1981 0.00573228
R18928 VDD.n1982 VDD.n1980 0.00573228
R18929 VDD.n1540 VDD.n1539 0.00564706
R18930 VDD.n582 VDD.n581 0.00563158
R18931 VDD.n665 VDD.n637 0.00563158
R18932 VDD.n686 VDD 0.00563158
R18933 VDD.n932 VDD.n931 0.00563158
R18934 VDD.n1015 VDD.n987 0.00563158
R18935 VDD.n1036 VDD 0.00563158
R18936 VDD.n1376 VDD.n1374 0.00552129
R18937 VDD.n1603 VDD.n1602 0.00542857
R18938 VDD.n378 VDD.n376 0.00536842
R18939 VDD.n335 VDD.n331 0.00536842
R18940 VDD.n1617 VDD.n1615 0.0051875
R18941 VDD.n193 VDD.n189 0.00510526
R18942 VDD.n236 VDD.n234 0.00510526
R18943 VDD.n260 VDD.n236 0.00510526
R18944 VDD.n281 VDD 0.00510526
R18945 VDD.n1913 VDD.n1912 0.00505015
R18946 VDD.t277 VDD.n1913 0.00505015
R18947 VDD.t277 VDD.n1894 0.00505015
R18948 VDD.n1909 VDD.n1894 0.00505015
R18949 VDD.n1824 VDD.n1823 0.00505015
R18950 VDD.n1861 VDD.n1848 0.00505015
R18951 VDD.t466 VDD.n1848 0.00505015
R18952 VDD.n1868 VDD.n1867 0.00505015
R18953 VDD.t466 VDD.n1868 0.00505015
R18954 VDD.n2182 VDD.n2169 0.00505015
R18955 VDD.t592 VDD.n2169 0.00505015
R18956 VDD.n2189 VDD.n2188 0.00505015
R18957 VDD.t592 VDD.n2189 0.00505015
R18958 VDD.n2145 VDD.n2144 0.00505015
R18959 VDD.n2234 VDD.n2233 0.00505015
R18960 VDD.t494 VDD.n2234 0.00505015
R18961 VDD.t494 VDD.n2215 0.00505015
R18962 VDD.n2230 VDD.n2215 0.00505015
R18963 VDD.n2440 VDD.n2427 0.00505015
R18964 VDD.t521 VDD.n2427 0.00505015
R18965 VDD.n2447 VDD.n2446 0.00505015
R18966 VDD.t521 VDD.n2447 0.00505015
R18967 VDD.n2403 VDD.n2402 0.00505015
R18968 VDD.n2492 VDD.n2491 0.00505015
R18969 VDD.t505 VDD.n2492 0.00505015
R18970 VDD.t505 VDD.n2473 0.00505015
R18971 VDD.n2488 VDD.n2473 0.00505015
R18972 VDD.n2698 VDD.n2685 0.00505015
R18973 VDD.t278 VDD.n2685 0.00505015
R18974 VDD.n2705 VDD.n2704 0.00505015
R18975 VDD.t278 VDD.n2705 0.00505015
R18976 VDD.n2661 VDD.n2660 0.00505015
R18977 VDD.n2750 VDD.n2749 0.00505015
R18978 VDD.t1023 VDD.n2750 0.00505015
R18979 VDD.t1023 VDD.n2731 0.00505015
R18980 VDD.n2746 VDD.n2731 0.00505015
R18981 VDD.n2956 VDD.n2943 0.00505015
R18982 VDD.t368 VDD.n2943 0.00505015
R18983 VDD.n2963 VDD.n2962 0.00505015
R18984 VDD.t368 VDD.n2963 0.00505015
R18985 VDD.n2919 VDD.n2918 0.00505015
R18986 VDD.n3008 VDD.n3007 0.00505015
R18987 VDD.t524 VDD.n3008 0.00505015
R18988 VDD.t524 VDD.n2989 0.00505015
R18989 VDD.n3004 VDD.n2989 0.00505015
R18990 VDD.n3214 VDD.n3201 0.00505015
R18991 VDD.t1087 VDD.n3201 0.00505015
R18992 VDD.n3221 VDD.n3220 0.00505015
R18993 VDD.t1087 VDD.n3221 0.00505015
R18994 VDD.n3177 VDD.n3176 0.00505015
R18995 VDD.n3266 VDD.n3265 0.00505015
R18996 VDD.t282 VDD.n3266 0.00505015
R18997 VDD.t282 VDD.n3247 0.00505015
R18998 VDD.n3262 VDD.n3247 0.00505015
R18999 VDD.n3472 VDD.n3459 0.00505015
R19000 VDD.t1093 VDD.n3459 0.00505015
R19001 VDD.n3479 VDD.n3478 0.00505015
R19002 VDD.t1093 VDD.n3479 0.00505015
R19003 VDD.n3435 VDD.n3434 0.00505015
R19004 VDD.n3524 VDD.n3523 0.00505015
R19005 VDD.t419 VDD.n3524 0.00505015
R19006 VDD.t419 VDD.n3505 0.00505015
R19007 VDD.n3520 VDD.n3505 0.00505015
R19008 VDD.n5792 VDD.n5779 0.00505015
R19009 VDD.t514 VDD.n5779 0.00505015
R19010 VDD.n5799 VDD.n5798 0.00505015
R19011 VDD.t514 VDD.n5799 0.00505015
R19012 VDD.n5755 VDD.n5754 0.00505015
R19013 VDD.n5844 VDD.n5843 0.00505015
R19014 VDD.t1075 VDD.n5844 0.00505015
R19015 VDD.t1075 VDD.n5825 0.00505015
R19016 VDD.n5840 VDD.n5825 0.00505015
R19017 VDD.n5538 VDD.n5525 0.00505015
R19018 VDD.t507 VDD.n5525 0.00505015
R19019 VDD.n5545 VDD.n5544 0.00505015
R19020 VDD.t507 VDD.n5545 0.00505015
R19021 VDD.n5501 VDD.n5500 0.00505015
R19022 VDD.n5590 VDD.n5589 0.00505015
R19023 VDD.t393 VDD.n5590 0.00505015
R19024 VDD.t393 VDD.n5571 0.00505015
R19025 VDD.n5586 VDD.n5571 0.00505015
R19026 VDD.n3730 VDD.n3717 0.00505015
R19027 VDD.t251 VDD.n3717 0.00505015
R19028 VDD.n3737 VDD.n3736 0.00505015
R19029 VDD.t251 VDD.n3737 0.00505015
R19030 VDD.n3693 VDD.n3692 0.00505015
R19031 VDD.n3782 VDD.n3781 0.00505015
R19032 VDD.t262 VDD.n3782 0.00505015
R19033 VDD.t262 VDD.n3763 0.00505015
R19034 VDD.n3778 VDD.n3763 0.00505015
R19035 VDD.n3988 VDD.n3975 0.00505015
R19036 VDD.t266 VDD.n3975 0.00505015
R19037 VDD.n3995 VDD.n3994 0.00505015
R19038 VDD.t266 VDD.n3995 0.00505015
R19039 VDD.n3951 VDD.n3950 0.00505015
R19040 VDD.n4040 VDD.n4039 0.00505015
R19041 VDD.t1084 VDD.n4040 0.00505015
R19042 VDD.t1084 VDD.n4021 0.00505015
R19043 VDD.n4036 VDD.n4021 0.00505015
R19044 VDD.n4246 VDD.n4233 0.00505015
R19045 VDD.t13 VDD.n4233 0.00505015
R19046 VDD.n4253 VDD.n4252 0.00505015
R19047 VDD.t13 VDD.n4253 0.00505015
R19048 VDD.n4209 VDD.n4208 0.00505015
R19049 VDD.n4298 VDD.n4297 0.00505015
R19050 VDD.t1021 VDD.n4298 0.00505015
R19051 VDD.t1021 VDD.n4279 0.00505015
R19052 VDD.n4294 VDD.n4279 0.00505015
R19053 VDD.n4504 VDD.n4491 0.00505015
R19054 VDD.t415 VDD.n4491 0.00505015
R19055 VDD.n4511 VDD.n4510 0.00505015
R19056 VDD.t415 VDD.n4511 0.00505015
R19057 VDD.n4467 VDD.n4466 0.00505015
R19058 VDD.n4556 VDD.n4555 0.00505015
R19059 VDD.t531 VDD.n4556 0.00505015
R19060 VDD.t531 VDD.n4537 0.00505015
R19061 VDD.n4552 VDD.n4537 0.00505015
R19062 VDD.n4762 VDD.n4749 0.00505015
R19063 VDD.t527 VDD.n4749 0.00505015
R19064 VDD.n4769 VDD.n4768 0.00505015
R19065 VDD.t527 VDD.n4769 0.00505015
R19066 VDD.n4725 VDD.n4724 0.00505015
R19067 VDD.n4814 VDD.n4813 0.00505015
R19068 VDD.t401 VDD.n4814 0.00505015
R19069 VDD.t401 VDD.n4795 0.00505015
R19070 VDD.n4810 VDD.n4795 0.00505015
R19071 VDD.n5020 VDD.n5007 0.00505015
R19072 VDD.t815 VDD.n5007 0.00505015
R19073 VDD.n5027 VDD.n5026 0.00505015
R19074 VDD.t815 VDD.n5027 0.00505015
R19075 VDD.n4983 VDD.n4982 0.00505015
R19076 VDD.n5072 VDD.n5071 0.00505015
R19077 VDD.t416 VDD.n5072 0.00505015
R19078 VDD.t416 VDD.n5053 0.00505015
R19079 VDD.n5068 VDD.n5053 0.00505015
R19080 VDD.n5278 VDD.n5265 0.00505015
R19081 VDD.t265 VDD.n5265 0.00505015
R19082 VDD.n5285 VDD.n5284 0.00505015
R19083 VDD.t265 VDD.n5285 0.00505015
R19084 VDD.n5241 VDD.n5240 0.00505015
R19085 VDD.n5330 VDD.n5329 0.00505015
R19086 VDD.t407 VDD.n5330 0.00505015
R19087 VDD.t407 VDD.n5311 0.00505015
R19088 VDD.n5326 VDD.n5311 0.00505015
R19089 VDD.n1311 VDD 0.00502128
R19090 VDD.n1340 VDD 0.00502128
R19091 VDD VDD.n1346 0.00502128
R19092 VDD.n1363 VDD 0.00502128
R19093 VDD.n1510 VDD 0.00502128
R19094 VDD.n379 VDD.n378 0.00484211
R19095 VDD.n336 VDD.n335 0.00484211
R19096 VDD.n278 VDD.n277 0.00484211
R19097 VDD.n1324 VDD.n1319 0.00475532
R19098 VDD VDD.n1509 0.00475532
R19099 VDD.n1504 VDD.n1261 0.00475532
R19100 VDD.n1287 VDD.n1286 0.00475532
R19101 VDD.n1751 VDD.n1722 0.00466667
R19102 VDD.n1703 VDD.n1702 0.00466667
R19103 VDD.n1692 VDD.n1691 0.00466667
R19104 VDD.n2100 VDD.n2071 0.00466667
R19105 VDD.n2052 VDD.n2051 0.00466667
R19106 VDD.n2041 VDD.n2040 0.00466667
R19107 VDD.n2330 VDD.n2301 0.00466667
R19108 VDD.n2282 VDD.n2281 0.00466667
R19109 VDD.n2271 VDD.n2270 0.00466667
R19110 VDD.n2588 VDD.n2559 0.00466667
R19111 VDD.n2540 VDD.n2539 0.00466667
R19112 VDD.n2529 VDD.n2528 0.00466667
R19113 VDD.n2846 VDD.n2817 0.00466667
R19114 VDD.n2798 VDD.n2797 0.00466667
R19115 VDD.n2787 VDD.n2786 0.00466667
R19116 VDD.n3104 VDD.n3075 0.00466667
R19117 VDD.n3056 VDD.n3055 0.00466667
R19118 VDD.n3045 VDD.n3044 0.00466667
R19119 VDD.n3362 VDD.n3333 0.00466667
R19120 VDD.n3314 VDD.n3313 0.00466667
R19121 VDD.n3303 VDD.n3302 0.00466667
R19122 VDD.n5685 VDD.n5656 0.00466667
R19123 VDD.n5637 VDD.n5636 0.00466667
R19124 VDD.n5626 VDD.n5625 0.00466667
R19125 VDD.n5431 VDD.n5402 0.00466667
R19126 VDD.n5383 VDD.n5382 0.00466667
R19127 VDD.n5372 VDD.n5371 0.00466667
R19128 VDD.n3620 VDD.n3591 0.00466667
R19129 VDD.n3572 VDD.n3571 0.00466667
R19130 VDD.n3561 VDD.n3560 0.00466667
R19131 VDD.n3878 VDD.n3849 0.00466667
R19132 VDD.n3830 VDD.n3829 0.00466667
R19133 VDD.n3819 VDD.n3818 0.00466667
R19134 VDD.n4136 VDD.n4107 0.00466667
R19135 VDD.n4088 VDD.n4087 0.00466667
R19136 VDD.n4077 VDD.n4076 0.00466667
R19137 VDD.n4394 VDD.n4365 0.00466667
R19138 VDD.n4346 VDD.n4345 0.00466667
R19139 VDD.n4335 VDD.n4334 0.00466667
R19140 VDD.n4652 VDD.n4623 0.00466667
R19141 VDD.n4604 VDD.n4603 0.00466667
R19142 VDD.n4593 VDD.n4592 0.00466667
R19143 VDD.n4910 VDD.n4881 0.00466667
R19144 VDD.n4862 VDD.n4861 0.00466667
R19145 VDD.n4851 VDD.n4850 0.00466667
R19146 VDD.n5168 VDD.n5139 0.00466667
R19147 VDD.n5120 VDD.n5119 0.00466667
R19148 VDD.n5109 VDD.n5108 0.00466667
R19149 VDD VDD.n35 0.00460833
R19150 VDD.n581 VDD.n577 0.00457895
R19151 VDD.n594 VDD.n590 0.00457895
R19152 VDD.n637 VDD.n635 0.00457895
R19153 VDD.n931 VDD.n927 0.00457895
R19154 VDD.n944 VDD.n940 0.00457895
R19155 VDD.n987 VDD.n985 0.00457895
R19156 VDD.n1547 VDD.n1546 0.00451563
R19157 VDD.n784 VDD.n783 0.00431579
R19158 VDD.n741 VDD.n740 0.00431579
R19159 VDD.n683 VDD.n682 0.00431579
R19160 VDD.n1134 VDD.n1133 0.00431579
R19161 VDD.n1091 VDD.n1090 0.00431579
R19162 VDD.n1033 VDD.n1032 0.00431579
R19163 VDD.n1406 VDD.n1405 0.0042234
R19164 VDD.n1304 VDD.n1303 0.00412319
R19165 VDD VDD.n809 0.00411272
R19166 VDD VDD.n1192 0.00411272
R19167 VDD.n1611 VDD.n1610 0.00410577
R19168 VDD.n180 VDD.n176 0.00405263
R19169 VDD.n512 VDD 0.00400806
R19170 VDD.n2125 VDD.n2013 0.00390318
R19171 VDD.n809 VDD 0.00378947
R19172 VDD.n1192 VDD 0.00378947
R19173 VDD.n1526 VDD.n1525 0.00369149
R19174 VDD.n1816 VDD.n1809 0.00364862
R19175 VDD.n2137 VDD.n2130 0.00364862
R19176 VDD.n2395 VDD.n2388 0.00364862
R19177 VDD.n2653 VDD.n2646 0.00364862
R19178 VDD.n2911 VDD.n2904 0.00364862
R19179 VDD.n3169 VDD.n3162 0.00364862
R19180 VDD.n3427 VDD.n3420 0.00364862
R19181 VDD.n5747 VDD.n5740 0.00364862
R19182 VDD.n5493 VDD.n5486 0.00364862
R19183 VDD.n3685 VDD.n3678 0.00364862
R19184 VDD.n3943 VDD.n3936 0.00364862
R19185 VDD.n4201 VDD.n4194 0.00364862
R19186 VDD.n4459 VDD.n4452 0.00364862
R19187 VDD.n4717 VDD.n4710 0.00364862
R19188 VDD.n4975 VDD.n4968 0.00364862
R19189 VDD.n5233 VDD.n5226 0.00364862
R19190 VDD.n1289 VDD 0.00342553
R19191 VDD.n1609 VDD.n1604 0.00339649
R19192 VDD VDD.n796 0.00330645
R19193 VDD.n139 VDD.n137 0.00326316
R19194 VDD.n1934 VDD.n1926 0.00317113
R19195 VDD.n1955 VDD.n1944 0.00317113
R19196 VDD.n1359 VDD.n1358 0.00315957
R19197 VDD.n1600 VDD 0.00304286
R19198 VDD.n780 VDD.n776 0.003
R19199 VDD.n735 VDD.n733 0.003
R19200 VDD.n1130 VDD.n1126 0.003
R19201 VDD.n1085 VDD.n1083 0.003
R19202 VDD.n1743 VDD.t441 0.00289124
R19203 VDD.n2092 VDD.t80 0.00289124
R19204 VDD.n2322 VDD.t1446 0.00289124
R19205 VDD.n2580 VDD.t567 0.00289124
R19206 VDD.n2838 VDD.t978 0.00289124
R19207 VDD.n3096 VDD.t545 0.00289124
R19208 VDD.n3354 VDD.t582 0.00289124
R19209 VDD.n5677 VDD.t1468 0.00289124
R19210 VDD.n5423 VDD.t995 0.00289124
R19211 VDD.n3612 VDD.t1336 0.00289124
R19212 VDD.n3870 VDD.t485 0.00289124
R19213 VDD.n4128 VDD.t5 0.00289124
R19214 VDD.n4386 VDD.t1052 0.00289124
R19215 VDD.n4644 VDD.t21 0.00289124
R19216 VDD.n4902 VDD.t563 0.00289124
R19217 VDD.n5160 VDD.t1008 0.00289124
R19218 VDD.n540 VDD.n538 0.00273684
R19219 VDD.n552 VDD 0.00273684
R19220 VDD.n619 VDD 0.00273684
R19221 VDD.n664 VDD.n660 0.00273684
R19222 VDD.n792 VDD 0.00273684
R19223 VDD.n745 VDD 0.00273684
R19224 VDD.n698 VDD 0.00273684
R19225 VDD.n680 VDD 0.00273684
R19226 VDD.n890 VDD.n888 0.00273684
R19227 VDD.n902 VDD 0.00273684
R19228 VDD.n969 VDD 0.00273684
R19229 VDD.n1014 VDD.n1010 0.00273684
R19230 VDD.n1142 VDD 0.00273684
R19231 VDD.n1095 VDD 0.00273684
R19232 VDD.n1048 VDD 0.00273684
R19233 VDD.n1030 VDD 0.00273684
R19234 VDD.n151 VDD 0.00273684
R19235 VDD.n218 VDD 0.00273684
R19236 VDD.n387 VDD 0.00273684
R19237 VDD.n340 VDD 0.00273684
R19238 VDD.n293 VDD 0.00273684
R19239 VDD.n275 VDD 0.00273684
R19240 VDD.n188 VDD.n186 0.00271053
R19241 VDD.n1926 VDD.n1925 0.00267116
R19242 VDD.n1956 VDD.n1955 0.00267116
R19243 VDD.n1506 VDD 0.00262766
R19244 VDD.n689 VDD.n688 0.00247368
R19245 VDD.n1039 VDD.n1038 0.00247368
R19246 VDD.n375 VDD.n371 0.00247368
R19247 VDD.n330 VDD.n328 0.00247368
R19248 VDD.n5859 VDD.n5858 0.00240789
R19249 VDD.n1838 VDD.n1837 0.00240766
R19250 VDD.n2159 VDD.n2158 0.00240766
R19251 VDD.n2417 VDD.n2416 0.00240766
R19252 VDD.n2675 VDD.n2674 0.00240766
R19253 VDD.n2933 VDD.n2932 0.00240766
R19254 VDD.n3191 VDD.n3190 0.00240766
R19255 VDD.n3449 VDD.n3448 0.00240766
R19256 VDD.n5769 VDD.n5768 0.00240766
R19257 VDD.n5515 VDD.n5514 0.00240766
R19258 VDD.n3707 VDD.n3706 0.00240766
R19259 VDD.n3965 VDD.n3964 0.00240766
R19260 VDD.n4223 VDD.n4222 0.00240766
R19261 VDD.n4481 VDD.n4480 0.00240766
R19262 VDD.n4739 VDD.n4738 0.00240766
R19263 VDD.n4997 VDD.n4996 0.00240766
R19264 VDD.n5255 VDD.n5254 0.00240766
R19265 VDD.n1601 VDD.n1600 0.00237143
R19266 VDD.n1359 VDD 0.0023617
R19267 VDD.n1369 VDD.n1368 0.0023617
R19268 VDD.n1829 VDD.n1825 0.00233824
R19269 VDD.n1831 VDD 0.00233824
R19270 VDD.n2150 VDD.n2146 0.00233824
R19271 VDD.n2152 VDD 0.00233824
R19272 VDD.n2408 VDD.n2404 0.00233824
R19273 VDD.n2410 VDD 0.00233824
R19274 VDD.n2666 VDD.n2662 0.00233824
R19275 VDD.n2668 VDD 0.00233824
R19276 VDD.n2924 VDD.n2920 0.00233824
R19277 VDD.n2926 VDD 0.00233824
R19278 VDD.n3182 VDD.n3178 0.00233824
R19279 VDD.n3184 VDD 0.00233824
R19280 VDD.n3440 VDD.n3436 0.00233824
R19281 VDD.n3442 VDD 0.00233824
R19282 VDD.n5760 VDD.n5756 0.00233824
R19283 VDD.n5762 VDD 0.00233824
R19284 VDD.n5506 VDD.n5502 0.00233824
R19285 VDD.n5508 VDD 0.00233824
R19286 VDD.n3698 VDD.n3694 0.00233824
R19287 VDD.n3700 VDD 0.00233824
R19288 VDD.n3956 VDD.n3952 0.00233824
R19289 VDD.n3958 VDD 0.00233824
R19290 VDD.n4214 VDD.n4210 0.00233824
R19291 VDD.n4216 VDD 0.00233824
R19292 VDD.n4472 VDD.n4468 0.00233824
R19293 VDD.n4474 VDD 0.00233824
R19294 VDD.n4730 VDD.n4726 0.00233824
R19295 VDD.n4732 VDD 0.00233824
R19296 VDD.n4988 VDD.n4984 0.00233824
R19297 VDD.n4990 VDD 0.00233824
R19298 VDD.n5246 VDD.n5242 0.00233824
R19299 VDD.n5248 VDD 0.00233824
R19300 VDD.n1454 VDD.n1317 0.00232979
R19301 VDD.n1431 VDD.n1319 0.00232979
R19302 VDD.n1879 VDD.t274 0.00231811
R19303 VDD.n2200 VDD.t511 0.00231811
R19304 VDD.n2458 VDD.t528 0.00231811
R19305 VDD.n2716 VDD.t1381 0.00231811
R19306 VDD.n2974 VDD.t414 0.00231811
R19307 VDD.n3232 VDD.t591 0.00231811
R19308 VDD.n3490 VDD.t1086 0.00231811
R19309 VDD.n5810 VDD.t276 0.00231811
R19310 VDD.n5556 VDD.t512 0.00231811
R19311 VDD.n3748 VDD.t1085 0.00231811
R19312 VDD.n4006 VDD.t526 0.00231811
R19313 VDD.n4264 VDD.t525 0.00231811
R19314 VDD.n4522 VDD.t264 0.00231811
R19315 VDD.n4780 VDD.t590 0.00231811
R19316 VDD.n5038 VDD.t1024 0.00231811
R19317 VDD.n5296 VDD.t275 0.00231811
R19318 VDD.n1270 VDD.n1246 0.00231159
R19319 VDD.n1726 VDD.n1724 0.00228571
R19320 VDD.n2075 VDD.n2073 0.00228571
R19321 VDD.n2305 VDD.n2303 0.00228571
R19322 VDD.n2563 VDD.n2561 0.00228571
R19323 VDD.n2821 VDD.n2819 0.00228571
R19324 VDD.n3079 VDD.n3077 0.00228571
R19325 VDD.n3337 VDD.n3335 0.00228571
R19326 VDD.n5660 VDD.n5658 0.00228571
R19327 VDD.n5406 VDD.n5404 0.00228571
R19328 VDD.n3595 VDD.n3593 0.00228571
R19329 VDD.n3853 VDD.n3851 0.00228571
R19330 VDD.n4111 VDD.n4109 0.00228571
R19331 VDD.n4369 VDD.n4367 0.00228571
R19332 VDD.n4627 VDD.n4625 0.00228571
R19333 VDD.n4885 VDD.n4883 0.00228571
R19334 VDD.n5143 VDD.n5141 0.00228571
R19335 VDD.n1694 VDD.n1693 0.00221302
R19336 VDD.n1695 VDD.n1694 0.00221302
R19337 VDD.n2043 VDD.n2042 0.00221302
R19338 VDD.n2044 VDD.n2043 0.00221302
R19339 VDD.n2273 VDD.n2272 0.00221302
R19340 VDD.n2274 VDD.n2273 0.00221302
R19341 VDD.n2531 VDD.n2530 0.00221302
R19342 VDD.n2532 VDD.n2531 0.00221302
R19343 VDD.n2789 VDD.n2788 0.00221302
R19344 VDD.n2790 VDD.n2789 0.00221302
R19345 VDD.n3047 VDD.n3046 0.00221302
R19346 VDD.n3048 VDD.n3047 0.00221302
R19347 VDD.n3305 VDD.n3304 0.00221302
R19348 VDD.n3306 VDD.n3305 0.00221302
R19349 VDD.n5628 VDD.n5627 0.00221302
R19350 VDD.n5629 VDD.n5628 0.00221302
R19351 VDD.n5374 VDD.n5373 0.00221302
R19352 VDD.n5375 VDD.n5374 0.00221302
R19353 VDD.n3563 VDD.n3562 0.00221302
R19354 VDD.n3564 VDD.n3563 0.00221302
R19355 VDD.n3821 VDD.n3820 0.00221302
R19356 VDD.n3822 VDD.n3821 0.00221302
R19357 VDD.n4079 VDD.n4078 0.00221302
R19358 VDD.n4080 VDD.n4079 0.00221302
R19359 VDD.n4337 VDD.n4336 0.00221302
R19360 VDD.n4338 VDD.n4337 0.00221302
R19361 VDD.n4595 VDD.n4594 0.00221302
R19362 VDD.n4596 VDD.n4595 0.00221302
R19363 VDD.n4853 VDD.n4852 0.00221302
R19364 VDD.n4854 VDD.n4853 0.00221302
R19365 VDD.n5111 VDD.n5110 0.00221302
R19366 VDD.n5112 VDD.n5111 0.00221302
R19367 VDD.n1693 VDD.n1692 0.00221271
R19368 VDD.n2042 VDD.n2041 0.00221271
R19369 VDD.n2272 VDD.n2271 0.00221271
R19370 VDD.n2530 VDD.n2529 0.00221271
R19371 VDD.n2788 VDD.n2787 0.00221271
R19372 VDD.n3046 VDD.n3045 0.00221271
R19373 VDD.n3304 VDD.n3303 0.00221271
R19374 VDD.n5627 VDD.n5626 0.00221271
R19375 VDD.n5373 VDD.n5372 0.00221271
R19376 VDD.n3562 VDD.n3561 0.00221271
R19377 VDD.n3820 VDD.n3819 0.00221271
R19378 VDD.n4078 VDD.n4077 0.00221271
R19379 VDD.n4336 VDD.n4335 0.00221271
R19380 VDD.n4594 VDD.n4593 0.00221271
R19381 VDD.n4852 VDD.n4851 0.00221271
R19382 VDD.n5110 VDD.n5109 0.00221271
R19383 VDD.n259 VDD.n255 0.00221053
R19384 VDD.n1732 VDD.n1730 0.00220611
R19385 VDD.n2081 VDD.n2079 0.00220611
R19386 VDD.n2311 VDD.n2309 0.00220611
R19387 VDD.n2569 VDD.n2567 0.00220611
R19388 VDD.n2827 VDD.n2825 0.00220611
R19389 VDD.n3085 VDD.n3083 0.00220611
R19390 VDD.n3343 VDD.n3341 0.00220611
R19391 VDD.n5666 VDD.n5664 0.00220611
R19392 VDD.n5412 VDD.n5410 0.00220611
R19393 VDD.n3601 VDD.n3599 0.00220611
R19394 VDD.n3859 VDD.n3857 0.00220611
R19395 VDD.n4117 VDD.n4115 0.00220611
R19396 VDD.n4375 VDD.n4373 0.00220611
R19397 VDD.n4633 VDD.n4631 0.00220611
R19398 VDD.n4891 VDD.n4889 0.00220611
R19399 VDD.n5149 VDD.n5147 0.00220611
R19400 VDD.n1702 VDD.n1681 0.0022058
R19401 VDD.n2051 VDD.n2030 0.0022058
R19402 VDD.n2281 VDD.n2260 0.0022058
R19403 VDD.n2539 VDD.n2518 0.0022058
R19404 VDD.n2797 VDD.n2776 0.0022058
R19405 VDD.n3055 VDD.n3034 0.0022058
R19406 VDD.n3313 VDD.n3292 0.0022058
R19407 VDD.n5636 VDD.n5615 0.0022058
R19408 VDD.n5382 VDD.n5361 0.0022058
R19409 VDD.n3571 VDD.n3550 0.0022058
R19410 VDD.n3829 VDD.n3808 0.0022058
R19411 VDD.n4087 VDD.n4066 0.0022058
R19412 VDD.n4345 VDD.n4324 0.0022058
R19413 VDD.n4603 VDD.n4582 0.0022058
R19414 VDD.n4861 VDD.n4840 0.0022058
R19415 VDD.n5119 VDD.n5098 0.0022058
R19416 VDD.n1745 VDD.n1724 0.0022058
R19417 VDD.n2094 VDD.n2073 0.0022058
R19418 VDD.n2324 VDD.n2303 0.0022058
R19419 VDD.n2582 VDD.n2561 0.0022058
R19420 VDD.n2840 VDD.n2819 0.0022058
R19421 VDD.n3098 VDD.n3077 0.0022058
R19422 VDD.n3356 VDD.n3335 0.0022058
R19423 VDD.n5679 VDD.n5658 0.0022058
R19424 VDD.n5425 VDD.n5404 0.0022058
R19425 VDD.n3614 VDD.n3593 0.0022058
R19426 VDD.n3872 VDD.n3851 0.0022058
R19427 VDD.n4130 VDD.n4109 0.0022058
R19428 VDD.n4388 VDD.n4367 0.0022058
R19429 VDD.n4646 VDD.n4625 0.0022058
R19430 VDD.n4904 VDD.n4883 0.0022058
R19431 VDD.n5162 VDD.n5141 0.0022058
R19432 VDD.n589 VDD.n587 0.00218421
R19433 VDD.n939 VDD.n937 0.00218421
R19434 VDD.n1745 VDD.n1744 0.00212475
R19435 VDD.n1681 VDD.n1678 0.00212475
R19436 VDD.n1732 VDD.n1712 0.00212475
R19437 VDD.n2094 VDD.n2093 0.00212475
R19438 VDD.n2030 VDD.n2027 0.00212475
R19439 VDD.n2081 VDD.n2061 0.00212475
R19440 VDD.n2324 VDD.n2323 0.00212475
R19441 VDD.n2260 VDD.n2257 0.00212475
R19442 VDD.n2311 VDD.n2291 0.00212475
R19443 VDD.n2582 VDD.n2581 0.00212475
R19444 VDD.n2518 VDD.n2515 0.00212475
R19445 VDD.n2569 VDD.n2549 0.00212475
R19446 VDD.n2840 VDD.n2839 0.00212475
R19447 VDD.n2776 VDD.n2773 0.00212475
R19448 VDD.n2827 VDD.n2807 0.00212475
R19449 VDD.n3098 VDD.n3097 0.00212475
R19450 VDD.n3034 VDD.n3031 0.00212475
R19451 VDD.n3085 VDD.n3065 0.00212475
R19452 VDD.n3356 VDD.n3355 0.00212475
R19453 VDD.n3292 VDD.n3289 0.00212475
R19454 VDD.n3343 VDD.n3323 0.00212475
R19455 VDD.n5679 VDD.n5678 0.00212475
R19456 VDD.n5615 VDD.n5612 0.00212475
R19457 VDD.n5666 VDD.n5646 0.00212475
R19458 VDD.n5425 VDD.n5424 0.00212475
R19459 VDD.n5361 VDD.n5358 0.00212475
R19460 VDD.n5412 VDD.n5392 0.00212475
R19461 VDD.n3614 VDD.n3613 0.00212475
R19462 VDD.n3550 VDD.n3547 0.00212475
R19463 VDD.n3601 VDD.n3581 0.00212475
R19464 VDD.n3872 VDD.n3871 0.00212475
R19465 VDD.n3808 VDD.n3805 0.00212475
R19466 VDD.n3859 VDD.n3839 0.00212475
R19467 VDD.n4130 VDD.n4129 0.00212475
R19468 VDD.n4066 VDD.n4063 0.00212475
R19469 VDD.n4117 VDD.n4097 0.00212475
R19470 VDD.n4388 VDD.n4387 0.00212475
R19471 VDD.n4324 VDD.n4321 0.00212475
R19472 VDD.n4375 VDD.n4355 0.00212475
R19473 VDD.n4646 VDD.n4645 0.00212475
R19474 VDD.n4582 VDD.n4579 0.00212475
R19475 VDD.n4633 VDD.n4613 0.00212475
R19476 VDD.n4904 VDD.n4903 0.00212475
R19477 VDD.n4840 VDD.n4837 0.00212475
R19478 VDD.n4891 VDD.n4871 0.00212475
R19479 VDD.n5162 VDD.n5161 0.00212475
R19480 VDD.n5098 VDD.n5095 0.00212475
R19481 VDD.n5149 VDD.n5129 0.00212475
R19482 VDD VDD.n1599 0.00202016
R19483 VDD.n22 VDD.n3 0.00195349
R19484 VDD.n21 VDD.n4 0.00195349
R19485 VDD.n17 VDD.n16 0.00195349
R19486 VDD.n15 VDD.n14 0.00195349
R19487 VDD.n11 VDD.n10 0.00195349
R19488 VDD.n1166 VDD.n1147 0.00195349
R19489 VDD.n1165 VDD.n1148 0.00195349
R19490 VDD.n1161 VDD.n1160 0.00195349
R19491 VDD.n1159 VDD.n1158 0.00195349
R19492 VDD.n1155 VDD.n1154 0.00195349
R19493 VDD.n284 VDD.n283 0.00194737
R19494 VDD.n281 VDD.n280 0.00194737
R19495 VDD.n1757 VDD.n1756 0.00194704
R19496 VDD.n2106 VDD.n2105 0.00194704
R19497 VDD.n2336 VDD.n2335 0.00194704
R19498 VDD.n2594 VDD.n2593 0.00194704
R19499 VDD.n2852 VDD.n2851 0.00194704
R19500 VDD.n3110 VDD.n3109 0.00194704
R19501 VDD.n3368 VDD.n3367 0.00194704
R19502 VDD.n5691 VDD.n5690 0.00194704
R19503 VDD.n5437 VDD.n5436 0.00194704
R19504 VDD.n3626 VDD.n3625 0.00194704
R19505 VDD.n3884 VDD.n3883 0.00194704
R19506 VDD.n4142 VDD.n4141 0.00194704
R19507 VDD.n4400 VDD.n4399 0.00194704
R19508 VDD.n4658 VDD.n4657 0.00194704
R19509 VDD.n4916 VDD.n4915 0.00194704
R19510 VDD.n5174 VDD.n5173 0.00194704
R19511 VDD.n795 VDD.n794 0.00190323
R19512 VDD.n1735 VDD.n1730 0.00188889
R19513 VDD.n2084 VDD.n2079 0.00188889
R19514 VDD.n2314 VDD.n2309 0.00188889
R19515 VDD.n2572 VDD.n2567 0.00188889
R19516 VDD.n2830 VDD.n2825 0.00188889
R19517 VDD.n3088 VDD.n3083 0.00188889
R19518 VDD.n3346 VDD.n3341 0.00188889
R19519 VDD.n5669 VDD.n5664 0.00188889
R19520 VDD.n5415 VDD.n5410 0.00188889
R19521 VDD.n3604 VDD.n3599 0.00188889
R19522 VDD.n3862 VDD.n3857 0.00188889
R19523 VDD.n4120 VDD.n4115 0.00188889
R19524 VDD.n4378 VDD.n4373 0.00188889
R19525 VDD.n4636 VDD.n4631 0.00188889
R19526 VDD.n4894 VDD.n4889 0.00188889
R19527 VDD.n5152 VDD.n5147 0.00188889
R19528 VDD.n1426 VDD.n1345 0.00182979
R19529 VDD.n1401 VDD.n1399 0.00182979
R19530 VDD.n1369 VDD.n1361 0.00182979
R19531 VDD.n1509 VDD.n1506 0.00182979
R19532 VDD.n1459 VDD.n1289 0.00182979
R19533 VDD.n1599 VDD.n1598 0.00178629
R19534 VDD.n1803 VDD.n1777 0.00175592
R19535 VDD.n1802 VDD.n1777 0.00175592
R19536 VDD.n2011 VDD.n1985 0.00175592
R19537 VDD.n2010 VDD.n1985 0.00175592
R19538 VDD.n2382 VDD.n2356 0.00175592
R19539 VDD.n2381 VDD.n2356 0.00175592
R19540 VDD.n2640 VDD.n2614 0.00175592
R19541 VDD.n2639 VDD.n2614 0.00175592
R19542 VDD.n2898 VDD.n2872 0.00175592
R19543 VDD.n2897 VDD.n2872 0.00175592
R19544 VDD.n3156 VDD.n3130 0.00175592
R19545 VDD.n3155 VDD.n3130 0.00175592
R19546 VDD.n3414 VDD.n3388 0.00175592
R19547 VDD.n3413 VDD.n3388 0.00175592
R19548 VDD.n5737 VDD.n5711 0.00175592
R19549 VDD.n5736 VDD.n5711 0.00175592
R19550 VDD.n5483 VDD.n5457 0.00175592
R19551 VDD.n5482 VDD.n5457 0.00175592
R19552 VDD.n3672 VDD.n3646 0.00175592
R19553 VDD.n3671 VDD.n3646 0.00175592
R19554 VDD.n3930 VDD.n3904 0.00175592
R19555 VDD.n3929 VDD.n3904 0.00175592
R19556 VDD.n4188 VDD.n4162 0.00175592
R19557 VDD.n4187 VDD.n4162 0.00175592
R19558 VDD.n4446 VDD.n4420 0.00175592
R19559 VDD.n4445 VDD.n4420 0.00175592
R19560 VDD.n4704 VDD.n4678 0.00175592
R19561 VDD.n4703 VDD.n4678 0.00175592
R19562 VDD.n4962 VDD.n4936 0.00175592
R19563 VDD.n4961 VDD.n4936 0.00175592
R19564 VDD.n5220 VDD.n5194 0.00175592
R19565 VDD.n5219 VDD.n5194 0.00175592
R19566 VDD.n1838 VDD.n1825 0.00162613
R19567 VDD.n2159 VDD.n2146 0.00162613
R19568 VDD.n2417 VDD.n2404 0.00162613
R19569 VDD.n2675 VDD.n2662 0.00162613
R19570 VDD.n2933 VDD.n2920 0.00162613
R19571 VDD.n3191 VDD.n3178 0.00162613
R19572 VDD.n3449 VDD.n3436 0.00162613
R19573 VDD.n5769 VDD.n5756 0.00162613
R19574 VDD.n5515 VDD.n5502 0.00162613
R19575 VDD.n3707 VDD.n3694 0.00162613
R19576 VDD.n3965 VDD.n3952 0.00162613
R19577 VDD.n4223 VDD.n4210 0.00162613
R19578 VDD.n4481 VDD.n4468 0.00162613
R19579 VDD.n4739 VDD.n4726 0.00162613
R19580 VDD.n4997 VDD.n4984 0.00162613
R19581 VDD.n5255 VDD.n5242 0.00162613
R19582 VDD.n1921 VDD.n1664 0.00162258
R19583 VDD.n2242 VDD.n1983 0.00162258
R19584 VDD.n2500 VDD.n2243 0.00162258
R19585 VDD.n2758 VDD.n2501 0.00162258
R19586 VDD.n3016 VDD.n2759 0.00162258
R19587 VDD.n3274 VDD.n3017 0.00162258
R19588 VDD.n3532 VDD.n3275 0.00162258
R19589 VDD.n3790 VDD.n3533 0.00162258
R19590 VDD.n4048 VDD.n3791 0.00162258
R19591 VDD.n4306 VDD.n4049 0.00162258
R19592 VDD.n4564 VDD.n4307 0.00162258
R19593 VDD.n4822 VDD.n4565 0.00162258
R19594 VDD.n5080 VDD.n4823 0.00162258
R19595 VDD.n5338 VDD.n5081 0.00162258
R19596 VDD.n1815 VDD.n1810 0.00161113
R19597 VDD.n2136 VDD.n2131 0.00161113
R19598 VDD.n2394 VDD.n2389 0.00161113
R19599 VDD.n2652 VDD.n2647 0.00161113
R19600 VDD.n2910 VDD.n2905 0.00161113
R19601 VDD.n3168 VDD.n3163 0.00161113
R19602 VDD.n3426 VDD.n3421 0.00161113
R19603 VDD.n5746 VDD.n5741 0.00161113
R19604 VDD.n5492 VDD.n5487 0.00161113
R19605 VDD.n3684 VDD.n3679 0.00161113
R19606 VDD.n3942 VDD.n3937 0.00161113
R19607 VDD.n4200 VDD.n4195 0.00161113
R19608 VDD.n4458 VDD.n4453 0.00161113
R19609 VDD.n4716 VDD.n4711 0.00161113
R19610 VDD.n4974 VDD.n4969 0.00161113
R19611 VDD.n5232 VDD.n5227 0.00161113
R19612 VDD.n1808 VDD.n1664 0.00160808
R19613 VDD.n2129 VDD.n1983 0.00160808
R19614 VDD.n2387 VDD.n2243 0.00160808
R19615 VDD.n2645 VDD.n2501 0.00160808
R19616 VDD.n2903 VDD.n2759 0.00160808
R19617 VDD.n3161 VDD.n3017 0.00160808
R19618 VDD.n3419 VDD.n3275 0.00160808
R19619 VDD.n3677 VDD.n3533 0.00160808
R19620 VDD.n3935 VDD.n3791 0.00160808
R19621 VDD.n4193 VDD.n4049 0.00160808
R19622 VDD.n4451 VDD.n4307 0.00160808
R19623 VDD.n4709 VDD.n4565 0.00160808
R19624 VDD.n4967 VDD.n4823 0.00160808
R19625 VDD.n5225 VDD.n5081 0.00160808
R19626 VDD.n1949 VDD.n1942 0.00158558
R19627 VDD.n1931 VDD.n1930 0.00158558
R19628 VDD.n1807 VDD.n1775 0.00157581
R19629 VDD.n2127 VDD.n2124 0.00157581
R19630 VDD.n2386 VDD.n2354 0.00157581
R19631 VDD.n2644 VDD.n2612 0.00157581
R19632 VDD.n2902 VDD.n2870 0.00157581
R19633 VDD.n3160 VDD.n3128 0.00157581
R19634 VDD.n3418 VDD.n3386 0.00157581
R19635 VDD.n3676 VDD.n3644 0.00157581
R19636 VDD.n3934 VDD.n3902 0.00157581
R19637 VDD.n4192 VDD.n4160 0.00157581
R19638 VDD.n4450 VDD.n4418 0.00157581
R19639 VDD.n4708 VDD.n4676 0.00157581
R19640 VDD.n4966 VDD.n4934 0.00157581
R19641 VDD.n5224 VDD.n5192 0.00157581
R19642 VDD.n1801 VDD.n1800 0.00151809
R19643 VDD.n2009 VDD.n2008 0.00151809
R19644 VDD.n2380 VDD.n2379 0.00151809
R19645 VDD.n2638 VDD.n2637 0.00151809
R19646 VDD.n2896 VDD.n2895 0.00151809
R19647 VDD.n3154 VDD.n3153 0.00151809
R19648 VDD.n3412 VDD.n3411 0.00151809
R19649 VDD.n5735 VDD.n5734 0.00151809
R19650 VDD.n5481 VDD.n5480 0.00151809
R19651 VDD.n3670 VDD.n3669 0.00151809
R19652 VDD.n3928 VDD.n3927 0.00151809
R19653 VDD.n4186 VDD.n4185 0.00151809
R19654 VDD.n4444 VDD.n4443 0.00151809
R19655 VDD.n4702 VDD.n4701 0.00151809
R19656 VDD.n4960 VDD.n4959 0.00151809
R19657 VDD.n5218 VDD.n5217 0.00151809
R19658 VDD.n1801 VDD.n1777 0.00149567
R19659 VDD.n2009 VDD.n1985 0.00149567
R19660 VDD.n2380 VDD.n2356 0.00149567
R19661 VDD.n2638 VDD.n2614 0.00149567
R19662 VDD.n2896 VDD.n2872 0.00149567
R19663 VDD.n3154 VDD.n3130 0.00149567
R19664 VDD.n3412 VDD.n3388 0.00149567
R19665 VDD.n5735 VDD.n5711 0.00149567
R19666 VDD.n5481 VDD.n5457 0.00149567
R19667 VDD.n3670 VDD.n3646 0.00149567
R19668 VDD.n3928 VDD.n3904 0.00149567
R19669 VDD.n4186 VDD.n4162 0.00149567
R19670 VDD.n4444 VDD.n4420 0.00149567
R19671 VDD.n4702 VDD.n4678 0.00149567
R19672 VDD.n4960 VDD.n4936 0.00149567
R19673 VDD.n5218 VDD.n5194 0.00149567
R19674 VDD.n1917 VDD.n1916 0.00148913
R19675 VDD.n2238 VDD.n2237 0.00148913
R19676 VDD.n2496 VDD.n2495 0.00148913
R19677 VDD.n2754 VDD.n2753 0.00148913
R19678 VDD.n3012 VDD.n3011 0.00148913
R19679 VDD.n3270 VDD.n3269 0.00148913
R19680 VDD.n3528 VDD.n3527 0.00148913
R19681 VDD.n5848 VDD.n5847 0.00148913
R19682 VDD.n5594 VDD.n5593 0.00148913
R19683 VDD.n3786 VDD.n3785 0.00148913
R19684 VDD.n4044 VDD.n4043 0.00148913
R19685 VDD.n4302 VDD.n4301 0.00148913
R19686 VDD.n4560 VDD.n4559 0.00148913
R19687 VDD.n4818 VDD.n4817 0.00148913
R19688 VDD.n5076 VDD.n5075 0.00148913
R19689 VDD.n5334 VDD.n5333 0.00148913
R19690 VDD.n1602 VDD.n1601 0.00147143
R19691 VDD.n1806 VDD.n1805 0.00147065
R19692 VDD.n2126 VDD.n2125 0.00147065
R19693 VDD.n2385 VDD.n2384 0.00147065
R19694 VDD.n2643 VDD.n2642 0.00147065
R19695 VDD.n2901 VDD.n2900 0.00147065
R19696 VDD.n3159 VDD.n3158 0.00147065
R19697 VDD.n3417 VDD.n3416 0.00147065
R19698 VDD.n3675 VDD.n3674 0.00147065
R19699 VDD.n3933 VDD.n3932 0.00147065
R19700 VDD.n4191 VDD.n4190 0.00147065
R19701 VDD.n4449 VDD.n4448 0.00147065
R19702 VDD.n4707 VDD.n4706 0.00147065
R19703 VDD.n4965 VDD.n4964 0.00147065
R19704 VDD.n5223 VDD.n5222 0.00147065
R19705 VDD.n1769 VDD.n1670 0.00145131
R19706 VDD.n1711 VDD.n1670 0.00145131
R19707 VDD.n2118 VDD.n2019 0.00145131
R19708 VDD.n2060 VDD.n2019 0.00145131
R19709 VDD.n2348 VDD.n2249 0.00145131
R19710 VDD.n2290 VDD.n2249 0.00145131
R19711 VDD.n2606 VDD.n2507 0.00145131
R19712 VDD.n2548 VDD.n2507 0.00145131
R19713 VDD.n2864 VDD.n2765 0.00145131
R19714 VDD.n2806 VDD.n2765 0.00145131
R19715 VDD.n3122 VDD.n3023 0.00145131
R19716 VDD.n3064 VDD.n3023 0.00145131
R19717 VDD.n3380 VDD.n3281 0.00145131
R19718 VDD.n3322 VDD.n3281 0.00145131
R19719 VDD.n5703 VDD.n5604 0.00145131
R19720 VDD.n5645 VDD.n5604 0.00145131
R19721 VDD.n5449 VDD.n5350 0.00145131
R19722 VDD.n5391 VDD.n5350 0.00145131
R19723 VDD.n3638 VDD.n3539 0.00145131
R19724 VDD.n3580 VDD.n3539 0.00145131
R19725 VDD.n3896 VDD.n3797 0.00145131
R19726 VDD.n3838 VDD.n3797 0.00145131
R19727 VDD.n4154 VDD.n4055 0.00145131
R19728 VDD.n4096 VDD.n4055 0.00145131
R19729 VDD.n4412 VDD.n4313 0.00145131
R19730 VDD.n4354 VDD.n4313 0.00145131
R19731 VDD.n4670 VDD.n4571 0.00145131
R19732 VDD.n4612 VDD.n4571 0.00145131
R19733 VDD.n4928 VDD.n4829 0.00145131
R19734 VDD.n4870 VDD.n4829 0.00145131
R19735 VDD.n5186 VDD.n5087 0.00145131
R19736 VDD.n5128 VDD.n5087 0.00145131
R19737 VDD.n1770 VDD.n1769 0.00145112
R19738 VDD.n2119 VDD.n2118 0.00145112
R19739 VDD.n2349 VDD.n2348 0.00145112
R19740 VDD.n2607 VDD.n2606 0.00145112
R19741 VDD.n2865 VDD.n2864 0.00145112
R19742 VDD.n3123 VDD.n3122 0.00145112
R19743 VDD.n3381 VDD.n3380 0.00145112
R19744 VDD.n5704 VDD.n5703 0.00145112
R19745 VDD.n5450 VDD.n5449 0.00145112
R19746 VDD.n3639 VDD.n3638 0.00145112
R19747 VDD.n3897 VDD.n3896 0.00145112
R19748 VDD.n4155 VDD.n4154 0.00145112
R19749 VDD.n4413 VDD.n4412 0.00145112
R19750 VDD.n4671 VDD.n4670 0.00145112
R19751 VDD.n4929 VDD.n4928 0.00145112
R19752 VDD.n5187 VDD.n5186 0.00145112
R19753 VDD.n1756 VDD.n1755 0.00144714
R19754 VDD.n2105 VDD.n2104 0.00144714
R19755 VDD.n2335 VDD.n2334 0.00144714
R19756 VDD.n2593 VDD.n2592 0.00144714
R19757 VDD.n2851 VDD.n2850 0.00144714
R19758 VDD.n3109 VDD.n3108 0.00144714
R19759 VDD.n3367 VDD.n3366 0.00144714
R19760 VDD.n5690 VDD.n5689 0.00144714
R19761 VDD.n5436 VDD.n5435 0.00144714
R19762 VDD.n3625 VDD.n3624 0.00144714
R19763 VDD.n3883 VDD.n3882 0.00144714
R19764 VDD.n4141 VDD.n4140 0.00144714
R19765 VDD.n4399 VDD.n4398 0.00144714
R19766 VDD.n4657 VDD.n4656 0.00144714
R19767 VDD.n4915 VDD.n4914 0.00144714
R19768 VDD.n5173 VDD.n5172 0.00144714
R19769 VDD.n1755 VDD.n1754 0.00144695
R19770 VDD.n2104 VDD.n2103 0.00144695
R19771 VDD.n2334 VDD.n2333 0.00144695
R19772 VDD.n2592 VDD.n2591 0.00144695
R19773 VDD.n2850 VDD.n2849 0.00144695
R19774 VDD.n3108 VDD.n3107 0.00144695
R19775 VDD.n3366 VDD.n3365 0.00144695
R19776 VDD.n5689 VDD.n5688 0.00144695
R19777 VDD.n5435 VDD.n5434 0.00144695
R19778 VDD.n3624 VDD.n3623 0.00144695
R19779 VDD.n3882 VDD.n3881 0.00144695
R19780 VDD.n4140 VDD.n4139 0.00144695
R19781 VDD.n4398 VDD.n4397 0.00144695
R19782 VDD.n4656 VDD.n4655 0.00144695
R19783 VDD.n4914 VDD.n4913 0.00144695
R19784 VDD.n5172 VDD.n5171 0.00144695
R19785 VDD.n798 VDD.n797 0.00143548
R19786 VDD.n686 VDD.n685 0.00142105
R19787 VDD.n1036 VDD.n1035 0.00142105
R19788 VDD.n1978 VDD.n1924 0.00139286
R19789 VDD.n1719 VDD.n1668 0.00139286
R19790 VDD.n2068 VDD.n2017 0.00139286
R19791 VDD.n2298 VDD.n2247 0.00139286
R19792 VDD.n2556 VDD.n2505 0.00139286
R19793 VDD.n2814 VDD.n2763 0.00139286
R19794 VDD.n3072 VDD.n3021 0.00139286
R19795 VDD.n3330 VDD.n3279 0.00139286
R19796 VDD.n5653 VDD.n5602 0.00139286
R19797 VDD.n5399 VDD.n5348 0.00139286
R19798 VDD.n3588 VDD.n3537 0.00139286
R19799 VDD.n3846 VDD.n3795 0.00139286
R19800 VDD.n4104 VDD.n4053 0.00139286
R19801 VDD.n4362 VDD.n4311 0.00139286
R19802 VDD.n4620 VDD.n4569 0.00139286
R19803 VDD.n4878 VDD.n4827 0.00139286
R19804 VDD.n5136 VDD.n5085 0.00139286
R19805 VDD.t1036 VDD.n1941 0.00134143
R19806 VDD.n1885 VDD.n1819 0.00133663
R19807 VDD.n1821 VDD.n1819 0.00133663
R19808 VDD.n2206 VDD.n2140 0.00133663
R19809 VDD.n2142 VDD.n2140 0.00133663
R19810 VDD.n2464 VDD.n2398 0.00133663
R19811 VDD.n2400 VDD.n2398 0.00133663
R19812 VDD.n2722 VDD.n2656 0.00133663
R19813 VDD.n2658 VDD.n2656 0.00133663
R19814 VDD.n2980 VDD.n2914 0.00133663
R19815 VDD.n2916 VDD.n2914 0.00133663
R19816 VDD.n3238 VDD.n3172 0.00133663
R19817 VDD.n3174 VDD.n3172 0.00133663
R19818 VDD.n3496 VDD.n3430 0.00133663
R19819 VDD.n3432 VDD.n3430 0.00133663
R19820 VDD.n5816 VDD.n5750 0.00133663
R19821 VDD.n5752 VDD.n5750 0.00133663
R19822 VDD.n5562 VDD.n5496 0.00133663
R19823 VDD.n5498 VDD.n5496 0.00133663
R19824 VDD.n3754 VDD.n3688 0.00133663
R19825 VDD.n3690 VDD.n3688 0.00133663
R19826 VDD.n4012 VDD.n3946 0.00133663
R19827 VDD.n3948 VDD.n3946 0.00133663
R19828 VDD.n4270 VDD.n4204 0.00133663
R19829 VDD.n4206 VDD.n4204 0.00133663
R19830 VDD.n4528 VDD.n4462 0.00133663
R19831 VDD.n4464 VDD.n4462 0.00133663
R19832 VDD.n4786 VDD.n4720 0.00133663
R19833 VDD.n4722 VDD.n4720 0.00133663
R19834 VDD.n5044 VDD.n4978 0.00133663
R19835 VDD.n4980 VDD.n4978 0.00133663
R19836 VDD.n5302 VDD.n5236 0.00133663
R19837 VDD.n5238 VDD.n5236 0.00133663
R19838 VDD.n1981 VDD 0.00130357
R19839 VDD.n283 VDD 0.00128947
R19840 VDD.n1805 VDD.n1775 0.00120516
R19841 VDD.n2125 VDD.n2124 0.00120516
R19842 VDD.n2384 VDD.n2354 0.00120516
R19843 VDD.n2642 VDD.n2612 0.00120516
R19844 VDD.n2900 VDD.n2870 0.00120516
R19845 VDD.n3158 VDD.n3128 0.00120516
R19846 VDD.n3416 VDD.n3386 0.00120516
R19847 VDD.n3674 VDD.n3644 0.00120516
R19848 VDD.n3932 VDD.n3902 0.00120516
R19849 VDD.n4190 VDD.n4160 0.00120516
R19850 VDD.n4448 VDD.n4418 0.00120516
R19851 VDD.n4706 VDD.n4676 0.00120516
R19852 VDD.n4964 VDD.n4934 0.00120516
R19853 VDD.n5222 VDD.n5192 0.00120516
R19854 VDD.n855 VDD.n821 0.00116652
R19855 VDD.n1238 VDD.n1204 0.00116652
R19856 VDD.n859 VDD.n858 0.00114708
R19857 VDD.n858 VDD.n856 0.00114708
R19858 VDD.n1242 VDD.n1241 0.00114708
R19859 VDD.n1241 VDD.n1239 0.00114708
R19860 VDD.n1871 VDD.n1844 0.00114565
R19861 VDD.n1847 VDD.n1844 0.00114565
R19862 VDD.n2192 VDD.n2165 0.00114565
R19863 VDD.n2168 VDD.n2165 0.00114565
R19864 VDD.n2450 VDD.n2423 0.00114565
R19865 VDD.n2426 VDD.n2423 0.00114565
R19866 VDD.n2708 VDD.n2681 0.00114565
R19867 VDD.n2684 VDD.n2681 0.00114565
R19868 VDD.n2966 VDD.n2939 0.00114565
R19869 VDD.n2942 VDD.n2939 0.00114565
R19870 VDD.n3224 VDD.n3197 0.00114565
R19871 VDD.n3200 VDD.n3197 0.00114565
R19872 VDD.n3482 VDD.n3455 0.00114565
R19873 VDD.n3458 VDD.n3455 0.00114565
R19874 VDD.n5802 VDD.n5775 0.00114565
R19875 VDD.n5778 VDD.n5775 0.00114565
R19876 VDD.n5548 VDD.n5521 0.00114565
R19877 VDD.n5524 VDD.n5521 0.00114565
R19878 VDD.n3740 VDD.n3713 0.00114565
R19879 VDD.n3716 VDD.n3713 0.00114565
R19880 VDD.n3998 VDD.n3971 0.00114565
R19881 VDD.n3974 VDD.n3971 0.00114565
R19882 VDD.n4256 VDD.n4229 0.00114565
R19883 VDD.n4232 VDD.n4229 0.00114565
R19884 VDD.n4514 VDD.n4487 0.00114565
R19885 VDD.n4490 VDD.n4487 0.00114565
R19886 VDD.n4772 VDD.n4745 0.00114565
R19887 VDD.n4748 VDD.n4745 0.00114565
R19888 VDD.n5030 VDD.n5003 0.00114565
R19889 VDD.n5006 VDD.n5003 0.00114565
R19890 VDD.n5288 VDD.n5261 0.00114565
R19891 VDD.n5264 VDD.n5261 0.00114565
R19892 VDD.n1739 VDD.n1738 0.00113805
R19893 VDD.n2088 VDD.n2087 0.00113805
R19894 VDD.n2318 VDD.n2317 0.00113805
R19895 VDD.n2576 VDD.n2575 0.00113805
R19896 VDD.n2834 VDD.n2833 0.00113805
R19897 VDD.n3092 VDD.n3091 0.00113805
R19898 VDD.n3350 VDD.n3349 0.00113805
R19899 VDD.n5673 VDD.n5672 0.00113805
R19900 VDD.n5419 VDD.n5418 0.00113805
R19901 VDD.n3608 VDD.n3607 0.00113805
R19902 VDD.n3866 VDD.n3865 0.00113805
R19903 VDD.n4124 VDD.n4123 0.00113805
R19904 VDD.n4382 VDD.n4381 0.00113805
R19905 VDD.n4640 VDD.n4639 0.00113805
R19906 VDD.n4898 VDD.n4897 0.00113805
R19907 VDD.n5156 VDD.n5155 0.00113805
R19908 VDD.n1621 VDD.n1620 0.00111657
R19909 VDD.n1976 VDD.n1975 0.00111635
R19910 VDD.t1038 VDD.n1969 0.0010973
R19911 VDD.n1798 VDD.n1797 0.00108642
R19912 VDD.n2006 VDD.n2005 0.00108642
R19913 VDD.n2377 VDD.n2376 0.00108642
R19914 VDD.n2635 VDD.n2634 0.00108642
R19915 VDD.n2893 VDD.n2892 0.00108642
R19916 VDD.n3151 VDD.n3150 0.00108642
R19917 VDD.n3409 VDD.n3408 0.00108642
R19918 VDD.n5732 VDD.n5731 0.00108642
R19919 VDD.n5478 VDD.n5477 0.00108642
R19920 VDD.n3667 VDD.n3666 0.00108642
R19921 VDD.n3925 VDD.n3924 0.00108642
R19922 VDD.n4183 VDD.n4182 0.00108642
R19923 VDD.n4441 VDD.n4440 0.00108642
R19924 VDD.n4699 VDD.n4698 0.00108642
R19925 VDD.n4957 VDD.n4956 0.00108642
R19926 VDD.n5215 VDD.n5214 0.00108642
R19927 VDD.n860 VDD.n859 0.00107711
R19928 VDD.n1243 VDD.n1242 0.00107711
R19929 VDD.n1642 VDD.n1641 0.00107006
R19930 VDD.n1613 VDD.n1612 0.00106596
R19931 VDD.n1752 VDD.n1720 0.00105202
R19932 VDD.n2101 VDD.n2069 0.00105202
R19933 VDD.n2331 VDD.n2299 0.00105202
R19934 VDD.n2589 VDD.n2557 0.00105202
R19935 VDD.n2847 VDD.n2815 0.00105202
R19936 VDD.n3105 VDD.n3073 0.00105202
R19937 VDD.n3363 VDD.n3331 0.00105202
R19938 VDD.n5686 VDD.n5654 0.00105202
R19939 VDD.n5432 VDD.n5400 0.00105202
R19940 VDD.n3621 VDD.n3589 0.00105202
R19941 VDD.n3879 VDD.n3847 0.00105202
R19942 VDD.n4137 VDD.n4105 0.00105202
R19943 VDD.n4395 VDD.n4363 0.00105202
R19944 VDD.n4653 VDD.n4621 0.00105202
R19945 VDD.n4911 VDD.n4879 0.00105202
R19946 VDD.n5169 VDD.n5137 0.00105202
R19947 VDD.n1431 VDD.n1430 0.00100344
R19948 VDD.n1455 VDD.n1454 0.00100344
R19949 VDD.n1374 VDD.n1373 0.00100342
R19950 VDD.n1711 VDD.n1710 0.00100293
R19951 VDD.n2060 VDD.n2059 0.00100293
R19952 VDD.n2290 VDD.n2289 0.00100293
R19953 VDD.n2548 VDD.n2547 0.00100293
R19954 VDD.n2806 VDD.n2805 0.00100293
R19955 VDD.n3064 VDD.n3063 0.00100293
R19956 VDD.n3322 VDD.n3321 0.00100293
R19957 VDD.n5645 VDD.n5644 0.00100293
R19958 VDD.n5391 VDD.n5390 0.00100293
R19959 VDD.n3580 VDD.n3579 0.00100293
R19960 VDD.n3838 VDD.n3837 0.00100293
R19961 VDD.n4096 VDD.n4095 0.00100293
R19962 VDD.n4354 VDD.n4353 0.00100293
R19963 VDD.n4612 VDD.n4611 0.00100293
R19964 VDD.n4870 VDD.n4869 0.00100293
R19965 VDD.n5128 VDD.n5127 0.00100293
R19966 VDD.n464 VDD.n463 0.00100258
R19967 VDD.n61 VDD.n60 0.00100258
R19968 VDD.n1837 VDD.n1826 0.00100132
R19969 VDD.n2158 VDD.n2147 0.00100132
R19970 VDD.n2416 VDD.n2405 0.00100132
R19971 VDD.n2674 VDD.n2663 0.00100132
R19972 VDD.n2932 VDD.n2921 0.00100132
R19973 VDD.n3190 VDD.n3179 0.00100132
R19974 VDD.n3448 VDD.n3437 0.00100132
R19975 VDD.n5768 VDD.n5757 0.00100132
R19976 VDD.n5514 VDD.n5503 0.00100132
R19977 VDD.n3706 VDD.n3695 0.00100132
R19978 VDD.n3964 VDD.n3953 0.00100132
R19979 VDD.n4222 VDD.n4211 0.00100132
R19980 VDD.n4480 VDD.n4469 0.00100132
R19981 VDD.n4738 VDD.n4727 0.00100132
R19982 VDD.n4996 VDD.n4985 0.00100132
R19983 VDD.n5254 VDD.n5243 0.00100132
R19984 VDD.n587 VDD.n586 0.00100097
R19985 VDD.n937 VDD.n936 0.00100097
R19986 VDD.n186 VDD.n185 0.00100097
R19987 VDD.n1547 VDD.n1541 0.00100097
R19988 VDD.n1620 VDD.n1614 0.00100057
R19989 VDD.n1798 VDD.n1777 0.00100033
R19990 VDD.n2006 VDD.n1985 0.00100033
R19991 VDD.n2377 VDD.n2356 0.00100033
R19992 VDD.n2635 VDD.n2614 0.00100033
R19993 VDD.n2893 VDD.n2872 0.00100033
R19994 VDD.n3151 VDD.n3130 0.00100033
R19995 VDD.n3409 VDD.n3388 0.00100033
R19996 VDD.n5732 VDD.n5711 0.00100033
R19997 VDD.n5478 VDD.n5457 0.00100033
R19998 VDD.n3667 VDD.n3646 0.00100033
R19999 VDD.n3925 VDD.n3904 0.00100033
R20000 VDD.n4183 VDD.n4162 0.00100033
R20001 VDD.n4441 VDD.n4420 0.00100033
R20002 VDD.n4699 VDD.n4678 0.00100033
R20003 VDD.n4957 VDD.n4936 0.00100033
R20004 VDD.n5215 VDD.n5194 0.00100033
R20005 VDD.n1882 VDD.n1821 0.00100021
R20006 VDD.n2203 VDD.n2142 0.00100021
R20007 VDD.n2461 VDD.n2400 0.00100021
R20008 VDD.n2719 VDD.n2658 0.00100021
R20009 VDD.n2977 VDD.n2916 0.00100021
R20010 VDD.n3235 VDD.n3174 0.00100021
R20011 VDD.n3493 VDD.n3432 0.00100021
R20012 VDD.n5813 VDD.n5752 0.00100021
R20013 VDD.n5559 VDD.n5498 0.00100021
R20014 VDD.n3751 VDD.n3690 0.00100021
R20015 VDD.n4009 VDD.n3948 0.00100021
R20016 VDD.n4267 VDD.n4206 0.00100021
R20017 VDD.n4525 VDD.n4464 0.00100021
R20018 VDD.n4783 VDD.n4722 0.00100021
R20019 VDD.n5041 VDD.n4980 0.00100021
R20020 VDD.n5299 VDD.n5238 0.00100021
R20021 VDD.n860 VDD.n855 0.00100013
R20022 VDD.n1243 VDD.n1238 0.00100013
R20023 VDD.n1757 VDD.n1711 0.0010001
R20024 VDD.n2106 VDD.n2060 0.0010001
R20025 VDD.n2336 VDD.n2290 0.0010001
R20026 VDD.n2594 VDD.n2548 0.0010001
R20027 VDD.n2852 VDD.n2806 0.0010001
R20028 VDD.n3110 VDD.n3064 0.0010001
R20029 VDD.n3368 VDD.n3322 0.0010001
R20030 VDD.n5691 VDD.n5645 0.0010001
R20031 VDD.n5437 VDD.n5391 0.0010001
R20032 VDD.n3626 VDD.n3580 0.0010001
R20033 VDD.n3884 VDD.n3838 0.0010001
R20034 VDD.n4142 VDD.n4096 0.0010001
R20035 VDD.n4400 VDD.n4354 0.0010001
R20036 VDD.n4658 VDD.n4612 0.0010001
R20037 VDD.n4916 VDD.n4870 0.0010001
R20038 VDD.n5174 VDD.n5128 0.0010001
R20039 VDD.n1641 VDD.n1640 0.00100008
R20040 VDD.n1952 VDD.n1944 0.00100003
R20041 VDD.n1934 VDD.n1927 0.00100003
R20042 VDD.n1920 VDD.n1808 0.00100002
R20043 VDD.n2241 VDD.n2129 0.00100002
R20044 VDD.n2499 VDD.n2387 0.00100002
R20045 VDD.n2757 VDD.n2645 0.00100002
R20046 VDD.n3015 VDD.n2903 0.00100002
R20047 VDD.n3273 VDD.n3161 0.00100002
R20048 VDD.n3531 VDD.n3419 0.00100002
R20049 VDD.n3789 VDD.n3677 0.00100002
R20050 VDD.n4047 VDD.n3935 0.00100002
R20051 VDD.n4305 VDD.n4193 0.00100002
R20052 VDD.n4563 VDD.n4451 0.00100002
R20053 VDD.n4821 VDD.n4709 0.00100002
R20054 VDD.n5079 VDD.n4967 0.00100002
R20055 VDD.n5337 VDD.n5225 0.00100002
R20056 VDD.n1317 VDD.n1315 0.001
R20057 VDD.n1975 VDD.n1927 0.001
R20058 VDD.n1979 VDD.n1923 0.001
R20059 VDD.n858 VDD.n857 0.001
R20060 VDD.n1241 VDD.n1240 0.001
R20061 VDD.n390 VDD.n389 0.000894737
R20062 VDD.n1640 VDD.n1638 0.000834423
R20063 VDD.n1460 VDD.n1459 0.000765957
R20064 VDD.n688 VDD 0.000763158
R20065 VDD.n1038 VDD 0.000763158
R20066 VDD.n793 VDD.n515 0.000631579
R20067 VDD.n1143 VDD.n865 0.000631579
R20068 VDD.n1621 VDD.n1615 0.000625544
R20069 VDD.n1619 VDD.n1615 0.000625542
R20070 VDD.n1977 VDD.n1976 0.00061635
R20071 VDD.n1978 VDD.n1977 0.000616347
R20072 VDD.n1736 VDD.n1729 0.000594432
R20073 VDD.n2085 VDD.n2078 0.000594432
R20074 VDD.n2315 VDD.n2308 0.000594432
R20075 VDD.n2573 VDD.n2566 0.000594432
R20076 VDD.n2831 VDD.n2824 0.000594432
R20077 VDD.n3089 VDD.n3082 0.000594432
R20078 VDD.n3347 VDD.n3340 0.000594432
R20079 VDD.n5670 VDD.n5663 0.000594432
R20080 VDD.n5416 VDD.n5409 0.000594432
R20081 VDD.n3605 VDD.n3598 0.000594432
R20082 VDD.n3863 VDD.n3856 0.000594432
R20083 VDD.n4121 VDD.n4114 0.000594432
R20084 VDD.n4379 VDD.n4372 0.000594432
R20085 VDD.n4637 VDD.n4630 0.000594432
R20086 VDD.n4895 VDD.n4888 0.000594432
R20087 VDD.n5153 VDD.n5146 0.000594432
R20088 VDD.n1773 VDD.n1772 0.000558569
R20089 VDD.n2122 VDD.n2121 0.000558569
R20090 VDD.n2352 VDD.n2351 0.000558569
R20091 VDD.n2610 VDD.n2609 0.000558569
R20092 VDD.n2868 VDD.n2867 0.000558569
R20093 VDD.n3126 VDD.n3125 0.000558569
R20094 VDD.n3384 VDD.n3383 0.000558569
R20095 VDD.n5707 VDD.n5706 0.000558569
R20096 VDD.n5453 VDD.n5452 0.000558569
R20097 VDD.n3642 VDD.n3641 0.000558569
R20098 VDD.n3900 VDD.n3899 0.000558569
R20099 VDD.n4158 VDD.n4157 0.000558569
R20100 VDD.n4416 VDD.n4415 0.000558569
R20101 VDD.n4674 VDD.n4673 0.000558569
R20102 VDD.n4932 VDD.n4931 0.000558569
R20103 VDD.n5190 VDD.n5189 0.000558569
R20104 VDD.n1740 VDD.n1739 0.000555817
R20105 VDD.n2089 VDD.n2088 0.000555817
R20106 VDD.n2319 VDD.n2318 0.000555817
R20107 VDD.n2577 VDD.n2576 0.000555817
R20108 VDD.n2835 VDD.n2834 0.000555817
R20109 VDD.n3093 VDD.n3092 0.000555817
R20110 VDD.n3351 VDD.n3350 0.000555817
R20111 VDD.n5674 VDD.n5673 0.000555817
R20112 VDD.n5420 VDD.n5419 0.000555817
R20113 VDD.n3609 VDD.n3608 0.000555817
R20114 VDD.n3867 VDD.n3866 0.000555817
R20115 VDD.n4125 VDD.n4124 0.000555817
R20116 VDD.n4383 VDD.n4382 0.000555817
R20117 VDD.n4641 VDD.n4640 0.000555817
R20118 VDD.n4899 VDD.n4898 0.000555817
R20119 VDD.n5157 VDD.n5156 0.000555817
R20120 VDD.n1768 VDD.n1668 0.000534058
R20121 VDD.n2117 VDD.n2017 0.000534058
R20122 VDD.n2347 VDD.n2247 0.000534058
R20123 VDD.n2605 VDD.n2505 0.000534058
R20124 VDD.n2863 VDD.n2763 0.000534058
R20125 VDD.n3121 VDD.n3021 0.000534058
R20126 VDD.n3379 VDD.n3279 0.000534058
R20127 VDD.n5702 VDD.n5602 0.000534058
R20128 VDD.n5448 VDD.n5348 0.000534058
R20129 VDD.n3637 VDD.n3537 0.000534058
R20130 VDD.n3895 VDD.n3795 0.000534058
R20131 VDD.n4153 VDD.n4053 0.000534058
R20132 VDD.n4411 VDD.n4311 0.000534058
R20133 VDD.n4669 VDD.n4569 0.000534058
R20134 VDD.n4927 VDD.n4827 0.000534058
R20135 VDD.n5185 VDD.n5085 0.000534058
R20136 VDD.n1886 VDD.n1885 0.000523376
R20137 VDD.n2207 VDD.n2206 0.000523376
R20138 VDD.n2465 VDD.n2464 0.000523376
R20139 VDD.n2723 VDD.n2722 0.000523376
R20140 VDD.n2981 VDD.n2980 0.000523376
R20141 VDD.n3239 VDD.n3238 0.000523376
R20142 VDD.n3497 VDD.n3496 0.000523376
R20143 VDD.n5817 VDD.n5816 0.000523376
R20144 VDD.n5563 VDD.n5562 0.000523376
R20145 VDD.n3755 VDD.n3754 0.000523376
R20146 VDD.n4013 VDD.n4012 0.000523376
R20147 VDD.n4271 VDD.n4270 0.000523376
R20148 VDD.n4529 VDD.n4528 0.000523376
R20149 VDD.n4787 VDD.n4786 0.000523376
R20150 VDD.n5045 VDD.n5044 0.000523376
R20151 VDD.n5303 VDD.n5302 0.000523376
R20152 VDD.n1704 VDD.n1703 0.000516232
R20153 VDD.n1691 VDD.n1685 0.000516232
R20154 VDD.n2053 VDD.n2052 0.000516232
R20155 VDD.n2040 VDD.n2034 0.000516232
R20156 VDD.n2283 VDD.n2282 0.000516232
R20157 VDD.n2270 VDD.n2264 0.000516232
R20158 VDD.n2541 VDD.n2540 0.000516232
R20159 VDD.n2528 VDD.n2522 0.000516232
R20160 VDD.n2799 VDD.n2798 0.000516232
R20161 VDD.n2786 VDD.n2780 0.000516232
R20162 VDD.n3057 VDD.n3056 0.000516232
R20163 VDD.n3044 VDD.n3038 0.000516232
R20164 VDD.n3315 VDD.n3314 0.000516232
R20165 VDD.n3302 VDD.n3296 0.000516232
R20166 VDD.n5638 VDD.n5637 0.000516232
R20167 VDD.n5625 VDD.n5619 0.000516232
R20168 VDD.n5384 VDD.n5383 0.000516232
R20169 VDD.n5371 VDD.n5365 0.000516232
R20170 VDD.n3573 VDD.n3572 0.000516232
R20171 VDD.n3560 VDD.n3554 0.000516232
R20172 VDD.n3831 VDD.n3830 0.000516232
R20173 VDD.n3818 VDD.n3812 0.000516232
R20174 VDD.n4089 VDD.n4088 0.000516232
R20175 VDD.n4076 VDD.n4070 0.000516232
R20176 VDD.n4347 VDD.n4346 0.000516232
R20177 VDD.n4334 VDD.n4328 0.000516232
R20178 VDD.n4605 VDD.n4604 0.000516232
R20179 VDD.n4592 VDD.n4586 0.000516232
R20180 VDD.n4863 VDD.n4862 0.000516232
R20181 VDD.n4850 VDD.n4844 0.000516232
R20182 VDD.n5121 VDD.n5120 0.000516232
R20183 VDD.n5108 VDD.n5102 0.000516232
R20184 VDD.n1735 VDD.n1734 0.000515622
R20185 VDD.n2084 VDD.n2083 0.000515622
R20186 VDD.n2314 VDD.n2313 0.000515622
R20187 VDD.n2572 VDD.n2571 0.000515622
R20188 VDD.n2830 VDD.n2829 0.000515622
R20189 VDD.n3088 VDD.n3087 0.000515622
R20190 VDD.n3346 VDD.n3345 0.000515622
R20191 VDD.n5669 VDD.n5668 0.000515622
R20192 VDD.n5415 VDD.n5414 0.000515622
R20193 VDD.n3604 VDD.n3603 0.000515622
R20194 VDD.n3862 VDD.n3861 0.000515622
R20195 VDD.n4120 VDD.n4119 0.000515622
R20196 VDD.n4378 VDD.n4377 0.000515622
R20197 VDD.n4636 VDD.n4635 0.000515622
R20198 VDD.n4894 VDD.n4893 0.000515622
R20199 VDD.n5152 VDD.n5151 0.000515622
R20200 VDD.n1876 VDD.n1875 0.000514451
R20201 VDD.n2197 VDD.n2196 0.000514451
R20202 VDD.n2455 VDD.n2454 0.000514451
R20203 VDD.n2713 VDD.n2712 0.000514451
R20204 VDD.n2971 VDD.n2970 0.000514451
R20205 VDD.n3229 VDD.n3228 0.000514451
R20206 VDD.n3487 VDD.n3486 0.000514451
R20207 VDD.n5807 VDD.n5806 0.000514451
R20208 VDD.n5553 VDD.n5552 0.000514451
R20209 VDD.n3745 VDD.n3744 0.000514451
R20210 VDD.n4003 VDD.n4002 0.000514451
R20211 VDD.n4261 VDD.n4260 0.000514451
R20212 VDD.n4519 VDD.n4518 0.000514451
R20213 VDD.n4777 VDD.n4776 0.000514451
R20214 VDD.n5035 VDD.n5034 0.000514451
R20215 VDD.n5293 VDD.n5292 0.000514451
R20216 VDD.n669 VDD.n521 0.000506553
R20217 VDD.n668 VDD.n518 0.000506553
R20218 VDD.n667 VDD.n666 0.000506553
R20219 VDD.n586 VDD.n585 0.000506553
R20220 VDD.n584 VDD.n583 0.000506553
R20221 VDD.n687 VDD.n670 0.000506553
R20222 VDD.n1019 VDD.n871 0.000506553
R20223 VDD.n1018 VDD.n868 0.000506553
R20224 VDD.n1017 VDD.n1016 0.000506553
R20225 VDD.n936 VDD.n935 0.000506553
R20226 VDD.n934 VDD.n933 0.000506553
R20227 VDD.n1037 VDD.n1020 0.000506553
R20228 VDD.n264 VDD.n120 0.000506553
R20229 VDD.n263 VDD.n117 0.000506553
R20230 VDD.n262 VDD.n261 0.000506553
R20231 VDD.n185 VDD.n184 0.000506553
R20232 VDD.n183 VDD.n182 0.000506553
R20233 VDD.n282 VDD.n265 0.000506553
R20234 VDD.n1458 VDD.n1457 0.000506553
R20235 VDD.n1508 VDD.n1507 0.000506553
R20236 VDD.n1456 VDD.n1455 0.000506553
R20237 VDD.n1430 VDD.n1429 0.000506553
R20238 VDD.n1398 VDD.n1397 0.000506553
R20239 VDD.n1373 VDD.n1372 0.000506553
R20240 VDD.n1371 VDD.n1370 0.000506553
R20241 VDD.n1428 VDD.n1427 0.000506553
R20242 VDD.n1726 VDD.n1725 0.000505865
R20243 VDD.n2075 VDD.n2074 0.000505865
R20244 VDD.n2305 VDD.n2304 0.000505865
R20245 VDD.n2563 VDD.n2562 0.000505865
R20246 VDD.n2821 VDD.n2820 0.000505865
R20247 VDD.n3079 VDD.n3078 0.000505865
R20248 VDD.n3337 VDD.n3336 0.000505865
R20249 VDD.n5660 VDD.n5659 0.000505865
R20250 VDD.n5406 VDD.n5405 0.000505865
R20251 VDD.n3595 VDD.n3594 0.000505865
R20252 VDD.n3853 VDD.n3852 0.000505865
R20253 VDD.n4111 VDD.n4110 0.000505865
R20254 VDD.n4369 VDD.n4368 0.000505865
R20255 VDD.n4627 VDD.n4626 0.000505865
R20256 VDD.n4885 VDD.n4884 0.000505865
R20257 VDD.n5143 VDD.n5142 0.000505865
R20258 VDD.n1839 VDD.n1838 0.000504381
R20259 VDD.n2160 VDD.n2159 0.000504381
R20260 VDD.n2418 VDD.n2417 0.000504381
R20261 VDD.n2676 VDD.n2675 0.000504381
R20262 VDD.n2934 VDD.n2933 0.000504381
R20263 VDD.n3192 VDD.n3191 0.000504381
R20264 VDD.n3450 VDD.n3449 0.000504381
R20265 VDD.n5770 VDD.n5769 0.000504381
R20266 VDD.n5516 VDD.n5515 0.000504381
R20267 VDD.n3708 VDD.n3707 0.000504381
R20268 VDD.n3966 VDD.n3965 0.000504381
R20269 VDD.n4224 VDD.n4223 0.000504381
R20270 VDD.n4482 VDD.n4481 0.000504381
R20271 VDD.n4740 VDD.n4739 0.000504381
R20272 VDD.n4998 VDD.n4997 0.000504381
R20273 VDD.n5256 VDD.n5255 0.000504381
R20274 VDD.n1719 VDD.n1671 0.000503792
R20275 VDD.n2068 VDD.n2020 0.000503792
R20276 VDD.n2298 VDD.n2250 0.000503792
R20277 VDD.n2556 VDD.n2508 0.000503792
R20278 VDD.n2814 VDD.n2766 0.000503792
R20279 VDD.n3072 VDD.n3024 0.000503792
R20280 VDD.n3330 VDD.n3282 0.000503792
R20281 VDD.n5653 VDD.n5605 0.000503792
R20282 VDD.n5399 VDD.n5351 0.000503792
R20283 VDD.n3588 VDD.n3540 0.000503792
R20284 VDD.n3846 VDD.n3798 0.000503792
R20285 VDD.n4104 VDD.n4056 0.000503792
R20286 VDD.n4362 VDD.n4314 0.000503792
R20287 VDD.n4620 VDD.n4572 0.000503792
R20288 VDD.n4878 VDD.n4830 0.000503792
R20289 VDD.n5136 VDD.n5088 0.000503792
R20290 VDD.n1427 VDD.n1426 0.000503441
R20291 VDD.n1399 VDD.n1398 0.000503441
R20292 VDD.n1370 VDD.n1369 0.000503441
R20293 VDD.n1459 VDD.n1458 0.000503441
R20294 VDD.n1509 VDD.n1508 0.000503441
R20295 VDD.n1345 VDD.n1344 0.000501258
R20296 VDD.n1319 VDD.n1318 0.000501258
R20297 VDD.n1401 VDD.n1400 0.000501258
R20298 VDD.n1361 VDD.n1360 0.000501258
R20299 VDD.n1289 VDD.n1288 0.000501258
R20300 VDD.n1506 VDD.n1505 0.000501258
R20301 VDD.n1818 VDD.n1817 0.000501164
R20302 VDD.n2139 VDD.n2138 0.000501164
R20303 VDD.n2397 VDD.n2396 0.000501164
R20304 VDD.n2655 VDD.n2654 0.000501164
R20305 VDD.n2913 VDD.n2912 0.000501164
R20306 VDD.n3171 VDD.n3170 0.000501164
R20307 VDD.n3429 VDD.n3428 0.000501164
R20308 VDD.n5749 VDD.n5748 0.000501164
R20309 VDD.n5495 VDD.n5494 0.000501164
R20310 VDD.n3687 VDD.n3686 0.000501164
R20311 VDD.n3945 VDD.n3944 0.000501164
R20312 VDD.n4203 VDD.n4202 0.000501164
R20313 VDD.n4461 VDD.n4460 0.000501164
R20314 VDD.n4719 VDD.n4718 0.000501164
R20315 VDD.n4977 VDD.n4976 0.000501164
R20316 VDD.n5235 VDD.n5234 0.000501164
R20317 VDD.n736 VDD.n521 0.00050097
R20318 VDD.n781 VDD.n518 0.00050097
R20319 VDD.n666 VDD.n665 0.00050097
R20320 VDD.n583 VDD.n582 0.00050097
R20321 VDD.n1086 VDD.n871 0.00050097
R20322 VDD.n1131 VDD.n868 0.00050097
R20323 VDD.n1016 VDD.n1015 0.00050097
R20324 VDD.n933 VDD.n932 0.00050097
R20325 VDD.n331 VDD.n120 0.00050097
R20326 VDD.n376 VDD.n117 0.00050097
R20327 VDD.n261 VDD.n260 0.00050097
R20328 VDD.n182 VDD.n181 0.00050097
R20329 VDD.n687 VDD.n686 0.00050097
R20330 VDD.n1037 VDD.n1036 0.00050097
R20331 VDD.n282 VDD.n281 0.00050097
R20332 VDD.n2193 VDD.n2192 0.000500414
R20333 VDD.n2451 VDD.n2450 0.000500414
R20334 VDD.n2709 VDD.n2708 0.000500414
R20335 VDD.n2967 VDD.n2966 0.000500414
R20336 VDD.n3225 VDD.n3224 0.000500414
R20337 VDD.n3483 VDD.n3482 0.000500414
R20338 VDD.n5803 VDD.n5802 0.000500414
R20339 VDD.n5549 VDD.n5548 0.000500414
R20340 VDD.n3741 VDD.n3740 0.000500414
R20341 VDD.n3999 VDD.n3998 0.000500414
R20342 VDD.n4257 VDD.n4256 0.000500414
R20343 VDD.n4515 VDD.n4514 0.000500414
R20344 VDD.n4773 VDD.n4772 0.000500414
R20345 VDD.n5031 VDD.n5030 0.000500414
R20346 VDD.n5289 VDD.n5288 0.000500414
R20347 VDD.n1872 VDD.n1871 0.000500414
R20348 VDD.n863 VDD.n862 0.000500259
R20349 VDD.n1920 VDD.n1919 0.000500184
R20350 VDD.n2241 VDD.n2240 0.000500184
R20351 VDD.n2499 VDD.n2498 0.000500184
R20352 VDD.n2757 VDD.n2756 0.000500184
R20353 VDD.n3015 VDD.n3014 0.000500184
R20354 VDD.n3273 VDD.n3272 0.000500184
R20355 VDD.n3531 VDD.n3530 0.000500184
R20356 VDD.n3789 VDD.n3788 0.000500184
R20357 VDD.n4047 VDD.n4046 0.000500184
R20358 VDD.n4305 VDD.n4304 0.000500184
R20359 VDD.n4563 VDD.n4562 0.000500184
R20360 VDD.n4821 VDD.n4820 0.000500184
R20361 VDD.n5079 VDD.n5078 0.000500184
R20362 VDD.n5337 VDD.n5336 0.000500184
R20363 VDD.n1775 VDD.n1774 0.000500121
R20364 VDD.n2124 VDD.n2123 0.000500121
R20365 VDD.n2354 VDD.n2353 0.000500121
R20366 VDD.n2612 VDD.n2611 0.000500121
R20367 VDD.n2870 VDD.n2869 0.000500121
R20368 VDD.n3128 VDD.n3127 0.000500121
R20369 VDD.n3386 VDD.n3385 0.000500121
R20370 VDD.n3644 VDD.n3643 0.000500121
R20371 VDD.n3902 VDD.n3901 0.000500121
R20372 VDD.n4160 VDD.n4159 0.000500121
R20373 VDD.n4418 VDD.n4417 0.000500121
R20374 VDD.n4676 VDD.n4675 0.000500121
R20375 VDD.n4934 VDD.n4933 0.000500121
R20376 VDD.n5192 VDD.n5191 0.000500121
R20377 VDD.n2162 VDD.n1983 0.000500117
R20378 VDD.n2420 VDD.n2243 0.000500117
R20379 VDD.n2678 VDD.n2501 0.000500117
R20380 VDD.n2936 VDD.n2759 0.000500117
R20381 VDD.n3194 VDD.n3017 0.000500117
R20382 VDD.n3452 VDD.n3275 0.000500117
R20383 VDD.n5772 VDD.n5709 0.000500117
R20384 VDD.n5518 VDD.n5455 0.000500117
R20385 VDD.n3710 VDD.n3533 0.000500117
R20386 VDD.n3968 VDD.n3791 0.000500117
R20387 VDD.n4226 VDD.n4049 0.000500117
R20388 VDD.n4484 VDD.n4307 0.000500117
R20389 VDD.n4742 VDD.n4565 0.000500117
R20390 VDD.n5000 VDD.n4823 0.000500117
R20391 VDD.n5258 VDD.n5081 0.000500117
R20392 VDD.n1841 VDD.n1664 0.000500117
R20393 VDD.n1602 VDD.n1246 0.000500071
R20394 VDD.n1601 VDD.n1540 0.000500071
R20395 OUT3.n142 OUT3.n140 145.809
R20396 OUT3.n91 OUT3.n89 145.809
R20397 OUT3.n53 OUT3.n51 145.809
R20398 OUT3.n7 OUT3.n5 145.809
R20399 OUT3.n91 OUT3.n90 107.409
R20400 OUT3.n93 OUT3.n92 107.409
R20401 OUT3.n95 OUT3.n94 107.409
R20402 OUT3.n97 OUT3.n96 107.409
R20403 OUT3.n99 OUT3.n98 107.409
R20404 OUT3.n101 OUT3.n100 107.409
R20405 OUT3.n53 OUT3.n52 107.409
R20406 OUT3.n55 OUT3.n54 107.409
R20407 OUT3.n57 OUT3.n56 107.409
R20408 OUT3.n59 OUT3.n58 107.409
R20409 OUT3.n61 OUT3.n60 107.409
R20410 OUT3.n63 OUT3.n62 107.409
R20411 OUT3.n7 OUT3.n6 107.409
R20412 OUT3.n9 OUT3.n8 107.409
R20413 OUT3.n11 OUT3.n10 107.409
R20414 OUT3.n13 OUT3.n12 107.409
R20415 OUT3.n15 OUT3.n14 107.409
R20416 OUT3.n17 OUT3.n16 107.409
R20417 OUT3.n142 OUT3.n141 107.407
R20418 OUT3.n144 OUT3.n143 107.407
R20419 OUT3.n146 OUT3.n145 107.407
R20420 OUT3.n148 OUT3.n147 107.407
R20421 OUT3.n150 OUT3.n149 107.407
R20422 OUT3.n152 OUT3.n151 107.407
R20423 OUT3.n160 OUT3.n158 87.1779
R20424 OUT3.n114 OUT3.n112 87.1779
R20425 OUT3.n72 OUT3.n70 87.1779
R20426 OUT3.n26 OUT3.n24 87.1779
R20427 OUT3.n160 OUT3.n159 52.82
R20428 OUT3.n162 OUT3.n161 52.82
R20429 OUT3.n164 OUT3.n163 52.82
R20430 OUT3.n166 OUT3.n165 52.82
R20431 OUT3.n168 OUT3.n167 52.82
R20432 OUT3.n170 OUT3.n169 52.82
R20433 OUT3.n114 OUT3.n113 52.82
R20434 OUT3.n116 OUT3.n115 52.82
R20435 OUT3.n118 OUT3.n117 52.82
R20436 OUT3.n120 OUT3.n119 52.82
R20437 OUT3.n122 OUT3.n121 52.82
R20438 OUT3.n124 OUT3.n123 52.82
R20439 OUT3.n72 OUT3.n71 52.82
R20440 OUT3.n74 OUT3.n73 52.82
R20441 OUT3.n76 OUT3.n75 52.82
R20442 OUT3.n78 OUT3.n77 52.82
R20443 OUT3.n80 OUT3.n79 52.82
R20444 OUT3.n82 OUT3.n81 52.82
R20445 OUT3.n26 OUT3.n25 52.82
R20446 OUT3.n28 OUT3.n27 52.82
R20447 OUT3.n30 OUT3.n29 52.82
R20448 OUT3.n32 OUT3.n31 52.82
R20449 OUT3.n34 OUT3.n33 52.82
R20450 OUT3.n36 OUT3.n35 52.82
R20451 OUT3.n144 OUT3.n142 38.4005
R20452 OUT3.n146 OUT3.n144 38.4005
R20453 OUT3.n148 OUT3.n146 38.4005
R20454 OUT3.n150 OUT3.n148 38.4005
R20455 OUT3.n152 OUT3.n150 38.4005
R20456 OUT3.n153 OUT3.n152 38.4005
R20457 OUT3.n93 OUT3.n91 38.4005
R20458 OUT3.n95 OUT3.n93 38.4005
R20459 OUT3.n97 OUT3.n95 38.4005
R20460 OUT3.n99 OUT3.n97 38.4005
R20461 OUT3.n101 OUT3.n99 38.4005
R20462 OUT3.n102 OUT3.n101 38.4005
R20463 OUT3.n55 OUT3.n53 38.4005
R20464 OUT3.n57 OUT3.n55 38.4005
R20465 OUT3.n59 OUT3.n57 38.4005
R20466 OUT3.n61 OUT3.n59 38.4005
R20467 OUT3.n63 OUT3.n61 38.4005
R20468 OUT3.n64 OUT3.n63 38.4005
R20469 OUT3.n9 OUT3.n7 38.4005
R20470 OUT3.n11 OUT3.n9 38.4005
R20471 OUT3.n13 OUT3.n11 38.4005
R20472 OUT3.n15 OUT3.n13 38.4005
R20473 OUT3.n17 OUT3.n15 38.4005
R20474 OUT3.n18 OUT3.n17 38.4005
R20475 OUT3.n162 OUT3.n160 34.3584
R20476 OUT3.n164 OUT3.n162 34.3584
R20477 OUT3.n166 OUT3.n164 34.3584
R20478 OUT3.n168 OUT3.n166 34.3584
R20479 OUT3.n170 OUT3.n168 34.3584
R20480 OUT3.n174 OUT3.n170 34.3584
R20481 OUT3.n116 OUT3.n114 34.3584
R20482 OUT3.n118 OUT3.n116 34.3584
R20483 OUT3.n120 OUT3.n118 34.3584
R20484 OUT3.n122 OUT3.n120 34.3584
R20485 OUT3.n124 OUT3.n122 34.3584
R20486 OUT3.n129 OUT3.n124 34.3584
R20487 OUT3.n74 OUT3.n72 34.3584
R20488 OUT3.n76 OUT3.n74 34.3584
R20489 OUT3.n78 OUT3.n76 34.3584
R20490 OUT3.n80 OUT3.n78 34.3584
R20491 OUT3.n82 OUT3.n80 34.3584
R20492 OUT3.n83 OUT3.n82 34.3584
R20493 OUT3.n28 OUT3.n26 34.3584
R20494 OUT3.n30 OUT3.n28 34.3584
R20495 OUT3.n32 OUT3.n30 34.3584
R20496 OUT3.n34 OUT3.n32 34.3584
R20497 OUT3.n36 OUT3.n34 34.3584
R20498 OUT3.n40 OUT3.n36 34.3584
R20499 OUT3.n135 OUT3.t75 26.5955
R20500 OUT3.n135 OUT3.t101 26.5955
R20501 OUT3.n140 OUT3.t85 26.5955
R20502 OUT3.n140 OUT3.t124 26.5955
R20503 OUT3.n141 OUT3.t99 26.5955
R20504 OUT3.n141 OUT3.t72 26.5955
R20505 OUT3.n143 OUT3.t70 26.5955
R20506 OUT3.n143 OUT3.t83 26.5955
R20507 OUT3.n145 OUT3.t91 26.5955
R20508 OUT3.n145 OUT3.t107 26.5955
R20509 OUT3.n147 OUT3.t105 26.5955
R20510 OUT3.n147 OUT3.t127 26.5955
R20511 OUT3.n149 OUT3.t125 26.5955
R20512 OUT3.n149 OUT3.t89 26.5955
R20513 OUT3.n151 OUT3.t116 26.5955
R20514 OUT3.n151 OUT3.t77 26.5955
R20515 OUT3.n89 OUT3.t86 26.5955
R20516 OUT3.n89 OUT3.t112 26.5955
R20517 OUT3.n90 OUT3.t110 26.5955
R20518 OUT3.n90 OUT3.t73 26.5955
R20519 OUT3.n92 OUT3.t64 26.5955
R20520 OUT3.n92 OUT3.t94 26.5955
R20521 OUT3.n94 OUT3.t65 26.5955
R20522 OUT3.n94 OUT3.t81 26.5955
R20523 OUT3.n96 OUT3.t79 26.5955
R20524 OUT3.n96 OUT3.t97 26.5955
R20525 OUT3.n98 OUT3.t104 26.5955
R20526 OUT3.n98 OUT3.t118 26.5955
R20527 OUT3.n100 OUT3.t123 26.5955
R20528 OUT3.n100 OUT3.t88 26.5955
R20529 OUT3.n51 OUT3.t68 26.5955
R20530 OUT3.n51 OUT3.t113 26.5955
R20531 OUT3.n52 OUT3.t84 26.5955
R20532 OUT3.n52 OUT3.t100 26.5955
R20533 OUT3.n54 OUT3.t108 26.5955
R20534 OUT3.n54 OUT3.t71 26.5955
R20535 OUT3.n56 OUT3.t120 26.5955
R20536 OUT3.n56 OUT3.t82 26.5955
R20537 OUT3.n58 OUT3.t90 26.5955
R20538 OUT3.n58 OUT3.t106 26.5955
R20539 OUT3.n60 OUT3.t114 26.5955
R20540 OUT3.n60 OUT3.t126 26.5955
R20541 OUT3.n62 OUT3.t93 26.5955
R20542 OUT3.n62 OUT3.t69 26.5955
R20543 OUT3.n1 OUT3.t122 26.5955
R20544 OUT3.n1 OUT3.t67 26.5955
R20545 OUT3.n5 OUT3.t74 26.5955
R20546 OUT3.n5 OUT3.t87 26.5955
R20547 OUT3.n6 OUT3.t95 26.5955
R20548 OUT3.n6 OUT3.t111 26.5955
R20549 OUT3.n8 OUT3.t109 26.5955
R20550 OUT3.n8 OUT3.t121 26.5955
R20551 OUT3.n10 OUT3.t98 26.5955
R20552 OUT3.n10 OUT3.t92 26.5955
R20553 OUT3.n12 OUT3.t119 26.5955
R20554 OUT3.n12 OUT3.t80 26.5955
R20555 OUT3.n14 OUT3.t78 26.5955
R20556 OUT3.n14 OUT3.t96 26.5955
R20557 OUT3.n16 OUT3.t103 26.5955
R20558 OUT3.n16 OUT3.t117 26.5955
R20559 OUT3.n46 OUT3.t115 25.6105
R20560 OUT3.n171 OUT3.t27 24.9236
R20561 OUT3.n171 OUT3.t53 24.9236
R20562 OUT3.n158 OUT3.t37 24.9236
R20563 OUT3.n158 OUT3.t12 24.9236
R20564 OUT3.n159 OUT3.t51 24.9236
R20565 OUT3.n159 OUT3.t24 24.9236
R20566 OUT3.n161 OUT3.t22 24.9236
R20567 OUT3.n161 OUT3.t35 24.9236
R20568 OUT3.n163 OUT3.t43 24.9236
R20569 OUT3.n163 OUT3.t59 24.9236
R20570 OUT3.n165 OUT3.t57 24.9236
R20571 OUT3.n165 OUT3.t15 24.9236
R20572 OUT3.n167 OUT3.t13 24.9236
R20573 OUT3.n167 OUT3.t41 24.9236
R20574 OUT3.n169 OUT3.t4 24.9236
R20575 OUT3.n169 OUT3.t29 24.9236
R20576 OUT3.n112 OUT3.t38 24.9236
R20577 OUT3.n112 OUT3.t0 24.9236
R20578 OUT3.n113 OUT3.t62 24.9236
R20579 OUT3.n113 OUT3.t25 24.9236
R20580 OUT3.n115 OUT3.t16 24.9236
R20581 OUT3.n115 OUT3.t46 24.9236
R20582 OUT3.n117 OUT3.t17 24.9236
R20583 OUT3.n117 OUT3.t33 24.9236
R20584 OUT3.n119 OUT3.t31 24.9236
R20585 OUT3.n119 OUT3.t49 24.9236
R20586 OUT3.n121 OUT3.t56 24.9236
R20587 OUT3.n121 OUT3.t6 24.9236
R20588 OUT3.n123 OUT3.t11 24.9236
R20589 OUT3.n123 OUT3.t40 24.9236
R20590 OUT3.n70 OUT3.t20 24.9236
R20591 OUT3.n70 OUT3.t1 24.9236
R20592 OUT3.n71 OUT3.t36 24.9236
R20593 OUT3.n71 OUT3.t52 24.9236
R20594 OUT3.n73 OUT3.t60 24.9236
R20595 OUT3.n73 OUT3.t23 24.9236
R20596 OUT3.n75 OUT3.t8 24.9236
R20597 OUT3.n75 OUT3.t34 24.9236
R20598 OUT3.n77 OUT3.t42 24.9236
R20599 OUT3.n77 OUT3.t58 24.9236
R20600 OUT3.n79 OUT3.t2 24.9236
R20601 OUT3.n79 OUT3.t14 24.9236
R20602 OUT3.n81 OUT3.t45 24.9236
R20603 OUT3.n81 OUT3.t21 24.9236
R20604 OUT3.n37 OUT3.t10 24.9236
R20605 OUT3.n37 OUT3.t19 24.9236
R20606 OUT3.n24 OUT3.t26 24.9236
R20607 OUT3.n24 OUT3.t39 24.9236
R20608 OUT3.n25 OUT3.t47 24.9236
R20609 OUT3.n25 OUT3.t63 24.9236
R20610 OUT3.n27 OUT3.t61 24.9236
R20611 OUT3.n27 OUT3.t9 24.9236
R20612 OUT3.n29 OUT3.t50 24.9236
R20613 OUT3.n29 OUT3.t44 24.9236
R20614 OUT3.n31 OUT3.t7 24.9236
R20615 OUT3.n31 OUT3.t32 24.9236
R20616 OUT3.n33 OUT3.t30 24.9236
R20617 OUT3.n33 OUT3.t48 24.9236
R20618 OUT3.n35 OUT3.t55 24.9236
R20619 OUT3.n35 OUT3.t5 24.9236
R20620 OUT3.n68 OUT3.t3 24.7196
R20621 OUT3.n105 OUT3.t66 24.6255
R20622 OUT3.n68 OUT3.t28 23.9564
R20623 OUT3.n127 OUT3.t18 23.1655
R20624 OUT3.n103 OUT3.t102 19.1164
R20625 OUT3.n126 OUT3.n125 13.8467
R20626 OUT3 OUT3.n174 11.4429
R20627 OUT3 OUT3.n129 11.4429
R20628 OUT3 OUT3.n83 11.4429
R20629 OUT3 OUT3.n40 11.4429
R20630 OUT3.n125 OUT3.t54 11.0774
R20631 OUT3.n47 OUT3.t76 10.8355
R20632 OUT3.n106 OUT3.n105 9.3005
R20633 OUT3.n110 OUT3.n109 9.3005
R20634 OUT3.n128 OUT3.n127 8.77252
R20635 OUT3.n136 OUT3.n135 8.76605
R20636 OUT3.n2 OUT3.n1 8.76605
R20637 OUT3.n50 OUT3.n49 8.70762
R20638 OUT3.n49 OUT3.n48 8.69892
R20639 OUT3.n172 OUT3.n171 7.87147
R20640 OUT3.n38 OUT3.n37 7.87147
R20641 OUT3.n48 OUT3.n47 7.77627
R20642 OUT3.n104 OUT3.n103 7.29637
R20643 OUT3.n69 OUT3.n68 6.88889
R20644 OUT3.n85 OUT3.n69 4.758
R20645 OUT3.n128 OUT3.n111 4.6505
R20646 OUT3.n107 OUT3.n106 4.6505
R20647 OUT3.n39 OUT3.n23 4.6505
R20648 OUT3.n20 OUT3.n19 4.6505
R20649 OUT3.n3 OUT3.n2 4.26717
R20650 OUT3.n175 OUT3 3.10353
R20651 OUT3.n130 OUT3 3.10353
R20652 OUT3.n84 OUT3 3.10353
R20653 OUT3.n41 OUT3 3.10353
R20654 OUT3.n173 OUT3.n157 3.1005
R20655 OUT3.n137 OUT3.n136 3.1005
R20656 OUT3.n155 OUT3.n154 3.1005
R20657 OUT3.n66 OUT3.n65 2.75
R20658 OUT3.n154 OUT3.n153 2.71565
R20659 OUT3.n106 OUT3.n102 2.71565
R20660 OUT3.n65 OUT3.n64 2.71565
R20661 OUT3.n19 OUT3.n18 2.71565
R20662 OUT3.n66 OUT3.n50 2.69896
R20663 OUT3.n105 OUT3.n104 1.9705
R20664 OUT3.n174 OUT3 1.74595
R20665 OUT3 OUT3.n173 1.74595
R20666 OUT3.n129 OUT3 1.74595
R20667 OUT3 OUT3.n128 1.74595
R20668 OUT3.n83 OUT3 1.74595
R20669 OUT3.n40 OUT3 1.74595
R20670 OUT3 OUT3.n39 1.74595
R20671 OUT3.n127 OUT3.n126 1.74224
R20672 OUT3.n181 OUT3.n180 0.810582
R20673 OUT3 OUT3.n183 0.597838
R20674 OUT3.n183 OUT3.n182 0.531962
R20675 OUT3.n182 OUT3.n181 0.531962
R20676 OUT3.n182 OUT3.n86 0.475506
R20677 OUT3 OUT3.n69 0.388379
R20678 OUT3.n173 OUT3.n172 0.300854
R20679 OUT3.n39 OUT3.n38 0.300854
R20680 OUT3.n183 OUT3.n45 0.275505
R20681 OUT3.n181 OUT3.n134 0.263005
R20682 OUT3.n180 OUT3.n179 0.1755
R20683 OUT3.n134 OUT3.n133 0.1755
R20684 OUT3.n45 OUT3.n44 0.1755
R20685 OUT3.n176 OUT3.n157 0.11675
R20686 OUT3.n131 OUT3.n111 0.11675
R20687 OUT3.n42 OUT3.n23 0.11675
R20688 OUT3.n132 OUT3.n107 0.10425
R20689 OUT3.n178 OUT3.n155 0.09175
R20690 OUT3.n43 OUT3.n20 0.09175
R20691 OUT3.n86 OUT3.n66 0.0855244
R20692 OUT3.n49 OUT3.n46 0.0578287
R20693 OUT3.n86 OUT3.n85 0.0505
R20694 OUT3.n155 OUT3.n139 0.04425
R20695 OUT3.n20 OUT3.n4 0.04425
R20696 OUT3.n107 OUT3.n88 0.043
R20697 OUT3.n111 OUT3.n110 0.03175
R20698 OUT3.n139 OUT3.n137 0.028
R20699 OUT3.n4 OUT3.n0 0.028
R20700 OUT3.n178 OUT3.n176 0.0255
R20701 OUT3.n157 OUT3.n156 0.0255
R20702 OUT3.n43 OUT3.n42 0.0255
R20703 OUT3.n23 OUT3.n22 0.0255
R20704 OUT3.n132 OUT3.n131 0.013
R20705 OUT3.n88 OUT3.n87 0.00450862
R20706 OUT3.n139 OUT3.n138 0.0025557
R20707 OUT3.n4 OUT3.n3 0.0025557
R20708 OUT3.n176 OUT3.n175 0.00053521
R20709 OUT3.n131 OUT3.n130 0.00053521
R20710 OUT3.n85 OUT3.n84 0.00053521
R20711 OUT3.n42 OUT3.n41 0.00053521
R20712 OUT3.n178 OUT3.n177 0.00050852
R20713 OUT3.n132 OUT3.n108 0.00050852
R20714 OUT3.n86 OUT3.n67 0.00050852
R20715 OUT3.n43 OUT3.n21 0.00050852
R20716 OUT3.n179 OUT3.n178 0.000500999
R20717 OUT3.n133 OUT3.n132 0.000500999
R20718 OUT3.n44 OUT3.n43 0.000500999
R20719 frontAnalog_v0p0p1_15.x63.A.n2 frontAnalog_v0p0p1_15.x63.A.t4 260.322
R20720 frontAnalog_v0p0p1_15.x63.A.n4 frontAnalog_v0p0p1_15.x63.A.t5 233.888
R20721 frontAnalog_v0p0p1_15.x63.A.n2 frontAnalog_v0p0p1_15.x63.A.t6 175.169
R20722 frontAnalog_v0p0p1_15.x63.A.n3 frontAnalog_v0p0p1_15.x63.A.t7 159.725
R20723 frontAnalog_v0p0p1_15.x63.A.n1 frontAnalog_v0p0p1_15.x63.A.t3 17.4109
R20724 frontAnalog_v0p0p1_15.x63.A.n0 frontAnalog_v0p0p1_15.x63.A.n2 9.75129
R20725 frontAnalog_v0p0p1_15.x63.A.n1 frontAnalog_v0p0p1_15.x63.A.t2 9.6037
R20726 frontAnalog_v0p0p1_15.x63.A.n0 frontAnalog_v0p0p1_15.x63.A 2.33338
R20727 frontAnalog_v0p0p1_15.x63.A.n5 frontAnalog_v0p0p1_15.x63.A.t1 8.40929
R20728 frontAnalog_v0p0p1_15.x63.A.n3 frontAnalog_v0p0p1_15.x63.A.t0 8.06629
R20729 frontAnalog_v0p0p1_15.x63.A.n4 frontAnalog_v0p0p1_15.x63.A.n3 1.73501
R20730 frontAnalog_v0p0p1_15.x63.A.n1 frontAnalog_v0p0p1_15.x63.A.n4 0.99025
R20731 frontAnalog_v0p0p1_15.x63.A.n5 frontAnalog_v0p0p1_15.x63.A.n1 0.853186
R20732 frontAnalog_v0p0p1_15.x63.A frontAnalog_v0p0p1_15.x63.A.n0 0.349517
R20733 frontAnalog_v0p0p1_15.x63.A frontAnalog_v0p0p1_15.x63.A.n5 0.24425
R20734 OUT0.n122 OUT0.n120 145.809
R20735 OUT0.n65 OUT0.n63 145.809
R20736 OUT0.n25 OUT0.n23 145.809
R20737 OUT0.n102 OUT0.n100 145.808
R20738 OUT0.n65 OUT0.n64 107.409
R20739 OUT0.n67 OUT0.n66 107.409
R20740 OUT0.n69 OUT0.n68 107.409
R20741 OUT0.n71 OUT0.n70 107.409
R20742 OUT0.n73 OUT0.n72 107.409
R20743 OUT0.n75 OUT0.n74 107.409
R20744 OUT0.n25 OUT0.n24 107.409
R20745 OUT0.n27 OUT0.n26 107.409
R20746 OUT0.n29 OUT0.n28 107.409
R20747 OUT0.n31 OUT0.n30 107.409
R20748 OUT0.n33 OUT0.n32 107.409
R20749 OUT0.n35 OUT0.n34 107.409
R20750 OUT0.n122 OUT0.n121 107.407
R20751 OUT0.n124 OUT0.n123 107.407
R20752 OUT0.n126 OUT0.n125 107.407
R20753 OUT0.n128 OUT0.n127 107.407
R20754 OUT0.n130 OUT0.n129 107.407
R20755 OUT0.n132 OUT0.n131 107.407
R20756 OUT0.n102 OUT0.n101 107.407
R20757 OUT0.n104 OUT0.n103 107.407
R20758 OUT0.n106 OUT0.n105 107.407
R20759 OUT0.n108 OUT0.n107 107.407
R20760 OUT0.n110 OUT0.n109 107.407
R20761 OUT0.n112 OUT0.n111 107.407
R20762 OUT0.n138 OUT0.n136 87.1779
R20763 OUT0.n83 OUT0.n81 87.1779
R20764 OUT0.n44 OUT0.n42 87.1779
R20765 OUT0.n4 OUT0.n2 87.1779
R20766 OUT0.n54 OUT0.n53 52.82
R20767 OUT0.n14 OUT0.n13 52.82
R20768 OUT0.n138 OUT0.n137 52.82
R20769 OUT0.n140 OUT0.n139 52.82
R20770 OUT0.n142 OUT0.n141 52.82
R20771 OUT0.n144 OUT0.n143 52.82
R20772 OUT0.n146 OUT0.n145 52.82
R20773 OUT0.n148 OUT0.n147 52.82
R20774 OUT0.n83 OUT0.n82 52.82
R20775 OUT0.n85 OUT0.n84 52.82
R20776 OUT0.n87 OUT0.n86 52.82
R20777 OUT0.n89 OUT0.n88 52.82
R20778 OUT0.n91 OUT0.n90 52.82
R20779 OUT0.n93 OUT0.n92 52.82
R20780 OUT0.n44 OUT0.n43 52.82
R20781 OUT0.n46 OUT0.n45 52.82
R20782 OUT0.n48 OUT0.n47 52.82
R20783 OUT0.n50 OUT0.n49 52.82
R20784 OUT0.n52 OUT0.n51 52.82
R20785 OUT0.n4 OUT0.n3 52.82
R20786 OUT0.n6 OUT0.n5 52.82
R20787 OUT0.n8 OUT0.n7 52.82
R20788 OUT0.n10 OUT0.n9 52.82
R20789 OUT0.n12 OUT0.n11 52.82
R20790 OUT0 OUT0.n149 51.0745
R20791 OUT0 OUT0.n94 51.0745
R20792 OUT0.n124 OUT0.n122 38.4005
R20793 OUT0.n126 OUT0.n124 38.4005
R20794 OUT0.n128 OUT0.n126 38.4005
R20795 OUT0.n130 OUT0.n128 38.4005
R20796 OUT0.n132 OUT0.n130 38.4005
R20797 OUT0.n133 OUT0.n132 38.4005
R20798 OUT0.n104 OUT0.n102 38.4005
R20799 OUT0.n106 OUT0.n104 38.4005
R20800 OUT0.n108 OUT0.n106 38.4005
R20801 OUT0.n110 OUT0.n108 38.4005
R20802 OUT0.n112 OUT0.n110 38.4005
R20803 OUT0.n113 OUT0.n112 38.4005
R20804 OUT0.n67 OUT0.n65 38.4005
R20805 OUT0.n69 OUT0.n67 38.4005
R20806 OUT0.n71 OUT0.n69 38.4005
R20807 OUT0.n73 OUT0.n71 38.4005
R20808 OUT0.n75 OUT0.n73 38.4005
R20809 OUT0.n76 OUT0.n75 38.4005
R20810 OUT0.n27 OUT0.n25 38.4005
R20811 OUT0.n29 OUT0.n27 38.4005
R20812 OUT0.n31 OUT0.n29 38.4005
R20813 OUT0.n33 OUT0.n31 38.4005
R20814 OUT0.n35 OUT0.n33 38.4005
R20815 OUT0.n36 OUT0.n35 38.4005
R20816 OUT0.n140 OUT0.n138 34.3584
R20817 OUT0.n142 OUT0.n140 34.3584
R20818 OUT0.n144 OUT0.n142 34.3584
R20819 OUT0.n146 OUT0.n144 34.3584
R20820 OUT0.n148 OUT0.n146 34.3584
R20821 OUT0.n150 OUT0.n148 34.3584
R20822 OUT0.n85 OUT0.n83 34.3584
R20823 OUT0.n87 OUT0.n85 34.3584
R20824 OUT0.n89 OUT0.n87 34.3584
R20825 OUT0.n91 OUT0.n89 34.3584
R20826 OUT0.n93 OUT0.n91 34.3584
R20827 OUT0.n95 OUT0.n93 34.3584
R20828 OUT0.n46 OUT0.n44 34.3584
R20829 OUT0.n48 OUT0.n46 34.3584
R20830 OUT0.n50 OUT0.n48 34.3584
R20831 OUT0.n52 OUT0.n50 34.3584
R20832 OUT0.n54 OUT0.n52 34.3584
R20833 OUT0.n58 OUT0.n54 34.3584
R20834 OUT0.n6 OUT0.n4 34.3584
R20835 OUT0.n8 OUT0.n6 34.3584
R20836 OUT0.n10 OUT0.n8 34.3584
R20837 OUT0.n12 OUT0.n10 34.3584
R20838 OUT0.n14 OUT0.n12 34.3584
R20839 OUT0.n18 OUT0.n14 34.3584
R20840 OUT0.n118 OUT0.t105 26.5955
R20841 OUT0.n118 OUT0.t118 26.5955
R20842 OUT0.n120 OUT0.t103 26.5955
R20843 OUT0.n120 OUT0.t75 26.5955
R20844 OUT0.n121 OUT0.t125 26.5955
R20845 OUT0.n121 OUT0.t91 26.5955
R20846 OUT0.n123 OUT0.t70 26.5955
R20847 OUT0.n123 OUT0.t111 26.5955
R20848 OUT0.n125 OUT0.t81 26.5955
R20849 OUT0.n125 OUT0.t99 26.5955
R20850 OUT0.n127 OUT0.t97 26.5955
R20851 OUT0.n127 OUT0.t114 26.5955
R20852 OUT0.n129 OUT0.t120 26.5955
R20853 OUT0.n129 OUT0.t86 26.5955
R20854 OUT0.n131 OUT0.t67 26.5955
R20855 OUT0.n131 OUT0.t107 26.5955
R20856 OUT0.n99 OUT0.t66 26.5955
R20857 OUT0.n99 OUT0.t95 26.5955
R20858 OUT0.n100 OUT0.t85 26.5955
R20859 OUT0.n100 OUT0.t94 26.5955
R20860 OUT0.n101 OUT0.t101 26.5955
R20861 OUT0.n101 OUT0.t74 26.5955
R20862 OUT0.n103 OUT0.t116 26.5955
R20863 OUT0.n103 OUT0.t88 26.5955
R20864 OUT0.n105 OUT0.t87 26.5955
R20865 OUT0.n105 OUT0.t100 26.5955
R20866 OUT0.n107 OUT0.t108 26.5955
R20867 OUT0.n107 OUT0.t122 26.5955
R20868 OUT0.n109 OUT0.t121 26.5955
R20869 OUT0.n109 OUT0.t76 26.5955
R20870 OUT0.n111 OUT0.t110 26.5955
R20871 OUT0.n111 OUT0.t78 26.5955
R20872 OUT0.n62 OUT0.t72 26.5955
R20873 OUT0.n62 OUT0.t106 26.5955
R20874 OUT0.n63 OUT0.t92 26.5955
R20875 OUT0.n63 OUT0.t104 26.5955
R20876 OUT0.n64 OUT0.t102 26.5955
R20877 OUT0.n64 OUT0.t126 26.5955
R20878 OUT0.n66 OUT0.t123 26.5955
R20879 OUT0.n66 OUT0.t89 26.5955
R20880 OUT0.n68 OUT0.t115 26.5955
R20881 OUT0.n68 OUT0.t83 26.5955
R20882 OUT0.n70 OUT0.t79 26.5955
R20883 OUT0.n70 OUT0.t98 26.5955
R20884 OUT0.n72 OUT0.t96 26.5955
R20885 OUT0.n72 OUT0.t113 26.5955
R20886 OUT0.n74 OUT0.t119 26.5955
R20887 OUT0.n74 OUT0.t68 26.5955
R20888 OUT0.n22 OUT0.t71 26.5955
R20889 OUT0.n22 OUT0.t84 26.5955
R20890 OUT0.n23 OUT0.t90 26.5955
R20891 OUT0.n23 OUT0.t112 26.5955
R20892 OUT0.n24 OUT0.t109 26.5955
R20893 OUT0.n24 OUT0.t124 26.5955
R20894 OUT0.n26 OUT0.t65 26.5955
R20895 OUT0.n26 OUT0.t77 26.5955
R20896 OUT0.n28 OUT0.t82 26.5955
R20897 OUT0.n28 OUT0.t117 26.5955
R20898 OUT0.n30 OUT0.t93 26.5955
R20899 OUT0.n30 OUT0.t64 26.5955
R20900 OUT0.n32 OUT0.t69 26.5955
R20901 OUT0.n32 OUT0.t80 26.5955
R20902 OUT0.n34 OUT0.t127 26.5955
R20903 OUT0.n34 OUT0.t73 26.5955
R20904 OUT0.n149 OUT0.t41 24.9236
R20905 OUT0.n149 OUT0.t54 24.9236
R20906 OUT0.n136 OUT0.t39 24.9236
R20907 OUT0.n136 OUT0.t11 24.9236
R20908 OUT0.n137 OUT0.t61 24.9236
R20909 OUT0.n137 OUT0.t27 24.9236
R20910 OUT0.n139 OUT0.t6 24.9236
R20911 OUT0.n139 OUT0.t47 24.9236
R20912 OUT0.n141 OUT0.t17 24.9236
R20913 OUT0.n141 OUT0.t35 24.9236
R20914 OUT0.n143 OUT0.t33 24.9236
R20915 OUT0.n143 OUT0.t50 24.9236
R20916 OUT0.n145 OUT0.t56 24.9236
R20917 OUT0.n145 OUT0.t22 24.9236
R20918 OUT0.n147 OUT0.t3 24.9236
R20919 OUT0.n147 OUT0.t43 24.9236
R20920 OUT0.n94 OUT0.t2 24.9236
R20921 OUT0.n94 OUT0.t31 24.9236
R20922 OUT0.n81 OUT0.t21 24.9236
R20923 OUT0.n81 OUT0.t30 24.9236
R20924 OUT0.n82 OUT0.t37 24.9236
R20925 OUT0.n82 OUT0.t10 24.9236
R20926 OUT0.n84 OUT0.t52 24.9236
R20927 OUT0.n84 OUT0.t24 24.9236
R20928 OUT0.n86 OUT0.t23 24.9236
R20929 OUT0.n86 OUT0.t36 24.9236
R20930 OUT0.n88 OUT0.t44 24.9236
R20931 OUT0.n88 OUT0.t58 24.9236
R20932 OUT0.n90 OUT0.t57 24.9236
R20933 OUT0.n90 OUT0.t12 24.9236
R20934 OUT0.n92 OUT0.t46 24.9236
R20935 OUT0.n92 OUT0.t14 24.9236
R20936 OUT0.n55 OUT0.t8 24.9236
R20937 OUT0.n55 OUT0.t42 24.9236
R20938 OUT0.n42 OUT0.t28 24.9236
R20939 OUT0.n42 OUT0.t40 24.9236
R20940 OUT0.n43 OUT0.t38 24.9236
R20941 OUT0.n43 OUT0.t62 24.9236
R20942 OUT0.n45 OUT0.t59 24.9236
R20943 OUT0.n45 OUT0.t25 24.9236
R20944 OUT0.n47 OUT0.t51 24.9236
R20945 OUT0.n47 OUT0.t19 24.9236
R20946 OUT0.n49 OUT0.t15 24.9236
R20947 OUT0.n49 OUT0.t34 24.9236
R20948 OUT0.n51 OUT0.t32 24.9236
R20949 OUT0.n51 OUT0.t49 24.9236
R20950 OUT0.n53 OUT0.t55 24.9236
R20951 OUT0.n53 OUT0.t4 24.9236
R20952 OUT0.n15 OUT0.t7 24.9236
R20953 OUT0.n15 OUT0.t20 24.9236
R20954 OUT0.n2 OUT0.t26 24.9236
R20955 OUT0.n2 OUT0.t48 24.9236
R20956 OUT0.n3 OUT0.t45 24.9236
R20957 OUT0.n3 OUT0.t60 24.9236
R20958 OUT0.n5 OUT0.t1 24.9236
R20959 OUT0.n5 OUT0.t13 24.9236
R20960 OUT0.n7 OUT0.t18 24.9236
R20961 OUT0.n7 OUT0.t53 24.9236
R20962 OUT0.n9 OUT0.t29 24.9236
R20963 OUT0.n9 OUT0.t0 24.9236
R20964 OUT0.n11 OUT0.t5 24.9236
R20965 OUT0.n11 OUT0.t16 24.9236
R20966 OUT0.n13 OUT0.t63 24.9236
R20967 OUT0.n13 OUT0.t9 24.9236
R20968 OUT0 OUT0.n150 11.4429
R20969 OUT0 OUT0.n95 11.4429
R20970 OUT0 OUT0.n58 11.4429
R20971 OUT0 OUT0.n18 11.4429
R20972 OUT0.n77 OUT0.n62 8.55118
R20973 OUT0.n37 OUT0.n22 8.55118
R20974 OUT0.n114 OUT0.n99 8.55117
R20975 OUT0.n119 OUT0.n118 8.47293
R20976 OUT0.n56 OUT0.n55 7.80093
R20977 OUT0.n16 OUT0.n15 7.80093
R20978 OUT0.n78 OUT0.n77 3.20954
R20979 OUT0.n38 OUT0.n37 3.20953
R20980 OUT0.n115 OUT0.n114 3.20289
R20981 OUT0.n151 OUT0 3.10353
R20982 OUT0.n96 OUT0 3.10353
R20983 OUT0.n59 OUT0 3.10353
R20984 OUT0.n19 OUT0 3.10353
R20985 OUT0.n135 OUT0.n134 3.1005
R20986 OUT0.n57 OUT0.n41 3.1005
R20987 OUT0.n17 OUT0.n1 3.1005
R20988 OUT0.n134 OUT0.n133 2.71565
R20989 OUT0.n114 OUT0.n113 2.13383
R20990 OUT0.n77 OUT0.n76 2.13383
R20991 OUT0.n37 OUT0.n36 2.13383
R20992 OUT0.n150 OUT0 1.74595
R20993 OUT0.n95 OUT0 1.74595
R20994 OUT0.n58 OUT0.n57 1.16414
R20995 OUT0.n18 OUT0.n17 1.16414
R20996 OUT0.n157 OUT0.n156 1.07337
R20997 OUT0.n158 OUT0.n157 0.69375
R20998 OUT0.n159 OUT0.n158 0.68905
R20999 OUT0.n56 OUT0 0.488972
R21000 OUT0.n16 OUT0 0.488972
R21001 OUT0.n158 OUT0.n79 0.414635
R21002 OUT0.n157 OUT0.n116 0.382465
R21003 OUT0.n159 OUT0.n39 0.368576
R21004 OUT0 OUT0.n159 0.281623
R21005 OUT0.n134 OUT0.n119 0.196887
R21006 OUT0.n79 OUT0.n78 0.157252
R21007 OUT0.n39 OUT0.n38 0.139891
R21008 OUT0.n156 OUT0.n155 0.139389
R21009 OUT0.n116 OUT0.n115 0.132946
R21010 OUT0.n60 OUT0.n41 0.113
R21011 OUT0.n20 OUT0.n1 0.113
R21012 OUT0.n154 OUT0.n135 0.101889
R21013 OUT0.n57 OUT0.n56 0.0893205
R21014 OUT0.n17 OUT0.n16 0.0893205
R21015 OUT0.n154 OUT0.n152 0.0282778
R21016 OUT0.n135 OUT0.n117 0.0268889
R21017 OUT0.n98 OUT0.n97 0.0213333
R21018 OUT0.n61 OUT0.n60 0.0143889
R21019 OUT0.n21 OUT0.n20 0.0143889
R21020 OUT0.n115 OUT0.n98 0.00100004
R21021 OUT0.n38 OUT0.n21 0.00100004
R21022 OUT0.n78 OUT0.n61 0.00100004
R21023 OUT0.n152 OUT0.n151 0.000513335
R21024 OUT0.n97 OUT0.n96 0.000513335
R21025 OUT0.n60 OUT0.n59 0.000513218
R21026 OUT0.n20 OUT0.n19 0.000513218
R21027 OUT0.n98 OUT0.n80 0.00050517
R21028 OUT0.n154 OUT0.n153 0.000504838
R21029 OUT0.n61 OUT0.n40 0.000504838
R21030 OUT0.n21 OUT0.n0 0.000504838
R21031 OUT0.n155 OUT0.n154 0.000501713
R21032 I5.t11 I5.t13 618.109
R21033 I5.n12 I5.t6 259.74
R21034 I5 I5.t11 253.56
R21035 I5.n3 I5.t9 228.899
R21036 I5.n18 I5.t7 180.286
R21037 I5.n3 I5.t8 159.411
R21038 I5.n12 I5.t10 157.083
R21039 I5.n20 I5.n19 152
R21040 I5.n26 I5.t5 117.314
R21041 I5.n20 I5.t14 111.091
R21042 I5.n26 I5.t12 110.853
R21043 I5.n18 I5.n17 74.4551
R21044 I5.n24 I5 37.6855
R21045 I5.n28 I5.t2 17.6181
R21046 I5.n29 I5.t4 14.2865
R21047 I5.n31 I5.t1 14.283
R21048 I5.n31 I5.t0 14.283
R21049 I5.n6 I5.n2 9.3005
R21050 I5.n6 I5.n5 9.3005
R21051 I5.n21 I5.n20 9.3005
R21052 I5.n14 I5 9.3005
R21053 I5.n33 I5.t3 8.77744
R21054 I5.n22 I5.n21 7.80966
R21055 I5.n13 I5.n12 7.57248
R21056 I5.n5 I5.n3 7.36978
R21057 I5.n20 I5.n18 6.53562
R21058 I5 I5.n13 4.8645
R21059 I5.n14 I5.n10 4.50988
R21060 I5.n4 I5.n2 3.46717
R21061 I5 I5.n34 3.14231
R21062 I5.n4 I5.n1 3.03286
R21063 I5.n19 I5.n17 2.32777
R21064 I5.n8 I5.n0 2.26553
R21065 I5.n7 I5.n1 2.26468
R21066 I5.n16 I5.n15 2.251
R21067 I5.n22 I5.n16 2.19001
R21068 I5.n19 I5 1.4966
R21069 I5.n23 I5.n9 1.36032
R21070 I5.n33 I5.n32 1.20426
R21071 I5.n23 I5.n22 1.07639
R21072 I5.n5 I5.n4 1.06717
R21073 I5.n2 I5 1.06717
R21074 I5.n9 I5.n8 0.71595
R21075 I5.n35 I5 0.588
R21076 I5 I5.n25 0.577033
R21077 I5.n21 I5.n17 0.499201
R21078 I5 I5.n35 0.441125
R21079 I5.n25 I5.n24 0.435179
R21080 I5.n34 I5.n33 0.32511
R21081 I5.n29 I5.n28 0.314673
R21082 I5.n30 I5.n29 0.299251
R21083 I5.n9 I5 0.221483
R21084 I5.n25 I5 0.20675
R21085 I5.n27 I5.n26 0.159555
R21086 I5.n32 I5.n31 0.106617
R21087 I5.n30 I5.n27 0.0796167
R21088 I5.n32 I5.n30 0.0480595
R21089 I5.n34 I5 0.046937
R21090 I5.n15 I5.n14 0.0301875
R21091 I5.n16 I5.n10 0.0205312
R21092 I5.n35 I5 0.0161667
R21093 I5.n35 I5 0.01225
R21094 I5.n6 I5.n0 0.00618182
R21095 I5.n1 I5.n0 0.00555107
R21096 I5.n7 I5.n6 0.00530477
R21097 I5.n11 I5.n10 0.00210765
R21098 I5.n13 I5.n11 0.00133438
R21099 I5.n8 I5.n7 0.00101192
R21100 I5.n15 I5.n11 0.00100001
R21101 I5.n24 I5.n23 0.000507778
R21102 I5.n28 I5.n27 0.000504658
R21103 OUT2.n122 OUT2.n120 145.809
R21104 OUT2.n65 OUT2.n63 145.809
R21105 OUT2.n25 OUT2.n23 145.809
R21106 OUT2.n102 OUT2.n100 145.808
R21107 OUT2.n65 OUT2.n64 107.409
R21108 OUT2.n67 OUT2.n66 107.409
R21109 OUT2.n69 OUT2.n68 107.409
R21110 OUT2.n71 OUT2.n70 107.409
R21111 OUT2.n73 OUT2.n72 107.409
R21112 OUT2.n75 OUT2.n74 107.409
R21113 OUT2.n25 OUT2.n24 107.409
R21114 OUT2.n27 OUT2.n26 107.409
R21115 OUT2.n29 OUT2.n28 107.409
R21116 OUT2.n31 OUT2.n30 107.409
R21117 OUT2.n33 OUT2.n32 107.409
R21118 OUT2.n35 OUT2.n34 107.409
R21119 OUT2.n122 OUT2.n121 107.407
R21120 OUT2.n124 OUT2.n123 107.407
R21121 OUT2.n126 OUT2.n125 107.407
R21122 OUT2.n128 OUT2.n127 107.407
R21123 OUT2.n130 OUT2.n129 107.407
R21124 OUT2.n132 OUT2.n131 107.407
R21125 OUT2.n102 OUT2.n101 107.407
R21126 OUT2.n104 OUT2.n103 107.407
R21127 OUT2.n106 OUT2.n105 107.407
R21128 OUT2.n108 OUT2.n107 107.407
R21129 OUT2.n110 OUT2.n109 107.407
R21130 OUT2.n112 OUT2.n111 107.407
R21131 OUT2.n138 OUT2.n136 87.1779
R21132 OUT2.n83 OUT2.n81 87.1779
R21133 OUT2.n44 OUT2.n42 87.1779
R21134 OUT2.n4 OUT2.n2 87.1779
R21135 OUT2.n54 OUT2.n53 52.82
R21136 OUT2.n14 OUT2.n13 52.82
R21137 OUT2.n138 OUT2.n137 52.82
R21138 OUT2.n140 OUT2.n139 52.82
R21139 OUT2.n142 OUT2.n141 52.82
R21140 OUT2.n144 OUT2.n143 52.82
R21141 OUT2.n146 OUT2.n145 52.82
R21142 OUT2.n148 OUT2.n147 52.82
R21143 OUT2.n83 OUT2.n82 52.82
R21144 OUT2.n85 OUT2.n84 52.82
R21145 OUT2.n87 OUT2.n86 52.82
R21146 OUT2.n89 OUT2.n88 52.82
R21147 OUT2.n91 OUT2.n90 52.82
R21148 OUT2.n93 OUT2.n92 52.82
R21149 OUT2.n44 OUT2.n43 52.82
R21150 OUT2.n46 OUT2.n45 52.82
R21151 OUT2.n48 OUT2.n47 52.82
R21152 OUT2.n50 OUT2.n49 52.82
R21153 OUT2.n52 OUT2.n51 52.82
R21154 OUT2.n4 OUT2.n3 52.82
R21155 OUT2.n6 OUT2.n5 52.82
R21156 OUT2.n8 OUT2.n7 52.82
R21157 OUT2.n10 OUT2.n9 52.82
R21158 OUT2.n12 OUT2.n11 52.82
R21159 OUT2 OUT2.n149 51.0745
R21160 OUT2 OUT2.n94 51.0745
R21161 OUT2.n124 OUT2.n122 38.4005
R21162 OUT2.n126 OUT2.n124 38.4005
R21163 OUT2.n128 OUT2.n126 38.4005
R21164 OUT2.n130 OUT2.n128 38.4005
R21165 OUT2.n132 OUT2.n130 38.4005
R21166 OUT2.n133 OUT2.n132 38.4005
R21167 OUT2.n104 OUT2.n102 38.4005
R21168 OUT2.n106 OUT2.n104 38.4005
R21169 OUT2.n108 OUT2.n106 38.4005
R21170 OUT2.n110 OUT2.n108 38.4005
R21171 OUT2.n112 OUT2.n110 38.4005
R21172 OUT2.n113 OUT2.n112 38.4005
R21173 OUT2.n67 OUT2.n65 38.4005
R21174 OUT2.n69 OUT2.n67 38.4005
R21175 OUT2.n71 OUT2.n69 38.4005
R21176 OUT2.n73 OUT2.n71 38.4005
R21177 OUT2.n75 OUT2.n73 38.4005
R21178 OUT2.n76 OUT2.n75 38.4005
R21179 OUT2.n27 OUT2.n25 38.4005
R21180 OUT2.n29 OUT2.n27 38.4005
R21181 OUT2.n31 OUT2.n29 38.4005
R21182 OUT2.n33 OUT2.n31 38.4005
R21183 OUT2.n35 OUT2.n33 38.4005
R21184 OUT2.n36 OUT2.n35 38.4005
R21185 OUT2.n140 OUT2.n138 34.3584
R21186 OUT2.n142 OUT2.n140 34.3584
R21187 OUT2.n144 OUT2.n142 34.3584
R21188 OUT2.n146 OUT2.n144 34.3584
R21189 OUT2.n148 OUT2.n146 34.3584
R21190 OUT2.n150 OUT2.n148 34.3584
R21191 OUT2.n85 OUT2.n83 34.3584
R21192 OUT2.n87 OUT2.n85 34.3584
R21193 OUT2.n89 OUT2.n87 34.3584
R21194 OUT2.n91 OUT2.n89 34.3584
R21195 OUT2.n93 OUT2.n91 34.3584
R21196 OUT2.n95 OUT2.n93 34.3584
R21197 OUT2.n46 OUT2.n44 34.3584
R21198 OUT2.n48 OUT2.n46 34.3584
R21199 OUT2.n50 OUT2.n48 34.3584
R21200 OUT2.n52 OUT2.n50 34.3584
R21201 OUT2.n54 OUT2.n52 34.3584
R21202 OUT2.n58 OUT2.n54 34.3584
R21203 OUT2.n6 OUT2.n4 34.3584
R21204 OUT2.n8 OUT2.n6 34.3584
R21205 OUT2.n10 OUT2.n8 34.3584
R21206 OUT2.n12 OUT2.n10 34.3584
R21207 OUT2.n14 OUT2.n12 34.3584
R21208 OUT2.n18 OUT2.n14 34.3584
R21209 OUT2.n118 OUT2.t116 26.5955
R21210 OUT2.n118 OUT2.t65 26.5955
R21211 OUT2.n120 OUT2.t114 26.5955
R21212 OUT2.n120 OUT2.t86 26.5955
R21213 OUT2.n121 OUT2.t72 26.5955
R21214 OUT2.n121 OUT2.t102 26.5955
R21215 OUT2.n123 OUT2.t81 26.5955
R21216 OUT2.n123 OUT2.t122 26.5955
R21217 OUT2.n125 OUT2.t92 26.5955
R21218 OUT2.n125 OUT2.t110 26.5955
R21219 OUT2.n127 OUT2.t108 26.5955
R21220 OUT2.n127 OUT2.t125 26.5955
R21221 OUT2.n129 OUT2.t67 26.5955
R21222 OUT2.n129 OUT2.t97 26.5955
R21223 OUT2.n131 OUT2.t78 26.5955
R21224 OUT2.n131 OUT2.t118 26.5955
R21225 OUT2.n99 OUT2.t77 26.5955
R21226 OUT2.n99 OUT2.t106 26.5955
R21227 OUT2.n100 OUT2.t96 26.5955
R21228 OUT2.n100 OUT2.t105 26.5955
R21229 OUT2.n101 OUT2.t112 26.5955
R21230 OUT2.n101 OUT2.t85 26.5955
R21231 OUT2.n103 OUT2.t127 26.5955
R21232 OUT2.n103 OUT2.t99 26.5955
R21233 OUT2.n105 OUT2.t98 26.5955
R21234 OUT2.n105 OUT2.t111 26.5955
R21235 OUT2.n107 OUT2.t119 26.5955
R21236 OUT2.n107 OUT2.t69 26.5955
R21237 OUT2.n109 OUT2.t68 26.5955
R21238 OUT2.n109 OUT2.t87 26.5955
R21239 OUT2.n111 OUT2.t121 26.5955
R21240 OUT2.n111 OUT2.t89 26.5955
R21241 OUT2.n62 OUT2.t83 26.5955
R21242 OUT2.n62 OUT2.t117 26.5955
R21243 OUT2.n63 OUT2.t103 26.5955
R21244 OUT2.n63 OUT2.t115 26.5955
R21245 OUT2.n64 OUT2.t113 26.5955
R21246 OUT2.n64 OUT2.t73 26.5955
R21247 OUT2.n66 OUT2.t70 26.5955
R21248 OUT2.n66 OUT2.t100 26.5955
R21249 OUT2.n68 OUT2.t126 26.5955
R21250 OUT2.n68 OUT2.t94 26.5955
R21251 OUT2.n70 OUT2.t91 26.5955
R21252 OUT2.n70 OUT2.t109 26.5955
R21253 OUT2.n72 OUT2.t107 26.5955
R21254 OUT2.n72 OUT2.t124 26.5955
R21255 OUT2.n74 OUT2.t66 26.5955
R21256 OUT2.n74 OUT2.t79 26.5955
R21257 OUT2.n22 OUT2.t82 26.5955
R21258 OUT2.n22 OUT2.t95 26.5955
R21259 OUT2.n23 OUT2.t101 26.5955
R21260 OUT2.n23 OUT2.t123 26.5955
R21261 OUT2.n24 OUT2.t120 26.5955
R21262 OUT2.n24 OUT2.t71 26.5955
R21263 OUT2.n26 OUT2.t76 26.5955
R21264 OUT2.n26 OUT2.t88 26.5955
R21265 OUT2.n28 OUT2.t93 26.5955
R21266 OUT2.n28 OUT2.t64 26.5955
R21267 OUT2.n30 OUT2.t104 26.5955
R21268 OUT2.n30 OUT2.t75 26.5955
R21269 OUT2.n32 OUT2.t80 26.5955
R21270 OUT2.n32 OUT2.t90 26.5955
R21271 OUT2.n34 OUT2.t74 26.5955
R21272 OUT2.n34 OUT2.t84 26.5955
R21273 OUT2.n149 OUT2.t6 24.9236
R21274 OUT2.n149 OUT2.t19 24.9236
R21275 OUT2.n136 OUT2.t4 24.9236
R21276 OUT2.n136 OUT2.t40 24.9236
R21277 OUT2.n137 OUT2.t26 24.9236
R21278 OUT2.n137 OUT2.t56 24.9236
R21279 OUT2.n139 OUT2.t35 24.9236
R21280 OUT2.n139 OUT2.t12 24.9236
R21281 OUT2.n141 OUT2.t46 24.9236
R21282 OUT2.n141 OUT2.t0 24.9236
R21283 OUT2.n143 OUT2.t62 24.9236
R21284 OUT2.n143 OUT2.t15 24.9236
R21285 OUT2.n145 OUT2.t21 24.9236
R21286 OUT2.n145 OUT2.t51 24.9236
R21287 OUT2.n147 OUT2.t32 24.9236
R21288 OUT2.n147 OUT2.t8 24.9236
R21289 OUT2.n94 OUT2.t31 24.9236
R21290 OUT2.n94 OUT2.t60 24.9236
R21291 OUT2.n81 OUT2.t50 24.9236
R21292 OUT2.n81 OUT2.t59 24.9236
R21293 OUT2.n82 OUT2.t2 24.9236
R21294 OUT2.n82 OUT2.t39 24.9236
R21295 OUT2.n84 OUT2.t17 24.9236
R21296 OUT2.n84 OUT2.t53 24.9236
R21297 OUT2.n86 OUT2.t52 24.9236
R21298 OUT2.n86 OUT2.t1 24.9236
R21299 OUT2.n88 OUT2.t9 24.9236
R21300 OUT2.n88 OUT2.t23 24.9236
R21301 OUT2.n90 OUT2.t22 24.9236
R21302 OUT2.n90 OUT2.t41 24.9236
R21303 OUT2.n92 OUT2.t11 24.9236
R21304 OUT2.n92 OUT2.t43 24.9236
R21305 OUT2.n55 OUT2.t37 24.9236
R21306 OUT2.n55 OUT2.t7 24.9236
R21307 OUT2.n42 OUT2.t57 24.9236
R21308 OUT2.n42 OUT2.t5 24.9236
R21309 OUT2.n43 OUT2.t3 24.9236
R21310 OUT2.n43 OUT2.t27 24.9236
R21311 OUT2.n45 OUT2.t24 24.9236
R21312 OUT2.n45 OUT2.t54 24.9236
R21313 OUT2.n47 OUT2.t16 24.9236
R21314 OUT2.n47 OUT2.t48 24.9236
R21315 OUT2.n49 OUT2.t44 24.9236
R21316 OUT2.n49 OUT2.t63 24.9236
R21317 OUT2.n51 OUT2.t61 24.9236
R21318 OUT2.n51 OUT2.t14 24.9236
R21319 OUT2.n53 OUT2.t20 24.9236
R21320 OUT2.n53 OUT2.t33 24.9236
R21321 OUT2.n15 OUT2.t36 24.9236
R21322 OUT2.n15 OUT2.t49 24.9236
R21323 OUT2.n2 OUT2.t55 24.9236
R21324 OUT2.n2 OUT2.t13 24.9236
R21325 OUT2.n3 OUT2.t10 24.9236
R21326 OUT2.n3 OUT2.t25 24.9236
R21327 OUT2.n5 OUT2.t30 24.9236
R21328 OUT2.n5 OUT2.t42 24.9236
R21329 OUT2.n7 OUT2.t47 24.9236
R21330 OUT2.n7 OUT2.t18 24.9236
R21331 OUT2.n9 OUT2.t58 24.9236
R21332 OUT2.n9 OUT2.t29 24.9236
R21333 OUT2.n11 OUT2.t34 24.9236
R21334 OUT2.n11 OUT2.t45 24.9236
R21335 OUT2.n13 OUT2.t28 24.9236
R21336 OUT2.n13 OUT2.t38 24.9236
R21337 OUT2 OUT2.n150 11.4429
R21338 OUT2 OUT2.n95 11.4429
R21339 OUT2 OUT2.n58 11.4429
R21340 OUT2 OUT2.n18 11.4429
R21341 OUT2.n77 OUT2.n62 8.55118
R21342 OUT2.n37 OUT2.n22 8.55118
R21343 OUT2.n114 OUT2.n99 8.55117
R21344 OUT2.n119 OUT2.n118 8.47293
R21345 OUT2.n56 OUT2.n55 7.80093
R21346 OUT2.n16 OUT2.n15 7.80093
R21347 OUT2.n78 OUT2.n77 3.20954
R21348 OUT2.n38 OUT2.n37 3.20953
R21349 OUT2.n115 OUT2.n114 3.20289
R21350 OUT2.n151 OUT2 3.10353
R21351 OUT2.n96 OUT2 3.10353
R21352 OUT2.n59 OUT2 3.10353
R21353 OUT2.n19 OUT2 3.10353
R21354 OUT2.n135 OUT2.n134 3.1005
R21355 OUT2.n57 OUT2.n41 3.1005
R21356 OUT2.n17 OUT2.n1 3.1005
R21357 OUT2.n134 OUT2.n133 2.71565
R21358 OUT2.n114 OUT2.n113 2.13383
R21359 OUT2.n77 OUT2.n76 2.13383
R21360 OUT2.n37 OUT2.n36 2.13383
R21361 OUT2.n150 OUT2 1.74595
R21362 OUT2.n95 OUT2 1.74595
R21363 OUT2.n58 OUT2.n57 1.16414
R21364 OUT2.n18 OUT2.n17 1.16414
R21365 OUT2.n157 OUT2.n156 1.07337
R21366 OUT2.n158 OUT2.n157 0.69375
R21367 OUT2.n159 OUT2.n158 0.68905
R21368 OUT2.n56 OUT2 0.488972
R21369 OUT2.n16 OUT2 0.488972
R21370 OUT2.n158 OUT2.n79 0.414635
R21371 OUT2.n157 OUT2.n116 0.382465
R21372 OUT2.n159 OUT2.n39 0.368576
R21373 OUT2 OUT2.n159 0.281623
R21374 OUT2.n134 OUT2.n119 0.196887
R21375 OUT2.n79 OUT2.n78 0.157252
R21376 OUT2.n39 OUT2.n38 0.139891
R21377 OUT2.n156 OUT2.n155 0.139389
R21378 OUT2.n116 OUT2.n115 0.132946
R21379 OUT2.n60 OUT2.n41 0.113
R21380 OUT2.n20 OUT2.n1 0.113
R21381 OUT2.n154 OUT2.n135 0.101889
R21382 OUT2.n57 OUT2.n56 0.0893205
R21383 OUT2.n17 OUT2.n16 0.0893205
R21384 OUT2.n154 OUT2.n152 0.0282778
R21385 OUT2.n135 OUT2.n117 0.0268889
R21386 OUT2.n98 OUT2.n97 0.0213333
R21387 OUT2.n61 OUT2.n60 0.0143889
R21388 OUT2.n21 OUT2.n20 0.0143889
R21389 OUT2.n115 OUT2.n98 0.00100004
R21390 OUT2.n38 OUT2.n21 0.00100004
R21391 OUT2.n78 OUT2.n61 0.00100004
R21392 OUT2.n152 OUT2.n151 0.000513335
R21393 OUT2.n97 OUT2.n96 0.000513335
R21394 OUT2.n60 OUT2.n59 0.000513218
R21395 OUT2.n20 OUT2.n19 0.000513218
R21396 OUT2.n98 OUT2.n80 0.00050517
R21397 OUT2.n154 OUT2.n153 0.000504838
R21398 OUT2.n61 OUT2.n40 0.000504838
R21399 OUT2.n21 OUT2.n0 0.000504838
R21400 OUT2.n155 OUT2.n154 0.000501713
R21401 VFS.n3 VFS 0.239679
R21402 VFS.n4 VFS.t2 0.0274553
R21403 VFS.n0 VFS.t0 0.0274553
R21404 VFS.n1 VFS.n0 0.0274531
R21405 VFS.n2 VFS.n1 0.0274531
R21406 VFS.n6 VFS.n5 0.0274531
R21407 VFS.n5 VFS.n4 0.0274531
R21408 VFS VFS.n6 0.014671
R21409 VFS.n3 VFS.n2 0.011546
R21410 VFS VFS.n3 0.00223611
R21411 VFS.n4 VFS.t5 0.000502142
R21412 VFS.n5 VFS.t3 0.000502142
R21413 VFS.n6 VFS.t7 0.000502142
R21414 VFS.n2 VFS.t1 0.000502142
R21415 VFS.n1 VFS.t4 0.000502142
R21416 VFS.n0 VFS.t6 0.000502142
R21417 VV16.n0 VV16.t17 167.365
R21418 VV16.n0 VV16.t16 92.4496
R21419 VV16.n1 VV16.n0 2.07493
R21420 VV16.n17 VV16 0.8559
R21421 VV16 VV16.n17 0.356917
R21422 VV16.n15 VV16.n14 0.141409
R21423 VV16.n13 VV16.n12 0.141409
R21424 VV16.n11 VV16.n10 0.141409
R21425 VV16.n9 VV16.n8 0.141409
R21426 VV16.n7 VV16.n6 0.141409
R21427 VV16.n5 VV16.n4 0.141409
R21428 VV16.n3 VV16.n2 0.141409
R21429 VV16.n1 VV16 0.12425
R21430 VV16 VV16.n16 0.105614
R21431 VV16 VV16.n1 0.05
R21432 VV16.n17 VV16 0.0193
R21433 VV16.n17 VV16 0.00833333
R21434 VV16.n2 VV16.t7 0.000729415
R21435 VV16.n16 VV16.n15 0.000727273
R21436 VV16.n14 VV16.n13 0.000727273
R21437 VV16.n12 VV16.n11 0.000727273
R21438 VV16.n10 VV16.n9 0.000727273
R21439 VV16.n8 VV16.n7 0.000727273
R21440 VV16.n6 VV16.n5 0.000727273
R21441 VV16.n4 VV16.n3 0.000727273
R21442 VV16.n3 VV16.t10 0.000502142
R21443 VV16.n5 VV16.t3 0.000502142
R21444 VV16.n7 VV16.t2 0.000502142
R21445 VV16.n9 VV16.t4 0.000502142
R21446 VV16.n11 VV16.t8 0.000502142
R21447 VV16.n13 VV16.t11 0.000502142
R21448 VV16.n15 VV16.t15 0.000502142
R21449 VV16.n16 VV16.t0 0.000502142
R21450 VV16.n14 VV16.t13 0.000502142
R21451 VV16.n12 VV16.t9 0.000502142
R21452 VV16.n10 VV16.t1 0.000502142
R21453 VV16.n8 VV16.t14 0.000502142
R21454 VV16.n6 VV16.t6 0.000502142
R21455 VV16.n4 VV16.t12 0.000502142
R21456 VV16.n2 VV16.t5 0.000502142
R21457 a_16599_n13205.n12 a_16599_n13205.t21 182.77
R21458 a_16599_n13205.n13 a_16599_n13205.t14 182.77
R21459 a_16599_n13205.n14 a_16599_n13205.t6 182.77
R21460 a_16599_n13205.n15 a_16599_n13205.t10 182.77
R21461 a_16599_n13205.n16 a_16599_n13205.t18 182.77
R21462 a_16599_n13205.n17 a_16599_n13205.t4 182.77
R21463 a_16599_n13205.n18 a_16599_n13205.t19 182.77
R21464 a_16599_n13205.n19 a_16599_n13205.t9 182.77
R21465 a_16599_n13205.n20 a_16599_n13205.t5 182.77
R21466 a_16599_n13205.n21 a_16599_n13205.t2 182.77
R21467 a_16599_n13205.n2 a_16599_n13205.t8 182.77
R21468 a_16599_n13205.n3 a_16599_n13205.t23 182.77
R21469 a_16599_n13205.n4 a_16599_n13205.t12 182.77
R21470 a_16599_n13205.n5 a_16599_n13205.t20 182.77
R21471 a_16599_n13205.n6 a_16599_n13205.t13 182.77
R21472 a_16599_n13205.n7 a_16599_n13205.t7 182.77
R21473 a_16599_n13205.n8 a_16599_n13205.t22 182.77
R21474 a_16599_n13205.n9 a_16599_n13205.t11 182.77
R21475 a_16599_n13205.n10 a_16599_n13205.t16 182.77
R21476 a_16599_n13205.n11 a_16599_n13205.t17 90.7933
R21477 a_16599_n13205.n1 a_16599_n13205.t15 90.7875
R21478 a_16599_n13205.n43 a_16599_n13205.t0 42.4202
R21479 a_16599_n13205.n0 a_16599_n13205.t3 4.35105
R21480 a_16599_n13205.t1 a_16599_n13205.n43 2.70045
R21481 a_16599_n13205.n2 a_16599_n13205.n1 2.03273
R21482 a_16599_n13205.n12 a_16599_n13205.n11 2.02124
R21483 a_16599_n13205.n41 a_16599_n13205.n40 0.835222
R21484 a_16599_n13205.n40 a_16599_n13205.n39 0.835222
R21485 a_16599_n13205.n39 a_16599_n13205.n38 0.835222
R21486 a_16599_n13205.n38 a_16599_n13205.n37 0.835222
R21487 a_16599_n13205.n37 a_16599_n13205.n36 0.835222
R21488 a_16599_n13205.n36 a_16599_n13205.n35 0.835222
R21489 a_16599_n13205.n35 a_16599_n13205.n34 0.835222
R21490 a_16599_n13205.n34 a_16599_n13205.n33 0.835222
R21491 a_16599_n13205.n33 a_16599_n13205.n32 0.835222
R21492 a_16599_n13205.n13 a_16599_n13205.n12 0.835222
R21493 a_16599_n13205.n14 a_16599_n13205.n13 0.835222
R21494 a_16599_n13205.n15 a_16599_n13205.n14 0.835222
R21495 a_16599_n13205.n16 a_16599_n13205.n15 0.835222
R21496 a_16599_n13205.n17 a_16599_n13205.n16 0.835222
R21497 a_16599_n13205.n18 a_16599_n13205.n17 0.835222
R21498 a_16599_n13205.n19 a_16599_n13205.n18 0.835222
R21499 a_16599_n13205.n20 a_16599_n13205.n19 0.835222
R21500 a_16599_n13205.n21 a_16599_n13205.n20 0.835222
R21501 a_16599_n13205.n10 a_16599_n13205.n9 0.835222
R21502 a_16599_n13205.n9 a_16599_n13205.n8 0.835222
R21503 a_16599_n13205.n8 a_16599_n13205.n7 0.835222
R21504 a_16599_n13205.n7 a_16599_n13205.n6 0.835222
R21505 a_16599_n13205.n6 a_16599_n13205.n5 0.835222
R21506 a_16599_n13205.n5 a_16599_n13205.n4 0.835222
R21507 a_16599_n13205.n4 a_16599_n13205.n3 0.835222
R21508 a_16599_n13205.n3 a_16599_n13205.n2 0.835222
R21509 a_16599_n13205.n24 a_16599_n13205.n23 0.835222
R21510 a_16599_n13205.n25 a_16599_n13205.n24 0.835222
R21511 a_16599_n13205.n26 a_16599_n13205.n25 0.835222
R21512 a_16599_n13205.n27 a_16599_n13205.n26 0.835222
R21513 a_16599_n13205.n28 a_16599_n13205.n27 0.835222
R21514 a_16599_n13205.n29 a_16599_n13205.n28 0.835222
R21515 a_16599_n13205.n30 a_16599_n13205.n29 0.835222
R21516 a_16599_n13205.n31 a_16599_n13205.n30 0.835222
R21517 a_16599_n13205.n0 a_16599_n13205.n42 0.750184
R21518 a_16599_n13205.n0 a_16599_n13205.n22 0.715064
R21519 a_16599_n13205.n22 a_16599_n13205.n10 0.553972
R21520 a_16599_n13205.n42 a_16599_n13205.n31 0.553972
R21521 a_16599_n13205.n43 a_16599_n13205.n0 0.403234
R21522 a_16599_n13205.n42 a_16599_n13205.n41 0.233139
R21523 a_16599_n13205.n22 a_16599_n13205.n21 0.233139
R21524 a_16541_n13117.n0 a_16541_n13117.t8 5.73525
R21525 a_16541_n13117.n18 a_16541_n13117.t20 5.34571
R21526 a_16541_n13117.n0 a_16541_n13117.t3 5.18362
R21527 a_16541_n13117.n1 a_16541_n13117.t14 5.18362
R21528 a_16541_n13117.n2 a_16541_n13117.t11 5.18362
R21529 a_16541_n13117.n3 a_16541_n13117.t17 5.18362
R21530 a_16541_n13117.n4 a_16541_n13117.t10 5.18362
R21531 a_16541_n13117.n5 a_16541_n13117.t4 5.18362
R21532 a_16541_n13117.n6 a_16541_n13117.t15 5.18362
R21533 a_16541_n13117.n7 a_16541_n13117.t12 5.18362
R21534 a_16541_n13117.n8 a_16541_n13117.t21 5.18362
R21535 a_16541_n13117.n9 a_16541_n13117.t6 5.18362
R21536 a_16541_n13117.n10 a_16541_n13117.t2 5.18362
R21537 a_16541_n13117.n11 a_16541_n13117.t18 5.18362
R21538 a_16541_n13117.n12 a_16541_n13117.t7 5.18362
R21539 a_16541_n13117.n13 a_16541_n13117.t19 5.18362
R21540 a_16541_n13117.n14 a_16541_n13117.t13 5.18362
R21541 a_16541_n13117.n15 a_16541_n13117.t5 5.18362
R21542 a_16541_n13117.n16 a_16541_n13117.t9 5.18362
R21543 a_16541_n13117.n17 a_16541_n13117.t16 5.18362
R21544 a_16541_n13117.t0 a_16541_n13117.n19 2.79552
R21545 a_16541_n13117.n19 a_16541_n13117.t1 2.38201
R21546 a_16541_n13117.n9 a_16541_n13117.n8 1.10376
R21547 a_16541_n13117.n1 a_16541_n13117.n0 0.55213
R21548 a_16541_n13117.n2 a_16541_n13117.n1 0.55213
R21549 a_16541_n13117.n3 a_16541_n13117.n2 0.55213
R21550 a_16541_n13117.n4 a_16541_n13117.n3 0.55213
R21551 a_16541_n13117.n5 a_16541_n13117.n4 0.55213
R21552 a_16541_n13117.n6 a_16541_n13117.n5 0.55213
R21553 a_16541_n13117.n7 a_16541_n13117.n6 0.55213
R21554 a_16541_n13117.n8 a_16541_n13117.n7 0.55213
R21555 a_16541_n13117.n10 a_16541_n13117.n9 0.55213
R21556 a_16541_n13117.n11 a_16541_n13117.n10 0.55213
R21557 a_16541_n13117.n12 a_16541_n13117.n11 0.55213
R21558 a_16541_n13117.n13 a_16541_n13117.n12 0.55213
R21559 a_16541_n13117.n14 a_16541_n13117.n13 0.55213
R21560 a_16541_n13117.n15 a_16541_n13117.n14 0.55213
R21561 a_16541_n13117.n16 a_16541_n13117.n15 0.55213
R21562 a_16541_n13117.n17 a_16541_n13117.n16 0.512683
R21563 a_16541_n13117.n19 a_16541_n13117.n18 0.168655
R21564 a_16541_n13117.n18 a_16541_n13117.n17 0.0581389
R21565 a_16719_n13117.n15 a_16719_n13117.t24 473.437
R21566 a_16719_n13117.n19 a_16719_n13117.t25 473.332
R21567 a_16719_n13117.n0 a_16719_n13117.t0 473.329
R21568 a_16719_n13117.n18 a_16719_n13117.t2 140.444
R21569 a_16719_n13117.n18 a_16719_n13117.t3 41.6504
R21570 a_16719_n13117.n2 a_16719_n13117.t12 5.95597
R21571 a_16719_n13117.n26 a_16719_n13117.t10 5.95597
R21572 a_16719_n13117.n8 a_16719_n13117.t5 5.32159
R21573 a_16719_n13117.n7 a_16719_n13117.t20 5.32159
R21574 a_16719_n13117.n6 a_16719_n13117.t14 5.32159
R21575 a_16719_n13117.n5 a_16719_n13117.t7 5.32159
R21576 a_16719_n13117.n4 a_16719_n13117.t15 5.32159
R21577 a_16719_n13117.n3 a_16719_n13117.t4 5.32159
R21578 a_16719_n13117.n2 a_16719_n13117.t19 5.32159
R21579 a_16719_n13117.n1 a_16719_n13117.t11 5.32159
R21580 a_16719_n13117.n11 a_16719_n13117.t16 5.32159
R21581 a_16719_n13117.n26 a_16719_n13117.t6 5.32159
R21582 a_16719_n13117.n27 a_16719_n13117.t13 5.32159
R21583 a_16719_n13117.n28 a_16719_n13117.t21 5.32159
R21584 a_16719_n13117.n29 a_16719_n13117.t17 5.32159
R21585 a_16719_n13117.n30 a_16719_n13117.t9 5.32159
R21586 a_16719_n13117.n25 a_16719_n13117.t8 5.32159
R21587 a_16719_n13117.n24 a_16719_n13117.t18 5.32159
R21588 a_16719_n13117.n23 a_16719_n13117.t22 5.32159
R21589 a_16719_n13117.t23 a_16719_n13117.n31 5.32059
R21590 a_16719_n13117.n14 a_16719_n13117.n13 2.75606
R21591 a_16719_n13117.n17 a_16719_n13117.n14 2.75328
R21592 a_16719_n13117.n14 a_16719_n13117.t1 1.50409
R21593 a_16719_n13117.n19 a_16719_n13117.n18 1.23545
R21594 a_16719_n13117.n23 a_16719_n13117.n22 1.02772
R21595 a_16719_n13117.n3 a_16719_n13117.n2 0.634875
R21596 a_16719_n13117.n4 a_16719_n13117.n3 0.634875
R21597 a_16719_n13117.n5 a_16719_n13117.n4 0.634875
R21598 a_16719_n13117.n6 a_16719_n13117.n5 0.634875
R21599 a_16719_n13117.n7 a_16719_n13117.n6 0.634875
R21600 a_16719_n13117.n8 a_16719_n13117.n7 0.634875
R21601 a_16719_n13117.n24 a_16719_n13117.n23 0.634875
R21602 a_16719_n13117.n25 a_16719_n13117.n24 0.634875
R21603 a_16719_n13117.n31 a_16719_n13117.n25 0.634875
R21604 a_16719_n13117.n31 a_16719_n13117.n30 0.634875
R21605 a_16719_n13117.n30 a_16719_n13117.n29 0.634875
R21606 a_16719_n13117.n29 a_16719_n13117.n28 0.634875
R21607 a_16719_n13117.n28 a_16719_n13117.n27 0.634875
R21608 a_16719_n13117.n27 a_16719_n13117.n26 0.634875
R21609 a_16719_n13117.n0 a_16719_n13117.n21 0.376529
R21610 a_16719_n13117.n16 a_16719_n13117.n15 0.271346
R21611 a_16719_n13117.n21 a_16719_n13117.n20 0.253053
R21612 a_16719_n13117.n9 a_16719_n13117.n8 0.202227
R21613 a_16719_n13117.n20 a_16719_n13117.n19 0.124538
R21614 a_16719_n13117.n17 a_16719_n13117.n16 0.119076
R21615 a_16719_n13117.n13 a_16719_n13117.n12 0.113872
R21616 a_16719_n13117.n0 a_16719_n13117.n17 0.10111
R21617 a_16719_n13117.n1 a_16719_n13117.n0 0.0537895
R21618 a_16719_n13117.n10 a_16719_n13117.n9 0.0386579
R21619 a_16719_n13117.n22 a_16719_n13117.n1 0.0360263
R21620 a_16719_n13117.n0 a_16719_n13117.n11 0.035794
R21621 a_16719_n13117.n11 a_16719_n13117.n10 0.0202368
R21622 CLK.t85 CLK.t89 344.122
R21623 CLK.t72 CLK.t34 344.122
R21624 CLK.t60 CLK.t16 344.122
R21625 CLK.t7 CLK.t57 344.122
R21626 CLK.t87 CLK.t36 344.122
R21627 CLK.t28 CLK.t80 344.122
R21628 CLK.t13 CLK.t70 344.122
R21629 CLK.t51 CLK.t6 344.122
R21630 CLK.t39 CLK.t95 344.122
R21631 CLK.t74 CLK.t71 344.122
R21632 CLK.t64 CLK.t18 344.122
R21633 CLK.t47 CLK.t5 344.122
R21634 CLK.t90 CLK.t38 344.122
R21635 CLK.t73 CLK.t27 344.122
R21636 CLK.t14 CLK.t63 344.122
R21637 CLK.t48 CLK.t46 344.122
R21638 CLK.n1 CLK.t50 232.299
R21639 CLK.n114 CLK.t42 232.299
R21640 CLK.n106 CLK.t84 232.299
R21641 CLK.n98 CLK.t67 232.299
R21642 CLK.n90 CLK.t52 232.299
R21643 CLK.n82 CLK.t1 232.299
R21644 CLK.n74 CLK.t75 232.299
R21645 CLK.n66 CLK.t21 232.299
R21646 CLK.n58 CLK.t3 232.299
R21647 CLK.n50 CLK.t43 232.299
R21648 CLK.n42 CLK.t31 232.299
R21649 CLK.n34 CLK.t68 232.299
R21650 CLK.n26 CLK.t55 232.299
R21651 CLK.n18 CLK.t93 232.299
R21652 CLK.n10 CLK.t77 232.299
R21653 CLK.n137 CLK.t22 232.299
R21654 CLK.n5 CLK.t94 182.915
R21655 CLK.n118 CLK.t81 182.915
R21656 CLK.n110 CLK.t61 182.915
R21657 CLK.n102 CLK.t8 182.915
R21658 CLK.n94 CLK.t88 182.915
R21659 CLK.n86 CLK.t29 182.915
R21660 CLK.n78 CLK.t19 182.915
R21661 CLK.n70 CLK.t53 182.915
R21662 CLK.n62 CLK.t40 182.915
R21663 CLK.n54 CLK.t76 182.915
R21664 CLK.n46 CLK.t65 182.915
R21665 CLK.n38 CLK.t10 182.915
R21666 CLK.n30 CLK.t91 182.915
R21667 CLK.n22 CLK.t32 182.915
R21668 CLK.n14 CLK.t15 182.915
R21669 CLK.n140 CLK.t49 182.915
R21670 CLK.n5 CLK.t85 182.91
R21671 CLK.n118 CLK.t72 182.91
R21672 CLK.n110 CLK.t60 182.91
R21673 CLK.n102 CLK.t7 182.91
R21674 CLK.n94 CLK.t87 182.91
R21675 CLK.n86 CLK.t28 182.91
R21676 CLK.n78 CLK.t13 182.91
R21677 CLK.n70 CLK.t51 182.91
R21678 CLK.n62 CLK.t39 182.91
R21679 CLK.n54 CLK.t74 182.91
R21680 CLK.n46 CLK.t64 182.91
R21681 CLK.n38 CLK.t47 182.91
R21682 CLK.n30 CLK.t90 182.91
R21683 CLK.n22 CLK.t73 182.91
R21684 CLK.n14 CLK.t14 182.91
R21685 CLK.n140 CLK.t48 182.91
R21686 CLK.t94 CLK.n4 182.769
R21687 CLK.t81 CLK.n117 182.769
R21688 CLK.t61 CLK.n109 182.769
R21689 CLK.t8 CLK.n101 182.769
R21690 CLK.t88 CLK.n93 182.769
R21691 CLK.t29 CLK.n85 182.769
R21692 CLK.t19 CLK.n77 182.769
R21693 CLK.t53 CLK.n69 182.769
R21694 CLK.t40 CLK.n61 182.769
R21695 CLK.t76 CLK.n53 182.769
R21696 CLK.t65 CLK.n45 182.769
R21697 CLK.t10 CLK.n37 182.769
R21698 CLK.t91 CLK.n29 182.769
R21699 CLK.t32 CLK.n21 182.769
R21700 CLK.t15 CLK.n13 182.769
R21701 CLK.t49 CLK.n139 182.769
R21702 CLK.n2 CLK.t26 161.262
R21703 CLK.n115 CLK.t59 161.262
R21704 CLK.n107 CLK.t37 161.262
R21705 CLK.n99 CLK.t82 161.262
R21706 CLK.n91 CLK.t62 161.262
R21707 CLK.n83 CLK.t9 161.262
R21708 CLK.n75 CLK.t0 161.262
R21709 CLK.n67 CLK.t30 161.262
R21710 CLK.n59 CLK.t20 161.262
R21711 CLK.n51 CLK.t54 161.262
R21712 CLK.n43 CLK.t41 161.262
R21713 CLK.n35 CLK.t83 161.262
R21714 CLK.n27 CLK.t66 161.262
R21715 CLK.n19 CLK.t11 161.262
R21716 CLK.n11 CLK.t92 161.262
R21717 CLK.n135 CLK.t86 161.262
R21718 CLK.n6 CLK.t23 159.958
R21719 CLK.n119 CLK.t24 159.958
R21720 CLK.n111 CLK.t12 159.958
R21721 CLK.n103 CLK.t44 159.958
R21722 CLK.n95 CLK.t33 159.958
R21723 CLK.n87 CLK.t69 159.958
R21724 CLK.n79 CLK.t56 159.958
R21725 CLK.n71 CLK.t2 159.958
R21726 CLK.n63 CLK.t79 159.958
R21727 CLK.n55 CLK.t25 159.958
R21728 CLK.n47 CLK.t4 159.958
R21729 CLK.n39 CLK.t45 159.958
R21730 CLK.n31 CLK.t35 159.958
R21731 CLK.n23 CLK.t17 159.958
R21732 CLK.n15 CLK.t58 159.958
R21733 CLK.n141 CLK.t78 159.958
R21734 CLK.n121 CLK 4.70942
R21735 CLK.n3 CLK.n2 4.5005
R21736 CLK.n116 CLK.n115 4.5005
R21737 CLK.n108 CLK.n107 4.5005
R21738 CLK.n100 CLK.n99 4.5005
R21739 CLK.n92 CLK.n91 4.5005
R21740 CLK.n84 CLK.n83 4.5005
R21741 CLK.n76 CLK.n75 4.5005
R21742 CLK.n68 CLK.n67 4.5005
R21743 CLK.n60 CLK.n59 4.5005
R21744 CLK.n52 CLK.n51 4.5005
R21745 CLK.n44 CLK.n43 4.5005
R21746 CLK.n36 CLK.n35 4.5005
R21747 CLK.n28 CLK.n27 4.5005
R21748 CLK.n20 CLK.n19 4.5005
R21749 CLK.n12 CLK.n11 4.5005
R21750 CLK.n122 CLK 4.19834
R21751 CLK.n124 CLK 4.19834
R21752 CLK.n127 CLK 4.19834
R21753 CLK.n123 CLK 4.18793
R21754 CLK.n126 CLK 4.18793
R21755 CLK.n125 CLK 4.17751
R21756 CLK.n132 CLK 4.17751
R21757 CLK.n128 CLK 4.16709
R21758 CLK.n129 CLK 4.16709
R21759 CLK.n131 CLK 4.16709
R21760 CLK.n133 CLK 4.16709
R21761 CLK CLK.n134 4.16709
R21762 CLK.n8 CLK 4.15668
R21763 CLK.n121 CLK 4.14654
R21764 CLK.n130 CLK 4.12571
R21765 CLK.n8 CLK 0.757091
R21766 CLK.n128 CLK.n127 0.620955
R21767 CLK.n125 CLK.n124 0.618682
R21768 CLK.n134 CLK.n8 0.616409
R21769 CLK.n133 CLK.n132 0.616409
R21770 CLK.n130 CLK.n129 0.616409
R21771 CLK.n123 CLK.n122 0.616409
R21772 CLK.n134 CLK.n133 0.614136
R21773 CLK.n129 CLK.n128 0.614136
R21774 CLK.n132 CLK.n131 0.611864
R21775 CLK.n131 CLK.n130 0.611864
R21776 CLK.n127 CLK.n126 0.611864
R21777 CLK.n126 CLK.n125 0.611864
R21778 CLK.n124 CLK.n123 0.611864
R21779 CLK.n122 CLK.n121 0.609591
R21780 CLK.n6 CLK.n5 0.56781
R21781 CLK.n119 CLK.n118 0.56781
R21782 CLK.n111 CLK.n110 0.56781
R21783 CLK.n103 CLK.n102 0.56781
R21784 CLK.n95 CLK.n94 0.56781
R21785 CLK.n87 CLK.n86 0.56781
R21786 CLK.n79 CLK.n78 0.56781
R21787 CLK.n71 CLK.n70 0.56781
R21788 CLK.n63 CLK.n62 0.56781
R21789 CLK.n55 CLK.n54 0.56781
R21790 CLK.n47 CLK.n46 0.56781
R21791 CLK.n39 CLK.n38 0.56781
R21792 CLK.n31 CLK.n30 0.56781
R21793 CLK.n23 CLK.n22 0.56781
R21794 CLK.n15 CLK.n14 0.56781
R21795 CLK.n141 CLK.n140 0.56781
R21796 CLK.n7 CLK.n6 0.428385
R21797 CLK.n120 CLK.n119 0.428385
R21798 CLK.n112 CLK.n111 0.428385
R21799 CLK.n104 CLK.n103 0.428385
R21800 CLK.n96 CLK.n95 0.428385
R21801 CLK.n88 CLK.n87 0.428385
R21802 CLK.n80 CLK.n79 0.428385
R21803 CLK.n72 CLK.n71 0.428385
R21804 CLK.n64 CLK.n63 0.428385
R21805 CLK.n56 CLK.n55 0.428385
R21806 CLK.n48 CLK.n47 0.428385
R21807 CLK.n40 CLK.n39 0.428385
R21808 CLK.n32 CLK.n31 0.428385
R21809 CLK.n24 CLK.n23 0.428385
R21810 CLK.n16 CLK.n15 0.428385
R21811 CLK.n142 CLK.n141 0.428385
R21812 CLK.n7 CLK 0.0573182
R21813 CLK.n104 CLK 0.0573182
R21814 CLK.n96 CLK 0.0573182
R21815 CLK.n88 CLK 0.0573182
R21816 CLK.n80 CLK 0.0573182
R21817 CLK.n72 CLK 0.0573182
R21818 CLK.n64 CLK 0.0573182
R21819 CLK.n56 CLK 0.0573182
R21820 CLK.n48 CLK 0.0573182
R21821 CLK.n32 CLK 0.0573182
R21822 CLK.n24 CLK 0.0573182
R21823 CLK.n16 CLK 0.0573182
R21824 CLK.n142 CLK 0.0573182
R21825 CLK.n120 CLK 0.0525833
R21826 CLK.n112 CLK 0.0525833
R21827 CLK.n40 CLK 0.0525833
R21828 CLK CLK.n7 0.0436818
R21829 CLK CLK.n104 0.0436818
R21830 CLK CLK.n96 0.0436818
R21831 CLK CLK.n88 0.0436818
R21832 CLK CLK.n80 0.0436818
R21833 CLK CLK.n72 0.0436818
R21834 CLK CLK.n64 0.0436818
R21835 CLK CLK.n56 0.0436818
R21836 CLK CLK.n48 0.0436818
R21837 CLK CLK.n32 0.0436818
R21838 CLK CLK.n24 0.0436818
R21839 CLK CLK.n16 0.0436818
R21840 CLK CLK.n142 0.0436818
R21841 CLK CLK.n120 0.0400833
R21842 CLK CLK.n112 0.0400833
R21843 CLK CLK.n40 0.0400833
R21844 CLK.n1 CLK.n0 0.0211923
R21845 CLK.n114 CLK.n113 0.0211923
R21846 CLK.n106 CLK.n105 0.0211923
R21847 CLK.n98 CLK.n97 0.0211923
R21848 CLK.n90 CLK.n89 0.0211923
R21849 CLK.n82 CLK.n81 0.0211923
R21850 CLK.n74 CLK.n73 0.0211923
R21851 CLK.n66 CLK.n65 0.0211923
R21852 CLK.n58 CLK.n57 0.0211923
R21853 CLK.n50 CLK.n49 0.0211923
R21854 CLK.n42 CLK.n41 0.0211923
R21855 CLK.n34 CLK.n33 0.0211923
R21856 CLK.n26 CLK.n25 0.0211923
R21857 CLK.n18 CLK.n17 0.0211923
R21858 CLK.n10 CLK.n9 0.0211923
R21859 CLK.n2 CLK.n0 0.0178077
R21860 CLK.n115 CLK.n113 0.0178077
R21861 CLK.n107 CLK.n105 0.0178077
R21862 CLK.n99 CLK.n97 0.0178077
R21863 CLK.n91 CLK.n89 0.0178077
R21864 CLK.n83 CLK.n81 0.0178077
R21865 CLK.n75 CLK.n73 0.0178077
R21866 CLK.n67 CLK.n65 0.0178077
R21867 CLK.n59 CLK.n57 0.0178077
R21868 CLK.n51 CLK.n49 0.0178077
R21869 CLK.n43 CLK.n41 0.0178077
R21870 CLK.n35 CLK.n33 0.0178077
R21871 CLK.n27 CLK.n25 0.0178077
R21872 CLK.n19 CLK.n17 0.0178077
R21873 CLK.n11 CLK.n9 0.0178077
R21874 CLK.n136 CLK.n135 0.0178077
R21875 CLK.n4 CLK.n0 0.00531334
R21876 CLK.n117 CLK.n113 0.00531334
R21877 CLK.n109 CLK.n105 0.00531334
R21878 CLK.n101 CLK.n97 0.00531334
R21879 CLK.n93 CLK.n89 0.00531334
R21880 CLK.n85 CLK.n81 0.00531334
R21881 CLK.n77 CLK.n73 0.00531334
R21882 CLK.n69 CLK.n65 0.00531334
R21883 CLK.n61 CLK.n57 0.00531334
R21884 CLK.n53 CLK.n49 0.00531334
R21885 CLK.n45 CLK.n41 0.00531334
R21886 CLK.n37 CLK.n33 0.00531334
R21887 CLK.n29 CLK.n25 0.00531334
R21888 CLK.n21 CLK.n17 0.00531334
R21889 CLK.n13 CLK.n9 0.00531334
R21890 CLK.n139 CLK.n136 0.00531334
R21891 CLK.n4 CLK.n3 0.00224847
R21892 CLK.n117 CLK.n116 0.00224847
R21893 CLK.n109 CLK.n108 0.00224847
R21894 CLK.n101 CLK.n100 0.00224847
R21895 CLK.n93 CLK.n92 0.00224847
R21896 CLK.n85 CLK.n84 0.00224847
R21897 CLK.n77 CLK.n76 0.00224847
R21898 CLK.n69 CLK.n68 0.00224847
R21899 CLK.n61 CLK.n60 0.00224847
R21900 CLK.n53 CLK.n52 0.00224847
R21901 CLK.n45 CLK.n44 0.00224847
R21902 CLK.n37 CLK.n36 0.00224847
R21903 CLK.n29 CLK.n28 0.00224847
R21904 CLK.n21 CLK.n20 0.00224847
R21905 CLK.n13 CLK.n12 0.00224847
R21906 CLK.n139 CLK.n138 0.00224847
R21907 CLK.n3 CLK.n1 0.00100535
R21908 CLK.n116 CLK.n114 0.00100535
R21909 CLK.n108 CLK.n106 0.00100535
R21910 CLK.n100 CLK.n98 0.00100535
R21911 CLK.n92 CLK.n90 0.00100535
R21912 CLK.n84 CLK.n82 0.00100535
R21913 CLK.n76 CLK.n74 0.00100535
R21914 CLK.n68 CLK.n66 0.00100535
R21915 CLK.n60 CLK.n58 0.00100535
R21916 CLK.n52 CLK.n50 0.00100535
R21917 CLK.n44 CLK.n42 0.00100535
R21918 CLK.n36 CLK.n34 0.00100535
R21919 CLK.n28 CLK.n26 0.00100535
R21920 CLK.n20 CLK.n18 0.00100535
R21921 CLK.n12 CLK.n10 0.00100535
R21922 CLK.n138 CLK.n137 0.00100535
R21923 frontAnalog_v0p0p1_10.x65.A.n1 frontAnalog_v0p0p1_10.x65.A.t4 260.322
R21924 frontAnalog_v0p0p1_10.x65.A.n3 frontAnalog_v0p0p1_10.x65.A.t7 233.929
R21925 frontAnalog_v0p0p1_10.x65.A.n1 frontAnalog_v0p0p1_10.x65.A.t6 175.169
R21926 frontAnalog_v0p0p1_10.x65.A.n2 frontAnalog_v0p0p1_10.x65.A.t5 160.416
R21927 frontAnalog_v0p0p1_10.x65.A.n4 frontAnalog_v0p0p1_10.x65.A.t1 17.4109
R21928 frontAnalog_v0p0p1_10.x65.A.n4 frontAnalog_v0p0p1_10.x65.A.t0 10.2053
R21929 frontAnalog_v0p0p1_10.x65.A.n0 frontAnalog_v0p0p1_10.x65.A 2.78715
R21930 frontAnalog_v0p0p1_10.x65.A.n0 frontAnalog_v0p0p1_10.x65.A.n1 9.09103
R21931 frontAnalog_v0p0p1_10.x65.A.n6 frontAnalog_v0p0p1_10.x65.A.t2 7.94569
R21932 frontAnalog_v0p0p1_10.x65.A.n2 frontAnalog_v0p0p1_10.x65.A.t3 7.55846
R21933 frontAnalog_v0p0p1_10.x65.A.n5 frontAnalog_v0p0p1_10.x65.A.n3 1.4614
R21934 frontAnalog_v0p0p1_10.x65.A.n3 frontAnalog_v0p0p1_10.x65.A.n2 1.19626
R21935 frontAnalog_v0p0p1_10.x65.A.n6 frontAnalog_v0p0p1_10.x65.A.n5 0.836961
R21936 frontAnalog_v0p0p1_10.x65.A frontAnalog_v0p0p1_10.x65.A.n0 0.390342
R21937 frontAnalog_v0p0p1_10.x65.A.n5 frontAnalog_v0p0p1_10.x65.A.n4 0.154668
R21938 frontAnalog_v0p0p1_10.x65.A frontAnalog_v0p0p1_10.x65.A.n6 0.08175
R21939 VV4.n0 VV4.t17 167.365
R21940 VV4.n0 VV4.t16 92.4488
R21941 VV4.n1 VV4.n0 2.07493
R21942 VV4.n10 VV4 0.572333
R21943 VV4 VV4.n10 0.429375
R21944 VV4.n9 VV4.n8 0.141636
R21945 VV4.n8 VV4.n7 0.141636
R21946 VV4.n7 VV4.n6 0.141636
R21947 VV4.n6 VV4.n5 0.141636
R21948 VV4.n5 VV4.n4 0.141636
R21949 VV4.n4 VV4.n3 0.141636
R21950 VV4.n3 VV4.n2 0.141636
R21951 VV4.n1 VV4 0.12425
R21952 VV4 VV4.n9 0.103284
R21953 VV4 VV4.n1 0.0314375
R21954 VV4.n10 VV4 0.00833333
R21955 VV4.n10 VV4 0.006375
R21956 VV4.n3 VV4.t13 0.000502142
R21957 VV4.n4 VV4.t5 0.000502142
R21958 VV4.n5 VV4.t1 0.000502142
R21959 VV4.n6 VV4.t9 0.000502142
R21960 VV4.n7 VV4.t2 0.000502142
R21961 VV4.n8 VV4.t7 0.000502142
R21962 VV4.n9 VV4.t0 0.000502142
R21963 VV4.n2 VV4.t12 0.000502142
R21964 VV4.n3 VV4.t14 0.000502142
R21965 VV4.n4 VV4.t4 0.000502142
R21966 VV4.n5 VV4.t15 0.000502142
R21967 VV4.n6 VV4.t6 0.000502142
R21968 VV4.n7 VV4.t11 0.000502142
R21969 VV4.n8 VV4.t3 0.000502142
R21970 VV4.n9 VV4.t10 0.000502142
R21971 VV4.n2 VV4.t8 0.000502142
R21972 VV3.n0 VV3.t17 167.365
R21973 VV3.n0 VV3.t16 92.4488
R21974 VV3.n1 VV3.n0 2.07493
R21975 VV3.n17 VV3 0.607583
R21976 VV3 VV3.n17 0.455812
R21977 VV3.n15 VV3.n14 0.141409
R21978 VV3.n13 VV3.n12 0.141409
R21979 VV3.n11 VV3.n10 0.141409
R21980 VV3.n9 VV3.n8 0.141409
R21981 VV3.n7 VV3.n6 0.141409
R21982 VV3.n5 VV3.n4 0.141409
R21983 VV3.n3 VV3.n2 0.141409
R21984 VV3.n1 VV3 0.12425
R21985 VV3 VV3.n16 0.100973
R21986 VV3 VV3.n1 0.0314375
R21987 VV3.n17 VV3 0.00833333
R21988 VV3.n17 VV3 0.006375
R21989 VV3.n2 VV3.t13 0.000729415
R21990 VV3.n16 VV3.n15 0.000727273
R21991 VV3.n14 VV3.n13 0.000727273
R21992 VV3.n12 VV3.n11 0.000727273
R21993 VV3.n10 VV3.n9 0.000727273
R21994 VV3.n8 VV3.n7 0.000727273
R21995 VV3.n6 VV3.n5 0.000727273
R21996 VV3.n4 VV3.n3 0.000727273
R21997 VV3.n3 VV3.t14 0.000502142
R21998 VV3.n5 VV3.t5 0.000502142
R21999 VV3.n7 VV3.t15 0.000502142
R22000 VV3.n9 VV3.t9 0.000502142
R22001 VV3.n11 VV3.t12 0.000502142
R22002 VV3.n13 VV3.t3 0.000502142
R22003 VV3.n15 VV3.t11 0.000502142
R22004 VV3.n2 VV3.t6 0.000502142
R22005 VV3.n4 VV3.t1 0.000502142
R22006 VV3.n6 VV3.t0 0.000502142
R22007 VV3.n8 VV3.t4 0.000502142
R22008 VV3.n10 VV3.t8 0.000502142
R22009 VV3.n12 VV3.t2 0.000502142
R22010 VV3.n14 VV3.t10 0.000502142
R22011 VV3.n16 VV3.t7 0.000502142
R22012 frontAnalog_v0p0p1_14.x63.A.n2 frontAnalog_v0p0p1_14.x63.A.t7 260.322
R22013 frontAnalog_v0p0p1_14.x63.A.n4 frontAnalog_v0p0p1_14.x63.A.t4 233.888
R22014 frontAnalog_v0p0p1_14.x63.A.n2 frontAnalog_v0p0p1_14.x63.A.t5 175.169
R22015 frontAnalog_v0p0p1_14.x63.A.n3 frontAnalog_v0p0p1_14.x63.A.t6 159.725
R22016 frontAnalog_v0p0p1_14.x63.A.n1 frontAnalog_v0p0p1_14.x63.A.t2 17.4109
R22017 frontAnalog_v0p0p1_14.x63.A.n0 frontAnalog_v0p0p1_14.x63.A.n2 9.75129
R22018 frontAnalog_v0p0p1_14.x63.A.n1 frontAnalog_v0p0p1_14.x63.A.t3 9.6037
R22019 frontAnalog_v0p0p1_14.x63.A.n0 frontAnalog_v0p0p1_14.x63.A 2.33338
R22020 frontAnalog_v0p0p1_14.x63.A.n5 frontAnalog_v0p0p1_14.x63.A.t0 8.40929
R22021 frontAnalog_v0p0p1_14.x63.A.n3 frontAnalog_v0p0p1_14.x63.A.t1 8.06629
R22022 frontAnalog_v0p0p1_14.x63.A.n4 frontAnalog_v0p0p1_14.x63.A.n3 1.73501
R22023 frontAnalog_v0p0p1_14.x63.A.n1 frontAnalog_v0p0p1_14.x63.A.n4 0.99025
R22024 frontAnalog_v0p0p1_14.x63.A.n5 frontAnalog_v0p0p1_14.x63.A.n1 0.853186
R22025 frontAnalog_v0p0p1_14.x63.A frontAnalog_v0p0p1_14.x63.A.n0 0.349517
R22026 frontAnalog_v0p0p1_14.x63.A frontAnalog_v0p0p1_14.x63.A.n5 0.24425
R22027 frontAnalog_v0p0p1_14.x65.A.n1 frontAnalog_v0p0p1_14.x65.A.t7 260.322
R22028 frontAnalog_v0p0p1_14.x65.A.n3 frontAnalog_v0p0p1_14.x65.A.t5 233.929
R22029 frontAnalog_v0p0p1_14.x65.A.n1 frontAnalog_v0p0p1_14.x65.A.t4 175.169
R22030 frontAnalog_v0p0p1_14.x65.A.n2 frontAnalog_v0p0p1_14.x65.A.t6 160.416
R22031 frontAnalog_v0p0p1_14.x65.A.n4 frontAnalog_v0p0p1_14.x65.A.t2 17.4109
R22032 frontAnalog_v0p0p1_14.x65.A.n4 frontAnalog_v0p0p1_14.x65.A.t3 10.2053
R22033 frontAnalog_v0p0p1_14.x65.A.n0 frontAnalog_v0p0p1_14.x65.A 2.78715
R22034 frontAnalog_v0p0p1_14.x65.A.n0 frontAnalog_v0p0p1_14.x65.A.n1 9.09103
R22035 frontAnalog_v0p0p1_14.x65.A.n6 frontAnalog_v0p0p1_14.x65.A.t0 7.94569
R22036 frontAnalog_v0p0p1_14.x65.A.n2 frontAnalog_v0p0p1_14.x65.A.t1 7.55846
R22037 frontAnalog_v0p0p1_14.x65.A.n5 frontAnalog_v0p0p1_14.x65.A.n3 1.4614
R22038 frontAnalog_v0p0p1_14.x65.A.n3 frontAnalog_v0p0p1_14.x65.A.n2 1.19626
R22039 frontAnalog_v0p0p1_14.x65.A.n6 frontAnalog_v0p0p1_14.x65.A.n5 0.836961
R22040 frontAnalog_v0p0p1_14.x65.A frontAnalog_v0p0p1_14.x65.A.n0 0.390342
R22041 frontAnalog_v0p0p1_14.x65.A.n5 frontAnalog_v0p0p1_14.x65.A.n4 0.154668
R22042 frontAnalog_v0p0p1_14.x65.A frontAnalog_v0p0p1_14.x65.A.n6 0.08175
R22043 frontAnalog_v0p0p1_5.RSfetsym_0.QN.n1 frontAnalog_v0p0p1_5.RSfetsym_0.QN.t6 117.511
R22044 frontAnalog_v0p0p1_5.RSfetsym_0.QN.n1 frontAnalog_v0p0p1_5.RSfetsym_0.QN.t5 110.698
R22045 frontAnalog_v0p0p1_5.RSfetsym_0.QN.n2 frontAnalog_v0p0p1_5.RSfetsym_0.QN.t2 19.1963
R22046 frontAnalog_v0p0p1_5.RSfetsym_0.QN.n3 frontAnalog_v0p0p1_5.RSfetsym_0.QN.t1 14.5206
R22047 frontAnalog_v0p0p1_5.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_5.RSfetsym_0.QN.t4 14.283
R22048 frontAnalog_v0p0p1_5.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_5.RSfetsym_0.QN.t3 14.283
R22049 frontAnalog_v0p0p1_5.RSfetsym_0.QN frontAnalog_v0p0p1_5.RSfetsym_0.QN.t0 9.14075
R22050 frontAnalog_v0p0p1_5.RSfetsym_0.QN.n2 frontAnalog_v0p0p1_5.RSfetsym_0.QN.n1 0.826818
R22051 frontAnalog_v0p0p1_5.RSfetsym_0.QN frontAnalog_v0p0p1_5.RSfetsym_0.QN.n0 0.74645
R22052 frontAnalog_v0p0p1_5.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_5.RSfetsym_0.QN.n3 0.249509
R22053 frontAnalog_v0p0p1_5.RSfetsym_0.QN.n3 frontAnalog_v0p0p1_5.RSfetsym_0.QN.n2 0.0968646
R22054 VV11.n0 VV11.t17 167.365
R22055 VV11.n0 VV11.t16 92.4496
R22056 VV11.n1 VV11.n0 2.07493
R22057 VV11.n17 VV11 0.5175
R22058 VV11 VV11.n17 0.38825
R22059 VV11.n15 VV11.n14 0.141409
R22060 VV11.n13 VV11.n12 0.141409
R22061 VV11.n11 VV11.n10 0.141409
R22062 VV11.n9 VV11.n8 0.141409
R22063 VV11.n7 VV11.n6 0.141409
R22064 VV11.n5 VV11.n4 0.141409
R22065 VV11.n3 VV11.n2 0.141409
R22066 VV11.n1 VV11 0.12425
R22067 VV11 VV11.n16 0.104098
R22068 VV11 VV11.n1 0.0314375
R22069 VV11.n17 VV11 0.00833333
R22070 VV11.n17 VV11 0.006375
R22071 VV11.n2 VV11.t9 0.000729415
R22072 VV11.n16 VV11.n15 0.000727273
R22073 VV11.n14 VV11.n13 0.000727273
R22074 VV11.n12 VV11.n11 0.000727273
R22075 VV11.n10 VV11.n9 0.000727273
R22076 VV11.n8 VV11.n7 0.000727273
R22077 VV11.n6 VV11.n5 0.000727273
R22078 VV11.n4 VV11.n3 0.000727273
R22079 VV11.n3 VV11.t10 0.000502142
R22080 VV11.n5 VV11.t15 0.000502142
R22081 VV11.n7 VV11.t2 0.000502142
R22082 VV11.n9 VV11.t6 0.000502142
R22083 VV11.n11 VV11.t13 0.000502142
R22084 VV11.n13 VV11.t11 0.000502142
R22085 VV11.n15 VV11.t3 0.000502142
R22086 VV11.n16 VV11.t1 0.000502142
R22087 VV11.n14 VV11.t14 0.000502142
R22088 VV11.n12 VV11.t5 0.000502142
R22089 VV11.n10 VV11.t8 0.000502142
R22090 VV11.n8 VV11.t4 0.000502142
R22091 VV11.n6 VV11.t0 0.000502142
R22092 VV11.n4 VV11.t12 0.000502142
R22093 VV11.n2 VV11.t7 0.000502142
R22094 VV10.n0 VV10.t16 167.365
R22095 VV10.n0 VV10.t17 92.4496
R22096 VV10.n1 VV10.n0 2.07493
R22097 VV10.n10 VV10 0.474417
R22098 VV10 VV10.n10 0.355937
R22099 VV10.n9 VV10.n8 0.141636
R22100 VV10.n8 VV10.n7 0.141636
R22101 VV10.n7 VV10.n6 0.141636
R22102 VV10.n6 VV10.n5 0.141636
R22103 VV10.n5 VV10.n4 0.141636
R22104 VV10.n4 VV10.n3 0.141636
R22105 VV10.n3 VV10.n2 0.141636
R22106 VV10.n1 VV10 0.12425
R22107 VV10 VV10.n9 0.104326
R22108 VV10 VV10.n1 0.028
R22109 VV10.n10 VV10 0.00833333
R22110 VV10.n10 VV10 0.006375
R22111 VV10.n2 VV10.t8 0.000502142
R22112 VV10.n3 VV10.t7 0.000502142
R22113 VV10.n4 VV10.t0 0.000502142
R22114 VV10.n5 VV10.t13 0.000502142
R22115 VV10.n6 VV10.t6 0.000502142
R22116 VV10.n7 VV10.t4 0.000502142
R22117 VV10.n8 VV10.t9 0.000502142
R22118 VV10.n9 VV10.t5 0.000502142
R22119 VV10.n9 VV10.t2 0.000502142
R22120 VV10.n8 VV10.t12 0.000502142
R22121 VV10.n7 VV10.t14 0.000502142
R22122 VV10.n6 VV10.t3 0.000502142
R22123 VV10.n5 VV10.t1 0.000502142
R22124 VV10.n4 VV10.t15 0.000502142
R22125 VV10.n3 VV10.t11 0.000502142
R22126 VV10.n2 VV10.t10 0.000502142
R22127 VV2.n0 VV2.t16 167.365
R22128 VV2.n0 VV2.t17 92.4488
R22129 VV2.n1 VV2.n0 2.07493
R22130 VV2.n17 VV2 0.64675
R22131 VV2 VV2.n17 0.485188
R22132 VV2.n15 VV2.n14 0.141409
R22133 VV2.n13 VV2.n12 0.141409
R22134 VV2.n11 VV2.n10 0.141409
R22135 VV2.n9 VV2.n8 0.141409
R22136 VV2.n7 VV2.n6 0.141409
R22137 VV2.n5 VV2.n4 0.141409
R22138 VV2.n3 VV2.n2 0.141409
R22139 VV2.n1 VV2 0.12425
R22140 VV2 VV2.n16 0.0968068
R22141 VV2 VV2.n1 0.028
R22142 VV2.n17 VV2 0.00833333
R22143 VV2.n17 VV2 0.006375
R22144 VV2.n2 VV2.t10 0.000729415
R22145 VV2.n16 VV2.n15 0.000727273
R22146 VV2.n14 VV2.n13 0.000727273
R22147 VV2.n12 VV2.n11 0.000727273
R22148 VV2.n10 VV2.n9 0.000727273
R22149 VV2.n8 VV2.n7 0.000727273
R22150 VV2.n6 VV2.n5 0.000727273
R22151 VV2.n4 VV2.n3 0.000727273
R22152 VV2.n4 VV2.t1 0.000502142
R22153 VV2.n6 VV2.t0 0.000502142
R22154 VV2.n8 VV2.t4 0.000502142
R22155 VV2.n10 VV2.t8 0.000502142
R22156 VV2.n12 VV2.t3 0.000502142
R22157 VV2.n14 VV2.t9 0.000502142
R22158 VV2.n16 VV2.t7 0.000502142
R22159 VV2.n3 VV2.t11 0.000502142
R22160 VV2.n5 VV2.t14 0.000502142
R22161 VV2.n7 VV2.t2 0.000502142
R22162 VV2.n9 VV2.t13 0.000502142
R22163 VV2.n11 VV2.t15 0.000502142
R22164 VV2.n13 VV2.t12 0.000502142
R22165 VV2.n15 VV2.t5 0.000502142
R22166 VV2.n2 VV2.t6 0.000502142
R22167 VV1.n0 VV1.t17 167.365
R22168 VV1.n0 VV1.t16 92.4488
R22169 VV1.n1 VV1.n0 2.07493
R22170 VV1.n10 VV1 0.8277
R22171 VV1 VV1.n10 0.591357
R22172 VV1.n9 VV1.n8 0.141636
R22173 VV1.n8 VV1.n7 0.141636
R22174 VV1.n7 VV1.n6 0.141636
R22175 VV1.n6 VV1.n5 0.141636
R22176 VV1.n5 VV1.n4 0.141636
R22177 VV1.n4 VV1.n3 0.141636
R22178 VV1.n3 VV1.n2 0.141636
R22179 VV1.n1 VV1 0.12425
R22180 VV1 VV1.n9 0.0980758
R22181 VV1 VV1.n1 0.0314375
R22182 VV1.n10 VV1 0.0099
R22183 VV1.n10 VV1 0.00721429
R22184 VV1.n3 VV1.t10 0.000502142
R22185 VV1.n4 VV1.t13 0.000502142
R22186 VV1.n5 VV1.t0 0.000502142
R22187 VV1.n6 VV1.t12 0.000502142
R22188 VV1.n7 VV1.t15 0.000502142
R22189 VV1.n8 VV1.t11 0.000502142
R22190 VV1.n9 VV1.t2 0.000502142
R22191 VV1.n2 VV1.t4 0.000502142
R22192 VV1.n3 VV1.t1 0.000502142
R22193 VV1.n4 VV1.t6 0.000502142
R22194 VV1.n5 VV1.t5 0.000502142
R22195 VV1.n6 VV1.t14 0.000502142
R22196 VV1.n7 VV1.t9 0.000502142
R22197 VV1.n8 VV1.t3 0.000502142
R22198 VV1.n9 VV1.t8 0.000502142
R22199 VV1.n2 VV1.t7 0.000502142
R22200 I0.n0 I0.t5 196.549
R22201 I0.n0 I0.t7 148.35
R22202 I0.n4 I0.t8 117.314
R22203 I0.n4 I0.t6 110.853
R22204 I0.n6 I0.t3 17.6181
R22205 I0.n7 I0.t1 14.2865
R22206 I0.n9 I0.t2 14.283
R22207 I0.n9 I0.t0 14.283
R22208 I0 I0.n12 9.77614
R22209 I0.n1 I0.n0 9.49592
R22210 I0.n11 I0.t4 8.77744
R22211 I0.n2 I0.n1 7.58085
R22212 I0.n1 I0 6.44187
R22213 I0.n3 I0.n2 2.50858
R22214 I0.n11 I0.n10 1.20426
R22215 I0.n2 I0 0.88934
R22216 I0.n12 I0.n11 0.32511
R22217 I0.n7 I0.n6 0.314673
R22218 I0.n8 I0.n7 0.299251
R22219 I0.n13 I0 0.204167
R22220 I0.n3 I0 0.2005
R22221 I0 I0.n3 0.1932
R22222 I0.n5 I0.n4 0.159555
R22223 I0 I0.n13 0.15325
R22224 I0.n10 I0.n9 0.106617
R22225 I0.n8 I0.n5 0.0796167
R22226 I0.n10 I0.n8 0.0480595
R22227 I0.n12 I0 0.046937
R22228 I0.n13 I0 0.0161667
R22229 I0.n13 I0 0.01225
R22230 I0.n6 I0.n5 0.000504658
R22231 R1 R1.t1 451.853
R22232 R1.n45 R1.t1 440.25
R22233 R1.n0 R1.t4 258.584
R22234 R1.n38 R1.t8 258.58
R22235 R1.n11 R1.t2 212.081
R22236 R1.n5 R1.t3 212.081
R22237 R1.n4 R1.t7 212.081
R22238 R1.n24 R1.t9 212.081
R22239 R1.n11 R1.t11 139.78
R22240 R1.n5 R1.t12 139.78
R22241 R1.n4 R1.t5 139.78
R22242 R1.n24 R1.t6 139.78
R22243 R1 R1.t0 126.855
R22244 R1.n34 R1.t10 110.734
R22245 R1.n46 R1.n45 50.2399
R22246 R1.n26 R1.n24 30.6732
R22247 R1.n6 R1.n4 30.6732
R22248 R1.n6 R1.n5 30.6732
R22249 R1.n12 R1.n11 30.6732
R22250 R1.n46 R1 25.4148
R22251 R1.n23 R1.n22 12.8005
R22252 R1.n26 R1.n25 12.4157
R22253 R1.n18 R1.n17 9.3005
R22254 R1.n32 R1.n31 9.3005
R22255 R1.n13 R1.n12 8.28655
R22256 R1.n21 R1.n6 8.28655
R22257 R1.n27 R1.n26 8.28655
R22258 R1.n22 R1.n21 4.3525
R22259 R1.n14 R1.n9 4.3525
R22260 R1.n10 R1 4.10569
R22261 R1.n28 R1.n3 4.0965
R22262 R1.n20 R1 3.8405
R22263 R1.n45 R1 2.84494
R22264 R1 R1.n1 2.3045
R22265 R1.n31 R1 2.3045
R22266 R1.n27 R1 2.3045
R22267 R1 R1.n23 2.0485
R22268 R1 R1.n46 1.94081
R22269 R1.n43 R1.n33 1.59023
R22270 R1.n13 R1.n10 1.15386
R22271 R1.n28 R1.n27 1.0245
R22272 R1.n17 R1 0.7685
R22273 R1.n21 R1.n20 0.5125
R22274 R1.n14 R1.n13 0.5125
R22275 R1.n33 R1.n1 0.462934
R22276 R1.n44 R1.n43 0.44229
R22277 R1.n44 R1.n0 0.179314
R22278 R1.n43 R1.n42 0.14376
R22279 R1.n7 R1.n2 0.105187
R22280 R1.n32 R1.n30 0.084875
R22281 R1.n18 R1.n16 0.0708125
R22282 R1.n47 R1.n44 0.0699392
R22283 R1.n42 R1.n41 0.0475
R22284 R1.n19 R1.n18 0.028625
R22285 R1.n8 R1.n7 0.0270625
R22286 R1.n16 R1.n15 0.0270625
R22287 R1.n30 R1.n29 0.0255
R22288 R1.n47 R1 0.0251063
R22289 R1.n33 R1.n32 0.0239512
R22290 R1.n36 R1.n35 0.0174119
R22291 R1.n37 R1.n34 0.0133182
R22292 R1 R1.n47 0.00738976
R22293 R1.n29 R1.n2 0.00675
R22294 R1.n19 R1.n8 0.003625
R22295 R1.n41 R1.n37 0.00263636
R22296 R1.n39 R1.n38 0.0020625
R22297 R1.n29 R1.n28 0.00119114
R22298 R1.n20 R1.n19 0.00119114
R22299 R1.n15 R1.n14 0.00119114
R22300 R1.n37 R1.n36 0.000747155
R22301 R1.n41 R1.n40 0.000588765
R22302 R1.n40 R1.n39 0.000588763
R22303 I2.n6 I2.t5 323.342
R22304 I2.n0 I2.t9 228.927
R22305 I2.n3 I2.t7 196.549
R22306 I2.n6 I2.t8 194.809
R22307 I2.n0 I2.t6 159.391
R22308 I2.n3 I2.t11 148.35
R22309 I2.n10 I2.t12 117.314
R22310 I2.n10 I2.t10 110.853
R22311 I2.n7 I2.n6 76.0005
R22312 I2.n4 I2.n3 76.0005
R22313 I2.n8 I2.n7 29.2624
R22314 I2.n12 I2.t0 17.6181
R22315 I2.n13 I2.t3 14.2865
R22316 I2.n15 I2.t1 14.283
R22317 I2.n15 I2.t2 14.283
R22318 I2.n5 I2 9.11
R22319 I2.n17 I2.t4 8.77744
R22320 I2.n1 I2.n0 8.68501
R22321 I2 I2.n18 7.11948
R22322 I2.n4 I2 5.78114
R22323 I2.n2 I2.n1 4.26764
R22324 I2 I2.n4 3.71663
R22325 I2.n1 I2 1.99697
R22326 I2.n7 I2 1.92927
R22327 I2.n8 I2.n5 1.79514
R22328 I2.n17 I2.n16 1.20426
R22329 I2.n5 I2.n2 0.570143
R22330 I2.n19 I2 0.360833
R22331 I2 I2.n9 0.349867
R22332 I2.n18 I2.n17 0.32511
R22333 I2.n13 I2.n12 0.314673
R22334 I2.n14 I2.n13 0.299251
R22335 I2 I2.n19 0.27075
R22336 I2.n9 I2.n8 0.226885
R22337 I2.n2 I2 0.221483
R22338 I2.n9 I2 0.20675
R22339 I2.n11 I2.n10 0.159555
R22340 I2.n16 I2.n15 0.106617
R22341 I2.n14 I2.n11 0.0796167
R22342 I2.n16 I2.n14 0.0480595
R22343 I2.n18 I2 0.046937
R22344 I2.n19 I2 0.0161667
R22345 I2.n19 I2 0.01225
R22346 I2.n12 I2.n11 0.000504658
R22347 OUT1.n122 OUT1.n120 145.809
R22348 OUT1.n65 OUT1.n63 145.809
R22349 OUT1.n25 OUT1.n23 145.809
R22350 OUT1.n102 OUT1.n100 145.808
R22351 OUT1.n65 OUT1.n64 107.409
R22352 OUT1.n67 OUT1.n66 107.409
R22353 OUT1.n69 OUT1.n68 107.409
R22354 OUT1.n71 OUT1.n70 107.409
R22355 OUT1.n73 OUT1.n72 107.409
R22356 OUT1.n75 OUT1.n74 107.409
R22357 OUT1.n25 OUT1.n24 107.409
R22358 OUT1.n27 OUT1.n26 107.409
R22359 OUT1.n29 OUT1.n28 107.409
R22360 OUT1.n31 OUT1.n30 107.409
R22361 OUT1.n33 OUT1.n32 107.409
R22362 OUT1.n35 OUT1.n34 107.409
R22363 OUT1.n122 OUT1.n121 107.407
R22364 OUT1.n124 OUT1.n123 107.407
R22365 OUT1.n126 OUT1.n125 107.407
R22366 OUT1.n128 OUT1.n127 107.407
R22367 OUT1.n130 OUT1.n129 107.407
R22368 OUT1.n132 OUT1.n131 107.407
R22369 OUT1.n102 OUT1.n101 107.407
R22370 OUT1.n104 OUT1.n103 107.407
R22371 OUT1.n106 OUT1.n105 107.407
R22372 OUT1.n108 OUT1.n107 107.407
R22373 OUT1.n110 OUT1.n109 107.407
R22374 OUT1.n112 OUT1.n111 107.407
R22375 OUT1.n138 OUT1.n136 87.1779
R22376 OUT1.n83 OUT1.n81 87.1779
R22377 OUT1.n44 OUT1.n42 87.1779
R22378 OUT1.n4 OUT1.n2 87.1779
R22379 OUT1.n54 OUT1.n53 52.82
R22380 OUT1.n14 OUT1.n13 52.82
R22381 OUT1.n138 OUT1.n137 52.82
R22382 OUT1.n140 OUT1.n139 52.82
R22383 OUT1.n142 OUT1.n141 52.82
R22384 OUT1.n144 OUT1.n143 52.82
R22385 OUT1.n146 OUT1.n145 52.82
R22386 OUT1.n148 OUT1.n147 52.82
R22387 OUT1.n83 OUT1.n82 52.82
R22388 OUT1.n85 OUT1.n84 52.82
R22389 OUT1.n87 OUT1.n86 52.82
R22390 OUT1.n89 OUT1.n88 52.82
R22391 OUT1.n91 OUT1.n90 52.82
R22392 OUT1.n93 OUT1.n92 52.82
R22393 OUT1.n44 OUT1.n43 52.82
R22394 OUT1.n46 OUT1.n45 52.82
R22395 OUT1.n48 OUT1.n47 52.82
R22396 OUT1.n50 OUT1.n49 52.82
R22397 OUT1.n52 OUT1.n51 52.82
R22398 OUT1.n4 OUT1.n3 52.82
R22399 OUT1.n6 OUT1.n5 52.82
R22400 OUT1.n8 OUT1.n7 52.82
R22401 OUT1.n10 OUT1.n9 52.82
R22402 OUT1.n12 OUT1.n11 52.82
R22403 OUT1 OUT1.n149 51.0745
R22404 OUT1 OUT1.n94 51.0745
R22405 OUT1.n124 OUT1.n122 38.4005
R22406 OUT1.n126 OUT1.n124 38.4005
R22407 OUT1.n128 OUT1.n126 38.4005
R22408 OUT1.n130 OUT1.n128 38.4005
R22409 OUT1.n132 OUT1.n130 38.4005
R22410 OUT1.n133 OUT1.n132 38.4005
R22411 OUT1.n104 OUT1.n102 38.4005
R22412 OUT1.n106 OUT1.n104 38.4005
R22413 OUT1.n108 OUT1.n106 38.4005
R22414 OUT1.n110 OUT1.n108 38.4005
R22415 OUT1.n112 OUT1.n110 38.4005
R22416 OUT1.n113 OUT1.n112 38.4005
R22417 OUT1.n67 OUT1.n65 38.4005
R22418 OUT1.n69 OUT1.n67 38.4005
R22419 OUT1.n71 OUT1.n69 38.4005
R22420 OUT1.n73 OUT1.n71 38.4005
R22421 OUT1.n75 OUT1.n73 38.4005
R22422 OUT1.n76 OUT1.n75 38.4005
R22423 OUT1.n27 OUT1.n25 38.4005
R22424 OUT1.n29 OUT1.n27 38.4005
R22425 OUT1.n31 OUT1.n29 38.4005
R22426 OUT1.n33 OUT1.n31 38.4005
R22427 OUT1.n35 OUT1.n33 38.4005
R22428 OUT1.n36 OUT1.n35 38.4005
R22429 OUT1.n140 OUT1.n138 34.3584
R22430 OUT1.n142 OUT1.n140 34.3584
R22431 OUT1.n144 OUT1.n142 34.3584
R22432 OUT1.n146 OUT1.n144 34.3584
R22433 OUT1.n148 OUT1.n146 34.3584
R22434 OUT1.n150 OUT1.n148 34.3584
R22435 OUT1.n85 OUT1.n83 34.3584
R22436 OUT1.n87 OUT1.n85 34.3584
R22437 OUT1.n89 OUT1.n87 34.3584
R22438 OUT1.n91 OUT1.n89 34.3584
R22439 OUT1.n93 OUT1.n91 34.3584
R22440 OUT1.n95 OUT1.n93 34.3584
R22441 OUT1.n46 OUT1.n44 34.3584
R22442 OUT1.n48 OUT1.n46 34.3584
R22443 OUT1.n50 OUT1.n48 34.3584
R22444 OUT1.n52 OUT1.n50 34.3584
R22445 OUT1.n54 OUT1.n52 34.3584
R22446 OUT1.n58 OUT1.n54 34.3584
R22447 OUT1.n6 OUT1.n4 34.3584
R22448 OUT1.n8 OUT1.n6 34.3584
R22449 OUT1.n10 OUT1.n8 34.3584
R22450 OUT1.n12 OUT1.n10 34.3584
R22451 OUT1.n14 OUT1.n12 34.3584
R22452 OUT1.n18 OUT1.n14 34.3584
R22453 OUT1.n118 OUT1.t99 26.5955
R22454 OUT1.n118 OUT1.t112 26.5955
R22455 OUT1.n120 OUT1.t97 26.5955
R22456 OUT1.n120 OUT1.t69 26.5955
R22457 OUT1.n121 OUT1.t119 26.5955
R22458 OUT1.n121 OUT1.t85 26.5955
R22459 OUT1.n123 OUT1.t64 26.5955
R22460 OUT1.n123 OUT1.t105 26.5955
R22461 OUT1.n125 OUT1.t75 26.5955
R22462 OUT1.n125 OUT1.t93 26.5955
R22463 OUT1.n127 OUT1.t91 26.5955
R22464 OUT1.n127 OUT1.t108 26.5955
R22465 OUT1.n129 OUT1.t114 26.5955
R22466 OUT1.n129 OUT1.t80 26.5955
R22467 OUT1.n131 OUT1.t125 26.5955
R22468 OUT1.n131 OUT1.t101 26.5955
R22469 OUT1.n99 OUT1.t124 26.5955
R22470 OUT1.n99 OUT1.t89 26.5955
R22471 OUT1.n100 OUT1.t79 26.5955
R22472 OUT1.n100 OUT1.t88 26.5955
R22473 OUT1.n101 OUT1.t95 26.5955
R22474 OUT1.n101 OUT1.t68 26.5955
R22475 OUT1.n103 OUT1.t110 26.5955
R22476 OUT1.n103 OUT1.t82 26.5955
R22477 OUT1.n105 OUT1.t81 26.5955
R22478 OUT1.n105 OUT1.t94 26.5955
R22479 OUT1.n107 OUT1.t102 26.5955
R22480 OUT1.n107 OUT1.t116 26.5955
R22481 OUT1.n109 OUT1.t115 26.5955
R22482 OUT1.n109 OUT1.t70 26.5955
R22483 OUT1.n111 OUT1.t104 26.5955
R22484 OUT1.n111 OUT1.t72 26.5955
R22485 OUT1.n62 OUT1.t66 26.5955
R22486 OUT1.n62 OUT1.t100 26.5955
R22487 OUT1.n63 OUT1.t86 26.5955
R22488 OUT1.n63 OUT1.t98 26.5955
R22489 OUT1.n64 OUT1.t96 26.5955
R22490 OUT1.n64 OUT1.t120 26.5955
R22491 OUT1.n66 OUT1.t117 26.5955
R22492 OUT1.n66 OUT1.t83 26.5955
R22493 OUT1.n68 OUT1.t109 26.5955
R22494 OUT1.n68 OUT1.t76 26.5955
R22495 OUT1.n70 OUT1.t74 26.5955
R22496 OUT1.n70 OUT1.t92 26.5955
R22497 OUT1.n72 OUT1.t90 26.5955
R22498 OUT1.n72 OUT1.t107 26.5955
R22499 OUT1.n74 OUT1.t113 26.5955
R22500 OUT1.n74 OUT1.t126 26.5955
R22501 OUT1.n22 OUT1.t65 26.5955
R22502 OUT1.n22 OUT1.t78 26.5955
R22503 OUT1.n23 OUT1.t84 26.5955
R22504 OUT1.n23 OUT1.t106 26.5955
R22505 OUT1.n24 OUT1.t103 26.5955
R22506 OUT1.n24 OUT1.t118 26.5955
R22507 OUT1.n26 OUT1.t123 26.5955
R22508 OUT1.n26 OUT1.t71 26.5955
R22509 OUT1.n28 OUT1.t77 26.5955
R22510 OUT1.n28 OUT1.t111 26.5955
R22511 OUT1.n30 OUT1.t87 26.5955
R22512 OUT1.n30 OUT1.t122 26.5955
R22513 OUT1.n32 OUT1.t127 26.5955
R22514 OUT1.n32 OUT1.t73 26.5955
R22515 OUT1.n34 OUT1.t121 26.5955
R22516 OUT1.n34 OUT1.t67 26.5955
R22517 OUT1.n149 OUT1.t46 24.9236
R22518 OUT1.n149 OUT1.t59 24.9236
R22519 OUT1.n136 OUT1.t44 24.9236
R22520 OUT1.n136 OUT1.t16 24.9236
R22521 OUT1.n137 OUT1.t2 24.9236
R22522 OUT1.n137 OUT1.t32 24.9236
R22523 OUT1.n139 OUT1.t11 24.9236
R22524 OUT1.n139 OUT1.t52 24.9236
R22525 OUT1.n141 OUT1.t22 24.9236
R22526 OUT1.n141 OUT1.t40 24.9236
R22527 OUT1.n143 OUT1.t38 24.9236
R22528 OUT1.n143 OUT1.t55 24.9236
R22529 OUT1.n145 OUT1.t61 24.9236
R22530 OUT1.n145 OUT1.t27 24.9236
R22531 OUT1.n147 OUT1.t8 24.9236
R22532 OUT1.n147 OUT1.t48 24.9236
R22533 OUT1.n94 OUT1.t7 24.9236
R22534 OUT1.n94 OUT1.t36 24.9236
R22535 OUT1.n81 OUT1.t26 24.9236
R22536 OUT1.n81 OUT1.t35 24.9236
R22537 OUT1.n82 OUT1.t42 24.9236
R22538 OUT1.n82 OUT1.t15 24.9236
R22539 OUT1.n84 OUT1.t57 24.9236
R22540 OUT1.n84 OUT1.t29 24.9236
R22541 OUT1.n86 OUT1.t28 24.9236
R22542 OUT1.n86 OUT1.t41 24.9236
R22543 OUT1.n88 OUT1.t49 24.9236
R22544 OUT1.n88 OUT1.t63 24.9236
R22545 OUT1.n90 OUT1.t62 24.9236
R22546 OUT1.n90 OUT1.t17 24.9236
R22547 OUT1.n92 OUT1.t51 24.9236
R22548 OUT1.n92 OUT1.t19 24.9236
R22549 OUT1.n55 OUT1.t13 24.9236
R22550 OUT1.n55 OUT1.t47 24.9236
R22551 OUT1.n42 OUT1.t33 24.9236
R22552 OUT1.n42 OUT1.t45 24.9236
R22553 OUT1.n43 OUT1.t43 24.9236
R22554 OUT1.n43 OUT1.t3 24.9236
R22555 OUT1.n45 OUT1.t0 24.9236
R22556 OUT1.n45 OUT1.t30 24.9236
R22557 OUT1.n47 OUT1.t56 24.9236
R22558 OUT1.n47 OUT1.t24 24.9236
R22559 OUT1.n49 OUT1.t20 24.9236
R22560 OUT1.n49 OUT1.t39 24.9236
R22561 OUT1.n51 OUT1.t37 24.9236
R22562 OUT1.n51 OUT1.t54 24.9236
R22563 OUT1.n53 OUT1.t60 24.9236
R22564 OUT1.n53 OUT1.t9 24.9236
R22565 OUT1.n15 OUT1.t12 24.9236
R22566 OUT1.n15 OUT1.t25 24.9236
R22567 OUT1.n2 OUT1.t31 24.9236
R22568 OUT1.n2 OUT1.t53 24.9236
R22569 OUT1.n3 OUT1.t50 24.9236
R22570 OUT1.n3 OUT1.t1 24.9236
R22571 OUT1.n5 OUT1.t6 24.9236
R22572 OUT1.n5 OUT1.t18 24.9236
R22573 OUT1.n7 OUT1.t23 24.9236
R22574 OUT1.n7 OUT1.t58 24.9236
R22575 OUT1.n9 OUT1.t34 24.9236
R22576 OUT1.n9 OUT1.t5 24.9236
R22577 OUT1.n11 OUT1.t10 24.9236
R22578 OUT1.n11 OUT1.t21 24.9236
R22579 OUT1.n13 OUT1.t4 24.9236
R22580 OUT1.n13 OUT1.t14 24.9236
R22581 OUT1 OUT1.n150 11.4429
R22582 OUT1 OUT1.n95 11.4429
R22583 OUT1 OUT1.n58 11.4429
R22584 OUT1 OUT1.n18 11.4429
R22585 OUT1.n77 OUT1.n62 8.55024
R22586 OUT1.n37 OUT1.n22 8.55024
R22587 OUT1.n114 OUT1.n99 8.55024
R22588 OUT1.n119 OUT1.n118 8.46262
R22589 OUT1.n56 OUT1.n55 7.77479
R22590 OUT1.n16 OUT1.n15 7.77479
R22591 OUT1.n135 OUT1.n134 4.6505
R22592 OUT1.n151 OUT1 3.29747
R22593 OUT1.n96 OUT1 3.29747
R22594 OUT1.n78 OUT1.n77 3.20821
R22595 OUT1.n38 OUT1.n37 3.2082
R22596 OUT1.n115 OUT1.n114 3.20156
R22597 OUT1.n59 OUT1 3.10353
R22598 OUT1.n19 OUT1 3.10353
R22599 OUT1.n57 OUT1.n41 3.1005
R22600 OUT1.n17 OUT1.n1 3.1005
R22601 OUT1.n134 OUT1.n133 2.71565
R22602 OUT1.n114 OUT1.n113 2.32777
R22603 OUT1.n77 OUT1.n76 2.32777
R22604 OUT1.n37 OUT1.n36 2.32777
R22605 OUT1.n150 OUT1 1.74595
R22606 OUT1.n95 OUT1 1.74595
R22607 OUT1.n157 OUT1.n156 1.07337
R22608 OUT1.n58 OUT1.n57 0.970197
R22609 OUT1.n18 OUT1.n17 0.970197
R22610 OUT1.n158 OUT1.n157 0.69375
R22611 OUT1.n159 OUT1.n158 0.68905
R22612 OUT1.n56 OUT1 0.649449
R22613 OUT1.n16 OUT1 0.649449
R22614 OUT1.n158 OUT1.n79 0.414635
R22615 OUT1.n157 OUT1.n116 0.382465
R22616 OUT1.n159 OUT1.n39 0.368576
R22617 OUT1 OUT1.n159 0.279743
R22618 OUT1.n134 OUT1.n119 0.207197
R22619 OUT1.n79 OUT1.n78 0.157252
R22620 OUT1.n39 OUT1.n38 0.139891
R22621 OUT1.n156 OUT1.n155 0.139389
R22622 OUT1.n116 OUT1.n115 0.132946
R22623 OUT1.n57 OUT1.n56 0.118507
R22624 OUT1.n17 OUT1.n16 0.118507
R22625 OUT1.n60 OUT1.n41 0.111611
R22626 OUT1.n20 OUT1.n1 0.111611
R22627 OUT1.n154 OUT1.n135 0.0991111
R22628 OUT1.n154 OUT1.n152 0.0296667
R22629 OUT1.n135 OUT1.n117 0.0282778
R22630 OUT1.n98 OUT1.n97 0.0227222
R22631 OUT1.n61 OUT1.n60 0.0171667
R22632 OUT1.n21 OUT1.n20 0.0171667
R22633 OUT1.n115 OUT1.n98 0.00100004
R22634 OUT1.n38 OUT1.n21 0.00100004
R22635 OUT1.n78 OUT1.n61 0.00100004
R22636 OUT1.n152 OUT1.n151 0.000513563
R22637 OUT1.n97 OUT1.n96 0.000513563
R22638 OUT1.n60 OUT1.n59 0.000513218
R22639 OUT1.n20 OUT1.n19 0.000513218
R22640 OUT1.n98 OUT1.n80 0.00050517
R22641 OUT1.n154 OUT1.n153 0.000504838
R22642 OUT1.n61 OUT1.n40 0.000504838
R22643 OUT1.n21 OUT1.n0 0.000504838
R22644 OUT1.n155 OUT1.n154 0.000501713
R22645 frontAnalog_v0p0p1_8.RSfetsym_0.QN.n1 frontAnalog_v0p0p1_8.RSfetsym_0.QN.t5 117.511
R22646 frontAnalog_v0p0p1_8.RSfetsym_0.QN.n1 frontAnalog_v0p0p1_8.RSfetsym_0.QN.t6 110.698
R22647 frontAnalog_v0p0p1_8.RSfetsym_0.QN.n2 frontAnalog_v0p0p1_8.RSfetsym_0.QN.t4 19.1963
R22648 frontAnalog_v0p0p1_8.RSfetsym_0.QN.n3 frontAnalog_v0p0p1_8.RSfetsym_0.QN.t0 14.5206
R22649 frontAnalog_v0p0p1_8.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_8.RSfetsym_0.QN.t2 14.283
R22650 frontAnalog_v0p0p1_8.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_8.RSfetsym_0.QN.t3 14.283
R22651 frontAnalog_v0p0p1_8.RSfetsym_0.QN frontAnalog_v0p0p1_8.RSfetsym_0.QN.t1 9.14075
R22652 frontAnalog_v0p0p1_8.RSfetsym_0.QN.n2 frontAnalog_v0p0p1_8.RSfetsym_0.QN.n1 0.826818
R22653 frontAnalog_v0p0p1_8.RSfetsym_0.QN frontAnalog_v0p0p1_8.RSfetsym_0.QN.n0 0.74645
R22654 frontAnalog_v0p0p1_8.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_8.RSfetsym_0.QN.n3 0.249509
R22655 frontAnalog_v0p0p1_8.RSfetsym_0.QN.n3 frontAnalog_v0p0p1_8.RSfetsym_0.QN.n2 0.0968646
R22656 VV9.n0 VV9.t17 167.365
R22657 VV9.n0 VV9.t16 92.4496
R22658 VV9.n1 VV9.n0 2.07493
R22659 VV9.n10 VV9 0.431333
R22660 VV9 VV9.n10 0.287722
R22661 VV9.n9 VV9.n8 0.141636
R22662 VV9.n8 VV9.n7 0.141636
R22663 VV9.n7 VV9.n6 0.141636
R22664 VV9.n6 VV9.n5 0.141636
R22665 VV9.n5 VV9.n4 0.141636
R22666 VV9.n4 VV9.n3 0.141636
R22667 VV9.n3 VV9.n2 0.141636
R22668 VV9.n1 VV9 0.12425
R22669 VV9 VV9.n9 0.102242
R22670 VV9 VV9.n1 0.0314375
R22671 VV9.n10 VV9 0.00833333
R22672 VV9.n10 VV9 0.00572222
R22673 VV9.n2 VV9.t8 0.000502142
R22674 VV9.n3 VV9.t0 0.000502142
R22675 VV9.n4 VV9.t3 0.000502142
R22676 VV9.n5 VV9.t4 0.000502142
R22677 VV9.n6 VV9.t12 0.000502142
R22678 VV9.n7 VV9.t9 0.000502142
R22679 VV9.n8 VV9.t13 0.000502142
R22680 VV9.n9 VV9.t15 0.000502142
R22681 VV9.n9 VV9.t5 0.000502142
R22682 VV9.n8 VV9.t11 0.000502142
R22683 VV9.n7 VV9.t2 0.000502142
R22684 VV9.n6 VV9.t6 0.000502142
R22685 VV9.n5 VV9.t14 0.000502142
R22686 VV9.n4 VV9.t1 0.000502142
R22687 VV9.n3 VV9.t7 0.000502142
R22688 VV9.n2 VV9.t10 0.000502142
R22689 VV15.n0 VV15.t16 167.365
R22690 VV15.n0 VV15.t17 92.4496
R22691 VV15.n1 VV15.n0 2.07493
R22692 VV15.n9 VV15.n8 0.141636
R22693 VV15.n8 VV15.n7 0.141636
R22694 VV15.n7 VV15.n6 0.141636
R22695 VV15.n6 VV15.n5 0.141636
R22696 VV15.n5 VV15.n4 0.141636
R22697 VV15.n4 VV15.n3 0.141636
R22698 VV15.n3 VV15.n2 0.141636
R22699 VV15.n1 VV15 0.12425
R22700 VV15 VV15.n9 0.100159
R22701 VV15 VV15.n1 0.0358571
R22702 VV15.n2 VV15.t1 0.000502142
R22703 VV15.n3 VV15.t15 0.000502142
R22704 VV15.n4 VV15.t11 0.000502142
R22705 VV15.n5 VV15.t13 0.000502142
R22706 VV15.n6 VV15.t6 0.000502142
R22707 VV15.n7 VV15.t5 0.000502142
R22708 VV15.n8 VV15.t4 0.000502142
R22709 VV15.n9 VV15.t10 0.000502142
R22710 VV15.n9 VV15.t14 0.000502142
R22711 VV15.n8 VV15.t12 0.000502142
R22712 VV15.n7 VV15.t8 0.000502142
R22713 VV15.n6 VV15.t3 0.000502142
R22714 VV15.n5 VV15.t0 0.000502142
R22715 VV15.n4 VV15.t2 0.000502142
R22716 VV15.n3 VV15.t9 0.000502142
R22717 VV15.n2 VV15.t7 0.000502142
R22718 frontAnalog_v0p0p1_2.x63.A.n2 frontAnalog_v0p0p1_2.x63.A.t5 260.322
R22719 frontAnalog_v0p0p1_2.x63.A.n4 frontAnalog_v0p0p1_2.x63.A.t4 233.888
R22720 frontAnalog_v0p0p1_2.x63.A.n2 frontAnalog_v0p0p1_2.x63.A.t6 175.169
R22721 frontAnalog_v0p0p1_2.x63.A.n3 frontAnalog_v0p0p1_2.x63.A.t7 159.725
R22722 frontAnalog_v0p0p1_2.x63.A.n1 frontAnalog_v0p0p1_2.x63.A.t0 17.4109
R22723 frontAnalog_v0p0p1_2.x63.A.n0 frontAnalog_v0p0p1_2.x63.A.n2 9.75129
R22724 frontAnalog_v0p0p1_2.x63.A.n1 frontAnalog_v0p0p1_2.x63.A.t1 9.6027
R22725 frontAnalog_v0p0p1_2.x63.A.n0 frontAnalog_v0p0p1_2.x63.A 2.33338
R22726 frontAnalog_v0p0p1_2.x63.A.n5 frontAnalog_v0p0p1_2.x63.A.t2 8.40929
R22727 frontAnalog_v0p0p1_2.x63.A.n3 frontAnalog_v0p0p1_2.x63.A.t3 8.06629
R22728 frontAnalog_v0p0p1_2.x63.A.n4 frontAnalog_v0p0p1_2.x63.A.n3 1.73501
R22729 frontAnalog_v0p0p1_2.x63.A.n1 frontAnalog_v0p0p1_2.x63.A.n4 0.99025
R22730 frontAnalog_v0p0p1_2.x63.A.n5 frontAnalog_v0p0p1_2.x63.A.n1 0.853186
R22731 frontAnalog_v0p0p1_2.x63.A frontAnalog_v0p0p1_2.x63.A.n0 0.349517
R22732 frontAnalog_v0p0p1_2.x63.A frontAnalog_v0p0p1_2.x63.A.n5 0.24425
R22733 frontAnalog_v0p0p1_2.x65.A.n1 frontAnalog_v0p0p1_2.x65.A.t4 260.322
R22734 frontAnalog_v0p0p1_2.x65.A.n4 frontAnalog_v0p0p1_2.x65.A.t6 233.929
R22735 frontAnalog_v0p0p1_2.x65.A.n1 frontAnalog_v0p0p1_2.x65.A.t5 175.169
R22736 frontAnalog_v0p0p1_2.x65.A.n3 frontAnalog_v0p0p1_2.x65.A.t7 160.416
R22737 frontAnalog_v0p0p1_2.x65.A.n2 frontAnalog_v0p0p1_2.x65.A.t3 17.4109
R22738 frontAnalog_v0p0p1_2.x65.A.n2 frontAnalog_v0p0p1_2.x65.A.t2 10.2053
R22739 frontAnalog_v0p0p1_2.x65.A.n0 frontAnalog_v0p0p1_2.x65.A 2.78715
R22740 frontAnalog_v0p0p1_2.x65.A.n0 frontAnalog_v0p0p1_2.x65.A.n1 9.09103
R22741 frontAnalog_v0p0p1_2.x65.A.n6 frontAnalog_v0p0p1_2.x65.A.t1 7.94569
R22742 frontAnalog_v0p0p1_2.x65.A.n3 frontAnalog_v0p0p1_2.x65.A.t0 7.55846
R22743 frontAnalog_v0p0p1_2.x65.A.n5 frontAnalog_v0p0p1_2.x65.A.n4 1.4614
R22744 frontAnalog_v0p0p1_2.x65.A.n4 frontAnalog_v0p0p1_2.x65.A.n3 1.19626
R22745 frontAnalog_v0p0p1_2.x65.A.n6 frontAnalog_v0p0p1_2.x65.A.n5 0.836961
R22746 frontAnalog_v0p0p1_2.x65.A frontAnalog_v0p0p1_2.x65.A.n0 0.390342
R22747 frontAnalog_v0p0p1_2.x65.A.n5 frontAnalog_v0p0p1_2.x65.A.n2 0.154668
R22748 frontAnalog_v0p0p1_2.x65.A frontAnalog_v0p0p1_2.x65.A.n6 0.08175
R22749 S0.n5 S0.t8 259.192
R22750 S0.n39 S0.t2 258.584
R22751 S0.n0 S0.t1 222.243
R22752 S0.n18 S0.t5 212.081
R22753 S0.n17 S0.t6 212.081
R22754 S0.n14 S0.t10 212.081
R22755 S0.n11 S0.t11 212.081
R22756 S0.n13 S0.n10 152
R22757 S0.n18 S0.t7 139.78
R22758 S0.n17 S0.t9 139.78
R22759 S0.n14 S0.t3 139.78
R22760 S0.n11 S0.t4 139.78
R22761 S0.n1 S0.t0 123.654
R22762 S0.n40 S0.t12 117.346
R22763 S0.n11 S0.n6 44.8017
R22764 S0.n2 S0.n1 43.0815
R22765 S0.n2 S0 32.4695
R22766 S0.n12 S0.n11 30.6732
R22767 S0.n15 S0.n14 30.6732
R22768 S0.n17 S0.n15 30.6732
R22769 S0.n19 S0.n17 30.6732
R22770 S0.n19 S0.n18 30.6732
R22771 S0.n14 S0.n13 18.2581
R22772 S0.n36 S0.n35 13.8245
R22773 S0.n30 S0.n10 12.8005
R22774 S0.n13 S0.n12 12.4157
R22775 S0.n25 S0.n24 11.5205
R22776 S0 S0.n0 10.4848
R22777 S0.n37 S0.n36 9.3005
R22778 S0.n35 S0.n7 9.3005
R22779 S0.n31 S0.n30 9.3005
R22780 S0.n26 S0.n25 9.3005
R22781 S0.n24 S0.n16 9.3005
R22782 S0.n29 S0.n15 8.28655
R22783 S0.n20 S0.n19 8.28655
R22784 S0.n12 S0.n8 8.28655
R22785 S0.n0 S0 5.50526
R22786 S0.n1 S0 5.16973
R22787 S0.n32 S0.n8 4.6505
R22788 S0.n29 S0.n9 4.6505
R22789 S0.n30 S0.n29 4.3525
R22790 S0.n24 S0.n23 4.3525
R22791 S0.n21 S0 4.10475
R22792 S0.n35 S0.n34 4.0965
R22793 S0.n28 S0 3.8405
R22794 S0.n22 S0.n21 2.33609
R22795 S0 S0.n6 2.3045
R22796 S0.n36 S0 2.3045
R22797 S0 S0.n8 2.3045
R22798 S0.n10 S0 2.0485
R22799 S0 S0.n2 1.98623
R22800 S0.n41 S0.n38 1.85764
R22801 S0.n39 S0.n5 1.60126
R22802 S0.n21 S0.n20 1.15434
R22803 S0.n34 S0.n8 1.0245
R22804 S0.n25 S0 0.7685
R22805 S0.n29 S0.n28 0.5125
R22806 S0.n23 S0.n20 0.5125
R22807 S0.n38 S0.n6 0.462934
R22808 S0.n42 S0.n41 0.429669
R22809 S0.n3 S0 0.232242
R22810 S0.n42 S0.n5 0.230918
R22811 S0.n3 S0 0.212579
R22812 S0.n40 S0.n39 0.12975
R22813 S0.n3 S0 0.129406
R22814 S0.n32 S0.n31 0.0766364
R22815 S0.n37 S0.n7 0.0618636
R22816 S0.n43 S0.n42 0.0592506
R22817 S0.n4 S0.n3 0.0590938
R22818 S0.n26 S0.n16 0.0516364
R22819 S0 S0.n43 0.0395625
R22820 S0.n38 S0.n37 0.0239512
R22821 S0.n27 S0.n26 0.0209545
R22822 S0.n43 S0.n4 0.0200312
R22823 S0.n31 S0.n9 0.0198182
R22824 S0.n22 S0.n16 0.0198182
R22825 S0.n33 S0.n7 0.0186818
R22826 S0.n4 S0 0.0156515
R22827 S0.n33 S0.n32 0.00504545
R22828 S0.n41 S0.n40 0.0028536
R22829 S0.n27 S0.n9 0.00277273
R22830 S0.n34 S0.n33 0.00119114
R22831 S0.n28 S0.n27 0.00119114
R22832 S0.n23 S0.n22 0.00119114
R22833 frontAnalog_v0p0p1_15.RSfetsym_0.QN.n1 frontAnalog_v0p0p1_15.RSfetsym_0.QN.t6 117.511
R22834 frontAnalog_v0p0p1_15.RSfetsym_0.QN.n1 frontAnalog_v0p0p1_15.RSfetsym_0.QN.t5 110.698
R22835 frontAnalog_v0p0p1_15.RSfetsym_0.QN.n2 frontAnalog_v0p0p1_15.RSfetsym_0.QN.t2 19.1963
R22836 frontAnalog_v0p0p1_15.RSfetsym_0.QN.n3 frontAnalog_v0p0p1_15.RSfetsym_0.QN.t1 14.5206
R22837 frontAnalog_v0p0p1_15.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_15.RSfetsym_0.QN.t4 14.283
R22838 frontAnalog_v0p0p1_15.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_15.RSfetsym_0.QN.t3 14.283
R22839 frontAnalog_v0p0p1_15.RSfetsym_0.QN frontAnalog_v0p0p1_15.RSfetsym_0.QN.t0 9.14075
R22840 frontAnalog_v0p0p1_15.RSfetsym_0.QN.n2 frontAnalog_v0p0p1_15.RSfetsym_0.QN.n1 0.826818
R22841 frontAnalog_v0p0p1_15.RSfetsym_0.QN frontAnalog_v0p0p1_15.RSfetsym_0.QN.n0 0.74645
R22842 frontAnalog_v0p0p1_15.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_15.RSfetsym_0.QN.n3 0.249509
R22843 frontAnalog_v0p0p1_15.RSfetsym_0.QN.n3 frontAnalog_v0p0p1_15.RSfetsym_0.QN.n2 0.0968646
R22844 I10.n6 I10.t12 323.342
R22845 I10.n0 I10.t11 228.927
R22846 I10.n3 I10.t6 196.549
R22847 I10.n6 I10.t10 194.809
R22848 I10.n0 I10.t8 159.391
R22849 I10.n3 I10.t9 148.35
R22850 I10.n10 I10.t7 117.314
R22851 I10.n10 I10.t5 110.852
R22852 I10.n7 I10.n6 76.0005
R22853 I10.n4 I10.n3 76.0005
R22854 I10.n8 I10.n7 29.3651
R22855 I10.n12 I10.t1 17.6181
R22856 I10.n13 I10.t0 14.2865
R22857 I10.n15 I10.t2 14.283
R22858 I10.n15 I10.t3 14.283
R22859 I10.n5 I10 9.11
R22860 I10.n17 I10.t4 8.77592
R22861 I10.n1 I10.n0 8.6846
R22862 I10.n4 I10 5.78114
R22863 I10.n2 I10.n1 4.26809
R22864 I10 I10.n4 3.71663
R22865 I10 I10.n18 2.22491
R22866 I10.n1 I10 1.99652
R22867 I10.n7 I10 1.92927
R22868 I10.n8 I10.n5 1.69246
R22869 I10.n17 I10.n16 1.20426
R22870 I10.n19 I10 0.760333
R22871 I10 I10.n9 0.7337
R22872 I10.n5 I10.n2 0.570143
R22873 I10 I10.n19 0.4564
R22874 I10.n18 I10.n17 0.336084
R22875 I10.n13 I10.n12 0.314673
R22876 I10.n14 I10.n13 0.300251
R22877 I10.n9 I10.n8 0.224535
R22878 I10.n2 I10 0.221483
R22879 I10.n9 I10 0.2005
R22880 I10.n11 I10.n10 0.159555
R22881 I10.n16 I10.n15 0.106617
R22882 I10.n14 I10.n11 0.0796167
R22883 I10.n16 I10.n14 0.0480595
R22884 I10.n19 I10 0.0161667
R22885 I10.n19 I10 0.0099
R22886 I10.n18 I10 0.00658123
R22887 I10.n12 I10.n11 0.000504658
R22888 frontAnalog_v0p0p1_6.RSfetsym_0.QN.n1 frontAnalog_v0p0p1_6.RSfetsym_0.QN.t6 117.511
R22889 frontAnalog_v0p0p1_6.RSfetsym_0.QN.n1 frontAnalog_v0p0p1_6.RSfetsym_0.QN.t5 110.698
R22890 frontAnalog_v0p0p1_6.RSfetsym_0.QN.n2 frontAnalog_v0p0p1_6.RSfetsym_0.QN.t2 19.1963
R22891 frontAnalog_v0p0p1_6.RSfetsym_0.QN.n3 frontAnalog_v0p0p1_6.RSfetsym_0.QN.t3 14.5206
R22892 frontAnalog_v0p0p1_6.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_6.RSfetsym_0.QN.t0 14.283
R22893 frontAnalog_v0p0p1_6.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_6.RSfetsym_0.QN.t1 14.283
R22894 frontAnalog_v0p0p1_6.RSfetsym_0.QN frontAnalog_v0p0p1_6.RSfetsym_0.QN.t4 9.14075
R22895 frontAnalog_v0p0p1_6.RSfetsym_0.QN.n2 frontAnalog_v0p0p1_6.RSfetsym_0.QN.n1 0.826818
R22896 frontAnalog_v0p0p1_6.RSfetsym_0.QN frontAnalog_v0p0p1_6.RSfetsym_0.QN.n0 0.74645
R22897 frontAnalog_v0p0p1_6.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_6.RSfetsym_0.QN.n3 0.249509
R22898 frontAnalog_v0p0p1_6.RSfetsym_0.QN.n3 frontAnalog_v0p0p1_6.RSfetsym_0.QN.n2 0.0968646
R22899 I13.t9 I13.t13 618.109
R22900 I13.n12 I13.t14 259.74
R22901 I13 I13.t9 253.56
R22902 I13.n0 I13.t11 228.899
R22903 I13.n19 I13.t6 180.286
R22904 I13.n0 I13.t10 159.411
R22905 I13.n12 I13.t8 157.083
R22906 I13.n29 I13.t5 117.314
R22907 I13.n20 I13.t7 111.091
R22908 I13.n29 I13.t12 110.852
R22909 I13.n23 I13 37.7071
R22910 I13.n31 I13.t4 17.6181
R22911 I13.n32 I13.t1 14.2865
R22912 I13.n34 I13.t2 14.283
R22913 I13.n34 I13.t3 14.283
R22914 I13.n21 I13.n20 9.3005
R22915 I13 I13.n11 9.3005
R22916 I13.n36 I13.t0 8.77592
R22917 I13.n22 I13.n21 7.80966
R22918 I13.n13 I13.n12 7.57248
R22919 I13.n1 I13.n0 7.36885
R22920 I13.n20 I13.n19 6.53562
R22921 I13 I13.n37 4.95588
R22922 I13.n13 I13 4.8645
R22923 I13.n3 I13.n2 3.46717
R22924 I13.n4 I13.n3 3.03286
R22925 I13.n18 I13.n17 2.32777
R22926 I13.n22 I13.n16 2.19001
R22927 I13.n17 I13 1.4966
R22928 I13.n36 I13.n35 1.20426
R22929 I13.n24 I13.n9 1.16836
R22930 I13.n23 I13.n22 1.07639
R22931 I13.n3 I13.n1 1.06717
R22932 I13.n2 I13 1.06717
R22933 I13.n25 I13 0.823
R22934 I13.n9 I13.n8 0.71595
R22935 I13.n27 I13 0.68435
R22936 I13.n28 I13 0.653017
R22937 I13 I13.n28 0.649412
R22938 I13.n21 I13.n18 0.499201
R22939 I13.n25 I13.n24 0.430355
R22940 I13.n37 I13.n36 0.336084
R22941 I13.n32 I13.n31 0.314673
R22942 I13.n33 I13.n32 0.300251
R22943 I13.n9 I13 0.221483
R22944 I13.n26 I13 0.2005
R22945 I13.n24 I13.n23 0.192464
R22946 I13.n30 I13.n29 0.159555
R22947 I13.n28 I13.n27 0.107817
R22948 I13.n35 I13.n34 0.106617
R22949 I13.n33 I13.n30 0.0796167
R22950 I13.n35 I13.n33 0.0480595
R22951 I13.n11 I13.n10 0.0301875
R22952 I13.n26 I13.n25 0.0287
R22953 I13.n27 I13.n26 0.0287
R22954 I13.n16 I13.n15 0.0205312
R22955 I13.n37 I13 0.00658123
R22956 I13.n6 I13.n5 0.00618182
R22957 I13.n5 I13.n4 0.00555107
R22958 I13.n7 I13.n6 0.00430477
R22959 I13.n15 I13.n14 0.00210765
R22960 I13.n14 I13.n13 0.00133438
R22961 I13.n8 I13.n7 0.00101192
R22962 I13.n14 I13.n10 0.00100001
R22963 I13.n31 I13.n30 0.000504658
R22964 frontAnalog_v0p0p1_10.IB.n0 frontAnalog_v0p0p1_10.IB.t1 182.794
R22965 frontAnalog_v0p0p1_10.IB.n1 frontAnalog_v0p0p1_10.IB.t12 91.7714
R22966 frontAnalog_v0p0p1_10.IB.n17 frontAnalog_v0p0p1_10.IB.t17 91.7714
R22967 frontAnalog_v0p0p1_10.IB.n16 frontAnalog_v0p0p1_10.IB.t14 91.7714
R22968 frontAnalog_v0p0p1_10.IB.n15 frontAnalog_v0p0p1_10.IB.t27 91.7714
R22969 frontAnalog_v0p0p1_10.IB.n14 frontAnalog_v0p0p1_10.IB.t21 91.7714
R22970 frontAnalog_v0p0p1_10.IB.n13 frontAnalog_v0p0p1_10.IB.t4 91.7714
R22971 frontAnalog_v0p0p1_10.IB.n12 frontAnalog_v0p0p1_10.IB.t31 91.7714
R22972 frontAnalog_v0p0p1_10.IB.n11 frontAnalog_v0p0p1_10.IB.t10 91.7714
R22973 frontAnalog_v0p0p1_10.IB.n10 frontAnalog_v0p0p1_10.IB.t7 91.7714
R22974 frontAnalog_v0p0p1_10.IB.n9 frontAnalog_v0p0p1_10.IB.t18 91.7714
R22975 frontAnalog_v0p0p1_10.IB.n8 frontAnalog_v0p0p1_10.IB.t15 91.7714
R22976 frontAnalog_v0p0p1_10.IB.n7 frontAnalog_v0p0p1_10.IB.t26 91.7714
R22977 frontAnalog_v0p0p1_10.IB.n6 frontAnalog_v0p0p1_10.IB.t22 91.7714
R22978 frontAnalog_v0p0p1_10.IB.n5 frontAnalog_v0p0p1_10.IB.t5 91.7714
R22979 frontAnalog_v0p0p1_10.IB.n4 frontAnalog_v0p0p1_10.IB.t32 91.7714
R22980 frontAnalog_v0p0p1_10.IB.n2 frontAnalog_v0p0p1_10.IB.t3 91.7714
R22981 frontAnalog_v0p0p1_10.IB.n17 frontAnalog_v0p0p1_10.IB.t28 91.3136
R22982 frontAnalog_v0p0p1_10.IB.n16 frontAnalog_v0p0p1_10.IB.t24 91.3136
R22983 frontAnalog_v0p0p1_10.IB.n15 frontAnalog_v0p0p1_10.IB.t6 91.3136
R22984 frontAnalog_v0p0p1_10.IB.n14 frontAnalog_v0p0p1_10.IB.t33 91.3136
R22985 frontAnalog_v0p0p1_10.IB.n13 frontAnalog_v0p0p1_10.IB.t13 91.3136
R22986 frontAnalog_v0p0p1_10.IB.n12 frontAnalog_v0p0p1_10.IB.t8 91.3136
R22987 frontAnalog_v0p0p1_10.IB.n11 frontAnalog_v0p0p1_10.IB.t20 91.3136
R22988 frontAnalog_v0p0p1_10.IB.n10 frontAnalog_v0p0p1_10.IB.t16 91.3136
R22989 frontAnalog_v0p0p1_10.IB.n9 frontAnalog_v0p0p1_10.IB.t30 91.3136
R22990 frontAnalog_v0p0p1_10.IB.n8 frontAnalog_v0p0p1_10.IB.t25 91.3136
R22991 frontAnalog_v0p0p1_10.IB.n7 frontAnalog_v0p0p1_10.IB.t19 91.3136
R22992 frontAnalog_v0p0p1_10.IB.n6 frontAnalog_v0p0p1_10.IB.t34 91.3136
R22993 frontAnalog_v0p0p1_10.IB.n5 frontAnalog_v0p0p1_10.IB.t29 91.3136
R22994 frontAnalog_v0p0p1_10.IB.n4 frontAnalog_v0p0p1_10.IB.t9 91.3136
R22995 frontAnalog_v0p0p1_10.IB.n2 frontAnalog_v0p0p1_10.IB.t11 91.3136
R22996 frontAnalog_v0p0p1_10.IB.n1 frontAnalog_v0p0p1_10.IB.t23 91.3136
R22997 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_10.IB.n17 45.9747
R22998 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_10.IB.n16 45.9747
R22999 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_10.IB.n15 45.9747
R23000 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_10.IB.n14 45.9747
R23001 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_10.IB.n13 45.9747
R23002 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_10.IB.n12 45.9747
R23003 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_10.IB.n11 45.9747
R23004 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_10.IB.n10 45.9747
R23005 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_10.IB.n9 45.9747
R23006 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_10.IB.n8 45.9747
R23007 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_10.IB.n7 45.9747
R23008 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_10.IB.n6 45.9747
R23009 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_10.IB.n5 45.9747
R23010 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_10.IB.n4 45.9747
R23011 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_10.IB.n2 45.9747
R23012 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_10.IB.n1 45.973
R23013 frontAnalog_v0p0p1_10.IB.n34 frontAnalog_v0p0p1_10.IB.t0 5.91044
R23014 frontAnalog_v0p0p1_10.IB.n32 frontAnalog_v0p0p1_10.IB.t2 4.35136
R23015 frontAnalog_v0p0p1_10.IB.n18 frontAnalog_v0p0p1_10.IB 1.53808
R23016 frontAnalog_v0p0p1_10.IB.n34 frontAnalog_v0p0p1_10.IB.n31 1.41054
R23017 frontAnalog_v0p0p1_10.IB.n3 frontAnalog_v0p0p1_10.IB 1.28321
R23018 frontAnalog_v0p0p1_10.IB.n29 frontAnalog_v0p0p1_10.IB 1.15021
R23019 frontAnalog_v0p0p1_10.IB.n28 frontAnalog_v0p0p1_10.IB 1.14904
R23020 frontAnalog_v0p0p1_10.IB.n26 frontAnalog_v0p0p1_10.IB 1.14883
R23021 frontAnalog_v0p0p1_10.IB.n30 frontAnalog_v0p0p1_10.IB 1.14802
R23022 frontAnalog_v0p0p1_10.IB.n19 frontAnalog_v0p0p1_10.IB 1.14536
R23023 frontAnalog_v0p0p1_10.IB.n25 frontAnalog_v0p0p1_10.IB 1.14495
R23024 frontAnalog_v0p0p1_10.IB.n27 frontAnalog_v0p0p1_10.IB 1.14447
R23025 frontAnalog_v0p0p1_10.IB.n21 frontAnalog_v0p0p1_10.IB 1.14439
R23026 frontAnalog_v0p0p1_10.IB.n22 frontAnalog_v0p0p1_10.IB 1.14419
R23027 frontAnalog_v0p0p1_10.IB.n24 frontAnalog_v0p0p1_10.IB 1.14189
R23028 frontAnalog_v0p0p1_10.IB.n23 frontAnalog_v0p0p1_10.IB 1.14114
R23029 frontAnalog_v0p0p1_10.IB.n18 frontAnalog_v0p0p1_10.IB 1.13988
R23030 frontAnalog_v0p0p1_10.IB.n20 frontAnalog_v0p0p1_10.IB 1.13929
R23031 frontAnalog_v0p0p1_10.IB.n3 frontAnalog_v0p0p1_10.IB 0.957022
R23032 frontAnalog_v0p0p1_10.IB.n33 frontAnalog_v0p0p1_10.IB.n32 0.807781
R23033 frontAnalog_v0p0p1_10.IB.n34 frontAnalog_v0p0p1_10.IB.n0 0.504831
R23034 frontAnalog_v0p0p1_10.IB.n30 frontAnalog_v0p0p1_10.IB.n29 0.399765
R23035 frontAnalog_v0p0p1_10.IB.n28 frontAnalog_v0p0p1_10.IB.n27 0.399029
R23036 frontAnalog_v0p0p1_10.IB.n25 frontAnalog_v0p0p1_10.IB.n24 0.399029
R23037 frontAnalog_v0p0p1_10.IB.n23 frontAnalog_v0p0p1_10.IB.n22 0.398294
R23038 frontAnalog_v0p0p1_10.IB.n21 frontAnalog_v0p0p1_10.IB.n20 0.398294
R23039 frontAnalog_v0p0p1_10.IB.n26 frontAnalog_v0p0p1_10.IB.n25 0.397559
R23040 frontAnalog_v0p0p1_10.IB.n22 frontAnalog_v0p0p1_10.IB.n21 0.396824
R23041 frontAnalog_v0p0p1_10.IB.n20 frontAnalog_v0p0p1_10.IB.n19 0.396824
R23042 frontAnalog_v0p0p1_10.IB.n19 frontAnalog_v0p0p1_10.IB.n18 0.396824
R23043 frontAnalog_v0p0p1_10.IB.n27 frontAnalog_v0p0p1_10.IB.n26 0.396088
R23044 frontAnalog_v0p0p1_10.IB.n24 frontAnalog_v0p0p1_10.IB.n23 0.396088
R23045 frontAnalog_v0p0p1_10.IB.n29 frontAnalog_v0p0p1_10.IB.n28 0.395353
R23046 frontAnalog_v0p0p1_10.IB.n31 frontAnalog_v0p0p1_10.IB.n30 0.249029
R23047 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_10.IB.n34 0.168769
R23048 frontAnalog_v0p0p1_10.IB.n31 frontAnalog_v0p0p1_10.IB.n3 0.151971
R23049 frontAnalog_v0p0p1_10.IB.n0 frontAnalog_v0p0p1_10.IB.n33 0.0762967
R23050 VV14.n0 VV14.t17 167.365
R23051 VV14.n0 VV14.t16 92.4496
R23052 VV14.n1 VV14.n0 2.07493
R23053 VV14.n10 VV14 0.638917
R23054 VV14 VV14.n10 0.479312
R23055 VV14.n9 VV14.n8 0.141636
R23056 VV14.n8 VV14.n7 0.141636
R23057 VV14.n7 VV14.n6 0.141636
R23058 VV14.n6 VV14.n5 0.141636
R23059 VV14.n5 VV14.n4 0.141636
R23060 VV14.n4 VV14.n3 0.141636
R23061 VV14.n3 VV14.n2 0.141636
R23062 VV14.n1 VV14 0.12425
R23063 VV14 VV14.n9 0.102242
R23064 VV14 VV14.n1 0.0358571
R23065 VV14.n10 VV14 0.00833333
R23066 VV14.n10 VV14 0.006375
R23067 VV14.n2 VV14.t14 0.000502142
R23068 VV14.n3 VV14.t6 0.000502142
R23069 VV14.n4 VV14.t2 0.000502142
R23070 VV14.n5 VV14.t8 0.000502142
R23071 VV14.n6 VV14.t10 0.000502142
R23072 VV14.n7 VV14.t11 0.000502142
R23073 VV14.n8 VV14.t7 0.000502142
R23074 VV14.n9 VV14.t0 0.000502142
R23075 VV14.n9 VV14.t9 0.000502142
R23076 VV14.n8 VV14.t3 0.000502142
R23077 VV14.n7 VV14.t4 0.000502142
R23078 VV14.n6 VV14.t5 0.000502142
R23079 VV14.n5 VV14.t13 0.000502142
R23080 VV14.n4 VV14.t12 0.000502142
R23081 VV14.n3 VV14.t15 0.000502142
R23082 VV14.n2 VV14.t1 0.000502142
R23083 VV13.n0 VV13.t16 167.365
R23084 VV13.n0 VV13.t17 92.4496
R23085 VV13.n1 VV13.n0 2.07493
R23086 VV13.n10 VV13 0.59975
R23087 VV13 VV13.n10 0.449937
R23088 VV13.n9 VV13.n8 0.141636
R23089 VV13.n8 VV13.n7 0.141636
R23090 VV13.n7 VV13.n6 0.141636
R23091 VV13.n6 VV13.n5 0.141636
R23092 VV13.n5 VV13.n4 0.141636
R23093 VV13.n4 VV13.n3 0.141636
R23094 VV13.n3 VV13.n2 0.141636
R23095 VV13.n1 VV13 0.12425
R23096 VV13 VV13.n9 0.0991174
R23097 VV13 VV13.n1 0.0314375
R23098 VV13.n10 VV13 0.00833333
R23099 VV13.n10 VV13 0.006375
R23100 VV13.n2 VV13.t7 0.000502142
R23101 VV13.n3 VV13.t10 0.000502142
R23102 VV13.n4 VV13.t2 0.000502142
R23103 VV13.n5 VV13.t13 0.000502142
R23104 VV13.n6 VV13.t9 0.000502142
R23105 VV13.n7 VV13.t8 0.000502142
R23106 VV13.n8 VV13.t14 0.000502142
R23107 VV13.n9 VV13.t0 0.000502142
R23108 VV13.n9 VV13.t1 0.000502142
R23109 VV13.n8 VV13.t5 0.000502142
R23110 VV13.n7 VV13.t12 0.000502142
R23111 VV13.n6 VV13.t11 0.000502142
R23112 VV13.n5 VV13.t6 0.000502142
R23113 VV13.n4 VV13.t3 0.000502142
R23114 VV13.n3 VV13.t4 0.000502142
R23115 VV13.n2 VV13.t15 0.000502142
R23116 VIN.n3 VIN.t19 167.326
R23117 VIN.n18 VIN.t11 167.326
R23118 VIN.n17 VIN.t5 167.326
R23119 VIN.n16 VIN.t20 167.326
R23120 VIN.n15 VIN.t15 167.326
R23121 VIN.n14 VIN.t26 167.326
R23122 VIN.n13 VIN.t23 167.326
R23123 VIN.n12 VIN.t1 167.326
R23124 VIN.n11 VIN.t28 167.326
R23125 VIN.n10 VIN.t13 167.326
R23126 VIN.n9 VIN.t6 167.326
R23127 VIN.n8 VIN.t31 167.326
R23128 VIN.n7 VIN.t16 167.326
R23129 VIN.n6 VIN.t10 167.326
R23130 VIN.n5 VIN.t24 167.326
R23131 VIN.n0 VIN.t4 167.326
R23132 VIN.n3 VIN.t17 92.4649
R23133 VIN.n18 VIN.t7 92.4649
R23134 VIN.n17 VIN.t0 92.4649
R23135 VIN.n16 VIN.t18 92.4649
R23136 VIN.n15 VIN.t12 92.4649
R23137 VIN.n14 VIN.t25 92.4649
R23138 VIN.n13 VIN.t21 92.4649
R23139 VIN.n12 VIN.t30 92.4649
R23140 VIN.n11 VIN.t27 92.4649
R23141 VIN.n10 VIN.t9 92.4649
R23142 VIN.n9 VIN.t2 92.4649
R23143 VIN.n8 VIN.t29 92.4649
R23144 VIN.n7 VIN.t14 92.4649
R23145 VIN.n6 VIN.t8 92.4649
R23146 VIN.n5 VIN.t22 92.4649
R23147 VIN.n0 VIN.t3 92.4649
R23148 VIN.n1 VIN 4.6255
R23149 VIN.n2 VIN.n1 1.6255
R23150 VIN VIN.n18 1.49913
R23151 VIN VIN.n17 1.49913
R23152 VIN VIN.n16 1.49913
R23153 VIN VIN.n15 1.49913
R23154 VIN VIN.n14 1.49913
R23155 VIN VIN.n13 1.49913
R23156 VIN VIN.n12 1.49913
R23157 VIN VIN.n11 1.49913
R23158 VIN VIN.n10 1.49913
R23159 VIN VIN.n9 1.49913
R23160 VIN VIN.n8 1.49913
R23161 VIN VIN.n7 1.49913
R23162 VIN VIN.n5 1.49913
R23163 VIN.n1 VIN.n0 1.49913
R23164 VIN VIN.n3 1.46056
R23165 VIN VIN.n6 1.46056
R23166 VIN.n19 VIN 1.04323
R23167 VIN.n32 VIN.n4 0.573417
R23168 VIN.n32 VIN.n31 0.563
R23169 VIN.n31 VIN.n30 0.563
R23170 VIN.n30 VIN.n29 0.563
R23171 VIN.n29 VIN.n28 0.563
R23172 VIN.n28 VIN.n27 0.563
R23173 VIN.n27 VIN.n26 0.563
R23174 VIN.n26 VIN.n25 0.563
R23175 VIN.n25 VIN.n24 0.563
R23176 VIN.n24 VIN.n23 0.563
R23177 VIN.n23 VIN.n22 0.563
R23178 VIN.n22 VIN.n21 0.563
R23179 VIN.n21 VIN.n20 0.563
R23180 VIN.n20 VIN.n19 0.563
R23181 VIN.n4 VIN 0.517333
R23182 VIN.n25 VIN 0.496386
R23183 VIN.n20 VIN 0.484963
R23184 VIN.n22 VIN 0.484963
R23185 VIN.n23 VIN 0.484963
R23186 VIN.n24 VIN 0.484963
R23187 VIN.n26 VIN 0.484963
R23188 VIN.n27 VIN 0.484963
R23189 VIN.n28 VIN 0.484963
R23190 VIN.n21 VIN 0.480732
R23191 VIN.n29 VIN 0.480732
R23192 VIN.n33 VIN.n32 0.47425
R23193 VIN.n19 VIN 0.473007
R23194 VIN.n31 VIN 0.473007
R23195 VIN.n30 VIN 0.45875
R23196 VIN.n2 VIN 0.316289
R23197 VIN.n4 VIN 0.169571
R23198 VIN VIN.n33 0.01
R23199 VIN.n33 VIN.n2 0.00707895
R23200 R0 R0.t1 451.853
R23201 R0.n45 R0.t1 440.25
R23202 R0.n0 R0.t5 258.584
R23203 R0.n38 R0.t9 258.58
R23204 R0.n11 R0.t3 212.081
R23205 R0.n5 R0.t4 212.081
R23206 R0.n4 R0.t8 212.081
R23207 R0.n24 R0.t10 212.081
R23208 R0.n11 R0.t12 139.78
R23209 R0.n5 R0.t2 139.78
R23210 R0.n4 R0.t6 139.78
R23211 R0.n24 R0.t7 139.78
R23212 R0 R0.t0 126.855
R23213 R0.n34 R0.t11 110.734
R23214 R0.n46 R0.n45 50.2399
R23215 R0.n26 R0.n24 30.6732
R23216 R0.n6 R0.n4 30.6732
R23217 R0.n6 R0.n5 30.6732
R23218 R0.n12 R0.n11 30.6732
R23219 R0.n46 R0 25.4148
R23220 R0.n23 R0.n22 12.8005
R23221 R0.n26 R0.n25 12.4157
R23222 R0.n18 R0.n17 9.3005
R23223 R0.n32 R0.n31 9.3005
R23224 R0.n13 R0.n12 8.28655
R23225 R0.n21 R0.n6 8.28655
R23226 R0.n27 R0.n26 8.28655
R23227 R0.n22 R0.n21 4.3525
R23228 R0.n14 R0.n9 4.3525
R23229 R0.n10 R0 4.10569
R23230 R0.n28 R0.n3 4.0965
R23231 R0.n20 R0 3.8405
R23232 R0.n45 R0 2.84494
R23233 R0 R0.n1 2.3045
R23234 R0.n31 R0 2.3045
R23235 R0.n27 R0 2.3045
R23236 R0 R0.n46 2.07932
R23237 R0 R0.n23 2.0485
R23238 R0.n43 R0.n33 1.59023
R23239 R0.n13 R0.n10 1.15386
R23240 R0.n28 R0.n27 1.0245
R23241 R0.n17 R0 0.7685
R23242 R0.n21 R0.n20 0.5125
R23243 R0.n14 R0.n13 0.5125
R23244 R0.n33 R0.n1 0.462934
R23245 R0.n44 R0.n43 0.44229
R23246 R0.n44 R0.n0 0.179314
R23247 R0.n43 R0.n42 0.14376
R23248 R0.n7 R0.n2 0.105187
R23249 R0.n32 R0.n30 0.084875
R23250 R0.n18 R0.n16 0.0708125
R23251 R0.n47 R0.n44 0.0699392
R23252 R0.n42 R0.n41 0.0475
R23253 R0.n19 R0.n18 0.028625
R23254 R0.n8 R0.n7 0.0270625
R23255 R0.n16 R0.n15 0.0270625
R23256 R0.n47 R0 0.0268713
R23257 R0.n30 R0.n29 0.0255
R23258 R0.n33 R0.n32 0.0239512
R23259 R0.n36 R0.n35 0.0174119
R23260 R0.n37 R0.n34 0.0133182
R23261 R0.n29 R0.n2 0.00675
R23262 R0 R0.n47 0.00419198
R23263 R0.n19 R0.n8 0.003625
R23264 R0.n41 R0.n37 0.00263636
R23265 R0.n39 R0.n38 0.0020625
R23266 R0.n29 R0.n28 0.00119114
R23267 R0.n20 R0.n19 0.00119114
R23268 R0.n15 R0.n14 0.00119114
R23269 R0.n37 R0.n36 0.000747155
R23270 R0.n41 R0.n40 0.000588765
R23271 R0.n40 R0.n39 0.000588763
R23272 frontAnalog_v0p0p1_4.x65.A.n1 frontAnalog_v0p0p1_4.x65.A.t4 260.322
R23273 frontAnalog_v0p0p1_4.x65.A.n3 frontAnalog_v0p0p1_4.x65.A.t7 233.929
R23274 frontAnalog_v0p0p1_4.x65.A.n1 frontAnalog_v0p0p1_4.x65.A.t5 175.169
R23275 frontAnalog_v0p0p1_4.x65.A.n2 frontAnalog_v0p0p1_4.x65.A.t6 160.416
R23276 frontAnalog_v0p0p1_4.x65.A.n4 frontAnalog_v0p0p1_4.x65.A.t2 17.4109
R23277 frontAnalog_v0p0p1_4.x65.A.n4 frontAnalog_v0p0p1_4.x65.A.t3 10.2053
R23278 frontAnalog_v0p0p1_4.x65.A.n0 frontAnalog_v0p0p1_4.x65.A 2.78715
R23279 frontAnalog_v0p0p1_4.x65.A.n0 frontAnalog_v0p0p1_4.x65.A.n1 9.09103
R23280 frontAnalog_v0p0p1_4.x65.A.n6 frontAnalog_v0p0p1_4.x65.A.t0 7.94569
R23281 frontAnalog_v0p0p1_4.x65.A.n2 frontAnalog_v0p0p1_4.x65.A.t1 7.55846
R23282 frontAnalog_v0p0p1_4.x65.A.n5 frontAnalog_v0p0p1_4.x65.A.n3 1.4614
R23283 frontAnalog_v0p0p1_4.x65.A.n3 frontAnalog_v0p0p1_4.x65.A.n2 1.19626
R23284 frontAnalog_v0p0p1_4.x65.A.n6 frontAnalog_v0p0p1_4.x65.A.n5 0.836961
R23285 frontAnalog_v0p0p1_4.x65.A frontAnalog_v0p0p1_4.x65.A.n0 0.390342
R23286 frontAnalog_v0p0p1_4.x65.A.n5 frontAnalog_v0p0p1_4.x65.A.n4 0.154668
R23287 frontAnalog_v0p0p1_4.x65.A frontAnalog_v0p0p1_4.x65.A.n6 0.08175
R23288 VV12.n0 VV12.t17 167.365
R23289 VV12.n0 VV12.t16 92.4496
R23290 VV12.n1 VV12.n0 2.07493
R23291 VV12.n17 VV12 0.560583
R23292 VV12 VV12.n17 0.420563
R23293 VV12.n15 VV12.n14 0.141409
R23294 VV12.n13 VV12.n12 0.141409
R23295 VV12.n11 VV12.n10 0.141409
R23296 VV12.n9 VV12.n8 0.141409
R23297 VV12.n7 VV12.n6 0.141409
R23298 VV12.n5 VV12.n4 0.141409
R23299 VV12.n3 VV12.n2 0.141409
R23300 VV12.n1 VV12 0.12425
R23301 VV12 VV12.n16 0.100973
R23302 VV12 VV12.n1 0.0314375
R23303 VV12.n17 VV12 0.00833333
R23304 VV12.n17 VV12 0.006375
R23305 VV12.n2 VV12.t7 0.000729415
R23306 VV12.n16 VV12.n15 0.000727273
R23307 VV12.n14 VV12.n13 0.000727273
R23308 VV12.n12 VV12.n11 0.000727273
R23309 VV12.n10 VV12.n9 0.000727273
R23310 VV12.n8 VV12.n7 0.000727273
R23311 VV12.n6 VV12.n5 0.000727273
R23312 VV12.n4 VV12.n3 0.000727273
R23313 VV12.n2 VV12.t6 0.000502142
R23314 VV12.n4 VV12.t12 0.000502142
R23315 VV12.n6 VV12.t1 0.000502142
R23316 VV12.n8 VV12.t4 0.000502142
R23317 VV12.n10 VV12.t8 0.000502142
R23318 VV12.n12 VV12.t5 0.000502142
R23319 VV12.n14 VV12.t15 0.000502142
R23320 VV12.n16 VV12.t2 0.000502142
R23321 VV12.n15 VV12.t0 0.000502142
R23322 VV12.n13 VV12.t14 0.000502142
R23323 VV12.n11 VV12.t9 0.000502142
R23324 VV12.n9 VV12.t10 0.000502142
R23325 VV12.n7 VV12.t13 0.000502142
R23326 VV12.n5 VV12.t3 0.000502142
R23327 VV12.n3 VV12.t11 0.000502142
R23328 frontAnalog_v0p0p1_9.x63.A.n2 frontAnalog_v0p0p1_9.x63.A.t5 260.322
R23329 frontAnalog_v0p0p1_9.x63.A.n4 frontAnalog_v0p0p1_9.x63.A.t6 233.888
R23330 frontAnalog_v0p0p1_9.x63.A.n2 frontAnalog_v0p0p1_9.x63.A.t7 175.169
R23331 frontAnalog_v0p0p1_9.x63.A.n3 frontAnalog_v0p0p1_9.x63.A.t4 159.725
R23332 frontAnalog_v0p0p1_9.x63.A.n1 frontAnalog_v0p0p1_9.x63.A.t0 17.4109
R23333 frontAnalog_v0p0p1_9.x63.A.n0 frontAnalog_v0p0p1_9.x63.A.n2 9.75129
R23334 frontAnalog_v0p0p1_9.x63.A.n1 frontAnalog_v0p0p1_9.x63.A.t1 9.6027
R23335 frontAnalog_v0p0p1_9.x63.A.n0 frontAnalog_v0p0p1_9.x63.A 2.33338
R23336 frontAnalog_v0p0p1_9.x63.A.n5 frontAnalog_v0p0p1_9.x63.A.t2 8.40929
R23337 frontAnalog_v0p0p1_9.x63.A.n3 frontAnalog_v0p0p1_9.x63.A.t3 8.06629
R23338 frontAnalog_v0p0p1_9.x63.A.n4 frontAnalog_v0p0p1_9.x63.A.n3 1.73501
R23339 frontAnalog_v0p0p1_9.x63.A.n1 frontAnalog_v0p0p1_9.x63.A.n4 0.99025
R23340 frontAnalog_v0p0p1_9.x63.A.n5 frontAnalog_v0p0p1_9.x63.A.n1 0.853186
R23341 frontAnalog_v0p0p1_9.x63.A frontAnalog_v0p0p1_9.x63.A.n0 0.349517
R23342 frontAnalog_v0p0p1_9.x63.A frontAnalog_v0p0p1_9.x63.A.n5 0.24425
R23343 frontAnalog_v0p0p1_9.x65.A.n1 frontAnalog_v0p0p1_9.x65.A.t6 260.322
R23344 frontAnalog_v0p0p1_9.x65.A.n3 frontAnalog_v0p0p1_9.x65.A.t5 233.929
R23345 frontAnalog_v0p0p1_9.x65.A.n1 frontAnalog_v0p0p1_9.x65.A.t4 175.169
R23346 frontAnalog_v0p0p1_9.x65.A.n2 frontAnalog_v0p0p1_9.x65.A.t7 160.416
R23347 frontAnalog_v0p0p1_9.x65.A.n4 frontAnalog_v0p0p1_9.x65.A.t0 17.4109
R23348 frontAnalog_v0p0p1_9.x65.A.n4 frontAnalog_v0p0p1_9.x65.A.t1 10.2053
R23349 frontAnalog_v0p0p1_9.x65.A.n0 frontAnalog_v0p0p1_9.x65.A 2.78715
R23350 frontAnalog_v0p0p1_9.x65.A.n0 frontAnalog_v0p0p1_9.x65.A.n1 9.09103
R23351 frontAnalog_v0p0p1_9.x65.A.n6 frontAnalog_v0p0p1_9.x65.A.t2 7.94569
R23352 frontAnalog_v0p0p1_9.x65.A.n2 frontAnalog_v0p0p1_9.x65.A.t3 7.55846
R23353 frontAnalog_v0p0p1_9.x65.A.n5 frontAnalog_v0p0p1_9.x65.A.n3 1.4614
R23354 frontAnalog_v0p0p1_9.x65.A.n3 frontAnalog_v0p0p1_9.x65.A.n2 1.19626
R23355 frontAnalog_v0p0p1_9.x65.A.n6 frontAnalog_v0p0p1_9.x65.A.n5 0.836961
R23356 frontAnalog_v0p0p1_9.x65.A frontAnalog_v0p0p1_9.x65.A.n0 0.390342
R23357 frontAnalog_v0p0p1_9.x65.A.n5 frontAnalog_v0p0p1_9.x65.A.n4 0.154668
R23358 frontAnalog_v0p0p1_9.x65.A frontAnalog_v0p0p1_9.x65.A.n6 0.08175
R23359 I1.t8 I1.t9 618.109
R23360 I1.n1 I1.t7 334.723
R23361 I1 I1.t8 253.56
R23362 I1.n1 I1.t6 206.19
R23363 I1.n5 I1.t10 117.314
R23364 I1.n5 I1.t5 110.853
R23365 I1 I1.n1 90.4462
R23366 I1.n0 I1 39.0702
R23367 I1.n7 I1.t2 17.6181
R23368 I1.n8 I1.t4 14.2865
R23369 I1.n10 I1.t0 14.283
R23370 I1.n10 I1.t1 14.283
R23371 I1.n12 I1.t3 8.77744
R23372 I1 I1.n13 8.44781
R23373 I1.n2 I1 7.13193
R23374 I1.n2 I1 5.30336
R23375 I1.n3 I1.n2 5.16688
R23376 I1.n3 I1.n0 2.29514
R23377 I1.n12 I1.n11 1.20426
R23378 I1.n0 I1 0.692911
R23379 I1.n13 I1.n12 0.32511
R23380 I1.n8 I1.n7 0.314673
R23381 I1.n9 I1.n8 0.299251
R23382 I1 I1.n14 0.2825
R23383 I1.n14 I1 0.212
R23384 I1.n4 I1 0.20675
R23385 I1.n6 I1.n5 0.159555
R23386 I1.n4 I1.n3 0.153447
R23387 I1.n11 I1.n10 0.106617
R23388 I1.n9 I1.n6 0.0796167
R23389 I1 I1.n4 0.0522
R23390 I1.n11 I1.n9 0.0480595
R23391 I1.n13 I1 0.046937
R23392 I1.n14 I1 0.0161667
R23393 I1.n14 I1 0.01225
R23394 I1.n7 I1.n6 0.000504658
R23395 frontAnalog_v0p0p1_9.RSfetsym_0.QN.n1 frontAnalog_v0p0p1_9.RSfetsym_0.QN.t6 117.511
R23396 frontAnalog_v0p0p1_9.RSfetsym_0.QN.n1 frontAnalog_v0p0p1_9.RSfetsym_0.QN.t5 110.698
R23397 frontAnalog_v0p0p1_9.RSfetsym_0.QN.n2 frontAnalog_v0p0p1_9.RSfetsym_0.QN.t1 19.1963
R23398 frontAnalog_v0p0p1_9.RSfetsym_0.QN.n3 frontAnalog_v0p0p1_9.RSfetsym_0.QN.t4 14.5206
R23399 frontAnalog_v0p0p1_9.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_9.RSfetsym_0.QN.t2 14.283
R23400 frontAnalog_v0p0p1_9.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_9.RSfetsym_0.QN.t3 14.283
R23401 frontAnalog_v0p0p1_9.RSfetsym_0.QN frontAnalog_v0p0p1_9.RSfetsym_0.QN.t0 9.14075
R23402 frontAnalog_v0p0p1_9.RSfetsym_0.QN.n2 frontAnalog_v0p0p1_9.RSfetsym_0.QN.n1 0.826818
R23403 frontAnalog_v0p0p1_9.RSfetsym_0.QN frontAnalog_v0p0p1_9.RSfetsym_0.QN.n0 0.74645
R23404 frontAnalog_v0p0p1_9.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_9.RSfetsym_0.QN.n3 0.249509
R23405 frontAnalog_v0p0p1_9.RSfetsym_0.QN.n3 frontAnalog_v0p0p1_9.RSfetsym_0.QN.n2 0.0968646
R23406 I6.n17 I6.t6 260.435
R23407 I6.n2 I6.t10 229.433
R23408 I6.n12 I6.t11 196.549
R23409 I6.n2 I6.t7 158.885
R23410 I6.n17 I6.t8 156.403
R23411 I6.n12 I6.t12 148.35
R23412 I6.n25 I6.t9 117.314
R23413 I6.n25 I6.t5 110.853
R23414 I6.n13 I6.n12 76.0005
R23415 I6.n27 I6.t4 17.6181
R23416 I6.n28 I6.t1 14.2865
R23417 I6.n30 I6.t2 14.283
R23418 I6.n30 I6.t3 14.283
R23419 I6.n5 I6.n4 9.3005
R23420 I6.n9 I6.n8 9.3005
R23421 I6.n5 I6.n3 9.3005
R23422 I6 I6.n16 9.3005
R23423 I6.n32 I6.t0 8.77744
R23424 I6.n18 I6.n17 7.60183
R23425 I6.n3 I6.n2 7.39171
R23426 I6.n22 I6.n14 6.24391
R23427 I6.n13 I6 5.78114
R23428 I6.n18 I6 4.8645
R23429 I6.n19 I6.n15 4.54557
R23430 I6.n10 I6.n9 4.51698
R23431 I6.n16 I6.n15 4.51121
R23432 I6.n8 I6.n7 4.5005
R23433 I6.n22 I6.n21 3.53643
R23434 I6.n14 I6.n13 3.51018
R23435 I6.n8 I6.n4 3.46717
R23436 I6 I6.n33 1.82181
R23437 I6.n32 I6.n31 1.20426
R23438 I6.n6 I6.n0 1.13339
R23439 I6.n11 I6.n10 1.11384
R23440 I6.n8 I6.n3 1.06717
R23441 I6.n4 I6 1.06717
R23442 I6.n23 I6.n11 0.874607
R23443 I6.n34 I6 0.6585
R23444 I6 I6.n24 0.647533
R23445 I6.n24 I6.n23 0.520635
R23446 I6 I6.n34 0.494
R23447 I6.n11 I6 0.372375
R23448 I6.n33 I6.n32 0.32511
R23449 I6.n28 I6.n27 0.314673
R23450 I6.n29 I6.n28 0.299251
R23451 I6.n23 I6.n22 0.214786
R23452 I6.n14 I6 0.206952
R23453 I6.n24 I6 0.20675
R23454 I6.n26 I6.n25 0.159555
R23455 I6.n31 I6.n30 0.106617
R23456 I6.n29 I6.n26 0.0796167
R23457 I6.n31 I6.n29 0.0480595
R23458 I6.n33 I6 0.046937
R23459 I6.n20 I6.n16 0.0344286
R23460 I6.n10 I6.n0 0.028
R23461 I6.n34 I6 0.0161667
R23462 I6.n9 I6.n1 0.0142363
R23463 I6.n34 I6 0.01225
R23464 I6.n7 I6.n1 0.00599451
R23465 I6.n6 I6.n5 0.00484776
R23466 I6.n7 I6.n6 0.00226981
R23467 I6.n21 I6.n15 0.00182856
R23468 I6.n21 I6.n20 0.00149885
R23469 I6.n19 I6.n18 0.00133362
R23470 I6.n20 I6.n19 0.00100077
R23471 I6.n1 I6.n0 0.000617139
R23472 I6.n27 I6.n26 0.000504658
R23473 frontAnalog_v0p0p1_13.RSfetsym_0.QN.n1 frontAnalog_v0p0p1_13.RSfetsym_0.QN.t6 117.511
R23474 frontAnalog_v0p0p1_13.RSfetsym_0.QN.n1 frontAnalog_v0p0p1_13.RSfetsym_0.QN.t5 110.698
R23475 frontAnalog_v0p0p1_13.RSfetsym_0.QN.n2 frontAnalog_v0p0p1_13.RSfetsym_0.QN.t2 19.1963
R23476 frontAnalog_v0p0p1_13.RSfetsym_0.QN.n3 frontAnalog_v0p0p1_13.RSfetsym_0.QN.t1 14.5206
R23477 frontAnalog_v0p0p1_13.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_13.RSfetsym_0.QN.t4 14.283
R23478 frontAnalog_v0p0p1_13.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_13.RSfetsym_0.QN.t3 14.283
R23479 frontAnalog_v0p0p1_13.RSfetsym_0.QN frontAnalog_v0p0p1_13.RSfetsym_0.QN.t0 9.14075
R23480 frontAnalog_v0p0p1_13.RSfetsym_0.QN.n2 frontAnalog_v0p0p1_13.RSfetsym_0.QN.n1 0.826818
R23481 frontAnalog_v0p0p1_13.RSfetsym_0.QN frontAnalog_v0p0p1_13.RSfetsym_0.QN.n0 0.74645
R23482 frontAnalog_v0p0p1_13.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_13.RSfetsym_0.QN.n3 0.249509
R23483 frontAnalog_v0p0p1_13.RSfetsym_0.QN.n3 frontAnalog_v0p0p1_13.RSfetsym_0.QN.n2 0.0968646
R23484 frontAnalog_v0p0p1_7.x65.A.n1 frontAnalog_v0p0p1_7.x65.A.t7 260.322
R23485 frontAnalog_v0p0p1_7.x65.A.n4 frontAnalog_v0p0p1_7.x65.A.t6 233.929
R23486 frontAnalog_v0p0p1_7.x65.A.n1 frontAnalog_v0p0p1_7.x65.A.t5 175.169
R23487 frontAnalog_v0p0p1_7.x65.A.n3 frontAnalog_v0p0p1_7.x65.A.t4 160.416
R23488 frontAnalog_v0p0p1_7.x65.A.n2 frontAnalog_v0p0p1_7.x65.A.t0 17.4109
R23489 frontAnalog_v0p0p1_7.x65.A.n2 frontAnalog_v0p0p1_7.x65.A.t3 10.2053
R23490 frontAnalog_v0p0p1_7.x65.A.n0 frontAnalog_v0p0p1_7.x65.A 2.78715
R23491 frontAnalog_v0p0p1_7.x65.A.n0 frontAnalog_v0p0p1_7.x65.A.n1 9.09103
R23492 frontAnalog_v0p0p1_7.x65.A.n6 frontAnalog_v0p0p1_7.x65.A.t2 7.94569
R23493 frontAnalog_v0p0p1_7.x65.A.n3 frontAnalog_v0p0p1_7.x65.A.t1 7.55846
R23494 frontAnalog_v0p0p1_7.x65.A.n5 frontAnalog_v0p0p1_7.x65.A.n4 1.4614
R23495 frontAnalog_v0p0p1_7.x65.A.n4 frontAnalog_v0p0p1_7.x65.A.n3 1.19626
R23496 frontAnalog_v0p0p1_7.x65.A.n6 frontAnalog_v0p0p1_7.x65.A.n5 0.836961
R23497 frontAnalog_v0p0p1_7.x65.A frontAnalog_v0p0p1_7.x65.A.n0 0.390342
R23498 frontAnalog_v0p0p1_7.x65.A.n5 frontAnalog_v0p0p1_7.x65.A.n2 0.154668
R23499 frontAnalog_v0p0p1_7.x65.A frontAnalog_v0p0p1_7.x65.A.n6 0.08175
R23500 frontAnalog_v0p0p1_7.x63.A.n2 frontAnalog_v0p0p1_7.x63.A.t6 260.322
R23501 frontAnalog_v0p0p1_7.x63.A.n4 frontAnalog_v0p0p1_7.x63.A.t7 233.888
R23502 frontAnalog_v0p0p1_7.x63.A.n2 frontAnalog_v0p0p1_7.x63.A.t4 175.169
R23503 frontAnalog_v0p0p1_7.x63.A.n3 frontAnalog_v0p0p1_7.x63.A.t5 159.725
R23504 frontAnalog_v0p0p1_7.x63.A.n1 frontAnalog_v0p0p1_7.x63.A.t0 17.4109
R23505 frontAnalog_v0p0p1_7.x63.A.n0 frontAnalog_v0p0p1_7.x63.A.n2 9.75129
R23506 frontAnalog_v0p0p1_7.x63.A.n1 frontAnalog_v0p0p1_7.x63.A.t1 9.6027
R23507 frontAnalog_v0p0p1_7.x63.A.n0 frontAnalog_v0p0p1_7.x63.A 2.33338
R23508 frontAnalog_v0p0p1_7.x63.A.n5 frontAnalog_v0p0p1_7.x63.A.t2 8.40929
R23509 frontAnalog_v0p0p1_7.x63.A.n3 frontAnalog_v0p0p1_7.x63.A.t3 8.06629
R23510 frontAnalog_v0p0p1_7.x63.A.n4 frontAnalog_v0p0p1_7.x63.A.n3 1.73501
R23511 frontAnalog_v0p0p1_7.x63.A.n1 frontAnalog_v0p0p1_7.x63.A.n4 0.99025
R23512 frontAnalog_v0p0p1_7.x63.A.n5 frontAnalog_v0p0p1_7.x63.A.n1 0.853186
R23513 frontAnalog_v0p0p1_7.x63.A frontAnalog_v0p0p1_7.x63.A.n0 0.349517
R23514 frontAnalog_v0p0p1_7.x63.A frontAnalog_v0p0p1_7.x63.A.n5 0.24425
R23515 I9.t7 I9.t9 618.109
R23516 I9.n1 I9.t8 334.723
R23517 I9 I9.t7 253.56
R23518 I9.n1 I9.t5 206.19
R23519 I9.n5 I9.t10 117.314
R23520 I9.n5 I9.t6 110.852
R23521 I9 I9.n1 90.4462
R23522 I9.n0 I9 39.0702
R23523 I9.n7 I9.t2 17.6181
R23524 I9.n8 I9.t4 14.2865
R23525 I9.n10 I9.t0 14.283
R23526 I9.n10 I9.t1 14.283
R23527 I9.n12 I9.t3 8.77592
R23528 I9.n2 I9 7.13193
R23529 I9.n2 I9 5.30336
R23530 I9.n3 I9.n2 5.27402
R23531 I9.n3 I9.n0 2.188
R23532 I9.n14 I9 1.2225
R23533 I9 I9.n4 1.20605
R23534 I9.n12 I9.n11 1.20426
R23535 I9 I9.n13 1.08107
R23536 I9.n0 I9 0.692911
R23537 I9 I9.n14 0.6115
R23538 I9.n13 I9.n12 0.338241
R23539 I9.n8 I9.n7 0.314673
R23540 I9.n9 I9.n8 0.300251
R23541 I9.n4 I9 0.2005
R23542 I9.n4 I9.n3 0.166764
R23543 I9.n6 I9.n5 0.159555
R23544 I9.n11 I9.n10 0.106617
R23545 I9.n9 I9.n6 0.0796167
R23546 I9.n11 I9.n9 0.0480595
R23547 I9.n14 I9 0.024
R23548 I9.n14 I9 0.01225
R23549 I9.n13 I9 0.00440792
R23550 I9.n7 I9.n6 0.000504658
R23551 VV7.n0 VV7.t16 167.365
R23552 VV7.n0 VV7.t17 92.4488
R23553 VV7.n1 VV7.n0 2.07493
R23554 VV7.n10 VV7 0.462667
R23555 VV7 VV7.n10 0.347125
R23556 VV7.n9 VV7.n8 0.141636
R23557 VV7.n8 VV7.n7 0.141636
R23558 VV7.n7 VV7.n6 0.141636
R23559 VV7.n6 VV7.n5 0.141636
R23560 VV7.n5 VV7.n4 0.141636
R23561 VV7.n4 VV7.n3 0.141636
R23562 VV7.n3 VV7.n2 0.141636
R23563 VV7.n1 VV7 0.12425
R23564 VV7 VV7.n9 0.101201
R23565 VV7 VV7.n1 0.028
R23566 VV7.n10 VV7 0.00833333
R23567 VV7.n10 VV7 0.006375
R23568 VV7.n3 VV7.t10 0.000502142
R23569 VV7.n4 VV7.t4 0.000502142
R23570 VV7.n5 VV7.t11 0.000502142
R23571 VV7.n6 VV7.t1 0.000502142
R23572 VV7.n7 VV7.t12 0.000502142
R23573 VV7.n8 VV7.t13 0.000502142
R23574 VV7.n9 VV7.t9 0.000502142
R23575 VV7.n2 VV7.t7 0.000502142
R23576 VV7.n3 VV7.t14 0.000502142
R23577 VV7.n4 VV7.t3 0.000502142
R23578 VV7.n5 VV7.t5 0.000502142
R23579 VV7.n6 VV7.t0 0.000502142
R23580 VV7.n7 VV7.t8 0.000502142
R23581 VV7.n8 VV7.t15 0.000502142
R23582 VV7.n9 VV7.t6 0.000502142
R23583 VV7.n2 VV7.t2 0.000502142
R23584 VV6.n0 VV6.t17 167.365
R23585 VV6.n0 VV6.t16 92.4488
R23586 VV6.n1 VV6.n0 2.07493
R23587 VV6.n17 VV6 0.501833
R23588 VV6 VV6.n17 0.3765
R23589 VV6.n15 VV6.n14 0.141409
R23590 VV6.n13 VV6.n12 0.141409
R23591 VV6.n11 VV6.n10 0.141409
R23592 VV6.n9 VV6.n8 0.141409
R23593 VV6.n7 VV6.n6 0.141409
R23594 VV6.n5 VV6.n4 0.141409
R23595 VV6.n3 VV6.n2 0.141409
R23596 VV6.n1 VV6 0.12425
R23597 VV6 VV6.n16 0.0988902
R23598 VV6 VV6.n1 0.0314375
R23599 VV6.n17 VV6 0.00833333
R23600 VV6.n17 VV6 0.006375
R23601 VV6.n2 VV6.t9 0.000729415
R23602 VV6.n16 VV6.n15 0.000727273
R23603 VV6.n14 VV6.n13 0.000727273
R23604 VV6.n12 VV6.n11 0.000727273
R23605 VV6.n10 VV6.n9 0.000727273
R23606 VV6.n8 VV6.n7 0.000727273
R23607 VV6.n6 VV6.n5 0.000727273
R23608 VV6.n4 VV6.n3 0.000727273
R23609 VV6.n3 VV6.t14 0.000502142
R23610 VV6.n5 VV6.t4 0.000502142
R23611 VV6.n7 VV6.t6 0.000502142
R23612 VV6.n9 VV6.t0 0.000502142
R23613 VV6.n11 VV6.t11 0.000502142
R23614 VV6.n13 VV6.t15 0.000502142
R23615 VV6.n15 VV6.t7 0.000502142
R23616 VV6.n2 VV6.t13 0.000502142
R23617 VV6.n4 VV6.t8 0.000502142
R23618 VV6.n6 VV6.t2 0.000502142
R23619 VV6.n8 VV6.t10 0.000502142
R23620 VV6.n10 VV6.t12 0.000502142
R23621 VV6.n12 VV6.t1 0.000502142
R23622 VV6.n14 VV6.t3 0.000502142
R23623 VV6.n16 VV6.t5 0.000502142
R23624 VV5.n0 VV5.t17 167.365
R23625 VV5.n0 VV5.t16 92.4488
R23626 VV5.n1 VV5.n0 2.07493
R23627 VV5.n17 VV5 0.537083
R23628 VV5 VV5.n17 0.402938
R23629 VV5.n15 VV5.n14 0.141409
R23630 VV5.n13 VV5.n12 0.141409
R23631 VV5.n11 VV5.n10 0.141409
R23632 VV5.n9 VV5.n8 0.141409
R23633 VV5.n7 VV5.n6 0.141409
R23634 VV5.n5 VV5.n4 0.141409
R23635 VV5.n3 VV5.n2 0.141409
R23636 VV5.n1 VV5 0.12425
R23637 VV5 VV5.n16 0.103057
R23638 VV5 VV5.n1 0.0314375
R23639 VV5.n17 VV5 0.00833333
R23640 VV5.n17 VV5 0.006375
R23641 VV5.n2 VV5.t11 0.000729415
R23642 VV5.n16 VV5.n15 0.000727273
R23643 VV5.n14 VV5.n13 0.000727273
R23644 VV5.n12 VV5.n11 0.000727273
R23645 VV5.n10 VV5.n9 0.000727273
R23646 VV5.n8 VV5.n7 0.000727273
R23647 VV5.n6 VV5.n5 0.000727273
R23648 VV5.n4 VV5.n3 0.000727273
R23649 VV5.n4 VV5.t8 0.000502142
R23650 VV5.n6 VV5.t4 0.000502142
R23651 VV5.n8 VV5.t10 0.000502142
R23652 VV5.n10 VV5.t13 0.000502142
R23653 VV5.n12 VV5.t0 0.000502142
R23654 VV5.n14 VV5.t5 0.000502142
R23655 VV5.n16 VV5.t7 0.000502142
R23656 VV5.n3 VV5.t14 0.000502142
R23657 VV5.n5 VV5.t6 0.000502142
R23658 VV5.n7 VV5.t2 0.000502142
R23659 VV5.n9 VV5.t12 0.000502142
R23660 VV5.n11 VV5.t3 0.000502142
R23661 VV5.n13 VV5.t9 0.000502142
R23662 VV5.n15 VV5.t1 0.000502142
R23663 VV5.n2 VV5.t15 0.000502142
R23664 frontAnalog_v0p0p1_13.x63.A.n2 frontAnalog_v0p0p1_13.x63.A.t4 260.322
R23665 frontAnalog_v0p0p1_13.x63.A.n4 frontAnalog_v0p0p1_13.x63.A.t5 233.888
R23666 frontAnalog_v0p0p1_13.x63.A.n2 frontAnalog_v0p0p1_13.x63.A.t6 175.169
R23667 frontAnalog_v0p0p1_13.x63.A.n3 frontAnalog_v0p0p1_13.x63.A.t7 159.725
R23668 frontAnalog_v0p0p1_13.x63.A.n1 frontAnalog_v0p0p1_13.x63.A.t3 17.4109
R23669 frontAnalog_v0p0p1_13.x63.A.n0 frontAnalog_v0p0p1_13.x63.A.n2 9.75129
R23670 frontAnalog_v0p0p1_13.x63.A.n1 frontAnalog_v0p0p1_13.x63.A.t0 9.6027
R23671 frontAnalog_v0p0p1_13.x63.A.n0 frontAnalog_v0p0p1_13.x63.A 2.33338
R23672 frontAnalog_v0p0p1_13.x63.A.n5 frontAnalog_v0p0p1_13.x63.A.t1 8.40929
R23673 frontAnalog_v0p0p1_13.x63.A.n3 frontAnalog_v0p0p1_13.x63.A.t2 8.06629
R23674 frontAnalog_v0p0p1_13.x63.A.n4 frontAnalog_v0p0p1_13.x63.A.n3 1.73501
R23675 frontAnalog_v0p0p1_13.x63.A.n1 frontAnalog_v0p0p1_13.x63.A.n4 0.99025
R23676 frontAnalog_v0p0p1_13.x63.A.n5 frontAnalog_v0p0p1_13.x63.A.n1 0.853186
R23677 frontAnalog_v0p0p1_13.x63.A frontAnalog_v0p0p1_13.x63.A.n0 0.349517
R23678 frontAnalog_v0p0p1_13.x63.A frontAnalog_v0p0p1_13.x63.A.n5 0.24425
R23679 frontAnalog_v0p0p1_10.x63.A.n2 frontAnalog_v0p0p1_10.x63.A.t5 260.322
R23680 frontAnalog_v0p0p1_10.x63.A.n4 frontAnalog_v0p0p1_10.x63.A.t6 233.888
R23681 frontAnalog_v0p0p1_10.x63.A.n2 frontAnalog_v0p0p1_10.x63.A.t7 175.169
R23682 frontAnalog_v0p0p1_10.x63.A.n3 frontAnalog_v0p0p1_10.x63.A.t4 159.725
R23683 frontAnalog_v0p0p1_10.x63.A.n1 frontAnalog_v0p0p1_10.x63.A.t0 17.4109
R23684 frontAnalog_v0p0p1_10.x63.A.n0 frontAnalog_v0p0p1_10.x63.A.n2 9.75129
R23685 frontAnalog_v0p0p1_10.x63.A.n1 frontAnalog_v0p0p1_10.x63.A.t1 9.6027
R23686 frontAnalog_v0p0p1_10.x63.A.n0 frontAnalog_v0p0p1_10.x63.A 2.33338
R23687 frontAnalog_v0p0p1_10.x63.A.n5 frontAnalog_v0p0p1_10.x63.A.t2 8.40929
R23688 frontAnalog_v0p0p1_10.x63.A.n3 frontAnalog_v0p0p1_10.x63.A.t3 8.06629
R23689 frontAnalog_v0p0p1_10.x63.A.n4 frontAnalog_v0p0p1_10.x63.A.n3 1.73501
R23690 frontAnalog_v0p0p1_10.x63.A.n1 frontAnalog_v0p0p1_10.x63.A.n4 0.99025
R23691 frontAnalog_v0p0p1_10.x63.A.n5 frontAnalog_v0p0p1_10.x63.A.n1 0.853186
R23692 frontAnalog_v0p0p1_10.x63.A frontAnalog_v0p0p1_10.x63.A.n0 0.349517
R23693 frontAnalog_v0p0p1_10.x63.A frontAnalog_v0p0p1_10.x63.A.n5 0.24425
R23694 frontAnalog_v0p0p1_5.x63.A.n2 frontAnalog_v0p0p1_5.x63.A.t4 260.322
R23695 frontAnalog_v0p0p1_5.x63.A.n4 frontAnalog_v0p0p1_5.x63.A.t5 233.888
R23696 frontAnalog_v0p0p1_5.x63.A.n2 frontAnalog_v0p0p1_5.x63.A.t6 175.169
R23697 frontAnalog_v0p0p1_5.x63.A.n3 frontAnalog_v0p0p1_5.x63.A.t7 159.725
R23698 frontAnalog_v0p0p1_5.x63.A.n1 frontAnalog_v0p0p1_5.x63.A.t0 17.4109
R23699 frontAnalog_v0p0p1_5.x63.A.n0 frontAnalog_v0p0p1_5.x63.A.n2 9.75129
R23700 frontAnalog_v0p0p1_5.x63.A.n1 frontAnalog_v0p0p1_5.x63.A.t1 9.6027
R23701 frontAnalog_v0p0p1_5.x63.A.n0 frontAnalog_v0p0p1_5.x63.A 2.33338
R23702 frontAnalog_v0p0p1_5.x63.A.n5 frontAnalog_v0p0p1_5.x63.A.t3 8.40929
R23703 frontAnalog_v0p0p1_5.x63.A.n3 frontAnalog_v0p0p1_5.x63.A.t2 8.06629
R23704 frontAnalog_v0p0p1_5.x63.A.n4 frontAnalog_v0p0p1_5.x63.A.n3 1.73501
R23705 frontAnalog_v0p0p1_5.x63.A.n1 frontAnalog_v0p0p1_5.x63.A.n4 0.99025
R23706 frontAnalog_v0p0p1_5.x63.A.n5 frontAnalog_v0p0p1_5.x63.A.n1 0.853186
R23707 frontAnalog_v0p0p1_5.x63.A frontAnalog_v0p0p1_5.x63.A.n0 0.349517
R23708 frontAnalog_v0p0p1_5.x63.A frontAnalog_v0p0p1_5.x63.A.n5 0.24425
R23709 frontAnalog_v0p0p1_3.x63.A.n2 frontAnalog_v0p0p1_3.x63.A.t5 260.322
R23710 frontAnalog_v0p0p1_3.x63.A.n4 frontAnalog_v0p0p1_3.x63.A.t6 233.888
R23711 frontAnalog_v0p0p1_3.x63.A.n2 frontAnalog_v0p0p1_3.x63.A.t7 175.169
R23712 frontAnalog_v0p0p1_3.x63.A.n3 frontAnalog_v0p0p1_3.x63.A.t4 159.725
R23713 frontAnalog_v0p0p1_3.x63.A.n1 frontAnalog_v0p0p1_3.x63.A.t1 17.4109
R23714 frontAnalog_v0p0p1_3.x63.A.n0 frontAnalog_v0p0p1_3.x63.A.n2 9.75129
R23715 frontAnalog_v0p0p1_3.x63.A.n1 frontAnalog_v0p0p1_3.x63.A.t0 9.6027
R23716 frontAnalog_v0p0p1_3.x63.A.n0 frontAnalog_v0p0p1_3.x63.A 2.33338
R23717 frontAnalog_v0p0p1_3.x63.A.n5 frontAnalog_v0p0p1_3.x63.A.t2 8.40929
R23718 frontAnalog_v0p0p1_3.x63.A.n3 frontAnalog_v0p0p1_3.x63.A.t3 8.06629
R23719 frontAnalog_v0p0p1_3.x63.A.n4 frontAnalog_v0p0p1_3.x63.A.n3 1.73501
R23720 frontAnalog_v0p0p1_3.x63.A.n1 frontAnalog_v0p0p1_3.x63.A.n4 0.99025
R23721 frontAnalog_v0p0p1_3.x63.A.n5 frontAnalog_v0p0p1_3.x63.A.n1 0.853186
R23722 frontAnalog_v0p0p1_3.x63.A frontAnalog_v0p0p1_3.x63.A.n0 0.349517
R23723 frontAnalog_v0p0p1_3.x63.A frontAnalog_v0p0p1_3.x63.A.n5 0.24425
R23724 frontAnalog_v0p0p1_3.x65.A.n1 frontAnalog_v0p0p1_3.x65.A.t4 260.322
R23725 frontAnalog_v0p0p1_3.x65.A.n3 frontAnalog_v0p0p1_3.x65.A.t7 233.929
R23726 frontAnalog_v0p0p1_3.x65.A.n1 frontAnalog_v0p0p1_3.x65.A.t6 175.169
R23727 frontAnalog_v0p0p1_3.x65.A.n2 frontAnalog_v0p0p1_3.x65.A.t5 160.416
R23728 frontAnalog_v0p0p1_3.x65.A.n4 frontAnalog_v0p0p1_3.x65.A.t1 17.4109
R23729 frontAnalog_v0p0p1_3.x65.A.n4 frontAnalog_v0p0p1_3.x65.A.t0 10.2053
R23730 frontAnalog_v0p0p1_3.x65.A.n0 frontAnalog_v0p0p1_3.x65.A 2.78715
R23731 frontAnalog_v0p0p1_3.x65.A.n0 frontAnalog_v0p0p1_3.x65.A.n1 9.09103
R23732 frontAnalog_v0p0p1_3.x65.A.n6 frontAnalog_v0p0p1_3.x65.A.t2 7.94569
R23733 frontAnalog_v0p0p1_3.x65.A.n2 frontAnalog_v0p0p1_3.x65.A.t3 7.55846
R23734 frontAnalog_v0p0p1_3.x65.A.n5 frontAnalog_v0p0p1_3.x65.A.n3 1.4614
R23735 frontAnalog_v0p0p1_3.x65.A.n3 frontAnalog_v0p0p1_3.x65.A.n2 1.19626
R23736 frontAnalog_v0p0p1_3.x65.A.n6 frontAnalog_v0p0p1_3.x65.A.n5 0.836961
R23737 frontAnalog_v0p0p1_3.x65.A frontAnalog_v0p0p1_3.x65.A.n0 0.390342
R23738 frontAnalog_v0p0p1_3.x65.A.n5 frontAnalog_v0p0p1_3.x65.A.n4 0.154668
R23739 frontAnalog_v0p0p1_3.x65.A frontAnalog_v0p0p1_3.x65.A.n6 0.08175
R23740 frontAnalog_v0p0p1_15.x65.A.n1 frontAnalog_v0p0p1_15.x65.A.t4 260.322
R23741 frontAnalog_v0p0p1_15.x65.A.n4 frontAnalog_v0p0p1_15.x65.A.t7 233.929
R23742 frontAnalog_v0p0p1_15.x65.A.n1 frontAnalog_v0p0p1_15.x65.A.t6 175.169
R23743 frontAnalog_v0p0p1_15.x65.A.n3 frontAnalog_v0p0p1_15.x65.A.t5 160.416
R23744 frontAnalog_v0p0p1_15.x65.A.n2 frontAnalog_v0p0p1_15.x65.A.t3 17.4109
R23745 frontAnalog_v0p0p1_15.x65.A.n2 frontAnalog_v0p0p1_15.x65.A.t2 10.2053
R23746 frontAnalog_v0p0p1_15.x65.A.n0 frontAnalog_v0p0p1_15.x65.A 2.78715
R23747 frontAnalog_v0p0p1_15.x65.A.n0 frontAnalog_v0p0p1_15.x65.A.n1 9.09103
R23748 frontAnalog_v0p0p1_15.x65.A.n6 frontAnalog_v0p0p1_15.x65.A.t1 7.94569
R23749 frontAnalog_v0p0p1_15.x65.A.n3 frontAnalog_v0p0p1_15.x65.A.t0 7.55846
R23750 frontAnalog_v0p0p1_15.x65.A.n5 frontAnalog_v0p0p1_15.x65.A.n4 1.4614
R23751 frontAnalog_v0p0p1_15.x65.A.n4 frontAnalog_v0p0p1_15.x65.A.n3 1.19626
R23752 frontAnalog_v0p0p1_15.x65.A.n6 frontAnalog_v0p0p1_15.x65.A.n5 0.836961
R23753 frontAnalog_v0p0p1_15.x65.A frontAnalog_v0p0p1_15.x65.A.n0 0.390342
R23754 frontAnalog_v0p0p1_15.x65.A.n5 frontAnalog_v0p0p1_15.x65.A.n2 0.154668
R23755 frontAnalog_v0p0p1_15.x65.A frontAnalog_v0p0p1_15.x65.A.n6 0.08175
R23756 frontAnalog_v0p0p1_4.x63.A.n2 frontAnalog_v0p0p1_4.x63.A.t6 260.322
R23757 frontAnalog_v0p0p1_4.x63.A.n4 frontAnalog_v0p0p1_4.x63.A.t4 233.888
R23758 frontAnalog_v0p0p1_4.x63.A.n2 frontAnalog_v0p0p1_4.x63.A.t5 175.169
R23759 frontAnalog_v0p0p1_4.x63.A.n3 frontAnalog_v0p0p1_4.x63.A.t7 159.725
R23760 frontAnalog_v0p0p1_4.x63.A.n1 frontAnalog_v0p0p1_4.x63.A.t3 17.4109
R23761 frontAnalog_v0p0p1_4.x63.A.n0 frontAnalog_v0p0p1_4.x63.A.n2 9.75129
R23762 frontAnalog_v0p0p1_4.x63.A.n1 frontAnalog_v0p0p1_4.x63.A.t2 9.6037
R23763 frontAnalog_v0p0p1_4.x63.A.n0 frontAnalog_v0p0p1_4.x63.A 2.33338
R23764 frontAnalog_v0p0p1_4.x63.A.n5 frontAnalog_v0p0p1_4.x63.A.t1 8.40929
R23765 frontAnalog_v0p0p1_4.x63.A.n3 frontAnalog_v0p0p1_4.x63.A.t0 8.06629
R23766 frontAnalog_v0p0p1_4.x63.A.n4 frontAnalog_v0p0p1_4.x63.A.n3 1.73501
R23767 frontAnalog_v0p0p1_4.x63.A.n1 frontAnalog_v0p0p1_4.x63.A.n4 0.99025
R23768 frontAnalog_v0p0p1_4.x63.A.n5 frontAnalog_v0p0p1_4.x63.A.n1 0.853186
R23769 frontAnalog_v0p0p1_4.x63.A frontAnalog_v0p0p1_4.x63.A.n0 0.349517
R23770 frontAnalog_v0p0p1_4.x63.A frontAnalog_v0p0p1_4.x63.A.n5 0.24425
R23771 frontAnalog_v0p0p1_1.x65.A.n1 frontAnalog_v0p0p1_1.x65.A.t4 260.322
R23772 frontAnalog_v0p0p1_1.x65.A.n3 frontAnalog_v0p0p1_1.x65.A.t7 233.929
R23773 frontAnalog_v0p0p1_1.x65.A.n1 frontAnalog_v0p0p1_1.x65.A.t6 175.169
R23774 frontAnalog_v0p0p1_1.x65.A.n2 frontAnalog_v0p0p1_1.x65.A.t5 160.416
R23775 frontAnalog_v0p0p1_1.x65.A.n4 frontAnalog_v0p0p1_1.x65.A.t0 17.4109
R23776 frontAnalog_v0p0p1_1.x65.A.n4 frontAnalog_v0p0p1_1.x65.A.t1 10.2053
R23777 frontAnalog_v0p0p1_1.x65.A.n0 frontAnalog_v0p0p1_1.x65.A 2.78715
R23778 frontAnalog_v0p0p1_1.x65.A.n0 frontAnalog_v0p0p1_1.x65.A.n1 9.09103
R23779 frontAnalog_v0p0p1_1.x65.A.n6 frontAnalog_v0p0p1_1.x65.A.t2 7.94569
R23780 frontAnalog_v0p0p1_1.x65.A.n2 frontAnalog_v0p0p1_1.x65.A.t3 7.55846
R23781 frontAnalog_v0p0p1_1.x65.A.n5 frontAnalog_v0p0p1_1.x65.A.n3 1.4614
R23782 frontAnalog_v0p0p1_1.x65.A.n3 frontAnalog_v0p0p1_1.x65.A.n2 1.19626
R23783 frontAnalog_v0p0p1_1.x65.A.n6 frontAnalog_v0p0p1_1.x65.A.n5 0.836961
R23784 frontAnalog_v0p0p1_1.x65.A frontAnalog_v0p0p1_1.x65.A.n0 0.390342
R23785 frontAnalog_v0p0p1_1.x65.A.n5 frontAnalog_v0p0p1_1.x65.A.n4 0.154668
R23786 frontAnalog_v0p0p1_1.x65.A frontAnalog_v0p0p1_1.x65.A.n6 0.08175
R23787 frontAnalog_v0p0p1_10.RSfetsym_0.QN.n1 frontAnalog_v0p0p1_10.RSfetsym_0.QN.t6 117.511
R23788 frontAnalog_v0p0p1_10.RSfetsym_0.QN.n1 frontAnalog_v0p0p1_10.RSfetsym_0.QN.t5 110.698
R23789 frontAnalog_v0p0p1_10.RSfetsym_0.QN.n2 frontAnalog_v0p0p1_10.RSfetsym_0.QN.t2 19.1963
R23790 frontAnalog_v0p0p1_10.RSfetsym_0.QN.n3 frontAnalog_v0p0p1_10.RSfetsym_0.QN.t0 14.5206
R23791 frontAnalog_v0p0p1_10.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_10.RSfetsym_0.QN.t3 14.283
R23792 frontAnalog_v0p0p1_10.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_10.RSfetsym_0.QN.t4 14.283
R23793 frontAnalog_v0p0p1_10.RSfetsym_0.QN frontAnalog_v0p0p1_10.RSfetsym_0.QN.t1 9.14075
R23794 frontAnalog_v0p0p1_10.RSfetsym_0.QN.n2 frontAnalog_v0p0p1_10.RSfetsym_0.QN.n1 0.826818
R23795 frontAnalog_v0p0p1_10.RSfetsym_0.QN frontAnalog_v0p0p1_10.RSfetsym_0.QN.n0 0.74645
R23796 frontAnalog_v0p0p1_10.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_10.RSfetsym_0.QN.n3 0.249509
R23797 frontAnalog_v0p0p1_10.RSfetsym_0.QN.n3 frontAnalog_v0p0p1_10.RSfetsym_0.QN.n2 0.0968646
R23798 I4.n2 I4.t5 260.435
R23799 I4.n7 I4.t11 230.576
R23800 I4.n10 I4.t7 196.549
R23801 I4.n7 I4.t8 158.275
R23802 I4.n2 I4.t10 156.403
R23803 I4.n10 I4.t9 148.35
R23804 I4.n15 I4.t6 117.314
R23805 I4.n15 I4.t12 110.853
R23806 I4.n17 I4.t0 17.6181
R23807 I4.n18 I4.t3 14.2865
R23808 I4.n20 I4.t2 14.283
R23809 I4.n20 I4.t1 14.283
R23810 I4.n11 I4.n10 9.49829
R23811 I4 I4.n1 9.3005
R23812 I4.n22 I4.t4 8.77744
R23813 I4.n8 I4.n7 8.76429
R23814 I4.n12 I4.n11 7.9582
R23815 I4.n9 I4.n8 7.74345
R23816 I4.n3 I4.n2 7.60183
R23817 I4.n8 I4 6.66717
R23818 I4.n11 I4 6.44139
R23819 I4.n3 I4 4.8645
R23820 I4.n4 I4.n0 4.54557
R23821 I4.n1 I4.n0 4.51121
R23822 I4 I4.n23 4.47065
R23823 I4.n13 I4.n6 2.33148
R23824 I4.n22 I4.n21 1.20426
R23825 I4.n12 I4.n9 1.0005
R23826 I4.n24 I4 0.509667
R23827 I4 I4.n14 0.4987
R23828 I4.n13 I4.n12 0.446956
R23829 I4 I4.n24 0.382375
R23830 I4.n9 I4 0.380411
R23831 I4.n14 I4.n13 0.368862
R23832 I4.n23 I4.n22 0.32511
R23833 I4.n18 I4.n17 0.314673
R23834 I4.n19 I4.n18 0.299251
R23835 I4.n14 I4 0.20675
R23836 I4.n16 I4.n15 0.159555
R23837 I4.n21 I4.n20 0.106617
R23838 I4.n19 I4.n16 0.0796167
R23839 I4.n21 I4.n19 0.0480595
R23840 I4.n23 I4 0.046937
R23841 I4.n5 I4.n1 0.0344286
R23842 I4.n24 I4 0.0161667
R23843 I4.n24 I4 0.01225
R23844 I4.n6 I4.n0 0.00182856
R23845 I4.n6 I4.n5 0.00149885
R23846 I4.n4 I4.n3 0.00133362
R23847 I4.n5 I4.n4 0.00100077
R23848 I4.n17 I4.n16 0.000504658
R23849 frontAnalog_v0p0p1_3.RSfetsym_0.QN.n1 frontAnalog_v0p0p1_3.RSfetsym_0.QN.t6 117.511
R23850 frontAnalog_v0p0p1_3.RSfetsym_0.QN.n1 frontAnalog_v0p0p1_3.RSfetsym_0.QN.t5 110.698
R23851 frontAnalog_v0p0p1_3.RSfetsym_0.QN.n2 frontAnalog_v0p0p1_3.RSfetsym_0.QN.t2 19.1963
R23852 frontAnalog_v0p0p1_3.RSfetsym_0.QN.n3 frontAnalog_v0p0p1_3.RSfetsym_0.QN.t0 14.5206
R23853 frontAnalog_v0p0p1_3.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_3.RSfetsym_0.QN.t3 14.283
R23854 frontAnalog_v0p0p1_3.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_3.RSfetsym_0.QN.t4 14.283
R23855 frontAnalog_v0p0p1_3.RSfetsym_0.QN frontAnalog_v0p0p1_3.RSfetsym_0.QN.t1 9.14075
R23856 frontAnalog_v0p0p1_3.RSfetsym_0.QN.n2 frontAnalog_v0p0p1_3.RSfetsym_0.QN.n1 0.826818
R23857 frontAnalog_v0p0p1_3.RSfetsym_0.QN frontAnalog_v0p0p1_3.RSfetsym_0.QN.n0 0.74645
R23858 frontAnalog_v0p0p1_3.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_3.RSfetsym_0.QN.n3 0.249509
R23859 frontAnalog_v0p0p1_3.RSfetsym_0.QN.n3 frontAnalog_v0p0p1_3.RSfetsym_0.QN.n2 0.0968646
R23860 frontAnalog_v0p0p1_6.x63.A.n2 frontAnalog_v0p0p1_6.x63.A.t4 260.322
R23861 frontAnalog_v0p0p1_6.x63.A.n4 frontAnalog_v0p0p1_6.x63.A.t7 233.888
R23862 frontAnalog_v0p0p1_6.x63.A.n2 frontAnalog_v0p0p1_6.x63.A.t6 175.169
R23863 frontAnalog_v0p0p1_6.x63.A.n3 frontAnalog_v0p0p1_6.x63.A.t5 159.725
R23864 frontAnalog_v0p0p1_6.x63.A.n1 frontAnalog_v0p0p1_6.x63.A.t1 17.4109
R23865 frontAnalog_v0p0p1_6.x63.A.n0 frontAnalog_v0p0p1_6.x63.A.n2 9.75129
R23866 frontAnalog_v0p0p1_6.x63.A.n1 frontAnalog_v0p0p1_6.x63.A.t0 9.6027
R23867 frontAnalog_v0p0p1_6.x63.A.n0 frontAnalog_v0p0p1_6.x63.A 2.33338
R23868 frontAnalog_v0p0p1_6.x63.A.n5 frontAnalog_v0p0p1_6.x63.A.t3 8.40929
R23869 frontAnalog_v0p0p1_6.x63.A.n3 frontAnalog_v0p0p1_6.x63.A.t2 8.06629
R23870 frontAnalog_v0p0p1_6.x63.A.n4 frontAnalog_v0p0p1_6.x63.A.n3 1.73501
R23871 frontAnalog_v0p0p1_6.x63.A.n1 frontAnalog_v0p0p1_6.x63.A.n4 0.99025
R23872 frontAnalog_v0p0p1_6.x63.A.n5 frontAnalog_v0p0p1_6.x63.A.n1 0.853186
R23873 frontAnalog_v0p0p1_6.x63.A frontAnalog_v0p0p1_6.x63.A.n0 0.349517
R23874 frontAnalog_v0p0p1_6.x63.A frontAnalog_v0p0p1_6.x63.A.n5 0.24425
R23875 frontAnalog_v0p0p1_12.RSfetsym_0.QN.n1 frontAnalog_v0p0p1_12.RSfetsym_0.QN.t6 117.511
R23876 frontAnalog_v0p0p1_12.RSfetsym_0.QN.n1 frontAnalog_v0p0p1_12.RSfetsym_0.QN.t5 110.698
R23877 frontAnalog_v0p0p1_12.RSfetsym_0.QN.n2 frontAnalog_v0p0p1_12.RSfetsym_0.QN.t0 19.1963
R23878 frontAnalog_v0p0p1_12.RSfetsym_0.QN.n3 frontAnalog_v0p0p1_12.RSfetsym_0.QN.t4 14.5206
R23879 frontAnalog_v0p0p1_12.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_12.RSfetsym_0.QN.t2 14.283
R23880 frontAnalog_v0p0p1_12.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_12.RSfetsym_0.QN.t1 14.283
R23881 frontAnalog_v0p0p1_12.RSfetsym_0.QN frontAnalog_v0p0p1_12.RSfetsym_0.QN.t3 9.14075
R23882 frontAnalog_v0p0p1_12.RSfetsym_0.QN.n2 frontAnalog_v0p0p1_12.RSfetsym_0.QN.n1 0.826818
R23883 frontAnalog_v0p0p1_12.RSfetsym_0.QN frontAnalog_v0p0p1_12.RSfetsym_0.QN.n0 0.74645
R23884 frontAnalog_v0p0p1_12.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_12.RSfetsym_0.QN.n3 0.249509
R23885 frontAnalog_v0p0p1_12.RSfetsym_0.QN.n3 frontAnalog_v0p0p1_12.RSfetsym_0.QN.n2 0.0968646
R23886 VL.n6 VL 0.23241
R23887 VL.n3 VL.t2 0.0203551
R23888 VL.n0 VL.t5 0.0203551
R23889 VL.n1 VL.n0 0.0203529
R23890 VL.n2 VL.n1 0.0203529
R23891 VL.n5 VL.n4 0.0203529
R23892 VL.n4 VL.n3 0.0203529
R23893 VL VL.n2 0.0111618
R23894 VL VL.n6 0.00913171
R23895 VL.n6 VL.n5 0.00105946
R23896 VL.n3 VL.t0 0.000502142
R23897 VL.n4 VL.t4 0.000502142
R23898 VL.n5 VL.t3 0.000502142
R23899 VL.n2 VL.t7 0.000502142
R23900 VL.n1 VL.t6 0.000502142
R23901 VL.n0 VL.t1 0.000502142
R23902 frontAnalog_v0p0p1_11.x65.A.n1 frontAnalog_v0p0p1_11.x65.A.t4 260.322
R23903 frontAnalog_v0p0p1_11.x65.A.n3 frontAnalog_v0p0p1_11.x65.A.t7 233.929
R23904 frontAnalog_v0p0p1_11.x65.A.n1 frontAnalog_v0p0p1_11.x65.A.t6 175.169
R23905 frontAnalog_v0p0p1_11.x65.A.n2 frontAnalog_v0p0p1_11.x65.A.t5 160.416
R23906 frontAnalog_v0p0p1_11.x65.A.n4 frontAnalog_v0p0p1_11.x65.A.t1 17.4109
R23907 frontAnalog_v0p0p1_11.x65.A.n4 frontAnalog_v0p0p1_11.x65.A.t0 10.2053
R23908 frontAnalog_v0p0p1_11.x65.A.n0 frontAnalog_v0p0p1_11.x65.A 2.78715
R23909 frontAnalog_v0p0p1_11.x65.A.n0 frontAnalog_v0p0p1_11.x65.A.n1 9.09103
R23910 frontAnalog_v0p0p1_11.x65.A.n6 frontAnalog_v0p0p1_11.x65.A.t2 7.94569
R23911 frontAnalog_v0p0p1_11.x65.A.n2 frontAnalog_v0p0p1_11.x65.A.t3 7.55846
R23912 frontAnalog_v0p0p1_11.x65.A.n5 frontAnalog_v0p0p1_11.x65.A.n3 1.4614
R23913 frontAnalog_v0p0p1_11.x65.A.n3 frontAnalog_v0p0p1_11.x65.A.n2 1.19626
R23914 frontAnalog_v0p0p1_11.x65.A.n6 frontAnalog_v0p0p1_11.x65.A.n5 0.836961
R23915 frontAnalog_v0p0p1_11.x65.A frontAnalog_v0p0p1_11.x65.A.n0 0.390342
R23916 frontAnalog_v0p0p1_11.x65.A.n5 frontAnalog_v0p0p1_11.x65.A.n4 0.154668
R23917 frontAnalog_v0p0p1_11.x65.A frontAnalog_v0p0p1_11.x65.A.n6 0.08175
R23918 VV8.n0 VV8.t17 167.365
R23919 VV8.n0 VV8.t16 92.4488
R23920 VV8.n1 VV8.n0 2.07493
R23921 VV8.n10 VV8 0.431333
R23922 VV8 VV8.n10 0.323625
R23923 VV8.n9 VV8.n8 0.141636
R23924 VV8.n8 VV8.n7 0.141636
R23925 VV8.n7 VV8.n6 0.141636
R23926 VV8.n6 VV8.n5 0.141636
R23927 VV8.n5 VV8.n4 0.141636
R23928 VV8.n4 VV8.n3 0.141636
R23929 VV8.n3 VV8.n2 0.141636
R23930 VV8.n1 VV8 0.12425
R23931 VV8 VV8.n9 0.100159
R23932 VV8 VV8.n1 0.0314375
R23933 VV8.n10 VV8 0.00833333
R23934 VV8.n10 VV8 0.006375
R23935 VV8.n3 VV8.t0 0.000502142
R23936 VV8.n4 VV8.t3 0.000502142
R23937 VV8.n5 VV8.t4 0.000502142
R23938 VV8.n6 VV8.t8 0.000502142
R23939 VV8.n7 VV8.t7 0.000502142
R23940 VV8.n8 VV8.t9 0.000502142
R23941 VV8.n9 VV8.t15 0.000502142
R23942 VV8.n2 VV8.t2 0.000502142
R23943 VV8.n3 VV8.t11 0.000502142
R23944 VV8.n4 VV8.t5 0.000502142
R23945 VV8.n5 VV8.t12 0.000502142
R23946 VV8.n6 VV8.t1 0.000502142
R23947 VV8.n7 VV8.t13 0.000502142
R23948 VV8.n8 VV8.t14 0.000502142
R23949 VV8.n9 VV8.t10 0.000502142
R23950 VV8.n2 VV8.t6 0.000502142
R23951 I12.n2 I12.t11 260.435
R23952 I12.n7 I12.t12 230.576
R23953 I12.n10 I12.t6 196.549
R23954 I12.n7 I12.t9 158.275
R23955 I12.n2 I12.t8 156.403
R23956 I12.n10 I12.t5 148.35
R23957 I12.n17 I12.t10 117.314
R23958 I12.n17 I12.t7 110.852
R23959 I12.n19 I12.t1 17.6181
R23960 I12.n20 I12.t4 14.2865
R23961 I12.n22 I12.t3 14.283
R23962 I12.n22 I12.t2 14.283
R23963 I12.n11 I12.n10 9.49829
R23964 I12 I12.n1 9.3005
R23965 I12.n24 I12.t0 8.77592
R23966 I12.n8 I12.n7 8.76429
R23967 I12.n12 I12.n11 7.9582
R23968 I12.n9 I12.n8 7.74345
R23969 I12.n3 I12.n2 7.60183
R23970 I12.n8 I12 6.66717
R23971 I12.n11 I12 6.44139
R23972 I12.n3 I12 4.8645
R23973 I12.n4 I12.n0 4.54557
R23974 I12.n1 I12.n0 4.51121
R23975 I12 I12.n25 3.93116
R23976 I12.n13 I12.n6 2.33638
R23977 I12.n24 I12.n23 1.20426
R23978 I12.n12 I12.n9 1.0005
R23979 I12.n26 I12 0.992722
R23980 I12.n14 I12 0.979667
R23981 I12 I12.n16 0.917
R23982 I12.n16 I12 0.82535
R23983 I12 I12.n26 0.447
R23984 I12.n13 I12.n12 0.446956
R23985 I12.n9 I12 0.380411
R23986 I12.n14 I12.n13 0.356917
R23987 I12.n25 I12.n24 0.336084
R23988 I12.n20 I12.n19 0.314673
R23989 I12.n21 I12.n20 0.300251
R23990 I12.n15 I12 0.2005
R23991 I12.n18 I12.n17 0.159555
R23992 I12.n23 I12.n22 0.106617
R23993 I12.n21 I12.n18 0.0796167
R23994 I12.n23 I12.n21 0.0480595
R23995 I12.n5 I12.n1 0.0344286
R23996 I12.n15 I12.n14 0.0287
R23997 I12.n16 I12.n15 0.0287
R23998 I12.n26 I12 0.0266111
R23999 I12.n26 I12 0.01225
R24000 I12.n25 I12 0.00658123
R24001 I12.n6 I12.n0 0.00182856
R24002 I12.n6 I12.n5 0.00149885
R24003 I12.n4 I12.n3 0.00133362
R24004 I12.n5 I12.n4 0.00100077
R24005 I12.n19 I12.n18 0.000504658
R24006 frontAnalog_v0p0p1_1.x63.A.n2 frontAnalog_v0p0p1_1.x63.A.t7 260.322
R24007 frontAnalog_v0p0p1_1.x63.A.n4 frontAnalog_v0p0p1_1.x63.A.t4 233.888
R24008 frontAnalog_v0p0p1_1.x63.A.n2 frontAnalog_v0p0p1_1.x63.A.t6 175.169
R24009 frontAnalog_v0p0p1_1.x63.A.n3 frontAnalog_v0p0p1_1.x63.A.t5 159.725
R24010 frontAnalog_v0p0p1_1.x63.A.n1 frontAnalog_v0p0p1_1.x63.A.t0 17.4109
R24011 frontAnalog_v0p0p1_1.x63.A.n0 frontAnalog_v0p0p1_1.x63.A.n2 9.75129
R24012 frontAnalog_v0p0p1_1.x63.A.n1 frontAnalog_v0p0p1_1.x63.A.t1 9.6027
R24013 frontAnalog_v0p0p1_1.x63.A.n0 frontAnalog_v0p0p1_1.x63.A 2.33338
R24014 frontAnalog_v0p0p1_1.x63.A.n5 frontAnalog_v0p0p1_1.x63.A.t2 8.40929
R24015 frontAnalog_v0p0p1_1.x63.A.n3 frontAnalog_v0p0p1_1.x63.A.t3 8.06629
R24016 frontAnalog_v0p0p1_1.x63.A.n4 frontAnalog_v0p0p1_1.x63.A.n3 1.73501
R24017 frontAnalog_v0p0p1_1.x63.A.n1 frontAnalog_v0p0p1_1.x63.A.n4 0.99025
R24018 frontAnalog_v0p0p1_1.x63.A.n5 frontAnalog_v0p0p1_1.x63.A.n1 0.853186
R24019 frontAnalog_v0p0p1_1.x63.A frontAnalog_v0p0p1_1.x63.A.n0 0.349517
R24020 frontAnalog_v0p0p1_1.x63.A frontAnalog_v0p0p1_1.x63.A.n5 0.24425
R24021 frontAnalog_v0p0p1_5.x65.A.n1 frontAnalog_v0p0p1_5.x65.A.t4 260.322
R24022 frontAnalog_v0p0p1_5.x65.A.n4 frontAnalog_v0p0p1_5.x65.A.t7 233.929
R24023 frontAnalog_v0p0p1_5.x65.A.n1 frontAnalog_v0p0p1_5.x65.A.t6 175.169
R24024 frontAnalog_v0p0p1_5.x65.A.n3 frontAnalog_v0p0p1_5.x65.A.t5 160.416
R24025 frontAnalog_v0p0p1_5.x65.A.n2 frontAnalog_v0p0p1_5.x65.A.t3 17.4109
R24026 frontAnalog_v0p0p1_5.x65.A.n2 frontAnalog_v0p0p1_5.x65.A.t2 10.2053
R24027 frontAnalog_v0p0p1_5.x65.A.n0 frontAnalog_v0p0p1_5.x65.A 2.78715
R24028 frontAnalog_v0p0p1_5.x65.A.n0 frontAnalog_v0p0p1_5.x65.A.n1 9.09103
R24029 frontAnalog_v0p0p1_5.x65.A.n6 frontAnalog_v0p0p1_5.x65.A.t1 7.94569
R24030 frontAnalog_v0p0p1_5.x65.A.n3 frontAnalog_v0p0p1_5.x65.A.t0 7.55846
R24031 frontAnalog_v0p0p1_5.x65.A.n5 frontAnalog_v0p0p1_5.x65.A.n4 1.4614
R24032 frontAnalog_v0p0p1_5.x65.A.n4 frontAnalog_v0p0p1_5.x65.A.n3 1.19626
R24033 frontAnalog_v0p0p1_5.x65.A.n6 frontAnalog_v0p0p1_5.x65.A.n5 0.836961
R24034 frontAnalog_v0p0p1_5.x65.A frontAnalog_v0p0p1_5.x65.A.n0 0.390342
R24035 frontAnalog_v0p0p1_5.x65.A.n5 frontAnalog_v0p0p1_5.x65.A.n2 0.154668
R24036 frontAnalog_v0p0p1_5.x65.A frontAnalog_v0p0p1_5.x65.A.n6 0.08175
R24037 frontAnalog_v0p0p1_14.RSfetsym_0.QN.n2 frontAnalog_v0p0p1_14.RSfetsym_0.QN.t6 117.511
R24038 frontAnalog_v0p0p1_14.RSfetsym_0.QN.n2 frontAnalog_v0p0p1_14.RSfetsym_0.QN.t5 110.698
R24039 frontAnalog_v0p0p1_14.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_14.RSfetsym_0.QN.t3 19.1963
R24040 frontAnalog_v0p0p1_14.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_14.RSfetsym_0.QN.t0 14.5206
R24041 frontAnalog_v0p0p1_14.RSfetsym_0.QN.n1 frontAnalog_v0p0p1_14.RSfetsym_0.QN.t4 14.283
R24042 frontAnalog_v0p0p1_14.RSfetsym_0.QN.n1 frontAnalog_v0p0p1_14.RSfetsym_0.QN.t1 14.283
R24043 frontAnalog_v0p0p1_14.RSfetsym_0.QN frontAnalog_v0p0p1_14.RSfetsym_0.QN.t2 9.13975
R24044 frontAnalog_v0p0p1_14.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_14.RSfetsym_0.QN.n2 0.826818
R24045 frontAnalog_v0p0p1_14.RSfetsym_0.QN frontAnalog_v0p0p1_14.RSfetsym_0.QN.n1 0.74645
R24046 frontAnalog_v0p0p1_14.RSfetsym_0.QN.n1 frontAnalog_v0p0p1_14.RSfetsym_0.QN.n0 0.34588
R24047 frontAnalog_v0p0p1_7.RSfetsym_0.QN.n1 frontAnalog_v0p0p1_7.RSfetsym_0.QN.t6 117.511
R24048 frontAnalog_v0p0p1_7.RSfetsym_0.QN.n1 frontAnalog_v0p0p1_7.RSfetsym_0.QN.t5 110.698
R24049 frontAnalog_v0p0p1_7.RSfetsym_0.QN.n2 frontAnalog_v0p0p1_7.RSfetsym_0.QN.t1 19.1963
R24050 frontAnalog_v0p0p1_7.RSfetsym_0.QN.n3 frontAnalog_v0p0p1_7.RSfetsym_0.QN.t4 14.5206
R24051 frontAnalog_v0p0p1_7.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_7.RSfetsym_0.QN.t2 14.283
R24052 frontAnalog_v0p0p1_7.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_7.RSfetsym_0.QN.t3 14.283
R24053 frontAnalog_v0p0p1_7.RSfetsym_0.QN frontAnalog_v0p0p1_7.RSfetsym_0.QN.t0 9.14075
R24054 frontAnalog_v0p0p1_7.RSfetsym_0.QN.n2 frontAnalog_v0p0p1_7.RSfetsym_0.QN.n1 0.826818
R24055 frontAnalog_v0p0p1_7.RSfetsym_0.QN frontAnalog_v0p0p1_7.RSfetsym_0.QN.n0 0.74645
R24056 frontAnalog_v0p0p1_7.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_7.RSfetsym_0.QN.n3 0.249509
R24057 frontAnalog_v0p0p1_7.RSfetsym_0.QN.n3 frontAnalog_v0p0p1_7.RSfetsym_0.QN.n2 0.0968646
R24058 frontAnalog_v0p0p1_0.RSfetsym_0.QN.n1 frontAnalog_v0p0p1_0.RSfetsym_0.QN.t5 117.511
R24059 frontAnalog_v0p0p1_0.RSfetsym_0.QN.n1 frontAnalog_v0p0p1_0.RSfetsym_0.QN.t6 110.698
R24060 frontAnalog_v0p0p1_0.RSfetsym_0.QN.n2 frontAnalog_v0p0p1_0.RSfetsym_0.QN.t1 19.1963
R24061 frontAnalog_v0p0p1_0.RSfetsym_0.QN.n3 frontAnalog_v0p0p1_0.RSfetsym_0.QN.t4 14.5206
R24062 frontAnalog_v0p0p1_0.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_0.RSfetsym_0.QN.t3 14.283
R24063 frontAnalog_v0p0p1_0.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_0.RSfetsym_0.QN.t2 14.283
R24064 frontAnalog_v0p0p1_0.RSfetsym_0.QN frontAnalog_v0p0p1_0.RSfetsym_0.QN.t0 9.14075
R24065 frontAnalog_v0p0p1_0.RSfetsym_0.QN.n2 frontAnalog_v0p0p1_0.RSfetsym_0.QN.n1 0.826818
R24066 frontAnalog_v0p0p1_0.RSfetsym_0.QN frontAnalog_v0p0p1_0.RSfetsym_0.QN.n0 0.74645
R24067 frontAnalog_v0p0p1_0.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_0.RSfetsym_0.QN.n3 0.249509
R24068 frontAnalog_v0p0p1_0.RSfetsym_0.QN.n3 frontAnalog_v0p0p1_0.RSfetsym_0.QN.n2 0.0968646
R24069 I8.n0 I8.t8 196.549
R24070 I8.n0 I8.t6 148.35
R24071 I8.n4 I8.t7 117.314
R24072 I8.n4 I8.t5 110.853
R24073 I8.n6 I8.t2 17.6181
R24074 I8.n7 I8.t1 14.2865
R24075 I8.n9 I8.t3 14.283
R24076 I8.n9 I8.t4 14.283
R24077 I8.n1 I8.n0 9.49592
R24078 I8.n11 I8.t0 8.77744
R24079 I8.n2 I8.n1 7.58085
R24080 I8.n1 I8 6.44187
R24081 I8.n3 I8.n2 2.34543
R24082 I8.n11 I8.n10 1.20426
R24083 I8.n2 I8 0.88934
R24084 I8 I8.n11 0.357737
R24085 I8 I8.n3 0.336158
R24086 I8.n7 I8.n6 0.314673
R24087 I8.n8 I8.n7 0.299251
R24088 I8.n3 I8 0.200892
R24089 I8.n5 I8.n4 0.159555
R24090 I8.n10 I8.n9 0.106617
R24091 I8.n8 I8.n5 0.0796167
R24092 I8.n10 I8.n8 0.0480595
R24093 I8.n6 I8.n5 0.000504658
R24094 S1.n0 S1.t5 259.192
R24095 S1.n34 S1.t10 258.584
R24096 S1.n39 S1.t1 222.243
R24097 S1.n13 S1.t2 212.081
R24098 S1.n8 S1.t3 212.081
R24099 S1.n7 S1.t7 212.081
R24100 S1.n4 S1.t8 212.081
R24101 S1.n13 S1.t4 139.78
R24102 S1.n8 S1.t6 139.78
R24103 S1.n7 S1.t11 139.78
R24104 S1.n4 S1.t12 139.78
R24105 S1.n40 S1.t0 123.654
R24106 S1.n35 S1.t9 117.346
R24107 S1.n41 S1.n40 43.0815
R24108 S1.n41 S1 32.4695
R24109 S1.n6 S1.n4 30.6732
R24110 S1.n9 S1.n7 30.6732
R24111 S1.n9 S1.n8 30.6732
R24112 S1.n14 S1.n13 30.6732
R24113 S1.n26 S1.n25 12.8005
R24114 S1.n6 S1.n5 12.4157
R24115 S1 S1.n39 10.4848
R24116 S1.n32 S1.n31 9.3005
R24117 S1.n21 S1.n20 9.3005
R24118 S1.n24 S1.n9 8.28655
R24119 S1.n16 S1.n14 8.28655
R24120 S1.n27 S1.n6 8.28655
R24121 S1.n39 S1 5.50526
R24122 S1.n40 S1 5.16973
R24123 S1.n25 S1.n24 4.3525
R24124 S1.n17 S1.n12 4.3525
R24125 S1.n15 S1 4.10475
R24126 S1.n28 S1.n3 4.0965
R24127 S1.n23 S1 3.8405
R24128 S1 S1.n1 2.3045
R24129 S1.n31 S1 2.3045
R24130 S1.n27 S1 2.3045
R24131 S1 S1.n26 2.0485
R24132 S1.n42 S1.n41 1.94684
R24133 S1.n36 S1.n33 1.85764
R24134 S1.n16 S1.n15 1.15434
R24135 S1.n28 S1.n27 1.0245
R24136 S1.n20 S1 0.7685
R24137 S1.n24 S1.n23 0.5125
R24138 S1.n17 S1.n16 0.5125
R24139 S1.n33 S1.n1 0.462934
R24140 S1.n37 S1.n36 0.429669
R24141 S1.n37 S1.n0 0.230918
R24142 S1 S1.n43 0.207965
R24143 S1.n35 S1.n34 0.12975
R24144 S1.n43 S1 0.101429
R24145 S1.n43 S1.n42 0.0907778
R24146 S1.n42 S1 0.0847014
R24147 S1.n10 S1.n2 0.0766364
R24148 S1.n32 S1.n30 0.0618636
R24149 S1.n38 S1.n37 0.0592506
R24150 S1.n43 S1.n38 0.0591993
R24151 S1.n21 S1.n19 0.0516364
R24152 S1.n38 S1 0.0266824
R24153 S1.n33 S1.n32 0.0239512
R24154 S1.n22 S1.n21 0.0209545
R24155 S1.n11 S1.n10 0.0198182
R24156 S1.n19 S1.n18 0.0198182
R24157 S1.n30 S1.n29 0.0186818
R24158 S1.n29 S1.n2 0.00504545
R24159 S1.n36 S1.n35 0.0028536
R24160 S1.n22 S1.n11 0.00277273
R24161 S1.n29 S1.n28 0.00119114
R24162 S1.n23 S1.n22 0.00119114
R24163 S1.n18 S1.n17 0.00119114
R24164 frontAnalog_v0p0p1_13.x65.A.n1 frontAnalog_v0p0p1_13.x65.A.t4 260.322
R24165 frontAnalog_v0p0p1_13.x65.A.n4 frontAnalog_v0p0p1_13.x65.A.t7 233.929
R24166 frontAnalog_v0p0p1_13.x65.A.n1 frontAnalog_v0p0p1_13.x65.A.t6 175.169
R24167 frontAnalog_v0p0p1_13.x65.A.n3 frontAnalog_v0p0p1_13.x65.A.t5 160.416
R24168 frontAnalog_v0p0p1_13.x65.A.n2 frontAnalog_v0p0p1_13.x65.A.t3 17.4109
R24169 frontAnalog_v0p0p1_13.x65.A.n2 frontAnalog_v0p0p1_13.x65.A.t2 10.2053
R24170 frontAnalog_v0p0p1_13.x65.A.n0 frontAnalog_v0p0p1_13.x65.A 2.78715
R24171 frontAnalog_v0p0p1_13.x65.A.n0 frontAnalog_v0p0p1_13.x65.A.n1 9.09103
R24172 frontAnalog_v0p0p1_13.x65.A.n6 frontAnalog_v0p0p1_13.x65.A.t1 7.94569
R24173 frontAnalog_v0p0p1_13.x65.A.n3 frontAnalog_v0p0p1_13.x65.A.t0 7.55846
R24174 frontAnalog_v0p0p1_13.x65.A.n5 frontAnalog_v0p0p1_13.x65.A.n4 1.4614
R24175 frontAnalog_v0p0p1_13.x65.A.n4 frontAnalog_v0p0p1_13.x65.A.n3 1.19626
R24176 frontAnalog_v0p0p1_13.x65.A.n6 frontAnalog_v0p0p1_13.x65.A.n5 0.836961
R24177 frontAnalog_v0p0p1_13.x65.A frontAnalog_v0p0p1_13.x65.A.n0 0.390342
R24178 frontAnalog_v0p0p1_13.x65.A.n5 frontAnalog_v0p0p1_13.x65.A.n2 0.154668
R24179 frontAnalog_v0p0p1_13.x65.A frontAnalog_v0p0p1_13.x65.A.n6 0.08175
R24180 frontAnalog_v0p0p1_11.RSfetsym_0.QN.n1 frontAnalog_v0p0p1_11.RSfetsym_0.QN.t6 117.511
R24181 frontAnalog_v0p0p1_11.RSfetsym_0.QN.n1 frontAnalog_v0p0p1_11.RSfetsym_0.QN.t5 110.698
R24182 frontAnalog_v0p0p1_11.RSfetsym_0.QN.n2 frontAnalog_v0p0p1_11.RSfetsym_0.QN.t2 19.1963
R24183 frontAnalog_v0p0p1_11.RSfetsym_0.QN.n3 frontAnalog_v0p0p1_11.RSfetsym_0.QN.t4 14.5206
R24184 frontAnalog_v0p0p1_11.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_11.RSfetsym_0.QN.t0 14.283
R24185 frontAnalog_v0p0p1_11.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_11.RSfetsym_0.QN.t1 14.283
R24186 frontAnalog_v0p0p1_11.RSfetsym_0.QN frontAnalog_v0p0p1_11.RSfetsym_0.QN.t3 9.14075
R24187 frontAnalog_v0p0p1_11.RSfetsym_0.QN.n2 frontAnalog_v0p0p1_11.RSfetsym_0.QN.n1 0.826818
R24188 frontAnalog_v0p0p1_11.RSfetsym_0.QN frontAnalog_v0p0p1_11.RSfetsym_0.QN.n0 0.74645
R24189 frontAnalog_v0p0p1_11.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_11.RSfetsym_0.QN.n3 0.249509
R24190 frontAnalog_v0p0p1_11.RSfetsym_0.QN.n3 frontAnalog_v0p0p1_11.RSfetsym_0.QN.n2 0.0968646
R24191 frontAnalog_v0p0p1_12.x63.A.n2 frontAnalog_v0p0p1_12.x63.A.t4 260.322
R24192 frontAnalog_v0p0p1_12.x63.A.n4 frontAnalog_v0p0p1_12.x63.A.t5 233.888
R24193 frontAnalog_v0p0p1_12.x63.A.n2 frontAnalog_v0p0p1_12.x63.A.t6 175.169
R24194 frontAnalog_v0p0p1_12.x63.A.n3 frontAnalog_v0p0p1_12.x63.A.t7 159.725
R24195 frontAnalog_v0p0p1_12.x63.A.n1 frontAnalog_v0p0p1_12.x63.A.t1 17.4109
R24196 frontAnalog_v0p0p1_12.x63.A.n0 frontAnalog_v0p0p1_12.x63.A.n2 9.75129
R24197 frontAnalog_v0p0p1_12.x63.A.n1 frontAnalog_v0p0p1_12.x63.A.t0 9.6027
R24198 frontAnalog_v0p0p1_12.x63.A.n0 frontAnalog_v0p0p1_12.x63.A 2.33338
R24199 frontAnalog_v0p0p1_12.x63.A.n5 frontAnalog_v0p0p1_12.x63.A.t3 8.40929
R24200 frontAnalog_v0p0p1_12.x63.A.n3 frontAnalog_v0p0p1_12.x63.A.t2 8.06629
R24201 frontAnalog_v0p0p1_12.x63.A.n4 frontAnalog_v0p0p1_12.x63.A.n3 1.73501
R24202 frontAnalog_v0p0p1_12.x63.A.n1 frontAnalog_v0p0p1_12.x63.A.n4 0.99025
R24203 frontAnalog_v0p0p1_12.x63.A.n5 frontAnalog_v0p0p1_12.x63.A.n1 0.853186
R24204 frontAnalog_v0p0p1_12.x63.A frontAnalog_v0p0p1_12.x63.A.n0 0.349517
R24205 frontAnalog_v0p0p1_12.x63.A frontAnalog_v0p0p1_12.x63.A.n5 0.24425
R24206 frontAnalog_v0p0p1_4.RSfetsym_0.QN.n1 frontAnalog_v0p0p1_4.RSfetsym_0.QN.t6 117.511
R24207 frontAnalog_v0p0p1_4.RSfetsym_0.QN.n1 frontAnalog_v0p0p1_4.RSfetsym_0.QN.t5 110.698
R24208 frontAnalog_v0p0p1_4.RSfetsym_0.QN.n2 frontAnalog_v0p0p1_4.RSfetsym_0.QN.t4 19.1963
R24209 frontAnalog_v0p0p1_4.RSfetsym_0.QN.n3 frontAnalog_v0p0p1_4.RSfetsym_0.QN.t1 14.5206
R24210 frontAnalog_v0p0p1_4.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_4.RSfetsym_0.QN.t2 14.283
R24211 frontAnalog_v0p0p1_4.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_4.RSfetsym_0.QN.t3 14.283
R24212 frontAnalog_v0p0p1_4.RSfetsym_0.QN frontAnalog_v0p0p1_4.RSfetsym_0.QN.t0 9.14075
R24213 frontAnalog_v0p0p1_4.RSfetsym_0.QN.n2 frontAnalog_v0p0p1_4.RSfetsym_0.QN.n1 0.826818
R24214 frontAnalog_v0p0p1_4.RSfetsym_0.QN frontAnalog_v0p0p1_4.RSfetsym_0.QN.n0 0.74645
R24215 frontAnalog_v0p0p1_4.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_4.RSfetsym_0.QN.n3 0.249509
R24216 frontAnalog_v0p0p1_4.RSfetsym_0.QN.n3 frontAnalog_v0p0p1_4.RSfetsym_0.QN.n2 0.0968646
R24217 I7.n4 I7.t5 261.116
R24218 I7.n0 I7.t7 186.03
R24219 I7.n4 I7.t10 155.746
R24220 I7.n0 I7.t8 137.829
R24221 I7.n12 I7.t6 117.314
R24222 I7.n12 I7.t9 110.852
R24223 I7 I7.n0 78.5605
R24224 I7.n9 I7 47.2619
R24225 I7.n14 I7.t1 17.6181
R24226 I7.n15 I7.t0 14.2865
R24227 I7.n17 I7.t3 14.283
R24228 I7.n17 I7.t2 14.283
R24229 I7.n6 I7.n5 9.3005
R24230 I7.n19 I7.t4 8.77592
R24231 I7.n5 I7.n4 7.65549
R24232 I7.n5 I7.n2 4.64342
R24233 I7.n2 I7.n1 4.52687
R24234 I7.n6 I7.n1 4.513
R24235 I7.n9 I7.n8 4.04922
R24236 I7.n3 I7 2.46419
R24237 I7.n19 I7.n18 1.20426
R24238 I7.n10 I7 0.808983
R24239 I7.n5 I7.n3 0.754023
R24240 I7 I7.n11 0.748897
R24241 I7.n21 I7 0.713803
R24242 I7 I7.n21 0.711434
R24243 I7.n11 I7.n10 0.674526
R24244 I7.n10 I7.n9 0.478179
R24245 I7 I7.n20 0.462023
R24246 I7.n20 I7.n19 0.32511
R24247 I7.n15 I7.n14 0.314673
R24248 I7.n16 I7.n15 0.300251
R24249 I7.n11 I7 0.20675
R24250 I7.n13 I7.n12 0.159555
R24251 I7.n18 I7.n17 0.106617
R24252 I7.n16 I7.n13 0.0796167
R24253 I7.n21 I7 0.0626967
R24254 I7.n21 I7 0.06249
R24255 I7.n18 I7.n16 0.0480595
R24256 I7.n20 I7 0.046937
R24257 I7.n7 I7.n6 0.0326429
R24258 I7.n7 I7.n2 0.0197253
R24259 I7.n8 I7.n1 0.00182856
R24260 I7.n8 I7.n7 0.00149885
R24261 I7.n7 I7.n3 0.00125261
R24262 I7.n14 I7.n13 0.000504658
R24263 frontAnalog_v0p0p1_11.x63.A.n2 frontAnalog_v0p0p1_11.x63.A.t5 260.322
R24264 frontAnalog_v0p0p1_11.x63.A.n4 frontAnalog_v0p0p1_11.x63.A.t6 233.888
R24265 frontAnalog_v0p0p1_11.x63.A.n2 frontAnalog_v0p0p1_11.x63.A.t7 175.169
R24266 frontAnalog_v0p0p1_11.x63.A.n3 frontAnalog_v0p0p1_11.x63.A.t4 159.725
R24267 frontAnalog_v0p0p1_11.x63.A.n1 frontAnalog_v0p0p1_11.x63.A.t0 17.4109
R24268 frontAnalog_v0p0p1_11.x63.A.n0 frontAnalog_v0p0p1_11.x63.A.n2 9.75129
R24269 frontAnalog_v0p0p1_11.x63.A.n1 frontAnalog_v0p0p1_11.x63.A.t1 9.6027
R24270 frontAnalog_v0p0p1_11.x63.A.n0 frontAnalog_v0p0p1_11.x63.A 2.33338
R24271 frontAnalog_v0p0p1_11.x63.A.n5 frontAnalog_v0p0p1_11.x63.A.t3 8.40929
R24272 frontAnalog_v0p0p1_11.x63.A.n3 frontAnalog_v0p0p1_11.x63.A.t2 8.06629
R24273 frontAnalog_v0p0p1_11.x63.A.n4 frontAnalog_v0p0p1_11.x63.A.n3 1.73501
R24274 frontAnalog_v0p0p1_11.x63.A.n1 frontAnalog_v0p0p1_11.x63.A.n4 0.99025
R24275 frontAnalog_v0p0p1_11.x63.A.n5 frontAnalog_v0p0p1_11.x63.A.n1 0.853186
R24276 frontAnalog_v0p0p1_11.x63.A frontAnalog_v0p0p1_11.x63.A.n0 0.349517
R24277 frontAnalog_v0p0p1_11.x63.A frontAnalog_v0p0p1_11.x63.A.n5 0.24425
R24278 frontAnalog_v0p0p1_8.x65.A.n1 frontAnalog_v0p0p1_8.x65.A.t4 260.322
R24279 frontAnalog_v0p0p1_8.x65.A.n3 frontAnalog_v0p0p1_8.x65.A.t7 233.929
R24280 frontAnalog_v0p0p1_8.x65.A.n1 frontAnalog_v0p0p1_8.x65.A.t6 175.169
R24281 frontAnalog_v0p0p1_8.x65.A.n2 frontAnalog_v0p0p1_8.x65.A.t5 160.416
R24282 frontAnalog_v0p0p1_8.x65.A.n4 frontAnalog_v0p0p1_8.x65.A.t0 17.4109
R24283 frontAnalog_v0p0p1_8.x65.A.n4 frontAnalog_v0p0p1_8.x65.A.t1 10.2053
R24284 frontAnalog_v0p0p1_8.x65.A.n0 frontAnalog_v0p0p1_8.x65.A 2.78715
R24285 frontAnalog_v0p0p1_8.x65.A.n0 frontAnalog_v0p0p1_8.x65.A.n1 9.09103
R24286 frontAnalog_v0p0p1_8.x65.A.n6 frontAnalog_v0p0p1_8.x65.A.t2 7.94569
R24287 frontAnalog_v0p0p1_8.x65.A.n2 frontAnalog_v0p0p1_8.x65.A.t3 7.55846
R24288 frontAnalog_v0p0p1_8.x65.A.n5 frontAnalog_v0p0p1_8.x65.A.n3 1.4614
R24289 frontAnalog_v0p0p1_8.x65.A.n3 frontAnalog_v0p0p1_8.x65.A.n2 1.19626
R24290 frontAnalog_v0p0p1_8.x65.A.n6 frontAnalog_v0p0p1_8.x65.A.n5 0.836961
R24291 frontAnalog_v0p0p1_8.x65.A frontAnalog_v0p0p1_8.x65.A.n0 0.390342
R24292 frontAnalog_v0p0p1_8.x65.A.n5 frontAnalog_v0p0p1_8.x65.A.n4 0.154668
R24293 frontAnalog_v0p0p1_8.x65.A frontAnalog_v0p0p1_8.x65.A.n6 0.08175
R24294 I14.n17 I14.t11 260.435
R24295 I14.n2 I14.t12 229.433
R24296 I14.n12 I14.t9 196.549
R24297 I14.n2 I14.t6 158.886
R24298 I14.n17 I14.t5 156.403
R24299 I14.n12 I14.t7 148.35
R24300 I14.n27 I14.t10 117.314
R24301 I14.n27 I14.t8 110.852
R24302 I14.n13 I14.n12 76.0005
R24303 I14.n29 I14.t0 17.6181
R24304 I14.n30 I14.t3 14.2865
R24305 I14.n32 I14.t1 14.283
R24306 I14.n32 I14.t2 14.283
R24307 I14 I14.n16 9.3005
R24308 I14.n5 I14.n3 9.3005
R24309 I14.n5 I14.n4 9.3005
R24310 I14.n9 I14.n8 9.3005
R24311 I14.n34 I14.t4 8.77592
R24312 I14.n18 I14.n17 7.60183
R24313 I14.n3 I14.n2 7.39078
R24314 I14.n22 I14.n14 6.24391
R24315 I14.n13 I14 5.78114
R24316 I14.n18 I14 4.8645
R24317 I14.n19 I14.n15 4.54557
R24318 I14.n10 I14.n9 4.51698
R24319 I14.n16 I14.n15 4.51121
R24320 I14.n8 I14.n7 4.5005
R24321 I14.n22 I14.n21 3.53643
R24322 I14.n14 I14.n13 3.51018
R24323 I14.n8 I14.n4 3.46717
R24324 I14.n34 I14.n33 1.20426
R24325 I14.n6 I14.n0 1.13339
R24326 I14.n11 I14.n10 1.11384
R24327 I14.n8 I14.n3 1.06717
R24328 I14.n4 I14 1.06717
R24329 I14.n23 I14.n11 0.767464
R24330 I14.n35 I14 0.731611
R24331 I14.n24 I14 0.718556
R24332 I14 I14.n26 0.655889
R24333 I14.n26 I14 0.59035
R24334 I14.n24 I14.n23 0.503793
R24335 I14.n11 I14 0.372375
R24336 I14 I14.n34 0.370547
R24337 I14.n23 I14.n22 0.321929
R24338 I14.n30 I14.n29 0.314673
R24339 I14.n31 I14.n30 0.300251
R24340 I14 I14.n35 0.299591
R24341 I14.n14 I14 0.206952
R24342 I14.n25 I14 0.2005
R24343 I14.n28 I14.n27 0.159555
R24344 I14.n33 I14.n32 0.106617
R24345 I14.n31 I14.n28 0.0796167
R24346 I14.n33 I14.n31 0.0480595
R24347 I14.n20 I14.n16 0.0344286
R24348 I14.n25 I14.n24 0.0287
R24349 I14.n26 I14.n25 0.0287
R24350 I14.n10 I14.n0 0.028
R24351 I14.n35 I14 0.0266111
R24352 I14.n9 I14.n1 0.0142363
R24353 I14.n35 I14 0.0111818
R24354 I14.n7 I14.n1 0.00599451
R24355 I14.n6 I14.n5 0.00409723
R24356 I14.n7 I14.n6 0.00202085
R24357 I14.n21 I14.n15 0.00182856
R24358 I14.n21 I14.n20 0.00149885
R24359 I14.n19 I14.n18 0.00133362
R24360 I14.n20 I14.n19 0.00100077
R24361 I14.n1 I14.n0 0.000617139
R24362 I14.n29 I14.n28 0.000504658
R24363 I15.n4 I15.t5 261.116
R24364 I15.n0 I15.t7 186.03
R24365 I15.n4 I15.t9 155.746
R24366 I15.n0 I15.t6 137.829
R24367 I15.n14 I15.t10 117.314
R24368 I15.n14 I15.t8 110.852
R24369 I15 I15.n0 78.5605
R24370 I15.n9 I15 47.2619
R24371 I15.n16 I15.t0 17.6181
R24372 I15.n17 I15.t4 14.2865
R24373 I15.n19 I15.t2 14.283
R24374 I15.n19 I15.t1 14.283
R24375 I15.n6 I15.n5 9.3005
R24376 I15.n21 I15.t3 8.77592
R24377 I15.n5 I15.n4 7.65549
R24378 I15.n5 I15.n2 4.64342
R24379 I15.n2 I15.n1 4.52687
R24380 I15.n6 I15.n1 4.513
R24381 I15.n9 I15.n8 4.04922
R24382 I15.n3 I15 2.46419
R24383 I15.n21 I15.n20 1.20426
R24384 I15.n5 I15.n3 0.754023
R24385 I15.n10 I15 0.70184
R24386 I15.n11 I15.n10 0.662978
R24387 I15.n10 I15.n9 0.585321
R24388 I15.n11 I15 0.577556
R24389 I15.n22 I15 0.559278
R24390 I15 I15.n13 0.514889
R24391 I15.n13 I15 0.46345
R24392 I15 I15.n21 0.370547
R24393 I15.n17 I15.n16 0.314673
R24394 I15.n18 I15.n17 0.300251
R24395 I15 I15.n22 0.25195
R24396 I15.n12 I15 0.2005
R24397 I15.n15 I15.n14 0.159555
R24398 I15.n20 I15.n19 0.106617
R24399 I15.n18 I15.n15 0.0796167
R24400 I15.n20 I15.n18 0.0480595
R24401 I15.n7 I15.n6 0.0326429
R24402 I15.n12 I15.n11 0.0287
R24403 I15.n13 I15.n12 0.0287
R24404 I15.n22 I15 0.0266111
R24405 I15.n7 I15.n2 0.0197253
R24406 I15.n22 I15 0.01225
R24407 I15.n8 I15.n1 0.00182856
R24408 I15.n8 I15.n7 0.00149885
R24409 I15.n7 I15.n3 0.00125261
R24410 I15.n16 I15.n15 0.000504658
R24411 I3.n4 I3.t7 334.723
R24412 I3.n3 I3.t10 323.342
R24413 I3.n4 I3.t9 206.19
R24414 I3.n3 I3.t6 194.809
R24415 I3.n0 I3.t5 186.03
R24416 I3.n0 I3.t11 137.829
R24417 I3.n8 I3.t12 117.314
R24418 I3.n8 I3.t8 110.853
R24419 I3 I3.n4 84.2291
R24420 I3 I3.n3 82.1338
R24421 I3.n1 I3.n0 76.0005
R24422 I3.n2 I3 66.7187
R24423 I3.n5 I3 26.4877
R24424 I3.n10 I3.t0 17.6181
R24425 I3.n11 I3.t3 14.2865
R24426 I3.n13 I3.t1 14.283
R24427 I3.n13 I3.t2 14.283
R24428 I3.n15 I3.t4 8.77744
R24429 I3.n1 I3 7.31479
R24430 I3 I3.n16 5.79898
R24431 I3.n5 I3 4.36044
R24432 I3 I3.n1 4.02336
R24433 I3.n6 I3.n5 2.61211
R24434 I3.n6 I3.n2 1.25943
R24435 I3.n15 I3.n14 1.20426
R24436 I3.n2 I3 0.969697
R24437 I3.n17 I3 0.431333
R24438 I3 I3.n7 0.420367
R24439 I3.n16 I3.n15 0.32511
R24440 I3 I3.n17 0.323625
R24441 I3.n11 I3.n10 0.314673
R24442 I3.n7 I3.n6 0.300322
R24443 I3.n12 I3.n11 0.299251
R24444 I3.n7 I3 0.20675
R24445 I3.n9 I3.n8 0.159555
R24446 I3.n14 I3.n13 0.106617
R24447 I3.n12 I3.n9 0.0796167
R24448 I3.n14 I3.n12 0.0480595
R24449 I3.n16 I3 0.046937
R24450 I3.n17 I3 0.0161667
R24451 I3.n17 I3 0.01225
R24452 I3.n10 I3.n9 0.000504658
R24453 frontAnalog_v0p0p1_1.RSfetsym_0.QN.n1 frontAnalog_v0p0p1_1.RSfetsym_0.QN.t6 117.511
R24454 frontAnalog_v0p0p1_1.RSfetsym_0.QN.n1 frontAnalog_v0p0p1_1.RSfetsym_0.QN.t5 110.698
R24455 frontAnalog_v0p0p1_1.RSfetsym_0.QN.n2 frontAnalog_v0p0p1_1.RSfetsym_0.QN.t2 19.1963
R24456 frontAnalog_v0p0p1_1.RSfetsym_0.QN.n3 frontAnalog_v0p0p1_1.RSfetsym_0.QN.t0 14.5206
R24457 frontAnalog_v0p0p1_1.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_1.RSfetsym_0.QN.t4 14.283
R24458 frontAnalog_v0p0p1_1.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_1.RSfetsym_0.QN.t3 14.283
R24459 frontAnalog_v0p0p1_1.RSfetsym_0.QN frontAnalog_v0p0p1_1.RSfetsym_0.QN.t1 9.14075
R24460 frontAnalog_v0p0p1_1.RSfetsym_0.QN.n2 frontAnalog_v0p0p1_1.RSfetsym_0.QN.n1 0.826818
R24461 frontAnalog_v0p0p1_1.RSfetsym_0.QN frontAnalog_v0p0p1_1.RSfetsym_0.QN.n0 0.74645
R24462 frontAnalog_v0p0p1_1.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_1.RSfetsym_0.QN.n3 0.249509
R24463 frontAnalog_v0p0p1_1.RSfetsym_0.QN.n3 frontAnalog_v0p0p1_1.RSfetsym_0.QN.n2 0.0968646
R24464 I11.n4 I11.t7 334.723
R24465 I11.n3 I11.t9 323.342
R24466 I11.n4 I11.t11 206.19
R24467 I11.n3 I11.t6 194.809
R24468 I11.n0 I11.t5 186.03
R24469 I11.n0 I11.t10 137.829
R24470 I11.n10 I11.t12 117.314
R24471 I11.n10 I11.t8 110.852
R24472 I11 I11.n4 84.2291
R24473 I11 I11.n3 82.1338
R24474 I11.n1 I11.n0 76.0005
R24475 I11.n2 I11 66.7187
R24476 I11.n5 I11 26.4877
R24477 I11.n12 I11.t1 17.6181
R24478 I11.n13 I11.t0 14.2865
R24479 I11.n15 I11.t2 14.283
R24480 I11.n15 I11.t3 14.283
R24481 I11.n17 I11.t4 8.77592
R24482 I11.n1 I11 7.31479
R24483 I11.n5 I11 4.36044
R24484 I11 I11.n1 4.02336
R24485 I11 I11.n18 3.30508
R24486 I11.n6 I11.n5 2.71925
R24487 I11.n17 I11.n16 1.20426
R24488 I11.n19 I11 1.17028
R24489 I11.n6 I11.n2 1.15229
R24490 I11.n7 I11 1.14156
R24491 I11 I11.n9 1.07889
R24492 I11.n9 I11 0.97105
R24493 I11.n2 I11 0.969697
R24494 I11 I11.n19 0.957591
R24495 I11.n18 I11.n17 0.33431
R24496 I11.n13 I11.n12 0.314673
R24497 I11.n14 I11.n13 0.300251
R24498 I11.n7 I11.n6 0.28348
R24499 I11.n8 I11 0.2005
R24500 I11.n11 I11.n10 0.159555
R24501 I11.n16 I11.n15 0.106617
R24502 I11.n14 I11.n11 0.0796167
R24503 I11.n16 I11.n14 0.0480595
R24504 I11.n8 I11.n7 0.0287
R24505 I11.n9 I11.n8 0.0287
R24506 I11.n19 I11 0.0109444
R24507 I11.n19 I11 0.00904545
R24508 I11.n18 I11 0.0087668
R24509 I11.n12 I11.n11 0.000504658
R24510 frontAnalog_v0p0p1_8.x63.A.n2 frontAnalog_v0p0p1_8.x63.A.t5 260.322
R24511 frontAnalog_v0p0p1_8.x63.A.n4 frontAnalog_v0p0p1_8.x63.A.t6 233.888
R24512 frontAnalog_v0p0p1_8.x63.A.n2 frontAnalog_v0p0p1_8.x63.A.t7 175.169
R24513 frontAnalog_v0p0p1_8.x63.A.n3 frontAnalog_v0p0p1_8.x63.A.t4 159.725
R24514 frontAnalog_v0p0p1_8.x63.A.n1 frontAnalog_v0p0p1_8.x63.A.t1 17.4109
R24515 frontAnalog_v0p0p1_8.x63.A.n0 frontAnalog_v0p0p1_8.x63.A.n2 9.75129
R24516 frontAnalog_v0p0p1_8.x63.A.n1 frontAnalog_v0p0p1_8.x63.A.t0 9.6027
R24517 frontAnalog_v0p0p1_8.x63.A.n0 frontAnalog_v0p0p1_8.x63.A 2.33338
R24518 frontAnalog_v0p0p1_8.x63.A.n5 frontAnalog_v0p0p1_8.x63.A.t2 8.40929
R24519 frontAnalog_v0p0p1_8.x63.A.n3 frontAnalog_v0p0p1_8.x63.A.t3 8.06629
R24520 frontAnalog_v0p0p1_8.x63.A.n4 frontAnalog_v0p0p1_8.x63.A.n3 1.73501
R24521 frontAnalog_v0p0p1_8.x63.A.n1 frontAnalog_v0p0p1_8.x63.A.n4 0.99025
R24522 frontAnalog_v0p0p1_8.x63.A.n5 frontAnalog_v0p0p1_8.x63.A.n1 0.853186
R24523 frontAnalog_v0p0p1_8.x63.A frontAnalog_v0p0p1_8.x63.A.n0 0.349517
R24524 frontAnalog_v0p0p1_8.x63.A frontAnalog_v0p0p1_8.x63.A.n5 0.24425
R24525 frontAnalog_v0p0p1_2.RSfetsym_0.QN.n1 frontAnalog_v0p0p1_2.RSfetsym_0.QN.t5 117.511
R24526 frontAnalog_v0p0p1_2.RSfetsym_0.QN.n1 frontAnalog_v0p0p1_2.RSfetsym_0.QN.t6 110.698
R24527 frontAnalog_v0p0p1_2.RSfetsym_0.QN.n2 frontAnalog_v0p0p1_2.RSfetsym_0.QN.t2 19.1963
R24528 frontAnalog_v0p0p1_2.RSfetsym_0.QN.n3 frontAnalog_v0p0p1_2.RSfetsym_0.QN.t0 14.5206
R24529 frontAnalog_v0p0p1_2.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_2.RSfetsym_0.QN.t3 14.283
R24530 frontAnalog_v0p0p1_2.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_2.RSfetsym_0.QN.t4 14.283
R24531 frontAnalog_v0p0p1_2.RSfetsym_0.QN frontAnalog_v0p0p1_2.RSfetsym_0.QN.t1 9.14075
R24532 frontAnalog_v0p0p1_2.RSfetsym_0.QN.n2 frontAnalog_v0p0p1_2.RSfetsym_0.QN.n1 0.826818
R24533 frontAnalog_v0p0p1_2.RSfetsym_0.QN frontAnalog_v0p0p1_2.RSfetsym_0.QN.n0 0.74645
R24534 frontAnalog_v0p0p1_2.RSfetsym_0.QN.n0 frontAnalog_v0p0p1_2.RSfetsym_0.QN.n3 0.249509
R24535 frontAnalog_v0p0p1_2.RSfetsym_0.QN.n3 frontAnalog_v0p0p1_2.RSfetsym_0.QN.n2 0.0968646
R24536 frontAnalog_v0p0p1_12.x65.A.n1 frontAnalog_v0p0p1_12.x65.A.t4 260.322
R24537 frontAnalog_v0p0p1_12.x65.A.n3 frontAnalog_v0p0p1_12.x65.A.t7 233.929
R24538 frontAnalog_v0p0p1_12.x65.A.n1 frontAnalog_v0p0p1_12.x65.A.t6 175.169
R24539 frontAnalog_v0p0p1_12.x65.A.n2 frontAnalog_v0p0p1_12.x65.A.t5 160.416
R24540 frontAnalog_v0p0p1_12.x65.A.n4 frontAnalog_v0p0p1_12.x65.A.t1 17.4109
R24541 frontAnalog_v0p0p1_12.x65.A.n4 frontAnalog_v0p0p1_12.x65.A.t0 10.2053
R24542 frontAnalog_v0p0p1_12.x65.A.n0 frontAnalog_v0p0p1_12.x65.A 2.78715
R24543 frontAnalog_v0p0p1_12.x65.A.n0 frontAnalog_v0p0p1_12.x65.A.n1 9.09103
R24544 frontAnalog_v0p0p1_12.x65.A.n6 frontAnalog_v0p0p1_12.x65.A.t3 7.94569
R24545 frontAnalog_v0p0p1_12.x65.A.n2 frontAnalog_v0p0p1_12.x65.A.t2 7.55846
R24546 frontAnalog_v0p0p1_12.x65.A.n5 frontAnalog_v0p0p1_12.x65.A.n3 1.4614
R24547 frontAnalog_v0p0p1_12.x65.A.n3 frontAnalog_v0p0p1_12.x65.A.n2 1.19626
R24548 frontAnalog_v0p0p1_12.x65.A.n6 frontAnalog_v0p0p1_12.x65.A.n5 0.836961
R24549 frontAnalog_v0p0p1_12.x65.A frontAnalog_v0p0p1_12.x65.A.n0 0.390342
R24550 frontAnalog_v0p0p1_12.x65.A.n5 frontAnalog_v0p0p1_12.x65.A.n4 0.154668
R24551 frontAnalog_v0p0p1_12.x65.A frontAnalog_v0p0p1_12.x65.A.n6 0.08175
R24552 frontAnalog_v0p0p1_6.x65.A.n1 frontAnalog_v0p0p1_6.x65.A.t6 260.322
R24553 frontAnalog_v0p0p1_6.x65.A.n3 frontAnalog_v0p0p1_6.x65.A.t5 233.929
R24554 frontAnalog_v0p0p1_6.x65.A.n1 frontAnalog_v0p0p1_6.x65.A.t7 175.169
R24555 frontAnalog_v0p0p1_6.x65.A.n2 frontAnalog_v0p0p1_6.x65.A.t4 160.416
R24556 frontAnalog_v0p0p1_6.x65.A.n4 frontAnalog_v0p0p1_6.x65.A.t0 17.4109
R24557 frontAnalog_v0p0p1_6.x65.A.n4 frontAnalog_v0p0p1_6.x65.A.t1 10.2053
R24558 frontAnalog_v0p0p1_6.x65.A.n0 frontAnalog_v0p0p1_6.x65.A 2.78715
R24559 frontAnalog_v0p0p1_6.x65.A.n0 frontAnalog_v0p0p1_6.x65.A.n1 9.09103
R24560 frontAnalog_v0p0p1_6.x65.A.n6 frontAnalog_v0p0p1_6.x65.A.t2 7.94569
R24561 frontAnalog_v0p0p1_6.x65.A.n2 frontAnalog_v0p0p1_6.x65.A.t3 7.55846
R24562 frontAnalog_v0p0p1_6.x65.A.n5 frontAnalog_v0p0p1_6.x65.A.n3 1.4614
R24563 frontAnalog_v0p0p1_6.x65.A.n3 frontAnalog_v0p0p1_6.x65.A.n2 1.19626
R24564 frontAnalog_v0p0p1_6.x65.A.n6 frontAnalog_v0p0p1_6.x65.A.n5 0.836961
R24565 frontAnalog_v0p0p1_6.x65.A frontAnalog_v0p0p1_6.x65.A.n0 0.390342
R24566 frontAnalog_v0p0p1_6.x65.A.n5 frontAnalog_v0p0p1_6.x65.A.n4 0.154668
R24567 frontAnalog_v0p0p1_6.x65.A frontAnalog_v0p0p1_6.x65.A.n6 0.08175
R24568 frontAnalog_v0p0p1_0.x65.A.n1 frontAnalog_v0p0p1_0.x65.A.t5 260.322
R24569 frontAnalog_v0p0p1_0.x65.A.n3 frontAnalog_v0p0p1_0.x65.A.t7 233.929
R24570 frontAnalog_v0p0p1_0.x65.A.n1 frontAnalog_v0p0p1_0.x65.A.t6 175.169
R24571 frontAnalog_v0p0p1_0.x65.A.n2 frontAnalog_v0p0p1_0.x65.A.t4 160.416
R24572 frontAnalog_v0p0p1_0.x65.A.n4 frontAnalog_v0p0p1_0.x65.A.t0 17.4109
R24573 frontAnalog_v0p0p1_0.x65.A.n4 frontAnalog_v0p0p1_0.x65.A.t3 10.2053
R24574 frontAnalog_v0p0p1_0.x65.A.n0 frontAnalog_v0p0p1_0.x65.A 2.78715
R24575 frontAnalog_v0p0p1_0.x65.A.n0 frontAnalog_v0p0p1_0.x65.A.n1 9.09103
R24576 frontAnalog_v0p0p1_0.x65.A.n6 frontAnalog_v0p0p1_0.x65.A.t1 7.94569
R24577 frontAnalog_v0p0p1_0.x65.A.n2 frontAnalog_v0p0p1_0.x65.A.t2 7.55846
R24578 frontAnalog_v0p0p1_0.x65.A.n5 frontAnalog_v0p0p1_0.x65.A.n3 1.4614
R24579 frontAnalog_v0p0p1_0.x65.A.n3 frontAnalog_v0p0p1_0.x65.A.n2 1.19626
R24580 frontAnalog_v0p0p1_0.x65.A.n6 frontAnalog_v0p0p1_0.x65.A.n5 0.836961
R24581 frontAnalog_v0p0p1_0.x65.A frontAnalog_v0p0p1_0.x65.A.n0 0.390342
R24582 frontAnalog_v0p0p1_0.x65.A.n5 frontAnalog_v0p0p1_0.x65.A.n4 0.154668
R24583 frontAnalog_v0p0p1_0.x65.A frontAnalog_v0p0p1_0.x65.A.n6 0.08175
R24584 frontAnalog_v0p0p1_0.x63.A.n2 frontAnalog_v0p0p1_0.x63.A.t5 260.322
R24585 frontAnalog_v0p0p1_0.x63.A.n4 frontAnalog_v0p0p1_0.x63.A.t4 233.888
R24586 frontAnalog_v0p0p1_0.x63.A.n2 frontAnalog_v0p0p1_0.x63.A.t6 175.169
R24587 frontAnalog_v0p0p1_0.x63.A.n3 frontAnalog_v0p0p1_0.x63.A.t7 159.725
R24588 frontAnalog_v0p0p1_0.x63.A.n1 frontAnalog_v0p0p1_0.x63.A.t0 17.4109
R24589 frontAnalog_v0p0p1_0.x63.A.n0 frontAnalog_v0p0p1_0.x63.A.n2 9.75129
R24590 frontAnalog_v0p0p1_0.x63.A.n1 frontAnalog_v0p0p1_0.x63.A.t1 9.6027
R24591 frontAnalog_v0p0p1_0.x63.A.n0 frontAnalog_v0p0p1_0.x63.A 2.33338
R24592 frontAnalog_v0p0p1_0.x63.A.n5 frontAnalog_v0p0p1_0.x63.A.t2 8.40929
R24593 frontAnalog_v0p0p1_0.x63.A.n3 frontAnalog_v0p0p1_0.x63.A.t3 8.06629
R24594 frontAnalog_v0p0p1_0.x63.A.n4 frontAnalog_v0p0p1_0.x63.A.n3 1.73501
R24595 frontAnalog_v0p0p1_0.x63.A.n1 frontAnalog_v0p0p1_0.x63.A.n4 0.99025
R24596 frontAnalog_v0p0p1_0.x63.A.n5 frontAnalog_v0p0p1_0.x63.A.n1 0.853186
R24597 frontAnalog_v0p0p1_0.x63.A frontAnalog_v0p0p1_0.x63.A.n0 0.349517
R24598 frontAnalog_v0p0p1_0.x63.A frontAnalog_v0p0p1_0.x63.A.n5 0.24425
C0 frontAnalog_v0p0p1_13.RSfetsym_0.QN I4 0.0512f
C1 a_57123_n9479# VDD 0.222f
C2 16to4_PriorityEncoder_v0p0p1_0.x3.x14.A 16to4_PriorityEncoder_v0p0p1_0.x3.x11.X 0.0721f
C3 frontAnalog_v0p0p1_14.RSfetsym_0.QN VDD 2.56f
C4 frontAnalog_v0p0p1_0.x63.X I14 1.78f
C5 a_77639_n42341# VDD 0.318f
C6 w_55000_n83928# w_55000_n84550# 0.327f
C7 w_55000_n68350# a_55268_n68736# 0.12f
C8 I9 I8 3.07f
C9 frontAnalog_v0p0p1_0.RSfetsym_0.QN frontAnalog_v0p0p1_0.RSfetsym_0.x1.Y 0.17f
C10 16to4_PriorityEncoder_v0p0p1_0.x5.x19.C I13 0.407f
C11 a_57123_n61959# frontAnalog_v0p0p1_11.x65.X 0.119f
C12 a_59578_n19170# I12 0.42f
C13 a_77605_n52819# I3 0.15f
C14 VV1 VL 1.96f
C15 a_53630_n14796# a_55268_n14736# 0.015f
C16 frontAnalog_v0p0p1_2.x65.A frontAnalog_v0p0p1_2.x65.X 0.0236f
C17 a_59577_n79083# VDD 0.0173f
C18 frontAnalog_v0p0p1_0.RSfetsym_0.QN VDD 2.56f
C19 w_55000_n35950# VIN 0.737f
C20 frontAnalog_v0p0p1_11.x65.A VIN 0.655f
C21 a_77605_n48109# I6 0.214f
C22 16to4_PriorityEncoder_v0p0p1_0.x3.A1 16to4_PriorityEncoder_v0p0p1_0.x3.x17.A 0.115f
C23 16to4_PriorityEncoder_v0p0p1_0.x5.x18.C I9 0.495f
C24 w_55000_n8328# frontAnalog_v0p0p1_0.x63.A 0.0792f
C25 w_55000_n30550# frontAnalog_v0p0p1_6.x65.A 0.0988f
C26 frontAnalog_v0p0p1_3.x65.A VIN 0.655f
C27 a_55268_n84936# VIN 0.177f
C28 frontAnalog_v0p0p1_5.x63.X I11 1.93f
C29 frontAnalog_v0p0p1_13.RSfetsym_0.x1.Y VDD 0.733f
C30 a_55268_n52536# VV7 0.215f
C31 w_55000_n2928# frontAnalog_v0p0p1_2.x65.A 0.658f
C32 16to4_PriorityEncoder_v0p0p1_0.x5.x17.A 16to4_PriorityEncoder_v0p0p1_0.x5.x15.X 0.0789f
C33 a_53630_n68796# CLK 0.0136f
C34 frontAnalog_v0p0p1_9.x63.X I6 1.85f
C35 a_53630_n84996# VV1 0.28f
C36 w_55000_n51528# frontAnalog_v0p0p1_9.x65.A 0.658f
C37 m3_58396_n4350# I15 0.0416f
C38 16to4_PriorityEncoder_v0p0p1_0.x5.x19.X 16to4_PriorityEncoder_v0p0p1_0.x5.x20.X 0.145f
C39 frontAnalog_v0p0p1_5.x63.A frontAnalog_v0p0p1_5.x63.X 0.0301f
C40 frontAnalog_v0p0p1_0.RSfetsym_0.x1.Y frontAnalog_v0p0p1_0.RSfetsym_0.x2.Y 0.0254f
C41 frontAnalog_v0p0p1_14.RSfetsym_0.QN a_59577_n79083# 0.418f
C42 16to4_PriorityEncoder_v0p0p1_0.x3.x16.C I1 0.0914f
C43 frontAnalog_v0p0p1_11.x65.X a_59578_n62370# 0.436f
C44 16to4_PriorityEncoder_v0p0p1_0.x5.x21.B 16to4_PriorityEncoder_v0p0p1_0.x5.x19.X 0.262f
C45 16to4_PriorityEncoder_v0p0p1_0.x3.x19.D 16to4_PriorityEncoder_v0p0p1_0.x3.x19.X 0.0195f
C46 w_55000_n3550# frontAnalog_v0p0p1_2.x63.A 0.659f
C47 w_55000_n46128# w_55000_n46750# 0.327f
C48 w_55000_n67728# VDD 0.854f
C49 frontAnalog_v0p0p1_12.x65.X frontAnalog_v0p0p1_12.RSfetsym_0.x1.Y 0.182f
C50 frontAnalog_v0p0p1_10.x65.X VDD 3.55f
C51 16to4_PriorityEncoder_v0p0p1_0.x3.x22.A I7 0.0853f
C52 frontAnalog_v0p0p1_0.RSfetsym_0.x2.Y VDD 0.926f
C53 w_55000_n52150# frontAnalog_v0p0p1_9.x63.A 0.659f
C54 frontAnalog_v0p0p1_10.IB a_53630_n63396# 0.473f
C55 a_57123_n68879# VDD 0.222f
C56 frontAnalog_v0p0p1_4.x63.A a_57123_n20279# 0.212f
C57 16to4_PriorityEncoder_v0p0p1_0.x3.x16.C I7 0.26f
C58 a_77605_n39305# 16to4_PriorityEncoder_v0p0p1_0.x5.x1.X 0.0991f
C59 I13 I8 0.331f
C60 frontAnalog_v0p0p1_4.RSfetsym_0.x1.Y I12 0.0436f
C61 a_53630_n74196# VIN 0.265f
C62 16to4_PriorityEncoder_v0p0p1_0.x5.x22.A 16to4_PriorityEncoder_v0p0p1_0.x5.x16.X 0.0732f
C63 16to4_PriorityEncoder_v0p0p1_0.x3.A1 16to4_PriorityEncoder_v0p0p1_0.x3.x15.X 0.0206f
C64 VIN VV8 2.62f
C65 m3_58396_n47550# VDD 1.3f
C66 frontAnalog_v0p0p1_7.x65.A VDD 3.45f
C67 w_55000_n57550# frontAnalog_v0p0p1_10.x65.A 0.0988f
C68 frontAnalog_v0p0p1_13.RSfetsym_0.QN a_59578_n67770# 0.255f
C69 frontAnalog_v0p0p1_4.x63.A CLK 1.81f
C70 16to4_PriorityEncoder_v0p0p1_0.x5.x22.A 16to4_PriorityEncoder_v0p0p1_0.x5.x21.B 0.064f
C71 frontAnalog_v0p0p1_1.x65.X CLK 0.0393f
C72 w_55000_n19750# CLK 0.535f
C73 frontAnalog_v0p0p1_8.x65.X VDD 3.55f
C74 w_55000_n40728# frontAnalog_v0p0p1_10.IB 0.0216f
C75 16to4_PriorityEncoder_v0p0p1_0.x3.EI 16to4_PriorityEncoder_v0p0p1_0.x3.x21.B 0.187f
C76 frontAnalog_v0p0p1_13.RSfetsym_0.QN VDD 2.56f
C77 16to4_PriorityEncoder_v0p0p1_0.x5.x18.C I13 0.3f
C78 frontAnalog_v0p0p1_12.RSfetsym_0.x1.Y frontAnalog_v0p0p1_12.x63.X 0.883f
C79 frontAnalog_v0p0p1_10.x63.X VDD 3.16f
C80 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_9.x63.A 0.0926f
C81 w_55000_n78528# frontAnalog_v0p0p1_14.x65.A 0.658f
C82 w_55000_n78528# VIN 0.866f
C83 w_55000_n8328# w_55000_n8950# 0.327f
C84 a_78159_n47589# 16to4_PriorityEncoder_v0p0p1_0.x3.x2.X 0.121f
C85 a_59577_n8883# I14 0.29f
C86 16to4_PriorityEncoder_v0p0p1_0.x5.x2.X a_77605_n40069# 0.134f
C87 frontAnalog_v0p0p1_10.x63.A a_55268_n57936# 1.24f
C88 frontAnalog_v0p0p1_0.RSfetsym_0.QN frontAnalog_v0p0p1_0.RSfetsym_0.x2.Y 0.018f
C89 frontAnalog_v0p0p1_11.x65.X frontAnalog_v0p0p1_11.RSfetsym_0.x1.Y 0.182f
C90 frontAnalog_v0p0p1_4.x65.A frontAnalog_v0p0p1_4.x65.X 0.0236f
C91 a_53630_n30996# a_55268_n30936# 0.015f
C92 a_55268_n79536# CLK 0.236f
C93 frontAnalog_v0p0p1_12.x65.X frontAnalog_v0p0p1_12.RSfetsym_0.QN 2.28f
C94 frontAnalog_v0p0p1_5.x63.A VIN 0.188f
C95 w_55000_n79150# frontAnalog_v0p0p1_14.x63.A 0.659f
C96 frontAnalog_v0p0p1_1.x65.A frontAnalog_v0p0p1_1.x65.X 0.0236f
C97 frontAnalog_v0p0p1_6.RSfetsym_0.QN I11 0.0512f
C98 frontAnalog_v0p0p1_13.x65.X frontAnalog_v0p0p1_13.x63.X 0.136f
C99 frontAnalog_v0p0p1_0.x63.X a_59577_n8883# 0.28f
C100 a_59577_n25083# I11 0.29f
C101 VV10 VV9 2.78f
C102 frontAnalog_v0p0p1_1.RSfetsym_0.x1.Y I8 0.0439f
C103 CLK I12 0.01f
C104 frontAnalog_v0p0p1_8.x63.X a_57123_n47279# 0.121f
C105 frontAnalog_v0p0p1_13.RSfetsym_0.x2.Y VDD 0.926f
C106 frontAnalog_v0p0p1_0.x63.A frontAnalog_v0p0p1_0.x65.A 3.16f
C107 frontAnalog_v0p0p1_4.RSfetsym_0.QN I12 2.02f
C108 frontAnalog_v0p0p1_12.x63.X a_57123_n74279# 0.121f
C109 a_57123_n18759# VDD 0.224f
C110 frontAnalog_v0p0p1_6.x65.A CLK 2.62f
C111 frontAnalog_v0p0p1_10.RSfetsym_0.QN a_59578_n56970# 0.255f
C112 frontAnalog_v0p0p1_10.IB a_55268_n74136# 0.0848f
C113 16to4_PriorityEncoder_v0p0p1_0.x3.x22.A 16to4_PriorityEncoder_v0p0p1_0.x3.x19.X 0.418f
C114 frontAnalog_v0p0p1_13.RSfetsym_0.QN frontAnalog_v0p0p1_13.RSfetsym_0.x1.Y 0.17f
C115 16to4_PriorityEncoder_v0p0p1_0.x3.A1 16to4_PriorityEncoder_v0p0p1_0.x3.x22.A 0.519f
C116 w_55000_n2928# VIN 0.867f
C117 frontAnalog_v0p0p1_11.RSfetsym_0.x1.Y frontAnalog_v0p0p1_11.x63.X 0.883f
C118 frontAnalog_v0p0p1_8.RSfetsym_0.x2.Y I7 0.198f
C119 frontAnalog_v0p0p1_12.x65.X frontAnalog_v0p0p1_12.RSfetsym_0.x2.Y 0.526f
C120 frontAnalog_v0p0p1_12.RSfetsym_0.QN frontAnalog_v0p0p1_12.x63.X 0.378f
C121 m3_58396_n25950# I11 0.0416f
C122 16to4_PriorityEncoder_v0p0p1_0.x5.x22.A 16to4_PriorityEncoder_v0p0p1_0.x5.x15.X 0.209f
C123 w_55000_n13728# a_53630_n14796# 0.359f
C124 16to4_PriorityEncoder_v0p0p1_0.x5.x19.X 16to4_PriorityEncoder_v0p0p1_0.x5.x21.X 0.131f
C125 w_55000_n62328# CLK 0.571f
C126 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_5.x65.A 0.0352f
C127 w_55000_n79150# frontAnalog_v0p0p1_10.IB 0.0217f
C128 a_55268_n57936# CLK 0.236f
C129 frontAnalog_v0p0p1_11.x65.X frontAnalog_v0p0p1_11.RSfetsym_0.QN 2.28f
C130 CLK I0 0.0103f
C131 frontAnalog_v0p0p1_4.RSfetsym_0.x2.Y I12 0.196f
C132 16to4_PriorityEncoder_v0p0p1_0.x5.A2 16to4_PriorityEncoder_v0p0p1_0.x1.A 0.38f
C133 a_59578_n19170# VDD 0.0213f
C134 w_55000_n41350# a_55268_n41736# 0.12f
C135 w_55000_n30550# VDD 0.829f
C136 frontAnalog_v0p0p1_10.x65.X frontAnalog_v0p0p1_10.x63.X 0.136f
C137 frontAnalog_v0p0p1_3.x65.X I13 0.446f
C138 a_78159_n47589# 16to4_PriorityEncoder_v0p0p1_0.x3.x1.X 0.192f
C139 frontAnalog_v0p0p1_13.RSfetsym_0.x1.Y frontAnalog_v0p0p1_13.RSfetsym_0.x2.Y 0.0254f
C140 frontAnalog_v0p0p1_1.x63.X I8 1.86f
C141 a_59578_n56970# I5 0.42f
C142 a_78097_n45737# VDD 0.332f
C143 frontAnalog_v0p0p1_11.x63.X a_57123_n63479# 0.121f
C144 16to4_PriorityEncoder_v0p0p1_0.x3.x19.C I1 0.347f
C145 frontAnalog_v0p0p1_8.x63.X frontAnalog_v0p0p1_8.RSfetsym_0.x2.Y 0.0923f
C146 16to4_PriorityEncoder_v0p0p1_0.x3.x21.B VDD 0.721f
C147 VDD VV10 4.56f
C148 frontAnalog_v0p0p1_12.x63.X frontAnalog_v0p0p1_12.RSfetsym_0.x2.Y 0.0923f
C149 frontAnalog_v0p0p1_9.x63.A VV7 0.587f
C150 CLK I4 0.01f
C151 frontAnalog_v0p0p1_9.RSfetsym_0.QN frontAnalog_v0p0p1_9.x63.X 0.378f
C152 16to4_PriorityEncoder_v0p0p1_0.x5.x22.A 16to4_PriorityEncoder_v0p0p1_0.x5.x21.X 0.0749f
C153 a_59577_n57483# VDD 0.0173f
C154 frontAnalog_v0p0p1_10.RSfetsym_0.QN frontAnalog_v0p0p1_10.RSfetsym_0.x1.Y 0.17f
C155 a_55268_n47136# CLK 0.236f
C156 I0 R0 1.89f
C157 frontAnalog_v0p0p1_15.x65.A VDD 3.45f
C158 a_55268_n63336# VIN 0.177f
C159 a_77605_n43295# VDD 0.551f
C160 w_55000_n8950# frontAnalog_v0p0p1_0.x65.A 0.0988f
C161 m3_58396_n74550# I2 0.0416f
C162 frontAnalog_v0p0p1_11.x65.X frontAnalog_v0p0p1_11.RSfetsym_0.x2.Y 0.526f
C163 frontAnalog_v0p0p1_11.RSfetsym_0.QN frontAnalog_v0p0p1_11.x63.X 0.378f
C164 frontAnalog_v0p0p1_9.x65.A VIN 0.655f
C165 w_55000_n3550# frontAnalog_v0p0p1_10.IB 0.0217f
C166 16to4_PriorityEncoder_v0p0p1_0.x3.x19.C I7 0.239f
C167 frontAnalog_v0p0p1_3.x63.X I13 1.85f
C168 a_78159_n47589# 16to4_PriorityEncoder_v0p0p1_0.x3.EO 0.128f
C169 CLK VV9 6.38f
C170 a_53630_n52596# VDD 0.134f
C171 frontAnalog_v0p0p1_10.x63.A VDD 3.67f
C172 w_55000_n41350# VIN 0.737f
C173 frontAnalog_v0p0p1_4.RSfetsym_0.x1.Y VDD 0.733f
C174 w_55000_n73128# VV3 0.798f
C175 frontAnalog_v0p0p1_10.RSfetsym_0.x1.Y frontAnalog_v0p0p1_10.RSfetsym_0.x2.Y 0.0254f
C176 16to4_PriorityEncoder_v0p0p1_0.x3.A2 VDD 1.79f
C177 frontAnalog_v0p0p1_13.RSfetsym_0.QN frontAnalog_v0p0p1_13.RSfetsym_0.x2.Y 0.018f
C178 16to4_PriorityEncoder_v0p0p1_0.x1.A a_82906_n47995# 0.206f
C179 16to4_PriorityEncoder_v0p0p1_0.x2.A 16to4_PriorityEncoder_v0p0p1_0.x3.GS 0.0652f
C180 a_53630_n20196# CLK 0.0136f
C181 frontAnalog_v0p0p1_10.RSfetsym_0.x1.Y I5 0.0436f
C182 16to4_PriorityEncoder_v0p0p1_0.x5.x2.X I14 0.0177f
C183 frontAnalog_v0p0p1_11.x63.X frontAnalog_v0p0p1_11.RSfetsym_0.x2.Y 0.0923f
C184 frontAnalog_v0p0p1_12.x63.A VV3 0.587f
C185 w_55000_n62328# frontAnalog_v0p0p1_11.x65.A 0.658f
C186 w_55000_n73128# VDD 0.854f
C187 frontAnalog_v0p0p1_12.RSfetsym_0.QN a_59577_n73683# 0.418f
C188 frontAnalog_v0p0p1_1.x65.A VV9 0.253f
C189 VDD VV14 4.05f
C190 16to4_PriorityEncoder_v0p0p1_0.x3.x22.A a_78525_n53555# 0.209f
C191 frontAnalog_v0p0p1_13.x63.X a_59577_n68283# 0.28f
C192 frontAnalog_v0p0p1_1.x63.X a_59577_n41283# 0.28f
C193 16to4_PriorityEncoder_v0p0p1_0.x5.x19.D 16to4_PriorityEncoder_v0p0p1_0.x5.x19.X 0.0195f
C194 frontAnalog_v0p0p1_12.x63.A VDD 3.67f
C195 16to4_PriorityEncoder_v0p0p1_0.x3.x18.C I1 0.495f
C196 CLK VV3 5.47f
C197 frontAnalog_v0p0p1_10.IB a_53630_n14796# 0.473f
C198 a_57123_n20279# VDD 0.222f
C199 w_55000_n62950# frontAnalog_v0p0p1_11.x63.A 0.659f
C200 S1 R1 0.136f
C201 m3_58396_n58350# VDD 1.3f
C202 16to4_PriorityEncoder_v0p0p1_0.x5.x4.A a_78159_n39549# 0.299f
C203 a_53630_n25596# VIN 0.265f
C204 w_55000_n78528# a_55268_n79536# 0.149f
C205 w_55000_n79150# a_53630_n79596# 0.394f
C206 frontAnalog_v0p0p1_10.x65.A a_57123_n56559# 0.214f
C207 frontAnalog_v0p0p1_14.x65.A VV2 0.253f
C208 VIN VV2 2.58f
C209 w_55000_n25150# CLK 0.535f
C210 VDD CLK 73.4f
C211 a_55268_n3936# VDD 0.565f
C212 w_55000_n46128# frontAnalog_v0p0p1_10.IB 0.0216f
C213 16to4_PriorityEncoder_v0p0p1_0.x3.x2.X I7 0.0129f
C214 frontAnalog_v0p0p1_7.x65.A VV10 0.252f
C215 16to4_PriorityEncoder_v0p0p1_0.x3.x18.C I7 0.229f
C216 frontAnalog_v0p0p1_4.RSfetsym_0.QN VDD 2.56f
C217 m3_58396_n79950# R1 0.14f
C218 I12 I11 5.01f
C219 w_55000_n35328# frontAnalog_v0p0p1_7.x63.A 0.0792f
C220 frontAnalog_v0p0p1_10.RSfetsym_0.QN frontAnalog_v0p0p1_10.RSfetsym_0.x2.Y 0.018f
C221 w_55000_n83928# VIN 0.866f
C222 16to4_PriorityEncoder_v0p0p1_0.x5.x19.D 16to4_PriorityEncoder_v0p0p1_0.x5.x22.A 0.0292f
C223 a_77605_n39305# I9 0.159f
C224 frontAnalog_v0p0p1_14.x65.A S1 0.0236f
C225 frontAnalog_v0p0p1_10.RSfetsym_0.QN I5 2.02f
C226 frontAnalog_v0p0p1_11.RSfetsym_0.QN a_59577_n62883# 0.418f
C227 I6 I0 0.364f
C228 I1 I3 1.73f
C229 a_78649_n39527# 16to4_PriorityEncoder_v0p0p1_0.x5.EO 0.135f
C230 w_55000_n46128# frontAnalog_v0p0p1_8.x65.A 0.658f
C231 frontAnalog_v0p0p1_10.x63.X a_59577_n57483# 0.28f
C232 VDD R0 3.16f
C233 w_55000_n62950# VV5 0.751f
C234 a_59577_n14283# I13 0.29f
C235 frontAnalog_v0p0p1_10.IB a_53630_n30996# 0.473f
C236 frontAnalog_v0p0p1_8.x63.A a_57123_n47279# 0.212f
C237 frontAnalog_v0p0p1_1.x65.A VDD 3.45f
C238 16to4_PriorityEncoder_v0p0p1_0.x3.EI I6 2.13f
C239 16to4_PriorityEncoder_v0p0p1_0.x5.x16.X VDD 0.556f
C240 a_77605_n47345# I0 0.211f
C241 16to4_PriorityEncoder_v0p0p1_0.x5.x20.X VDD 0.473f
C242 w_55000_n46750# frontAnalog_v0p0p1_8.x63.A 0.659f
C243 frontAnalog_v0p0p1_4.RSfetsym_0.x2.Y VDD 0.926f
C244 I7 I3 1.25f
C245 I4 I6 2.39f
C246 I2 I1 8.04f
C247 16to4_PriorityEncoder_v0p0p1_0.x5.x21.B VDD 0.923f
C248 frontAnalog_v0p0p1_9.RSfetsym_0.x1.Y frontAnalog_v0p0p1_9.x63.X 0.883f
C249 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_0.x63.A 0.0858f
C250 a_55268_n47136# VV8 0.215f
C251 w_55000_n8328# VV15 0.798f
C252 frontAnalog_v0p0p1_10.x63.A frontAnalog_v0p0p1_10.x63.X 0.0301f
C253 frontAnalog_v0p0p1_10.IB a_55268_n25536# 0.0848f
C254 16to4_PriorityEncoder_v0p0p1_0.x2.A 16to4_PriorityEncoder_v0p0p1_0.x3.EO 0.02f
C255 frontAnalog_v0p0p1_1.RSfetsym_0.x2.Y I8 0.199f
C256 a_59578_n83970# I0 0.42f
C257 frontAnalog_v0p0p1_10.RSfetsym_0.x2.Y I5 0.198f
C258 w_55000_n8328# VIN 0.866f
C259 a_78649_n39527# 16to4_PriorityEncoder_v0p0p1_0.x5.GS 0.136f
C260 frontAnalog_v0p0p1_12.x65.X I2 0.446f
C261 I7 I2 0.468f
C262 w_55000_n14350# a_55268_n14736# 0.12f
C263 w_55000_n67728# CLK 0.571f
C264 VV9 VV8 3.01f
C265 a_57123_n24159# frontAnalog_v0p0p1_5.x65.X 0.119f
C266 w_55000_n84550# frontAnalog_v0p0p1_10.IB 0.0217f
C267 frontAnalog_v0p0p1_10.x65.X CLK 0.0402f
C268 frontAnalog_v0p0p1_11.x65.A VDD 3.45f
C269 w_55000_n35950# VDD 0.829f
C270 frontAnalog_v0p0p1_3.x65.A VDD 3.45f
C271 a_55268_n84936# VDD 0.565f
C272 a_55268_n30936# VV11 0.215f
C273 frontAnalog_v0p0p1_2.x63.A frontAnalog_v0p0p1_2.x65.A 3.16f
C274 w_55000_n8328# a_53630_n9396# 0.359f
C275 16to4_PriorityEncoder_v0p0p1_0.x43.A 16to4_PriorityEncoder_v0p0p1_0.x43.Y 1.52f
C276 frontAnalog_v0p0p1_8.RSfetsym_0.x1.Y VDD 0.733f
C277 frontAnalog_v0p0p1_7.x65.A CLK 2.61f
C278 16to4_PriorityEncoder_v0p0p1_0.x5.x19.D I12 0.206f
C279 frontAnalog_v0p0p1_10.x63.X m3_58396_n58350# 0.139f
C280 frontAnalog_v0p0p1_12.x63.X I2 1.85f
C281 frontAnalog_v0p0p1_8.x65.X CLK 0.0393f
C282 frontAnalog_v0p0p1_9.RSfetsym_0.x2.Y I6 0.198f
C283 frontAnalog_v0p0p1_5.x65.X a_59578_n24570# 0.436f
C284 frontAnalog_v0p0p1_15.RSfetsym_0.x1.Y I0 0.0436f
C285 16to4_PriorityEncoder_v0p0p1_0.x5.x15.X VDD 0.272f
C286 a_55268_n14736# VIN 0.177f
C287 frontAnalog_v0p0p1_10.x63.X CLK 0.785f
C288 frontAnalog_v0p0p1_7.x65.X I9 0.445f
C289 a_53630_n74196# VV3 0.28f
C290 w_55000_n8950# frontAnalog_v0p0p1_10.IB 0.0217f
C291 16to4_PriorityEncoder_v0p0p1_0.x3.EI a_77605_n51335# 0.122f
C292 a_57123_n13359# frontAnalog_v0p0p1_3.x65.X 0.119f
C293 16to4_PriorityEncoder_v0p0p1_0.x3.EI 16to4_PriorityEncoder_v0p0p1_0.x3.x4.A 0.547f
C294 a_57123_n51159# VDD 0.224f
C295 16to4_PriorityEncoder_v0p0p1_0.x3.A0 16to4_PriorityEncoder_v0p0p1_0.x3.x20.X 0.0149f
C296 w_55000_n46750# VIN 0.737f
C297 VDD I6 5.5f
C298 a_53630_n74196# VDD 0.134f
C299 16to4_PriorityEncoder_v0p0p1_0.x5.x4.A VDD 1.92f
C300 VDD VV8 4.18f
C301 w_55000_n62328# a_55268_n63336# 0.149f
C302 w_55000_n62950# a_53630_n63396# 0.394f
C303 a_59577_n52083# I6 0.29f
C304 a_77605_n47345# VDD 0.152f
C305 16to4_PriorityEncoder_v0p0p1_0.x5.x14.A 16to4_PriorityEncoder_v0p0p1_0.x5.A2 0.074f
C306 16to4_PriorityEncoder_v0p0p1_0.x5.x21.X VDD 0.514f
C307 frontAnalog_v0p0p1_0.x65.A VV15 0.253f
C308 frontAnalog_v0p0p1_7.x63.X I9 1.73f
C309 frontAnalog_v0p0p1_0.x65.A VIN 0.655f
C310 w_55000_n24528# frontAnalog_v0p0p1_5.x65.A 0.658f
C311 w_55000_n51528# w_55000_n52150# 0.327f
C312 a_55268_n30936# VIN 0.177f
C313 w_55000_n78528# VDD 0.854f
C314 VDD I11 9.86f
C315 frontAnalog_v0p0p1_3.x65.X a_59578_n13770# 0.436f
C316 a_57123_n83559# S0 0.119f
C317 a_59578_n83970# VDD 0.0213f
C318 frontAnalog_v0p0p1_5.x65.X frontAnalog_v0p0p1_5.RSfetsym_0.x1.Y 0.182f
C319 a_55268_n79536# VV2 0.215f
C320 frontAnalog_v0p0p1_15.RSfetsym_0.QN I0 2.02f
C321 w_55000_n25150# frontAnalog_v0p0p1_5.x63.A 0.659f
C322 frontAnalog_v0p0p1_5.x63.A VDD 3.67f
C323 frontAnalog_v0p0p1_10.IB VV4 3.7f
C324 m3_58396_n69150# VDD 1.3f
C325 w_55000_n35950# frontAnalog_v0p0p1_7.x65.A 0.0988f
C326 16to4_PriorityEncoder_v0p0p1_0.x3.EI 16to4_PriorityEncoder_v0p0p1_0.x3.x16.X 0.076f
C327 a_77605_n40069# I13 0.16f
C328 VDD OUT0 6.72f
C329 16to4_PriorityEncoder_v0p0p1_0.x2.A 16to4_PriorityEncoder_v0p0p1_0.x21.A 0.0121f
C330 a_59577_n84483# I0 0.29f
C331 w_55000_n30550# CLK 0.535f
C332 w_55000_n46128# a_53630_n47196# 0.359f
C333 frontAnalog_v0p0p1_2.x65.X VDD 3.55f
C334 w_55000_n51528# frontAnalog_v0p0p1_10.IB 0.0216f
C335 16to4_PriorityEncoder_v0p0p1_0.x5.x16.C I12 0.202f
C336 I10 I9 7.73f
C337 frontAnalog_v0p0p1_4.RSfetsym_0.QN a_59578_n19170# 0.255f
C338 16to4_PriorityEncoder_v0p0p1_0.x5.x22.A I15 0.0853f
C339 a_59577_n73683# I2 0.29f
C340 frontAnalog_v0p0p1_3.x63.X m3_58396_n15150# 0.139f
C341 a_53630_n41796# a_55268_n41736# 0.015f
C342 frontAnalog_v0p0p1_8.x65.X frontAnalog_v0p0p1_8.RSfetsym_0.x1.Y 0.182f
C343 frontAnalog_v0p0p1_2.x63.A VIN 0.187f
C344 w_55000_n13728# w_55000_n14350# 0.327f
C345 w_55000_n2928# VDD 0.854f
C346 frontAnalog_v0p0p1_5.RSfetsym_0.x1.Y frontAnalog_v0p0p1_5.x63.X 0.883f
C347 CLK VV10 6.39f
C348 16to4_PriorityEncoder_v0p0p1_0.x3.EI 16to4_PriorityEncoder_v0p0p1_0.x3.x17.A 0.02f
C349 a_78065_n49349# VDD 0.156f
C350 16to4_PriorityEncoder_v0p0p1_0.x3.EI a_77637_n49127# 0.0829f
C351 w_55000_n41350# VV9 0.751f
C352 frontAnalog_v0p0p1_0.x63.A a_55268_n9336# 1.24f
C353 frontAnalog_v0p0p1_1.x65.X a_59578_n40770# 0.436f
C354 frontAnalog_v0p0p1_15.x65.A CLK 2.62f
C355 a_57123_n29559# frontAnalog_v0p0p1_6.x65.X 0.119f
C356 w_55000_n84550# VV1 0.751f
C357 a_82906_n47995# 16to4_PriorityEncoder_v0p0p1_0.x3.A1 0.121f
C358 frontAnalog_v0p0p1_3.x65.X frontAnalog_v0p0p1_3.RSfetsym_0.x1.Y 0.182f
C359 a_77605_n51335# VDD 0.435f
C360 frontAnalog_v0p0p1_15.RSfetsym_0.x1.Y VDD 0.733f
C361 16to4_PriorityEncoder_v0p0p1_0.x3.x4.A VDD 1.55f
C362 frontAnalog_v0p0p1_5.x65.X frontAnalog_v0p0p1_5.RSfetsym_0.QN 2.28f
C363 VIN VV13 2.58f
C364 16to4_PriorityEncoder_v0p0p1_0.x3.x19.D I0 0.122f
C365 frontAnalog_v0p0p1_2.x63.X VDD 3.16f
C366 frontAnalog_v0p0p1_4.x65.X frontAnalog_v0p0p1_4.x63.X 0.136f
C367 a_53630_n52596# CLK 0.0136f
C368 frontAnalog_v0p0p1_10.x63.A CLK 1.81f
C369 frontAnalog_v0p0p1_10.x65.A VV6 0.253f
C370 frontAnalog_v0p0p1_13.x65.A VV4 0.253f
C371 a_78097_n45737# 16to4_PriorityEncoder_v0p0p1_0.x5.x20.X 0.137f
C372 frontAnalog_v0p0p1_15.RSfetsym_0.x2.Y S0 0.526f
C373 16to4_PriorityEncoder_v0p0p1_0.x3.EI a_78649_n47567# 0.181f
C374 16to4_PriorityEncoder_v0p0p1_0.x3.EI 16to4_PriorityEncoder_v0p0p1_0.x3.x19.D 1.93f
C375 frontAnalog_v0p0p1_5.x63.X a_57123_n25679# 0.121f
C376 w_55000_n73128# frontAnalog_v0p0p1_12.x63.A 0.0792f
C377 frontAnalog_v0p0p1_2.x65.A frontAnalog_v0p0p1_10.IB 0.0352f
C378 16to4_PriorityEncoder_v0p0p1_0.x42.A 16to4_PriorityEncoder_v0p0p1_0.x43.A 0.392f
C379 a_53630_n41796# VIN 0.265f
C380 w_55000_n13728# VIN 0.866f
C381 16to4_PriorityEncoder_v0p0p1_0.x5.x21.B a_78097_n45737# 0.186f
C382 a_59577_n35883# I9 0.29f
C383 16to4_PriorityEncoder_v0p0p1_0.x5.x19.D VDD 3.27f
C384 16to4_PriorityEncoder_v0p0p1_0.x3.x19.D I4 0.206f
C385 frontAnalog_v0p0p1_4.RSfetsym_0.QN frontAnalog_v0p0p1_4.RSfetsym_0.x1.Y 0.17f
C386 frontAnalog_v0p0p1_6.x65.X a_59578_n29970# 0.436f
C387 a_77605_n43295# 16to4_PriorityEncoder_v0p0p1_0.x5.x16.X 0.0121f
C388 16to4_PriorityEncoder_v0p0p1_0.x36.Y OUT2 8.68f
C389 I14 I9 0.258f
C390 I13 I10 0.644f
C391 a_55268_n63336# VDD 0.565f
C392 frontAnalog_v0p0p1_9.RSfetsym_0.QN frontAnalog_v0p0p1_9.RSfetsym_0.x2.Y 0.018f
C393 frontAnalog_v0p0p1_3.RSfetsym_0.x1.Y frontAnalog_v0p0p1_3.x63.X 0.883f
C394 a_78065_n41309# 16to4_PriorityEncoder_v0p0p1_0.x5.A2 0.144f
C395 16to4_PriorityEncoder_v0p0p1_0.x3.x2.X a_77605_n48109# 0.134f
C396 16to4_PriorityEncoder_v0p0p1_0.x3.EI 16to4_PriorityEncoder_v0p0p1_0.x3.x15.X 0.0245f
C397 frontAnalog_v0p0p1_5.RSfetsym_0.QN frontAnalog_v0p0p1_5.x63.X 0.378f
C398 frontAnalog_v0p0p1_5.x65.X frontAnalog_v0p0p1_5.RSfetsym_0.x2.Y 0.526f
C399 a_59578_n78570# S1 0.436f
C400 w_55000_n73128# CLK 0.571f
C401 16to4_PriorityEncoder_v0p0p1_0.x2.A 16to4_PriorityEncoder_v0p0p1_0.x2.X 0.0402f
C402 frontAnalog_v0p0p1_9.x65.A VDD 3.45f
C403 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_8.x63.A 0.0926f
C404 frontAnalog_v0p0p1_10.IB a_53630_n36396# 0.473f
C405 CLK VV14 6.32f
C406 VV6 VV5 4.54f
C407 w_55000_n41350# VDD 0.829f
C408 frontAnalog_v0p0p1_3.x65.X frontAnalog_v0p0p1_3.RSfetsym_0.QN 2.28f
C409 frontAnalog_v0p0p1_12.x63.A CLK 1.81f
C410 16to4_PriorityEncoder_v0p0p1_0.x3.x16.X VDD 0.505f
C411 frontAnalog_v0p0p1_15.RSfetsym_0.QN VDD 2.56f
C412 frontAnalog_v0p0p1_9.RSfetsym_0.QN VDD 2.56f
C413 I15 I12 0.786f
C414 frontAnalog_v0p0p1_14.x63.A R1 0.0301f
C415 w_55000_n8950# a_55268_n9336# 0.12f
C416 w_55000_n51528# VV7 0.798f
C417 frontAnalog_v0p0p1_10.IB VV11 3.7f
C418 frontAnalog_v0p0p1_4.RSfetsym_0.x1.Y frontAnalog_v0p0p1_4.RSfetsym_0.x2.Y 0.0254f
C419 frontAnalog_v0p0p1_8.x63.A frontAnalog_v0p0p1_8.x65.A 3.16f
C420 16to4_PriorityEncoder_v0p0p1_0.x5.x1.X 16to4_PriorityEncoder_v0p0p1_0.x5.x2.X 0.129f
C421 w_55000_n35950# VV10 0.751f
C422 a_53630_n3996# VV16 0.28f
C423 frontAnalog_v0p0p1_9.RSfetsym_0.QN a_59577_n52083# 0.418f
C424 frontAnalog_v0p0p1_3.x63.X a_57123_n14879# 0.121f
C425 a_55268_n3936# CLK 0.236f
C426 a_59577_n84483# VDD 0.0173f
C427 frontAnalog_v0p0p1_5.x63.X frontAnalog_v0p0p1_5.RSfetsym_0.x2.Y 0.0923f
C428 frontAnalog_v0p0p1_15.x65.A a_55268_n84936# 0.461f
C429 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_13.x63.A 0.0926f
C430 16to4_PriorityEncoder_v0p0p1_0.x3.x17.A VDD 1.34f
C431 a_77637_n49127# VDD 0.218f
C432 frontAnalog_v0p0p1_6.x65.X frontAnalog_v0p0p1_6.RSfetsym_0.x1.Y 0.182f
C433 frontAnalog_v0p0p1_10.IB a_55268_n41736# 0.0848f
C434 w_55000_n14350# frontAnalog_v0p0p1_10.IB 0.0217f
C435 frontAnalog_v0p0p1_14.x63.A frontAnalog_v0p0p1_14.x65.A 3.16f
C436 frontAnalog_v0p0p1_14.x63.A VIN 0.19f
C437 a_53630_n36396# a_55268_n36336# 0.015f
C438 frontAnalog_v0p0p1_3.RSfetsym_0.QN frontAnalog_v0p0p1_3.x63.X 0.378f
C439 frontAnalog_v0p0p1_3.x65.X frontAnalog_v0p0p1_3.RSfetsym_0.x2.Y 0.526f
C440 VV3 VV2 4.95f
C441 I14 I13 10.5f
C442 w_55000_n52150# VIN 0.737f
C443 frontAnalog_v0p0p1_14.RSfetsym_0.x1.Y S1 0.182f
C444 a_59577_n3483# VDD 0.0173f
C445 CLK R0 0.786f
C446 16to4_PriorityEncoder_v0p0p1_0.x3.x16.C I0 0.12f
C447 a_57123_n72759# VDD 0.224f
C448 16to4_PriorityEncoder_v0p0p1_0.x3.EI 16to4_PriorityEncoder_v0p0p1_0.x3.x22.A 0.0483f
C449 16to4_PriorityEncoder_v0p0p1_0.x5.x19.C I12 0.405f
C450 16to4_PriorityEncoder_v0p0p1_0.x5.x2.X 16to4_PriorityEncoder_v0p0p1_0.x5.EO 0.0749f
C451 w_55000_n24528# a_55268_n25536# 0.149f
C452 w_55000_n25150# a_53630_n25596# 0.394f
C453 a_53630_n25596# VDD 0.134f
C454 frontAnalog_v0p0p1_1.x65.A CLK 2.61f
C455 a_77605_n43295# 16to4_PriorityEncoder_v0p0p1_0.x5.x15.X 0.0951f
C456 VDD VV2 4.22f
C457 a_78649_n47567# VDD 0.235f
C458 16to4_PriorityEncoder_v0p0p1_0.x3.EI 16to4_PriorityEncoder_v0p0p1_0.x3.x16.C 2.08f
C459 16to4_PriorityEncoder_v0p0p1_0.x3.x19.D VDD 1.32f
C460 frontAnalog_v0p0p1_15.x63.A a_57123_n85079# 0.212f
C461 16to4_PriorityEncoder_v0p0p1_0.x5.GS 16to4_PriorityEncoder_v0p0p1_0.x43.A 0.0166f
C462 frontAnalog_v0p0p1_4.RSfetsym_0.QN frontAnalog_v0p0p1_4.RSfetsym_0.x2.Y 0.018f
C463 16to4_PriorityEncoder_v0p0p1_0.x5.x16.C VDD 2.83f
C464 frontAnalog_v0p0p1_6.RSfetsym_0.x1.Y frontAnalog_v0p0p1_6.x63.X 0.883f
C465 16to4_PriorityEncoder_v0p0p1_0.x3.x16.C I4 0.202f
C466 frontAnalog_v0p0p1_1.x65.X I8 0.445f
C467 w_55000_n83928# VDD 0.854f
C468 frontAnalog_v0p0p1_10.IB VV15 4.34f
C469 a_78097_n45737# 16to4_PriorityEncoder_v0p0p1_0.x5.x21.X 0.109f
C470 frontAnalog_v0p0p1_6.x65.A a_55268_n30936# 0.461f
C471 frontAnalog_v0p0p1_3.x63.X frontAnalog_v0p0p1_3.RSfetsym_0.x2.Y 0.0923f
C472 VDD S1 3.55f
C473 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_14.x65.A 0.0352f
C474 frontAnalog_v0p0p1_10.IB VIN 32.9f
C475 16to4_PriorityEncoder_v0p0p1_0.x5.x17.A 16to4_PriorityEncoder_v0p0p1_0.x5.A2 0.047f
C476 frontAnalog_v0p0p1_11.x63.A VV5 0.587f
C477 16to4_PriorityEncoder_v0p0p1_0.x3.x15.X VDD 0.26f
C478 frontAnalog_v0p0p1_5.RSfetsym_0.QN a_59577_n25083# 0.418f
C479 frontAnalog_v0p0p1_3.x65.A VV14 0.253f
C480 frontAnalog_v0p0p1_11.x65.X I4 0.446f
C481 a_59578_n46170# VDD 0.0213f
C482 a_59578_n73170# VDD 0.0213f
C483 frontAnalog_v0p0p1_13.x63.A frontAnalog_v0p0p1_13.x65.A 3.16f
C484 frontAnalog_v0p0p1_4.x63.X a_59577_n19683# 0.28f
C485 frontAnalog_v0p0p1_1.RSfetsym_0.QN a_59578_n40770# 0.255f
C486 frontAnalog_v0p0p1_5.x65.A VV12 0.253f
C487 frontAnalog_v0p0p1_6.x65.X frontAnalog_v0p0p1_6.RSfetsym_0.QN 2.28f
C488 m3_58396_n79950# VDD 1.3f
C489 frontAnalog_v0p0p1_4.x63.A VV13 0.587f
C490 w_55000_n19750# VV13 0.751f
C491 16to4_PriorityEncoder_v0p0p1_0.x2.A 16to4_PriorityEncoder_v0p0p1_0.x3.A0 0.398f
C492 frontAnalog_v0p0p1_8.x65.A VIN 0.654f
C493 frontAnalog_v0p0p1_14.RSfetsym_0.QN S1 2.28f
C494 16to4_PriorityEncoder_v0p0p1_0.x5.x16.X 16to4_PriorityEncoder_v0p0p1_0.x5.x21.B 0.0218f
C495 16to4_PriorityEncoder_v0p0p1_0.x5.x21.B 16to4_PriorityEncoder_v0p0p1_0.x5.x20.X 0.0561f
C496 frontAnalog_v0p0p1_11.x65.A CLK 2.61f
C497 w_55000_n35950# CLK 0.535f
C498 w_55000_n46750# a_55268_n47136# 0.12f
C499 w_55000_n56928# frontAnalog_v0p0p1_10.IB 0.0216f
C500 frontAnalog_v0p0p1_6.x63.X a_57123_n31079# 0.121f
C501 frontAnalog_v0p0p1_0.x65.A a_57123_n7959# 0.214f
C502 frontAnalog_v0p0p1_3.x65.A CLK 2.61f
C503 a_55268_n84936# CLK 0.236f
C504 I12 I8 0.558f
C505 frontAnalog_v0p0p1_9.RSfetsym_0.x1.Y frontAnalog_v0p0p1_9.RSfetsym_0.x2.Y 0.0254f
C506 frontAnalog_v0p0p1_10.IB a_53630_n9396# 0.473f
C507 w_55000_n8328# VDD 0.854f
C508 a_55268_n36336# VIN 0.177f
C509 frontAnalog_v0p0p1_11.x63.X I4 1.85f
C510 w_55000_n73128# a_53630_n74196# 0.359f
C511 frontAnalog_v0p0p1_14.RSfetsym_0.x2.Y I1 0.198f
C512 frontAnalog_v0p0p1_6.x65.X frontAnalog_v0p0p1_6.RSfetsym_0.x2.Y 0.526f
C513 frontAnalog_v0p0p1_6.RSfetsym_0.QN frontAnalog_v0p0p1_6.x63.X 0.378f
C514 16to4_PriorityEncoder_v0p0p1_0.x5.x18.C I12 0.432f
C515 a_59578_n40770# VDD 0.0213f
C516 a_55268_n68736# VV4 0.215f
C517 frontAnalog_v0p0p1_3.RSfetsym_0.QN a_59577_n14283# 0.418f
C518 frontAnalog_v0p0p1_13.x65.A VIN 0.655f
C519 frontAnalog_v0p0p1_9.RSfetsym_0.x1.Y VDD 0.733f
C520 w_55000_n73750# frontAnalog_v0p0p1_12.x65.A 0.0988f
C521 16to4_PriorityEncoder_v0p0p1_0.x5.GS 16to4_PriorityEncoder_v0p0p1_0.x42.A 0.098f
C522 frontAnalog_v0p0p1_12.RSfetsym_0.x1.Y VDD 0.733f
C523 16to4_PriorityEncoder_v0p0p1_0.x3.EI a_78097_n53777# 0.106f
C524 a_77605_n45765# I13 0.193f
C525 16to4_PriorityEncoder_v0p0p1_0.x3.x22.A VDD 3.23f
C526 frontAnalog_v0p0p1_1.x63.X m3_58396_n42150# 0.139f
C527 CLK I6 0.01f
C528 a_53630_n74196# CLK 0.0136f
C529 CLK VV8 5.47f
C530 VDD I15 9.55f
C531 w_55000_n40728# frontAnalog_v0p0p1_1.x63.A 0.0792f
C532 16to4_PriorityEncoder_v0p0p1_0.x3.x16.C VDD 0.834f
C533 a_77605_n43545# VDD 0.571f
C534 w_55000_n19128# VIN 0.868f
C535 frontAnalog_v0p0p1_6.x63.A VV11 0.587f
C536 frontAnalog_v0p0p1_0.x63.A frontAnalog_v0p0p1_0.x63.X 0.0301f
C537 frontAnalog_v0p0p1_6.x63.X frontAnalog_v0p0p1_6.RSfetsym_0.x2.Y 0.0923f
C538 16to4_PriorityEncoder_v0p0p1_0.x5.x15.X 16to4_PriorityEncoder_v0p0p1_0.x5.x16.X 0.253f
C539 frontAnalog_v0p0p1_11.x65.X VDD 3.55f
C540 VIN VV7 2.61f
C541 a_55268_n14736# VDD 0.565f
C542 w_55000_n78528# CLK 0.571f
C543 a_57123_n47279# VDD 0.222f
C544 frontAnalog_v0p0p1_10.IB a_53630_n68796# 0.473f
C545 a_57123_n74279# VDD 0.222f
C546 CLK I11 0.01f
C547 16to4_PriorityEncoder_v0p0p1_0.x3.x19.C I0 0.12f
C548 16to4_PriorityEncoder_v0p0p1_0.x3.A2 a_78065_n49349# 0.144f
C549 a_77639_n42341# I15 0.192f
C550 a_53630_n79596# VIN 0.265f
C551 frontAnalog_v0p0p1_8.x65.X a_59578_n46170# 0.436f
C552 w_55000_n46750# VDD 0.829f
C553 16to4_PriorityEncoder_v0p0p1_0.x5.x22.A 16to4_PriorityEncoder_v0p0p1_0.x5.A2 0.0408f
C554 16to4_PriorityEncoder_v0p0p1_0.x3.EI 16to4_PriorityEncoder_v0p0p1_0.x3.x19.C 1.71f
C555 frontAnalog_v0p0p1_5.x63.A CLK 1.81f
C556 frontAnalog_v0p0p1_0.RSfetsym_0.QN I15 0.0512f
C557 frontAnalog_v0p0p1_12.RSfetsym_0.QN VDD 2.56f
C558 16to4_PriorityEncoder_v0p0p1_0.x5.EO 16to4_PriorityEncoder_v0p0p1_0.x5.GS 0.927f
C559 16to4_PriorityEncoder_v0p0p1_0.x5.x19.C VDD 2.86f
C560 16to4_PriorityEncoder_v0p0p1_0.x5.A2 16to4_PriorityEncoder_v0p0p1_0.x35.A 0.0138f
C561 16to4_PriorityEncoder_v0p0p1_0.x3.x19.C I4 0.405f
C562 frontAnalog_v0p0p1_14.x63.A a_55268_n79536# 1.24f
C563 16to4_PriorityEncoder_v0p0p1_0.x3.x16.X 16to4_PriorityEncoder_v0p0p1_0.x3.x21.B 0.0218f
C564 frontAnalog_v0p0p1_11.x63.X VDD 3.16f
C565 16to4_PriorityEncoder_v0p0p1_0.x5.x20.X 16to4_PriorityEncoder_v0p0p1_0.x5.x21.X 0.122f
C566 frontAnalog_v0p0p1_2.x65.X CLK 0.0302f
C567 m3_58396_n9750# VDD 1.3f
C568 a_59577_n62883# I4 0.29f
C569 16to4_PriorityEncoder_v0p0p1_0.x5.x16.X I11 0.0148f
C570 16to4_PriorityEncoder_v0p0p1_0.x5.x21.B 16to4_PriorityEncoder_v0p0p1_0.x5.x21.X 0.0197f
C571 frontAnalog_v0p0p1_0.x65.A VDD 3.45f
C572 w_55000_n29928# a_53630_n30996# 0.359f
C573 a_55268_n30936# VDD 0.565f
C574 VIN VV1 2.01f
C575 16to4_PriorityEncoder_v0p0p1_0.x3.EI a_77637_n50057# 0.0878f
C576 I13 I5 0.0641f
C577 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_4.x63.A 0.0926f
C578 w_55000_n2928# CLK 0.57f
C579 frontAnalog_v0p0p1_6.RSfetsym_0.QN a_59577_n30483# 0.418f
C580 w_55000_n3550# a_53630_n3996# 0.394f
C581 16to4_PriorityEncoder_v0p0p1_0.x3.x11.X VDD 0.507f
C582 w_55000_n2928# a_55268_n3936# 0.149f
C583 frontAnalog_v0p0p1_1.RSfetsym_0.QN I8 2.02f
C584 w_55000_n19750# frontAnalog_v0p0p1_10.IB 0.0217f
C585 a_77605_n44527# I9 0.147f
C586 frontAnalog_v0p0p1_6.x63.A a_57123_n31079# 0.212f
C587 16to4_PriorityEncoder_v0p0p1_0.x3.EI a_77605_n51585# 0.14f
C588 frontAnalog_v0p0p1_6.x63.A VIN 0.187f
C589 16to4_PriorityEncoder_v0p0p1_0.x5.x21.B I11 0.0112f
C590 a_77605_n52567# I1 0.147f
C591 a_53630_n63396# VV5 0.28f
C592 w_55000_n57550# VIN 0.737f
C593 frontAnalog_v0p0p1_8.RSfetsym_0.x2.Y VDD 0.926f
C594 16to4_PriorityEncoder_v0p0p1_0.x3.A0 16to4_PriorityEncoder_v0p0p1_0.x3.x19.X 0.0123f
C595 frontAnalog_v0p0p1_12.RSfetsym_0.x2.Y VDD 0.926f
C596 a_55268_n9336# VV15 0.215f
C597 a_53630_n57996# VIN 0.265f
C598 frontAnalog_v0p0p1_9.x63.A a_55268_n52536# 1.24f
C599 a_78097_n53777# VDD 0.219f
C600 a_55268_n9336# VIN 0.177f
C601 a_57123_n24159# VDD 0.224f
C602 a_53630_n41796# VV9 0.28f
C603 a_53630_n20196# VV13 0.28f
C604 frontAnalog_v0p0p1_2.x63.X CLK 0.785f
C605 frontAnalog_v0p0p1_10.IB a_55268_n79536# 0.0848f
C606 m3_58396_n20550# I12 0.0416f
C607 16to4_PriorityEncoder_v0p0p1_0.x3.x2.X I0 0.0265f
C608 frontAnalog_v0p0p1_13.x63.A a_55268_n68736# 1.24f
C609 16to4_PriorityEncoder_v0p0p1_0.x3.x18.C I0 0.119f
C610 a_55268_n25536# VV12 0.215f
C611 w_55000_n56928# w_55000_n57550# 0.327f
C612 frontAnalog_v0p0p1_2.x63.A VDD 3.67f
C613 VDD I8 7.79f
C614 16to4_PriorityEncoder_v0p0p1_0.x3.x19.D 16to4_PriorityEncoder_v0p0p1_0.x3.x21.B 0.151f
C615 frontAnalog_v0p0p1_6.x65.A frontAnalog_v0p0p1_6.x65.X 0.0236f
C616 a_53630_n47196# VIN 0.265f
C617 w_55000_n56928# a_53630_n57996# 0.359f
C618 frontAnalog_v0p0p1_15.RSfetsym_0.x1.Y R0 0.883f
C619 16to4_PriorityEncoder_v0p0p1_0.x3.EI 16to4_PriorityEncoder_v0p0p1_0.x3.x18.C 1.56f
C620 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_6.x65.A 0.0352f
C621 a_55268_n63336# CLK 0.236f
C622 16to4_PriorityEncoder_v0p0p1_0.x3.x2.X I4 0.0262f
C623 16to4_PriorityEncoder_v0p0p1_0.x3.A2 16to4_PriorityEncoder_v0p0p1_0.x3.x17.A 0.047f
C624 a_59578_n24570# VDD 0.0213f
C625 a_53630_n9396# a_55268_n9336# 0.015f
C626 16to4_PriorityEncoder_v0p0p1_0.x5.x18.C VDD 2.22f
C627 a_78349_n43045# 16to4_PriorityEncoder_v0p0p1_0.x1.A 0.151f
C628 16to4_PriorityEncoder_v0p0p1_0.x5.A2 16to4_PriorityEncoder_v0p0p1_0.x34.A 0.0422f
C629 16to4_PriorityEncoder_v0p0p1_0.x3.x18.C I4 0.432f
C630 frontAnalog_v0p0p1_9.x65.A CLK 2.61f
C631 w_55000_n83928# frontAnalog_v0p0p1_15.x65.A 0.658f
C632 16to4_PriorityEncoder_v0p0p1_0.x3.EI 16to4_PriorityEncoder_v0p0p1_0.x3.GS 0.123f
C633 16to4_PriorityEncoder_v0p0p1_0.x5.x16.C a_77605_n43295# 0.0949f
C634 VDD VV13 4.13f
C635 a_59578_n29970# I10 0.42f
C636 16to4_PriorityEncoder_v0p0p1_0.x3.x19.C VDD 1.19f
C637 w_55000_n41350# CLK 0.535f
C638 w_55000_n62328# frontAnalog_v0p0p1_10.IB 0.0216f
C639 I3 I0 0.677f
C640 frontAnalog_v0p0p1_1.RSfetsym_0.QN a_59577_n41283# 0.418f
C641 I5 I1 0.378f
C642 frontAnalog_v0p0p1_10.IB a_55268_n57936# 0.0848f
C643 a_59577_n62883# VDD 0.0173f
C644 a_82906_n47995# 16to4_PriorityEncoder_v0p0p1_0.x1.X 0.12f
C645 w_55000_n19128# frontAnalog_v0p0p1_4.x63.A 0.0792f
C646 w_55000_n84550# frontAnalog_v0p0p1_15.x63.A 0.659f
C647 a_57123_n40359# frontAnalog_v0p0p1_1.x65.X 0.119f
C648 w_55000_n19128# w_55000_n19750# 0.327f
C649 a_53630_n41796# VDD 0.134f
C650 frontAnalog_v0p0p1_12.x65.A a_55268_n74136# 0.461f
C651 w_55000_n13728# VDD 0.854f
C652 frontAnalog_v0p0p1_8.RSfetsym_0.QN I7 2.02f
C653 a_55268_n68736# VIN 0.177f
C654 16to4_PriorityEncoder_v0p0p1_0.x3.EI I3 1.97f
C655 w_55000_n73750# a_55268_n74136# 0.12f
C656 16to4_PriorityEncoder_v0p0p1_0.x5.x4.A I11 0.0406f
C657 a_77637_n50057# VDD 0.234f
C658 16to4_PriorityEncoder_v0p0p1_0.x5.x19.D 16to4_PriorityEncoder_v0p0p1_0.x5.x21.B 0.151f
C659 I4 I3 5.52f
C660 I2 I0 2.46f
C661 a_77605_n51585# VDD 0.432f
C662 I7 I5 1.12f
C663 a_77605_n53805# I5 0.193f
C664 frontAnalog_v0p0p1_15.RSfetsym_0.QN R0 0.378f
C665 w_55000_n41350# frontAnalog_v0p0p1_1.x65.A 0.0988f
C666 frontAnalog_v0p0p1_10.IB a_55268_n47136# 0.0848f
C667 frontAnalog_v0p0p1_4.x65.A VIN 0.657f
C668 16to4_PriorityEncoder_v0p0p1_0.x3.EI 16to4_PriorityEncoder_v0p0p1_0.x5.A2 0.507f
C669 16to4_PriorityEncoder_v0p0p1_0.x3.EI I2 1.27f
C670 a_59577_n41283# VDD 0.0173f
C671 frontAnalog_v0p0p1_5.RSfetsym_0.x1.Y VDD 0.733f
C672 frontAnalog_v0p0p1_8.x65.X frontAnalog_v0p0p1_8.RSfetsym_0.x2.Y 0.526f
C673 frontAnalog_v0p0p1_8.RSfetsym_0.QN frontAnalog_v0p0p1_8.x63.X 0.378f
C674 I2 I4 0.848f
C675 a_59577_n84483# R0 0.28f
C676 frontAnalog_v0p0p1_6.RSfetsym_0.x1.Y I10 0.0436f
C677 a_53630_n25596# CLK 0.0136f
C678 16to4_PriorityEncoder_v0p0p1_0.x3.x22.A 16to4_PriorityEncoder_v0p0p1_0.x3.x21.B 0.064f
C679 16to4_PriorityEncoder_v0p0p1_0.x3.A0 a_78525_n53555# 0.149f
C680 frontAnalog_v0p0p1_10.IB VV9 3.69f
C681 w_55000_n24528# VIN 0.866f
C682 frontAnalog_v0p0p1_8.x65.A a_55268_n47136# 0.461f
C683 CLK VV2 6.06f
C684 VDD OUT2 6.68f
C685 a_53630_n79596# a_55268_n79536# 0.015f
C686 frontAnalog_v0p0p1_11.x65.A a_55268_n63336# 0.461f
C687 16to4_PriorityEncoder_v0p0p1_0.x3.x20.X 16to4_PriorityEncoder_v0p0p1_0.x3.x21.X 0.122f
C688 16to4_PriorityEncoder_v0p0p1_0.x3.x2.X VDD 0.371f
C689 frontAnalog_v0p0p1_3.x65.X VDD 3.55f
C690 a_57123_n79679# R1 0.121f
C691 w_55000_n83928# CLK 0.571f
C692 16to4_PriorityEncoder_v0p0p1_0.x3.x18.C VDD 0.691f
C693 frontAnalog_v0p0p1_8.x65.X I8 0.0353f
C694 frontAnalog_v0p0p1_14.x63.A VDD 3.67f
C695 CLK S1 0.0415f
C696 frontAnalog_v0p0p1_10.IB a_53630_n20196# 0.473f
C697 a_57123_n25679# VDD 0.222f
C698 frontAnalog_v0p0p1_14.x65.A a_57123_n78159# 0.214f
C699 a_78525_n45515# 16to4_PriorityEncoder_v0p0p1_0.x2.A 0.148f
C700 w_55000_n52150# VDD 0.829f
C701 16to4_PriorityEncoder_v0p0p1_0.x3.EI 16to4_PriorityEncoder_v0p0p1_0.x3.EO 0.187f
C702 16to4_PriorityEncoder_v0p0p1_0.x3.GS VDD 0.608f
C703 16to4_PriorityEncoder_v0p0p1_0.x3.x4.A a_77605_n47345# 0.0112f
C704 a_82906_n43855# 16to4_PriorityEncoder_v0p0p1_0.x34.A 0.12f
C705 16to4_PriorityEncoder_v0p0p1_0.x3.A2 16to4_PriorityEncoder_v0p0p1_0.x3.x22.A 0.0408f
C706 frontAnalog_v0p0p1_5.RSfetsym_0.QN VDD 2.56f
C707 frontAnalog_v0p0p1_10.IB VV3 3.7f
C708 frontAnalog_v0p0p1_2.RSfetsym_0.QN a_59578_n2970# 0.255f
C709 a_59578_n67770# I3 0.42f
C710 frontAnalog_v0p0p1_1.x63.A frontAnalog_v0p0p1_1.x63.X 0.0301f
C711 16to4_PriorityEncoder_v0p0p1_0.x5.x16.C 16to4_PriorityEncoder_v0p0p1_0.x5.x16.X 0.07f
C712 frontAnalog_v0p0p1_3.x63.X VDD 3.16f
C713 m3_58396_n20550# VDD 1.3f
C714 16to4_PriorityEncoder_v0p0p1_0.x5.x19.D 16to4_PriorityEncoder_v0p0p1_0.x5.x4.A 0.0516f
C715 frontAnalog_v0p0p1_6.RSfetsym_0.QN I10 2.02f
C716 frontAnalog_v0p0p1_11.RSfetsym_0.QN I5 0.0512f
C717 VDD I3 3.87f
C718 w_55000_n3550# VV16 0.751f
C719 w_55000_n30550# a_55268_n30936# 0.12f
C720 frontAnalog_v0p0p1_6.x65.X VDD 3.55f
C721 a_53630_n68796# a_55268_n68736# 0.015f
C722 frontAnalog_v0p0p1_9.x65.A a_57123_n51159# 0.214f
C723 w_55000_n8328# CLK 0.571f
C724 w_55000_n25150# frontAnalog_v0p0p1_10.IB 0.0217f
C725 frontAnalog_v0p0p1_10.IB VDD 47.1f
C726 a_57123_n34959# frontAnalog_v0p0p1_7.x65.X 0.119f
C727 frontAnalog_v0p0p1_6.x63.A frontAnalog_v0p0p1_6.x65.A 3.16f
C728 16to4_PriorityEncoder_v0p0p1_0.x5.x19.C a_77605_n43295# 0.173f
C729 frontAnalog_v0p0p1_3.RSfetsym_0.QN I14 0.0554f
C730 w_55000_n62950# VIN 0.737f
C731 frontAnalog_v0p0p1_14.RSfetsym_0.x2.Y R1 0.0923f
C732 frontAnalog_v0p0p1_13.x65.A a_57123_n67359# 0.214f
C733 16to4_PriorityEncoder_v0p0p1_0.x5.x19.D I11 1.27f
C734 frontAnalog_v0p0p1_9.RSfetsym_0.QN I6 2.02f
C735 16to4_PriorityEncoder_v0p0p1_0.x5.A2 VDD 3.08f
C736 VDD I2 4.22f
C737 frontAnalog_v0p0p1_5.RSfetsym_0.x2.Y VDD 0.926f
C738 16to4_PriorityEncoder_v0p0p1_0.x5.x17.A I14 0.0474f
C739 frontAnalog_v0p0p1_8.RSfetsym_0.QN a_59577_n46683# 0.418f
C740 frontAnalog_v0p0p1_8.x65.A VDD 3.45f
C741 frontAnalog_v0p0p1_2.x65.X frontAnalog_v0p0p1_2.x63.X 0.136f
C742 w_55000_n68350# VV4 0.751f
C743 16to4_PriorityEncoder_v0p0p1_0.x3.x1.X VDD 0.393f
C744 frontAnalog_v0p0p1_6.RSfetsym_0.x2.Y I10 0.196f
C745 a_55268_n14736# VV14 0.215f
C746 16to4_PriorityEncoder_v0p0p1_0.x3.x21.B a_78097_n53777# 0.186f
C747 frontAnalog_v0p0p1_6.x63.X VDD 3.16f
C748 frontAnalog_v0p0p1_7.x65.X a_59578_n35370# 0.436f
C749 CLK I15 0.01f
C750 frontAnalog_v0p0p1_14.RSfetsym_0.QN I2 0.0512f
C751 frontAnalog_v0p0p1_2.RSfetsym_0.QN frontAnalog_v0p0p1_2.RSfetsym_0.x1.Y 0.17f
C752 w_55000_n83928# a_55268_n84936# 0.149f
C753 a_55268_n36336# VDD 0.565f
C754 w_55000_n19128# a_53630_n20196# 0.359f
C755 w_55000_n84550# a_53630_n84996# 0.394f
C756 16to4_PriorityEncoder_v0p0p1_0.x22.Y VDD 17f
C757 16to4_PriorityEncoder_v0p0p1_0.x3.x17.A I6 0.0474f
C758 frontAnalog_v0p0p1_12.x63.A a_57123_n74279# 0.212f
C759 frontAnalog_v0p0p1_13.RSfetsym_0.x1.Y I3 0.0436f
C760 w_55000_n57550# a_55268_n57936# 0.12f
C761 a_53630_n57996# a_55268_n57936# 0.015f
C762 frontAnalog_v0p0p1_15.RSfetsym_0.QN a_59578_n83970# 0.255f
C763 frontAnalog_v0p0p1_11.x65.X CLK 0.0398f
C764 frontAnalog_v0p0p1_7.x63.A VIN 0.187f
C765 a_55268_n14736# CLK 0.236f
C766 frontAnalog_v0p0p1_13.x65.A VDD 3.45f
C767 frontAnalog_v0p0p1_4.x63.A frontAnalog_v0p0p1_4.x65.A 3.16f
C768 w_55000_n29928# VV11 0.798f
C769 w_55000_n19750# frontAnalog_v0p0p1_4.x65.A 0.0988f
C770 16to4_PriorityEncoder_v0p0p1_0.x5.x16.C 16to4_PriorityEncoder_v0p0p1_0.x5.x15.X 0.0319f
C771 16to4_PriorityEncoder_v0p0p1_0.x3.EO VDD 0.761f
C772 frontAnalog_v0p0p1_13.x63.A frontAnalog_v0p0p1_13.x63.X 0.0301f
C773 w_55000_n46750# CLK 0.535f
C774 w_55000_n67728# frontAnalog_v0p0p1_10.IB 0.0216f
C775 16to4_PriorityEncoder_v0p0p1_0.x3.x19.D I6 0.464f
C776 16to4_PriorityEncoder_v0p0p1_0.x5.x16.X a_77605_n43545# 0.102f
C777 VV12 VV11 3.43f
C778 frontAnalog_v0p0p1_2.RSfetsym_0.x1.Y frontAnalog_v0p0p1_2.RSfetsym_0.x2.Y 0.0254f
C779 a_82906_n51645# 16to4_PriorityEncoder_v0p0p1_0.x2.X 0.12f
C780 frontAnalog_v0p0p1_1.x63.A a_57123_n41879# 0.212f
C781 16to4_PriorityEncoder_v0p0p1_0.x3.x19.C 16to4_PriorityEncoder_v0p0p1_0.x3.x21.B 0.0127f
C782 a_82906_n47995# VDD 0.179f
C783 a_77605_n40069# I12 0.208f
C784 a_59577_n14283# VDD 0.0173f
C785 a_57123_n40359# VDD 0.224f
C786 frontAnalog_v0p0p1_12.x65.A frontAnalog_v0p0p1_12.x65.X 0.0236f
C787 w_55000_n19128# VDD 0.854f
C788 a_55268_n20136# VIN 0.177f
C789 frontAnalog_v0p0p1_11.x63.X CLK 0.785f
C790 VDD VV7 4.76f
C791 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_7.x65.A 0.0352f
C792 frontAnalog_v0p0p1_7.x65.X frontAnalog_v0p0p1_7.RSfetsym_0.x1.Y 0.182f
C793 frontAnalog_v0p0p1_11.x63.A a_57123_n63479# 0.212f
C794 w_55000_n78528# VV2 0.798f
C795 frontAnalog_v0p0p1_0.x65.A CLK 2.61f
C796 a_55268_n30936# CLK 0.236f
C797 frontAnalog_v0p0p1_13.RSfetsym_0.QN I3 2.02f
C798 a_53630_n47196# a_55268_n47136# 0.015f
C799 a_77605_n51335# 16to4_PriorityEncoder_v0p0p1_0.x3.x16.X 0.0121f
C800 frontAnalog_v0p0p1_15.RSfetsym_0.QN frontAnalog_v0p0p1_15.RSfetsym_0.x1.Y 0.17f
C801 a_53630_n79596# VDD 0.134f
C802 16to4_PriorityEncoder_v0p0p1_0.x5.x16.C I11 0.132f
C803 16to4_PriorityEncoder_v0p0p1_0.x22.A VDD 1.52f
C804 VV16 VFS 4.16f
C805 16to4_PriorityEncoder_v0p0p1_0.x3.x17.A a_78065_n49349# 0.2f
C806 a_82906_n43855# VDD 0.181f
C807 a_59577_n30483# VDD 0.0173f
C808 w_55000_n29928# VIN 0.866f
C809 frontAnalog_v0p0p1_8.x65.A frontAnalog_v0p0p1_8.x65.X 0.0236f
C810 a_77605_n39305# VDD 0.149f
C811 w_55000_n67728# frontAnalog_v0p0p1_13.x65.A 0.658f
C812 16to4_PriorityEncoder_v0p0p1_0.x5.x19.C 16to4_PriorityEncoder_v0p0p1_0.x5.x21.B 0.0127f
C813 frontAnalog_v0p0p1_7.RSfetsym_0.x1.Y frontAnalog_v0p0p1_7.x63.X 0.883f
C814 16to4_PriorityEncoder_v0p0p1_0.x5.x22.A I14 0.0536f
C815 frontAnalog_v0p0p1_11.x65.A frontAnalog_v0p0p1_11.x65.X 0.0236f
C816 frontAnalog_v0p0p1_2.RSfetsym_0.QN frontAnalog_v0p0p1_2.RSfetsym_0.x2.Y 0.018f
C817 frontAnalog_v0p0p1_13.RSfetsym_0.x2.Y I3 0.198f
C818 frontAnalog_v0p0p1_7.x65.A a_55268_n36336# 0.461f
C819 a_77605_n53805# 16to4_PriorityEncoder_v0p0p1_0.x3.x20.X 0.0895f
C820 16to4_PriorityEncoder_v0p0p1_0.x29.Y OUT1 8.67f
C821 VDD VV1 2.06f
C822 VV14 VV13 4.07f
C823 frontAnalog_v0p0p1_3.x65.A a_55268_n14736# 0.461f
C824 frontAnalog_v0p0p1_2.x63.A a_55268_n3936# 1.24f
C825 frontAnalog_v0p0p1_2.x63.A CLK 1.8f
C826 CLK I8 0.01f
C827 VIN VV12 2.55f
C828 frontAnalog_v0p0p1_9.RSfetsym_0.x1.Y I6 0.0436f
C829 w_55000_n68350# frontAnalog_v0p0p1_13.x63.A 0.659f
C830 frontAnalog_v0p0p1_6.x63.A VDD 3.67f
C831 frontAnalog_v0p0p1_7.x65.X frontAnalog_v0p0p1_7.RSfetsym_0.QN 2.28f
C832 frontAnalog_v0p0p1_2.x63.X a_59577_n3483# 0.28f
C833 I12 I10 0.849f
C834 w_55000_n57550# VDD 0.829f
C835 16to4_PriorityEncoder_v0p0p1_0.x3.x22.A I6 0.0536f
C836 16to4_PriorityEncoder_v0p0p1_0.x3.x18.C 16to4_PriorityEncoder_v0p0p1_0.x3.x21.B 0.014f
C837 a_53630_n57996# VDD 0.134f
C838 w_55000_n13728# VV14 0.798f
C839 a_55268_n9336# VDD 0.565f
C840 16to4_PriorityEncoder_v0p0p1_0.x3.x19.D 16to4_PriorityEncoder_v0p0p1_0.x3.x4.A 0.0516f
C841 a_77605_n48109# I5 0.16f
C842 CLK VV13 6.01f
C843 frontAnalog_v0p0p1_15.x63.A VIN 0.188f
C844 16to4_PriorityEncoder_v0p0p1_0.x3.x16.C I6 0.491f
C845 frontAnalog_v0p0p1_7.x63.X a_57123_n36479# 0.121f
C846 frontAnalog_v0p0p1_7.x63.X m3_58396_n36750# 0.139f
C847 I13 I9 0.376f
C848 m3_58396_n31350# VDD 1.3f
C849 frontAnalog_v0p0p1_15.RSfetsym_0.QN a_59577_n84483# 0.418f
C850 a_77605_n51335# 16to4_PriorityEncoder_v0p0p1_0.x3.x15.X 0.0951f
C851 a_53630_n41796# CLK 0.0136f
C852 w_55000_n13728# CLK 0.571f
C853 a_53630_n47196# VDD 0.134f
C854 frontAnalog_v0p0p1_7.RSfetsym_0.QN frontAnalog_v0p0p1_7.x63.X 0.378f
C855 w_55000_n30550# frontAnalog_v0p0p1_10.IB 0.0217f
C856 frontAnalog_v0p0p1_7.x65.X frontAnalog_v0p0p1_7.RSfetsym_0.x2.Y 0.526f
C857 16to4_PriorityEncoder_v0p0p1_0.x3.x17.A 16to4_PriorityEncoder_v0p0p1_0.x3.x16.X 0.0198f
C858 a_82906_n51645# 16to4_PriorityEncoder_v0p0p1_0.x3.A0 0.119f
C859 frontAnalog_v0p0p1_9.x63.X m3_58396_n52950# 0.139f
C860 16to4_PriorityEncoder_v0p0p1_0.x21.A VDD 0.539f
C861 16to4_PriorityEncoder_v0p0p1_0.x3.x21.B I3 0.0112f
C862 w_55000_n52150# a_53630_n52596# 0.394f
C863 w_55000_n51528# a_55268_n52536# 0.149f
C864 I15 I11 1.03f
C865 16to4_PriorityEncoder_v0p0p1_0.x5.x16.C 16to4_PriorityEncoder_v0p0p1_0.x5.x19.D 1.24f
C866 a_77605_n43545# I11 0.162f
C867 w_55000_n68350# VIN 0.737f
C868 VV5 VV4 5.09f
C869 frontAnalog_v0p0p1_10.IB VV10 3.7f
C870 w_55000_n46750# VV8 0.751f
C871 16to4_PriorityEncoder_v0p0p1_0.x5.x18.C 16to4_PriorityEncoder_v0p0p1_0.x5.x21.B 0.014f
C872 a_77637_n42017# I14 0.186f
C873 16to4_PriorityEncoder_v0p0p1_0.x1.A 16to4_PriorityEncoder_v0p0p1_0.x2.A 0.304f
C874 frontAnalog_v0p0p1_8.RSfetsym_0.x1.Y frontAnalog_v0p0p1_8.RSfetsym_0.x2.Y 0.0254f
C875 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_15.x65.A 0.0352f
C876 16to4_PriorityEncoder_v0p0p1_0.x3.x19.X 16to4_PriorityEncoder_v0p0p1_0.x3.x20.X 0.145f
C877 I14 I12 2.36f
C878 a_77605_n52819# 16to4_PriorityEncoder_v0p0p1_0.x3.x19.X 0.0873f
C879 frontAnalog_v0p0p1_7.x63.X frontAnalog_v0p0p1_7.RSfetsym_0.x2.Y 0.0923f
C880 w_55000_n62328# w_55000_n62950# 0.327f
C881 frontAnalog_v0p0p1_2.x65.X I15 0.445f
C882 a_55268_n68736# VDD 0.565f
C883 frontAnalog_v0p0p1_4.x63.A a_55268_n20136# 1.24f
C884 frontAnalog_v0p0p1_10.IB a_53630_n52596# 0.473f
C885 w_55000_n35328# a_53630_n36396# 0.359f
C886 a_53630_n3996# VIN 0.265f
C887 frontAnalog_v0p0p1_7.x65.X VDD 3.55f
C888 w_55000_n19750# a_55268_n20136# 0.12f
C889 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_10.x63.A 0.0926f
C890 a_77605_n40069# VDD 0.156f
C891 16to4_PriorityEncoder_v0p0p1_0.x3.x22.A a_78065_n49349# 0.077f
C892 16to4_PriorityEncoder_v0p0p1_0.x3.x15.X 16to4_PriorityEncoder_v0p0p1_0.x3.x16.X 0.253f
C893 I0 S0 0.446f
C894 frontAnalog_v0p0p1_1.x63.A a_55268_n41736# 1.24f
C895 16to4_PriorityEncoder_v0p0p1_0.x5.x19.C I11 0.921f
C896 a_57123_n7959# frontAnalog_v0p0p1_0.x65.X 0.119f
C897 frontAnalog_v0p0p1_3.x65.X CLK 0.0393f
C898 a_55268_n36336# VV10 0.215f
C899 16to4_PriorityEncoder_v0p0p1_0.x3.x22.A a_77605_n51335# 0.0116f
C900 frontAnalog_v0p0p1_14.x63.A CLK 1.81f
C901 VIN VV6 2.58f
C902 frontAnalog_v0p0p1_4.x65.A VDD 3.45f
C903 16to4_PriorityEncoder_v0p0p1_0.x3.x16.C a_77605_n51335# 0.0949f
C904 w_55000_n52150# CLK 0.535f
C905 w_55000_n73128# frontAnalog_v0p0p1_10.IB 0.0216f
C906 16to4_PriorityEncoder_v0p0p1_0.x5.A2 16to4_PriorityEncoder_v0p0p1_0.x3.A2 0.358f
C907 frontAnalog_v0p0p1_2.x63.X I15 1.78f
C908 16to4_PriorityEncoder_v0p0p1_0.x3.x17.A 16to4_PriorityEncoder_v0p0p1_0.x3.x15.X 0.0789f
C909 frontAnalog_v0p0p1_10.IB VV14 3.7f
C910 frontAnalog_v0p0p1_7.x63.X VDD 3.16f
C911 16to4_PriorityEncoder_v0p0p1_0.x2.X VDD 0.351f
C912 w_55000_n24528# w_55000_n25150# 0.327f
C913 w_55000_n24528# VDD 0.854f
C914 w_55000_n13728# frontAnalog_v0p0p1_3.x65.A 0.658f
C915 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_12.x63.A 0.0926f
C916 frontAnalog_v0p0p1_5.x65.A a_55268_n25536# 0.461f
C917 w_55000_n56928# VV6 0.798f
C918 frontAnalog_v0p0p1_1.x63.X I9 0.015f
C919 frontAnalog_v0p0p1_0.x65.X a_59578_n8370# 0.436f
C920 frontAnalog_v0p0p1_3.x63.X CLK 0.785f
C921 frontAnalog_v0p0p1_7.RSfetsym_0.QN a_59577_n35883# 0.418f
C922 frontAnalog_v0p0p1_1.x63.A VIN 0.187f
C923 16to4_PriorityEncoder_v0p0p1_0.x5.x19.D I15 0.244f
C924 frontAnalog_v0p0p1_7.x63.A a_57123_n36479# 0.212f
C925 CLK I3 0.01f
C926 frontAnalog_v0p0p1_6.x65.X CLK 0.0402f
C927 frontAnalog_v0p0p1_3.x63.A a_57123_n14879# 0.212f
C928 frontAnalog_v0p0p1_10.IB a_55268_n3936# 0.0848f
C929 frontAnalog_v0p0p1_10.IB CLK 33.4f
C930 w_55000_n14350# frontAnalog_v0p0p1_3.x63.A 0.659f
C931 frontAnalog_v0p0p1_9.RSfetsym_0.QN frontAnalog_v0p0p1_9.RSfetsym_0.x1.Y 0.17f
C932 a_57123_n78159# VDD 0.224f
C933 a_59578_n8370# I14 0.42f
C934 w_55000_n67728# a_55268_n68736# 0.149f
C935 w_55000_n68350# a_53630_n68796# 0.394f
C936 16to4_PriorityEncoder_v0p0p1_0.x3.x19.C I6 0.304f
C937 16to4_PriorityEncoder_v0p0p1_0.x3.x22.A 16to4_PriorityEncoder_v0p0p1_0.x3.x16.X 0.0732f
C938 I11 I8 0.672f
C939 VDD I10 7.98f
C940 16to4_PriorityEncoder_v0p0p1_0.x43.Y OUT3 7.92f
C941 frontAnalog_v0p0p1_2.x65.A VV16 0.252f
C942 16to4_PriorityEncoder_v0p0p1_0.x3.A2 16to4_PriorityEncoder_v0p0p1_0.x3.EO 0.162f
C943 CLK I2 0.01f
C944 16to4_PriorityEncoder_v0p0p1_0.x3.x11.X a_78065_n49349# 0.202f
C945 frontAnalog_v0p0p1_9.x65.X a_59578_n51570# 0.436f
C946 frontAnalog_v0p0p1_2.x65.A a_57123_n2559# 0.214f
C947 a_57123_n79679# VDD 0.222f
C948 16to4_PriorityEncoder_v0p0p1_0.x3.x16.C 16to4_PriorityEncoder_v0p0p1_0.x3.x16.X 0.07f
C949 frontAnalog_v0p0p1_8.x65.A CLK 2.61f
C950 w_55000_n35328# VIN 0.866f
C951 a_78649_n39527# VDD 0.414f
C952 w_55000_n29928# frontAnalog_v0p0p1_6.x65.A 0.658f
C953 a_53630_n84996# VIN 0.265f
C954 a_59578_n24570# I11 0.42f
C955 16to4_PriorityEncoder_v0p0p1_0.x5.x18.C I11 0.251f
C956 a_53630_n52596# VV7 0.28f
C957 frontAnalog_v0p0p1_6.x63.X CLK 0.785f
C958 a_77637_n50057# I6 0.186f
C959 frontAnalog_v0p0p1_7.x65.A frontAnalog_v0p0p1_7.x65.X 0.0236f
C960 16to4_PriorityEncoder_v0p0p1_0.x5.x17.A a_78349_n43045# 0.213f
C961 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_1.x65.A 0.0352f
C962 16to4_PriorityEncoder_v0p0p1_0.x3.x19.X 16to4_PriorityEncoder_v0p0p1_0.x3.x21.X 0.131f
C963 a_78525_n53555# 16to4_PriorityEncoder_v0p0p1_0.x3.x20.X 0.0765f
C964 frontAnalog_v0p0p1_3.x65.A frontAnalog_v0p0p1_3.x65.X 0.0236f
C965 16to4_PriorityEncoder_v0p0p1_0.x3.x22.A 16to4_PriorityEncoder_v0p0p1_0.x3.x17.A 1.27f
C966 16to4_PriorityEncoder_v0p0p1_0.x5.x19.C 16to4_PriorityEncoder_v0p0p1_0.x5.x19.D 0.996f
C967 a_77637_n49127# 16to4_PriorityEncoder_v0p0p1_0.x3.x22.A 0.0288f
C968 frontAnalog_v0p0p1_11.x63.A VIN 0.187f
C969 frontAnalog_v0p0p1_12.x63.X m3_58396_n74550# 0.139f
C970 a_55268_n36336# CLK 0.236f
C971 w_55000_n30550# frontAnalog_v0p0p1_6.x63.A 0.659f
C972 frontAnalog_v0p0p1_0.x65.X frontAnalog_v0p0p1_0.RSfetsym_0.x1.Y 0.182f
C973 frontAnalog_v0p0p1_3.x63.A VIN 0.19f
C974 frontAnalog_v0p0p1_14.RSfetsym_0.x1.Y frontAnalog_v0p0p1_14.RSfetsym_0.x2.Y 0.0254f
C975 frontAnalog_v0p0p1_10.x65.A VIN 0.655f
C976 w_55000_n2928# frontAnalog_v0p0p1_2.x63.A 0.0792f
C977 w_55000_n62950# VDD 0.829f
C978 VDD S0 3.55f
C979 a_57123_n56559# VDD 0.224f
C980 16to4_PriorityEncoder_v0p0p1_0.x1.A 16to4_PriorityEncoder_v0p0p1_0.x3.A1 0.426f
C981 frontAnalog_v0p0p1_15.x65.A VV1 0.252f
C982 w_55000_n51528# frontAnalog_v0p0p1_9.x63.A 0.0792f
C983 frontAnalog_v0p0p1_13.x65.A CLK 2.61f
C984 frontAnalog_v0p0p1_0.x65.X VDD 3.55f
C985 frontAnalog_v0p0p1_0.RSfetsym_0.x1.Y I14 0.0432f
C986 a_55268_n52536# VIN 0.177f
C987 a_59577_n3483# I15 0.29f
C988 16to4_PriorityEncoder_v0p0p1_0.x3.x19.D 16to4_PriorityEncoder_v0p0p1_0.x3.x22.A 0.0292f
C989 a_59577_n35883# VDD 0.0173f
C990 a_77639_n50381# I7 0.192f
C991 m3_58396_n42150# VDD 1.3f
C992 w_55000_n56928# frontAnalog_v0p0p1_10.x65.A 0.658f
C993 VDD I14 7.95f
C994 frontAnalog_v0p0p1_2.x63.A frontAnalog_v0p0p1_2.x63.X 0.0301f
C995 a_82906_n43855# 16to4_PriorityEncoder_v0p0p1_0.x3.A2 0.119f
C996 frontAnalog_v0p0p1_14.RSfetsym_0.x2.Y VDD 0.926f
C997 a_57123_n67359# frontAnalog_v0p0p1_13.x65.X 0.119f
C998 16to4_PriorityEncoder_v0p0p1_0.x3.x16.C 16to4_PriorityEncoder_v0p0p1_0.x3.x19.D 1.24f
C999 16to4_PriorityEncoder_v0p0p1_0.x3.x2.X I6 0.0177f
C1000 frontAnalog_v0p0p1_0.RSfetsym_0.x1.Y frontAnalog_v0p0p1_0.x63.X 0.883f
C1001 VIN VV5 2.63f
C1002 w_55000_n19128# CLK 0.571f
C1003 frontAnalog_v0p0p1_5.RSfetsym_0.x1.Y I11 0.0436f
C1004 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_11.x65.A 0.0352f
C1005 a_57123_n45759# VDD 0.224f
C1006 w_55000_n35950# frontAnalog_v0p0p1_10.IB 0.0217f
C1007 16to4_PriorityEncoder_v0p0p1_0.x3.x18.C I6 0.3f
C1008 16to4_PriorityEncoder_v0p0p1_0.x3.x22.A 16to4_PriorityEncoder_v0p0p1_0.x3.x15.X 0.209f
C1009 a_53630_n20196# a_55268_n20136# 0.015f
C1010 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_3.x65.A 0.0352f
C1011 16to4_PriorityEncoder_v0p0p1_0.x5.x16.C I15 0.26f
C1012 16to4_PriorityEncoder_v0p0p1_0.x3.A0 VDD 0.829f
C1013 frontAnalog_v0p0p1_10.IB a_55268_n84936# 0.0848f
C1014 16to4_PriorityEncoder_v0p0p1_0.x5.x16.C a_77605_n43545# 0.0677f
C1015 frontAnalog_v0p0p1_12.x65.A VIN 0.655f
C1016 a_59578_n56970# VDD 0.0213f
C1017 w_55000_n57550# frontAnalog_v0p0p1_10.x63.A 0.659f
C1018 frontAnalog_v0p0p1_7.x63.A VDD 3.67f
C1019 CLK VV7 5.72f
C1020 w_55000_n73750# VIN 0.737f
C1021 a_77605_n47345# 16to4_PriorityEncoder_v0p0p1_0.x3.x2.X 0.0313f
C1022 frontAnalog_v0p0p1_0.x63.X VDD 3.16f
C1023 16to4_PriorityEncoder_v0p0p1_0.x5.x19.X a_78525_n45515# 0.193f
C1024 16to4_PriorityEncoder_v0p0p1_0.x3.x16.C 16to4_PriorityEncoder_v0p0p1_0.x3.x15.X 0.0319f
C1025 16to4_PriorityEncoder_v0p0p1_0.x5.x19.D I8 0.122f
C1026 16to4_PriorityEncoder_v0p0p1_0.x3.x19.C a_77605_n51335# 0.173f
C1027 frontAnalog_v0p0p1_1.RSfetsym_0.x1.Y frontAnalog_v0p0p1_1.x63.X 0.883f
C1028 frontAnalog_v0p0p1_0.x65.X frontAnalog_v0p0p1_0.RSfetsym_0.QN 2.28f
C1029 frontAnalog_v0p0p1_14.RSfetsym_0.QN frontAnalog_v0p0p1_14.RSfetsym_0.x2.Y 0.018f
C1030 frontAnalog_v0p0p1_4.x65.A a_57123_n18759# 0.214f
C1031 a_53630_n79596# CLK 0.0136f
C1032 w_55000_n78528# frontAnalog_v0p0p1_14.x63.A 0.0792f
C1033 16to4_PriorityEncoder_v0p0p1_0.x3.x11.X 16to4_PriorityEncoder_v0p0p1_0.x3.x17.A 0.125f
C1034 a_77637_n49127# 16to4_PriorityEncoder_v0p0p1_0.x3.x11.X 0.109f
C1035 16to4_PriorityEncoder_v0p0p1_0.x5.x18.C 16to4_PriorityEncoder_v0p0p1_0.x5.x19.D 0.491f
C1036 frontAnalog_v0p0p1_1.x65.A a_57123_n40359# 0.214f
C1037 frontAnalog_v0p0p1_13.x65.X a_59578_n67770# 0.436f
C1038 VV16 VV15 4.68f
C1039 frontAnalog_v0p0p1_0.RSfetsym_0.QN I14 2.02f
C1040 frontAnalog_v0p0p1_0.x63.X a_57123_n9479# 0.121f
C1041 a_77637_n40777# 16to4_PriorityEncoder_v0p0p1_0.x5.x14.A 0.135f
C1042 VIN VV16 2.34f
C1043 I6 I3 0.602f
C1044 frontAnalog_v0p0p1_13.x65.X VDD 3.55f
C1045 w_55000_n35950# a_55268_n36336# 0.12f
C1046 I7 I1 0.244f
C1047 a_55268_n20136# VDD 0.565f
C1048 16to4_PriorityEncoder_v0p0p1_0.x3.A1 a_78349_n51085# 0.151f
C1049 16to4_PriorityEncoder_v0p0p1_0.x5.x22.A a_78525_n45515# 0.209f
C1050 a_57123_n56559# frontAnalog_v0p0p1_10.x65.X 0.119f
C1051 frontAnalog_v0p0p1_10.IB a_53630_n74196# 0.473f
C1052 16to4_PriorityEncoder_v0p0p1_0.x5.x19.C 16to4_PriorityEncoder_v0p0p1_0.x5.x16.C 1.95f
C1053 frontAnalog_v0p0p1_5.x63.A a_57123_n25679# 0.212f
C1054 frontAnalog_v0p0p1_10.IB VV8 3.7f
C1055 frontAnalog_v0p0p1_1.RSfetsym_0.x2.Y I9 0.0165f
C1056 a_77605_n47345# I3 0.0597f
C1057 frontAnalog_v0p0p1_0.x65.X frontAnalog_v0p0p1_0.RSfetsym_0.x2.Y 0.526f
C1058 frontAnalog_v0p0p1_0.RSfetsym_0.QN frontAnalog_v0p0p1_0.x63.X 0.378f
C1059 CLK VV1 5.44f
C1060 frontAnalog_v0p0p1_5.RSfetsym_0.QN I11 2.02f
C1061 I5 I0 0.344f
C1062 I2 I6 0.441f
C1063 frontAnalog_v0p0p1_12.RSfetsym_0.QN a_59578_n73170# 0.255f
C1064 16to4_PriorityEncoder_v0p0p1_0.x5.x22.A a_78349_n43045# 0.17f
C1065 a_78525_n53555# 16to4_PriorityEncoder_v0p0p1_0.x3.x21.X 0.202f
C1066 frontAnalog_v0p0p1_10.RSfetsym_0.x1.Y VDD 0.733f
C1067 frontAnalog_v0p0p1_6.x63.A CLK 1.81f
C1068 frontAnalog_v0p0p1_0.RSfetsym_0.x2.Y I14 0.195f
C1069 w_55000_n57550# CLK 0.535f
C1070 16to4_PriorityEncoder_v0p0p1_0.x3.EI I5 3.69f
C1071 w_55000_n78528# frontAnalog_v0p0p1_10.IB 0.0216f
C1072 frontAnalog_v0p0p1_8.x65.A VV8 0.253f
C1073 a_53630_n57996# CLK 0.0136f
C1074 frontAnalog_v0p0p1_13.x63.X VDD 3.16f
C1075 a_77605_n47345# I2 0.216f
C1076 frontAnalog_v0p0p1_4.x63.A frontAnalog_v0p0p1_4.x63.X 0.0301f
C1077 a_55268_n9336# CLK 0.236f
C1078 I4 I5 6.86f
C1079 frontAnalog_v0p0p1_4.x65.X I12 0.446f
C1080 w_55000_n41350# a_53630_n41796# 0.394f
C1081 w_55000_n40728# a_55268_n41736# 0.149f
C1082 w_55000_n29928# VDD 0.854f
C1083 frontAnalog_v0p0p1_10.x65.X a_59578_n56970# 0.436f
C1084 16to4_PriorityEncoder_v0p0p1_0.x2.A 16to4_PriorityEncoder_v0p0p1_0.x3.A1 1.21f
C1085 m3_58396_n69150# I3 0.0416f
C1086 16to4_PriorityEncoder_v0p0p1_0.x3.x4.A 16to4_PriorityEncoder_v0p0p1_0.x3.x2.X 0.125f
C1087 a_77605_n47345# 16to4_PriorityEncoder_v0p0p1_0.x3.x1.X 0.0991f
C1088 16to4_PriorityEncoder_v0p0p1_0.x5.x2.X I12 0.0262f
C1089 frontAnalog_v0p0p1_13.x65.X frontAnalog_v0p0p1_13.RSfetsym_0.x1.Y 0.182f
C1090 frontAnalog_v0p0p1_5.x65.A frontAnalog_v0p0p1_5.x65.X 0.0236f
C1091 frontAnalog_v0p0p1_0.x63.X frontAnalog_v0p0p1_0.RSfetsym_0.x2.Y 0.0923f
C1092 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_5.x63.A 0.0926f
C1093 frontAnalog_v0p0p1_5.RSfetsym_0.x2.Y I11 0.198f
C1094 a_77605_n45765# VDD 0.552f
C1095 a_55268_n57936# VV6 0.215f
C1096 a_78159_n39549# 16to4_PriorityEncoder_v0p0p1_0.x5.x2.X 0.121f
C1097 a_77605_n52567# VDD 0.432f
C1098 frontAnalog_v0p0p1_8.x63.X I7 1.85f
C1099 frontAnalog_v0p0p1_12.x65.X frontAnalog_v0p0p1_12.x63.X 0.136f
C1100 16to4_PriorityEncoder_v0p0p1_0.x3.x16.X a_77605_n51585# 0.102f
C1101 w_55000_n25150# VV12 0.751f
C1102 VDD VV12 4.13f
C1103 a_57123_n58079# VDD 0.222f
C1104 frontAnalog_v0p0p1_7.x63.A frontAnalog_v0p0p1_7.x65.A 3.16f
C1105 a_57123_n45759# frontAnalog_v0p0p1_8.x65.X 0.119f
C1106 a_53630_n47196# CLK 0.0136f
C1107 a_59577_n8883# VDD 0.0173f
C1108 frontAnalog_v0p0p1_9.x63.A frontAnalog_v0p0p1_9.x63.X 0.0301f
C1109 a_53630_n63396# VIN 0.265f
C1110 16to4_PriorityEncoder_v0p0p1_0.x5.x16.C I8 0.12f
C1111 w_55000_n8328# frontAnalog_v0p0p1_0.x65.A 0.658f
C1112 frontAnalog_v0p0p1_11.RSfetsym_0.QN a_59578_n62370# 0.255f
C1113 frontAnalog_v0p0p1_4.x63.X I12 1.85f
C1114 w_55000_n2928# frontAnalog_v0p0p1_10.IB 0.0216f
C1115 frontAnalog_v0p0p1_12.RSfetsym_0.QN frontAnalog_v0p0p1_12.RSfetsym_0.x1.Y 0.17f
C1116 a_59578_n13770# I13 0.42f
C1117 16to4_PriorityEncoder_v0p0p1_0.x3.x17.A a_77637_n50057# 0.14f
C1118 frontAnalog_v0p0p1_10.RSfetsym_0.QN VDD 2.56f
C1119 m3_58396_n15150# I13 0.0416f
C1120 frontAnalog_v0p0p1_15.x63.A VDD 3.67f
C1121 frontAnalog_v0p0p1_13.RSfetsym_0.x1.Y frontAnalog_v0p0p1_13.x63.X 0.883f
C1122 w_55000_n40728# VIN 0.866f
C1123 16to4_PriorityEncoder_v0p0p1_0.x3.x19.C 16to4_PriorityEncoder_v0p0p1_0.x3.x19.D 0.996f
C1124 w_55000_n8950# frontAnalog_v0p0p1_0.x63.A 0.659f
C1125 16to4_PriorityEncoder_v0p0p1_0.x3.x4.A I3 0.0406f
C1126 frontAnalog_v0p0p1_9.x63.A VIN 0.187f
C1127 w_55000_n3550# frontAnalog_v0p0p1_2.x65.A 0.0988f
C1128 16to4_PriorityEncoder_v0p0p1_0.x5.x19.C I15 0.239f
C1129 16to4_PriorityEncoder_v0p0p1_0.x5.x19.C a_77605_n43545# 0.176f
C1130 16to4_PriorityEncoder_v0p0p1_0.x22.Y OUT0 8.68f
C1131 frontAnalog_v0p0p1_9.x65.X frontAnalog_v0p0p1_9.x63.X 0.136f
C1132 frontAnalog_v0p0p1_10.x65.X frontAnalog_v0p0p1_10.RSfetsym_0.x1.Y 0.182f
C1133 16to4_PriorityEncoder_v0p0p1_0.x43.Y VDD 11.4f
C1134 16to4_PriorityEncoder_v0p0p1_0.x3.x11.X 16to4_PriorityEncoder_v0p0p1_0.x3.x22.A 0.0936f
C1135 a_55268_n84936# VV1 0.214f
C1136 VV8 VV7 3.46f
C1137 w_55000_n52150# frontAnalog_v0p0p1_9.x65.A 0.0988f
C1138 a_55268_n68736# CLK 0.236f
C1139 a_77605_n43295# I10 0.167f
C1140 frontAnalog_v0p0p1_7.x65.X CLK 0.0389f
C1141 frontAnalog_v0p0p1_13.x65.X frontAnalog_v0p0p1_13.RSfetsym_0.QN 2.28f
C1142 frontAnalog_v0p0p1_0.RSfetsym_0.QN a_59577_n8883# 0.418f
C1143 frontAnalog_v0p0p1_8.RSfetsym_0.QN VDD 2.56f
C1144 a_77605_n51335# I2 0.167f
C1145 16to4_PriorityEncoder_v0p0p1_0.x3.x4.A I2 0.0109f
C1146 frontAnalog_v0p0p1_11.x65.X frontAnalog_v0p0p1_11.x63.X 0.136f
C1147 w_55000_n68350# VDD 0.829f
C1148 frontAnalog_v0p0p1_12.RSfetsym_0.x1.Y frontAnalog_v0p0p1_12.RSfetsym_0.x2.Y 0.0254f
C1149 frontAnalog_v0p0p1_10.RSfetsym_0.x2.Y VDD 0.926f
C1150 16to4_PriorityEncoder_v0p0p1_0.x3.x4.A 16to4_PriorityEncoder_v0p0p1_0.x3.x1.X 0.118f
C1151 frontAnalog_v0p0p1_13.x63.X a_57123_n68879# 0.121f
C1152 frontAnalog_v0p0p1_1.x63.X a_57123_n41879# 0.121f
C1153 frontAnalog_v0p0p1_1.RSfetsym_0.x1.Y frontAnalog_v0p0p1_1.RSfetsym_0.x2.Y 0.0254f
C1154 frontAnalog_v0p0p1_4.x65.A CLK 2.61f
C1155 VDD I5 5.32f
C1156 a_59578_n40770# I8 0.42f
C1157 frontAnalog_v0p0p1_10.IB a_55268_n63336# 0.0848f
C1158 a_59577_n68283# VDD 0.0173f
C1159 frontAnalog_v0p0p1_11.RSfetsym_0.QN frontAnalog_v0p0p1_11.RSfetsym_0.x1.Y 0.17f
C1160 a_78159_n39549# 16to4_PriorityEncoder_v0p0p1_0.x5.x1.X 0.192f
C1161 w_55000_n62328# frontAnalog_v0p0p1_11.x63.A 0.0792f
C1162 16to4_PriorityEncoder_v0p0p1_0.x5.x17.A 16to4_PriorityEncoder_v0p0p1_0.x1.A 0.115f
C1163 a_55268_n74136# VIN 0.177f
C1164 frontAnalog_v0p0p1_1.x63.A VV9 0.587f
C1165 m3_58396_n52950# VDD 1.3f
C1166 16to4_PriorityEncoder_v0p0p1_0.x5.x4.A a_77605_n39305# 0.0112f
C1167 frontAnalog_v0p0p1_10.RSfetsym_0.x1.Y frontAnalog_v0p0p1_10.x63.X 0.883f
C1168 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_9.x65.A 0.0352f
C1169 frontAnalog_v0p0p1_3.RSfetsym_0.x1.Y I13 0.0436f
C1170 w_55000_n78528# a_53630_n79596# 0.359f
C1171 frontAnalog_v0p0p1_15.x65.A S0 0.0236f
C1172 VDD OUT1 6.71f
C1173 frontAnalog_v0p0p1_10.x65.A a_55268_n57936# 0.461f
C1174 frontAnalog_v0p0p1_13.RSfetsym_0.QN frontAnalog_v0p0p1_13.x63.X 0.378f
C1175 frontAnalog_v0p0p1_7.x63.X CLK 0.785f
C1176 frontAnalog_v0p0p1_13.x65.X frontAnalog_v0p0p1_13.RSfetsym_0.x2.Y 0.526f
C1177 16to4_PriorityEncoder_v0p0p1_0.x3.x16.X I3 0.0148f
C1178 w_55000_n24528# CLK 0.571f
C1179 a_53630_n3996# VDD 0.134f
C1180 w_55000_n41350# frontAnalog_v0p0p1_10.IB 0.0217f
C1181 a_59577_n46683# I7 0.29f
C1182 I15 I8 0.342f
C1183 frontAnalog_v0p0p1_5.x65.A VIN 0.655f
C1184 w_55000_n79150# frontAnalog_v0p0p1_14.x65.A 0.0988f
C1185 frontAnalog_v0p0p1_10.x65.X frontAnalog_v0p0p1_10.RSfetsym_0.QN 2.28f
C1186 w_55000_n79150# VIN 0.737f
C1187 16to4_PriorityEncoder_v0p0p1_0.x3.x4.A 16to4_PriorityEncoder_v0p0p1_0.x3.EO 0.0491f
C1188 16to4_PriorityEncoder_v0p0p1_0.x3.x19.D 16to4_PriorityEncoder_v0p0p1_0.x3.x2.X 0.014f
C1189 a_77605_n39305# I11 0.0597f
C1190 frontAnalog_v0p0p1_14.x63.A VV2 0.587f
C1191 16to4_PriorityEncoder_v0p0p1_0.x3.x18.C 16to4_PriorityEncoder_v0p0p1_0.x3.x19.D 0.491f
C1192 VDD VV6 4.67f
C1193 frontAnalog_v0p0p1_11.RSfetsym_0.x1.Y frontAnalog_v0p0p1_11.RSfetsym_0.x2.Y 0.0254f
C1194 a_78159_n39549# 16to4_PriorityEncoder_v0p0p1_0.x5.EO 0.128f
C1195 a_59577_n19683# I12 0.29f
C1196 frontAnalog_v0p0p1_7.x63.A VV10 0.587f
C1197 16to4_PriorityEncoder_v0p0p1_0.x5.x18.C I15 0.229f
C1198 frontAnalog_v0p0p1_12.RSfetsym_0.QN frontAnalog_v0p0p1_12.RSfetsym_0.x2.Y 0.018f
C1199 frontAnalog_v0p0p1_10.x63.X a_57123_n58079# 0.121f
C1200 w_55000_n62328# VV5 0.798f
C1201 a_78649_n47567# 16to4_PriorityEncoder_v0p0p1_0.x3.GS 0.136f
C1202 frontAnalog_v0p0p1_13.x63.X frontAnalog_v0p0p1_13.RSfetsym_0.x2.Y 0.0923f
C1203 16to4_PriorityEncoder_v0p0p1_0.x43.A VDD 1.46f
C1204 frontAnalog_v0p0p1_1.x63.X frontAnalog_v0p0p1_1.RSfetsym_0.x2.Y 0.0923f
C1205 CLK I10 0.0103f
C1206 16to4_PriorityEncoder_v0p0p1_0.x3.x19.C 16to4_PriorityEncoder_v0p0p1_0.x3.x16.C 1.95f
C1207 frontAnalog_v0p0p1_8.x63.X a_59577_n46683# 0.28f
C1208 w_55000_n67728# w_55000_n68350# 0.327f
C1209 w_55000_n46128# frontAnalog_v0p0p1_8.x63.A 0.0792f
C1210 frontAnalog_v0p0p1_12.x63.X a_59577_n73683# 0.28f
C1211 frontAnalog_v0p0p1_4.x65.X VDD 3.55f
C1212 a_77605_n44527# VDD 0.439f
C1213 frontAnalog_v0p0p1_10.x65.X frontAnalog_v0p0p1_10.RSfetsym_0.x2.Y 0.526f
C1214 frontAnalog_v0p0p1_10.RSfetsym_0.QN frontAnalog_v0p0p1_10.x63.X 0.378f
C1215 frontAnalog_v0p0p1_3.RSfetsym_0.QN I13 2.02f
C1216 a_53630_n47196# VV8 0.28f
C1217 frontAnalog_v0p0p1_1.x63.A VDD 3.67f
C1218 16to4_PriorityEncoder_v0p0p1_0.x5.x19.C I8 0.12f
C1219 frontAnalog_v0p0p1_10.IB a_53630_n25596# 0.473f
C1220 16to4_PriorityEncoder_v0p0p1_0.x5.x2.X VDD 0.367f
C1221 w_55000_n3550# VIN 0.735f
C1222 16to4_PriorityEncoder_v0p0p1_0.x3.x19.D I3 1.27f
C1223 frontAnalog_v0p0p1_10.x65.X I5 0.446f
C1224 a_77637_n41087# I13 0.194f
C1225 frontAnalog_v0p0p1_10.IB VV2 3.69f
C1226 frontAnalog_v0p0p1_8.x65.X frontAnalog_v0p0p1_8.RSfetsym_0.QN 2.28f
C1227 16to4_PriorityEncoder_v0p0p1_0.x3.x16.C a_77605_n51585# 0.0677f
C1228 w_55000_n13728# a_55268_n14736# 0.149f
C1229 w_55000_n14350# a_53630_n14796# 0.394f
C1230 16to4_PriorityEncoder_v0p0p1_0.x1.A 16to4_PriorityEncoder_v0p0p1_0.x28.A 0.0126f
C1231 16to4_PriorityEncoder_v0p0p1_0.x5.EO 16to4_PriorityEncoder_v0p0p1_0.x3.EI 0.644f
C1232 16to4_PriorityEncoder_v0p0p1_0.x5.x18.C 16to4_PriorityEncoder_v0p0p1_0.x5.x19.C 2.6f
C1233 w_55000_n62950# CLK 0.535f
C1234 w_55000_n83928# frontAnalog_v0p0p1_10.IB 0.0216f
C1235 CLK S0 0.0406f
C1236 frontAnalog_v0p0p1_11.RSfetsym_0.QN frontAnalog_v0p0p1_11.RSfetsym_0.x2.Y 0.018f
C1237 a_77605_n44779# 16to4_PriorityEncoder_v0p0p1_0.x5.x19.X 0.0873f
C1238 16to4_PriorityEncoder_v0p0p1_0.x3.x19.D I2 0.196f
C1239 frontAnalog_v0p0p1_0.x65.X CLK 0.0389f
C1240 frontAnalog_v0p0p1_4.x63.X VDD 3.16f
C1241 frontAnalog_v0p0p1_9.x65.A VV7 0.252f
C1242 w_55000_n29928# w_55000_n30550# 0.327f
C1243 frontAnalog_v0p0p1_10.x63.X frontAnalog_v0p0p1_10.RSfetsym_0.x2.Y 0.0923f
C1244 w_55000_n35328# VDD 0.854f
C1245 frontAnalog_v0p0p1_3.RSfetsym_0.x2.Y I13 0.196f
C1246 a_53630_n84996# VDD 0.134f
C1247 frontAnalog_v0p0p1_13.RSfetsym_0.QN a_59577_n68283# 0.418f
C1248 a_53630_n30996# VV11 0.28f
C1249 m3_58396_n63750# I4 0.0416f
C1250 frontAnalog_v0p0p1_10.x63.X I5 1.85f
C1251 a_78525_n45515# VDD 0.165f
C1252 frontAnalog_v0p0p1_11.x63.X a_59577_n62883# 0.28f
C1253 CLK I14 0.01f
C1254 S0 R0 0.136f
C1255 16to4_PriorityEncoder_v0p0p1_0.x5.x22.A 16to4_PriorityEncoder_v0p0p1_0.x1.A 0.492f
C1256 a_59578_n73170# I2 0.42f
C1257 frontAnalog_v0p0p1_11.x63.A VDD 3.67f
C1258 frontAnalog_v0p0p1_3.x63.A VDD 3.67f
C1259 16to4_PriorityEncoder_v0p0p1_0.x42.A VDD 0.536f
C1260 frontAnalog_v0p0p1_10.x65.A VDD 3.45f
C1261 16to4_PriorityEncoder_v0p0p1_0.x3.EI 16to4_PriorityEncoder_v0p0p1_0.x3.x20.X 0.208f
C1262 a_78349_n43045# VDD 0.164f
C1263 a_53630_n14796# VIN 0.265f
C1264 a_77637_n48817# 16to4_PriorityEncoder_v0p0p1_0.x3.x14.A 0.135f
C1265 a_77605_n52567# 16to4_PriorityEncoder_v0p0p1_0.x3.x21.B 0.116f
C1266 frontAnalog_v0p0p1_7.x63.A CLK 1.81f
C1267 16to4_PriorityEncoder_v0p0p1_0.x3.EI a_77605_n52819# 0.175f
C1268 frontAnalog_v0p0p1_0.x63.X CLK 0.785f
C1269 w_55000_n8328# frontAnalog_v0p0p1_10.IB 0.0216f
C1270 a_78649_n47567# 16to4_PriorityEncoder_v0p0p1_0.x3.EO 0.135f
C1271 frontAnalog_v0p0p1_8.x63.A frontAnalog_v0p0p1_8.x63.X 0.0301f
C1272 a_55268_n52536# VDD 0.565f
C1273 w_55000_n46128# VIN 0.866f
C1274 I1 R1 1.9f
C1275 16to4_PriorityEncoder_v0p0p1_0.x5.x1.X VDD 0.39f
C1276 16to4_PriorityEncoder_v0p0p1_0.x5.x18.C I8 0.119f
C1277 a_77605_n48109# I7 0.0614f
C1278 frontAnalog_v0p0p1_12.x65.A VV3 0.253f
C1279 w_55000_n62328# a_53630_n63396# 0.359f
C1280 w_55000_n73750# VV3 0.751f
C1281 frontAnalog_v0p0p1_10.RSfetsym_0.QN a_59577_n57483# 0.418f
C1282 16to4_PriorityEncoder_v0p0p1_0.x3.x19.X a_78525_n53555# 0.193f
C1283 frontAnalog_v0p0p1_10.x63.A a_57123_n58079# 0.212f
C1284 VDD VV5 4.19f
C1285 frontAnalog_v0p0p1_13.x65.X CLK 0.0407f
C1286 16to4_PriorityEncoder_v0p0p1_0.x5.x14.A a_78065_n41309# 0.197f
C1287 16to4_PriorityEncoder_v0p0p1_0.x1.A 16to4_PriorityEncoder_v0p0p1_0.x1.X 0.0412f
C1288 a_55268_n20136# CLK 0.236f
C1289 frontAnalog_v0p0p1_15.x63.A frontAnalog_v0p0p1_15.x65.A 3.16f
C1290 16to4_PriorityEncoder_v0p0p1_0.x3.x16.C I3 0.132f
C1291 frontAnalog_v0p0p1_12.x65.A VDD 3.45f
C1292 a_59578_n35370# I9 0.42f
C1293 w_55000_n62950# frontAnalog_v0p0p1_11.x65.A 0.0988f
C1294 frontAnalog_v0p0p1_1.x65.X I9 0.0396f
C1295 a_53630_n30996# VIN 0.265f
C1296 w_55000_n73750# VDD 0.829f
C1297 frontAnalog_v0p0p1_12.RSfetsym_0.x1.Y I2 0.0436f
C1298 16to4_PriorityEncoder_v0p0p1_0.x5.EO VDD 1.06f
C1299 16to4_PriorityEncoder_v0p0p1_0.x5.x4.A I10 0.0109f
C1300 a_53630_n79596# VV2 0.28f
C1301 frontAnalog_v0p0p1_0.x63.A VV15 0.587f
C1302 16to4_PriorityEncoder_v0p0p1_0.x5.x22.A I13 0.066f
C1303 16to4_PriorityEncoder_v0p0p1_0.x3.x16.C I2 0.925f
C1304 w_55000_n24528# frontAnalog_v0p0p1_5.x63.A 0.0792f
C1305 frontAnalog_v0p0p1_10.IB a_55268_n14736# 0.0848f
C1306 frontAnalog_v0p0p1_0.x63.A VIN 0.19f
C1307 a_59577_n19683# VDD 0.0173f
C1308 m3_58396_n63750# VDD 1.3f
C1309 w_55000_n35328# frontAnalog_v0p0p1_7.x65.A 0.658f
C1310 a_55268_n25536# VIN 0.177f
C1311 w_55000_n79150# a_55268_n79536# 0.12f
C1312 frontAnalog_v0p0p1_13.x63.X CLK 0.785f
C1313 16to4_PriorityEncoder_v0p0p1_0.x5.x19.X 16to4_PriorityEncoder_v0p0p1_0.x2.A 0.0122f
C1314 VDD VV16 4.5f
C1315 frontAnalog_v0p0p1_10.x65.A frontAnalog_v0p0p1_10.x65.X 0.0236f
C1316 a_59577_n41283# I8 0.29f
C1317 a_59577_n57483# I5 0.29f
C1318 w_55000_n29928# CLK 0.571f
C1319 a_57123_n2559# VDD 0.224f
C1320 w_55000_n46750# frontAnalog_v0p0p1_10.IB 0.0217f
C1321 a_57123_n18759# frontAnalog_v0p0p1_4.x65.X 0.119f
C1322 frontAnalog_v0p0p1_12.RSfetsym_0.QN I3 0.0512f
C1323 I12 I9 0.43f
C1324 I11 I10 7.54f
C1325 w_55000_n35950# frontAnalog_v0p0p1_7.x63.A 0.659f
C1326 w_55000_n84550# VIN 0.737f
C1327 16to4_PriorityEncoder_v0p0p1_0.x3.x19.C a_77605_n51585# 0.176f
C1328 VV2 VV1 4.46f
C1329 frontAnalog_v0p0p1_9.x63.A a_57123_n52679# 0.212f
C1330 16to4_PriorityEncoder_v0p0p1_0.x5.GS VDD 0.771f
C1331 CLK VV12 6.38f
C1332 16to4_PriorityEncoder_v0p0p1_0.x3.x20.X VDD 0.242f
C1333 frontAnalog_v0p0p1_7.RSfetsym_0.x1.Y I9 0.0433f
C1334 w_55000_n40728# VV9 0.798f
C1335 a_77605_n52819# VDD 0.435f
C1336 w_55000_n46750# frontAnalog_v0p0p1_8.x65.A 0.0988f
C1337 w_55000_n83928# VV1 0.798f
C1338 16to4_PriorityEncoder_v0p0p1_0.x5.x22.A 16to4_PriorityEncoder_v0p0p1_0.x2.A 0.132f
C1339 frontAnalog_v0p0p1_12.RSfetsym_0.QN I2 2.02f
C1340 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_0.x65.A 0.0352f
C1341 frontAnalog_v0p0p1_10.IB a_55268_n30936# 0.0848f
C1342 a_59578_n2970# VDD 0.0213f
C1343 frontAnalog_v0p0p1_4.x65.X a_59578_n19170# 0.436f
C1344 frontAnalog_v0p0p1_15.x63.A CLK 1.81f
C1345 a_77605_n45765# 16to4_PriorityEncoder_v0p0p1_0.x5.x20.X 0.0895f
C1346 a_59578_n83970# S0 0.436f
C1347 w_55000_n8950# VV15 0.751f
C1348 16to4_PriorityEncoder_v0p0p1_0.x5.x14.A 16to4_PriorityEncoder_v0p0p1_0.x5.x17.A 0.105f
C1349 16to4_PriorityEncoder_v0p0p1_0.x3.EI 16to4_PriorityEncoder_v0p0p1_0.x1.A 0.534f
C1350 frontAnalog_v0p0p1_15.RSfetsym_0.x2.Y I0 0.198f
C1351 w_55000_n8950# VIN 0.737f
C1352 16to4_PriorityEncoder_v0p0p1_0.x3.x18.C 16to4_PriorityEncoder_v0p0p1_0.x3.x19.C 2.6f
C1353 16to4_PriorityEncoder_v0p0p1_0.x5.x11.X I13 0.0201f
C1354 a_77637_n40777# I12 0.188f
C1355 frontAnalog_v0p0p1_10.x63.A VV6 0.587f
C1356 m3_58396_n36750# I9 0.0416f
C1357 frontAnalog_v0p0p1_12.RSfetsym_0.x2.Y I2 0.198f
C1358 a_53630_n63396# VDD 0.134f
C1359 frontAnalog_v0p0p1_13.x63.A VV4 0.587f
C1360 I13 I12 7.14f
C1361 I14 I11 0.782f
C1362 frontAnalog_v0p0p1_15.x63.A R0 0.0301f
C1363 frontAnalog_v0p0p1_5.RSfetsym_0.QN a_59578_n24570# 0.255f
C1364 w_55000_n68350# CLK 0.535f
C1365 16to4_PriorityEncoder_v0p0p1_0.x2.A a_82906_n51645# 0.207f
C1366 frontAnalog_v0p0p1_2.x63.A frontAnalog_v0p0p1_10.IB 0.0784f
C1367 m3_58396_n58350# I5 0.0416f
C1368 frontAnalog_v0p0p1_7.RSfetsym_0.QN I9 2.02f
C1369 frontAnalog_v0p0p1_1.x65.X frontAnalog_v0p0p1_1.RSfetsym_0.x1.Y 0.182f
C1370 CLK I5 0.01f
C1371 w_55000_n40728# VDD 0.854f
C1372 a_57123_n83559# VDD 0.224f
C1373 w_55000_n8950# a_53630_n9396# 0.394f
C1374 frontAnalog_v0p0p1_9.x63.A VDD 3.67f
C1375 w_55000_n8328# a_55268_n9336# 0.149f
C1376 16to4_PriorityEncoder_v0p0p1_0.x5.x19.D I10 0.196f
C1377 frontAnalog_v0p0p1_2.RSfetsym_0.x1.Y VDD 0.733f
C1378 16to4_PriorityEncoder_v0p0p1_0.x3.x19.C I3 0.921f
C1379 16to4_PriorityEncoder_v0p0p1_0.x3.EI 16to4_PriorityEncoder_v0p0p1_0.x3.x14.A 0.0111f
C1380 frontAnalog_v0p0p1_4.x65.X frontAnalog_v0p0p1_4.RSfetsym_0.x1.Y 0.182f
C1381 frontAnalog_v0p0p1_10.IB VV13 3.7f
C1382 w_55000_n35328# VV10 0.798f
C1383 frontAnalog_v0p0p1_9.x65.X frontAnalog_v0p0p1_9.RSfetsym_0.x2.Y 0.526f
C1384 a_53630_n3996# CLK 0.0136f
C1385 a_53630_n3996# a_55268_n3936# 0.015f
C1386 16to4_PriorityEncoder_v0p0p1_0.x3.x14.A I4 0.0493f
C1387 a_57123_n85079# VDD 0.222f
C1388 frontAnalog_v0p0p1_15.RSfetsym_0.x1.Y S0 0.182f
C1389 frontAnalog_v0p0p1_5.x65.X frontAnalog_v0p0p1_5.x63.X 0.136f
C1390 VIN VV4 2.6f
C1391 frontAnalog_v0p0p1_7.RSfetsym_0.x2.Y I9 0.192f
C1392 a_55268_n74136# VV3 0.215f
C1393 frontAnalog_v0p0p1_10.IB a_53630_n41796# 0.473f
C1394 16to4_PriorityEncoder_v0p0p1_0.x3.x19.C I2 0.447f
C1395 w_55000_n13728# frontAnalog_v0p0p1_10.IB 0.0216f
C1396 frontAnalog_v0p0p1_3.RSfetsym_0.QN a_59578_n13770# 0.255f
C1397 CLK VV6 6.01f
C1398 a_77605_n51585# I3 0.162f
C1399 frontAnalog_v0p0p1_9.x65.X VDD 3.55f
C1400 frontAnalog_v0p0p1_5.RSfetsym_0.QN frontAnalog_v0p0p1_5.RSfetsym_0.x1.Y 0.17f
C1401 w_55000_n51528# VIN 0.866f
C1402 frontAnalog_v0p0p1_15.x63.A a_55268_n84936# 1.24f
C1403 a_57123_n4079# VDD 0.222f
C1404 16to4_PriorityEncoder_v0p0p1_0.x3.x21.X VDD 0.501f
C1405 a_55268_n74136# VDD 0.565f
C1406 frontAnalog_v0p0p1_4.RSfetsym_0.x1.Y frontAnalog_v0p0p1_4.x63.X 0.883f
C1407 frontAnalog_v0p0p1_1.x65.X frontAnalog_v0p0p1_1.x63.X 0.136f
C1408 w_55000_n24528# a_53630_n25596# 0.359f
C1409 w_55000_n62950# a_55268_n63336# 0.12f
C1410 a_78159_n47589# VDD 0.152f
C1411 16to4_PriorityEncoder_v0p0p1_0.x3.EI a_77639_n50381# 0.088f
C1412 16to4_PriorityEncoder_v0p0p1_0.x1.A VDD 2.17f
C1413 frontAnalog_v0p0p1_4.x65.X CLK 0.0393f
C1414 frontAnalog_v0p0p1_10.x63.A frontAnalog_v0p0p1_10.x65.A 3.16f
C1415 frontAnalog_v0p0p1_2.RSfetsym_0.QN VDD 2.56f
C1416 frontAnalog_v0p0p1_4.x65.X frontAnalog_v0p0p1_4.RSfetsym_0.QN 2.28f
C1417 w_55000_n25150# frontAnalog_v0p0p1_5.x65.A 0.0988f
C1418 16to4_PriorityEncoder_v0p0p1_0.x5.x19.D I14 0.464f
C1419 frontAnalog_v0p0p1_5.x65.A VDD 3.45f
C1420 frontAnalog_v0p0p1_1.x63.A CLK 1.81f
C1421 w_55000_n79150# VDD 0.829f
C1422 VDD I9 6.66f
C1423 a_77605_n44779# VDD 0.614f
C1424 frontAnalog_v0p0p1_8.RSfetsym_0.QN frontAnalog_v0p0p1_8.RSfetsym_0.x1.Y 0.17f
C1425 frontAnalog_v0p0p1_3.x65.X frontAnalog_v0p0p1_3.x63.X 0.136f
C1426 16to4_PriorityEncoder_v0p0p1_0.x5.x17.A a_78065_n41309# 0.2f
C1427 frontAnalog_v0p0p1_15.RSfetsym_0.QN S0 2.28f
C1428 frontAnalog_v0p0p1_15.RSfetsym_0.x2.Y VDD 0.926f
C1429 frontAnalog_v0p0p1_5.RSfetsym_0.x1.Y frontAnalog_v0p0p1_5.RSfetsym_0.x2.Y 0.0254f
C1430 16to4_PriorityEncoder_v0p0p1_0.x5.x14.A 16to4_PriorityEncoder_v0p0p1_0.x5.x22.A 0.0179f
C1431 16to4_PriorityEncoder_v0p0p1_0.x3.EI 16to4_PriorityEncoder_v0p0p1_0.x2.A 0.645f
C1432 frontAnalog_v0p0p1_10.RSfetsym_0.QN I6 0.0512f
C1433 a_53630_n52596# a_55268_n52536# 0.015f
C1434 frontAnalog_v0p0p1_13.x63.X m3_58396_n69150# 0.139f
C1435 16to4_PriorityEncoder_v0p0p1_0.x3.x18.C I3 0.251f
C1436 frontAnalog_v0p0p1_4.x63.X a_57123_n20279# 0.121f
C1437 m3_58396_n74550# VDD 1.3f
C1438 frontAnalog_v0p0p1_6.x63.A a_55268_n30936# 1.24f
C1439 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_14.x63.A 0.0926f
C1440 frontAnalog_v0p0p1_3.RSfetsym_0.QN frontAnalog_v0p0p1_3.RSfetsym_0.x1.Y 0.17f
C1441 w_55000_n19128# VV13 0.798f
C1442 frontAnalog_v0p0p1_2.x65.A VIN 0.653f
C1443 frontAnalog_v0p0p1_3.x63.A VV14 0.587f
C1444 a_57123_n78159# S1 0.119f
C1445 frontAnalog_v0p0p1_4.x63.X CLK 0.785f
C1446 16to4_PriorityEncoder_v0p0p1_0.x5.x16.C I10 0.925f
C1447 frontAnalog_v0p0p1_2.RSfetsym_0.x2.Y VDD 0.926f
C1448 w_55000_n46750# a_53630_n47196# 0.394f
C1449 w_55000_n35328# CLK 0.571f
C1450 w_55000_n46128# a_55268_n47136# 0.149f
C1451 frontAnalog_v0p0p1_1.x63.A frontAnalog_v0p0p1_1.x65.A 3.16f
C1452 w_55000_n52150# frontAnalog_v0p0p1_10.IB 0.0217f
C1453 I1 I0 6.2f
C1454 frontAnalog_v0p0p1_4.RSfetsym_0.QN frontAnalog_v0p0p1_4.x63.X 0.378f
C1455 frontAnalog_v0p0p1_4.x65.X frontAnalog_v0p0p1_4.RSfetsym_0.x2.Y 0.526f
C1456 frontAnalog_v0p0p1_0.x65.A a_55268_n9336# 0.461f
C1457 frontAnalog_v0p0p1_5.x63.A VV12 0.587f
C1458 a_53630_n84996# CLK 0.0136f
C1459 16to4_PriorityEncoder_v0p0p1_0.x3.x14.A VDD 0.462f
C1460 16to4_PriorityEncoder_v0p0p1_0.x3.x18.C I2 0.341f
C1461 16to4_PriorityEncoder_v0p0p1_0.x29.A 16to4_PriorityEncoder_v0p0p1_0.x29.Y 1.51f
C1462 a_77605_n44527# 16to4_PriorityEncoder_v0p0p1_0.x5.x21.B 0.116f
C1463 w_55000_n3550# VDD 0.829f
C1464 16to4_PriorityEncoder_v0p0p1_0.x3.x1.X 16to4_PriorityEncoder_v0p0p1_0.x3.x2.X 0.129f
C1465 a_77605_n39305# I8 0.211f
C1466 a_77605_n40069# I15 0.0614f
C1467 frontAnalog_v0p0p1_8.x63.A VIN 0.186f
C1468 a_53630_n36396# VIN 0.265f
C1469 16to4_PriorityEncoder_v0p0p1_0.x3.EI I1 0.437f
C1470 a_59578_n62370# I4 0.42f
C1471 frontAnalog_v0p0p1_11.x63.A CLK 1.81f
C1472 a_59578_n78570# I1 0.42f
C1473 frontAnalog_v0p0p1_3.x63.A CLK 1.81f
C1474 frontAnalog_v0p0p1_6.RSfetsym_0.QN a_59578_n29970# 0.255f
C1475 frontAnalog_v0p0p1_10.x65.A CLK 2.61f
C1476 a_77637_n40777# VDD 0.318f
C1477 I4 I1 0.432f
C1478 I5 I6 8.44f
C1479 I7 I0 0.403f
C1480 a_53630_n68796# VV4 0.28f
C1481 frontAnalog_v0p0p1_3.RSfetsym_0.x1.Y frontAnalog_v0p0p1_3.RSfetsym_0.x2.Y 0.0254f
C1482 VDD I13 12.2f
C1483 a_78349_n51085# VDD 0.164f
C1484 16to4_PriorityEncoder_v0p0p1_0.x3.x21.B 16to4_PriorityEncoder_v0p0p1_0.x3.x20.X 0.0561f
C1485 frontAnalog_v0p0p1_5.RSfetsym_0.QN frontAnalog_v0p0p1_5.RSfetsym_0.x2.Y 0.018f
C1486 VIN VV11 2.52f
C1487 w_55000_n73128# frontAnalog_v0p0p1_12.x65.A 0.658f
C1488 m3_58396_n52950# I6 0.0416f
C1489 16to4_PriorityEncoder_v0p0p1_0.x3.x21.B a_77605_n52819# 0.0141f
C1490 16to4_PriorityEncoder_v0p0p1_0.x3.EI I7 4.79f
C1491 16to4_PriorityEncoder_v0p0p1_0.x3.EI a_77605_n53805# 0.343f
C1492 w_55000_n73128# w_55000_n73750# 0.327f
C1493 frontAnalog_v0p0p1_4.x63.X frontAnalog_v0p0p1_4.RSfetsym_0.x2.Y 0.0923f
C1494 frontAnalog_v0p0p1_1.RSfetsym_0.QN frontAnalog_v0p0p1_1.RSfetsym_0.x1.Y 0.17f
C1495 a_55268_n52536# CLK 0.236f
C1496 I2 I3 7.24f
C1497 a_78525_n45515# 16to4_PriorityEncoder_v0p0p1_0.x5.x20.X 0.0765f
C1498 I7 I4 0.77f
C1499 16to4_PriorityEncoder_v0p0p1_0.x3.x2.X 16to4_PriorityEncoder_v0p0p1_0.x3.EO 0.0749f
C1500 frontAnalog_v0p0p1_13.x63.A VIN 0.188f
C1501 frontAnalog_v0p0p1_12.x63.A frontAnalog_v0p0p1_12.x65.A 3.16f
C1502 frontAnalog_v0p0p1_5.x63.X a_59577_n25083# 0.28f
C1503 16to4_PriorityEncoder_v0p0p1_0.x5.x14.A 16to4_PriorityEncoder_v0p0p1_0.x5.x11.X 0.0721f
C1504 w_55000_n73750# frontAnalog_v0p0p1_12.x63.A 0.659f
C1505 a_77639_n50381# VDD 0.23f
C1506 a_55268_n41736# VIN 0.177f
C1507 w_55000_n14350# VIN 0.737f
C1508 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_8.x65.A 0.0352f
C1509 frontAnalog_v0p0p1_6.x65.X frontAnalog_v0p0p1_6.x63.X 0.136f
C1510 CLK VV5 5.47f
C1511 16to4_PriorityEncoder_v0p0p1_0.x5.x14.A I12 0.0493f
C1512 16to4_PriorityEncoder_v0p0p1_0.x5.x16.C I14 0.491f
C1513 a_78349_n43045# 16to4_PriorityEncoder_v0p0p1_0.x5.x16.X 0.0673f
C1514 a_57123_n61959# VDD 0.224f
C1515 16to4_PriorityEncoder_v0p0p1_0.x3.EO 16to4_PriorityEncoder_v0p0p1_0.x3.GS 0.9f
C1516 frontAnalog_v0p0p1_12.x65.A CLK 2.61f
C1517 16to4_PriorityEncoder_v0p0p1_0.x5.x19.D a_77605_n45765# 0.0838f
C1518 a_53630_n14796# VDD 0.134f
C1519 m3_58396_n85350# I0 0.0416f
C1520 frontAnalog_v0p0p1_14.RSfetsym_0.x2.Y S1 0.526f
C1521 frontAnalog_v0p0p1_11.RSfetsym_0.x1.Y I4 0.0436f
C1522 w_55000_n73750# CLK 0.535f
C1523 16to4_PriorityEncoder_v0p0p1_0.x2.A VDD 1.89f
C1524 frontAnalog_v0p0p1_10.IB a_55268_n36336# 0.0848f
C1525 frontAnalog_v0p0p1_14.RSfetsym_0.x1.Y I1 0.0436f
C1526 frontAnalog_v0p0p1_5.x63.X m3_58396_n25950# 0.139f
C1527 frontAnalog_v0p0p1_6.RSfetsym_0.QN frontAnalog_v0p0p1_6.RSfetsym_0.x1.Y 0.17f
C1528 frontAnalog_v0p0p1_1.RSfetsym_0.x1.Y VDD 0.733f
C1529 w_55000_n46128# VDD 0.854f
C1530 w_55000_n35328# w_55000_n35950# 0.327f
C1531 frontAnalog_v0p0p1_3.RSfetsym_0.QN frontAnalog_v0p0p1_3.RSfetsym_0.x2.Y 0.018f
C1532 I15 I10 0.444f
C1533 16to4_PriorityEncoder_v0p0p1_0.x5.x22.A a_78065_n41309# 0.077f
C1534 16to4_PriorityEncoder_v0p0p1_0.x36.A 16to4_PriorityEncoder_v0p0p1_0.x36.Y 1.51f
C1535 a_53630_n84996# a_55268_n84936# 0.015f
C1536 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_13.x65.A 0.0352f
C1537 w_55000_n52150# VV7 0.751f
C1538 VIN VV15 2.56f
C1539 frontAnalog_v0p0p1_4.RSfetsym_0.QN a_59577_n19683# 0.418f
C1540 frontAnalog_v0p0p1_1.x65.X frontAnalog_v0p0p1_1.RSfetsym_0.x2.Y 0.526f
C1541 frontAnalog_v0p0p1_1.RSfetsym_0.QN frontAnalog_v0p0p1_1.x63.X 0.378f
C1542 frontAnalog_v0p0p1_14.x65.A VIN 0.655f
C1543 CLK VV16 4.89f
C1544 a_55268_n3936# VV16 0.214f
C1545 a_59578_n62370# VDD 0.0213f
C1546 16to4_PriorityEncoder_v0p0p1_0.x5.x4.A 16to4_PriorityEncoder_v0p0p1_0.x5.x2.X 0.125f
C1547 frontAnalog_v0p0p1_11.x63.A frontAnalog_v0p0p1_11.x65.A 3.16f
C1548 frontAnalog_v0p0p1_3.x63.X a_59577_n14283# 0.28f
C1549 m3_58396_n4350# VDD 1.3f
C1550 frontAnalog_v0p0p1_3.x63.A frontAnalog_v0p0p1_3.x65.A 3.16f
C1551 VDD I1 5.08f
C1552 frontAnalog_v0p0p1_15.x65.A a_57123_n83559# 0.214f
C1553 a_53630_n30996# VDD 0.134f
C1554 16to4_PriorityEncoder_v0p0p1_0.x3.EI 16to4_PriorityEncoder_v0p0p1_0.x3.x19.X 0.0149f
C1555 16to4_PriorityEncoder_v0p0p1_0.x3.x4.A I5 0.0107f
C1556 frontAnalog_v0p0p1_6.RSfetsym_0.x1.Y frontAnalog_v0p0p1_6.RSfetsym_0.x2.Y 0.0254f
C1557 16to4_PriorityEncoder_v0p0p1_0.x3.EI 16to4_PriorityEncoder_v0p0p1_0.x5.x14.A 0.0145f
C1558 w_55000_n2928# a_53630_n3996# 0.359f
C1559 w_55000_n19128# frontAnalog_v0p0p1_10.IB 0.0216f
C1560 w_55000_n56928# VIN 0.866f
C1561 frontAnalog_v0p0p1_10.IB VV7 3.69f
C1562 frontAnalog_v0p0p1_11.RSfetsym_0.QN I4 2.02f
C1563 frontAnalog_v0p0p1_0.x63.A VDD 3.67f
C1564 16to4_PriorityEncoder_v0p0p1_0.x5.x19.C I10 0.447f
C1565 a_53630_n9396# VV15 0.28f
C1566 frontAnalog_v0p0p1_12.x65.X VDD 3.55f
C1567 VDD I7 5.83f
C1568 frontAnalog_v0p0p1_14.RSfetsym_0.QN I1 2.02f
C1569 a_77605_n53805# VDD 0.201f
C1570 a_53630_n9396# VIN 0.265f
C1571 w_55000_n25150# a_55268_n25536# 0.12f
C1572 a_55268_n25536# VDD 0.565f
C1573 frontAnalog_v0p0p1_1.x63.X VDD 3.16f
C1574 a_78349_n43045# 16to4_PriorityEncoder_v0p0p1_0.x5.x15.X 0.219f
C1575 frontAnalog_v0p0p1_10.IB a_53630_n79596# 0.473f
C1576 frontAnalog_v0p0p1_11.x65.A VV5 0.253f
C1577 16to4_PriorityEncoder_v0p0p1_0.x3.x21.B 16to4_PriorityEncoder_v0p0p1_0.x3.x21.X 0.0197f
C1578 I15 I14 5.72f
C1579 16to4_PriorityEncoder_v0p0p1_0.x3.x22.A 16to4_PriorityEncoder_v0p0p1_0.x3.A0 0.132f
C1580 a_59577_n79083# I1 0.29f
C1581 frontAnalog_v0p0p1_0.x63.A a_57123_n9479# 0.212f
C1582 a_53630_n25596# VV12 0.28f
C1583 w_55000_n84550# VDD 0.829f
C1584 16to4_PriorityEncoder_v0p0p1_0.x28.A 16to4_PriorityEncoder_v0p0p1_0.x29.A 0.392f
C1585 frontAnalog_v0p0p1_11.RSfetsym_0.x1.Y VDD 0.733f
C1586 a_78525_n45515# 16to4_PriorityEncoder_v0p0p1_0.x5.x21.X 0.202f
C1587 frontAnalog_v0p0p1_6.x65.A a_57123_n29559# 0.214f
C1588 16to4_PriorityEncoder_v0p0p1_0.x3.x19.D a_77605_n52567# 0.14f
C1589 frontAnalog_v0p0p1_4.x65.A VV13 0.253f
C1590 16to4_PriorityEncoder_v0p0p1_0.x5.x11.X a_78065_n41309# 0.202f
C1591 frontAnalog_v0p0p1_11.RSfetsym_0.x2.Y I4 0.198f
C1592 frontAnalog_v0p0p1_8.x63.X VDD 3.16f
C1593 a_53630_n63396# CLK 0.0136f
C1594 frontAnalog_v0p0p1_12.x63.X VDD 3.16f
C1595 frontAnalog_v0p0p1_6.RSfetsym_0.QN frontAnalog_v0p0p1_6.RSfetsym_0.x2.Y 0.018f
C1596 16to4_PriorityEncoder_v0p0p1_0.x5.A2 a_82906_n43855# 0.208f
C1597 frontAnalog_v0p0p1_10.IB VV1 0.0595f
C1598 m3_58396_n85350# VDD 1.3f
C1599 16to4_PriorityEncoder_v0p0p1_0.x5.x4.A 16to4_PriorityEncoder_v0p0p1_0.x5.x1.X 0.118f
C1600 16to4_PriorityEncoder_v0p0p1_0.x5.x22.A 16to4_PriorityEncoder_v0p0p1_0.x5.x17.A 1.27f
C1601 a_77637_n41087# 16to4_PriorityEncoder_v0p0p1_0.x5.x22.A 0.0288f
C1602 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_6.x63.A 0.0926f
C1603 w_55000_n40728# CLK 0.571f
C1604 w_55000_n57550# frontAnalog_v0p0p1_10.IB 0.0217f
C1605 frontAnalog_v0p0p1_6.x63.X a_59577_n30483# 0.28f
C1606 I10 I8 2.5f
C1607 frontAnalog_v0p0p1_0.x65.A frontAnalog_v0p0p1_0.x65.X 0.0236f
C1608 frontAnalog_v0p0p1_10.IB a_53630_n57996# 0.473f
C1609 16to4_PriorityEncoder_v0p0p1_0.x5.x19.C I14 0.305f
C1610 a_57123_n63479# VDD 0.222f
C1611 16to4_PriorityEncoder_v0p0p1_0.x22.A 16to4_PriorityEncoder_v0p0p1_0.x22.Y 1.51f
C1612 frontAnalog_v0p0p1_9.x63.A CLK 1.81f
C1613 w_55000_n83928# frontAnalog_v0p0p1_15.x63.A 0.0792f
C1614 frontAnalog_v0p0p1_10.IB a_55268_n9336# 0.0848f
C1615 a_59578_n51570# VDD 0.0213f
C1616 a_77637_n49127# I5 0.194f
C1617 a_53630_n68796# VIN 0.265f
C1618 w_55000_n8950# VDD 0.829f
C1619 m3_58396_n9750# I14 0.0416f
C1620 16to4_PriorityEncoder_v0p0p1_0.x1.A 16to4_PriorityEncoder_v0p0p1_0.x3.A2 1.46f
C1621 w_55000_n73128# a_55268_n74136# 0.149f
C1622 w_55000_n73750# a_53630_n74196# 0.394f
C1623 16to4_PriorityEncoder_v0p0p1_0.x5.x18.C I10 0.341f
C1624 16to4_PriorityEncoder_v0p0p1_0.x5.x19.D a_77605_n44527# 0.14f
C1625 16to4_PriorityEncoder_v0p0p1_0.x3.x19.X VDD 0.892f
C1626 16to4_PriorityEncoder_v0p0p1_0.x5.x14.A VDD 0.487f
C1627 frontAnalog_v0p0p1_6.x63.A frontAnalog_v0p0p1_6.x63.X 0.0301f
C1628 16to4_PriorityEncoder_v0p0p1_0.x5.x4.A 16to4_PriorityEncoder_v0p0p1_0.x5.EO 0.0491f
C1629 frontAnalog_v0p0p1_11.RSfetsym_0.QN VDD 2.56f
C1630 16to4_PriorityEncoder_v0p0p1_0.x3.A1 VDD 1.93f
C1631 16to4_PriorityEncoder_v0p0p1_0.x5.x19.D 16to4_PriorityEncoder_v0p0p1_0.x5.x2.X 0.014f
C1632 frontAnalog_v0p0p1_12.x63.A a_55268_n74136# 1.24f
C1633 w_55000_n40728# frontAnalog_v0p0p1_1.x65.A 0.658f
C1634 frontAnalog_v0p0p1_0.x63.X m3_58396_n9750# 0.139f
C1635 frontAnalog_v0p0p1_10.IB a_53630_n47196# 0.473f
C1636 frontAnalog_v0p0p1_6.x65.A VV11 0.253f
C1637 m3_58396_n47550# I7 0.0416f
C1638 16to4_PriorityEncoder_v0p0p1_0.x3.x19.D I5 0.551f
C1639 a_57123_n41879# VDD 0.222f
C1640 frontAnalog_v0p0p1_9.x65.X CLK 0.0407f
C1641 frontAnalog_v0p0p1_8.RSfetsym_0.QN a_59578_n46170# 0.255f
C1642 a_55268_n74136# CLK 0.236f
C1643 a_57123_n85079# R0 0.121f
C1644 frontAnalog_v0p0p1_8.x65.X I7 0.446f
C1645 w_55000_n41350# frontAnalog_v0p0p1_1.x63.A 0.659f
C1646 VV4 VV3 5.64f
C1647 frontAnalog_v0p0p1_4.x63.A VIN 0.194f
C1648 16to4_PriorityEncoder_v0p0p1_0.x35.A 16to4_PriorityEncoder_v0p0p1_0.x36.A 0.392f
C1649 frontAnalog_v0p0p1_6.x63.X m3_58396_n31350# 0.139f
C1650 w_55000_n19750# VIN 0.737f
C1651 frontAnalog_v0p0p1_1.RSfetsym_0.QN frontAnalog_v0p0p1_1.RSfetsym_0.x2.Y 0.018f
C1652 16to4_PriorityEncoder_v0p0p1_0.x3.A2 16to4_PriorityEncoder_v0p0p1_0.x3.x14.A 0.074f
C1653 m3_58396_n42150# I8 0.0416f
C1654 frontAnalog_v0p0p1_11.RSfetsym_0.x2.Y VDD 0.926f
C1655 I14 I8 0.358f
C1656 16to4_PriorityEncoder_v0p0p1_0.x5.x17.A a_77637_n42017# 0.14f
C1657 a_57123_n13359# VDD 0.224f
C1658 16to4_PriorityEncoder_v0p0p1_0.x5.x11.X 16to4_PriorityEncoder_v0p0p1_0.x5.x17.A 0.125f
C1659 VDD VV4 4.13f
C1660 a_77637_n41087# 16to4_PriorityEncoder_v0p0p1_0.x5.x11.X 0.109f
C1661 frontAnalog_v0p0p1_5.x65.A CLK 2.61f
C1662 w_55000_n79150# CLK 0.535f
C1663 frontAnalog_v0p0p1_8.x63.X m3_58396_n47550# 0.139f
C1664 CLK I9 0.01f
C1665 a_59577_n46683# VDD 0.0173f
C1666 16to4_PriorityEncoder_v0p0p1_0.x5.x22.A 16to4_PriorityEncoder_v0p0p1_0.x5.x19.X 0.418f
C1667 frontAnalog_v0p0p1_10.IB a_55268_n68736# 0.0848f
C1668 frontAnalog_v0p0p1_8.x63.A a_55268_n47136# 1.24f
C1669 a_59577_n73683# VDD 0.0173f
C1670 a_55268_n79536# VIN 0.177f
C1671 frontAnalog_v0p0p1_14.x65.A a_55268_n79536# 0.461f
C1672 16to4_PriorityEncoder_v0p0p1_0.x5.x18.C I14 0.301f
C1673 frontAnalog_v0p0p1_11.x63.A a_55268_n63336# 1.24f
C1674 frontAnalog_v0p0p1_8.x65.X frontAnalog_v0p0p1_8.x63.X 0.136f
C1675 w_55000_n51528# VDD 0.854f
C1676 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_4.x65.A 0.0352f
C1677 frontAnalog_v0p0p1_1.RSfetsym_0.x2.Y VDD 0.926f
C1678 16to4_PriorityEncoder_v0p0p1_0.x5.x16.X 16to4_PriorityEncoder_v0p0p1_0.x1.A 0.0159f
C1679 frontAnalog_v0p0p1_6.x65.A VIN 0.655f
C1680 a_57123_n2559# frontAnalog_v0p0p1_2.x65.X 0.119f
C1681 a_59578_n13770# VDD 0.0213f
C1682 frontAnalog_v0p0p1_15.RSfetsym_0.x2.Y R0 0.0923f
C1683 m3_58396_n15150# VDD 1.3f
C1684 w_55000_n2928# VV16 0.798f
C1685 w_55000_n29928# a_55268_n30936# 0.149f
C1686 w_55000_n30550# a_53630_n30996# 0.394f
C1687 a_57123_n29559# VDD 0.224f
C1688 a_77605_n48109# I4 0.208f
C1689 frontAnalog_v0p0p1_9.x65.A a_55268_n52536# 0.461f
C1690 w_55000_n3550# a_55268_n3936# 0.12f
C1691 w_55000_n3550# CLK 0.535f
C1692 frontAnalog_v0p0p1_14.x63.A a_57123_n79679# 0.212f
C1693 w_55000_n24528# frontAnalog_v0p0p1_10.IB 0.0216f
C1694 16to4_PriorityEncoder_v0p0p1_0.x5.x21.B a_77605_n44779# 0.0141f
C1695 16to4_PriorityEncoder_v0p0p1_0.x1.X 16to4_PriorityEncoder_v0p0p1_0.x28.A 0.0747f
C1696 16to4_PriorityEncoder_v0p0p1_0.x3.x22.A I5 0.066f
C1697 a_55268_n63336# VV5 0.215f
C1698 w_55000_n62328# VIN 0.866f
C1699 16to4_PriorityEncoder_v0p0p1_0.x3.A2 16to4_PriorityEncoder_v0p0p1_0.x2.A 0.401f
C1700 frontAnalog_v0p0p1_13.x65.A a_55268_n68736# 0.461f
C1701 a_55268_n57936# VIN 0.177f
C1702 16to4_PriorityEncoder_v0p0p1_0.x3.EI 16to4_PriorityEncoder_v0p0p1_0.x5.x17.A 0.0296f
C1703 a_78065_n41309# VDD 0.161f
C1704 CLK I13 0.01f
C1705 a_78525_n53555# VDD 0.151f
C1706 16to4_PriorityEncoder_v0p0p1_0.x3.x16.C I5 0.415f
C1707 frontAnalog_v0p0p1_9.x63.X a_57123_n52679# 0.121f
C1708 a_55268_n41736# VV9 0.215f
C1709 frontAnalog_v0p0p1_5.x65.X VDD 3.55f
C1710 frontAnalog_v0p0p1_2.x65.A VDD 3.45f
C1711 a_55268_n20136# VV13 0.215f
C1712 frontAnalog_v0p0p1_2.x65.X a_59578_n2970# 0.436f
C1713 w_55000_n67728# VV4 0.798f
C1714 a_53630_n14796# VV14 0.28f
C1715 frontAnalog_v0p0p1_6.x65.X I10 0.446f
C1716 a_59578_n29970# VDD 0.0213f
C1717 16to4_PriorityEncoder_v0p0p1_0.x21.A 16to4_PriorityEncoder_v0p0p1_0.x22.A 0.392f
C1718 frontAnalog_v0p0p1_8.x63.A VDD 3.67f
C1719 16to4_PriorityEncoder_v0p0p1_0.x29.Y VDD 16.6f
C1720 w_55000_n83928# a_53630_n84996# 0.359f
C1721 a_53630_n36396# VDD 0.134f
C1722 w_55000_n56928# a_55268_n57936# 0.149f
C1723 w_55000_n57550# a_53630_n57996# 0.394f
C1724 a_55268_n47136# VIN 0.177f
C1725 frontAnalog_v0p0p1_3.RSfetsym_0.x1.Y VDD 0.733f
C1726 a_57123_n51159# frontAnalog_v0p0p1_9.x65.X 0.119f
C1727 frontAnalog_v0p0p1_9.x65.X I6 0.446f
C1728 a_53630_n14796# CLK 0.0136f
C1729 frontAnalog_v0p0p1_5.x63.X VDD 3.16f
C1730 16to4_PriorityEncoder_v0p0p1_0.x5.x15.X 16to4_PriorityEncoder_v0p0p1_0.x1.A 0.0206f
C1731 VDD VV11 4.38f
C1732 w_55000_n84550# frontAnalog_v0p0p1_15.x65.A 0.0988f
C1733 w_55000_n19128# frontAnalog_v0p0p1_4.x65.A 0.658f
C1734 VIN VV9 2.55f
C1735 a_53630_n74196# a_55268_n74136# 0.015f
C1736 frontAnalog_v0p0p1_6.x63.X I10 1.85f
C1737 16to4_PriorityEncoder_v0p0p1_0.x5.x11.X 16to4_PriorityEncoder_v0p0p1_0.x5.x22.A 0.0936f
C1738 frontAnalog_v0p0p1_14.RSfetsym_0.x1.Y R1 0.883f
C1739 w_55000_n46128# CLK 0.571f
C1740 w_55000_n62950# frontAnalog_v0p0p1_10.IB 0.0217f
C1741 frontAnalog_v0p0p1_9.x63.X frontAnalog_v0p0p1_9.RSfetsym_0.x2.Y 0.0923f
C1742 frontAnalog_v0p0p1_13.x63.A VDD 3.67f
C1743 frontAnalog_v0p0p1_8.RSfetsym_0.QN frontAnalog_v0p0p1_8.RSfetsym_0.x2.Y 0.018f
C1744 frontAnalog_v0p0p1_2.x65.X frontAnalog_v0p0p1_2.RSfetsym_0.x1.Y 0.182f
C1745 w_55000_n19750# frontAnalog_v0p0p1_4.x63.A 0.659f
C1746 a_57123_n14879# VDD 0.222f
C1747 a_77605_n48109# VDD 0.154f
C1748 VV13 VV12 4.41f
C1749 16to4_PriorityEncoder_v0p0p1_0.x3.x19.C a_77605_n52567# 0.157f
C1750 16to4_PriorityEncoder_v0p0p1_0.x3.x11.X I5 0.0201f
C1751 frontAnalog_v0p0p1_12.x65.A a_57123_n72759# 0.214f
C1752 a_55268_n41736# VDD 0.565f
C1753 w_55000_n14350# VDD 0.829f
C1754 16to4_PriorityEncoder_v0p0p1_0.x36.Y VDD 16.6f
C1755 a_53630_n20196# VIN 0.265f
C1756 16to4_PriorityEncoder_v0p0p1_0.x5.x4.A I9 0.0154f
C1757 frontAnalog_v0p0p1_6.RSfetsym_0.x1.Y VDD 0.733f
C1758 16to4_PriorityEncoder_v0p0p1_0.x34.A 16to4_PriorityEncoder_v0p0p1_0.x35.A 0.0737f
C1759 16to4_PriorityEncoder_v0p0p1_0.x5.x2.X I15 0.0129f
C1760 16to4_PriorityEncoder_v0p0p1_0.x3.EI a_77637_n48817# 0.0883f
C1761 16to4_PriorityEncoder_v0p0p1_0.x5.x20.X 16to4_PriorityEncoder_v0p0p1_0.x2.A 0.0148f
C1762 CLK I1 0.0103f
C1763 frontAnalog_v0p0p1_9.x63.X VDD 3.16f
C1764 a_53630_n30996# CLK 0.0136f
C1765 VDD R1 3.16f
C1766 frontAnalog_v0p0p1_3.RSfetsym_0.QN VDD 2.56f
C1767 a_77637_n48817# I4 0.188f
C1768 frontAnalog_v0p0p1_8.RSfetsym_0.QN I8 0.0774f
C1769 16to4_PriorityEncoder_v0p0p1_0.x3.x21.B 16to4_PriorityEncoder_v0p0p1_0.x3.x19.X 0.262f
C1770 VIN VV3 2.63f
C1771 w_55000_n78528# w_55000_n79150# 0.327f
C1772 16to4_PriorityEncoder_v0p0p1_0.x5.x17.A VDD 1.36f
C1773 frontAnalog_v0p0p1_9.x63.X a_59577_n52083# 0.28f
C1774 a_77637_n41087# VDD 0.307f
C1775 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_7.x63.A 0.0926f
C1776 I11 I9 1.73f
C1777 a_53630_n63396# a_55268_n63336# 0.015f
C1778 a_77605_n44779# I11 0.15f
C1779 frontAnalog_v0p0p1_2.RSfetsym_0.x1.Y frontAnalog_v0p0p1_2.x63.X 0.883f
C1780 frontAnalog_v0p0p1_0.x63.A CLK 1.8f
C1781 16to4_PriorityEncoder_v0p0p1_0.x29.A VDD 1.52f
C1782 frontAnalog_v0p0p1_12.x65.X CLK 0.0402f
C1783 CLK I7 0.01f
C1784 VDD VV15 4.05f
C1785 a_55268_n25536# CLK 0.236f
C1786 frontAnalog_v0p0p1_1.x63.X CLK 0.785f
C1787 a_57123_n31079# VDD 0.222f
C1788 frontAnalog_v0p0p1_14.RSfetsym_0.QN R1 0.378f
C1789 w_55000_n25150# VIN 0.737f
C1790 VDD VIN 32.7f
C1791 frontAnalog_v0p0p1_8.x65.A a_57123_n45759# 0.214f
C1792 frontAnalog_v0p0p1_14.x65.A VDD 3.45f
C1793 frontAnalog_v0p0p1_5.x63.A frontAnalog_v0p0p1_5.x65.A 3.16f
C1794 16to4_PriorityEncoder_v0p0p1_0.x3.EI 16to4_PriorityEncoder_v0p0p1_0.x5.x22.A 0.208f
C1795 16to4_PriorityEncoder_v0p0p1_0.x5.x19.C a_77605_n44527# 0.157f
C1796 frontAnalog_v0p0p1_11.x65.A a_57123_n61959# 0.214f
C1797 frontAnalog_v0p0p1_2.x65.X frontAnalog_v0p0p1_2.RSfetsym_0.QN 2.28f
C1798 frontAnalog_v0p0p1_12.x63.A frontAnalog_v0p0p1_12.x63.X 0.0301f
C1799 frontAnalog_v0p0p1_13.x65.X I3 0.446f
C1800 frontAnalog_v0p0p1_3.RSfetsym_0.x2.Y VDD 0.926f
C1801 a_59577_n79083# R1 0.28f
C1802 w_55000_n84550# CLK 0.535f
C1803 frontAnalog_v0p0p1_6.RSfetsym_0.QN VDD 2.56f
C1804 frontAnalog_v0p0p1_10.IB a_55268_n20136# 0.0848f
C1805 a_59577_n25083# VDD 0.0173f
C1806 w_55000_n67728# frontAnalog_v0p0p1_13.x63.A 0.0792f
C1807 16to4_PriorityEncoder_v0p0p1_0.x5.x4.A I13 0.0107f
C1808 16to4_PriorityEncoder_v0p0p1_0.x3.x19.C I5 0.407f
C1809 frontAnalog_v0p0p1_9.x63.A frontAnalog_v0p0p1_9.x65.A 3.16f
C1810 frontAnalog_v0p0p1_2.x63.X a_57123_n4079# 0.121f
C1811 frontAnalog_v0p0p1_8.x63.X CLK 0.785f
C1812 16to4_PriorityEncoder_v0p0p1_0.x3.x19.D a_77605_n52819# 0.148f
C1813 w_55000_n40728# w_55000_n41350# 0.327f
C1814 16to4_PriorityEncoder_v0p0p1_0.x3.A2 16to4_PriorityEncoder_v0p0p1_0.x3.A1 0.787f
C1815 w_55000_n56928# VDD 0.854f
C1816 frontAnalog_v0p0p1_7.x63.A a_55268_n36336# 1.24f
C1817 frontAnalog_v0p0p1_12.x63.X CLK 0.785f
C1818 16to4_PriorityEncoder_v0p0p1_0.x3.x18.C a_77605_n52567# 0.117f
C1819 a_59577_n30483# I10 0.29f
C1820 16to4_PriorityEncoder_v0p0p1_0.x36.A VDD 1.52f
C1821 frontAnalog_v0p0p1_3.x63.A a_55268_n14736# 1.24f
C1822 a_77605_n39305# I10 0.216f
C1823 16to4_PriorityEncoder_v0p0p1_0.x3.x4.A a_78159_n47589# 0.299f
C1824 frontAnalog_v0p0p1_13.x63.A a_57123_n68879# 0.212f
C1825 a_53630_n9396# VDD 0.134f
C1826 frontAnalog_v0p0p1_2.x65.X frontAnalog_v0p0p1_2.RSfetsym_0.x2.Y 0.526f
C1827 frontAnalog_v0p0p1_2.RSfetsym_0.QN frontAnalog_v0p0p1_2.x63.X 0.378f
C1828 frontAnalog_v0p0p1_13.x63.X I3 1.85f
C1829 I13 I11 1.27f
C1830 m3_58396_n25950# VDD 1.3f
C1831 frontAnalog_v0p0p1_15.RSfetsym_0.x1.Y frontAnalog_v0p0p1_15.RSfetsym_0.x2.Y 0.0254f
C1832 frontAnalog_v0p0p1_6.RSfetsym_0.x2.Y VDD 0.926f
C1833 frontAnalog_v0p0p1_9.x65.A frontAnalog_v0p0p1_9.x65.X 0.0236f
C1834 w_55000_n8950# CLK 0.535f
C1835 w_55000_n29928# frontAnalog_v0p0p1_10.IB 0.0216f
C1836 frontAnalog_v0p0p1_7.RSfetsym_0.QN a_59578_n35370# 0.255f
C1837 frontAnalog_v0p0p1_11.x63.A frontAnalog_v0p0p1_11.x63.X 0.0301f
C1838 a_77637_n48817# VDD 0.23f
C1839 16to4_PriorityEncoder_v0p0p1_0.x5.x19.X VDD 0.938f
C1840 m3_58396_n85350# R0 0.14f
C1841 16to4_PriorityEncoder_v0p0p1_0.x2.X 16to4_PriorityEncoder_v0p0p1_0.x21.A 0.0749f
C1842 16to4_PriorityEncoder_v0p0p1_0.x28.A VDD 0.538f
C1843 16to4_PriorityEncoder_v0p0p1_0.x5.x2.X I8 0.0265f
C1844 w_55000_n51528# a_53630_n52596# 0.359f
C1845 w_55000_n67728# VIN 0.866f
C1846 w_55000_n2928# w_55000_n3550# 0.327f
C1847 16to4_PriorityEncoder_v0p0p1_0.x3.x14.A a_78065_n49349# 0.197f
C1848 frontAnalog_v0p0p1_9.x65.X frontAnalog_v0p0p1_9.RSfetsym_0.QN 2.28f
C1849 16to4_PriorityEncoder_v0p0p1_0.x5.x19.D I9 0.937f
C1850 frontAnalog_v0p0p1_13.x65.A frontAnalog_v0p0p1_13.x65.X 0.0236f
C1851 16to4_PriorityEncoder_v0p0p1_0.x5.x19.D a_77605_n44779# 0.148f
C1852 w_55000_n46128# VV8 0.798f
C1853 16to4_PriorityEncoder_v0p0p1_0.x5.x18.C a_77605_n44527# 0.117f
C1854 frontAnalog_v0p0p1_10.IB VV12 3.69f
C1855 frontAnalog_v0p0p1_2.x63.X frontAnalog_v0p0p1_2.RSfetsym_0.x2.Y 0.0923f
C1856 m3_58396_n31350# I10 0.0416f
C1857 frontAnalog_v0p0p1_8.RSfetsym_0.x1.Y I7 0.0436f
C1858 frontAnalog_v0p0p1_7.x65.A VIN 0.655f
C1859 16to4_PriorityEncoder_v0p0p1_0.x5.x22.A VDD 3.25f
C1860 frontAnalog_v0p0p1_7.x65.X frontAnalog_v0p0p1_7.x63.X 0.136f
C1861 16to4_PriorityEncoder_v0p0p1_0.x3.x18.C I5 0.299f
C1862 I6 I1 0.26f
C1863 a_53630_n68796# VDD 0.134f
C1864 w_55000_n19750# a_53630_n20196# 0.394f
C1865 a_57123_n34959# VDD 0.224f
C1866 w_55000_n19128# a_55268_n20136# 0.149f
C1867 w_55000_n84550# a_55268_n84936# 0.12f
C1868 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_15.x63.A 0.0926f
C1869 frontAnalog_v0p0p1_1.x65.X frontAnalog_v0p0p1_1.RSfetsym_0.QN 2.28f
C1870 16to4_PriorityEncoder_v0p0p1_0.x35.A VDD 0.539f
C1871 frontAnalog_v0p0p1_15.RSfetsym_0.QN frontAnalog_v0p0p1_15.RSfetsym_0.x2.Y 0.018f
C1872 a_77605_n47345# I1 0.159f
C1873 frontAnalog_v0p0p1_7.RSfetsym_0.QN frontAnalog_v0p0p1_7.RSfetsym_0.x1.Y 0.17f
C1874 CLK VV4 5.72f
C1875 a_53630_n36396# VV10 0.28f
C1876 VDD OUT3 7.1f
C1877 frontAnalog_v0p0p1_8.RSfetsym_0.x1.Y frontAnalog_v0p0p1_8.x63.X 0.883f
C1878 w_55000_n30550# VV11 0.751f
C1879 I7 I6 5.92f
C1880 16to4_PriorityEncoder_v0p0p1_0.x5.x22.A a_77639_n42341# 0.155f
C1881 16to4_PriorityEncoder_v0p0p1_0.x3.EI I0 0.365f
C1882 w_55000_n51528# CLK 0.571f
C1883 w_55000_n68350# frontAnalog_v0p0p1_10.IB 0.0217f
C1884 16to4_PriorityEncoder_v0p0p1_0.x5.x19.D I13 0.551f
C1885 a_59578_n2970# I15 0.42f
C1886 VV11 VV10 3.38f
C1887 16to4_PriorityEncoder_v0p0p1_0.x43.Y 16to4_PriorityEncoder_v0p0p1_0.x5.A2 0.0114f
C1888 I5 I3 1.27f
C1889 I4 I0 0.575f
C1890 frontAnalog_v0p0p1_11.x63.X m3_58396_n63750# 0.139f
C1891 a_59577_n68283# I3 0.29f
C1892 a_59578_n35370# VDD 0.0213f
C1893 frontAnalog_v0p0p1_2.RSfetsym_0.QN a_59577_n3483# 0.418f
C1894 frontAnalog_v0p0p1_4.x63.A VDD 3.67f
C1895 16to4_PriorityEncoder_v0p0p1_0.x1.X VDD 0.347f
C1896 a_82906_n51645# VDD 0.18f
C1897 frontAnalog_v0p0p1_1.x65.X VDD 3.55f
C1898 w_55000_n19750# VDD 0.829f
C1899 16to4_PriorityEncoder_v0p0p1_0.x3.EI I4 1.8f
C1900 frontAnalog_v0p0p1_7.RSfetsym_0.x1.Y frontAnalog_v0p0p1_7.RSfetsym_0.x2.Y 0.0254f
C1901 w_55000_n79150# VV2 0.751f
C1902 I2 I5 0.649f
C1903 frontAnalog_v0p0p1_10.IB a_53630_n3996# 0.472f
C1904 a_78349_n51085# 16to4_PriorityEncoder_v0p0p1_0.x3.x16.X 0.0673f
C1905 w_55000_n13728# frontAnalog_v0p0p1_3.x63.A 0.0792f
C1906 16to4_PriorityEncoder_v0p0p1_0.x3.x14.A 16to4_PriorityEncoder_v0p0p1_0.x3.x17.A 0.105f
C1907 a_55268_n79536# VDD 0.565f
C1908 16to4_PriorityEncoder_v0p0p1_0.x5.x16.C I9 0.0914f
C1909 frontAnalog_v0p0p1_5.x63.A a_55268_n25536# 1.24f
C1910 a_77637_n42017# VDD 0.322f
C1911 w_55000_n67728# a_53630_n68796# 0.359f
C1912 16to4_PriorityEncoder_v0p0p1_0.x5.x11.X VDD 0.514f
C1913 VDD I12 11.5f
C1914 frontAnalog_v0p0p1_5.x65.X CLK 0.0398f
C1915 16to4_PriorityEncoder_v0p0p1_0.x34.A VDD 0.347f
C1916 frontAnalog_v0p0p1_2.x65.A CLK 2.61f
C1917 frontAnalog_v0p0p1_2.x65.A a_55268_n3936# 0.461f
C1918 frontAnalog_v0p0p1_10.IB VV6 3.7f
C1919 w_55000_n30550# VIN 0.737f
C1920 a_59578_n51570# I6 0.42f
C1921 a_78159_n39549# VDD 0.155f
C1922 16to4_PriorityEncoder_v0p0p1_0.x3.x4.A I1 0.0154f
C1923 w_55000_n68350# frontAnalog_v0p0p1_13.x65.A 0.0988f
C1924 frontAnalog_v0p0p1_2.x63.X m3_58396_n4350# 0.139f
C1925 frontAnalog_v0p0p1_6.x65.A VDD 3.45f
C1926 frontAnalog_v0p0p1_2.RSfetsym_0.x1.Y I15 0.0432f
C1927 16to4_PriorityEncoder_v0p0p1_0.x3.x17.A a_78349_n51085# 0.213f
C1928 frontAnalog_v0p0p1_7.RSfetsym_0.x1.Y VDD 0.733f
C1929 frontAnalog_v0p0p1_7.x65.A a_57123_n34959# 0.214f
C1930 frontAnalog_v0p0p1_2.x63.A VV16 0.587f
C1931 a_78097_n53777# 16to4_PriorityEncoder_v0p0p1_0.x3.x20.X 0.137f
C1932 a_77605_n40069# I14 0.214f
C1933 frontAnalog_v0p0p1_3.x65.A a_57123_n13359# 0.214f
C1934 VIN VV10 2.56f
C1935 frontAnalog_v0p0p1_9.x65.X frontAnalog_v0p0p1_9.RSfetsym_0.x1.Y 0.182f
C1936 frontAnalog_v0p0p1_8.x63.A CLK 1.81f
C1937 a_53630_n36396# CLK 0.0136f
C1938 w_55000_n29928# frontAnalog_v0p0p1_6.x63.A 0.0792f
C1939 frontAnalog_v0p0p1_15.x65.A VIN 0.655f
C1940 frontAnalog_v0p0p1_7.RSfetsym_0.QN frontAnalog_v0p0p1_7.RSfetsym_0.x2.Y 0.018f
C1941 w_55000_n62328# VDD 0.854f
C1942 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_1.x63.A 0.0926f
C1943 16to4_PriorityEncoder_v0p0p1_0.x3.x22.A 16to4_PriorityEncoder_v0p0p1_0.x3.x21.X 0.0749f
C1944 frontAnalog_v0p0p1_5.x63.X CLK 0.785f
C1945 a_55268_n57936# VDD 0.565f
C1946 w_55000_n14350# VV14 0.751f
C1947 VDD I0 4.37f
C1948 a_57123_n7959# VDD 0.224f
C1949 CLK VV11 6.86f
C1950 frontAnalog_v0p0p1_7.x63.X a_59577_n35883# 0.28f
C1951 a_53630_n52596# VIN 0.265f
C1952 frontAnalog_v0p0p1_10.x63.A VIN 0.187f
C1953 16to4_PriorityEncoder_v0p0p1_0.x5.x16.C I13 0.415f
C1954 a_57123_n36479# VDD 0.222f
C1955 frontAnalog_v0p0p1_4.x63.X m3_58396_n20550# 0.139f
C1956 16to4_PriorityEncoder_v0p0p1_0.x3.EI VDD 7.86f
C1957 m3_58396_n36750# VDD 1.3f
C1958 a_78349_n51085# 16to4_PriorityEncoder_v0p0p1_0.x3.x15.X 0.219f
C1959 frontAnalog_v0p0p1_13.x63.A CLK 1.81f
C1960 frontAnalog_v0p0p1_15.x63.A VV1 0.587f
C1961 a_59578_n78570# VDD 0.0213f
C1962 frontAnalog_v0p0p1_15.RSfetsym_0.QN I1 0.0512f
C1963 VDD I4 4.33f
C1964 a_55268_n41736# CLK 0.236f
C1965 w_55000_n14350# CLK 0.535f
C1966 a_55268_n47136# VDD 0.565f
C1967 w_55000_n35328# frontAnalog_v0p0p1_10.IB 0.0216f
C1968 frontAnalog_v0p0p1_2.RSfetsym_0.QN I15 2.02f
C1969 a_57123_n52679# VDD 0.222f
C1970 frontAnalog_v0p0p1_10.IB a_53630_n84996# 0.473f
C1971 frontAnalog_v0p0p1_7.x63.A frontAnalog_v0p0p1_7.x63.X 0.0301f
C1972 frontAnalog_v0p0p1_7.RSfetsym_0.QN VDD 2.56f
C1973 16to4_PriorityEncoder_v0p0p1_0.x3.x19.C a_77605_n52819# 0.102f
C1974 I15 I9 0.29f
C1975 w_55000_n52150# a_55268_n52536# 0.12f
C1976 w_55000_n56928# frontAnalog_v0p0p1_10.x63.A 0.0792f
C1977 frontAnalog_v0p0p1_3.x63.A frontAnalog_v0p0p1_3.x63.X 0.0301f
C1978 w_55000_n73128# VIN 0.866f
C1979 a_59578_n8370# VDD 0.0213f
C1980 VV15 VV14 5.48f
C1981 frontAnalog_v0p0p1_9.x63.X CLK 0.785f
C1982 VIN VV14 2.56f
C1983 CLK R1 0.786f
C1984 frontAnalog_v0p0p1_14.RSfetsym_0.QN a_59578_n78570# 0.255f
C1985 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_11.x63.A 0.0926f
C1986 frontAnalog_v0p0p1_9.RSfetsym_0.QN I7 0.0512f
C1987 VDD VV9 4.76f
C1988 frontAnalog_v0p0p1_4.x65.A a_55268_n20136# 0.461f
C1989 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_3.x63.A 0.0926f
C1990 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_10.x65.A 0.0352f
C1991 frontAnalog_v0p0p1_12.x63.A VIN 0.187f
C1992 I14 I10 0.443f
C1993 VV7 VV6 4.01f
C1994 frontAnalog_v0p0p1_1.x65.A a_55268_n41736# 0.461f
C1995 16to4_PriorityEncoder_v0p0p1_0.x3.x14.A 16to4_PriorityEncoder_v0p0p1_0.x3.x22.A 0.0179f
C1996 frontAnalog_v0p0p1_2.RSfetsym_0.x2.Y I15 0.194f
C1997 CLK VV15 6.32f
C1998 a_57123_n67359# VDD 0.224f
C1999 frontAnalog_v0p0p1_7.RSfetsym_0.x2.Y VDD 0.926f
C2000 frontAnalog_v0p0p1_14.x65.A CLK 2.62f
C2001 CLK VIN 46f
C2002 w_55000_n35950# a_53630_n36396# 0.394f
C2003 w_55000_n35328# a_55268_n36336# 0.149f
C2004 frontAnalog_v0p0p1_10.IB a_55268_n52536# 0.0848f
C2005 a_55268_n3936# VIN 0.177f
C2006 a_53630_n20196# VDD 0.134f
C2007 frontAnalog_v0p0p1_1.RSfetsym_0.QN VDD 2.56f
C2008 frontAnalog_v0p0p1_14.RSfetsym_0.x1.Y VDD 0.733f
C2009 16to4_PriorityEncoder_v0p0p1_0.x5.x19.C I9 0.347f
C2010 frontAnalog_v0p0p1_0.RSfetsym_0.QN a_59578_n8370# 0.255f
C2011 16to4_PriorityEncoder_v0p0p1_0.x3.x19.D I1 0.937f
C2012 16to4_PriorityEncoder_v0p0p1_0.x5.x19.C a_77605_n44779# 0.102f
C2013 16to4_PriorityEncoder_v0p0p1_0.x3.x22.A a_78349_n51085# 0.17f
C2014 frontAnalog_v0p0p1_9.RSfetsym_0.x2.Y VDD 0.926f
C2015 frontAnalog_v0p0p1_10.IB VV5 3.69f
C2016 16to4_PriorityEncoder_v0p0p1_0.x5.x17.A 16to4_PriorityEncoder_v0p0p1_0.x5.x16.X 0.0198f
C2017 16to4_PriorityEncoder_v0p0p1_0.x5.x22.A a_77605_n43295# 0.0116f
C2018 a_57123_n72759# frontAnalog_v0p0p1_12.x65.X 0.119f
C2019 a_78097_n53777# 16to4_PriorityEncoder_v0p0p1_0.x3.x21.X 0.109f
C2020 VDD VV3 4.13f
C2021 frontAnalog_v0p0p1_10.IB frontAnalog_v0p0p1_12.x65.A 0.0352f
C2022 I15 I13 1.14f
C2023 frontAnalog_v0p0p1_0.RSfetsym_0.x1.Y VDD 0.733f
C2024 I1 S1 0.446f
C2025 a_53630_n25596# a_55268_n25536# 0.015f
C2026 w_55000_n56928# CLK 0.571f
C2027 frontAnalog_v0p0p1_0.x65.X I14 0.445f
C2028 w_55000_n73750# frontAnalog_v0p0p1_10.IB 0.0217f
C2029 frontAnalog_v0p0p1_14.RSfetsym_0.QN frontAnalog_v0p0p1_14.RSfetsym_0.x1.Y 0.17f
C2030 frontAnalog_v0p0p1_1.x65.A VIN 0.655f
C2031 a_59578_n67770# VDD 0.0213f
C2032 16to4_PriorityEncoder_v0p0p1_0.x3.x19.D I7 0.244f
C2033 16to4_PriorityEncoder_v0p0p1_0.x3.x19.D a_77605_n53805# 0.0838f
C2034 a_53630_n9396# CLK 0.0136f
C2035 16to4_PriorityEncoder_v0p0p1_0.x3.x22.A a_77639_n50381# 0.155f
C2036 w_55000_n40728# a_53630_n41796# 0.359f
C2037 w_55000_n25150# VDD 0.829f
C2038 frontAnalog_v0p0p1_2.x63.A a_57123_n4079# 0.212f
C2039 w_55000_n14350# frontAnalog_v0p0p1_3.x65.A 0.0988f
C2040 frontAnalog_v0p0p1_9.RSfetsym_0.QN a_59578_n51570# 0.255f
C2041 m3_58396_n79950# I1 0.0416f
C2042 frontAnalog_v0p0p1_5.x65.A a_57123_n24159# 0.214f
C2043 w_55000_n57550# VV6 0.751f
C2044 frontAnalog_v0p0p1_8.x63.A VV8 0.587f
C2045 frontAnalog_v0p0p1_0.x65.X frontAnalog_v0p0p1_0.x63.X 0.136f
C2046 frontAnalog_v0p0p1_5.x65.X I11 0.446f
C2047 a_53630_n57996# VV6 0.28f
C2048 a_77605_n39305# 16to4_PriorityEncoder_v0p0p1_0.x5.x2.X 0.0313f
C2049 a_59577_n52083# VDD 0.0173f
C2050 16to4_PriorityEncoder_v0p0p1_0.x5.EO 16to4_PriorityEncoder_v0p0p1_0.x5.A2 0.136f
C2051 a_59578_n46170# I7 0.42f
C2052 frontAnalog_v0p0p1_10.IB VV16 6.01f
C2053 16to4_PriorityEncoder_v0p0p1_0.x3.A1 16to4_PriorityEncoder_v0p0p1_0.x3.x16.X 0.0159f
C2054 frontAnalog_v0p0p1_12.x65.X a_59578_n73170# 0.436f
C2055 w_55000_n24528# VV12 0.798f
C2056 R0 GND 6.13f
C2057 S0 GND 6.15f
C2058 R1 GND 6.18f
C2059 S1 GND 5.54f
C2060 VL GND 0.131p
C2061 VV1 GND 71.7f
C2062 VV2 GND 80.7f
C2063 OUT0 GND 30.2f
C2064 VV3 GND 76.1f
C2065 VV4 GND 72.1f
C2066 VV5 GND 71.2f
C2067 OUT1 GND 30.3f
C2068 I0 GND 42f
C2069 I3 GND 36.7f
C2070 I1 GND 40.1f
C2071 I6 GND 25.8f
C2072 I5 GND 31f
C2073 I4 GND 30.9f
C2074 I2 GND 38.8f
C2075 I7 GND 23.9f
C2076 VV6 GND 69.4f
C2077 VV7 GND 66.9f
C2078 OUT2 GND 30.2f
C2079 VV8 GND 64.2f
C2080 VV9 GND 60.7f
C2081 OUT3 GND 31.9f
C2082 I8 GND 36.5f
C2083 I9 GND 24f
C2084 VV10 GND 63.8f
C2085 I10 GND 27.6f
C2086 VV11 GND 68.1f
C2087 VFS GND 0.114p
C2088 I11 GND 30.8f
C2089 VV12 GND 72.9f
C2090 I12 GND 34.8f
C2091 VV13 GND 74.3f
C2092 I13 GND 42.8f
C2093 VV14 GND 73.4f
C2094 I14 GND 67.5f
C2095 VV15 GND 76f
C2096 I15 GND 72.7f
C2097 VV16 GND 76.5f
C2098 VIN GND 0.208p
C2099 CLK GND 0.279p
C2100 VDD GND 2.19p
C2101 m3_58396_n85350# GND 0.214f $ **FLOATING
C2102 m3_58396_n79950# GND 0.215f $ **FLOATING
C2103 m3_58396_n74550# GND 0.216f $ **FLOATING
C2104 m3_58396_n69150# GND 0.216f $ **FLOATING
C2105 m3_58396_n63750# GND 0.216f $ **FLOATING
C2106 m3_58396_n58350# GND 0.216f $ **FLOATING
C2107 m3_58396_n52950# GND 0.216f $ **FLOATING
C2108 m3_58396_n47550# GND 0.216f $ **FLOATING
C2109 m3_58396_n42150# GND 0.216f $ **FLOATING
C2110 m3_58396_n36750# GND 0.216f $ **FLOATING
C2111 m3_58396_n31350# GND 0.216f $ **FLOATING
C2112 m3_58396_n25950# GND 0.216f $ **FLOATING
C2113 m3_58396_n20550# GND 0.216f $ **FLOATING
C2114 m3_58396_n15150# GND 0.216f $ **FLOATING
C2115 m3_58396_n9750# GND 0.216f $ **FLOATING
C2116 m3_58396_n4350# GND 0.216f $ **FLOATING
C2117 a_59577_n84483# GND 0.561f
C2118 a_57123_n85079# GND 0.319f
C2119 frontAnalog_v0p0p1_15.RSfetsym_0.x2.Y GND 1.53f
C2120 a_59578_n83970# GND 0.555f
C2121 frontAnalog_v0p0p1_15.RSfetsym_0.x1.Y GND 1.93f
C2122 frontAnalog_v0p0p1_15.RSfetsym_0.QN GND 6.31f
C2123 a_57123_n83559# GND 0.318f
C2124 a_55268_n84936# GND 1.17f
C2125 a_53630_n84996# GND 2.61f
C2126 frontAnalog_v0p0p1_15.x65.A GND 2.63f
C2127 frontAnalog_v0p0p1_15.x63.A GND 2.46f
C2128 a_59577_n79083# GND 0.561f
C2129 a_57123_n79679# GND 0.319f
C2130 frontAnalog_v0p0p1_14.RSfetsym_0.x2.Y GND 1.53f
C2131 a_59578_n78570# GND 0.555f
C2132 frontAnalog_v0p0p1_14.RSfetsym_0.x1.Y GND 1.93f
C2133 frontAnalog_v0p0p1_14.RSfetsym_0.QN GND 6.32f
C2134 a_57123_n78159# GND 0.318f
C2135 a_55268_n79536# GND 1.17f
C2136 a_53630_n79596# GND 2.61f
C2137 frontAnalog_v0p0p1_14.x65.A GND 2.63f
C2138 frontAnalog_v0p0p1_14.x63.A GND 2.46f
C2139 a_59577_n73683# GND 0.561f
C2140 a_57123_n74279# GND 0.319f
C2141 frontAnalog_v0p0p1_12.RSfetsym_0.x2.Y GND 1.53f
C2142 frontAnalog_v0p0p1_12.x63.X GND 5.15f
C2143 a_59578_n73170# GND 0.555f
C2144 frontAnalog_v0p0p1_12.RSfetsym_0.x1.Y GND 1.93f
C2145 frontAnalog_v0p0p1_12.RSfetsym_0.QN GND 6.32f
C2146 frontAnalog_v0p0p1_12.x65.X GND 5.07f
C2147 a_57123_n72759# GND 0.318f
C2148 a_55268_n74136# GND 1.17f
C2149 a_53630_n74196# GND 2.61f
C2150 frontAnalog_v0p0p1_12.x65.A GND 2.64f
C2151 frontAnalog_v0p0p1_12.x63.A GND 2.46f
C2152 a_59577_n68283# GND 0.561f
C2153 a_57123_n68879# GND 0.319f
C2154 frontAnalog_v0p0p1_13.RSfetsym_0.x2.Y GND 1.53f
C2155 frontAnalog_v0p0p1_13.x63.X GND 5.15f
C2156 a_59578_n67770# GND 0.555f
C2157 frontAnalog_v0p0p1_13.RSfetsym_0.x1.Y GND 1.93f
C2158 frontAnalog_v0p0p1_13.RSfetsym_0.QN GND 6.32f
C2159 frontAnalog_v0p0p1_13.x65.X GND 5.07f
C2160 a_57123_n67359# GND 0.318f
C2161 a_55268_n68736# GND 1.17f
C2162 a_53630_n68796# GND 2.61f
C2163 frontAnalog_v0p0p1_13.x65.A GND 2.64f
C2164 frontAnalog_v0p0p1_13.x63.A GND 2.46f
C2165 a_59577_n62883# GND 0.561f
C2166 a_57123_n63479# GND 0.319f
C2167 frontAnalog_v0p0p1_11.RSfetsym_0.x2.Y GND 1.53f
C2168 frontAnalog_v0p0p1_11.x63.X GND 5.15f
C2169 a_59578_n62370# GND 0.555f
C2170 frontAnalog_v0p0p1_11.RSfetsym_0.x1.Y GND 1.93f
C2171 frontAnalog_v0p0p1_11.RSfetsym_0.QN GND 6.32f
C2172 frontAnalog_v0p0p1_11.x65.X GND 5.07f
C2173 a_57123_n61959# GND 0.318f
C2174 a_55268_n63336# GND 1.17f
C2175 a_53630_n63396# GND 2.61f
C2176 frontAnalog_v0p0p1_11.x65.A GND 2.64f
C2177 frontAnalog_v0p0p1_11.x63.A GND 2.46f
C2178 a_59577_n57483# GND 0.561f
C2179 a_57123_n58079# GND 0.319f
C2180 frontAnalog_v0p0p1_10.RSfetsym_0.x2.Y GND 1.53f
C2181 frontAnalog_v0p0p1_10.x63.X GND 5.15f
C2182 a_59578_n56970# GND 0.555f
C2183 frontAnalog_v0p0p1_10.RSfetsym_0.x1.Y GND 1.93f
C2184 frontAnalog_v0p0p1_10.RSfetsym_0.QN GND 6.32f
C2185 frontAnalog_v0p0p1_10.x65.X GND 5.07f
C2186 a_57123_n56559# GND 0.318f
C2187 a_55268_n57936# GND 1.17f
C2188 a_53630_n57996# GND 2.61f
C2189 frontAnalog_v0p0p1_10.x65.A GND 2.64f
C2190 frontAnalog_v0p0p1_10.x63.A GND 2.46f
C2191 16to4_PriorityEncoder_v0p0p1_0.x3.x21.X GND 0.245f
C2192 16to4_PriorityEncoder_v0p0p1_0.x3.x20.X GND 0.69f
C2193 a_78525_n53555# GND 0.366f
C2194 a_78097_n53777# GND 0.22f
C2195 a_77605_n53805# GND 0.296f
C2196 16to4_PriorityEncoder_v0p0p1_0.x3.x19.X GND 0.443f
C2197 a_77605_n52819# GND 0.295f
C2198 16to4_PriorityEncoder_v0p0p1_0.x3.x21.B GND 0.662f
C2199 a_77605_n52567# GND 0.295f
C2200 a_59577_n52083# GND 0.561f
C2201 16to4_PriorityEncoder_v0p0p1_0.x3.A0 GND 7.55f
C2202 a_57123_n52679# GND 0.319f
C2203 frontAnalog_v0p0p1_9.RSfetsym_0.x2.Y GND 1.53f
C2204 frontAnalog_v0p0p1_9.x63.X GND 5.15f
C2205 a_77605_n51585# GND 0.297f
C2206 16to4_PriorityEncoder_v0p0p1_0.x22.Y GND 9.85f
C2207 16to4_PriorityEncoder_v0p0p1_0.x22.A GND 2.13f
C2208 16to4_PriorityEncoder_v0p0p1_0.x21.A GND 0.663f
C2209 16to4_PriorityEncoder_v0p0p1_0.x2.X GND 0.382f
C2210 a_82906_n51645# GND 0.263f
C2211 a_59578_n51570# GND 0.555f
C2212 16to4_PriorityEncoder_v0p0p1_0.x3.x16.X GND 0.871f
C2213 16to4_PriorityEncoder_v0p0p1_0.x3.x15.X GND 0.334f
C2214 frontAnalog_v0p0p1_9.RSfetsym_0.x1.Y GND 1.93f
C2215 a_78349_n51085# GND 0.369f
C2216 a_77605_n51335# GND 0.296f
C2217 frontAnalog_v0p0p1_9.RSfetsym_0.QN GND 6.32f
C2218 frontAnalog_v0p0p1_9.x65.X GND 5.07f
C2219 a_57123_n51159# GND 0.318f
C2220 a_55268_n52536# GND 1.17f
C2221 a_53630_n52596# GND 2.61f
C2222 a_77639_n50381# GND 0.286f
C2223 frontAnalog_v0p0p1_9.x65.A GND 2.64f
C2224 frontAnalog_v0p0p1_9.x63.A GND 2.46f
C2225 a_77637_n50057# GND 0.288f
C2226 a_78065_n49349# GND 0.367f
C2227 16to4_PriorityEncoder_v0p0p1_0.x3.x17.A GND 0.917f
C2228 16to4_PriorityEncoder_v0p0p1_0.x3.x22.A GND 2.02f
C2229 16to4_PriorityEncoder_v0p0p1_0.x3.x11.X GND 0.263f
C2230 a_77637_n49127# GND 0.28f
C2231 16to4_PriorityEncoder_v0p0p1_0.x3.x14.A GND 0.978f
C2232 a_77637_n48817# GND 0.289f
C2233 16to4_PriorityEncoder_v0p0p1_0.x3.A1 GND 5.12f
C2234 16to4_PriorityEncoder_v0p0p1_0.x29.Y GND 9.86f
C2235 16to4_PriorityEncoder_v0p0p1_0.x29.A GND 2.13f
C2236 16to4_PriorityEncoder_v0p0p1_0.x28.A GND 0.665f
C2237 16to4_PriorityEncoder_v0p0p1_0.x1.X GND 0.383f
C2238 a_82906_n47995# GND 0.265f
C2239 a_77605_n48109# GND 0.388f
C2240 16to4_PriorityEncoder_v0p0p1_0.x3.GS GND 2.06f
C2241 16to4_PriorityEncoder_v0p0p1_0.x3.EO GND 2.32f
C2242 16to4_PriorityEncoder_v0p0p1_0.x3.x2.X GND 0.676f
C2243 16to4_PriorityEncoder_v0p0p1_0.x3.x1.X GND 0.162f
C2244 a_78649_n47567# GND 0.258f
C2245 a_78159_n47589# GND 0.343f
C2246 a_77605_n47345# GND 0.379f
C2247 16to4_PriorityEncoder_v0p0p1_0.x3.x4.A GND 1.07f
C2248 16to4_PriorityEncoder_v0p0p1_0.x3.x19.D GND 4.1f
C2249 16to4_PriorityEncoder_v0p0p1_0.x3.x16.C GND 1.84f
C2250 16to4_PriorityEncoder_v0p0p1_0.x3.x19.C GND 4.41f
C2251 16to4_PriorityEncoder_v0p0p1_0.x3.x18.C GND 1.88f
C2252 a_59577_n46683# GND 0.561f
C2253 a_57123_n47279# GND 0.319f
C2254 frontAnalog_v0p0p1_8.RSfetsym_0.x2.Y GND 1.53f
C2255 frontAnalog_v0p0p1_8.x63.X GND 5.15f
C2256 a_59578_n46170# GND 0.555f
C2257 16to4_PriorityEncoder_v0p0p1_0.x2.A GND 6.65f
C2258 16to4_PriorityEncoder_v0p0p1_0.x5.x21.X GND 0.242f
C2259 16to4_PriorityEncoder_v0p0p1_0.x5.x20.X GND 0.684f
C2260 frontAnalog_v0p0p1_8.RSfetsym_0.x1.Y GND 1.93f
C2261 a_78525_n45515# GND 0.364f
C2262 a_78097_n45737# GND 0.217f
C2263 a_77605_n45765# GND 0.291f
C2264 frontAnalog_v0p0p1_8.RSfetsym_0.QN GND 6.29f
C2265 frontAnalog_v0p0p1_8.x65.X GND 5.03f
C2266 a_57123_n45759# GND 0.318f
C2267 a_55268_n47136# GND 1.17f
C2268 a_53630_n47196# GND 2.61f
C2269 16to4_PriorityEncoder_v0p0p1_0.x5.x19.X GND 0.434f
C2270 frontAnalog_v0p0p1_8.x65.A GND 2.64f
C2271 frontAnalog_v0p0p1_8.x63.A GND 2.46f
C2272 a_77605_n44779# GND 0.293f
C2273 16to4_PriorityEncoder_v0p0p1_0.x5.x21.B GND 0.652f
C2274 a_77605_n44527# GND 0.295f
C2275 16to4_PriorityEncoder_v0p0p1_0.x3.A2 GND 7.64f
C2276 16to4_PriorityEncoder_v0p0p1_0.x36.Y GND 9.83f
C2277 16to4_PriorityEncoder_v0p0p1_0.x36.A GND 2.12f
C2278 16to4_PriorityEncoder_v0p0p1_0.x35.A GND 0.662f
C2279 16to4_PriorityEncoder_v0p0p1_0.x34.A GND 0.379f
C2280 a_82906_n43855# GND 0.263f
C2281 a_77605_n43545# GND 0.297f
C2282 16to4_PriorityEncoder_v0p0p1_0.x1.A GND 5.67f
C2283 16to4_PriorityEncoder_v0p0p1_0.x5.x16.X GND 0.871f
C2284 16to4_PriorityEncoder_v0p0p1_0.x5.x15.X GND 0.334f
C2285 a_78349_n43045# GND 0.369f
C2286 a_77605_n43295# GND 0.296f
C2287 a_77639_n42341# GND 0.286f
C2288 a_77637_n42017# GND 0.288f
C2289 16to4_PriorityEncoder_v0p0p1_0.x5.A2 GND 5.29f
C2290 a_78065_n41309# GND 0.367f
C2291 16to4_PriorityEncoder_v0p0p1_0.x5.x17.A GND 0.876f
C2292 16to4_PriorityEncoder_v0p0p1_0.x5.x22.A GND 1.77f
C2293 16to4_PriorityEncoder_v0p0p1_0.x5.x11.X GND 0.263f
C2294 a_77637_n41087# GND 0.28f
C2295 a_59577_n41283# GND 0.561f
C2296 a_57123_n41879# GND 0.319f
C2297 frontAnalog_v0p0p1_1.RSfetsym_0.x2.Y GND 1.51f
C2298 frontAnalog_v0p0p1_1.x63.X GND 5.14f
C2299 16to4_PriorityEncoder_v0p0p1_0.x5.x14.A GND 0.958f
C2300 a_59578_n40770# GND 0.555f
C2301 a_77637_n40777# GND 0.289f
C2302 frontAnalog_v0p0p1_1.RSfetsym_0.x1.Y GND 1.92f
C2303 16to4_PriorityEncoder_v0p0p1_0.x3.EI GND 18.6f
C2304 frontAnalog_v0p0p1_1.RSfetsym_0.QN GND 6.38f
C2305 a_77605_n40069# GND 0.391f
C2306 frontAnalog_v0p0p1_1.x65.X GND 5f
C2307 a_57123_n40359# GND 0.318f
C2308 a_55268_n41736# GND 1.17f
C2309 a_53630_n41796# GND 2.61f
C2310 16to4_PriorityEncoder_v0p0p1_0.x43.Y GND 9.88f
C2311 16to4_PriorityEncoder_v0p0p1_0.x43.A GND 2.02f
C2312 16to4_PriorityEncoder_v0p0p1_0.x42.A GND 0.633f
C2313 16to4_PriorityEncoder_v0p0p1_0.x5.GS GND 2.51f
C2314 frontAnalog_v0p0p1_1.x65.A GND 2.64f
C2315 frontAnalog_v0p0p1_1.x63.A GND 2.46f
C2316 16to4_PriorityEncoder_v0p0p1_0.x5.EO GND 2.62f
C2317 16to4_PriorityEncoder_v0p0p1_0.x5.x2.X GND 0.684f
C2318 16to4_PriorityEncoder_v0p0p1_0.x5.x1.X GND 0.167f
C2319 a_78649_n39527# GND 0.262f
C2320 a_78159_n39549# GND 0.347f
C2321 a_77605_n39305# GND 0.384f
C2322 16to4_PriorityEncoder_v0p0p1_0.x5.x4.A GND 1.5f
C2323 16to4_PriorityEncoder_v0p0p1_0.x5.x19.D GND 4.1f
C2324 16to4_PriorityEncoder_v0p0p1_0.x5.x16.C GND 1.85f
C2325 16to4_PriorityEncoder_v0p0p1_0.x5.x19.C GND 4.42f
C2326 16to4_PriorityEncoder_v0p0p1_0.x5.x18.C GND 1.89f
C2327 a_59577_n35883# GND 0.561f
C2328 a_57123_n36479# GND 0.319f
C2329 frontAnalog_v0p0p1_7.RSfetsym_0.x2.Y GND 1.53f
C2330 frontAnalog_v0p0p1_7.x63.X GND 5.23f
C2331 a_59578_n35370# GND 0.555f
C2332 frontAnalog_v0p0p1_7.RSfetsym_0.x1.Y GND 1.93f
C2333 frontAnalog_v0p0p1_7.RSfetsym_0.QN GND 6.38f
C2334 frontAnalog_v0p0p1_7.x65.X GND 5.07f
C2335 a_57123_n34959# GND 0.318f
C2336 a_55268_n36336# GND 1.17f
C2337 a_53630_n36396# GND 2.61f
C2338 frontAnalog_v0p0p1_7.x65.A GND 2.64f
C2339 frontAnalog_v0p0p1_7.x63.A GND 2.46f
C2340 a_59577_n30483# GND 0.561f
C2341 a_57123_n31079# GND 0.319f
C2342 frontAnalog_v0p0p1_6.RSfetsym_0.x2.Y GND 1.53f
C2343 frontAnalog_v0p0p1_6.x63.X GND 5.17f
C2344 a_59578_n29970# GND 0.555f
C2345 frontAnalog_v0p0p1_6.RSfetsym_0.x1.Y GND 1.93f
C2346 frontAnalog_v0p0p1_6.RSfetsym_0.QN GND 6.32f
C2347 frontAnalog_v0p0p1_6.x65.X GND 5.07f
C2348 a_57123_n29559# GND 0.318f
C2349 a_55268_n30936# GND 1.17f
C2350 a_53630_n30996# GND 2.61f
C2351 frontAnalog_v0p0p1_6.x65.A GND 2.63f
C2352 frontAnalog_v0p0p1_6.x63.A GND 2.46f
C2353 a_59577_n25083# GND 0.561f
C2354 a_57123_n25679# GND 0.319f
C2355 frontAnalog_v0p0p1_5.RSfetsym_0.x2.Y GND 1.53f
C2356 frontAnalog_v0p0p1_5.x63.X GND 5.13f
C2357 a_59578_n24570# GND 0.555f
C2358 frontAnalog_v0p0p1_5.RSfetsym_0.x1.Y GND 1.93f
C2359 frontAnalog_v0p0p1_5.RSfetsym_0.QN GND 6.38f
C2360 frontAnalog_v0p0p1_5.x65.X GND 5.07f
C2361 a_57123_n24159# GND 0.318f
C2362 a_55268_n25536# GND 1.17f
C2363 a_53630_n25596# GND 2.61f
C2364 frontAnalog_v0p0p1_5.x65.A GND 2.64f
C2365 frontAnalog_v0p0p1_5.x63.A GND 2.46f
C2366 a_59577_n19683# GND 0.561f
C2367 a_57123_n20279# GND 0.319f
C2368 frontAnalog_v0p0p1_4.RSfetsym_0.x2.Y GND 1.53f
C2369 frontAnalog_v0p0p1_4.x63.X GND 5.17f
C2370 a_59578_n19170# GND 0.555f
C2371 frontAnalog_v0p0p1_4.RSfetsym_0.x1.Y GND 1.93f
C2372 frontAnalog_v0p0p1_4.RSfetsym_0.QN GND 6.38f
C2373 frontAnalog_v0p0p1_4.x65.X GND 5.07f
C2374 a_57123_n18759# GND 0.318f
C2375 a_55268_n20136# GND 1.17f
C2376 a_53630_n20196# GND 2.61f
C2377 frontAnalog_v0p0p1_4.x65.A GND 2.63f
C2378 frontAnalog_v0p0p1_4.x63.A GND 2.46f
C2379 a_59577_n14283# GND 0.561f
C2380 a_57123_n14879# GND 0.319f
C2381 frontAnalog_v0p0p1_3.RSfetsym_0.x2.Y GND 1.53f
C2382 frontAnalog_v0p0p1_3.x63.X GND 5.17f
C2383 a_59578_n13770# GND 0.555f
C2384 frontAnalog_v0p0p1_3.RSfetsym_0.x1.Y GND 1.93f
C2385 frontAnalog_v0p0p1_3.RSfetsym_0.QN GND 6.31f
C2386 frontAnalog_v0p0p1_3.x65.X GND 5.07f
C2387 a_57123_n13359# GND 0.318f
C2388 a_55268_n14736# GND 1.17f
C2389 a_53630_n14796# GND 2.61f
C2390 frontAnalog_v0p0p1_3.x65.A GND 2.64f
C2391 frontAnalog_v0p0p1_3.x63.A GND 2.46f
C2392 a_59577_n8883# GND 0.561f
C2393 a_57123_n9479# GND 0.319f
C2394 frontAnalog_v0p0p1_0.RSfetsym_0.x2.Y GND 1.53f
C2395 frontAnalog_v0p0p1_0.x63.X GND 5.18f
C2396 a_59578_n8370# GND 0.555f
C2397 frontAnalog_v0p0p1_0.RSfetsym_0.x1.Y GND 1.93f
C2398 frontAnalog_v0p0p1_0.RSfetsym_0.QN GND 6.32f
C2399 frontAnalog_v0p0p1_0.x65.X GND 5.07f
C2400 a_57123_n7959# GND 0.318f
C2401 a_55268_n9336# GND 1.17f
C2402 a_53630_n9396# GND 2.61f
C2403 frontAnalog_v0p0p1_0.x65.A GND 2.64f
C2404 frontAnalog_v0p0p1_0.x63.A GND 2.46f
C2405 a_59577_n3483# GND 0.561f
C2406 a_57123_n4079# GND 0.319f
C2407 frontAnalog_v0p0p1_2.RSfetsym_0.x2.Y GND 1.53f
C2408 frontAnalog_v0p0p1_2.x63.X GND 5.18f
C2409 a_59578_n2970# GND 0.555f
C2410 frontAnalog_v0p0p1_2.RSfetsym_0.x1.Y GND 1.93f
C2411 frontAnalog_v0p0p1_2.RSfetsym_0.QN GND 6.38f
C2412 frontAnalog_v0p0p1_2.x65.X GND 5.07f
C2413 a_57123_n2559# GND 0.318f
C2414 a_55268_n3936# GND 1.17f
C2415 a_53630_n3996# GND 2.61f
C2416 frontAnalog_v0p0p1_10.IB GND 0.288p
C2417 frontAnalog_v0p0p1_2.x65.A GND 2.63f
C2418 frontAnalog_v0p0p1_2.x63.A GND 2.46f
C2419 w_55000_n84550# GND 2.69f
C2420 w_55000_n83928# GND 2.69f
C2421 w_55000_n79150# GND 2.69f
C2422 w_55000_n78528# GND 2.69f
C2423 w_55000_n73750# GND 2.69f
C2424 w_55000_n73128# GND 2.69f
C2425 w_55000_n68350# GND 2.69f
C2426 w_55000_n67728# GND 2.69f
C2427 w_55000_n62950# GND 2.69f
C2428 w_55000_n62328# GND 2.69f
C2429 w_55000_n57550# GND 2.69f
C2430 w_55000_n56928# GND 2.69f
C2431 w_55000_n52150# GND 2.69f
C2432 w_55000_n51528# GND 2.69f
C2433 w_55000_n46750# GND 2.69f
C2434 w_55000_n46128# GND 2.69f
C2435 w_55000_n41350# GND 2.69f
C2436 w_55000_n40728# GND 2.69f
C2437 w_55000_n35950# GND 2.69f
C2438 w_55000_n35328# GND 2.69f
C2439 w_55000_n30550# GND 2.69f
C2440 w_55000_n29928# GND 2.69f
C2441 w_55000_n25150# GND 2.69f
C2442 w_55000_n24528# GND 2.69f
C2443 w_55000_n19750# GND 2.69f
C2444 w_55000_n19128# GND 2.68f
C2445 w_55000_n14350# GND 2.69f
C2446 w_55000_n13728# GND 2.69f
C2447 w_55000_n8950# GND 2.69f
C2448 w_55000_n8328# GND 2.69f
C2449 w_55000_n3550# GND 2.69f
C2450 w_55000_n2928# GND 2.68f
C2451 frontAnalog_v0p0p1_0.x63.A.n0 GND 0.12f
C2452 frontAnalog_v0p0p1_0.x63.A.n1 GND 2.22f
C2453 frontAnalog_v0p0p1_0.x63.A.t6 GND 0.014f
C2454 frontAnalog_v0p0p1_0.x63.A.t5 GND 0.0225f
C2455 frontAnalog_v0p0p1_0.x63.A.n2 GND 0.0465f
C2456 frontAnalog_v0p0p1_0.x63.A.t2 GND 0.151f
C2457 frontAnalog_v0p0p1_0.x63.A.t4 GND 0.0256f
C2458 frontAnalog_v0p0p1_0.x63.A.t3 GND 0.173f
C2459 frontAnalog_v0p0p1_0.x63.A.t7 GND 0.175f
C2460 frontAnalog_v0p0p1_0.x63.A.n3 GND 1f
C2461 frontAnalog_v0p0p1_0.x63.A.n4 GND 0.953f
C2462 frontAnalog_v0p0p1_0.x63.A.t0 GND 0.0156f
C2463 frontAnalog_v0p0p1_0.x63.A.t1 GND 0.334f
C2464 frontAnalog_v0p0p1_0.x63.A.n5 GND 1.25f
C2465 frontAnalog_v0p0p1_0.x65.A.n0 GND 0.139f
C2466 frontAnalog_v0p0p1_0.x65.A.t5 GND 0.028f
C2467 frontAnalog_v0p0p1_0.x65.A.t6 GND 0.0175f
C2468 frontAnalog_v0p0p1_0.x65.A.n1 GND 0.0568f
C2469 frontAnalog_v0p0p1_0.x65.A.t7 GND 0.0318f
C2470 frontAnalog_v0p0p1_0.x65.A.t2 GND 0.141f
C2471 frontAnalog_v0p0p1_0.x65.A.t4 GND 0.219f
C2472 frontAnalog_v0p0p1_0.x65.A.n2 GND 1.37f
C2473 frontAnalog_v0p0p1_0.x65.A.n3 GND 0.898f
C2474 frontAnalog_v0p0p1_0.x65.A.t3 GND 0.463f
C2475 frontAnalog_v0p0p1_0.x65.A.t0 GND 0.0194f
C2476 frontAnalog_v0p0p1_0.x65.A.n4 GND 1.6f
C2477 frontAnalog_v0p0p1_0.x65.A.n5 GND 2.01f
C2478 frontAnalog_v0p0p1_0.x65.A.t1 GND 0.149f
C2479 frontAnalog_v0p0p1_0.x65.A.n6 GND 1.72f
C2480 frontAnalog_v0p0p1_6.x65.A.n0 GND 0.139f
C2481 frontAnalog_v0p0p1_6.x65.A.t6 GND 0.028f
C2482 frontAnalog_v0p0p1_6.x65.A.t7 GND 0.0175f
C2483 frontAnalog_v0p0p1_6.x65.A.n1 GND 0.0568f
C2484 frontAnalog_v0p0p1_6.x65.A.t2 GND 0.149f
C2485 frontAnalog_v0p0p1_6.x65.A.t5 GND 0.0318f
C2486 frontAnalog_v0p0p1_6.x65.A.t3 GND 0.141f
C2487 frontAnalog_v0p0p1_6.x65.A.t4 GND 0.219f
C2488 frontAnalog_v0p0p1_6.x65.A.n2 GND 1.37f
C2489 frontAnalog_v0p0p1_6.x65.A.n3 GND 0.898f
C2490 frontAnalog_v0p0p1_6.x65.A.t1 GND 0.463f
C2491 frontAnalog_v0p0p1_6.x65.A.t0 GND 0.0194f
C2492 frontAnalog_v0p0p1_6.x65.A.n4 GND 1.6f
C2493 frontAnalog_v0p0p1_6.x65.A.n5 GND 2.01f
C2494 frontAnalog_v0p0p1_6.x65.A.n6 GND 1.72f
C2495 frontAnalog_v0p0p1_12.x65.A.n0 GND 0.139f
C2496 frontAnalog_v0p0p1_12.x65.A.t4 GND 0.028f
C2497 frontAnalog_v0p0p1_12.x65.A.t6 GND 0.0175f
C2498 frontAnalog_v0p0p1_12.x65.A.n1 GND 0.0568f
C2499 frontAnalog_v0p0p1_12.x65.A.t3 GND 0.149f
C2500 frontAnalog_v0p0p1_12.x65.A.t7 GND 0.0318f
C2501 frontAnalog_v0p0p1_12.x65.A.t2 GND 0.141f
C2502 frontAnalog_v0p0p1_12.x65.A.t5 GND 0.219f
C2503 frontAnalog_v0p0p1_12.x65.A.n2 GND 1.37f
C2504 frontAnalog_v0p0p1_12.x65.A.n3 GND 0.898f
C2505 frontAnalog_v0p0p1_12.x65.A.t0 GND 0.463f
C2506 frontAnalog_v0p0p1_12.x65.A.t1 GND 0.0194f
C2507 frontAnalog_v0p0p1_12.x65.A.n4 GND 1.6f
C2508 frontAnalog_v0p0p1_12.x65.A.n5 GND 2.01f
C2509 frontAnalog_v0p0p1_12.x65.A.n6 GND 1.72f
C2510 frontAnalog_v0p0p1_2.RSfetsym_0.QN.n0 GND 1.01f
C2511 frontAnalog_v0p0p1_2.RSfetsym_0.QN.t5 GND 0.0321f
C2512 frontAnalog_v0p0p1_2.RSfetsym_0.QN.t6 GND 0.0947f
C2513 frontAnalog_v0p0p1_2.RSfetsym_0.QN.n1 GND 1.49f
C2514 frontAnalog_v0p0p1_2.RSfetsym_0.QN.n2 GND 0.595f
C2515 frontAnalog_v0p0p1_2.RSfetsym_0.QN.t0 GND 0.0368f
C2516 frontAnalog_v0p0p1_2.RSfetsym_0.QN.n3 GND 0.631f
C2517 frontAnalog_v0p0p1_2.RSfetsym_0.QN.t3 GND 0.0322f
C2518 frontAnalog_v0p0p1_2.RSfetsym_0.QN.t4 GND 0.0322f
C2519 frontAnalog_v0p0p1_2.RSfetsym_0.QN.t1 GND 0.0566f
C2520 frontAnalog_v0p0p1_8.x63.A.n0 GND 0.12f
C2521 frontAnalog_v0p0p1_8.x63.A.n1 GND 2.22f
C2522 frontAnalog_v0p0p1_8.x63.A.t7 GND 0.014f
C2523 frontAnalog_v0p0p1_8.x63.A.t5 GND 0.0225f
C2524 frontAnalog_v0p0p1_8.x63.A.n2 GND 0.0465f
C2525 frontAnalog_v0p0p1_8.x63.A.t2 GND 0.151f
C2526 frontAnalog_v0p0p1_8.x63.A.t6 GND 0.0256f
C2527 frontAnalog_v0p0p1_8.x63.A.t3 GND 0.173f
C2528 frontAnalog_v0p0p1_8.x63.A.t4 GND 0.175f
C2529 frontAnalog_v0p0p1_8.x63.A.n3 GND 1f
C2530 frontAnalog_v0p0p1_8.x63.A.n4 GND 0.953f
C2531 frontAnalog_v0p0p1_8.x63.A.t1 GND 0.0156f
C2532 frontAnalog_v0p0p1_8.x63.A.t0 GND 0.334f
C2533 frontAnalog_v0p0p1_8.x63.A.n5 GND 1.25f
C2534 I11.n0 GND 0.0104f
C2535 I11.n2 GND 0.656f
C2536 I11.n3 GND 0.0139f
C2537 I11.n4 GND 0.0107f
C2538 I11.n5 GND 1.18f
C2539 I11.n6 GND 0.54f
C2540 I11.n7 GND 0.672f
C2541 I11.n8 GND 0.176f
C2542 I11.n9 GND 1.1f
C2543 I11.t8 GND 0.0238f
C2544 I11.n10 GND 0.373f
C2545 I11.n11 GND 0.0495f
C2546 I11.n12 GND 0.112f
C2547 I11.n13 GND 0.0744f
C2548 I11.n14 GND 0.0795f
C2549 I11.n15 GND 0.11f
C2550 I11.n16 GND 0.104f
C2551 I11.n17 GND 0.25f
C2552 I11.n18 GND 10.7f
C2553 I11.n19 GND 1.25f
C2554 frontAnalog_v0p0p1_1.RSfetsym_0.QN.n0 GND 1.01f
C2555 frontAnalog_v0p0p1_1.RSfetsym_0.QN.t6 GND 0.0321f
C2556 frontAnalog_v0p0p1_1.RSfetsym_0.QN.t5 GND 0.0947f
C2557 frontAnalog_v0p0p1_1.RSfetsym_0.QN.n1 GND 1.49f
C2558 frontAnalog_v0p0p1_1.RSfetsym_0.QN.n2 GND 0.595f
C2559 frontAnalog_v0p0p1_1.RSfetsym_0.QN.t0 GND 0.0368f
C2560 frontAnalog_v0p0p1_1.RSfetsym_0.QN.n3 GND 0.631f
C2561 frontAnalog_v0p0p1_1.RSfetsym_0.QN.t4 GND 0.0322f
C2562 frontAnalog_v0p0p1_1.RSfetsym_0.QN.t3 GND 0.0322f
C2563 frontAnalog_v0p0p1_1.RSfetsym_0.QN.t1 GND 0.0566f
C2564 I3.n2 GND 0.415f
C2565 I3.n5 GND 0.725f
C2566 I3.n6 GND 0.341f
C2567 I3.n7 GND 0.534f
C2568 I3.t8 GND 0.0148f
C2569 I3.n8 GND 0.232f
C2570 I3.n9 GND 0.0307f
C2571 I3.n10 GND 0.0697f
C2572 I3.n11 GND 0.0462f
C2573 I3.n12 GND 0.0494f
C2574 I3.n13 GND 0.0681f
C2575 I3.n14 GND 0.0644f
C2576 I3.n15 GND 0.148f
C2577 I3.n16 GND 8.61f
C2578 I3.n17 GND 0.854f
C2579 I15.n8 GND 0.145f
C2580 I15.n9 GND 0.314f
C2581 I15.n10 GND 0.13f
C2582 I15.n11 GND 0.181f
C2583 I15.n12 GND 0.0659f
C2584 I15.n13 GND 0.199f
C2585 I15.n14 GND 0.14f
C2586 I15.n15 GND 0.0185f
C2587 I15.n16 GND 0.0419f
C2588 I15.n17 GND 0.0278f
C2589 I15.n18 GND 0.0297f
C2590 I15.n19 GND 0.041f
C2591 I15.n20 GND 0.0388f
C2592 I15.n21 GND 0.101f
C2593 I15.n22 GND 0.335f
C2594 I14.n10 GND 0.0698f
C2595 I14.n11 GND 0.169f
C2596 I14.n14 GND 0.0912f
C2597 I14.n21 GND 0.219f
C2598 I14.n22 GND 0.364f
C2599 I14.n23 GND 0.218f
C2600 I14.n24 GND 0.375f
C2601 I14.n25 GND 0.12f
C2602 I14.n26 GND 0.456f
C2603 I14.t8 GND 0.0161f
C2604 I14.n27 GND 0.253f
C2605 I14.n28 GND 0.0335f
C2606 I14.n29 GND 0.076f
C2607 I14.n30 GND 0.0504f
C2608 I14.n31 GND 0.0539f
C2609 I14.n32 GND 0.0742f
C2610 I14.n33 GND 0.0703f
C2611 I14.n34 GND 0.184f
C2612 I14.n35 GND 0.839f
C2613 frontAnalog_v0p0p1_8.x65.A.n0 GND 0.139f
C2614 frontAnalog_v0p0p1_8.x65.A.t4 GND 0.028f
C2615 frontAnalog_v0p0p1_8.x65.A.t6 GND 0.0175f
C2616 frontAnalog_v0p0p1_8.x65.A.n1 GND 0.0568f
C2617 frontAnalog_v0p0p1_8.x65.A.t2 GND 0.149f
C2618 frontAnalog_v0p0p1_8.x65.A.t7 GND 0.0318f
C2619 frontAnalog_v0p0p1_8.x65.A.t3 GND 0.141f
C2620 frontAnalog_v0p0p1_8.x65.A.t5 GND 0.219f
C2621 frontAnalog_v0p0p1_8.x65.A.n2 GND 1.37f
C2622 frontAnalog_v0p0p1_8.x65.A.n3 GND 0.898f
C2623 frontAnalog_v0p0p1_8.x65.A.t1 GND 0.463f
C2624 frontAnalog_v0p0p1_8.x65.A.t0 GND 0.0194f
C2625 frontAnalog_v0p0p1_8.x65.A.n4 GND 1.6f
C2626 frontAnalog_v0p0p1_8.x65.A.n5 GND 2.01f
C2627 frontAnalog_v0p0p1_8.x65.A.n6 GND 1.72f
C2628 frontAnalog_v0p0p1_11.x63.A.n0 GND 0.12f
C2629 frontAnalog_v0p0p1_11.x63.A.n1 GND 2.22f
C2630 frontAnalog_v0p0p1_11.x63.A.t7 GND 0.014f
C2631 frontAnalog_v0p0p1_11.x63.A.t5 GND 0.0225f
C2632 frontAnalog_v0p0p1_11.x63.A.n2 GND 0.0465f
C2633 frontAnalog_v0p0p1_11.x63.A.t3 GND 0.151f
C2634 frontAnalog_v0p0p1_11.x63.A.t6 GND 0.0256f
C2635 frontAnalog_v0p0p1_11.x63.A.t2 GND 0.173f
C2636 frontAnalog_v0p0p1_11.x63.A.t4 GND 0.175f
C2637 frontAnalog_v0p0p1_11.x63.A.n3 GND 1f
C2638 frontAnalog_v0p0p1_11.x63.A.n4 GND 0.953f
C2639 frontAnalog_v0p0p1_11.x63.A.t0 GND 0.0156f
C2640 frontAnalog_v0p0p1_11.x63.A.t1 GND 0.334f
C2641 frontAnalog_v0p0p1_11.x63.A.n5 GND 1.25f
C2642 I7.n0 GND 0.0144f
C2643 I7.n4 GND 0.0134f
C2644 I7.n8 GND 0.524f
C2645 I7.n9 GND 1.12f
C2646 I7.n10 GND 0.477f
C2647 I7.n11 GND 1.87f
C2648 I7.t6 GND 0.0105f
C2649 I7.t9 GND 0.0322f
C2650 I7.n12 GND 0.505f
C2651 I7.n13 GND 0.0669f
C2652 I7.t0 GND 0.0108f
C2653 I7.n14 GND 0.152f
C2654 I7.n15 GND 0.101f
C2655 I7.n16 GND 0.108f
C2656 I7.t3 GND 0.0108f
C2657 I7.t2 GND 0.0108f
C2658 I7.n17 GND 0.148f
C2659 I7.n18 GND 0.14f
C2660 I7.t4 GND 0.0119f
C2661 I7.n19 GND 0.323f
C2662 I7.n20 GND 4.75f
C2663 I7.n21 GND 2.77f
C2664 frontAnalog_v0p0p1_4.RSfetsym_0.QN.n0 GND 1.01f
C2665 frontAnalog_v0p0p1_4.RSfetsym_0.QN.t6 GND 0.0321f
C2666 frontAnalog_v0p0p1_4.RSfetsym_0.QN.t5 GND 0.0947f
C2667 frontAnalog_v0p0p1_4.RSfetsym_0.QN.n1 GND 1.49f
C2668 frontAnalog_v0p0p1_4.RSfetsym_0.QN.n2 GND 0.595f
C2669 frontAnalog_v0p0p1_4.RSfetsym_0.QN.t1 GND 0.0368f
C2670 frontAnalog_v0p0p1_4.RSfetsym_0.QN.n3 GND 0.631f
C2671 frontAnalog_v0p0p1_4.RSfetsym_0.QN.t2 GND 0.0322f
C2672 frontAnalog_v0p0p1_4.RSfetsym_0.QN.t3 GND 0.0322f
C2673 frontAnalog_v0p0p1_4.RSfetsym_0.QN.t0 GND 0.0566f
C2674 frontAnalog_v0p0p1_12.x63.A.n0 GND 0.12f
C2675 frontAnalog_v0p0p1_12.x63.A.n1 GND 2.22f
C2676 frontAnalog_v0p0p1_12.x63.A.t6 GND 0.014f
C2677 frontAnalog_v0p0p1_12.x63.A.t4 GND 0.0225f
C2678 frontAnalog_v0p0p1_12.x63.A.n2 GND 0.0465f
C2679 frontAnalog_v0p0p1_12.x63.A.t3 GND 0.151f
C2680 frontAnalog_v0p0p1_12.x63.A.t5 GND 0.0256f
C2681 frontAnalog_v0p0p1_12.x63.A.t2 GND 0.173f
C2682 frontAnalog_v0p0p1_12.x63.A.t7 GND 0.175f
C2683 frontAnalog_v0p0p1_12.x63.A.n3 GND 1f
C2684 frontAnalog_v0p0p1_12.x63.A.n4 GND 0.953f
C2685 frontAnalog_v0p0p1_12.x63.A.t1 GND 0.0156f
C2686 frontAnalog_v0p0p1_12.x63.A.t0 GND 0.334f
C2687 frontAnalog_v0p0p1_12.x63.A.n5 GND 1.25f
C2688 frontAnalog_v0p0p1_11.RSfetsym_0.QN.n0 GND 1.01f
C2689 frontAnalog_v0p0p1_11.RSfetsym_0.QN.t6 GND 0.0321f
C2690 frontAnalog_v0p0p1_11.RSfetsym_0.QN.t5 GND 0.0947f
C2691 frontAnalog_v0p0p1_11.RSfetsym_0.QN.n1 GND 1.49f
C2692 frontAnalog_v0p0p1_11.RSfetsym_0.QN.n2 GND 0.595f
C2693 frontAnalog_v0p0p1_11.RSfetsym_0.QN.t4 GND 0.0368f
C2694 frontAnalog_v0p0p1_11.RSfetsym_0.QN.n3 GND 0.631f
C2695 frontAnalog_v0p0p1_11.RSfetsym_0.QN.t0 GND 0.0322f
C2696 frontAnalog_v0p0p1_11.RSfetsym_0.QN.t1 GND 0.0322f
C2697 frontAnalog_v0p0p1_11.RSfetsym_0.QN.t3 GND 0.0566f
C2698 frontAnalog_v0p0p1_13.x65.A.n0 GND 0.139f
C2699 frontAnalog_v0p0p1_13.x65.A.t4 GND 0.028f
C2700 frontAnalog_v0p0p1_13.x65.A.t6 GND 0.0175f
C2701 frontAnalog_v0p0p1_13.x65.A.n1 GND 0.0568f
C2702 frontAnalog_v0p0p1_13.x65.A.t1 GND 0.149f
C2703 frontAnalog_v0p0p1_13.x65.A.t2 GND 0.463f
C2704 frontAnalog_v0p0p1_13.x65.A.t3 GND 0.0194f
C2705 frontAnalog_v0p0p1_13.x65.A.n2 GND 1.6f
C2706 frontAnalog_v0p0p1_13.x65.A.t7 GND 0.0318f
C2707 frontAnalog_v0p0p1_13.x65.A.t0 GND 0.141f
C2708 frontAnalog_v0p0p1_13.x65.A.t5 GND 0.219f
C2709 frontAnalog_v0p0p1_13.x65.A.n3 GND 1.37f
C2710 frontAnalog_v0p0p1_13.x65.A.n4 GND 0.898f
C2711 frontAnalog_v0p0p1_13.x65.A.n5 GND 2.01f
C2712 frontAnalog_v0p0p1_13.x65.A.n6 GND 1.72f
C2713 S1.t5 GND 0.055f
C2714 S1.n0 GND 0.184f
C2715 S1.n1 GND 0.0119f
C2716 S1.n2 GND 0.0137f
C2717 S1.t8 GND 0.0148f
C2718 S1.n4 GND 0.0247f
C2719 S1.t7 GND 0.0148f
C2720 S1.n7 GND 0.0193f
C2721 S1.t3 GND 0.0148f
C2722 S1.n8 GND 0.0213f
C2723 S1.n10 GND 0.0162f
C2724 S1.t2 GND 0.0148f
C2725 S1.n13 GND 0.0199f
C2726 S1.n18 GND 0.0187f
C2727 S1.n19 GND 0.012f
C2728 S1.n21 GND 0.0122f
C2729 S1.n30 GND 0.0135f
C2730 S1.n32 GND 0.0145f
C2731 S1.n33 GND 0.795f
C2732 S1.t9 GND 0.02f
C2733 S1.t10 GND 0.0549f
C2734 S1.n34 GND 0.23f
C2735 S1.n35 GND 0.564f
C2736 S1.n36 GND 0.815f
C2737 S1.n37 GND 0.383f
C2738 S1.n38 GND 0.381f
C2739 S1.t1 GND 0.0217f
C2740 S1.t0 GND 0.0155f
C2741 S1.n40 GND 0.017f
C2742 S1.n41 GND 0.407f
C2743 S1.n42 GND 0.93f
C2744 S1.n43 GND 0.274f
C2745 I8.n1 GND 0.148f
C2746 I8.n2 GND 0.382f
C2747 I8.n3 GND 3f
C2748 I8.t5 GND 0.0145f
C2749 I8.n4 GND 0.228f
C2750 I8.n5 GND 0.0302f
C2751 I8.n6 GND 0.0684f
C2752 I8.n7 GND 0.0454f
C2753 I8.n8 GND 0.0485f
C2754 I8.n9 GND 0.0668f
C2755 I8.n10 GND 0.0632f
C2756 I8.n11 GND 0.165f
C2757 frontAnalog_v0p0p1_0.RSfetsym_0.QN.n0 GND 1.01f
C2758 frontAnalog_v0p0p1_0.RSfetsym_0.QN.t5 GND 0.0321f
C2759 frontAnalog_v0p0p1_0.RSfetsym_0.QN.t6 GND 0.0947f
C2760 frontAnalog_v0p0p1_0.RSfetsym_0.QN.n1 GND 1.49f
C2761 frontAnalog_v0p0p1_0.RSfetsym_0.QN.n2 GND 0.595f
C2762 frontAnalog_v0p0p1_0.RSfetsym_0.QN.t4 GND 0.0368f
C2763 frontAnalog_v0p0p1_0.RSfetsym_0.QN.n3 GND 0.631f
C2764 frontAnalog_v0p0p1_0.RSfetsym_0.QN.t3 GND 0.0322f
C2765 frontAnalog_v0p0p1_0.RSfetsym_0.QN.t2 GND 0.0322f
C2766 frontAnalog_v0p0p1_0.RSfetsym_0.QN.t0 GND 0.0566f
C2767 frontAnalog_v0p0p1_7.RSfetsym_0.QN.n0 GND 1.01f
C2768 frontAnalog_v0p0p1_7.RSfetsym_0.QN.t6 GND 0.0321f
C2769 frontAnalog_v0p0p1_7.RSfetsym_0.QN.t5 GND 0.0947f
C2770 frontAnalog_v0p0p1_7.RSfetsym_0.QN.n1 GND 1.49f
C2771 frontAnalog_v0p0p1_7.RSfetsym_0.QN.n2 GND 0.595f
C2772 frontAnalog_v0p0p1_7.RSfetsym_0.QN.t4 GND 0.0368f
C2773 frontAnalog_v0p0p1_7.RSfetsym_0.QN.n3 GND 0.631f
C2774 frontAnalog_v0p0p1_7.RSfetsym_0.QN.t2 GND 0.0322f
C2775 frontAnalog_v0p0p1_7.RSfetsym_0.QN.t3 GND 0.0322f
C2776 frontAnalog_v0p0p1_7.RSfetsym_0.QN.t0 GND 0.0566f
C2777 frontAnalog_v0p0p1_14.RSfetsym_0.QN.n0 GND 1.23f
C2778 frontAnalog_v0p0p1_14.RSfetsym_0.QN.n1 GND 1.01f
C2779 frontAnalog_v0p0p1_14.RSfetsym_0.QN.t2 GND 0.0566f
C2780 frontAnalog_v0p0p1_14.RSfetsym_0.QN.t4 GND 0.0322f
C2781 frontAnalog_v0p0p1_14.RSfetsym_0.QN.t1 GND 0.0322f
C2782 frontAnalog_v0p0p1_14.RSfetsym_0.QN.t6 GND 0.0321f
C2783 frontAnalog_v0p0p1_14.RSfetsym_0.QN.t5 GND 0.0947f
C2784 frontAnalog_v0p0p1_14.RSfetsym_0.QN.n2 GND 1.49f
C2785 frontAnalog_v0p0p1_14.RSfetsym_0.QN.t0 GND 0.0368f
C2786 frontAnalog_v0p0p1_5.x65.A.n0 GND 0.139f
C2787 frontAnalog_v0p0p1_5.x65.A.t4 GND 0.028f
C2788 frontAnalog_v0p0p1_5.x65.A.t6 GND 0.0175f
C2789 frontAnalog_v0p0p1_5.x65.A.n1 GND 0.0568f
C2790 frontAnalog_v0p0p1_5.x65.A.t1 GND 0.149f
C2791 frontAnalog_v0p0p1_5.x65.A.t2 GND 0.463f
C2792 frontAnalog_v0p0p1_5.x65.A.t3 GND 0.0194f
C2793 frontAnalog_v0p0p1_5.x65.A.n2 GND 1.6f
C2794 frontAnalog_v0p0p1_5.x65.A.t7 GND 0.0318f
C2795 frontAnalog_v0p0p1_5.x65.A.t0 GND 0.141f
C2796 frontAnalog_v0p0p1_5.x65.A.t5 GND 0.219f
C2797 frontAnalog_v0p0p1_5.x65.A.n3 GND 1.37f
C2798 frontAnalog_v0p0p1_5.x65.A.n4 GND 0.898f
C2799 frontAnalog_v0p0p1_5.x65.A.n5 GND 2.01f
C2800 frontAnalog_v0p0p1_5.x65.A.n6 GND 1.72f
C2801 frontAnalog_v0p0p1_1.x63.A.n0 GND 0.12f
C2802 frontAnalog_v0p0p1_1.x63.A.n1 GND 2.22f
C2803 frontAnalog_v0p0p1_1.x63.A.t6 GND 0.014f
C2804 frontAnalog_v0p0p1_1.x63.A.t7 GND 0.0225f
C2805 frontAnalog_v0p0p1_1.x63.A.n2 GND 0.0465f
C2806 frontAnalog_v0p0p1_1.x63.A.t2 GND 0.151f
C2807 frontAnalog_v0p0p1_1.x63.A.t4 GND 0.0256f
C2808 frontAnalog_v0p0p1_1.x63.A.t3 GND 0.173f
C2809 frontAnalog_v0p0p1_1.x63.A.t5 GND 0.175f
C2810 frontAnalog_v0p0p1_1.x63.A.n3 GND 1f
C2811 frontAnalog_v0p0p1_1.x63.A.n4 GND 0.953f
C2812 frontAnalog_v0p0p1_1.x63.A.t0 GND 0.0156f
C2813 frontAnalog_v0p0p1_1.x63.A.t1 GND 0.334f
C2814 frontAnalog_v0p0p1_1.x63.A.n5 GND 1.25f
C2815 I12.n6 GND 0.185f
C2816 I12.n7 GND 0.0109f
C2817 I12.n8 GND 0.03f
C2818 I12.n9 GND 0.325f
C2819 I12.n11 GND 0.142f
C2820 I12.n12 GND 0.302f
C2821 I12.n13 GND 0.398f
C2822 I12.n14 GND 0.59f
C2823 I12.n15 GND 0.167f
C2824 I12.n16 GND 0.886f
C2825 I12.t7 GND 0.0226f
C2826 I12.n17 GND 0.354f
C2827 I12.n18 GND 0.0469f
C2828 I12.n19 GND 0.106f
C2829 I12.n20 GND 0.0705f
C2830 I12.n21 GND 0.0753f
C2831 I12.n22 GND 0.104f
C2832 I12.n23 GND 0.0983f
C2833 I12.n24 GND 0.236f
C2834 I12.n25 GND 12.4f
C2835 I12.n26 GND 1.48f
C2836 VV8.t16 GND 0.022f
C2837 VV8.n0 GND 0.18f
C2838 VV8.n1 GND 0.0872f
C2839 VV8.t15 GND 0.288f
C2840 VV8.t10 GND 0.288f
C2841 VV8.t9 GND 0.288f
C2842 VV8.t14 GND 0.288f
C2843 VV8.t7 GND 0.288f
C2844 VV8.t13 GND 0.288f
C2845 VV8.t8 GND 0.288f
C2846 VV8.t1 GND 0.288f
C2847 VV8.t4 GND 0.288f
C2848 VV8.t12 GND 0.288f
C2849 VV8.t3 GND 0.288f
C2850 VV8.t5 GND 0.288f
C2851 VV8.t0 GND 0.288f
C2852 VV8.t11 GND 0.288f
C2853 VV8.t2 GND 0.288f
C2854 VV8.t6 GND 0.288f
C2855 VV8.n2 GND 0.688f
C2856 VV8.n3 GND 0.707f
C2857 VV8.n4 GND 0.707f
C2858 VV8.n5 GND 0.707f
C2859 VV8.n6 GND 0.707f
C2860 VV8.n7 GND 0.707f
C2861 VV8.n8 GND 0.707f
C2862 VV8.n9 GND 0.63f
C2863 VV8.n10 GND 1.5f
C2864 frontAnalog_v0p0p1_11.x65.A.n0 GND 0.139f
C2865 frontAnalog_v0p0p1_11.x65.A.t4 GND 0.028f
C2866 frontAnalog_v0p0p1_11.x65.A.t6 GND 0.0175f
C2867 frontAnalog_v0p0p1_11.x65.A.n1 GND 0.0568f
C2868 frontAnalog_v0p0p1_11.x65.A.t2 GND 0.149f
C2869 frontAnalog_v0p0p1_11.x65.A.t7 GND 0.0318f
C2870 frontAnalog_v0p0p1_11.x65.A.t3 GND 0.141f
C2871 frontAnalog_v0p0p1_11.x65.A.t5 GND 0.219f
C2872 frontAnalog_v0p0p1_11.x65.A.n2 GND 1.37f
C2873 frontAnalog_v0p0p1_11.x65.A.n3 GND 0.898f
C2874 frontAnalog_v0p0p1_11.x65.A.t0 GND 0.463f
C2875 frontAnalog_v0p0p1_11.x65.A.t1 GND 0.0194f
C2876 frontAnalog_v0p0p1_11.x65.A.n4 GND 1.6f
C2877 frontAnalog_v0p0p1_11.x65.A.n5 GND 2.01f
C2878 frontAnalog_v0p0p1_11.x65.A.n6 GND 1.72f
C2879 frontAnalog_v0p0p1_12.RSfetsym_0.QN.n0 GND 1.01f
C2880 frontAnalog_v0p0p1_12.RSfetsym_0.QN.t6 GND 0.0321f
C2881 frontAnalog_v0p0p1_12.RSfetsym_0.QN.t5 GND 0.0947f
C2882 frontAnalog_v0p0p1_12.RSfetsym_0.QN.n1 GND 1.49f
C2883 frontAnalog_v0p0p1_12.RSfetsym_0.QN.n2 GND 0.595f
C2884 frontAnalog_v0p0p1_12.RSfetsym_0.QN.t4 GND 0.0368f
C2885 frontAnalog_v0p0p1_12.RSfetsym_0.QN.n3 GND 0.631f
C2886 frontAnalog_v0p0p1_12.RSfetsym_0.QN.t2 GND 0.0322f
C2887 frontAnalog_v0p0p1_12.RSfetsym_0.QN.t1 GND 0.0322f
C2888 frontAnalog_v0p0p1_12.RSfetsym_0.QN.t3 GND 0.0566f
C2889 frontAnalog_v0p0p1_6.x63.A.n0 GND 0.12f
C2890 frontAnalog_v0p0p1_6.x63.A.n1 GND 2.22f
C2891 frontAnalog_v0p0p1_6.x63.A.t6 GND 0.014f
C2892 frontAnalog_v0p0p1_6.x63.A.t4 GND 0.0225f
C2893 frontAnalog_v0p0p1_6.x63.A.n2 GND 0.0465f
C2894 frontAnalog_v0p0p1_6.x63.A.t3 GND 0.151f
C2895 frontAnalog_v0p0p1_6.x63.A.t7 GND 0.0256f
C2896 frontAnalog_v0p0p1_6.x63.A.t2 GND 0.173f
C2897 frontAnalog_v0p0p1_6.x63.A.t5 GND 0.175f
C2898 frontAnalog_v0p0p1_6.x63.A.n3 GND 1f
C2899 frontAnalog_v0p0p1_6.x63.A.n4 GND 0.953f
C2900 frontAnalog_v0p0p1_6.x63.A.t1 GND 0.0156f
C2901 frontAnalog_v0p0p1_6.x63.A.t0 GND 0.334f
C2902 frontAnalog_v0p0p1_6.x63.A.n5 GND 1.25f
C2903 frontAnalog_v0p0p1_3.RSfetsym_0.QN.n0 GND 1.01f
C2904 frontAnalog_v0p0p1_3.RSfetsym_0.QN.t6 GND 0.0321f
C2905 frontAnalog_v0p0p1_3.RSfetsym_0.QN.t5 GND 0.0947f
C2906 frontAnalog_v0p0p1_3.RSfetsym_0.QN.n1 GND 1.49f
C2907 frontAnalog_v0p0p1_3.RSfetsym_0.QN.n2 GND 0.595f
C2908 frontAnalog_v0p0p1_3.RSfetsym_0.QN.t0 GND 0.0368f
C2909 frontAnalog_v0p0p1_3.RSfetsym_0.QN.n3 GND 0.631f
C2910 frontAnalog_v0p0p1_3.RSfetsym_0.QN.t3 GND 0.0322f
C2911 frontAnalog_v0p0p1_3.RSfetsym_0.QN.t4 GND 0.0322f
C2912 frontAnalog_v0p0p1_3.RSfetsym_0.QN.t1 GND 0.0566f
C2913 I4.n6 GND 0.166f
C2914 I4.n8 GND 0.0269f
C2915 I4.n9 GND 0.292f
C2916 I4.n11 GND 0.127f
C2917 I4.n12 GND 0.271f
C2918 I4.n13 GND 0.373f
C2919 I4.n14 GND 0.84f
C2920 I4.t12 GND 0.0202f
C2921 I4.n15 GND 0.317f
C2922 I4.n16 GND 0.042f
C2923 I4.n17 GND 0.0953f
C2924 I4.n18 GND 0.0632f
C2925 I4.n19 GND 0.0676f
C2926 I4.n20 GND 0.0931f
C2927 I4.n21 GND 0.0881f
C2928 I4.n22 GND 0.203f
C2929 I4.n23 GND 9.7f
C2930 I4.n24 GND 1.37f
C2931 frontAnalog_v0p0p1_10.RSfetsym_0.QN.n0 GND 1.01f
C2932 frontAnalog_v0p0p1_10.RSfetsym_0.QN.t6 GND 0.0321f
C2933 frontAnalog_v0p0p1_10.RSfetsym_0.QN.t5 GND 0.0947f
C2934 frontAnalog_v0p0p1_10.RSfetsym_0.QN.n1 GND 1.49f
C2935 frontAnalog_v0p0p1_10.RSfetsym_0.QN.n2 GND 0.595f
C2936 frontAnalog_v0p0p1_10.RSfetsym_0.QN.t0 GND 0.0368f
C2937 frontAnalog_v0p0p1_10.RSfetsym_0.QN.n3 GND 0.631f
C2938 frontAnalog_v0p0p1_10.RSfetsym_0.QN.t3 GND 0.0322f
C2939 frontAnalog_v0p0p1_10.RSfetsym_0.QN.t4 GND 0.0322f
C2940 frontAnalog_v0p0p1_10.RSfetsym_0.QN.t1 GND 0.0566f
C2941 frontAnalog_v0p0p1_1.x65.A.n0 GND 0.139f
C2942 frontAnalog_v0p0p1_1.x65.A.t4 GND 0.028f
C2943 frontAnalog_v0p0p1_1.x65.A.t6 GND 0.0175f
C2944 frontAnalog_v0p0p1_1.x65.A.n1 GND 0.0568f
C2945 frontAnalog_v0p0p1_1.x65.A.t2 GND 0.149f
C2946 frontAnalog_v0p0p1_1.x65.A.t7 GND 0.0318f
C2947 frontAnalog_v0p0p1_1.x65.A.t3 GND 0.141f
C2948 frontAnalog_v0p0p1_1.x65.A.t5 GND 0.219f
C2949 frontAnalog_v0p0p1_1.x65.A.n2 GND 1.37f
C2950 frontAnalog_v0p0p1_1.x65.A.n3 GND 0.898f
C2951 frontAnalog_v0p0p1_1.x65.A.t1 GND 0.463f
C2952 frontAnalog_v0p0p1_1.x65.A.t0 GND 0.0194f
C2953 frontAnalog_v0p0p1_1.x65.A.n4 GND 1.6f
C2954 frontAnalog_v0p0p1_1.x65.A.n5 GND 2.01f
C2955 frontAnalog_v0p0p1_1.x65.A.n6 GND 1.72f
C2956 frontAnalog_v0p0p1_4.x63.A.n0 GND 0.12f
C2957 frontAnalog_v0p0p1_4.x63.A.n1 GND 2.22f
C2958 frontAnalog_v0p0p1_4.x63.A.t5 GND 0.014f
C2959 frontAnalog_v0p0p1_4.x63.A.t6 GND 0.0225f
C2960 frontAnalog_v0p0p1_4.x63.A.n2 GND 0.0465f
C2961 frontAnalog_v0p0p1_4.x63.A.t1 GND 0.151f
C2962 frontAnalog_v0p0p1_4.x63.A.t3 GND 0.0156f
C2963 frontAnalog_v0p0p1_4.x63.A.t2 GND 0.335f
C2964 frontAnalog_v0p0p1_4.x63.A.t4 GND 0.0256f
C2965 frontAnalog_v0p0p1_4.x63.A.t0 GND 0.173f
C2966 frontAnalog_v0p0p1_4.x63.A.t7 GND 0.175f
C2967 frontAnalog_v0p0p1_4.x63.A.n3 GND 1f
C2968 frontAnalog_v0p0p1_4.x63.A.n4 GND 0.953f
C2969 frontAnalog_v0p0p1_4.x63.A.n5 GND 1.25f
C2970 frontAnalog_v0p0p1_15.x65.A.n0 GND 0.139f
C2971 frontAnalog_v0p0p1_15.x65.A.t4 GND 0.028f
C2972 frontAnalog_v0p0p1_15.x65.A.t6 GND 0.0175f
C2973 frontAnalog_v0p0p1_15.x65.A.n1 GND 0.0568f
C2974 frontAnalog_v0p0p1_15.x65.A.t1 GND 0.149f
C2975 frontAnalog_v0p0p1_15.x65.A.t2 GND 0.463f
C2976 frontAnalog_v0p0p1_15.x65.A.t3 GND 0.0194f
C2977 frontAnalog_v0p0p1_15.x65.A.n2 GND 1.6f
C2978 frontAnalog_v0p0p1_15.x65.A.t7 GND 0.0318f
C2979 frontAnalog_v0p0p1_15.x65.A.t0 GND 0.141f
C2980 frontAnalog_v0p0p1_15.x65.A.t5 GND 0.219f
C2981 frontAnalog_v0p0p1_15.x65.A.n3 GND 1.37f
C2982 frontAnalog_v0p0p1_15.x65.A.n4 GND 0.898f
C2983 frontAnalog_v0p0p1_15.x65.A.n5 GND 2.01f
C2984 frontAnalog_v0p0p1_15.x65.A.n6 GND 1.72f
C2985 frontAnalog_v0p0p1_3.x65.A.n0 GND 0.139f
C2986 frontAnalog_v0p0p1_3.x65.A.t4 GND 0.028f
C2987 frontAnalog_v0p0p1_3.x65.A.t6 GND 0.0175f
C2988 frontAnalog_v0p0p1_3.x65.A.n1 GND 0.0568f
C2989 frontAnalog_v0p0p1_3.x65.A.t2 GND 0.149f
C2990 frontAnalog_v0p0p1_3.x65.A.t7 GND 0.0318f
C2991 frontAnalog_v0p0p1_3.x65.A.t3 GND 0.141f
C2992 frontAnalog_v0p0p1_3.x65.A.t5 GND 0.219f
C2993 frontAnalog_v0p0p1_3.x65.A.n2 GND 1.37f
C2994 frontAnalog_v0p0p1_3.x65.A.n3 GND 0.898f
C2995 frontAnalog_v0p0p1_3.x65.A.t0 GND 0.463f
C2996 frontAnalog_v0p0p1_3.x65.A.t1 GND 0.0194f
C2997 frontAnalog_v0p0p1_3.x65.A.n4 GND 1.6f
C2998 frontAnalog_v0p0p1_3.x65.A.n5 GND 2.01f
C2999 frontAnalog_v0p0p1_3.x65.A.n6 GND 1.72f
C3000 frontAnalog_v0p0p1_3.x63.A.n0 GND 0.12f
C3001 frontAnalog_v0p0p1_3.x63.A.n1 GND 2.22f
C3002 frontAnalog_v0p0p1_3.x63.A.t7 GND 0.014f
C3003 frontAnalog_v0p0p1_3.x63.A.t5 GND 0.0225f
C3004 frontAnalog_v0p0p1_3.x63.A.n2 GND 0.0465f
C3005 frontAnalog_v0p0p1_3.x63.A.t2 GND 0.151f
C3006 frontAnalog_v0p0p1_3.x63.A.t6 GND 0.0256f
C3007 frontAnalog_v0p0p1_3.x63.A.t3 GND 0.173f
C3008 frontAnalog_v0p0p1_3.x63.A.t4 GND 0.175f
C3009 frontAnalog_v0p0p1_3.x63.A.n3 GND 1f
C3010 frontAnalog_v0p0p1_3.x63.A.n4 GND 0.953f
C3011 frontAnalog_v0p0p1_3.x63.A.t1 GND 0.0156f
C3012 frontAnalog_v0p0p1_3.x63.A.t0 GND 0.334f
C3013 frontAnalog_v0p0p1_3.x63.A.n5 GND 1.25f
C3014 frontAnalog_v0p0p1_5.x63.A.n0 GND 0.12f
C3015 frontAnalog_v0p0p1_5.x63.A.n1 GND 2.22f
C3016 frontAnalog_v0p0p1_5.x63.A.t6 GND 0.014f
C3017 frontAnalog_v0p0p1_5.x63.A.t4 GND 0.0225f
C3018 frontAnalog_v0p0p1_5.x63.A.n2 GND 0.0465f
C3019 frontAnalog_v0p0p1_5.x63.A.t3 GND 0.151f
C3020 frontAnalog_v0p0p1_5.x63.A.t5 GND 0.0256f
C3021 frontAnalog_v0p0p1_5.x63.A.t2 GND 0.173f
C3022 frontAnalog_v0p0p1_5.x63.A.t7 GND 0.175f
C3023 frontAnalog_v0p0p1_5.x63.A.n3 GND 1f
C3024 frontAnalog_v0p0p1_5.x63.A.n4 GND 0.953f
C3025 frontAnalog_v0p0p1_5.x63.A.t0 GND 0.0156f
C3026 frontAnalog_v0p0p1_5.x63.A.t1 GND 0.334f
C3027 frontAnalog_v0p0p1_5.x63.A.n5 GND 1.25f
C3028 frontAnalog_v0p0p1_10.x63.A.n0 GND 0.12f
C3029 frontAnalog_v0p0p1_10.x63.A.n1 GND 2.22f
C3030 frontAnalog_v0p0p1_10.x63.A.t7 GND 0.014f
C3031 frontAnalog_v0p0p1_10.x63.A.t5 GND 0.0225f
C3032 frontAnalog_v0p0p1_10.x63.A.n2 GND 0.0465f
C3033 frontAnalog_v0p0p1_10.x63.A.t2 GND 0.151f
C3034 frontAnalog_v0p0p1_10.x63.A.t6 GND 0.0256f
C3035 frontAnalog_v0p0p1_10.x63.A.t3 GND 0.173f
C3036 frontAnalog_v0p0p1_10.x63.A.t4 GND 0.175f
C3037 frontAnalog_v0p0p1_10.x63.A.n3 GND 1f
C3038 frontAnalog_v0p0p1_10.x63.A.n4 GND 0.953f
C3039 frontAnalog_v0p0p1_10.x63.A.t0 GND 0.0156f
C3040 frontAnalog_v0p0p1_10.x63.A.t1 GND 0.334f
C3041 frontAnalog_v0p0p1_10.x63.A.n5 GND 1.25f
C3042 frontAnalog_v0p0p1_13.x63.A.n0 GND 0.12f
C3043 frontAnalog_v0p0p1_13.x63.A.n1 GND 2.22f
C3044 frontAnalog_v0p0p1_13.x63.A.t6 GND 0.014f
C3045 frontAnalog_v0p0p1_13.x63.A.t4 GND 0.0225f
C3046 frontAnalog_v0p0p1_13.x63.A.n2 GND 0.0465f
C3047 frontAnalog_v0p0p1_13.x63.A.t1 GND 0.151f
C3048 frontAnalog_v0p0p1_13.x63.A.t5 GND 0.0256f
C3049 frontAnalog_v0p0p1_13.x63.A.t2 GND 0.173f
C3050 frontAnalog_v0p0p1_13.x63.A.t7 GND 0.175f
C3051 frontAnalog_v0p0p1_13.x63.A.n3 GND 1f
C3052 frontAnalog_v0p0p1_13.x63.A.n4 GND 0.953f
C3053 frontAnalog_v0p0p1_13.x63.A.t3 GND 0.0156f
C3054 frontAnalog_v0p0p1_13.x63.A.t0 GND 0.334f
C3055 frontAnalog_v0p0p1_13.x63.A.n5 GND 1.25f
C3056 VV5.t16 GND 0.0238f
C3057 VV5.n0 GND 0.195f
C3058 VV5.n1 GND 0.0942f
C3059 VV5.t7 GND 0.311f
C3060 VV5.t1 GND 0.311f
C3061 VV5.t5 GND 0.311f
C3062 VV5.t9 GND 0.311f
C3063 VV5.t0 GND 0.311f
C3064 VV5.t3 GND 0.311f
C3065 VV5.t13 GND 0.311f
C3066 VV5.t12 GND 0.311f
C3067 VV5.t10 GND 0.311f
C3068 VV5.t2 GND 0.311f
C3069 VV5.t4 GND 0.311f
C3070 VV5.t6 GND 0.311f
C3071 VV5.t8 GND 0.311f
C3072 VV5.t14 GND 0.311f
C3073 VV5.t11 GND 0.67f
C3074 VV5.t15 GND 0.311f
C3075 VV5.n2 GND 0.385f
C3076 VV5.n3 GND 0.382f
C3077 VV5.n4 GND 0.382f
C3078 VV5.n5 GND 0.382f
C3079 VV5.n6 GND 0.382f
C3080 VV5.n7 GND 0.382f
C3081 VV5.n8 GND 0.382f
C3082 VV5.n9 GND 0.382f
C3083 VV5.n10 GND 0.382f
C3084 VV5.n11 GND 0.382f
C3085 VV5.n12 GND 0.382f
C3086 VV5.n13 GND 0.382f
C3087 VV5.n14 GND 0.382f
C3088 VV5.n15 GND 0.382f
C3089 VV5.n16 GND 0.306f
C3090 VV5.n17 GND 2.01f
C3091 VV6.t16 GND 0.0241f
C3092 VV6.n0 GND 0.197f
C3093 VV6.n1 GND 0.0955f
C3094 VV6.t5 GND 0.315f
C3095 VV6.t7 GND 0.315f
C3096 VV6.t3 GND 0.315f
C3097 VV6.t15 GND 0.315f
C3098 VV6.t1 GND 0.315f
C3099 VV6.t11 GND 0.315f
C3100 VV6.t12 GND 0.315f
C3101 VV6.t0 GND 0.315f
C3102 VV6.t10 GND 0.315f
C3103 VV6.t6 GND 0.315f
C3104 VV6.t2 GND 0.315f
C3105 VV6.t4 GND 0.315f
C3106 VV6.t8 GND 0.315f
C3107 VV6.t14 GND 0.315f
C3108 VV6.t13 GND 0.315f
C3109 VV6.t9 GND 0.679f
C3110 VV6.n2 GND 0.39f
C3111 VV6.n3 GND 0.387f
C3112 VV6.n4 GND 0.387f
C3113 VV6.n5 GND 0.387f
C3114 VV6.n6 GND 0.387f
C3115 VV6.n7 GND 0.387f
C3116 VV6.n8 GND 0.387f
C3117 VV6.n9 GND 0.387f
C3118 VV6.n10 GND 0.387f
C3119 VV6.n11 GND 0.387f
C3120 VV6.n12 GND 0.387f
C3121 VV6.n13 GND 0.387f
C3122 VV6.n14 GND 0.387f
C3123 VV6.n15 GND 0.387f
C3124 VV6.n16 GND 0.301f
C3125 VV6.n17 GND 1.91f
C3126 VV7.t17 GND 0.0233f
C3127 VV7.n0 GND 0.191f
C3128 VV7.n1 GND 0.0964f
C3129 VV7.t9 GND 0.305f
C3130 VV7.t6 GND 0.305f
C3131 VV7.t13 GND 0.305f
C3132 VV7.t15 GND 0.305f
C3133 VV7.t12 GND 0.305f
C3134 VV7.t8 GND 0.305f
C3135 VV7.t1 GND 0.305f
C3136 VV7.t0 GND 0.305f
C3137 VV7.t11 GND 0.305f
C3138 VV7.t5 GND 0.305f
C3139 VV7.t4 GND 0.305f
C3140 VV7.t3 GND 0.305f
C3141 VV7.t10 GND 0.305f
C3142 VV7.t14 GND 0.305f
C3143 VV7.t7 GND 0.305f
C3144 VV7.t2 GND 0.305f
C3145 VV7.n2 GND 0.73f
C3146 VV7.n3 GND 0.749f
C3147 VV7.n4 GND 0.749f
C3148 VV7.n5 GND 0.749f
C3149 VV7.n6 GND 0.749f
C3150 VV7.n7 GND 0.749f
C3151 VV7.n8 GND 0.749f
C3152 VV7.n9 GND 0.67f
C3153 VV7.n10 GND 1.7f
C3154 I9.t7 GND 0.0147f
C3155 I9.n0 GND 0.872f
C3156 I9.n1 GND 0.0157f
C3157 I9.n2 GND 0.674f
C3158 I9.n3 GND 1.18f
C3159 I9.n4 GND 1.29f
C3160 I9.t10 GND 0.0108f
C3161 I9.t6 GND 0.0331f
C3162 I9.n5 GND 0.519f
C3163 I9.n6 GND 0.0687f
C3164 I9.t4 GND 0.0111f
C3165 I9.n7 GND 0.156f
C3166 I9.n8 GND 0.103f
C3167 I9.n9 GND 0.11f
C3168 I9.t0 GND 0.0111f
C3169 I9.t1 GND 0.0111f
C3170 I9.n10 GND 0.152f
C3171 I9.n11 GND 0.144f
C3172 I9.t3 GND 0.0122f
C3173 I9.n12 GND 0.345f
C3174 I9.n13 GND 5.19f
C3175 I9.n14 GND 3.04f
C3176 frontAnalog_v0p0p1_7.x63.A.n0 GND 0.12f
C3177 frontAnalog_v0p0p1_7.x63.A.n1 GND 2.22f
C3178 frontAnalog_v0p0p1_7.x63.A.t4 GND 0.014f
C3179 frontAnalog_v0p0p1_7.x63.A.t6 GND 0.0225f
C3180 frontAnalog_v0p0p1_7.x63.A.n2 GND 0.0465f
C3181 frontAnalog_v0p0p1_7.x63.A.t2 GND 0.151f
C3182 frontAnalog_v0p0p1_7.x63.A.t7 GND 0.0256f
C3183 frontAnalog_v0p0p1_7.x63.A.t3 GND 0.173f
C3184 frontAnalog_v0p0p1_7.x63.A.t5 GND 0.175f
C3185 frontAnalog_v0p0p1_7.x63.A.n3 GND 1f
C3186 frontAnalog_v0p0p1_7.x63.A.n4 GND 0.953f
C3187 frontAnalog_v0p0p1_7.x63.A.t0 GND 0.0156f
C3188 frontAnalog_v0p0p1_7.x63.A.t1 GND 0.334f
C3189 frontAnalog_v0p0p1_7.x63.A.n5 GND 1.25f
C3190 frontAnalog_v0p0p1_7.x65.A.n0 GND 0.139f
C3191 frontAnalog_v0p0p1_7.x65.A.t7 GND 0.028f
C3192 frontAnalog_v0p0p1_7.x65.A.t5 GND 0.0175f
C3193 frontAnalog_v0p0p1_7.x65.A.n1 GND 0.0568f
C3194 frontAnalog_v0p0p1_7.x65.A.t2 GND 0.149f
C3195 frontAnalog_v0p0p1_7.x65.A.t3 GND 0.463f
C3196 frontAnalog_v0p0p1_7.x65.A.t0 GND 0.0194f
C3197 frontAnalog_v0p0p1_7.x65.A.n2 GND 1.6f
C3198 frontAnalog_v0p0p1_7.x65.A.t6 GND 0.0318f
C3199 frontAnalog_v0p0p1_7.x65.A.t1 GND 0.141f
C3200 frontAnalog_v0p0p1_7.x65.A.t4 GND 0.219f
C3201 frontAnalog_v0p0p1_7.x65.A.n3 GND 1.37f
C3202 frontAnalog_v0p0p1_7.x65.A.n4 GND 0.898f
C3203 frontAnalog_v0p0p1_7.x65.A.n5 GND 2.01f
C3204 frontAnalog_v0p0p1_7.x65.A.n6 GND 1.72f
C3205 frontAnalog_v0p0p1_13.RSfetsym_0.QN.n0 GND 1.01f
C3206 frontAnalog_v0p0p1_13.RSfetsym_0.QN.t6 GND 0.0321f
C3207 frontAnalog_v0p0p1_13.RSfetsym_0.QN.t5 GND 0.0947f
C3208 frontAnalog_v0p0p1_13.RSfetsym_0.QN.n1 GND 1.49f
C3209 frontAnalog_v0p0p1_13.RSfetsym_0.QN.n2 GND 0.595f
C3210 frontAnalog_v0p0p1_13.RSfetsym_0.QN.t1 GND 0.0368f
C3211 frontAnalog_v0p0p1_13.RSfetsym_0.QN.n3 GND 0.631f
C3212 frontAnalog_v0p0p1_13.RSfetsym_0.QN.t4 GND 0.0322f
C3213 frontAnalog_v0p0p1_13.RSfetsym_0.QN.t3 GND 0.0322f
C3214 frontAnalog_v0p0p1_13.RSfetsym_0.QN.t0 GND 0.0566f
C3215 I6.n0 GND 0.0126f
C3216 I6.n2 GND 0.0175f
C3217 I6.n10 GND 0.155f
C3218 I6.n11 GND 0.393f
C3219 I6.n12 GND 0.0114f
C3220 I6.n13 GND 0.0116f
C3221 I6.n14 GND 0.203f
C3222 I6.n17 GND 0.0149f
C3223 I6.n21 GND 0.487f
C3224 I6.n22 GND 0.793f
C3225 I6.n23 GND 0.497f
C3226 I6.n24 GND 1.87f
C3227 I6.t9 GND 0.0117f
C3228 I6.t5 GND 0.0359f
C3229 I6.n25 GND 0.563f
C3230 I6.n26 GND 0.0746f
C3231 I6.t1 GND 0.0121f
C3232 I6.n27 GND 0.169f
C3233 I6.n28 GND 0.112f
C3234 I6.n29 GND 0.12f
C3235 I6.t2 GND 0.0121f
C3236 I6.t3 GND 0.0121f
C3237 I6.n30 GND 0.165f
C3238 I6.n31 GND 0.156f
C3239 I6.t0 GND 0.0132f
C3240 I6.n32 GND 0.36f
C3241 I6.n33 GND 9.83f
C3242 I6.n34 GND 3.13f
C3243 frontAnalog_v0p0p1_9.RSfetsym_0.QN.n0 GND 1.01f
C3244 frontAnalog_v0p0p1_9.RSfetsym_0.QN.t6 GND 0.0321f
C3245 frontAnalog_v0p0p1_9.RSfetsym_0.QN.t5 GND 0.0947f
C3246 frontAnalog_v0p0p1_9.RSfetsym_0.QN.n1 GND 1.49f
C3247 frontAnalog_v0p0p1_9.RSfetsym_0.QN.n2 GND 0.595f
C3248 frontAnalog_v0p0p1_9.RSfetsym_0.QN.t4 GND 0.0368f
C3249 frontAnalog_v0p0p1_9.RSfetsym_0.QN.n3 GND 0.631f
C3250 frontAnalog_v0p0p1_9.RSfetsym_0.QN.t2 GND 0.0322f
C3251 frontAnalog_v0p0p1_9.RSfetsym_0.QN.t3 GND 0.0322f
C3252 frontAnalog_v0p0p1_9.RSfetsym_0.QN.t0 GND 0.0566f
C3253 I1.n0 GND 0.369f
C3254 I1.n2 GND 0.274f
C3255 I1.n3 GND 0.487f
C3256 I1.n4 GND 0.183f
C3257 I1.t5 GND 0.0138f
C3258 I1.n5 GND 0.216f
C3259 I1.n6 GND 0.0286f
C3260 I1.n7 GND 0.0648f
C3261 I1.n8 GND 0.043f
C3262 I1.n9 GND 0.046f
C3263 I1.n10 GND 0.0634f
C3264 I1.n11 GND 0.0599f
C3265 I1.n12 GND 0.138f
C3266 I1.n13 GND 10.8f
C3267 I1.n14 GND 0.53f
C3268 frontAnalog_v0p0p1_9.x65.A.n0 GND 0.139f
C3269 frontAnalog_v0p0p1_9.x65.A.t6 GND 0.028f
C3270 frontAnalog_v0p0p1_9.x65.A.t4 GND 0.0175f
C3271 frontAnalog_v0p0p1_9.x65.A.n1 GND 0.0568f
C3272 frontAnalog_v0p0p1_9.x65.A.t2 GND 0.149f
C3273 frontAnalog_v0p0p1_9.x65.A.t5 GND 0.0318f
C3274 frontAnalog_v0p0p1_9.x65.A.t3 GND 0.141f
C3275 frontAnalog_v0p0p1_9.x65.A.t7 GND 0.219f
C3276 frontAnalog_v0p0p1_9.x65.A.n2 GND 1.37f
C3277 frontAnalog_v0p0p1_9.x65.A.n3 GND 0.898f
C3278 frontAnalog_v0p0p1_9.x65.A.t1 GND 0.463f
C3279 frontAnalog_v0p0p1_9.x65.A.t0 GND 0.0194f
C3280 frontAnalog_v0p0p1_9.x65.A.n4 GND 1.6f
C3281 frontAnalog_v0p0p1_9.x65.A.n5 GND 2.01f
C3282 frontAnalog_v0p0p1_9.x65.A.n6 GND 1.72f
C3283 frontAnalog_v0p0p1_9.x63.A.n0 GND 0.12f
C3284 frontAnalog_v0p0p1_9.x63.A.n1 GND 2.22f
C3285 frontAnalog_v0p0p1_9.x63.A.t7 GND 0.014f
C3286 frontAnalog_v0p0p1_9.x63.A.t5 GND 0.0225f
C3287 frontAnalog_v0p0p1_9.x63.A.n2 GND 0.0465f
C3288 frontAnalog_v0p0p1_9.x63.A.t2 GND 0.151f
C3289 frontAnalog_v0p0p1_9.x63.A.t6 GND 0.0256f
C3290 frontAnalog_v0p0p1_9.x63.A.t3 GND 0.173f
C3291 frontAnalog_v0p0p1_9.x63.A.t4 GND 0.175f
C3292 frontAnalog_v0p0p1_9.x63.A.n3 GND 1f
C3293 frontAnalog_v0p0p1_9.x63.A.n4 GND 0.953f
C3294 frontAnalog_v0p0p1_9.x63.A.t0 GND 0.0156f
C3295 frontAnalog_v0p0p1_9.x63.A.t1 GND 0.334f
C3296 frontAnalog_v0p0p1_9.x63.A.n5 GND 1.25f
C3297 VV12.t16 GND 0.0235f
C3298 VV12.n0 GND 0.193f
C3299 VV12.n1 GND 0.0932f
C3300 VV12.t2 GND 0.308f
C3301 VV12.t0 GND 0.308f
C3302 VV12.t15 GND 0.308f
C3303 VV12.t14 GND 0.308f
C3304 VV12.t5 GND 0.308f
C3305 VV12.t9 GND 0.308f
C3306 VV12.t8 GND 0.308f
C3307 VV12.t10 GND 0.308f
C3308 VV12.t4 GND 0.308f
C3309 VV12.t13 GND 0.308f
C3310 VV12.t1 GND 0.308f
C3311 VV12.t3 GND 0.308f
C3312 VV12.t12 GND 0.308f
C3313 VV12.t11 GND 0.308f
C3314 VV12.t6 GND 0.308f
C3315 VV12.t7 GND 0.664f
C3316 VV12.n2 GND 0.381f
C3317 VV12.n3 GND 0.378f
C3318 VV12.n4 GND 0.378f
C3319 VV12.n5 GND 0.378f
C3320 VV12.n6 GND 0.378f
C3321 VV12.n7 GND 0.378f
C3322 VV12.n8 GND 0.378f
C3323 VV12.n9 GND 0.378f
C3324 VV12.n10 GND 0.378f
C3325 VV12.n11 GND 0.378f
C3326 VV12.n12 GND 0.378f
C3327 VV12.n13 GND 0.378f
C3328 VV12.n14 GND 0.378f
C3329 VV12.n15 GND 0.378f
C3330 VV12.n16 GND 0.298f
C3331 VV12.n17 GND 2.08f
C3332 frontAnalog_v0p0p1_4.x65.A.n0 GND 0.139f
C3333 frontAnalog_v0p0p1_4.x65.A.t4 GND 0.028f
C3334 frontAnalog_v0p0p1_4.x65.A.t5 GND 0.0175f
C3335 frontAnalog_v0p0p1_4.x65.A.n1 GND 0.0568f
C3336 frontAnalog_v0p0p1_4.x65.A.t7 GND 0.0318f
C3337 frontAnalog_v0p0p1_4.x65.A.t1 GND 0.141f
C3338 frontAnalog_v0p0p1_4.x65.A.t6 GND 0.219f
C3339 frontAnalog_v0p0p1_4.x65.A.n2 GND 1.37f
C3340 frontAnalog_v0p0p1_4.x65.A.n3 GND 0.898f
C3341 frontAnalog_v0p0p1_4.x65.A.t3 GND 0.463f
C3342 frontAnalog_v0p0p1_4.x65.A.t2 GND 0.0194f
C3343 frontAnalog_v0p0p1_4.x65.A.n4 GND 1.6f
C3344 frontAnalog_v0p0p1_4.x65.A.n5 GND 2.01f
C3345 frontAnalog_v0p0p1_4.x65.A.t0 GND 0.149f
C3346 frontAnalog_v0p0p1_4.x65.A.n6 GND 1.72f
C3347 R0.t5 GND 0.0312f
C3348 R0.n0 GND 0.109f
C3349 R0.n4 GND 0.011f
C3350 R0.n5 GND 0.0121f
C3351 R0.n11 GND 0.0113f
C3352 R0.n24 GND 0.0141f
C3353 R0.n33 GND 0.425f
C3354 R0.t11 GND 0.0104f
C3355 R0.n34 GND 0.215f
C3356 R0.t9 GND 0.0312f
C3357 R0.n38 GND 0.0288f
C3358 R0.n41 GND 0.0127f
C3359 R0.n42 GND 0.0859f
C3360 R0.n43 GND 0.447f
C3361 R0.n44 GND 0.157f
C3362 R0.t1 GND 0.0122f
C3363 R0.n45 GND 0.0113f
C3364 R0.n46 GND 0.311f
C3365 R0.n47 GND 0.216f
C3366 VIN.t3 GND 0.0561f
C3367 VIN.n0 GND 0.453f
C3368 VIN.n1 GND 0.127f
C3369 VIN.t17 GND 0.0561f
C3370 VIN.n3 GND 0.45f
C3371 VIN.n4 GND 5.68f
C3372 VIN.t22 GND 0.0561f
C3373 VIN.n5 GND 0.453f
C3374 VIN.t8 GND 0.0561f
C3375 VIN.n6 GND 0.45f
C3376 VIN.t14 GND 0.0561f
C3377 VIN.n7 GND 0.453f
C3378 VIN.t29 GND 0.0561f
C3379 VIN.n8 GND 0.453f
C3380 VIN.t2 GND 0.0561f
C3381 VIN.n9 GND 0.453f
C3382 VIN.t9 GND 0.0561f
C3383 VIN.n10 GND 0.453f
C3384 VIN.t27 GND 0.0561f
C3385 VIN.n11 GND 0.453f
C3386 VIN.t30 GND 0.0561f
C3387 VIN.n12 GND 0.453f
C3388 VIN.t21 GND 0.0561f
C3389 VIN.n13 GND 0.453f
C3390 VIN.t25 GND 0.0561f
C3391 VIN.n14 GND 0.453f
C3392 VIN.t12 GND 0.0561f
C3393 VIN.n15 GND 0.453f
C3394 VIN.t18 GND 0.0561f
C3395 VIN.n16 GND 0.453f
C3396 VIN.t0 GND 0.0561f
C3397 VIN.n17 GND 0.453f
C3398 VIN.t7 GND 0.0561f
C3399 VIN.n18 GND 0.453f
C3400 VIN.n19 GND 11.9f
C3401 VIN.n20 GND 7.41f
C3402 VIN.n21 GND 7.41f
C3403 VIN.n22 GND 7.41f
C3404 VIN.n23 GND 7.41f
C3405 VIN.n24 GND 7.41f
C3406 VIN.n25 GND 7.42f
C3407 VIN.n26 GND 7.41f
C3408 VIN.n27 GND 7.41f
C3409 VIN.n28 GND 7.41f
C3410 VIN.n29 GND 7.41f
C3411 VIN.n30 GND 7.38f
C3412 VIN.n31 GND 7.41f
C3413 VIN.n32 GND 7.49f
C3414 VIN.n33 GND 1.18f
C3415 VV13.t17 GND 0.024f
C3416 VV13.n0 GND 0.196f
C3417 VV13.n1 GND 0.095f
C3418 VV13.t0 GND 0.313f
C3419 VV13.t1 GND 0.313f
C3420 VV13.t14 GND 0.313f
C3421 VV13.t5 GND 0.313f
C3422 VV13.t8 GND 0.313f
C3423 VV13.t12 GND 0.313f
C3424 VV13.t9 GND 0.313f
C3425 VV13.t11 GND 0.313f
C3426 VV13.t13 GND 0.313f
C3427 VV13.t6 GND 0.313f
C3428 VV13.t2 GND 0.313f
C3429 VV13.t3 GND 0.313f
C3430 VV13.t10 GND 0.313f
C3431 VV13.t4 GND 0.313f
C3432 VV13.t7 GND 0.313f
C3433 VV13.t15 GND 0.313f
C3434 VV13.n2 GND 0.75f
C3435 VV13.n3 GND 0.77f
C3436 VV13.n4 GND 0.77f
C3437 VV13.n5 GND 0.77f
C3438 VV13.n6 GND 0.77f
C3439 VV13.n7 GND 0.77f
C3440 VV13.n8 GND 0.77f
C3441 VV13.n9 GND 0.684f
C3442 VV13.n10 GND 2.26f
C3443 VV14.t16 GND 0.0249f
C3444 VV14.n0 GND 0.204f
C3445 VV14.n1 GND 0.0945f
C3446 VV14.t0 GND 0.326f
C3447 VV14.t9 GND 0.326f
C3448 VV14.t7 GND 0.326f
C3449 VV14.t3 GND 0.326f
C3450 VV14.t11 GND 0.326f
C3451 VV14.t4 GND 0.326f
C3452 VV14.t10 GND 0.326f
C3453 VV14.t5 GND 0.326f
C3454 VV14.t8 GND 0.326f
C3455 VV14.t13 GND 0.326f
C3456 VV14.t2 GND 0.326f
C3457 VV14.t12 GND 0.326f
C3458 VV14.t6 GND 0.326f
C3459 VV14.t15 GND 0.326f
C3460 VV14.t14 GND 0.326f
C3461 VV14.t1 GND 0.326f
C3462 VV14.n2 GND 0.781f
C3463 VV14.n3 GND 0.801f
C3464 VV14.n4 GND 0.801f
C3465 VV14.n5 GND 0.801f
C3466 VV14.n6 GND 0.801f
C3467 VV14.n7 GND 0.801f
C3468 VV14.n8 GND 0.801f
C3469 VV14.n9 GND 0.719f
C3470 VV14.n10 GND 2.51f
C3471 frontAnalog_v0p0p1_10.IB.n0 GND 0.0726f
C3472 frontAnalog_v0p0p1_10.IB.t12 GND 0.0832f
C3473 frontAnalog_v0p0p1_10.IB.t23 GND 0.0823f
C3474 frontAnalog_v0p0p1_10.IB.t3 GND 0.0832f
C3475 frontAnalog_v0p0p1_10.IB.t11 GND 0.0823f
C3476 frontAnalog_v0p0p1_10.IB.n3 GND 8.18f
C3477 frontAnalog_v0p0p1_10.IB.t32 GND 0.0832f
C3478 frontAnalog_v0p0p1_10.IB.t9 GND 0.0823f
C3479 frontAnalog_v0p0p1_10.IB.t5 GND 0.0832f
C3480 frontAnalog_v0p0p1_10.IB.t29 GND 0.0823f
C3481 frontAnalog_v0p0p1_10.IB.t22 GND 0.0832f
C3482 frontAnalog_v0p0p1_10.IB.t34 GND 0.0823f
C3483 frontAnalog_v0p0p1_10.IB.t26 GND 0.0832f
C3484 frontAnalog_v0p0p1_10.IB.t19 GND 0.0823f
C3485 frontAnalog_v0p0p1_10.IB.t15 GND 0.0832f
C3486 frontAnalog_v0p0p1_10.IB.t25 GND 0.0823f
C3487 frontAnalog_v0p0p1_10.IB.t18 GND 0.0832f
C3488 frontAnalog_v0p0p1_10.IB.t30 GND 0.0823f
C3489 frontAnalog_v0p0p1_10.IB.t7 GND 0.0832f
C3490 frontAnalog_v0p0p1_10.IB.t16 GND 0.0823f
C3491 frontAnalog_v0p0p1_10.IB.t10 GND 0.0832f
C3492 frontAnalog_v0p0p1_10.IB.t20 GND 0.0823f
C3493 frontAnalog_v0p0p1_10.IB.t31 GND 0.0832f
C3494 frontAnalog_v0p0p1_10.IB.t8 GND 0.0823f
C3495 frontAnalog_v0p0p1_10.IB.t4 GND 0.0832f
C3496 frontAnalog_v0p0p1_10.IB.t13 GND 0.0823f
C3497 frontAnalog_v0p0p1_10.IB.t21 GND 0.0832f
C3498 frontAnalog_v0p0p1_10.IB.t33 GND 0.0823f
C3499 frontAnalog_v0p0p1_10.IB.t27 GND 0.0832f
C3500 frontAnalog_v0p0p1_10.IB.t6 GND 0.0823f
C3501 frontAnalog_v0p0p1_10.IB.t14 GND 0.0832f
C3502 frontAnalog_v0p0p1_10.IB.t24 GND 0.0823f
C3503 frontAnalog_v0p0p1_10.IB.t17 GND 0.0832f
C3504 frontAnalog_v0p0p1_10.IB.t28 GND 0.0823f
C3505 frontAnalog_v0p0p1_10.IB.n18 GND 12.2f
C3506 frontAnalog_v0p0p1_10.IB.n19 GND 8.47f
C3507 frontAnalog_v0p0p1_10.IB.n20 GND 8.42f
C3508 frontAnalog_v0p0p1_10.IB.n21 GND 8.53f
C3509 frontAnalog_v0p0p1_10.IB.n22 GND 8.42f
C3510 frontAnalog_v0p0p1_10.IB.n23 GND 8.48f
C3511 frontAnalog_v0p0p1_10.IB.n24 GND 8.43f
C3512 frontAnalog_v0p0p1_10.IB.n25 GND 8.47f
C3513 frontAnalog_v0p0p1_10.IB.n26 GND 8.42f
C3514 frontAnalog_v0p0p1_10.IB.n27 GND 8.43f
C3515 frontAnalog_v0p0p1_10.IB.n28 GND 8.48f
C3516 frontAnalog_v0p0p1_10.IB.n29 GND 8.53f
C3517 frontAnalog_v0p0p1_10.IB.n30 GND 7.05f
C3518 frontAnalog_v0p0p1_10.IB.n31 GND 14.7f
C3519 frontAnalog_v0p0p1_10.IB.t1 GND 0.0463f
C3520 frontAnalog_v0p0p1_10.IB.n32 GND 0.124f
C3521 frontAnalog_v0p0p1_10.IB.n33 GND 0.0147f
C3522 frontAnalog_v0p0p1_10.IB.t0 GND 0.634f
C3523 frontAnalog_v0p0p1_10.IB.n34 GND 10.9f
C3524 I13.n0 GND 0.0101f
C3525 I13.n8 GND 0.113f
C3526 I13.n9 GND 0.263f
C3527 I13.n16 GND 0.16f
C3528 I13.n21 GND 0.425f
C3529 I13.n22 GND 1.01f
C3530 I13.n23 GND 0.47f
C3531 I13.n24 GND 0.282f
C3532 I13.n25 GND 0.501f
C3533 I13.n26 GND 0.153f
C3534 I13.n27 GND 0.407f
C3535 I13.n28 GND 0.585f
C3536 I13.t12 GND 0.0207f
C3537 I13.n29 GND 0.325f
C3538 I13.n30 GND 0.043f
C3539 I13.n31 GND 0.0975f
C3540 I13.n32 GND 0.0647f
C3541 I13.n33 GND 0.0691f
C3542 I13.n34 GND 0.0953f
C3543 I13.n35 GND 0.0902f
C3544 I13.n36 GND 0.217f
C3545 I13.n37 GND 14f
C3546 frontAnalog_v0p0p1_6.RSfetsym_0.QN.n0 GND 1.01f
C3547 frontAnalog_v0p0p1_6.RSfetsym_0.QN.t6 GND 0.0321f
C3548 frontAnalog_v0p0p1_6.RSfetsym_0.QN.t5 GND 0.0947f
C3549 frontAnalog_v0p0p1_6.RSfetsym_0.QN.n1 GND 1.49f
C3550 frontAnalog_v0p0p1_6.RSfetsym_0.QN.n2 GND 0.595f
C3551 frontAnalog_v0p0p1_6.RSfetsym_0.QN.t3 GND 0.0368f
C3552 frontAnalog_v0p0p1_6.RSfetsym_0.QN.n3 GND 0.631f
C3553 frontAnalog_v0p0p1_6.RSfetsym_0.QN.t0 GND 0.0322f
C3554 frontAnalog_v0p0p1_6.RSfetsym_0.QN.t1 GND 0.0322f
C3555 frontAnalog_v0p0p1_6.RSfetsym_0.QN.t4 GND 0.0566f
C3556 I10.n0 GND 0.0159f
C3557 I10.n1 GND 0.115f
C3558 I10.n2 GND 0.234f
C3559 I10.n3 GND 0.0102f
C3560 I10.n4 GND 0.0106f
C3561 I10.n5 GND 0.582f
C3562 I10.n6 GND 0.0182f
C3563 I10.n7 GND 0.0846f
C3564 I10.n8 GND 1.42f
C3565 I10.n9 GND 1.7f
C3566 I10.t7 GND 0.0105f
C3567 I10.t5 GND 0.0321f
C3568 I10.n10 GND 0.503f
C3569 I10.n11 GND 0.0666f
C3570 I10.t0 GND 0.0108f
C3571 I10.n12 GND 0.151f
C3572 I10.n13 GND 0.1f
C3573 I10.n14 GND 0.107f
C3574 I10.t2 GND 0.0108f
C3575 I10.t3 GND 0.0108f
C3576 I10.n15 GND 0.148f
C3577 I10.n16 GND 0.14f
C3578 I10.t4 GND 0.0118f
C3579 I10.n17 GND 0.336f
C3580 I10.n18 GND 9.3f
C3581 I10.n19 GND 3.68f
C3582 frontAnalog_v0p0p1_15.RSfetsym_0.QN.n0 GND 1.01f
C3583 frontAnalog_v0p0p1_15.RSfetsym_0.QN.t6 GND 0.0321f
C3584 frontAnalog_v0p0p1_15.RSfetsym_0.QN.t5 GND 0.0947f
C3585 frontAnalog_v0p0p1_15.RSfetsym_0.QN.n1 GND 1.49f
C3586 frontAnalog_v0p0p1_15.RSfetsym_0.QN.n2 GND 0.595f
C3587 frontAnalog_v0p0p1_15.RSfetsym_0.QN.t1 GND 0.0368f
C3588 frontAnalog_v0p0p1_15.RSfetsym_0.QN.n3 GND 0.631f
C3589 frontAnalog_v0p0p1_15.RSfetsym_0.QN.t4 GND 0.0322f
C3590 frontAnalog_v0p0p1_15.RSfetsym_0.QN.t3 GND 0.0322f
C3591 frontAnalog_v0p0p1_15.RSfetsym_0.QN.t0 GND 0.0566f
C3592 S0.t1 GND 0.0214f
C3593 S0.t0 GND 0.0152f
C3594 S0.n1 GND 0.0168f
C3595 S0.n2 GND 0.419f
C3596 S0.n3 GND 0.461f
C3597 S0.n4 GND 0.134f
C3598 S0.t8 GND 0.0542f
C3599 S0.n5 GND 0.181f
C3600 S0.n6 GND 0.0118f
C3601 S0.n7 GND 0.0133f
C3602 S0.t10 GND 0.0146f
C3603 S0.t11 GND 0.0146f
C3604 S0.n11 GND 0.0244f
C3605 S0.n14 GND 0.0191f
C3606 S0.n16 GND 0.0118f
C3607 S0.t6 GND 0.0146f
C3608 S0.n17 GND 0.021f
C3609 S0.t5 GND 0.0146f
C3610 S0.n18 GND 0.0196f
C3611 S0.n22 GND 0.0185f
C3612 S0.n26 GND 0.012f
C3613 S0.n31 GND 0.016f
C3614 S0.n32 GND 0.0135f
C3615 S0.n37 GND 0.0143f
C3616 S0.n38 GND 0.784f
C3617 S0.t12 GND 0.0197f
C3618 S0.t2 GND 0.0541f
C3619 S0.n39 GND 0.227f
C3620 S0.n40 GND 0.556f
C3621 S0.n41 GND 0.804f
C3622 S0.n42 GND 0.377f
C3623 S0.n43 GND 0.372f
C3624 frontAnalog_v0p0p1_2.x65.A.n0 GND 0.139f
C3625 frontAnalog_v0p0p1_2.x65.A.t4 GND 0.028f
C3626 frontAnalog_v0p0p1_2.x65.A.t5 GND 0.0175f
C3627 frontAnalog_v0p0p1_2.x65.A.n1 GND 0.0568f
C3628 frontAnalog_v0p0p1_2.x65.A.t1 GND 0.149f
C3629 frontAnalog_v0p0p1_2.x65.A.t2 GND 0.463f
C3630 frontAnalog_v0p0p1_2.x65.A.t3 GND 0.0194f
C3631 frontAnalog_v0p0p1_2.x65.A.n2 GND 1.6f
C3632 frontAnalog_v0p0p1_2.x65.A.t6 GND 0.0318f
C3633 frontAnalog_v0p0p1_2.x65.A.t0 GND 0.141f
C3634 frontAnalog_v0p0p1_2.x65.A.t7 GND 0.219f
C3635 frontAnalog_v0p0p1_2.x65.A.n3 GND 1.37f
C3636 frontAnalog_v0p0p1_2.x65.A.n4 GND 0.898f
C3637 frontAnalog_v0p0p1_2.x65.A.n5 GND 2.01f
C3638 frontAnalog_v0p0p1_2.x65.A.n6 GND 1.72f
C3639 frontAnalog_v0p0p1_2.x63.A.n0 GND 0.12f
C3640 frontAnalog_v0p0p1_2.x63.A.n1 GND 2.22f
C3641 frontAnalog_v0p0p1_2.x63.A.t6 GND 0.014f
C3642 frontAnalog_v0p0p1_2.x63.A.t5 GND 0.0225f
C3643 frontAnalog_v0p0p1_2.x63.A.n2 GND 0.0465f
C3644 frontAnalog_v0p0p1_2.x63.A.t2 GND 0.151f
C3645 frontAnalog_v0p0p1_2.x63.A.t4 GND 0.0256f
C3646 frontAnalog_v0p0p1_2.x63.A.t3 GND 0.173f
C3647 frontAnalog_v0p0p1_2.x63.A.t7 GND 0.175f
C3648 frontAnalog_v0p0p1_2.x63.A.n3 GND 1f
C3649 frontAnalog_v0p0p1_2.x63.A.n4 GND 0.953f
C3650 frontAnalog_v0p0p1_2.x63.A.t0 GND 0.0156f
C3651 frontAnalog_v0p0p1_2.x63.A.t1 GND 0.334f
C3652 frontAnalog_v0p0p1_2.x63.A.n5 GND 1.25f
C3653 VV15.t17 GND 0.0258f
C3654 VV15.n0 GND 0.212f
C3655 VV15.n1 GND 0.0979f
C3656 VV15.t10 GND 0.338f
C3657 VV15.t14 GND 0.338f
C3658 VV15.t4 GND 0.338f
C3659 VV15.t12 GND 0.338f
C3660 VV15.t5 GND 0.338f
C3661 VV15.t8 GND 0.338f
C3662 VV15.t6 GND 0.338f
C3663 VV15.t3 GND 0.338f
C3664 VV15.t13 GND 0.338f
C3665 VV15.t0 GND 0.338f
C3666 VV15.t11 GND 0.338f
C3667 VV15.t2 GND 0.338f
C3668 VV15.t15 GND 0.338f
C3669 VV15.t9 GND 0.338f
C3670 VV15.t1 GND 0.338f
C3671 VV15.t7 GND 0.338f
C3672 VV15.n2 GND 0.808f
C3673 VV15.n3 GND 0.829f
C3674 VV15.n4 GND 0.829f
C3675 VV15.n5 GND 0.829f
C3676 VV15.n6 GND 0.829f
C3677 VV15.n7 GND 0.829f
C3678 VV15.n8 GND 0.829f
C3679 VV15.n9 GND 0.74f
C3680 VV9.t16 GND 0.0231f
C3681 VV9.n0 GND 0.189f
C3682 VV9.n1 GND 0.0915f
C3683 VV9.t15 GND 0.302f
C3684 VV9.t5 GND 0.302f
C3685 VV9.t13 GND 0.302f
C3686 VV9.t11 GND 0.302f
C3687 VV9.t9 GND 0.302f
C3688 VV9.t2 GND 0.302f
C3689 VV9.t12 GND 0.302f
C3690 VV9.t6 GND 0.302f
C3691 VV9.t4 GND 0.302f
C3692 VV9.t14 GND 0.302f
C3693 VV9.t3 GND 0.302f
C3694 VV9.t1 GND 0.302f
C3695 VV9.t0 GND 0.302f
C3696 VV9.t7 GND 0.302f
C3697 VV9.t8 GND 0.302f
C3698 VV9.t10 GND 0.302f
C3699 VV9.n2 GND 0.723f
C3700 VV9.n3 GND 0.742f
C3701 VV9.n4 GND 0.742f
C3702 VV9.n5 GND 0.742f
C3703 VV9.n6 GND 0.742f
C3704 VV9.n7 GND 0.742f
C3705 VV9.n8 GND 0.742f
C3706 VV9.n9 GND 0.666f
C3707 VV9.n10 GND 1.69f
C3708 frontAnalog_v0p0p1_8.RSfetsym_0.QN.n0 GND 1.01f
C3709 frontAnalog_v0p0p1_8.RSfetsym_0.QN.t5 GND 0.0321f
C3710 frontAnalog_v0p0p1_8.RSfetsym_0.QN.t6 GND 0.0947f
C3711 frontAnalog_v0p0p1_8.RSfetsym_0.QN.n1 GND 1.49f
C3712 frontAnalog_v0p0p1_8.RSfetsym_0.QN.n2 GND 0.595f
C3713 frontAnalog_v0p0p1_8.RSfetsym_0.QN.t0 GND 0.0368f
C3714 frontAnalog_v0p0p1_8.RSfetsym_0.QN.n3 GND 0.631f
C3715 frontAnalog_v0p0p1_8.RSfetsym_0.QN.t2 GND 0.0322f
C3716 frontAnalog_v0p0p1_8.RSfetsym_0.QN.t3 GND 0.0322f
C3717 frontAnalog_v0p0p1_8.RSfetsym_0.QN.t1 GND 0.0566f
C3718 OUT1.n2 GND 0.0114f
C3719 OUT1.n4 GND 0.0242f
C3720 OUT1.n6 GND 0.0161f
C3721 OUT1.n8 GND 0.0161f
C3722 OUT1.n10 GND 0.0161f
C3723 OUT1.n12 GND 0.0161f
C3724 OUT1.n14 GND 0.0161f
C3725 OUT1.n23 GND 0.014f
C3726 OUT1.n25 GND 0.0348f
C3727 OUT1.n27 GND 0.021f
C3728 OUT1.n29 GND 0.021f
C3729 OUT1.n31 GND 0.021f
C3730 OUT1.n33 GND 0.021f
C3731 OUT1.n35 GND 0.021f
C3732 OUT1.n37 GND 0.0147f
C3733 OUT1.n38 GND 0.0297f
C3734 OUT1.n39 GND 0.0229f
C3735 OUT1.n42 GND 0.0114f
C3736 OUT1.n44 GND 0.0242f
C3737 OUT1.n46 GND 0.0161f
C3738 OUT1.n48 GND 0.0161f
C3739 OUT1.n50 GND 0.0161f
C3740 OUT1.n52 GND 0.0161f
C3741 OUT1.n54 GND 0.0161f
C3742 OUT1.n63 GND 0.014f
C3743 OUT1.n65 GND 0.0348f
C3744 OUT1.n67 GND 0.021f
C3745 OUT1.n69 GND 0.021f
C3746 OUT1.n71 GND 0.021f
C3747 OUT1.n73 GND 0.021f
C3748 OUT1.n75 GND 0.021f
C3749 OUT1.n77 GND 0.0147f
C3750 OUT1.n78 GND 0.0274f
C3751 OUT1.n79 GND 0.0203f
C3752 OUT1.n81 GND 0.0114f
C3753 OUT1.n83 GND 0.0242f
C3754 OUT1.n85 GND 0.0161f
C3755 OUT1.n87 GND 0.0161f
C3756 OUT1.n89 GND 0.0161f
C3757 OUT1.n91 GND 0.0161f
C3758 OUT1.n93 GND 0.0161f
C3759 OUT1.n97 GND 0.0126f
C3760 OUT1.n100 GND 0.014f
C3761 OUT1.n102 GND 0.0348f
C3762 OUT1.n104 GND 0.021f
C3763 OUT1.n106 GND 0.021f
C3764 OUT1.n108 GND 0.021f
C3765 OUT1.n110 GND 0.021f
C3766 OUT1.n112 GND 0.021f
C3767 OUT1.n114 GND 0.0147f
C3768 OUT1.n115 GND 0.0284f
C3769 OUT1.n116 GND 0.0234f
C3770 OUT1.n120 GND 0.014f
C3771 OUT1.n122 GND 0.0348f
C3772 OUT1.n124 GND 0.021f
C3773 OUT1.n126 GND 0.021f
C3774 OUT1.n128 GND 0.021f
C3775 OUT1.n130 GND 0.021f
C3776 OUT1.n132 GND 0.021f
C3777 OUT1.n136 GND 0.0114f
C3778 OUT1.n138 GND 0.0242f
C3779 OUT1.n140 GND 0.0161f
C3780 OUT1.n142 GND 0.0161f
C3781 OUT1.n144 GND 0.0161f
C3782 OUT1.n146 GND 0.0161f
C3783 OUT1.n148 GND 0.0161f
C3784 OUT1.n152 GND 0.0129f
C3785 OUT1.n155 GND 0.0204f
C3786 OUT1.n156 GND 0.108f
C3787 OUT1.n157 GND 0.275f
C3788 OUT1.n158 GND 0.224f
C3789 OUT1.n159 GND 0.228f
C3790 I2.n1 GND 0.0619f
C3791 I2.n2 GND 0.126f
C3792 I2.n5 GND 0.321f
C3793 I2.n7 GND 0.0436f
C3794 I2.n8 GND 0.762f
C3795 I2.n9 GND 0.536f
C3796 I2.t10 GND 0.0173f
C3797 I2.n10 GND 0.271f
C3798 I2.n11 GND 0.0359f
C3799 I2.n12 GND 0.0814f
C3800 I2.n13 GND 0.054f
C3801 I2.n14 GND 0.0577f
C3802 I2.n15 GND 0.0795f
C3803 I2.n16 GND 0.0752f
C3804 I2.n17 GND 0.173f
C3805 I2.n18 GND 11.8f
C3806 I2.n19 GND 0.84f
C3807 R1.t4 GND 0.0309f
C3808 R1.n0 GND 0.108f
C3809 R1.n4 GND 0.0109f
C3810 R1.n5 GND 0.012f
C3811 R1.n11 GND 0.0112f
C3812 R1.n24 GND 0.0139f
C3813 R1.n33 GND 0.421f
C3814 R1.t10 GND 0.0103f
C3815 R1.n34 GND 0.213f
C3816 R1.t8 GND 0.0309f
C3817 R1.n38 GND 0.0285f
C3818 R1.n41 GND 0.0125f
C3819 R1.n42 GND 0.0851f
C3820 R1.n43 GND 0.442f
C3821 R1.n44 GND 0.155f
C3822 R1.t1 GND 0.0121f
C3823 R1.n45 GND 0.0112f
C3824 R1.n46 GND 0.276f
C3825 R1.n47 GND 0.225f
C3826 I0.n1 GND 0.0918f
C3827 I0.n2 GND 0.245f
C3828 I0.n3 GND 0.301f
C3829 I0.n4 GND 0.142f
C3830 I0.n5 GND 0.0187f
C3831 I0.n6 GND 0.0425f
C3832 I0.n7 GND 0.0282f
C3833 I0.n8 GND 0.0301f
C3834 I0.n9 GND 0.0415f
C3835 I0.n10 GND 0.0393f
C3836 I0.n11 GND 0.0905f
C3837 I0.n12 GND 7.99f
C3838 I0.n13 GND 0.256f
C3839 VV1.t16 GND 0.0127f
C3840 VV1.n0 GND 0.104f
C3841 VV1.n1 GND 0.0503f
C3842 VV1.t2 GND 0.166f
C3843 VV1.t8 GND 0.166f
C3844 VV1.t11 GND 0.166f
C3845 VV1.t3 GND 0.166f
C3846 VV1.t15 GND 0.166f
C3847 VV1.t9 GND 0.166f
C3848 VV1.t12 GND 0.166f
C3849 VV1.t14 GND 0.166f
C3850 VV1.t0 GND 0.166f
C3851 VV1.t5 GND 0.166f
C3852 VV1.t13 GND 0.166f
C3853 VV1.t6 GND 0.166f
C3854 VV1.t10 GND 0.166f
C3855 VV1.t1 GND 0.166f
C3856 VV1.t4 GND 0.166f
C3857 VV1.t7 GND 0.166f
C3858 VV1.n2 GND 0.398f
C3859 VV1.n3 GND 0.408f
C3860 VV1.n4 GND 0.408f
C3861 VV1.n5 GND 0.408f
C3862 VV1.n6 GND 0.408f
C3863 VV1.n7 GND 0.408f
C3864 VV1.n8 GND 0.408f
C3865 VV1.n9 GND 0.361f
C3866 VV1.n10 GND 1.18f
C3867 VV2.t17 GND 0.023f
C3868 VV2.n0 GND 0.188f
C3869 VV2.n1 GND 0.0951f
C3870 VV2.t7 GND 0.301f
C3871 VV2.t5 GND 0.301f
C3872 VV2.t9 GND 0.301f
C3873 VV2.t12 GND 0.301f
C3874 VV2.t3 GND 0.301f
C3875 VV2.t15 GND 0.301f
C3876 VV2.t8 GND 0.301f
C3877 VV2.t13 GND 0.301f
C3878 VV2.t4 GND 0.301f
C3879 VV2.t2 GND 0.301f
C3880 VV2.t0 GND 0.301f
C3881 VV2.t14 GND 0.301f
C3882 VV2.t1 GND 0.301f
C3883 VV2.t11 GND 0.301f
C3884 VV2.t10 GND 0.648f
C3885 VV2.t6 GND 0.301f
C3886 VV2.n2 GND 0.372f
C3887 VV2.n3 GND 0.369f
C3888 VV2.n4 GND 0.369f
C3889 VV2.n5 GND 0.369f
C3890 VV2.n6 GND 0.369f
C3891 VV2.n7 GND 0.369f
C3892 VV2.n8 GND 0.369f
C3893 VV2.n9 GND 0.369f
C3894 VV2.n10 GND 0.369f
C3895 VV2.n11 GND 0.369f
C3896 VV2.n12 GND 0.369f
C3897 VV2.n13 GND 0.369f
C3898 VV2.n14 GND 0.369f
C3899 VV2.n15 GND 0.369f
C3900 VV2.n16 GND 0.283f
C3901 VV2.n17 GND 2.34f
C3902 VV10.t17 GND 0.0223f
C3903 VV10.n0 GND 0.183f
C3904 VV10.n1 GND 0.0923f
C3905 VV10.t5 GND 0.292f
C3906 VV10.t2 GND 0.292f
C3907 VV10.t9 GND 0.292f
C3908 VV10.t12 GND 0.292f
C3909 VV10.t4 GND 0.292f
C3910 VV10.t14 GND 0.292f
C3911 VV10.t6 GND 0.292f
C3912 VV10.t3 GND 0.292f
C3913 VV10.t13 GND 0.292f
C3914 VV10.t1 GND 0.292f
C3915 VV10.t0 GND 0.292f
C3916 VV10.t15 GND 0.292f
C3917 VV10.t7 GND 0.292f
C3918 VV10.t11 GND 0.292f
C3919 VV10.t8 GND 0.292f
C3920 VV10.t10 GND 0.292f
C3921 VV10.n2 GND 0.699f
C3922 VV10.n3 GND 0.717f
C3923 VV10.n4 GND 0.717f
C3924 VV10.n5 GND 0.717f
C3925 VV10.n6 GND 0.717f
C3926 VV10.n7 GND 0.717f
C3927 VV10.n8 GND 0.717f
C3928 VV10.n9 GND 0.648f
C3929 VV10.n10 GND 1.67f
C3930 VV11.t16 GND 0.0237f
C3931 VV11.n0 GND 0.194f
C3932 VV11.n1 GND 0.0938f
C3933 VV11.t1 GND 0.309f
C3934 VV11.t3 GND 0.309f
C3935 VV11.t14 GND 0.309f
C3936 VV11.t11 GND 0.309f
C3937 VV11.t5 GND 0.309f
C3938 VV11.t13 GND 0.309f
C3939 VV11.t8 GND 0.309f
C3940 VV11.t6 GND 0.309f
C3941 VV11.t4 GND 0.309f
C3942 VV11.t2 GND 0.309f
C3943 VV11.t0 GND 0.309f
C3944 VV11.t15 GND 0.309f
C3945 VV11.t12 GND 0.309f
C3946 VV11.t10 GND 0.309f
C3947 VV11.t7 GND 0.309f
C3948 VV11.t9 GND 0.666f
C3949 VV11.n2 GND 0.383f
C3950 VV11.n3 GND 0.38f
C3951 VV11.n4 GND 0.38f
C3952 VV11.n5 GND 0.38f
C3953 VV11.n6 GND 0.38f
C3954 VV11.n7 GND 0.38f
C3955 VV11.n8 GND 0.38f
C3956 VV11.n9 GND 0.38f
C3957 VV11.n10 GND 0.38f
C3958 VV11.n11 GND 0.38f
C3959 VV11.n12 GND 0.38f
C3960 VV11.n13 GND 0.38f
C3961 VV11.n14 GND 0.38f
C3962 VV11.n15 GND 0.38f
C3963 VV11.n16 GND 0.307f
C3964 VV11.n17 GND 1.93f
C3965 frontAnalog_v0p0p1_5.RSfetsym_0.QN.n0 GND 1.01f
C3966 frontAnalog_v0p0p1_5.RSfetsym_0.QN.t6 GND 0.0321f
C3967 frontAnalog_v0p0p1_5.RSfetsym_0.QN.t5 GND 0.0947f
C3968 frontAnalog_v0p0p1_5.RSfetsym_0.QN.n1 GND 1.49f
C3969 frontAnalog_v0p0p1_5.RSfetsym_0.QN.n2 GND 0.595f
C3970 frontAnalog_v0p0p1_5.RSfetsym_0.QN.t1 GND 0.0368f
C3971 frontAnalog_v0p0p1_5.RSfetsym_0.QN.n3 GND 0.631f
C3972 frontAnalog_v0p0p1_5.RSfetsym_0.QN.t4 GND 0.0322f
C3973 frontAnalog_v0p0p1_5.RSfetsym_0.QN.t3 GND 0.0322f
C3974 frontAnalog_v0p0p1_5.RSfetsym_0.QN.t0 GND 0.0566f
C3975 frontAnalog_v0p0p1_14.x65.A.n0 GND 0.139f
C3976 frontAnalog_v0p0p1_14.x65.A.t7 GND 0.028f
C3977 frontAnalog_v0p0p1_14.x65.A.t4 GND 0.0175f
C3978 frontAnalog_v0p0p1_14.x65.A.n1 GND 0.0568f
C3979 frontAnalog_v0p0p1_14.x65.A.t5 GND 0.0318f
C3980 frontAnalog_v0p0p1_14.x65.A.t1 GND 0.141f
C3981 frontAnalog_v0p0p1_14.x65.A.t6 GND 0.219f
C3982 frontAnalog_v0p0p1_14.x65.A.n2 GND 1.37f
C3983 frontAnalog_v0p0p1_14.x65.A.n3 GND 0.898f
C3984 frontAnalog_v0p0p1_14.x65.A.t3 GND 0.463f
C3985 frontAnalog_v0p0p1_14.x65.A.t2 GND 0.0194f
C3986 frontAnalog_v0p0p1_14.x65.A.n4 GND 1.6f
C3987 frontAnalog_v0p0p1_14.x65.A.n5 GND 2.01f
C3988 frontAnalog_v0p0p1_14.x65.A.t0 GND 0.149f
C3989 frontAnalog_v0p0p1_14.x65.A.n6 GND 1.72f
C3990 frontAnalog_v0p0p1_14.x63.A.n0 GND 0.12f
C3991 frontAnalog_v0p0p1_14.x63.A.n1 GND 2.22f
C3992 frontAnalog_v0p0p1_14.x63.A.t5 GND 0.014f
C3993 frontAnalog_v0p0p1_14.x63.A.t7 GND 0.0225f
C3994 frontAnalog_v0p0p1_14.x63.A.n2 GND 0.0465f
C3995 frontAnalog_v0p0p1_14.x63.A.t4 GND 0.0256f
C3996 frontAnalog_v0p0p1_14.x63.A.t1 GND 0.173f
C3997 frontAnalog_v0p0p1_14.x63.A.t6 GND 0.175f
C3998 frontAnalog_v0p0p1_14.x63.A.n3 GND 1f
C3999 frontAnalog_v0p0p1_14.x63.A.n4 GND 0.953f
C4000 frontAnalog_v0p0p1_14.x63.A.t2 GND 0.0156f
C4001 frontAnalog_v0p0p1_14.x63.A.t3 GND 0.335f
C4002 frontAnalog_v0p0p1_14.x63.A.t0 GND 0.151f
C4003 frontAnalog_v0p0p1_14.x63.A.n5 GND 1.25f
C4004 VV3.t16 GND 0.0237f
C4005 VV3.n0 GND 0.194f
C4006 VV3.n1 GND 0.094f
C4007 VV3.t7 GND 0.31f
C4008 VV3.t11 GND 0.31f
C4009 VV3.t10 GND 0.31f
C4010 VV3.t3 GND 0.31f
C4011 VV3.t2 GND 0.31f
C4012 VV3.t12 GND 0.31f
C4013 VV3.t8 GND 0.31f
C4014 VV3.t9 GND 0.31f
C4015 VV3.t4 GND 0.31f
C4016 VV3.t15 GND 0.31f
C4017 VV3.t0 GND 0.31f
C4018 VV3.t5 GND 0.31f
C4019 VV3.t1 GND 0.31f
C4020 VV3.t14 GND 0.31f
C4021 VV3.t6 GND 0.31f
C4022 VV3.t13 GND 0.669f
C4023 VV3.n2 GND 0.384f
C4024 VV3.n3 GND 0.381f
C4025 VV3.n4 GND 0.381f
C4026 VV3.n5 GND 0.381f
C4027 VV3.n6 GND 0.381f
C4028 VV3.n7 GND 0.381f
C4029 VV3.n8 GND 0.381f
C4030 VV3.n9 GND 0.381f
C4031 VV3.n10 GND 0.381f
C4032 VV3.n11 GND 0.381f
C4033 VV3.n12 GND 0.381f
C4034 VV3.n13 GND 0.381f
C4035 VV3.n14 GND 0.381f
C4036 VV3.n15 GND 0.381f
C4037 VV3.n16 GND 0.301f
C4038 VV3.n17 GND 2.27f
C4039 VV4.t16 GND 0.0245f
C4040 VV4.n0 GND 0.201f
C4041 VV4.n1 GND 0.097f
C4042 VV4.t0 GND 0.32f
C4043 VV4.t10 GND 0.32f
C4044 VV4.t7 GND 0.32f
C4045 VV4.t3 GND 0.32f
C4046 VV4.t2 GND 0.32f
C4047 VV4.t11 GND 0.32f
C4048 VV4.t9 GND 0.32f
C4049 VV4.t6 GND 0.32f
C4050 VV4.t1 GND 0.32f
C4051 VV4.t15 GND 0.32f
C4052 VV4.t5 GND 0.32f
C4053 VV4.t4 GND 0.32f
C4054 VV4.t13 GND 0.32f
C4055 VV4.t14 GND 0.32f
C4056 VV4.t12 GND 0.32f
C4057 VV4.t8 GND 0.32f
C4058 VV4.n2 GND 0.766f
C4059 VV4.n3 GND 0.786f
C4060 VV4.n4 GND 0.786f
C4061 VV4.n5 GND 0.786f
C4062 VV4.n6 GND 0.786f
C4063 VV4.n7 GND 0.786f
C4064 VV4.n8 GND 0.786f
C4065 VV4.n9 GND 0.708f
C4066 VV4.n10 GND 2.21f
C4067 frontAnalog_v0p0p1_10.x65.A.n0 GND 0.139f
C4068 frontAnalog_v0p0p1_10.x65.A.t4 GND 0.028f
C4069 frontAnalog_v0p0p1_10.x65.A.t6 GND 0.0175f
C4070 frontAnalog_v0p0p1_10.x65.A.n1 GND 0.0568f
C4071 frontAnalog_v0p0p1_10.x65.A.t2 GND 0.149f
C4072 frontAnalog_v0p0p1_10.x65.A.t7 GND 0.0318f
C4073 frontAnalog_v0p0p1_10.x65.A.t3 GND 0.141f
C4074 frontAnalog_v0p0p1_10.x65.A.t5 GND 0.219f
C4075 frontAnalog_v0p0p1_10.x65.A.n2 GND 1.37f
C4076 frontAnalog_v0p0p1_10.x65.A.n3 GND 0.898f
C4077 frontAnalog_v0p0p1_10.x65.A.t0 GND 0.463f
C4078 frontAnalog_v0p0p1_10.x65.A.t1 GND 0.0194f
C4079 frontAnalog_v0p0p1_10.x65.A.n4 GND 1.6f
C4080 frontAnalog_v0p0p1_10.x65.A.n5 GND 2.01f
C4081 frontAnalog_v0p0p1_10.x65.A.n6 GND 1.72f
C4082 CLK.t23 GND 0.0562f
C4083 CLK.t89 GND 0.325f
C4084 CLK.t85 GND 0.329f
C4085 CLK.n1 GND 0.286f
C4086 CLK.t26 GND 0.0592f
C4087 CLK.n2 GND 0.463f
C4088 CLK.n4 GND 0.0676f
C4089 CLK.t94 GND 0.0942f
C4090 CLK.n5 GND 0.395f
C4091 CLK.n6 GND 0.36f
C4092 CLK.n7 GND 0.1f
C4093 CLK.n8 GND 14.1f
C4094 CLK.t58 GND 0.0562f
C4095 CLK.t63 GND 0.325f
C4096 CLK.t14 GND 0.329f
C4097 CLK.n10 GND 0.286f
C4098 CLK.t92 GND 0.0592f
C4099 CLK.n11 GND 0.463f
C4100 CLK.n13 GND 0.0676f
C4101 CLK.t15 GND 0.0942f
C4102 CLK.n14 GND 0.395f
C4103 CLK.n15 GND 0.36f
C4104 CLK.n16 GND 0.1f
C4105 CLK.t17 GND 0.0562f
C4106 CLK.t27 GND 0.325f
C4107 CLK.t73 GND 0.329f
C4108 CLK.n18 GND 0.286f
C4109 CLK.t11 GND 0.0592f
C4110 CLK.n19 GND 0.463f
C4111 CLK.n21 GND 0.0676f
C4112 CLK.t32 GND 0.0942f
C4113 CLK.n22 GND 0.395f
C4114 CLK.n23 GND 0.36f
C4115 CLK.n24 GND 0.1f
C4116 CLK.t35 GND 0.0562f
C4117 CLK.t38 GND 0.325f
C4118 CLK.t90 GND 0.329f
C4119 CLK.n26 GND 0.286f
C4120 CLK.t66 GND 0.0592f
C4121 CLK.n27 GND 0.463f
C4122 CLK.n29 GND 0.0676f
C4123 CLK.t91 GND 0.0942f
C4124 CLK.n30 GND 0.395f
C4125 CLK.n31 GND 0.36f
C4126 CLK.n32 GND 0.1f
C4127 CLK.t45 GND 0.0562f
C4128 CLK.t5 GND 0.325f
C4129 CLK.t47 GND 0.329f
C4130 CLK.n34 GND 0.286f
C4131 CLK.t83 GND 0.0592f
C4132 CLK.n35 GND 0.463f
C4133 CLK.n37 GND 0.0676f
C4134 CLK.t10 GND 0.0942f
C4135 CLK.n38 GND 0.395f
C4136 CLK.n39 GND 0.36f
C4137 CLK.n40 GND 0.104f
C4138 CLK.t4 GND 0.0562f
C4139 CLK.t18 GND 0.325f
C4140 CLK.t64 GND 0.329f
C4141 CLK.n42 GND 0.286f
C4142 CLK.t41 GND 0.0592f
C4143 CLK.n43 GND 0.463f
C4144 CLK.n45 GND 0.0676f
C4145 CLK.t65 GND 0.0942f
C4146 CLK.n46 GND 0.395f
C4147 CLK.n47 GND 0.36f
C4148 CLK.n48 GND 0.1f
C4149 CLK.t25 GND 0.0562f
C4150 CLK.t71 GND 0.325f
C4151 CLK.t74 GND 0.329f
C4152 CLK.n50 GND 0.286f
C4153 CLK.t54 GND 0.0592f
C4154 CLK.n51 GND 0.463f
C4155 CLK.n53 GND 0.0676f
C4156 CLK.t76 GND 0.0942f
C4157 CLK.n54 GND 0.395f
C4158 CLK.n55 GND 0.36f
C4159 CLK.n56 GND 0.1f
C4160 CLK.t79 GND 0.0562f
C4161 CLK.t95 GND 0.325f
C4162 CLK.t39 GND 0.329f
C4163 CLK.n58 GND 0.286f
C4164 CLK.t20 GND 0.0592f
C4165 CLK.n59 GND 0.463f
C4166 CLK.n61 GND 0.0676f
C4167 CLK.t40 GND 0.0942f
C4168 CLK.n62 GND 0.395f
C4169 CLK.n63 GND 0.36f
C4170 CLK.n64 GND 0.1f
C4171 CLK.t2 GND 0.0562f
C4172 CLK.t6 GND 0.325f
C4173 CLK.t51 GND 0.329f
C4174 CLK.n66 GND 0.286f
C4175 CLK.t30 GND 0.0592f
C4176 CLK.n67 GND 0.463f
C4177 CLK.n69 GND 0.0676f
C4178 CLK.t53 GND 0.0942f
C4179 CLK.n70 GND 0.395f
C4180 CLK.n71 GND 0.36f
C4181 CLK.n72 GND 0.1f
C4182 CLK.t56 GND 0.0562f
C4183 CLK.t70 GND 0.325f
C4184 CLK.t13 GND 0.329f
C4185 CLK.n74 GND 0.286f
C4186 CLK.t0 GND 0.0592f
C4187 CLK.n75 GND 0.463f
C4188 CLK.n77 GND 0.0676f
C4189 CLK.t19 GND 0.0942f
C4190 CLK.n78 GND 0.395f
C4191 CLK.n79 GND 0.36f
C4192 CLK.n80 GND 0.1f
C4193 CLK.t69 GND 0.0562f
C4194 CLK.t80 GND 0.325f
C4195 CLK.t28 GND 0.329f
C4196 CLK.n82 GND 0.286f
C4197 CLK.t9 GND 0.0592f
C4198 CLK.n83 GND 0.463f
C4199 CLK.n85 GND 0.0676f
C4200 CLK.t29 GND 0.0942f
C4201 CLK.n86 GND 0.395f
C4202 CLK.n87 GND 0.36f
C4203 CLK.n88 GND 0.1f
C4204 CLK.t33 GND 0.0562f
C4205 CLK.t36 GND 0.325f
C4206 CLK.t87 GND 0.329f
C4207 CLK.n90 GND 0.286f
C4208 CLK.t62 GND 0.0592f
C4209 CLK.n91 GND 0.463f
C4210 CLK.n93 GND 0.0676f
C4211 CLK.t88 GND 0.0942f
C4212 CLK.n94 GND 0.395f
C4213 CLK.n95 GND 0.36f
C4214 CLK.n96 GND 0.1f
C4215 CLK.t44 GND 0.0562f
C4216 CLK.t57 GND 0.325f
C4217 CLK.t7 GND 0.329f
C4218 CLK.n98 GND 0.286f
C4219 CLK.t82 GND 0.0592f
C4220 CLK.n99 GND 0.463f
C4221 CLK.n101 GND 0.0676f
C4222 CLK.t8 GND 0.0942f
C4223 CLK.n102 GND 0.395f
C4224 CLK.n103 GND 0.36f
C4225 CLK.n104 GND 0.1f
C4226 CLK.t12 GND 0.0562f
C4227 CLK.t16 GND 0.325f
C4228 CLK.t60 GND 0.329f
C4229 CLK.n106 GND 0.286f
C4230 CLK.t37 GND 0.0592f
C4231 CLK.n107 GND 0.463f
C4232 CLK.n109 GND 0.0676f
C4233 CLK.t61 GND 0.0942f
C4234 CLK.n110 GND 0.395f
C4235 CLK.n111 GND 0.36f
C4236 CLK.n112 GND 0.104f
C4237 CLK.t24 GND 0.0562f
C4238 CLK.t34 GND 0.325f
C4239 CLK.t72 GND 0.329f
C4240 CLK.n114 GND 0.286f
C4241 CLK.t59 GND 0.0592f
C4242 CLK.n115 GND 0.463f
C4243 CLK.n117 GND 0.0676f
C4244 CLK.t81 GND 0.0942f
C4245 CLK.n118 GND 0.395f
C4246 CLK.n119 GND 0.36f
C4247 CLK.n120 GND 0.104f
C4248 CLK.n121 GND 19.3f
C4249 CLK.n122 GND 12.7f
C4250 CLK.n123 GND 12.8f
C4251 CLK.n124 GND 12.8f
C4252 CLK.n125 GND 12.8f
C4253 CLK.n126 GND 12.7f
C4254 CLK.n127 GND 12.8f
C4255 CLK.n128 GND 12.8f
C4256 CLK.n129 GND 12.8f
C4257 CLK.n130 GND 12.7f
C4258 CLK.n131 GND 12.7f
C4259 CLK.n132 GND 12.8f
C4260 CLK.n133 GND 12.8f
C4261 CLK.n134 GND 12.8f
C4262 CLK.t78 GND 0.0562f
C4263 CLK.t46 GND 0.325f
C4264 CLK.t48 GND 0.329f
C4265 CLK.t86 GND 0.0592f
C4266 CLK.n135 GND 0.463f
C4267 CLK.n137 GND 0.286f
C4268 CLK.n139 GND 0.0676f
C4269 CLK.t49 GND 0.0942f
C4270 CLK.n140 GND 0.395f
C4271 CLK.n141 GND 0.36f
C4272 CLK.n142 GND 0.1f
C4273 a_16719_n13117.n0 GND 1.47f
C4274 a_16719_n13117.n1 GND 1.14f
C4275 a_16719_n13117.t8 GND 0.177f
C4276 a_16719_n13117.t18 GND 0.177f
C4277 a_16719_n13117.t22 GND 0.177f
C4278 a_16719_n13117.t11 GND 0.177f
C4279 a_16719_n13117.t16 GND 0.177f
C4280 a_16719_n13117.t5 GND 0.177f
C4281 a_16719_n13117.t20 GND 0.177f
C4282 a_16719_n13117.t14 GND 0.177f
C4283 a_16719_n13117.t7 GND 0.177f
C4284 a_16719_n13117.t15 GND 0.177f
C4285 a_16719_n13117.t4 GND 0.177f
C4286 a_16719_n13117.t19 GND 0.177f
C4287 a_16719_n13117.t12 GND 0.252f
C4288 a_16719_n13117.n2 GND 1.4f
C4289 a_16719_n13117.n3 GND 0.768f
C4290 a_16719_n13117.n4 GND 0.768f
C4291 a_16719_n13117.n5 GND 0.768f
C4292 a_16719_n13117.n6 GND 0.768f
C4293 a_16719_n13117.n7 GND 0.768f
C4294 a_16719_n13117.n8 GND 0.72f
C4295 a_16719_n13117.n9 GND 0.273f
C4296 a_16719_n13117.n10 GND 0.325f
C4297 a_16719_n13117.n11 GND 0.912f
C4298 a_16719_n13117.n12 GND 2.03f
C4299 a_16719_n13117.n13 GND 1.47f
C4300 a_16719_n13117.t1 GND 0.238f
C4301 a_16719_n13117.n14 GND 2.05f
C4302 a_16719_n13117.t24 GND 1.7f
C4303 a_16719_n13117.n15 GND 0.991f
C4304 a_16719_n13117.n16 GND 0.0433f
C4305 a_16719_n13117.n17 GND 0.426f
C4306 a_16719_n13117.t0 GND 1.7f
C4307 a_16719_n13117.t2 GND 0.0103f
C4308 a_16719_n13117.n18 GND 0.213f
C4309 a_16719_n13117.t25 GND 1.7f
C4310 a_16719_n13117.n19 GND 1.05f
C4311 a_16719_n13117.n20 GND 0.0503f
C4312 a_16719_n13117.n21 GND 0.0699f
C4313 a_16719_n13117.n22 GND 0.308f
C4314 a_16719_n13117.n23 GND 0.811f
C4315 a_16719_n13117.n24 GND 0.768f
C4316 a_16719_n13117.n25 GND 0.768f
C4317 a_16719_n13117.t9 GND 0.177f
C4318 a_16719_n13117.t17 GND 0.177f
C4319 a_16719_n13117.t21 GND 0.177f
C4320 a_16719_n13117.t13 GND 0.177f
C4321 a_16719_n13117.t6 GND 0.177f
C4322 a_16719_n13117.t10 GND 0.252f
C4323 a_16719_n13117.n26 GND 1.4f
C4324 a_16719_n13117.n27 GND 0.768f
C4325 a_16719_n13117.n28 GND 0.768f
C4326 a_16719_n13117.n29 GND 0.768f
C4327 a_16719_n13117.n30 GND 0.768f
C4328 a_16719_n13117.n31 GND 0.768f
C4329 a_16719_n13117.t23 GND 0.177f
C4330 a_16541_n13117.t16 GND 0.112f
C4331 a_16541_n13117.t9 GND 0.112f
C4332 a_16541_n13117.t5 GND 0.112f
C4333 a_16541_n13117.t13 GND 0.112f
C4334 a_16541_n13117.t19 GND 0.112f
C4335 a_16541_n13117.t7 GND 0.112f
C4336 a_16541_n13117.t18 GND 0.112f
C4337 a_16541_n13117.t2 GND 0.112f
C4338 a_16541_n13117.t6 GND 0.112f
C4339 a_16541_n13117.t21 GND 0.112f
C4340 a_16541_n13117.t12 GND 0.112f
C4341 a_16541_n13117.t15 GND 0.112f
C4342 a_16541_n13117.t4 GND 0.112f
C4343 a_16541_n13117.t10 GND 0.112f
C4344 a_16541_n13117.t17 GND 0.112f
C4345 a_16541_n13117.t11 GND 0.112f
C4346 a_16541_n13117.t14 GND 0.112f
C4347 a_16541_n13117.t3 GND 0.112f
C4348 a_16541_n13117.t8 GND 0.161f
C4349 a_16541_n13117.n0 GND 1.02f
C4350 a_16541_n13117.n1 GND 0.558f
C4351 a_16541_n13117.n2 GND 0.558f
C4352 a_16541_n13117.n3 GND 0.558f
C4353 a_16541_n13117.n4 GND 0.558f
C4354 a_16541_n13117.n5 GND 0.558f
C4355 a_16541_n13117.n6 GND 0.558f
C4356 a_16541_n13117.n7 GND 0.558f
C4357 a_16541_n13117.n8 GND 0.614f
C4358 a_16541_n13117.n9 GND 0.614f
C4359 a_16541_n13117.n10 GND 0.558f
C4360 a_16541_n13117.n11 GND 0.558f
C4361 a_16541_n13117.n12 GND 0.558f
C4362 a_16541_n13117.n13 GND 0.558f
C4363 a_16541_n13117.n14 GND 0.558f
C4364 a_16541_n13117.n15 GND 0.558f
C4365 a_16541_n13117.n16 GND 0.554f
C4366 a_16541_n13117.n17 GND 0.627f
C4367 a_16541_n13117.t20 GND 0.127f
C4368 a_16541_n13117.n18 GND 1.13f
C4369 a_16541_n13117.t1 GND 0.376f
C4370 a_16541_n13117.n19 GND 10.1f
C4371 a_16541_n13117.t0 GND 1.21f
C4372 a_16599_n13205.n0 GND 0.681f
C4373 a_16599_n13205.t15 GND 0.179f
C4374 a_16599_n13205.n1 GND 0.251f
C4375 a_16599_n13205.t8 GND 0.179f
C4376 a_16599_n13205.n2 GND 0.378f
C4377 a_16599_n13205.t23 GND 0.179f
C4378 a_16599_n13205.n3 GND 0.197f
C4379 a_16599_n13205.t12 GND 0.179f
C4380 a_16599_n13205.n4 GND 0.197f
C4381 a_16599_n13205.t20 GND 0.179f
C4382 a_16599_n13205.n5 GND 0.197f
C4383 a_16599_n13205.t13 GND 0.179f
C4384 a_16599_n13205.n6 GND 0.197f
C4385 a_16599_n13205.t7 GND 0.179f
C4386 a_16599_n13205.n7 GND 0.197f
C4387 a_16599_n13205.t22 GND 0.179f
C4388 a_16599_n13205.n8 GND 0.197f
C4389 a_16599_n13205.t11 GND 0.179f
C4390 a_16599_n13205.n9 GND 0.197f
C4391 a_16599_n13205.t16 GND 0.179f
C4392 a_16599_n13205.n10 GND 0.184f
C4393 a_16599_n13205.t2 GND 0.179f
C4394 a_16599_n13205.t5 GND 0.179f
C4395 a_16599_n13205.t9 GND 0.179f
C4396 a_16599_n13205.t19 GND 0.179f
C4397 a_16599_n13205.t4 GND 0.179f
C4398 a_16599_n13205.t18 GND 0.179f
C4399 a_16599_n13205.t10 GND 0.179f
C4400 a_16599_n13205.t6 GND 0.179f
C4401 a_16599_n13205.t14 GND 0.179f
C4402 a_16599_n13205.t21 GND 0.179f
C4403 a_16599_n13205.t17 GND 0.179f
C4404 a_16599_n13205.n11 GND 0.252f
C4405 a_16599_n13205.n12 GND 0.376f
C4406 a_16599_n13205.n13 GND 0.197f
C4407 a_16599_n13205.n14 GND 0.197f
C4408 a_16599_n13205.n15 GND 0.197f
C4409 a_16599_n13205.n16 GND 0.197f
C4410 a_16599_n13205.n17 GND 0.197f
C4411 a_16599_n13205.n18 GND 0.197f
C4412 a_16599_n13205.n19 GND 0.197f
C4413 a_16599_n13205.n20 GND 0.197f
C4414 a_16599_n13205.n21 GND 0.169f
C4415 a_16599_n13205.n22 GND 0.102f
C4416 a_16599_n13205.n23 GND 0.377f
C4417 a_16599_n13205.n24 GND 0.197f
C4418 a_16599_n13205.n25 GND 0.197f
C4419 a_16599_n13205.n26 GND 0.197f
C4420 a_16599_n13205.n27 GND 0.197f
C4421 a_16599_n13205.n28 GND 0.197f
C4422 a_16599_n13205.n29 GND 0.197f
C4423 a_16599_n13205.n30 GND 0.197f
C4424 a_16599_n13205.n31 GND 0.184f
C4425 a_16599_n13205.n32 GND 0.376f
C4426 a_16599_n13205.n33 GND 0.197f
C4427 a_16599_n13205.n34 GND 0.197f
C4428 a_16599_n13205.n35 GND 0.197f
C4429 a_16599_n13205.n36 GND 0.197f
C4430 a_16599_n13205.n37 GND 0.197f
C4431 a_16599_n13205.n38 GND 0.197f
C4432 a_16599_n13205.n39 GND 0.197f
C4433 a_16599_n13205.n40 GND 0.197f
C4434 a_16599_n13205.n41 GND 0.169f
C4435 a_16599_n13205.n42 GND 0.108f
C4436 a_16599_n13205.t3 GND 0.0381f
C4437 a_16599_n13205.n43 GND 2.83f
C4438 a_16599_n13205.t1 GND 1.94f
C4439 VV16.t16 GND 0.0223f
C4440 VV16.n0 GND 0.183f
C4441 VV16.n1 GND 0.077f
C4442 VV16.t0 GND 0.292f
C4443 VV16.t15 GND 0.292f
C4444 VV16.t13 GND 0.292f
C4445 VV16.t11 GND 0.292f
C4446 VV16.t9 GND 0.292f
C4447 VV16.t8 GND 0.292f
C4448 VV16.t1 GND 0.292f
C4449 VV16.t4 GND 0.292f
C4450 VV16.t14 GND 0.292f
C4451 VV16.t2 GND 0.292f
C4452 VV16.t6 GND 0.292f
C4453 VV16.t3 GND 0.292f
C4454 VV16.t12 GND 0.292f
C4455 VV16.t10 GND 0.292f
C4456 VV16.t5 GND 0.292f
C4457 VV16.t7 GND 0.629f
C4458 VV16.n2 GND 0.362f
C4459 VV16.n3 GND 0.359f
C4460 VV16.n4 GND 0.359f
C4461 VV16.n5 GND 0.359f
C4462 VV16.n6 GND 0.359f
C4463 VV16.n7 GND 0.359f
C4464 VV16.n8 GND 0.359f
C4465 VV16.n9 GND 0.359f
C4466 VV16.n10 GND 0.359f
C4467 VV16.n11 GND 0.359f
C4468 VV16.n12 GND 0.359f
C4469 VV16.n13 GND 0.359f
C4470 VV16.n14 GND 0.359f
C4471 VV16.n15 GND 0.359f
C4472 VV16.n16 GND 0.291f
C4473 VV16.n17 GND 3.07f
C4474 VFS.t0 GND 0.108f
C4475 VFS.n0 GND 0.0961f
C4476 VFS.n1 GND 0.0961f
C4477 VFS.n2 GND 0.0687f
C4478 VFS.n3 GND 2.49f
C4479 VFS.t2 GND 0.0898f
C4480 VFS.n4 GND 0.0961f
C4481 VFS.n5 GND 0.0961f
C4482 VFS.n6 GND 0.0741f
C4483 OUT2.n2 GND 0.0114f
C4484 OUT2.n4 GND 0.0241f
C4485 OUT2.n6 GND 0.0161f
C4486 OUT2.n8 GND 0.0161f
C4487 OUT2.n10 GND 0.0161f
C4488 OUT2.n12 GND 0.0161f
C4489 OUT2.n14 GND 0.0161f
C4490 OUT2.n23 GND 0.014f
C4491 OUT2.n25 GND 0.0348f
C4492 OUT2.n27 GND 0.021f
C4493 OUT2.n29 GND 0.021f
C4494 OUT2.n31 GND 0.021f
C4495 OUT2.n33 GND 0.021f
C4496 OUT2.n35 GND 0.021f
C4497 OUT2.n37 GND 0.0147f
C4498 OUT2.n38 GND 0.0296f
C4499 OUT2.n39 GND 0.0229f
C4500 OUT2.n42 GND 0.0114f
C4501 OUT2.n44 GND 0.0241f
C4502 OUT2.n46 GND 0.0161f
C4503 OUT2.n48 GND 0.0161f
C4504 OUT2.n50 GND 0.0161f
C4505 OUT2.n52 GND 0.0161f
C4506 OUT2.n54 GND 0.0161f
C4507 OUT2.n63 GND 0.014f
C4508 OUT2.n65 GND 0.0348f
C4509 OUT2.n67 GND 0.021f
C4510 OUT2.n69 GND 0.021f
C4511 OUT2.n71 GND 0.021f
C4512 OUT2.n73 GND 0.021f
C4513 OUT2.n75 GND 0.021f
C4514 OUT2.n77 GND 0.0147f
C4515 OUT2.n78 GND 0.0273f
C4516 OUT2.n79 GND 0.0203f
C4517 OUT2.n81 GND 0.0114f
C4518 OUT2.n83 GND 0.0241f
C4519 OUT2.n85 GND 0.0161f
C4520 OUT2.n87 GND 0.0161f
C4521 OUT2.n89 GND 0.0161f
C4522 OUT2.n91 GND 0.0161f
C4523 OUT2.n93 GND 0.0161f
C4524 OUT2.n97 GND 0.0126f
C4525 OUT2.n100 GND 0.014f
C4526 OUT2.n102 GND 0.0348f
C4527 OUT2.n104 GND 0.021f
C4528 OUT2.n106 GND 0.021f
C4529 OUT2.n108 GND 0.021f
C4530 OUT2.n110 GND 0.021f
C4531 OUT2.n112 GND 0.021f
C4532 OUT2.n114 GND 0.0147f
C4533 OUT2.n115 GND 0.0284f
C4534 OUT2.n116 GND 0.0234f
C4535 OUT2.n120 GND 0.014f
C4536 OUT2.n122 GND 0.0348f
C4537 OUT2.n124 GND 0.021f
C4538 OUT2.n126 GND 0.021f
C4539 OUT2.n128 GND 0.021f
C4540 OUT2.n130 GND 0.021f
C4541 OUT2.n132 GND 0.021f
C4542 OUT2.n136 GND 0.0114f
C4543 OUT2.n138 GND 0.0241f
C4544 OUT2.n140 GND 0.0161f
C4545 OUT2.n142 GND 0.0161f
C4546 OUT2.n144 GND 0.0161f
C4547 OUT2.n146 GND 0.0161f
C4548 OUT2.n148 GND 0.0161f
C4549 OUT2.n152 GND 0.013f
C4550 OUT2.n155 GND 0.0204f
C4551 OUT2.n156 GND 0.108f
C4552 OUT2.n157 GND 0.275f
C4553 OUT2.n158 GND 0.224f
C4554 OUT2.n159 GND 0.228f
C4555 I5.t11 GND 0.0123f
C4556 I5.n3 GND 0.0135f
C4557 I5.n8 GND 0.15f
C4558 I5.n9 GND 0.374f
C4559 I5.n12 GND 0.0114f
C4560 I5.n16 GND 0.213f
C4561 I5.n21 GND 0.567f
C4562 I5.n22 GND 1.34f
C4563 I5.n23 GND 0.305f
C4564 I5.n24 GND 0.686f
C4565 I5.n25 GND 1.29f
C4566 I5.t12 GND 0.0276f
C4567 I5.n26 GND 0.432f
C4568 I5.n27 GND 0.0573f
C4569 I5.n28 GND 0.13f
C4570 I5.n29 GND 0.0861f
C4571 I5.n30 GND 0.0921f
C4572 I5.n31 GND 0.127f
C4573 I5.n32 GND 0.12f
C4574 I5.t3 GND 0.0102f
C4575 I5.n33 GND 0.276f
C4576 I5.n34 GND 10.4f
C4577 I5.n35 GND 2.15f
C4578 OUT0.n2 GND 0.0114f
C4579 OUT0.n4 GND 0.0241f
C4580 OUT0.n6 GND 0.0161f
C4581 OUT0.n8 GND 0.0161f
C4582 OUT0.n10 GND 0.0161f
C4583 OUT0.n12 GND 0.0161f
C4584 OUT0.n14 GND 0.0161f
C4585 OUT0.n23 GND 0.014f
C4586 OUT0.n25 GND 0.0348f
C4587 OUT0.n27 GND 0.021f
C4588 OUT0.n29 GND 0.021f
C4589 OUT0.n31 GND 0.021f
C4590 OUT0.n33 GND 0.021f
C4591 OUT0.n35 GND 0.021f
C4592 OUT0.n37 GND 0.0147f
C4593 OUT0.n38 GND 0.0296f
C4594 OUT0.n39 GND 0.0229f
C4595 OUT0.n42 GND 0.0114f
C4596 OUT0.n44 GND 0.0241f
C4597 OUT0.n46 GND 0.0161f
C4598 OUT0.n48 GND 0.0161f
C4599 OUT0.n50 GND 0.0161f
C4600 OUT0.n52 GND 0.0161f
C4601 OUT0.n54 GND 0.0161f
C4602 OUT0.n63 GND 0.014f
C4603 OUT0.n65 GND 0.0348f
C4604 OUT0.n67 GND 0.021f
C4605 OUT0.n69 GND 0.021f
C4606 OUT0.n71 GND 0.021f
C4607 OUT0.n73 GND 0.021f
C4608 OUT0.n75 GND 0.021f
C4609 OUT0.n77 GND 0.0147f
C4610 OUT0.n78 GND 0.0273f
C4611 OUT0.n79 GND 0.0203f
C4612 OUT0.n81 GND 0.0114f
C4613 OUT0.n83 GND 0.0241f
C4614 OUT0.n85 GND 0.0161f
C4615 OUT0.n87 GND 0.0161f
C4616 OUT0.n89 GND 0.0161f
C4617 OUT0.n91 GND 0.0161f
C4618 OUT0.n93 GND 0.0161f
C4619 OUT0.n97 GND 0.0126f
C4620 OUT0.n100 GND 0.014f
C4621 OUT0.n102 GND 0.0348f
C4622 OUT0.n104 GND 0.021f
C4623 OUT0.n106 GND 0.021f
C4624 OUT0.n108 GND 0.021f
C4625 OUT0.n110 GND 0.021f
C4626 OUT0.n112 GND 0.021f
C4627 OUT0.n114 GND 0.0147f
C4628 OUT0.n115 GND 0.0284f
C4629 OUT0.n116 GND 0.0234f
C4630 OUT0.n120 GND 0.014f
C4631 OUT0.n122 GND 0.0348f
C4632 OUT0.n124 GND 0.021f
C4633 OUT0.n126 GND 0.021f
C4634 OUT0.n128 GND 0.021f
C4635 OUT0.n130 GND 0.021f
C4636 OUT0.n132 GND 0.021f
C4637 OUT0.n136 GND 0.0114f
C4638 OUT0.n138 GND 0.0241f
C4639 OUT0.n140 GND 0.0161f
C4640 OUT0.n142 GND 0.0161f
C4641 OUT0.n144 GND 0.0161f
C4642 OUT0.n146 GND 0.0161f
C4643 OUT0.n148 GND 0.0161f
C4644 OUT0.n152 GND 0.013f
C4645 OUT0.n155 GND 0.0204f
C4646 OUT0.n156 GND 0.108f
C4647 OUT0.n157 GND 0.275f
C4648 OUT0.n158 GND 0.224f
C4649 OUT0.n159 GND 0.228f
C4650 frontAnalog_v0p0p1_15.x63.A.n0 GND 0.12f
C4651 frontAnalog_v0p0p1_15.x63.A.n1 GND 2.22f
C4652 frontAnalog_v0p0p1_15.x63.A.t6 GND 0.014f
C4653 frontAnalog_v0p0p1_15.x63.A.t4 GND 0.0225f
C4654 frontAnalog_v0p0p1_15.x63.A.n2 GND 0.0465f
C4655 frontAnalog_v0p0p1_15.x63.A.t1 GND 0.151f
C4656 frontAnalog_v0p0p1_15.x63.A.t3 GND 0.0156f
C4657 frontAnalog_v0p0p1_15.x63.A.t2 GND 0.335f
C4658 frontAnalog_v0p0p1_15.x63.A.t5 GND 0.0256f
C4659 frontAnalog_v0p0p1_15.x63.A.t0 GND 0.173f
C4660 frontAnalog_v0p0p1_15.x63.A.t7 GND 0.175f
C4661 frontAnalog_v0p0p1_15.x63.A.n3 GND 1f
C4662 frontAnalog_v0p0p1_15.x63.A.n4 GND 0.953f
C4663 frontAnalog_v0p0p1_15.x63.A.n5 GND 1.25f
C4664 OUT3.n5 GND 0.0122f
C4665 OUT3.n7 GND 0.0305f
C4666 OUT3.n9 GND 0.0184f
C4667 OUT3.n11 GND 0.0184f
C4668 OUT3.n13 GND 0.0184f
C4669 OUT3.n15 GND 0.0184f
C4670 OUT3.n17 GND 0.0184f
C4671 OUT3.n26 GND 0.0212f
C4672 OUT3.n28 GND 0.0141f
C4673 OUT3.n30 GND 0.0141f
C4674 OUT3.n32 GND 0.0141f
C4675 OUT3.n34 GND 0.0141f
C4676 OUT3.n36 GND 0.0141f
C4677 OUT3.n44 GND 0.027f
C4678 OUT3.n45 GND 0.0219f
C4679 OUT3.n51 GND 0.0122f
C4680 OUT3.n53 GND 0.0305f
C4681 OUT3.n55 GND 0.0184f
C4682 OUT3.n57 GND 0.0184f
C4683 OUT3.n59 GND 0.0184f
C4684 OUT3.n61 GND 0.0184f
C4685 OUT3.n63 GND 0.0184f
C4686 OUT3.n66 GND 0.0157f
C4687 OUT3.n72 GND 0.0212f
C4688 OUT3.n74 GND 0.0141f
C4689 OUT3.n76 GND 0.0141f
C4690 OUT3.n78 GND 0.0141f
C4691 OUT3.n80 GND 0.0141f
C4692 OUT3.n82 GND 0.0141f
C4693 OUT3.n85 GND 0.015f
C4694 OUT3.n86 GND 0.0477f
C4695 OUT3.n87 GND 0.0111f
C4696 OUT3.n89 GND 0.0122f
C4697 OUT3.n91 GND 0.0305f
C4698 OUT3.n93 GND 0.0184f
C4699 OUT3.n95 GND 0.0184f
C4700 OUT3.n97 GND 0.0184f
C4701 OUT3.n99 GND 0.0184f
C4702 OUT3.n101 GND 0.0184f
C4703 OUT3.n114 GND 0.0212f
C4704 OUT3.n116 GND 0.0141f
C4705 OUT3.n118 GND 0.0141f
C4706 OUT3.n120 GND 0.0141f
C4707 OUT3.n122 GND 0.0141f
C4708 OUT3.n124 GND 0.0141f
C4709 OUT3.n133 GND 0.0282f
C4710 OUT3.n134 GND 0.0213f
C4711 OUT3.n140 GND 0.0122f
C4712 OUT3.n142 GND 0.0305f
C4713 OUT3.n144 GND 0.0184f
C4714 OUT3.n146 GND 0.0184f
C4715 OUT3.n148 GND 0.0184f
C4716 OUT3.n150 GND 0.0184f
C4717 OUT3.n152 GND 0.0184f
C4718 OUT3.n160 GND 0.0212f
C4719 OUT3.n162 GND 0.0141f
C4720 OUT3.n164 GND 0.0141f
C4721 OUT3.n166 GND 0.0141f
C4722 OUT3.n168 GND 0.0141f
C4723 OUT3.n170 GND 0.0141f
C4724 OUT3.n179 GND 0.027f
C4725 OUT3.n180 GND 0.119f
C4726 OUT3.n181 GND 0.304f
C4727 OUT3.n182 GND 0.264f
C4728 OUT3.n183 GND 0.577f
C4729 VDD.t1064 GND 0.0126f
C4730 VDD.t358 GND 0.0124f
C4731 VDD.t69 GND 0.0105f
C4732 VDD.t455 GND 0.0129f
C4733 VDD.t1122 GND 0.0134f
C4734 VDD.t449 GND 0.0107f
C4735 VDD.t360 GND 0.0281f
C4736 VDD.t974 GND 0.0485f
C4737 VDD.t836 GND 0.0199f
C4738 VDD.t605 GND 0.0209f
C4739 VDD.t471 GND 0.0209f
C4740 VDD.t1464 GND 0.0241f
C4741 VDD.t1454 GND 0.0392f
C4742 VDD.n0 GND 0.0192f
C4743 VDD.n26 GND 0.0309f
C4744 VDD.n28 GND 0.013f
C4745 VDD.n33 GND 0.0119f
C4746 VDD.n34 GND 0.119f
C4747 VDD.n35 GND 0.374f
C4748 VDD.n59 GND 0.0109f
C4749 VDD.t17 GND 0.116f
C4750 VDD.t426 GND 0.0557f
C4751 VDD.t635 GND 0.117f
C4752 VDD.t285 GND 0.0442f
C4753 VDD.n60 GND 0.0473f
C4754 VDD.n61 GND 0.0682f
C4755 VDD.n62 GND 0.734f
C4756 VDD.t804 GND 0.0191f
C4757 VDD.t1486 GND 0.0128f
C4758 VDD.t645 GND 0.0119f
C4759 VDD.t785 GND 0.0133f
C4760 VDD.t629 GND 0.0122f
C4761 VDD.t1452 GND 0.011f
C4762 VDD.t1489 GND 0.0158f
C4763 VDD.t431 GND 0.0129f
C4764 VDD.t801 GND 0.0159f
C4765 VDD.t1376 GND 0.0246f
C4766 VDD.t502 GND 0.0354f
C4767 VDD.t1443 GND 0.0205f
C4768 VDD.t457 GND 0.0215f
C4769 VDD.t595 GND 0.0215f
C4770 VDD.t287 GND 0.0249f
C4771 VDD.t429 GND 0.0409f
C4772 VDD.n79 GND 0.0137f
C4773 VDD.n108 GND 0.0126f
C4774 VDD.n109 GND 0.0862f
C4775 VDD.n110 GND 0.735f
C4776 VDD.n114 GND 0.0334f
C4777 VDD.n117 GND 0.0144f
C4778 VDD.n120 GND 0.0144f
C4779 VDD.t664 GND 0.0109f
C4780 VDD.n127 GND 0.0327f
C4781 VDD.t654 GND 0.0428f
C4782 VDD.t680 GND 0.0183f
C4783 VDD.t766 GND 0.0183f
C4784 VDD.t658 GND 0.0183f
C4785 VDD.t778 GND 0.0183f
C4786 VDD.t670 GND 0.0124f
C4787 VDD.n130 GND 0.0218f
C4788 VDD.n132 GND 0.136f
C4789 VDD.n136 GND 0.0301f
C4790 VDD.n137 GND 0.0182f
C4791 VDD.n139 GND 0.0129f
C4792 VDD.n143 GND 0.0339f
C4793 VDD.n147 GND 0.0339f
C4794 VDD.n149 GND 0.0339f
C4795 VDD.n150 GND 0.0255f
C4796 VDD.n151 GND 0.0201f
C4797 VDD.n153 GND 0.0339f
C4798 VDD.n157 GND 0.0339f
C4799 VDD.n159 GND 0.0339f
C4800 VDD.n163 GND 0.0339f
C4801 VDD.n165 GND 0.0339f
C4802 VDD.n169 GND 0.0339f
C4803 VDD.n171 GND 0.0339f
C4804 VDD.n175 GND 0.029f
C4805 VDD.n176 GND 0.0182f
C4806 VDD.n180 GND 0.0129f
C4807 VDD.n181 GND 0.017f
C4808 VDD.n182 GND 0.0144f
C4809 VDD.n183 GND 0.0147f
C4810 VDD.t698 GND 0.015f
C4811 VDD.t768 GND 0.0183f
C4812 VDD.t678 GND 0.0183f
C4813 VDD.t746 GND 0.0183f
C4814 VDD.t770 GND 0.0183f
C4815 VDD.t666 GND 0.0183f
C4816 VDD.t730 GND 0.0183f
C4817 VDD.t760 GND 0.0183f
C4818 VDD.t692 GND 0.0183f
C4819 VDD.t736 GND 0.0176f
C4820 VDD.t656 GND 0.0237f
C4821 VDD.t724 GND 0.0183f
C4822 VDD.t750 GND 0.0183f
C4823 VDD.t776 GND 0.0183f
C4824 VDD.t704 GND 0.0148f
C4825 VDD.t754 GND 0.0183f
C4826 VDD.t668 GND 0.0183f
C4827 VDD.t732 GND 0.0183f
C4828 VDD.t702 GND 0.0183f
C4829 VDD.t772 GND 0.0237f
C4830 VDD.t720 GND 0.0176f
C4831 VDD.t696 GND 0.0183f
C4832 VDD.t764 GND 0.0183f
C4833 VDD.t716 GND 0.0183f
C4834 VDD.t690 GND 0.0183f
C4835 VDD.t758 GND 0.0183f
C4836 VDD.t676 GND 0.0183f
C4837 VDD.t742 GND 0.0183f
C4838 VDD.t708 GND 0.0183f
C4839 VDD.t672 GND 0.0183f
C4840 VDD.t738 GND 0.0126f
C4841 VDD.n184 GND 0.0147f
C4842 VDD.n185 GND 0.0144f
C4843 VDD.n186 GND 0.0136f
C4844 VDD.n188 GND 0.0164f
C4845 VDD.n189 GND 0.0182f
C4846 VDD.n193 GND 0.0234f
C4847 VDD.n197 GND 0.0339f
C4848 VDD.n199 GND 0.0339f
C4849 VDD.n203 GND 0.0339f
C4850 VDD.n205 GND 0.0339f
C4851 VDD.n209 GND 0.0339f
C4852 VDD.n211 GND 0.0339f
C4853 VDD.n215 GND 0.0339f
C4854 VDD.n217 GND 0.0339f
C4855 VDD.n218 GND 0.0201f
C4856 VDD.n221 GND 0.0255f
C4857 VDD.n223 GND 0.0339f
C4858 VDD.n227 GND 0.0339f
C4859 VDD.n229 GND 0.0339f
C4860 VDD.n233 GND 0.0275f
C4861 VDD.n234 GND 0.0182f
C4862 VDD.n236 GND 0.0129f
C4863 VDD.n238 GND 0.0339f
C4864 VDD.n242 GND 0.0339f
C4865 VDD.n244 GND 0.0339f
C4866 VDD.n248 GND 0.0339f
C4867 VDD.n250 GND 0.0339f
C4868 VDD.n254 GND 0.0315f
C4869 VDD.n255 GND 0.0182f
C4870 VDD.n259 GND 0.0129f
C4871 VDD.n260 GND 0.017f
C4872 VDD.n261 GND 0.0144f
C4873 VDD.n262 GND 0.0147f
C4874 VDD.t728 GND 0.0165f
C4875 VDD.t756 GND 0.0183f
C4876 VDD.t686 GND 0.0183f
C4877 VDD.t712 GND 0.0183f
C4878 VDD.t744 GND 0.0183f
C4879 VDD.t688 GND 0.0183f
C4880 VDD.t714 GND 0.0183f
C4881 VDD.t660 GND 0.0183f
C4882 VDD.t682 GND 0.0183f
C4883 VDD.t700 GND 0.0176f
C4884 VDD.t722 GND 0.0237f
C4885 VDD.t748 GND 0.0183f
C4886 VDD.t774 GND 0.0183f
C4887 VDD.n263 GND 0.0147f
C4888 VDD.t752 GND 0.018f
C4889 VDD.t684 GND 0.0183f
C4890 VDD.t706 GND 0.0183f
C4891 VDD.t740 GND 0.0183f
C4892 VDD.t674 GND 0.0183f
C4893 VDD.t710 GND 0.0183f
C4894 VDD.t652 GND 0.0183f
C4895 VDD.t734 GND 0.0183f
C4896 VDD.t762 GND 0.0183f
C4897 VDD.t694 GND 0.0183f
C4898 VDD.t718 GND 0.0183f
C4899 VDD.t662 GND 0.0176f
C4900 VDD.t227 GND 0.0237f
C4901 VDD.t241 GND 0.0176f
C4902 VDD.n264 GND 0.0147f
C4903 VDD.t229 GND 0.0183f
C4904 VDD.t239 GND 0.0183f
C4905 VDD.t235 GND 0.0183f
C4906 VDD.t243 GND 0.0183f
C4907 VDD.t223 GND 0.0183f
C4908 VDD.t237 GND 0.0183f
C4909 VDD.t245 GND 0.0183f
C4910 VDD.t225 GND 0.0183f
C4911 VDD.t231 GND 0.0183f
C4912 VDD.t215 GND 0.0183f
C4913 VDD.t219 GND 0.0183f
C4914 VDD.t233 GND 0.0183f
C4915 VDD.t217 GND 0.0176f
C4916 VDD.t986 GND 0.0236f
C4917 VDD.t988 GND 0.0183f
C4918 VDD.t990 GND 0.0183f
C4919 VDD.t992 GND 0.0173f
C4920 VDD.t1290 GND 0.0194f
C4921 VDD.t1356 GND 0.0184f
C4922 VDD.t596 GND 0.0307f
C4923 VDD.t379 GND 0.0231f
C4924 VDD.n265 GND 0.0241f
C4925 VDD.n269 GND 0.0508f
C4926 VDD.n271 GND 0.0395f
C4927 VDD.n272 GND 0.0255f
C4928 VDD.n275 GND 0.0201f
C4929 VDD.n277 GND 0.0231f
C4930 VDD.n278 GND 0.0182f
C4931 VDD.n280 GND 0.0129f
C4932 VDD.n282 GND 0.0144f
C4933 VDD.n284 GND 0.019f
C4934 VDD.n286 GND 0.0339f
C4935 VDD.n289 GND 0.0339f
C4936 VDD.n291 GND 0.0339f
C4937 VDD.n292 GND 0.0255f
C4938 VDD.n293 GND 0.0201f
C4939 VDD.n295 GND 0.0339f
C4940 VDD.n299 GND 0.0339f
C4941 VDD.n301 GND 0.0339f
C4942 VDD.n305 GND 0.0339f
C4943 VDD.n307 GND 0.0339f
C4944 VDD.n311 GND 0.0339f
C4945 VDD.n313 GND 0.0339f
C4946 VDD.n317 GND 0.0339f
C4947 VDD.n321 GND 0.0339f
C4948 VDD.n323 GND 0.0339f
C4949 VDD.n327 GND 0.0312f
C4950 VDD.n328 GND 0.0182f
C4951 VDD.n330 GND 0.0129f
C4952 VDD.n331 GND 0.017f
C4953 VDD.n335 GND 0.0129f
C4954 VDD.n336 GND 0.0182f
C4955 VDD.n338 GND 0.0279f
C4956 VDD.n339 GND 0.0255f
C4957 VDD.n340 GND 0.0201f
C4958 VDD.n342 GND 0.0339f
C4959 VDD.n346 GND 0.0339f
C4960 VDD.n348 GND 0.0339f
C4961 VDD.n352 GND 0.0339f
C4962 VDD.n354 GND 0.0339f
C4963 VDD.n358 GND 0.0339f
C4964 VDD.n360 GND 0.0339f
C4965 VDD.n364 GND 0.0339f
C4966 VDD.n368 GND 0.0339f
C4967 VDD.n370 GND 0.0312f
C4968 VDD.n371 GND 0.0182f
C4969 VDD.n375 GND 0.0129f
C4970 VDD.n376 GND 0.017f
C4971 VDD.n378 GND 0.0129f
C4972 VDD.n379 GND 0.0182f
C4973 VDD.n383 GND 0.0279f
C4974 VDD.n385 GND 0.0339f
C4975 VDD.n386 GND 0.0255f
C4976 VDD.n387 GND 0.0201f
C4977 VDD.n389 GND 0.0175f
C4978 VDD.n390 GND 11.9f
C4979 VDD.t257 GND 0.0126f
C4980 VDD.t347 GND 0.0121f
C4981 VDD.t1321 GND 0.0106f
C4982 VDD.t1316 GND 0.0134f
C4983 VDD.t1441 GND 0.0121f
C4984 VDD.t1341 GND 0.0169f
C4985 VDD.t611 GND 0.0466f
C4986 VDD.n406 GND 0.0153f
C4987 VDD.n407 GND 0.257f
C4988 VDD.t470 GND 0.0452f
C4989 VDD.t967 GND 0.0156f
C4990 VDD.t326 GND 0.0346f
C4991 VDD.t364 GND 0.0646f
C4992 VDD.t362 GND 0.0275f
C4993 VDD.n408 GND 0.0207f
C4994 VDD.n437 GND 0.0116f
C4995 VDD.n438 GND 0.16f
C4996 VDD.n462 GND 0.0109f
C4997 VDD.t553 GND 0.116f
C4998 VDD.t73 GND 0.0557f
C4999 VDD.t460 GND 0.117f
C5000 VDD.t75 GND 0.0442f
C5001 VDD.n463 GND 0.0473f
C5002 VDD.n464 GND 0.0682f
C5003 VDD.t328 GND 0.0191f
C5004 VDD.t1493 GND 0.0128f
C5005 VDD.t491 GND 0.0119f
C5006 VDD.t345 GND 0.0133f
C5007 VDD.t71 GND 0.0122f
C5008 VDD.t1103 GND 0.011f
C5009 VDD.t1495 GND 0.0158f
C5010 VDD.t637 GND 0.0129f
C5011 VDD.t351 GND 0.0159f
C5012 VDD.t557 GND 0.0246f
C5013 VDD.t335 GND 0.0354f
C5014 VDD.t559 GND 0.0205f
C5015 VDD.t1066 GND 0.0215f
C5016 VDD.t598 GND 0.0215f
C5017 VDD.t468 GND 0.0249f
C5018 VDD.t411 GND 0.0409f
C5019 VDD.n481 GND 0.0137f
C5020 VDD.n510 GND 0.0126f
C5021 VDD.n511 GND 0.0862f
C5022 VDD.n512 GND 0.468f
C5023 VDD.n513 GND 0.59f
C5024 VDD.n515 GND 0.0172f
C5025 VDD.n518 GND 0.0144f
C5026 VDD.n521 GND 0.0144f
C5027 VDD.t111 GND 0.0113f
C5028 VDD.n528 GND 0.0334f
C5029 VDD.t101 GND 0.042f
C5030 VDD.t127 GND 0.0183f
C5031 VDD.t213 GND 0.0183f
C5032 VDD.t105 GND 0.0183f
C5033 VDD.t97 GND 0.0183f
C5034 VDD.t119 GND 0.0128f
C5035 VDD.n531 GND 0.0216f
C5036 VDD.n533 GND 0.135f
C5037 VDD.n537 GND 0.0308f
C5038 VDD.n538 GND 0.0182f
C5039 VDD.n540 GND 0.0129f
C5040 VDD.n544 GND 0.0339f
C5041 VDD.n548 GND 0.0339f
C5042 VDD.n550 GND 0.0339f
C5043 VDD.n551 GND 0.0255f
C5044 VDD.n552 GND 0.0201f
C5045 VDD.n554 GND 0.0339f
C5046 VDD.n558 GND 0.0339f
C5047 VDD.n560 GND 0.0339f
C5048 VDD.n564 GND 0.0339f
C5049 VDD.n566 GND 0.0339f
C5050 VDD.n570 GND 0.0339f
C5051 VDD.n572 GND 0.0339f
C5052 VDD.n576 GND 0.0282f
C5053 VDD.n577 GND 0.0182f
C5054 VDD.n581 GND 0.0129f
C5055 VDD.n582 GND 0.017f
C5056 VDD.n583 GND 0.0144f
C5057 VDD.n584 GND 0.0147f
C5058 VDD.t145 GND 0.0146f
C5059 VDD.t87 GND 0.0183f
C5060 VDD.t123 GND 0.0183f
C5061 VDD.t193 GND 0.0183f
C5062 VDD.t89 GND 0.0183f
C5063 VDD.t113 GND 0.0183f
C5064 VDD.t177 GND 0.0183f
C5065 VDD.t207 GND 0.0183f
C5066 VDD.t139 GND 0.0183f
C5067 VDD.t183 GND 0.0176f
C5068 VDD.t103 GND 0.0237f
C5069 VDD.t171 GND 0.0183f
C5070 VDD.t197 GND 0.0183f
C5071 VDD.t95 GND 0.0183f
C5072 VDD.t151 GND 0.0152f
C5073 VDD.t201 GND 0.0183f
C5074 VDD.t115 GND 0.0183f
C5075 VDD.t179 GND 0.0183f
C5076 VDD.t149 GND 0.0183f
C5077 VDD.t91 GND 0.0237f
C5078 VDD.t167 GND 0.0176f
C5079 VDD.t143 GND 0.0183f
C5080 VDD.t211 GND 0.0183f
C5081 VDD.t163 GND 0.0183f
C5082 VDD.t137 GND 0.0183f
C5083 VDD.t205 GND 0.0183f
C5084 VDD.t125 GND 0.0183f
C5085 VDD.t189 GND 0.0183f
C5086 VDD.t155 GND 0.0183f
C5087 VDD.t117 GND 0.0183f
C5088 VDD.t185 GND 0.0122f
C5089 VDD.n585 GND 0.0147f
C5090 VDD.n586 GND 0.0144f
C5091 VDD.n587 GND 0.0127f
C5092 VDD.n589 GND 0.0172f
C5093 VDD.n590 GND 0.0182f
C5094 VDD.n594 GND 0.0227f
C5095 VDD.n598 GND 0.0339f
C5096 VDD.n600 GND 0.0339f
C5097 VDD.n604 GND 0.0339f
C5098 VDD.n606 GND 0.0339f
C5099 VDD.n610 GND 0.0339f
C5100 VDD.n612 GND 0.0339f
C5101 VDD.n616 GND 0.0339f
C5102 VDD.n618 GND 0.0339f
C5103 VDD.n619 GND 0.0201f
C5104 VDD.n622 GND 0.0255f
C5105 VDD.n624 GND 0.0339f
C5106 VDD.n628 GND 0.0339f
C5107 VDD.n630 GND 0.0339f
C5108 VDD.n634 GND 0.0282f
C5109 VDD.n635 GND 0.0182f
C5110 VDD.n637 GND 0.0129f
C5111 VDD.n641 GND 0.0339f
C5112 VDD.n643 GND 0.0339f
C5113 VDD.n647 GND 0.0339f
C5114 VDD.n649 GND 0.0339f
C5115 VDD.n653 GND 0.0339f
C5116 VDD.n655 GND 0.0339f
C5117 VDD.n659 GND 0.0308f
C5118 VDD.n660 GND 0.0182f
C5119 VDD.n664 GND 0.0129f
C5120 VDD.n665 GND 0.017f
C5121 VDD.n666 GND 0.0144f
C5122 VDD.n667 GND 0.0147f
C5123 VDD.t175 GND 0.0161f
C5124 VDD.t203 GND 0.0183f
C5125 VDD.t133 GND 0.0183f
C5126 VDD.t159 GND 0.0183f
C5127 VDD.t191 GND 0.0183f
C5128 VDD.t135 GND 0.0183f
C5129 VDD.t161 GND 0.0183f
C5130 VDD.t107 GND 0.0183f
C5131 VDD.t129 GND 0.0183f
C5132 VDD.t147 GND 0.0176f
C5133 VDD.t169 GND 0.0237f
C5134 VDD.t195 GND 0.0183f
C5135 VDD.t93 GND 0.0183f
C5136 VDD.n668 GND 0.0147f
C5137 VDD.t199 GND 0.0176f
C5138 VDD.t131 GND 0.0183f
C5139 VDD.t153 GND 0.0183f
C5140 VDD.t187 GND 0.0183f
C5141 VDD.t121 GND 0.0183f
C5142 VDD.t157 GND 0.0183f
C5143 VDD.t99 GND 0.0183f
C5144 VDD.t181 GND 0.0183f
C5145 VDD.t209 GND 0.0183f
C5146 VDD.t141 GND 0.0183f
C5147 VDD.t165 GND 0.0183f
C5148 VDD.t109 GND 0.0176f
C5149 VDD.t1397 GND 0.0237f
C5150 VDD.t1411 GND 0.018f
C5151 VDD.n669 GND 0.0147f
C5152 VDD.t1399 GND 0.0183f
C5153 VDD.t1409 GND 0.0183f
C5154 VDD.t1405 GND 0.0183f
C5155 VDD.t1413 GND 0.0183f
C5156 VDD.t1393 GND 0.0183f
C5157 VDD.t1407 GND 0.0183f
C5158 VDD.t1415 GND 0.0183f
C5159 VDD.t1395 GND 0.0183f
C5160 VDD.t1401 GND 0.0183f
C5161 VDD.t1385 GND 0.0183f
C5162 VDD.t1389 GND 0.0183f
C5163 VDD.t1403 GND 0.0183f
C5164 VDD.t1387 GND 0.0176f
C5165 VDD.t339 GND 0.0236f
C5166 VDD.t341 GND 0.0183f
C5167 VDD.t343 GND 0.0183f
C5168 VDD.t337 GND 0.0173f
C5169 VDD.t1045 GND 0.0194f
C5170 VDD.t603 GND 0.0184f
C5171 VDD.t1046 GND 0.0307f
C5172 VDD.t780 GND 0.0226f
C5173 VDD.n670 GND 0.0241f
C5174 VDD.n674 GND 0.0508f
C5175 VDD.n676 GND 0.0395f
C5176 VDD.n677 GND 0.0255f
C5177 VDD.n680 GND 0.0201f
C5178 VDD.n682 GND 0.0223f
C5179 VDD.n683 GND 0.0182f
C5180 VDD.n685 GND 0.0129f
C5181 VDD.n687 GND 0.0144f
C5182 VDD.n689 GND 0.0197f
C5183 VDD.n691 GND 0.0339f
C5184 VDD.n694 GND 0.0339f
C5185 VDD.n696 GND 0.0339f
C5186 VDD.n697 GND 0.0255f
C5187 VDD.n698 GND 0.0201f
C5188 VDD.n700 GND 0.0339f
C5189 VDD.n704 GND 0.0339f
C5190 VDD.n706 GND 0.0339f
C5191 VDD.n710 GND 0.0339f
C5192 VDD.n712 GND 0.0339f
C5193 VDD.n716 GND 0.0339f
C5194 VDD.n718 GND 0.0339f
C5195 VDD.n722 GND 0.0339f
C5196 VDD.n726 GND 0.0339f
C5197 VDD.n728 GND 0.0339f
C5198 VDD.n732 GND 0.0304f
C5199 VDD.n733 GND 0.0182f
C5200 VDD.n735 GND 0.0129f
C5201 VDD.n736 GND 0.017f
C5202 VDD.n740 GND 0.0129f
C5203 VDD.n741 GND 0.0182f
C5204 VDD.n743 GND 0.0286f
C5205 VDD.n744 GND 0.0255f
C5206 VDD.n745 GND 0.0201f
C5207 VDD.n747 GND 0.0339f
C5208 VDD.n751 GND 0.0339f
C5209 VDD.n753 GND 0.0339f
C5210 VDD.n757 GND 0.0339f
C5211 VDD.n759 GND 0.0339f
C5212 VDD.n763 GND 0.0339f
C5213 VDD.n765 GND 0.0339f
C5214 VDD.n769 GND 0.0339f
C5215 VDD.n773 GND 0.0339f
C5216 VDD.n775 GND 0.0304f
C5217 VDD.n776 GND 0.0182f
C5218 VDD.n780 GND 0.0129f
C5219 VDD.n781 GND 0.017f
C5220 VDD.n783 GND 0.0129f
C5221 VDD.n784 GND 0.0182f
C5222 VDD.n788 GND 0.0286f
C5223 VDD.n790 GND 0.0339f
C5224 VDD.n791 GND 0.0255f
C5225 VDD.n792 GND 0.0199f
C5226 VDD.n793 GND 11.9f
C5227 VDD.n794 GND 3.73f
C5228 VDD.n795 GND 0.519f
C5229 VDD.n796 GND 0.596f
C5230 VDD.n797 GND 2.81f
C5231 VDD.n798 GND 1.01f
C5232 VDD.n799 GND 0.0114f
C5233 VDD.n802 GND 0.0124f
C5234 VDD.n807 GND 0.0138f
C5235 VDD.n808 GND 0.0561f
C5236 VDD.n814 GND 0.0124f
C5237 VDD.n815 GND 0.0124f
C5238 VDD.n820 GND 0.0323f
C5239 VDD.n853 GND 0.0239f
C5240 VDD.t551 GND 0.0103f
C5241 VDD.t356 GND 0.0258f
C5242 VDD.t613 GND 0.0248f
C5243 VDD.t621 GND 0.0302f
C5244 VDD.t1090 GND 0.026f
C5245 VDD.t1110 GND 0.0225f
C5246 VDD.t1345 GND 0.0188f
C5247 VDD.t588 GND 0.0298f
C5248 VDD.t1096 GND 0.026f
C5249 VDD.t1107 GND 0.0225f
C5250 VDD.t334 GND 0.0225f
C5251 VDD.t782 GND 0.0215f
C5252 VDD.t330 GND 0.0231f
C5253 VDD.t1343 GND 0.0229f
C5254 VDD.t1314 GND 0.0231f
C5255 VDD.t1319 GND 0.0231f
C5256 VDD.t354 GND 0.0291f
C5257 VDD.n857 GND 0.0705f
C5258 VDD.n861 GND 0.0196f
C5259 VDD.n862 GND 0.0687f
C5260 VDD.n863 GND 4.84f
C5261 VDD.n865 GND 0.0172f
C5262 VDD.n868 GND 0.0144f
C5263 VDD.n871 GND 0.0144f
C5264 VDD.t884 GND 0.0113f
C5265 VDD.n878 GND 0.0334f
C5266 VDD.t874 GND 0.042f
C5267 VDD.t900 GND 0.0183f
C5268 VDD.t858 GND 0.0183f
C5269 VDD.t878 GND 0.0183f
C5270 VDD.t870 GND 0.0183f
C5271 VDD.t890 GND 0.0128f
C5272 VDD.n881 GND 0.0216f
C5273 VDD.n883 GND 0.135f
C5274 VDD.n887 GND 0.0308f
C5275 VDD.n888 GND 0.0182f
C5276 VDD.n890 GND 0.0129f
C5277 VDD.n894 GND 0.0339f
C5278 VDD.n898 GND 0.0339f
C5279 VDD.n900 GND 0.0339f
C5280 VDD.n901 GND 0.0255f
C5281 VDD.n902 GND 0.0201f
C5282 VDD.n904 GND 0.0339f
C5283 VDD.n908 GND 0.0339f
C5284 VDD.n910 GND 0.0339f
C5285 VDD.n914 GND 0.0339f
C5286 VDD.n916 GND 0.0339f
C5287 VDD.n920 GND 0.0339f
C5288 VDD.n922 GND 0.0339f
C5289 VDD.n926 GND 0.0282f
C5290 VDD.n927 GND 0.0182f
C5291 VDD.n931 GND 0.0129f
C5292 VDD.n932 GND 0.017f
C5293 VDD.n933 GND 0.0144f
C5294 VDD.n934 GND 0.0147f
C5295 VDD.t918 GND 0.0146f
C5296 VDD.t860 GND 0.0183f
C5297 VDD.t896 GND 0.0183f
C5298 VDD.t838 GND 0.0183f
C5299 VDD.t862 GND 0.0183f
C5300 VDD.t886 GND 0.0183f
C5301 VDD.t950 GND 0.0183f
C5302 VDD.t852 GND 0.0183f
C5303 VDD.t912 GND 0.0183f
C5304 VDD.t956 GND 0.0176f
C5305 VDD.t876 GND 0.0237f
C5306 VDD.t932 GND 0.0183f
C5307 VDD.t842 GND 0.0183f
C5308 VDD.t868 GND 0.0183f
C5309 VDD.t924 GND 0.0152f
C5310 VDD.t846 GND 0.0183f
C5311 VDD.t888 GND 0.0183f
C5312 VDD.t952 GND 0.0183f
C5313 VDD.t922 GND 0.0183f
C5314 VDD.t864 GND 0.0237f
C5315 VDD.t942 GND 0.0176f
C5316 VDD.t916 GND 0.0183f
C5317 VDD.t856 GND 0.0183f
C5318 VDD.t938 GND 0.0183f
C5319 VDD.t910 GND 0.0183f
C5320 VDD.t850 GND 0.0183f
C5321 VDD.t898 GND 0.0183f
C5322 VDD.t962 GND 0.0183f
C5323 VDD.t928 GND 0.0183f
C5324 VDD.t892 GND 0.0183f
C5325 VDD.t958 GND 0.0122f
C5326 VDD.n935 GND 0.0147f
C5327 VDD.n936 GND 0.0144f
C5328 VDD.n937 GND 0.0127f
C5329 VDD.n939 GND 0.0172f
C5330 VDD.n940 GND 0.0182f
C5331 VDD.n944 GND 0.0227f
C5332 VDD.n948 GND 0.0339f
C5333 VDD.n950 GND 0.0339f
C5334 VDD.n954 GND 0.0339f
C5335 VDD.n956 GND 0.0339f
C5336 VDD.n960 GND 0.0339f
C5337 VDD.n962 GND 0.0339f
C5338 VDD.n966 GND 0.0339f
C5339 VDD.n968 GND 0.0339f
C5340 VDD.n969 GND 0.0201f
C5341 VDD.n972 GND 0.0255f
C5342 VDD.n974 GND 0.0339f
C5343 VDD.n978 GND 0.0339f
C5344 VDD.n980 GND 0.0339f
C5345 VDD.n984 GND 0.0282f
C5346 VDD.n985 GND 0.0182f
C5347 VDD.n987 GND 0.0129f
C5348 VDD.n991 GND 0.0339f
C5349 VDD.n993 GND 0.0339f
C5350 VDD.n997 GND 0.0339f
C5351 VDD.n999 GND 0.0339f
C5352 VDD.n1003 GND 0.0339f
C5353 VDD.n1005 GND 0.0339f
C5354 VDD.n1009 GND 0.0308f
C5355 VDD.n1010 GND 0.0182f
C5356 VDD.n1014 GND 0.0129f
C5357 VDD.n1015 GND 0.017f
C5358 VDD.n1016 GND 0.0144f
C5359 VDD.n1017 GND 0.0147f
C5360 VDD.t948 GND 0.0161f
C5361 VDD.t848 GND 0.0183f
C5362 VDD.t902 GND 0.0183f
C5363 VDD.t934 GND 0.0183f
C5364 VDD.t964 GND 0.0183f
C5365 VDD.t908 GND 0.0183f
C5366 VDD.t936 GND 0.0183f
C5367 VDD.t880 GND 0.0183f
C5368 VDD.t904 GND 0.0183f
C5369 VDD.t920 GND 0.0176f
C5370 VDD.t944 GND 0.0237f
C5371 VDD.t840 GND 0.0183f
C5372 VDD.t866 GND 0.0183f
C5373 VDD.n1018 GND 0.0147f
C5374 VDD.t844 GND 0.0176f
C5375 VDD.t906 GND 0.0183f
C5376 VDD.t926 GND 0.0183f
C5377 VDD.t960 GND 0.0183f
C5378 VDD.t894 GND 0.0183f
C5379 VDD.t930 GND 0.0183f
C5380 VDD.t872 GND 0.0183f
C5381 VDD.t954 GND 0.0183f
C5382 VDD.t854 GND 0.0183f
C5383 VDD.t914 GND 0.0183f
C5384 VDD.t940 GND 0.0183f
C5385 VDD.t882 GND 0.0176f
C5386 VDD.t53 GND 0.0237f
C5387 VDD.t35 GND 0.018f
C5388 VDD.n1019 GND 0.0147f
C5389 VDD.t55 GND 0.0183f
C5390 VDD.t65 GND 0.0183f
C5391 VDD.t61 GND 0.0183f
C5392 VDD.t37 GND 0.0183f
C5393 VDD.t49 GND 0.0183f
C5394 VDD.t63 GND 0.0183f
C5395 VDD.t39 GND 0.0183f
C5396 VDD.t51 GND 0.0183f
C5397 VDD.t57 GND 0.0183f
C5398 VDD.t41 GND 0.0183f
C5399 VDD.t45 GND 0.0183f
C5400 VDD.t59 GND 0.0183f
C5401 VDD.t43 GND 0.0176f
C5402 VDD.t1080 GND 0.0236f
C5403 VDD.t1082 GND 0.0183f
C5404 VDD.t1076 GND 0.0183f
C5405 VDD.t1078 GND 0.0173f
C5406 VDD.t819 GND 0.0194f
C5407 VDD.t1351 GND 0.0184f
C5408 VDD.t1431 GND 0.0307f
C5409 VDD.t1484 GND 0.0226f
C5410 VDD.n1020 GND 0.0241f
C5411 VDD.n1024 GND 0.0508f
C5412 VDD.n1026 GND 0.0395f
C5413 VDD.n1027 GND 0.0255f
C5414 VDD.n1030 GND 0.0201f
C5415 VDD.n1032 GND 0.0223f
C5416 VDD.n1033 GND 0.0182f
C5417 VDD.n1035 GND 0.0129f
C5418 VDD.n1037 GND 0.0144f
C5419 VDD.n1039 GND 0.0197f
C5420 VDD.n1041 GND 0.0339f
C5421 VDD.n1044 GND 0.0339f
C5422 VDD.n1046 GND 0.0339f
C5423 VDD.n1047 GND 0.0255f
C5424 VDD.n1048 GND 0.0201f
C5425 VDD.n1050 GND 0.0339f
C5426 VDD.n1054 GND 0.0339f
C5427 VDD.n1056 GND 0.0339f
C5428 VDD.n1060 GND 0.0339f
C5429 VDD.n1062 GND 0.0339f
C5430 VDD.n1066 GND 0.0339f
C5431 VDD.n1068 GND 0.0339f
C5432 VDD.n1072 GND 0.0339f
C5433 VDD.n1076 GND 0.0339f
C5434 VDD.n1078 GND 0.0339f
C5435 VDD.n1082 GND 0.0304f
C5436 VDD.n1083 GND 0.0182f
C5437 VDD.n1085 GND 0.0129f
C5438 VDD.n1086 GND 0.017f
C5439 VDD.n1090 GND 0.0129f
C5440 VDD.n1091 GND 0.0182f
C5441 VDD.n1093 GND 0.0286f
C5442 VDD.n1094 GND 0.0255f
C5443 VDD.n1095 GND 0.0201f
C5444 VDD.n1097 GND 0.0339f
C5445 VDD.n1101 GND 0.0339f
C5446 VDD.n1103 GND 0.0339f
C5447 VDD.n1107 GND 0.0339f
C5448 VDD.n1109 GND 0.0339f
C5449 VDD.n1113 GND 0.0339f
C5450 VDD.n1115 GND 0.0339f
C5451 VDD.n1119 GND 0.0339f
C5452 VDD.n1123 GND 0.0339f
C5453 VDD.n1125 GND 0.0304f
C5454 VDD.n1126 GND 0.0182f
C5455 VDD.n1130 GND 0.0129f
C5456 VDD.n1131 GND 0.017f
C5457 VDD.n1133 GND 0.0129f
C5458 VDD.n1134 GND 0.0182f
C5459 VDD.n1138 GND 0.0286f
C5460 VDD.n1140 GND 0.0339f
C5461 VDD.n1141 GND 0.0255f
C5462 VDD.n1142 GND 0.0199f
C5463 VDD.n1143 GND 13.2f
C5464 VDD.t971 GND 0.0126f
C5465 VDD.t810 GND 0.0124f
C5466 VDD.t627 GND 0.0105f
C5467 VDD.t462 GND 0.0129f
C5468 VDD.t1457 GND 0.0134f
C5469 VDD.t565 GND 0.0107f
C5470 VDD.t813 GND 0.0281f
C5471 VDD.t381 GND 0.0485f
C5472 VDD.t538 GND 0.0199f
C5473 VDD.t651 GND 0.0209f
C5474 VDD.t289 GND 0.0209f
C5475 VDD.t451 GND 0.0241f
C5476 VDD.t498 GND 0.0392f
C5477 VDD.n1144 GND 0.0192f
C5478 VDD.n1170 GND 0.0309f
C5479 VDD.n1172 GND 0.013f
C5480 VDD.n1177 GND 0.0119f
C5481 VDD.n1178 GND 0.119f
C5482 VDD.n1179 GND 0.593f
C5483 VDD.n1180 GND 3.2f
C5484 VDD.n1181 GND 4.85f
C5485 VDD.n1182 GND 0.0114f
C5486 VDD.n1185 GND 0.0124f
C5487 VDD.n1190 GND 0.0138f
C5488 VDD.n1191 GND 0.0561f
C5489 VDD.n1197 GND 0.0124f
C5490 VDD.n1198 GND 0.0124f
C5491 VDD.n1203 GND 0.0323f
C5492 VDD.n1236 GND 0.0239f
C5493 VDD.t606 GND 0.0103f
C5494 VDD.t807 GND 0.0258f
C5495 VDD.t534 GND 0.0248f
C5496 VDD.t578 GND 0.0302f
C5497 VDD.t1282 GND 0.026f
C5498 VDD.t1005 GND 0.0225f
C5499 VDD.t577 GND 0.0188f
C5500 VDD.t403 GND 0.0298f
C5501 VDD.t258 GND 0.026f
C5502 VDD.t1426 GND 0.0225f
C5503 VDD.t837 GND 0.0225f
C5504 VDD.t428 GND 0.0215f
C5505 VDD.t969 GND 0.0231f
C5506 VDD.t1374 GND 0.0229f
C5507 VDD.t1360 GND 0.0231f
C5508 VDD.t1311 GND 0.0231f
C5509 VDD.t798 GND 0.0291f
C5510 VDD.n1240 GND 0.0705f
C5511 VDD.n1244 GND 0.0196f
C5512 VDD.n1245 GND 0.599f
C5513 VDD.n1246 GND 0.414f
C5514 VDD.n1249 GND 0.0195f
C5515 VDD.n1251 GND 0.133f
C5516 VDD.n1255 GND 0.0281f
C5517 VDD.n1270 GND 0.03f
C5518 VDD.n1274 GND 0.0493f
C5519 VDD.n1276 GND 0.0493f
C5520 VDD.n1280 GND 0.0493f
C5521 VDD.n1282 GND 0.0493f
C5522 VDD.n1283 GND 0.146f
C5523 VDD.n1285 GND 0.0168f
C5524 VDD.t1236 GND 0.0238f
C5525 VDD.t1160 GND 0.0238f
C5526 VDD.t1212 GND 0.0238f
C5527 VDD.t1138 GND 0.0238f
C5528 VDD.t1164 GND 0.0238f
C5529 VDD.t1196 GND 0.0238f
C5530 VDD.t1132 GND 0.0238f
C5531 VDD.t1222 GND 0.0207f
C5532 VDD.n1291 GND 0.0439f
C5533 VDD.n1295 GND 0.0493f
C5534 VDD.n1297 GND 0.0493f
C5535 VDD.n1301 GND 0.0493f
C5536 VDD.n1303 GND 0.0354f
C5537 VDD.n1304 GND 0.091f
C5538 VDD.n1308 GND 0.0131f
C5539 VDD.n1310 GND 0.0168f
C5540 VDD.n1314 GND 0.0154f
C5541 VDD.t1174 GND 0.0238f
C5542 VDD.t1206 GND 0.0238f
C5543 VDD.t1250 GND 0.0238f
C5544 VDD.t1178 GND 0.0227f
C5545 VDD.t312 GND 0.0238f
C5546 VDD.t302 GND 0.0238f
C5547 VDD.t324 GND 0.0238f
C5548 VDD.t318 GND 0.0125f
C5549 VDD.n1325 GND 0.012f
C5550 VDD.n1327 GND 0.0119f
C5551 VDD.n1331 GND 0.0168f
C5552 VDD.n1333 GND 0.0168f
C5553 VDD.n1337 GND 0.0168f
C5554 VDD.n1339 GND 0.0168f
C5555 VDD.n1346 GND 0.0124f
C5556 VDD.t298 GND 0.0238f
C5557 VDD.t308 GND 0.0238f
C5558 VDD.t316 GND 0.0218f
C5559 VDD.n1349 GND 0.0126f
C5560 VDD.n1351 GND 0.0168f
C5561 VDD.n1354 GND 0.0168f
C5562 VDD.n1356 GND 0.0168f
C5563 VDD.n1363 GND 0.0104f
C5564 VDD.n1365 GND 0.011f
C5565 VDD.n1370 GND 0.0105f
C5566 VDD.t1482 GND 0.0295f
C5567 VDD.n1371 GND 0.03f
C5568 VDD.t1278 GND 0.0225f
C5569 VDD.t1274 GND 0.0238f
C5570 VDD.t1272 GND 0.0238f
C5571 VDD.t1276 GND 0.0308f
C5572 VDD.t296 GND 0.013f
C5573 VDD.n1372 GND 0.0178f
C5574 VDD.n1373 GND 0.0105f
C5575 VDD.n1374 GND 0.0101f
C5576 VDD.n1381 GND 0.012f
C5577 VDD.n1383 GND 0.0168f
C5578 VDD.n1387 GND 0.0168f
C5579 VDD.n1389 GND 0.0168f
C5580 VDD.n1393 GND 0.0132f
C5581 VDD.t322 GND 0.0238f
C5582 VDD.t304 GND 0.0238f
C5583 VDD.t314 GND 0.0238f
C5584 VDD.t294 GND 0.0201f
C5585 VDD.t320 GND 0.0238f
C5586 VDD.t306 GND 0.0238f
C5587 VDD.t310 GND 0.0238f
C5588 VDD.t300 GND 0.0156f
C5589 VDD.n1397 GND 0.0178f
C5590 VDD.n1398 GND 0.0105f
C5591 VDD.n1406 GND 0.012f
C5592 VDD.n1410 GND 0.0155f
C5593 VDD.n1412 GND 0.0168f
C5594 VDD.n1416 GND 0.0168f
C5595 VDD.n1418 GND 0.0168f
C5596 VDD.n1422 GND 0.0138f
C5597 VDD.n1427 GND 0.0105f
C5598 VDD.n1428 GND 0.0249f
C5599 VDD.t1244 GND 0.023f
C5600 VDD.t1166 GND 0.0238f
C5601 VDD.t1140 GND 0.0238f
C5602 VDD.t1194 GND 0.0238f
C5603 VDD.t1162 GND 0.0238f
C5604 VDD.t1136 GND 0.0238f
C5605 VDD.t1210 GND 0.013f
C5606 VDD.n1429 GND 0.0178f
C5607 VDD.n1430 GND 0.0105f
C5608 VDD.n1433 GND 0.0161f
C5609 VDD.n1437 GND 0.0168f
C5610 VDD.n1441 GND 0.0168f
C5611 VDD.n1443 GND 0.0168f
C5612 VDD.n1447 GND 0.0168f
C5613 VDD.n1449 GND 0.0168f
C5614 VDD.n1453 GND 0.0173f
C5615 VDD.n1455 GND 0.0105f
C5616 VDD.t1246 GND 0.0238f
C5617 VDD.t1150 GND 0.0238f
C5618 VDD.t1228 GND 0.0238f
C5619 VDD.t1198 GND 0.0184f
C5620 VDD.n1456 GND 0.0178f
C5621 VDD.t1146 GND 0.0244f
C5622 VDD.t1220 GND 0.023f
C5623 VDD.t1168 GND 0.0238f
C5624 VDD.t1142 GND 0.0365f
C5625 VDD.t1216 GND 0.0523f
C5626 VDD.t1184 GND 0.0528f
C5627 VDD.t1124 GND 0.0528f
C5628 VDD.t1158 GND 0.0528f
C5629 VDD.t1126 GND 0.0528f
C5630 VDD.t1190 GND 0.0528f
C5631 VDD.t1154 GND 0.0528f
C5632 VDD.t1232 GND 0.0528f
C5633 VDD.t1204 GND 0.0528f
C5634 VDD.t1172 GND 0.0528f
C5635 VDD.t1242 GND 0.0531f
C5636 VDD.t1200 GND 0.0239f
C5637 VDD.t1128 GND 0.0309f
C5638 VDD.n1457 GND 0.017f
C5639 VDD.n1458 GND 0.0105f
C5640 VDD.n1463 GND 0.0105f
C5641 VDD.n1467 GND 0.0168f
C5642 VDD.n1469 GND 0.0168f
C5643 VDD.n1473 GND 0.0168f
C5644 VDD.n1475 GND 0.0168f
C5645 VDD.n1479 GND 0.0168f
C5646 VDD.n1481 GND 0.0168f
C5647 VDD.n1485 GND 0.0168f
C5648 VDD.n1489 GND 0.0168f
C5649 VDD.n1491 GND 0.0168f
C5650 VDD.n1495 GND 0.0168f
C5651 VDD.n1497 GND 0.0168f
C5652 VDD.n1501 GND 0.0168f
C5653 VDD.n1503 GND 0.0153f
C5654 VDD.n1504 GND 0.012f
C5655 VDD.t1240 GND 0.0547f
C5656 VDD.t1130 GND 0.0238f
C5657 VDD.t1202 GND 0.0238f
C5658 VDD.t1230 GND 0.0238f
C5659 VDD.t1152 GND 0.0238f
C5660 VDD.t1188 GND 0.0238f
C5661 VDD.t1234 GND 0.0238f
C5662 VDD.t1156 GND 0.0238f
C5663 VDD.t1192 GND 0.0238f
C5664 VDD.t1180 GND 0.0238f
C5665 VDD.t1214 GND 0.0238f
C5666 VDD.t1238 GND 0.0238f
C5667 VDD.t1186 GND 0.0238f
C5668 VDD.t1218 GND 0.0238f
C5669 VDD.t1144 GND 0.0238f
C5670 VDD.t1170 GND 0.023f
C5671 VDD.t1208 GND 0.0238f
C5672 VDD.t1176 GND 0.0238f
C5673 VDD.t1248 GND 0.0238f
C5674 VDD.t1224 GND 0.0238f
C5675 VDD.t1134 GND 0.0238f
C5676 VDD.t1182 GND 0.0238f
C5677 VDD.t1148 GND 0.0238f
C5678 VDD.t1226 GND 0.0286f
C5679 VDD.n1507 GND 0.0249f
C5680 VDD.n1508 GND 0.0105f
C5681 VDD.n1513 GND 0.0134f
C5682 VDD.n1517 GND 0.0168f
C5683 VDD.n1519 GND 0.0168f
C5684 VDD.n1523 GND 0.0168f
C5685 VDD.n1526 GND 0.12f
C5686 VDD.n1527 GND 0.0341f
C5687 VDD.n1529 GND 0.0364f
C5688 VDD.n1533 GND 0.0364f
C5689 VDD.n1537 GND 0.0364f
C5690 VDD.n1539 GND 0.0265f
C5691 VDD.n1540 GND 0.407f
C5692 VDD.t536 GND 0.0326f
C5693 VDD.n1541 GND 0.0471f
C5694 VDD.n1548 GND 0.116f
C5695 VDD.t1013 GND 0.0126f
C5696 VDD.t788 GND 0.0121f
C5697 VDD.t1303 GND 0.0106f
C5698 VDD.t1359 GND 0.0134f
C5699 VDD.t539 GND 0.0121f
C5700 VDD.t823 GND 0.0169f
C5701 VDD.t1491 GND 0.0466f
C5702 VDD.n1564 GND 0.0153f
C5703 VDD.n1565 GND 0.257f
C5704 VDD.t290 GND 0.0452f
C5705 VDD.t649 GND 0.0156f
C5706 VDD.t791 GND 0.0346f
C5707 VDD.t1119 GND 0.0646f
C5708 VDD.t509 GND 0.0275f
C5709 VDD.n1566 GND 0.0207f
C5710 VDD.n1595 GND 0.0116f
C5711 VDD.n1596 GND 0.16f
C5712 VDD.n1597 GND 0.601f
C5713 VDD.n1598 GND 0.581f
C5714 VDD.n1599 GND 0.446f
C5715 VDD.n1600 GND 3.26f
C5716 VDD.n1601 GND 2.59f
C5717 VDD.n1602 GND 4.7f
C5718 VDD.n1603 GND 13.5f
C5719 VDD.n1613 GND 0.0244f
C5720 VDD.n1622 GND 0.0743f
C5721 VDD.n1623 GND 0.0594f
C5722 VDD.n1642 GND 0.046f
C5723 VDD.n1646 GND 0.0396f
C5724 VDD.n1652 GND 0.0351f
C5725 VDD.n1653 GND 0.156f
C5726 VDD.n1654 GND 0.13f
C5727 VDD.n1655 GND 0.0932f
C5728 VDD.n1656 GND 0.12f
C5729 VDD.n1657 GND 0.148f
C5730 VDD.n1658 GND 0.146f
C5731 VDD.n1659 GND 0.133f
C5732 VDD.n1660 GND 0.152f
C5733 VDD.n1661 GND 0.114f
C5734 VDD.n1662 GND 0.299f
C5735 VDD.n1663 GND 11.5f
C5736 VDD.n1664 GND 0.275f
C5737 VDD.n1665 GND 0.0237f
C5738 VDD.n1666 GND 0.0462f
C5739 VDD.t1031 GND 0.0597f
C5740 VDD.n1678 GND 0.0351f
C5741 VDD.n1686 GND 0.0437f
C5742 VDD.n1687 GND 0.0152f
C5743 VDD.n1688 GND 0.0128f
C5744 VDD.n1695 GND 0.0504f
C5745 VDD.n1711 GND 0.0735f
C5746 VDD.t441 GND 0.0597f
C5747 VDD.n1712 GND 0.0351f
C5748 VDD.n1721 GND 0.0491f
C5749 VDD.n1723 GND 0.0135f
C5750 VDD.n1737 GND 0.0484f
C5751 VDD.n1738 GND 0.0582f
C5752 VDD.n1744 GND 0.0584f
C5753 VDD.n1748 GND 0.0134f
C5754 VDD.n1749 GND 0.047f
C5755 VDD.n1753 GND 0.0289f
C5756 VDD.n1754 GND 0.0135f
C5757 VDD.t1014 GND 0.169f
C5758 VDD.n1764 GND 0.0735f
C5759 VDD.n1770 GND 0.0135f
C5760 VDD.n1771 GND 0.0287f
C5761 VDD.n1773 GND 0.0248f
C5762 VDD.n1774 GND 0.13f
C5763 VDD.n1775 GND 0.427f
C5764 VDD.n1801 GND 0.0444f
C5765 VDD.t443 GND 0.0187f
C5766 VDD.n1802 GND 0.0194f
C5767 VDD.n1803 GND 0.0239f
C5768 VDD.t1028 GND 0.0185f
C5769 VDD.n1804 GND 0.16f
C5770 VDD.n1805 GND 0.967f
C5771 VDD.n1806 GND 0.103f
C5772 VDD.n1807 GND 1.15f
C5773 VDD.n1808 GND 0.921f
C5774 VDD.t1498 GND 0.0383f
C5775 VDD.t464 GND 0.0134f
C5776 VDD.n1809 GND 0.0699f
C5777 VDD.n1816 GND 0.058f
C5778 VDD.n1817 GND 0.0223f
C5779 VDD.n1821 GND 0.0683f
C5780 VDD.n1823 GND 0.078f
C5781 VDD.n1825 GND 0.0106f
C5782 VDD.t1088 GND 0.0288f
C5783 VDD.t599 GND 0.0109f
C5784 VDD.n1836 GND 0.0397f
C5785 VDD.n1839 GND 0.0201f
C5786 VDD.n1840 GND 0.0133f
C5787 VDD.n1841 GND 0.114f
C5788 VDD.n1842 GND 0.0382f
C5789 VDD.n1847 GND 0.0681f
C5790 VDD.n1849 GND 0.0899f
C5791 VDD.n1857 GND 0.0866f
C5792 VDD.n1858 GND 0.0386f
C5793 VDD.n1863 GND 0.0419f
C5794 VDD.t466 GND 0.0681f
C5795 VDD.n1872 GND 0.295f
C5796 VDD.n1873 GND 0.165f
C5797 VDD.n1874 GND 0.0664f
C5798 VDD.n1875 GND 0.0216f
C5799 VDD.t274 GND 0.0856f
C5800 VDD.n1886 GND 0.0455f
C5801 VDD.n1887 GND 0.112f
C5802 VDD.n1889 GND 0.0121f
C5803 VDD.n1892 GND 0.0858f
C5804 VDD.n1893 GND 0.0899f
C5805 VDD.n1901 GND 0.0427f
C5806 VDD.n1905 GND 0.0386f
C5807 VDD.t277 GND 0.0681f
C5808 VDD.n1914 GND 0.0681f
C5809 VDD.n1916 GND 0.0876f
C5810 VDD.n1917 GND 0.28f
C5811 VDD.n1918 GND 0.166f
C5812 VDD.n1919 GND 0.196f
C5813 VDD.n1920 GND 0.0783f
C5814 VDD.n1921 GND 6.12f
C5815 VDD.n1922 GND 0.159f
C5816 VDD.n1923 GND 0.138f
C5817 VDD.t1027 GND 0.0214f
C5818 VDD.t1039 GND 0.0214f
C5819 VDD.n1924 GND 0.326f
C5820 VDD.n1925 GND 0.0174f
C5821 VDD.n1926 GND 0.0127f
C5822 VDD.n1927 GND 0.4f
C5823 VDD.n1930 GND 0.0303f
C5824 VDD.n1931 GND 0.317f
C5825 VDD.n1933 GND 0.127f
C5826 VDD.n1935 GND 0.0135f
C5827 VDD.n1939 GND 0.2f
C5828 VDD.n1940 GND 0.0135f
C5829 VDD.n1942 GND 0.0303f
C5830 VDD.n1943 GND 0.0182f
C5831 VDD.t1037 GND 0.0214f
C5832 VDD.n1945 GND 0.163f
C5833 VDD.n1946 GND 0.0852f
C5834 VDD.n1948 GND 0.0135f
C5835 VDD.n1949 GND 0.317f
C5836 VDD.n1950 GND 0.0169f
C5837 VDD.n1951 GND 0.0169f
C5838 VDD.t1036 GND 0.399f
C5839 VDD.n1952 GND 0.014f
C5840 VDD.n1953 GND 0.2f
C5841 VDD.n1954 GND 0.0127f
C5842 VDD.n1955 GND 0.0127f
C5843 VDD.n1957 GND 0.0884f
C5844 VDD.n1960 GND 0.0169f
C5845 VDD.n1961 GND 0.0169f
C5846 VDD.t1026 GND 0.387f
C5847 VDD.n1967 GND 0.0169f
C5848 VDD.n1968 GND 0.0169f
C5849 VDD.t1038 GND 0.4f
C5850 VDD.n1970 GND 0.0169f
C5851 VDD.n1971 GND 0.0169f
C5852 VDD.n1974 GND 0.0135f
C5853 VDD.n1976 GND 0.0127f
C5854 VDD.n1979 GND 0.202f
C5855 VDD.n1980 GND 0.127f
C5856 VDD.n1981 GND 0.0329f
C5857 VDD.n1982 GND 9.56f
C5858 VDD.n1983 GND 0.275f
C5859 VDD.n2009 GND 0.0444f
C5860 VDD.t77 GND 0.0187f
C5861 VDD.n2010 GND 0.0194f
C5862 VDD.n2011 GND 0.0239f
C5863 VDD.t1266 GND 0.0185f
C5864 VDD.n2012 GND 0.612f
C5865 VDD.n2013 GND 0.462f
C5866 VDD.n2014 GND 0.0237f
C5867 VDD.n2015 GND 0.0462f
C5868 VDD.t1264 GND 0.0597f
C5869 VDD.n2027 GND 0.0351f
C5870 VDD.n2035 GND 0.0437f
C5871 VDD.n2036 GND 0.0152f
C5872 VDD.n2037 GND 0.0128f
C5873 VDD.n2044 GND 0.0504f
C5874 VDD.n2060 GND 0.0735f
C5875 VDD.t80 GND 0.0597f
C5876 VDD.n2061 GND 0.0351f
C5877 VDD.n2070 GND 0.0491f
C5878 VDD.n2072 GND 0.0135f
C5879 VDD.n2086 GND 0.0484f
C5880 VDD.n2087 GND 0.0582f
C5881 VDD.n2093 GND 0.0584f
C5882 VDD.n2097 GND 0.0134f
C5883 VDD.n2098 GND 0.047f
C5884 VDD.n2102 GND 0.0289f
C5885 VDD.n2103 GND 0.0135f
C5886 VDD.t623 GND 0.169f
C5887 VDD.n2113 GND 0.0735f
C5888 VDD.n2119 GND 0.0135f
C5889 VDD.n2120 GND 0.0287f
C5890 VDD.n2122 GND 0.0248f
C5891 VDD.n2123 GND 0.13f
C5892 VDD.n2124 GND 0.427f
C5893 VDD.n2125 GND 0.0484f
C5894 VDD.n2126 GND 0.103f
C5895 VDD.n2127 GND 0.584f
C5896 VDD.n2128 GND 1.1f
C5897 VDD.n2129 GND 0.436f
C5898 VDD.t625 GND 0.0383f
C5899 VDD.t255 GND 0.0134f
C5900 VDD.n2130 GND 0.0699f
C5901 VDD.n2137 GND 0.058f
C5902 VDD.n2138 GND 0.0223f
C5903 VDD.n2142 GND 0.0683f
C5904 VDD.n2144 GND 0.078f
C5905 VDD.n2146 GND 0.0106f
C5906 VDD.t555 GND 0.0288f
C5907 VDD.t1011 GND 0.0109f
C5908 VDD.n2157 GND 0.0397f
C5909 VDD.n2160 GND 0.0201f
C5910 VDD.n2161 GND 0.0133f
C5911 VDD.n2162 GND 0.114f
C5912 VDD.n2163 GND 0.0382f
C5913 VDD.n2168 GND 0.0681f
C5914 VDD.n2170 GND 0.0899f
C5915 VDD.n2178 GND 0.0866f
C5916 VDD.n2179 GND 0.0386f
C5917 VDD.n2184 GND 0.0419f
C5918 VDD.t592 GND 0.0681f
C5919 VDD.n2193 GND 0.295f
C5920 VDD.n2194 GND 0.165f
C5921 VDD.n2195 GND 0.0664f
C5922 VDD.n2196 GND 0.0216f
C5923 VDD.t511 GND 0.0856f
C5924 VDD.n2207 GND 0.0455f
C5925 VDD.n2208 GND 0.112f
C5926 VDD.n2210 GND 0.0121f
C5927 VDD.n2213 GND 0.0858f
C5928 VDD.n2214 GND 0.0899f
C5929 VDD.n2222 GND 0.0427f
C5930 VDD.n2226 GND 0.0386f
C5931 VDD.t494 GND 0.0681f
C5932 VDD.n2235 GND 0.0681f
C5933 VDD.n2237 GND 0.0876f
C5934 VDD.n2238 GND 0.28f
C5935 VDD.n2239 GND 0.166f
C5936 VDD.n2240 GND 0.196f
C5937 VDD.n2241 GND 0.0783f
C5938 VDD.n2242 GND 6.12f
C5939 VDD.n2243 GND 0.275f
C5940 VDD.n2244 GND 0.0237f
C5941 VDD.n2245 GND 0.0462f
C5942 VDD.t831 GND 0.0597f
C5943 VDD.n2257 GND 0.0351f
C5944 VDD.n2265 GND 0.0437f
C5945 VDD.n2266 GND 0.0152f
C5946 VDD.n2267 GND 0.0128f
C5947 VDD.n2274 GND 0.0504f
C5948 VDD.n2290 GND 0.0735f
C5949 VDD.t1446 GND 0.0597f
C5950 VDD.n2291 GND 0.0351f
C5951 VDD.n2300 GND 0.0491f
C5952 VDD.n2302 GND 0.0135f
C5953 VDD.n2316 GND 0.0484f
C5954 VDD.n2317 GND 0.0582f
C5955 VDD.n2323 GND 0.0584f
C5956 VDD.n2327 GND 0.0134f
C5957 VDD.n2328 GND 0.047f
C5958 VDD.n2332 GND 0.0289f
C5959 VDD.n2333 GND 0.0135f
C5960 VDD.t1331 GND 0.169f
C5961 VDD.n2343 GND 0.0735f
C5962 VDD.n2349 GND 0.0135f
C5963 VDD.n2350 GND 0.0287f
C5964 VDD.n2352 GND 0.0248f
C5965 VDD.n2353 GND 0.13f
C5966 VDD.n2354 GND 0.427f
C5967 VDD.n2380 GND 0.0444f
C5968 VDD.t1444 GND 0.0187f
C5969 VDD.n2381 GND 0.0194f
C5970 VDD.n2382 GND 0.0239f
C5971 VDD.t828 GND 0.0185f
C5972 VDD.n2383 GND 0.16f
C5973 VDD.n2384 GND 0.967f
C5974 VDD.n2385 GND 0.103f
C5975 VDD.n2386 GND 1.15f
C5976 VDD.n2387 GND 0.921f
C5977 VDD.t1284 GND 0.0383f
C5978 VDD.t1017 GND 0.0134f
C5979 VDD.n2388 GND 0.0699f
C5980 VDD.n2395 GND 0.058f
C5981 VDD.n2396 GND 0.0223f
C5982 VDD.n2400 GND 0.0683f
C5983 VDD.n2402 GND 0.078f
C5984 VDD.n2404 GND 0.0106f
C5985 VDD.t1383 GND 0.0288f
C5986 VDD.t615 GND 0.0109f
C5987 VDD.n2415 GND 0.0397f
C5988 VDD.n2418 GND 0.0201f
C5989 VDD.n2419 GND 0.0133f
C5990 VDD.n2420 GND 0.114f
C5991 VDD.n2421 GND 0.0382f
C5992 VDD.n2426 GND 0.0681f
C5993 VDD.n2428 GND 0.0899f
C5994 VDD.n2436 GND 0.0866f
C5995 VDD.n2437 GND 0.0386f
C5996 VDD.n2442 GND 0.0419f
C5997 VDD.t521 GND 0.0681f
C5998 VDD.n2451 GND 0.295f
C5999 VDD.n2452 GND 0.165f
C6000 VDD.n2453 GND 0.0664f
C6001 VDD.n2454 GND 0.0216f
C6002 VDD.t528 GND 0.0856f
C6003 VDD.n2465 GND 0.0455f
C6004 VDD.n2466 GND 0.112f
C6005 VDD.n2468 GND 0.0121f
C6006 VDD.n2471 GND 0.0858f
C6007 VDD.n2472 GND 0.0899f
C6008 VDD.n2480 GND 0.0427f
C6009 VDD.n2484 GND 0.0386f
C6010 VDD.t505 GND 0.0681f
C6011 VDD.n2493 GND 0.0681f
C6012 VDD.n2495 GND 0.0876f
C6013 VDD.n2496 GND 0.28f
C6014 VDD.n2497 GND 0.166f
C6015 VDD.n2498 GND 0.196f
C6016 VDD.n2499 GND 0.0783f
C6017 VDD.n2500 GND 6.12f
C6018 VDD.n2501 GND 0.275f
C6019 VDD.n2502 GND 0.0237f
C6020 VDD.n2503 GND 0.0462f
C6021 VDD.t1417 GND 0.0597f
C6022 VDD.n2515 GND 0.0351f
C6023 VDD.n2523 GND 0.0437f
C6024 VDD.n2524 GND 0.0152f
C6025 VDD.n2525 GND 0.0128f
C6026 VDD.n2532 GND 0.0504f
C6027 VDD.n2548 GND 0.0735f
C6028 VDD.t567 GND 0.0597f
C6029 VDD.n2549 GND 0.0351f
C6030 VDD.n2558 GND 0.0491f
C6031 VDD.n2560 GND 0.0135f
C6032 VDD.n2574 GND 0.0484f
C6033 VDD.n2575 GND 0.0582f
C6034 VDD.n2581 GND 0.0584f
C6035 VDD.n2585 GND 0.0134f
C6036 VDD.n2586 GND 0.047f
C6037 VDD.n2590 GND 0.0289f
C6038 VDD.n2591 GND 0.0135f
C6039 VDD.t825 GND 0.169f
C6040 VDD.n2601 GND 0.0735f
C6041 VDD.n2607 GND 0.0135f
C6042 VDD.n2608 GND 0.0287f
C6043 VDD.n2610 GND 0.0248f
C6044 VDD.n2611 GND 0.13f
C6045 VDD.n2612 GND 0.427f
C6046 VDD.n2638 GND 0.0444f
C6047 VDD.t569 GND 0.0187f
C6048 VDD.n2639 GND 0.0194f
C6049 VDD.n2640 GND 0.0239f
C6050 VDD.t1419 GND 0.0185f
C6051 VDD.n2641 GND 0.16f
C6052 VDD.n2642 GND 0.967f
C6053 VDD.n2643 GND 0.103f
C6054 VDD.n2644 GND 1.15f
C6055 VDD.n2645 GND 0.921f
C6056 VDD.t85 GND 0.0383f
C6057 VDD.t1323 GND 0.0134f
C6058 VDD.n2646 GND 0.0699f
C6059 VDD.n2653 GND 0.058f
C6060 VDD.n2654 GND 0.0223f
C6061 VDD.n2658 GND 0.0683f
C6062 VDD.n2660 GND 0.078f
C6063 VDD.n2662 GND 0.0106f
C6064 VDD.t575 GND 0.0288f
C6065 VDD.t247 GND 0.0109f
C6066 VDD.n2673 GND 0.0397f
C6067 VDD.n2676 GND 0.0201f
C6068 VDD.n2677 GND 0.0133f
C6069 VDD.n2678 GND 0.114f
C6070 VDD.n2679 GND 0.0382f
C6071 VDD.n2684 GND 0.0681f
C6072 VDD.n2686 GND 0.0899f
C6073 VDD.n2694 GND 0.0866f
C6074 VDD.n2695 GND 0.0386f
C6075 VDD.n2700 GND 0.0419f
C6076 VDD.t278 GND 0.0681f
C6077 VDD.n2709 GND 0.295f
C6078 VDD.n2710 GND 0.165f
C6079 VDD.n2711 GND 0.0664f
C6080 VDD.n2712 GND 0.0216f
C6081 VDD.t1381 GND 0.0856f
C6082 VDD.n2723 GND 0.0455f
C6083 VDD.n2724 GND 0.112f
C6084 VDD.n2726 GND 0.0121f
C6085 VDD.n2729 GND 0.0858f
C6086 VDD.n2730 GND 0.0899f
C6087 VDD.n2738 GND 0.0427f
C6088 VDD.n2742 GND 0.0386f
C6089 VDD.t1023 GND 0.0681f
C6090 VDD.n2751 GND 0.0681f
C6091 VDD.n2753 GND 0.0876f
C6092 VDD.n2754 GND 0.28f
C6093 VDD.n2755 GND 0.166f
C6094 VDD.n2756 GND 0.196f
C6095 VDD.n2757 GND 0.0783f
C6096 VDD.n2758 GND 6.12f
C6097 VDD.n2759 GND 0.275f
C6098 VDD.n2760 GND 0.0237f
C6099 VDD.n2761 GND 0.0462f
C6100 VDD.t436 GND 0.0597f
C6101 VDD.n2773 GND 0.0351f
C6102 VDD.n2781 GND 0.0437f
C6103 VDD.n2782 GND 0.0152f
C6104 VDD.n2783 GND 0.0128f
C6105 VDD.n2790 GND 0.0504f
C6106 VDD.n2806 GND 0.0735f
C6107 VDD.t978 GND 0.0597f
C6108 VDD.n2807 GND 0.0351f
C6109 VDD.n2816 GND 0.0491f
C6110 VDD.n2818 GND 0.0135f
C6111 VDD.n2832 GND 0.0484f
C6112 VDD.n2833 GND 0.0582f
C6113 VDD.n2839 GND 0.0584f
C6114 VDD.n2843 GND 0.0134f
C6115 VDD.n2844 GND 0.047f
C6116 VDD.n2848 GND 0.0289f
C6117 VDD.n2849 GND 0.0135f
C6118 VDD.t424 GND 0.169f
C6119 VDD.n2859 GND 0.0735f
C6120 VDD.n2865 GND 0.0135f
C6121 VDD.n2866 GND 0.0287f
C6122 VDD.n2868 GND 0.0248f
C6123 VDD.n2869 GND 0.13f
C6124 VDD.n2870 GND 0.427f
C6125 VDD.n2896 GND 0.0444f
C6126 VDD.t976 GND 0.0187f
C6127 VDD.n2897 GND 0.0194f
C6128 VDD.n2898 GND 0.0239f
C6129 VDD.t433 GND 0.0185f
C6130 VDD.n2899 GND 0.16f
C6131 VDD.n2900 GND 0.967f
C6132 VDD.n2901 GND 0.103f
C6133 VDD.n2902 GND 1.15f
C6134 VDD.n2903 GND 0.921f
C6135 VDD.t272 GND 0.0383f
C6136 VDD.t366 GND 0.0134f
C6137 VDD.n2904 GND 0.0699f
C6138 VDD.n2911 GND 0.058f
C6139 VDD.n2912 GND 0.0223f
C6140 VDD.n2916 GND 0.0683f
C6141 VDD.n2918 GND 0.078f
C6142 VDD.n2920 GND 0.0106f
C6143 VDD.t1479 GND 0.0288f
C6144 VDD.t618 GND 0.0109f
C6145 VDD.n2931 GND 0.0397f
C6146 VDD.n2934 GND 0.0201f
C6147 VDD.n2935 GND 0.0133f
C6148 VDD.n2936 GND 0.114f
C6149 VDD.n2937 GND 0.0382f
C6150 VDD.n2942 GND 0.0681f
C6151 VDD.n2944 GND 0.0899f
C6152 VDD.n2952 GND 0.0866f
C6153 VDD.n2953 GND 0.0386f
C6154 VDD.n2958 GND 0.0419f
C6155 VDD.t368 GND 0.0681f
C6156 VDD.n2967 GND 0.295f
C6157 VDD.n2968 GND 0.165f
C6158 VDD.n2969 GND 0.0664f
C6159 VDD.n2970 GND 0.0216f
C6160 VDD.t414 GND 0.0856f
C6161 VDD.n2981 GND 0.0455f
C6162 VDD.n2982 GND 0.112f
C6163 VDD.n2984 GND 0.0121f
C6164 VDD.n2987 GND 0.0858f
C6165 VDD.n2988 GND 0.0899f
C6166 VDD.n2996 GND 0.0427f
C6167 VDD.n3000 GND 0.0386f
C6168 VDD.t524 GND 0.0681f
C6169 VDD.n3009 GND 0.0681f
C6170 VDD.n3011 GND 0.0876f
C6171 VDD.n3012 GND 0.28f
C6172 VDD.n3013 GND 0.166f
C6173 VDD.n3014 GND 0.196f
C6174 VDD.n3015 GND 0.0783f
C6175 VDD.n3016 GND 6.12f
C6176 VDD.n3017 GND 0.275f
C6177 VDD.n3018 GND 0.0237f
C6178 VDD.n3019 GND 0.0462f
C6179 VDD.t383 GND 0.0597f
C6180 VDD.n3031 GND 0.0351f
C6181 VDD.n3039 GND 0.0437f
C6182 VDD.n3040 GND 0.0152f
C6183 VDD.n3041 GND 0.0128f
C6184 VDD.n3048 GND 0.0504f
C6185 VDD.n3064 GND 0.0735f
C6186 VDD.t545 GND 0.0597f
C6187 VDD.n3065 GND 0.0351f
C6188 VDD.n3074 GND 0.0491f
C6189 VDD.n3076 GND 0.0135f
C6190 VDD.n3090 GND 0.0484f
C6191 VDD.n3091 GND 0.0582f
C6192 VDD.n3097 GND 0.0584f
C6193 VDD.n3101 GND 0.0134f
C6194 VDD.n3102 GND 0.047f
C6195 VDD.n3106 GND 0.0289f
C6196 VDD.n3107 GND 0.0135f
C6197 VDD.t395 GND 0.169f
C6198 VDD.n3117 GND 0.0735f
C6199 VDD.n3123 GND 0.0135f
C6200 VDD.n3124 GND 0.0287f
C6201 VDD.n3126 GND 0.0248f
C6202 VDD.n3127 GND 0.13f
C6203 VDD.n3128 GND 0.427f
C6204 VDD.n3154 GND 0.0444f
C6205 VDD.t543 GND 0.0187f
C6206 VDD.n3155 GND 0.0194f
C6207 VDD.n3156 GND 0.0239f
C6208 VDD.t385 GND 0.0185f
C6209 VDD.n3157 GND 0.16f
C6210 VDD.n3158 GND 0.967f
C6211 VDD.n3159 GND 0.103f
C6212 VDD.n3160 GND 1.15f
C6213 VDD.n3161 GND 0.921f
C6214 VDD.t541 GND 0.0383f
C6215 VDD.t1459 GND 0.0134f
C6216 VDD.n3162 GND 0.0699f
C6217 VDD.n3169 GND 0.058f
C6218 VDD.n3170 GND 0.0223f
C6219 VDD.n3174 GND 0.0683f
C6220 VDD.n3176 GND 0.078f
C6221 VDD.n3178 GND 0.0106f
C6222 VDD.t1003 GND 0.0288f
C6223 VDD.t647 GND 0.0109f
C6224 VDD.n3189 GND 0.0397f
C6225 VDD.n3192 GND 0.0201f
C6226 VDD.n3193 GND 0.0133f
C6227 VDD.n3194 GND 0.114f
C6228 VDD.n3195 GND 0.0382f
C6229 VDD.n3200 GND 0.0681f
C6230 VDD.n3202 GND 0.0899f
C6231 VDD.n3210 GND 0.0866f
C6232 VDD.n3211 GND 0.0386f
C6233 VDD.n3216 GND 0.0419f
C6234 VDD.t1087 GND 0.0681f
C6235 VDD.n3225 GND 0.295f
C6236 VDD.n3226 GND 0.165f
C6237 VDD.n3227 GND 0.0664f
C6238 VDD.n3228 GND 0.0216f
C6239 VDD.t591 GND 0.0856f
C6240 VDD.n3239 GND 0.0455f
C6241 VDD.n3240 GND 0.112f
C6242 VDD.n3242 GND 0.0121f
C6243 VDD.n3245 GND 0.0858f
C6244 VDD.n3246 GND 0.0899f
C6245 VDD.n3254 GND 0.0427f
C6246 VDD.n3258 GND 0.0386f
C6247 VDD.t282 GND 0.0681f
C6248 VDD.n3267 GND 0.0681f
C6249 VDD.n3269 GND 0.0876f
C6250 VDD.n3270 GND 0.28f
C6251 VDD.n3271 GND 0.166f
C6252 VDD.n3272 GND 0.196f
C6253 VDD.n3273 GND 0.0783f
C6254 VDD.n3274 GND 6.12f
C6255 VDD.n3275 GND 0.275f
C6256 VDD.n3276 GND 0.0237f
C6257 VDD.n3277 GND 0.0462f
C6258 VDD.t1295 GND 0.0597f
C6259 VDD.n3289 GND 0.0351f
C6260 VDD.n3297 GND 0.0437f
C6261 VDD.n3298 GND 0.0152f
C6262 VDD.n3299 GND 0.0128f
C6263 VDD.n3306 GND 0.0504f
C6264 VDD.n3322 GND 0.0735f
C6265 VDD.t582 GND 0.0597f
C6266 VDD.n3323 GND 0.0351f
C6267 VDD.n3332 GND 0.0491f
C6268 VDD.n3334 GND 0.0135f
C6269 VDD.n3348 GND 0.0484f
C6270 VDD.n3349 GND 0.0582f
C6271 VDD.n3355 GND 0.0584f
C6272 VDD.n3359 GND 0.0134f
C6273 VDD.n3360 GND 0.047f
C6274 VDD.n3364 GND 0.0289f
C6275 VDD.n3365 GND 0.0135f
C6276 VDD.t639 GND 0.169f
C6277 VDD.n3375 GND 0.0735f
C6278 VDD.n3381 GND 0.0135f
C6279 VDD.n3382 GND 0.0287f
C6280 VDD.n3384 GND 0.0248f
C6281 VDD.n3385 GND 0.13f
C6282 VDD.n3386 GND 0.427f
C6283 VDD.n3412 GND 0.0444f
C6284 VDD.t580 GND 0.0187f
C6285 VDD.n3413 GND 0.0194f
C6286 VDD.n3414 GND 0.0239f
C6287 VDD.t1297 GND 0.0185f
C6288 VDD.n3415 GND 0.16f
C6289 VDD.n3416 GND 0.967f
C6290 VDD.n3417 GND 0.103f
C6291 VDD.n3418 GND 1.15f
C6292 VDD.n3419 GND 0.921f
C6293 VDD.t1280 GND 0.0383f
C6294 VDD.t1293 GND 0.0134f
C6295 VDD.n3420 GND 0.0699f
C6296 VDD.n3427 GND 0.058f
C6297 VDD.n3428 GND 0.0223f
C6298 VDD.n3432 GND 0.0683f
C6299 VDD.n3434 GND 0.078f
C6300 VDD.n3436 GND 0.0106f
C6301 VDD.t397 GND 0.0288f
C6302 VDD.t532 GND 0.0109f
C6303 VDD.n3447 GND 0.0397f
C6304 VDD.n3450 GND 0.0201f
C6305 VDD.n3451 GND 0.0133f
C6306 VDD.n3452 GND 0.114f
C6307 VDD.n3453 GND 0.0382f
C6308 VDD.n3458 GND 0.0681f
C6309 VDD.n3460 GND 0.0899f
C6310 VDD.n3468 GND 0.0866f
C6311 VDD.n3469 GND 0.0386f
C6312 VDD.n3474 GND 0.0419f
C6313 VDD.t1093 GND 0.0681f
C6314 VDD.n3483 GND 0.295f
C6315 VDD.n3484 GND 0.165f
C6316 VDD.n3485 GND 0.0664f
C6317 VDD.n3486 GND 0.0216f
C6318 VDD.t1086 GND 0.0856f
C6319 VDD.n3497 GND 0.0455f
C6320 VDD.n3498 GND 0.112f
C6321 VDD.n3500 GND 0.0121f
C6322 VDD.n3503 GND 0.0858f
C6323 VDD.n3504 GND 0.0899f
C6324 VDD.n3512 GND 0.0427f
C6325 VDD.n3516 GND 0.0386f
C6326 VDD.t419 GND 0.0681f
C6327 VDD.n3525 GND 0.0681f
C6328 VDD.n3527 GND 0.0876f
C6329 VDD.n3528 GND 0.28f
C6330 VDD.n3529 GND 0.166f
C6331 VDD.n3530 GND 0.196f
C6332 VDD.n3531 GND 0.0783f
C6333 VDD.n3532 GND 6.12f
C6334 VDD.n3533 GND 0.275f
C6335 VDD.n3534 GND 0.0237f
C6336 VDD.n3535 GND 0.0462f
C6337 VDD.t1366 GND 0.0597f
C6338 VDD.n3547 GND 0.0351f
C6339 VDD.n3555 GND 0.0437f
C6340 VDD.n3556 GND 0.0152f
C6341 VDD.n3557 GND 0.0128f
C6342 VDD.n3564 GND 0.0504f
C6343 VDD.n3580 GND 0.0735f
C6344 VDD.t1336 GND 0.0597f
C6345 VDD.n3581 GND 0.0351f
C6346 VDD.n3590 GND 0.0491f
C6347 VDD.n3592 GND 0.0135f
C6348 VDD.n3606 GND 0.0484f
C6349 VDD.n3607 GND 0.0582f
C6350 VDD.n3613 GND 0.0584f
C6351 VDD.n3617 GND 0.0134f
C6352 VDD.n3618 GND 0.047f
C6353 VDD.n3622 GND 0.0289f
C6354 VDD.n3623 GND 0.0135f
C6355 VDD.t249 GND 0.169f
C6356 VDD.n3633 GND 0.0735f
C6357 VDD.n3639 GND 0.0135f
C6358 VDD.n3640 GND 0.0287f
C6359 VDD.n3642 GND 0.0248f
C6360 VDD.n3643 GND 0.13f
C6361 VDD.n3644 GND 0.427f
C6362 VDD.n3670 GND 0.0444f
C6363 VDD.t1333 GND 0.0187f
C6364 VDD.n3671 GND 0.0194f
C6365 VDD.n3672 GND 0.0239f
C6366 VDD.t1368 GND 0.0185f
C6367 VDD.n3673 GND 0.16f
C6368 VDD.n3674 GND 0.967f
C6369 VDD.n3675 GND 0.103f
C6370 VDD.n3676 GND 1.15f
C6371 VDD.n3677 GND 0.921f
C6372 VDD.t1101 GND 0.0383f
C6373 VDD.t253 GND 0.0134f
C6374 VDD.n3678 GND 0.0699f
C6375 VDD.n3685 GND 0.058f
C6376 VDD.n3686 GND 0.0223f
C6377 VDD.n3690 GND 0.0683f
C6378 VDD.n3692 GND 0.078f
C6379 VDD.n3694 GND 0.0106f
C6380 VDD.t1070 GND 0.0288f
C6381 VDD.t291 GND 0.0109f
C6382 VDD.n3705 GND 0.0397f
C6383 VDD.n3708 GND 0.0201f
C6384 VDD.n3709 GND 0.0133f
C6385 VDD.n3710 GND 0.114f
C6386 VDD.n3711 GND 0.0382f
C6387 VDD.n3716 GND 0.0681f
C6388 VDD.n3718 GND 0.0899f
C6389 VDD.n3726 GND 0.0866f
C6390 VDD.n3727 GND 0.0386f
C6391 VDD.n3732 GND 0.0419f
C6392 VDD.t251 GND 0.0681f
C6393 VDD.n3741 GND 0.295f
C6394 VDD.n3742 GND 0.165f
C6395 VDD.n3743 GND 0.0664f
C6396 VDD.n3744 GND 0.0216f
C6397 VDD.t1085 GND 0.0856f
C6398 VDD.n3755 GND 0.0455f
C6399 VDD.n3756 GND 0.112f
C6400 VDD.n3758 GND 0.0121f
C6401 VDD.n3761 GND 0.0858f
C6402 VDD.n3762 GND 0.0899f
C6403 VDD.n3770 GND 0.0427f
C6404 VDD.n3774 GND 0.0386f
C6405 VDD.t262 GND 0.0681f
C6406 VDD.n3783 GND 0.0681f
C6407 VDD.n3785 GND 0.0876f
C6408 VDD.n3786 GND 0.28f
C6409 VDD.n3787 GND 0.166f
C6410 VDD.n3788 GND 0.196f
C6411 VDD.n3789 GND 0.0783f
C6412 VDD.n3790 GND 6.12f
C6413 VDD.n3791 GND 0.275f
C6414 VDD.n3792 GND 0.0237f
C6415 VDD.n3793 GND 0.0462f
C6416 VDD.t1114 GND 0.0597f
C6417 VDD.n3805 GND 0.0351f
C6418 VDD.n3813 GND 0.0437f
C6419 VDD.n3814 GND 0.0152f
C6420 VDD.n3815 GND 0.0128f
C6421 VDD.n3822 GND 0.0504f
C6422 VDD.n3838 GND 0.0735f
C6423 VDD.t485 GND 0.0597f
C6424 VDD.n3839 GND 0.0351f
C6425 VDD.n3848 GND 0.0491f
C6426 VDD.n3850 GND 0.0135f
C6427 VDD.n3864 GND 0.0484f
C6428 VDD.n3865 GND 0.0582f
C6429 VDD.n3871 GND 0.0584f
C6430 VDD.n3875 GND 0.0134f
C6431 VDD.n3876 GND 0.047f
C6432 VDD.n3880 GND 0.0289f
C6433 VDD.n3881 GND 0.0135f
C6434 VDD.t1317 GND 0.169f
C6435 VDD.n3891 GND 0.0735f
C6436 VDD.n3897 GND 0.0135f
C6437 VDD.n3898 GND 0.0287f
C6438 VDD.n3900 GND 0.0248f
C6439 VDD.n3901 GND 0.13f
C6440 VDD.n3902 GND 0.427f
C6441 VDD.n3928 GND 0.0444f
C6442 VDD.t483 GND 0.0187f
C6443 VDD.n3929 GND 0.0194f
C6444 VDD.n3930 GND 0.0239f
C6445 VDD.t1111 GND 0.0185f
C6446 VDD.n3931 GND 0.16f
C6447 VDD.n3932 GND 0.967f
C6448 VDD.n3933 GND 0.103f
C6449 VDD.n3934 GND 1.15f
C6450 VDD.n3935 GND 0.921f
C6451 VDD.t1048 GND 0.0383f
C6452 VDD.t268 GND 0.0134f
C6453 VDD.n3936 GND 0.0699f
C6454 VDD.n3943 GND 0.058f
C6455 VDD.n3944 GND 0.0223f
C6456 VDD.n3948 GND 0.0683f
C6457 VDD.n3950 GND 0.078f
C6458 VDD.n3952 GND 0.0106f
C6459 VDD.t1062 GND 0.0288f
C6460 VDD.t1348 GND 0.0109f
C6461 VDD.n3963 GND 0.0397f
C6462 VDD.n3966 GND 0.0201f
C6463 VDD.n3967 GND 0.0133f
C6464 VDD.n3968 GND 0.114f
C6465 VDD.n3969 GND 0.0382f
C6466 VDD.n3974 GND 0.0681f
C6467 VDD.n3976 GND 0.0899f
C6468 VDD.n3984 GND 0.0866f
C6469 VDD.n3985 GND 0.0386f
C6470 VDD.n3990 GND 0.0419f
C6471 VDD.t266 GND 0.0681f
C6472 VDD.n3999 GND 0.295f
C6473 VDD.n4000 GND 0.165f
C6474 VDD.n4001 GND 0.0664f
C6475 VDD.n4002 GND 0.0216f
C6476 VDD.t526 GND 0.0856f
C6477 VDD.n4013 GND 0.0455f
C6478 VDD.n4014 GND 0.112f
C6479 VDD.n4016 GND 0.0121f
C6480 VDD.n4019 GND 0.0858f
C6481 VDD.n4020 GND 0.0899f
C6482 VDD.n4028 GND 0.0427f
C6483 VDD.n4032 GND 0.0386f
C6484 VDD.t1084 GND 0.0681f
C6485 VDD.n4041 GND 0.0681f
C6486 VDD.n4043 GND 0.0876f
C6487 VDD.n4044 GND 0.28f
C6488 VDD.n4045 GND 0.166f
C6489 VDD.n4046 GND 0.196f
C6490 VDD.n4047 GND 0.0783f
C6491 VDD.n4048 GND 6.12f
C6492 VDD.n4049 GND 0.275f
C6493 VDD.n4050 GND 0.0237f
C6494 VDD.n4051 GND 0.0462f
C6495 VDD.t30 GND 0.0597f
C6496 VDD.n4063 GND 0.0351f
C6497 VDD.n4071 GND 0.0437f
C6498 VDD.n4072 GND 0.0152f
C6499 VDD.n4073 GND 0.0128f
C6500 VDD.n4080 GND 0.0504f
C6501 VDD.n4096 GND 0.0735f
C6502 VDD.t5 GND 0.0597f
C6503 VDD.n4097 GND 0.0351f
C6504 VDD.n4106 GND 0.0491f
C6505 VDD.n4108 GND 0.0135f
C6506 VDD.n4122 GND 0.0484f
C6507 VDD.n4123 GND 0.0582f
C6508 VDD.n4129 GND 0.0584f
C6509 VDD.n4133 GND 0.0134f
C6510 VDD.n4134 GND 0.047f
C6511 VDD.n4138 GND 0.0289f
C6512 VDD.n4139 GND 0.0135f
C6513 VDD.t409 GND 0.169f
C6514 VDD.n4149 GND 0.0735f
C6515 VDD.n4155 GND 0.0135f
C6516 VDD.n4156 GND 0.0287f
C6517 VDD.n4158 GND 0.0248f
C6518 VDD.n4159 GND 0.13f
C6519 VDD.n4160 GND 0.427f
C6520 VDD.n4186 GND 0.0444f
C6521 VDD.t7 GND 0.0187f
C6522 VDD.n4187 GND 0.0194f
C6523 VDD.n4188 GND 0.0239f
C6524 VDD.t27 GND 0.0185f
C6525 VDD.n4189 GND 0.16f
C6526 VDD.n4190 GND 0.967f
C6527 VDD.n4191 GND 0.103f
C6528 VDD.n4192 GND 1.15f
C6529 VDD.n4193 GND 0.921f
C6530 VDD.t1462 GND 0.0383f
C6531 VDD.t15 GND 0.0134f
C6532 VDD.n4194 GND 0.0699f
C6533 VDD.n4201 GND 0.058f
C6534 VDD.n4202 GND 0.0223f
C6535 VDD.n4206 GND 0.0683f
C6536 VDD.n4208 GND 0.078f
C6537 VDD.n4210 GND 0.0106f
C6538 VDD.t984 GND 0.0288f
C6539 VDD.t1363 GND 0.0109f
C6540 VDD.n4221 GND 0.0397f
C6541 VDD.n4224 GND 0.0201f
C6542 VDD.n4225 GND 0.0133f
C6543 VDD.n4226 GND 0.114f
C6544 VDD.n4227 GND 0.0382f
C6545 VDD.n4232 GND 0.0681f
C6546 VDD.n4234 GND 0.0899f
C6547 VDD.n4242 GND 0.0866f
C6548 VDD.n4243 GND 0.0386f
C6549 VDD.n4248 GND 0.0419f
C6550 VDD.t13 GND 0.0681f
C6551 VDD.n4257 GND 0.295f
C6552 VDD.n4258 GND 0.165f
C6553 VDD.n4259 GND 0.0664f
C6554 VDD.n4260 GND 0.0216f
C6555 VDD.t525 GND 0.0856f
C6556 VDD.n4271 GND 0.0455f
C6557 VDD.n4272 GND 0.112f
C6558 VDD.n4274 GND 0.0121f
C6559 VDD.n4277 GND 0.0858f
C6560 VDD.n4278 GND 0.0899f
C6561 VDD.n4286 GND 0.0427f
C6562 VDD.n4290 GND 0.0386f
C6563 VDD.t1021 GND 0.0681f
C6564 VDD.n4299 GND 0.0681f
C6565 VDD.n4301 GND 0.0876f
C6566 VDD.n4302 GND 0.28f
C6567 VDD.n4303 GND 0.166f
C6568 VDD.n4304 GND 0.196f
C6569 VDD.n4305 GND 0.0783f
C6570 VDD.n4306 GND 6.12f
C6571 VDD.n4307 GND 0.275f
C6572 VDD.n4308 GND 0.0237f
C6573 VDD.n4309 GND 0.0462f
C6574 VDD.t1436 GND 0.0597f
C6575 VDD.n4321 GND 0.0351f
C6576 VDD.n4329 GND 0.0437f
C6577 VDD.n4330 GND 0.0152f
C6578 VDD.n4331 GND 0.0128f
C6579 VDD.n4338 GND 0.0504f
C6580 VDD.n4354 GND 0.0735f
C6581 VDD.t1052 GND 0.0597f
C6582 VDD.n4355 GND 0.0351f
C6583 VDD.n4364 GND 0.0491f
C6584 VDD.n4366 GND 0.0135f
C6585 VDD.n4380 GND 0.0484f
C6586 VDD.n4381 GND 0.0582f
C6587 VDD.n4387 GND 0.0584f
C6588 VDD.n4391 GND 0.0134f
C6589 VDD.n4392 GND 0.047f
C6590 VDD.n4396 GND 0.0289f
C6591 VDD.n4397 GND 0.0135f
C6592 VDD.t1108 GND 0.169f
C6593 VDD.n4407 GND 0.0735f
C6594 VDD.n4413 GND 0.0135f
C6595 VDD.n4414 GND 0.0287f
C6596 VDD.n4416 GND 0.0248f
C6597 VDD.n4417 GND 0.13f
C6598 VDD.n4418 GND 0.427f
C6599 VDD.n4444 GND 0.0444f
C6600 VDD.t1050 GND 0.0187f
C6601 VDD.n4445 GND 0.0194f
C6602 VDD.n4446 GND 0.0239f
C6603 VDD.t1433 GND 0.0185f
C6604 VDD.n4447 GND 0.16f
C6605 VDD.n4448 GND 0.967f
C6606 VDD.n4449 GND 0.103f
C6607 VDD.n4450 GND 1.15f
C6608 VDD.n4451 GND 0.921f
C6609 VDD.t1105 GND 0.0383f
C6610 VDD.t1067 GND 0.0134f
C6611 VDD.n4452 GND 0.0699f
C6612 VDD.n4459 GND 0.058f
C6613 VDD.n4460 GND 0.0223f
C6614 VDD.n4464 GND 0.0683f
C6615 VDD.n4466 GND 0.078f
C6616 VDD.n4468 GND 0.0106f
C6617 VDD.t458 GND 0.0288f
C6618 VDD.t608 GND 0.0109f
C6619 VDD.n4479 GND 0.0397f
C6620 VDD.n4482 GND 0.0201f
C6621 VDD.n4483 GND 0.0133f
C6622 VDD.n4484 GND 0.114f
C6623 VDD.n4485 GND 0.0382f
C6624 VDD.n4490 GND 0.0681f
C6625 VDD.n4492 GND 0.0899f
C6626 VDD.n4500 GND 0.0866f
C6627 VDD.n4501 GND 0.0386f
C6628 VDD.n4506 GND 0.0419f
C6629 VDD.t415 GND 0.0681f
C6630 VDD.n4515 GND 0.295f
C6631 VDD.n4516 GND 0.165f
C6632 VDD.n4517 GND 0.0664f
C6633 VDD.n4518 GND 0.0216f
C6634 VDD.t264 GND 0.0856f
C6635 VDD.n4529 GND 0.0455f
C6636 VDD.n4530 GND 0.112f
C6637 VDD.n4532 GND 0.0121f
C6638 VDD.n4535 GND 0.0858f
C6639 VDD.n4536 GND 0.0899f
C6640 VDD.n4544 GND 0.0427f
C6641 VDD.n4548 GND 0.0386f
C6642 VDD.t531 GND 0.0681f
C6643 VDD.n4557 GND 0.0681f
C6644 VDD.n4559 GND 0.0876f
C6645 VDD.n4560 GND 0.28f
C6646 VDD.n4561 GND 0.166f
C6647 VDD.n4562 GND 0.196f
C6648 VDD.n4563 GND 0.0783f
C6649 VDD.n4564 GND 6.12f
C6650 VDD.n4565 GND 0.275f
C6651 VDD.n4566 GND 0.0237f
C6652 VDD.n4567 GND 0.0462f
C6653 VDD.t370 GND 0.0597f
C6654 VDD.n4579 GND 0.0351f
C6655 VDD.n4587 GND 0.0437f
C6656 VDD.n4588 GND 0.0152f
C6657 VDD.n4589 GND 0.0128f
C6658 VDD.n4596 GND 0.0504f
C6659 VDD.n4612 GND 0.0735f
C6660 VDD.t21 GND 0.0597f
C6661 VDD.n4613 GND 0.0351f
C6662 VDD.n4622 GND 0.0491f
C6663 VDD.n4624 GND 0.0135f
C6664 VDD.n4638 GND 0.0484f
C6665 VDD.n4639 GND 0.0582f
C6666 VDD.n4645 GND 0.0584f
C6667 VDD.n4649 GND 0.0134f
C6668 VDD.n4650 GND 0.047f
C6669 VDD.n4654 GND 0.0289f
C6670 VDD.n4655 GND 0.0135f
C6671 VDD.t332 GND 0.169f
C6672 VDD.n4665 GND 0.0735f
C6673 VDD.n4671 GND 0.0135f
C6674 VDD.n4672 GND 0.0287f
C6675 VDD.n4674 GND 0.0248f
C6676 VDD.n4675 GND 0.13f
C6677 VDD.n4676 GND 0.427f
C6678 VDD.n4702 GND 0.0444f
C6679 VDD.t19 GND 0.0187f
C6680 VDD.n4703 GND 0.0194f
C6681 VDD.n4704 GND 0.0239f
C6682 VDD.t372 GND 0.0185f
C6683 VDD.n4705 GND 0.16f
C6684 VDD.n4706 GND 0.967f
C6685 VDD.n4707 GND 0.103f
C6686 VDD.n4708 GND 1.15f
C6687 VDD.n4709 GND 0.921f
C6688 VDD.t1500 GND 0.0383f
C6689 VDD.t1309 GND 0.0134f
C6690 VDD.n4710 GND 0.0699f
C6691 VDD.n4717 GND 0.058f
C6692 VDD.n4718 GND 0.0223f
C6693 VDD.n4722 GND 0.0683f
C6694 VDD.n4724 GND 0.078f
C6695 VDD.n4726 GND 0.0106f
C6696 VDD.t1474 GND 0.0288f
C6697 VDD.t399 GND 0.0109f
C6698 VDD.n4737 GND 0.0397f
C6699 VDD.n4740 GND 0.0201f
C6700 VDD.n4741 GND 0.0133f
C6701 VDD.n4742 GND 0.114f
C6702 VDD.n4743 GND 0.0382f
C6703 VDD.n4748 GND 0.0681f
C6704 VDD.n4750 GND 0.0899f
C6705 VDD.n4758 GND 0.0866f
C6706 VDD.n4759 GND 0.0386f
C6707 VDD.n4764 GND 0.0419f
C6708 VDD.t527 GND 0.0681f
C6709 VDD.n4773 GND 0.295f
C6710 VDD.n4774 GND 0.165f
C6711 VDD.n4775 GND 0.0664f
C6712 VDD.n4776 GND 0.0216f
C6713 VDD.t590 GND 0.0856f
C6714 VDD.n4787 GND 0.0455f
C6715 VDD.n4788 GND 0.112f
C6716 VDD.n4790 GND 0.0121f
C6717 VDD.n4793 GND 0.0858f
C6718 VDD.n4794 GND 0.0899f
C6719 VDD.n4802 GND 0.0427f
C6720 VDD.n4806 GND 0.0386f
C6721 VDD.t401 GND 0.0681f
C6722 VDD.n4815 GND 0.0681f
C6723 VDD.n4817 GND 0.0876f
C6724 VDD.n4818 GND 0.28f
C6725 VDD.n4819 GND 0.166f
C6726 VDD.n4820 GND 0.196f
C6727 VDD.n4821 GND 0.0783f
C6728 VDD.n4822 GND 6.12f
C6729 VDD.n4823 GND 0.275f
C6730 VDD.n4824 GND 0.0237f
C6731 VDD.n4825 GND 0.0462f
C6732 VDD.t422 GND 0.0597f
C6733 VDD.n4837 GND 0.0351f
C6734 VDD.n4845 GND 0.0437f
C6735 VDD.n4846 GND 0.0152f
C6736 VDD.n4847 GND 0.0128f
C6737 VDD.n4854 GND 0.0504f
C6738 VDD.n4870 GND 0.0735f
C6739 VDD.t563 GND 0.0597f
C6740 VDD.n4871 GND 0.0351f
C6741 VDD.n4880 GND 0.0491f
C6742 VDD.n4882 GND 0.0135f
C6743 VDD.n4896 GND 0.0484f
C6744 VDD.n4897 GND 0.0582f
C6745 VDD.n4903 GND 0.0584f
C6746 VDD.n4907 GND 0.0134f
C6747 VDD.n4908 GND 0.047f
C6748 VDD.n4912 GND 0.0289f
C6749 VDD.n4913 GND 0.0135f
C6750 VDD.t279 GND 0.169f
C6751 VDD.n4923 GND 0.0735f
C6752 VDD.n4929 GND 0.0135f
C6753 VDD.n4930 GND 0.0287f
C6754 VDD.n4932 GND 0.0248f
C6755 VDD.n4933 GND 0.13f
C6756 VDD.n4934 GND 0.427f
C6757 VDD.n4960 GND 0.0444f
C6758 VDD.t560 GND 0.0187f
C6759 VDD.n4961 GND 0.0194f
C6760 VDD.n4962 GND 0.0239f
C6761 VDD.t420 GND 0.0185f
C6762 VDD.n4963 GND 0.16f
C6763 VDD.n4964 GND 0.967f
C6764 VDD.n4965 GND 0.103f
C6765 VDD.n4966 GND 1.15f
C6766 VDD.n4967 GND 0.921f
C6767 VDD.t1288 GND 0.0383f
C6768 VDD.t817 GND 0.0134f
C6769 VDD.n4968 GND 0.0699f
C6770 VDD.n4975 GND 0.058f
C6771 VDD.n4976 GND 0.0223f
C6772 VDD.n4980 GND 0.0683f
C6773 VDD.n4982 GND 0.078f
C6774 VDD.n4984 GND 0.0106f
C6775 VDD.t1042 GND 0.0288f
C6776 VDD.t1099 GND 0.0109f
C6777 VDD.n4995 GND 0.0397f
C6778 VDD.n4998 GND 0.0201f
C6779 VDD.n4999 GND 0.0133f
C6780 VDD.n5000 GND 0.114f
C6781 VDD.n5001 GND 0.0382f
C6782 VDD.n5006 GND 0.0681f
C6783 VDD.n5008 GND 0.0899f
C6784 VDD.n5016 GND 0.0866f
C6785 VDD.n5017 GND 0.0386f
C6786 VDD.n5022 GND 0.0419f
C6787 VDD.t815 GND 0.0681f
C6788 VDD.n5031 GND 0.295f
C6789 VDD.n5032 GND 0.165f
C6790 VDD.n5033 GND 0.0664f
C6791 VDD.n5034 GND 0.0216f
C6792 VDD.t1024 GND 0.0856f
C6793 VDD.n5045 GND 0.0455f
C6794 VDD.n5046 GND 0.112f
C6795 VDD.n5048 GND 0.0121f
C6796 VDD.n5051 GND 0.0858f
C6797 VDD.n5052 GND 0.0899f
C6798 VDD.n5060 GND 0.0427f
C6799 VDD.n5064 GND 0.0386f
C6800 VDD.t416 GND 0.0681f
C6801 VDD.n5073 GND 0.0681f
C6802 VDD.n5075 GND 0.0876f
C6803 VDD.n5076 GND 0.28f
C6804 VDD.n5077 GND 0.166f
C6805 VDD.n5078 GND 0.196f
C6806 VDD.n5079 GND 0.0783f
C6807 VDD.n5080 GND 6.12f
C6808 VDD.n5081 GND 0.275f
C6809 VDD.n5082 GND 0.0237f
C6810 VDD.n5083 GND 0.0462f
C6811 VDD.t0 GND 0.0597f
C6812 VDD.n5095 GND 0.0351f
C6813 VDD.n5103 GND 0.0437f
C6814 VDD.n5104 GND 0.0152f
C6815 VDD.n5105 GND 0.0128f
C6816 VDD.n5112 GND 0.0504f
C6817 VDD.n5128 GND 0.0735f
C6818 VDD.t1008 GND 0.0597f
C6819 VDD.n5129 GND 0.0351f
C6820 VDD.n5138 GND 0.0491f
C6821 VDD.n5140 GND 0.0135f
C6822 VDD.n5154 GND 0.0484f
C6823 VDD.n5155 GND 0.0582f
C6824 VDD.n5161 GND 0.0584f
C6825 VDD.n5165 GND 0.0134f
C6826 VDD.n5166 GND 0.047f
C6827 VDD.n5170 GND 0.0289f
C6828 VDD.n5171 GND 0.0135f
C6829 VDD.t1060 GND 0.169f
C6830 VDD.n5181 GND 0.0735f
C6831 VDD.n5187 GND 0.0135f
C6832 VDD.n5188 GND 0.0287f
C6833 VDD.n5190 GND 0.0248f
C6834 VDD.n5191 GND 0.13f
C6835 VDD.n5192 GND 0.427f
C6836 VDD.n5218 GND 0.0444f
C6837 VDD.t1006 GND 0.0187f
C6838 VDD.n5219 GND 0.0194f
C6839 VDD.n5220 GND 0.0239f
C6840 VDD.t2 GND 0.0185f
C6841 VDD.n5221 GND 0.16f
C6842 VDD.n5222 GND 0.967f
C6843 VDD.n5223 GND 0.103f
C6844 VDD.n5224 GND 1.15f
C6845 VDD.n5225 GND 0.921f
C6846 VDD.t481 GND 0.0383f
C6847 VDD.t1058 GND 0.0134f
C6848 VDD.n5226 GND 0.0699f
C6849 VDD.n5233 GND 0.058f
C6850 VDD.n5234 GND 0.0223f
C6851 VDD.n5238 GND 0.0683f
C6852 VDD.n5240 GND 0.078f
C6853 VDD.n5242 GND 0.0106f
C6854 VDD.t633 GND 0.0288f
C6855 VDD.t405 GND 0.0109f
C6856 VDD.n5253 GND 0.0397f
C6857 VDD.n5256 GND 0.0201f
C6858 VDD.n5257 GND 0.0133f
C6859 VDD.n5258 GND 0.114f
C6860 VDD.n5259 GND 0.0382f
C6861 VDD.n5264 GND 0.0681f
C6862 VDD.n5266 GND 0.0899f
C6863 VDD.n5274 GND 0.0866f
C6864 VDD.n5275 GND 0.0386f
C6865 VDD.n5280 GND 0.0419f
C6866 VDD.t265 GND 0.0681f
C6867 VDD.n5289 GND 0.295f
C6868 VDD.n5290 GND 0.165f
C6869 VDD.n5291 GND 0.0664f
C6870 VDD.n5292 GND 0.0216f
C6871 VDD.t275 GND 0.0856f
C6872 VDD.n5303 GND 0.0455f
C6873 VDD.n5304 GND 0.112f
C6874 VDD.n5306 GND 0.0121f
C6875 VDD.n5309 GND 0.0858f
C6876 VDD.n5310 GND 0.0899f
C6877 VDD.n5318 GND 0.0427f
C6878 VDD.n5322 GND 0.0386f
C6879 VDD.t407 GND 0.0681f
C6880 VDD.n5331 GND 0.0681f
C6881 VDD.n5333 GND 0.0876f
C6882 VDD.n5334 GND 0.28f
C6883 VDD.n5335 GND 0.166f
C6884 VDD.n5336 GND 0.196f
C6885 VDD.n5337 GND 0.0783f
C6886 VDD.n5338 GND 9.87f
C6887 VDD.n5339 GND 22.6f
C6888 VDD.n5340 GND 14f
C6889 VDD.n5341 GND 14f
C6890 VDD.n5342 GND 14f
C6891 VDD.n5343 GND 14f
C6892 VDD.n5344 GND 14.5f
C6893 VDD.n5345 GND 0.0237f
C6894 VDD.n5346 GND 0.0462f
C6895 VDD.t1258 GND 0.0597f
C6896 VDD.n5358 GND 0.0351f
C6897 VDD.n5366 GND 0.0437f
C6898 VDD.n5367 GND 0.0152f
C6899 VDD.n5368 GND 0.0128f
C6900 VDD.n5375 GND 0.0504f
C6901 VDD.n5391 GND 0.0735f
C6902 VDD.t995 GND 0.0597f
C6903 VDD.n5392 GND 0.0351f
C6904 VDD.n5401 GND 0.0491f
C6905 VDD.n5403 GND 0.0135f
C6906 VDD.n5417 GND 0.0484f
C6907 VDD.n5418 GND 0.0582f
C6908 VDD.n5424 GND 0.0584f
C6909 VDD.n5428 GND 0.0134f
C6910 VDD.n5429 GND 0.047f
C6911 VDD.n5433 GND 0.0289f
C6912 VDD.n5434 GND 0.0135f
C6913 VDD.t270 GND 0.169f
C6914 VDD.n5444 GND 0.0735f
C6915 VDD.n5450 GND 0.0135f
C6916 VDD.n5451 GND 0.0287f
C6917 VDD.n5453 GND 0.0248f
C6918 VDD.n5454 GND 0.927f
C6919 VDD.n5455 GND 1.67f
C6920 VDD.n5481 GND 0.0444f
C6921 VDD.t997 GND 0.0187f
C6922 VDD.n5482 GND 0.0194f
C6923 VDD.n5483 GND 0.0239f
C6924 VDD.t1256 GND 0.0185f
C6925 VDD.n5484 GND 0.17f
C6926 VDD.n5485 GND 1.7f
C6927 VDD.t453 GND 0.0383f
C6928 VDD.t643 GND 0.0134f
C6929 VDD.n5486 GND 0.0699f
C6930 VDD.n5493 GND 0.058f
C6931 VDD.n5494 GND 0.0223f
C6932 VDD.n5498 GND 0.0683f
C6933 VDD.n5500 GND 0.078f
C6934 VDD.n5502 GND 0.0106f
C6935 VDD.t1305 GND 0.0288f
C6936 VDD.t391 GND 0.0109f
C6937 VDD.n5513 GND 0.0397f
C6938 VDD.n5516 GND 0.0201f
C6939 VDD.n5517 GND 0.0133f
C6940 VDD.n5518 GND 0.114f
C6941 VDD.n5519 GND 0.0382f
C6942 VDD.n5524 GND 0.0681f
C6943 VDD.n5526 GND 0.0899f
C6944 VDD.n5534 GND 0.0866f
C6945 VDD.n5535 GND 0.0386f
C6946 VDD.n5540 GND 0.0419f
C6947 VDD.t507 GND 0.0681f
C6948 VDD.n5549 GND 0.295f
C6949 VDD.n5550 GND 0.165f
C6950 VDD.n5551 GND 0.0664f
C6951 VDD.n5552 GND 0.0216f
C6952 VDD.t512 GND 0.0856f
C6953 VDD.n5563 GND 0.0455f
C6954 VDD.n5564 GND 0.112f
C6955 VDD.n5566 GND 0.0121f
C6956 VDD.n5569 GND 0.0858f
C6957 VDD.n5570 GND 0.0899f
C6958 VDD.n5578 GND 0.0427f
C6959 VDD.n5582 GND 0.0386f
C6960 VDD.t393 GND 0.0681f
C6961 VDD.n5591 GND 0.0681f
C6962 VDD.n5593 GND 0.0876f
C6963 VDD.n5594 GND 0.28f
C6964 VDD.n5595 GND 0.166f
C6965 VDD.n5596 GND 1.98f
C6966 VDD.n5597 GND 6.4f
C6967 VDD.n5598 GND 11.2f
C6968 VDD.n5599 GND 0.0237f
C6969 VDD.n5600 GND 0.0462f
C6970 VDD.t476 GND 0.0597f
C6971 VDD.n5612 GND 0.0351f
C6972 VDD.n5620 GND 0.0437f
C6973 VDD.n5621 GND 0.0152f
C6974 VDD.n5622 GND 0.0128f
C6975 VDD.n5629 GND 0.0504f
C6976 VDD.n5645 GND 0.0735f
C6977 VDD.t1468 GND 0.0597f
C6978 VDD.n5646 GND 0.0351f
C6979 VDD.n5655 GND 0.0491f
C6980 VDD.n5657 GND 0.0135f
C6981 VDD.n5671 GND 0.0484f
C6982 VDD.n5672 GND 0.0582f
C6983 VDD.n5678 GND 0.0584f
C6984 VDD.n5682 GND 0.0134f
C6985 VDD.n5683 GND 0.047f
C6986 VDD.n5687 GND 0.0289f
C6987 VDD.n5688 GND 0.0135f
C6988 VDD.t1307 GND 0.169f
C6989 VDD.n5698 GND 0.0735f
C6990 VDD.n5704 GND 0.0135f
C6991 VDD.n5705 GND 0.0287f
C6992 VDD.n5707 GND 0.0248f
C6993 VDD.n5708 GND 0.927f
C6994 VDD.n5709 GND 1.67f
C6995 VDD.n5735 GND 0.0444f
C6996 VDD.t1466 GND 0.0187f
C6997 VDD.n5736 GND 0.0194f
C6998 VDD.n5737 GND 0.0239f
C6999 VDD.t473 GND 0.0185f
C7000 VDD.n5738 GND 0.17f
C7001 VDD.n5739 GND 1.7f
C7002 VDD.t519 GND 0.0383f
C7003 VDD.t601 GND 0.0134f
C7004 VDD.n5740 GND 0.0699f
C7005 VDD.n5747 GND 0.058f
C7006 VDD.n5748 GND 0.0223f
C7007 VDD.n5752 GND 0.0683f
C7008 VDD.n5754 GND 0.078f
C7009 VDD.n5756 GND 0.0106f
C7010 VDD.t67 GND 0.0288f
C7011 VDD.t1353 GND 0.0109f
C7012 VDD.n5767 GND 0.0397f
C7013 VDD.n5770 GND 0.0201f
C7014 VDD.n5771 GND 0.0133f
C7015 VDD.n5772 GND 0.114f
C7016 VDD.n5773 GND 0.0382f
C7017 VDD.n5778 GND 0.0681f
C7018 VDD.n5780 GND 0.0899f
C7019 VDD.n5788 GND 0.0866f
C7020 VDD.n5789 GND 0.0386f
C7021 VDD.n5794 GND 0.0419f
C7022 VDD.t514 GND 0.0681f
C7023 VDD.n5803 GND 0.295f
C7024 VDD.n5804 GND 0.165f
C7025 VDD.n5805 GND 0.0664f
C7026 VDD.n5806 GND 0.0216f
C7027 VDD.t276 GND 0.0856f
C7028 VDD.n5817 GND 0.0455f
C7029 VDD.n5818 GND 0.112f
C7030 VDD.n5820 GND 0.0121f
C7031 VDD.n5823 GND 0.0858f
C7032 VDD.n5824 GND 0.0899f
C7033 VDD.n5832 GND 0.0427f
C7034 VDD.n5836 GND 0.0386f
C7035 VDD.t1075 GND 0.0681f
C7036 VDD.n5845 GND 0.0681f
C7037 VDD.n5847 GND 0.0876f
C7038 VDD.n5848 GND 0.28f
C7039 VDD.n5849 GND 0.166f
C7040 VDD.n5850 GND 1.98f
C7041 VDD.n5851 GND 6.4f
C7042 VDD.n5852 GND 11.2f
C7043 VDD.n5853 GND 14.5f
C7044 VDD.n5854 GND 14f
C7045 VDD.n5855 GND 14f
C7046 VDD.n5856 GND 14f
C7047 VDD.n5857 GND 14f
C7048 VDD.n5858 GND 10.2f
C7049 VDD.n5859 GND 7.31f
C7050 VDD.n5860 GND 20.4f
C7051 VDD.n5861 GND 34.2f
C7052 VDD.n5862 GND 10.2f
C7053 VDD.n5863 GND 14.2f
.ends

