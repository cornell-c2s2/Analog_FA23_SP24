magic
tech sky130A
magscale 1 2
timestamp 1717119771
<< error_p >>
rect -372 5072 -314 5078
rect -176 5072 -118 5078
rect 20 5072 78 5078
rect 216 5072 274 5078
rect 412 5072 470 5078
rect -372 5038 -360 5072
rect -176 5038 -164 5072
rect 20 5038 32 5072
rect 216 5038 228 5072
rect 412 5038 424 5072
rect -372 5032 -314 5038
rect -176 5032 -118 5038
rect 20 5032 78 5038
rect 216 5032 274 5038
rect 412 5032 470 5038
rect -470 -5038 -412 -5032
rect -274 -5038 -216 -5032
rect -78 -5038 -20 -5032
rect 118 -5038 176 -5032
rect 314 -5038 372 -5032
rect -470 -5072 -458 -5038
rect -274 -5072 -262 -5038
rect -78 -5072 -66 -5038
rect 118 -5072 130 -5038
rect 314 -5072 326 -5038
rect -470 -5078 -412 -5072
rect -274 -5078 -216 -5072
rect -78 -5078 -20 -5072
rect 118 -5078 176 -5072
rect 314 -5078 372 -5072
<< pwell >>
rect -657 -5210 657 5210
<< nmos >>
rect -461 -5000 -421 5000
rect -363 -5000 -323 5000
rect -265 -5000 -225 5000
rect -167 -5000 -127 5000
rect -69 -5000 -29 5000
rect 29 -5000 69 5000
rect 127 -5000 167 5000
rect 225 -5000 265 5000
rect 323 -5000 363 5000
rect 421 -5000 461 5000
<< ndiff >>
rect -519 4988 -461 5000
rect -519 -4988 -507 4988
rect -473 -4988 -461 4988
rect -519 -5000 -461 -4988
rect -421 4988 -363 5000
rect -421 -4988 -409 4988
rect -375 -4988 -363 4988
rect -421 -5000 -363 -4988
rect -323 4988 -265 5000
rect -323 -4988 -311 4988
rect -277 -4988 -265 4988
rect -323 -5000 -265 -4988
rect -225 4988 -167 5000
rect -225 -4988 -213 4988
rect -179 -4988 -167 4988
rect -225 -5000 -167 -4988
rect -127 4988 -69 5000
rect -127 -4988 -115 4988
rect -81 -4988 -69 4988
rect -127 -5000 -69 -4988
rect -29 4988 29 5000
rect -29 -4988 -17 4988
rect 17 -4988 29 4988
rect -29 -5000 29 -4988
rect 69 4988 127 5000
rect 69 -4988 81 4988
rect 115 -4988 127 4988
rect 69 -5000 127 -4988
rect 167 4988 225 5000
rect 167 -4988 179 4988
rect 213 -4988 225 4988
rect 167 -5000 225 -4988
rect 265 4988 323 5000
rect 265 -4988 277 4988
rect 311 -4988 323 4988
rect 265 -5000 323 -4988
rect 363 4988 421 5000
rect 363 -4988 375 4988
rect 409 -4988 421 4988
rect 363 -5000 421 -4988
rect 461 4988 519 5000
rect 461 -4988 473 4988
rect 507 -4988 519 4988
rect 461 -5000 519 -4988
<< ndiffc >>
rect -507 -4988 -473 4988
rect -409 -4988 -375 4988
rect -311 -4988 -277 4988
rect -213 -4988 -179 4988
rect -115 -4988 -81 4988
rect -17 -4988 17 4988
rect 81 -4988 115 4988
rect 179 -4988 213 4988
rect 277 -4988 311 4988
rect 375 -4988 409 4988
rect 473 -4988 507 4988
<< psubdiff >>
rect -621 5140 621 5174
rect -621 5078 -587 5140
rect 587 5078 621 5140
rect -621 -5140 -587 -5078
rect 587 -5140 621 -5078
rect -621 -5174 -525 -5140
rect 525 -5174 621 -5140
<< psubdiffcont >>
rect -621 -5078 -587 5078
rect 587 -5078 621 5078
rect -525 -5174 525 -5140
<< poly >>
rect -376 5072 -310 5088
rect -376 5038 -360 5072
rect -326 5038 -310 5072
rect -461 5000 -421 5026
rect -376 5022 -310 5038
rect -180 5072 -114 5088
rect -180 5038 -164 5072
rect -130 5038 -114 5072
rect -363 5000 -323 5022
rect -265 5000 -225 5026
rect -180 5022 -114 5038
rect 16 5072 82 5088
rect 16 5038 32 5072
rect 66 5038 82 5072
rect -167 5000 -127 5022
rect -69 5000 -29 5026
rect 16 5022 82 5038
rect 212 5072 278 5088
rect 212 5038 228 5072
rect 262 5038 278 5072
rect 29 5000 69 5022
rect 127 5000 167 5026
rect 212 5022 278 5038
rect 408 5072 474 5088
rect 408 5038 424 5072
rect 458 5038 474 5072
rect 225 5000 265 5022
rect 323 5000 363 5026
rect 408 5022 474 5038
rect 421 5000 461 5022
rect -461 -5022 -421 -5000
rect -474 -5038 -408 -5022
rect -363 -5026 -323 -5000
rect -265 -5022 -225 -5000
rect -474 -5072 -458 -5038
rect -424 -5072 -408 -5038
rect -474 -5088 -408 -5072
rect -278 -5038 -212 -5022
rect -167 -5026 -127 -5000
rect -69 -5022 -29 -5000
rect -278 -5072 -262 -5038
rect -228 -5072 -212 -5038
rect -278 -5088 -212 -5072
rect -82 -5038 -16 -5022
rect 29 -5026 69 -5000
rect 127 -5022 167 -5000
rect -82 -5072 -66 -5038
rect -32 -5072 -16 -5038
rect -82 -5088 -16 -5072
rect 114 -5038 180 -5022
rect 225 -5026 265 -5000
rect 323 -5022 363 -5000
rect 114 -5072 130 -5038
rect 164 -5072 180 -5038
rect 114 -5088 180 -5072
rect 310 -5038 376 -5022
rect 421 -5026 461 -5000
rect 310 -5072 326 -5038
rect 360 -5072 376 -5038
rect 310 -5088 376 -5072
<< polycont >>
rect -360 5038 -326 5072
rect -164 5038 -130 5072
rect 32 5038 66 5072
rect 228 5038 262 5072
rect 424 5038 458 5072
rect -458 -5072 -424 -5038
rect -262 -5072 -228 -5038
rect -66 -5072 -32 -5038
rect 130 -5072 164 -5038
rect 326 -5072 360 -5038
<< locali >>
rect -621 5140 621 5174
rect -621 5078 -587 5140
rect 587 5078 621 5140
rect -376 5038 -360 5072
rect -326 5038 -310 5072
rect -180 5038 -164 5072
rect -130 5038 -114 5072
rect 16 5038 32 5072
rect 66 5038 82 5072
rect 212 5038 228 5072
rect 262 5038 278 5072
rect 408 5038 424 5072
rect 458 5038 474 5072
rect -507 4988 -473 5004
rect -507 -5004 -473 -4988
rect -409 4988 -375 5004
rect -409 -5004 -375 -4988
rect -311 4988 -277 5004
rect -311 -5004 -277 -4988
rect -213 4988 -179 5004
rect -213 -5004 -179 -4988
rect -115 4988 -81 5004
rect -115 -5004 -81 -4988
rect -17 4988 17 5004
rect -17 -5004 17 -4988
rect 81 4988 115 5004
rect 81 -5004 115 -4988
rect 179 4988 213 5004
rect 179 -5004 213 -4988
rect 277 4988 311 5004
rect 277 -5004 311 -4988
rect 375 4988 409 5004
rect 375 -5004 409 -4988
rect 473 4988 507 5004
rect 473 -5004 507 -4988
rect -474 -5072 -458 -5038
rect -424 -5072 -408 -5038
rect -278 -5072 -262 -5038
rect -228 -5072 -212 -5038
rect -82 -5072 -66 -5038
rect -32 -5072 -16 -5038
rect 114 -5072 130 -5038
rect 164 -5072 180 -5038
rect 310 -5072 326 -5038
rect 360 -5072 376 -5038
rect -621 -5140 -587 -5078
rect 587 -5140 621 -5078
rect -621 -5174 -525 -5140
rect 525 -5174 621 -5140
<< viali >>
rect -360 5038 -326 5072
rect -164 5038 -130 5072
rect 32 5038 66 5072
rect 228 5038 262 5072
rect 424 5038 458 5072
rect -621 -2570 -587 2570
rect -507 -4988 -473 4988
rect -409 -4988 -375 4988
rect -311 -4988 -277 4988
rect -213 -4988 -179 4988
rect -115 -4988 -81 4988
rect -17 -4988 17 4988
rect 81 -4988 115 4988
rect 179 -4988 213 4988
rect 277 -4988 311 4988
rect 375 -4988 409 4988
rect 473 -4988 507 4988
rect 587 -2570 621 2570
rect -458 -5072 -424 -5038
rect -262 -5072 -228 -5038
rect -66 -5072 -32 -5038
rect 130 -5072 164 -5038
rect 326 -5072 360 -5038
rect -293 -5174 293 -5140
<< metal1 >>
rect -372 5072 -314 5078
rect -372 5038 -360 5072
rect -326 5038 -314 5072
rect -372 5032 -314 5038
rect -176 5072 -118 5078
rect -176 5038 -164 5072
rect -130 5038 -118 5072
rect -176 5032 -118 5038
rect 20 5072 78 5078
rect 20 5038 32 5072
rect 66 5038 78 5072
rect 20 5032 78 5038
rect 216 5072 274 5078
rect 216 5038 228 5072
rect 262 5038 274 5072
rect 216 5032 274 5038
rect 412 5072 470 5078
rect 412 5038 424 5072
rect 458 5038 470 5072
rect 412 5032 470 5038
rect -513 4988 -467 5000
rect -627 2570 -581 2582
rect -627 -2570 -621 2570
rect -587 -2570 -581 2570
rect -627 -2582 -581 -2570
rect -513 -4988 -507 4988
rect -473 -4988 -467 4988
rect -513 -5000 -467 -4988
rect -415 4988 -369 5000
rect -415 -4988 -409 4988
rect -375 -4988 -369 4988
rect -415 -5000 -369 -4988
rect -317 4988 -271 5000
rect -317 -4988 -311 4988
rect -277 -4988 -271 4988
rect -317 -5000 -271 -4988
rect -219 4988 -173 5000
rect -219 -4988 -213 4988
rect -179 -4988 -173 4988
rect -219 -5000 -173 -4988
rect -121 4988 -75 5000
rect -121 -4988 -115 4988
rect -81 -4988 -75 4988
rect -121 -5000 -75 -4988
rect -23 4988 23 5000
rect -23 -4988 -17 4988
rect 17 -4988 23 4988
rect -23 -5000 23 -4988
rect 75 4988 121 5000
rect 75 -4988 81 4988
rect 115 -4988 121 4988
rect 75 -5000 121 -4988
rect 173 4988 219 5000
rect 173 -4988 179 4988
rect 213 -4988 219 4988
rect 173 -5000 219 -4988
rect 271 4988 317 5000
rect 271 -4988 277 4988
rect 311 -4988 317 4988
rect 271 -5000 317 -4988
rect 369 4988 415 5000
rect 369 -4988 375 4988
rect 409 -4988 415 4988
rect 369 -5000 415 -4988
rect 467 4988 513 5000
rect 467 -4988 473 4988
rect 507 -4988 513 4988
rect 581 2570 627 2582
rect 581 -2570 587 2570
rect 621 -2570 627 2570
rect 581 -2582 627 -2570
rect 467 -5000 513 -4988
rect -470 -5038 -412 -5032
rect -470 -5072 -458 -5038
rect -424 -5072 -412 -5038
rect -470 -5078 -412 -5072
rect -274 -5038 -216 -5032
rect -274 -5072 -262 -5038
rect -228 -5072 -216 -5038
rect -274 -5078 -216 -5072
rect -78 -5038 -20 -5032
rect -78 -5072 -66 -5038
rect -32 -5072 -20 -5038
rect -78 -5078 -20 -5072
rect 118 -5038 176 -5032
rect 118 -5072 130 -5038
rect 164 -5072 176 -5038
rect 118 -5078 176 -5072
rect 314 -5038 372 -5032
rect 314 -5072 326 -5038
rect 360 -5072 372 -5038
rect 314 -5078 372 -5072
rect -305 -5140 305 -5134
rect -305 -5174 -293 -5140
rect 293 -5174 305 -5140
rect -305 -5180 305 -5174
<< properties >>
string FIXED_BBOX -604 -5157 604 5157
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 50 l 0.2 m 1 nf 10 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 0 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 50 viagr 50 viagl 50 viagt 0
<< end >>
