** sch_path: /foss/designs/Analog_FA23_SP24/SP24_caravel_user_project_analog/xschem/user_analog_project_wrapper.sch
.subckt user_analog_project_wrapper vdda1 vdda2 vssa1 vssa2 vccd1 vccd2 vssd1 vssd2 wb_clk_i wb_rst_i wbs_stb_i wbs_cyc_i wbs_we_i
+ wbs_sel_i[3] wbs_sel_i[2] wbs_sel_i[1] wbs_sel_i[0] wbs_dat_i[31] wbs_dat_i[30] wbs_dat_i[29] wbs_dat_i[28] wbs_dat_i[27] wbs_dat_i[26]
+ wbs_dat_i[25] wbs_dat_i[24] wbs_dat_i[23] wbs_dat_i[22] wbs_dat_i[21] wbs_dat_i[20] wbs_dat_i[19] wbs_dat_i[18] wbs_dat_i[17] wbs_dat_i[16]
+ wbs_dat_i[15] wbs_dat_i[14] wbs_dat_i[13] wbs_dat_i[12] wbs_dat_i[11] wbs_dat_i[10] wbs_dat_i[9] wbs_dat_i[8] wbs_dat_i[7] wbs_dat_i[6]
+ wbs_dat_i[5] wbs_dat_i[4] wbs_dat_i[3] wbs_dat_i[2] wbs_dat_i[1] wbs_dat_i[0] wbs_adr_i[31] wbs_adr_i[30] wbs_adr_i[29] wbs_adr_i[28]
+ wbs_adr_i[27] wbs_adr_i[26] wbs_adr_i[25] wbs_adr_i[24] wbs_adr_i[23] wbs_adr_i[22] wbs_adr_i[21] wbs_adr_i[20] wbs_adr_i[19] wbs_adr_i[18]
+ wbs_adr_i[17] wbs_adr_i[16] wbs_adr_i[15] wbs_adr_i[14] wbs_adr_i[13] wbs_adr_i[12] wbs_adr_i[11] wbs_adr_i[10] wbs_adr_i[9] wbs_adr_i[8]
+ wbs_adr_i[7] wbs_adr_i[6] wbs_adr_i[5] wbs_adr_i[4] wbs_adr_i[3] wbs_adr_i[2] wbs_adr_i[1] wbs_adr_i[0] wbs_ack_o wbs_dat_o[31] wbs_dat_o[30]
+ wbs_dat_o[29] wbs_dat_o[28] wbs_dat_o[27] wbs_dat_o[26] wbs_dat_o[25] wbs_dat_o[24] wbs_dat_o[23] wbs_dat_o[22] wbs_dat_o[21] wbs_dat_o[20]
+ wbs_dat_o[19] wbs_dat_o[18] wbs_dat_o[17] wbs_dat_o[16] wbs_dat_o[15] wbs_dat_o[14] wbs_dat_o[13] wbs_dat_o[12] wbs_dat_o[11] wbs_dat_o[10]
+ wbs_dat_o[9] wbs_dat_o[8] wbs_dat_o[7] wbs_dat_o[6] wbs_dat_o[5] wbs_dat_o[4] wbs_dat_o[3] wbs_dat_o[2] wbs_dat_o[1] wbs_dat_o[0]
+ la_data_in[127] la_data_in[126] la_data_in[125] la_data_in[124] la_data_in[123] la_data_in[122] la_data_in[121] la_data_in[120] la_data_in[119]
+ la_data_in[118] la_data_in[117] la_data_in[116] la_data_in[115] la_data_in[114] la_data_in[113] la_data_in[112] la_data_in[111] la_data_in[110]
+ la_data_in[109] la_data_in[108] la_data_in[107] la_data_in[106] la_data_in[105] la_data_in[104] la_data_in[103] la_data_in[102] la_data_in[101]
+ la_data_in[100] la_data_in[99] la_data_in[98] la_data_in[97] la_data_in[96] la_data_in[95] la_data_in[94] la_data_in[93] la_data_in[92]
+ la_data_in[91] la_data_in[90] la_data_in[89] la_data_in[88] la_data_in[87] la_data_in[86] la_data_in[85] la_data_in[84] la_data_in[83]
+ la_data_in[82] la_data_in[81] la_data_in[80] la_data_in[79] la_data_in[78] la_data_in[77] la_data_in[76] la_data_in[75] la_data_in[74]
+ la_data_in[73] la_data_in[72] la_data_in[71] la_data_in[70] la_data_in[69] la_data_in[68] la_data_in[67] la_data_in[66] la_data_in[65]
+ la_data_in[64] la_data_in[63] la_data_in[62] la_data_in[61] la_data_in[60] la_data_in[59] la_data_in[58] la_data_in[57] la_data_in[56]
+ la_data_in[55] la_data_in[54] la_data_in[53] la_data_in[52] la_data_in[51] la_data_in[50] la_data_in[49] la_data_in[48] la_data_in[47]
+ la_data_in[46] la_data_in[45] la_data_in[44] la_data_in[43] la_data_in[42] la_data_in[41] la_data_in[40] la_data_in[39] la_data_in[38]
+ la_data_in[37] la_data_in[36] la_data_in[35] la_data_in[34] la_data_in[33] la_data_in[32] la_data_in[31] la_data_in[30] la_data_in[29]
+ la_data_in[28] la_data_in[27] la_data_in[26] la_data_in[25] la_data_in[24] la_data_in[23] la_data_in[22] la_data_in[21] la_data_in[20]
+ la_data_in[19] la_data_in[18] la_data_in[17] la_data_in[16] la_data_in[15] la_data_in[14] la_data_in[13] la_data_in[12] la_data_in[11]
+ la_data_in[10] la_data_in[9] la_data_in[8] la_data_in[7] la_data_in[6] la_data_in[5] la_data_in[4] la_data_in[3] la_data_in[2] la_data_in[1]
+ la_data_in[0] la_data_out[127] la_data_out[126] la_data_out[125] la_data_out[124] la_data_out[123] la_data_out[122] la_data_out[121]
+ la_data_out[120] la_data_out[119] la_data_out[118] la_data_out[117] la_data_out[116] la_data_out[115] la_data_out[114] la_data_out[113]
+ la_data_out[112] la_data_out[111] la_data_out[110] la_data_out[109] la_data_out[108] la_data_out[107] la_data_out[106] la_data_out[105]
+ la_data_out[104] la_data_out[103] la_data_out[102] la_data_out[101] la_data_out[100] la_data_out[99] la_data_out[98] la_data_out[97]
+ la_data_out[96] la_data_out[95] la_data_out[94] la_data_out[93] la_data_out[92] la_data_out[91] la_data_out[90] la_data_out[89] la_data_out[88]
+ la_data_out[87] la_data_out[86] la_data_out[85] la_data_out[84] la_data_out[83] la_data_out[82] la_data_out[81] la_data_out[80] la_data_out[79]
+ la_data_out[78] la_data_out[77] la_data_out[76] la_data_out[75] la_data_out[74] la_data_out[73] la_data_out[72] la_data_out[71] la_data_out[70]
+ la_data_out[69] la_data_out[68] la_data_out[67] la_data_out[66] la_data_out[65] la_data_out[64] la_data_out[63] la_data_out[62] la_data_out[61]
+ la_data_out[60] la_data_out[59] la_data_out[58] la_data_out[57] la_data_out[56] la_data_out[55] la_data_out[54] la_data_out[53] la_data_out[52]
+ la_data_out[51] la_data_out[50] la_data_out[49] la_data_out[48] la_data_out[47] la_data_out[46] la_data_out[45] la_data_out[44] la_data_out[43]
+ la_data_out[42] la_data_out[41] la_data_out[40] la_data_out[39] la_data_out[38] la_data_out[37] la_data_out[36] la_data_out[35] la_data_out[34]
+ la_data_out[33] la_data_out[32] la_data_out[31] la_data_out[30] la_data_out[29] la_data_out[28] la_data_out[27] la_data_out[26] la_data_out[25]
+ la_data_out[24] la_data_out[23] la_data_out[22] la_data_out[21] la_data_out[20] la_data_out[19] la_data_out[18] la_data_out[17] la_data_out[16]
+ la_data_out[15] la_data_out[14] la_data_out[13] la_data_out[12] la_data_out[11] la_data_out[10] la_data_out[9] la_data_out[8] la_data_out[7]
+ la_data_out[6] la_data_out[5] la_data_out[4] la_data_out[3] la_data_out[2] la_data_out[1] la_data_out[0] la_oenb[127] la_oenb[126] la_oenb[125]
+ la_oenb[124] la_oenb[123] la_oenb[122] la_oenb[121] la_oenb[120] la_oenb[119] la_oenb[118] la_oenb[117] la_oenb[116] la_oenb[115] la_oenb[114]
+ la_oenb[113] la_oenb[112] la_oenb[111] la_oenb[110] la_oenb[109] la_oenb[108] la_oenb[107] la_oenb[106] la_oenb[105] la_oenb[104] la_oenb[103]
+ la_oenb[102] la_oenb[101] la_oenb[100] la_oenb[99] la_oenb[98] la_oenb[97] la_oenb[96] la_oenb[95] la_oenb[94] la_oenb[93] la_oenb[92]
+ la_oenb[91] la_oenb[90] la_oenb[89] la_oenb[88] la_oenb[87] la_oenb[86] la_oenb[85] la_oenb[84] la_oenb[83] la_oenb[82] la_oenb[81]
+ la_oenb[80] la_oenb[79] la_oenb[78] la_oenb[77] la_oenb[76] la_oenb[75] la_oenb[74] la_oenb[73] la_oenb[72] la_oenb[71] la_oenb[70]
+ la_oenb[69] la_oenb[68] la_oenb[67] la_oenb[66] la_oenb[65] la_oenb[64] la_oenb[63] la_oenb[62] la_oenb[61] la_oenb[60] la_oenb[59]
+ la_oenb[58] la_oenb[57] la_oenb[56] la_oenb[55] la_oenb[54] la_oenb[53] la_oenb[52] la_oenb[51] la_oenb[50] la_oenb[49] la_oenb[48]
+ la_oenb[47] la_oenb[46] la_oenb[45] la_oenb[44] la_oenb[43] la_oenb[42] la_oenb[41] la_oenb[40] la_oenb[39] la_oenb[38] la_oenb[37]
+ la_oenb[36] la_oenb[35] la_oenb[34] la_oenb[33] la_oenb[32] la_oenb[31] la_oenb[30] la_oenb[29] la_oenb[28] la_oenb[27] la_oenb[26]
+ la_oenb[25] la_oenb[24] la_oenb[23] la_oenb[22] la_oenb[21] la_oenb[20] la_oenb[19] la_oenb[18] la_oenb[17] la_oenb[16] la_oenb[15]
+ la_oenb[14] la_oenb[13] la_oenb[12] la_oenb[11] la_oenb[10] la_oenb[9] la_oenb[8] la_oenb[7] la_oenb[6] la_oenb[5] la_oenb[4] la_oenb[3]
+ la_oenb[2] la_oenb[1] la_oenb[0] io_in[26] io_in[25] io_in[24] io_in[23] io_in[22] io_in[21] io_in[20] io_in[19] io_in[18] io_in[17]
+ io_in[16] io_in[15] io_in[14] io_in[13] io_in[12] io_in[11] io_in[10] io_in[9] io_in[8] io_in[7] io_in[6] io_in[5] io_in[4] io_in[3]
+ io_in[2] io_in[1] io_in[0] io_in_3v3[26] io_in_3v3[25] io_in_3v3[24] io_in_3v3[23] io_in_3v3[22] io_in_3v3[21] io_in_3v3[20] io_in_3v3[19]
+ io_in_3v3[18] io_in_3v3[17] io_in_3v3[16] io_in_3v3[15] io_in_3v3[14] io_in_3v3[13] io_in_3v3[12] io_in_3v3[11] io_in_3v3[10] io_in_3v3[9]
+ io_in_3v3[8] io_in_3v3[7] io_in_3v3[6] io_in_3v3[5] io_in_3v3[4] io_in_3v3[3] io_in_3v3[2] io_in_3v3[1] io_in_3v3[0] io_out[26] io_out[25]
+ io_out[24] io_out[23] io_out[22] io_out[21] io_out[20] io_out[19] io_out[18] io_out[17] io_out[16] io_out[15] io_out[14] io_out[13]
+ io_out[12] io_out[11] io_out[10] io_out[9] io_out[8] io_out[7] io_out[6] io_out[5] io_out[4] io_out[3] io_out[2] io_out[1] io_out[0]
+ io_oeb[26] io_oeb[25] io_oeb[24] io_oeb[23] io_oeb[22] io_oeb[21] io_oeb[20] io_oeb[19] io_oeb[18] io_oeb[17] io_oeb[16] io_oeb[15]
+ io_oeb[14] io_oeb[13] io_oeb[12] io_oeb[11] io_oeb[10] io_oeb[9] io_oeb[8] io_oeb[7] io_oeb[6] io_oeb[5] io_oeb[4] io_oeb[3] io_oeb[2]
+ io_oeb[1] io_oeb[0] gpio_analog[17] gpio_analog[16] gpio_analog[15] gpio_analog[14] gpio_analog[13] gpio_analog[12] gpio_analog[11]
+ gpio_analog[10] gpio_analog[9] gpio_analog[8] gpio_analog[7] gpio_analog[6] gpio_analog[5] gpio_analog[4] gpio_analog[3] gpio_analog[2]
+ gpio_analog[1] gpio_analog[0] gpio_noesd[17] gpio_noesd[16] gpio_noesd[15] gpio_noesd[14] gpio_noesd[13] gpio_noesd[12] gpio_noesd[11]
+ gpio_noesd[10] gpio_noesd[9] gpio_noesd[8] gpio_noesd[7] gpio_noesd[6] gpio_noesd[5] gpio_noesd[4] gpio_noesd[3] gpio_noesd[2] gpio_noesd[1]
+ gpio_noesd[0] io_analog[10] io_analog[9] io_analog[8] io_analog[7] io_analog[6] io_analog[5] io_analog[4] io_analog[3] io_analog[2]
+ io_analog[1] io_analog[0] io_clamp_high[2] io_clamp_high[1] io_clamp_high[0] io_clamp_low[2] io_clamp_low[1] io_clamp_low[0] user_clock2
+ user_irq[2] user_irq[1] user_irq[0]
*.PININFO vdda1:B vdda2:B vssa1:B vssa2:B vccd1:B vccd2:B vssd1:B vssd2:B wb_clk_i:I wb_rst_i:I wbs_stb_i:I wbs_cyc_i:I wbs_we_i:I
*+ wbs_sel_i[3:0]:I wbs_dat_i[31:0]:I wbs_adr_i[31:0]:I wbs_ack_o:O wbs_dat_o[31:0]:O la_data_in[127:0]:I la_data_out[127:0]:O io_in[26:0]:I
*+ io_in_3v3[26:0]:I user_clock2:I io_out[26:0]:O io_oeb[26:0]:O gpio_analog[17:0]:B gpio_noesd[17:0]:B io_analog[10:0]:B io_clamp_high[2:0]:B
*+ io_clamp_low[2:0]:B user_irq[2:0]:O la_oenb[127:0]:I
x1 vccd1 io_analog[5] io_analog[3] io_analog[4] io_analog[1] net1 io_analog[0] io_analog[2] DS_2024_3p0
x2 vccd2 net1 io_analog[9] io_analog[10] gpio_analog[7] io_analog[8] gpio_analog[8] io_analog[7] gpio_analog[9] gpio_analog[10]
+ flashADC
x4 vccd1 io_analog[0] net1 ESD
x5 vccd1 io_analog[2] net1 ESD
x6 vccd1 io_analog[1] net1 ESD
x7 vccd1 io_analog[4] net1 ESD
x8 vccd1 io_analog[5] net1 ESD
x3 vccd1 io_analog[3] net1 ESD
x9 vccd2 io_analog[8] net1 ESD
x10 vccd2 io_analog[7] net1 ESD
x11 vccd2 io_analog[10] net1 ESD
x12 vccd2 io_analog[9] net1 ESD
R1 vssa2 net1 sky130_fd_pr__res_generic_m3 W=10 L=23.5 m=1
R2 vssa1 net1 sky130_fd_pr__res_generic_m3 W=10 L=24 m=1
.ends

* expanding   symbol:  /foss/designs/Analog_FA23_SP24/SP24_caravel_user_project_analog/xschem/xschem_DeltaSigma/DS_2024_3p0.sym #
*+ of pins=8
** sym_path: /foss/designs/Analog_FA23_SP24/SP24_caravel_user_project_analog/xschem/xschem_DeltaSigma/DS_2024_3p0.sym
** sch_path: /foss/designs/Analog_FA23_SP24/SP24_caravel_user_project_analog/xschem/xschem_DeltaSigma/DS_2024_3p0.sch
.subckt DS_2024_3p0 VDD VMID OUT VREFP VREFN GND SIG CLK
*.PININFO SIG:I CLK:I VDD:I VMID:I VREFP:I OUT:O VREFN:I GND:I
x1 VDD VMID net1 INTOUT1 GND C2S2_Amp_F_I
x2 VDD VMID net2 INTOUT2 GND C2S2_Amp_F_I
x5 VREFP VDD net3 OUT GND VREFN 1Bit_DAC_Inv
x4 VREFP VDD DACOUT OUT GND VREFN 1Bit_DAC
x3 VDD INTOUT2 OUT CLK GND VMID 1Bit_Clk_ADC
XR5 net1 SIG GND sky130_fd_pr__res_xhigh_po_5p73 L=286.5 mult=1 m=1
XR1 net2 INTOUT1 GND sky130_fd_pr__res_xhigh_po_5p73 L=286.5 mult=1 m=1
XR2 net1 net3 GND sky130_fd_pr__res_xhigh_po_5p73 L=286.5 mult=1 m=1
XR3 net2 DACOUT GND sky130_fd_pr__res_xhigh_po_5p73 L=286.5 mult=1 m=1
XC3 net2 INTOUT2 sky130_fd_pr__cap_mim_m3_1 W=15.7 L=15.7 m=12
XC1 net1 INTOUT1 sky130_fd_pr__cap_mim_m3_1 W=15.7 L=15.7 m=12
.ends


* expanding   symbol:  /foss/designs/Analog_FA23_SP24/flashADC/xschem/flashADC.sym # of pins=10
** sym_path: /foss/designs/Analog_FA23_SP24/flashADC/xschem/flashADC.sym
** sch_path: /foss/designs/Analog_FA23_SP24/flashADC/xschem/flashADC.sch
.subckt flashADC VDD GND VIN CLK OUT3 VFS OUT2 VL OUT1 OUT0
*.PININFO VDD:I GND:I VIN:I CLK:I VFS:I VL:I OUT3:O OUT2:O OUT1:O OUT0:O
XR1 VL net2 GND sky130_fd_pr__res_xhigh_po_5p73 L=2.667 mult=8 m=8
XR2 net2 net1 GND sky130_fd_pr__res_xhigh_po_5p73 L=2.667 mult=8 m=8
XR3 net1 net3 GND sky130_fd_pr__res_xhigh_po_5p73 L=2.667 mult=8 m=8
XR4 net3 net4 GND sky130_fd_pr__res_xhigh_po_5p73 L=2.667 mult=8 m=8
XR5 net4 net5 GND sky130_fd_pr__res_xhigh_po_5p73 L=2.667 mult=8 m=8
XR6 net5 net6 GND sky130_fd_pr__res_xhigh_po_5p73 L=2.667 mult=8 m=8
XR7 net6 net7 GND sky130_fd_pr__res_xhigh_po_5p73 L=2.667 mult=8 m=8
XR8 net7 net8 GND sky130_fd_pr__res_xhigh_po_5p73 L=2.667 mult=8 m=8
XR9 net8 net9 GND sky130_fd_pr__res_xhigh_po_5p73 L=2.667 mult=8 m=8
XR10 net9 net10 GND sky130_fd_pr__res_xhigh_po_5p73 L=2.667 mult=8 m=8
XR11 net10 net11 GND sky130_fd_pr__res_xhigh_po_5p73 L=2.667 mult=8 m=8
XR12 net11 net12 GND sky130_fd_pr__res_xhigh_po_5p73 L=2.667 mult=8 m=8
XR13 net12 net13 GND sky130_fd_pr__res_xhigh_po_5p73 L=2.667 mult=8 m=8
XR14 net13 net14 GND sky130_fd_pr__res_xhigh_po_5p73 L=2.667 mult=8 m=8
XR15 net14 net15 GND sky130_fd_pr__res_xhigh_po_5p73 L=2.667 mult=8 m=8
XR16 net15 net16 GND sky130_fd_pr__res_xhigh_po_5p73 L=2.667 mult=8 m=8
XR18 net16 VFS GND sky130_fd_pr__res_xhigh_po_5p73 L=2.667 mult=8 m=8
x1 OUT3 VDD net17 net18 net19 net20 net21 net22 OUT2 net23 net24 VDD net25 net26 net27 net28 OUT1 net29 net30 GND net31 net32 OUT0
+ 16to4_PriorityEncoder_v0p0p1
x18 VDD IB GND PTAT_v0p0p0
x2 VDD GND net15 VIN CLK net18 IB frontAnalog_v0p0p1
x3 VDD GND net14 VIN CLK net19 IB frontAnalog_v0p0p1
x4 VDD GND net13 VIN CLK net20 IB frontAnalog_v0p0p1
x5 VDD GND net12 VIN CLK net21 IB frontAnalog_v0p0p1
x6 VDD GND net11 VIN CLK net22 IB frontAnalog_v0p0p1
x7 VDD GND net10 VIN CLK net23 IB frontAnalog_v0p0p1
x8 VDD GND net9 VIN CLK net24 IB frontAnalog_v0p0p1
x9 VDD GND net8 VIN CLK net25 IB frontAnalog_v0p0p1
x10 VDD GND net7 VIN CLK net26 IB frontAnalog_v0p0p1
x11 VDD GND net6 VIN CLK net27 IB frontAnalog_v0p0p1
x12 VDD GND net5 VIN CLK net28 IB frontAnalog_v0p0p1
x13 VDD GND net4 VIN CLK net29 IB frontAnalog_v0p0p1
x14 VDD GND net3 VIN CLK net30 IB frontAnalog_v0p0p1
x15 VDD GND net1 VIN CLK net31 IB frontAnalog_v0p0p1
x16 VDD GND net2 VIN CLK net32 IB frontAnalog_v0p0p1
x17 VDD GND net16 VIN CLK net17 IB frontAnalog_v0p0p1
XC1 IB GND sky130_fd_pr__cap_mim_m3_2 W=30 L=30 m=72
.ends


* expanding   symbol:  /foss/designs/Analog_FA23_SP24/flashADC/xschem/ESD.sym # of pins=3
** sym_path: /foss/designs/Analog_FA23_SP24/flashADC/xschem/ESD.sym
** sch_path: /foss/designs/Analog_FA23_SP24/flashADC/xschem/ESD.sch
.subckt ESD VDD VIO VSS
*.PININFO VSS:I VDD:I VIO:B
XM24 VSS VSS VIO VSS sky130_fd_pr__nfet_01v8 L=0.2 W=500 nf=10 m=1
XM25 VIO VIO VDD VSS sky130_fd_pr__nfet_01v8 L=0.2 W=500 nf=10 m=1
.ends


* expanding   symbol:  /foss/designs/Analog_FA23_SP24/DeltaSigma/xschem/C2S2_Amp_F_I.sym # of pins=5
** sym_path: /foss/designs/Analog_FA23_SP24/DeltaSigma/xschem/C2S2_Amp_F_I.sym
** sch_path: /foss/designs/Analog_FA23_SP24/DeltaSigma/xschem/C2S2_Amp_F_I.sch
.subckt C2S2_Amp_F_I VDD VP VN OUT VSS
*.PININFO VN:I VDD:I VSS:I VP:I OUT:O
XM28 net1 net4 VSS VSS sky130_fd_pr__nfet_01v8 L=1 W=70 nf=14 m=1
XM29 net2 VN net1 VSS sky130_fd_pr__nfet_01v8 L=0.5 W=35 nf=7 m=1
XM30 net3 VP net1 VSS sky130_fd_pr__nfet_01v8 L=0.5 W=35 nf=7 m=1
XM31 net2 net2 VDD VDD sky130_fd_pr__pfet_01v8 L=0.5 W=105 nf=21 m=1
XM32 net3 net2 VDD VDD sky130_fd_pr__pfet_01v8 L=0.5 W=105 nf=21 m=1
XM38 OUT net3 VDD VDD sky130_fd_pr__pfet_01v8 L=0.5 W=200 nf=40 m=1
XM39 OUT net4 VSS VSS sky130_fd_pr__nfet_01v8 L=1 W=60 nf=12 m=1
XC2 OUT net5 sky130_fd_pr__cap_mim_m3_1 W=16 L=16 m=4
XR6 net5 net3 VSS sky130_fd_pr__res_xhigh_po_5p73 L=10.1 mult=4 m=4
XM40 net4 net6 VDD VDD sky130_fd_pr__pfet_01v8 L=1 W=30 nf=6 m=1
XM41 net6 net6 VDD VDD sky130_fd_pr__pfet_01v8 L=1 W=30 nf=6 m=1
XM42 net6 net4 net7 VSS sky130_fd_pr__nfet_01v8 L=1 W=30 nf=6 m=1
XM43 net4 net4 VSS VSS sky130_fd_pr__nfet_01v8 L=1 W=5 nf=4 m=1
XM44 net6 net6 net4 VSS sky130_fd_pr__nfet_01v8 L=0.5 W=5 nf=2 m=1
XR8 VSS net7 VSS sky130_fd_pr__res_xhigh_po_5p73 L=69 mult=4 m=4
.ends


* expanding   symbol:  /foss/designs/Analog_FA23_SP24/DeltaSigma/xschem/1Bit_DAC_Inv.sym # of pins=6
** sym_path: /foss/designs/Analog_FA23_SP24/DeltaSigma/xschem/1Bit_DAC_Inv.sym
** sch_path: /foss/designs/Analog_FA23_SP24/DeltaSigma/xschem/1Bit_DAC_Inv.sch
.subckt 1Bit_DAC_Inv VREF_P VDD OUT VIN VSS VREF_N
*.PININFO VREF_P:B VREF_N:B VSS:B VDD:B VIN:I OUT:O
XM1 VREF_N net1 OUT VDD sky130_fd_pr__pfet_01v8 L=0.15 W=95 nf=19 m=1
XM2 VREF_N VIN OUT VSS sky130_fd_pr__nfet_01v8 L=0.15 W=45 nf=9 m=1
XM3 VREF_P VIN OUT VDD sky130_fd_pr__pfet_01v8 L=0.15 W=95 nf=19 m=1
XM4 VREF_P net1 OUT VSS sky130_fd_pr__nfet_01v8 L=0.15 W=45 nf=9 m=1
XM8 net1 VIN VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=20 nf=4 m=1
XM5 net1 VIN VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=10 nf=2 m=1
.ends


* expanding   symbol:  /foss/designs/Analog_FA23_SP24/DeltaSigma/xschem/1Bit_DAC.sym # of pins=6
** sym_path: /foss/designs/Analog_FA23_SP24/DeltaSigma/xschem/1Bit_DAC.sym
** sch_path: /foss/designs/Analog_FA23_SP24/DeltaSigma/xschem/1Bit_DAC.sch
.subckt 1Bit_DAC VREF_P VDD OUT VIN VSS VREF_N
*.PININFO VREF_P:B VREF_N:B VSS:B VDD:B VIN:I OUT:O
XM1 VREF_N VIN OUT VDD sky130_fd_pr__pfet_01v8 L=0.15 W=95 nf=19 m=1
XM2 VREF_N net1 OUT VSS sky130_fd_pr__nfet_01v8 L=0.15 W=45 nf=9 m=1
XM3 VREF_P net1 OUT VDD sky130_fd_pr__pfet_01v8 L=0.15 W=95 nf=19 m=1
XM4 VREF_P VIN OUT VSS sky130_fd_pr__nfet_01v8 L=0.15 W=45 nf=9 m=1
XM8 net1 VIN VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=20 nf=4 m=1
XM5 net1 VIN VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=10 nf=2 m=1
.ends


* expanding   symbol:  /foss/designs/Analog_FA23_SP24/DeltaSigma/xschem/1Bit_Clk_ADC.sym # of pins=6
** sym_path: /foss/designs/Analog_FA23_SP24/DeltaSigma/xschem/1Bit_Clk_ADC.sym
** sch_path: /foss/designs/Analog_FA23_SP24/DeltaSigma/xschem/1Bit_Clk_ADC.sch
.subckt 1Bit_Clk_ADC VDD SIG OUT CLK VSS VMID
*.PININFO SIG:I VDD:I VSS:I CLK:I OUT:O VMID:I
x3 net4 net1 VSS VSS VDD VDD net2 sky130_fd_sc_hd__nand2_4
x4 net2 net3 VSS VSS VDD VDD net1 sky130_fd_sc_hd__nand2_4
x5 net5 CLK VSS VSS VDD VDD net4 sky130_fd_sc_hd__nand2_4
x6 CLK COMP VSS VSS VDD VDD net3 sky130_fd_sc_hd__nand2_4
x8 COMP VSS VSS VDD VDD net5 sky130_fd_sc_hd__inv_4
x9 net8 net6 VSS VSS VDD VDD OUT sky130_fd_sc_hd__nand2_4
x10 OUT net7 VSS VSS VDD VDD net6 sky130_fd_sc_hd__nand2_4
x11 net10 net9 VSS VSS VDD VDD net8 sky130_fd_sc_hd__nand2_4
x12 net9 net1 VSS VSS VDD VDD net7 sky130_fd_sc_hd__nand2_4
x14 CLK VSS VSS VDD VDD net9 sky130_fd_sc_hd__clkinv_1
x13 net1 VSS VSS VDD VDD net10 sky130_fd_sc_hd__inv_4
x1 VDD VMID SIG COMP VSS C2S2_Amp_F
.ends


* expanding   symbol:  /foss/designs/Analog_FA23_SP24/PriorityEncoder/xschem/16to4_PriorityEncoder_v0p0p1.sym # of pins=23
** sym_path: /foss/designs/Analog_FA23_SP24/PriorityEncoder/xschem/16to4_PriorityEncoder_v0p0p1.sym
** sch_path: /foss/designs/Analog_FA23_SP24/PriorityEncoder/xschem/16to4_PriorityEncoder_v0p0p1.sch
.subckt 16to4_PriorityEncoder_v0p0p1 A3 EI I15 I14 I13 I12 I11 I10 A2 I9 I8 VDD I7 I6 I5 I4 A1 I3 I2 GND I1 I0 A0
*.PININFO I14:I I13:I I12:I I11:I I10:I I9:I I8:I I7:I I6:I I5:I I4:I I3:I I2:I I1:I I0:I A3:O I15:I EI:I A2:O A1:O A0:O VDD:I
*+ GND:I
x11 net4 net5 GND GND VDD VDD net14 sky130_fd_sc_hd__or2_1
x20 net15 GND GND VDD VDD net16 sky130_fd_sc_hd__inv_1
x21 net16 GND GND VDD VDD net17 sky130_fd_sc_hd__inv_4
x22 net17 GND GND VDD VDD net13 sky130_fd_sc_hd__inv_16
x27 net18 GND GND VDD VDD net19 sky130_fd_sc_hd__inv_1
x28 net19 GND GND VDD VDD net20 sky130_fd_sc_hd__inv_4
x29 net20 GND GND VDD VDD net12 sky130_fd_sc_hd__inv_16
x34 net14 GND GND VDD VDD net21 sky130_fd_sc_hd__inv_1
x35 net21 GND GND VDD VDD net22 sky130_fd_sc_hd__inv_4
x36 net22 GND GND VDD VDD net11 sky130_fd_sc_hd__inv_16
x41 net3 GND GND VDD VDD net23 sky130_fd_sc_hd__inv_1
x42 net23 GND GND VDD VDD net24 sky130_fd_sc_hd__inv_4
x43 net24 GND GND VDD VDD net10 sky130_fd_sc_hd__inv_16
x7 net2 GND GND VDD VDD net1 sky130_fd_sc_hd__inv_1
x1 net6 net7 GND GND VDD VDD net18 sky130_fd_sc_hd__or2_1
x2 net8 net9 GND GND VDD VDD net15 sky130_fd_sc_hd__or2_1
* noconn #net25
* noconn #net26
x5 I9 I13 I11 I8 I10 I14 I15 I12 net2 net3 net4 net6 net8 EI VDD GND 8to3_Priority_Encoder_v0p2p0
x3 I1 I5 I3 I0 I2 I6 I7 I4 net25 net26 net5 net7 net9 net1 VDD GND 8to3_Priority_Encoder_v0p2p0
x6 net10 GND GND VDD VDD A3 sky130_fd_sc_hd__inv_16
x4 net10 GND GND VDD VDD A3 sky130_fd_sc_hd__inv_16
x8 net10 GND GND VDD VDD A3 sky130_fd_sc_hd__inv_16
x9 net10 GND GND VDD VDD A3 sky130_fd_sc_hd__inv_16
x10 net11 GND GND VDD VDD A2 sky130_fd_sc_hd__inv_16
x12 net11 GND GND VDD VDD A2 sky130_fd_sc_hd__inv_16
x13 net11 GND GND VDD VDD A2 sky130_fd_sc_hd__inv_16
x14 net11 GND GND VDD VDD A2 sky130_fd_sc_hd__inv_16
x15 net12 GND GND VDD VDD A1 sky130_fd_sc_hd__inv_16
x16 net12 GND GND VDD VDD A1 sky130_fd_sc_hd__inv_16
x17 net12 GND GND VDD VDD A1 sky130_fd_sc_hd__inv_16
x18 net12 GND GND VDD VDD A1 sky130_fd_sc_hd__inv_16
x19 net13 GND GND VDD VDD A0 sky130_fd_sc_hd__inv_16
x23 net13 GND GND VDD VDD A0 sky130_fd_sc_hd__inv_16
x24 net13 GND GND VDD VDD A0 sky130_fd_sc_hd__inv_16
x25 net13 GND GND VDD VDD A0 sky130_fd_sc_hd__inv_16
.ends


* expanding   symbol:  /foss/designs/Analog_FA23_SP24/PTAT/xschem/PTAT_v0p0p0.sym # of pins=3
** sym_path: /foss/designs/Analog_FA23_SP24/PTAT/xschem/PTAT_v0p0p0.sym
** sch_path: /foss/designs/Analog_FA23_SP24/PTAT/xschem/PTAT_v0p0p0.sch
.subckt PTAT_v0p0p0 VDD VOUT VSS
*.PININFO VSS:I VDD:I VOUT:O
XM1 net1 net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt L=1 W=19 nf=1 m=1
XM2 net2 net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt L=1 W=19 nf=1 m=1
XM3 VOUT net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt L=1 W=19 nf=1 m=1
XM4 net1 net1 VSS VSS sky130_fd_pr__nfet_01v8_lvt L=0.6 W=4 nf=1 m=1
XM5 net2 net1 net3 VSS sky130_fd_pr__nfet_01v8_lvt L=0.6 W=4 nf=1 m=20
XM6 net2 net2 net1 VSS sky130_fd_pr__nfet_01v8_lvt L=0.15 W=0.42 nf=1 m=1
XM7 VOUT VOUT VSS VSS sky130_fd_pr__nfet_01v8_lvt L=0.6 W=4 nf=1 m=1
XR1 VSS net3 VSS sky130_fd_pr__res_xhigh_po_5p73 L=85.94 mult=1 m=1
XR2 VSS net3 VSS sky130_fd_pr__res_xhigh_po_5p73 L=85.94 mult=1 m=1
.ends


* expanding   symbol:  /foss/designs/Analog_FA23_SP24/flashADC/xschem/frontAnalog_v0p0p1.sym # of pins=7
** sym_path: /foss/designs/Analog_FA23_SP24/flashADC/xschem/frontAnalog_v0p0p1.sym
** sch_path: /foss/designs/Analog_FA23_SP24/flashADC/xschem/frontAnalog_v0p0p1.sch
.subckt frontAnalog_v0p0p1 VDD GND VN VIN CLK Q IB
*.PININFO VDD:I GND:I VN:I VIN:I IB:I CLK:I Q:O
x63 net1 GND GND VDD VDD net3 sky130_fd_sc_hd__buf_1
x65 net2 GND GND VDD VDD net4 sky130_fd_sc_hd__buf_1
* noconn #net5
x1 VDD net3 net4 Q net5 GND RSfetsym
x2 VDD net2 net1 VN VIN CLK IB GND class_AB_v4_sym
.ends


* expanding   symbol:  /foss/designs/Analog_FA23_SP24/DeltaSigma/xschem/C2S2_Amp_F.sym # of pins=5
** sym_path: /foss/designs/Analog_FA23_SP24/DeltaSigma/xschem/C2S2_Amp_F.sym
** sch_path: /foss/designs/Analog_FA23_SP24/DeltaSigma/xschem/C2S2_Amp_F.sch
.subckt C2S2_Amp_F VDD VP VN OUT VSS
*.PININFO VN:I VDD:I VSS:I VP:I OUT:O
XM28 net1 net4 VSS VSS sky130_fd_pr__nfet_01v8 L=1 W=70 nf=14 m=1
XM29 net2 VN net1 VSS sky130_fd_pr__nfet_01v8 L=0.5 W=35 nf=7 m=1
XM30 net3 VP net1 VSS sky130_fd_pr__nfet_01v8 L=0.5 W=35 nf=7 m=1
XM31 net2 net2 VDD VDD sky130_fd_pr__pfet_01v8 L=0.5 W=105 nf=21 m=1
XM32 net3 net2 VDD VDD sky130_fd_pr__pfet_01v8 L=0.5 W=105 nf=21 m=1
XM38 OUT net3 VDD VDD sky130_fd_pr__pfet_01v8 L=0.5 W=200 nf=40 m=1
XM39 OUT net4 VSS VSS sky130_fd_pr__nfet_01v8 L=1 W=60 nf=12 m=1
XC2 OUT net5 sky130_fd_pr__cap_mim_m3_1 W=16 L=16 m=4
XR6 net5 net3 VSS sky130_fd_pr__res_xhigh_po_5p73 L=10.1 mult=4 m=4
XM40 net4 net6 VDD VDD sky130_fd_pr__pfet_01v8 L=1 W=30 nf=6 m=1
XM41 net6 net6 VDD VDD sky130_fd_pr__pfet_01v8 L=1 W=30 nf=6 m=1
XM42 net6 net4 net7 VSS sky130_fd_pr__nfet_01v8 L=1 W=30 nf=6 m=1
XM43 net4 net4 VSS VSS sky130_fd_pr__nfet_01v8 L=1 W=5 nf=4 m=1
XM44 net6 net6 net4 VSS sky130_fd_pr__nfet_01v8 L=0.5 W=5 nf=2 m=1
XR8 VSS net7 VSS sky130_fd_pr__res_xhigh_po_5p73 L=69 mult=4 m=4
.ends


* expanding   symbol:  /foss/designs/Analog_FA23_SP24/PriorityEncoder/xschem/8to3_Priority_Encoder_v0p2p0.sym # of pins=16
** sym_path: /foss/designs/Analog_FA23_SP24/PriorityEncoder/xschem/8to3_Priority_Encoder_v0p2p0.sym
** sch_path: /foss/designs/Analog_FA23_SP24/PriorityEncoder/xschem/8to3_Priority_Encoder_v0p2p0.sch
.subckt 8to3_Priority_Encoder_v0p2p0 I1 I5 I3 I0 I2 I6 I7 I4 EO GS A2 A1 A0 EI VDD GND
*.PININFO I0:I I1:I I2:I I3:I I4:I I5:I I6:I I7:I EI:I EO:O GS:O A2:O A1:O A0:O VDD:I GND:I
x9 EI GND GND VDD VDD net5 sky130_fd_sc_hd__inv_1
x1 I0 I1 I2 I3 GND GND VDD VDD net7 sky130_fd_sc_hd__or4_1
x2 I4 I5 I6 I7 GND GND VDD VDD net6 sky130_fd_sc_hd__or4_1
x4 net5 net7 net6 GND GND VDD VDD EO sky130_fd_sc_hd__or3_1
x8 EO EI GND GND VDD VDD GS sky130_fd_sc_hd__and2_1
x10 EI I4 GND GND VDD VDD net8 sky130_fd_sc_hd__and2_1
x11 EI I5 GND GND VDD VDD net9 sky130_fd_sc_hd__and2_1
x12 EI I6 GND GND VDD VDD net10 sky130_fd_sc_hd__and2_1
x13 EI I7 GND GND VDD VDD net11 sky130_fd_sc_hd__and2_1
x14 net8 net9 net10 net11 GND GND VDD VDD A2 sky130_fd_sc_hd__or4_1
x17 net10 net11 net13 net12 GND GND VDD VDD A1 sky130_fd_sc_hd__or4_1
x15 I2 net2 net3 EI GND GND VDD VDD net13 sky130_fd_sc_hd__and4_1
x16 I3 net2 net3 EI GND GND VDD VDD net12 sky130_fd_sc_hd__and4_1
x18 net2 I1 net1 net4 GND GND VDD VDD net14 sky130_fd_sc_hd__and4_1
x19 EI I3 net2 net4 GND GND VDD VDD net15 sky130_fd_sc_hd__and4_1
x20 I5 net4 EI GND GND VDD VDD net17 sky130_fd_sc_hd__and3_1
x21 EI net14 GND GND VDD VDD net16 sky130_fd_sc_hd__and2_1
x22 net11 net16 net15 net17 GND GND VDD VDD A0 sky130_fd_sc_hd__or4_1
x3 I6 GND GND VDD VDD net4 sky130_fd_sc_hd__inv_1
x5 I5 GND GND VDD VDD net3 sky130_fd_sc_hd__inv_1
x6 I4 GND GND VDD VDD net2 sky130_fd_sc_hd__inv_1
x7 I2 GND GND VDD VDD net1 sky130_fd_sc_hd__inv_1
.ends


* expanding   symbol:  /foss/designs/Analog_FA23_SP24/RSlatch/xschem/RSfetsym.sym # of pins=6
** sym_path: /foss/designs/Analog_FA23_SP24/RSlatch/xschem/RSfetsym.sym
** sch_path: /foss/designs/Analog_FA23_SP24/RSlatch/xschem/RSfetsym.sch
.subckt RSfetsym VDD S R Q QN GND
*.PININFO Q:O QN:O S:I R:I VDD:B GND:B
XM1 QN S net1 GND sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM2 net1 Q GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM3 Q R net2 GND sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM4 net2 QN GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM5 QN Q VDD VDD sky130_fd_pr__pfet_01v8 L=0.30 W=2 nf=1 m=1
XM6 Q QN VDD VDD sky130_fd_pr__pfet_01v8 L=0.30 W=2 nf=1 m=1
XM7 QN S VDD VDD sky130_fd_pr__pfet_01v8 L=0.25 W=4 nf=2 m=1
XM8 Q R VDD VDD sky130_fd_pr__pfet_01v8 L=0.25 W=4 nf=2 m=1
XM9 QN net3 GND GND sky130_fd_pr__nfet_01v8 L=0.25 W=2 nf=1 m=1
XM10 Q net4 GND GND sky130_fd_pr__nfet_01v8 L=0.25 W=2 nf=1 m=1
x2 R GND GND VDD VDD net3 sky130_fd_sc_hd__inv_4
x1 S GND GND VDD VDD net4 sky130_fd_sc_hd__inv_4
.ends


* expanding   symbol:  /foss/designs/Analog_FA23_SP24/strongARM/class_AB_v4_sym.sym # of pins=8
** sym_path: /foss/designs/Analog_FA23_SP24/strongARM/class_AB_v4_sym.sym
** sch_path: /foss/designs/Analog_FA23_SP24/strongARM/class_AB_v4_sym.sch
.subckt class_AB_v4_sym VDD VON VOP VIN VIP CLK IB VSS
*.PININFO VDD:B IB:I VSS:B VIP:I VIN:I VON:O VOP:O CLK:I
XM17 net3 VIP VIR VSS sky130_fd_pr__nfet_01v8_lvt L=0.6 W=4 nf=1 m=1
XM15 net2 VIN VIR VSS sky130_fd_pr__nfet_01v8_lvt L=0.6 W=4 nf=1 m=1
XM13 VIR IB VSS VSS sky130_fd_pr__nfet_01v8_lvt L=0.6 W=4 nf=1 m=2
XM6 VON VOP VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4 nf=1 m=1
XM7 VOP VON VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4 nf=1 m=1
XM10 VOP VON net1 VSS sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 nf=1 m=1
XM11 VON VOP net1 VSS sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 nf=1 m=1
XM1 net1 CLK VSS VSS sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 nf=1 m=1
XM2 VOP CLK VON VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4 nf=1 m=1
XM9 net2 CLK VOP VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4 nf=1 m=1
XM14 net3 CLK VON VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4 nf=1 m=1
XM3 VDD CLK net3 VSS sky130_fd_pr__nfet_01v8_lvt L=0.6 W=4 nf=1 m=1
XM4 VDD CLK net2 VSS sky130_fd_pr__nfet_01v8_lvt L=0.6 W=4 nf=1 m=1
XC1 VIP net2 VSS sky130_fd_pr__cap_var_lvt W=2 L=0.18 m=1
XC2 VIN net3 VSS sky130_fd_pr__cap_var_lvt W=2 L=0.18 m=1
.ends

.GLOBAL VDD
.GLOBAL GND
.GLOBAL VMID
.GLOBAL VREFP
.GLOBAL VREFN
.end
