* NGSPICE file created from DS_flat.ext - technology: sky130A

.subckt DS_flat GND VREFP VREFN SIG VMID OUT CLK VDD
X0 VDD.t450 a_156330_n13996.t49 a_153429_n11365.t26 VDD.t437 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X1 VDD.t159 a_216625_n11375.t32 1Bit_Clk_ADC_0.x6.B VDD.t158 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X2 a_219526_n14006.t41 a_219526_n14006.t40 VDD.t523 VDD.t46 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X3 1Bit_Clk_ADC_0.sky130_fd_sc_hd__nand2_4_0.Y 1Bit_Clk_ADC_0.x14.Y.t3 a_232253_n27658# GND.t148 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 1Bit_Clk_ADC_0.x3.B.t7 1Bit_Clk_ADC_0.x3.Y a_230965_n27658# GND.t318 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 a_216435_n47946.t1 OUT.t12 GND.t349 GND.t348 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=1.55 ps=10.62 w=5 l=0.15
X6 a_155026_n27776.t9 GND.t380 GND.t379 sky130_fd_pr__res_xhigh_po_5p73 l=69.16
X7 VREFP.t55 a_216435_n47946.t6 1Bit_DAC_0.OUT.t52 VDD.t467 sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=0.15
X8 a_156330_n13996.t45 a_156330_n13996.t44 VDD.t449 VDD.t402 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=0.5
X9 a_219318_n20038.t24 C2S2_Amp_F_I_0.OUT a_219526_n14006.t42 GND.t238 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X10 a_188130_n13996.t45 a_188130_n13996.t44 VDD.t178 VDD.t81 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X11 GND.t396 1Bit_Clk_ADC_0.x6.B 1Bit_Clk_ADC_0.x5.A GND.t395 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 1Bit_Clk_ADC_0.x11.A 1Bit_Clk_ADC_0.x3.B.t12 VDD.t133 VDD.t132 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X13 a_231797_n27343# 1Bit_Clk_ADC_0.x14.Y.t4 GND.t147 GND.t146 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X14 a_230137_n27658# CLK.t0 1Bit_Clk_ADC_0.x4.B GND.t346 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X15 a_232253_n27658# 1Bit_Clk_ADC_0.x14.Y.t5 1Bit_Clk_ADC_0.sky130_fd_sc_hd__nand2_4_0.Y GND.t145 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X16 VREFP.t54 a_216435_n47946.t7 1Bit_DAC_0.OUT.t39 VDD.t33 sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=0.15
X17 VDD.t32 a_188937_n26928.t19 a_188937_n26928.t20 VDD.t31 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X18 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t7 a_157137_n26928.t22 VDD.t74 VDD.t73 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=1
X19 1Bit_Clk_ADC_0.x6.B a_214193_n11375.t6 sky130_fd_pr__cap_mim_m3_1 l=16 w=16
X20 GND.t15 1Bit_Clk_ADC_0.x3.B.t13 1Bit_Clk_ADC_0.x11.A GND.t14 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X21 VDD.t376 a_216625_n11375.t33 1Bit_Clk_ADC_0.x6.B VDD.t375 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X22 GND.t254 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t16 a_156122_n20028.t23 GND.t253 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X23 1Bit_Clk_ADC_0.x6.B a_216625_n11375.t34 VDD.t182 VDD.t181 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X24 1Bit_Clk_ADC_0.x9.A 1Bit_Clk_ADC_0.x11.A a_231797_n27343# GND.t374 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X25 GND.t182 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t16 a_187922_n20028.t21 GND.t181 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X26 VREFP.t28 OUT.t13 1Bit_DAC_0.OUT.t5 GND.t350 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=0.15
X27 1Bit_Clk_ADC_0.x6.B a_216625_n11375.t35 VDD.t319 VDD.t318 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X28 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t7 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t6 GND.t356 GND.t355 sky130_fd_pr__nfet_01v8 ad=0.18125 pd=1.54 as=0.18125 ps=1.54 w=1.25 l=1
X29 GND.t256 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t17 C2S2_Amp_F_I_1.OUT.t24 GND.t255 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X30 VDD.t362 a_220333_n26938.t15 a_220333_n26938.t16 VDD.t212 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X31 GND.t172 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t17 a_187922_n20028.t20 GND.t171 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X32 1Bit_Clk_ADC_0.x3.A CLK.t1 VDD.t173 VDD.t172 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X33 GND.t328 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t18 C2S2_Amp_F_I_1.OUT.t23 GND.t327 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X34 a_218222_n27786.t8 GND.t378 GND.t377 sky130_fd_pr__res_xhigh_po_5p73 l=69.16
X35 a_157137_n26928.t21 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t19 a_155026_n27776.t8 GND.t329 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X36 a_216435_n47946.t5 OUT.t14 VDD.t554 VDD.t553 sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=0.15
X37 GND.t178 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t18 C2S2_Amp_F_I_0.OUT GND.t177 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X38 a_216625_n11375.t5 a_219526_n14006.t49 VDD.t47 VDD.t46 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X39 a_156330_n13996.t43 a_156330_n13996.t42 VDD.t448 VDD.t400 sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=0.5
X40 1Bit_Clk_ADC_0.x3.Y 1Bit_Clk_ADC_0.x3.B.t14 VDD.t66 VDD.t65 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X41 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t7 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t6 GND.t402 GND.t401 sky130_fd_pr__nfet_01v8 ad=0.18125 pd=1.54 as=0.3625 ps=3.08 w=1.25 l=1
X42 1Bit_Clk_ADC_0.x6.B a_216625_n11375.t36 VDD.t180 VDD.t179 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=0.5
X43 a_219526_n14006.t48 C2S2_Amp_F_I_0.OUT a_219318_n20038.t23 GND.t44 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=0.5
X44 C2S2_Amp_F_I_1.OUT.t64 a_153429_n11365.t32 VDD.t668 VDD.t667 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X45 1Bit_DAC_0.OUT.t30 a_216435_n47946.t8 VREFP.t53 VDD.t354 sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=0.15
X46 OUT.t3 1Bit_Clk_ADC_0.x9.B VDD.t239 VDD.t238 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X47 VDD.t162 a_220333_n26938.t22 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t15 VDD.t161 sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=1
X48 1Bit_DAC_Inv_0.OUT.t38 OUT.t15 VREFP.t14 VDD.t716 sky130_fd_pr__pfet_01v8 ad=1.55 pd=10.62 as=0.825 ps=5.33 w=5 l=0.15
X49 a_153429_n11365.t25 a_156330_n13996.t50 VDD.t447 VDD.t433 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X50 VDD.t282 a_219526_n14006.t38 a_219526_n14006.t39 VDD.t48 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X51 GND.t220 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t16 1Bit_Clk_ADC_0.x6.B GND.t219 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X52 GND.t222 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t17 a_219318_n20038.t13 GND.t221 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X53 VREFN.t46 a_181475_n46496.t6 1Bit_DAC_Inv_0.OUT.t43 VDD.t386 sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=0.15
X54 VDD.t196 a_188130_n13996.t49 a_185229_n11365.t23 VDD.t195 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X55 GND.t36 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t19 a_187922_n20028.t19 GND.t35 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X56 1Bit_DAC_0.OUT.t31 a_216435_n47946.t9 VREFP.t52 VDD.t372 sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=0.15
X57 VDD.t446 a_156330_n13996.t51 a_153429_n11365.t24 VDD.t431 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X58 a_156330_n13996.t41 a_156330_n13996.t40 VDD.t445 VDD.t398 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X59 1Bit_Clk_ADC_0.x3.B.t3 1Bit_Clk_ADC_0.x4.B VDD.t497 VDD.t496 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X60 VDD.t377 a_188130_n13996.t42 a_188130_n13996.t43 VDD.t83 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X61 VDD.t465 a_188130_n13996.t40 a_188130_n13996.t41 VDD.t464 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X62 GND.t411 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t18 1Bit_Clk_ADC_0.x6.B GND.t410 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X63 C2S2_Amp_F_I_0.VN.t1 a_208326_n43908# GND.t69 sky130_fd_pr__res_xhigh_po_5p73 l=57.3
X64 1Bit_Clk_ADC_0.x5.A 1Bit_Clk_ADC_0.x6.B VDD.t696 VDD.t695 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X65 a_185229_n11365.t22 a_188130_n13996.t50 VDD.t197 VDD.t89 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X66 a_185229_n11365.t0 VMID.t0 a_187922_n20028.t3 GND.t40 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X67 1Bit_DAC_0.OUT.t45 a_216435_n47946.t10 VREFP.t51 VDD.t209 sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=0.15
X68 a_156122_n20028.t4 VMID.t1 a_153429_n11365.t3 GND.t41 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X69 a_172166_n12474# C2S2_Amp_F_I_1.OUT.t0 GND.t20 sky130_fd_pr__res_xhigh_po_5p73 l=57.3
X70 a_188130_n13996.t0 C2S2_Amp_F_I_0.VN.t2 a_187922_n20028.t0 GND.t5 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X71 VDD.t321 1Bit_Clk_ADC_0.x3.B.t15 1Bit_Clk_ADC_0.sky130_fd_sc_hd__nand2_4_0.Y VDD.t320 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X72 1Bit_Clk_ADC_0.x6.B a_216625_n11375.t37 VDD.t9 VDD.t8 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X73 VDD.t495 1Bit_Clk_ADC_0.x4.B 1Bit_Clk_ADC_0.x3.B.t2 VDD.t494 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X74 a_157137_n26928.t4 a_157137_n26928.t3 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t1 GND.t32 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.58 as=0.3625 ps=2.79 w=2.5 l=0.5
X75 VDD.t694 1Bit_Clk_ADC_0.x6.B 1Bit_Clk_ADC_0.x5.A VDD.t693 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X76 1Bit_Clk_ADC_0.x6.B a_216625_n11375.t38 VDD.t139 VDD.t138 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X77 VDD.t718 OUT.t16 a_216435_n47946.t4 VDD.t717 sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=0.15
X78 VDD.t666 a_153429_n11365.t33 C2S2_Amp_F_I_1.OUT.t63 VDD.t665 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X79 a_214193_n11375.t0 a_216625_n11375.t0 GND.t4 sky130_fd_pr__res_xhigh_po_5p73 l=10.16
X80 a_150997_n11365.t6 a_153429_n11365.t29 GND.t310 sky130_fd_pr__res_xhigh_po_5p73 l=10.16
X81 C2S2_Amp_F_I_0.VN.t3 C2S2_Amp_F_I_0.OUT sky130_fd_pr__cap_mim_m3_1 l=15.7 w=15.7
X82 VDD.t49 a_219526_n14006.t50 a_216625_n11375.t6 VDD.t48 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X83 a_233081_n27658# 1Bit_Clk_ADC_0.sky130_fd_sc_hd__nand2_4_0.Y GND.t136 GND.t135 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X84 VREFP.t29 OUT.t17 1Bit_DAC_Inv_0.OUT.t37 VDD.t719 sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=0.15
X85 VDD.t508 a_216625_n11375.t39 1Bit_Clk_ADC_0.x6.B VDD.t507 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X86 GND.t394 1Bit_Clk_ADC_0.x6.B a_230137_n27658# GND.t393 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X87 a_156330_n13996.t39 a_156330_n13996.t38 VDD.t444 VDD.t396 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X88 a_188130_n13996.t39 a_188130_n13996.t38 VDD.t88 VDD.t87 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X89 1Bit_DAC_Inv_0.OUT.t45 a_181475_n46496.t7 VREFN.t45 VDD.t456 sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=0.15
X90 C2S2_Amp_F_I_1.OUT.t62 a_153429_n11365.t34 VDD.t664 VDD.t663 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X91 VDD.t274 a_185229_n11365.t32 C2S2_Amp_F_I_0.OUT VDD.t273 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X92 VREFP.t50 a_216435_n47946.t11 1Bit_DAC_0.OUT.t33 VDD.t500 sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=0.15
X93 a_153429_n11365.t1 a_150997_n11365.t0 GND.t6 sky130_fd_pr__res_xhigh_po_5p73 l=10.16
X94 VDD.t347 a_185229_n11365.t33 C2S2_Amp_F_I_0.OUT VDD.t346 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X95 a_153429_n11365.t0 VMID.t2 a_156122_n20028.t1 GND.t2 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X96 1Bit_Clk_ADC_0.x9.B OUT.t18 a_233081_n27658# GND.t339 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X97 1Bit_DAC_Inv_0.OUT.t10 a_181475_n46496.t8 VREFN.t44 VDD.t192 sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=0.15
X98 VDD.t135 1Bit_Clk_ADC_0.x14.Y.t6 1Bit_Clk_ADC_0.x9.A VDD.t134 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X99 a_188937_n26928.t18 a_188937_n26928.t17 VDD.t30 VDD.t29 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X100 a_219526_n14006.t37 a_219526_n14006.t36 VDD.t279 VDD.t38 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X101 VREFP.t49 a_216435_n47946.t12 1Bit_DAC_0.OUT.t44 VDD.t355 sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=0.15
X102 GND.t307 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t20 a_156122_n20028.t22 GND.t306 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X103 a_218222_n27786.t2 GND.t83 GND.t82 sky130_fd_pr__res_xhigh_po_5p73 l=69.16
X104 1Bit_DAC_Inv_0.OUT.t50 a_181475_n46496.t9 VREFN.t43 VDD.t518 sky130_fd_pr__pfet_01v8 ad=1.55 pd=10.62 as=0.825 ps=5.33 w=5 l=0.15
X105 a_153429_n11365.t23 a_156330_n13996.t52 VDD.t443 VDD.t429 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X106 VDD.t442 a_156330_n13996.t36 a_156330_n13996.t37 VDD.t392 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X107 VDD.t662 a_153429_n11365.t35 C2S2_Amp_F_I_1.OUT.t61 VDD.t661 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X108 GND.t413 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t19 a_219318_n20038.t25 GND.t412 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X109 VDD.t151 CLK.t2 1Bit_Clk_ADC_0.x14.Y.t0 VDD.t150 sky130_fd_pr__pfet_01v8_hvt ad=0.2352 pd=2.24 as=0.1134 ps=1.11 w=0.84 l=0.15
X110 a_196466_n47634# 1Bit_DAC_0.OUT.t28 GND.t224 sky130_fd_pr__res_xhigh_po_5p73 l=57.3
X111 1Bit_DAC_Inv_0.OUT.t18 OUT.t19 VREFN.t8 GND.t340 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=0.15
X112 GND.t176 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t4 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t5 GND.t175 sky130_fd_pr__nfet_01v8 ad=0.18125 pd=1.54 as=0.18125 ps=1.54 w=1.25 l=1
X113 GND.t309 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t21 C2S2_Amp_F_I_1.OUT.t22 GND.t308 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X114 a_187922_n20028.t18 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t20 GND.t170 GND.t169 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X115 VDD.t473 a_220333_n26938.t13 a_220333_n26938.t14 VDD.t200 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X116 a_220333_n26938.t12 a_220333_n26938.t11 VDD.t698 VDD.t198 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=1
X117 a_219526_n14006.t35 a_219526_n14006.t34 VDD.t19 VDD.t18 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X118 1Bit_Clk_ADC_0.x4.B CLK.t3 VDD.t521 VDD.t520 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X119 VDD.t588 1Bit_Clk_ADC_0.x3.A 1Bit_Clk_ADC_0.x3.Y VDD.t587 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X120 C2S2_Amp_F_I_0.OUT C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t21 GND.t34 GND.t33 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X121 a_231021_n27343# 1Bit_Clk_ADC_0.x3.B.t16 GND.t113 GND.t112 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X122 VDD.t441 a_156330_n13996.t53 a_153429_n11365.t22 VDD.t427 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X123 1Bit_Clk_ADC_0.x11.A 1Bit_Clk_ADC_0.x3.B.t17 VDD.t224 VDD.t223 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X124 a_185229_n11365.t21 a_188130_n13996.t51 VDD.t308 VDD.t228 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=0.5
X125 1Bit_Clk_ADC_0.x6.B a_216625_n11375.t40 VDD.t129 VDD.t128 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X126 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t5 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t4 GND.t80 GND.t79 sky130_fd_pr__nfet_01v8 ad=0.18125 pd=1.54 as=0.18125 ps=1.54 w=1.25 l=1
X127 1Bit_Clk_ADC_0.x6.B a_216625_n11375.t41 VDD.t131 VDD.t130 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X128 C2S2_Amp_F_I_0.OUT C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t22 GND.t174 GND.t173 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X129 1Bit_Clk_ADC_0.x9.B OUT.t20 VDD.t551 VDD.t550 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X130 a_216625_n11375.t13 VMID.t3 a_219318_n20038.t4 GND.t74 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X131 1Bit_DAC_Inv_0.OUT.t36 OUT.t21 VREFP.t31 VDD.t720 sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=0.15
X132 GND.t9 CLK.t4 a_230193_n27343# GND.t8 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X133 VDD.t71 CLK.t5 1Bit_Clk_ADC_0.x4.B VDD.t70 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X134 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t14 a_220333_n26938.t23 VDD.t164 VDD.t163 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X135 VREFN.t42 a_181475_n46496.t10 1Bit_DAC_Inv_0.OUT.t40 VDD.t294 sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=0.15
X136 VDD.t3 a_219526_n14006.t32 a_219526_n14006.t33 VDD.t2 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X137 GND.t119 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t20 a_219318_n20038.t8 GND.t118 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X138 a_186826_n27776.t7 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t23 a_188937_n26928.t21 GND.t338 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X139 a_216625_n11375.t2 a_219526_n14006.t51 VDD.t39 VDD.t38 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X140 1Bit_DAC_Inv_0.OUT.t35 OUT.t22 VREFP.t6 VDD.t721 sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=0.15
X141 VREFN.t41 a_181475_n46496.t11 1Bit_DAC_Inv_0.OUT.t1 VDD.t26 sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=0.15
X142 VDD.t660 a_153429_n11365.t36 C2S2_Amp_F_I_1.OUT.t60 VDD.t659 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X143 a_186826_n27776.t6 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t24 a_188937_n26928.t2 GND.t185 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=1
X144 VDD.t658 a_153429_n11365.t37 C2S2_Amp_F_I_1.OUT.t59 VDD.t657 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X145 a_156330_n13996.t35 a_156330_n13996.t34 VDD.t440 VDD.t390 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X146 C2S2_Amp_F_I_0.OUT a_185229_n11365.t34 VDD.t453 VDD.t452 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X147 C2S2_Amp_F_I_0.OUT a_185229_n11365.t35 VDD.t13 VDD.t12 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X148 VDD.t227 a_188130_n13996.t36 a_188130_n13996.t37 VDD.t193 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X149 VREFN.t40 a_181475_n46496.t12 1Bit_DAC_Inv_0.OUT.t48 VDD.t514 sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=0.15
X150 1Bit_Clk_ADC_0.x6.B 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t21 GND.t121 GND.t120 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X151 VDD.t122 a_188937_n26928.t22 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t15 VDD.t121 sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=1
X152 VREFN.t7 OUT.t23 1Bit_DAC_Inv_0.OUT.t12 GND.t431 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=0.15
X153 a_232253_n27658# 1Bit_Clk_ADC_0.x14.Y.t7 1Bit_Clk_ADC_0.sky130_fd_sc_hd__nand2_4_0.Y GND.t144 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X154 a_230965_n27658# 1Bit_Clk_ADC_0.x3.Y 1Bit_Clk_ADC_0.x3.B.t6 GND.t317 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X155 a_216625_n11375.t18 a_219526_n14006.t52 VDD.t275 VDD.t18 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X156 C2S2_Amp_F_I_0.OUT C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t25 GND.t429 GND.t428 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X157 a_187922_n20028.t17 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t26 GND.t162 GND.t161 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X158 1Bit_Clk_ADC_0.x6.B a_214193_n11375.t5 sky130_fd_pr__cap_mim_m3_1 l=16 w=16
X159 VREFN.t39 a_181475_n46496.t13 1Bit_DAC_Inv_0.OUT.t52 VDD.t522 sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=0.15
X160 1Bit_DAC_0.OUT.t36 a_216435_n47946.t13 VREFP.t48 VDD.t387 sky130_fd_pr__pfet_01v8 ad=1.55 pd=10.62 as=0.825 ps=5.33 w=5 l=0.15
X161 a_153429_n11365.t21 a_156330_n13996.t54 VDD.t439 VDD.t424 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X162 VDD.t438 a_156330_n13996.t32 a_156330_n13996.t33 VDD.t437 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X163 C2S2_Amp_F_I_1.OUT.t58 a_153429_n11365.t38 VDD.t656 VDD.t655 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X164 C2S2_Amp_F_I_0.OUT a_185229_n11365.t36 VDD.t351 VDD.t350 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X165 a_216625_n11375.t23 VMID.t4 a_219318_n20038.t14 GND.t238 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X166 VDD.t291 1Bit_Clk_ADC_0.x3.B.t18 1Bit_Clk_ADC_0.x11.A VDD.t290 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X167 VREFN.t27 OUT.t24 1Bit_DAC_0.OUT.t2 VDD.t552 sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=0.15
X168 VDD.t358 a_185229_n11365.t37 C2S2_Amp_F_I_0.OUT VDD.t357 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X169 VDD.t489 a_219526_n14006.t30 a_219526_n14006.t31 VDD.t43 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X170 a_188130_n13996.t2 C2S2_Amp_F_I_0.VN.t4 a_187922_n20028.t2 GND.t13 sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=0.5
X171 VDD.t436 a_156330_n13996.t55 a_153429_n11365.t20 VDD.t421 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X172 a_231797_n27343# 1Bit_Clk_ADC_0.x11.A 1Bit_Clk_ADC_0.x9.A GND.t373 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X173 VDD.t570 1Bit_Clk_ADC_0.x9.A OUT.t11 VDD.t569 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X174 1Bit_Clk_ADC_0.x3.A 1Bit_Clk_ADC_0.x5.A VDD.t578 VDD.t577 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X175 VDD.t155 a_216625_n11375.t42 1Bit_Clk_ADC_0.x6.B VDD.t154 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X176 VDD.t143 a_219526_n14006.t53 a_216625_n11375.t9 VDD.t2 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X177 VDD.t41 a_216625_n11375.t43 1Bit_Clk_ADC_0.x6.B VDD.t40 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X178 GND.t342 OUT.t25 a_181475_n46496.t1 GND.t341 sky130_fd_pr__nfet_01v8 ad=1.55 pd=10.62 as=0.825 ps=5.33 w=5 l=0.15
X179 VDD.t499 a_185229_n11365.t38 C2S2_Amp_F_I_0.OUT VDD.t498 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X180 VDD.t382 CLK.t6 1Bit_Clk_ADC_0.x3.A VDD.t381 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X181 a_174650_n12474# a_175892_n24334# GND.t57 sky130_fd_pr__res_xhigh_po_5p73 l=57.3
X182 1Bit_DAC_Inv_0.OUT.t44 a_181475_n46496.t14 VREFN.t38 VDD.t451 sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=0.15
X183 C2S2_Amp_F_I_0.OUT a_182797_n11365.t5 sky130_fd_pr__cap_mim_m3_1 l=16 w=16
X184 1Bit_Clk_ADC_0.x6.B a_216625_n11375.t44 VDD.t203 VDD.t202 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X185 1Bit_DAC_Inv_0.OUT.t11 OUT.t26 VREFN.t6 GND.t343 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=0.15
X186 C2S2_Amp_F_I_1.OUT.t57 a_153429_n11365.t39 VDD.t654 VDD.t653 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X187 a_219318_n20038.t3 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t22 GND.t66 GND.t65 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X188 VDD.t652 a_153429_n11365.t40 C2S2_Amp_F_I_1.OUT.t56 VDD.t651 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X189 a_219318_n20038.t1 VMID.t5 a_216625_n11375.t7 GND.t44 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=0.5
X190 1Bit_Clk_ADC_0.x9.B 1Bit_Clk_ADC_0.sky130_fd_sc_hd__nand2_4_0.Y VDD.t306 VDD.t305 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X191 1Bit_DAC_Inv_0.OUT.t4 a_181475_n46496.t15 VREFN.t37 VDD.t72 sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=0.15
X192 C2S2_Amp_F_I_0.OUT a_185229_n11365.t39 VDD.t37 VDD.t36 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X193 VDD.t76 a_157137_n26928.t23 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t6 VDD.t75 sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=1
X194 VREFP.t47 a_216435_n47946.t14 1Bit_DAC_0.OUT.t32 VDD.t383 sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=0.15
X195 1Bit_Clk_ADC_0.x3.A 1Bit_Clk_ADC_0.x5.A a_230193_n27343# GND.t365 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X196 a_143150_n12474# a_144392_n24334# GND.t163 sky130_fd_pr__res_xhigh_po_5p73 l=57.3
X197 VDD.t692 1Bit_Clk_ADC_0.x6.B 1Bit_Clk_ADC_0.x4.B VDD.t691 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X198 GND.t335 CLK.t7 1Bit_Clk_ADC_0.x14.Y.t1 GND.t334 sky130_fd_pr__nfet_01v8 ad=0.1197 pd=1.41 as=0.1092 ps=1.36 w=0.42 l=0.15
X199 C2S2_Amp_F_I_1.OUT.t21 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t22 GND.t258 GND.t257 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X200 1Bit_DAC_0.OUT.t0 OUT.t27 VREFN.t26 VDD.t57 sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=0.15
X201 VDD.t504 a_157137_n26928.t24 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t5 VDD.t503 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X202 VDD.t44 a_219526_n14006.t54 a_216625_n11375.t3 VDD.t43 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X203 a_219526_n14006.t29 a_219526_n14006.t28 VDD.t1 VDD.t0 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X204 C2S2_Amp_F_I_1.OUT.t55 a_153429_n11365.t41 VDD.t650 VDD.t649 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X205 GND.t260 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t23 C2S2_Amp_F_I_1.OUT.t20 GND.t259 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=1
X206 1Bit_Clk_ADC_0.x6.B 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t23 GND.t68 GND.t67 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X207 1Bit_DAC_0.OUT.t10 OUT.t28 VREFN.t25 VDD.t58 sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=0.15
X208 VDD.t304 1Bit_Clk_ADC_0.sky130_fd_sc_hd__nand2_4_0.Y 1Bit_Clk_ADC_0.x9.B VDD.t303 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X209 C2S2_Amp_F_I_1.OUT.t54 a_153429_n11365.t42 VDD.t648 VDD.t647 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X210 VDD.t435 a_156330_n13996.t56 a_153429_n11365.t19 VDD.t419 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X211 a_156330_n13996.t31 a_156330_n13996.t30 VDD.t434 VDD.t433 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X212 VDD.t471 a_185229_n11365.t40 C2S2_Amp_F_I_0.OUT VDD.t470 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X213 a_230193_n27343# 1Bit_Clk_ADC_0.x5.A 1Bit_Clk_ADC_0.x3.A GND.t364 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X214 VDD.t690 1Bit_Clk_ADC_0.x6.B 1Bit_Clk_ADC_0.x5.A VDD.t689 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X215 a_155026_n27776.t7 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t24 a_157137_n26928.t20 GND.t264 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=1
X216 a_185229_n11365.t20 a_188130_n13996.t52 VDD.t309 VDD.t111 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X217 VDD.t466 a_188130_n13996.t34 a_188130_n13996.t35 VDD.t195 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X218 a_187922_n20028.t16 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t27 GND.t184 GND.t183 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X219 VDD.t60 OUT.t29 a_181475_n46496.t5 VDD.t59 sky130_fd_pr__pfet_01v8 ad=1.55 pd=10.62 as=0.825 ps=5.33 w=5 l=0.15
X220 VDD.t241 a_185229_n11365.t41 C2S2_Amp_F_I_0.OUT VDD.t240 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X221 VDD.t432 a_156330_n13996.t28 a_156330_n13996.t29 VDD.t431 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X222 1Bit_DAC_0.OUT.t11 OUT.t30 VREFN.t24 VDD.t487 sky130_fd_pr__pfet_01v8 ad=1.55 pd=10.62 as=0.825 ps=5.33 w=5 l=0.15
X223 VDD.t108 1Bit_Clk_ADC_0.x14.Y.t8 1Bit_Clk_ADC_0.x9.A VDD.t107 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X224 a_188130_n13996.t33 a_188130_n13996.t32 VDD.t90 VDD.t89 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X225 GND.t195 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t28 a_187922_n20028.t15 GND.t194 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=1
X226 a_156330_n13996.t3 C2S2_Amp_F_I_1.VN.t2 a_156122_n20028.t6 GND.t43 sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=0.5
X227 a_187922_n20028.t6 VMID.t6 a_185229_n11365.t24 GND.t5 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X228 1Bit_DAC_0.OUT.t54 a_216435_n47946.t15 VREFN.t55 GND.t42 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=0.15
X229 C2S2_Amp_F_I_1.VN.t0 a_177926_n43908# GND.t3 sky130_fd_pr__res_xhigh_po_5p73 l=57.3
X230 a_230965_n27658# 1Bit_Clk_ADC_0.x4.B GND.t299 GND.t298 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X231 a_181475_n46496.t0 OUT.t31 GND.t291 GND.t290 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=1.55 ps=10.62 w=5 l=0.15
X232 a_172166_n12474# a_173408_n24334# GND.t427 sky130_fd_pr__res_xhigh_po_5p73 l=57.3
X233 a_187922_n20028.t27 C2S2_Amp_F_I_0.VN.t5 a_188130_n13996.t48 GND.t415 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X234 C2S2_Amp_F_I_1.VN.t3 C2S2_Amp_F_I_1.OUT.t10 sky130_fd_pr__cap_mim_m3_1 l=15.7 w=15.7
X235 VDD.t558 a_216625_n11375.t45 1Bit_Clk_ADC_0.x6.B VDD.t557 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X236 1Bit_Clk_ADC_0.x9.A 1Bit_Clk_ADC_0.x11.A VDD.t676 VDD.t675 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X237 VDD.t646 a_153429_n11365.t43 C2S2_Amp_F_I_1.OUT.t53 VDD.t645 sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=0.5
X238 a_219318_n20038.t5 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t24 GND.t76 GND.t75 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X239 a_186826_n27776.t9 GND.t426 GND.t425 sky130_fd_pr__res_xhigh_po_5p73 l=69.16
X240 1Bit_DAC_Inv_0.OUT.t2 a_181475_n46496.t16 VREFP.t1 GND.t12 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=0.15
X241 C2S2_Amp_F_I_1.VN.t4 C2S2_Amp_F_I_1.OUT.t8 sky130_fd_pr__cap_mim_m3_1 l=15.7 w=15.7
X242 GND.t85 1Bit_Clk_ADC_0.x3.B.t19 a_232253_n27658# GND.t84 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X243 1Bit_Clk_ADC_0.x3.B.t5 1Bit_Clk_ADC_0.x3.Y a_230965_n27658# GND.t316 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X244 1Bit_Clk_ADC_0.x6.B 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t25 GND.t78 GND.t77 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X245 C2S2_Amp_F_I_1.OUT.t65 a_150997_n11365.t5 sky130_fd_pr__cap_mim_m3_1 l=16 w=16
X246 1Bit_DAC_Inv_0.OUT.t3 a_181475_n46496.t17 VREFP.t2 GND.t31 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=0.15
X247 a_187922_n20028.t14 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t29 GND.t277 GND.t276 sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=1
X248 1Bit_DAC_0.OUT.t37 a_216435_n47946.t16 VREFP.t46 VDD.t328 sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=0.15
X249 1Bit_Clk_ADC_0.x6.B a_216625_n11375.t46 VDD.t704 VDD.t703 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X250 a_216625_n11375.t4 a_219526_n14006.t55 VDD.t45 VDD.t0 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X251 a_153429_n11365.t5 a_150997_n11365.t1 GND.t6 sky130_fd_pr__res_xhigh_po_5p73 l=10.16
X252 a_218222_n27786.t1 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t26 a_220333_n26938.t0 GND.t58 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=1
X253 1Bit_Clk_ADC_0.x6.B a_216625_n11375.t47 VDD.t215 VDD.t214 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X254 VREFN.t23 OUT.t32 1Bit_DAC_0.OUT.t12 VDD.t488 sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=0.15
X255 C2S2_Amp_F_I_0.OUT a_185229_n11365.t42 VDD.t243 VDD.t242 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X256 VREFN.t22 OUT.t33 1Bit_DAC_0.OUT.t22 VDD.t483 sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=0.15
X257 1Bit_DAC_0.OUT.t40 a_216435_n47946.t17 VREFP.t45 VDD.t711 sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=0.15
X258 a_219526_n14006.t47 C2S2_Amp_F_I_0.OUT a_219318_n20038.t22 GND.t239 sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=0.5
X259 1Bit_Clk_ADC_0.x9.A 1Bit_Clk_ADC_0.x11.A a_231797_n27343# GND.t372 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X260 a_181475_n46496.t4 OUT.t34 VDD.t485 VDD.t484 sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=0.15
X261 VREFN.t21 OUT.t35 1Bit_DAC_0.OUT.t9 VDD.t486 sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=0.15
X262 VDD.t644 a_153429_n11365.t44 C2S2_Amp_F_I_1.OUT.t52 VDD.t643 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X263 VREFN.t54 a_216435_n47946.t18 1Bit_DAC_0.OUT.t34 GND.t354 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=0.15
X264 C2S2_Amp_F_I_1.VN.t5 C2S2_Amp_F_I_1.OUT.t3 sky130_fd_pr__cap_mim_m3_1 l=15.7 w=15.7
X265 1Bit_Clk_ADC_0.sky130_fd_sc_hd__nand2_4_0.Y 1Bit_Clk_ADC_0.x14.Y.t9 VDD.t339 VDD.t338 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X266 1Bit_Clk_ADC_0.x3.B.t11 1Bit_Clk_ADC_0.x3.Y VDD.t531 VDD.t530 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X267 a_155026_n27776.t0 GND.t56 GND.t55 sky130_fd_pr__res_xhigh_po_5p73 l=69.16
X268 a_156330_n13996.t27 a_156330_n13996.t26 VDD.t430 VDD.t429 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X269 VREFN.t20 OUT.t36 1Bit_DAC_0.OUT.t1 VDD.t712 sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=0.15
X270 C2S2_Amp_F_I_1.OUT.t51 a_153429_n11365.t45 VDD.t642 VDD.t641 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X271 1Bit_Clk_ADC_0.x6.B a_214193_n11375.t4 sky130_fd_pr__cap_mim_m3_1 l=16 w=16
X272 a_232625_n27343# 1Bit_Clk_ADC_0.x9.B GND.t95 GND.t94 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X273 VREFP.t34 a_181475_n46496.t18 1Bit_DAC_Inv_0.OUT.t53 GND.t351 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=0.15
X274 VDD.t258 CLK.t8 1Bit_Clk_ADC_0.x4.B VDD.t257 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X275 a_166066_n47634# 1Bit_DAC_Inv_0.OUT.t41 GND.t153 sky130_fd_pr__res_xhigh_po_5p73 l=57.3
X276 C2S2_Amp_F_I_0.VN.t6 C2S2_Amp_F_I_0.OUT sky130_fd_pr__cap_mim_m3_1 l=15.7 w=15.7
X277 VDD.t556 1Bit_Clk_ADC_0.x14.Y.t10 1Bit_Clk_ADC_0.sky130_fd_sc_hd__nand2_4_0.Y VDD.t555 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X278 VDD.t344 a_188937_n26928.t15 a_188937_n26928.t16 VDD.t343 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X279 VDD.t359 a_188130_n13996.t53 a_185229_n11365.t19 VDD.t334 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X280 VDD.t709 1Bit_Clk_ADC_0.x3.B.t20 1Bit_Clk_ADC_0.x11.A VDD.t708 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X281 GND.t143 1Bit_Clk_ADC_0.x14.Y.t11 a_231797_n27343# GND.t142 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X282 VDD.t361 a_188130_n13996.t54 a_185229_n11365.t18 VDD.t360 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X283 VREFP.t32 a_181475_n46496.t19 1Bit_DAC_Inv_0.OUT.t42 GND.t154 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=0.15
X284 VDD.t428 a_156330_n13996.t24 a_156330_n13996.t25 VDD.t427 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X285 VDD.t371 a_216625_n11375.t48 1Bit_Clk_ADC_0.x6.B VDD.t370 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X286 a_188130_n13996.t31 a_188130_n13996.t30 VDD.t229 VDD.t228 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=0.5
X287 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t15 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t14 GND.t262 GND.t261 sky130_fd_pr__nfet_01v8 ad=0.18125 pd=1.54 as=0.3625 ps=3.08 w=1.25 l=1
X288 a_156330_n13996.t0 C2S2_Amp_F_I_1.VN.t6 a_156122_n20028.t0 GND.t1 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=0.5
X289 GND.t266 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t25 a_156122_n20028.t21 GND.t265 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=1
X290 a_156122_n20028.t20 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t26 GND.t251 GND.t250 sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=1
X291 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t4 a_157137_n26928.t25 VDD.t506 VDD.t505 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X292 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t14 a_188937_n26928.t23 VDD.t252 VDD.t123 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=1
X293 C2S2_Amp_F_I_1.VN.t7 C2S2_Amp_F_I_1.OUT.t12 sky130_fd_pr__cap_mim_m3_1 l=15.7 w=15.7
X294 C2S2_Amp_F_I_1.OUT.t50 a_153429_n11365.t46 VDD.t640 VDD.t639 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X295 GND.t60 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t27 1Bit_Clk_ADC_0.x6.B GND.t59 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=1
X296 a_233081_n27658# OUT.t37 1Bit_Clk_ADC_0.x9.B GND.t430 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X297 VDD.t714 OUT.t38 a_181475_n46496.t3 VDD.t713 sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=0.15
X298 C2S2_Amp_F_I_1.OUT.t49 a_153429_n11365.t47 VDD.t638 VDD.t637 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X299 VDD.t98 a_185229_n11365.t43 C2S2_Amp_F_I_0.OUT VDD.t97 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X300 1Bit_DAC_0.OUT.t14 OUT.t39 VREFN.t19 VDD.t204 sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=0.15
X301 a_155026_n27776.t3 GND.t214 GND.t213 sky130_fd_pr__res_xhigh_po_5p73 l=69.16
X302 GND.t158 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t30 a_187922_n20028.t13 GND.t157 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X303 VDD.t11 a_185229_n11365.t44 C2S2_Amp_F_I_0.OUT VDD.t10 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X304 1Bit_DAC_0.OUT.t35 a_216435_n47946.t19 VREFN.t53 GND.t159 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=0.15
X305 1Bit_DAC_Inv_0.OUT.t34 OUT.t40 VREFP.t10 VDD.t205 sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=1.55 ps=10.62 w=5 l=0.15
X306 1Bit_Clk_ADC_0.sky130_fd_sc_hd__nand2_4_0.Y 1Bit_Clk_ADC_0.x14.Y.t12 a_232253_n27658# GND.t141 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X307 1Bit_DAC_0.OUT.t24 OUT.t41 VREFN.t18 VDD.t206 sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=0.15
X308 1Bit_DAC_Inv_0.OUT.t33 OUT.t42 VREFP.t7 VDD.t56 sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=0.15
X309 a_157137_n26928.t19 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t27 a_155026_n27776.t6 GND.t252 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X310 GND.t406 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t31 C2S2_Amp_F_I_0.OUT GND.t405 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X311 GND.t107 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t28 a_219318_n20038.t6 GND.t106 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X312 a_219318_n20038.t7 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t29 GND.t109 GND.t108 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X313 a_188937_n26928.t0 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t32 a_186826_n27776.t5 GND.t21 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X314 a_182797_n11365.t0 a_185229_n11365.t2 GND.t151 sky130_fd_pr__res_xhigh_po_5p73 l=10.16
X315 VDD.t636 a_153429_n11365.t48 C2S2_Amp_F_I_1.OUT.t48 VDD.t635 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X316 VDD.t426 a_156330_n13996.t57 a_153429_n11365.t18 VDD.t415 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X317 a_156330_n13996.t23 a_156330_n13996.t22 VDD.t425 VDD.t424 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X318 a_219318_n20038.t21 C2S2_Amp_F_I_0.OUT a_219526_n14006.t46 GND.t210 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X319 C2S2_Amp_F_I_0.OUT a_185229_n11365.t45 VDD.t539 VDD.t538 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X320 a_219318_n20038.t12 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t30 GND.t216 GND.t215 sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=1
X321 1Bit_DAC_Inv_0.OUT.t5 a_181475_n46496.t20 VREFP.t3 GND.t53 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=0.15
X322 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t13 a_220333_n26938.t24 VDD.t211 VDD.t210 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X323 GND.t392 1Bit_Clk_ADC_0.x6.B a_230137_n27658# GND.t391 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X324 a_187922_n20028.t24 VMID.t7 a_185229_n11365.t27 GND.t13 sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=0.5
X325 GND.t218 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t31 1Bit_Clk_ADC_0.x6.B GND.t217 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X326 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t13 a_188937_n26928.t24 VDD.t253 VDD.t105 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X327 VDD.t423 a_156330_n13996.t58 a_153429_n11365.t17 VDD.t413 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X328 a_219526_n14006.t27 a_219526_n14006.t26 VDD.t145 VDD.t144 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X329 C2S2_Amp_F_I_0.VN.t7 C2S2_Amp_F_I_0.OUT sky130_fd_pr__cap_mim_m3_1 l=15.7 w=15.7
X330 VDD.t353 1Bit_Clk_ADC_0.x3.B.t21 1Bit_Clk_ADC_0.x3.Y VDD.t352 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X331 a_218222_n27786.t0 GND.t19 GND.t18 sky130_fd_pr__res_xhigh_po_5p73 l=69.16
X332 a_185229_n11365.t17 a_188130_n13996.t55 VDD.t285 VDD.t266 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X333 C2S2_Amp_F_I_1.VN.t8 C2S2_Amp_F_I_1.OUT.t9 sky130_fd_pr__cap_mim_m3_1 l=15.7 w=15.7
X334 VDD.t422 a_156330_n13996.t20 a_156330_n13996.t21 VDD.t421 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X335 1Bit_Clk_ADC_0.x3.A CLK.t9 VDD.t15 VDD.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X336 1Bit_DAC_0.OUT.t17 OUT.t43 VREFP.t27 GND.t27 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=0.15
X337 1Bit_Clk_ADC_0.x3.Y 1Bit_Clk_ADC_0.x3.A a_231021_n27343# GND.t369 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X338 VDD.t62 a_219526_n14006.t24 a_219526_n14006.t25 VDD.t61 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X339 a_188937_n26928.t4 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t33 a_186826_n27776.t4 GND.t196 sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=1
X340 1Bit_DAC_0.OUT.t4 OUT.t44 VREFP.t26 GND.t28 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=0.15
X341 VREFP.t13 OUT.t45 1Bit_DAC_Inv_0.OUT.t32 VDD.t367 sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=0.15
X342 1Bit_Clk_ADC_0.x6.B a_216625_n11375.t49 VDD.t560 VDD.t559 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X343 VDD.t302 1Bit_Clk_ADC_0.sky130_fd_sc_hd__nand2_4_0.Y 1Bit_Clk_ADC_0.x9.B VDD.t301 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X344 a_188937_n26928.t8 a_188937_n26928.t7 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t9 GND.t51 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.58 as=0.3625 ps=2.79 w=2.5 l=0.5
X345 a_230193_n27343# 1Bit_Clk_ADC_0.x5.A 1Bit_Clk_ADC_0.x3.A GND.t363 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X346 C2S2_Amp_F_I_1.OUT.t66 a_150997_n11365.t4 sky130_fd_pr__cap_mim_m3_1 l=16 w=16
X347 1Bit_Clk_ADC_0.x4.B 1Bit_Clk_ADC_0.x6.B VDD.t688 VDD.t687 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X348 C2S2_Amp_F_I_1.OUT.t47 a_153429_n11365.t49 VDD.t634 VDD.t633 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X349 a_231021_n27343# 1Bit_Clk_ADC_0.x3.B.t22 GND.t111 GND.t110 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X350 VDD.t127 a_185229_n11365.t46 C2S2_Amp_F_I_0.OUT VDD.t126 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X351 a_157137_n26928.t16 a_157137_n26928.t15 VDD.t533 VDD.t73 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=1
X352 C2S2_Amp_F_I_1.VN.t1 a_144392_n24334# GND.t357 sky130_fd_pr__res_xhigh_po_5p73 l=57.3
X353 1Bit_Clk_ADC_0.x9.B OUT.t46 VDD.t369 VDD.t368 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X354 a_182797_n11365.t1 a_185229_n11365.t25 GND.t151 sky130_fd_pr__res_xhigh_po_5p73 l=10.16
X355 a_219526_n14006.t23 a_219526_n14006.t22 VDD.t580 VDD.t579 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X356 a_216625_n11375.t21 a_219526_n14006.t56 VDD.t340 VDD.t144 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X357 VDD.t632 a_153429_n11365.t50 C2S2_Amp_F_I_1.OUT.t46 VDD.t631 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X358 VDD.t420 a_156330_n13996.t18 a_156330_n13996.t19 VDD.t419 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X359 VDD.t630 a_153429_n11365.t51 C2S2_Amp_F_I_1.OUT.t45 VDD.t629 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X360 a_153429_n11365.t16 a_156330_n13996.t59 VDD.t418 VDD.t410 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X361 C2S2_Amp_F_I_0.OUT a_185229_n11365.t47 VDD.t469 VDD.t468 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X362 a_188130_n13996.t29 a_188130_n13996.t28 VDD.t112 VDD.t111 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X363 C2S2_Amp_F_I_0.OUT a_185229_n11365.t48 VDD.t35 VDD.t34 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X364 GND.t23 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t32 a_219318_n20038.t0 GND.t22 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=1
X365 GND.t279 1Bit_Clk_ADC_0.x3.B.t23 a_232253_n27658# GND.t278 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X366 a_156122_n20028.t27 VMID.t8 a_153429_n11365.t30 GND.t43 sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=0.5
X367 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t3 a_157137_n26928.t26 VDD.t68 VDD.t67 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X368 a_185229_n11365.t31 VMID.t9 a_187922_n20028.t26 GND.t415 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X369 VDD.t674 1Bit_Clk_ADC_0.x11.A 1Bit_Clk_ADC_0.x9.A VDD.t673 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X370 VDD.t313 a_219526_n14006.t57 a_216625_n11375.t19 VDD.t61 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X371 VREFP.t25 OUT.t47 1Bit_DAC_0.OUT.t23 GND.t205 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=0.15
X372 1Bit_Clk_ADC_0.x6.B a_216625_n11375.t50 VDD.t265 VDD.t264 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X373 a_232253_n27658# 1Bit_Clk_ADC_0.x3.B.t24 GND.t417 GND.t416 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X374 a_156122_n20028.t19 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t28 GND.t324 GND.t323 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X375 a_230965_n27658# 1Bit_Clk_ADC_0.x3.Y 1Bit_Clk_ADC_0.x3.B.t4 GND.t315 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X376 VDD.t222 a_185229_n11365.t49 C2S2_Amp_F_I_0.OUT VDD.t221 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X377 VREFP.t24 OUT.t48 1Bit_DAC_0.OUT.t3 GND.t289 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=0.15
X378 a_196466_n45150# a_208326_n46392# GND.t69 sky130_fd_pr__res_xhigh_po_5p73 l=57.3
X379 1Bit_DAC_Inv_0.OUT.t31 OUT.t49 VREFP.t12 VDD.t480 sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=0.15
X380 VDD.t710 a_220333_n26938.t9 a_220333_n26938.t10 VDD.t161 sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=1
X381 a_216435_n47946.t3 OUT.t50 VDD.t482 VDD.t481 sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=1.55 ps=10.62 w=5 l=0.15
X382 C2S2_Amp_F_I_1.OUT.t19 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t29 GND.t326 GND.t325 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X383 GND.t140 1Bit_Clk_ADC_0.x14.Y.t13 a_231797_n27343# GND.t139 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X384 OUT.t7 1Bit_Clk_ADC_0.x9.A a_232625_n27343# GND.t361 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X385 a_157137_n26928.t18 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t30 a_155026_n27776.t5 GND.t247 sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=1
X386 VDD.t317 a_216625_n11375.t51 1Bit_Clk_ADC_0.x6.B VDD.t316 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X387 a_216625_n11375.t29 a_219526_n14006.t58 VDD.t679 VDD.t579 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X388 C2S2_Amp_F_I_1.VN.t9 C2S2_Amp_F_I_1.OUT.t7 sky130_fd_pr__cap_mim_m3_1 l=15.7 w=15.7
X389 VDD.t342 a_216625_n11375.t52 1Bit_Clk_ADC_0.x6.B VDD.t341 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X390 VDD.t628 a_153429_n11365.t52 C2S2_Amp_F_I_1.OUT.t44 VDD.t627 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X391 a_231797_n27343# 1Bit_Clk_ADC_0.x11.A 1Bit_Clk_ADC_0.x9.A GND.t371 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X392 1Bit_Clk_ADC_0.x3.A 1Bit_Clk_ADC_0.x5.A VDD.t576 VDD.t575 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X393 a_219318_n20038.t15 VMID.t10 a_216625_n11375.t24 GND.t239 sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=0.5
X394 C2S2_Amp_F_I_0.OUT a_185229_n11365.t50 VDD.t337 VDD.t336 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X395 GND.t25 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t33 1Bit_Clk_ADC_0.x6.B GND.t24 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X396 GND.t202 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t34 a_219318_n20038.t10 GND.t201 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X397 1Bit_DAC_0.OUT.t43 a_216435_n47946.t20 VREFP.t44 VDD.t548 sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=1.55 ps=10.62 w=5 l=0.15
X398 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t0 a_157137_n26928.t1 a_157137_n26928.t2 GND.t280 sky130_fd_pr__nfet_01v8 ad=0.3625 pd=2.79 as=0.725 ps=5.58 w=2.5 l=0.5
X399 a_219526_n14006.t21 a_219526_n14006.t20 VDD.t298 VDD.t297 sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=0.5
X400 VDD.t186 1Bit_Clk_ADC_0.x14.Y.t14 1Bit_Clk_ADC_0.sky130_fd_sc_hd__nand2_4_0.Y VDD.t185 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X401 VDD.t529 1Bit_Clk_ADC_0.x3.Y 1Bit_Clk_ADC_0.x3.B.t10 VDD.t528 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X402 GND.t123 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t34 a_187922_n20028.t12 GND.t122 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X403 C2S2_Amp_F_I_0.VN.t8 C2S2_Amp_F_I_0.OUT sky130_fd_pr__cap_mim_m3_1 l=15.7 w=15.7
X404 VDD.t574 1Bit_Clk_ADC_0.x5.A 1Bit_Clk_ADC_0.x3.A VDD.t573 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X405 1Bit_DAC_0.OUT.t41 a_216435_n47946.t21 VREFP.t43 VDD.t191 sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=0.15
X406 C2S2_Amp_F_I_1.OUT.t43 a_153429_n11365.t53 VDD.t626 VDD.t625 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X407 C2S2_Amp_F_I_1.OUT.t42 a_153429_n11365.t54 VDD.t624 VDD.t623 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=0.5
X408 VDD.t78 a_185229_n11365.t51 C2S2_Amp_F_I_0.OUT VDD.t77 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X409 GND.t93 1Bit_Clk_ADC_0.x9.B a_232625_n27343# GND.t92 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X410 a_218222_n27786.t6 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t35 a_220333_n26938.t19 GND.t203 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X411 a_220333_n26938.t20 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t36 a_218222_n27786.t7 GND.t283 sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=1
X412 VDD.t25 a_219526_n14006.t18 a_219526_n14006.t19 VDD.t24 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X413 1Bit_DAC_0.OUT.t25 OUT.t51 VREFP.t23 GND.t204 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=0.15
X414 a_186826_n27776.t3 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t35 a_188937_n26928.t1 GND.t86 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X415 1Bit_Clk_ADC_0.x5.A 1Bit_Clk_ADC_0.x6.B GND.t390 GND.t389 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X416 VDD.t620 a_153429_n11365.t55 C2S2_Amp_F_I_1.OUT.t41 VDD.t619 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X417 VDD.t417 a_156330_n13996.t60 a_153429_n11365.t15 VDD.t408 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X418 a_185229_n11365.t16 a_188130_n13996.t56 VDD.t286 VDD.t91 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X419 VDD.t335 a_188130_n13996.t26 a_188130_n13996.t27 VDD.t334 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X420 C2S2_Amp_F_I_0.OUT a_185229_n11365.t52 VDD.t272 VDD.t271 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X421 a_156122_n20028.t3 C2S2_Amp_F_I_1.VN.t10 a_156330_n13996.t1 GND.t39 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X422 a_185229_n11365.t15 a_188130_n13996.t57 VDD.t147 VDD.t146 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X423 VDD.t519 a_188130_n13996.t24 a_188130_n13996.t25 VDD.t360 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X424 C2S2_Amp_F_I_1.VN.t11 C2S2_Amp_F_I_1.OUT.t11 sky130_fd_pr__cap_mim_m3_1 l=15.7 w=15.7
X425 a_156122_n20028.t7 VMID.t11 a_153429_n11365.t4 GND.t1 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=0.5
X426 a_214193_n11375.t2 a_216625_n11375.t12 GND.t62 sky130_fd_pr__res_xhigh_po_5p73 l=10.16
X427 VREFP.t8 OUT.t52 1Bit_DAC_Inv_0.OUT.t30 VDD.t365 sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=0.15
X428 a_220333_n26938.t4 a_220333_n26938.t3 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t9 GND.t87 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.58 as=0.3625 ps=2.79 w=2.5 l=0.5
X429 1Bit_Clk_ADC_0.x6.B a_216625_n11375.t53 VDD.t168 VDD.t167 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X430 a_216625_n11375.t20 a_219526_n14006.t59 VDD.t331 VDD.t297 sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=0.5
X431 1Bit_DAC_Inv_0.OUT.t46 a_181475_n46496.t21 VREFN.t36 VDD.t457 sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=1.55 ps=10.62 w=5 l=0.15
X432 VDD.t622 a_153429_n11365.t56 C2S2_Amp_F_I_1.OUT.t40 VDD.t621 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X433 C2S2_Amp_F_I_1.OUT.t39 a_153429_n11365.t57 VDD.t618 VDD.t617 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X434 C2S2_Amp_F_I_0.OUT a_185229_n11365.t53 VDD.t543 VDD.t542 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X435 VREFP.t16 OUT.t53 1Bit_DAC_Inv_0.OUT.t29 VDD.t366 sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=0.15
X436 1Bit_DAC_Inv_0.OUT.t7 a_181475_n46496.t22 VREFN.t35 VDD.t137 sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=0.15
X437 VREFP.t42 a_216435_n47946.t22 1Bit_DAC_0.OUT.t53 VDD.t312 sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=0.15
X438 1Bit_Clk_ADC_0.x9.A 1Bit_Clk_ADC_0.x11.A VDD.t672 VDD.t671 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X439 GND.t297 1Bit_Clk_ADC_0.x4.B a_230965_n27658# GND.t296 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X440 GND.t249 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t31 a_156122_n20028.t18 GND.t248 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X441 VDD.t69 a_157137_n26928.t27 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t2 VDD.t63 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X442 VDD.t511 a_219526_n14006.t60 a_216625_n11375.t27 VDD.t24 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X443 a_216625_n11375.t31 a_214193_n11375.t7 GND.t414 sky130_fd_pr__res_xhigh_po_5p73 l=10.16
X444 C2S2_Amp_F_I_1.OUT.t67 a_150997_n11365.t3 sky130_fd_pr__cap_mim_m3_1 l=16 w=16
X445 a_196466_n47634# a_208326_n46392# GND.t376 sky130_fd_pr__res_xhigh_po_5p73 l=57.3
X446 VDD.t510 a_216625_n11375.t54 1Bit_Clk_ADC_0.x6.B VDD.t509 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X447 C2S2_Amp_F_I_1.OUT.t38 a_153429_n11365.t58 VDD.t616 VDD.t615 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X448 a_156122_n20028.t17 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t32 GND.t245 GND.t244 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X449 a_216625_n11375.t22 VMID.t12 a_219318_n20038.t11 GND.t210 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X450 VDD.t237 1Bit_Clk_ADC_0.x9.B OUT.t2 VDD.t236 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X451 VDD.t249 a_185229_n11365.t54 C2S2_Amp_F_I_0.OUT VDD.t248 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X452 VDD.t416 a_156330_n13996.t16 a_156330_n13996.t17 VDD.t415 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X453 a_219526_n14006.t45 C2S2_Amp_F_I_0.OUT a_219318_n20038.t20 GND.t300 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X454 a_220333_n26938.t8 a_220333_n26938.t7 VDD.t356 VDD.t163 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X455 C2S2_Amp_F_I_1.OUT.t37 a_153429_n11365.t59 VDD.t614 VDD.t613 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X456 VDD.t21 a_219526_n14006.t16 a_219526_n14006.t17 VDD.t20 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X457 a_155026_n27776.t4 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t33 a_157137_n26928.t17 GND.t246 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X458 a_219526_n14006.t15 a_219526_n14006.t14 VDD.t260 VDD.t22 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X459 VDD.t493 1Bit_Clk_ADC_0.x4.B 1Bit_Clk_ADC_0.x3.B.t1 VDD.t492 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X460 VDD.t254 a_188937_n26928.t25 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t12 VDD.t31 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X461 VDD.t414 a_156330_n13996.t14 a_156330_n13996.t15 VDD.t413 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X462 GND.t241 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t34 C2S2_Amp_F_I_1.OUT.t18 GND.t240 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X463 1Bit_Clk_ADC_0.x9.A 1Bit_Clk_ADC_0.x14.Y.t15 VDD.t188 VDD.t187 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X464 a_153429_n11365.t14 a_156330_n13996.t61 VDD.t412 VDD.t405 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X465 C2S2_Amp_F_I_0.OUT a_185229_n11365.t55 VDD.t5 VDD.t4 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X466 VDD.t28 a_216625_n11375.t55 1Bit_Clk_ADC_0.x6.B VDD.t27 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X467 a_188130_n13996.t23 a_188130_n13996.t22 VDD.t267 VDD.t266 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X468 GND.t275 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t36 C2S2_Amp_F_I_0.OUT GND.t274 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=1
X469 VDD.t149 a_188130_n13996.t58 a_185229_n11365.t14 VDD.t148 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X470 a_186826_n27776.t0 GND.t71 GND.t70 sky130_fd_pr__res_xhigh_po_5p73 l=69.16
X471 VDD.t125 a_188937_n26928.t13 a_188937_n26928.t14 VDD.t121 sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=1
X472 1Bit_Clk_ADC_0.sky130_fd_sc_hd__nand2_4_0.Y 1Bit_Clk_ADC_0.x3.B.t25 VDD.t281 VDD.t280 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X473 1Bit_Clk_ADC_0.x3.B.t9 1Bit_Clk_ADC_0.x3.Y VDD.t527 VDD.t526 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X474 a_231021_n27343# 1Bit_Clk_ADC_0.x3.A 1Bit_Clk_ADC_0.x3.Y GND.t368 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X475 GND.t285 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t37 a_219318_n20038.t16 GND.t284 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X476 1Bit_DAC_Inv_0.OUT.t28 OUT.t54 VREFP.t4 VDD.t42 sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=0.15
X477 VREFN.t34 a_181475_n46496.t23 1Bit_DAC_Inv_0.OUT.t6 VDD.t136 sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=0.15
X478 VDD.t213 a_220333_n26938.t25 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t12 VDD.t212 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X479 1Bit_DAC_0.OUT.t51 a_216435_n47946.t23 VREFP.t41 VDD.t532 sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=0.15
X480 C2S2_Amp_F_I_1.OUT.t36 a_153429_n11365.t60 VDD.t612 VDD.t611 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X481 VDD.t80 a_185229_n11365.t56 C2S2_Amp_F_I_0.OUT VDD.t79 sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=0.5
X482 VREFN.t33 a_181475_n46496.t24 1Bit_DAC_Inv_0.OUT.t49 VDD.t515 sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=0.15
X483 GND.t273 1Bit_Clk_ADC_0.x3.B.t26 a_231021_n27343# GND.t272 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X484 VREFN.t5 OUT.t55 1Bit_DAC_Inv_0.OUT.t17 GND.t16 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=1.55 ps=10.62 w=5 l=0.15
X485 a_187922_n20028.t1 C2S2_Amp_F_I_0.VN.t9 a_188130_n13996.t1 GND.t11 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X486 1Bit_Clk_ADC_0.x6.B 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t38 GND.t399 GND.t398 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X487 a_196466_n45150# a_208326_n43908# GND.t69 sky130_fd_pr__res_xhigh_po_5p73 l=57.3
X488 VREFN.t32 a_181475_n46496.t25 1Bit_DAC_Inv_0.OUT.t47 VDD.t472 sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=0.15
X489 a_218222_n27786.t9 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t39 a_220333_n26938.t21 GND.t400 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X490 C2S2_Amp_F_I_0.OUT C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t37 GND.t404 GND.t403 sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=1
X491 VREFN.t4 OUT.t56 1Bit_DAC_Inv_0.OUT.t16 GND.t17 sky130_fd_pr__nfet_01v8 ad=1.55 pd=10.62 as=0.825 ps=5.33 w=5 l=0.15
X492 GND.t134 1Bit_Clk_ADC_0.sky130_fd_sc_hd__nand2_4_0.Y a_233081_n27658# GND.t133 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X493 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t8 a_220333_n26938.t1 a_220333_n26938.t2 GND.t160 sky130_fd_pr__nfet_01v8 ad=0.3625 pd=2.79 as=0.725 ps=5.58 w=2.5 l=0.5
X494 VDD.t261 a_219526_n14006.t61 a_216625_n11375.t16 VDD.t20 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X495 a_230137_n27658# 1Bit_Clk_ADC_0.x6.B GND.t388 GND.t387 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X496 a_150997_n11365.t7 a_153429_n11365.t31 GND.t310 sky130_fd_pr__res_xhigh_po_5p73 l=10.16
X497 C2S2_Amp_F_I_1.OUT.t35 a_153429_n11365.t61 VDD.t610 VDD.t609 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X498 a_216625_n11375.t1 a_219526_n14006.t62 VDD.t23 VDD.t22 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X499 VDD.t608 a_153429_n11365.t62 C2S2_Amp_F_I_1.OUT.t34 VDD.t607 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X500 VDD.t349 a_185229_n11365.t57 C2S2_Amp_F_I_0.OUT VDD.t348 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X501 a_185229_n11365.t13 a_188130_n13996.t59 VDD.t100 VDD.t99 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X502 a_185229_n11365.t29 a_182797_n11365.t6 GND.t370 sky130_fd_pr__res_xhigh_po_5p73 l=10.16
X503 C2S2_Amp_F_I_0.OUT a_185229_n11365.t58 VDD.t247 VDD.t246 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X504 a_156330_n13996.t13 a_156330_n13996.t12 VDD.t411 VDD.t410 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X505 a_233081_n27658# OUT.t57 1Bit_Clk_ADC_0.x9.B GND.t149 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X506 GND.t198 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t38 C2S2_Amp_F_I_0.OUT GND.t197 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X507 1Bit_Clk_ADC_0.x4.B CLK.t10 a_230137_n27658# GND.t397 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X508 C2S2_Amp_F_I_1.VN.t12 C2S2_Amp_F_I_1.OUT.t2 sky130_fd_pr__cap_mim_m3_1 l=15.7 w=15.7
X509 OUT.t6 1Bit_Clk_ADC_0.x9.A a_232625_n27343# GND.t360 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X510 C2S2_Amp_F_I_0.OUT a_182797_n11365.t4 sky130_fd_pr__cap_mim_m3_1 l=16 w=16
X511 VREFP.t17 OUT.t58 1Bit_DAC_Inv_0.OUT.t27 VDD.t307 sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=0.15
X512 1Bit_DAC_Inv_0.OUT.t56 a_181475_n46496.t26 VREFN.t31 VDD.t707 sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=0.15
X513 a_140666_n12474# SIG.t0 GND.t152 sky130_fd_pr__res_xhigh_po_5p73 l=57.3
X514 VDD.t345 a_157137_n26928.t13 a_157137_n26928.t14 VDD.t75 sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=1
X515 a_186826_n27776.t1 GND.t168 GND.t167 sky130_fd_pr__res_xhigh_po_5p73 l=69.16
X516 VDD.t715 a_157137_n26928.t11 a_157137_n26928.t12 VDD.t503 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X517 1Bit_DAC_Inv_0.OUT.t8 a_181475_n46496.t27 VREFN.t30 VDD.t140 sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=0.15
X518 a_232625_n27343# 1Bit_Clk_ADC_0.x9.A OUT.t5 GND.t359 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X519 1Bit_Clk_ADC_0.x3.Y 1Bit_Clk_ADC_0.x3.A VDD.t586 VDD.t585 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X520 a_156122_n20028.t16 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t35 GND.t243 GND.t242 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X521 a_166066_n45150# a_177926_n46392# GND.t3 sky130_fd_pr__res_xhigh_po_5p73 l=57.3
X522 1Bit_Clk_ADC_0.x6.B a_216625_n11375.t56 VDD.t177 VDD.t176 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X523 1Bit_DAC_Inv_0.OUT.t14 OUT.t59 VREFN.t3 GND.t150 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=0.15
X524 1Bit_DAC_Inv_0.OUT.t39 a_181475_n46496.t28 VREFN.t29 VDD.t289 sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=0.15
X525 GND.t234 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t36 a_156122_n20028.t15 GND.t233 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X526 VREFP.t40 a_216435_n47946.t24 1Bit_DAC_0.OUT.t56 VDD.t722 sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=0.15
X527 VDD.t119 OUT.t60 1Bit_Clk_ADC_0.x9.B VDD.t118 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X528 a_155026_n27776.t2 GND.t125 GND.t124 sky130_fd_pr__res_xhigh_po_5p73 l=69.16
X529 VDD.t572 1Bit_Clk_ADC_0.x5.A 1Bit_Clk_ADC_0.x3.A VDD.t571 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X530 1Bit_Clk_ADC_0.x6.B a_216625_n11375.t57 VDD.t364 VDD.t363 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X531 1Bit_Clk_ADC_0.x11.A 1Bit_Clk_ADC_0.x3.B.t27 GND.t46 GND.t45 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X532 a_230193_n27343# CLK.t11 GND.t333 GND.t332 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X533 VDD.t541 1Bit_Clk_ADC_0.x3.B.t28 1Bit_Clk_ADC_0.x3.Y VDD.t540 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X534 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t13 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t12 GND.t268 GND.t267 sky130_fd_pr__nfet_01v8 ad=0.18125 pd=1.54 as=0.18125 ps=1.54 w=1.25 l=1
X535 a_156122_n20028.t8 C2S2_Amp_F_I_1.VN.t13 a_156330_n13996.t46 GND.t237 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X536 1Bit_DAC_0.OUT.t8 OUT.t61 VREFN.t17 VDD.t120 sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=1.55 ps=10.62 w=5 l=0.15
X537 GND.t236 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t37 a_156122_n20028.t14 GND.t235 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X538 a_188130_n13996.t3 C2S2_Amp_F_I_0.VN.t10 a_187922_n20028.t4 GND.t54 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=0.5
X539 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t3 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t2 GND.t282 GND.t281 sky130_fd_pr__nfet_01v8 ad=0.18125 pd=1.54 as=0.3625 ps=3.08 w=1.25 l=1
X540 C2S2_Amp_F_I_1.OUT.t17 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t38 GND.t320 GND.t319 sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=1
X541 VREFP.t39 a_216435_n47946.t25 1Bit_DAC_0.OUT.t38 VDD.t697 sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=0.15
X542 1Bit_DAC_Inv_0.OUT.t13 OUT.t62 VREFN.t2 GND.t49 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=0.15
X543 1Bit_DAC_0.OUT.t16 OUT.t63 VREFN.t16 VDD.t460 sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=0.15
X544 1Bit_Clk_ADC_0.sky130_fd_sc_hd__nand2_4_0.Y 1Bit_Clk_ADC_0.x14.Y.t16 VDD.t288 VDD.t287 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X545 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t11 a_188937_n26928.t26 VDD.t705 VDD.t29 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X546 GND.t322 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t39 C2S2_Amp_F_I_1.OUT.t16 GND.t321 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X547 VDD.t606 a_153429_n11365.t63 C2S2_Amp_F_I_1.OUT.t33 VDD.t605 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X548 C2S2_Amp_F_I_0.OUT a_185229_n11365.t59 VDD.t296 VDD.t295 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X549 a_232625_n27343# 1Bit_Clk_ADC_0.x9.B GND.t91 GND.t90 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X550 C2S2_Amp_F_I_0.VN.t11 C2S2_Amp_F_I_0.OUT sky130_fd_pr__cap_mim_m3_1 l=15.7 w=15.7
X551 1Bit_Clk_ADC_0.x3.Y 1Bit_Clk_ADC_0.x3.A a_231021_n27343# GND.t367 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X552 VDD.t604 a_153429_n11365.t64 C2S2_Amp_F_I_1.OUT.t32 VDD.t603 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X553 a_219318_n20038.t26 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t40 GND.t420 GND.t419 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X554 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t11 a_220333_n26938.t26 VDD.t199 VDD.t198 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=1
X555 1Bit_Clk_ADC_0.x4.B 1Bit_Clk_ADC_0.x6.B VDD.t686 VDD.t685 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X556 VDD.t201 a_220333_n26938.t27 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t10 VDD.t200 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X557 a_219526_n14006.t13 a_219526_n14006.t12 VDD.t536 VDD.t165 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X558 VDD.t101 a_188130_n13996.t60 a_185229_n11365.t12 VDD.t95 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X559 a_219318_n20038.t27 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t41 GND.t422 GND.t421 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X560 a_188937_n26928.t3 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t39 a_186826_n27776.t2 GND.t186 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X561 VDD.t409 a_156330_n13996.t10 a_156330_n13996.t11 VDD.t408 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X562 C2S2_Amp_F_I_1.OUT.t31 a_153429_n11365.t65 VDD.t602 VDD.t601 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X563 a_153429_n11365.t13 a_156330_n13996.t62 VDD.t407 VDD.t394 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X564 VDD.t109 a_188130_n13996.t61 a_185229_n11365.t11 VDD.t93 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X565 a_188130_n13996.t21 a_188130_n13996.t20 VDD.t92 VDD.t91 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X566 a_153429_n11365.t27 VMID.t13 a_156122_n20028.t9 GND.t39 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X567 a_188130_n13996.t19 a_188130_n13996.t18 VDD.t378 VDD.t146 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X568 VREFN.t1 OUT.t64 1Bit_DAC_Inv_0.OUT.t19 GND.t263 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=0.15
X569 VREFN.t28 a_181475_n46496.t29 1Bit_DAC_Inv_0.OUT.t9 VDD.t171 sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=0.15
X570 VDD.t190 a_185229_n11365.t60 C2S2_Amp_F_I_0.OUT VDD.t189 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X571 a_156330_n13996.t2 C2S2_Amp_F_I_1.VN.t14 a_156122_n20028.t5 GND.t10 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X572 VDD.t110 a_188130_n13996.t62 a_185229_n11365.t10 VDD.t16 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X573 1Bit_Clk_ADC_0.x6.B 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t42 GND.t188 GND.t187 sky130_fd_pr__nfet_01v8 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=1
X574 1Bit_Clk_ADC_0.x9.A 1Bit_Clk_ADC_0.x14.Y.t17 VDD.t220 VDD.t219 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X575 OUT.t10 1Bit_Clk_ADC_0.x9.A VDD.t568 VDD.t567 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X576 a_216625_n11375.t10 a_214193_n11375.t1 GND.t61 sky130_fd_pr__res_xhigh_po_5p73 l=10.16
X577 a_220333_n26938.t18 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t43 a_218222_n27786.t4 GND.t189 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X578 VDD.t208 a_216625_n11375.t58 1Bit_Clk_ADC_0.x6.B VDD.t207 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X579 C2S2_Amp_F_I_1.VN.t15 C2S2_Amp_F_I_1.OUT.t6 sky130_fd_pr__cap_mim_m3_1 l=15.7 w=15.7
X580 GND.t73 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t40 a_187922_n20028.t11 GND.t72 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X581 VREFN.t15 OUT.t65 1Bit_DAC_0.OUT.t20 VDD.t461 sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=0.15
X582 1Bit_DAC_0.OUT.t50 a_216435_n47946.t26 VREFP.t38 VDD.t270 sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=0.15
X583 GND.t295 1Bit_Clk_ADC_0.x4.B a_230965_n27658# GND.t294 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X584 VREFN.t0 OUT.t66 1Bit_DAC_Inv_0.OUT.t15 GND.t48 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=0.15
X585 C2S2_Amp_F_I_1.OUT.t68 a_150997_n11365.t2 sky130_fd_pr__cap_mim_m3_1 l=16 w=16
X586 VDD.t562 a_216625_n11375.t59 1Bit_Clk_ADC_0.x6.B VDD.t561 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X587 a_181475_n46496.t2 OUT.t67 VDD.t116 VDD.t115 sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=1.55 ps=10.62 w=5 l=0.15
X588 VDD.t670 1Bit_Clk_ADC_0.x11.A 1Bit_Clk_ADC_0.x9.A VDD.t669 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X589 VREFN.t14 OUT.t68 1Bit_DAC_0.OUT.t13 VDD.t117 sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=0.15
X590 VREFN.t52 a_216435_n47946.t27 1Bit_DAC_0.OUT.t42 GND.t314 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=1.55 ps=10.62 w=5 l=0.15
X591 a_232253_n27658# 1Bit_Clk_ADC_0.x3.B.t29 GND.t97 GND.t96 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X592 a_230965_n27658# 1Bit_Clk_ADC_0.x4.B GND.t293 GND.t292 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X593 VREFN.t13 OUT.t69 1Bit_DAC_0.OUT.t21 VDD.t102 sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=0.15
X594 a_218222_n27786.t5 GND.t193 GND.t192 sky130_fd_pr__res_xhigh_po_5p73 l=69.16
X595 VREFN.t51 a_216435_n47946.t28 1Bit_DAC_0.OUT.t29 GND.t0 sky130_fd_pr__nfet_01v8 ad=1.55 pd=10.62 as=0.825 ps=5.33 w=5 l=0.15
X596 VDD.t327 a_216625_n11375.t60 1Bit_Clk_ADC_0.x6.B VDD.t326 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X597 a_216625_n11375.t11 a_219526_n14006.t63 VDD.t166 VDD.t165 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X598 OUT.t1 1Bit_Clk_ADC_0.x9.B VDD.t235 VDD.t234 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X599 1Bit_Clk_ADC_0.x6.B a_216625_n11375.t61 VDD.t284 VDD.t283 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X600 a_219526_n14006.t44 C2S2_Amp_F_I_0.OUT a_219318_n20038.t19 GND.t52 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X601 VDD.t600 a_153429_n11365.t66 C2S2_Amp_F_I_1.OUT.t30 VDD.t599 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X602 C2S2_Amp_F_I_0.VN.t12 C2S2_Amp_F_I_0.OUT sky130_fd_pr__cap_mim_m3_1 l=15.7 w=15.7
X603 a_166066_n47634# a_177926_n46392# GND.t81 sky130_fd_pr__res_xhigh_po_5p73 l=57.3
X604 a_157137_n26928.t10 a_157137_n26928.t9 VDD.t544 VDD.t505 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X605 a_219318_n20038.t17 VMID.t14 a_216625_n11375.t26 GND.t300 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X606 C2S2_Amp_F_I_0.OUT a_182797_n11365.t3 sky130_fd_pr__cap_mim_m3_1 l=16 w=16
X607 C2S2_Amp_F_I_0.OUT a_185229_n11365.t61 VDD.t502 VDD.t501 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X608 1Bit_Clk_ADC_0.sky130_fd_sc_hd__nand2_4_0.Y 1Bit_Clk_ADC_0.x3.B.t30 VDD.t459 VDD.t458 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X609 a_188937_n26928.t12 a_188937_n26928.t11 VDD.t124 VDD.t123 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=1
X610 VREFP.t0 a_181475_n46496.t30 1Bit_DAC_Inv_0.OUT.t0 GND.t7 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=1.55 ps=10.62 w=5 l=0.15
X611 VDD.t678 a_219526_n14006.t10 a_219526_n14006.t11 VDD.t262 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X612 GND.t345 CLK.t12 a_230193_n27343# GND.t344 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X613 1Bit_Clk_ADC_0.x5.A 1Bit_Clk_ADC_0.x6.B VDD.t684 VDD.t683 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X614 VDD.t315 a_219526_n14006.t8 a_219526_n14006.t9 VDD.t314 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X615 a_156330_n13996.t9 a_156330_n13996.t8 VDD.t406 VDD.t405 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X616 VREFP.t33 a_181475_n46496.t31 1Bit_DAC_Inv_0.OUT.t51 GND.t311 sky130_fd_pr__nfet_01v8 ad=1.55 pd=10.62 as=0.825 ps=5.33 w=5 l=0.15
X617 VDD.t404 a_156330_n13996.t63 a_153429_n11365.t12 VDD.t388 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X618 a_185229_n11365.t9 a_188130_n13996.t63 VDD.t51 VDD.t50 sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=0.5
X619 C2S2_Amp_F_I_0.VN.t13 C2S2_Amp_F_I_0.OUT sky130_fd_pr__cap_mim_m3_1 l=15.7 w=15.7
X620 GND.t313 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t10 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t11 GND.t312 sky130_fd_pr__nfet_01v8 ad=0.18125 pd=1.54 as=0.18125 ps=1.54 w=1.25 l=1
X621 a_156122_n20028.t13 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t40 GND.t230 GND.t229 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X622 VDD.t259 a_188130_n13996.t16 a_188130_n13996.t17 VDD.t148 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X623 VDD.t245 1Bit_Clk_ADC_0.x3.B.t31 1Bit_Clk_ADC_0.sky130_fd_sc_hd__nand2_4_0.Y VDD.t244 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X624 GND.t200 1Bit_Clk_ADC_0.x3.B.t32 a_231021_n27343# GND.t199 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X625 a_185229_n11365.t8 a_188130_n13996.t64 VDD.t53 VDD.t52 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X626 1Bit_DAC_0.OUT.t27 OUT.t70 VREFN.t12 VDD.t103 sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=0.15
X627 VREFP.t37 a_216435_n47946.t29 1Bit_DAC_0.OUT.t48 VDD.t545 sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=0.15
X628 VDD.t525 1Bit_Clk_ADC_0.x3.Y 1Bit_Clk_ADC_0.x3.B.t8 VDD.t524 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X629 a_188130_n13996.t47 C2S2_Amp_F_I_0.VN.t14 a_187922_n20028.t22 GND.t305 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X630 GND.t89 1Bit_Clk_ADC_0.x9.B a_232625_n27343# GND.t88 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X631 VDD.t218 a_219526_n14006.t6 a_219526_n14006.t7 VDD.t216 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X632 C2S2_Amp_F_I_1.OUT.t15 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t41 GND.t232 GND.t231 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X633 GND.t226 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t42 a_156122_n20028.t12 GND.t225 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X634 1Bit_DAC_0.OUT.t19 OUT.t71 VREFN.t11 VDD.t104 sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=0.15
X635 a_153429_n11365.t11 a_156330_n13996.t64 VDD.t403 VDD.t402 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=0.5
X636 C2S2_Amp_F_I_1.OUT.t14 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t43 GND.t228 GND.t227 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X637 a_185229_n11365.t7 a_188130_n13996.t65 VDD.t82 VDD.t81 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X638 VDD.t256 a_216625_n11375.t62 1Bit_Clk_ADC_0.x6.B VDD.t255 sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=0.5
X639 a_187922_n20028.t10 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t41 GND.t30 GND.t29 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X640 1Bit_DAC_0.OUT.t15 OUT.t72 VREFN.t10 VDD.t113 sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=0.15
X641 a_220333_n26938.t6 a_220333_n26938.t5 VDD.t278 VDD.t210 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X642 1Bit_DAC_0.OUT.t49 a_216435_n47946.t30 VREFN.t50 GND.t336 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=0.15
X643 a_185229_n11365.t28 VMID.t15 a_187922_n20028.t25 GND.t11 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X644 1Bit_Clk_ADC_0.x5.A 1Bit_Clk_ADC_0.x6.B GND.t386 GND.t385 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X645 a_188937_n26928.t10 a_188937_n26928.t9 VDD.t106 VDD.t105 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X646 1Bit_Clk_ADC_0.x4.B CLK.t13 a_230137_n27658# GND.t347 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X647 a_155026_n27776.t1 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t44 a_157137_n26928.t0 GND.t98 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X648 C2S2_Amp_F_I_0.OUT C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t42 GND.t165 GND.t164 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X649 a_166066_n45150# a_177926_n43908# GND.t3 sky130_fd_pr__res_xhigh_po_5p73 l=57.3
X650 VDD.t263 a_219526_n14006.t64 a_216625_n11375.t17 VDD.t262 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X651 1Bit_DAC_0.OUT.t46 a_216435_n47946.t31 VREFN.t49 GND.t166 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=0.15
X652 1Bit_Clk_ADC_0.x11.A 1Bit_Clk_ADC_0.x3.B.t33 GND.t103 GND.t102 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X653 1Bit_Clk_ADC_0.x6.B a_216625_n11375.t63 VDD.t86 VDD.t85 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X654 GND.t191 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t2 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t3 GND.t190 sky130_fd_pr__nfet_01v8 ad=0.18125 pd=1.54 as=0.18125 ps=1.54 w=1.25 l=1
X655 VDD.t479 a_219526_n14006.t65 a_216625_n11375.t25 VDD.t314 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X656 GND.t384 1Bit_Clk_ADC_0.x6.B 1Bit_Clk_ADC_0.x5.A GND.t383 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X657 a_188130_n13996.t15 a_188130_n13996.t14 VDD.t160 VDD.t99 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X658 1Bit_Clk_ADC_0.x14.Y.t2 CLK.t14 VDD.t547 VDD.t546 sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.11 as=0.2184 ps=2.2 w=0.84 l=0.15
X659 1Bit_Clk_ADC_0.x9.B OUT.t73 a_233081_n27658# GND.t47 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X660 C2S2_Amp_F_I_1.OUT.t29 a_153429_n11365.t67 VDD.t598 VDD.t597 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X661 VDD.t535 a_185229_n11365.t62 C2S2_Amp_F_I_0.OUT VDD.t534 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X662 GND.t115 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t44 1Bit_Clk_ADC_0.x6.B GND.t114 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X663 GND.t304 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t0 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t1 GND.t303 sky130_fd_pr__nfet_01v8 ad=0.3625 pd=3.08 as=0.18125 ps=1.54 w=1.25 l=1
X664 a_230137_n27658# CLK.t15 1Bit_Clk_ADC_0.x4.B GND.t269 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X665 VDD.t251 a_185229_n11365.t63 C2S2_Amp_F_I_0.OUT VDD.t250 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X666 1Bit_DAC_Inv_0.OUT.t54 a_181475_n46496.t32 VREFP.t35 GND.t352 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=0.15
X667 1Bit_Clk_ADC_0.x6.B 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t45 GND.t117 GND.t116 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X668 a_220333_n26938.t17 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t46 a_218222_n27786.t3 GND.t126 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X669 a_187922_n20028.t9 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t43 GND.t271 GND.t270 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X670 VDD.t217 a_219526_n14006.t66 a_216625_n11375.t14 VDD.t216 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X671 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t8 a_188937_n26928.t5 a_188937_n26928.t6 GND.t50 sky130_fd_pr__nfet_01v8 ad=0.3625 pd=2.79 as=0.725 ps=5.58 w=2.5 l=0.5
X672 a_153429_n11365.t10 a_156330_n13996.t65 VDD.t401 VDD.t400 sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=0.5
X673 C2S2_Amp_F_I_0.VN.t0 a_175892_n24334# GND.t105 sky130_fd_pr__res_xhigh_po_5p73 l=57.3
X674 VDD.t596 a_153429_n11365.t68 C2S2_Amp_F_I_1.OUT.t28 VDD.t595 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X675 C2S2_Amp_F_I_0.OUT a_185229_n11365.t64 VDD.t517 VDD.t516 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=0.5
X676 C2S2_Amp_F_I_0.VN.t15 C2S2_Amp_F_I_0.OUT sky130_fd_pr__cap_mim_m3_1 l=15.7 w=15.7
X677 VDD.t584 1Bit_Clk_ADC_0.x3.A 1Bit_Clk_ADC_0.x3.Y VDD.t583 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X678 a_140666_n12474# a_141908_n24334# GND.t409 sky130_fd_pr__res_xhigh_po_5p73 l=57.3
X679 a_185229_n11365.t30 a_182797_n11365.t7 GND.t375 sky130_fd_pr__res_xhigh_po_5p73 l=10.16
X680 a_219526_n14006.t5 a_219526_n14006.t4 VDD.t537 VDD.t230 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X681 C2S2_Amp_F_I_0.OUT C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t44 GND.t180 GND.t179 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X682 VREFN.t9 OUT.t74 1Bit_DAC_0.OUT.t18 VDD.t114 sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=0.15
X683 VREFN.t48 a_216435_n47946.t32 1Bit_DAC_0.OUT.t55 GND.t337 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=0.15
X684 VREFP.t5 OUT.t75 1Bit_DAC_Inv_0.OUT.t26 VDD.t54 sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=0.15
X685 a_231797_n27343# 1Bit_Clk_ADC_0.x14.Y.t18 GND.t138 GND.t137 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X686 a_219526_n14006.t3 a_219526_n14006.t2 VDD.t153 VDD.t152 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=0.5
X687 a_153429_n11365.t9 a_156330_n13996.t66 VDD.t399 VDD.t398 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X688 VDD.t84 a_188130_n13996.t66 a_185229_n11365.t6 VDD.t83 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X689 GND.t64 1Bit_Clk_ADC_0.x3.B.t34 1Bit_Clk_ADC_0.x11.A GND.t63 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X690 1Bit_Clk_ADC_0.x3.Y 1Bit_Clk_ADC_0.x3.B.t35 VDD.t277 VDD.t276 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X691 1Bit_Clk_ADC_0.x6.B a_216625_n11375.t64 VDD.t184 VDD.t183 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X692 1Bit_Clk_ADC_0.x6.B a_214193_n11375.t3 sky130_fd_pr__cap_mim_m3_1 l=16 w=16
X693 C2S2_Amp_F_I_1.VN.t16 C2S2_Amp_F_I_1.OUT.t4 sky130_fd_pr__cap_mim_m3_1 l=15.7 w=15.7
X694 VDD.t325 a_185229_n11365.t65 C2S2_Amp_F_I_0.OUT VDD.t324 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X695 VDD.t512 a_188130_n13996.t67 a_185229_n11365.t5 VDD.t464 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X696 1Bit_Clk_ADC_0.x6.B a_216625_n11375.t65 VDD.t269 VDD.t268 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X697 VREFN.t47 a_216435_n47946.t33 1Bit_DAC_0.OUT.t47 GND.t101 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=0.15
X698 VREFP.t18 OUT.t76 1Bit_DAC_Inv_0.OUT.t25 VDD.t55 sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=0.15
X699 a_153429_n11365.t28 VMID.t16 a_156122_n20028.t24 GND.t237 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X700 a_157137_n26928.t8 a_157137_n26928.t7 VDD.t549 VDD.t67 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X701 a_187922_n20028.t7 C2S2_Amp_F_I_0.VN.t16 a_188130_n13996.t46 GND.t40 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X702 a_156330_n13996.t48 C2S2_Amp_F_I_1.VN.t17 a_156122_n20028.t26 GND.t41 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X703 C2S2_Amp_F_I_0.VN.t17 C2S2_Amp_F_I_0.OUT sky130_fd_pr__cap_mim_m3_1 l=15.7 w=15.7
X704 a_187922_n20028.t5 VMID.t17 a_185229_n11365.t1 GND.t54 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=0.5
X705 VREFP.t36 a_181475_n46496.t33 1Bit_DAC_Inv_0.OUT.t55 GND.t353 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=0.15
X706 VDD.t157 a_216625_n11375.t66 1Bit_Clk_ADC_0.x6.B VDD.t156 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X707 1Bit_Clk_ADC_0.x3.B.t0 1Bit_Clk_ADC_0.x4.B VDD.t491 VDD.t490 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X708 a_231021_n27343# 1Bit_Clk_ADC_0.x3.A 1Bit_Clk_ADC_0.x3.Y GND.t366 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X709 VDD.t594 a_153429_n11365.t69 C2S2_Amp_F_I_1.OUT.t27 VDD.t593 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X710 GND.t331 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t8 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t9 GND.t330 sky130_fd_pr__nfet_01v8 ad=0.3625 pd=3.08 as=0.18125 ps=1.54 w=1.25 l=1
X711 VDD.t7 a_185229_n11365.t66 C2S2_Amp_F_I_0.OUT VDD.t6 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X712 C2S2_Amp_F_I_1.VN.t18 C2S2_Amp_F_I_1.OUT.t5 sky130_fd_pr__cap_mim_m3_1 l=15.7 w=15.7
X713 C2S2_Amp_F_I_0.OUT a_185229_n11365.t67 VDD.t385 VDD.t384 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X714 a_156122_n20028.t11 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t45 GND.t100 GND.t99 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X715 VDD.t142 a_219526_n14006.t0 a_219526_n14006.t1 VDD.t141 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X716 OUT.t9 1Bit_Clk_ADC_0.x9.A VDD.t566 VDD.t565 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X717 a_216625_n11375.t15 a_219526_n14006.t67 VDD.t231 VDD.t230 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X718 a_216625_n11375.t30 a_219526_n14006.t68 VDD.t680 VDD.t152 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=1.45 ps=10.58 w=5 l=0.5
X719 VDD.t706 a_188937_n26928.t27 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t10 VDD.t343 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X720 a_153429_n11365.t8 a_156330_n13996.t67 VDD.t397 VDD.t396 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X721 a_156122_n20028.t10 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t46 GND.t207 GND.t206 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X722 VDD.t96 a_188130_n13996.t12 a_188130_n13996.t13 VDD.t95 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X723 VREFP.t22 OUT.t77 1Bit_DAC_0.OUT.t6 GND.t26 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=1.55 ps=10.62 w=5 l=0.15
X724 C2S2_Amp_F_I_0.OUT a_182797_n11365.t2 sky130_fd_pr__cap_mim_m3_1 l=16 w=16
X725 VDD.t592 a_153429_n11365.t70 C2S2_Amp_F_I_1.OUT.t26 VDD.t591 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X726 C2S2_Amp_F_I_0.OUT a_185229_n11365.t68 VDD.t702 VDD.t701 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X727 a_185229_n11365.t4 a_188130_n13996.t68 VDD.t513 VDD.t87 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X728 GND.t132 1Bit_Clk_ADC_0.sky130_fd_sc_hd__nand2_4_0.Y a_233081_n27658# GND.t131 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X729 1Bit_DAC_Inv_0.OUT.t24 OUT.t78 VREFP.t9 VDD.t477 sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=0.15
X730 a_174650_n12474# a_173408_n24334# GND.t418 sky130_fd_pr__res_xhigh_po_5p73 l=57.3
X731 a_187922_n20028.t8 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t45 GND.t212 GND.t211 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X732 C2S2_Amp_F_I_0.OUT a_185229_n11365.t69 VDD.t455 VDD.t454 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X733 a_156330_n13996.t7 a_156330_n13996.t6 VDD.t395 VDD.t394 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X734 a_230137_n27658# 1Bit_Clk_ADC_0.x6.B GND.t382 GND.t381 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X735 a_156122_n20028.t2 VMID.t18 a_153429_n11365.t2 GND.t10 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X736 VDD.t94 a_188130_n13996.t10 a_188130_n13996.t11 VDD.t93 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X737 VREFP.t21 OUT.t79 1Bit_DAC_0.OUT.t26 GND.t288 sky130_fd_pr__nfet_01v8 ad=1.55 pd=10.62 as=0.825 ps=5.33 w=5 l=0.15
X738 VDD.t564 1Bit_Clk_ADC_0.x9.A OUT.t8 VDD.t563 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X739 C2S2_Amp_F_I_1.OUT.t13 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t47 GND.t209 GND.t208 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X740 VDD.t17 a_188130_n13996.t8 a_188130_n13996.t9 VDD.t16 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X741 C2S2_Amp_F_I_0.VN.t18 C2S2_Amp_F_I_0.OUT sky130_fd_pr__cap_mim_m3_1 l=15.7 w=15.7
X742 a_156122_n20028.t25 C2S2_Amp_F_I_1.VN.t19 a_156330_n13996.t47 GND.t2 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X743 1Bit_DAC_Inv_0.OUT.t23 OUT.t80 VREFP.t11 VDD.t478 sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=0.15
X744 a_233081_n27658# 1Bit_Clk_ADC_0.sky130_fd_sc_hd__nand2_4_0.Y GND.t130 GND.t129 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X745 VDD.t393 a_156330_n13996.t68 a_153429_n11365.t7 VDD.t392 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X746 a_143150_n12474# a_141908_n24334# GND.t104 sky130_fd_pr__res_xhigh_po_5p73 l=57.3
X747 1Bit_DAC_Inv_0.OUT.t22 OUT.t81 VREFP.t15 VDD.t474 sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=0.15
X748 GND.t424 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t0 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t1 GND.t423 sky130_fd_pr__nfet_01v8 ad=0.3625 pd=3.08 as=0.18125 ps=1.54 w=1.25 l=1
X749 1Bit_Clk_ADC_0.x6.B a_216625_n11375.t67 VDD.t374 VDD.t373 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X750 GND.t302 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t46 C2S2_Amp_F_I_0.OUT GND.t301 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X751 a_219318_n20038.t9 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t47 GND.t128 GND.t127 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X752 a_186826_n27776.t8 GND.t408 GND.t407 sky130_fd_pr__res_xhigh_po_5p73 l=69.16
X753 VDD.t311 CLK.t16 1Bit_Clk_ADC_0.x3.A VDD.t310 sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X754 C2S2_Amp_F_I_1.VN.t20 C2S2_Amp_F_I_1.OUT.t1 sky130_fd_pr__cap_mim_m3_1 l=15.7 w=15.7
X755 GND.t287 OUT.t82 a_216435_n47946.t0 GND.t286 sky130_fd_pr__nfet_01v8 ad=1.55 pd=10.62 as=0.825 ps=5.33 w=5 l=0.15
X756 VDD.t677 a_219526_n14006.t69 a_216625_n11375.t28 VDD.t141 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X757 1Bit_Clk_ADC_0.x9.B 1Bit_Clk_ADC_0.sky130_fd_sc_hd__nand2_4_0.Y VDD.t300 VDD.t299 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X758 VDD.t233 1Bit_Clk_ADC_0.x9.B OUT.t0 VDD.t232 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X759 VDD.t226 a_216625_n11375.t68 1Bit_Clk_ADC_0.x6.B VDD.t225 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X760 VDD.t682 1Bit_Clk_ADC_0.x6.B 1Bit_Clk_ADC_0.x4.B VDD.t681 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X761 a_232625_n27343# 1Bit_Clk_ADC_0.x9.A OUT.t4 GND.t358 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X762 1Bit_Clk_ADC_0.x3.A 1Bit_Clk_ADC_0.x5.A a_230193_n27343# GND.t362 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X763 1Bit_Clk_ADC_0.x3.Y 1Bit_Clk_ADC_0.x3.A VDD.t582 VDD.t581 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X764 VDD.t323 a_216625_n11375.t69 1Bit_Clk_ADC_0.x6.B VDD.t322 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X765 VDD.t330 a_216625_n11375.t70 1Bit_Clk_ADC_0.x6.B VDD.t329 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X766 a_219318_n20038.t2 VMID.t19 a_216625_n11375.t8 GND.t52 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X767 VDD.t170 a_216625_n11375.t71 1Bit_Clk_ADC_0.x6.B VDD.t169 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X768 a_219318_n20038.t18 C2S2_Amp_F_I_0.OUT a_219526_n14006.t43 GND.t74 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X769 C2S2_Amp_F_I_0.VN.t19 C2S2_Amp_F_I_0.OUT sky130_fd_pr__cap_mim_m3_1 l=15.7 w=15.7
X770 VDD.t476 OUT.t83 1Bit_Clk_ADC_0.x9.B VDD.t475 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X771 GND.t156 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t47 C2S2_Amp_F_I_0.OUT GND.t155 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X772 a_230193_n27343# CLK.t17 GND.t38 GND.t37 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X773 1Bit_Clk_ADC_0.x4.B CLK.t18 VDD.t463 VDD.t462 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X774 1Bit_DAC_0.OUT.t7 OUT.t84 VREFP.t20 GND.t223 sky130_fd_pr__nfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=0.15
X775 a_153429_n11365.t6 a_156330_n13996.t69 VDD.t391 VDD.t390 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X776 C2S2_Amp_F_I_1.OUT.t25 a_153429_n11365.t71 VDD.t590 VDD.t589 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X777 C2S2_Amp_F_I_0.OUT a_185229_n11365.t70 VDD.t175 VDD.t174 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X778 VREFP.t19 OUT.t85 1Bit_DAC_Inv_0.OUT.t21 VDD.t379 sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=0.15
X779 VDD.t194 a_188130_n13996.t69 a_185229_n11365.t3 VDD.t193 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X780 VDD.t293 a_185229_n11365.t71 C2S2_Amp_F_I_0.OUT VDD.t292 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X781 VDD.t389 a_156330_n13996.t4 a_156330_n13996.t5 VDD.t388 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X782 a_188130_n13996.t7 a_188130_n13996.t6 VDD.t333 VDD.t50 sky130_fd_pr__pfet_01v8 ad=1.45 pd=10.58 as=0.725 ps=5.29 w=5 l=0.5
X783 VREFP.t30 OUT.t86 1Bit_DAC_Inv_0.OUT.t20 VDD.t380 sky130_fd_pr__pfet_01v8 ad=0.825 pd=5.33 as=0.825 ps=5.33 w=5 l=0.15
X784 a_188130_n13996.t5 a_188130_n13996.t4 VDD.t332 VDD.t52 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X785 a_187922_n20028.t23 VMID.t20 a_185229_n11365.t26 GND.t305 sky130_fd_pr__nfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=0.5
X786 VDD.t700 OUT.t87 a_216435_n47946.t2 VDD.t699 sky130_fd_pr__pfet_01v8 ad=1.55 pd=10.62 as=0.825 ps=5.33 w=5 l=0.15
X787 VDD.t64 a_157137_n26928.t5 a_157137_n26928.t6 VDD.t63 sky130_fd_pr__pfet_01v8 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=1
X788 C2S2_Amp_F_I_0.VN.t20 C2S2_Amp_F_I_0.OUT sky130_fd_pr__cap_mim_m3_1 l=15.7 w=15.7
R0 a_156330_n13996.n80 a_156330_n13996.n62 585
R1 a_156330_n13996.n80 a_156330_n13996.n61 585
R2 a_156330_n13996.n80 a_156330_n13996.n60 585
R3 a_156330_n13996.n80 a_156330_n13996.n58 585
R4 a_156330_n13996.n80 a_156330_n13996.n57 585
R5 a_156330_n13996.n80 a_156330_n13996.n56 585
R6 a_156330_n13996.n80 a_156330_n13996.n53 585
R7 a_156330_n13996.n80 a_156330_n13996.n28 291.375
R8 a_156330_n13996.n95 a_156330_n13996.n51 585
R9 a_156330_n13996.n95 a_156330_n13996.n50 585
R10 a_156330_n13996.n95 a_156330_n13996.n49 585
R11 a_156330_n13996.n95 a_156330_n13996.n47 585
R12 a_156330_n13996.n95 a_156330_n13996.n46 585
R13 a_156330_n13996.n95 a_156330_n13996.n45 585
R14 a_156330_n13996.n95 a_156330_n13996.n44 585
R15 a_156330_n13996.n95 a_156330_n13996.n29 291.375
R16 a_156330_n13996.n108 a_156330_n13996.n107 585
R17 a_156330_n13996.n108 a_156330_n13996.n43 585
R18 a_156330_n13996.n108 a_156330_n13996.n42 585
R19 a_156330_n13996.n108 a_156330_n13996.n41 585
R20 a_156330_n13996.n108 a_156330_n13996.n40 585
R21 a_156330_n13996.n108 a_156330_n13996.n39 585
R22 a_156330_n13996.n108 a_156330_n13996.n37 585
R23 a_156330_n13996.n108 a_156330_n13996.n36 585
R24 a_156330_n13996.n108 a_156330_n13996.n35 585
R25 a_156330_n13996.n108 a_156330_n13996.n34 585
R26 a_156330_n13996.n108 a_156330_n13996.n30 291.375
R27 a_156330_n13996.n72 a_156330_n13996.n22 116.999
R28 a_156330_n13996.n72 a_156330_n13996.n65 585
R29 a_156330_n13996.n72 a_156330_n13996.n63 585
R30 a_156330_n13996.n72 a_156330_n13996.n20 116.999
R31 a_156330_n13996.n20 a_156330_n13996.n19 2.92
R32 a_156330_n13996.t44 a_156330_n13996.n2 433.543
R33 a_156330_n13996.t42 a_156330_n13996.n19 433.543
R34 a_156330_n13996.n12 a_156330_n13996.t42 433.351
R35 a_156330_n13996.n1 a_156330_n13996.t30 433.149
R36 a_156330_n13996.t20 a_156330_n13996.n19 433.149
R37 a_156330_n13996.n0 a_156330_n13996.t20 433.149
R38 a_156330_n13996.n19 a_156330_n13996.t26 433.149
R39 a_156330_n13996.t26 a_156330_n13996.n0 433.149
R40 a_156330_n13996.n1 a_156330_n13996.t28 433.149
R41 a_156330_n13996.t28 a_156330_n13996.n4 433.149
R42 a_156330_n13996.t40 a_156330_n13996.n1 433.149
R43 a_156330_n13996.n3 a_156330_n13996.t40 433.149
R44 a_156330_n13996.t4 a_156330_n13996.n1 433.149
R45 a_156330_n13996.n3 a_156330_n13996.t4 433.149
R46 a_156330_n13996.n1 a_156330_n13996.t8 433.149
R47 a_156330_n13996.t8 a_156330_n13996.n3 433.149
R48 a_156330_n13996.n1 a_156330_n13996.t14 433.149
R49 a_156330_n13996.t14 a_156330_n13996.n3 433.149
R50 a_156330_n13996.t34 a_156330_n13996.n0 433.149
R51 a_156330_n13996.n19 a_156330_n13996.t34 433.149
R52 a_156330_n13996.n2 a_156330_n13996.t24 433.149
R53 a_156330_n13996.t24 a_156330_n13996.n5 433.149
R54 a_156330_n13996.t6 a_156330_n13996.n2 433.149
R55 a_156330_n13996.n5 a_156330_n13996.t6 433.149
R56 a_156330_n13996.t10 a_156330_n13996.n2 433.149
R57 a_156330_n13996.n5 a_156330_n13996.t10 433.149
R58 a_156330_n13996.n4 a_156330_n13996.t12 433.149
R59 a_156330_n13996.t12 a_156330_n13996.n5 433.149
R60 a_156330_n13996.n4 a_156330_n13996.t18 433.149
R61 a_156330_n13996.t18 a_156330_n13996.n1 433.149
R62 a_156330_n13996.n5 a_156330_n13996.t32 433.149
R63 a_156330_n13996.t32 a_156330_n13996.n2 433.149
R64 a_156330_n13996.t38 a_156330_n13996.n5 433.149
R65 a_156330_n13996.n2 a_156330_n13996.t38 433.149
R66 a_156330_n13996.n6 a_156330_n13996.t54 433.149
R67 a_156330_n13996.t54 a_156330_n13996.n13 433.149
R68 a_156330_n13996.t49 a_156330_n13996.n6 433.149
R69 a_156330_n13996.n13 a_156330_n13996.t49 433.149
R70 a_156330_n13996.t67 a_156330_n13996.n6 433.149
R71 a_156330_n13996.n14 a_156330_n13996.t67 433.149
R72 a_156330_n13996.n7 a_156330_n13996.t53 433.149
R73 a_156330_n13996.t53 a_156330_n13996.n14 433.149
R74 a_156330_n13996.n7 a_156330_n13996.t62 433.149
R75 a_156330_n13996.t62 a_156330_n13996.n14 433.149
R76 a_156330_n13996.t60 a_156330_n13996.n7 433.149
R77 a_156330_n13996.n14 a_156330_n13996.t60 433.149
R78 a_156330_n13996.t59 a_156330_n13996.n7 433.149
R79 a_156330_n13996.n14 a_156330_n13996.t59 433.149
R80 a_156330_n13996.t56 a_156330_n13996.n14 433.149
R81 a_156330_n13996.n8 a_156330_n13996.t56 433.149
R82 a_156330_n13996.t50 a_156330_n13996.n14 433.149
R83 a_156330_n13996.n8 a_156330_n13996.t50 433.149
R84 a_156330_n13996.t51 a_156330_n13996.n8 433.149
R85 a_156330_n13996.n14 a_156330_n13996.t51 433.149
R86 a_156330_n13996.t66 a_156330_n13996.n8 433.149
R87 a_156330_n13996.n14 a_156330_n13996.t66 433.149
R88 a_156330_n13996.n9 a_156330_n13996.t63 433.149
R89 a_156330_n13996.t63 a_156330_n13996.n11 433.149
R90 a_156330_n13996.n9 a_156330_n13996.t61 433.149
R91 a_156330_n13996.t61 a_156330_n13996.n11 433.149
R92 a_156330_n13996.t58 a_156330_n13996.n9 433.149
R93 a_156330_n13996.n12 a_156330_n13996.t58 433.149
R94 a_156330_n13996.t69 a_156330_n13996.n9 433.149
R95 a_156330_n13996.n12 a_156330_n13996.t69 433.149
R96 a_156330_n13996.n10 a_156330_n13996.t55 433.149
R97 a_156330_n13996.t55 a_156330_n13996.n12 433.149
R98 a_156330_n13996.n10 a_156330_n13996.t52 433.149
R99 a_156330_n13996.t52 a_156330_n13996.n12 433.149
R100 a_156330_n13996.n10 a_156330_n13996.t68 433.149
R101 a_156330_n13996.n12 a_156330_n13996.t68 433.149
R102 a_156330_n13996.t36 a_156330_n13996.n19 433.149
R103 a_156330_n13996.n0 a_156330_n13996.t36 433.149
R104 a_156330_n13996.n6 a_156330_n13996.t57 433.149
R105 a_156330_n13996.t57 a_156330_n13996.n13 433.149
R106 a_156330_n13996.n13 a_156330_n13996.t44 433.149
R107 a_156330_n13996.n2 a_156330_n13996.t16 433.149
R108 a_156330_n13996.n13 a_156330_n13996.t16 433.149
R109 a_156330_n13996.t22 a_156330_n13996.n13 433.149
R110 a_156330_n13996.n2 a_156330_n13996.t22 433.149
R111 a_156330_n13996.n4 a_156330_n13996.t30 433.149
R112 a_156330_n13996.n80 a_156330_n13996.n59 286.238
R113 a_156330_n13996.n95 a_156330_n13996.n48 286.238
R114 a_156330_n13996.n108 a_156330_n13996.n38 286.238
R115 a_156330_n13996.n72 a_156330_n13996.n64 286.238
R116 a_156330_n13996.n66 a_156330_n13996.t65 215.964
R117 a_156330_n13996.n26 a_156330_n13996.t64 215.963
R118 a_156330_n13996.n87 a_156330_n13996.n23 47.0484
R119 a_156330_n13996.n85 a_156330_n13996.n23 47.0484
R120 a_156330_n13996.n84 a_156330_n13996.n23 47.0484
R121 a_156330_n13996.n83 a_156330_n13996.n23 47.0484
R122 a_156330_n13996.n82 a_156330_n13996.n23 47.0484
R123 a_156330_n13996.n81 a_156330_n13996.n23 47.0484
R124 a_156330_n13996.n76 a_156330_n13996.n60 24.8476
R125 a_156330_n13996.n75 a_156330_n13996.n58 24.8476
R126 a_156330_n13996.n91 a_156330_n13996.n49 24.8476
R127 a_156330_n13996.n90 a_156330_n13996.n47 24.8476
R128 a_156330_n13996.n101 a_156330_n13996.n39 24.8476
R129 a_156330_n13996.n100 a_156330_n13996.n37 24.8476
R130 a_156330_n13996.n70 a_156330_n13996.n65 24.8476
R131 a_156330_n13996.n69 a_156330_n13996.n63 24.8476
R132 a_156330_n13996.n77 a_156330_n13996.n61 23.3417
R133 a_156330_n13996.n74 a_156330_n13996.n57 23.3417
R134 a_156330_n13996.n92 a_156330_n13996.n50 23.3417
R135 a_156330_n13996.n89 a_156330_n13996.n46 23.3417
R136 a_156330_n13996.n102 a_156330_n13996.n40 23.3417
R137 a_156330_n13996.n99 a_156330_n13996.n36 23.3417
R138 a_156330_n13996.n68 a_156330_n13996.n20 31.3636
R139 a_156330_n13996.n78 a_156330_n13996.n62 21.8358
R140 a_156330_n13996.n73 a_156330_n13996.n56 21.8358
R141 a_156330_n13996.n93 a_156330_n13996.n51 21.8358
R142 a_156330_n13996.n88 a_156330_n13996.n45 21.8358
R143 a_156330_n13996.n103 a_156330_n13996.n41 21.8358
R144 a_156330_n13996.n98 a_156330_n13996.n35 21.8358
R145 a_156330_n13996.n79 a_156330_n13996.n24 28.1963
R146 a_156330_n13996.n55 a_156330_n13996.n53 20.3299
R147 a_156330_n13996.n94 a_156330_n13996.n25 28.1963
R148 a_156330_n13996.n52 a_156330_n13996.n44 20.3299
R149 a_156330_n13996.n104 a_156330_n13996.n42 20.3299
R150 a_156330_n13996.n97 a_156330_n13996.n34 20.3299
R151 a_156330_n13996.n107 a_156330_n13996.n13 19.0887
R152 a_156330_n13996.n54 a_156330_n13996.n28 24.6333
R153 a_156330_n13996.n86 a_156330_n13996.n29 24.6333
R154 a_156330_n13996.n105 a_156330_n13996.n43 18.824
R155 a_156330_n13996.n96 a_156330_n13996.n30 24.6333
R156 a_156330_n13996.n80 a_156330_n13996.n24 194.291
R157 a_156330_n13996.n28 a_156330_n13996.n19 9.76605
R158 a_156330_n13996.n95 a_156330_n13996.n25 194.291
R159 a_156330_n13996.n2 a_156330_n13996.n29 9.76605
R160 a_156330_n13996.n107 a_156330_n13996.n106 17.3181
R161 a_156330_n13996.n30 a_156330_n13996.n2 9.76605
R162 a_156330_n13996.n22 a_156330_n13996.n0 2.92
R163 a_156330_n13996.n76 a_156330_n13996.n59 13.2799
R164 a_156330_n13996.n75 a_156330_n13996.n59 13.2799
R165 a_156330_n13996.n91 a_156330_n13996.n48 13.2799
R166 a_156330_n13996.n90 a_156330_n13996.n48 13.2799
R167 a_156330_n13996.n101 a_156330_n13996.n38 13.2799
R168 a_156330_n13996.n100 a_156330_n13996.n38 13.2799
R169 a_156330_n13996.n70 a_156330_n13996.n64 13.2799
R170 a_156330_n13996.n69 a_156330_n13996.n64 13.2799
R171 a_156330_n13996.n21 a_156330_n13996.n70 9.3005
R172 a_156330_n13996.n21 a_156330_n13996.n71 9.3005
R173 a_156330_n13996.n21 a_156330_n13996.n69 9.3005
R174 a_156330_n13996.n21 a_156330_n13996.n68 9.3005
R175 a_156330_n13996.n15 a_156330_n13996.n97 9.3005
R176 a_156330_n13996.n15 a_156330_n13996.n96 9.3005
R177 a_156330_n13996.n15 a_156330_n13996.n98 9.3005
R178 a_156330_n13996.n16 a_156330_n13996.n101 9.3005
R179 a_156330_n13996.n16 a_156330_n13996.n102 9.3005
R180 a_156330_n13996.n16 a_156330_n13996.n103 9.3005
R181 a_156330_n13996.n16 a_156330_n13996.n104 9.3005
R182 a_156330_n13996.n16 a_156330_n13996.n105 9.3005
R183 a_156330_n13996.n106 a_156330_n13996.n16 9.3005
R184 a_156330_n13996.n16 a_156330_n13996.n100 9.3005
R185 a_156330_n13996.n16 a_156330_n13996.n99 9.3005
R186 a_156330_n13996.n17 a_156330_n13996.n91 9.3005
R187 a_156330_n13996.n17 a_156330_n13996.n92 9.3005
R188 a_156330_n13996.n17 a_156330_n13996.n93 9.3005
R189 a_156330_n13996.n17 a_156330_n13996.n94 9.3005
R190 a_156330_n13996.n25 a_156330_n13996.n5 6.07169
R191 a_156330_n13996.n17 a_156330_n13996.n90 9.3005
R192 a_156330_n13996.n17 a_156330_n13996.n89 9.3005
R193 a_156330_n13996.n17 a_156330_n13996.n88 9.3005
R194 a_156330_n13996.n17 a_156330_n13996.n52 9.3005
R195 a_156330_n13996.n17 a_156330_n13996.n86 9.3005
R196 a_156330_n13996.n18 a_156330_n13996.n76 9.3005
R197 a_156330_n13996.n18 a_156330_n13996.n77 9.3005
R198 a_156330_n13996.n18 a_156330_n13996.n78 9.3005
R199 a_156330_n13996.n18 a_156330_n13996.n79 9.3005
R200 a_156330_n13996.n0 a_156330_n13996.n24 6.07169
R201 a_156330_n13996.n18 a_156330_n13996.n75 9.3005
R202 a_156330_n13996.n18 a_156330_n13996.n74 9.3005
R203 a_156330_n13996.n18 a_156330_n13996.n73 9.3005
R204 a_156330_n13996.n55 a_156330_n13996.n18 9.3005
R205 a_156330_n13996.n18 a_156330_n13996.n54 9.3005
R206 a_156330_n13996.n106 a_156330_n13996.n43 8.28285
R207 a_156330_n13996.n17 a_156330_n13996.n23 3.89414
R208 a_156330_n13996.n23 a_156330_n13996.n18 3.89414
R209 a_156330_n13996.n27 a_156330_n13996.n33 18.4327
R210 a_156330_n13996.n27 a_156330_n13996.n67 18.4327
R211 a_156330_n13996.n27 a_156330_n13996.n109 18.433
R212 a_156330_n13996.n54 a_156330_n13996.n53 6.77697
R213 a_156330_n13996.n86 a_156330_n13996.n44 6.77697
R214 a_156330_n13996.n105 a_156330_n13996.n42 6.77697
R215 a_156330_n13996.n96 a_156330_n13996.n34 6.77697
R216 a_156330_n13996.n80 a_156330_n13996.t21 5.7135
R217 a_156330_n13996.n80 a_156330_n13996.t35 5.7135
R218 a_156330_n13996.n95 a_156330_n13996.t25 5.7135
R219 a_156330_n13996.n95 a_156330_n13996.t39 5.7135
R220 a_156330_n13996.n87 a_156330_n13996.t17 5.7135
R221 a_156330_n13996.n87 a_156330_n13996.t45 5.7135
R222 a_156330_n13996.n85 a_156330_n13996.t11 5.7135
R223 a_156330_n13996.n85 a_156330_n13996.t7 5.7135
R224 a_156330_n13996.n84 a_156330_n13996.t19 5.7135
R225 a_156330_n13996.n84 a_156330_n13996.t13 5.7135
R226 a_156330_n13996.n83 a_156330_n13996.t29 5.7135
R227 a_156330_n13996.n83 a_156330_n13996.t31 5.7135
R228 a_156330_n13996.n82 a_156330_n13996.t5 5.7135
R229 a_156330_n13996.n82 a_156330_n13996.t41 5.7135
R230 a_156330_n13996.n81 a_156330_n13996.t15 5.7135
R231 a_156330_n13996.n81 a_156330_n13996.t9 5.7135
R232 a_156330_n13996.n108 a_156330_n13996.t33 5.7135
R233 a_156330_n13996.n108 a_156330_n13996.t23 5.7135
R234 a_156330_n13996.n72 a_156330_n13996.t37 5.7135
R235 a_156330_n13996.n72 a_156330_n13996.t27 5.7135
R236 a_156330_n13996.n27 a_156330_n13996.t3 94.44
R237 a_156330_n13996.n79 a_156330_n13996.n62 5.27109
R238 a_156330_n13996.n56 a_156330_n13996.n55 5.27109
R239 a_156330_n13996.n94 a_156330_n13996.n51 5.27109
R240 a_156330_n13996.n52 a_156330_n13996.n45 5.27109
R241 a_156330_n13996.n104 a_156330_n13996.n41 5.27109
R242 a_156330_n13996.n97 a_156330_n13996.n35 5.27109
R243 a_156330_n13996.n27 a_156330_n13996.n31 4.69006
R244 a_156330_n13996.n15 a_156330_n13996.n31 2.21422
R245 a_156330_n13996.n19 a_156330_n13996.n32 2.21422
R246 a_156330_n13996.n32 a_156330_n13996.n27 4.5738
R247 a_156330_n13996.n23 a_156330_n13996.t43 198.911
R248 a_156330_n13996.n78 a_156330_n13996.n61 3.76521
R249 a_156330_n13996.n73 a_156330_n13996.n57 3.76521
R250 a_156330_n13996.n93 a_156330_n13996.n50 3.76521
R251 a_156330_n13996.n88 a_156330_n13996.n46 3.76521
R252 a_156330_n13996.n103 a_156330_n13996.n40 3.76521
R253 a_156330_n13996.n98 a_156330_n13996.n36 3.76521
R254 a_156330_n13996.n22 a_156330_n13996.n71 31.3636
R255 a_156330_n13996.n33 a_156330_n13996.t1 3.4805
R256 a_156330_n13996.n33 a_156330_n13996.t2 3.4805
R257 a_156330_n13996.n67 a_156330_n13996.t46 3.4805
R258 a_156330_n13996.n67 a_156330_n13996.t48 3.4805
R259 a_156330_n13996.n109 a_156330_n13996.t47 3.4805
R260 a_156330_n13996.t0 a_156330_n13996.n109 3.4805
R261 a_156330_n13996.n7 a_156330_n13996.n6 2.3705
R262 a_156330_n13996.n77 a_156330_n13996.n60 2.25932
R263 a_156330_n13996.n74 a_156330_n13996.n58 2.25932
R264 a_156330_n13996.n92 a_156330_n13996.n49 2.25932
R265 a_156330_n13996.n89 a_156330_n13996.n47 2.25932
R266 a_156330_n13996.n102 a_156330_n13996.n39 2.25932
R267 a_156330_n13996.n99 a_156330_n13996.n37 2.25932
R268 a_156330_n13996.n71 a_156330_n13996.n65 2.25932
R269 a_156330_n13996.n68 a_156330_n13996.n63 2.25932
R270 a_156330_n13996.n23 a_156330_n13996.n31 2.2506
R271 a_156330_n13996.n32 a_156330_n13996.n23 1.75553
R272 a_156330_n13996.n15 a_156330_n13996.n2 1.75199
R273 a_156330_n13996.n0 a_156330_n13996.n18 1.64967
R274 a_156330_n13996.n5 a_156330_n13996.n17 1.64967
R275 a_156330_n13996.n13 a_156330_n13996.n5 1.63467
R276 a_156330_n13996.n6 a_156330_n13996.n26 1.62034
R277 a_156330_n13996.n66 a_156330_n13996.n10 1.61786
R278 a_156330_n13996.n14 a_156330_n13996.n1 1.60531
R279 a_156330_n13996.n11 a_156330_n13996.n14 1.5805
R280 a_156330_n13996.n14 a_156330_n13996.n13 1.5805
R281 a_156330_n13996.n12 a_156330_n13996.n11 1.5805
R282 a_156330_n13996.n10 a_156330_n13996.n9 1.5805
R283 a_156330_n13996.n9 a_156330_n13996.n8 1.5805
R284 a_156330_n13996.n8 a_156330_n13996.n7 1.5805
R285 a_156330_n13996.n4 a_156330_n13996.n3 1.5805
R286 a_156330_n13996.n4 a_156330_n13996.n2 1.5805
R287 a_156330_n13996.n1 a_156330_n13996.n0 1.53258
R288 a_156330_n13996.n16 a_156330_n13996.n15 1.42603
R289 a_156330_n13996.n21 a_156330_n13996.n19 1.39252
R290 a_156330_n13996.n13 a_156330_n13996.n26 1.22534
R291 a_156330_n13996.n12 a_156330_n13996.n66 1.22286
R292 a_156330_n13996.n3 a_156330_n13996.n19 1.1855
R293 a_156330_n13996.n5 a_156330_n13996.n1 1.1855
R294 a_156330_n13996.n0 a_156330_n13996.n21 1.1005
R295 a_156330_n13996.n17 a_156330_n13996.n2 1.09535
R296 a_156330_n13996.n18 a_156330_n13996.n19 1.09535
R297 a_156330_n13996.n0 a_156330_n13996.n12 1.01624
R298 a_156330_n13996.n16 a_156330_n13996.n13 1.00124
R299 a_153429_n11365.n141 a_153429_n11365.n140 815.966
R300 a_153429_n11365.n280 a_153429_n11365.n274 585
R301 a_153429_n11365.n280 a_153429_n11365.n273 585
R302 a_153429_n11365.n281 a_153429_n11365.n280 585
R303 a_153429_n11365.n266 a_153429_n11365.n260 585
R304 a_153429_n11365.n266 a_153429_n11365.n259 585
R305 a_153429_n11365.n267 a_153429_n11365.n266 585
R306 a_153429_n11365.n252 a_153429_n11365.n246 585
R307 a_153429_n11365.n252 a_153429_n11365.n245 585
R308 a_153429_n11365.n253 a_153429_n11365.n252 585
R309 a_153429_n11365.n238 a_153429_n11365.n232 585
R310 a_153429_n11365.n238 a_153429_n11365.n231 585
R311 a_153429_n11365.n239 a_153429_n11365.n238 585
R312 a_153429_n11365.n224 a_153429_n11365.n218 585
R313 a_153429_n11365.n224 a_153429_n11365.n217 585
R314 a_153429_n11365.n225 a_153429_n11365.n224 585
R315 a_153429_n11365.n210 a_153429_n11365.n204 585
R316 a_153429_n11365.n210 a_153429_n11365.n203 585
R317 a_153429_n11365.n211 a_153429_n11365.n210 585
R318 a_153429_n11365.n196 a_153429_n11365.n190 585
R319 a_153429_n11365.n196 a_153429_n11365.n189 585
R320 a_153429_n11365.n197 a_153429_n11365.n196 585
R321 a_153429_n11365.n182 a_153429_n11365.n176 585
R322 a_153429_n11365.n182 a_153429_n11365.n175 585
R323 a_153429_n11365.n183 a_153429_n11365.n182 585
R324 a_153429_n11365.n168 a_153429_n11365.n162 585
R325 a_153429_n11365.n168 a_153429_n11365.n161 585
R326 a_153429_n11365.n169 a_153429_n11365.n168 585
R327 a_153429_n11365.n154 a_153429_n11365.n148 585
R328 a_153429_n11365.n154 a_153429_n11365.n147 585
R329 a_153429_n11365.n155 a_153429_n11365.n154 585
R330 a_153429_n11365.n125 a_153429_n11365.n124 585
R331 a_153429_n11365.n122 a_153429_n11365.n121 585
R332 a_153429_n11365.n132 a_153429_n11365.n131 585
R333 a_153429_n11365.n134 a_153429_n11365.n133 585
R334 a_153429_n11365.n119 a_153429_n11365.n118 585
R335 a_153429_n11365.n140 a_153429_n11365.n139 585
R336 a_153429_n11365.n24 a_153429_n11365.t54 433.149
R337 a_153429_n11365.t54 a_153429_n11365.n23 433.149
R338 a_153429_n11365.n25 a_153429_n11365.t33 433.149
R339 a_153429_n11365.t33 a_153429_n11365.n20 433.149
R340 a_153429_n11365.t45 a_153429_n11365.n26 433.149
R341 a_153429_n11365.n27 a_153429_n11365.t45 433.149
R342 a_153429_n11365.t35 a_153429_n11365.n19 433.149
R343 a_153429_n11365.n28 a_153429_n11365.t35 433.149
R344 a_153429_n11365.n30 a_153429_n11365.t32 433.149
R345 a_153429_n11365.t32 a_153429_n11365.n29 433.149
R346 a_153429_n11365.n31 a_153429_n11365.t68 433.149
R347 a_153429_n11365.t68 a_153429_n11365.n18 433.149
R348 a_153429_n11365.t49 a_153429_n11365.n32 433.149
R349 a_153429_n11365.n33 a_153429_n11365.t49 433.149
R350 a_153429_n11365.t40 a_153429_n11365.n17 433.149
R351 a_153429_n11365.n286 a_153429_n11365.t40 433.149
R352 a_153429_n11365.n288 a_153429_n11365.t59 433.149
R353 a_153429_n11365.t59 a_153429_n11365.n287 433.149
R354 a_153429_n11365.n289 a_153429_n11365.t48 433.149
R355 a_153429_n11365.t48 a_153429_n11365.n16 433.149
R356 a_153429_n11365.t38 a_153429_n11365.n290 433.149
R357 a_153429_n11365.n291 a_153429_n11365.t38 433.149
R358 a_153429_n11365.t66 a_153429_n11365.n15 433.149
R359 a_153429_n11365.n292 a_153429_n11365.t66 433.149
R360 a_153429_n11365.n294 a_153429_n11365.t58 433.149
R361 a_153429_n11365.t58 a_153429_n11365.n293 433.149
R362 a_153429_n11365.n295 a_153429_n11365.t52 433.149
R363 a_153429_n11365.t52 a_153429_n11365.n14 433.149
R364 a_153429_n11365.t65 a_153429_n11365.n296 433.149
R365 a_153429_n11365.n297 a_153429_n11365.t65 433.149
R366 a_153429_n11365.t55 a_153429_n11365.n13 433.149
R367 a_153429_n11365.n298 a_153429_n11365.t55 433.149
R368 a_153429_n11365.n300 a_153429_n11365.t34 433.149
R369 a_153429_n11365.t34 a_153429_n11365.n299 433.149
R370 a_153429_n11365.n301 a_153429_n11365.t70 433.149
R371 a_153429_n11365.t70 a_153429_n11365.n12 433.149
R372 a_153429_n11365.t67 a_153429_n11365.n302 433.149
R373 a_153429_n11365.n303 a_153429_n11365.t67 433.149
R374 a_153429_n11365.t62 a_153429_n11365.n11 433.149
R375 a_153429_n11365.n304 a_153429_n11365.t62 433.149
R376 a_153429_n11365.n306 a_153429_n11365.t57 433.149
R377 a_153429_n11365.t57 a_153429_n11365.n305 433.149
R378 a_153429_n11365.n307 a_153429_n11365.t51 433.149
R379 a_153429_n11365.t51 a_153429_n11365.n10 433.149
R380 a_153429_n11365.t42 a_153429_n11365.n308 433.149
R381 a_153429_n11365.n309 a_153429_n11365.t42 433.149
R382 a_153429_n11365.t37 a_153429_n11365.n9 433.149
R383 a_153429_n11365.n310 a_153429_n11365.t37 433.149
R384 a_153429_n11365.n312 a_153429_n11365.t71 433.149
R385 a_153429_n11365.t71 a_153429_n11365.n311 433.149
R386 a_153429_n11365.n313 a_153429_n11365.t69 433.149
R387 a_153429_n11365.t69 a_153429_n11365.n8 433.149
R388 a_153429_n11365.t47 a_153429_n11365.n314 433.149
R389 a_153429_n11365.n315 a_153429_n11365.t47 433.149
R390 a_153429_n11365.t64 a_153429_n11365.n7 433.149
R391 a_153429_n11365.n316 a_153429_n11365.t64 433.149
R392 a_153429_n11365.n318 a_153429_n11365.t53 433.149
R393 a_153429_n11365.t53 a_153429_n11365.n317 433.149
R394 a_153429_n11365.n319 a_153429_n11365.t44 433.149
R395 a_153429_n11365.t44 a_153429_n11365.n6 433.149
R396 a_153429_n11365.t39 a_153429_n11365.n320 433.149
R397 a_153429_n11365.n321 a_153429_n11365.t39 433.149
R398 a_153429_n11365.t63 a_153429_n11365.n4 433.149
R399 a_153429_n11365.n322 a_153429_n11365.t63 433.149
R400 a_153429_n11365.n324 a_153429_n11365.t60 433.149
R401 a_153429_n11365.t60 a_153429_n11365.n323 433.149
R402 a_153429_n11365.n325 a_153429_n11365.t50 433.149
R403 a_153429_n11365.t50 a_153429_n11365.n3 433.149
R404 a_153429_n11365.t41 a_153429_n11365.n326 433.149
R405 a_153429_n11365.n327 a_153429_n11365.t41 433.149
R406 a_153429_n11365.t36 a_153429_n11365.n2 433.149
R407 a_153429_n11365.n328 a_153429_n11365.t36 433.149
R408 a_153429_n11365.n330 a_153429_n11365.t61 433.149
R409 a_153429_n11365.t61 a_153429_n11365.n329 433.149
R410 a_153429_n11365.n331 a_153429_n11365.t56 433.149
R411 a_153429_n11365.t56 a_153429_n11365.n1 433.149
R412 a_153429_n11365.t46 a_153429_n11365.n332 433.149
R413 a_153429_n11365.n333 a_153429_n11365.t46 433.149
R414 a_153429_n11365.t43 a_153429_n11365.n0 433.149
R415 a_153429_n11365.n334 a_153429_n11365.t43 433.149
R416 a_153429_n11365.t10 a_153429_n11365.n123 384.339
R417 a_153429_n11365.n44 a_153429_n11365.n43 325.69
R418 a_153429_n11365.n124 a_153429_n11365.n121 230.966
R419 a_153429_n11365.n132 a_153429_n11365.n121 230.966
R420 a_153429_n11365.n133 a_153429_n11365.n132 230.966
R421 a_153429_n11365.n133 a_153429_n11365.n118 230.966
R422 a_153429_n11365.n140 a_153429_n11365.n118 230.966
R423 a_153429_n11365.n45 a_153429_n11365.n44 185
R424 a_153429_n11365.n40 a_153429_n11365.n39 185
R425 a_153429_n11365.n52 a_153429_n11365.n51 185
R426 a_153429_n11365.n53 a_153429_n11365.n37 185
R427 a_153429_n11365.n58 a_153429_n11365.n57 185
R428 a_153429_n11365.n56 a_153429_n11365.n55 185
R429 a_153429_n11365.n70 a_153429_n11365.n67 185
R430 a_153429_n11365.n72 a_153429_n11365.n67 185
R431 a_153429_n11365.n68 a_153429_n11365.n67 185
R432 a_153429_n11365.n77 a_153429_n11365.n67 185
R433 a_153429_n11365.n86 a_153429_n11365.n83 185
R434 a_153429_n11365.n88 a_153429_n11365.n83 185
R435 a_153429_n11365.n84 a_153429_n11365.n83 185
R436 a_153429_n11365.n93 a_153429_n11365.n83 185
R437 a_153429_n11365.n102 a_153429_n11365.n99 185
R438 a_153429_n11365.n104 a_153429_n11365.n99 185
R439 a_153429_n11365.n100 a_153429_n11365.n99 185
R440 a_153429_n11365.n109 a_153429_n11365.n99 185
R441 a_153429_n11365.n54 a_153429_n11365.t4 174.857
R442 a_153429_n11365.n44 a_153429_n11365.n39 140.69
R443 a_153429_n11365.n52 a_153429_n11365.n39 140.69
R444 a_153429_n11365.n53 a_153429_n11365.n52 140.69
R445 a_153429_n11365.n57 a_153429_n11365.n53 140.69
R446 a_153429_n11365.n57 a_153429_n11365.n56 140.69
R447 a_153429_n11365.n124 a_153429_n11365.t10 115.484
R448 a_153429_n11365.n56 a_153429_n11365.t4 70.3453
R449 a_153429_n11365.n280 a_153429_n11365.n279 51.6891
R450 a_153429_n11365.n266 a_153429_n11365.n265 51.6891
R451 a_153429_n11365.n252 a_153429_n11365.n251 51.6891
R452 a_153429_n11365.n238 a_153429_n11365.n237 51.6891
R453 a_153429_n11365.n224 a_153429_n11365.n223 51.6891
R454 a_153429_n11365.n210 a_153429_n11365.n209 51.6891
R455 a_153429_n11365.n196 a_153429_n11365.n195 51.6891
R456 a_153429_n11365.n182 a_153429_n11365.n181 51.6891
R457 a_153429_n11365.n168 a_153429_n11365.n167 51.6891
R458 a_153429_n11365.n154 a_153429_n11365.n153 51.6891
R459 a_153429_n11365.n279 a_153429_n11365.n278 29.8062
R460 a_153429_n11365.n265 a_153429_n11365.n264 29.8062
R461 a_153429_n11365.n251 a_153429_n11365.n250 29.8062
R462 a_153429_n11365.n237 a_153429_n11365.n236 29.8062
R463 a_153429_n11365.n223 a_153429_n11365.n222 29.8062
R464 a_153429_n11365.n209 a_153429_n11365.n208 29.8062
R465 a_153429_n11365.n195 a_153429_n11365.n194 29.8062
R466 a_153429_n11365.n181 a_153429_n11365.n180 29.8062
R467 a_153429_n11365.n167 a_153429_n11365.n166 29.8062
R468 a_153429_n11365.n153 a_153429_n11365.n152 29.8062
R469 a_153429_n11365.n125 a_153429_n11365.n123 29.3167
R470 a_153429_n11365.n55 a_153429_n11365.n54 28.4333
R471 a_153429_n11365.n79 a_153429_n11365.n78 26.8428
R472 a_153429_n11365.n95 a_153429_n11365.n94 26.8428
R473 a_153429_n11365.n111 a_153429_n11365.n110 26.8428
R474 a_153429_n11365.n126 a_153429_n11365.n122 24.8476
R475 a_153429_n11365.n58 a_153429_n11365.n38 24.8476
R476 a_153429_n11365.n131 a_153429_n11365.n130 23.3417
R477 a_153429_n11365.n59 a_153429_n11365.n37 23.3417
R478 a_153429_n11365.n134 a_153429_n11365.n120 21.8358
R479 a_153429_n11365.n51 a_153429_n11365.n50 21.8358
R480 a_153429_n11365.n78 a_153429_n11365.n77 21.8358
R481 a_153429_n11365.n94 a_153429_n11365.n93 21.8358
R482 a_153429_n11365.n110 a_153429_n11365.n109 21.8358
R483 a_153429_n11365.n278 a_153429_n11365.n274 20.3299
R484 a_153429_n11365.n264 a_153429_n11365.n260 20.3299
R485 a_153429_n11365.n250 a_153429_n11365.n246 20.3299
R486 a_153429_n11365.n236 a_153429_n11365.n232 20.3299
R487 a_153429_n11365.n222 a_153429_n11365.n218 20.3299
R488 a_153429_n11365.n208 a_153429_n11365.n204 20.3299
R489 a_153429_n11365.n194 a_153429_n11365.n190 20.3299
R490 a_153429_n11365.n180 a_153429_n11365.n176 20.3299
R491 a_153429_n11365.n166 a_153429_n11365.n162 20.3299
R492 a_153429_n11365.n152 a_153429_n11365.n148 20.3299
R493 a_153429_n11365.n135 a_153429_n11365.n119 20.3299
R494 a_153429_n11365.n49 a_153429_n11365.n40 20.3299
R495 a_153429_n11365.n76 a_153429_n11365.n68 20.3299
R496 a_153429_n11365.n92 a_153429_n11365.n84 20.3299
R497 a_153429_n11365.n108 a_153429_n11365.n100 20.3299
R498 a_153429_n11365.n282 a_153429_n11365.n281 19.1618
R499 a_153429_n11365.n268 a_153429_n11365.n267 19.1618
R500 a_153429_n11365.n254 a_153429_n11365.n253 19.1618
R501 a_153429_n11365.n240 a_153429_n11365.n239 19.1618
R502 a_153429_n11365.n226 a_153429_n11365.n225 19.1618
R503 a_153429_n11365.n212 a_153429_n11365.n211 19.1618
R504 a_153429_n11365.n198 a_153429_n11365.n197 19.1618
R505 a_153429_n11365.n184 a_153429_n11365.n183 19.1618
R506 a_153429_n11365.n170 a_153429_n11365.n169 19.1618
R507 a_153429_n11365.n156 a_153429_n11365.n155 19.1618
R508 a_153429_n11365.n142 a_153429_n11365.n141 19.1618
R509 a_153429_n11365.n43 a_153429_n11365.n34 19.1618
R510 a_153429_n11365.n70 a_153429_n11365.n65 19.1618
R511 a_153429_n11365.n86 a_153429_n11365.n64 19.1618
R512 a_153429_n11365.n102 a_153429_n11365.n63 19.1618
R513 a_153429_n11365.n275 a_153429_n11365.n273 18.824
R514 a_153429_n11365.n261 a_153429_n11365.n259 18.824
R515 a_153429_n11365.n247 a_153429_n11365.n245 18.824
R516 a_153429_n11365.n233 a_153429_n11365.n231 18.824
R517 a_153429_n11365.n219 a_153429_n11365.n217 18.824
R518 a_153429_n11365.n205 a_153429_n11365.n203 18.824
R519 a_153429_n11365.n191 a_153429_n11365.n189 18.824
R520 a_153429_n11365.n177 a_153429_n11365.n175 18.824
R521 a_153429_n11365.n163 a_153429_n11365.n161 18.824
R522 a_153429_n11365.n149 a_153429_n11365.n147 18.824
R523 a_153429_n11365.n139 a_153429_n11365.n138 18.824
R524 a_153429_n11365.n46 a_153429_n11365.n45 18.824
R525 a_153429_n11365.n73 a_153429_n11365.n72 18.824
R526 a_153429_n11365.n89 a_153429_n11365.n88 18.824
R527 a_153429_n11365.n105 a_153429_n11365.n104 18.824
R528 a_153429_n11365.n281 a_153429_n11365.n272 17.3181
R529 a_153429_n11365.n267 a_153429_n11365.n258 17.3181
R530 a_153429_n11365.n253 a_153429_n11365.n244 17.3181
R531 a_153429_n11365.n239 a_153429_n11365.n230 17.3181
R532 a_153429_n11365.n225 a_153429_n11365.n216 17.3181
R533 a_153429_n11365.n211 a_153429_n11365.n202 17.3181
R534 a_153429_n11365.n197 a_153429_n11365.n188 17.3181
R535 a_153429_n11365.n183 a_153429_n11365.n174 17.3181
R536 a_153429_n11365.n169 a_153429_n11365.n160 17.3181
R537 a_153429_n11365.n155 a_153429_n11365.n146 17.3181
R538 a_153429_n11365.n141 a_153429_n11365.n117 17.3181
R539 a_153429_n11365.n43 a_153429_n11365.n42 17.3181
R540 a_153429_n11365.n71 a_153429_n11365.n70 17.3181
R541 a_153429_n11365.n87 a_153429_n11365.n86 17.3181
R542 a_153429_n11365.n103 a_153429_n11365.n102 17.3181
R543 a_153429_n11365.n79 a_153429_n11365.n67 16.7801
R544 a_153429_n11365.n95 a_153429_n11365.n83 16.7801
R545 a_153429_n11365.n111 a_153429_n11365.n99 16.7801
R546 a_153429_n11365.n272 a_153429_n11365.n271 9.3005
R547 a_153429_n11365.n278 a_153429_n11365.n277 9.3005
R548 a_153429_n11365.n276 a_153429_n11365.n275 9.3005
R549 a_153429_n11365.n258 a_153429_n11365.n257 9.3005
R550 a_153429_n11365.n264 a_153429_n11365.n263 9.3005
R551 a_153429_n11365.n262 a_153429_n11365.n261 9.3005
R552 a_153429_n11365.n244 a_153429_n11365.n243 9.3005
R553 a_153429_n11365.n250 a_153429_n11365.n249 9.3005
R554 a_153429_n11365.n248 a_153429_n11365.n247 9.3005
R555 a_153429_n11365.n230 a_153429_n11365.n229 9.3005
R556 a_153429_n11365.n236 a_153429_n11365.n235 9.3005
R557 a_153429_n11365.n234 a_153429_n11365.n233 9.3005
R558 a_153429_n11365.n216 a_153429_n11365.n215 9.3005
R559 a_153429_n11365.n222 a_153429_n11365.n221 9.3005
R560 a_153429_n11365.n220 a_153429_n11365.n219 9.3005
R561 a_153429_n11365.n202 a_153429_n11365.n201 9.3005
R562 a_153429_n11365.n208 a_153429_n11365.n207 9.3005
R563 a_153429_n11365.n206 a_153429_n11365.n205 9.3005
R564 a_153429_n11365.n188 a_153429_n11365.n187 9.3005
R565 a_153429_n11365.n194 a_153429_n11365.n193 9.3005
R566 a_153429_n11365.n192 a_153429_n11365.n191 9.3005
R567 a_153429_n11365.n174 a_153429_n11365.n173 9.3005
R568 a_153429_n11365.n180 a_153429_n11365.n179 9.3005
R569 a_153429_n11365.n178 a_153429_n11365.n177 9.3005
R570 a_153429_n11365.n160 a_153429_n11365.n159 9.3005
R571 a_153429_n11365.n166 a_153429_n11365.n165 9.3005
R572 a_153429_n11365.n164 a_153429_n11365.n163 9.3005
R573 a_153429_n11365.n146 a_153429_n11365.n145 9.3005
R574 a_153429_n11365.n152 a_153429_n11365.n151 9.3005
R575 a_153429_n11365.n150 a_153429_n11365.n149 9.3005
R576 a_153429_n11365.n127 a_153429_n11365.n126 9.3005
R577 a_153429_n11365.n130 a_153429_n11365.n129 9.3005
R578 a_153429_n11365.n117 a_153429_n11365.n116 9.3005
R579 a_153429_n11365.n136 a_153429_n11365.n135 9.3005
R580 a_153429_n11365.n138 a_153429_n11365.n137 9.3005
R581 a_153429_n11365.n128 a_153429_n11365.n120 9.3005
R582 a_153429_n11365.n38 a_153429_n11365.n36 9.3005
R583 a_153429_n11365.n60 a_153429_n11365.n59 9.3005
R584 a_153429_n11365.n50 a_153429_n11365.n35 9.3005
R585 a_153429_n11365.n49 a_153429_n11365.n48 9.3005
R586 a_153429_n11365.n47 a_153429_n11365.n46 9.3005
R587 a_153429_n11365.n42 a_153429_n11365.n41 9.3005
R588 a_153429_n11365.n78 a_153429_n11365.n66 9.3005
R589 a_153429_n11365.n76 a_153429_n11365.n75 9.3005
R590 a_153429_n11365.n74 a_153429_n11365.n73 9.3005
R591 a_153429_n11365.n71 a_153429_n11365.n69 9.3005
R592 a_153429_n11365.n94 a_153429_n11365.n82 9.3005
R593 a_153429_n11365.n92 a_153429_n11365.n91 9.3005
R594 a_153429_n11365.n90 a_153429_n11365.n89 9.3005
R595 a_153429_n11365.n87 a_153429_n11365.n85 9.3005
R596 a_153429_n11365.n110 a_153429_n11365.n98 9.3005
R597 a_153429_n11365.n108 a_153429_n11365.n107 9.3005
R598 a_153429_n11365.n106 a_153429_n11365.n105 9.3005
R599 a_153429_n11365.n103 a_153429_n11365.n101 9.3005
R600 a_153429_n11365.n273 a_153429_n11365.n272 8.28285
R601 a_153429_n11365.n259 a_153429_n11365.n258 8.28285
R602 a_153429_n11365.n245 a_153429_n11365.n244 8.28285
R603 a_153429_n11365.n231 a_153429_n11365.n230 8.28285
R604 a_153429_n11365.n217 a_153429_n11365.n216 8.28285
R605 a_153429_n11365.n203 a_153429_n11365.n202 8.28285
R606 a_153429_n11365.n189 a_153429_n11365.n188 8.28285
R607 a_153429_n11365.n175 a_153429_n11365.n174 8.28285
R608 a_153429_n11365.n161 a_153429_n11365.n160 8.28285
R609 a_153429_n11365.n147 a_153429_n11365.n146 8.28285
R610 a_153429_n11365.n139 a_153429_n11365.n117 8.28285
R611 a_153429_n11365.n45 a_153429_n11365.n42 8.28285
R612 a_153429_n11365.n72 a_153429_n11365.n71 8.28285
R613 a_153429_n11365.n88 a_153429_n11365.n87 8.28285
R614 a_153429_n11365.n104 a_153429_n11365.n103 8.28285
R615 a_153429_n11365.n283 a_153429_n11365.n270 7.9105
R616 a_153429_n11365.n269 a_153429_n11365.n256 7.9105
R617 a_153429_n11365.n255 a_153429_n11365.n242 7.9105
R618 a_153429_n11365.n241 a_153429_n11365.n228 7.9105
R619 a_153429_n11365.n227 a_153429_n11365.n214 7.9105
R620 a_153429_n11365.n213 a_153429_n11365.n200 7.9105
R621 a_153429_n11365.n199 a_153429_n11365.n186 7.9105
R622 a_153429_n11365.n185 a_153429_n11365.n172 7.9105
R623 a_153429_n11365.n171 a_153429_n11365.n158 7.9105
R624 a_153429_n11365.n157 a_153429_n11365.n144 7.9105
R625 a_153429_n11365.n143 a_153429_n11365.n115 7.9105
R626 a_153429_n11365.n62 a_153429_n11365.n34 7.9105
R627 a_153429_n11365.n81 a_153429_n11365.n65 7.9105
R628 a_153429_n11365.n97 a_153429_n11365.n64 7.9105
R629 a_153429_n11365.n113 a_153429_n11365.n63 7.9105
R630 a_153429_n11365.n113 a_153429_n11365.n112 7.9105
R631 a_153429_n11365.n97 a_153429_n11365.n96 7.9105
R632 a_153429_n11365.n81 a_153429_n11365.n80 7.9105
R633 a_153429_n11365.n62 a_153429_n11365.n61 7.9105
R634 a_153429_n11365.n143 a_153429_n11365.n142 7.9105
R635 a_153429_n11365.n157 a_153429_n11365.n156 7.9105
R636 a_153429_n11365.n171 a_153429_n11365.n170 7.9105
R637 a_153429_n11365.n185 a_153429_n11365.n184 7.9105
R638 a_153429_n11365.n199 a_153429_n11365.n198 7.9105
R639 a_153429_n11365.n213 a_153429_n11365.n212 7.9105
R640 a_153429_n11365.n227 a_153429_n11365.n226 7.9105
R641 a_153429_n11365.n241 a_153429_n11365.n240 7.9105
R642 a_153429_n11365.n255 a_153429_n11365.n254 7.9105
R643 a_153429_n11365.n269 a_153429_n11365.n268 7.9105
R644 a_153429_n11365.n283 a_153429_n11365.n282 7.9105
R645 a_153429_n11365.n275 a_153429_n11365.n274 6.77697
R646 a_153429_n11365.n261 a_153429_n11365.n260 6.77697
R647 a_153429_n11365.n247 a_153429_n11365.n246 6.77697
R648 a_153429_n11365.n233 a_153429_n11365.n232 6.77697
R649 a_153429_n11365.n219 a_153429_n11365.n218 6.77697
R650 a_153429_n11365.n205 a_153429_n11365.n204 6.77697
R651 a_153429_n11365.n191 a_153429_n11365.n190 6.77697
R652 a_153429_n11365.n177 a_153429_n11365.n176 6.77697
R653 a_153429_n11365.n163 a_153429_n11365.n162 6.77697
R654 a_153429_n11365.n149 a_153429_n11365.n148 6.77697
R655 a_153429_n11365.n138 a_153429_n11365.n119 6.77697
R656 a_153429_n11365.n46 a_153429_n11365.n40 6.77697
R657 a_153429_n11365.n73 a_153429_n11365.n68 6.77697
R658 a_153429_n11365.n89 a_153429_n11365.n84 6.77697
R659 a_153429_n11365.n105 a_153429_n11365.n100 6.77697
R660 a_153429_n11365.n280 a_153429_n11365.t18 5.7135
R661 a_153429_n11365.n280 a_153429_n11365.t11 5.7135
R662 a_153429_n11365.n266 a_153429_n11365.t26 5.7135
R663 a_153429_n11365.n266 a_153429_n11365.t21 5.7135
R664 a_153429_n11365.n252 a_153429_n11365.t22 5.7135
R665 a_153429_n11365.n252 a_153429_n11365.t8 5.7135
R666 a_153429_n11365.n238 a_153429_n11365.t15 5.7135
R667 a_153429_n11365.n238 a_153429_n11365.t13 5.7135
R668 a_153429_n11365.n224 a_153429_n11365.t19 5.7135
R669 a_153429_n11365.n224 a_153429_n11365.t16 5.7135
R670 a_153429_n11365.n210 a_153429_n11365.t24 5.7135
R671 a_153429_n11365.n210 a_153429_n11365.t25 5.7135
R672 a_153429_n11365.n196 a_153429_n11365.t12 5.7135
R673 a_153429_n11365.n196 a_153429_n11365.t9 5.7135
R674 a_153429_n11365.n182 a_153429_n11365.t17 5.7135
R675 a_153429_n11365.n182 a_153429_n11365.t14 5.7135
R676 a_153429_n11365.n168 a_153429_n11365.t20 5.7135
R677 a_153429_n11365.n168 a_153429_n11365.t6 5.7135
R678 a_153429_n11365.n154 a_153429_n11365.t7 5.7135
R679 a_153429_n11365.n154 a_153429_n11365.t23 5.7135
R680 a_153429_n11365.n285 a_153429_n11365.n284 5.58552
R681 a_153429_n11365.n114 a_153429_n11365.n5 5.58552
R682 a_153429_n11365.n54 a_153429_n11365.n36 5.33935
R683 a_153429_n11365.n135 a_153429_n11365.n134 5.27109
R684 a_153429_n11365.n51 a_153429_n11365.n49 5.27109
R685 a_153429_n11365.n77 a_153429_n11365.n76 5.27109
R686 a_153429_n11365.n93 a_153429_n11365.n92 5.27109
R687 a_153429_n11365.n109 a_153429_n11365.n108 5.27109
R688 a_153429_n11365.n127 a_153429_n11365.n123 4.51911
R689 a_153429_n11365.n114 a_153429_n11365.n113 3.82472
R690 a_153429_n11365.n284 a_153429_n11365.n62 3.80493
R691 a_153429_n11365.n131 a_153429_n11365.n120 3.76521
R692 a_153429_n11365.n50 a_153429_n11365.n37 3.76521
R693 a_153429_n11365.n80 a_153429_n11365.n79 3.75827
R694 a_153429_n11365.n96 a_153429_n11365.n95 3.75827
R695 a_153429_n11365.n112 a_153429_n11365.n111 3.75827
R696 a_153429_n11365.n67 a_153429_n11365.t2 3.4805
R697 a_153429_n11365.n67 a_153429_n11365.t0 3.4805
R698 a_153429_n11365.n83 a_153429_n11365.t3 3.4805
R699 a_153429_n11365.n83 a_153429_n11365.t27 3.4805
R700 a_153429_n11365.n99 a_153429_n11365.t30 3.4805
R701 a_153429_n11365.n99 a_153429_n11365.t28 3.4805
R702 a_153429_n11365.n279 a_153429_n11365.n270 3.43565
R703 a_153429_n11365.n265 a_153429_n11365.n256 3.43565
R704 a_153429_n11365.n251 a_153429_n11365.n242 3.43565
R705 a_153429_n11365.n237 a_153429_n11365.n228 3.43565
R706 a_153429_n11365.n223 a_153429_n11365.n214 3.43565
R707 a_153429_n11365.n209 a_153429_n11365.n200 3.43565
R708 a_153429_n11365.n195 a_153429_n11365.n186 3.43565
R709 a_153429_n11365.n181 a_153429_n11365.n172 3.43565
R710 a_153429_n11365.n167 a_153429_n11365.n158 3.43565
R711 a_153429_n11365.n153 a_153429_n11365.n144 3.43565
R712 a_153429_n11365.t1 a_153429_n11365.n336 2.84983
R713 a_153429_n11365.n21 a_153429_n11365.t31 2.83311
R714 a_153429_n11365.n336 a_153429_n11365.t5 2.7853
R715 a_153429_n11365.n21 a_153429_n11365.t29 2.77004
R716 a_153429_n11365.n130 a_153429_n11365.n122 2.25932
R717 a_153429_n11365.n59 a_153429_n11365.n58 2.25932
R718 a_153429_n11365.n284 a_153429_n11365.n283 1.75537
R719 a_153429_n11365.n143 a_153429_n11365.n114 1.72874
R720 a_153429_n11365.n335 a_153429_n11365.n334 1.11019
R721 a_153429_n11365.n23 a_153429_n11365.n22 1.09519
R722 a_153429_n11365.n335 a_153429_n11365.n0 1.06331
R723 a_153429_n11365.n24 a_153429_n11365.n22 1.04831
R724 a_153429_n11365.n126 a_153429_n11365.n125 0.753441
R725 a_153429_n11365.n55 a_153429_n11365.n38 0.753441
R726 a_153429_n11365.n334 a_153429_n11365.n333 0.3955
R727 a_153429_n11365.n333 a_153429_n11365.n1 0.3955
R728 a_153429_n11365.n329 a_153429_n11365.n1 0.3955
R729 a_153429_n11365.n329 a_153429_n11365.n328 0.3955
R730 a_153429_n11365.n328 a_153429_n11365.n327 0.3955
R731 a_153429_n11365.n327 a_153429_n11365.n3 0.3955
R732 a_153429_n11365.n322 a_153429_n11365.n321 0.3955
R733 a_153429_n11365.n321 a_153429_n11365.n6 0.3955
R734 a_153429_n11365.n317 a_153429_n11365.n6 0.3955
R735 a_153429_n11365.n317 a_153429_n11365.n316 0.3955
R736 a_153429_n11365.n316 a_153429_n11365.n315 0.3955
R737 a_153429_n11365.n315 a_153429_n11365.n8 0.3955
R738 a_153429_n11365.n311 a_153429_n11365.n8 0.3955
R739 a_153429_n11365.n311 a_153429_n11365.n310 0.3955
R740 a_153429_n11365.n310 a_153429_n11365.n309 0.3955
R741 a_153429_n11365.n309 a_153429_n11365.n10 0.3955
R742 a_153429_n11365.n305 a_153429_n11365.n10 0.3955
R743 a_153429_n11365.n305 a_153429_n11365.n304 0.3955
R744 a_153429_n11365.n304 a_153429_n11365.n303 0.3955
R745 a_153429_n11365.n303 a_153429_n11365.n12 0.3955
R746 a_153429_n11365.n299 a_153429_n11365.n12 0.3955
R747 a_153429_n11365.n299 a_153429_n11365.n298 0.3955
R748 a_153429_n11365.n298 a_153429_n11365.n297 0.3955
R749 a_153429_n11365.n297 a_153429_n11365.n14 0.3955
R750 a_153429_n11365.n293 a_153429_n11365.n14 0.3955
R751 a_153429_n11365.n293 a_153429_n11365.n292 0.3955
R752 a_153429_n11365.n292 a_153429_n11365.n291 0.3955
R753 a_153429_n11365.n291 a_153429_n11365.n16 0.3955
R754 a_153429_n11365.n287 a_153429_n11365.n16 0.3955
R755 a_153429_n11365.n33 a_153429_n11365.n18 0.3955
R756 a_153429_n11365.n29 a_153429_n11365.n18 0.3955
R757 a_153429_n11365.n29 a_153429_n11365.n28 0.3955
R758 a_153429_n11365.n28 a_153429_n11365.n27 0.3955
R759 a_153429_n11365.n27 a_153429_n11365.n20 0.3955
R760 a_153429_n11365.n23 a_153429_n11365.n20 0.3955
R761 a_153429_n11365.n332 a_153429_n11365.n0 0.3955
R762 a_153429_n11365.n332 a_153429_n11365.n331 0.3955
R763 a_153429_n11365.n331 a_153429_n11365.n330 0.3955
R764 a_153429_n11365.n330 a_153429_n11365.n2 0.3955
R765 a_153429_n11365.n326 a_153429_n11365.n2 0.3955
R766 a_153429_n11365.n326 a_153429_n11365.n325 0.3955
R767 a_153429_n11365.n325 a_153429_n11365.n324 0.3955
R768 a_153429_n11365.n324 a_153429_n11365.n4 0.3955
R769 a_153429_n11365.n320 a_153429_n11365.n4 0.3955
R770 a_153429_n11365.n320 a_153429_n11365.n319 0.3955
R771 a_153429_n11365.n319 a_153429_n11365.n318 0.3955
R772 a_153429_n11365.n318 a_153429_n11365.n7 0.3955
R773 a_153429_n11365.n314 a_153429_n11365.n7 0.3955
R774 a_153429_n11365.n314 a_153429_n11365.n313 0.3955
R775 a_153429_n11365.n313 a_153429_n11365.n312 0.3955
R776 a_153429_n11365.n312 a_153429_n11365.n9 0.3955
R777 a_153429_n11365.n308 a_153429_n11365.n9 0.3955
R778 a_153429_n11365.n308 a_153429_n11365.n307 0.3955
R779 a_153429_n11365.n307 a_153429_n11365.n306 0.3955
R780 a_153429_n11365.n306 a_153429_n11365.n11 0.3955
R781 a_153429_n11365.n302 a_153429_n11365.n11 0.3955
R782 a_153429_n11365.n302 a_153429_n11365.n301 0.3955
R783 a_153429_n11365.n301 a_153429_n11365.n300 0.3955
R784 a_153429_n11365.n300 a_153429_n11365.n13 0.3955
R785 a_153429_n11365.n296 a_153429_n11365.n13 0.3955
R786 a_153429_n11365.n296 a_153429_n11365.n295 0.3955
R787 a_153429_n11365.n295 a_153429_n11365.n294 0.3955
R788 a_153429_n11365.n294 a_153429_n11365.n15 0.3955
R789 a_153429_n11365.n290 a_153429_n11365.n15 0.3955
R790 a_153429_n11365.n290 a_153429_n11365.n289 0.3955
R791 a_153429_n11365.n289 a_153429_n11365.n288 0.3955
R792 a_153429_n11365.n288 a_153429_n11365.n17 0.3955
R793 a_153429_n11365.n32 a_153429_n11365.n17 0.3955
R794 a_153429_n11365.n32 a_153429_n11365.n31 0.3955
R795 a_153429_n11365.n31 a_153429_n11365.n30 0.3955
R796 a_153429_n11365.n30 a_153429_n11365.n19 0.3955
R797 a_153429_n11365.n26 a_153429_n11365.n19 0.3955
R798 a_153429_n11365.n26 a_153429_n11365.n25 0.3955
R799 a_153429_n11365.n25 a_153429_n11365.n24 0.3955
R800 a_153429_n11365.n287 a_153429_n11365.n286 0.370955
R801 a_153429_n11365.n323 a_153429_n11365.n322 0.351864
R802 a_153429_n11365.n22 a_153429_n11365.n21 0.349638
R803 a_153429_n11365.n336 a_153429_n11365.n335 0.349638
R804 a_153429_n11365.n277 a_153429_n11365.n276 0.196152
R805 a_153429_n11365.n263 a_153429_n11365.n262 0.196152
R806 a_153429_n11365.n249 a_153429_n11365.n248 0.196152
R807 a_153429_n11365.n235 a_153429_n11365.n234 0.196152
R808 a_153429_n11365.n221 a_153429_n11365.n220 0.196152
R809 a_153429_n11365.n207 a_153429_n11365.n206 0.196152
R810 a_153429_n11365.n193 a_153429_n11365.n192 0.196152
R811 a_153429_n11365.n179 a_153429_n11365.n178 0.196152
R812 a_153429_n11365.n165 a_153429_n11365.n164 0.196152
R813 a_153429_n11365.n151 a_153429_n11365.n150 0.196152
R814 a_153429_n11365.n129 a_153429_n11365.n127 0.196152
R815 a_153429_n11365.n137 a_153429_n11365.n136 0.196152
R816 a_153429_n11365.n48 a_153429_n11365.n47 0.196152
R817 a_153429_n11365.n48 a_153429_n11365.n35 0.196152
R818 a_153429_n11365.n75 a_153429_n11365.n74 0.196152
R819 a_153429_n11365.n75 a_153429_n11365.n66 0.196152
R820 a_153429_n11365.n91 a_153429_n11365.n90 0.196152
R821 a_153429_n11365.n91 a_153429_n11365.n82 0.196152
R822 a_153429_n11365.n107 a_153429_n11365.n106 0.196152
R823 a_153429_n11365.n107 a_153429_n11365.n98 0.196152
R824 a_153429_n11365.n129 a_153429_n11365.n128 0.194824
R825 a_153429_n11365.n276 a_153429_n11365.n271 0.186853
R826 a_153429_n11365.n262 a_153429_n11365.n257 0.186853
R827 a_153429_n11365.n248 a_153429_n11365.n243 0.186853
R828 a_153429_n11365.n234 a_153429_n11365.n229 0.186853
R829 a_153429_n11365.n220 a_153429_n11365.n215 0.186853
R830 a_153429_n11365.n206 a_153429_n11365.n201 0.186853
R831 a_153429_n11365.n192 a_153429_n11365.n187 0.186853
R832 a_153429_n11365.n178 a_153429_n11365.n173 0.186853
R833 a_153429_n11365.n164 a_153429_n11365.n159 0.186853
R834 a_153429_n11365.n150 a_153429_n11365.n145 0.186853
R835 a_153429_n11365.n137 a_153429_n11365.n116 0.186853
R836 a_153429_n11365.n47 a_153429_n11365.n41 0.186853
R837 a_153429_n11365.n74 a_153429_n11365.n69 0.186853
R838 a_153429_n11365.n90 a_153429_n11365.n85 0.186853
R839 a_153429_n11365.n106 a_153429_n11365.n101 0.186853
R840 a_153429_n11365.n60 a_153429_n11365.n36 0.184196
R841 a_153429_n11365.n5 a_153429_n11365.n3 0.166409
R842 a_153429_n11365.n285 a_153429_n11365.n33 0.131409
R843 a_153429_n11365.n61 a_153429_n11365.n35 0.0790024
R844 a_153429_n11365.n80 a_153429_n11365.n66 0.0790024
R845 a_153429_n11365.n96 a_153429_n11365.n82 0.0790024
R846 a_153429_n11365.n112 a_153429_n11365.n98 0.0790024
R847 a_153429_n11365.n286 a_153429_n11365.n285 0.0709545
R848 a_153429_n11365.n277 a_153429_n11365.n270 0.0572633
R849 a_153429_n11365.n263 a_153429_n11365.n256 0.0572633
R850 a_153429_n11365.n249 a_153429_n11365.n242 0.0572633
R851 a_153429_n11365.n235 a_153429_n11365.n228 0.0572633
R852 a_153429_n11365.n221 a_153429_n11365.n214 0.0572633
R853 a_153429_n11365.n207 a_153429_n11365.n200 0.0572633
R854 a_153429_n11365.n193 a_153429_n11365.n186 0.0572633
R855 a_153429_n11365.n179 a_153429_n11365.n172 0.0572633
R856 a_153429_n11365.n165 a_153429_n11365.n158 0.0572633
R857 a_153429_n11365.n151 a_153429_n11365.n144 0.0572633
R858 a_153429_n11365.n136 a_153429_n11365.n115 0.0572633
R859 a_153429_n11365.n323 a_153429_n11365.n5 0.0550455
R860 a_153429_n11365.n171 a_153429_n11365.n157 0.0506333
R861 a_153429_n11365.n185 a_153429_n11365.n171 0.0506333
R862 a_153429_n11365.n213 a_153429_n11365.n199 0.0506333
R863 a_153429_n11365.n241 a_153429_n11365.n227 0.0506333
R864 a_153429_n11365.n255 a_153429_n11365.n241 0.0506333
R865 a_153429_n11365.n283 a_153429_n11365.n269 0.0506333
R866 a_153429_n11365.n157 a_153429_n11365.n143 0.0490667
R867 a_153429_n11365.n199 a_153429_n11365.n185 0.0490667
R868 a_153429_n11365.n227 a_153429_n11365.n213 0.0490667
R869 a_153429_n11365.n269 a_153429_n11365.n255 0.0490667
R870 a_153429_n11365.n128 a_153429_n11365.n115 0.0477222
R871 a_153429_n11365.n113 a_153429_n11365.n97 0.0400789
R872 a_153429_n11365.n81 a_153429_n11365.n62 0.0400789
R873 a_153429_n11365.n282 a_153429_n11365.n271 0.0393889
R874 a_153429_n11365.n268 a_153429_n11365.n257 0.0393889
R875 a_153429_n11365.n254 a_153429_n11365.n243 0.0393889
R876 a_153429_n11365.n240 a_153429_n11365.n229 0.0393889
R877 a_153429_n11365.n226 a_153429_n11365.n215 0.0393889
R878 a_153429_n11365.n212 a_153429_n11365.n201 0.0393889
R879 a_153429_n11365.n198 a_153429_n11365.n187 0.0393889
R880 a_153429_n11365.n184 a_153429_n11365.n173 0.0393889
R881 a_153429_n11365.n170 a_153429_n11365.n159 0.0393889
R882 a_153429_n11365.n156 a_153429_n11365.n145 0.0393889
R883 a_153429_n11365.n142 a_153429_n11365.n116 0.0393889
R884 a_153429_n11365.n41 a_153429_n11365.n34 0.0393889
R885 a_153429_n11365.n69 a_153429_n11365.n65 0.0393889
R886 a_153429_n11365.n85 a_153429_n11365.n64 0.0393889
R887 a_153429_n11365.n101 a_153429_n11365.n63 0.0393889
R888 a_153429_n11365.n97 a_153429_n11365.n81 0.0388421
R889 a_153429_n11365.n61 a_153429_n11365.n60 0.0366111
R890 VDD.n5240 VDD.n5192 5911.77
R891 VDD.n5240 VDD.n5193 5911.77
R892 VDD.n5239 VDD.n5192 5911.77
R893 VDD.n5239 VDD.n5193 5911.77
R894 VDD.n5229 VDD.n5194 5911.77
R895 VDD.n5229 VDD.n5195 5911.77
R896 VDD.n5225 VDD.n5195 5911.77
R897 VDD.n5225 VDD.n5194 5911.77
R898 VDD.n5296 VDD.n5251 5911.77
R899 VDD.n5298 VDD.n5251 5911.77
R900 VDD.n5296 VDD.n5252 5911.77
R901 VDD.n5298 VDD.n5252 5911.77
R902 VDD.n5285 VDD.n5258 5911.77
R903 VDD.n5285 VDD.n5284 5911.77
R904 VDD.n5284 VDD.n5283 5911.77
R905 VDD.n5283 VDD.n5258 5911.77
R906 VDD.n5212 VDD.n5203 3370.59
R907 VDD.n5212 VDD.n5204 3370.59
R908 VDD.n5210 VDD.n5204 3370.59
R909 VDD.n5210 VDD.n5203 3370.59
R910 VDD.n5272 VDD.n5263 3370.59
R911 VDD.n5272 VDD.n5264 3370.59
R912 VDD.n5270 VDD.n5264 3370.59
R913 VDD.n5270 VDD.n5263 3370.59
R914 VDD.n5456 VDD.t694 877.144
R915 VDD.n5332 VDD.t709 877.144
R916 VDD.n3127 VDD.n3125 815.966
R917 VDD.n3202 VDD.n3180 815.966
R918 VDD.n3623 VDD.n3601 815.966
R919 VDD.n3483 VDD.n3461 815.966
R920 VDD.n533 VDD.n531 815.966
R921 VDD.n608 VDD.n586 815.966
R922 VDD.n1029 VDD.n1007 815.966
R923 VDD.n889 VDD.n867 815.966
R924 VDD.n6096 VDD.n6094 815.966
R925 VDD.n6171 VDD.n6149 815.966
R926 VDD.n6592 VDD.n6570 815.966
R927 VDD.n6452 VDD.n6430 815.966
R928 VDD.n4243 VDD.n4201 765.883
R929 VDD.n4900 VDD.n4834 765.883
R930 VDD.n4869 VDD.n4836 765.883
R931 VDD.n4240 VDD.n4199 765.883
R932 VDD.n1649 VDD.n1607 765.883
R933 VDD.n2306 VDD.n2240 765.883
R934 VDD.n2275 VDD.n2242 765.883
R935 VDD.n1646 VDD.n1605 765.883
R936 VDD.n7212 VDD.n7170 765.883
R937 VDD.n7869 VDD.n7803 765.883
R938 VDD.n7838 VDD.n7805 765.883
R939 VDD.n7209 VDD.n7168 765.883
R940 VDD.n4422 VDD.n4387 748.236
R941 VDD.n5074 VDD.n3885 748.236
R942 VDD.n4390 VDD.n4137 748.236
R943 VDD.n5034 VDD.n3887 748.236
R944 VDD.n4385 VDD.n4143 748.236
R945 VDD.n5072 VDD.n3890 748.236
R946 VDD.n4425 VDD.n4139 748.236
R947 VDD.n3907 VDD.n3888 748.236
R948 VDD.n1828 VDD.n1793 748.236
R949 VDD.n2480 VDD.n1291 748.236
R950 VDD.n1796 VDD.n1543 748.236
R951 VDD.n2440 VDD.n1293 748.236
R952 VDD.n1791 VDD.n1549 748.236
R953 VDD.n2478 VDD.n1296 748.236
R954 VDD.n1831 VDD.n1545 748.236
R955 VDD.n1313 VDD.n1294 748.236
R956 VDD.n7391 VDD.n7356 748.236
R957 VDD.n8043 VDD.n6854 748.236
R958 VDD.n7359 VDD.n7106 748.236
R959 VDD.n8003 VDD.n6856 748.236
R960 VDD.n7354 VDD.n7112 748.236
R961 VDD.n8041 VDD.n6859 748.236
R962 VDD.n7394 VDD.n7108 748.236
R963 VDD.n6876 VDD.n6857 748.236
R964 VDD.n2671 VDD.n2670 744.707
R965 VDD.n3015 VDD.n2734 744.707
R966 VDD.n3087 VDD.n2629 744.707
R967 VDD.n2978 VDD.n2732 744.707
R968 VDD.n2803 VDD.n2636 744.707
R969 VDD.n3017 VDD.n2730 744.707
R970 VDD.n2886 VDD.n2731 744.707
R971 VDD.n2849 VDD.n2848 744.707
R972 VDD.n77 VDD.n76 744.707
R973 VDD.n421 VDD.n140 744.707
R974 VDD.n493 VDD.n35 744.707
R975 VDD.n384 VDD.n138 744.707
R976 VDD.n209 VDD.n42 744.707
R977 VDD.n423 VDD.n136 744.707
R978 VDD.n292 VDD.n137 744.707
R979 VDD.n255 VDD.n254 744.707
R980 VDD.n5640 VDD.n5639 744.707
R981 VDD.n5984 VDD.n5703 744.707
R982 VDD.n6056 VDD.n5598 744.707
R983 VDD.n5947 VDD.n5701 744.707
R984 VDD.n5772 VDD.n5605 744.707
R985 VDD.n5986 VDD.n5699 744.707
R986 VDD.n5855 VDD.n5700 744.707
R987 VDD.n5818 VDD.n5817 744.707
R988 VDD.n5238 VDD.n5190 630.588
R989 VDD.n5238 VDD.n5237 630.588
R990 VDD.n5228 VDD.n5227 630.588
R991 VDD.n5227 VDD.n5226 630.588
R992 VDD.n5295 VDD.n5250 630.588
R993 VDD.n5299 VDD.n5250 630.588
R994 VDD.n5286 VDD.n5257 630.588
R995 VDD.n5282 VDD.n5257 630.588
R996 VDD.n2615 VDD.n2614 585
R997 VDD.n2613 VDD.n2612 585
R998 VDD.n2604 VDD.n2603 585
R999 VDD.n2607 VDD.n2606 585
R1000 VDD.n2934 VDD.n2933 585
R1001 VDD.n2932 VDD.n2931 585
R1002 VDD.n2923 VDD.n2922 585
R1003 VDD.n2926 VDD.n2925 585
R1004 VDD.n2909 VDD.n2908 585
R1005 VDD.n2907 VDD.n2906 585
R1006 VDD.n2746 VDD.n2745 585
R1007 VDD.n2751 VDD.n2750 585
R1008 VDD.n2787 VDD.n2786 585
R1009 VDD.n2828 VDD.n2827 585
R1010 VDD.n2830 VDD.n2829 585
R1011 VDD.n2831 VDD.n2784 585
R1012 VDD.n3126 VDD.n3125 585
R1013 VDD.n3134 VDD.n3133 585
R1014 VDD.n3135 VDD.n3123 585
R1015 VDD.n3144 VDD.n3143 585
R1016 VDD.n3142 VDD.n3141 585
R1017 VDD.n3137 VDD.n3136 585
R1018 VDD.n3152 VDD.n3150 585
R1019 VDD.n3151 VDD.n3150 585
R1020 VDD.n3157 VDD.n3150 585
R1021 VDD.n3385 VDD.n3383 585
R1022 VDD.n3384 VDD.n3383 585
R1023 VDD.n3390 VDD.n3383 585
R1024 VDD.n3398 VDD.n3396 585
R1025 VDD.n3397 VDD.n3396 585
R1026 VDD.n3403 VDD.n3396 585
R1027 VDD.n3411 VDD.n3409 585
R1028 VDD.n3410 VDD.n3409 585
R1029 VDD.n3416 VDD.n3409 585
R1030 VDD.n3424 VDD.n3422 585
R1031 VDD.n3423 VDD.n3422 585
R1032 VDD.n3429 VDD.n3422 585
R1033 VDD.n3368 VDD.n3366 585
R1034 VDD.n3367 VDD.n3366 585
R1035 VDD.n3373 VDD.n3366 585
R1036 VDD.n3354 VDD.n3352 585
R1037 VDD.n3353 VDD.n3352 585
R1038 VDD.n3359 VDD.n3352 585
R1039 VDD.n3340 VDD.n3338 585
R1040 VDD.n3339 VDD.n3338 585
R1041 VDD.n3345 VDD.n3338 585
R1042 VDD.n3108 VDD.n3106 585
R1043 VDD.n3107 VDD.n3106 585
R1044 VDD.n3113 VDD.n3106 585
R1045 VDD.n5165 VDD.n5163 585
R1046 VDD.n5164 VDD.n5163 585
R1047 VDD.n5170 VDD.n5163 585
R1048 VDD.n3203 VDD.n3202 585
R1049 VDD.n3201 VDD.n3200 585
R1050 VDD.n3197 VDD.n3183 585
R1051 VDD.n3187 VDD.n3184 585
R1052 VDD.n3192 VDD.n3191 585
R1053 VDD.n3190 VDD.n3189 585
R1054 VDD.n3215 VDD.n3208 585
R1055 VDD.n3216 VDD.n3215 585
R1056 VDD.n3215 VDD.n3214 585
R1057 VDD.n3289 VDD.n3282 585
R1058 VDD.n3290 VDD.n3289 585
R1059 VDD.n3289 VDD.n3288 585
R1060 VDD.n3302 VDD.n3295 585
R1061 VDD.n3303 VDD.n3302 585
R1062 VDD.n3302 VDD.n3301 585
R1063 VDD.n3315 VDD.n3308 585
R1064 VDD.n3316 VDD.n3315 585
R1065 VDD.n3315 VDD.n3314 585
R1066 VDD.n3328 VDD.n3321 585
R1067 VDD.n3329 VDD.n3328 585
R1068 VDD.n3328 VDD.n3327 585
R1069 VDD.n3272 VDD.n3265 585
R1070 VDD.n3273 VDD.n3272 585
R1071 VDD.n3272 VDD.n3271 585
R1072 VDD.n3258 VDD.n3251 585
R1073 VDD.n3259 VDD.n3258 585
R1074 VDD.n3258 VDD.n3257 585
R1075 VDD.n3244 VDD.n3237 585
R1076 VDD.n3245 VDD.n3244 585
R1077 VDD.n3244 VDD.n3243 585
R1078 VDD.n3230 VDD.n3223 585
R1079 VDD.n3231 VDD.n3230 585
R1080 VDD.n3230 VDD.n3229 585
R1081 VDD.n3171 VDD.n3164 585
R1082 VDD.n3172 VDD.n3171 585
R1083 VDD.n3171 VDD.n3170 585
R1084 VDD.n3624 VDD.n3623 585
R1085 VDD.n3622 VDD.n3621 585
R1086 VDD.n3618 VDD.n3604 585
R1087 VDD.n3608 VDD.n3605 585
R1088 VDD.n3613 VDD.n3612 585
R1089 VDD.n3611 VDD.n3610 585
R1090 VDD.n3636 VDD.n3629 585
R1091 VDD.n3637 VDD.n3636 585
R1092 VDD.n3636 VDD.n3635 585
R1093 VDD.n3650 VDD.n3643 585
R1094 VDD.n3651 VDD.n3650 585
R1095 VDD.n3650 VDD.n3649 585
R1096 VDD.n3663 VDD.n3656 585
R1097 VDD.n3664 VDD.n3663 585
R1098 VDD.n3663 VDD.n3662 585
R1099 VDD.n3676 VDD.n3669 585
R1100 VDD.n3677 VDD.n3676 585
R1101 VDD.n3676 VDD.n3675 585
R1102 VDD.n3689 VDD.n3682 585
R1103 VDD.n3690 VDD.n3689 585
R1104 VDD.n3689 VDD.n3688 585
R1105 VDD.n3702 VDD.n3695 585
R1106 VDD.n3703 VDD.n3702 585
R1107 VDD.n3702 VDD.n3701 585
R1108 VDD.n3715 VDD.n3708 585
R1109 VDD.n3716 VDD.n3715 585
R1110 VDD.n3715 VDD.n3714 585
R1111 VDD.n3729 VDD.n3722 585
R1112 VDD.n3730 VDD.n3729 585
R1113 VDD.n3729 VDD.n3728 585
R1114 VDD.n3742 VDD.n3735 585
R1115 VDD.n3743 VDD.n3742 585
R1116 VDD.n3742 VDD.n3741 585
R1117 VDD.n3755 VDD.n3748 585
R1118 VDD.n3756 VDD.n3755 585
R1119 VDD.n3755 VDD.n3754 585
R1120 VDD.n3768 VDD.n3761 585
R1121 VDD.n3769 VDD.n3768 585
R1122 VDD.n3768 VDD.n3767 585
R1123 VDD.n3781 VDD.n3774 585
R1124 VDD.n3782 VDD.n3781 585
R1125 VDD.n3781 VDD.n3780 585
R1126 VDD.n3582 VDD.n3575 585
R1127 VDD.n3583 VDD.n3582 585
R1128 VDD.n3582 VDD.n3581 585
R1129 VDD.n3568 VDD.n3561 585
R1130 VDD.n3569 VDD.n3568 585
R1131 VDD.n3568 VDD.n3567 585
R1132 VDD.n3554 VDD.n3547 585
R1133 VDD.n3555 VDD.n3554 585
R1134 VDD.n3554 VDD.n3553 585
R1135 VDD.n3540 VDD.n3533 585
R1136 VDD.n3541 VDD.n3540 585
R1137 VDD.n3540 VDD.n3539 585
R1138 VDD.n3526 VDD.n3519 585
R1139 VDD.n3527 VDD.n3526 585
R1140 VDD.n3526 VDD.n3525 585
R1141 VDD.n3512 VDD.n3505 585
R1142 VDD.n3513 VDD.n3512 585
R1143 VDD.n3512 VDD.n3511 585
R1144 VDD.n3497 VDD.n3490 585
R1145 VDD.n3498 VDD.n3497 585
R1146 VDD.n3497 VDD.n3496 585
R1147 VDD.n3484 VDD.n3483 585
R1148 VDD.n3482 VDD.n3481 585
R1149 VDD.n3478 VDD.n3464 585
R1150 VDD.n3468 VDD.n3465 585
R1151 VDD.n3473 VDD.n3472 585
R1152 VDD.n3471 VDD.n3470 585
R1153 VDD.n21 VDD.n20 585
R1154 VDD.n19 VDD.n18 585
R1155 VDD.n10 VDD.n9 585
R1156 VDD.n13 VDD.n12 585
R1157 VDD.n340 VDD.n339 585
R1158 VDD.n338 VDD.n337 585
R1159 VDD.n329 VDD.n328 585
R1160 VDD.n332 VDD.n331 585
R1161 VDD.n315 VDD.n314 585
R1162 VDD.n313 VDD.n312 585
R1163 VDD.n152 VDD.n151 585
R1164 VDD.n157 VDD.n156 585
R1165 VDD.n193 VDD.n192 585
R1166 VDD.n234 VDD.n233 585
R1167 VDD.n236 VDD.n235 585
R1168 VDD.n237 VDD.n190 585
R1169 VDD.n532 VDD.n531 585
R1170 VDD.n540 VDD.n539 585
R1171 VDD.n541 VDD.n529 585
R1172 VDD.n550 VDD.n549 585
R1173 VDD.n548 VDD.n547 585
R1174 VDD.n543 VDD.n542 585
R1175 VDD.n558 VDD.n556 585
R1176 VDD.n557 VDD.n556 585
R1177 VDD.n563 VDD.n556 585
R1178 VDD.n791 VDD.n789 585
R1179 VDD.n790 VDD.n789 585
R1180 VDD.n796 VDD.n789 585
R1181 VDD.n804 VDD.n802 585
R1182 VDD.n803 VDD.n802 585
R1183 VDD.n809 VDD.n802 585
R1184 VDD.n817 VDD.n815 585
R1185 VDD.n816 VDD.n815 585
R1186 VDD.n822 VDD.n815 585
R1187 VDD.n830 VDD.n828 585
R1188 VDD.n829 VDD.n828 585
R1189 VDD.n835 VDD.n828 585
R1190 VDD.n774 VDD.n772 585
R1191 VDD.n773 VDD.n772 585
R1192 VDD.n779 VDD.n772 585
R1193 VDD.n760 VDD.n758 585
R1194 VDD.n759 VDD.n758 585
R1195 VDD.n765 VDD.n758 585
R1196 VDD.n746 VDD.n744 585
R1197 VDD.n745 VDD.n744 585
R1198 VDD.n751 VDD.n744 585
R1199 VDD.n514 VDD.n512 585
R1200 VDD.n513 VDD.n512 585
R1201 VDD.n519 VDD.n512 585
R1202 VDD.n2571 VDD.n2569 585
R1203 VDD.n2570 VDD.n2569 585
R1204 VDD.n2576 VDD.n2569 585
R1205 VDD.n609 VDD.n608 585
R1206 VDD.n607 VDD.n606 585
R1207 VDD.n603 VDD.n589 585
R1208 VDD.n593 VDD.n590 585
R1209 VDD.n598 VDD.n597 585
R1210 VDD.n596 VDD.n595 585
R1211 VDD.n621 VDD.n614 585
R1212 VDD.n622 VDD.n621 585
R1213 VDD.n621 VDD.n620 585
R1214 VDD.n695 VDD.n688 585
R1215 VDD.n696 VDD.n695 585
R1216 VDD.n695 VDD.n694 585
R1217 VDD.n708 VDD.n701 585
R1218 VDD.n709 VDD.n708 585
R1219 VDD.n708 VDD.n707 585
R1220 VDD.n721 VDD.n714 585
R1221 VDD.n722 VDD.n721 585
R1222 VDD.n721 VDD.n720 585
R1223 VDD.n734 VDD.n727 585
R1224 VDD.n735 VDD.n734 585
R1225 VDD.n734 VDD.n733 585
R1226 VDD.n678 VDD.n671 585
R1227 VDD.n679 VDD.n678 585
R1228 VDD.n678 VDD.n677 585
R1229 VDD.n664 VDD.n657 585
R1230 VDD.n665 VDD.n664 585
R1231 VDD.n664 VDD.n663 585
R1232 VDD.n650 VDD.n643 585
R1233 VDD.n651 VDD.n650 585
R1234 VDD.n650 VDD.n649 585
R1235 VDD.n636 VDD.n629 585
R1236 VDD.n637 VDD.n636 585
R1237 VDD.n636 VDD.n635 585
R1238 VDD.n577 VDD.n570 585
R1239 VDD.n578 VDD.n577 585
R1240 VDD.n577 VDD.n576 585
R1241 VDD.n1030 VDD.n1029 585
R1242 VDD.n1028 VDD.n1027 585
R1243 VDD.n1024 VDD.n1010 585
R1244 VDD.n1014 VDD.n1011 585
R1245 VDD.n1019 VDD.n1018 585
R1246 VDD.n1017 VDD.n1016 585
R1247 VDD.n1042 VDD.n1035 585
R1248 VDD.n1043 VDD.n1042 585
R1249 VDD.n1042 VDD.n1041 585
R1250 VDD.n1056 VDD.n1049 585
R1251 VDD.n1057 VDD.n1056 585
R1252 VDD.n1056 VDD.n1055 585
R1253 VDD.n1069 VDD.n1062 585
R1254 VDD.n1070 VDD.n1069 585
R1255 VDD.n1069 VDD.n1068 585
R1256 VDD.n1082 VDD.n1075 585
R1257 VDD.n1083 VDD.n1082 585
R1258 VDD.n1082 VDD.n1081 585
R1259 VDD.n1095 VDD.n1088 585
R1260 VDD.n1096 VDD.n1095 585
R1261 VDD.n1095 VDD.n1094 585
R1262 VDD.n1108 VDD.n1101 585
R1263 VDD.n1109 VDD.n1108 585
R1264 VDD.n1108 VDD.n1107 585
R1265 VDD.n1121 VDD.n1114 585
R1266 VDD.n1122 VDD.n1121 585
R1267 VDD.n1121 VDD.n1120 585
R1268 VDD.n1135 VDD.n1128 585
R1269 VDD.n1136 VDD.n1135 585
R1270 VDD.n1135 VDD.n1134 585
R1271 VDD.n1148 VDD.n1141 585
R1272 VDD.n1149 VDD.n1148 585
R1273 VDD.n1148 VDD.n1147 585
R1274 VDD.n1161 VDD.n1154 585
R1275 VDD.n1162 VDD.n1161 585
R1276 VDD.n1161 VDD.n1160 585
R1277 VDD.n1174 VDD.n1167 585
R1278 VDD.n1175 VDD.n1174 585
R1279 VDD.n1174 VDD.n1173 585
R1280 VDD.n1187 VDD.n1180 585
R1281 VDD.n1188 VDD.n1187 585
R1282 VDD.n1187 VDD.n1186 585
R1283 VDD.n988 VDD.n981 585
R1284 VDD.n989 VDD.n988 585
R1285 VDD.n988 VDD.n987 585
R1286 VDD.n974 VDD.n967 585
R1287 VDD.n975 VDD.n974 585
R1288 VDD.n974 VDD.n973 585
R1289 VDD.n960 VDD.n953 585
R1290 VDD.n961 VDD.n960 585
R1291 VDD.n960 VDD.n959 585
R1292 VDD.n946 VDD.n939 585
R1293 VDD.n947 VDD.n946 585
R1294 VDD.n946 VDD.n945 585
R1295 VDD.n932 VDD.n925 585
R1296 VDD.n933 VDD.n932 585
R1297 VDD.n932 VDD.n931 585
R1298 VDD.n918 VDD.n911 585
R1299 VDD.n919 VDD.n918 585
R1300 VDD.n918 VDD.n917 585
R1301 VDD.n903 VDD.n896 585
R1302 VDD.n904 VDD.n903 585
R1303 VDD.n903 VDD.n902 585
R1304 VDD.n890 VDD.n889 585
R1305 VDD.n888 VDD.n887 585
R1306 VDD.n884 VDD.n870 585
R1307 VDD.n874 VDD.n871 585
R1308 VDD.n879 VDD.n878 585
R1309 VDD.n877 VDD.n876 585
R1310 VDD.n5584 VDD.n5583 585
R1311 VDD.n5582 VDD.n5581 585
R1312 VDD.n5573 VDD.n5572 585
R1313 VDD.n5576 VDD.n5575 585
R1314 VDD.n5903 VDD.n5902 585
R1315 VDD.n5901 VDD.n5900 585
R1316 VDD.n5892 VDD.n5891 585
R1317 VDD.n5895 VDD.n5894 585
R1318 VDD.n5878 VDD.n5877 585
R1319 VDD.n5876 VDD.n5875 585
R1320 VDD.n5715 VDD.n5714 585
R1321 VDD.n5720 VDD.n5719 585
R1322 VDD.n5756 VDD.n5755 585
R1323 VDD.n5797 VDD.n5796 585
R1324 VDD.n5799 VDD.n5798 585
R1325 VDD.n5800 VDD.n5753 585
R1326 VDD.n6095 VDD.n6094 585
R1327 VDD.n6103 VDD.n6102 585
R1328 VDD.n6104 VDD.n6092 585
R1329 VDD.n6113 VDD.n6112 585
R1330 VDD.n6111 VDD.n6110 585
R1331 VDD.n6106 VDD.n6105 585
R1332 VDD.n6121 VDD.n6119 585
R1333 VDD.n6120 VDD.n6119 585
R1334 VDD.n6126 VDD.n6119 585
R1335 VDD.n6354 VDD.n6352 585
R1336 VDD.n6353 VDD.n6352 585
R1337 VDD.n6359 VDD.n6352 585
R1338 VDD.n6367 VDD.n6365 585
R1339 VDD.n6366 VDD.n6365 585
R1340 VDD.n6372 VDD.n6365 585
R1341 VDD.n6380 VDD.n6378 585
R1342 VDD.n6379 VDD.n6378 585
R1343 VDD.n6385 VDD.n6378 585
R1344 VDD.n6393 VDD.n6391 585
R1345 VDD.n6392 VDD.n6391 585
R1346 VDD.n6398 VDD.n6391 585
R1347 VDD.n6337 VDD.n6335 585
R1348 VDD.n6336 VDD.n6335 585
R1349 VDD.n6342 VDD.n6335 585
R1350 VDD.n6323 VDD.n6321 585
R1351 VDD.n6322 VDD.n6321 585
R1352 VDD.n6328 VDD.n6321 585
R1353 VDD.n6309 VDD.n6307 585
R1354 VDD.n6308 VDD.n6307 585
R1355 VDD.n6314 VDD.n6307 585
R1356 VDD.n6077 VDD.n6075 585
R1357 VDD.n6076 VDD.n6075 585
R1358 VDD.n6082 VDD.n6075 585
R1359 VDD.n8134 VDD.n8132 585
R1360 VDD.n8133 VDD.n8132 585
R1361 VDD.n8139 VDD.n8132 585
R1362 VDD.n6172 VDD.n6171 585
R1363 VDD.n6170 VDD.n6169 585
R1364 VDD.n6166 VDD.n6152 585
R1365 VDD.n6156 VDD.n6153 585
R1366 VDD.n6161 VDD.n6160 585
R1367 VDD.n6159 VDD.n6158 585
R1368 VDD.n6184 VDD.n6177 585
R1369 VDD.n6185 VDD.n6184 585
R1370 VDD.n6184 VDD.n6183 585
R1371 VDD.n6258 VDD.n6251 585
R1372 VDD.n6259 VDD.n6258 585
R1373 VDD.n6258 VDD.n6257 585
R1374 VDD.n6271 VDD.n6264 585
R1375 VDD.n6272 VDD.n6271 585
R1376 VDD.n6271 VDD.n6270 585
R1377 VDD.n6284 VDD.n6277 585
R1378 VDD.n6285 VDD.n6284 585
R1379 VDD.n6284 VDD.n6283 585
R1380 VDD.n6297 VDD.n6290 585
R1381 VDD.n6298 VDD.n6297 585
R1382 VDD.n6297 VDD.n6296 585
R1383 VDD.n6241 VDD.n6234 585
R1384 VDD.n6242 VDD.n6241 585
R1385 VDD.n6241 VDD.n6240 585
R1386 VDD.n6227 VDD.n6220 585
R1387 VDD.n6228 VDD.n6227 585
R1388 VDD.n6227 VDD.n6226 585
R1389 VDD.n6213 VDD.n6206 585
R1390 VDD.n6214 VDD.n6213 585
R1391 VDD.n6213 VDD.n6212 585
R1392 VDD.n6199 VDD.n6192 585
R1393 VDD.n6200 VDD.n6199 585
R1394 VDD.n6199 VDD.n6198 585
R1395 VDD.n6140 VDD.n6133 585
R1396 VDD.n6141 VDD.n6140 585
R1397 VDD.n6140 VDD.n6139 585
R1398 VDD.n6593 VDD.n6592 585
R1399 VDD.n6591 VDD.n6590 585
R1400 VDD.n6587 VDD.n6573 585
R1401 VDD.n6577 VDD.n6574 585
R1402 VDD.n6582 VDD.n6581 585
R1403 VDD.n6580 VDD.n6579 585
R1404 VDD.n6605 VDD.n6598 585
R1405 VDD.n6606 VDD.n6605 585
R1406 VDD.n6605 VDD.n6604 585
R1407 VDD.n6619 VDD.n6612 585
R1408 VDD.n6620 VDD.n6619 585
R1409 VDD.n6619 VDD.n6618 585
R1410 VDD.n6632 VDD.n6625 585
R1411 VDD.n6633 VDD.n6632 585
R1412 VDD.n6632 VDD.n6631 585
R1413 VDD.n6645 VDD.n6638 585
R1414 VDD.n6646 VDD.n6645 585
R1415 VDD.n6645 VDD.n6644 585
R1416 VDD.n6658 VDD.n6651 585
R1417 VDD.n6659 VDD.n6658 585
R1418 VDD.n6658 VDD.n6657 585
R1419 VDD.n6671 VDD.n6664 585
R1420 VDD.n6672 VDD.n6671 585
R1421 VDD.n6671 VDD.n6670 585
R1422 VDD.n6684 VDD.n6677 585
R1423 VDD.n6685 VDD.n6684 585
R1424 VDD.n6684 VDD.n6683 585
R1425 VDD.n6698 VDD.n6691 585
R1426 VDD.n6699 VDD.n6698 585
R1427 VDD.n6698 VDD.n6697 585
R1428 VDD.n6711 VDD.n6704 585
R1429 VDD.n6712 VDD.n6711 585
R1430 VDD.n6711 VDD.n6710 585
R1431 VDD.n6724 VDD.n6717 585
R1432 VDD.n6725 VDD.n6724 585
R1433 VDD.n6724 VDD.n6723 585
R1434 VDD.n6737 VDD.n6730 585
R1435 VDD.n6738 VDD.n6737 585
R1436 VDD.n6737 VDD.n6736 585
R1437 VDD.n6750 VDD.n6743 585
R1438 VDD.n6751 VDD.n6750 585
R1439 VDD.n6750 VDD.n6749 585
R1440 VDD.n6551 VDD.n6544 585
R1441 VDD.n6552 VDD.n6551 585
R1442 VDD.n6551 VDD.n6550 585
R1443 VDD.n6537 VDD.n6530 585
R1444 VDD.n6538 VDD.n6537 585
R1445 VDD.n6537 VDD.n6536 585
R1446 VDD.n6523 VDD.n6516 585
R1447 VDD.n6524 VDD.n6523 585
R1448 VDD.n6523 VDD.n6522 585
R1449 VDD.n6509 VDD.n6502 585
R1450 VDD.n6510 VDD.n6509 585
R1451 VDD.n6509 VDD.n6508 585
R1452 VDD.n6495 VDD.n6488 585
R1453 VDD.n6496 VDD.n6495 585
R1454 VDD.n6495 VDD.n6494 585
R1455 VDD.n6481 VDD.n6474 585
R1456 VDD.n6482 VDD.n6481 585
R1457 VDD.n6481 VDD.n6480 585
R1458 VDD.n6466 VDD.n6459 585
R1459 VDD.n6467 VDD.n6466 585
R1460 VDD.n6466 VDD.n6465 585
R1461 VDD.n6453 VDD.n6452 585
R1462 VDD.n6451 VDD.n6450 585
R1463 VDD.n6447 VDD.n6433 585
R1464 VDD.n6437 VDD.n6434 585
R1465 VDD.n6442 VDD.n6441 585
R1466 VDD.n6440 VDD.n6439 585
R1467 VDD.t575 VDD.t693 582.109
R1468 VDD.n2614 VDD.n2600 518.284
R1469 VDD.n2933 VDD.n2919 518.284
R1470 VDD.n20 VDD.n6 518.284
R1471 VDD.n339 VDD.n325 518.284
R1472 VDD.n5583 VDD.n5569 518.284
R1473 VDD.n5902 VDD.n5888 518.284
R1474 VDD.n2908 VDD.n2742 504.488
R1475 VDD.n2794 VDD.n2786 504.488
R1476 VDD.n314 VDD.n148 504.488
R1477 VDD.n200 VDD.n192 504.488
R1478 VDD.n5877 VDD.n5711 504.488
R1479 VDD.n5763 VDD.n5755 504.488
R1480 VDD.n2753 VDD.n2750 499.86
R1481 VDD.n2833 VDD.n2784 499.86
R1482 VDD.n159 VDD.n156 499.86
R1483 VDD.n239 VDD.n190 499.86
R1484 VDD.n5722 VDD.n5719 499.86
R1485 VDD.n5802 VDD.n5753 499.86
R1486 VDD.t581 VDD 488.971
R1487 VDD.n5427 VDD.t547 414.087
R1488 VDD.n5431 VDD.t151 405.404
R1489 VDD.t673 VDD.n5512 393.505
R1490 VDD.t345 VDD.n2605 384.339
R1491 VDD.t533 VDD.n2924 384.339
R1492 VDD.n3138 VDD.t449 384.339
R1493 VDD.n3188 VDD.t403 384.339
R1494 VDD.n3609 VDD.t624 384.339
R1495 VDD.n3469 VDD.t646 384.339
R1496 VDD.t125 VDD.n11 384.339
R1497 VDD.t124 VDD.n330 384.339
R1498 VDD.n544 VDD.t229 384.339
R1499 VDD.n594 VDD.t308 384.339
R1500 VDD.n1015 VDD.t517 384.339
R1501 VDD.n875 VDD.t80 384.339
R1502 VDD.t710 VDD.n5574 384.339
R1503 VDD.t698 VDD.n5893 384.339
R1504 VDD.n6107 VDD.t153 384.339
R1505 VDD.n6157 VDD.t680 384.339
R1506 VDD.n6578 VDD.t180 384.339
R1507 VDD.n6438 VDD.t256 384.339
R1508 VDD.n5228 VDD.n5198 375.954
R1509 VDD.n5287 VDD.n5286 375.954
R1510 VDD.n5425 VDD.n5424 372.646
R1511 VDD.n5384 VDD.n5383 372.646
R1512 VDD.n5382 VDD.n5381 372.646
R1513 VDD.n5360 VDD.n5359 371.964
R1514 VDD VDD.t70 371.557
R1515 VDD.n5559 VDD.n5558 371.195
R1516 VDD.n5536 VDD.n5535 371.195
R1517 VDD.n5491 VDD.n5486 371.195
R1518 VDD.n5512 VDD.n5511 370
R1519 VDD.n5514 VDD.n5513 370
R1520 VDD.n5538 VDD.n5537 370
R1521 VDD.n5561 VDD.n5560 370
R1522 VDD.n5362 VDD.n5361 370
R1523 VDD.n5404 VDD.n5403 370
R1524 VDD.n5406 VDD.n5405 370
R1525 VDD.n5423 VDD.n5422 370
R1526 VDD.n5243 VDD.n5190 369.93
R1527 VDD.n5295 VDD.n5294 369.93
R1528 VDD.n5404 VDD 367.334
R1529 VDD.n5213 VDD.n5202 359.529
R1530 VDD.n5209 VDD.n5202 359.529
R1531 VDD.n5273 VDD.n5262 359.529
R1532 VDD.n5269 VDD.n5262 359.529
R1533 VDD.n5488 VDD.t564 350.045
R1534 VDD.n5346 VDD.t119 350.043
R1535 VDD.n5445 VDD.t576 342.841
R1536 VDD.n5544 VDD.t582 342.841
R1537 VDD.n5481 VDD.t674 342.841
R1538 VDD.n5412 VDD.t71 342.839
R1539 VDD.n5391 VDD.t529 338.488
R1540 VDD.n5340 VDD.t556 338.488
R1541 VDD.n5452 VDD.n5448 320.976
R1542 VDD.n5562 VDD.n5443 320.976
R1543 VDD.n5552 VDD.n5551 320.976
R1544 VDD.n5464 VDD.n5463 320.976
R1545 VDD.n5467 VDD.n5466 320.976
R1546 VDD.n5529 VDD.n5528 320.976
R1547 VDD.n5472 VDD.n5471 320.976
R1548 VDD.n5520 VDD.n5474 320.976
R1549 VDD.n5479 VDD.n5478 320.976
R1550 VDD.n5505 VDD.n5504 320.976
R1551 VDD.n5499 VDD.n5483 320.976
R1552 VDD.n5493 VDD.n5492 320.976
R1553 VDD.n5489 VDD.n5487 320.976
R1554 VDD.n5330 VDD.n5329 320.976
R1555 VDD.n5345 VDD.n5344 320.976
R1556 VDD.n5313 VDD.n5312 320.976
R1557 VDD.n5315 VDD.n5314 320.976
R1558 VDD.n5319 VDD.n5318 320.976
R1559 VDD.n5322 VDD.n5321 320.976
R1560 VDD.n5327 VDD.n5326 320.976
R1561 VDD.n5397 VDD.n5396 320.976
R1562 VDD.n5335 VDD.n5334 320.976
R1563 VDD.n5368 VDD.n5337 320.976
R1564 VDD.n5371 VDD.n5370 320.976
R1565 VDD.n5343 VDD.n5342 320.976
R1566 VDD.n5353 VDD.n5349 320.976
R1567 VDD VDD.t150 299.068
R1568 VDD.n5237 VDD.n5236 297.036
R1569 VDD.n5300 VDD.n5299 297.036
R1570 VDD.t708 VDD 282.889
R1571 VDD.n5226 VDD.n5224 275.812
R1572 VDD.n5282 VDD.n5281 275.812
R1573 VDD.n5209 VDD.n5208 273.108
R1574 VDD.n5269 VDD.n5268 273.108
R1575 VDD.n5214 VDD.n5213 272.356
R1576 VDD.n5274 VDD.n5273 272.356
R1577 VDD.n5432 VDD.t686 249.901
R1578 VDD.n5411 VDD.t497 249.901
R1579 VDD.n5376 VDD.t459 249.901
R1580 VDD.n5339 VDD.t306 249.901
R1581 VDD.n5450 VDD.t696 248.843
R1582 VDD.n5390 VDD.t133 248.843
R1583 VDD.t150 VDD.t546 248.599
R1584 VDD.n5545 VDD.t311 245.636
R1585 VDD.n5522 VDD.t353 245.636
R1586 VDD.n5523 VDD.t188 245.636
R1587 VDD.n5480 VDD.t239 245.636
R1588 VDD.n2671 VDD.n2635 240
R1589 VDD.n2644 VDD.n2635 240
R1590 VDD.n3075 VDD.n2644 240
R1591 VDD.n3075 VDD.n2645 240
R1592 VDD.n3071 VDD.n2645 240
R1593 VDD.n3071 VDD.n2676 240
R1594 VDD.n3063 VDD.n2676 240
R1595 VDD.n3063 VDD.n2686 240
R1596 VDD.n3059 VDD.n2686 240
R1597 VDD.n3059 VDD.n2688 240
R1598 VDD.n3051 VDD.n2688 240
R1599 VDD.n3051 VDD.n2698 240
R1600 VDD.n3047 VDD.n2698 240
R1601 VDD.n3047 VDD.n2700 240
R1602 VDD.n3039 VDD.n2700 240
R1603 VDD.n3039 VDD.n2710 240
R1604 VDD.n3035 VDD.n2710 240
R1605 VDD.n3035 VDD.n2712 240
R1606 VDD.n3027 VDD.n2712 240
R1607 VDD.n3027 VDD.n2722 240
R1608 VDD.n3023 VDD.n2722 240
R1609 VDD.n3023 VDD.n2724 240
R1610 VDD.n3015 VDD.n2724 240
R1611 VDD.n2670 VDD.n2669 240
R1612 VDD.n2667 VDD.n2648 240
R1613 VDD.n2663 VDD.n2662 240
R1614 VDD.n2660 VDD.n2651 240
R1615 VDD.n2655 VDD.n2654 240
R1616 VDD.n3097 VDD.n3096 240
R1617 VDD.n3094 VDD.n2626 240
R1618 VDD.n3090 VDD.n3089 240
R1619 VDD.n3083 VDD.n2629 240
R1620 VDD.n3083 VDD.n2631 240
R1621 VDD.n2642 VDD.n2631 240
R1622 VDD.n2947 VDD.n2642 240
R1623 VDD.n2947 VDD.n2678 240
R1624 VDD.n2950 VDD.n2678 240
R1625 VDD.n2950 VDD.n2684 240
R1626 VDD.n2953 VDD.n2684 240
R1627 VDD.n2953 VDD.n2690 240
R1628 VDD.n2956 VDD.n2690 240
R1629 VDD.n2956 VDD.n2696 240
R1630 VDD.n2959 VDD.n2696 240
R1631 VDD.n2959 VDD.n2702 240
R1632 VDD.n2962 VDD.n2702 240
R1633 VDD.n2962 VDD.n2708 240
R1634 VDD.n2965 VDD.n2708 240
R1635 VDD.n2965 VDD.n2714 240
R1636 VDD.n2968 VDD.n2714 240
R1637 VDD.n2968 VDD.n2720 240
R1638 VDD.n2971 VDD.n2720 240
R1639 VDD.n2971 VDD.n2726 240
R1640 VDD.n2974 VDD.n2726 240
R1641 VDD.n2974 VDD.n2732 240
R1642 VDD.n3011 VDD.n3009 240
R1643 VDD.n3007 VDD.n2736 240
R1644 VDD.n3003 VDD.n3001 240
R1645 VDD.n2999 VDD.n2738 240
R1646 VDD.n2992 VDD.n2990 240
R1647 VDD.n2987 VDD.n2986 240
R1648 VDD.n2984 VDD.n2945 240
R1649 VDD.n2980 VDD.n2978 240
R1650 VDD.n3081 VDD.n2636 240
R1651 VDD.n3081 VDD.n2637 240
R1652 VDD.n3077 VDD.n2637 240
R1653 VDD.n3077 VDD.n2640 240
R1654 VDD.n3069 VDD.n2640 240
R1655 VDD.n3069 VDD.n2679 240
R1656 VDD.n3065 VDD.n2679 240
R1657 VDD.n3065 VDD.n2681 240
R1658 VDD.n3057 VDD.n2681 240
R1659 VDD.n3057 VDD.n2691 240
R1660 VDD.n3053 VDD.n2691 240
R1661 VDD.n3053 VDD.n2693 240
R1662 VDD.n3045 VDD.n2693 240
R1663 VDD.n3045 VDD.n2703 240
R1664 VDD.n3041 VDD.n2703 240
R1665 VDD.n3041 VDD.n2705 240
R1666 VDD.n3033 VDD.n2705 240
R1667 VDD.n3033 VDD.n2715 240
R1668 VDD.n3029 VDD.n2715 240
R1669 VDD.n3029 VDD.n2717 240
R1670 VDD.n3021 VDD.n2717 240
R1671 VDD.n3021 VDD.n2728 240
R1672 VDD.n3017 VDD.n2728 240
R1673 VDD.n2760 VDD.n2758 240
R1674 VDD.n2764 VDD.n2758 240
R1675 VDD.n2768 VDD.n2766 240
R1676 VDD.n2772 VDD.n2756 240
R1677 VDD.n2900 VDD.n2774 240
R1678 VDD.n2898 VDD.n2775 240
R1679 VDD.n2894 VDD.n2892 240
R1680 VDD.n2890 VDD.n2777 240
R1681 VDD.n2849 VDD.n2633 240
R1682 VDD.n2852 VDD.n2633 240
R1683 VDD.n2852 VDD.n2641 240
R1684 VDD.n2855 VDD.n2641 240
R1685 VDD.n2855 VDD.n2677 240
R1686 VDD.n2858 VDD.n2677 240
R1687 VDD.n2858 VDD.n2683 240
R1688 VDD.n2861 VDD.n2683 240
R1689 VDD.n2861 VDD.n2689 240
R1690 VDD.n2864 VDD.n2689 240
R1691 VDD.n2864 VDD.n2695 240
R1692 VDD.n2867 VDD.n2695 240
R1693 VDD.n2867 VDD.n2701 240
R1694 VDD.n2870 VDD.n2701 240
R1695 VDD.n2870 VDD.n2707 240
R1696 VDD.n2873 VDD.n2707 240
R1697 VDD.n2873 VDD.n2713 240
R1698 VDD.n2876 VDD.n2713 240
R1699 VDD.n2876 VDD.n2719 240
R1700 VDD.n2879 VDD.n2719 240
R1701 VDD.n2879 VDD.n2725 240
R1702 VDD.n2882 VDD.n2725 240
R1703 VDD.n2882 VDD.n2731 240
R1704 VDD.n2807 VDD.n2805 240
R1705 VDD.n2811 VDD.n2800 240
R1706 VDD.n2814 VDD.n2813 240
R1707 VDD.n2815 VDD.n2814 240
R1708 VDD.n2821 VDD.n2819 240
R1709 VDD.n2838 VDD.n2781 240
R1710 VDD.n2842 VDD.n2840 240
R1711 VDD.n2846 VDD.n2779 240
R1712 VDD.n4387 VDD.n4120 240
R1713 VDD.n4466 VDD.n4120 240
R1714 VDD.n4466 VDD.n4117 240
R1715 VDD.n4471 VDD.n4117 240
R1716 VDD.n4471 VDD.n4118 240
R1717 VDD.n4118 VDD.n4093 240
R1718 VDD.n4500 VDD.n4093 240
R1719 VDD.n4500 VDD.n4090 240
R1720 VDD.n4505 VDD.n4090 240
R1721 VDD.n4505 VDD.n4091 240
R1722 VDD.n4091 VDD.n4068 240
R1723 VDD.n4535 VDD.n4068 240
R1724 VDD.n4535 VDD.n3442 240
R1725 VDD.n5155 VDD.n3442 240
R1726 VDD.n5155 VDD.n3443 240
R1727 VDD.n4550 VDD.n3443 240
R1728 VDD.n4576 VDD.n4550 240
R1729 VDD.n4576 VDD.n4030 240
R1730 VDD.n4618 VDD.n4030 240
R1731 VDD.n4618 VDD.n4031 240
R1732 VDD.n4031 VDD.n4005 240
R1733 VDD.n4653 VDD.n4005 240
R1734 VDD.n4653 VDD.n3996 240
R1735 VDD.n4670 VDD.n3996 240
R1736 VDD.n4670 VDD.n3997 240
R1737 VDD.n3997 VDD.n3967 240
R1738 VDD.n4697 VDD.n3967 240
R1739 VDD.n4697 VDD.n3968 240
R1740 VDD.n3968 VDD.n3936 240
R1741 VDD.n4724 VDD.n3936 240
R1742 VDD.n4724 VDD.n3937 240
R1743 VDD.n3937 VDD.n3800 240
R1744 VDD.n5132 VDD.n3800 240
R1745 VDD.n5132 VDD.n3801 240
R1746 VDD.n4756 VDD.n3801 240
R1747 VDD.n4756 VDD.n3821 240
R1748 VDD.n5113 VDD.n3821 240
R1749 VDD.n5113 VDD.n3822 240
R1750 VDD.n5109 VDD.n3822 240
R1751 VDD.n5109 VDD.n3825 240
R1752 VDD.n3862 VDD.n3825 240
R1753 VDD.n3862 VDD.n3860 240
R1754 VDD.n5090 VDD.n3860 240
R1755 VDD.n5090 VDD.n3861 240
R1756 VDD.n5086 VDD.n3861 240
R1757 VDD.n5086 VDD.n3866 240
R1758 VDD.n5078 VDD.n3866 240
R1759 VDD.n5078 VDD.n3883 240
R1760 VDD.n5074 VDD.n3883 240
R1761 VDD.n4422 VDD.n4388 240
R1762 VDD.n4418 VDD.n4417 240
R1763 VDD.n4414 VDD.n4413 240
R1764 VDD.n4410 VDD.n4409 240
R1765 VDD.n4406 VDD.n4405 240
R1766 VDD.n4402 VDD.n4401 240
R1767 VDD.n4398 VDD.n4397 240
R1768 VDD.n4394 VDD.n4393 240
R1769 VDD.n4432 VDD.n4137 240
R1770 VDD.n4432 VDD.n4122 240
R1771 VDD.n4437 VDD.n4122 240
R1772 VDD.n4437 VDD.n4115 240
R1773 VDD.n4115 VDD.n4109 240
R1774 VDD.n4479 VDD.n4109 240
R1775 VDD.n4479 VDD.n4095 240
R1776 VDD.n4483 VDD.n4095 240
R1777 VDD.n4483 VDD.n4087 240
R1778 VDD.n4492 VDD.n4087 240
R1779 VDD.n4492 VDD.n4103 240
R1780 VDD.n4103 VDD.n4067 240
R1781 VDD.n4067 VDD.n3438 240
R1782 VDD.n5157 VDD.n3438 240
R1783 VDD.n5157 VDD.n3439 240
R1784 VDD.n4056 VDD.n3439 240
R1785 VDD.n4578 VDD.n4056 240
R1786 VDD.n4578 VDD.n4051 240
R1787 VDD.n4051 VDD.n4028 240
R1788 VDD.n4028 VDD.n4022 240
R1789 VDD.n4625 VDD.n4022 240
R1790 VDD.n4625 VDD.n4007 240
R1791 VDD.n4638 VDD.n4007 240
R1792 VDD.n4638 VDD.n3993 240
R1793 VDD.n4018 VDD.n3993 240
R1794 VDD.n4633 VDD.n4018 240
R1795 VDD.n4633 VDD.n3965 240
R1796 VDD.n4630 VDD.n3965 240
R1797 VDD.n4630 VDD.n3960 240
R1798 VDD.n3960 VDD.n3934 240
R1799 VDD.n3951 VDD.n3934 240
R1800 VDD.n3951 VDD.n3928 240
R1801 VDD.n3928 VDD.n3797 240
R1802 VDD.n4740 VDD.n3797 240
R1803 VDD.n4741 VDD.n4740 240
R1804 VDD.n4741 VDD.n3921 240
R1805 VDD.n3921 VDD.n3818 240
R1806 VDD.n4977 VDD.n3818 240
R1807 VDD.n4977 VDD.n3827 240
R1808 VDD.n5103 VDD.n3827 240
R1809 VDD.n5103 VDD.n3834 240
R1810 VDD.n3914 VDD.n3834 240
R1811 VDD.n3914 VDD.n3857 240
R1812 VDD.n4991 VDD.n3857 240
R1813 VDD.n4991 VDD.n3868 240
R1814 VDD.n4995 VDD.n3868 240
R1815 VDD.n4995 VDD.n3881 240
R1816 VDD.n5031 VDD.n3881 240
R1817 VDD.n5031 VDD.n3887 240
R1818 VDD.n5064 VDD.n3909 240
R1819 VDD.n5060 VDD.n3909 240
R1820 VDD.n5058 VDD.n5057 240
R1821 VDD.n5054 VDD.n5053 240
R1822 VDD.n5050 VDD.n5049 240
R1823 VDD.n5046 VDD.n5045 240
R1824 VDD.n5042 VDD.n5041 240
R1825 VDD.n5038 VDD.n5037 240
R1826 VDD.n4385 VDD.n4124 240
R1827 VDD.n4464 VDD.n4124 240
R1828 VDD.n4464 VDD.n4125 240
R1829 VDD.n4125 VDD.n4116 240
R1830 VDD.n4459 VDD.n4116 240
R1831 VDD.n4459 VDD.n4097 240
R1832 VDD.n4498 VDD.n4097 240
R1833 VDD.n4498 VDD.n4098 240
R1834 VDD.n4098 VDD.n4089 240
R1835 VDD.n4101 VDD.n4089 240
R1836 VDD.n4101 VDD.n4064 240
R1837 VDD.n4537 VDD.n4064 240
R1838 VDD.n4538 VDD.n4537 240
R1839 VDD.n4538 VDD.n3436 240
R1840 VDD.n4547 VDD.n3436 240
R1841 VDD.n4548 VDD.n4547 240
R1842 VDD.n4548 VDD.n4052 240
R1843 VDD.n4585 VDD.n4052 240
R1844 VDD.n4585 VDD.n4029 240
R1845 VDD.n4581 VDD.n4029 240
R1846 VDD.n4581 VDD.n4009 240
R1847 VDD.n4651 VDD.n4009 240
R1848 VDD.n4651 VDD.n4010 240
R1849 VDD.n4010 VDD.n3995 240
R1850 VDD.n4646 VDD.n3995 240
R1851 VDD.n4646 VDD.n4016 240
R1852 VDD.n4016 VDD.n3966 240
R1853 VDD.n4012 VDD.n3966 240
R1854 VDD.n4012 VDD.n3932 240
R1855 VDD.n4726 VDD.n3932 240
R1856 VDD.n4726 VDD.n3929 240
R1857 VDD.n4732 VDD.n3929 240
R1858 VDD.n4732 VDD.n3799 240
R1859 VDD.n3922 VDD.n3799 240
R1860 VDD.n4743 VDD.n3922 240
R1861 VDD.n4746 VDD.n4743 240
R1862 VDD.n4746 VDD.n3820 240
R1863 VDD.n3829 VDD.n3820 240
R1864 VDD.n5107 VDD.n3829 240
R1865 VDD.n5107 VDD.n3830 240
R1866 VDD.n3873 VDD.n3830 240
R1867 VDD.n3874 VDD.n3873 240
R1868 VDD.n3874 VDD.n3859 240
R1869 VDD.n3870 VDD.n3859 240
R1870 VDD.n5084 VDD.n3870 240
R1871 VDD.n5084 VDD.n3871 240
R1872 VDD.n5080 VDD.n3871 240
R1873 VDD.n5080 VDD.n3879 240
R1874 VDD.n5072 VDD.n3879 240
R1875 VDD.n4381 VDD.n4143 240
R1876 VDD.n4379 VDD.n4378 240
R1877 VDD.n4375 VDD.n4374 240
R1878 VDD.n4371 VDD.n4370 240
R1879 VDD.n4367 VDD.n4366 240
R1880 VDD.n4363 VDD.n4362 240
R1881 VDD.n4359 VDD.n4358 240
R1882 VDD.n4355 VDD.n4141 240
R1883 VDD.n4430 VDD.n4139 240
R1884 VDD.n4430 VDD.n4123 240
R1885 VDD.n4123 VDD.n4113 240
R1886 VDD.n4473 VDD.n4113 240
R1887 VDD.n4473 VDD.n4111 240
R1888 VDD.n4477 VDD.n4111 240
R1889 VDD.n4477 VDD.n4096 240
R1890 VDD.n4485 VDD.n4096 240
R1891 VDD.n4485 VDD.n4088 240
R1892 VDD.n4490 VDD.n4088 240
R1893 VDD.n4490 VDD.n4105 240
R1894 VDD.n4105 VDD.n4062 240
R1895 VDD.n4540 VDD.n4062 240
R1896 VDD.n4540 VDD.n3441 240
R1897 VDD.n4060 VDD.n3441 240
R1898 VDD.n4546 VDD.n4060 240
R1899 VDD.n4546 VDD.n4058 240
R1900 VDD.n4058 VDD.n4026 240
R1901 VDD.n4620 VDD.n4026 240
R1902 VDD.n4620 VDD.n4024 240
R1903 VDD.n4624 VDD.n4024 240
R1904 VDD.n4624 VDD.n4008 240
R1905 VDD.n4640 VDD.n4008 240
R1906 VDD.n4640 VDD.n3994 240
R1907 VDD.n4644 VDD.n3994 240
R1908 VDD.n4644 VDD.n3963 240
R1909 VDD.n4699 VDD.n3963 240
R1910 VDD.n4699 VDD.n3961 240
R1911 VDD.n4704 VDD.n3961 240
R1912 VDD.n4704 VDD.n3935 240
R1913 VDD.n3935 VDD.n3926 240
R1914 VDD.n4734 VDD.n3926 240
R1915 VDD.n4734 VDD.n3798 240
R1916 VDD.n4738 VDD.n3798 240
R1917 VDD.n4738 VDD.n3919 240
R1918 VDD.n4748 VDD.n3919 240
R1919 VDD.n4748 VDD.n3819 240
R1920 VDD.n4979 VDD.n3819 240
R1921 VDD.n4979 VDD.n3828 240
R1922 VDD.n3836 VDD.n3828 240
R1923 VDD.n4984 VDD.n3836 240
R1924 VDD.n4985 VDD.n4984 240
R1925 VDD.n4985 VDD.n3858 240
R1926 VDD.n4989 VDD.n3858 240
R1927 VDD.n4989 VDD.n3869 240
R1928 VDD.n4997 VDD.n3869 240
R1929 VDD.n4997 VDD.n3882 240
R1930 VDD.n5029 VDD.n3882 240
R1931 VDD.n5029 VDD.n3888 240
R1932 VDD.n5068 VDD.n3892 240
R1933 VDD.n5002 VDD.n5001 240
R1934 VDD.n5006 VDD.n5005 240
R1935 VDD.n5010 VDD.n5009 240
R1936 VDD.n5014 VDD.n5013 240
R1937 VDD.n5018 VDD.n5017 240
R1938 VDD.n5022 VDD.n5021 240
R1939 VDD.n5024 VDD.n3907 240
R1940 VDD.n4247 VDD.n4201 240
R1941 VDD.n4247 VDD.n4195 240
R1942 VDD.n4255 VDD.n4195 240
R1943 VDD.n4255 VDD.n4193 240
R1944 VDD.n4259 VDD.n4193 240
R1945 VDD.n4259 VDD.n4187 240
R1946 VDD.n4268 VDD.n4187 240
R1947 VDD.n4268 VDD.n4185 240
R1948 VDD.n4272 VDD.n4185 240
R1949 VDD.n4272 VDD.n4180 240
R1950 VDD.n4281 VDD.n4180 240
R1951 VDD.n4281 VDD.n4178 240
R1952 VDD.n4285 VDD.n4178 240
R1953 VDD.n4285 VDD.n4173 240
R1954 VDD.n4293 VDD.n4173 240
R1955 VDD.n4293 VDD.n4171 240
R1956 VDD.n4298 VDD.n4171 240
R1957 VDD.n4298 VDD.n4164 240
R1958 VDD.n4345 VDD.n4164 240
R1959 VDD.n4346 VDD.n4345 240
R1960 VDD.n4346 VDD.n4161 240
R1961 VDD.n4353 VDD.n4161 240
R1962 VDD.n4353 VDD.n4162 240
R1963 VDD.n4162 VDD.n4134 240
R1964 VDD.n4440 VDD.n4134 240
R1965 VDD.n4440 VDD.n4128 240
R1966 VDD.n4456 VDD.n4128 240
R1967 VDD.n4456 VDD.n4129 240
R1968 VDD.n4449 VDD.n4129 240
R1969 VDD.n4449 VDD.n4085 240
R1970 VDD.n4508 VDD.n4085 240
R1971 VDD.n4508 VDD.n4079 240
R1972 VDD.n4524 VDD.n4079 240
R1973 VDD.n4524 VDD.n4080 240
R1974 VDD.n4517 VDD.n4080 240
R1975 VDD.n4517 VDD.n3453 240
R1976 VDD.n5146 VDD.n3453 240
R1977 VDD.n5146 VDD.n3454 240
R1978 VDD.n4049 VDD.n3454 240
R1979 VDD.n4588 VDD.n4049 240
R1980 VDD.n4588 VDD.n4044 240
R1981 VDD.n4604 VDD.n4044 240
R1982 VDD.n4604 VDD.n4045 240
R1983 VDD.n4597 VDD.n4045 240
R1984 VDD.n4597 VDD.n3991 240
R1985 VDD.n4673 VDD.n3991 240
R1986 VDD.n4673 VDD.n3985 240
R1987 VDD.n4685 VDD.n3985 240
R1988 VDD.n4685 VDD.n3986 240
R1989 VDD.n3986 VDD.n3957 240
R1990 VDD.n4707 VDD.n3957 240
R1991 VDD.n4707 VDD.n3953 240
R1992 VDD.n4715 VDD.n3953 240
R1993 VDD.n4715 VDD.n3794 240
R1994 VDD.n5135 VDD.n3794 240
R1995 VDD.n5135 VDD.n3795 240
R1996 VDD.n5123 VDD.n3795 240
R1997 VDD.n5123 VDD.n3811 240
R1998 VDD.n5116 VDD.n3811 240
R1999 VDD.n5116 VDD.n3816 240
R2000 VDD.n3846 VDD.n3816 240
R2001 VDD.n3846 VDD.n3839 240
R2002 VDD.n5100 VDD.n3839 240
R2003 VDD.n5100 VDD.n3840 240
R2004 VDD.n5093 VDD.n3840 240
R2005 VDD.n5093 VDD.n3854 240
R2006 VDD.n4793 VDD.n3854 240
R2007 VDD.n4794 VDD.n4793 240
R2008 VDD.n4794 VDD.n4785 240
R2009 VDD.n4800 VDD.n4785 240
R2010 VDD.n4801 VDD.n4800 240
R2011 VDD.n4802 VDD.n4801 240
R2012 VDD.n4802 VDD.n4782 240
R2013 VDD.n4941 VDD.n4782 240
R2014 VDD.n4941 VDD.n4783 240
R2015 VDD.n4937 VDD.n4783 240
R2016 VDD.n4937 VDD.n4806 240
R2017 VDD.n4933 VDD.n4806 240
R2018 VDD.n4933 VDD.n4811 240
R2019 VDD.n4929 VDD.n4811 240
R2020 VDD.n4929 VDD.n4813 240
R2021 VDD.n4925 VDD.n4813 240
R2022 VDD.n4925 VDD.n4817 240
R2023 VDD.n4921 VDD.n4817 240
R2024 VDD.n4921 VDD.n4819 240
R2025 VDD.n4917 VDD.n4819 240
R2026 VDD.n4917 VDD.n4825 240
R2027 VDD.n4913 VDD.n4825 240
R2028 VDD.n4913 VDD.n4827 240
R2029 VDD.n4909 VDD.n4827 240
R2030 VDD.n4909 VDD.n4832 240
R2031 VDD.n4905 VDD.n4832 240
R2032 VDD.n4905 VDD.n4834 240
R2033 VDD.n4845 VDD.n4844 240
R2034 VDD.n4895 VDD.n4844 240
R2035 VDD.n4893 VDD.n4892 240
R2036 VDD.n4889 VDD.n4888 240
R2037 VDD.n4885 VDD.n4884 240
R2038 VDD.n4881 VDD.n4880 240
R2039 VDD.n4877 VDD.n4876 240
R2040 VDD.n4873 VDD.n4872 240
R2041 VDD.n4249 VDD.n4199 240
R2042 VDD.n4249 VDD.n4197 240
R2043 VDD.n4253 VDD.n4197 240
R2044 VDD.n4253 VDD.n4191 240
R2045 VDD.n4261 VDD.n4191 240
R2046 VDD.n4261 VDD.n4189 240
R2047 VDD.n4265 VDD.n4189 240
R2048 VDD.n4265 VDD.n4183 240
R2049 VDD.n4274 VDD.n4183 240
R2050 VDD.n4274 VDD.n4181 240
R2051 VDD.n4278 VDD.n4181 240
R2052 VDD.n4278 VDD.n4177 240
R2053 VDD.n4287 VDD.n4177 240
R2054 VDD.n4287 VDD.n4175 240
R2055 VDD.n4291 VDD.n4175 240
R2056 VDD.n4291 VDD.n4169 240
R2057 VDD.n4300 VDD.n4169 240
R2058 VDD.n4300 VDD.n4166 240
R2059 VDD.n4343 VDD.n4166 240
R2060 VDD.n4343 VDD.n4167 240
R2061 VDD.n4339 VDD.n4167 240
R2062 VDD.n4339 VDD.n4160 240
R2063 VDD.n4336 VDD.n4160 240
R2064 VDD.n4336 VDD.n4335 240
R2065 VDD.n4335 VDD.n4135 240
R2066 VDD.n4328 VDD.n4135 240
R2067 VDD.n4328 VDD.n4127 240
R2068 VDD.n4309 VDD.n4127 240
R2069 VDD.n4320 VDD.n4309 240
R2070 VDD.n4320 VDD.n4319 240
R2071 VDD.n4319 VDD.n4086 240
R2072 VDD.n4086 VDD.n4075 240
R2073 VDD.n4526 VDD.n4075 240
R2074 VDD.n4527 VDD.n4526 240
R2075 VDD.n4528 VDD.n4527 240
R2076 VDD.n4528 VDD.n3450 240
R2077 VDD.n5148 VDD.n3450 240
R2078 VDD.n5148 VDD.n3451 240
R2079 VDD.n4565 VDD.n3451 240
R2080 VDD.n4565 VDD.n4050 240
R2081 VDD.n4050 VDD.n4042 240
R2082 VDD.n4606 VDD.n4042 240
R2083 VDD.n4611 VDD.n4606 240
R2084 VDD.n4611 VDD.n4610 240
R2085 VDD.n4610 VDD.n4607 240
R2086 VDD.n4607 VDD.n3992 240
R2087 VDD.n3992 VDD.n3981 240
R2088 VDD.n4687 VDD.n3981 240
R2089 VDD.n4688 VDD.n4687 240
R2090 VDD.n4690 VDD.n4688 240
R2091 VDD.n4690 VDD.n3959 240
R2092 VDD.n3959 VDD.n3946 240
R2093 VDD.n4717 VDD.n3946 240
R2094 VDD.n4717 VDD.n3950 240
R2095 VDD.n3950 VDD.n3796 240
R2096 VDD.n3808 VDD.n3796 240
R2097 VDD.n5125 VDD.n3808 240
R2098 VDD.n5125 VDD.n3809 240
R2099 VDD.n3817 VDD.n3809 240
R2100 VDD.n4975 VDD.n3817 240
R2101 VDD.n4975 VDD.n4751 240
R2102 VDD.n4968 VDD.n4751 240
R2103 VDD.n4968 VDD.n3837 240
R2104 VDD.n4769 VDD.n3837 240
R2105 VDD.n4769 VDD.n3856 240
R2106 VDD.n4958 VDD.n3856 240
R2107 VDD.n4958 VDD.n4957 240
R2108 VDD.n4957 VDD.n4773 240
R2109 VDD.n4950 VDD.n4773 240
R2110 VDD.n4950 VDD.n4949 240
R2111 VDD.n4949 VDD.n4777 240
R2112 VDD.n4945 VDD.n4777 240
R2113 VDD.n4945 VDD.n4944 240
R2114 VDD.n4944 VDD.n4943 240
R2115 VDD.n4943 VDD.n4779 240
R2116 VDD.n4807 VDD.n4779 240
R2117 VDD.n4808 VDD.n4807 240
R2118 VDD.n4809 VDD.n4808 240
R2119 VDD.n4850 VDD.n4809 240
R2120 VDD.n4850 VDD.n4814 240
R2121 VDD.n4815 VDD.n4814 240
R2122 VDD.n4816 VDD.n4815 240
R2123 VDD.n4855 VDD.n4816 240
R2124 VDD.n4855 VDD.n4821 240
R2125 VDD.n4822 VDD.n4821 240
R2126 VDD.n4823 VDD.n4822 240
R2127 VDD.n4860 VDD.n4823 240
R2128 VDD.n4860 VDD.n4828 240
R2129 VDD.n4829 VDD.n4828 240
R2130 VDD.n4830 VDD.n4829 240
R2131 VDD.n4865 VDD.n4830 240
R2132 VDD.n4865 VDD.n4835 240
R2133 VDD.n4836 VDD.n4835 240
R2134 VDD.n4212 VDD.n4203 240
R2135 VDD.n4216 VDD.n4215 240
R2136 VDD.n4220 VDD.n4219 240
R2137 VDD.n4224 VDD.n4223 240
R2138 VDD.n4228 VDD.n4227 240
R2139 VDD.n4232 VDD.n4231 240
R2140 VDD.n4236 VDD.n4235 240
R2141 VDD.n4240 VDD.n4211 240
R2142 VDD.n77 VDD.n41 240
R2143 VDD.n50 VDD.n41 240
R2144 VDD.n481 VDD.n50 240
R2145 VDD.n481 VDD.n51 240
R2146 VDD.n477 VDD.n51 240
R2147 VDD.n477 VDD.n82 240
R2148 VDD.n469 VDD.n82 240
R2149 VDD.n469 VDD.n92 240
R2150 VDD.n465 VDD.n92 240
R2151 VDD.n465 VDD.n94 240
R2152 VDD.n457 VDD.n94 240
R2153 VDD.n457 VDD.n104 240
R2154 VDD.n453 VDD.n104 240
R2155 VDD.n453 VDD.n106 240
R2156 VDD.n445 VDD.n106 240
R2157 VDD.n445 VDD.n116 240
R2158 VDD.n441 VDD.n116 240
R2159 VDD.n441 VDD.n118 240
R2160 VDD.n433 VDD.n118 240
R2161 VDD.n433 VDD.n128 240
R2162 VDD.n429 VDD.n128 240
R2163 VDD.n429 VDD.n130 240
R2164 VDD.n421 VDD.n130 240
R2165 VDD.n76 VDD.n75 240
R2166 VDD.n73 VDD.n54 240
R2167 VDD.n69 VDD.n68 240
R2168 VDD.n66 VDD.n57 240
R2169 VDD.n61 VDD.n60 240
R2170 VDD.n503 VDD.n502 240
R2171 VDD.n500 VDD.n32 240
R2172 VDD.n496 VDD.n495 240
R2173 VDD.n489 VDD.n35 240
R2174 VDD.n489 VDD.n37 240
R2175 VDD.n48 VDD.n37 240
R2176 VDD.n353 VDD.n48 240
R2177 VDD.n353 VDD.n84 240
R2178 VDD.n356 VDD.n84 240
R2179 VDD.n356 VDD.n90 240
R2180 VDD.n359 VDD.n90 240
R2181 VDD.n359 VDD.n96 240
R2182 VDD.n362 VDD.n96 240
R2183 VDD.n362 VDD.n102 240
R2184 VDD.n365 VDD.n102 240
R2185 VDD.n365 VDD.n108 240
R2186 VDD.n368 VDD.n108 240
R2187 VDD.n368 VDD.n114 240
R2188 VDD.n371 VDD.n114 240
R2189 VDD.n371 VDD.n120 240
R2190 VDD.n374 VDD.n120 240
R2191 VDD.n374 VDD.n126 240
R2192 VDD.n377 VDD.n126 240
R2193 VDD.n377 VDD.n132 240
R2194 VDD.n380 VDD.n132 240
R2195 VDD.n380 VDD.n138 240
R2196 VDD.n417 VDD.n415 240
R2197 VDD.n413 VDD.n142 240
R2198 VDD.n409 VDD.n407 240
R2199 VDD.n405 VDD.n144 240
R2200 VDD.n398 VDD.n396 240
R2201 VDD.n393 VDD.n392 240
R2202 VDD.n390 VDD.n351 240
R2203 VDD.n386 VDD.n384 240
R2204 VDD.n487 VDD.n42 240
R2205 VDD.n487 VDD.n43 240
R2206 VDD.n483 VDD.n43 240
R2207 VDD.n483 VDD.n46 240
R2208 VDD.n475 VDD.n46 240
R2209 VDD.n475 VDD.n85 240
R2210 VDD.n471 VDD.n85 240
R2211 VDD.n471 VDD.n87 240
R2212 VDD.n463 VDD.n87 240
R2213 VDD.n463 VDD.n97 240
R2214 VDD.n459 VDD.n97 240
R2215 VDD.n459 VDD.n99 240
R2216 VDD.n451 VDD.n99 240
R2217 VDD.n451 VDD.n109 240
R2218 VDD.n447 VDD.n109 240
R2219 VDD.n447 VDD.n111 240
R2220 VDD.n439 VDD.n111 240
R2221 VDD.n439 VDD.n121 240
R2222 VDD.n435 VDD.n121 240
R2223 VDD.n435 VDD.n123 240
R2224 VDD.n427 VDD.n123 240
R2225 VDD.n427 VDD.n134 240
R2226 VDD.n423 VDD.n134 240
R2227 VDD.n166 VDD.n164 240
R2228 VDD.n170 VDD.n164 240
R2229 VDD.n174 VDD.n172 240
R2230 VDD.n178 VDD.n162 240
R2231 VDD.n306 VDD.n180 240
R2232 VDD.n304 VDD.n181 240
R2233 VDD.n300 VDD.n298 240
R2234 VDD.n296 VDD.n183 240
R2235 VDD.n255 VDD.n39 240
R2236 VDD.n258 VDD.n39 240
R2237 VDD.n258 VDD.n47 240
R2238 VDD.n261 VDD.n47 240
R2239 VDD.n261 VDD.n83 240
R2240 VDD.n264 VDD.n83 240
R2241 VDD.n264 VDD.n89 240
R2242 VDD.n267 VDD.n89 240
R2243 VDD.n267 VDD.n95 240
R2244 VDD.n270 VDD.n95 240
R2245 VDD.n270 VDD.n101 240
R2246 VDD.n273 VDD.n101 240
R2247 VDD.n273 VDD.n107 240
R2248 VDD.n276 VDD.n107 240
R2249 VDD.n276 VDD.n113 240
R2250 VDD.n279 VDD.n113 240
R2251 VDD.n279 VDD.n119 240
R2252 VDD.n282 VDD.n119 240
R2253 VDD.n282 VDD.n125 240
R2254 VDD.n285 VDD.n125 240
R2255 VDD.n285 VDD.n131 240
R2256 VDD.n288 VDD.n131 240
R2257 VDD.n288 VDD.n137 240
R2258 VDD.n213 VDD.n211 240
R2259 VDD.n217 VDD.n206 240
R2260 VDD.n220 VDD.n219 240
R2261 VDD.n221 VDD.n220 240
R2262 VDD.n227 VDD.n225 240
R2263 VDD.n244 VDD.n187 240
R2264 VDD.n248 VDD.n246 240
R2265 VDD.n252 VDD.n185 240
R2266 VDD.n1793 VDD.n1526 240
R2267 VDD.n1872 VDD.n1526 240
R2268 VDD.n1872 VDD.n1523 240
R2269 VDD.n1877 VDD.n1523 240
R2270 VDD.n1877 VDD.n1524 240
R2271 VDD.n1524 VDD.n1499 240
R2272 VDD.n1906 VDD.n1499 240
R2273 VDD.n1906 VDD.n1496 240
R2274 VDD.n1911 VDD.n1496 240
R2275 VDD.n1911 VDD.n1497 240
R2276 VDD.n1497 VDD.n1474 240
R2277 VDD.n1941 VDD.n1474 240
R2278 VDD.n1941 VDD.n848 240
R2279 VDD.n2561 VDD.n848 240
R2280 VDD.n2561 VDD.n849 240
R2281 VDD.n1956 VDD.n849 240
R2282 VDD.n1982 VDD.n1956 240
R2283 VDD.n1982 VDD.n1436 240
R2284 VDD.n2024 VDD.n1436 240
R2285 VDD.n2024 VDD.n1437 240
R2286 VDD.n1437 VDD.n1411 240
R2287 VDD.n2059 VDD.n1411 240
R2288 VDD.n2059 VDD.n1402 240
R2289 VDD.n2076 VDD.n1402 240
R2290 VDD.n2076 VDD.n1403 240
R2291 VDD.n1403 VDD.n1373 240
R2292 VDD.n2103 VDD.n1373 240
R2293 VDD.n2103 VDD.n1374 240
R2294 VDD.n1374 VDD.n1342 240
R2295 VDD.n2130 VDD.n1342 240
R2296 VDD.n2130 VDD.n1343 240
R2297 VDD.n1343 VDD.n1206 240
R2298 VDD.n2538 VDD.n1206 240
R2299 VDD.n2538 VDD.n1207 240
R2300 VDD.n2162 VDD.n1207 240
R2301 VDD.n2162 VDD.n1227 240
R2302 VDD.n2519 VDD.n1227 240
R2303 VDD.n2519 VDD.n1228 240
R2304 VDD.n2515 VDD.n1228 240
R2305 VDD.n2515 VDD.n1231 240
R2306 VDD.n1268 VDD.n1231 240
R2307 VDD.n1268 VDD.n1266 240
R2308 VDD.n2496 VDD.n1266 240
R2309 VDD.n2496 VDD.n1267 240
R2310 VDD.n2492 VDD.n1267 240
R2311 VDD.n2492 VDD.n1272 240
R2312 VDD.n2484 VDD.n1272 240
R2313 VDD.n2484 VDD.n1289 240
R2314 VDD.n2480 VDD.n1289 240
R2315 VDD.n1828 VDD.n1794 240
R2316 VDD.n1824 VDD.n1823 240
R2317 VDD.n1820 VDD.n1819 240
R2318 VDD.n1816 VDD.n1815 240
R2319 VDD.n1812 VDD.n1811 240
R2320 VDD.n1808 VDD.n1807 240
R2321 VDD.n1804 VDD.n1803 240
R2322 VDD.n1800 VDD.n1799 240
R2323 VDD.n1838 VDD.n1543 240
R2324 VDD.n1838 VDD.n1528 240
R2325 VDD.n1843 VDD.n1528 240
R2326 VDD.n1843 VDD.n1521 240
R2327 VDD.n1521 VDD.n1515 240
R2328 VDD.n1885 VDD.n1515 240
R2329 VDD.n1885 VDD.n1501 240
R2330 VDD.n1889 VDD.n1501 240
R2331 VDD.n1889 VDD.n1493 240
R2332 VDD.n1898 VDD.n1493 240
R2333 VDD.n1898 VDD.n1509 240
R2334 VDD.n1509 VDD.n1473 240
R2335 VDD.n1473 VDD.n844 240
R2336 VDD.n2563 VDD.n844 240
R2337 VDD.n2563 VDD.n845 240
R2338 VDD.n1462 VDD.n845 240
R2339 VDD.n1984 VDD.n1462 240
R2340 VDD.n1984 VDD.n1457 240
R2341 VDD.n1457 VDD.n1434 240
R2342 VDD.n1434 VDD.n1428 240
R2343 VDD.n2031 VDD.n1428 240
R2344 VDD.n2031 VDD.n1413 240
R2345 VDD.n2044 VDD.n1413 240
R2346 VDD.n2044 VDD.n1399 240
R2347 VDD.n1424 VDD.n1399 240
R2348 VDD.n2039 VDD.n1424 240
R2349 VDD.n2039 VDD.n1371 240
R2350 VDD.n2036 VDD.n1371 240
R2351 VDD.n2036 VDD.n1366 240
R2352 VDD.n1366 VDD.n1340 240
R2353 VDD.n1357 VDD.n1340 240
R2354 VDD.n1357 VDD.n1334 240
R2355 VDD.n1334 VDD.n1203 240
R2356 VDD.n2146 VDD.n1203 240
R2357 VDD.n2147 VDD.n2146 240
R2358 VDD.n2147 VDD.n1327 240
R2359 VDD.n1327 VDD.n1224 240
R2360 VDD.n2383 VDD.n1224 240
R2361 VDD.n2383 VDD.n1233 240
R2362 VDD.n2509 VDD.n1233 240
R2363 VDD.n2509 VDD.n1240 240
R2364 VDD.n1320 VDD.n1240 240
R2365 VDD.n1320 VDD.n1263 240
R2366 VDD.n2397 VDD.n1263 240
R2367 VDD.n2397 VDD.n1274 240
R2368 VDD.n2401 VDD.n1274 240
R2369 VDD.n2401 VDD.n1287 240
R2370 VDD.n2437 VDD.n1287 240
R2371 VDD.n2437 VDD.n1293 240
R2372 VDD.n2470 VDD.n1315 240
R2373 VDD.n2466 VDD.n1315 240
R2374 VDD.n2464 VDD.n2463 240
R2375 VDD.n2460 VDD.n2459 240
R2376 VDD.n2456 VDD.n2455 240
R2377 VDD.n2452 VDD.n2451 240
R2378 VDD.n2448 VDD.n2447 240
R2379 VDD.n2444 VDD.n2443 240
R2380 VDD.n1791 VDD.n1530 240
R2381 VDD.n1870 VDD.n1530 240
R2382 VDD.n1870 VDD.n1531 240
R2383 VDD.n1531 VDD.n1522 240
R2384 VDD.n1865 VDD.n1522 240
R2385 VDD.n1865 VDD.n1503 240
R2386 VDD.n1904 VDD.n1503 240
R2387 VDD.n1904 VDD.n1504 240
R2388 VDD.n1504 VDD.n1495 240
R2389 VDD.n1507 VDD.n1495 240
R2390 VDD.n1507 VDD.n1470 240
R2391 VDD.n1943 VDD.n1470 240
R2392 VDD.n1944 VDD.n1943 240
R2393 VDD.n1944 VDD.n842 240
R2394 VDD.n1953 VDD.n842 240
R2395 VDD.n1954 VDD.n1953 240
R2396 VDD.n1954 VDD.n1458 240
R2397 VDD.n1991 VDD.n1458 240
R2398 VDD.n1991 VDD.n1435 240
R2399 VDD.n1987 VDD.n1435 240
R2400 VDD.n1987 VDD.n1415 240
R2401 VDD.n2057 VDD.n1415 240
R2402 VDD.n2057 VDD.n1416 240
R2403 VDD.n1416 VDD.n1401 240
R2404 VDD.n2052 VDD.n1401 240
R2405 VDD.n2052 VDD.n1422 240
R2406 VDD.n1422 VDD.n1372 240
R2407 VDD.n1418 VDD.n1372 240
R2408 VDD.n1418 VDD.n1338 240
R2409 VDD.n2132 VDD.n1338 240
R2410 VDD.n2132 VDD.n1335 240
R2411 VDD.n2138 VDD.n1335 240
R2412 VDD.n2138 VDD.n1205 240
R2413 VDD.n1328 VDD.n1205 240
R2414 VDD.n2149 VDD.n1328 240
R2415 VDD.n2152 VDD.n2149 240
R2416 VDD.n2152 VDD.n1226 240
R2417 VDD.n1235 VDD.n1226 240
R2418 VDD.n2513 VDD.n1235 240
R2419 VDD.n2513 VDD.n1236 240
R2420 VDD.n1279 VDD.n1236 240
R2421 VDD.n1280 VDD.n1279 240
R2422 VDD.n1280 VDD.n1265 240
R2423 VDD.n1276 VDD.n1265 240
R2424 VDD.n2490 VDD.n1276 240
R2425 VDD.n2490 VDD.n1277 240
R2426 VDD.n2486 VDD.n1277 240
R2427 VDD.n2486 VDD.n1285 240
R2428 VDD.n2478 VDD.n1285 240
R2429 VDD.n1787 VDD.n1549 240
R2430 VDD.n1785 VDD.n1784 240
R2431 VDD.n1781 VDD.n1780 240
R2432 VDD.n1777 VDD.n1776 240
R2433 VDD.n1773 VDD.n1772 240
R2434 VDD.n1769 VDD.n1768 240
R2435 VDD.n1765 VDD.n1764 240
R2436 VDD.n1761 VDD.n1547 240
R2437 VDD.n1836 VDD.n1545 240
R2438 VDD.n1836 VDD.n1529 240
R2439 VDD.n1529 VDD.n1519 240
R2440 VDD.n1879 VDD.n1519 240
R2441 VDD.n1879 VDD.n1517 240
R2442 VDD.n1883 VDD.n1517 240
R2443 VDD.n1883 VDD.n1502 240
R2444 VDD.n1891 VDD.n1502 240
R2445 VDD.n1891 VDD.n1494 240
R2446 VDD.n1896 VDD.n1494 240
R2447 VDD.n1896 VDD.n1511 240
R2448 VDD.n1511 VDD.n1468 240
R2449 VDD.n1946 VDD.n1468 240
R2450 VDD.n1946 VDD.n847 240
R2451 VDD.n1466 VDD.n847 240
R2452 VDD.n1952 VDD.n1466 240
R2453 VDD.n1952 VDD.n1464 240
R2454 VDD.n1464 VDD.n1432 240
R2455 VDD.n2026 VDD.n1432 240
R2456 VDD.n2026 VDD.n1430 240
R2457 VDD.n2030 VDD.n1430 240
R2458 VDD.n2030 VDD.n1414 240
R2459 VDD.n2046 VDD.n1414 240
R2460 VDD.n2046 VDD.n1400 240
R2461 VDD.n2050 VDD.n1400 240
R2462 VDD.n2050 VDD.n1369 240
R2463 VDD.n2105 VDD.n1369 240
R2464 VDD.n2105 VDD.n1367 240
R2465 VDD.n2110 VDD.n1367 240
R2466 VDD.n2110 VDD.n1341 240
R2467 VDD.n1341 VDD.n1332 240
R2468 VDD.n2140 VDD.n1332 240
R2469 VDD.n2140 VDD.n1204 240
R2470 VDD.n2144 VDD.n1204 240
R2471 VDD.n2144 VDD.n1325 240
R2472 VDD.n2154 VDD.n1325 240
R2473 VDD.n2154 VDD.n1225 240
R2474 VDD.n2385 VDD.n1225 240
R2475 VDD.n2385 VDD.n1234 240
R2476 VDD.n1242 VDD.n1234 240
R2477 VDD.n2390 VDD.n1242 240
R2478 VDD.n2391 VDD.n2390 240
R2479 VDD.n2391 VDD.n1264 240
R2480 VDD.n2395 VDD.n1264 240
R2481 VDD.n2395 VDD.n1275 240
R2482 VDD.n2403 VDD.n1275 240
R2483 VDD.n2403 VDD.n1288 240
R2484 VDD.n2435 VDD.n1288 240
R2485 VDD.n2435 VDD.n1294 240
R2486 VDD.n2474 VDD.n1298 240
R2487 VDD.n2408 VDD.n2407 240
R2488 VDD.n2412 VDD.n2411 240
R2489 VDD.n2416 VDD.n2415 240
R2490 VDD.n2420 VDD.n2419 240
R2491 VDD.n2424 VDD.n2423 240
R2492 VDD.n2428 VDD.n2427 240
R2493 VDD.n2430 VDD.n1313 240
R2494 VDD.n1653 VDD.n1607 240
R2495 VDD.n1653 VDD.n1601 240
R2496 VDD.n1661 VDD.n1601 240
R2497 VDD.n1661 VDD.n1599 240
R2498 VDD.n1665 VDD.n1599 240
R2499 VDD.n1665 VDD.n1593 240
R2500 VDD.n1674 VDD.n1593 240
R2501 VDD.n1674 VDD.n1591 240
R2502 VDD.n1678 VDD.n1591 240
R2503 VDD.n1678 VDD.n1586 240
R2504 VDD.n1687 VDD.n1586 240
R2505 VDD.n1687 VDD.n1584 240
R2506 VDD.n1691 VDD.n1584 240
R2507 VDD.n1691 VDD.n1579 240
R2508 VDD.n1699 VDD.n1579 240
R2509 VDD.n1699 VDD.n1577 240
R2510 VDD.n1704 VDD.n1577 240
R2511 VDD.n1704 VDD.n1570 240
R2512 VDD.n1751 VDD.n1570 240
R2513 VDD.n1752 VDD.n1751 240
R2514 VDD.n1752 VDD.n1567 240
R2515 VDD.n1759 VDD.n1567 240
R2516 VDD.n1759 VDD.n1568 240
R2517 VDD.n1568 VDD.n1540 240
R2518 VDD.n1846 VDD.n1540 240
R2519 VDD.n1846 VDD.n1534 240
R2520 VDD.n1862 VDD.n1534 240
R2521 VDD.n1862 VDD.n1535 240
R2522 VDD.n1855 VDD.n1535 240
R2523 VDD.n1855 VDD.n1491 240
R2524 VDD.n1914 VDD.n1491 240
R2525 VDD.n1914 VDD.n1485 240
R2526 VDD.n1930 VDD.n1485 240
R2527 VDD.n1930 VDD.n1486 240
R2528 VDD.n1923 VDD.n1486 240
R2529 VDD.n1923 VDD.n859 240
R2530 VDD.n2552 VDD.n859 240
R2531 VDD.n2552 VDD.n860 240
R2532 VDD.n1455 VDD.n860 240
R2533 VDD.n1994 VDD.n1455 240
R2534 VDD.n1994 VDD.n1450 240
R2535 VDD.n2010 VDD.n1450 240
R2536 VDD.n2010 VDD.n1451 240
R2537 VDD.n2003 VDD.n1451 240
R2538 VDD.n2003 VDD.n1397 240
R2539 VDD.n2079 VDD.n1397 240
R2540 VDD.n2079 VDD.n1391 240
R2541 VDD.n2091 VDD.n1391 240
R2542 VDD.n2091 VDD.n1392 240
R2543 VDD.n1392 VDD.n1363 240
R2544 VDD.n2113 VDD.n1363 240
R2545 VDD.n2113 VDD.n1359 240
R2546 VDD.n2121 VDD.n1359 240
R2547 VDD.n2121 VDD.n1200 240
R2548 VDD.n2541 VDD.n1200 240
R2549 VDD.n2541 VDD.n1201 240
R2550 VDD.n2529 VDD.n1201 240
R2551 VDD.n2529 VDD.n1217 240
R2552 VDD.n2522 VDD.n1217 240
R2553 VDD.n2522 VDD.n1222 240
R2554 VDD.n1252 VDD.n1222 240
R2555 VDD.n1252 VDD.n1245 240
R2556 VDD.n2506 VDD.n1245 240
R2557 VDD.n2506 VDD.n1246 240
R2558 VDD.n2499 VDD.n1246 240
R2559 VDD.n2499 VDD.n1260 240
R2560 VDD.n2199 VDD.n1260 240
R2561 VDD.n2200 VDD.n2199 240
R2562 VDD.n2200 VDD.n2191 240
R2563 VDD.n2206 VDD.n2191 240
R2564 VDD.n2207 VDD.n2206 240
R2565 VDD.n2208 VDD.n2207 240
R2566 VDD.n2208 VDD.n2188 240
R2567 VDD.n2347 VDD.n2188 240
R2568 VDD.n2347 VDD.n2189 240
R2569 VDD.n2343 VDD.n2189 240
R2570 VDD.n2343 VDD.n2212 240
R2571 VDD.n2339 VDD.n2212 240
R2572 VDD.n2339 VDD.n2217 240
R2573 VDD.n2335 VDD.n2217 240
R2574 VDD.n2335 VDD.n2219 240
R2575 VDD.n2331 VDD.n2219 240
R2576 VDD.n2331 VDD.n2223 240
R2577 VDD.n2327 VDD.n2223 240
R2578 VDD.n2327 VDD.n2225 240
R2579 VDD.n2323 VDD.n2225 240
R2580 VDD.n2323 VDD.n2231 240
R2581 VDD.n2319 VDD.n2231 240
R2582 VDD.n2319 VDD.n2233 240
R2583 VDD.n2315 VDD.n2233 240
R2584 VDD.n2315 VDD.n2238 240
R2585 VDD.n2311 VDD.n2238 240
R2586 VDD.n2311 VDD.n2240 240
R2587 VDD.n2251 VDD.n2250 240
R2588 VDD.n2301 VDD.n2250 240
R2589 VDD.n2299 VDD.n2298 240
R2590 VDD.n2295 VDD.n2294 240
R2591 VDD.n2291 VDD.n2290 240
R2592 VDD.n2287 VDD.n2286 240
R2593 VDD.n2283 VDD.n2282 240
R2594 VDD.n2279 VDD.n2278 240
R2595 VDD.n1655 VDD.n1605 240
R2596 VDD.n1655 VDD.n1603 240
R2597 VDD.n1659 VDD.n1603 240
R2598 VDD.n1659 VDD.n1597 240
R2599 VDD.n1667 VDD.n1597 240
R2600 VDD.n1667 VDD.n1595 240
R2601 VDD.n1671 VDD.n1595 240
R2602 VDD.n1671 VDD.n1589 240
R2603 VDD.n1680 VDD.n1589 240
R2604 VDD.n1680 VDD.n1587 240
R2605 VDD.n1684 VDD.n1587 240
R2606 VDD.n1684 VDD.n1583 240
R2607 VDD.n1693 VDD.n1583 240
R2608 VDD.n1693 VDD.n1581 240
R2609 VDD.n1697 VDD.n1581 240
R2610 VDD.n1697 VDD.n1575 240
R2611 VDD.n1706 VDD.n1575 240
R2612 VDD.n1706 VDD.n1572 240
R2613 VDD.n1749 VDD.n1572 240
R2614 VDD.n1749 VDD.n1573 240
R2615 VDD.n1745 VDD.n1573 240
R2616 VDD.n1745 VDD.n1566 240
R2617 VDD.n1742 VDD.n1566 240
R2618 VDD.n1742 VDD.n1741 240
R2619 VDD.n1741 VDD.n1541 240
R2620 VDD.n1734 VDD.n1541 240
R2621 VDD.n1734 VDD.n1533 240
R2622 VDD.n1715 VDD.n1533 240
R2623 VDD.n1726 VDD.n1715 240
R2624 VDD.n1726 VDD.n1725 240
R2625 VDD.n1725 VDD.n1492 240
R2626 VDD.n1492 VDD.n1481 240
R2627 VDD.n1932 VDD.n1481 240
R2628 VDD.n1933 VDD.n1932 240
R2629 VDD.n1934 VDD.n1933 240
R2630 VDD.n1934 VDD.n856 240
R2631 VDD.n2554 VDD.n856 240
R2632 VDD.n2554 VDD.n857 240
R2633 VDD.n1971 VDD.n857 240
R2634 VDD.n1971 VDD.n1456 240
R2635 VDD.n1456 VDD.n1448 240
R2636 VDD.n2012 VDD.n1448 240
R2637 VDD.n2017 VDD.n2012 240
R2638 VDD.n2017 VDD.n2016 240
R2639 VDD.n2016 VDD.n2013 240
R2640 VDD.n2013 VDD.n1398 240
R2641 VDD.n1398 VDD.n1387 240
R2642 VDD.n2093 VDD.n1387 240
R2643 VDD.n2094 VDD.n2093 240
R2644 VDD.n2096 VDD.n2094 240
R2645 VDD.n2096 VDD.n1365 240
R2646 VDD.n1365 VDD.n1352 240
R2647 VDD.n2123 VDD.n1352 240
R2648 VDD.n2123 VDD.n1356 240
R2649 VDD.n1356 VDD.n1202 240
R2650 VDD.n1214 VDD.n1202 240
R2651 VDD.n2531 VDD.n1214 240
R2652 VDD.n2531 VDD.n1215 240
R2653 VDD.n1223 VDD.n1215 240
R2654 VDD.n2381 VDD.n1223 240
R2655 VDD.n2381 VDD.n2157 240
R2656 VDD.n2374 VDD.n2157 240
R2657 VDD.n2374 VDD.n1243 240
R2658 VDD.n2175 VDD.n1243 240
R2659 VDD.n2175 VDD.n1262 240
R2660 VDD.n2364 VDD.n1262 240
R2661 VDD.n2364 VDD.n2363 240
R2662 VDD.n2363 VDD.n2179 240
R2663 VDD.n2356 VDD.n2179 240
R2664 VDD.n2356 VDD.n2355 240
R2665 VDD.n2355 VDD.n2183 240
R2666 VDD.n2351 VDD.n2183 240
R2667 VDD.n2351 VDD.n2350 240
R2668 VDD.n2350 VDD.n2349 240
R2669 VDD.n2349 VDD.n2185 240
R2670 VDD.n2213 VDD.n2185 240
R2671 VDD.n2214 VDD.n2213 240
R2672 VDD.n2215 VDD.n2214 240
R2673 VDD.n2256 VDD.n2215 240
R2674 VDD.n2256 VDD.n2220 240
R2675 VDD.n2221 VDD.n2220 240
R2676 VDD.n2222 VDD.n2221 240
R2677 VDD.n2261 VDD.n2222 240
R2678 VDD.n2261 VDD.n2227 240
R2679 VDD.n2228 VDD.n2227 240
R2680 VDD.n2229 VDD.n2228 240
R2681 VDD.n2266 VDD.n2229 240
R2682 VDD.n2266 VDD.n2234 240
R2683 VDD.n2235 VDD.n2234 240
R2684 VDD.n2236 VDD.n2235 240
R2685 VDD.n2271 VDD.n2236 240
R2686 VDD.n2271 VDD.n2241 240
R2687 VDD.n2242 VDD.n2241 240
R2688 VDD.n1618 VDD.n1609 240
R2689 VDD.n1622 VDD.n1621 240
R2690 VDD.n1626 VDD.n1625 240
R2691 VDD.n1630 VDD.n1629 240
R2692 VDD.n1634 VDD.n1633 240
R2693 VDD.n1638 VDD.n1637 240
R2694 VDD.n1642 VDD.n1641 240
R2695 VDD.n1646 VDD.n1617 240
R2696 VDD.n5640 VDD.n5604 240
R2697 VDD.n5613 VDD.n5604 240
R2698 VDD.n6044 VDD.n5613 240
R2699 VDD.n6044 VDD.n5614 240
R2700 VDD.n6040 VDD.n5614 240
R2701 VDD.n6040 VDD.n5645 240
R2702 VDD.n6032 VDD.n5645 240
R2703 VDD.n6032 VDD.n5655 240
R2704 VDD.n6028 VDD.n5655 240
R2705 VDD.n6028 VDD.n5657 240
R2706 VDD.n6020 VDD.n5657 240
R2707 VDD.n6020 VDD.n5667 240
R2708 VDD.n6016 VDD.n5667 240
R2709 VDD.n6016 VDD.n5669 240
R2710 VDD.n6008 VDD.n5669 240
R2711 VDD.n6008 VDD.n5679 240
R2712 VDD.n6004 VDD.n5679 240
R2713 VDD.n6004 VDD.n5681 240
R2714 VDD.n5996 VDD.n5681 240
R2715 VDD.n5996 VDD.n5691 240
R2716 VDD.n5992 VDD.n5691 240
R2717 VDD.n5992 VDD.n5693 240
R2718 VDD.n5984 VDD.n5693 240
R2719 VDD.n5639 VDD.n5638 240
R2720 VDD.n5636 VDD.n5617 240
R2721 VDD.n5632 VDD.n5631 240
R2722 VDD.n5629 VDD.n5620 240
R2723 VDD.n5624 VDD.n5623 240
R2724 VDD.n6066 VDD.n6065 240
R2725 VDD.n6063 VDD.n5595 240
R2726 VDD.n6059 VDD.n6058 240
R2727 VDD.n6052 VDD.n5598 240
R2728 VDD.n6052 VDD.n5600 240
R2729 VDD.n5611 VDD.n5600 240
R2730 VDD.n5916 VDD.n5611 240
R2731 VDD.n5916 VDD.n5647 240
R2732 VDD.n5919 VDD.n5647 240
R2733 VDD.n5919 VDD.n5653 240
R2734 VDD.n5922 VDD.n5653 240
R2735 VDD.n5922 VDD.n5659 240
R2736 VDD.n5925 VDD.n5659 240
R2737 VDD.n5925 VDD.n5665 240
R2738 VDD.n5928 VDD.n5665 240
R2739 VDD.n5928 VDD.n5671 240
R2740 VDD.n5931 VDD.n5671 240
R2741 VDD.n5931 VDD.n5677 240
R2742 VDD.n5934 VDD.n5677 240
R2743 VDD.n5934 VDD.n5683 240
R2744 VDD.n5937 VDD.n5683 240
R2745 VDD.n5937 VDD.n5689 240
R2746 VDD.n5940 VDD.n5689 240
R2747 VDD.n5940 VDD.n5695 240
R2748 VDD.n5943 VDD.n5695 240
R2749 VDD.n5943 VDD.n5701 240
R2750 VDD.n5980 VDD.n5978 240
R2751 VDD.n5976 VDD.n5705 240
R2752 VDD.n5972 VDD.n5970 240
R2753 VDD.n5968 VDD.n5707 240
R2754 VDD.n5961 VDD.n5959 240
R2755 VDD.n5956 VDD.n5955 240
R2756 VDD.n5953 VDD.n5914 240
R2757 VDD.n5949 VDD.n5947 240
R2758 VDD.n6050 VDD.n5605 240
R2759 VDD.n6050 VDD.n5606 240
R2760 VDD.n6046 VDD.n5606 240
R2761 VDD.n6046 VDD.n5609 240
R2762 VDD.n6038 VDD.n5609 240
R2763 VDD.n6038 VDD.n5648 240
R2764 VDD.n6034 VDD.n5648 240
R2765 VDD.n6034 VDD.n5650 240
R2766 VDD.n6026 VDD.n5650 240
R2767 VDD.n6026 VDD.n5660 240
R2768 VDD.n6022 VDD.n5660 240
R2769 VDD.n6022 VDD.n5662 240
R2770 VDD.n6014 VDD.n5662 240
R2771 VDD.n6014 VDD.n5672 240
R2772 VDD.n6010 VDD.n5672 240
R2773 VDD.n6010 VDD.n5674 240
R2774 VDD.n6002 VDD.n5674 240
R2775 VDD.n6002 VDD.n5684 240
R2776 VDD.n5998 VDD.n5684 240
R2777 VDD.n5998 VDD.n5686 240
R2778 VDD.n5990 VDD.n5686 240
R2779 VDD.n5990 VDD.n5697 240
R2780 VDD.n5986 VDD.n5697 240
R2781 VDD.n5729 VDD.n5727 240
R2782 VDD.n5733 VDD.n5727 240
R2783 VDD.n5737 VDD.n5735 240
R2784 VDD.n5741 VDD.n5725 240
R2785 VDD.n5869 VDD.n5743 240
R2786 VDD.n5867 VDD.n5744 240
R2787 VDD.n5863 VDD.n5861 240
R2788 VDD.n5859 VDD.n5746 240
R2789 VDD.n5818 VDD.n5602 240
R2790 VDD.n5821 VDD.n5602 240
R2791 VDD.n5821 VDD.n5610 240
R2792 VDD.n5824 VDD.n5610 240
R2793 VDD.n5824 VDD.n5646 240
R2794 VDD.n5827 VDD.n5646 240
R2795 VDD.n5827 VDD.n5652 240
R2796 VDD.n5830 VDD.n5652 240
R2797 VDD.n5830 VDD.n5658 240
R2798 VDD.n5833 VDD.n5658 240
R2799 VDD.n5833 VDD.n5664 240
R2800 VDD.n5836 VDD.n5664 240
R2801 VDD.n5836 VDD.n5670 240
R2802 VDD.n5839 VDD.n5670 240
R2803 VDD.n5839 VDD.n5676 240
R2804 VDD.n5842 VDD.n5676 240
R2805 VDD.n5842 VDD.n5682 240
R2806 VDD.n5845 VDD.n5682 240
R2807 VDD.n5845 VDD.n5688 240
R2808 VDD.n5848 VDD.n5688 240
R2809 VDD.n5848 VDD.n5694 240
R2810 VDD.n5851 VDD.n5694 240
R2811 VDD.n5851 VDD.n5700 240
R2812 VDD.n5776 VDD.n5774 240
R2813 VDD.n5780 VDD.n5769 240
R2814 VDD.n5783 VDD.n5782 240
R2815 VDD.n5784 VDD.n5783 240
R2816 VDD.n5790 VDD.n5788 240
R2817 VDD.n5807 VDD.n5750 240
R2818 VDD.n5811 VDD.n5809 240
R2819 VDD.n5815 VDD.n5748 240
R2820 VDD.n7356 VDD.n7089 240
R2821 VDD.n7435 VDD.n7089 240
R2822 VDD.n7435 VDD.n7086 240
R2823 VDD.n7440 VDD.n7086 240
R2824 VDD.n7440 VDD.n7087 240
R2825 VDD.n7087 VDD.n7062 240
R2826 VDD.n7469 VDD.n7062 240
R2827 VDD.n7469 VDD.n7059 240
R2828 VDD.n7474 VDD.n7059 240
R2829 VDD.n7474 VDD.n7060 240
R2830 VDD.n7060 VDD.n7037 240
R2831 VDD.n7504 VDD.n7037 240
R2832 VDD.n7504 VDD.n6411 240
R2833 VDD.n8124 VDD.n6411 240
R2834 VDD.n8124 VDD.n6412 240
R2835 VDD.n7519 VDD.n6412 240
R2836 VDD.n7545 VDD.n7519 240
R2837 VDD.n7545 VDD.n6999 240
R2838 VDD.n7587 VDD.n6999 240
R2839 VDD.n7587 VDD.n7000 240
R2840 VDD.n7000 VDD.n6974 240
R2841 VDD.n7622 VDD.n6974 240
R2842 VDD.n7622 VDD.n6965 240
R2843 VDD.n7639 VDD.n6965 240
R2844 VDD.n7639 VDD.n6966 240
R2845 VDD.n6966 VDD.n6936 240
R2846 VDD.n7666 VDD.n6936 240
R2847 VDD.n7666 VDD.n6937 240
R2848 VDD.n6937 VDD.n6905 240
R2849 VDD.n7693 VDD.n6905 240
R2850 VDD.n7693 VDD.n6906 240
R2851 VDD.n6906 VDD.n6769 240
R2852 VDD.n8101 VDD.n6769 240
R2853 VDD.n8101 VDD.n6770 240
R2854 VDD.n7725 VDD.n6770 240
R2855 VDD.n7725 VDD.n6790 240
R2856 VDD.n8082 VDD.n6790 240
R2857 VDD.n8082 VDD.n6791 240
R2858 VDD.n8078 VDD.n6791 240
R2859 VDD.n8078 VDD.n6794 240
R2860 VDD.n6831 VDD.n6794 240
R2861 VDD.n6831 VDD.n6829 240
R2862 VDD.n8059 VDD.n6829 240
R2863 VDD.n8059 VDD.n6830 240
R2864 VDD.n8055 VDD.n6830 240
R2865 VDD.n8055 VDD.n6835 240
R2866 VDD.n8047 VDD.n6835 240
R2867 VDD.n8047 VDD.n6852 240
R2868 VDD.n8043 VDD.n6852 240
R2869 VDD.n7391 VDD.n7357 240
R2870 VDD.n7387 VDD.n7386 240
R2871 VDD.n7383 VDD.n7382 240
R2872 VDD.n7379 VDD.n7378 240
R2873 VDD.n7375 VDD.n7374 240
R2874 VDD.n7371 VDD.n7370 240
R2875 VDD.n7367 VDD.n7366 240
R2876 VDD.n7363 VDD.n7362 240
R2877 VDD.n7401 VDD.n7106 240
R2878 VDD.n7401 VDD.n7091 240
R2879 VDD.n7406 VDD.n7091 240
R2880 VDD.n7406 VDD.n7084 240
R2881 VDD.n7084 VDD.n7078 240
R2882 VDD.n7448 VDD.n7078 240
R2883 VDD.n7448 VDD.n7064 240
R2884 VDD.n7452 VDD.n7064 240
R2885 VDD.n7452 VDD.n7056 240
R2886 VDD.n7461 VDD.n7056 240
R2887 VDD.n7461 VDD.n7072 240
R2888 VDD.n7072 VDD.n7036 240
R2889 VDD.n7036 VDD.n6407 240
R2890 VDD.n8126 VDD.n6407 240
R2891 VDD.n8126 VDD.n6408 240
R2892 VDD.n7025 VDD.n6408 240
R2893 VDD.n7547 VDD.n7025 240
R2894 VDD.n7547 VDD.n7020 240
R2895 VDD.n7020 VDD.n6997 240
R2896 VDD.n6997 VDD.n6991 240
R2897 VDD.n7594 VDD.n6991 240
R2898 VDD.n7594 VDD.n6976 240
R2899 VDD.n7607 VDD.n6976 240
R2900 VDD.n7607 VDD.n6962 240
R2901 VDD.n6987 VDD.n6962 240
R2902 VDD.n7602 VDD.n6987 240
R2903 VDD.n7602 VDD.n6934 240
R2904 VDD.n7599 VDD.n6934 240
R2905 VDD.n7599 VDD.n6929 240
R2906 VDD.n6929 VDD.n6903 240
R2907 VDD.n6920 VDD.n6903 240
R2908 VDD.n6920 VDD.n6897 240
R2909 VDD.n6897 VDD.n6766 240
R2910 VDD.n7709 VDD.n6766 240
R2911 VDD.n7710 VDD.n7709 240
R2912 VDD.n7710 VDD.n6890 240
R2913 VDD.n6890 VDD.n6787 240
R2914 VDD.n7946 VDD.n6787 240
R2915 VDD.n7946 VDD.n6796 240
R2916 VDD.n8072 VDD.n6796 240
R2917 VDD.n8072 VDD.n6803 240
R2918 VDD.n6883 VDD.n6803 240
R2919 VDD.n6883 VDD.n6826 240
R2920 VDD.n7960 VDD.n6826 240
R2921 VDD.n7960 VDD.n6837 240
R2922 VDD.n7964 VDD.n6837 240
R2923 VDD.n7964 VDD.n6850 240
R2924 VDD.n8000 VDD.n6850 240
R2925 VDD.n8000 VDD.n6856 240
R2926 VDD.n8033 VDD.n6878 240
R2927 VDD.n8029 VDD.n6878 240
R2928 VDD.n8027 VDD.n8026 240
R2929 VDD.n8023 VDD.n8022 240
R2930 VDD.n8019 VDD.n8018 240
R2931 VDD.n8015 VDD.n8014 240
R2932 VDD.n8011 VDD.n8010 240
R2933 VDD.n8007 VDD.n8006 240
R2934 VDD.n7354 VDD.n7093 240
R2935 VDD.n7433 VDD.n7093 240
R2936 VDD.n7433 VDD.n7094 240
R2937 VDD.n7094 VDD.n7085 240
R2938 VDD.n7428 VDD.n7085 240
R2939 VDD.n7428 VDD.n7066 240
R2940 VDD.n7467 VDD.n7066 240
R2941 VDD.n7467 VDD.n7067 240
R2942 VDD.n7067 VDD.n7058 240
R2943 VDD.n7070 VDD.n7058 240
R2944 VDD.n7070 VDD.n7033 240
R2945 VDD.n7506 VDD.n7033 240
R2946 VDD.n7507 VDD.n7506 240
R2947 VDD.n7507 VDD.n6405 240
R2948 VDD.n7516 VDD.n6405 240
R2949 VDD.n7517 VDD.n7516 240
R2950 VDD.n7517 VDD.n7021 240
R2951 VDD.n7554 VDD.n7021 240
R2952 VDD.n7554 VDD.n6998 240
R2953 VDD.n7550 VDD.n6998 240
R2954 VDD.n7550 VDD.n6978 240
R2955 VDD.n7620 VDD.n6978 240
R2956 VDD.n7620 VDD.n6979 240
R2957 VDD.n6979 VDD.n6964 240
R2958 VDD.n7615 VDD.n6964 240
R2959 VDD.n7615 VDD.n6985 240
R2960 VDD.n6985 VDD.n6935 240
R2961 VDD.n6981 VDD.n6935 240
R2962 VDD.n6981 VDD.n6901 240
R2963 VDD.n7695 VDD.n6901 240
R2964 VDD.n7695 VDD.n6898 240
R2965 VDD.n7701 VDD.n6898 240
R2966 VDD.n7701 VDD.n6768 240
R2967 VDD.n6891 VDD.n6768 240
R2968 VDD.n7712 VDD.n6891 240
R2969 VDD.n7715 VDD.n7712 240
R2970 VDD.n7715 VDD.n6789 240
R2971 VDD.n6798 VDD.n6789 240
R2972 VDD.n8076 VDD.n6798 240
R2973 VDD.n8076 VDD.n6799 240
R2974 VDD.n6842 VDD.n6799 240
R2975 VDD.n6843 VDD.n6842 240
R2976 VDD.n6843 VDD.n6828 240
R2977 VDD.n6839 VDD.n6828 240
R2978 VDD.n8053 VDD.n6839 240
R2979 VDD.n8053 VDD.n6840 240
R2980 VDD.n8049 VDD.n6840 240
R2981 VDD.n8049 VDD.n6848 240
R2982 VDD.n8041 VDD.n6848 240
R2983 VDD.n7350 VDD.n7112 240
R2984 VDD.n7348 VDD.n7347 240
R2985 VDD.n7344 VDD.n7343 240
R2986 VDD.n7340 VDD.n7339 240
R2987 VDD.n7336 VDD.n7335 240
R2988 VDD.n7332 VDD.n7331 240
R2989 VDD.n7328 VDD.n7327 240
R2990 VDD.n7324 VDD.n7110 240
R2991 VDD.n7399 VDD.n7108 240
R2992 VDD.n7399 VDD.n7092 240
R2993 VDD.n7092 VDD.n7082 240
R2994 VDD.n7442 VDD.n7082 240
R2995 VDD.n7442 VDD.n7080 240
R2996 VDD.n7446 VDD.n7080 240
R2997 VDD.n7446 VDD.n7065 240
R2998 VDD.n7454 VDD.n7065 240
R2999 VDD.n7454 VDD.n7057 240
R3000 VDD.n7459 VDD.n7057 240
R3001 VDD.n7459 VDD.n7074 240
R3002 VDD.n7074 VDD.n7031 240
R3003 VDD.n7509 VDD.n7031 240
R3004 VDD.n7509 VDD.n6410 240
R3005 VDD.n7029 VDD.n6410 240
R3006 VDD.n7515 VDD.n7029 240
R3007 VDD.n7515 VDD.n7027 240
R3008 VDD.n7027 VDD.n6995 240
R3009 VDD.n7589 VDD.n6995 240
R3010 VDD.n7589 VDD.n6993 240
R3011 VDD.n7593 VDD.n6993 240
R3012 VDD.n7593 VDD.n6977 240
R3013 VDD.n7609 VDD.n6977 240
R3014 VDD.n7609 VDD.n6963 240
R3015 VDD.n7613 VDD.n6963 240
R3016 VDD.n7613 VDD.n6932 240
R3017 VDD.n7668 VDD.n6932 240
R3018 VDD.n7668 VDD.n6930 240
R3019 VDD.n7673 VDD.n6930 240
R3020 VDD.n7673 VDD.n6904 240
R3021 VDD.n6904 VDD.n6895 240
R3022 VDD.n7703 VDD.n6895 240
R3023 VDD.n7703 VDD.n6767 240
R3024 VDD.n7707 VDD.n6767 240
R3025 VDD.n7707 VDD.n6888 240
R3026 VDD.n7717 VDD.n6888 240
R3027 VDD.n7717 VDD.n6788 240
R3028 VDD.n7948 VDD.n6788 240
R3029 VDD.n7948 VDD.n6797 240
R3030 VDD.n6805 VDD.n6797 240
R3031 VDD.n7953 VDD.n6805 240
R3032 VDD.n7954 VDD.n7953 240
R3033 VDD.n7954 VDD.n6827 240
R3034 VDD.n7958 VDD.n6827 240
R3035 VDD.n7958 VDD.n6838 240
R3036 VDD.n7966 VDD.n6838 240
R3037 VDD.n7966 VDD.n6851 240
R3038 VDD.n7998 VDD.n6851 240
R3039 VDD.n7998 VDD.n6857 240
R3040 VDD.n8037 VDD.n6861 240
R3041 VDD.n7971 VDD.n7970 240
R3042 VDD.n7975 VDD.n7974 240
R3043 VDD.n7979 VDD.n7978 240
R3044 VDD.n7983 VDD.n7982 240
R3045 VDD.n7987 VDD.n7986 240
R3046 VDD.n7991 VDD.n7990 240
R3047 VDD.n7993 VDD.n6876 240
R3048 VDD.n7216 VDD.n7170 240
R3049 VDD.n7216 VDD.n7164 240
R3050 VDD.n7224 VDD.n7164 240
R3051 VDD.n7224 VDD.n7162 240
R3052 VDD.n7228 VDD.n7162 240
R3053 VDD.n7228 VDD.n7156 240
R3054 VDD.n7237 VDD.n7156 240
R3055 VDD.n7237 VDD.n7154 240
R3056 VDD.n7241 VDD.n7154 240
R3057 VDD.n7241 VDD.n7149 240
R3058 VDD.n7250 VDD.n7149 240
R3059 VDD.n7250 VDD.n7147 240
R3060 VDD.n7254 VDD.n7147 240
R3061 VDD.n7254 VDD.n7142 240
R3062 VDD.n7262 VDD.n7142 240
R3063 VDD.n7262 VDD.n7140 240
R3064 VDD.n7267 VDD.n7140 240
R3065 VDD.n7267 VDD.n7133 240
R3066 VDD.n7314 VDD.n7133 240
R3067 VDD.n7315 VDD.n7314 240
R3068 VDD.n7315 VDD.n7130 240
R3069 VDD.n7322 VDD.n7130 240
R3070 VDD.n7322 VDD.n7131 240
R3071 VDD.n7131 VDD.n7103 240
R3072 VDD.n7409 VDD.n7103 240
R3073 VDD.n7409 VDD.n7097 240
R3074 VDD.n7425 VDD.n7097 240
R3075 VDD.n7425 VDD.n7098 240
R3076 VDD.n7418 VDD.n7098 240
R3077 VDD.n7418 VDD.n7054 240
R3078 VDD.n7477 VDD.n7054 240
R3079 VDD.n7477 VDD.n7048 240
R3080 VDD.n7493 VDD.n7048 240
R3081 VDD.n7493 VDD.n7049 240
R3082 VDD.n7486 VDD.n7049 240
R3083 VDD.n7486 VDD.n6422 240
R3084 VDD.n8115 VDD.n6422 240
R3085 VDD.n8115 VDD.n6423 240
R3086 VDD.n7018 VDD.n6423 240
R3087 VDD.n7557 VDD.n7018 240
R3088 VDD.n7557 VDD.n7013 240
R3089 VDD.n7573 VDD.n7013 240
R3090 VDD.n7573 VDD.n7014 240
R3091 VDD.n7566 VDD.n7014 240
R3092 VDD.n7566 VDD.n6960 240
R3093 VDD.n7642 VDD.n6960 240
R3094 VDD.n7642 VDD.n6954 240
R3095 VDD.n7654 VDD.n6954 240
R3096 VDD.n7654 VDD.n6955 240
R3097 VDD.n6955 VDD.n6926 240
R3098 VDD.n7676 VDD.n6926 240
R3099 VDD.n7676 VDD.n6922 240
R3100 VDD.n7684 VDD.n6922 240
R3101 VDD.n7684 VDD.n6763 240
R3102 VDD.n8104 VDD.n6763 240
R3103 VDD.n8104 VDD.n6764 240
R3104 VDD.n8092 VDD.n6764 240
R3105 VDD.n8092 VDD.n6780 240
R3106 VDD.n8085 VDD.n6780 240
R3107 VDD.n8085 VDD.n6785 240
R3108 VDD.n6815 VDD.n6785 240
R3109 VDD.n6815 VDD.n6808 240
R3110 VDD.n8069 VDD.n6808 240
R3111 VDD.n8069 VDD.n6809 240
R3112 VDD.n8062 VDD.n6809 240
R3113 VDD.n8062 VDD.n6823 240
R3114 VDD.n7762 VDD.n6823 240
R3115 VDD.n7763 VDD.n7762 240
R3116 VDD.n7763 VDD.n7754 240
R3117 VDD.n7769 VDD.n7754 240
R3118 VDD.n7770 VDD.n7769 240
R3119 VDD.n7771 VDD.n7770 240
R3120 VDD.n7771 VDD.n7751 240
R3121 VDD.n7910 VDD.n7751 240
R3122 VDD.n7910 VDD.n7752 240
R3123 VDD.n7906 VDD.n7752 240
R3124 VDD.n7906 VDD.n7775 240
R3125 VDD.n7902 VDD.n7775 240
R3126 VDD.n7902 VDD.n7780 240
R3127 VDD.n7898 VDD.n7780 240
R3128 VDD.n7898 VDD.n7782 240
R3129 VDD.n7894 VDD.n7782 240
R3130 VDD.n7894 VDD.n7786 240
R3131 VDD.n7890 VDD.n7786 240
R3132 VDD.n7890 VDD.n7788 240
R3133 VDD.n7886 VDD.n7788 240
R3134 VDD.n7886 VDD.n7794 240
R3135 VDD.n7882 VDD.n7794 240
R3136 VDD.n7882 VDD.n7796 240
R3137 VDD.n7878 VDD.n7796 240
R3138 VDD.n7878 VDD.n7801 240
R3139 VDD.n7874 VDD.n7801 240
R3140 VDD.n7874 VDD.n7803 240
R3141 VDD.n7814 VDD.n7813 240
R3142 VDD.n7864 VDD.n7813 240
R3143 VDD.n7862 VDD.n7861 240
R3144 VDD.n7858 VDD.n7857 240
R3145 VDD.n7854 VDD.n7853 240
R3146 VDD.n7850 VDD.n7849 240
R3147 VDD.n7846 VDD.n7845 240
R3148 VDD.n7842 VDD.n7841 240
R3149 VDD.n7218 VDD.n7168 240
R3150 VDD.n7218 VDD.n7166 240
R3151 VDD.n7222 VDD.n7166 240
R3152 VDD.n7222 VDD.n7160 240
R3153 VDD.n7230 VDD.n7160 240
R3154 VDD.n7230 VDD.n7158 240
R3155 VDD.n7234 VDD.n7158 240
R3156 VDD.n7234 VDD.n7152 240
R3157 VDD.n7243 VDD.n7152 240
R3158 VDD.n7243 VDD.n7150 240
R3159 VDD.n7247 VDD.n7150 240
R3160 VDD.n7247 VDD.n7146 240
R3161 VDD.n7256 VDD.n7146 240
R3162 VDD.n7256 VDD.n7144 240
R3163 VDD.n7260 VDD.n7144 240
R3164 VDD.n7260 VDD.n7138 240
R3165 VDD.n7269 VDD.n7138 240
R3166 VDD.n7269 VDD.n7135 240
R3167 VDD.n7312 VDD.n7135 240
R3168 VDD.n7312 VDD.n7136 240
R3169 VDD.n7308 VDD.n7136 240
R3170 VDD.n7308 VDD.n7129 240
R3171 VDD.n7305 VDD.n7129 240
R3172 VDD.n7305 VDD.n7304 240
R3173 VDD.n7304 VDD.n7104 240
R3174 VDD.n7297 VDD.n7104 240
R3175 VDD.n7297 VDD.n7096 240
R3176 VDD.n7278 VDD.n7096 240
R3177 VDD.n7289 VDD.n7278 240
R3178 VDD.n7289 VDD.n7288 240
R3179 VDD.n7288 VDD.n7055 240
R3180 VDD.n7055 VDD.n7044 240
R3181 VDD.n7495 VDD.n7044 240
R3182 VDD.n7496 VDD.n7495 240
R3183 VDD.n7497 VDD.n7496 240
R3184 VDD.n7497 VDD.n6419 240
R3185 VDD.n8117 VDD.n6419 240
R3186 VDD.n8117 VDD.n6420 240
R3187 VDD.n7534 VDD.n6420 240
R3188 VDD.n7534 VDD.n7019 240
R3189 VDD.n7019 VDD.n7011 240
R3190 VDD.n7575 VDD.n7011 240
R3191 VDD.n7580 VDD.n7575 240
R3192 VDD.n7580 VDD.n7579 240
R3193 VDD.n7579 VDD.n7576 240
R3194 VDD.n7576 VDD.n6961 240
R3195 VDD.n6961 VDD.n6950 240
R3196 VDD.n7656 VDD.n6950 240
R3197 VDD.n7657 VDD.n7656 240
R3198 VDD.n7659 VDD.n7657 240
R3199 VDD.n7659 VDD.n6928 240
R3200 VDD.n6928 VDD.n6915 240
R3201 VDD.n7686 VDD.n6915 240
R3202 VDD.n7686 VDD.n6919 240
R3203 VDD.n6919 VDD.n6765 240
R3204 VDD.n6777 VDD.n6765 240
R3205 VDD.n8094 VDD.n6777 240
R3206 VDD.n8094 VDD.n6778 240
R3207 VDD.n6786 VDD.n6778 240
R3208 VDD.n7944 VDD.n6786 240
R3209 VDD.n7944 VDD.n7720 240
R3210 VDD.n7937 VDD.n7720 240
R3211 VDD.n7937 VDD.n6806 240
R3212 VDD.n7738 VDD.n6806 240
R3213 VDD.n7738 VDD.n6825 240
R3214 VDD.n7927 VDD.n6825 240
R3215 VDD.n7927 VDD.n7926 240
R3216 VDD.n7926 VDD.n7742 240
R3217 VDD.n7919 VDD.n7742 240
R3218 VDD.n7919 VDD.n7918 240
R3219 VDD.n7918 VDD.n7746 240
R3220 VDD.n7914 VDD.n7746 240
R3221 VDD.n7914 VDD.n7913 240
R3222 VDD.n7913 VDD.n7912 240
R3223 VDD.n7912 VDD.n7748 240
R3224 VDD.n7776 VDD.n7748 240
R3225 VDD.n7777 VDD.n7776 240
R3226 VDD.n7778 VDD.n7777 240
R3227 VDD.n7819 VDD.n7778 240
R3228 VDD.n7819 VDD.n7783 240
R3229 VDD.n7784 VDD.n7783 240
R3230 VDD.n7785 VDD.n7784 240
R3231 VDD.n7824 VDD.n7785 240
R3232 VDD.n7824 VDD.n7790 240
R3233 VDD.n7791 VDD.n7790 240
R3234 VDD.n7792 VDD.n7791 240
R3235 VDD.n7829 VDD.n7792 240
R3236 VDD.n7829 VDD.n7797 240
R3237 VDD.n7798 VDD.n7797 240
R3238 VDD.n7799 VDD.n7798 240
R3239 VDD.n7834 VDD.n7799 240
R3240 VDD.n7834 VDD.n7804 240
R3241 VDD.n7805 VDD.n7804 240
R3242 VDD.n7181 VDD.n7172 240
R3243 VDD.n7185 VDD.n7184 240
R3244 VDD.n7189 VDD.n7188 240
R3245 VDD.n7193 VDD.n7192 240
R3246 VDD.n7197 VDD.n7196 240
R3247 VDD.n7201 VDD.n7200 240
R3248 VDD.n7205 VDD.n7204 240
R3249 VDD.n7209 VDD.n7180 240
R3250 VDD.n5361 VDD 238.556
R3251 VDD.n2614 VDD.n2613 230.966
R3252 VDD.n2613 VDD.n2603 230.966
R3253 VDD.n2606 VDD.n2603 230.966
R3254 VDD.n2933 VDD.n2932 230.966
R3255 VDD.n2932 VDD.n2922 230.966
R3256 VDD.n2925 VDD.n2922 230.966
R3257 VDD.n2908 VDD.n2907 230.966
R3258 VDD.n2907 VDD.n2745 230.966
R3259 VDD.n2828 VDD.n2786 230.966
R3260 VDD.n2829 VDD.n2828 230.966
R3261 VDD.n3134 VDD.n3125 230.966
R3262 VDD.n3135 VDD.n3134 230.966
R3263 VDD.n3143 VDD.n3135 230.966
R3264 VDD.n3143 VDD.n3142 230.966
R3265 VDD.n3142 VDD.n3136 230.966
R3266 VDD.n3202 VDD.n3201 230.966
R3267 VDD.n3201 VDD.n3183 230.966
R3268 VDD.n3187 VDD.n3183 230.966
R3269 VDD.n3191 VDD.n3187 230.966
R3270 VDD.n3191 VDD.n3190 230.966
R3271 VDD.n3623 VDD.n3622 230.966
R3272 VDD.n3622 VDD.n3604 230.966
R3273 VDD.n3608 VDD.n3604 230.966
R3274 VDD.n3612 VDD.n3608 230.966
R3275 VDD.n3612 VDD.n3611 230.966
R3276 VDD.n3483 VDD.n3482 230.966
R3277 VDD.n3482 VDD.n3464 230.966
R3278 VDD.n3468 VDD.n3464 230.966
R3279 VDD.n3472 VDD.n3468 230.966
R3280 VDD.n3472 VDD.n3471 230.966
R3281 VDD.n20 VDD.n19 230.966
R3282 VDD.n19 VDD.n9 230.966
R3283 VDD.n12 VDD.n9 230.966
R3284 VDD.n339 VDD.n338 230.966
R3285 VDD.n338 VDD.n328 230.966
R3286 VDD.n331 VDD.n328 230.966
R3287 VDD.n314 VDD.n313 230.966
R3288 VDD.n313 VDD.n151 230.966
R3289 VDD.n234 VDD.n192 230.966
R3290 VDD.n235 VDD.n234 230.966
R3291 VDD.n540 VDD.n531 230.966
R3292 VDD.n541 VDD.n540 230.966
R3293 VDD.n549 VDD.n541 230.966
R3294 VDD.n549 VDD.n548 230.966
R3295 VDD.n548 VDD.n542 230.966
R3296 VDD.n608 VDD.n607 230.966
R3297 VDD.n607 VDD.n589 230.966
R3298 VDD.n593 VDD.n589 230.966
R3299 VDD.n597 VDD.n593 230.966
R3300 VDD.n597 VDD.n596 230.966
R3301 VDD.n1029 VDD.n1028 230.966
R3302 VDD.n1028 VDD.n1010 230.966
R3303 VDD.n1014 VDD.n1010 230.966
R3304 VDD.n1018 VDD.n1014 230.966
R3305 VDD.n1018 VDD.n1017 230.966
R3306 VDD.n889 VDD.n888 230.966
R3307 VDD.n888 VDD.n870 230.966
R3308 VDD.n874 VDD.n870 230.966
R3309 VDD.n878 VDD.n874 230.966
R3310 VDD.n878 VDD.n877 230.966
R3311 VDD.n5583 VDD.n5582 230.966
R3312 VDD.n5582 VDD.n5572 230.966
R3313 VDD.n5575 VDD.n5572 230.966
R3314 VDD.n5902 VDD.n5901 230.966
R3315 VDD.n5901 VDD.n5891 230.966
R3316 VDD.n5894 VDD.n5891 230.966
R3317 VDD.n5877 VDD.n5876 230.966
R3318 VDD.n5876 VDD.n5714 230.966
R3319 VDD.n5797 VDD.n5755 230.966
R3320 VDD.n5798 VDD.n5797 230.966
R3321 VDD.n6103 VDD.n6094 230.966
R3322 VDD.n6104 VDD.n6103 230.966
R3323 VDD.n6112 VDD.n6104 230.966
R3324 VDD.n6112 VDD.n6111 230.966
R3325 VDD.n6111 VDD.n6105 230.966
R3326 VDD.n6171 VDD.n6170 230.966
R3327 VDD.n6170 VDD.n6152 230.966
R3328 VDD.n6156 VDD.n6152 230.966
R3329 VDD.n6160 VDD.n6156 230.966
R3330 VDD.n6160 VDD.n6159 230.966
R3331 VDD.n6592 VDD.n6591 230.966
R3332 VDD.n6591 VDD.n6573 230.966
R3333 VDD.n6577 VDD.n6573 230.966
R3334 VDD.n6581 VDD.n6577 230.966
R3335 VDD.n6581 VDD.n6580 230.966
R3336 VDD.n6452 VDD.n6451 230.966
R3337 VDD.n6451 VDD.n6433 230.966
R3338 VDD.n6437 VDD.n6433 230.966
R3339 VDD.n6441 VDD.n6437 230.966
R3340 VDD.n6441 VDD.n6440 230.966
R3341 VDD.t567 VDD.t563 195.589
R3342 VDD.t569 VDD.t567 195.589
R3343 VDD.t565 VDD.t232 195.589
R3344 VDD.t232 VDD.t234 195.589
R3345 VDD.t234 VDD.t236 195.589
R3346 VDD.t236 VDD.t238 195.589
R3347 VDD.t675 VDD.t673 195.589
R3348 VDD.t669 VDD.t675 195.589
R3349 VDD.t671 VDD.t669 195.589
R3350 VDD.t107 VDD.t219 195.589
R3351 VDD.t219 VDD.t134 195.589
R3352 VDD.t134 VDD.t187 195.589
R3353 VDD.t276 VDD.t352 195.589
R3354 VDD.t540 VDD.t276 195.589
R3355 VDD.t65 VDD.t540 195.589
R3356 VDD.t583 VDD.t65 195.589
R3357 VDD.t585 VDD.t587 195.589
R3358 VDD.t587 VDD.t581 195.589
R3359 VDD.t381 VDD.t14 195.589
R3360 VDD.t172 VDD.t381 195.589
R3361 VDD.t573 VDD.t172 195.589
R3362 VDD.t577 VDD.t573 195.589
R3363 VDD.t571 VDD.t575 195.589
R3364 VDD.t693 VDD.t683 195.589
R3365 VDD.t683 VDD.t689 195.589
R3366 VDD.t689 VDD.t695 195.589
R3367 VDD.t546 VDD 192.369
R3368 VDD.n3013 VDD.n2734 185
R3369 VDD.n3012 VDD.n3011 185
R3370 VDD.n3009 VDD.n2735 185
R3371 VDD.n3007 VDD.n3006 185
R3372 VDD.n3005 VDD.n2736 185
R3373 VDD.n3004 VDD.n3003 185
R3374 VDD.n3001 VDD.n2737 185
R3375 VDD.n2999 VDD.n2998 185
R3376 VDD.n2739 VDD.n2738 185
R3377 VDD.n2993 VDD.n2992 185
R3378 VDD.n2990 VDD.n2989 185
R3379 VDD.n2988 VDD.n2987 185
R3380 VDD.n2986 VDD.n2944 185
R3381 VDD.n2984 VDD.n2983 185
R3382 VDD.n2982 VDD.n2945 185
R3383 VDD.n2981 VDD.n2980 185
R3384 VDD.n2978 VDD.n2977 185
R3385 VDD.n2978 VDD.n2733 185
R3386 VDD.n2976 VDD.n2732 185
R3387 VDD.n3016 VDD.n2732 185
R3388 VDD.n2975 VDD.n2974 185
R3389 VDD.n2974 VDD.n2727 185
R3390 VDD.n2973 VDD.n2726 185
R3391 VDD.n3022 VDD.n2726 185
R3392 VDD.n2972 VDD.n2971 185
R3393 VDD.n2971 VDD.n2721 185
R3394 VDD.n2970 VDD.n2720 185
R3395 VDD.n3028 VDD.n2720 185
R3396 VDD.n2969 VDD.n2968 185
R3397 VDD.n2968 VDD.n2718 185
R3398 VDD.n2967 VDD.n2714 185
R3399 VDD.n3034 VDD.n2714 185
R3400 VDD.n2966 VDD.n2965 185
R3401 VDD.n2965 VDD.n2709 185
R3402 VDD.n2964 VDD.n2708 185
R3403 VDD.n3040 VDD.n2708 185
R3404 VDD.n2963 VDD.n2962 185
R3405 VDD.n2962 VDD.n2706 185
R3406 VDD.n2961 VDD.n2702 185
R3407 VDD.n3046 VDD.n2702 185
R3408 VDD.n2960 VDD.n2959 185
R3409 VDD.n2959 VDD.n2697 185
R3410 VDD.n2958 VDD.n2696 185
R3411 VDD.n3052 VDD.n2696 185
R3412 VDD.n2957 VDD.n2956 185
R3413 VDD.n2956 VDD.n2694 185
R3414 VDD.n2955 VDD.n2690 185
R3415 VDD.n3058 VDD.n2690 185
R3416 VDD.n2954 VDD.n2953 185
R3417 VDD.n2953 VDD.n2685 185
R3418 VDD.n2952 VDD.n2684 185
R3419 VDD.n3064 VDD.n2684 185
R3420 VDD.n2951 VDD.n2950 185
R3421 VDD.n2950 VDD.n2682 185
R3422 VDD.n2949 VDD.n2678 185
R3423 VDD.n3070 VDD.n2678 185
R3424 VDD.n2948 VDD.n2947 185
R3425 VDD.n2947 VDD.n2643 185
R3426 VDD.n2946 VDD.n2642 185
R3427 VDD.n3076 VDD.n2642 185
R3428 VDD.n2631 VDD.n2630 185
R3429 VDD.n2634 VDD.n2631 185
R3430 VDD.n3084 VDD.n3083 185
R3431 VDD.n3083 VDD.n3082 185
R3432 VDD.n3085 VDD.n2629 185
R3433 VDD.n2632 VDD.n2629 185
R3434 VDD.n3087 VDD.n3086 185
R3435 VDD.n3089 VDD.n2627 185
R3436 VDD.n3091 VDD.n3090 185
R3437 VDD.n3092 VDD.n2626 185
R3438 VDD.n3094 VDD.n3093 185
R3439 VDD.n3096 VDD.n2623 185
R3440 VDD.n3098 VDD.n3097 185
R3441 VDD.n2654 VDD.n2622 185
R3442 VDD.n2656 VDD.n2655 185
R3443 VDD.n2658 VDD.n2651 185
R3444 VDD.n2660 VDD.n2659 185
R3445 VDD.n2662 VDD.n2649 185
R3446 VDD.n2664 VDD.n2663 185
R3447 VDD.n2665 VDD.n2648 185
R3448 VDD.n2667 VDD.n2666 185
R3449 VDD.n2669 VDD.n2647 185
R3450 VDD.n2670 VDD.n2646 185
R3451 VDD.n2670 VDD.n2625 185
R3452 VDD.n2672 VDD.n2671 185
R3453 VDD.n2671 VDD.n2632 185
R3454 VDD.n2673 VDD.n2635 185
R3455 VDD.n3082 VDD.n2635 185
R3456 VDD.n2674 VDD.n2644 185
R3457 VDD.n2644 VDD.n2634 185
R3458 VDD.n3075 VDD.n3074 185
R3459 VDD.n3076 VDD.n3075 185
R3460 VDD.n3073 VDD.n2645 185
R3461 VDD.n2645 VDD.n2643 185
R3462 VDD.n3072 VDD.n3071 185
R3463 VDD.n3071 VDD.n3070 185
R3464 VDD.n2676 VDD.n2675 185
R3465 VDD.n2682 VDD.n2676 185
R3466 VDD.n3063 VDD.n3062 185
R3467 VDD.n3064 VDD.n3063 185
R3468 VDD.n3061 VDD.n2686 185
R3469 VDD.n2686 VDD.n2685 185
R3470 VDD.n3060 VDD.n3059 185
R3471 VDD.n3059 VDD.n3058 185
R3472 VDD.n2688 VDD.n2687 185
R3473 VDD.n2694 VDD.n2688 185
R3474 VDD.n3051 VDD.n3050 185
R3475 VDD.n3052 VDD.n3051 185
R3476 VDD.n3049 VDD.n2698 185
R3477 VDD.n2698 VDD.n2697 185
R3478 VDD.n3048 VDD.n3047 185
R3479 VDD.n3047 VDD.n3046 185
R3480 VDD.n2700 VDD.n2699 185
R3481 VDD.n2706 VDD.n2700 185
R3482 VDD.n3039 VDD.n3038 185
R3483 VDD.n3040 VDD.n3039 185
R3484 VDD.n3037 VDD.n2710 185
R3485 VDD.n2710 VDD.n2709 185
R3486 VDD.n3036 VDD.n3035 185
R3487 VDD.n3035 VDD.n3034 185
R3488 VDD.n2712 VDD.n2711 185
R3489 VDD.n2718 VDD.n2712 185
R3490 VDD.n3027 VDD.n3026 185
R3491 VDD.n3028 VDD.n3027 185
R3492 VDD.n3025 VDD.n2722 185
R3493 VDD.n2722 VDD.n2721 185
R3494 VDD.n3024 VDD.n3023 185
R3495 VDD.n3023 VDD.n3022 185
R3496 VDD.n2724 VDD.n2723 185
R3497 VDD.n2727 VDD.n2724 185
R3498 VDD.n3015 VDD.n3014 185
R3499 VDD.n3016 VDD.n3015 185
R3500 VDD.n2814 VDD.n2798 185
R3501 VDD.n2814 VDD.n2625 185
R3502 VDD.n2813 VDD.n2799 185
R3503 VDD.n2811 VDD.n2810 185
R3504 VDD.n2809 VDD.n2800 185
R3505 VDD.n2808 VDD.n2807 185
R3506 VDD.n2805 VDD.n2801 185
R3507 VDD.n2803 VDD.n2802 185
R3508 VDD.n2638 VDD.n2636 185
R3509 VDD.n2636 VDD.n2632 185
R3510 VDD.n3081 VDD.n3080 185
R3511 VDD.n3082 VDD.n3081 185
R3512 VDD.n3079 VDD.n2637 185
R3513 VDD.n2637 VDD.n2634 185
R3514 VDD.n3078 VDD.n3077 185
R3515 VDD.n3077 VDD.n3076 185
R3516 VDD.n2640 VDD.n2639 185
R3517 VDD.n2643 VDD.n2640 185
R3518 VDD.n3069 VDD.n3068 185
R3519 VDD.n3070 VDD.n3069 185
R3520 VDD.n3067 VDD.n2679 185
R3521 VDD.n2682 VDD.n2679 185
R3522 VDD.n3066 VDD.n3065 185
R3523 VDD.n3065 VDD.n3064 185
R3524 VDD.n2681 VDD.n2680 185
R3525 VDD.n2685 VDD.n2681 185
R3526 VDD.n3057 VDD.n3056 185
R3527 VDD.n3058 VDD.n3057 185
R3528 VDD.n3055 VDD.n2691 185
R3529 VDD.n2694 VDD.n2691 185
R3530 VDD.n3054 VDD.n3053 185
R3531 VDD.n3053 VDD.n3052 185
R3532 VDD.n2693 VDD.n2692 185
R3533 VDD.n2697 VDD.n2693 185
R3534 VDD.n3045 VDD.n3044 185
R3535 VDD.n3046 VDD.n3045 185
R3536 VDD.n3043 VDD.n2703 185
R3537 VDD.n2706 VDD.n2703 185
R3538 VDD.n3042 VDD.n3041 185
R3539 VDD.n3041 VDD.n3040 185
R3540 VDD.n2705 VDD.n2704 185
R3541 VDD.n2709 VDD.n2705 185
R3542 VDD.n3033 VDD.n3032 185
R3543 VDD.n3034 VDD.n3033 185
R3544 VDD.n3031 VDD.n2715 185
R3545 VDD.n2718 VDD.n2715 185
R3546 VDD.n3030 VDD.n3029 185
R3547 VDD.n3029 VDD.n3028 185
R3548 VDD.n2717 VDD.n2716 185
R3549 VDD.n2721 VDD.n2717 185
R3550 VDD.n3021 VDD.n3020 185
R3551 VDD.n3022 VDD.n3021 185
R3552 VDD.n3019 VDD.n2728 185
R3553 VDD.n2728 VDD.n2727 185
R3554 VDD.n3018 VDD.n3017 185
R3555 VDD.n3017 VDD.n3016 185
R3556 VDD.n2730 VDD.n2729 185
R3557 VDD.n2761 VDD.n2760 185
R3558 VDD.n2762 VDD.n2758 185
R3559 VDD.n2758 VDD.n2733 185
R3560 VDD.n2764 VDD.n2763 185
R3561 VDD.n2766 VDD.n2757 185
R3562 VDD.n2769 VDD.n2768 185
R3563 VDD.n2770 VDD.n2756 185
R3564 VDD.n2772 VDD.n2771 185
R3565 VDD.n2774 VDD.n2749 185
R3566 VDD.n2901 VDD.n2900 185
R3567 VDD.n2898 VDD.n2897 185
R3568 VDD.n2896 VDD.n2775 185
R3569 VDD.n2895 VDD.n2894 185
R3570 VDD.n2892 VDD.n2776 185
R3571 VDD.n2890 VDD.n2889 185
R3572 VDD.n2888 VDD.n2777 185
R3573 VDD.n2887 VDD.n2886 185
R3574 VDD.n2884 VDD.n2731 185
R3575 VDD.n3016 VDD.n2731 185
R3576 VDD.n2883 VDD.n2882 185
R3577 VDD.n2882 VDD.n2727 185
R3578 VDD.n2881 VDD.n2725 185
R3579 VDD.n3022 VDD.n2725 185
R3580 VDD.n2880 VDD.n2879 185
R3581 VDD.n2879 VDD.n2721 185
R3582 VDD.n2878 VDD.n2719 185
R3583 VDD.n3028 VDD.n2719 185
R3584 VDD.n2877 VDD.n2876 185
R3585 VDD.n2876 VDD.n2718 185
R3586 VDD.n2875 VDD.n2713 185
R3587 VDD.n3034 VDD.n2713 185
R3588 VDD.n2874 VDD.n2873 185
R3589 VDD.n2873 VDD.n2709 185
R3590 VDD.n2872 VDD.n2707 185
R3591 VDD.n3040 VDD.n2707 185
R3592 VDD.n2871 VDD.n2870 185
R3593 VDD.n2870 VDD.n2706 185
R3594 VDD.n2869 VDD.n2701 185
R3595 VDD.n3046 VDD.n2701 185
R3596 VDD.n2868 VDD.n2867 185
R3597 VDD.n2867 VDD.n2697 185
R3598 VDD.n2866 VDD.n2695 185
R3599 VDD.n3052 VDD.n2695 185
R3600 VDD.n2865 VDD.n2864 185
R3601 VDD.n2864 VDD.n2694 185
R3602 VDD.n2863 VDD.n2689 185
R3603 VDD.n3058 VDD.n2689 185
R3604 VDD.n2862 VDD.n2861 185
R3605 VDD.n2861 VDD.n2685 185
R3606 VDD.n2860 VDD.n2683 185
R3607 VDD.n3064 VDD.n2683 185
R3608 VDD.n2859 VDD.n2858 185
R3609 VDD.n2858 VDD.n2682 185
R3610 VDD.n2857 VDD.n2677 185
R3611 VDD.n3070 VDD.n2677 185
R3612 VDD.n2856 VDD.n2855 185
R3613 VDD.n2855 VDD.n2643 185
R3614 VDD.n2854 VDD.n2641 185
R3615 VDD.n3076 VDD.n2641 185
R3616 VDD.n2853 VDD.n2852 185
R3617 VDD.n2852 VDD.n2634 185
R3618 VDD.n2851 VDD.n2633 185
R3619 VDD.n3082 VDD.n2633 185
R3620 VDD.n2850 VDD.n2849 185
R3621 VDD.n2849 VDD.n2632 185
R3622 VDD.n2848 VDD.n2778 185
R3623 VDD.n2846 VDD.n2845 185
R3624 VDD.n2844 VDD.n2779 185
R3625 VDD.n2843 VDD.n2842 185
R3626 VDD.n2840 VDD.n2780 185
R3627 VDD.n2838 VDD.n2837 185
R3628 VDD.n2836 VDD.n2781 185
R3629 VDD.n2819 VDD.n2782 185
R3630 VDD.n2822 VDD.n2821 185
R3631 VDD.n2823 VDD.n2815 185
R3632 VDD.n5070 VDD.n3890 185
R3633 VDD.n5069 VDD.n5068 185
R3634 VDD.n3892 VDD.n3891 185
R3635 VDD.n5001 VDD.n5000 185
R3636 VDD.n5003 VDD.n5002 185
R3637 VDD.n5005 VDD.n5004 185
R3638 VDD.n5007 VDD.n5006 185
R3639 VDD.n5009 VDD.n5008 185
R3640 VDD.n5011 VDD.n5010 185
R3641 VDD.n5013 VDD.n5012 185
R3642 VDD.n5015 VDD.n5014 185
R3643 VDD.n5017 VDD.n5016 185
R3644 VDD.n5019 VDD.n5018 185
R3645 VDD.n5021 VDD.n5020 185
R3646 VDD.n5023 VDD.n5022 185
R3647 VDD.n5025 VDD.n5024 185
R3648 VDD.n5026 VDD.n3907 185
R3649 VDD.n5066 VDD.n3907 185
R3650 VDD.n5027 VDD.n3888 185
R3651 VDD.n5073 VDD.n3888 185
R3652 VDD.n5029 VDD.n5028 185
R3653 VDD.n5030 VDD.n5029 185
R3654 VDD.n4999 VDD.n3882 185
R3655 VDD.n5079 VDD.n3882 185
R3656 VDD.n4998 VDD.n4997 185
R3657 VDD.n4997 VDD.n4996 185
R3658 VDD.n3912 VDD.n3869 185
R3659 VDD.n5085 VDD.n3869 185
R3660 VDD.n4989 VDD.n4988 185
R3661 VDD.n4990 VDD.n4989 185
R3662 VDD.n4987 VDD.n3858 185
R3663 VDD.n5091 VDD.n3858 185
R3664 VDD.n4986 VDD.n4985 185
R3665 VDD.n4985 VDD.n3855 185
R3666 VDD.n4984 VDD.n4983 185
R3667 VDD.n4984 VDD.n3838 185
R3668 VDD.n4982 VDD.n3836 185
R3669 VDD.n5102 VDD.n3836 185
R3670 VDD.n4981 VDD.n3828 185
R3671 VDD.n5108 VDD.n3828 185
R3672 VDD.n4980 VDD.n4979 185
R3673 VDD.n4979 VDD.n4978 185
R3674 VDD.n4750 VDD.n3819 185
R3675 VDD.n5114 VDD.n3819 185
R3676 VDD.n4749 VDD.n4748 185
R3677 VDD.n4748 VDD.n4747 185
R3678 VDD.n3919 VDD.n3918 185
R3679 VDD.n3919 VDD.n3810 185
R3680 VDD.n4738 VDD.n4737 185
R3681 VDD.n4739 VDD.n4738 185
R3682 VDD.n4736 VDD.n3798 185
R3683 VDD.n5133 VDD.n3798 185
R3684 VDD.n4735 VDD.n4734 185
R3685 VDD.n4734 VDD.n4733 185
R3686 VDD.n3926 VDD.n3925 185
R3687 VDD.n3952 VDD.n3926 185
R3688 VDD.n4702 VDD.n3935 185
R3689 VDD.n4725 VDD.n3935 185
R3690 VDD.n4704 VDD.n4703 185
R3691 VDD.n4705 VDD.n4704 185
R3692 VDD.n4701 VDD.n3961 185
R3693 VDD.n3961 VDD.n3958 185
R3694 VDD.n4700 VDD.n4699 185
R3695 VDD.n4699 VDD.n4698 185
R3696 VDD.n3963 VDD.n3962 185
R3697 VDD.n3984 VDD.n3963 185
R3698 VDD.n4644 VDD.n4643 185
R3699 VDD.n4645 VDD.n4644 185
R3700 VDD.n4642 VDD.n3994 185
R3701 VDD.n4671 VDD.n3994 185
R3702 VDD.n4641 VDD.n4640 185
R3703 VDD.n4640 VDD.n4639 185
R3704 VDD.n4019 VDD.n4008 185
R3705 VDD.n4652 VDD.n4008 185
R3706 VDD.n4624 VDD.n4623 185
R3707 VDD.t629 VDD.n4624 185
R3708 VDD.n4622 VDD.n4024 185
R3709 VDD.n4043 VDD.n4024 185
R3710 VDD.n4621 VDD.n4620 185
R3711 VDD.n4620 VDD.n4619 185
R3712 VDD.n4026 VDD.n4025 185
R3713 VDD.n4586 VDD.n4026 185
R3714 VDD.n4544 VDD.n4058 185
R3715 VDD.n4577 VDD.n4058 185
R3716 VDD.n4546 VDD.n4545 185
R3717 VDD.n4549 VDD.n4546 185
R3718 VDD.n4543 VDD.n4060 185
R3719 VDD.n4060 VDD.n3452 185
R3720 VDD.n4542 VDD.n3441 185
R3721 VDD.n5156 VDD.n3441 185
R3722 VDD.n4541 VDD.n4540 185
R3723 VDD.n4540 VDD.n4539 185
R3724 VDD.n4062 VDD.n4061 185
R3725 VDD.n4536 VDD.n4062 185
R3726 VDD.n4488 VDD.n4105 185
R3727 VDD.n4105 VDD.n4078 185
R3728 VDD.n4490 VDD.n4489 185
R3729 VDD.n4491 VDD.n4490 185
R3730 VDD.n4487 VDD.n4088 185
R3731 VDD.n4506 VDD.n4088 185
R3732 VDD.n4486 VDD.n4485 185
R3733 VDD.n4485 VDD.n4484 185
R3734 VDD.n4106 VDD.n4096 185
R3735 VDD.n4499 VDD.n4096 185
R3736 VDD.n4477 VDD.n4476 185
R3737 VDD.n4478 VDD.n4477 185
R3738 VDD.n4475 VDD.n4111 185
R3739 VDD.n4458 VDD.n4111 185
R3740 VDD.n4474 VDD.n4473 185
R3741 VDD.n4473 VDD.n4472 185
R3742 VDD.n4113 VDD.n4112 185
R3743 VDD.n4438 VDD.n4113 185
R3744 VDD.n4428 VDD.n4123 185
R3745 VDD.n4465 VDD.n4123 185
R3746 VDD.n4430 VDD.n4429 185
R3747 VDD.n4431 VDD.n4430 185
R3748 VDD.n4427 VDD.n4139 185
R3749 VDD.n4386 VDD.n4139 185
R3750 VDD.n4426 VDD.n4425 185
R3751 VDD.n4141 VDD.n4140 185
R3752 VDD.n4356 VDD.n4355 185
R3753 VDD.n4358 VDD.n4357 185
R3754 VDD.n4360 VDD.n4359 185
R3755 VDD.n4362 VDD.n4361 185
R3756 VDD.n4364 VDD.n4363 185
R3757 VDD.n4366 VDD.n4365 185
R3758 VDD.n4368 VDD.n4367 185
R3759 VDD.n4370 VDD.n4369 185
R3760 VDD.n4372 VDD.n4371 185
R3761 VDD.n4374 VDD.n4373 185
R3762 VDD.n4376 VDD.n4375 185
R3763 VDD.n4378 VDD.n4377 185
R3764 VDD.n4380 VDD.n4379 185
R3765 VDD.n4382 VDD.n4381 185
R3766 VDD.n4383 VDD.n4143 185
R3767 VDD.n4423 VDD.n4143 185
R3768 VDD.n4385 VDD.n4384 185
R3769 VDD.n4386 VDD.n4385 185
R3770 VDD.n4126 VDD.n4124 185
R3771 VDD.n4431 VDD.n4124 185
R3772 VDD.n4464 VDD.n4463 185
R3773 VDD.n4465 VDD.n4464 185
R3774 VDD.n4462 VDD.n4125 185
R3775 VDD.n4438 VDD.n4125 185
R3776 VDD.n4461 VDD.n4116 185
R3777 VDD.n4472 VDD.n4116 185
R3778 VDD.n4460 VDD.n4459 185
R3779 VDD.n4459 VDD.n4458 185
R3780 VDD.n4099 VDD.n4097 185
R3781 VDD.n4478 VDD.n4097 185
R3782 VDD.n4498 VDD.n4497 185
R3783 VDD.n4499 VDD.n4498 185
R3784 VDD.n4496 VDD.n4098 185
R3785 VDD.n4484 VDD.n4098 185
R3786 VDD.n4495 VDD.n4089 185
R3787 VDD.n4506 VDD.n4089 185
R3788 VDD.n4493 VDD.n4101 185
R3789 VDD.n4491 VDD.n4101 185
R3790 VDD.n4102 VDD.n4064 185
R3791 VDD.n4078 VDD.n4064 185
R3792 VDD.n4537 VDD.n4065 185
R3793 VDD.n4537 VDD.n4536 185
R3794 VDD.n4538 VDD.n3435 185
R3795 VDD.n4539 VDD.n4538 185
R3796 VDD.n5158 VDD.n3436 185
R3797 VDD.n5156 VDD.n3436 185
R3798 VDD.n4547 VDD.n3437 185
R3799 VDD.n4547 VDD.n3452 185
R3800 VDD.n4548 VDD.n4055 185
R3801 VDD.n4549 VDD.n4548 185
R3802 VDD.n4579 VDD.n4052 185
R3803 VDD.n4577 VDD.n4052 185
R3804 VDD.n4585 VDD.n4584 185
R3805 VDD.n4586 VDD.n4585 185
R3806 VDD.n4583 VDD.n4029 185
R3807 VDD.n4619 VDD.n4029 185
R3808 VDD.n4582 VDD.n4581 185
R3809 VDD.n4581 VDD.n4043 185
R3810 VDD.n4011 VDD.n4009 185
R3811 VDD.t629 VDD.n4009 185
R3812 VDD.n4651 VDD.n4650 185
R3813 VDD.n4652 VDD.n4651 185
R3814 VDD.n4649 VDD.n4010 185
R3815 VDD.n4639 VDD.n4010 185
R3816 VDD.n4648 VDD.n3995 185
R3817 VDD.n4671 VDD.n3995 185
R3818 VDD.n4647 VDD.n4646 185
R3819 VDD.n4646 VDD.n4645 185
R3820 VDD.n4016 VDD.n4015 185
R3821 VDD.n4016 VDD.n3984 185
R3822 VDD.n4014 VDD.n3966 185
R3823 VDD.n4698 VDD.n3966 185
R3824 VDD.n4013 VDD.n4012 185
R3825 VDD.n4012 VDD.n3958 185
R3826 VDD.n3932 VDD.n3931 185
R3827 VDD.n4705 VDD.n3932 185
R3828 VDD.n4727 VDD.n4726 185
R3829 VDD.n4726 VDD.n4725 185
R3830 VDD.n4728 VDD.n3929 185
R3831 VDD.n3952 VDD.n3929 185
R3832 VDD.n4732 VDD.n4731 185
R3833 VDD.n4733 VDD.n4732 185
R3834 VDD.n4730 VDD.n3799 185
R3835 VDD.n5133 VDD.n3799 185
R3836 VDD.n3923 VDD.n3922 185
R3837 VDD.n4739 VDD.n3922 185
R3838 VDD.n4743 VDD.n4742 185
R3839 VDD.n4743 VDD.n3810 185
R3840 VDD.n4746 VDD.n4745 185
R3841 VDD.n4747 VDD.n4746 185
R3842 VDD.n4744 VDD.n3820 185
R3843 VDD.n5114 VDD.n3820 185
R3844 VDD.n3831 VDD.n3829 185
R3845 VDD.n4978 VDD.n3829 185
R3846 VDD.n5107 VDD.n5106 185
R3847 VDD.n5108 VDD.n5107 185
R3848 VDD.n3832 VDD.n3830 185
R3849 VDD.n5102 VDD.n3830 185
R3850 VDD.n3873 VDD.n3872 185
R3851 VDD.n3873 VDD.n3838 185
R3852 VDD.n3875 VDD.n3874 185
R3853 VDD.n3874 VDD.n3855 185
R3854 VDD.n3876 VDD.n3859 185
R3855 VDD.n5091 VDD.n3859 185
R3856 VDD.n3877 VDD.n3870 185
R3857 VDD.n4990 VDD.n3870 185
R3858 VDD.n5084 VDD.n5083 185
R3859 VDD.n5085 VDD.n5084 185
R3860 VDD.n5082 VDD.n3871 185
R3861 VDD.n4996 VDD.n3871 185
R3862 VDD.n5081 VDD.n5080 185
R3863 VDD.n5080 VDD.n5079 185
R3864 VDD.n3879 VDD.n3878 185
R3865 VDD.n5030 VDD.n3879 185
R3866 VDD.n5072 VDD.n5071 185
R3867 VDD.n5073 VDD.n5072 185
R3868 VDD.n3885 VDD.n3884 185
R3869 VDD.n5064 VDD.n5063 185
R3870 VDD.n5062 VDD.n3909 185
R3871 VDD.n5066 VDD.n3909 185
R3872 VDD.n5061 VDD.n5060 185
R3873 VDD.n5059 VDD.n5058 185
R3874 VDD.n5057 VDD.n5056 185
R3875 VDD.n5055 VDD.n5054 185
R3876 VDD.n5053 VDD.n5052 185
R3877 VDD.n5051 VDD.n5050 185
R3878 VDD.n5049 VDD.n5048 185
R3879 VDD.n5047 VDD.n5046 185
R3880 VDD.n5045 VDD.n5044 185
R3881 VDD.n5043 VDD.n5042 185
R3882 VDD.n5041 VDD.n5040 185
R3883 VDD.n5039 VDD.n5038 185
R3884 VDD.n5037 VDD.n5036 185
R3885 VDD.n5035 VDD.n5034 185
R3886 VDD.n5033 VDD.n3887 185
R3887 VDD.n5073 VDD.n3887 185
R3888 VDD.n5032 VDD.n5031 185
R3889 VDD.n5031 VDD.n5030 185
R3890 VDD.n3910 VDD.n3881 185
R3891 VDD.n5079 VDD.n3881 185
R3892 VDD.n4995 VDD.n4994 185
R3893 VDD.n4996 VDD.n4995 185
R3894 VDD.n4993 VDD.n3868 185
R3895 VDD.n5085 VDD.n3868 185
R3896 VDD.n4992 VDD.n4991 185
R3897 VDD.n4991 VDD.n4990 185
R3898 VDD.n3916 VDD.n3857 185
R3899 VDD.n5091 VDD.n3857 185
R3900 VDD.n3915 VDD.n3914 185
R3901 VDD.n3914 VDD.n3855 185
R3902 VDD.n3834 VDD.n3833 185
R3903 VDD.n3838 VDD.n3834 185
R3904 VDD.n5104 VDD.n5103 185
R3905 VDD.n5103 VDD.n5102 185
R3906 VDD.n5106 VDD.n3827 185
R3907 VDD.n5108 VDD.n3827 185
R3908 VDD.n4977 VDD.n3831 185
R3909 VDD.n4978 VDD.n4977 185
R3910 VDD.n4744 VDD.n3818 185
R3911 VDD.n5114 VDD.n3818 185
R3912 VDD.n4745 VDD.n3921 185
R3913 VDD.n4747 VDD.n3921 185
R3914 VDD.n4742 VDD.n4741 185
R3915 VDD.n4741 VDD.n3810 185
R3916 VDD.n4740 VDD.n3923 185
R3917 VDD.n4740 VDD.n4739 185
R3918 VDD.n4730 VDD.n3797 185
R3919 VDD.n5133 VDD.n3797 185
R3920 VDD.n4731 VDD.n3928 185
R3921 VDD.n4733 VDD.n3928 185
R3922 VDD.n3951 VDD.n3930 185
R3923 VDD.n3952 VDD.n3951 185
R3924 VDD.n4628 VDD.n3934 185
R3925 VDD.n4725 VDD.n3934 185
R3926 VDD.n4629 VDD.n3960 185
R3927 VDD.n4705 VDD.n3960 185
R3928 VDD.n4631 VDD.n4630 185
R3929 VDD.n4630 VDD.n3958 185
R3930 VDD.n4632 VDD.n3965 185
R3931 VDD.n4698 VDD.n3965 185
R3932 VDD.n4634 VDD.n4633 185
R3933 VDD.n4633 VDD.n3984 185
R3934 VDD.n4635 VDD.n4018 185
R3935 VDD.n4645 VDD.n4018 185
R3936 VDD.n4636 VDD.n3993 185
R3937 VDD.n4671 VDD.n3993 185
R3938 VDD.n4638 VDD.n4637 185
R3939 VDD.n4639 VDD.n4638 185
R3940 VDD.n4627 VDD.n4007 185
R3941 VDD.n4652 VDD.n4007 185
R3942 VDD.n4626 VDD.n4625 185
R3943 VDD.n4625 VDD.t629 185
R3944 VDD.n4022 VDD.n4021 185
R3945 VDD.n4043 VDD.n4022 185
R3946 VDD.n4053 VDD.n4028 185
R3947 VDD.n4619 VDD.n4028 185
R3948 VDD.n4054 VDD.n4051 185
R3949 VDD.n4586 VDD.n4051 185
R3950 VDD.n4579 VDD.n4578 185
R3951 VDD.n4578 VDD.n4577 185
R3952 VDD.n4056 VDD.n4055 185
R3953 VDD.n4549 VDD.n4056 185
R3954 VDD.n3439 VDD.n3437 185
R3955 VDD.n3452 VDD.n3439 185
R3956 VDD.n5158 VDD.n5157 185
R3957 VDD.n5157 VDD.n5156 185
R3958 VDD.n3438 VDD.n3435 185
R3959 VDD.n4539 VDD.n3438 185
R3960 VDD.n4067 VDD.n4065 185
R3961 VDD.n4536 VDD.n4067 185
R3962 VDD.n4103 VDD.n4102 185
R3963 VDD.n4103 VDD.n4078 185
R3964 VDD.n4493 VDD.n4492 185
R3965 VDD.n4492 VDD.n4491 185
R3966 VDD.n4100 VDD.n4087 185
R3967 VDD.n4506 VDD.n4087 185
R3968 VDD.n4483 VDD.n4482 185
R3969 VDD.n4484 VDD.n4483 185
R3970 VDD.n4481 VDD.n4095 185
R3971 VDD.n4499 VDD.n4095 185
R3972 VDD.n4480 VDD.n4479 185
R3973 VDD.n4479 VDD.n4478 185
R3974 VDD.n4109 VDD.n4108 185
R3975 VDD.n4458 VDD.n4109 185
R3976 VDD.n4435 VDD.n4115 185
R3977 VDD.n4472 VDD.n4115 185
R3978 VDD.n4437 VDD.n4436 185
R3979 VDD.n4438 VDD.n4437 185
R3980 VDD.n4434 VDD.n4122 185
R3981 VDD.n4465 VDD.n4122 185
R3982 VDD.n4433 VDD.n4432 185
R3983 VDD.n4432 VDD.n4431 185
R3984 VDD.n4137 VDD.n4136 185
R3985 VDD.n4386 VDD.n4137 185
R3986 VDD.n4391 VDD.n4390 185
R3987 VDD.n4393 VDD.n4392 185
R3988 VDD.n4395 VDD.n4394 185
R3989 VDD.n4397 VDD.n4396 185
R3990 VDD.n4399 VDD.n4398 185
R3991 VDD.n4401 VDD.n4400 185
R3992 VDD.n4403 VDD.n4402 185
R3993 VDD.n4405 VDD.n4404 185
R3994 VDD.n4407 VDD.n4406 185
R3995 VDD.n4409 VDD.n4408 185
R3996 VDD.n4411 VDD.n4410 185
R3997 VDD.n4413 VDD.n4412 185
R3998 VDD.n4415 VDD.n4414 185
R3999 VDD.n4417 VDD.n4416 185
R4000 VDD.n4419 VDD.n4418 185
R4001 VDD.n4420 VDD.n4388 185
R4002 VDD.n4422 VDD.n4421 185
R4003 VDD.n4423 VDD.n4422 185
R4004 VDD.n4389 VDD.n4387 185
R4005 VDD.n4387 VDD.n4386 185
R4006 VDD.n4120 VDD.n4119 185
R4007 VDD.n4431 VDD.n4120 185
R4008 VDD.n4467 VDD.n4466 185
R4009 VDD.n4466 VDD.n4465 185
R4010 VDD.n4468 VDD.n4117 185
R4011 VDD.n4438 VDD.n4117 185
R4012 VDD.n4471 VDD.n4470 185
R4013 VDD.n4472 VDD.n4471 185
R4014 VDD.n4469 VDD.n4118 185
R4015 VDD.n4458 VDD.n4118 185
R4016 VDD.n4093 VDD.n4092 185
R4017 VDD.n4478 VDD.n4093 185
R4018 VDD.n4501 VDD.n4500 185
R4019 VDD.n4500 VDD.n4499 185
R4020 VDD.n4502 VDD.n4090 185
R4021 VDD.n4484 VDD.n4090 185
R4022 VDD.n4505 VDD.n4504 185
R4023 VDD.n4506 VDD.n4505 185
R4024 VDD.n4503 VDD.n4091 185
R4025 VDD.n4491 VDD.n4091 185
R4026 VDD.n4069 VDD.n4068 185
R4027 VDD.n4078 VDD.n4068 185
R4028 VDD.n4535 VDD.n4534 185
R4029 VDD.n4536 VDD.n4535 185
R4030 VDD.n4070 VDD.n3442 185
R4031 VDD.n4539 VDD.n3442 185
R4032 VDD.n5155 VDD.n5154 185
R4033 VDD.n5156 VDD.n5155 185
R4034 VDD.n3445 VDD.n3443 185
R4035 VDD.n3452 VDD.n3443 185
R4036 VDD.n4552 VDD.n4550 185
R4037 VDD.n4550 VDD.n4549 185
R4038 VDD.n4576 VDD.n4575 185
R4039 VDD.n4577 VDD.n4576 185
R4040 VDD.n4554 VDD.n4030 185
R4041 VDD.n4586 VDD.n4030 185
R4042 VDD.n4618 VDD.n4617 185
R4043 VDD.n4619 VDD.n4618 185
R4044 VDD.n4033 VDD.n4031 185
R4045 VDD.n4043 VDD.n4031 185
R4046 VDD.n4035 VDD.n4005 185
R4047 VDD.t629 VDD.n4005 185
R4048 VDD.n4654 VDD.n4653 185
R4049 VDD.n4653 VDD.n4652 185
R4050 VDD.n4655 VDD.n3996 185
R4051 VDD.n4639 VDD.n3996 185
R4052 VDD.n4670 VDD.n4669 185
R4053 VDD.n4671 VDD.n4670 185
R4054 VDD.n4668 VDD.n3997 185
R4055 VDD.n4645 VDD.n3997 185
R4056 VDD.n3999 VDD.n3967 185
R4057 VDD.n3984 VDD.n3967 185
R4058 VDD.n4697 VDD.n4696 185
R4059 VDD.n4698 VDD.n4697 185
R4060 VDD.n3970 VDD.n3968 185
R4061 VDD.n3968 VDD.n3958 185
R4062 VDD.n3972 VDD.n3936 185
R4063 VDD.n4705 VDD.n3936 185
R4064 VDD.n4724 VDD.n4723 185
R4065 VDD.n4725 VDD.n4724 185
R4066 VDD.n3939 VDD.n3937 185
R4067 VDD.n3952 VDD.n3937 185
R4068 VDD.n3941 VDD.n3800 185
R4069 VDD.n4733 VDD.n3800 185
R4070 VDD.n5132 VDD.n5131 185
R4071 VDD.n5133 VDD.n5132 185
R4072 VDD.n3803 VDD.n3801 185
R4073 VDD.n4739 VDD.n3801 185
R4074 VDD.n4757 VDD.n4756 185
R4075 VDD.n4756 VDD.n3810 185
R4076 VDD.n4758 VDD.n3821 185
R4077 VDD.n4747 VDD.n3821 185
R4078 VDD.n5113 VDD.n5112 185
R4079 VDD.n5114 VDD.n5113 185
R4080 VDD.n5111 VDD.n3822 185
R4081 VDD.n4978 VDD.n3822 185
R4082 VDD.n5110 VDD.n5109 185
R4083 VDD.n5109 VDD.n5108 185
R4084 VDD.n3825 VDD.n3824 185
R4085 VDD.n5102 VDD.n3825 185
R4086 VDD.n3863 VDD.n3862 185
R4087 VDD.n3862 VDD.n3838 185
R4088 VDD.n3864 VDD.n3860 185
R4089 VDD.n3860 VDD.n3855 185
R4090 VDD.n5090 VDD.n5089 185
R4091 VDD.n5091 VDD.n5090 185
R4092 VDD.n5088 VDD.n3861 185
R4093 VDD.n4990 VDD.n3861 185
R4094 VDD.n5087 VDD.n5086 185
R4095 VDD.n5086 VDD.n5085 185
R4096 VDD.n3866 VDD.n3865 185
R4097 VDD.n4996 VDD.n3866 185
R4098 VDD.n5078 VDD.n5077 185
R4099 VDD.n5079 VDD.n5078 185
R4100 VDD.n5076 VDD.n3883 185
R4101 VDD.n5030 VDD.n3883 185
R4102 VDD.n5075 VDD.n5074 185
R4103 VDD.n5074 VDD.n5073 185
R4104 VDD.n4240 VDD.n4239 185
R4105 VDD.n4241 VDD.n4240 185
R4106 VDD.n4238 VDD.n4211 185
R4107 VDD.n4237 VDD.n4236 185
R4108 VDD.n4235 VDD.n4234 185
R4109 VDD.n4233 VDD.n4232 185
R4110 VDD.n4231 VDD.n4230 185
R4111 VDD.n4229 VDD.n4228 185
R4112 VDD.n4227 VDD.n4226 185
R4113 VDD.n4225 VDD.n4224 185
R4114 VDD.n4223 VDD.n4222 185
R4115 VDD.n4221 VDD.n4220 185
R4116 VDD.n4219 VDD.n4218 185
R4117 VDD.n4217 VDD.n4216 185
R4118 VDD.n4215 VDD.n4214 185
R4119 VDD.n4213 VDD.n4212 185
R4120 VDD.n4203 VDD.n4202 185
R4121 VDD.n4244 VDD.n4243 185
R4122 VDD.n4245 VDD.n4201 185
R4123 VDD.n4201 VDD.n4200 185
R4124 VDD.n4247 VDD.n4246 185
R4125 VDD.n4248 VDD.n4247 185
R4126 VDD.n4195 VDD.n4194 185
R4127 VDD.n4196 VDD.n4195 185
R4128 VDD.n4256 VDD.n4255 185
R4129 VDD.n4255 VDD.n4254 185
R4130 VDD.n4257 VDD.n4193 185
R4131 VDD.n4193 VDD.n4192 185
R4132 VDD.n4259 VDD.n4258 185
R4133 VDD.n4260 VDD.n4259 185
R4134 VDD.n4187 VDD.n4186 185
R4135 VDD.n4188 VDD.n4187 185
R4136 VDD.n4269 VDD.n4268 185
R4137 VDD.n4268 VDD.n4267 185
R4138 VDD.n4270 VDD.n4185 185
R4139 VDD.n4266 VDD.n4185 185
R4140 VDD.n4272 VDD.n4271 185
R4141 VDD.n4273 VDD.n4272 185
R4142 VDD.n4180 VDD.n4179 185
R4143 VDD.n4184 VDD.n4180 185
R4144 VDD.n4282 VDD.n4281 185
R4145 VDD.n4281 VDD.n4280 185
R4146 VDD.n4283 VDD.n4178 185
R4147 VDD.n4279 VDD.n4178 185
R4148 VDD.n4285 VDD.n4284 185
R4149 VDD.n4286 VDD.n4285 185
R4150 VDD.n4173 VDD.n4172 185
R4151 VDD.n4174 VDD.n4173 185
R4152 VDD.n4294 VDD.n4293 185
R4153 VDD.n4293 VDD.n4292 185
R4154 VDD.n4295 VDD.n4171 185
R4155 VDD.n4171 VDD.n4170 185
R4156 VDD.n4298 VDD.n4297 185
R4157 VDD.n4299 VDD.n4298 185
R4158 VDD.n4296 VDD.n4164 185
R4159 VDD.n4165 VDD.n4164 185
R4160 VDD.n4345 VDD.n4163 185
R4161 VDD.n4345 VDD.n4344 185
R4162 VDD.n4347 VDD.n4346 185
R4163 VDD.n4346 VDD.n4142 185
R4164 VDD.n4348 VDD.n4161 185
R4165 VDD.n4161 VDD.n4151 185
R4166 VDD.n4353 VDD.n4352 185
R4167 VDD.n4354 VDD.n4353 185
R4168 VDD.n4351 VDD.n4162 185
R4169 VDD.n4162 VDD.n4138 185
R4170 VDD.n4349 VDD.n4134 185
R4171 VDD.n4134 VDD.n4121 185
R4172 VDD.n4441 VDD.n4440 185
R4173 VDD.n4440 VDD.n4439 185
R4174 VDD.n4442 VDD.n4128 185
R4175 VDD.n4128 VDD.n4114 185
R4176 VDD.n4456 VDD.n4455 185
R4177 VDD.n4457 VDD.n4456 185
R4178 VDD.n4131 VDD.n4129 185
R4179 VDD.n4129 VDD.n4110 185
R4180 VDD.n4450 VDD.n4449 185
R4181 VDD.n4449 VDD.n4094 185
R4182 VDD.n4447 VDD.n4085 185
R4183 VDD.n4107 VDD.n4085 185
R4184 VDD.n4509 VDD.n4508 185
R4185 VDD.n4508 VDD.n4507 185
R4186 VDD.n4510 VDD.n4079 185
R4187 VDD.n4104 VDD.n4079 185
R4188 VDD.n4524 VDD.n4523 185
R4189 VDD.n4525 VDD.n4524 185
R4190 VDD.n4082 VDD.n4080 185
R4191 VDD.n4080 VDD.n4066 185
R4192 VDD.n4518 VDD.n4517 185
R4193 VDD.n4517 VDD.n4063 185
R4194 VDD.n4515 VDD.n3453 185
R4195 VDD.n3453 VDD.n3440 185
R4196 VDD.n5146 VDD.n5145 185
R4197 VDD.n5147 VDD.n5146 185
R4198 VDD.n5144 VDD.n3454 185
R4199 VDD.n4059 VDD.n3454 185
R4200 VDD.n4049 VDD.n3456 185
R4201 VDD.n4057 VDD.n4049 185
R4202 VDD.n4589 VDD.n4588 185
R4203 VDD.n4588 VDD.n4587 185
R4204 VDD.n4590 VDD.n4044 185
R4205 VDD.n4044 VDD.n4027 185
R4206 VDD.n4604 VDD.n4603 185
R4207 VDD.n4605 VDD.n4604 185
R4208 VDD.n4047 VDD.n4045 185
R4209 VDD.n4045 VDD.n4023 185
R4210 VDD.n4598 VDD.n4597 185
R4211 VDD.n4597 VDD.n4006 185
R4212 VDD.n4595 VDD.n3991 185
R4213 VDD.n4020 VDD.n3991 185
R4214 VDD.n4674 VDD.n4673 185
R4215 VDD.n4673 VDD.n4672 185
R4216 VDD.n4675 VDD.n3985 185
R4217 VDD.n4017 VDD.n3985 185
R4218 VDD.n4685 VDD.n4684 185
R4219 VDD.n4686 VDD.n4685 185
R4220 VDD.n3988 VDD.n3986 185
R4221 VDD.n3986 VDD.n3964 185
R4222 VDD.n4679 VDD.n3957 185
R4223 VDD.n4689 VDD.n3957 185
R4224 VDD.n4708 VDD.n4707 185
R4225 VDD.n4707 VDD.n4706 185
R4226 VDD.n3954 VDD.n3953 185
R4227 VDD.n3953 VDD.n3933 185
R4228 VDD.n4715 VDD.n4714 185
R4229 VDD.n4716 VDD.n4715 185
R4230 VDD.n3794 VDD.n3792 185
R4231 VDD.n3927 VDD.n3794 185
R4232 VDD.n5136 VDD.n5135 185
R4233 VDD.n5135 VDD.n5134 185
R4234 VDD.n3795 VDD.n3793 185
R4235 VDD.n3924 VDD.n3795 185
R4236 VDD.n5123 VDD.n5122 185
R4237 VDD.n5124 VDD.n5123 185
R4238 VDD.n3813 VDD.n3811 185
R4239 VDD.n3920 VDD.n3811 185
R4240 VDD.n5117 VDD.n5116 185
R4241 VDD.n5116 VDD.n5115 185
R4242 VDD.n3844 VDD.n3816 185
R4243 VDD.n4976 VDD.n3816 185
R4244 VDD.n3847 VDD.n3846 185
R4245 VDD.n3846 VDD.n3826 185
R4246 VDD.n3848 VDD.n3839 185
R4247 VDD.n3839 VDD.n3835 185
R4248 VDD.n5100 VDD.n5099 185
R4249 VDD.n5101 VDD.n5100 185
R4250 VDD.n3842 VDD.n3840 185
R4251 VDD.n4768 VDD.n3840 185
R4252 VDD.n5094 VDD.n5093 185
R4253 VDD.n5093 VDD.n5092 185
R4254 VDD.n4789 VDD.n3854 185
R4255 VDD.n3917 VDD.n3854 185
R4256 VDD.n4793 VDD.n4792 185
R4257 VDD.n4793 VDD.n3867 185
R4258 VDD.n4795 VDD.n4794 185
R4259 VDD.n4794 VDD.n3913 185
R4260 VDD.n4786 VDD.n4785 185
R4261 VDD.n4785 VDD.n3880 185
R4262 VDD.n4800 VDD.n4799 185
R4263 VDD.n4800 VDD.n3911 185
R4264 VDD.n4801 VDD.n4784 185
R4265 VDD.n4801 VDD.n3886 185
R4266 VDD.n4803 VDD.n4802 185
R4267 VDD.n4802 VDD.n3889 185
R4268 VDD.n4804 VDD.n4782 185
R4269 VDD.n4782 VDD.n3908 185
R4270 VDD.n4941 VDD.n4940 185
R4271 VDD.n4942 VDD.n4941 185
R4272 VDD.n4939 VDD.n4783 185
R4273 VDD.n4783 VDD.n4781 185
R4274 VDD.n4938 VDD.n4937 185
R4275 VDD.n4937 VDD.n4936 185
R4276 VDD.n4806 VDD.n4805 185
R4277 VDD.n4935 VDD.n4806 185
R4278 VDD.n4933 VDD.n4932 185
R4279 VDD.n4934 VDD.n4933 185
R4280 VDD.n4931 VDD.n4811 185
R4281 VDD.n4811 VDD.n4810 185
R4282 VDD.n4930 VDD.n4929 185
R4283 VDD.n4929 VDD.n4928 185
R4284 VDD.n4813 VDD.n4812 185
R4285 VDD.n4927 VDD.n4813 185
R4286 VDD.n4925 VDD.n4924 185
R4287 VDD.n4926 VDD.n4925 185
R4288 VDD.n4923 VDD.n4817 185
R4289 VDD.n4820 VDD.n4817 185
R4290 VDD.n4922 VDD.n4921 185
R4291 VDD.n4921 VDD.n4920 185
R4292 VDD.n4819 VDD.n4818 185
R4293 VDD.n4919 VDD.n4819 185
R4294 VDD.n4917 VDD.n4916 185
R4295 VDD.n4918 VDD.n4917 185
R4296 VDD.n4915 VDD.n4825 185
R4297 VDD.n4825 VDD.n4824 185
R4298 VDD.n4914 VDD.n4913 185
R4299 VDD.n4913 VDD.n4912 185
R4300 VDD.n4827 VDD.n4826 185
R4301 VDD.n4911 VDD.n4827 185
R4302 VDD.n4909 VDD.n4908 185
R4303 VDD.n4910 VDD.n4909 185
R4304 VDD.n4907 VDD.n4832 185
R4305 VDD.n4832 VDD.n4831 185
R4306 VDD.n4906 VDD.n4905 185
R4307 VDD.n4905 VDD.n4904 185
R4308 VDD.n4834 VDD.n4833 185
R4309 VDD.n4903 VDD.n4834 185
R4310 VDD.n4900 VDD.n4899 185
R4311 VDD.n4898 VDD.n4845 185
R4312 VDD.n4897 VDD.n4844 185
R4313 VDD.n4902 VDD.n4844 185
R4314 VDD.n4896 VDD.n4895 185
R4315 VDD.n4894 VDD.n4893 185
R4316 VDD.n4892 VDD.n4891 185
R4317 VDD.n4890 VDD.n4889 185
R4318 VDD.n4888 VDD.n4887 185
R4319 VDD.n4886 VDD.n4885 185
R4320 VDD.n4884 VDD.n4883 185
R4321 VDD.n4882 VDD.n4881 185
R4322 VDD.n4880 VDD.n4879 185
R4323 VDD.n4878 VDD.n4877 185
R4324 VDD.n4876 VDD.n4875 185
R4325 VDD.n4874 VDD.n4873 185
R4326 VDD.n4872 VDD.n4871 185
R4327 VDD.n4870 VDD.n4869 185
R4328 VDD.n4868 VDD.n4836 185
R4329 VDD.n4903 VDD.n4836 185
R4330 VDD.n4867 VDD.n4835 185
R4331 VDD.n4904 VDD.n4835 185
R4332 VDD.n4866 VDD.n4865 185
R4333 VDD.n4865 VDD.n4831 185
R4334 VDD.n4864 VDD.n4830 185
R4335 VDD.n4910 VDD.n4830 185
R4336 VDD.n4863 VDD.n4829 185
R4337 VDD.n4911 VDD.n4829 185
R4338 VDD.n4862 VDD.n4828 185
R4339 VDD.n4912 VDD.n4828 185
R4340 VDD.n4861 VDD.n4860 185
R4341 VDD.n4860 VDD.n4824 185
R4342 VDD.n4859 VDD.n4823 185
R4343 VDD.n4918 VDD.n4823 185
R4344 VDD.n4858 VDD.n4822 185
R4345 VDD.n4919 VDD.n4822 185
R4346 VDD.n4857 VDD.n4821 185
R4347 VDD.n4920 VDD.n4821 185
R4348 VDD.n4856 VDD.n4855 185
R4349 VDD.n4855 VDD.n4820 185
R4350 VDD.n4854 VDD.n4816 185
R4351 VDD.n4926 VDD.n4816 185
R4352 VDD.n4853 VDD.n4815 185
R4353 VDD.n4927 VDD.n4815 185
R4354 VDD.n4852 VDD.n4814 185
R4355 VDD.n4928 VDD.n4814 185
R4356 VDD.n4851 VDD.n4850 185
R4357 VDD.n4850 VDD.n4810 185
R4358 VDD.n4849 VDD.n4809 185
R4359 VDD.n4934 VDD.n4809 185
R4360 VDD.n4848 VDD.n4808 185
R4361 VDD.n4935 VDD.n4808 185
R4362 VDD.n4847 VDD.n4807 185
R4363 VDD.n4936 VDD.n4807 185
R4364 VDD.n4846 VDD.n4779 185
R4365 VDD.n4781 VDD.n4779 185
R4366 VDD.n4943 VDD.n4780 185
R4367 VDD.n4943 VDD.n4942 185
R4368 VDD.n4944 VDD.n4778 185
R4369 VDD.n4944 VDD.n3908 185
R4370 VDD.n4946 VDD.n4945 185
R4371 VDD.n4945 VDD.n3889 185
R4372 VDD.n4947 VDD.n4777 185
R4373 VDD.n4777 VDD.n3886 185
R4374 VDD.n4949 VDD.n4948 185
R4375 VDD.n4949 VDD.n3911 185
R4376 VDD.n4951 VDD.n4950 185
R4377 VDD.n4950 VDD.n3880 185
R4378 VDD.n4774 VDD.n4773 185
R4379 VDD.n4773 VDD.n3913 185
R4380 VDD.n4957 VDD.n4956 185
R4381 VDD.n4957 VDD.n3867 185
R4382 VDD.n4959 VDD.n4958 185
R4383 VDD.n4958 VDD.n3917 185
R4384 VDD.n4961 VDD.n3856 185
R4385 VDD.n5092 VDD.n3856 185
R4386 VDD.n4770 VDD.n4769 185
R4387 VDD.n4769 VDD.n4768 185
R4388 VDD.n4966 VDD.n3837 185
R4389 VDD.n5101 VDD.n3837 185
R4390 VDD.n4969 VDD.n4968 185
R4391 VDD.n4968 VDD.n3835 185
R4392 VDD.n4753 VDD.n4751 185
R4393 VDD.n4751 VDD.n3826 185
R4394 VDD.n4975 VDD.n4974 185
R4395 VDD.n4976 VDD.n4975 185
R4396 VDD.n4762 VDD.n3817 185
R4397 VDD.n5115 VDD.n3817 185
R4398 VDD.n4761 VDD.n3809 185
R4399 VDD.n3920 VDD.n3809 185
R4400 VDD.n5126 VDD.n5125 185
R4401 VDD.n5125 VDD.n5124 185
R4402 VDD.n3808 VDD.n3806 185
R4403 VDD.n3924 VDD.n3808 185
R4404 VDD.n3947 VDD.n3796 185
R4405 VDD.n5134 VDD.n3796 185
R4406 VDD.n3950 VDD.n3949 185
R4407 VDD.n3950 VDD.n3927 185
R4408 VDD.n4718 VDD.n4717 185
R4409 VDD.n4717 VDD.n4716 185
R4410 VDD.n3946 VDD.n3944 185
R4411 VDD.n3946 VDD.n3933 185
R4412 VDD.n3977 VDD.n3959 185
R4413 VDD.n4706 VDD.n3959 185
R4414 VDD.n4691 VDD.n4690 185
R4415 VDD.n4690 VDD.n4689 185
R4416 VDD.n4688 VDD.n3975 185
R4417 VDD.n4688 VDD.n3964 185
R4418 VDD.n4687 VDD.n3983 185
R4419 VDD.n4687 VDD.n4686 185
R4420 VDD.n4663 VDD.n3981 185
R4421 VDD.n4017 VDD.n3981 185
R4422 VDD.n4661 VDD.n3992 185
R4423 VDD.n4672 VDD.n3992 185
R4424 VDD.n4607 VDD.n4002 185
R4425 VDD.n4607 VDD.n4020 185
R4426 VDD.n4610 VDD.n4609 185
R4427 VDD.n4610 VDD.n4006 185
R4428 VDD.n4612 VDD.n4611 185
R4429 VDD.n4611 VDD.n4023 185
R4430 VDD.n4606 VDD.n4038 185
R4431 VDD.n4606 VDD.n4605 185
R4432 VDD.n4570 VDD.n4042 185
R4433 VDD.n4042 VDD.n4027 185
R4434 VDD.n4568 VDD.n4050 185
R4435 VDD.n4587 VDD.n4050 185
R4436 VDD.n4566 VDD.n4565 185
R4437 VDD.n4565 VDD.n4057 185
R4438 VDD.n3451 VDD.n3449 185
R4439 VDD.n4059 VDD.n3451 185
R4440 VDD.n5149 VDD.n5148 185
R4441 VDD.n5148 VDD.n5147 185
R4442 VDD.n3450 VDD.n3448 185
R4443 VDD.n3450 VDD.n3440 185
R4444 VDD.n4529 VDD.n4528 185
R4445 VDD.n4528 VDD.n4063 185
R4446 VDD.n4527 VDD.n4073 185
R4447 VDD.n4527 VDD.n4066 185
R4448 VDD.n4526 VDD.n4077 185
R4449 VDD.n4526 VDD.n4525 185
R4450 VDD.n4313 VDD.n4075 185
R4451 VDD.n4104 VDD.n4075 185
R4452 VDD.n4310 VDD.n4086 185
R4453 VDD.n4507 VDD.n4086 185
R4454 VDD.n4319 VDD.n4318 185
R4455 VDD.n4319 VDD.n4107 185
R4456 VDD.n4321 VDD.n4320 185
R4457 VDD.n4320 VDD.n4094 185
R4458 VDD.n4309 VDD.n4306 185
R4459 VDD.n4309 VDD.n4110 185
R4460 VDD.n4326 VDD.n4127 185
R4461 VDD.n4457 VDD.n4127 185
R4462 VDD.n4329 VDD.n4328 185
R4463 VDD.n4328 VDD.n4114 185
R4464 VDD.n4304 VDD.n4135 185
R4465 VDD.n4439 VDD.n4135 185
R4466 VDD.n4335 VDD.n4334 185
R4467 VDD.n4335 VDD.n4121 185
R4468 VDD.n4337 VDD.n4336 185
R4469 VDD.n4336 VDD.n4138 185
R4470 VDD.n4338 VDD.n4160 185
R4471 VDD.n4354 VDD.n4160 185
R4472 VDD.n4340 VDD.n4339 185
R4473 VDD.n4339 VDD.n4151 185
R4474 VDD.n4341 VDD.n4167 185
R4475 VDD.n4167 VDD.n4142 185
R4476 VDD.n4343 VDD.n4342 185
R4477 VDD.n4344 VDD.n4343 185
R4478 VDD.n4302 VDD.n4166 185
R4479 VDD.n4166 VDD.n4165 185
R4480 VDD.n4301 VDD.n4300 185
R4481 VDD.n4300 VDD.n4299 185
R4482 VDD.n4169 VDD.n4168 185
R4483 VDD.n4170 VDD.n4169 185
R4484 VDD.n4291 VDD.n4290 185
R4485 VDD.n4292 VDD.n4291 185
R4486 VDD.n4289 VDD.n4175 185
R4487 VDD.n4175 VDD.n4174 185
R4488 VDD.n4288 VDD.n4287 185
R4489 VDD.n4287 VDD.n4286 185
R4490 VDD.n4177 VDD.n4176 185
R4491 VDD.n4279 VDD.n4177 185
R4492 VDD.n4278 VDD.n4277 185
R4493 VDD.n4280 VDD.n4278 185
R4494 VDD.n4276 VDD.n4181 185
R4495 VDD.n4184 VDD.n4181 185
R4496 VDD.n4275 VDD.n4274 185
R4497 VDD.n4274 VDD.n4273 185
R4498 VDD.n4183 VDD.n4182 185
R4499 VDD.n4266 VDD.n4183 185
R4500 VDD.n4265 VDD.n4264 185
R4501 VDD.n4267 VDD.n4265 185
R4502 VDD.n4263 VDD.n4189 185
R4503 VDD.n4189 VDD.n4188 185
R4504 VDD.n4262 VDD.n4261 185
R4505 VDD.n4261 VDD.n4260 185
R4506 VDD.n4191 VDD.n4190 185
R4507 VDD.n4192 VDD.n4191 185
R4508 VDD.n4253 VDD.n4252 185
R4509 VDD.n4254 VDD.n4253 185
R4510 VDD.n4251 VDD.n4197 185
R4511 VDD.n4197 VDD.n4196 185
R4512 VDD.n4250 VDD.n4249 185
R4513 VDD.n4249 VDD.n4248 185
R4514 VDD.n4199 VDD.n4198 185
R4515 VDD.n4200 VDD.n4199 185
R4516 VDD.n419 VDD.n140 185
R4517 VDD.n418 VDD.n417 185
R4518 VDD.n415 VDD.n141 185
R4519 VDD.n413 VDD.n412 185
R4520 VDD.n411 VDD.n142 185
R4521 VDD.n410 VDD.n409 185
R4522 VDD.n407 VDD.n143 185
R4523 VDD.n405 VDD.n404 185
R4524 VDD.n145 VDD.n144 185
R4525 VDD.n399 VDD.n398 185
R4526 VDD.n396 VDD.n395 185
R4527 VDD.n394 VDD.n393 185
R4528 VDD.n392 VDD.n350 185
R4529 VDD.n390 VDD.n389 185
R4530 VDD.n388 VDD.n351 185
R4531 VDD.n387 VDD.n386 185
R4532 VDD.n384 VDD.n383 185
R4533 VDD.n384 VDD.n139 185
R4534 VDD.n382 VDD.n138 185
R4535 VDD.n422 VDD.n138 185
R4536 VDD.n381 VDD.n380 185
R4537 VDD.n380 VDD.n133 185
R4538 VDD.n379 VDD.n132 185
R4539 VDD.n428 VDD.n132 185
R4540 VDD.n378 VDD.n377 185
R4541 VDD.n377 VDD.n127 185
R4542 VDD.n376 VDD.n126 185
R4543 VDD.n434 VDD.n126 185
R4544 VDD.n375 VDD.n374 185
R4545 VDD.n374 VDD.n124 185
R4546 VDD.n373 VDD.n120 185
R4547 VDD.n440 VDD.n120 185
R4548 VDD.n372 VDD.n371 185
R4549 VDD.n371 VDD.n115 185
R4550 VDD.n370 VDD.n114 185
R4551 VDD.n446 VDD.n114 185
R4552 VDD.n369 VDD.n368 185
R4553 VDD.n368 VDD.n112 185
R4554 VDD.n367 VDD.n108 185
R4555 VDD.n452 VDD.n108 185
R4556 VDD.n366 VDD.n365 185
R4557 VDD.n365 VDD.n103 185
R4558 VDD.n364 VDD.n102 185
R4559 VDD.n458 VDD.n102 185
R4560 VDD.n363 VDD.n362 185
R4561 VDD.n362 VDD.n100 185
R4562 VDD.n361 VDD.n96 185
R4563 VDD.n464 VDD.n96 185
R4564 VDD.n360 VDD.n359 185
R4565 VDD.n359 VDD.n91 185
R4566 VDD.n358 VDD.n90 185
R4567 VDD.n470 VDD.n90 185
R4568 VDD.n357 VDD.n356 185
R4569 VDD.n356 VDD.n88 185
R4570 VDD.n355 VDD.n84 185
R4571 VDD.n476 VDD.n84 185
R4572 VDD.n354 VDD.n353 185
R4573 VDD.n353 VDD.n49 185
R4574 VDD.n352 VDD.n48 185
R4575 VDD.n482 VDD.n48 185
R4576 VDD.n37 VDD.n36 185
R4577 VDD.n40 VDD.n37 185
R4578 VDD.n490 VDD.n489 185
R4579 VDD.n489 VDD.n488 185
R4580 VDD.n491 VDD.n35 185
R4581 VDD.n38 VDD.n35 185
R4582 VDD.n493 VDD.n492 185
R4583 VDD.n495 VDD.n33 185
R4584 VDD.n497 VDD.n496 185
R4585 VDD.n498 VDD.n32 185
R4586 VDD.n500 VDD.n499 185
R4587 VDD.n502 VDD.n29 185
R4588 VDD.n504 VDD.n503 185
R4589 VDD.n60 VDD.n28 185
R4590 VDD.n62 VDD.n61 185
R4591 VDD.n64 VDD.n57 185
R4592 VDD.n66 VDD.n65 185
R4593 VDD.n68 VDD.n55 185
R4594 VDD.n70 VDD.n69 185
R4595 VDD.n71 VDD.n54 185
R4596 VDD.n73 VDD.n72 185
R4597 VDD.n75 VDD.n53 185
R4598 VDD.n76 VDD.n52 185
R4599 VDD.n76 VDD.n31 185
R4600 VDD.n78 VDD.n77 185
R4601 VDD.n77 VDD.n38 185
R4602 VDD.n79 VDD.n41 185
R4603 VDD.n488 VDD.n41 185
R4604 VDD.n80 VDD.n50 185
R4605 VDD.n50 VDD.n40 185
R4606 VDD.n481 VDD.n480 185
R4607 VDD.n482 VDD.n481 185
R4608 VDD.n479 VDD.n51 185
R4609 VDD.n51 VDD.n49 185
R4610 VDD.n478 VDD.n477 185
R4611 VDD.n477 VDD.n476 185
R4612 VDD.n82 VDD.n81 185
R4613 VDD.n88 VDD.n82 185
R4614 VDD.n469 VDD.n468 185
R4615 VDD.n470 VDD.n469 185
R4616 VDD.n467 VDD.n92 185
R4617 VDD.n92 VDD.n91 185
R4618 VDD.n466 VDD.n465 185
R4619 VDD.n465 VDD.n464 185
R4620 VDD.n94 VDD.n93 185
R4621 VDD.n100 VDD.n94 185
R4622 VDD.n457 VDD.n456 185
R4623 VDD.n458 VDD.n457 185
R4624 VDD.n455 VDD.n104 185
R4625 VDD.n104 VDD.n103 185
R4626 VDD.n454 VDD.n453 185
R4627 VDD.n453 VDD.n452 185
R4628 VDD.n106 VDD.n105 185
R4629 VDD.n112 VDD.n106 185
R4630 VDD.n445 VDD.n444 185
R4631 VDD.n446 VDD.n445 185
R4632 VDD.n443 VDD.n116 185
R4633 VDD.n116 VDD.n115 185
R4634 VDD.n442 VDD.n441 185
R4635 VDD.n441 VDD.n440 185
R4636 VDD.n118 VDD.n117 185
R4637 VDD.n124 VDD.n118 185
R4638 VDD.n433 VDD.n432 185
R4639 VDD.n434 VDD.n433 185
R4640 VDD.n431 VDD.n128 185
R4641 VDD.n128 VDD.n127 185
R4642 VDD.n430 VDD.n429 185
R4643 VDD.n429 VDD.n428 185
R4644 VDD.n130 VDD.n129 185
R4645 VDD.n133 VDD.n130 185
R4646 VDD.n421 VDD.n420 185
R4647 VDD.n422 VDD.n421 185
R4648 VDD.n220 VDD.n204 185
R4649 VDD.n220 VDD.n31 185
R4650 VDD.n219 VDD.n205 185
R4651 VDD.n217 VDD.n216 185
R4652 VDD.n215 VDD.n206 185
R4653 VDD.n214 VDD.n213 185
R4654 VDD.n211 VDD.n207 185
R4655 VDD.n209 VDD.n208 185
R4656 VDD.n44 VDD.n42 185
R4657 VDD.n42 VDD.n38 185
R4658 VDD.n487 VDD.n486 185
R4659 VDD.n488 VDD.n487 185
R4660 VDD.n485 VDD.n43 185
R4661 VDD.n43 VDD.n40 185
R4662 VDD.n484 VDD.n483 185
R4663 VDD.n483 VDD.n482 185
R4664 VDD.n46 VDD.n45 185
R4665 VDD.n49 VDD.n46 185
R4666 VDD.n475 VDD.n474 185
R4667 VDD.n476 VDD.n475 185
R4668 VDD.n473 VDD.n85 185
R4669 VDD.n88 VDD.n85 185
R4670 VDD.n472 VDD.n471 185
R4671 VDD.n471 VDD.n470 185
R4672 VDD.n87 VDD.n86 185
R4673 VDD.n91 VDD.n87 185
R4674 VDD.n463 VDD.n462 185
R4675 VDD.n464 VDD.n463 185
R4676 VDD.n461 VDD.n97 185
R4677 VDD.n100 VDD.n97 185
R4678 VDD.n460 VDD.n459 185
R4679 VDD.n459 VDD.n458 185
R4680 VDD.n99 VDD.n98 185
R4681 VDD.n103 VDD.n99 185
R4682 VDD.n451 VDD.n450 185
R4683 VDD.n452 VDD.n451 185
R4684 VDD.n449 VDD.n109 185
R4685 VDD.n112 VDD.n109 185
R4686 VDD.n448 VDD.n447 185
R4687 VDD.n447 VDD.n446 185
R4688 VDD.n111 VDD.n110 185
R4689 VDD.n115 VDD.n111 185
R4690 VDD.n439 VDD.n438 185
R4691 VDD.n440 VDD.n439 185
R4692 VDD.n437 VDD.n121 185
R4693 VDD.n124 VDD.n121 185
R4694 VDD.n436 VDD.n435 185
R4695 VDD.n435 VDD.n434 185
R4696 VDD.n123 VDD.n122 185
R4697 VDD.n127 VDD.n123 185
R4698 VDD.n427 VDD.n426 185
R4699 VDD.n428 VDD.n427 185
R4700 VDD.n425 VDD.n134 185
R4701 VDD.n134 VDD.n133 185
R4702 VDD.n424 VDD.n423 185
R4703 VDD.n423 VDD.n422 185
R4704 VDD.n136 VDD.n135 185
R4705 VDD.n167 VDD.n166 185
R4706 VDD.n168 VDD.n164 185
R4707 VDD.n164 VDD.n139 185
R4708 VDD.n170 VDD.n169 185
R4709 VDD.n172 VDD.n163 185
R4710 VDD.n175 VDD.n174 185
R4711 VDD.n176 VDD.n162 185
R4712 VDD.n178 VDD.n177 185
R4713 VDD.n180 VDD.n155 185
R4714 VDD.n307 VDD.n306 185
R4715 VDD.n304 VDD.n303 185
R4716 VDD.n302 VDD.n181 185
R4717 VDD.n301 VDD.n300 185
R4718 VDD.n298 VDD.n182 185
R4719 VDD.n296 VDD.n295 185
R4720 VDD.n294 VDD.n183 185
R4721 VDD.n293 VDD.n292 185
R4722 VDD.n290 VDD.n137 185
R4723 VDD.n422 VDD.n137 185
R4724 VDD.n289 VDD.n288 185
R4725 VDD.n288 VDD.n133 185
R4726 VDD.n287 VDD.n131 185
R4727 VDD.n428 VDD.n131 185
R4728 VDD.n286 VDD.n285 185
R4729 VDD.n285 VDD.n127 185
R4730 VDD.n284 VDD.n125 185
R4731 VDD.n434 VDD.n125 185
R4732 VDD.n283 VDD.n282 185
R4733 VDD.n282 VDD.n124 185
R4734 VDD.n281 VDD.n119 185
R4735 VDD.n440 VDD.n119 185
R4736 VDD.n280 VDD.n279 185
R4737 VDD.n279 VDD.n115 185
R4738 VDD.n278 VDD.n113 185
R4739 VDD.n446 VDD.n113 185
R4740 VDD.n277 VDD.n276 185
R4741 VDD.n276 VDD.n112 185
R4742 VDD.n275 VDD.n107 185
R4743 VDD.n452 VDD.n107 185
R4744 VDD.n274 VDD.n273 185
R4745 VDD.n273 VDD.n103 185
R4746 VDD.n272 VDD.n101 185
R4747 VDD.n458 VDD.n101 185
R4748 VDD.n271 VDD.n270 185
R4749 VDD.n270 VDD.n100 185
R4750 VDD.n269 VDD.n95 185
R4751 VDD.n464 VDD.n95 185
R4752 VDD.n268 VDD.n267 185
R4753 VDD.n267 VDD.n91 185
R4754 VDD.n266 VDD.n89 185
R4755 VDD.n470 VDD.n89 185
R4756 VDD.n265 VDD.n264 185
R4757 VDD.n264 VDD.n88 185
R4758 VDD.n263 VDD.n83 185
R4759 VDD.n476 VDD.n83 185
R4760 VDD.n262 VDD.n261 185
R4761 VDD.n261 VDD.n49 185
R4762 VDD.n260 VDD.n47 185
R4763 VDD.n482 VDD.n47 185
R4764 VDD.n259 VDD.n258 185
R4765 VDD.n258 VDD.n40 185
R4766 VDD.n257 VDD.n39 185
R4767 VDD.n488 VDD.n39 185
R4768 VDD.n256 VDD.n255 185
R4769 VDD.n255 VDD.n38 185
R4770 VDD.n254 VDD.n184 185
R4771 VDD.n252 VDD.n251 185
R4772 VDD.n250 VDD.n185 185
R4773 VDD.n249 VDD.n248 185
R4774 VDD.n246 VDD.n186 185
R4775 VDD.n244 VDD.n243 185
R4776 VDD.n242 VDD.n187 185
R4777 VDD.n225 VDD.n188 185
R4778 VDD.n228 VDD.n227 185
R4779 VDD.n229 VDD.n221 185
R4780 VDD.n2476 VDD.n1296 185
R4781 VDD.n2475 VDD.n2474 185
R4782 VDD.n1298 VDD.n1297 185
R4783 VDD.n2407 VDD.n2406 185
R4784 VDD.n2409 VDD.n2408 185
R4785 VDD.n2411 VDD.n2410 185
R4786 VDD.n2413 VDD.n2412 185
R4787 VDD.n2415 VDD.n2414 185
R4788 VDD.n2417 VDD.n2416 185
R4789 VDD.n2419 VDD.n2418 185
R4790 VDD.n2421 VDD.n2420 185
R4791 VDD.n2423 VDD.n2422 185
R4792 VDD.n2425 VDD.n2424 185
R4793 VDD.n2427 VDD.n2426 185
R4794 VDD.n2429 VDD.n2428 185
R4795 VDD.n2431 VDD.n2430 185
R4796 VDD.n2432 VDD.n1313 185
R4797 VDD.n2472 VDD.n1313 185
R4798 VDD.n2433 VDD.n1294 185
R4799 VDD.n2479 VDD.n1294 185
R4800 VDD.n2435 VDD.n2434 185
R4801 VDD.n2436 VDD.n2435 185
R4802 VDD.n2405 VDD.n1288 185
R4803 VDD.n2485 VDD.n1288 185
R4804 VDD.n2404 VDD.n2403 185
R4805 VDD.n2403 VDD.n2402 185
R4806 VDD.n1318 VDD.n1275 185
R4807 VDD.n2491 VDD.n1275 185
R4808 VDD.n2395 VDD.n2394 185
R4809 VDD.n2396 VDD.n2395 185
R4810 VDD.n2393 VDD.n1264 185
R4811 VDD.n2497 VDD.n1264 185
R4812 VDD.n2392 VDD.n2391 185
R4813 VDD.n2391 VDD.n1261 185
R4814 VDD.n2390 VDD.n2389 185
R4815 VDD.n2390 VDD.n1244 185
R4816 VDD.n2388 VDD.n1242 185
R4817 VDD.n2508 VDD.n1242 185
R4818 VDD.n2387 VDD.n1234 185
R4819 VDD.n2514 VDD.n1234 185
R4820 VDD.n2386 VDD.n2385 185
R4821 VDD.n2385 VDD.n2384 185
R4822 VDD.n2156 VDD.n1225 185
R4823 VDD.n2520 VDD.n1225 185
R4824 VDD.n2155 VDD.n2154 185
R4825 VDD.n2154 VDD.n2153 185
R4826 VDD.n1325 VDD.n1324 185
R4827 VDD.n1325 VDD.n1216 185
R4828 VDD.n2144 VDD.n2143 185
R4829 VDD.n2145 VDD.n2144 185
R4830 VDD.n2142 VDD.n1204 185
R4831 VDD.n2539 VDD.n1204 185
R4832 VDD.n2141 VDD.n2140 185
R4833 VDD.n2140 VDD.n2139 185
R4834 VDD.n1332 VDD.n1331 185
R4835 VDD.n1358 VDD.n1332 185
R4836 VDD.n2108 VDD.n1341 185
R4837 VDD.n2131 VDD.n1341 185
R4838 VDD.n2110 VDD.n2109 185
R4839 VDD.n2111 VDD.n2110 185
R4840 VDD.n2107 VDD.n1367 185
R4841 VDD.n1367 VDD.n1364 185
R4842 VDD.n2106 VDD.n2105 185
R4843 VDD.n2105 VDD.n2104 185
R4844 VDD.n1369 VDD.n1368 185
R4845 VDD.n1390 VDD.n1369 185
R4846 VDD.n2050 VDD.n2049 185
R4847 VDD.n2051 VDD.n2050 185
R4848 VDD.n2048 VDD.n1400 185
R4849 VDD.n2077 VDD.n1400 185
R4850 VDD.n2047 VDD.n2046 185
R4851 VDD.n2046 VDD.n2045 185
R4852 VDD.n1425 VDD.n1414 185
R4853 VDD.n2058 VDD.n1414 185
R4854 VDD.n2030 VDD.n2029 185
R4855 VDD.t10 VDD.n2030 185
R4856 VDD.n2028 VDD.n1430 185
R4857 VDD.n1449 VDD.n1430 185
R4858 VDD.n2027 VDD.n2026 185
R4859 VDD.n2026 VDD.n2025 185
R4860 VDD.n1432 VDD.n1431 185
R4861 VDD.n1992 VDD.n1432 185
R4862 VDD.n1950 VDD.n1464 185
R4863 VDD.n1983 VDD.n1464 185
R4864 VDD.n1952 VDD.n1951 185
R4865 VDD.n1955 VDD.n1952 185
R4866 VDD.n1949 VDD.n1466 185
R4867 VDD.n1466 VDD.n858 185
R4868 VDD.n1948 VDD.n847 185
R4869 VDD.n2562 VDD.n847 185
R4870 VDD.n1947 VDD.n1946 185
R4871 VDD.n1946 VDD.n1945 185
R4872 VDD.n1468 VDD.n1467 185
R4873 VDD.n1942 VDD.n1468 185
R4874 VDD.n1894 VDD.n1511 185
R4875 VDD.n1511 VDD.n1484 185
R4876 VDD.n1896 VDD.n1895 185
R4877 VDD.n1897 VDD.n1896 185
R4878 VDD.n1893 VDD.n1494 185
R4879 VDD.n1912 VDD.n1494 185
R4880 VDD.n1892 VDD.n1891 185
R4881 VDD.n1891 VDD.n1890 185
R4882 VDD.n1512 VDD.n1502 185
R4883 VDD.n1905 VDD.n1502 185
R4884 VDD.n1883 VDD.n1882 185
R4885 VDD.n1884 VDD.n1883 185
R4886 VDD.n1881 VDD.n1517 185
R4887 VDD.n1864 VDD.n1517 185
R4888 VDD.n1880 VDD.n1879 185
R4889 VDD.n1879 VDD.n1878 185
R4890 VDD.n1519 VDD.n1518 185
R4891 VDD.n1844 VDD.n1519 185
R4892 VDD.n1834 VDD.n1529 185
R4893 VDD.n1871 VDD.n1529 185
R4894 VDD.n1836 VDD.n1835 185
R4895 VDD.n1837 VDD.n1836 185
R4896 VDD.n1833 VDD.n1545 185
R4897 VDD.n1792 VDD.n1545 185
R4898 VDD.n1832 VDD.n1831 185
R4899 VDD.n1547 VDD.n1546 185
R4900 VDD.n1762 VDD.n1761 185
R4901 VDD.n1764 VDD.n1763 185
R4902 VDD.n1766 VDD.n1765 185
R4903 VDD.n1768 VDD.n1767 185
R4904 VDD.n1770 VDD.n1769 185
R4905 VDD.n1772 VDD.n1771 185
R4906 VDD.n1774 VDD.n1773 185
R4907 VDD.n1776 VDD.n1775 185
R4908 VDD.n1778 VDD.n1777 185
R4909 VDD.n1780 VDD.n1779 185
R4910 VDD.n1782 VDD.n1781 185
R4911 VDD.n1784 VDD.n1783 185
R4912 VDD.n1786 VDD.n1785 185
R4913 VDD.n1788 VDD.n1787 185
R4914 VDD.n1789 VDD.n1549 185
R4915 VDD.n1829 VDD.n1549 185
R4916 VDD.n1791 VDD.n1790 185
R4917 VDD.n1792 VDD.n1791 185
R4918 VDD.n1532 VDD.n1530 185
R4919 VDD.n1837 VDD.n1530 185
R4920 VDD.n1870 VDD.n1869 185
R4921 VDD.n1871 VDD.n1870 185
R4922 VDD.n1868 VDD.n1531 185
R4923 VDD.n1844 VDD.n1531 185
R4924 VDD.n1867 VDD.n1522 185
R4925 VDD.n1878 VDD.n1522 185
R4926 VDD.n1866 VDD.n1865 185
R4927 VDD.n1865 VDD.n1864 185
R4928 VDD.n1505 VDD.n1503 185
R4929 VDD.n1884 VDD.n1503 185
R4930 VDD.n1904 VDD.n1903 185
R4931 VDD.n1905 VDD.n1904 185
R4932 VDD.n1902 VDD.n1504 185
R4933 VDD.n1890 VDD.n1504 185
R4934 VDD.n1901 VDD.n1495 185
R4935 VDD.n1912 VDD.n1495 185
R4936 VDD.n1899 VDD.n1507 185
R4937 VDD.n1897 VDD.n1507 185
R4938 VDD.n1508 VDD.n1470 185
R4939 VDD.n1484 VDD.n1470 185
R4940 VDD.n1943 VDD.n1471 185
R4941 VDD.n1943 VDD.n1942 185
R4942 VDD.n1944 VDD.n841 185
R4943 VDD.n1945 VDD.n1944 185
R4944 VDD.n2564 VDD.n842 185
R4945 VDD.n2562 VDD.n842 185
R4946 VDD.n1953 VDD.n843 185
R4947 VDD.n1953 VDD.n858 185
R4948 VDD.n1954 VDD.n1461 185
R4949 VDD.n1955 VDD.n1954 185
R4950 VDD.n1985 VDD.n1458 185
R4951 VDD.n1983 VDD.n1458 185
R4952 VDD.n1991 VDD.n1990 185
R4953 VDD.n1992 VDD.n1991 185
R4954 VDD.n1989 VDD.n1435 185
R4955 VDD.n2025 VDD.n1435 185
R4956 VDD.n1988 VDD.n1987 185
R4957 VDD.n1987 VDD.n1449 185
R4958 VDD.n1417 VDD.n1415 185
R4959 VDD.t10 VDD.n1415 185
R4960 VDD.n2057 VDD.n2056 185
R4961 VDD.n2058 VDD.n2057 185
R4962 VDD.n2055 VDD.n1416 185
R4963 VDD.n2045 VDD.n1416 185
R4964 VDD.n2054 VDD.n1401 185
R4965 VDD.n2077 VDD.n1401 185
R4966 VDD.n2053 VDD.n2052 185
R4967 VDD.n2052 VDD.n2051 185
R4968 VDD.n1422 VDD.n1421 185
R4969 VDD.n1422 VDD.n1390 185
R4970 VDD.n1420 VDD.n1372 185
R4971 VDD.n2104 VDD.n1372 185
R4972 VDD.n1419 VDD.n1418 185
R4973 VDD.n1418 VDD.n1364 185
R4974 VDD.n1338 VDD.n1337 185
R4975 VDD.n2111 VDD.n1338 185
R4976 VDD.n2133 VDD.n2132 185
R4977 VDD.n2132 VDD.n2131 185
R4978 VDD.n2134 VDD.n1335 185
R4979 VDD.n1358 VDD.n1335 185
R4980 VDD.n2138 VDD.n2137 185
R4981 VDD.n2139 VDD.n2138 185
R4982 VDD.n2136 VDD.n1205 185
R4983 VDD.n2539 VDD.n1205 185
R4984 VDD.n1329 VDD.n1328 185
R4985 VDD.n2145 VDD.n1328 185
R4986 VDD.n2149 VDD.n2148 185
R4987 VDD.n2149 VDD.n1216 185
R4988 VDD.n2152 VDD.n2151 185
R4989 VDD.n2153 VDD.n2152 185
R4990 VDD.n2150 VDD.n1226 185
R4991 VDD.n2520 VDD.n1226 185
R4992 VDD.n1237 VDD.n1235 185
R4993 VDD.n2384 VDD.n1235 185
R4994 VDD.n2513 VDD.n2512 185
R4995 VDD.n2514 VDD.n2513 185
R4996 VDD.n1238 VDD.n1236 185
R4997 VDD.n2508 VDD.n1236 185
R4998 VDD.n1279 VDD.n1278 185
R4999 VDD.n1279 VDD.n1244 185
R5000 VDD.n1281 VDD.n1280 185
R5001 VDD.n1280 VDD.n1261 185
R5002 VDD.n1282 VDD.n1265 185
R5003 VDD.n2497 VDD.n1265 185
R5004 VDD.n1283 VDD.n1276 185
R5005 VDD.n2396 VDD.n1276 185
R5006 VDD.n2490 VDD.n2489 185
R5007 VDD.n2491 VDD.n2490 185
R5008 VDD.n2488 VDD.n1277 185
R5009 VDD.n2402 VDD.n1277 185
R5010 VDD.n2487 VDD.n2486 185
R5011 VDD.n2486 VDD.n2485 185
R5012 VDD.n1285 VDD.n1284 185
R5013 VDD.n2436 VDD.n1285 185
R5014 VDD.n2478 VDD.n2477 185
R5015 VDD.n2479 VDD.n2478 185
R5016 VDD.n1291 VDD.n1290 185
R5017 VDD.n2470 VDD.n2469 185
R5018 VDD.n2468 VDD.n1315 185
R5019 VDD.n2472 VDD.n1315 185
R5020 VDD.n2467 VDD.n2466 185
R5021 VDD.n2465 VDD.n2464 185
R5022 VDD.n2463 VDD.n2462 185
R5023 VDD.n2461 VDD.n2460 185
R5024 VDD.n2459 VDD.n2458 185
R5025 VDD.n2457 VDD.n2456 185
R5026 VDD.n2455 VDD.n2454 185
R5027 VDD.n2453 VDD.n2452 185
R5028 VDD.n2451 VDD.n2450 185
R5029 VDD.n2449 VDD.n2448 185
R5030 VDD.n2447 VDD.n2446 185
R5031 VDD.n2445 VDD.n2444 185
R5032 VDD.n2443 VDD.n2442 185
R5033 VDD.n2441 VDD.n2440 185
R5034 VDD.n2439 VDD.n1293 185
R5035 VDD.n2479 VDD.n1293 185
R5036 VDD.n2438 VDD.n2437 185
R5037 VDD.n2437 VDD.n2436 185
R5038 VDD.n1316 VDD.n1287 185
R5039 VDD.n2485 VDD.n1287 185
R5040 VDD.n2401 VDD.n2400 185
R5041 VDD.n2402 VDD.n2401 185
R5042 VDD.n2399 VDD.n1274 185
R5043 VDD.n2491 VDD.n1274 185
R5044 VDD.n2398 VDD.n2397 185
R5045 VDD.n2397 VDD.n2396 185
R5046 VDD.n1322 VDD.n1263 185
R5047 VDD.n2497 VDD.n1263 185
R5048 VDD.n1321 VDD.n1320 185
R5049 VDD.n1320 VDD.n1261 185
R5050 VDD.n1240 VDD.n1239 185
R5051 VDD.n1244 VDD.n1240 185
R5052 VDD.n2510 VDD.n2509 185
R5053 VDD.n2509 VDD.n2508 185
R5054 VDD.n2512 VDD.n1233 185
R5055 VDD.n2514 VDD.n1233 185
R5056 VDD.n2383 VDD.n1237 185
R5057 VDD.n2384 VDD.n2383 185
R5058 VDD.n2150 VDD.n1224 185
R5059 VDD.n2520 VDD.n1224 185
R5060 VDD.n2151 VDD.n1327 185
R5061 VDD.n2153 VDD.n1327 185
R5062 VDD.n2148 VDD.n2147 185
R5063 VDD.n2147 VDD.n1216 185
R5064 VDD.n2146 VDD.n1329 185
R5065 VDD.n2146 VDD.n2145 185
R5066 VDD.n2136 VDD.n1203 185
R5067 VDD.n2539 VDD.n1203 185
R5068 VDD.n2137 VDD.n1334 185
R5069 VDD.n2139 VDD.n1334 185
R5070 VDD.n1357 VDD.n1336 185
R5071 VDD.n1358 VDD.n1357 185
R5072 VDD.n2034 VDD.n1340 185
R5073 VDD.n2131 VDD.n1340 185
R5074 VDD.n2035 VDD.n1366 185
R5075 VDD.n2111 VDD.n1366 185
R5076 VDD.n2037 VDD.n2036 185
R5077 VDD.n2036 VDD.n1364 185
R5078 VDD.n2038 VDD.n1371 185
R5079 VDD.n2104 VDD.n1371 185
R5080 VDD.n2040 VDD.n2039 185
R5081 VDD.n2039 VDD.n1390 185
R5082 VDD.n2041 VDD.n1424 185
R5083 VDD.n2051 VDD.n1424 185
R5084 VDD.n2042 VDD.n1399 185
R5085 VDD.n2077 VDD.n1399 185
R5086 VDD.n2044 VDD.n2043 185
R5087 VDD.n2045 VDD.n2044 185
R5088 VDD.n2033 VDD.n1413 185
R5089 VDD.n2058 VDD.n1413 185
R5090 VDD.n2032 VDD.n2031 185
R5091 VDD.n2031 VDD.t10 185
R5092 VDD.n1428 VDD.n1427 185
R5093 VDD.n1449 VDD.n1428 185
R5094 VDD.n1459 VDD.n1434 185
R5095 VDD.n2025 VDD.n1434 185
R5096 VDD.n1460 VDD.n1457 185
R5097 VDD.n1992 VDD.n1457 185
R5098 VDD.n1985 VDD.n1984 185
R5099 VDD.n1984 VDD.n1983 185
R5100 VDD.n1462 VDD.n1461 185
R5101 VDD.n1955 VDD.n1462 185
R5102 VDD.n845 VDD.n843 185
R5103 VDD.n858 VDD.n845 185
R5104 VDD.n2564 VDD.n2563 185
R5105 VDD.n2563 VDD.n2562 185
R5106 VDD.n844 VDD.n841 185
R5107 VDD.n1945 VDD.n844 185
R5108 VDD.n1473 VDD.n1471 185
R5109 VDD.n1942 VDD.n1473 185
R5110 VDD.n1509 VDD.n1508 185
R5111 VDD.n1509 VDD.n1484 185
R5112 VDD.n1899 VDD.n1898 185
R5113 VDD.n1898 VDD.n1897 185
R5114 VDD.n1506 VDD.n1493 185
R5115 VDD.n1912 VDD.n1493 185
R5116 VDD.n1889 VDD.n1888 185
R5117 VDD.n1890 VDD.n1889 185
R5118 VDD.n1887 VDD.n1501 185
R5119 VDD.n1905 VDD.n1501 185
R5120 VDD.n1886 VDD.n1885 185
R5121 VDD.n1885 VDD.n1884 185
R5122 VDD.n1515 VDD.n1514 185
R5123 VDD.n1864 VDD.n1515 185
R5124 VDD.n1841 VDD.n1521 185
R5125 VDD.n1878 VDD.n1521 185
R5126 VDD.n1843 VDD.n1842 185
R5127 VDD.n1844 VDD.n1843 185
R5128 VDD.n1840 VDD.n1528 185
R5129 VDD.n1871 VDD.n1528 185
R5130 VDD.n1839 VDD.n1838 185
R5131 VDD.n1838 VDD.n1837 185
R5132 VDD.n1543 VDD.n1542 185
R5133 VDD.n1792 VDD.n1543 185
R5134 VDD.n1797 VDD.n1796 185
R5135 VDD.n1799 VDD.n1798 185
R5136 VDD.n1801 VDD.n1800 185
R5137 VDD.n1803 VDD.n1802 185
R5138 VDD.n1805 VDD.n1804 185
R5139 VDD.n1807 VDD.n1806 185
R5140 VDD.n1809 VDD.n1808 185
R5141 VDD.n1811 VDD.n1810 185
R5142 VDD.n1813 VDD.n1812 185
R5143 VDD.n1815 VDD.n1814 185
R5144 VDD.n1817 VDD.n1816 185
R5145 VDD.n1819 VDD.n1818 185
R5146 VDD.n1821 VDD.n1820 185
R5147 VDD.n1823 VDD.n1822 185
R5148 VDD.n1825 VDD.n1824 185
R5149 VDD.n1826 VDD.n1794 185
R5150 VDD.n1828 VDD.n1827 185
R5151 VDD.n1829 VDD.n1828 185
R5152 VDD.n1795 VDD.n1793 185
R5153 VDD.n1793 VDD.n1792 185
R5154 VDD.n1526 VDD.n1525 185
R5155 VDD.n1837 VDD.n1526 185
R5156 VDD.n1873 VDD.n1872 185
R5157 VDD.n1872 VDD.n1871 185
R5158 VDD.n1874 VDD.n1523 185
R5159 VDD.n1844 VDD.n1523 185
R5160 VDD.n1877 VDD.n1876 185
R5161 VDD.n1878 VDD.n1877 185
R5162 VDD.n1875 VDD.n1524 185
R5163 VDD.n1864 VDD.n1524 185
R5164 VDD.n1499 VDD.n1498 185
R5165 VDD.n1884 VDD.n1499 185
R5166 VDD.n1907 VDD.n1906 185
R5167 VDD.n1906 VDD.n1905 185
R5168 VDD.n1908 VDD.n1496 185
R5169 VDD.n1890 VDD.n1496 185
R5170 VDD.n1911 VDD.n1910 185
R5171 VDD.n1912 VDD.n1911 185
R5172 VDD.n1909 VDD.n1497 185
R5173 VDD.n1897 VDD.n1497 185
R5174 VDD.n1475 VDD.n1474 185
R5175 VDD.n1484 VDD.n1474 185
R5176 VDD.n1941 VDD.n1940 185
R5177 VDD.n1942 VDD.n1941 185
R5178 VDD.n1476 VDD.n848 185
R5179 VDD.n1945 VDD.n848 185
R5180 VDD.n2561 VDD.n2560 185
R5181 VDD.n2562 VDD.n2561 185
R5182 VDD.n851 VDD.n849 185
R5183 VDD.n858 VDD.n849 185
R5184 VDD.n1958 VDD.n1956 185
R5185 VDD.n1956 VDD.n1955 185
R5186 VDD.n1982 VDD.n1981 185
R5187 VDD.n1983 VDD.n1982 185
R5188 VDD.n1960 VDD.n1436 185
R5189 VDD.n1992 VDD.n1436 185
R5190 VDD.n2024 VDD.n2023 185
R5191 VDD.n2025 VDD.n2024 185
R5192 VDD.n1439 VDD.n1437 185
R5193 VDD.n1449 VDD.n1437 185
R5194 VDD.n1441 VDD.n1411 185
R5195 VDD.t10 VDD.n1411 185
R5196 VDD.n2060 VDD.n2059 185
R5197 VDD.n2059 VDD.n2058 185
R5198 VDD.n2061 VDD.n1402 185
R5199 VDD.n2045 VDD.n1402 185
R5200 VDD.n2076 VDD.n2075 185
R5201 VDD.n2077 VDD.n2076 185
R5202 VDD.n2074 VDD.n1403 185
R5203 VDD.n2051 VDD.n1403 185
R5204 VDD.n1405 VDD.n1373 185
R5205 VDD.n1390 VDD.n1373 185
R5206 VDD.n2103 VDD.n2102 185
R5207 VDD.n2104 VDD.n2103 185
R5208 VDD.n1376 VDD.n1374 185
R5209 VDD.n1374 VDD.n1364 185
R5210 VDD.n1378 VDD.n1342 185
R5211 VDD.n2111 VDD.n1342 185
R5212 VDD.n2130 VDD.n2129 185
R5213 VDD.n2131 VDD.n2130 185
R5214 VDD.n1345 VDD.n1343 185
R5215 VDD.n1358 VDD.n1343 185
R5216 VDD.n1347 VDD.n1206 185
R5217 VDD.n2139 VDD.n1206 185
R5218 VDD.n2538 VDD.n2537 185
R5219 VDD.n2539 VDD.n2538 185
R5220 VDD.n1209 VDD.n1207 185
R5221 VDD.n2145 VDD.n1207 185
R5222 VDD.n2163 VDD.n2162 185
R5223 VDD.n2162 VDD.n1216 185
R5224 VDD.n2164 VDD.n1227 185
R5225 VDD.n2153 VDD.n1227 185
R5226 VDD.n2519 VDD.n2518 185
R5227 VDD.n2520 VDD.n2519 185
R5228 VDD.n2517 VDD.n1228 185
R5229 VDD.n2384 VDD.n1228 185
R5230 VDD.n2516 VDD.n2515 185
R5231 VDD.n2515 VDD.n2514 185
R5232 VDD.n1231 VDD.n1230 185
R5233 VDD.n2508 VDD.n1231 185
R5234 VDD.n1269 VDD.n1268 185
R5235 VDD.n1268 VDD.n1244 185
R5236 VDD.n1270 VDD.n1266 185
R5237 VDD.n1266 VDD.n1261 185
R5238 VDD.n2496 VDD.n2495 185
R5239 VDD.n2497 VDD.n2496 185
R5240 VDD.n2494 VDD.n1267 185
R5241 VDD.n2396 VDD.n1267 185
R5242 VDD.n2493 VDD.n2492 185
R5243 VDD.n2492 VDD.n2491 185
R5244 VDD.n1272 VDD.n1271 185
R5245 VDD.n2402 VDD.n1272 185
R5246 VDD.n2484 VDD.n2483 185
R5247 VDD.n2485 VDD.n2484 185
R5248 VDD.n2482 VDD.n1289 185
R5249 VDD.n2436 VDD.n1289 185
R5250 VDD.n2481 VDD.n2480 185
R5251 VDD.n2480 VDD.n2479 185
R5252 VDD.n1646 VDD.n1645 185
R5253 VDD.n1647 VDD.n1646 185
R5254 VDD.n1644 VDD.n1617 185
R5255 VDD.n1643 VDD.n1642 185
R5256 VDD.n1641 VDD.n1640 185
R5257 VDD.n1639 VDD.n1638 185
R5258 VDD.n1637 VDD.n1636 185
R5259 VDD.n1635 VDD.n1634 185
R5260 VDD.n1633 VDD.n1632 185
R5261 VDD.n1631 VDD.n1630 185
R5262 VDD.n1629 VDD.n1628 185
R5263 VDD.n1627 VDD.n1626 185
R5264 VDD.n1625 VDD.n1624 185
R5265 VDD.n1623 VDD.n1622 185
R5266 VDD.n1621 VDD.n1620 185
R5267 VDD.n1619 VDD.n1618 185
R5268 VDD.n1609 VDD.n1608 185
R5269 VDD.n1650 VDD.n1649 185
R5270 VDD.n1651 VDD.n1607 185
R5271 VDD.n1607 VDD.n1606 185
R5272 VDD.n1653 VDD.n1652 185
R5273 VDD.n1654 VDD.n1653 185
R5274 VDD.n1601 VDD.n1600 185
R5275 VDD.n1602 VDD.n1601 185
R5276 VDD.n1662 VDD.n1661 185
R5277 VDD.n1661 VDD.n1660 185
R5278 VDD.n1663 VDD.n1599 185
R5279 VDD.n1599 VDD.n1598 185
R5280 VDD.n1665 VDD.n1664 185
R5281 VDD.n1666 VDD.n1665 185
R5282 VDD.n1593 VDD.n1592 185
R5283 VDD.n1594 VDD.n1593 185
R5284 VDD.n1675 VDD.n1674 185
R5285 VDD.n1674 VDD.n1673 185
R5286 VDD.n1676 VDD.n1591 185
R5287 VDD.n1672 VDD.n1591 185
R5288 VDD.n1678 VDD.n1677 185
R5289 VDD.n1679 VDD.n1678 185
R5290 VDD.n1586 VDD.n1585 185
R5291 VDD.n1590 VDD.n1586 185
R5292 VDD.n1688 VDD.n1687 185
R5293 VDD.n1687 VDD.n1686 185
R5294 VDD.n1689 VDD.n1584 185
R5295 VDD.n1685 VDD.n1584 185
R5296 VDD.n1691 VDD.n1690 185
R5297 VDD.n1692 VDD.n1691 185
R5298 VDD.n1579 VDD.n1578 185
R5299 VDD.n1580 VDD.n1579 185
R5300 VDD.n1700 VDD.n1699 185
R5301 VDD.n1699 VDD.n1698 185
R5302 VDD.n1701 VDD.n1577 185
R5303 VDD.n1577 VDD.n1576 185
R5304 VDD.n1704 VDD.n1703 185
R5305 VDD.n1705 VDD.n1704 185
R5306 VDD.n1702 VDD.n1570 185
R5307 VDD.n1571 VDD.n1570 185
R5308 VDD.n1751 VDD.n1569 185
R5309 VDD.n1751 VDD.n1750 185
R5310 VDD.n1753 VDD.n1752 185
R5311 VDD.n1752 VDD.n1548 185
R5312 VDD.n1754 VDD.n1567 185
R5313 VDD.n1567 VDD.n1557 185
R5314 VDD.n1759 VDD.n1758 185
R5315 VDD.n1760 VDD.n1759 185
R5316 VDD.n1757 VDD.n1568 185
R5317 VDD.n1568 VDD.n1544 185
R5318 VDD.n1755 VDD.n1540 185
R5319 VDD.n1540 VDD.n1527 185
R5320 VDD.n1847 VDD.n1846 185
R5321 VDD.n1846 VDD.n1845 185
R5322 VDD.n1848 VDD.n1534 185
R5323 VDD.n1534 VDD.n1520 185
R5324 VDD.n1862 VDD.n1861 185
R5325 VDD.n1863 VDD.n1862 185
R5326 VDD.n1537 VDD.n1535 185
R5327 VDD.n1535 VDD.n1516 185
R5328 VDD.n1856 VDD.n1855 185
R5329 VDD.n1855 VDD.n1500 185
R5330 VDD.n1853 VDD.n1491 185
R5331 VDD.n1513 VDD.n1491 185
R5332 VDD.n1915 VDD.n1914 185
R5333 VDD.n1914 VDD.n1913 185
R5334 VDD.n1916 VDD.n1485 185
R5335 VDD.n1510 VDD.n1485 185
R5336 VDD.n1930 VDD.n1929 185
R5337 VDD.n1931 VDD.n1930 185
R5338 VDD.n1488 VDD.n1486 185
R5339 VDD.n1486 VDD.n1472 185
R5340 VDD.n1924 VDD.n1923 185
R5341 VDD.n1923 VDD.n1469 185
R5342 VDD.n1921 VDD.n859 185
R5343 VDD.n859 VDD.n846 185
R5344 VDD.n2552 VDD.n2551 185
R5345 VDD.n2553 VDD.n2552 185
R5346 VDD.n2550 VDD.n860 185
R5347 VDD.n1465 VDD.n860 185
R5348 VDD.n1455 VDD.n862 185
R5349 VDD.n1463 VDD.n1455 185
R5350 VDD.n1995 VDD.n1994 185
R5351 VDD.n1994 VDD.n1993 185
R5352 VDD.n1996 VDD.n1450 185
R5353 VDD.n1450 VDD.n1433 185
R5354 VDD.n2010 VDD.n2009 185
R5355 VDD.n2011 VDD.n2010 185
R5356 VDD.n1453 VDD.n1451 185
R5357 VDD.n1451 VDD.n1429 185
R5358 VDD.n2004 VDD.n2003 185
R5359 VDD.n2003 VDD.n1412 185
R5360 VDD.n2001 VDD.n1397 185
R5361 VDD.n1426 VDD.n1397 185
R5362 VDD.n2080 VDD.n2079 185
R5363 VDD.n2079 VDD.n2078 185
R5364 VDD.n2081 VDD.n1391 185
R5365 VDD.n1423 VDD.n1391 185
R5366 VDD.n2091 VDD.n2090 185
R5367 VDD.n2092 VDD.n2091 185
R5368 VDD.n1394 VDD.n1392 185
R5369 VDD.n1392 VDD.n1370 185
R5370 VDD.n2085 VDD.n1363 185
R5371 VDD.n2095 VDD.n1363 185
R5372 VDD.n2114 VDD.n2113 185
R5373 VDD.n2113 VDD.n2112 185
R5374 VDD.n1360 VDD.n1359 185
R5375 VDD.n1359 VDD.n1339 185
R5376 VDD.n2121 VDD.n2120 185
R5377 VDD.n2122 VDD.n2121 185
R5378 VDD.n1200 VDD.n1198 185
R5379 VDD.n1333 VDD.n1200 185
R5380 VDD.n2542 VDD.n2541 185
R5381 VDD.n2541 VDD.n2540 185
R5382 VDD.n1201 VDD.n1199 185
R5383 VDD.n1330 VDD.n1201 185
R5384 VDD.n2529 VDD.n2528 185
R5385 VDD.n2530 VDD.n2529 185
R5386 VDD.n1219 VDD.n1217 185
R5387 VDD.n1326 VDD.n1217 185
R5388 VDD.n2523 VDD.n2522 185
R5389 VDD.n2522 VDD.n2521 185
R5390 VDD.n1250 VDD.n1222 185
R5391 VDD.n2382 VDD.n1222 185
R5392 VDD.n1253 VDD.n1252 185
R5393 VDD.n1252 VDD.n1232 185
R5394 VDD.n1254 VDD.n1245 185
R5395 VDD.n1245 VDD.n1241 185
R5396 VDD.n2506 VDD.n2505 185
R5397 VDD.n2507 VDD.n2506 185
R5398 VDD.n1248 VDD.n1246 185
R5399 VDD.n2174 VDD.n1246 185
R5400 VDD.n2500 VDD.n2499 185
R5401 VDD.n2499 VDD.n2498 185
R5402 VDD.n2195 VDD.n1260 185
R5403 VDD.n1323 VDD.n1260 185
R5404 VDD.n2199 VDD.n2198 185
R5405 VDD.n2199 VDD.n1273 185
R5406 VDD.n2201 VDD.n2200 185
R5407 VDD.n2200 VDD.n1319 185
R5408 VDD.n2192 VDD.n2191 185
R5409 VDD.n2191 VDD.n1286 185
R5410 VDD.n2206 VDD.n2205 185
R5411 VDD.n2206 VDD.n1317 185
R5412 VDD.n2207 VDD.n2190 185
R5413 VDD.n2207 VDD.n1292 185
R5414 VDD.n2209 VDD.n2208 185
R5415 VDD.n2208 VDD.n1295 185
R5416 VDD.n2210 VDD.n2188 185
R5417 VDD.n2188 VDD.n1314 185
R5418 VDD.n2347 VDD.n2346 185
R5419 VDD.n2348 VDD.n2347 185
R5420 VDD.n2345 VDD.n2189 185
R5421 VDD.n2189 VDD.n2187 185
R5422 VDD.n2344 VDD.n2343 185
R5423 VDD.n2343 VDD.n2342 185
R5424 VDD.n2212 VDD.n2211 185
R5425 VDD.n2341 VDD.n2212 185
R5426 VDD.n2339 VDD.n2338 185
R5427 VDD.n2340 VDD.n2339 185
R5428 VDD.n2337 VDD.n2217 185
R5429 VDD.n2217 VDD.n2216 185
R5430 VDD.n2336 VDD.n2335 185
R5431 VDD.n2335 VDD.n2334 185
R5432 VDD.n2219 VDD.n2218 185
R5433 VDD.n2333 VDD.n2219 185
R5434 VDD.n2331 VDD.n2330 185
R5435 VDD.n2332 VDD.n2331 185
R5436 VDD.n2329 VDD.n2223 185
R5437 VDD.n2226 VDD.n2223 185
R5438 VDD.n2328 VDD.n2327 185
R5439 VDD.n2327 VDD.n2326 185
R5440 VDD.n2225 VDD.n2224 185
R5441 VDD.n2325 VDD.n2225 185
R5442 VDD.n2323 VDD.n2322 185
R5443 VDD.n2324 VDD.n2323 185
R5444 VDD.n2321 VDD.n2231 185
R5445 VDD.n2231 VDD.n2230 185
R5446 VDD.n2320 VDD.n2319 185
R5447 VDD.n2319 VDD.n2318 185
R5448 VDD.n2233 VDD.n2232 185
R5449 VDD.n2317 VDD.n2233 185
R5450 VDD.n2315 VDD.n2314 185
R5451 VDD.n2316 VDD.n2315 185
R5452 VDD.n2313 VDD.n2238 185
R5453 VDD.n2238 VDD.n2237 185
R5454 VDD.n2312 VDD.n2311 185
R5455 VDD.n2311 VDD.n2310 185
R5456 VDD.n2240 VDD.n2239 185
R5457 VDD.n2309 VDD.n2240 185
R5458 VDD.n2306 VDD.n2305 185
R5459 VDD.n2304 VDD.n2251 185
R5460 VDD.n2303 VDD.n2250 185
R5461 VDD.n2308 VDD.n2250 185
R5462 VDD.n2302 VDD.n2301 185
R5463 VDD.n2300 VDD.n2299 185
R5464 VDD.n2298 VDD.n2297 185
R5465 VDD.n2296 VDD.n2295 185
R5466 VDD.n2294 VDD.n2293 185
R5467 VDD.n2292 VDD.n2291 185
R5468 VDD.n2290 VDD.n2289 185
R5469 VDD.n2288 VDD.n2287 185
R5470 VDD.n2286 VDD.n2285 185
R5471 VDD.n2284 VDD.n2283 185
R5472 VDD.n2282 VDD.n2281 185
R5473 VDD.n2280 VDD.n2279 185
R5474 VDD.n2278 VDD.n2277 185
R5475 VDD.n2276 VDD.n2275 185
R5476 VDD.n2274 VDD.n2242 185
R5477 VDD.n2309 VDD.n2242 185
R5478 VDD.n2273 VDD.n2241 185
R5479 VDD.n2310 VDD.n2241 185
R5480 VDD.n2272 VDD.n2271 185
R5481 VDD.n2271 VDD.n2237 185
R5482 VDD.n2270 VDD.n2236 185
R5483 VDD.n2316 VDD.n2236 185
R5484 VDD.n2269 VDD.n2235 185
R5485 VDD.n2317 VDD.n2235 185
R5486 VDD.n2268 VDD.n2234 185
R5487 VDD.n2318 VDD.n2234 185
R5488 VDD.n2267 VDD.n2266 185
R5489 VDD.n2266 VDD.n2230 185
R5490 VDD.n2265 VDD.n2229 185
R5491 VDD.n2324 VDD.n2229 185
R5492 VDD.n2264 VDD.n2228 185
R5493 VDD.n2325 VDD.n2228 185
R5494 VDD.n2263 VDD.n2227 185
R5495 VDD.n2326 VDD.n2227 185
R5496 VDD.n2262 VDD.n2261 185
R5497 VDD.n2261 VDD.n2226 185
R5498 VDD.n2260 VDD.n2222 185
R5499 VDD.n2332 VDD.n2222 185
R5500 VDD.n2259 VDD.n2221 185
R5501 VDD.n2333 VDD.n2221 185
R5502 VDD.n2258 VDD.n2220 185
R5503 VDD.n2334 VDD.n2220 185
R5504 VDD.n2257 VDD.n2256 185
R5505 VDD.n2256 VDD.n2216 185
R5506 VDD.n2255 VDD.n2215 185
R5507 VDD.n2340 VDD.n2215 185
R5508 VDD.n2254 VDD.n2214 185
R5509 VDD.n2341 VDD.n2214 185
R5510 VDD.n2253 VDD.n2213 185
R5511 VDD.n2342 VDD.n2213 185
R5512 VDD.n2252 VDD.n2185 185
R5513 VDD.n2187 VDD.n2185 185
R5514 VDD.n2349 VDD.n2186 185
R5515 VDD.n2349 VDD.n2348 185
R5516 VDD.n2350 VDD.n2184 185
R5517 VDD.n2350 VDD.n1314 185
R5518 VDD.n2352 VDD.n2351 185
R5519 VDD.n2351 VDD.n1295 185
R5520 VDD.n2353 VDD.n2183 185
R5521 VDD.n2183 VDD.n1292 185
R5522 VDD.n2355 VDD.n2354 185
R5523 VDD.n2355 VDD.n1317 185
R5524 VDD.n2357 VDD.n2356 185
R5525 VDD.n2356 VDD.n1286 185
R5526 VDD.n2180 VDD.n2179 185
R5527 VDD.n2179 VDD.n1319 185
R5528 VDD.n2363 VDD.n2362 185
R5529 VDD.n2363 VDD.n1273 185
R5530 VDD.n2365 VDD.n2364 185
R5531 VDD.n2364 VDD.n1323 185
R5532 VDD.n2367 VDD.n1262 185
R5533 VDD.n2498 VDD.n1262 185
R5534 VDD.n2176 VDD.n2175 185
R5535 VDD.n2175 VDD.n2174 185
R5536 VDD.n2372 VDD.n1243 185
R5537 VDD.n2507 VDD.n1243 185
R5538 VDD.n2375 VDD.n2374 185
R5539 VDD.n2374 VDD.n1241 185
R5540 VDD.n2159 VDD.n2157 185
R5541 VDD.n2157 VDD.n1232 185
R5542 VDD.n2381 VDD.n2380 185
R5543 VDD.n2382 VDD.n2381 185
R5544 VDD.n2168 VDD.n1223 185
R5545 VDD.n2521 VDD.n1223 185
R5546 VDD.n2167 VDD.n1215 185
R5547 VDD.n1326 VDD.n1215 185
R5548 VDD.n2532 VDD.n2531 185
R5549 VDD.n2531 VDD.n2530 185
R5550 VDD.n1214 VDD.n1212 185
R5551 VDD.n1330 VDD.n1214 185
R5552 VDD.n1353 VDD.n1202 185
R5553 VDD.n2540 VDD.n1202 185
R5554 VDD.n1356 VDD.n1355 185
R5555 VDD.n1356 VDD.n1333 185
R5556 VDD.n2124 VDD.n2123 185
R5557 VDD.n2123 VDD.n2122 185
R5558 VDD.n1352 VDD.n1350 185
R5559 VDD.n1352 VDD.n1339 185
R5560 VDD.n1383 VDD.n1365 185
R5561 VDD.n2112 VDD.n1365 185
R5562 VDD.n2097 VDD.n2096 185
R5563 VDD.n2096 VDD.n2095 185
R5564 VDD.n2094 VDD.n1381 185
R5565 VDD.n2094 VDD.n1370 185
R5566 VDD.n2093 VDD.n1389 185
R5567 VDD.n2093 VDD.n2092 185
R5568 VDD.n2069 VDD.n1387 185
R5569 VDD.n1423 VDD.n1387 185
R5570 VDD.n2067 VDD.n1398 185
R5571 VDD.n2078 VDD.n1398 185
R5572 VDD.n2013 VDD.n1408 185
R5573 VDD.n2013 VDD.n1426 185
R5574 VDD.n2016 VDD.n2015 185
R5575 VDD.n2016 VDD.n1412 185
R5576 VDD.n2018 VDD.n2017 185
R5577 VDD.n2017 VDD.n1429 185
R5578 VDD.n2012 VDD.n1444 185
R5579 VDD.n2012 VDD.n2011 185
R5580 VDD.n1976 VDD.n1448 185
R5581 VDD.n1448 VDD.n1433 185
R5582 VDD.n1974 VDD.n1456 185
R5583 VDD.n1993 VDD.n1456 185
R5584 VDD.n1972 VDD.n1971 185
R5585 VDD.n1971 VDD.n1463 185
R5586 VDD.n857 VDD.n855 185
R5587 VDD.n1465 VDD.n857 185
R5588 VDD.n2555 VDD.n2554 185
R5589 VDD.n2554 VDD.n2553 185
R5590 VDD.n856 VDD.n854 185
R5591 VDD.n856 VDD.n846 185
R5592 VDD.n1935 VDD.n1934 185
R5593 VDD.n1934 VDD.n1469 185
R5594 VDD.n1933 VDD.n1479 185
R5595 VDD.n1933 VDD.n1472 185
R5596 VDD.n1932 VDD.n1483 185
R5597 VDD.n1932 VDD.n1931 185
R5598 VDD.n1719 VDD.n1481 185
R5599 VDD.n1510 VDD.n1481 185
R5600 VDD.n1716 VDD.n1492 185
R5601 VDD.n1913 VDD.n1492 185
R5602 VDD.n1725 VDD.n1724 185
R5603 VDD.n1725 VDD.n1513 185
R5604 VDD.n1727 VDD.n1726 185
R5605 VDD.n1726 VDD.n1500 185
R5606 VDD.n1715 VDD.n1712 185
R5607 VDD.n1715 VDD.n1516 185
R5608 VDD.n1732 VDD.n1533 185
R5609 VDD.n1863 VDD.n1533 185
R5610 VDD.n1735 VDD.n1734 185
R5611 VDD.n1734 VDD.n1520 185
R5612 VDD.n1710 VDD.n1541 185
R5613 VDD.n1845 VDD.n1541 185
R5614 VDD.n1741 VDD.n1740 185
R5615 VDD.n1741 VDD.n1527 185
R5616 VDD.n1743 VDD.n1742 185
R5617 VDD.n1742 VDD.n1544 185
R5618 VDD.n1744 VDD.n1566 185
R5619 VDD.n1760 VDD.n1566 185
R5620 VDD.n1746 VDD.n1745 185
R5621 VDD.n1745 VDD.n1557 185
R5622 VDD.n1747 VDD.n1573 185
R5623 VDD.n1573 VDD.n1548 185
R5624 VDD.n1749 VDD.n1748 185
R5625 VDD.n1750 VDD.n1749 185
R5626 VDD.n1708 VDD.n1572 185
R5627 VDD.n1572 VDD.n1571 185
R5628 VDD.n1707 VDD.n1706 185
R5629 VDD.n1706 VDD.n1705 185
R5630 VDD.n1575 VDD.n1574 185
R5631 VDD.n1576 VDD.n1575 185
R5632 VDD.n1697 VDD.n1696 185
R5633 VDD.n1698 VDD.n1697 185
R5634 VDD.n1695 VDD.n1581 185
R5635 VDD.n1581 VDD.n1580 185
R5636 VDD.n1694 VDD.n1693 185
R5637 VDD.n1693 VDD.n1692 185
R5638 VDD.n1583 VDD.n1582 185
R5639 VDD.n1685 VDD.n1583 185
R5640 VDD.n1684 VDD.n1683 185
R5641 VDD.n1686 VDD.n1684 185
R5642 VDD.n1682 VDD.n1587 185
R5643 VDD.n1590 VDD.n1587 185
R5644 VDD.n1681 VDD.n1680 185
R5645 VDD.n1680 VDD.n1679 185
R5646 VDD.n1589 VDD.n1588 185
R5647 VDD.n1672 VDD.n1589 185
R5648 VDD.n1671 VDD.n1670 185
R5649 VDD.n1673 VDD.n1671 185
R5650 VDD.n1669 VDD.n1595 185
R5651 VDD.n1595 VDD.n1594 185
R5652 VDD.n1668 VDD.n1667 185
R5653 VDD.n1667 VDD.n1666 185
R5654 VDD.n1597 VDD.n1596 185
R5655 VDD.n1598 VDD.n1597 185
R5656 VDD.n1659 VDD.n1658 185
R5657 VDD.n1660 VDD.n1659 185
R5658 VDD.n1657 VDD.n1603 185
R5659 VDD.n1603 VDD.n1602 185
R5660 VDD.n1656 VDD.n1655 185
R5661 VDD.n1655 VDD.n1654 185
R5662 VDD.n1605 VDD.n1604 185
R5663 VDD.n1606 VDD.n1605 185
R5664 VDD.n5982 VDD.n5703 185
R5665 VDD.n5981 VDD.n5980 185
R5666 VDD.n5978 VDD.n5704 185
R5667 VDD.n5976 VDD.n5975 185
R5668 VDD.n5974 VDD.n5705 185
R5669 VDD.n5973 VDD.n5972 185
R5670 VDD.n5970 VDD.n5706 185
R5671 VDD.n5968 VDD.n5967 185
R5672 VDD.n5708 VDD.n5707 185
R5673 VDD.n5962 VDD.n5961 185
R5674 VDD.n5959 VDD.n5958 185
R5675 VDD.n5957 VDD.n5956 185
R5676 VDD.n5955 VDD.n5913 185
R5677 VDD.n5953 VDD.n5952 185
R5678 VDD.n5951 VDD.n5914 185
R5679 VDD.n5950 VDD.n5949 185
R5680 VDD.n5947 VDD.n5946 185
R5681 VDD.n5947 VDD.n5702 185
R5682 VDD.n5945 VDD.n5701 185
R5683 VDD.n5985 VDD.n5701 185
R5684 VDD.n5944 VDD.n5943 185
R5685 VDD.n5943 VDD.n5696 185
R5686 VDD.n5942 VDD.n5695 185
R5687 VDD.n5991 VDD.n5695 185
R5688 VDD.n5941 VDD.n5940 185
R5689 VDD.n5940 VDD.n5690 185
R5690 VDD.n5939 VDD.n5689 185
R5691 VDD.n5997 VDD.n5689 185
R5692 VDD.n5938 VDD.n5937 185
R5693 VDD.n5937 VDD.n5687 185
R5694 VDD.n5936 VDD.n5683 185
R5695 VDD.n6003 VDD.n5683 185
R5696 VDD.n5935 VDD.n5934 185
R5697 VDD.n5934 VDD.n5678 185
R5698 VDD.n5933 VDD.n5677 185
R5699 VDD.n6009 VDD.n5677 185
R5700 VDD.n5932 VDD.n5931 185
R5701 VDD.n5931 VDD.n5675 185
R5702 VDD.n5930 VDD.n5671 185
R5703 VDD.n6015 VDD.n5671 185
R5704 VDD.n5929 VDD.n5928 185
R5705 VDD.n5928 VDD.n5666 185
R5706 VDD.n5927 VDD.n5665 185
R5707 VDD.n6021 VDD.n5665 185
R5708 VDD.n5926 VDD.n5925 185
R5709 VDD.n5925 VDD.n5663 185
R5710 VDD.n5924 VDD.n5659 185
R5711 VDD.n6027 VDD.n5659 185
R5712 VDD.n5923 VDD.n5922 185
R5713 VDD.n5922 VDD.n5654 185
R5714 VDD.n5921 VDD.n5653 185
R5715 VDD.n6033 VDD.n5653 185
R5716 VDD.n5920 VDD.n5919 185
R5717 VDD.n5919 VDD.n5651 185
R5718 VDD.n5918 VDD.n5647 185
R5719 VDD.n6039 VDD.n5647 185
R5720 VDD.n5917 VDD.n5916 185
R5721 VDD.n5916 VDD.n5612 185
R5722 VDD.n5915 VDD.n5611 185
R5723 VDD.n6045 VDD.n5611 185
R5724 VDD.n5600 VDD.n5599 185
R5725 VDD.n5603 VDD.n5600 185
R5726 VDD.n6053 VDD.n6052 185
R5727 VDD.n6052 VDD.n6051 185
R5728 VDD.n6054 VDD.n5598 185
R5729 VDD.n5601 VDD.n5598 185
R5730 VDD.n6056 VDD.n6055 185
R5731 VDD.n6058 VDD.n5596 185
R5732 VDD.n6060 VDD.n6059 185
R5733 VDD.n6061 VDD.n5595 185
R5734 VDD.n6063 VDD.n6062 185
R5735 VDD.n6065 VDD.n5592 185
R5736 VDD.n6067 VDD.n6066 185
R5737 VDD.n5623 VDD.n5591 185
R5738 VDD.n5625 VDD.n5624 185
R5739 VDD.n5627 VDD.n5620 185
R5740 VDD.n5629 VDD.n5628 185
R5741 VDD.n5631 VDD.n5618 185
R5742 VDD.n5633 VDD.n5632 185
R5743 VDD.n5634 VDD.n5617 185
R5744 VDD.n5636 VDD.n5635 185
R5745 VDD.n5638 VDD.n5616 185
R5746 VDD.n5639 VDD.n5615 185
R5747 VDD.n5639 VDD.n5594 185
R5748 VDD.n5641 VDD.n5640 185
R5749 VDD.n5640 VDD.n5601 185
R5750 VDD.n5642 VDD.n5604 185
R5751 VDD.n6051 VDD.n5604 185
R5752 VDD.n5643 VDD.n5613 185
R5753 VDD.n5613 VDD.n5603 185
R5754 VDD.n6044 VDD.n6043 185
R5755 VDD.n6045 VDD.n6044 185
R5756 VDD.n6042 VDD.n5614 185
R5757 VDD.n5614 VDD.n5612 185
R5758 VDD.n6041 VDD.n6040 185
R5759 VDD.n6040 VDD.n6039 185
R5760 VDD.n5645 VDD.n5644 185
R5761 VDD.n5651 VDD.n5645 185
R5762 VDD.n6032 VDD.n6031 185
R5763 VDD.n6033 VDD.n6032 185
R5764 VDD.n6030 VDD.n5655 185
R5765 VDD.n5655 VDD.n5654 185
R5766 VDD.n6029 VDD.n6028 185
R5767 VDD.n6028 VDD.n6027 185
R5768 VDD.n5657 VDD.n5656 185
R5769 VDD.n5663 VDD.n5657 185
R5770 VDD.n6020 VDD.n6019 185
R5771 VDD.n6021 VDD.n6020 185
R5772 VDD.n6018 VDD.n5667 185
R5773 VDD.n5667 VDD.n5666 185
R5774 VDD.n6017 VDD.n6016 185
R5775 VDD.n6016 VDD.n6015 185
R5776 VDD.n5669 VDD.n5668 185
R5777 VDD.n5675 VDD.n5669 185
R5778 VDD.n6008 VDD.n6007 185
R5779 VDD.n6009 VDD.n6008 185
R5780 VDD.n6006 VDD.n5679 185
R5781 VDD.n5679 VDD.n5678 185
R5782 VDD.n6005 VDD.n6004 185
R5783 VDD.n6004 VDD.n6003 185
R5784 VDD.n5681 VDD.n5680 185
R5785 VDD.n5687 VDD.n5681 185
R5786 VDD.n5996 VDD.n5995 185
R5787 VDD.n5997 VDD.n5996 185
R5788 VDD.n5994 VDD.n5691 185
R5789 VDD.n5691 VDD.n5690 185
R5790 VDD.n5993 VDD.n5992 185
R5791 VDD.n5992 VDD.n5991 185
R5792 VDD.n5693 VDD.n5692 185
R5793 VDD.n5696 VDD.n5693 185
R5794 VDD.n5984 VDD.n5983 185
R5795 VDD.n5985 VDD.n5984 185
R5796 VDD.n5783 VDD.n5767 185
R5797 VDD.n5783 VDD.n5594 185
R5798 VDD.n5782 VDD.n5768 185
R5799 VDD.n5780 VDD.n5779 185
R5800 VDD.n5778 VDD.n5769 185
R5801 VDD.n5777 VDD.n5776 185
R5802 VDD.n5774 VDD.n5770 185
R5803 VDD.n5772 VDD.n5771 185
R5804 VDD.n5607 VDD.n5605 185
R5805 VDD.n5605 VDD.n5601 185
R5806 VDD.n6050 VDD.n6049 185
R5807 VDD.n6051 VDD.n6050 185
R5808 VDD.n6048 VDD.n5606 185
R5809 VDD.n5606 VDD.n5603 185
R5810 VDD.n6047 VDD.n6046 185
R5811 VDD.n6046 VDD.n6045 185
R5812 VDD.n5609 VDD.n5608 185
R5813 VDD.n5612 VDD.n5609 185
R5814 VDD.n6038 VDD.n6037 185
R5815 VDD.n6039 VDD.n6038 185
R5816 VDD.n6036 VDD.n5648 185
R5817 VDD.n5651 VDD.n5648 185
R5818 VDD.n6035 VDD.n6034 185
R5819 VDD.n6034 VDD.n6033 185
R5820 VDD.n5650 VDD.n5649 185
R5821 VDD.n5654 VDD.n5650 185
R5822 VDD.n6026 VDD.n6025 185
R5823 VDD.n6027 VDD.n6026 185
R5824 VDD.n6024 VDD.n5660 185
R5825 VDD.n5663 VDD.n5660 185
R5826 VDD.n6023 VDD.n6022 185
R5827 VDD.n6022 VDD.n6021 185
R5828 VDD.n5662 VDD.n5661 185
R5829 VDD.n5666 VDD.n5662 185
R5830 VDD.n6014 VDD.n6013 185
R5831 VDD.n6015 VDD.n6014 185
R5832 VDD.n6012 VDD.n5672 185
R5833 VDD.n5675 VDD.n5672 185
R5834 VDD.n6011 VDD.n6010 185
R5835 VDD.n6010 VDD.n6009 185
R5836 VDD.n5674 VDD.n5673 185
R5837 VDD.n5678 VDD.n5674 185
R5838 VDD.n6002 VDD.n6001 185
R5839 VDD.n6003 VDD.n6002 185
R5840 VDD.n6000 VDD.n5684 185
R5841 VDD.n5687 VDD.n5684 185
R5842 VDD.n5999 VDD.n5998 185
R5843 VDD.n5998 VDD.n5997 185
R5844 VDD.n5686 VDD.n5685 185
R5845 VDD.n5690 VDD.n5686 185
R5846 VDD.n5990 VDD.n5989 185
R5847 VDD.n5991 VDD.n5990 185
R5848 VDD.n5988 VDD.n5697 185
R5849 VDD.n5697 VDD.n5696 185
R5850 VDD.n5987 VDD.n5986 185
R5851 VDD.n5986 VDD.n5985 185
R5852 VDD.n5699 VDD.n5698 185
R5853 VDD.n5730 VDD.n5729 185
R5854 VDD.n5731 VDD.n5727 185
R5855 VDD.n5727 VDD.n5702 185
R5856 VDD.n5733 VDD.n5732 185
R5857 VDD.n5735 VDD.n5726 185
R5858 VDD.n5738 VDD.n5737 185
R5859 VDD.n5739 VDD.n5725 185
R5860 VDD.n5741 VDD.n5740 185
R5861 VDD.n5743 VDD.n5718 185
R5862 VDD.n5870 VDD.n5869 185
R5863 VDD.n5867 VDD.n5866 185
R5864 VDD.n5865 VDD.n5744 185
R5865 VDD.n5864 VDD.n5863 185
R5866 VDD.n5861 VDD.n5745 185
R5867 VDD.n5859 VDD.n5858 185
R5868 VDD.n5857 VDD.n5746 185
R5869 VDD.n5856 VDD.n5855 185
R5870 VDD.n5853 VDD.n5700 185
R5871 VDD.n5985 VDD.n5700 185
R5872 VDD.n5852 VDD.n5851 185
R5873 VDD.n5851 VDD.n5696 185
R5874 VDD.n5850 VDD.n5694 185
R5875 VDD.n5991 VDD.n5694 185
R5876 VDD.n5849 VDD.n5848 185
R5877 VDD.n5848 VDD.n5690 185
R5878 VDD.n5847 VDD.n5688 185
R5879 VDD.n5997 VDD.n5688 185
R5880 VDD.n5846 VDD.n5845 185
R5881 VDD.n5845 VDD.n5687 185
R5882 VDD.n5844 VDD.n5682 185
R5883 VDD.n6003 VDD.n5682 185
R5884 VDD.n5843 VDD.n5842 185
R5885 VDD.n5842 VDD.n5678 185
R5886 VDD.n5841 VDD.n5676 185
R5887 VDD.n6009 VDD.n5676 185
R5888 VDD.n5840 VDD.n5839 185
R5889 VDD.n5839 VDD.n5675 185
R5890 VDD.n5838 VDD.n5670 185
R5891 VDD.n6015 VDD.n5670 185
R5892 VDD.n5837 VDD.n5836 185
R5893 VDD.n5836 VDD.n5666 185
R5894 VDD.n5835 VDD.n5664 185
R5895 VDD.n6021 VDD.n5664 185
R5896 VDD.n5834 VDD.n5833 185
R5897 VDD.n5833 VDD.n5663 185
R5898 VDD.n5832 VDD.n5658 185
R5899 VDD.n6027 VDD.n5658 185
R5900 VDD.n5831 VDD.n5830 185
R5901 VDD.n5830 VDD.n5654 185
R5902 VDD.n5829 VDD.n5652 185
R5903 VDD.n6033 VDD.n5652 185
R5904 VDD.n5828 VDD.n5827 185
R5905 VDD.n5827 VDD.n5651 185
R5906 VDD.n5826 VDD.n5646 185
R5907 VDD.n6039 VDD.n5646 185
R5908 VDD.n5825 VDD.n5824 185
R5909 VDD.n5824 VDD.n5612 185
R5910 VDD.n5823 VDD.n5610 185
R5911 VDD.n6045 VDD.n5610 185
R5912 VDD.n5822 VDD.n5821 185
R5913 VDD.n5821 VDD.n5603 185
R5914 VDD.n5820 VDD.n5602 185
R5915 VDD.n6051 VDD.n5602 185
R5916 VDD.n5819 VDD.n5818 185
R5917 VDD.n5818 VDD.n5601 185
R5918 VDD.n5817 VDD.n5747 185
R5919 VDD.n5815 VDD.n5814 185
R5920 VDD.n5813 VDD.n5748 185
R5921 VDD.n5812 VDD.n5811 185
R5922 VDD.n5809 VDD.n5749 185
R5923 VDD.n5807 VDD.n5806 185
R5924 VDD.n5805 VDD.n5750 185
R5925 VDD.n5788 VDD.n5751 185
R5926 VDD.n5791 VDD.n5790 185
R5927 VDD.n5792 VDD.n5784 185
R5928 VDD.n8039 VDD.n6859 185
R5929 VDD.n8038 VDD.n8037 185
R5930 VDD.n6861 VDD.n6860 185
R5931 VDD.n7970 VDD.n7969 185
R5932 VDD.n7972 VDD.n7971 185
R5933 VDD.n7974 VDD.n7973 185
R5934 VDD.n7976 VDD.n7975 185
R5935 VDD.n7978 VDD.n7977 185
R5936 VDD.n7980 VDD.n7979 185
R5937 VDD.n7982 VDD.n7981 185
R5938 VDD.n7984 VDD.n7983 185
R5939 VDD.n7986 VDD.n7985 185
R5940 VDD.n7988 VDD.n7987 185
R5941 VDD.n7990 VDD.n7989 185
R5942 VDD.n7992 VDD.n7991 185
R5943 VDD.n7994 VDD.n7993 185
R5944 VDD.n7995 VDD.n6876 185
R5945 VDD.n8035 VDD.n6876 185
R5946 VDD.n7996 VDD.n6857 185
R5947 VDD.n8042 VDD.n6857 185
R5948 VDD.n7998 VDD.n7997 185
R5949 VDD.n7999 VDD.n7998 185
R5950 VDD.n7968 VDD.n6851 185
R5951 VDD.n8048 VDD.n6851 185
R5952 VDD.n7967 VDD.n7966 185
R5953 VDD.n7966 VDD.n7965 185
R5954 VDD.n6881 VDD.n6838 185
R5955 VDD.n8054 VDD.n6838 185
R5956 VDD.n7958 VDD.n7957 185
R5957 VDD.n7959 VDD.n7958 185
R5958 VDD.n7956 VDD.n6827 185
R5959 VDD.n8060 VDD.n6827 185
R5960 VDD.n7955 VDD.n7954 185
R5961 VDD.n7954 VDD.n6824 185
R5962 VDD.n7953 VDD.n7952 185
R5963 VDD.n7953 VDD.n6807 185
R5964 VDD.n7951 VDD.n6805 185
R5965 VDD.n8071 VDD.n6805 185
R5966 VDD.n7950 VDD.n6797 185
R5967 VDD.n8077 VDD.n6797 185
R5968 VDD.n7949 VDD.n7948 185
R5969 VDD.n7948 VDD.n7947 185
R5970 VDD.n7719 VDD.n6788 185
R5971 VDD.n8083 VDD.n6788 185
R5972 VDD.n7718 VDD.n7717 185
R5973 VDD.n7717 VDD.n7716 185
R5974 VDD.n6888 VDD.n6887 185
R5975 VDD.n6888 VDD.n6779 185
R5976 VDD.n7707 VDD.n7706 185
R5977 VDD.n7708 VDD.n7707 185
R5978 VDD.n7705 VDD.n6767 185
R5979 VDD.n8102 VDD.n6767 185
R5980 VDD.n7704 VDD.n7703 185
R5981 VDD.n7703 VDD.n7702 185
R5982 VDD.n6895 VDD.n6894 185
R5983 VDD.n6921 VDD.n6895 185
R5984 VDD.n7671 VDD.n6904 185
R5985 VDD.n7694 VDD.n6904 185
R5986 VDD.n7673 VDD.n7672 185
R5987 VDD.n7674 VDD.n7673 185
R5988 VDD.n7670 VDD.n6930 185
R5989 VDD.n6930 VDD.n6927 185
R5990 VDD.n7669 VDD.n7668 185
R5991 VDD.n7668 VDD.n7667 185
R5992 VDD.n6932 VDD.n6931 185
R5993 VDD.n6953 VDD.n6932 185
R5994 VDD.n7613 VDD.n7612 185
R5995 VDD.n7614 VDD.n7613 185
R5996 VDD.n7611 VDD.n6963 185
R5997 VDD.n7640 VDD.n6963 185
R5998 VDD.n7610 VDD.n7609 185
R5999 VDD.n7609 VDD.n7608 185
R6000 VDD.n6988 VDD.n6977 185
R6001 VDD.n7621 VDD.n6977 185
R6002 VDD.n7593 VDD.n7592 185
R6003 VDD.t316 VDD.n7593 185
R6004 VDD.n7591 VDD.n6993 185
R6005 VDD.n7012 VDD.n6993 185
R6006 VDD.n7590 VDD.n7589 185
R6007 VDD.n7589 VDD.n7588 185
R6008 VDD.n6995 VDD.n6994 185
R6009 VDD.n7555 VDD.n6995 185
R6010 VDD.n7513 VDD.n7027 185
R6011 VDD.n7546 VDD.n7027 185
R6012 VDD.n7515 VDD.n7514 185
R6013 VDD.n7518 VDD.n7515 185
R6014 VDD.n7512 VDD.n7029 185
R6015 VDD.n7029 VDD.n6421 185
R6016 VDD.n7511 VDD.n6410 185
R6017 VDD.n8125 VDD.n6410 185
R6018 VDD.n7510 VDD.n7509 185
R6019 VDD.n7509 VDD.n7508 185
R6020 VDD.n7031 VDD.n7030 185
R6021 VDD.n7505 VDD.n7031 185
R6022 VDD.n7457 VDD.n7074 185
R6023 VDD.n7074 VDD.n7047 185
R6024 VDD.n7459 VDD.n7458 185
R6025 VDD.n7460 VDD.n7459 185
R6026 VDD.n7456 VDD.n7057 185
R6027 VDD.n7475 VDD.n7057 185
R6028 VDD.n7455 VDD.n7454 185
R6029 VDD.n7454 VDD.n7453 185
R6030 VDD.n7075 VDD.n7065 185
R6031 VDD.n7468 VDD.n7065 185
R6032 VDD.n7446 VDD.n7445 185
R6033 VDD.n7447 VDD.n7446 185
R6034 VDD.n7444 VDD.n7080 185
R6035 VDD.n7427 VDD.n7080 185
R6036 VDD.n7443 VDD.n7442 185
R6037 VDD.n7442 VDD.n7441 185
R6038 VDD.n7082 VDD.n7081 185
R6039 VDD.n7407 VDD.n7082 185
R6040 VDD.n7397 VDD.n7092 185
R6041 VDD.n7434 VDD.n7092 185
R6042 VDD.n7399 VDD.n7398 185
R6043 VDD.n7400 VDD.n7399 185
R6044 VDD.n7396 VDD.n7108 185
R6045 VDD.n7355 VDD.n7108 185
R6046 VDD.n7395 VDD.n7394 185
R6047 VDD.n7110 VDD.n7109 185
R6048 VDD.n7325 VDD.n7324 185
R6049 VDD.n7327 VDD.n7326 185
R6050 VDD.n7329 VDD.n7328 185
R6051 VDD.n7331 VDD.n7330 185
R6052 VDD.n7333 VDD.n7332 185
R6053 VDD.n7335 VDD.n7334 185
R6054 VDD.n7337 VDD.n7336 185
R6055 VDD.n7339 VDD.n7338 185
R6056 VDD.n7341 VDD.n7340 185
R6057 VDD.n7343 VDD.n7342 185
R6058 VDD.n7345 VDD.n7344 185
R6059 VDD.n7347 VDD.n7346 185
R6060 VDD.n7349 VDD.n7348 185
R6061 VDD.n7351 VDD.n7350 185
R6062 VDD.n7352 VDD.n7112 185
R6063 VDD.n7392 VDD.n7112 185
R6064 VDD.n7354 VDD.n7353 185
R6065 VDD.n7355 VDD.n7354 185
R6066 VDD.n7095 VDD.n7093 185
R6067 VDD.n7400 VDD.n7093 185
R6068 VDD.n7433 VDD.n7432 185
R6069 VDD.n7434 VDD.n7433 185
R6070 VDD.n7431 VDD.n7094 185
R6071 VDD.n7407 VDD.n7094 185
R6072 VDD.n7430 VDD.n7085 185
R6073 VDD.n7441 VDD.n7085 185
R6074 VDD.n7429 VDD.n7428 185
R6075 VDD.n7428 VDD.n7427 185
R6076 VDD.n7068 VDD.n7066 185
R6077 VDD.n7447 VDD.n7066 185
R6078 VDD.n7467 VDD.n7466 185
R6079 VDD.n7468 VDD.n7467 185
R6080 VDD.n7465 VDD.n7067 185
R6081 VDD.n7453 VDD.n7067 185
R6082 VDD.n7464 VDD.n7058 185
R6083 VDD.n7475 VDD.n7058 185
R6084 VDD.n7462 VDD.n7070 185
R6085 VDD.n7460 VDD.n7070 185
R6086 VDD.n7071 VDD.n7033 185
R6087 VDD.n7047 VDD.n7033 185
R6088 VDD.n7506 VDD.n7034 185
R6089 VDD.n7506 VDD.n7505 185
R6090 VDD.n7507 VDD.n6404 185
R6091 VDD.n7508 VDD.n7507 185
R6092 VDD.n8127 VDD.n6405 185
R6093 VDD.n8125 VDD.n6405 185
R6094 VDD.n7516 VDD.n6406 185
R6095 VDD.n7516 VDD.n6421 185
R6096 VDD.n7517 VDD.n7024 185
R6097 VDD.n7518 VDD.n7517 185
R6098 VDD.n7548 VDD.n7021 185
R6099 VDD.n7546 VDD.n7021 185
R6100 VDD.n7554 VDD.n7553 185
R6101 VDD.n7555 VDD.n7554 185
R6102 VDD.n7552 VDD.n6998 185
R6103 VDD.n7588 VDD.n6998 185
R6104 VDD.n7551 VDD.n7550 185
R6105 VDD.n7550 VDD.n7012 185
R6106 VDD.n6980 VDD.n6978 185
R6107 VDD.t316 VDD.n6978 185
R6108 VDD.n7620 VDD.n7619 185
R6109 VDD.n7621 VDD.n7620 185
R6110 VDD.n7618 VDD.n6979 185
R6111 VDD.n7608 VDD.n6979 185
R6112 VDD.n7617 VDD.n6964 185
R6113 VDD.n7640 VDD.n6964 185
R6114 VDD.n7616 VDD.n7615 185
R6115 VDD.n7615 VDD.n7614 185
R6116 VDD.n6985 VDD.n6984 185
R6117 VDD.n6985 VDD.n6953 185
R6118 VDD.n6983 VDD.n6935 185
R6119 VDD.n7667 VDD.n6935 185
R6120 VDD.n6982 VDD.n6981 185
R6121 VDD.n6981 VDD.n6927 185
R6122 VDD.n6901 VDD.n6900 185
R6123 VDD.n7674 VDD.n6901 185
R6124 VDD.n7696 VDD.n7695 185
R6125 VDD.n7695 VDD.n7694 185
R6126 VDD.n7697 VDD.n6898 185
R6127 VDD.n6921 VDD.n6898 185
R6128 VDD.n7701 VDD.n7700 185
R6129 VDD.n7702 VDD.n7701 185
R6130 VDD.n7699 VDD.n6768 185
R6131 VDD.n8102 VDD.n6768 185
R6132 VDD.n6892 VDD.n6891 185
R6133 VDD.n7708 VDD.n6891 185
R6134 VDD.n7712 VDD.n7711 185
R6135 VDD.n7712 VDD.n6779 185
R6136 VDD.n7715 VDD.n7714 185
R6137 VDD.n7716 VDD.n7715 185
R6138 VDD.n7713 VDD.n6789 185
R6139 VDD.n8083 VDD.n6789 185
R6140 VDD.n6800 VDD.n6798 185
R6141 VDD.n7947 VDD.n6798 185
R6142 VDD.n8076 VDD.n8075 185
R6143 VDD.n8077 VDD.n8076 185
R6144 VDD.n6801 VDD.n6799 185
R6145 VDD.n8071 VDD.n6799 185
R6146 VDD.n6842 VDD.n6841 185
R6147 VDD.n6842 VDD.n6807 185
R6148 VDD.n6844 VDD.n6843 185
R6149 VDD.n6843 VDD.n6824 185
R6150 VDD.n6845 VDD.n6828 185
R6151 VDD.n8060 VDD.n6828 185
R6152 VDD.n6846 VDD.n6839 185
R6153 VDD.n7959 VDD.n6839 185
R6154 VDD.n8053 VDD.n8052 185
R6155 VDD.n8054 VDD.n8053 185
R6156 VDD.n8051 VDD.n6840 185
R6157 VDD.n7965 VDD.n6840 185
R6158 VDD.n8050 VDD.n8049 185
R6159 VDD.n8049 VDD.n8048 185
R6160 VDD.n6848 VDD.n6847 185
R6161 VDD.n7999 VDD.n6848 185
R6162 VDD.n8041 VDD.n8040 185
R6163 VDD.n8042 VDD.n8041 185
R6164 VDD.n6854 VDD.n6853 185
R6165 VDD.n8033 VDD.n8032 185
R6166 VDD.n8031 VDD.n6878 185
R6167 VDD.n8035 VDD.n6878 185
R6168 VDD.n8030 VDD.n8029 185
R6169 VDD.n8028 VDD.n8027 185
R6170 VDD.n8026 VDD.n8025 185
R6171 VDD.n8024 VDD.n8023 185
R6172 VDD.n8022 VDD.n8021 185
R6173 VDD.n8020 VDD.n8019 185
R6174 VDD.n8018 VDD.n8017 185
R6175 VDD.n8016 VDD.n8015 185
R6176 VDD.n8014 VDD.n8013 185
R6177 VDD.n8012 VDD.n8011 185
R6178 VDD.n8010 VDD.n8009 185
R6179 VDD.n8008 VDD.n8007 185
R6180 VDD.n8006 VDD.n8005 185
R6181 VDD.n8004 VDD.n8003 185
R6182 VDD.n8002 VDD.n6856 185
R6183 VDD.n8042 VDD.n6856 185
R6184 VDD.n8001 VDD.n8000 185
R6185 VDD.n8000 VDD.n7999 185
R6186 VDD.n6879 VDD.n6850 185
R6187 VDD.n8048 VDD.n6850 185
R6188 VDD.n7964 VDD.n7963 185
R6189 VDD.n7965 VDD.n7964 185
R6190 VDD.n7962 VDD.n6837 185
R6191 VDD.n8054 VDD.n6837 185
R6192 VDD.n7961 VDD.n7960 185
R6193 VDD.n7960 VDD.n7959 185
R6194 VDD.n6885 VDD.n6826 185
R6195 VDD.n8060 VDD.n6826 185
R6196 VDD.n6884 VDD.n6883 185
R6197 VDD.n6883 VDD.n6824 185
R6198 VDD.n6803 VDD.n6802 185
R6199 VDD.n6807 VDD.n6803 185
R6200 VDD.n8073 VDD.n8072 185
R6201 VDD.n8072 VDD.n8071 185
R6202 VDD.n8075 VDD.n6796 185
R6203 VDD.n8077 VDD.n6796 185
R6204 VDD.n7946 VDD.n6800 185
R6205 VDD.n7947 VDD.n7946 185
R6206 VDD.n7713 VDD.n6787 185
R6207 VDD.n8083 VDD.n6787 185
R6208 VDD.n7714 VDD.n6890 185
R6209 VDD.n7716 VDD.n6890 185
R6210 VDD.n7711 VDD.n7710 185
R6211 VDD.n7710 VDD.n6779 185
R6212 VDD.n7709 VDD.n6892 185
R6213 VDD.n7709 VDD.n7708 185
R6214 VDD.n7699 VDD.n6766 185
R6215 VDD.n8102 VDD.n6766 185
R6216 VDD.n7700 VDD.n6897 185
R6217 VDD.n7702 VDD.n6897 185
R6218 VDD.n6920 VDD.n6899 185
R6219 VDD.n6921 VDD.n6920 185
R6220 VDD.n7597 VDD.n6903 185
R6221 VDD.n7694 VDD.n6903 185
R6222 VDD.n7598 VDD.n6929 185
R6223 VDD.n7674 VDD.n6929 185
R6224 VDD.n7600 VDD.n7599 185
R6225 VDD.n7599 VDD.n6927 185
R6226 VDD.n7601 VDD.n6934 185
R6227 VDD.n7667 VDD.n6934 185
R6228 VDD.n7603 VDD.n7602 185
R6229 VDD.n7602 VDD.n6953 185
R6230 VDD.n7604 VDD.n6987 185
R6231 VDD.n7614 VDD.n6987 185
R6232 VDD.n7605 VDD.n6962 185
R6233 VDD.n7640 VDD.n6962 185
R6234 VDD.n7607 VDD.n7606 185
R6235 VDD.n7608 VDD.n7607 185
R6236 VDD.n7596 VDD.n6976 185
R6237 VDD.n7621 VDD.n6976 185
R6238 VDD.n7595 VDD.n7594 185
R6239 VDD.n7594 VDD.t316 185
R6240 VDD.n6991 VDD.n6990 185
R6241 VDD.n7012 VDD.n6991 185
R6242 VDD.n7022 VDD.n6997 185
R6243 VDD.n7588 VDD.n6997 185
R6244 VDD.n7023 VDD.n7020 185
R6245 VDD.n7555 VDD.n7020 185
R6246 VDD.n7548 VDD.n7547 185
R6247 VDD.n7547 VDD.n7546 185
R6248 VDD.n7025 VDD.n7024 185
R6249 VDD.n7518 VDD.n7025 185
R6250 VDD.n6408 VDD.n6406 185
R6251 VDD.n6421 VDD.n6408 185
R6252 VDD.n8127 VDD.n8126 185
R6253 VDD.n8126 VDD.n8125 185
R6254 VDD.n6407 VDD.n6404 185
R6255 VDD.n7508 VDD.n6407 185
R6256 VDD.n7036 VDD.n7034 185
R6257 VDD.n7505 VDD.n7036 185
R6258 VDD.n7072 VDD.n7071 185
R6259 VDD.n7072 VDD.n7047 185
R6260 VDD.n7462 VDD.n7461 185
R6261 VDD.n7461 VDD.n7460 185
R6262 VDD.n7069 VDD.n7056 185
R6263 VDD.n7475 VDD.n7056 185
R6264 VDD.n7452 VDD.n7451 185
R6265 VDD.n7453 VDD.n7452 185
R6266 VDD.n7450 VDD.n7064 185
R6267 VDD.n7468 VDD.n7064 185
R6268 VDD.n7449 VDD.n7448 185
R6269 VDD.n7448 VDD.n7447 185
R6270 VDD.n7078 VDD.n7077 185
R6271 VDD.n7427 VDD.n7078 185
R6272 VDD.n7404 VDD.n7084 185
R6273 VDD.n7441 VDD.n7084 185
R6274 VDD.n7406 VDD.n7405 185
R6275 VDD.n7407 VDD.n7406 185
R6276 VDD.n7403 VDD.n7091 185
R6277 VDD.n7434 VDD.n7091 185
R6278 VDD.n7402 VDD.n7401 185
R6279 VDD.n7401 VDD.n7400 185
R6280 VDD.n7106 VDD.n7105 185
R6281 VDD.n7355 VDD.n7106 185
R6282 VDD.n7360 VDD.n7359 185
R6283 VDD.n7362 VDD.n7361 185
R6284 VDD.n7364 VDD.n7363 185
R6285 VDD.n7366 VDD.n7365 185
R6286 VDD.n7368 VDD.n7367 185
R6287 VDD.n7370 VDD.n7369 185
R6288 VDD.n7372 VDD.n7371 185
R6289 VDD.n7374 VDD.n7373 185
R6290 VDD.n7376 VDD.n7375 185
R6291 VDD.n7378 VDD.n7377 185
R6292 VDD.n7380 VDD.n7379 185
R6293 VDD.n7382 VDD.n7381 185
R6294 VDD.n7384 VDD.n7383 185
R6295 VDD.n7386 VDD.n7385 185
R6296 VDD.n7388 VDD.n7387 185
R6297 VDD.n7389 VDD.n7357 185
R6298 VDD.n7391 VDD.n7390 185
R6299 VDD.n7392 VDD.n7391 185
R6300 VDD.n7358 VDD.n7356 185
R6301 VDD.n7356 VDD.n7355 185
R6302 VDD.n7089 VDD.n7088 185
R6303 VDD.n7400 VDD.n7089 185
R6304 VDD.n7436 VDD.n7435 185
R6305 VDD.n7435 VDD.n7434 185
R6306 VDD.n7437 VDD.n7086 185
R6307 VDD.n7407 VDD.n7086 185
R6308 VDD.n7440 VDD.n7439 185
R6309 VDD.n7441 VDD.n7440 185
R6310 VDD.n7438 VDD.n7087 185
R6311 VDD.n7427 VDD.n7087 185
R6312 VDD.n7062 VDD.n7061 185
R6313 VDD.n7447 VDD.n7062 185
R6314 VDD.n7470 VDD.n7469 185
R6315 VDD.n7469 VDD.n7468 185
R6316 VDD.n7471 VDD.n7059 185
R6317 VDD.n7453 VDD.n7059 185
R6318 VDD.n7474 VDD.n7473 185
R6319 VDD.n7475 VDD.n7474 185
R6320 VDD.n7472 VDD.n7060 185
R6321 VDD.n7460 VDD.n7060 185
R6322 VDD.n7038 VDD.n7037 185
R6323 VDD.n7047 VDD.n7037 185
R6324 VDD.n7504 VDD.n7503 185
R6325 VDD.n7505 VDD.n7504 185
R6326 VDD.n7039 VDD.n6411 185
R6327 VDD.n7508 VDD.n6411 185
R6328 VDD.n8124 VDD.n8123 185
R6329 VDD.n8125 VDD.n8124 185
R6330 VDD.n6414 VDD.n6412 185
R6331 VDD.n6421 VDD.n6412 185
R6332 VDD.n7521 VDD.n7519 185
R6333 VDD.n7519 VDD.n7518 185
R6334 VDD.n7545 VDD.n7544 185
R6335 VDD.n7546 VDD.n7545 185
R6336 VDD.n7523 VDD.n6999 185
R6337 VDD.n7555 VDD.n6999 185
R6338 VDD.n7587 VDD.n7586 185
R6339 VDD.n7588 VDD.n7587 185
R6340 VDD.n7002 VDD.n7000 185
R6341 VDD.n7012 VDD.n7000 185
R6342 VDD.n7004 VDD.n6974 185
R6343 VDD.t316 VDD.n6974 185
R6344 VDD.n7623 VDD.n7622 185
R6345 VDD.n7622 VDD.n7621 185
R6346 VDD.n7624 VDD.n6965 185
R6347 VDD.n7608 VDD.n6965 185
R6348 VDD.n7639 VDD.n7638 185
R6349 VDD.n7640 VDD.n7639 185
R6350 VDD.n7637 VDD.n6966 185
R6351 VDD.n7614 VDD.n6966 185
R6352 VDD.n6968 VDD.n6936 185
R6353 VDD.n6953 VDD.n6936 185
R6354 VDD.n7666 VDD.n7665 185
R6355 VDD.n7667 VDD.n7666 185
R6356 VDD.n6939 VDD.n6937 185
R6357 VDD.n6937 VDD.n6927 185
R6358 VDD.n6941 VDD.n6905 185
R6359 VDD.n7674 VDD.n6905 185
R6360 VDD.n7693 VDD.n7692 185
R6361 VDD.n7694 VDD.n7693 185
R6362 VDD.n6908 VDD.n6906 185
R6363 VDD.n6921 VDD.n6906 185
R6364 VDD.n6910 VDD.n6769 185
R6365 VDD.n7702 VDD.n6769 185
R6366 VDD.n8101 VDD.n8100 185
R6367 VDD.n8102 VDD.n8101 185
R6368 VDD.n6772 VDD.n6770 185
R6369 VDD.n7708 VDD.n6770 185
R6370 VDD.n7726 VDD.n7725 185
R6371 VDD.n7725 VDD.n6779 185
R6372 VDD.n7727 VDD.n6790 185
R6373 VDD.n7716 VDD.n6790 185
R6374 VDD.n8082 VDD.n8081 185
R6375 VDD.n8083 VDD.n8082 185
R6376 VDD.n8080 VDD.n6791 185
R6377 VDD.n7947 VDD.n6791 185
R6378 VDD.n8079 VDD.n8078 185
R6379 VDD.n8078 VDD.n8077 185
R6380 VDD.n6794 VDD.n6793 185
R6381 VDD.n8071 VDD.n6794 185
R6382 VDD.n6832 VDD.n6831 185
R6383 VDD.n6831 VDD.n6807 185
R6384 VDD.n6833 VDD.n6829 185
R6385 VDD.n6829 VDD.n6824 185
R6386 VDD.n8059 VDD.n8058 185
R6387 VDD.n8060 VDD.n8059 185
R6388 VDD.n8057 VDD.n6830 185
R6389 VDD.n7959 VDD.n6830 185
R6390 VDD.n8056 VDD.n8055 185
R6391 VDD.n8055 VDD.n8054 185
R6392 VDD.n6835 VDD.n6834 185
R6393 VDD.n7965 VDD.n6835 185
R6394 VDD.n8047 VDD.n8046 185
R6395 VDD.n8048 VDD.n8047 185
R6396 VDD.n8045 VDD.n6852 185
R6397 VDD.n7999 VDD.n6852 185
R6398 VDD.n8044 VDD.n8043 185
R6399 VDD.n8043 VDD.n8042 185
R6400 VDD.n7209 VDD.n7208 185
R6401 VDD.n7210 VDD.n7209 185
R6402 VDD.n7207 VDD.n7180 185
R6403 VDD.n7206 VDD.n7205 185
R6404 VDD.n7204 VDD.n7203 185
R6405 VDD.n7202 VDD.n7201 185
R6406 VDD.n7200 VDD.n7199 185
R6407 VDD.n7198 VDD.n7197 185
R6408 VDD.n7196 VDD.n7195 185
R6409 VDD.n7194 VDD.n7193 185
R6410 VDD.n7192 VDD.n7191 185
R6411 VDD.n7190 VDD.n7189 185
R6412 VDD.n7188 VDD.n7187 185
R6413 VDD.n7186 VDD.n7185 185
R6414 VDD.n7184 VDD.n7183 185
R6415 VDD.n7182 VDD.n7181 185
R6416 VDD.n7172 VDD.n7171 185
R6417 VDD.n7213 VDD.n7212 185
R6418 VDD.n7214 VDD.n7170 185
R6419 VDD.n7170 VDD.n7169 185
R6420 VDD.n7216 VDD.n7215 185
R6421 VDD.n7217 VDD.n7216 185
R6422 VDD.n7164 VDD.n7163 185
R6423 VDD.n7165 VDD.n7164 185
R6424 VDD.n7225 VDD.n7224 185
R6425 VDD.n7224 VDD.n7223 185
R6426 VDD.n7226 VDD.n7162 185
R6427 VDD.n7162 VDD.n7161 185
R6428 VDD.n7228 VDD.n7227 185
R6429 VDD.n7229 VDD.n7228 185
R6430 VDD.n7156 VDD.n7155 185
R6431 VDD.n7157 VDD.n7156 185
R6432 VDD.n7238 VDD.n7237 185
R6433 VDD.n7237 VDD.n7236 185
R6434 VDD.n7239 VDD.n7154 185
R6435 VDD.n7235 VDD.n7154 185
R6436 VDD.n7241 VDD.n7240 185
R6437 VDD.n7242 VDD.n7241 185
R6438 VDD.n7149 VDD.n7148 185
R6439 VDD.n7153 VDD.n7149 185
R6440 VDD.n7251 VDD.n7250 185
R6441 VDD.n7250 VDD.n7249 185
R6442 VDD.n7252 VDD.n7147 185
R6443 VDD.n7248 VDD.n7147 185
R6444 VDD.n7254 VDD.n7253 185
R6445 VDD.n7255 VDD.n7254 185
R6446 VDD.n7142 VDD.n7141 185
R6447 VDD.n7143 VDD.n7142 185
R6448 VDD.n7263 VDD.n7262 185
R6449 VDD.n7262 VDD.n7261 185
R6450 VDD.n7264 VDD.n7140 185
R6451 VDD.n7140 VDD.n7139 185
R6452 VDD.n7267 VDD.n7266 185
R6453 VDD.n7268 VDD.n7267 185
R6454 VDD.n7265 VDD.n7133 185
R6455 VDD.n7134 VDD.n7133 185
R6456 VDD.n7314 VDD.n7132 185
R6457 VDD.n7314 VDD.n7313 185
R6458 VDD.n7316 VDD.n7315 185
R6459 VDD.n7315 VDD.n7111 185
R6460 VDD.n7317 VDD.n7130 185
R6461 VDD.n7130 VDD.n7120 185
R6462 VDD.n7322 VDD.n7321 185
R6463 VDD.n7323 VDD.n7322 185
R6464 VDD.n7320 VDD.n7131 185
R6465 VDD.n7131 VDD.n7107 185
R6466 VDD.n7318 VDD.n7103 185
R6467 VDD.n7103 VDD.n7090 185
R6468 VDD.n7410 VDD.n7409 185
R6469 VDD.n7409 VDD.n7408 185
R6470 VDD.n7411 VDD.n7097 185
R6471 VDD.n7097 VDD.n7083 185
R6472 VDD.n7425 VDD.n7424 185
R6473 VDD.n7426 VDD.n7425 185
R6474 VDD.n7100 VDD.n7098 185
R6475 VDD.n7098 VDD.n7079 185
R6476 VDD.n7419 VDD.n7418 185
R6477 VDD.n7418 VDD.n7063 185
R6478 VDD.n7416 VDD.n7054 185
R6479 VDD.n7076 VDD.n7054 185
R6480 VDD.n7478 VDD.n7477 185
R6481 VDD.n7477 VDD.n7476 185
R6482 VDD.n7479 VDD.n7048 185
R6483 VDD.n7073 VDD.n7048 185
R6484 VDD.n7493 VDD.n7492 185
R6485 VDD.n7494 VDD.n7493 185
R6486 VDD.n7051 VDD.n7049 185
R6487 VDD.n7049 VDD.n7035 185
R6488 VDD.n7487 VDD.n7486 185
R6489 VDD.n7486 VDD.n7032 185
R6490 VDD.n7484 VDD.n6422 185
R6491 VDD.n6422 VDD.n6409 185
R6492 VDD.n8115 VDD.n8114 185
R6493 VDD.n8116 VDD.n8115 185
R6494 VDD.n8113 VDD.n6423 185
R6495 VDD.n7028 VDD.n6423 185
R6496 VDD.n7018 VDD.n6425 185
R6497 VDD.n7026 VDD.n7018 185
R6498 VDD.n7558 VDD.n7557 185
R6499 VDD.n7557 VDD.n7556 185
R6500 VDD.n7559 VDD.n7013 185
R6501 VDD.n7013 VDD.n6996 185
R6502 VDD.n7573 VDD.n7572 185
R6503 VDD.n7574 VDD.n7573 185
R6504 VDD.n7016 VDD.n7014 185
R6505 VDD.n7014 VDD.n6992 185
R6506 VDD.n7567 VDD.n7566 185
R6507 VDD.n7566 VDD.n6975 185
R6508 VDD.n7564 VDD.n6960 185
R6509 VDD.n6989 VDD.n6960 185
R6510 VDD.n7643 VDD.n7642 185
R6511 VDD.n7642 VDD.n7641 185
R6512 VDD.n7644 VDD.n6954 185
R6513 VDD.n6986 VDD.n6954 185
R6514 VDD.n7654 VDD.n7653 185
R6515 VDD.n7655 VDD.n7654 185
R6516 VDD.n6957 VDD.n6955 185
R6517 VDD.n6955 VDD.n6933 185
R6518 VDD.n7648 VDD.n6926 185
R6519 VDD.n7658 VDD.n6926 185
R6520 VDD.n7677 VDD.n7676 185
R6521 VDD.n7676 VDD.n7675 185
R6522 VDD.n6923 VDD.n6922 185
R6523 VDD.n6922 VDD.n6902 185
R6524 VDD.n7684 VDD.n7683 185
R6525 VDD.n7685 VDD.n7684 185
R6526 VDD.n6763 VDD.n6761 185
R6527 VDD.n6896 VDD.n6763 185
R6528 VDD.n8105 VDD.n8104 185
R6529 VDD.n8104 VDD.n8103 185
R6530 VDD.n6764 VDD.n6762 185
R6531 VDD.n6893 VDD.n6764 185
R6532 VDD.n8092 VDD.n8091 185
R6533 VDD.n8093 VDD.n8092 185
R6534 VDD.n6782 VDD.n6780 185
R6535 VDD.n6889 VDD.n6780 185
R6536 VDD.n8086 VDD.n8085 185
R6537 VDD.n8085 VDD.n8084 185
R6538 VDD.n6813 VDD.n6785 185
R6539 VDD.n7945 VDD.n6785 185
R6540 VDD.n6816 VDD.n6815 185
R6541 VDD.n6815 VDD.n6795 185
R6542 VDD.n6817 VDD.n6808 185
R6543 VDD.n6808 VDD.n6804 185
R6544 VDD.n8069 VDD.n8068 185
R6545 VDD.n8070 VDD.n8069 185
R6546 VDD.n6811 VDD.n6809 185
R6547 VDD.n7737 VDD.n6809 185
R6548 VDD.n8063 VDD.n8062 185
R6549 VDD.n8062 VDD.n8061 185
R6550 VDD.n7758 VDD.n6823 185
R6551 VDD.n6886 VDD.n6823 185
R6552 VDD.n7762 VDD.n7761 185
R6553 VDD.n7762 VDD.n6836 185
R6554 VDD.n7764 VDD.n7763 185
R6555 VDD.n7763 VDD.n6882 185
R6556 VDD.n7755 VDD.n7754 185
R6557 VDD.n7754 VDD.n6849 185
R6558 VDD.n7769 VDD.n7768 185
R6559 VDD.n7769 VDD.n6880 185
R6560 VDD.n7770 VDD.n7753 185
R6561 VDD.n7770 VDD.n6855 185
R6562 VDD.n7772 VDD.n7771 185
R6563 VDD.n7771 VDD.n6858 185
R6564 VDD.n7773 VDD.n7751 185
R6565 VDD.n7751 VDD.n6877 185
R6566 VDD.n7910 VDD.n7909 185
R6567 VDD.n7911 VDD.n7910 185
R6568 VDD.n7908 VDD.n7752 185
R6569 VDD.n7752 VDD.n7750 185
R6570 VDD.n7907 VDD.n7906 185
R6571 VDD.n7906 VDD.n7905 185
R6572 VDD.n7775 VDD.n7774 185
R6573 VDD.n7904 VDD.n7775 185
R6574 VDD.n7902 VDD.n7901 185
R6575 VDD.n7903 VDD.n7902 185
R6576 VDD.n7900 VDD.n7780 185
R6577 VDD.n7780 VDD.n7779 185
R6578 VDD.n7899 VDD.n7898 185
R6579 VDD.n7898 VDD.n7897 185
R6580 VDD.n7782 VDD.n7781 185
R6581 VDD.n7896 VDD.n7782 185
R6582 VDD.n7894 VDD.n7893 185
R6583 VDD.n7895 VDD.n7894 185
R6584 VDD.n7892 VDD.n7786 185
R6585 VDD.n7789 VDD.n7786 185
R6586 VDD.n7891 VDD.n7890 185
R6587 VDD.n7890 VDD.n7889 185
R6588 VDD.n7788 VDD.n7787 185
R6589 VDD.n7888 VDD.n7788 185
R6590 VDD.n7886 VDD.n7885 185
R6591 VDD.n7887 VDD.n7886 185
R6592 VDD.n7884 VDD.n7794 185
R6593 VDD.n7794 VDD.n7793 185
R6594 VDD.n7883 VDD.n7882 185
R6595 VDD.n7882 VDD.n7881 185
R6596 VDD.n7796 VDD.n7795 185
R6597 VDD.n7880 VDD.n7796 185
R6598 VDD.n7878 VDD.n7877 185
R6599 VDD.n7879 VDD.n7878 185
R6600 VDD.n7876 VDD.n7801 185
R6601 VDD.n7801 VDD.n7800 185
R6602 VDD.n7875 VDD.n7874 185
R6603 VDD.n7874 VDD.n7873 185
R6604 VDD.n7803 VDD.n7802 185
R6605 VDD.n7872 VDD.n7803 185
R6606 VDD.n7869 VDD.n7868 185
R6607 VDD.n7867 VDD.n7814 185
R6608 VDD.n7866 VDD.n7813 185
R6609 VDD.n7871 VDD.n7813 185
R6610 VDD.n7865 VDD.n7864 185
R6611 VDD.n7863 VDD.n7862 185
R6612 VDD.n7861 VDD.n7860 185
R6613 VDD.n7859 VDD.n7858 185
R6614 VDD.n7857 VDD.n7856 185
R6615 VDD.n7855 VDD.n7854 185
R6616 VDD.n7853 VDD.n7852 185
R6617 VDD.n7851 VDD.n7850 185
R6618 VDD.n7849 VDD.n7848 185
R6619 VDD.n7847 VDD.n7846 185
R6620 VDD.n7845 VDD.n7844 185
R6621 VDD.n7843 VDD.n7842 185
R6622 VDD.n7841 VDD.n7840 185
R6623 VDD.n7839 VDD.n7838 185
R6624 VDD.n7837 VDD.n7805 185
R6625 VDD.n7872 VDD.n7805 185
R6626 VDD.n7836 VDD.n7804 185
R6627 VDD.n7873 VDD.n7804 185
R6628 VDD.n7835 VDD.n7834 185
R6629 VDD.n7834 VDD.n7800 185
R6630 VDD.n7833 VDD.n7799 185
R6631 VDD.n7879 VDD.n7799 185
R6632 VDD.n7832 VDD.n7798 185
R6633 VDD.n7880 VDD.n7798 185
R6634 VDD.n7831 VDD.n7797 185
R6635 VDD.n7881 VDD.n7797 185
R6636 VDD.n7830 VDD.n7829 185
R6637 VDD.n7829 VDD.n7793 185
R6638 VDD.n7828 VDD.n7792 185
R6639 VDD.n7887 VDD.n7792 185
R6640 VDD.n7827 VDD.n7791 185
R6641 VDD.n7888 VDD.n7791 185
R6642 VDD.n7826 VDD.n7790 185
R6643 VDD.n7889 VDD.n7790 185
R6644 VDD.n7825 VDD.n7824 185
R6645 VDD.n7824 VDD.n7789 185
R6646 VDD.n7823 VDD.n7785 185
R6647 VDD.n7895 VDD.n7785 185
R6648 VDD.n7822 VDD.n7784 185
R6649 VDD.n7896 VDD.n7784 185
R6650 VDD.n7821 VDD.n7783 185
R6651 VDD.n7897 VDD.n7783 185
R6652 VDD.n7820 VDD.n7819 185
R6653 VDD.n7819 VDD.n7779 185
R6654 VDD.n7818 VDD.n7778 185
R6655 VDD.n7903 VDD.n7778 185
R6656 VDD.n7817 VDD.n7777 185
R6657 VDD.n7904 VDD.n7777 185
R6658 VDD.n7816 VDD.n7776 185
R6659 VDD.n7905 VDD.n7776 185
R6660 VDD.n7815 VDD.n7748 185
R6661 VDD.n7750 VDD.n7748 185
R6662 VDD.n7912 VDD.n7749 185
R6663 VDD.n7912 VDD.n7911 185
R6664 VDD.n7913 VDD.n7747 185
R6665 VDD.n7913 VDD.n6877 185
R6666 VDD.n7915 VDD.n7914 185
R6667 VDD.n7914 VDD.n6858 185
R6668 VDD.n7916 VDD.n7746 185
R6669 VDD.n7746 VDD.n6855 185
R6670 VDD.n7918 VDD.n7917 185
R6671 VDD.n7918 VDD.n6880 185
R6672 VDD.n7920 VDD.n7919 185
R6673 VDD.n7919 VDD.n6849 185
R6674 VDD.n7743 VDD.n7742 185
R6675 VDD.n7742 VDD.n6882 185
R6676 VDD.n7926 VDD.n7925 185
R6677 VDD.n7926 VDD.n6836 185
R6678 VDD.n7928 VDD.n7927 185
R6679 VDD.n7927 VDD.n6886 185
R6680 VDD.n7930 VDD.n6825 185
R6681 VDD.n8061 VDD.n6825 185
R6682 VDD.n7739 VDD.n7738 185
R6683 VDD.n7738 VDD.n7737 185
R6684 VDD.n7935 VDD.n6806 185
R6685 VDD.n8070 VDD.n6806 185
R6686 VDD.n7938 VDD.n7937 185
R6687 VDD.n7937 VDD.n6804 185
R6688 VDD.n7722 VDD.n7720 185
R6689 VDD.n7720 VDD.n6795 185
R6690 VDD.n7944 VDD.n7943 185
R6691 VDD.n7945 VDD.n7944 185
R6692 VDD.n7731 VDD.n6786 185
R6693 VDD.n8084 VDD.n6786 185
R6694 VDD.n7730 VDD.n6778 185
R6695 VDD.n6889 VDD.n6778 185
R6696 VDD.n8095 VDD.n8094 185
R6697 VDD.n8094 VDD.n8093 185
R6698 VDD.n6777 VDD.n6775 185
R6699 VDD.n6893 VDD.n6777 185
R6700 VDD.n6916 VDD.n6765 185
R6701 VDD.n8103 VDD.n6765 185
R6702 VDD.n6919 VDD.n6918 185
R6703 VDD.n6919 VDD.n6896 185
R6704 VDD.n7687 VDD.n7686 185
R6705 VDD.n7686 VDD.n7685 185
R6706 VDD.n6915 VDD.n6913 185
R6707 VDD.n6915 VDD.n6902 185
R6708 VDD.n6946 VDD.n6928 185
R6709 VDD.n7675 VDD.n6928 185
R6710 VDD.n7660 VDD.n7659 185
R6711 VDD.n7659 VDD.n7658 185
R6712 VDD.n7657 VDD.n6944 185
R6713 VDD.n7657 VDD.n6933 185
R6714 VDD.n7656 VDD.n6952 185
R6715 VDD.n7656 VDD.n7655 185
R6716 VDD.n7632 VDD.n6950 185
R6717 VDD.n6986 VDD.n6950 185
R6718 VDD.n7630 VDD.n6961 185
R6719 VDD.n7641 VDD.n6961 185
R6720 VDD.n7576 VDD.n6971 185
R6721 VDD.n7576 VDD.n6989 185
R6722 VDD.n7579 VDD.n7578 185
R6723 VDD.n7579 VDD.n6975 185
R6724 VDD.n7581 VDD.n7580 185
R6725 VDD.n7580 VDD.n6992 185
R6726 VDD.n7575 VDD.n7007 185
R6727 VDD.n7575 VDD.n7574 185
R6728 VDD.n7539 VDD.n7011 185
R6729 VDD.n7011 VDD.n6996 185
R6730 VDD.n7537 VDD.n7019 185
R6731 VDD.n7556 VDD.n7019 185
R6732 VDD.n7535 VDD.n7534 185
R6733 VDD.n7534 VDD.n7026 185
R6734 VDD.n6420 VDD.n6418 185
R6735 VDD.n7028 VDD.n6420 185
R6736 VDD.n8118 VDD.n8117 185
R6737 VDD.n8117 VDD.n8116 185
R6738 VDD.n6419 VDD.n6417 185
R6739 VDD.n6419 VDD.n6409 185
R6740 VDD.n7498 VDD.n7497 185
R6741 VDD.n7497 VDD.n7032 185
R6742 VDD.n7496 VDD.n7042 185
R6743 VDD.n7496 VDD.n7035 185
R6744 VDD.n7495 VDD.n7046 185
R6745 VDD.n7495 VDD.n7494 185
R6746 VDD.n7282 VDD.n7044 185
R6747 VDD.n7073 VDD.n7044 185
R6748 VDD.n7279 VDD.n7055 185
R6749 VDD.n7476 VDD.n7055 185
R6750 VDD.n7288 VDD.n7287 185
R6751 VDD.n7288 VDD.n7076 185
R6752 VDD.n7290 VDD.n7289 185
R6753 VDD.n7289 VDD.n7063 185
R6754 VDD.n7278 VDD.n7275 185
R6755 VDD.n7278 VDD.n7079 185
R6756 VDD.n7295 VDD.n7096 185
R6757 VDD.n7426 VDD.n7096 185
R6758 VDD.n7298 VDD.n7297 185
R6759 VDD.n7297 VDD.n7083 185
R6760 VDD.n7273 VDD.n7104 185
R6761 VDD.n7408 VDD.n7104 185
R6762 VDD.n7304 VDD.n7303 185
R6763 VDD.n7304 VDD.n7090 185
R6764 VDD.n7306 VDD.n7305 185
R6765 VDD.n7305 VDD.n7107 185
R6766 VDD.n7307 VDD.n7129 185
R6767 VDD.n7323 VDD.n7129 185
R6768 VDD.n7309 VDD.n7308 185
R6769 VDD.n7308 VDD.n7120 185
R6770 VDD.n7310 VDD.n7136 185
R6771 VDD.n7136 VDD.n7111 185
R6772 VDD.n7312 VDD.n7311 185
R6773 VDD.n7313 VDD.n7312 185
R6774 VDD.n7271 VDD.n7135 185
R6775 VDD.n7135 VDD.n7134 185
R6776 VDD.n7270 VDD.n7269 185
R6777 VDD.n7269 VDD.n7268 185
R6778 VDD.n7138 VDD.n7137 185
R6779 VDD.n7139 VDD.n7138 185
R6780 VDD.n7260 VDD.n7259 185
R6781 VDD.n7261 VDD.n7260 185
R6782 VDD.n7258 VDD.n7144 185
R6783 VDD.n7144 VDD.n7143 185
R6784 VDD.n7257 VDD.n7256 185
R6785 VDD.n7256 VDD.n7255 185
R6786 VDD.n7146 VDD.n7145 185
R6787 VDD.n7248 VDD.n7146 185
R6788 VDD.n7247 VDD.n7246 185
R6789 VDD.n7249 VDD.n7247 185
R6790 VDD.n7245 VDD.n7150 185
R6791 VDD.n7153 VDD.n7150 185
R6792 VDD.n7244 VDD.n7243 185
R6793 VDD.n7243 VDD.n7242 185
R6794 VDD.n7152 VDD.n7151 185
R6795 VDD.n7235 VDD.n7152 185
R6796 VDD.n7234 VDD.n7233 185
R6797 VDD.n7236 VDD.n7234 185
R6798 VDD.n7232 VDD.n7158 185
R6799 VDD.n7158 VDD.n7157 185
R6800 VDD.n7231 VDD.n7230 185
R6801 VDD.n7230 VDD.n7229 185
R6802 VDD.n7160 VDD.n7159 185
R6803 VDD.n7161 VDD.n7160 185
R6804 VDD.n7222 VDD.n7221 185
R6805 VDD.n7223 VDD.n7222 185
R6806 VDD.n7220 VDD.n7166 185
R6807 VDD.n7166 VDD.n7165 185
R6808 VDD.n7219 VDD.n7218 185
R6809 VDD.n7218 VDD.n7217 185
R6810 VDD.n7168 VDD.n7167 185
R6811 VDD.n7169 VDD.n7168 185
R6812 VDD.n5536 VDD 183.946
R6813 VDD.t550 VDD.t118 177.333
R6814 VDD.t475 VDD.t550 177.333
R6815 VDD.t303 VDD.t368 177.333
R6816 VDD.t299 VDD.t303 177.333
R6817 VDD.t301 VDD.t299 177.333
R6818 VDD.t305 VDD.t301 177.333
R6819 VDD.t555 VDD.t287 177.333
R6820 VDD.t287 VDD.t185 177.333
R6821 VDD.t185 VDD.t338 177.333
R6822 VDD.t338 VDD.t244 177.333
R6823 VDD.t320 VDD.t280 177.333
R6824 VDD.t458 VDD.t320 177.333
R6825 VDD.t223 VDD.t290 177.333
R6826 VDD.t290 VDD.t132 177.333
R6827 VDD.t530 VDD.t528 177.333
R6828 VDD.t524 VDD.t530 177.333
R6829 VDD.t526 VDD.t524 177.333
R6830 VDD.t494 VDD.t526 177.333
R6831 VDD.t490 VDD.t494 177.333
R6832 VDD.t492 VDD.t496 177.333
R6833 VDD.t257 VDD.t462 177.333
R6834 VDD.t520 VDD.t257 177.333
R6835 VDD.t681 VDD.t520 177.333
R6836 VDD.t687 VDD.t681 177.333
R6837 VDD.t691 VDD.t687 177.333
R6838 VDD.t695 VDD 174.632
R6839 VDD.n5537 VDD.t583 160.662
R6840 VDD.t132 VDD 158.333
R6841 VDD.n5423 VDD.t70 149.889
R6842 VDD.t238 VDD 149.02
R6843 VDD.t187 VDD 149.02
R6844 VDD.n5232 VDD.n5191 143.53
R6845 VDD.n5243 VDD.n5242 143.53
R6846 VDD.n5224 VDD.n5199 143.53
R6847 VDD.n5218 VDD.n5198 143.53
R6848 VDD.n5290 VDD.n5249 143.53
R6849 VDD.n5294 VDD.n5254 143.53
R6850 VDD.n5281 VDD.n5259 143.53
R6851 VDD.n5287 VDD.n5256 143.53
R6852 VDD.n5220 VDD.n5199 143.469
R6853 VDD.n5277 VDD.n5259 143.469
R6854 VDD.n5424 VDD.t685 141.445
R6855 VDD.t368 VDD.n5360 137.222
R6856 VDD VDD.t305 135.112
R6857 VDD VDD.t458 135.112
R6858 VDD.t496 VDD 135.112
R6859 VDD.t685 VDD 135.112
R6860 VDD.n5361 VDD.t555 133
R6861 VDD.t14 VDD.n5559 132.721
R6862 VDD.n5560 VDD.t577 132.721
R6863 VDD.n5513 VDD.t107 128.065
R6864 VDD.n5236 VDD.n5232 127.859
R6865 VDD.n5300 VDD.n5249 127.859
R6866 VDD.n5225 VDD.t716 117.906
R6867 VDD.t457 VDD.n5193 117.906
R6868 VDD.t59 VDD.n5210 117.906
R6869 VDD.n5212 VDD.t115 117.906
R6870 VDD.t387 VDD.n5283 117.906
R6871 VDD.n5298 VDD.t120 117.906
R6872 VDD.t699 VDD.n5270 117.906
R6873 VDD.n5272 VDD.t481 117.906
R6874 VDD.n5405 VDD.t492 116.112
R6875 VDD.n2606 VDD.t345 115.484
R6876 VDD.n2925 VDD.t533 115.484
R6877 VDD.t74 VDD.n2745 115.484
R6878 VDD.n2750 VDD.t74 115.484
R6879 VDD.n2829 VDD.t76 115.484
R6880 VDD.t76 VDD.n2784 115.484
R6881 VDD.t449 VDD.n3136 115.484
R6882 VDD.n3190 VDD.t403 115.484
R6883 VDD.n3611 VDD.t624 115.484
R6884 VDD.n3471 VDD.t646 115.484
R6885 VDD.n12 VDD.t125 115.484
R6886 VDD.n331 VDD.t124 115.484
R6887 VDD.t252 VDD.n151 115.484
R6888 VDD.n156 VDD.t252 115.484
R6889 VDD.n235 VDD.t122 115.484
R6890 VDD.t122 VDD.n190 115.484
R6891 VDD.t229 VDD.n542 115.484
R6892 VDD.n596 VDD.t308 115.484
R6893 VDD.n1017 VDD.t517 115.484
R6894 VDD.n877 VDD.t80 115.484
R6895 VDD.n5575 VDD.t710 115.484
R6896 VDD.n5894 VDD.t698 115.484
R6897 VDD.t199 VDD.n5714 115.484
R6898 VDD.n5719 VDD.t199 115.484
R6899 VDD.n5798 VDD.t162 115.484
R6900 VDD.t162 VDD.n5753 115.484
R6901 VDD.t153 VDD.n6105 115.484
R6902 VDD.n6159 VDD.t680 115.484
R6903 VDD.n6580 VDD.t180 115.484
R6904 VDD.n6440 VDD.t256 115.484
R6905 VDD.n5382 VDD.t244 107.668
R6906 VDD.n5383 VDD.t708 107.668
R6907 VDD.n5230 VDD.t205 107.025
R6908 VDD.t518 VDD.n5231 107.025
R6909 VDD.t548 VDD.n5253 107.025
R6910 VDD.t487 VDD.n5297 107.025
R6911 VDD.n5242 VDD.n5241 103.013
R6912 VDD.n5289 VDD.n5254 103.013
R6913 VDD.n5486 VDD.t565 100.124
R6914 VDD.n5219 VDD.n5218 96.9887
R6915 VDD.n5276 VDD.n5256 96.9887
R6916 VDD.n5486 VDD.t569 95.4662
R6917 VDD.n4245 VDD.n4244 81.6946
R6918 VDD.n4239 VDD.n4198 81.6946
R6919 VDD.n4899 VDD.n4833 81.6946
R6920 VDD.n4870 VDD.n4868 81.6946
R6921 VDD.n1651 VDD.n1650 81.6946
R6922 VDD.n1645 VDD.n1604 81.6946
R6923 VDD.n2305 VDD.n2239 81.6946
R6924 VDD.n2276 VDD.n2274 81.6946
R6925 VDD.n7214 VDD.n7213 81.6946
R6926 VDD.n7208 VDD.n7167 81.6946
R6927 VDD.n7868 VDD.n7802 81.6946
R6928 VDD.n7839 VDD.n7837 81.6946
R6929 VDD.n4391 VDD.n4136 79.8123
R6930 VDD.n4421 VDD.n4389 79.8123
R6931 VDD.n5075 VDD.n3884 79.8123
R6932 VDD.n5035 VDD.n5033 79.8123
R6933 VDD.n5071 VDD.n5070 79.8123
R6934 VDD.n4384 VDD.n4383 79.8123
R6935 VDD.n4427 VDD.n4426 79.8123
R6936 VDD.n5027 VDD.n5026 79.8123
R6937 VDD.n1797 VDD.n1542 79.8123
R6938 VDD.n1827 VDD.n1795 79.8123
R6939 VDD.n2481 VDD.n1290 79.8123
R6940 VDD.n2441 VDD.n2439 79.8123
R6941 VDD.n2477 VDD.n2476 79.8123
R6942 VDD.n1790 VDD.n1789 79.8123
R6943 VDD.n1833 VDD.n1832 79.8123
R6944 VDD.n2433 VDD.n2432 79.8123
R6945 VDD.n7360 VDD.n7105 79.8123
R6946 VDD.n7390 VDD.n7358 79.8123
R6947 VDD.n8044 VDD.n6853 79.8123
R6948 VDD.n8004 VDD.n8002 79.8123
R6949 VDD.n8040 VDD.n8039 79.8123
R6950 VDD.n7353 VDD.n7352 79.8123
R6951 VDD.n7396 VDD.n7395 79.8123
R6952 VDD.n7996 VDD.n7995 79.8123
R6953 VDD.n2672 VDD.n2646 79.4358
R6954 VDD.n3014 VDD.n3013 79.4358
R6955 VDD.n3086 VDD.n3085 79.4358
R6956 VDD.n2977 VDD.n2976 79.4358
R6957 VDD.n2802 VDD.n2638 79.4358
R6958 VDD.n3018 VDD.n2729 79.4358
R6959 VDD.n2887 VDD.n2884 79.4358
R6960 VDD.n2850 VDD.n2778 79.4358
R6961 VDD.n78 VDD.n52 79.4358
R6962 VDD.n420 VDD.n419 79.4358
R6963 VDD.n492 VDD.n491 79.4358
R6964 VDD.n383 VDD.n382 79.4358
R6965 VDD.n208 VDD.n44 79.4358
R6966 VDD.n424 VDD.n135 79.4358
R6967 VDD.n293 VDD.n290 79.4358
R6968 VDD.n256 VDD.n184 79.4358
R6969 VDD.n5641 VDD.n5615 79.4358
R6970 VDD.n5983 VDD.n5982 79.4358
R6971 VDD.n6055 VDD.n6054 79.4358
R6972 VDD.n5946 VDD.n5945 79.4358
R6973 VDD.n5771 VDD.n5607 79.4358
R6974 VDD.n5987 VDD.n5698 79.4358
R6975 VDD.n5856 VDD.n5853 79.4358
R6976 VDD.n5819 VDD.n5747 79.4358
R6977 VDD.n5214 VDD.n5201 79.2266
R6978 VDD.n5274 VDD.n5261 79.2266
R6979 VDD.n5208 VDD.n5201 78.4737
R6980 VDD.n5268 VDD.n5261 78.4737
R6981 VDD.n2668 VDD.n2667 72.7879
R6982 VDD.n2663 VDD.n2650 72.7879
R6983 VDD.n2661 VDD.n2660 72.7879
R6984 VDD.n2655 VDD.n2653 72.7879
R6985 VDD.n3097 VDD.n2624 72.7879
R6986 VDD.n3095 VDD.n3094 72.7879
R6987 VDD.n3090 VDD.n2628 72.7879
R6988 VDD.n3088 VDD.n3087 72.7879
R6989 VDD.n3010 VDD.n2734 72.7879
R6990 VDD.n3009 VDD.n3008 72.7879
R6991 VDD.n3002 VDD.n2736 72.7879
R6992 VDD.n3001 VDD.n3000 72.7879
R6993 VDD.n2991 VDD.n2738 72.7879
R6994 VDD.n2990 VDD.n2943 72.7879
R6995 VDD.n2986 VDD.n2985 72.7879
R6996 VDD.n2979 VDD.n2945 72.7879
R6997 VDD.n3011 VDD.n3010 72.7879
R6998 VDD.n3008 VDD.n3007 72.7879
R6999 VDD.n3003 VDD.n3002 72.7879
R7000 VDD.n3000 VDD.n2999 72.7879
R7001 VDD.n2992 VDD.n2991 72.7879
R7002 VDD.n2987 VDD.n2943 72.7879
R7003 VDD.n2985 VDD.n2984 72.7879
R7004 VDD.n2980 VDD.n2979 72.7879
R7005 VDD.n3089 VDD.n3088 72.7879
R7006 VDD.n2628 VDD.n2626 72.7879
R7007 VDD.n3096 VDD.n3095 72.7879
R7008 VDD.n2654 VDD.n2624 72.7879
R7009 VDD.n2653 VDD.n2651 72.7879
R7010 VDD.n2662 VDD.n2661 72.7879
R7011 VDD.n2650 VDD.n2648 72.7879
R7012 VDD.n2669 VDD.n2668 72.7879
R7013 VDD.n2759 VDD.n2730 72.7879
R7014 VDD.n2765 VDD.n2764 72.7879
R7015 VDD.n2768 VDD.n2767 72.7879
R7016 VDD.n2773 VDD.n2772 72.7879
R7017 VDD.n2900 VDD.n2899 72.7879
R7018 VDD.n2893 VDD.n2775 72.7879
R7019 VDD.n2892 VDD.n2891 72.7879
R7020 VDD.n2885 VDD.n2777 72.7879
R7021 VDD.n2804 VDD.n2803 72.7879
R7022 VDD.n2807 VDD.n2806 72.7879
R7023 VDD.n2812 VDD.n2811 72.7879
R7024 VDD.n2820 VDD.n2815 72.7879
R7025 VDD.n2819 VDD.n2818 72.7879
R7026 VDD.n2839 VDD.n2838 72.7879
R7027 VDD.n2842 VDD.n2841 72.7879
R7028 VDD.n2847 VDD.n2846 72.7879
R7029 VDD.n2813 VDD.n2812 72.7879
R7030 VDD.n2806 VDD.n2800 72.7879
R7031 VDD.n2805 VDD.n2804 72.7879
R7032 VDD.n2760 VDD.n2759 72.7879
R7033 VDD.n2766 VDD.n2765 72.7879
R7034 VDD.n2767 VDD.n2756 72.7879
R7035 VDD.n2774 VDD.n2773 72.7879
R7036 VDD.n2899 VDD.n2898 72.7879
R7037 VDD.n2894 VDD.n2893 72.7879
R7038 VDD.n2891 VDD.n2890 72.7879
R7039 VDD.n2886 VDD.n2885 72.7879
R7040 VDD.n2848 VDD.n2847 72.7879
R7041 VDD.n2841 VDD.n2779 72.7879
R7042 VDD.n2840 VDD.n2839 72.7879
R7043 VDD.n2818 VDD.n2781 72.7879
R7044 VDD.n2821 VDD.n2820 72.7879
R7045 VDD.n4418 VDD.n4159 72.7879
R7046 VDD.n4414 VDD.n4158 72.7879
R7047 VDD.n4410 VDD.n4157 72.7879
R7048 VDD.n4406 VDD.n4156 72.7879
R7049 VDD.n4402 VDD.n4155 72.7879
R7050 VDD.n4398 VDD.n4154 72.7879
R7051 VDD.n4394 VDD.n4153 72.7879
R7052 VDD.n4390 VDD.n4152 72.7879
R7053 VDD.n5065 VDD.n3885 72.7879
R7054 VDD.n5060 VDD.n3893 72.7879
R7055 VDD.n5057 VDD.n3894 72.7879
R7056 VDD.n5053 VDD.n3895 72.7879
R7057 VDD.n5049 VDD.n3896 72.7879
R7058 VDD.n5045 VDD.n3897 72.7879
R7059 VDD.n5041 VDD.n3898 72.7879
R7060 VDD.n5037 VDD.n3899 72.7879
R7061 VDD.n4379 VDD.n4144 72.7879
R7062 VDD.n4375 VDD.n4145 72.7879
R7063 VDD.n4371 VDD.n4146 72.7879
R7064 VDD.n4367 VDD.n4147 72.7879
R7065 VDD.n4363 VDD.n4148 72.7879
R7066 VDD.n4359 VDD.n4149 72.7879
R7067 VDD.n4355 VDD.n4150 72.7879
R7068 VDD.n4425 VDD.n4424 72.7879
R7069 VDD.n5067 VDD.n3890 72.7879
R7070 VDD.n3900 VDD.n3892 72.7879
R7071 VDD.n5002 VDD.n3901 72.7879
R7072 VDD.n5006 VDD.n3902 72.7879
R7073 VDD.n5010 VDD.n3903 72.7879
R7074 VDD.n5014 VDD.n3904 72.7879
R7075 VDD.n5018 VDD.n3905 72.7879
R7076 VDD.n5022 VDD.n3906 72.7879
R7077 VDD.n5068 VDD.n5067 72.7879
R7078 VDD.n5001 VDD.n3900 72.7879
R7079 VDD.n5005 VDD.n3901 72.7879
R7080 VDD.n5009 VDD.n3902 72.7879
R7081 VDD.n5013 VDD.n3903 72.7879
R7082 VDD.n5017 VDD.n3904 72.7879
R7083 VDD.n5021 VDD.n3905 72.7879
R7084 VDD.n5024 VDD.n3906 72.7879
R7085 VDD.n4424 VDD.n4141 72.7879
R7086 VDD.n4358 VDD.n4150 72.7879
R7087 VDD.n4362 VDD.n4149 72.7879
R7088 VDD.n4366 VDD.n4148 72.7879
R7089 VDD.n4370 VDD.n4147 72.7879
R7090 VDD.n4374 VDD.n4146 72.7879
R7091 VDD.n4378 VDD.n4145 72.7879
R7092 VDD.n4381 VDD.n4144 72.7879
R7093 VDD.n5065 VDD.n5064 72.7879
R7094 VDD.n5058 VDD.n3893 72.7879
R7095 VDD.n5054 VDD.n3894 72.7879
R7096 VDD.n5050 VDD.n3895 72.7879
R7097 VDD.n5046 VDD.n3896 72.7879
R7098 VDD.n5042 VDD.n3897 72.7879
R7099 VDD.n5038 VDD.n3898 72.7879
R7100 VDD.n5034 VDD.n3899 72.7879
R7101 VDD.n4393 VDD.n4152 72.7879
R7102 VDD.n4397 VDD.n4153 72.7879
R7103 VDD.n4401 VDD.n4154 72.7879
R7104 VDD.n4405 VDD.n4155 72.7879
R7105 VDD.n4409 VDD.n4156 72.7879
R7106 VDD.n4413 VDD.n4157 72.7879
R7107 VDD.n4417 VDD.n4158 72.7879
R7108 VDD.n4388 VDD.n4159 72.7879
R7109 VDD.n4901 VDD.n4900 72.7879
R7110 VDD.n4895 VDD.n4837 72.7879
R7111 VDD.n4892 VDD.n4838 72.7879
R7112 VDD.n4888 VDD.n4839 72.7879
R7113 VDD.n4884 VDD.n4840 72.7879
R7114 VDD.n4880 VDD.n4841 72.7879
R7115 VDD.n4876 VDD.n4842 72.7879
R7116 VDD.n4872 VDD.n4843 72.7879
R7117 VDD.n4243 VDD.n4242 72.7879
R7118 VDD.n4212 VDD.n4204 72.7879
R7119 VDD.n4216 VDD.n4205 72.7879
R7120 VDD.n4220 VDD.n4206 72.7879
R7121 VDD.n4224 VDD.n4207 72.7879
R7122 VDD.n4228 VDD.n4208 72.7879
R7123 VDD.n4232 VDD.n4209 72.7879
R7124 VDD.n4236 VDD.n4210 72.7879
R7125 VDD.n4211 VDD.n4210 72.7879
R7126 VDD.n4235 VDD.n4209 72.7879
R7127 VDD.n4231 VDD.n4208 72.7879
R7128 VDD.n4227 VDD.n4207 72.7879
R7129 VDD.n4223 VDD.n4206 72.7879
R7130 VDD.n4219 VDD.n4205 72.7879
R7131 VDD.n4215 VDD.n4204 72.7879
R7132 VDD.n4242 VDD.n4203 72.7879
R7133 VDD.n4901 VDD.n4845 72.7879
R7134 VDD.n4893 VDD.n4837 72.7879
R7135 VDD.n4889 VDD.n4838 72.7879
R7136 VDD.n4885 VDD.n4839 72.7879
R7137 VDD.n4881 VDD.n4840 72.7879
R7138 VDD.n4877 VDD.n4841 72.7879
R7139 VDD.n4873 VDD.n4842 72.7879
R7140 VDD.n4869 VDD.n4843 72.7879
R7141 VDD.n74 VDD.n73 72.7879
R7142 VDD.n69 VDD.n56 72.7879
R7143 VDD.n67 VDD.n66 72.7879
R7144 VDD.n61 VDD.n59 72.7879
R7145 VDD.n503 VDD.n30 72.7879
R7146 VDD.n501 VDD.n500 72.7879
R7147 VDD.n496 VDD.n34 72.7879
R7148 VDD.n494 VDD.n493 72.7879
R7149 VDD.n416 VDD.n140 72.7879
R7150 VDD.n415 VDD.n414 72.7879
R7151 VDD.n408 VDD.n142 72.7879
R7152 VDD.n407 VDD.n406 72.7879
R7153 VDD.n397 VDD.n144 72.7879
R7154 VDD.n396 VDD.n349 72.7879
R7155 VDD.n392 VDD.n391 72.7879
R7156 VDD.n385 VDD.n351 72.7879
R7157 VDD.n417 VDD.n416 72.7879
R7158 VDD.n414 VDD.n413 72.7879
R7159 VDD.n409 VDD.n408 72.7879
R7160 VDD.n406 VDD.n405 72.7879
R7161 VDD.n398 VDD.n397 72.7879
R7162 VDD.n393 VDD.n349 72.7879
R7163 VDD.n391 VDD.n390 72.7879
R7164 VDD.n386 VDD.n385 72.7879
R7165 VDD.n495 VDD.n494 72.7879
R7166 VDD.n34 VDD.n32 72.7879
R7167 VDD.n502 VDD.n501 72.7879
R7168 VDD.n60 VDD.n30 72.7879
R7169 VDD.n59 VDD.n57 72.7879
R7170 VDD.n68 VDD.n67 72.7879
R7171 VDD.n56 VDD.n54 72.7879
R7172 VDD.n75 VDD.n74 72.7879
R7173 VDD.n165 VDD.n136 72.7879
R7174 VDD.n171 VDD.n170 72.7879
R7175 VDD.n174 VDD.n173 72.7879
R7176 VDD.n179 VDD.n178 72.7879
R7177 VDD.n306 VDD.n305 72.7879
R7178 VDD.n299 VDD.n181 72.7879
R7179 VDD.n298 VDD.n297 72.7879
R7180 VDD.n291 VDD.n183 72.7879
R7181 VDD.n210 VDD.n209 72.7879
R7182 VDD.n213 VDD.n212 72.7879
R7183 VDD.n218 VDD.n217 72.7879
R7184 VDD.n226 VDD.n221 72.7879
R7185 VDD.n225 VDD.n224 72.7879
R7186 VDD.n245 VDD.n244 72.7879
R7187 VDD.n248 VDD.n247 72.7879
R7188 VDD.n253 VDD.n252 72.7879
R7189 VDD.n219 VDD.n218 72.7879
R7190 VDD.n212 VDD.n206 72.7879
R7191 VDD.n211 VDD.n210 72.7879
R7192 VDD.n166 VDD.n165 72.7879
R7193 VDD.n172 VDD.n171 72.7879
R7194 VDD.n173 VDD.n162 72.7879
R7195 VDD.n180 VDD.n179 72.7879
R7196 VDD.n305 VDD.n304 72.7879
R7197 VDD.n300 VDD.n299 72.7879
R7198 VDD.n297 VDD.n296 72.7879
R7199 VDD.n292 VDD.n291 72.7879
R7200 VDD.n254 VDD.n253 72.7879
R7201 VDD.n247 VDD.n185 72.7879
R7202 VDD.n246 VDD.n245 72.7879
R7203 VDD.n224 VDD.n187 72.7879
R7204 VDD.n227 VDD.n226 72.7879
R7205 VDD.n1824 VDD.n1565 72.7879
R7206 VDD.n1820 VDD.n1564 72.7879
R7207 VDD.n1816 VDD.n1563 72.7879
R7208 VDD.n1812 VDD.n1562 72.7879
R7209 VDD.n1808 VDD.n1561 72.7879
R7210 VDD.n1804 VDD.n1560 72.7879
R7211 VDD.n1800 VDD.n1559 72.7879
R7212 VDD.n1796 VDD.n1558 72.7879
R7213 VDD.n2471 VDD.n1291 72.7879
R7214 VDD.n2466 VDD.n1299 72.7879
R7215 VDD.n2463 VDD.n1300 72.7879
R7216 VDD.n2459 VDD.n1301 72.7879
R7217 VDD.n2455 VDD.n1302 72.7879
R7218 VDD.n2451 VDD.n1303 72.7879
R7219 VDD.n2447 VDD.n1304 72.7879
R7220 VDD.n2443 VDD.n1305 72.7879
R7221 VDD.n1785 VDD.n1550 72.7879
R7222 VDD.n1781 VDD.n1551 72.7879
R7223 VDD.n1777 VDD.n1552 72.7879
R7224 VDD.n1773 VDD.n1553 72.7879
R7225 VDD.n1769 VDD.n1554 72.7879
R7226 VDD.n1765 VDD.n1555 72.7879
R7227 VDD.n1761 VDD.n1556 72.7879
R7228 VDD.n1831 VDD.n1830 72.7879
R7229 VDD.n2473 VDD.n1296 72.7879
R7230 VDD.n1306 VDD.n1298 72.7879
R7231 VDD.n2408 VDD.n1307 72.7879
R7232 VDD.n2412 VDD.n1308 72.7879
R7233 VDD.n2416 VDD.n1309 72.7879
R7234 VDD.n2420 VDD.n1310 72.7879
R7235 VDD.n2424 VDD.n1311 72.7879
R7236 VDD.n2428 VDD.n1312 72.7879
R7237 VDD.n2474 VDD.n2473 72.7879
R7238 VDD.n2407 VDD.n1306 72.7879
R7239 VDD.n2411 VDD.n1307 72.7879
R7240 VDD.n2415 VDD.n1308 72.7879
R7241 VDD.n2419 VDD.n1309 72.7879
R7242 VDD.n2423 VDD.n1310 72.7879
R7243 VDD.n2427 VDD.n1311 72.7879
R7244 VDD.n2430 VDD.n1312 72.7879
R7245 VDD.n1830 VDD.n1547 72.7879
R7246 VDD.n1764 VDD.n1556 72.7879
R7247 VDD.n1768 VDD.n1555 72.7879
R7248 VDD.n1772 VDD.n1554 72.7879
R7249 VDD.n1776 VDD.n1553 72.7879
R7250 VDD.n1780 VDD.n1552 72.7879
R7251 VDD.n1784 VDD.n1551 72.7879
R7252 VDD.n1787 VDD.n1550 72.7879
R7253 VDD.n2471 VDD.n2470 72.7879
R7254 VDD.n2464 VDD.n1299 72.7879
R7255 VDD.n2460 VDD.n1300 72.7879
R7256 VDD.n2456 VDD.n1301 72.7879
R7257 VDD.n2452 VDD.n1302 72.7879
R7258 VDD.n2448 VDD.n1303 72.7879
R7259 VDD.n2444 VDD.n1304 72.7879
R7260 VDD.n2440 VDD.n1305 72.7879
R7261 VDD.n1799 VDD.n1558 72.7879
R7262 VDD.n1803 VDD.n1559 72.7879
R7263 VDD.n1807 VDD.n1560 72.7879
R7264 VDD.n1811 VDD.n1561 72.7879
R7265 VDD.n1815 VDD.n1562 72.7879
R7266 VDD.n1819 VDD.n1563 72.7879
R7267 VDD.n1823 VDD.n1564 72.7879
R7268 VDD.n1794 VDD.n1565 72.7879
R7269 VDD.n2307 VDD.n2306 72.7879
R7270 VDD.n2301 VDD.n2243 72.7879
R7271 VDD.n2298 VDD.n2244 72.7879
R7272 VDD.n2294 VDD.n2245 72.7879
R7273 VDD.n2290 VDD.n2246 72.7879
R7274 VDD.n2286 VDD.n2247 72.7879
R7275 VDD.n2282 VDD.n2248 72.7879
R7276 VDD.n2278 VDD.n2249 72.7879
R7277 VDD.n1649 VDD.n1648 72.7879
R7278 VDD.n1618 VDD.n1610 72.7879
R7279 VDD.n1622 VDD.n1611 72.7879
R7280 VDD.n1626 VDD.n1612 72.7879
R7281 VDD.n1630 VDD.n1613 72.7879
R7282 VDD.n1634 VDD.n1614 72.7879
R7283 VDD.n1638 VDD.n1615 72.7879
R7284 VDD.n1642 VDD.n1616 72.7879
R7285 VDD.n1617 VDD.n1616 72.7879
R7286 VDD.n1641 VDD.n1615 72.7879
R7287 VDD.n1637 VDD.n1614 72.7879
R7288 VDD.n1633 VDD.n1613 72.7879
R7289 VDD.n1629 VDD.n1612 72.7879
R7290 VDD.n1625 VDD.n1611 72.7879
R7291 VDD.n1621 VDD.n1610 72.7879
R7292 VDD.n1648 VDD.n1609 72.7879
R7293 VDD.n2307 VDD.n2251 72.7879
R7294 VDD.n2299 VDD.n2243 72.7879
R7295 VDD.n2295 VDD.n2244 72.7879
R7296 VDD.n2291 VDD.n2245 72.7879
R7297 VDD.n2287 VDD.n2246 72.7879
R7298 VDD.n2283 VDD.n2247 72.7879
R7299 VDD.n2279 VDD.n2248 72.7879
R7300 VDD.n2275 VDD.n2249 72.7879
R7301 VDD.n5637 VDD.n5636 72.7879
R7302 VDD.n5632 VDD.n5619 72.7879
R7303 VDD.n5630 VDD.n5629 72.7879
R7304 VDD.n5624 VDD.n5622 72.7879
R7305 VDD.n6066 VDD.n5593 72.7879
R7306 VDD.n6064 VDD.n6063 72.7879
R7307 VDD.n6059 VDD.n5597 72.7879
R7308 VDD.n6057 VDD.n6056 72.7879
R7309 VDD.n5979 VDD.n5703 72.7879
R7310 VDD.n5978 VDD.n5977 72.7879
R7311 VDD.n5971 VDD.n5705 72.7879
R7312 VDD.n5970 VDD.n5969 72.7879
R7313 VDD.n5960 VDD.n5707 72.7879
R7314 VDD.n5959 VDD.n5912 72.7879
R7315 VDD.n5955 VDD.n5954 72.7879
R7316 VDD.n5948 VDD.n5914 72.7879
R7317 VDD.n5980 VDD.n5979 72.7879
R7318 VDD.n5977 VDD.n5976 72.7879
R7319 VDD.n5972 VDD.n5971 72.7879
R7320 VDD.n5969 VDD.n5968 72.7879
R7321 VDD.n5961 VDD.n5960 72.7879
R7322 VDD.n5956 VDD.n5912 72.7879
R7323 VDD.n5954 VDD.n5953 72.7879
R7324 VDD.n5949 VDD.n5948 72.7879
R7325 VDD.n6058 VDD.n6057 72.7879
R7326 VDD.n5597 VDD.n5595 72.7879
R7327 VDD.n6065 VDD.n6064 72.7879
R7328 VDD.n5623 VDD.n5593 72.7879
R7329 VDD.n5622 VDD.n5620 72.7879
R7330 VDD.n5631 VDD.n5630 72.7879
R7331 VDD.n5619 VDD.n5617 72.7879
R7332 VDD.n5638 VDD.n5637 72.7879
R7333 VDD.n5728 VDD.n5699 72.7879
R7334 VDD.n5734 VDD.n5733 72.7879
R7335 VDD.n5737 VDD.n5736 72.7879
R7336 VDD.n5742 VDD.n5741 72.7879
R7337 VDD.n5869 VDD.n5868 72.7879
R7338 VDD.n5862 VDD.n5744 72.7879
R7339 VDD.n5861 VDD.n5860 72.7879
R7340 VDD.n5854 VDD.n5746 72.7879
R7341 VDD.n5773 VDD.n5772 72.7879
R7342 VDD.n5776 VDD.n5775 72.7879
R7343 VDD.n5781 VDD.n5780 72.7879
R7344 VDD.n5789 VDD.n5784 72.7879
R7345 VDD.n5788 VDD.n5787 72.7879
R7346 VDD.n5808 VDD.n5807 72.7879
R7347 VDD.n5811 VDD.n5810 72.7879
R7348 VDD.n5816 VDD.n5815 72.7879
R7349 VDD.n5782 VDD.n5781 72.7879
R7350 VDD.n5775 VDD.n5769 72.7879
R7351 VDD.n5774 VDD.n5773 72.7879
R7352 VDD.n5729 VDD.n5728 72.7879
R7353 VDD.n5735 VDD.n5734 72.7879
R7354 VDD.n5736 VDD.n5725 72.7879
R7355 VDD.n5743 VDD.n5742 72.7879
R7356 VDD.n5868 VDD.n5867 72.7879
R7357 VDD.n5863 VDD.n5862 72.7879
R7358 VDD.n5860 VDD.n5859 72.7879
R7359 VDD.n5855 VDD.n5854 72.7879
R7360 VDD.n5817 VDD.n5816 72.7879
R7361 VDD.n5810 VDD.n5748 72.7879
R7362 VDD.n5809 VDD.n5808 72.7879
R7363 VDD.n5787 VDD.n5750 72.7879
R7364 VDD.n5790 VDD.n5789 72.7879
R7365 VDD.n7387 VDD.n7128 72.7879
R7366 VDD.n7383 VDD.n7127 72.7879
R7367 VDD.n7379 VDD.n7126 72.7879
R7368 VDD.n7375 VDD.n7125 72.7879
R7369 VDD.n7371 VDD.n7124 72.7879
R7370 VDD.n7367 VDD.n7123 72.7879
R7371 VDD.n7363 VDD.n7122 72.7879
R7372 VDD.n7359 VDD.n7121 72.7879
R7373 VDD.n8034 VDD.n6854 72.7879
R7374 VDD.n8029 VDD.n6862 72.7879
R7375 VDD.n8026 VDD.n6863 72.7879
R7376 VDD.n8022 VDD.n6864 72.7879
R7377 VDD.n8018 VDD.n6865 72.7879
R7378 VDD.n8014 VDD.n6866 72.7879
R7379 VDD.n8010 VDD.n6867 72.7879
R7380 VDD.n8006 VDD.n6868 72.7879
R7381 VDD.n7348 VDD.n7113 72.7879
R7382 VDD.n7344 VDD.n7114 72.7879
R7383 VDD.n7340 VDD.n7115 72.7879
R7384 VDD.n7336 VDD.n7116 72.7879
R7385 VDD.n7332 VDD.n7117 72.7879
R7386 VDD.n7328 VDD.n7118 72.7879
R7387 VDD.n7324 VDD.n7119 72.7879
R7388 VDD.n7394 VDD.n7393 72.7879
R7389 VDD.n8036 VDD.n6859 72.7879
R7390 VDD.n6869 VDD.n6861 72.7879
R7391 VDD.n7971 VDD.n6870 72.7879
R7392 VDD.n7975 VDD.n6871 72.7879
R7393 VDD.n7979 VDD.n6872 72.7879
R7394 VDD.n7983 VDD.n6873 72.7879
R7395 VDD.n7987 VDD.n6874 72.7879
R7396 VDD.n7991 VDD.n6875 72.7879
R7397 VDD.n8037 VDD.n8036 72.7879
R7398 VDD.n7970 VDD.n6869 72.7879
R7399 VDD.n7974 VDD.n6870 72.7879
R7400 VDD.n7978 VDD.n6871 72.7879
R7401 VDD.n7982 VDD.n6872 72.7879
R7402 VDD.n7986 VDD.n6873 72.7879
R7403 VDD.n7990 VDD.n6874 72.7879
R7404 VDD.n7993 VDD.n6875 72.7879
R7405 VDD.n7393 VDD.n7110 72.7879
R7406 VDD.n7327 VDD.n7119 72.7879
R7407 VDD.n7331 VDD.n7118 72.7879
R7408 VDD.n7335 VDD.n7117 72.7879
R7409 VDD.n7339 VDD.n7116 72.7879
R7410 VDD.n7343 VDD.n7115 72.7879
R7411 VDD.n7347 VDD.n7114 72.7879
R7412 VDD.n7350 VDD.n7113 72.7879
R7413 VDD.n8034 VDD.n8033 72.7879
R7414 VDD.n8027 VDD.n6862 72.7879
R7415 VDD.n8023 VDD.n6863 72.7879
R7416 VDD.n8019 VDD.n6864 72.7879
R7417 VDD.n8015 VDD.n6865 72.7879
R7418 VDD.n8011 VDD.n6866 72.7879
R7419 VDD.n8007 VDD.n6867 72.7879
R7420 VDD.n8003 VDD.n6868 72.7879
R7421 VDD.n7362 VDD.n7121 72.7879
R7422 VDD.n7366 VDD.n7122 72.7879
R7423 VDD.n7370 VDD.n7123 72.7879
R7424 VDD.n7374 VDD.n7124 72.7879
R7425 VDD.n7378 VDD.n7125 72.7879
R7426 VDD.n7382 VDD.n7126 72.7879
R7427 VDD.n7386 VDD.n7127 72.7879
R7428 VDD.n7357 VDD.n7128 72.7879
R7429 VDD.n7870 VDD.n7869 72.7879
R7430 VDD.n7864 VDD.n7806 72.7879
R7431 VDD.n7861 VDD.n7807 72.7879
R7432 VDD.n7857 VDD.n7808 72.7879
R7433 VDD.n7853 VDD.n7809 72.7879
R7434 VDD.n7849 VDD.n7810 72.7879
R7435 VDD.n7845 VDD.n7811 72.7879
R7436 VDD.n7841 VDD.n7812 72.7879
R7437 VDD.n7212 VDD.n7211 72.7879
R7438 VDD.n7181 VDD.n7173 72.7879
R7439 VDD.n7185 VDD.n7174 72.7879
R7440 VDD.n7189 VDD.n7175 72.7879
R7441 VDD.n7193 VDD.n7176 72.7879
R7442 VDD.n7197 VDD.n7177 72.7879
R7443 VDD.n7201 VDD.n7178 72.7879
R7444 VDD.n7205 VDD.n7179 72.7879
R7445 VDD.n7180 VDD.n7179 72.7879
R7446 VDD.n7204 VDD.n7178 72.7879
R7447 VDD.n7200 VDD.n7177 72.7879
R7448 VDD.n7196 VDD.n7176 72.7879
R7449 VDD.n7192 VDD.n7175 72.7879
R7450 VDD.n7188 VDD.n7174 72.7879
R7451 VDD.n7184 VDD.n7173 72.7879
R7452 VDD.n7211 VDD.n7172 72.7879
R7453 VDD.n7870 VDD.n7814 72.7879
R7454 VDD.n7862 VDD.n7806 72.7879
R7455 VDD.n7858 VDD.n7807 72.7879
R7456 VDD.n7854 VDD.n7808 72.7879
R7457 VDD.n7850 VDD.n7809 72.7879
R7458 VDD.n7846 VDD.n7810 72.7879
R7459 VDD.n7842 VDD.n7811 72.7879
R7460 VDD.n7838 VDD.n7812 72.7879
R7461 VDD.t352 VDD 69.8534
R7462 VDD VDD.t310 69.8534
R7463 VDD.t280 VDD.n5382 69.6672
R7464 VDD.n5383 VDD.t223 69.6672
R7465 VDD.n5513 VDD.t671 67.525
R7466 VDD.n5231 VDD.n5230 64.7432
R7467 VDD.n5297 VDD.n5253 64.7432
R7468 VDD.t716 VDD.t719 63.4219
R7469 VDD.t719 VDD.t720 63.4219
R7470 VDD.t720 VDD.t365 63.4219
R7471 VDD.t365 VDD.t721 63.4219
R7472 VDD.t721 VDD.t366 63.4219
R7473 VDD.t366 VDD.t42 63.4219
R7474 VDD.t42 VDD.t307 63.4219
R7475 VDD.t307 VDD.t474 63.4219
R7476 VDD.t474 VDD.t380 63.4219
R7477 VDD.t380 VDD.t56 63.4219
R7478 VDD.t56 VDD.t367 63.4219
R7479 VDD.t367 VDD.t480 63.4219
R7480 VDD.t480 VDD.t54 63.4219
R7481 VDD.t54 VDD.t477 63.4219
R7482 VDD.t477 VDD.t55 63.4219
R7483 VDD.t55 VDD.t478 63.4219
R7484 VDD.t478 VDD.t379 63.4219
R7485 VDD.t379 VDD.t205 63.4219
R7486 VDD.t514 VDD.t518 63.4219
R7487 VDD.t451 VDD.t514 63.4219
R7488 VDD.t522 VDD.t451 63.4219
R7489 VDD.t72 VDD.t522 63.4219
R7490 VDD.t472 VDD.t72 63.4219
R7491 VDD.t289 VDD.t472 63.4219
R7492 VDD.t171 VDD.t289 63.4219
R7493 VDD.t192 VDD.t171 63.4219
R7494 VDD.t26 VDD.t192 63.4219
R7495 VDD.t26 VDD.t137 63.4219
R7496 VDD.t137 VDD.t136 63.4219
R7497 VDD.t136 VDD.t707 63.4219
R7498 VDD.t707 VDD.t515 63.4219
R7499 VDD.t515 VDD.t140 63.4219
R7500 VDD.t140 VDD.t386 63.4219
R7501 VDD.t386 VDD.t456 63.4219
R7502 VDD.t456 VDD.t294 63.4219
R7503 VDD.t294 VDD.t457 63.4219
R7504 VDD.t484 VDD.t59 63.4219
R7505 VDD.t115 VDD.t713 63.4219
R7506 VDD.t383 VDD.t387 63.4219
R7507 VDD.t328 VDD.t383 63.4219
R7508 VDD.t722 VDD.t328 63.4219
R7509 VDD.t711 VDD.t722 63.4219
R7510 VDD.t697 VDD.t711 63.4219
R7511 VDD.t270 VDD.t697 63.4219
R7512 VDD.t545 VDD.t270 63.4219
R7513 VDD.t209 VDD.t545 63.4219
R7514 VDD.t355 VDD.t209 63.4219
R7515 VDD.t355 VDD.t191 63.4219
R7516 VDD.t191 VDD.t312 63.4219
R7517 VDD.t312 VDD.t532 63.4219
R7518 VDD.t532 VDD.t467 63.4219
R7519 VDD.t467 VDD.t354 63.4219
R7520 VDD.t354 VDD.t33 63.4219
R7521 VDD.t33 VDD.t372 63.4219
R7522 VDD.t372 VDD.t500 63.4219
R7523 VDD.t500 VDD.t548 63.4219
R7524 VDD.t486 VDD.t487 63.4219
R7525 VDD.t204 VDD.t486 63.4219
R7526 VDD.t712 VDD.t204 63.4219
R7527 VDD.t206 VDD.t712 63.4219
R7528 VDD.t102 VDD.t206 63.4219
R7529 VDD.t113 VDD.t102 63.4219
R7530 VDD.t114 VDD.t113 63.4219
R7531 VDD.t58 VDD.t114 63.4219
R7532 VDD.t483 VDD.t58 63.4219
R7533 VDD.t460 VDD.t483 63.4219
R7534 VDD.t461 VDD.t460 63.4219
R7535 VDD.t103 VDD.t461 63.4219
R7536 VDD.t117 VDD.t103 63.4219
R7537 VDD.t104 VDD.t117 63.4219
R7538 VDD.t552 VDD.t104 63.4219
R7539 VDD.t57 VDD.t552 63.4219
R7540 VDD.t488 VDD.t57 63.4219
R7541 VDD.t120 VDD.t488 63.4219
R7542 VDD.t553 VDD.t699 63.4219
R7543 VDD.t481 VDD.t717 63.4219
R7544 VDD.n5559 VDD.t310 62.8681
R7545 VDD.n5560 VDD.t571 62.8681
R7546 VDD.n5405 VDD.t490 61.2227
R7547 VDD.n5207 VDD.t60 59.5631
R7548 VDD.n5200 VDD.t116 59.5631
R7549 VDD.n5267 VDD.t700 59.5631
R7550 VDD.n5260 VDD.t482 59.5631
R7551 VDD.n3010 VDD.n2733 56.1076
R7552 VDD.n3008 VDD.n2733 56.1076
R7553 VDD.n3002 VDD.n2733 56.1076
R7554 VDD.n3000 VDD.n2733 56.1076
R7555 VDD.n2991 VDD.n2733 56.1076
R7556 VDD.n2943 VDD.n2733 56.1076
R7557 VDD.n2985 VDD.n2733 56.1076
R7558 VDD.n2979 VDD.n2733 56.1076
R7559 VDD.n3088 VDD.n2625 56.1076
R7560 VDD.n2628 VDD.n2625 56.1076
R7561 VDD.n3095 VDD.n2625 56.1076
R7562 VDD.n2625 VDD.n2624 56.1076
R7563 VDD.n2653 VDD.n2625 56.1076
R7564 VDD.n2661 VDD.n2625 56.1076
R7565 VDD.n2650 VDD.n2625 56.1076
R7566 VDD.n2668 VDD.n2625 56.1076
R7567 VDD.n2812 VDD.n2625 56.1076
R7568 VDD.n2806 VDD.n2625 56.1076
R7569 VDD.n2804 VDD.n2625 56.1076
R7570 VDD.n2759 VDD.n2733 56.1076
R7571 VDD.n2765 VDD.n2733 56.1076
R7572 VDD.n2767 VDD.n2733 56.1076
R7573 VDD.n2773 VDD.n2733 56.1076
R7574 VDD.n2899 VDD.n2733 56.1076
R7575 VDD.n2893 VDD.n2733 56.1076
R7576 VDD.n2891 VDD.n2733 56.1076
R7577 VDD.n2885 VDD.n2733 56.1076
R7578 VDD.n2847 VDD.n2625 56.1076
R7579 VDD.n2841 VDD.n2625 56.1076
R7580 VDD.n2839 VDD.n2625 56.1076
R7581 VDD.n2818 VDD.n2625 56.1076
R7582 VDD.n2820 VDD.n2625 56.1076
R7583 VDD.n5067 VDD.n5066 56.1076
R7584 VDD.n5066 VDD.n3900 56.1076
R7585 VDD.n5066 VDD.n3901 56.1076
R7586 VDD.n5066 VDD.n3902 56.1076
R7587 VDD.n5066 VDD.n3903 56.1076
R7588 VDD.n5066 VDD.n3904 56.1076
R7589 VDD.n5066 VDD.n3905 56.1076
R7590 VDD.n5066 VDD.n3906 56.1076
R7591 VDD.n4424 VDD.n4423 56.1076
R7592 VDD.n4423 VDD.n4150 56.1076
R7593 VDD.n4423 VDD.n4149 56.1076
R7594 VDD.n4423 VDD.n4148 56.1076
R7595 VDD.n4423 VDD.n4147 56.1076
R7596 VDD.n4423 VDD.n4146 56.1076
R7597 VDD.n4423 VDD.n4145 56.1076
R7598 VDD.n4423 VDD.n4144 56.1076
R7599 VDD.n5066 VDD.n5065 56.1076
R7600 VDD.n5066 VDD.n3893 56.1076
R7601 VDD.n5066 VDD.n3894 56.1076
R7602 VDD.n5066 VDD.n3895 56.1076
R7603 VDD.n5066 VDD.n3896 56.1076
R7604 VDD.n5066 VDD.n3897 56.1076
R7605 VDD.n5066 VDD.n3898 56.1076
R7606 VDD.n5066 VDD.n3899 56.1076
R7607 VDD.n4423 VDD.n4152 56.1076
R7608 VDD.n4423 VDD.n4153 56.1076
R7609 VDD.n4423 VDD.n4154 56.1076
R7610 VDD.n4423 VDD.n4155 56.1076
R7611 VDD.n4423 VDD.n4156 56.1076
R7612 VDD.n4423 VDD.n4157 56.1076
R7613 VDD.n4423 VDD.n4158 56.1076
R7614 VDD.n4423 VDD.n4159 56.1076
R7615 VDD.n4241 VDD.n4210 56.1076
R7616 VDD.n4241 VDD.n4209 56.1076
R7617 VDD.n4241 VDD.n4208 56.1076
R7618 VDD.n4241 VDD.n4207 56.1076
R7619 VDD.n4241 VDD.n4206 56.1076
R7620 VDD.n4241 VDD.n4205 56.1076
R7621 VDD.n4241 VDD.n4204 56.1076
R7622 VDD.n4242 VDD.n4241 56.1076
R7623 VDD.n4902 VDD.n4901 56.1076
R7624 VDD.n4902 VDD.n4837 56.1076
R7625 VDD.n4902 VDD.n4838 56.1076
R7626 VDD.n4902 VDD.n4839 56.1076
R7627 VDD.n4902 VDD.n4840 56.1076
R7628 VDD.n4902 VDD.n4841 56.1076
R7629 VDD.n4902 VDD.n4842 56.1076
R7630 VDD.n4902 VDD.n4843 56.1076
R7631 VDD.n416 VDD.n139 56.1076
R7632 VDD.n414 VDD.n139 56.1076
R7633 VDD.n408 VDD.n139 56.1076
R7634 VDD.n406 VDD.n139 56.1076
R7635 VDD.n397 VDD.n139 56.1076
R7636 VDD.n349 VDD.n139 56.1076
R7637 VDD.n391 VDD.n139 56.1076
R7638 VDD.n385 VDD.n139 56.1076
R7639 VDD.n494 VDD.n31 56.1076
R7640 VDD.n34 VDD.n31 56.1076
R7641 VDD.n501 VDD.n31 56.1076
R7642 VDD.n31 VDD.n30 56.1076
R7643 VDD.n59 VDD.n31 56.1076
R7644 VDD.n67 VDD.n31 56.1076
R7645 VDD.n56 VDD.n31 56.1076
R7646 VDD.n74 VDD.n31 56.1076
R7647 VDD.n218 VDD.n31 56.1076
R7648 VDD.n212 VDD.n31 56.1076
R7649 VDD.n210 VDD.n31 56.1076
R7650 VDD.n165 VDD.n139 56.1076
R7651 VDD.n171 VDD.n139 56.1076
R7652 VDD.n173 VDD.n139 56.1076
R7653 VDD.n179 VDD.n139 56.1076
R7654 VDD.n305 VDD.n139 56.1076
R7655 VDD.n299 VDD.n139 56.1076
R7656 VDD.n297 VDD.n139 56.1076
R7657 VDD.n291 VDD.n139 56.1076
R7658 VDD.n253 VDD.n31 56.1076
R7659 VDD.n247 VDD.n31 56.1076
R7660 VDD.n245 VDD.n31 56.1076
R7661 VDD.n224 VDD.n31 56.1076
R7662 VDD.n226 VDD.n31 56.1076
R7663 VDD.n2473 VDD.n2472 56.1076
R7664 VDD.n2472 VDD.n1306 56.1076
R7665 VDD.n2472 VDD.n1307 56.1076
R7666 VDD.n2472 VDD.n1308 56.1076
R7667 VDD.n2472 VDD.n1309 56.1076
R7668 VDD.n2472 VDD.n1310 56.1076
R7669 VDD.n2472 VDD.n1311 56.1076
R7670 VDD.n2472 VDD.n1312 56.1076
R7671 VDD.n1830 VDD.n1829 56.1076
R7672 VDD.n1829 VDD.n1556 56.1076
R7673 VDD.n1829 VDD.n1555 56.1076
R7674 VDD.n1829 VDD.n1554 56.1076
R7675 VDD.n1829 VDD.n1553 56.1076
R7676 VDD.n1829 VDD.n1552 56.1076
R7677 VDD.n1829 VDD.n1551 56.1076
R7678 VDD.n1829 VDD.n1550 56.1076
R7679 VDD.n2472 VDD.n2471 56.1076
R7680 VDD.n2472 VDD.n1299 56.1076
R7681 VDD.n2472 VDD.n1300 56.1076
R7682 VDD.n2472 VDD.n1301 56.1076
R7683 VDD.n2472 VDD.n1302 56.1076
R7684 VDD.n2472 VDD.n1303 56.1076
R7685 VDD.n2472 VDD.n1304 56.1076
R7686 VDD.n2472 VDD.n1305 56.1076
R7687 VDD.n1829 VDD.n1558 56.1076
R7688 VDD.n1829 VDD.n1559 56.1076
R7689 VDD.n1829 VDD.n1560 56.1076
R7690 VDD.n1829 VDD.n1561 56.1076
R7691 VDD.n1829 VDD.n1562 56.1076
R7692 VDD.n1829 VDD.n1563 56.1076
R7693 VDD.n1829 VDD.n1564 56.1076
R7694 VDD.n1829 VDD.n1565 56.1076
R7695 VDD.n1647 VDD.n1616 56.1076
R7696 VDD.n1647 VDD.n1615 56.1076
R7697 VDD.n1647 VDD.n1614 56.1076
R7698 VDD.n1647 VDD.n1613 56.1076
R7699 VDD.n1647 VDD.n1612 56.1076
R7700 VDD.n1647 VDD.n1611 56.1076
R7701 VDD.n1647 VDD.n1610 56.1076
R7702 VDD.n1648 VDD.n1647 56.1076
R7703 VDD.n2308 VDD.n2307 56.1076
R7704 VDD.n2308 VDD.n2243 56.1076
R7705 VDD.n2308 VDD.n2244 56.1076
R7706 VDD.n2308 VDD.n2245 56.1076
R7707 VDD.n2308 VDD.n2246 56.1076
R7708 VDD.n2308 VDD.n2247 56.1076
R7709 VDD.n2308 VDD.n2248 56.1076
R7710 VDD.n2308 VDD.n2249 56.1076
R7711 VDD.n5979 VDD.n5702 56.1076
R7712 VDD.n5977 VDD.n5702 56.1076
R7713 VDD.n5971 VDD.n5702 56.1076
R7714 VDD.n5969 VDD.n5702 56.1076
R7715 VDD.n5960 VDD.n5702 56.1076
R7716 VDD.n5912 VDD.n5702 56.1076
R7717 VDD.n5954 VDD.n5702 56.1076
R7718 VDD.n5948 VDD.n5702 56.1076
R7719 VDD.n6057 VDD.n5594 56.1076
R7720 VDD.n5597 VDD.n5594 56.1076
R7721 VDD.n6064 VDD.n5594 56.1076
R7722 VDD.n5594 VDD.n5593 56.1076
R7723 VDD.n5622 VDD.n5594 56.1076
R7724 VDD.n5630 VDD.n5594 56.1076
R7725 VDD.n5619 VDD.n5594 56.1076
R7726 VDD.n5637 VDD.n5594 56.1076
R7727 VDD.n5781 VDD.n5594 56.1076
R7728 VDD.n5775 VDD.n5594 56.1076
R7729 VDD.n5773 VDD.n5594 56.1076
R7730 VDD.n5728 VDD.n5702 56.1076
R7731 VDD.n5734 VDD.n5702 56.1076
R7732 VDD.n5736 VDD.n5702 56.1076
R7733 VDD.n5742 VDD.n5702 56.1076
R7734 VDD.n5868 VDD.n5702 56.1076
R7735 VDD.n5862 VDD.n5702 56.1076
R7736 VDD.n5860 VDD.n5702 56.1076
R7737 VDD.n5854 VDD.n5702 56.1076
R7738 VDD.n5816 VDD.n5594 56.1076
R7739 VDD.n5810 VDD.n5594 56.1076
R7740 VDD.n5808 VDD.n5594 56.1076
R7741 VDD.n5787 VDD.n5594 56.1076
R7742 VDD.n5789 VDD.n5594 56.1076
R7743 VDD.n8036 VDD.n8035 56.1076
R7744 VDD.n8035 VDD.n6869 56.1076
R7745 VDD.n8035 VDD.n6870 56.1076
R7746 VDD.n8035 VDD.n6871 56.1076
R7747 VDD.n8035 VDD.n6872 56.1076
R7748 VDD.n8035 VDD.n6873 56.1076
R7749 VDD.n8035 VDD.n6874 56.1076
R7750 VDD.n8035 VDD.n6875 56.1076
R7751 VDD.n7393 VDD.n7392 56.1076
R7752 VDD.n7392 VDD.n7119 56.1076
R7753 VDD.n7392 VDD.n7118 56.1076
R7754 VDD.n7392 VDD.n7117 56.1076
R7755 VDD.n7392 VDD.n7116 56.1076
R7756 VDD.n7392 VDD.n7115 56.1076
R7757 VDD.n7392 VDD.n7114 56.1076
R7758 VDD.n7392 VDD.n7113 56.1076
R7759 VDD.n8035 VDD.n8034 56.1076
R7760 VDD.n8035 VDD.n6862 56.1076
R7761 VDD.n8035 VDD.n6863 56.1076
R7762 VDD.n8035 VDD.n6864 56.1076
R7763 VDD.n8035 VDD.n6865 56.1076
R7764 VDD.n8035 VDD.n6866 56.1076
R7765 VDD.n8035 VDD.n6867 56.1076
R7766 VDD.n8035 VDD.n6868 56.1076
R7767 VDD.n7392 VDD.n7121 56.1076
R7768 VDD.n7392 VDD.n7122 56.1076
R7769 VDD.n7392 VDD.n7123 56.1076
R7770 VDD.n7392 VDD.n7124 56.1076
R7771 VDD.n7392 VDD.n7125 56.1076
R7772 VDD.n7392 VDD.n7126 56.1076
R7773 VDD.n7392 VDD.n7127 56.1076
R7774 VDD.n7392 VDD.n7128 56.1076
R7775 VDD.n7210 VDD.n7179 56.1076
R7776 VDD.n7210 VDD.n7178 56.1076
R7777 VDD.n7210 VDD.n7177 56.1076
R7778 VDD.n7210 VDD.n7176 56.1076
R7779 VDD.n7210 VDD.n7175 56.1076
R7780 VDD.n7210 VDD.n7174 56.1076
R7781 VDD.n7210 VDD.n7173 56.1076
R7782 VDD.n7211 VDD.n7210 56.1076
R7783 VDD.n7871 VDD.n7870 56.1076
R7784 VDD.n7871 VDD.n7806 56.1076
R7785 VDD.n7871 VDD.n7807 56.1076
R7786 VDD.n7871 VDD.n7808 56.1076
R7787 VDD.n7871 VDD.n7809 56.1076
R7788 VDD.n7871 VDD.n7810 56.1076
R7789 VDD.n7871 VDD.n7811 56.1076
R7790 VDD.n7871 VDD.n7812 56.1076
R7791 VDD.n5206 VDD.n5205 53.0621
R7792 VDD.n5266 VDD.n5265 53.0621
R7793 VDD.n3215 VDD.n3211 51.6897
R7794 VDD.n3289 VDD.n3285 51.6897
R7795 VDD.n3302 VDD.n3298 51.6897
R7796 VDD.n3315 VDD.n3311 51.6897
R7797 VDD.n3328 VDD.n3324 51.6897
R7798 VDD.n3272 VDD.n3268 51.6897
R7799 VDD.n3258 VDD.n3254 51.6897
R7800 VDD.n3244 VDD.n3240 51.6897
R7801 VDD.n3230 VDD.n3226 51.6897
R7802 VDD.n3171 VDD.n3167 51.6897
R7803 VDD.n621 VDD.n617 51.6897
R7804 VDD.n695 VDD.n691 51.6897
R7805 VDD.n708 VDD.n704 51.6897
R7806 VDD.n721 VDD.n717 51.6897
R7807 VDD.n734 VDD.n730 51.6897
R7808 VDD.n678 VDD.n674 51.6897
R7809 VDD.n664 VDD.n660 51.6897
R7810 VDD.n650 VDD.n646 51.6897
R7811 VDD.n636 VDD.n632 51.6897
R7812 VDD.n577 VDD.n573 51.6897
R7813 VDD.n6184 VDD.n6180 51.6897
R7814 VDD.n6258 VDD.n6254 51.6897
R7815 VDD.n6271 VDD.n6267 51.6897
R7816 VDD.n6284 VDD.n6280 51.6897
R7817 VDD.n6297 VDD.n6293 51.6897
R7818 VDD.n6241 VDD.n6237 51.6897
R7819 VDD.n6227 VDD.n6223 51.6897
R7820 VDD.n6213 VDD.n6209 51.6897
R7821 VDD.n6199 VDD.n6195 51.6897
R7822 VDD.n6140 VDD.n6136 51.6897
R7823 VDD.n3159 VDD.n3150 51.6837
R7824 VDD.n3392 VDD.n3383 51.6837
R7825 VDD.n3405 VDD.n3396 51.6837
R7826 VDD.n3418 VDD.n3409 51.6837
R7827 VDD.n3431 VDD.n3422 51.6837
R7828 VDD.n3375 VDD.n3366 51.6837
R7829 VDD.n3361 VDD.n3352 51.6837
R7830 VDD.n3347 VDD.n3338 51.6837
R7831 VDD.n3115 VDD.n3106 51.6837
R7832 VDD.n5172 VDD.n5163 51.6837
R7833 VDD.n565 VDD.n556 51.6837
R7834 VDD.n798 VDD.n789 51.6837
R7835 VDD.n811 VDD.n802 51.6837
R7836 VDD.n824 VDD.n815 51.6837
R7837 VDD.n837 VDD.n828 51.6837
R7838 VDD.n781 VDD.n772 51.6837
R7839 VDD.n767 VDD.n758 51.6837
R7840 VDD.n753 VDD.n744 51.6837
R7841 VDD.n521 VDD.n512 51.6837
R7842 VDD.n2578 VDD.n2569 51.6837
R7843 VDD.n6128 VDD.n6119 51.6837
R7844 VDD.n6361 VDD.n6352 51.6837
R7845 VDD.n6374 VDD.n6365 51.6837
R7846 VDD.n6387 VDD.n6378 51.6837
R7847 VDD.n6400 VDD.n6391 51.6837
R7848 VDD.n6344 VDD.n6335 51.6837
R7849 VDD.n6330 VDD.n6321 51.6837
R7850 VDD.n6316 VDD.n6307 51.6837
R7851 VDD.n6084 VDD.n6075 51.6837
R7852 VDD.n8141 VDD.n8132 51.6837
R7853 VDD.n3636 VDD.n3632 51.6704
R7854 VDD.n3650 VDD.n3646 51.6704
R7855 VDD.n3663 VDD.n3659 51.6704
R7856 VDD.n3676 VDD.n3672 51.6704
R7857 VDD.n3689 VDD.n3685 51.6704
R7858 VDD.n3702 VDD.n3698 51.6704
R7859 VDD.n3715 VDD.n3711 51.6704
R7860 VDD.n3729 VDD.n3725 51.6704
R7861 VDD.n3742 VDD.n3738 51.6704
R7862 VDD.n3755 VDD.n3751 51.6704
R7863 VDD.n3768 VDD.n3764 51.6704
R7864 VDD.n3781 VDD.n3777 51.6704
R7865 VDD.n3582 VDD.n3578 51.6704
R7866 VDD.n3568 VDD.n3564 51.6704
R7867 VDD.n3554 VDD.n3550 51.6704
R7868 VDD.n3540 VDD.n3536 51.6704
R7869 VDD.n3526 VDD.n3522 51.6704
R7870 VDD.n3512 VDD.n3508 51.6704
R7871 VDD.n3497 VDD.n3493 51.6704
R7872 VDD.n1042 VDD.n1038 51.6704
R7873 VDD.n1056 VDD.n1052 51.6704
R7874 VDD.n1069 VDD.n1065 51.6704
R7875 VDD.n1082 VDD.n1078 51.6704
R7876 VDD.n1095 VDD.n1091 51.6704
R7877 VDD.n1108 VDD.n1104 51.6704
R7878 VDD.n1121 VDD.n1117 51.6704
R7879 VDD.n1135 VDD.n1131 51.6704
R7880 VDD.n1148 VDD.n1144 51.6704
R7881 VDD.n1161 VDD.n1157 51.6704
R7882 VDD.n1174 VDD.n1170 51.6704
R7883 VDD.n1187 VDD.n1183 51.6704
R7884 VDD.n988 VDD.n984 51.6704
R7885 VDD.n974 VDD.n970 51.6704
R7886 VDD.n960 VDD.n956 51.6704
R7887 VDD.n946 VDD.n942 51.6704
R7888 VDD.n932 VDD.n928 51.6704
R7889 VDD.n918 VDD.n914 51.6704
R7890 VDD.n903 VDD.n899 51.6704
R7891 VDD.n6605 VDD.n6601 51.6704
R7892 VDD.n6619 VDD.n6615 51.6704
R7893 VDD.n6632 VDD.n6628 51.6704
R7894 VDD.n6645 VDD.n6641 51.6704
R7895 VDD.n6658 VDD.n6654 51.6704
R7896 VDD.n6671 VDD.n6667 51.6704
R7897 VDD.n6684 VDD.n6680 51.6704
R7898 VDD.n6698 VDD.n6694 51.6704
R7899 VDD.n6711 VDD.n6707 51.6704
R7900 VDD.n6724 VDD.n6720 51.6704
R7901 VDD.n6737 VDD.n6733 51.6704
R7902 VDD.n6750 VDD.n6746 51.6704
R7903 VDD.n6551 VDD.n6547 51.6704
R7904 VDD.n6537 VDD.n6533 51.6704
R7905 VDD.n6523 VDD.n6519 51.6704
R7906 VDD.n6509 VDD.n6505 51.6704
R7907 VDD.n6495 VDD.n6491 51.6704
R7908 VDD.n6481 VDD.n6477 51.6704
R7909 VDD.n6466 VDD.n6462 51.6704
R7910 VDD.n2918 VDD.n2917 51.0589
R7911 VDD.n2916 VDD.n2915 51.0589
R7912 VDD.n324 VDD.n323 51.0589
R7913 VDD.n322 VDD.n321 51.0589
R7914 VDD.n5887 VDD.n5886 51.0589
R7915 VDD.n5885 VDD.n5884 51.0589
R7916 VDD.n2741 VDD.n2740 51.0019
R7917 VDD.n2791 VDD.n2788 51.0019
R7918 VDD.n147 VDD.n146 51.0019
R7919 VDD.n197 VDD.n194 51.0019
R7920 VDD.n5710 VDD.n5709 51.0019
R7921 VDD.n5760 VDD.n5757 51.0019
R7922 VDD.n5220 VDD.n5219 46.4801
R7923 VDD.n5277 VDD.n5276 46.4801
R7924 VDD.n5241 VDD.n5191 40.5181
R7925 VDD.n5290 VDD.n5289 40.5181
R7926 VDD.n5360 VDD.t475 40.1116
R7927 VDD.n5424 VDD.t691 35.8894
R7928 VDD VDD.n5536 34.927
R7929 VDD.n5537 VDD.t585 34.927
R7930 VDD.n5452 VDD.n5446 34.6358
R7931 VDD.n5452 VDD.n5451 34.6358
R7932 VDD.n5554 VDD.n5553 34.6358
R7933 VDD.n5543 VDD.n5542 34.6358
R7934 VDD.n5531 VDD.n5530 34.6358
R7935 VDD.n5524 VDD.n5521 34.6358
R7936 VDD.n5519 VDD.n5475 34.6358
R7937 VDD.n5507 VDD.n5506 34.6358
R7938 VDD.n5498 VDD.n5484 34.6358
R7939 VDD.n5418 VDD.n5417 34.6358
R7940 VDD.n5437 VDD.n5436 34.6358
R7941 VDD.n5399 VDD.n5398 34.6358
R7942 VDD.n5389 VDD.n5330 34.6358
R7943 VDD.n5372 VDD.n5369 34.6358
R7944 VDD.n5355 VDD.n5354 34.6358
R7945 VDD.n2632 VDD.n2625 34.2522
R7946 VDD.n3016 VDD.n2733 34.2522
R7947 VDD.n38 VDD.n31 34.2522
R7948 VDD.n422 VDD.n139 34.2522
R7949 VDD.n5601 VDD.n5594 34.2522
R7950 VDD.n5985 VDD.n5702 34.2522
R7951 VDD.n5546 VDD.n5545 33.8829
R7952 VDD.n5535 VDD.n5534 33.5064
R7953 VDD.n5523 VDD.n5522 32.7534
R7954 VDD.n5563 VDD.n5442 32.164
R7955 VDD.n5211 VDD.t484 31.7112
R7956 VDD.t713 VDD.n5211 31.7112
R7957 VDD.n5271 VDD.t553 31.7112
R7958 VDD.t717 VDD.n5271 31.7112
R7959 VDD.n5457 VDD.n5456 31.2476
R7960 VDD.n5557 VDD.n5464 30.8711
R7961 VDD.n5534 VDD.n5472 30.8711
R7962 VDD.n5521 VDD.n5520 30.8711
R7963 VDD.n5500 VDD.n5499 30.8711
R7964 VDD.n5377 VDD.n5335 30.8711
R7965 VDD.n5353 VDD.n5352 30.8711
R7966 VDD.n5359 VDD.n5358 30.4946
R7967 VDD.n5367 VDD.n5338 30.2283
R7968 VDD.n3634 VDD.n3632 29.8117
R7969 VDD.n3648 VDD.n3646 29.8117
R7970 VDD.n3661 VDD.n3659 29.8117
R7971 VDD.n3674 VDD.n3672 29.8117
R7972 VDD.n3687 VDD.n3685 29.8117
R7973 VDD.n3700 VDD.n3698 29.8117
R7974 VDD.n3713 VDD.n3711 29.8117
R7975 VDD.n3727 VDD.n3725 29.8117
R7976 VDD.n3740 VDD.n3738 29.8117
R7977 VDD.n3753 VDD.n3751 29.8117
R7978 VDD.n3766 VDD.n3764 29.8117
R7979 VDD.n3779 VDD.n3777 29.8117
R7980 VDD.n3580 VDD.n3578 29.8117
R7981 VDD.n3566 VDD.n3564 29.8117
R7982 VDD.n3552 VDD.n3550 29.8117
R7983 VDD.n3538 VDD.n3536 29.8117
R7984 VDD.n3524 VDD.n3522 29.8117
R7985 VDD.n3510 VDD.n3508 29.8117
R7986 VDD.n3495 VDD.n3493 29.8117
R7987 VDD.n1040 VDD.n1038 29.8117
R7988 VDD.n1054 VDD.n1052 29.8117
R7989 VDD.n1067 VDD.n1065 29.8117
R7990 VDD.n1080 VDD.n1078 29.8117
R7991 VDD.n1093 VDD.n1091 29.8117
R7992 VDD.n1106 VDD.n1104 29.8117
R7993 VDD.n1119 VDD.n1117 29.8117
R7994 VDD.n1133 VDD.n1131 29.8117
R7995 VDD.n1146 VDD.n1144 29.8117
R7996 VDD.n1159 VDD.n1157 29.8117
R7997 VDD.n1172 VDD.n1170 29.8117
R7998 VDD.n1185 VDD.n1183 29.8117
R7999 VDD.n986 VDD.n984 29.8117
R8000 VDD.n972 VDD.n970 29.8117
R8001 VDD.n958 VDD.n956 29.8117
R8002 VDD.n944 VDD.n942 29.8117
R8003 VDD.n930 VDD.n928 29.8117
R8004 VDD.n916 VDD.n914 29.8117
R8005 VDD.n901 VDD.n899 29.8117
R8006 VDD.n6603 VDD.n6601 29.8117
R8007 VDD.n6617 VDD.n6615 29.8117
R8008 VDD.n6630 VDD.n6628 29.8117
R8009 VDD.n6643 VDD.n6641 29.8117
R8010 VDD.n6656 VDD.n6654 29.8117
R8011 VDD.n6669 VDD.n6667 29.8117
R8012 VDD.n6682 VDD.n6680 29.8117
R8013 VDD.n6696 VDD.n6694 29.8117
R8014 VDD.n6709 VDD.n6707 29.8117
R8015 VDD.n6722 VDD.n6720 29.8117
R8016 VDD.n6735 VDD.n6733 29.8117
R8017 VDD.n6748 VDD.n6746 29.8117
R8018 VDD.n6549 VDD.n6547 29.8117
R8019 VDD.n6535 VDD.n6533 29.8117
R8020 VDD.n6521 VDD.n6519 29.8117
R8021 VDD.n6507 VDD.n6505 29.8117
R8022 VDD.n6493 VDD.n6491 29.8117
R8023 VDD.n6479 VDD.n6477 29.8117
R8024 VDD.n6464 VDD.n6462 29.8117
R8025 VDD.n3159 VDD.n3158 29.8077
R8026 VDD.n3392 VDD.n3391 29.8077
R8027 VDD.n3405 VDD.n3404 29.8077
R8028 VDD.n3418 VDD.n3417 29.8077
R8029 VDD.n3431 VDD.n3430 29.8077
R8030 VDD.n3375 VDD.n3374 29.8077
R8031 VDD.n3361 VDD.n3360 29.8077
R8032 VDD.n3347 VDD.n3346 29.8077
R8033 VDD.n3115 VDD.n3114 29.8077
R8034 VDD.n5172 VDD.n5171 29.8077
R8035 VDD.n565 VDD.n564 29.8077
R8036 VDD.n798 VDD.n797 29.8077
R8037 VDD.n811 VDD.n810 29.8077
R8038 VDD.n824 VDD.n823 29.8077
R8039 VDD.n837 VDD.n836 29.8077
R8040 VDD.n781 VDD.n780 29.8077
R8041 VDD.n767 VDD.n766 29.8077
R8042 VDD.n753 VDD.n752 29.8077
R8043 VDD.n521 VDD.n520 29.8077
R8044 VDD.n2578 VDD.n2577 29.8077
R8045 VDD.n6128 VDD.n6127 29.8077
R8046 VDD.n6361 VDD.n6360 29.8077
R8047 VDD.n6374 VDD.n6373 29.8077
R8048 VDD.n6387 VDD.n6386 29.8077
R8049 VDD.n6400 VDD.n6399 29.8077
R8050 VDD.n6344 VDD.n6343 29.8077
R8051 VDD.n6330 VDD.n6329 29.8077
R8052 VDD.n6316 VDD.n6315 29.8077
R8053 VDD.n6084 VDD.n6083 29.8077
R8054 VDD.n8141 VDD.n8140 29.8077
R8055 VDD.n3213 VDD.n3211 29.806
R8056 VDD.n3287 VDD.n3285 29.806
R8057 VDD.n3300 VDD.n3298 29.806
R8058 VDD.n3313 VDD.n3311 29.806
R8059 VDD.n3326 VDD.n3324 29.806
R8060 VDD.n3270 VDD.n3268 29.806
R8061 VDD.n3256 VDD.n3254 29.806
R8062 VDD.n3242 VDD.n3240 29.806
R8063 VDD.n3228 VDD.n3226 29.806
R8064 VDD.n3169 VDD.n3167 29.806
R8065 VDD.n619 VDD.n617 29.806
R8066 VDD.n693 VDD.n691 29.806
R8067 VDD.n706 VDD.n704 29.806
R8068 VDD.n719 VDD.n717 29.806
R8069 VDD.n732 VDD.n730 29.806
R8070 VDD.n676 VDD.n674 29.806
R8071 VDD.n662 VDD.n660 29.806
R8072 VDD.n648 VDD.n646 29.806
R8073 VDD.n634 VDD.n632 29.806
R8074 VDD.n575 VDD.n573 29.806
R8075 VDD.n6182 VDD.n6180 29.806
R8076 VDD.n6256 VDD.n6254 29.806
R8077 VDD.n6269 VDD.n6267 29.806
R8078 VDD.n6282 VDD.n6280 29.806
R8079 VDD.n6295 VDD.n6293 29.806
R8080 VDD.n6239 VDD.n6237 29.806
R8081 VDD.n6225 VDD.n6223 29.806
R8082 VDD.n6211 VDD.n6209 29.806
R8083 VDD.n6197 VDD.n6195 29.806
R8084 VDD.n6138 VDD.n6136 29.806
R8085 VDD.n2607 VDD.n2605 29.3167
R8086 VDD.n2926 VDD.n2924 29.3167
R8087 VDD.n3138 VDD.n3137 29.3167
R8088 VDD.n3189 VDD.n3188 29.3167
R8089 VDD.n3610 VDD.n3609 29.3167
R8090 VDD.n3470 VDD.n3469 29.3167
R8091 VDD.n13 VDD.n11 29.3167
R8092 VDD.n332 VDD.n330 29.3167
R8093 VDD.n544 VDD.n543 29.3167
R8094 VDD.n595 VDD.n594 29.3167
R8095 VDD.n1016 VDD.n1015 29.3167
R8096 VDD.n876 VDD.n875 29.3167
R8097 VDD.n5576 VDD.n5574 29.3167
R8098 VDD.n5895 VDD.n5893 29.3167
R8099 VDD.n6107 VDD.n6106 29.3167
R8100 VDD.n6158 VDD.n6157 29.3167
R8101 VDD.n6579 VDD.n6578 29.3167
R8102 VDD.n6439 VDD.n6438 29.3167
R8103 VDD.n2753 VDD.n2752 29.2693
R8104 VDD.n2833 VDD.n2832 29.2693
R8105 VDD.n159 VDD.n158 29.2693
R8106 VDD.n239 VDD.n238 29.2693
R8107 VDD.n5722 VDD.n5721 29.2693
R8108 VDD.n5802 VDD.n5801 29.2693
R8109 VDD.n5558 VDD.n5462 28.2358
R8110 VDD.n5384 VDD.n5330 28.2358
R8111 VDD.n2910 VDD.n2742 27.5029
R8112 VDD.n2795 VDD.n2794 27.5029
R8113 VDD.n316 VDD.n148 27.5029
R8114 VDD.n201 VDD.n200 27.5029
R8115 VDD.n5879 VDD.n5711 27.5029
R8116 VDD.n5764 VDD.n5763 27.5029
R8117 VDD.t462 VDD.n5423 27.4449
R8118 VDD.n5392 VDD.n5390 27.1064
R8119 VDD.n5448 VDD.t684 26.5955
R8120 VDD.n5448 VDD.t690 26.5955
R8121 VDD.n5443 VDD.t578 26.5955
R8122 VDD.n5443 VDD.t572 26.5955
R8123 VDD.n5551 VDD.t173 26.5955
R8124 VDD.n5551 VDD.t574 26.5955
R8125 VDD.n5463 VDD.t15 26.5955
R8126 VDD.n5463 VDD.t382 26.5955
R8127 VDD.n5466 VDD.t586 26.5955
R8128 VDD.n5466 VDD.t588 26.5955
R8129 VDD.n5528 VDD.t66 26.5955
R8130 VDD.n5528 VDD.t584 26.5955
R8131 VDD.n5471 VDD.t277 26.5955
R8132 VDD.n5471 VDD.t541 26.5955
R8133 VDD.n5474 VDD.t220 26.5955
R8134 VDD.n5474 VDD.t135 26.5955
R8135 VDD.n5478 VDD.t672 26.5955
R8136 VDD.n5478 VDD.t108 26.5955
R8137 VDD.n5504 VDD.t676 26.5955
R8138 VDD.n5504 VDD.t670 26.5955
R8139 VDD.n5483 VDD.t235 26.5955
R8140 VDD.n5483 VDD.t237 26.5955
R8141 VDD.n5492 VDD.t566 26.5955
R8142 VDD.n5492 VDD.t233 26.5955
R8143 VDD.n5487 VDD.t568 26.5955
R8144 VDD.n5487 VDD.t570 26.5955
R8145 VDD.n5329 VDD.t224 26.5955
R8146 VDD.n5329 VDD.t291 26.5955
R8147 VDD.n5344 VDD.t551 26.5955
R8148 VDD.n5344 VDD.t476 26.5955
R8149 VDD.n5312 VDD.t521 26.5955
R8150 VDD.n5312 VDD.t682 26.5955
R8151 VDD.n5314 VDD.t688 26.5955
R8152 VDD.n5314 VDD.t692 26.5955
R8153 VDD.n5318 VDD.t463 26.5955
R8154 VDD.n5318 VDD.t258 26.5955
R8155 VDD.n5321 VDD.t491 26.5955
R8156 VDD.n5321 VDD.t493 26.5955
R8157 VDD.n5326 VDD.t531 26.5955
R8158 VDD.n5326 VDD.t525 26.5955
R8159 VDD.n5396 VDD.t527 26.5955
R8160 VDD.n5396 VDD.t495 26.5955
R8161 VDD.n5334 VDD.t281 26.5955
R8162 VDD.n5334 VDD.t321 26.5955
R8163 VDD.n5337 VDD.t288 26.5955
R8164 VDD.n5337 VDD.t186 26.5955
R8165 VDD.n5370 VDD.t339 26.5955
R8166 VDD.n5370 VDD.t245 26.5955
R8167 VDD.n5342 VDD.t369 26.5955
R8168 VDD.n5342 VDD.t304 26.5955
R8169 VDD.n5349 VDD.t300 26.5955
R8170 VDD.n5349 VDD.t302 26.5955
R8171 VDD.n5203 VDD.n5201 26.4291
R8172 VDD.n5211 VDD.n5203 26.4291
R8173 VDD.n5204 VDD.n5202 26.4291
R8174 VDD.n5211 VDD.n5204 26.4291
R8175 VDD.n5263 VDD.n5261 26.4291
R8176 VDD.n5271 VDD.n5263 26.4291
R8177 VDD.n5264 VDD.n5262 26.4291
R8178 VDD.n5271 VDD.n5264 26.4291
R8179 VDD.n2616 VDD.n2600 26.212
R8180 VDD.n2935 VDD.n2919 26.212
R8181 VDD.n22 VDD.n6 26.212
R8182 VDD.n341 VDD.n325 26.212
R8183 VDD.n5585 VDD.n5569 26.212
R8184 VDD.n5904 VDD.n5888 26.212
R8185 VDD.n5430 VDD.n5427 25.977
R8186 VDD.n5433 VDD.n5432 25.977
R8187 VDD.n5411 VDD.n5410 25.977
R8188 VDD.n5377 VDD.n5376 25.977
R8189 VDD.n5352 VDD.n5339 25.977
R8190 VDD.n2751 VDD.n2746 25.6005
R8191 VDD.n2673 VDD.n2672 25.6005
R8192 VDD.n2674 VDD.n2673 25.6005
R8193 VDD.n3074 VDD.n2674 25.6005
R8194 VDD.n3074 VDD.n3073 25.6005
R8195 VDD.n3073 VDD.n3072 25.6005
R8196 VDD.n3072 VDD.n2675 25.6005
R8197 VDD.n3062 VDD.n2675 25.6005
R8198 VDD.n3062 VDD.n3061 25.6005
R8199 VDD.n3061 VDD.n3060 25.6005
R8200 VDD.n3060 VDD.n2687 25.6005
R8201 VDD.n3050 VDD.n2687 25.6005
R8202 VDD.n3050 VDD.n3049 25.6005
R8203 VDD.n3049 VDD.n3048 25.6005
R8204 VDD.n3048 VDD.n2699 25.6005
R8205 VDD.n3038 VDD.n2699 25.6005
R8206 VDD.n3038 VDD.n3037 25.6005
R8207 VDD.n3037 VDD.n3036 25.6005
R8208 VDD.n3036 VDD.n2711 25.6005
R8209 VDD.n3026 VDD.n2711 25.6005
R8210 VDD.n3026 VDD.n3025 25.6005
R8211 VDD.n3025 VDD.n3024 25.6005
R8212 VDD.n3024 VDD.n2723 25.6005
R8213 VDD.n3014 VDD.n2723 25.6005
R8214 VDD.n2647 VDD.n2646 25.6005
R8215 VDD.n2666 VDD.n2647 25.6005
R8216 VDD.n2666 VDD.n2665 25.6005
R8217 VDD.n2665 VDD.n2664 25.6005
R8218 VDD.n2664 VDD.n2649 25.6005
R8219 VDD.n2659 VDD.n2649 25.6005
R8220 VDD.n3098 VDD.n2623 25.6005
R8221 VDD.n3093 VDD.n2623 25.6005
R8222 VDD.n3093 VDD.n3092 25.6005
R8223 VDD.n3092 VDD.n3091 25.6005
R8224 VDD.n3091 VDD.n2627 25.6005
R8225 VDD.n3086 VDD.n2627 25.6005
R8226 VDD.n3085 VDD.n3084 25.6005
R8227 VDD.n3084 VDD.n2630 25.6005
R8228 VDD.n2946 VDD.n2630 25.6005
R8229 VDD.n2948 VDD.n2946 25.6005
R8230 VDD.n2949 VDD.n2948 25.6005
R8231 VDD.n2951 VDD.n2949 25.6005
R8232 VDD.n2952 VDD.n2951 25.6005
R8233 VDD.n2954 VDD.n2952 25.6005
R8234 VDD.n2955 VDD.n2954 25.6005
R8235 VDD.n2957 VDD.n2955 25.6005
R8236 VDD.n2958 VDD.n2957 25.6005
R8237 VDD.n2960 VDD.n2958 25.6005
R8238 VDD.n2961 VDD.n2960 25.6005
R8239 VDD.n2963 VDD.n2961 25.6005
R8240 VDD.n2964 VDD.n2963 25.6005
R8241 VDD.n2966 VDD.n2964 25.6005
R8242 VDD.n2967 VDD.n2966 25.6005
R8243 VDD.n2969 VDD.n2967 25.6005
R8244 VDD.n2970 VDD.n2969 25.6005
R8245 VDD.n2972 VDD.n2970 25.6005
R8246 VDD.n2973 VDD.n2972 25.6005
R8247 VDD.n2975 VDD.n2973 25.6005
R8248 VDD.n2976 VDD.n2975 25.6005
R8249 VDD.n2989 VDD.n2988 25.6005
R8250 VDD.n2988 VDD.n2944 25.6005
R8251 VDD.n2983 VDD.n2944 25.6005
R8252 VDD.n2983 VDD.n2982 25.6005
R8253 VDD.n2982 VDD.n2981 25.6005
R8254 VDD.n2981 VDD.n2977 25.6005
R8255 VDD.n3013 VDD.n3012 25.6005
R8256 VDD.n3012 VDD.n2735 25.6005
R8257 VDD.n3006 VDD.n2735 25.6005
R8258 VDD.n3006 VDD.n3005 25.6005
R8259 VDD.n3005 VDD.n3004 25.6005
R8260 VDD.n3004 VDD.n2737 25.6005
R8261 VDD.n2802 VDD.n2801 25.6005
R8262 VDD.n2808 VDD.n2801 25.6005
R8263 VDD.n2809 VDD.n2808 25.6005
R8264 VDD.n2810 VDD.n2809 25.6005
R8265 VDD.n2810 VDD.n2799 25.6005
R8266 VDD.n2799 VDD.n2798 25.6005
R8267 VDD.n3080 VDD.n2638 25.6005
R8268 VDD.n3080 VDD.n3079 25.6005
R8269 VDD.n3079 VDD.n3078 25.6005
R8270 VDD.n3078 VDD.n2639 25.6005
R8271 VDD.n3068 VDD.n2639 25.6005
R8272 VDD.n3068 VDD.n3067 25.6005
R8273 VDD.n3067 VDD.n3066 25.6005
R8274 VDD.n3066 VDD.n2680 25.6005
R8275 VDD.n3056 VDD.n2680 25.6005
R8276 VDD.n3056 VDD.n3055 25.6005
R8277 VDD.n3055 VDD.n3054 25.6005
R8278 VDD.n3054 VDD.n2692 25.6005
R8279 VDD.n3044 VDD.n2692 25.6005
R8280 VDD.n3044 VDD.n3043 25.6005
R8281 VDD.n3043 VDD.n3042 25.6005
R8282 VDD.n3042 VDD.n2704 25.6005
R8283 VDD.n3032 VDD.n2704 25.6005
R8284 VDD.n3032 VDD.n3031 25.6005
R8285 VDD.n3031 VDD.n3030 25.6005
R8286 VDD.n3030 VDD.n2716 25.6005
R8287 VDD.n3020 VDD.n2716 25.6005
R8288 VDD.n3020 VDD.n3019 25.6005
R8289 VDD.n3019 VDD.n3018 25.6005
R8290 VDD.n2761 VDD.n2729 25.6005
R8291 VDD.n2762 VDD.n2761 25.6005
R8292 VDD.n2763 VDD.n2762 25.6005
R8293 VDD.n2763 VDD.n2757 25.6005
R8294 VDD.n2769 VDD.n2757 25.6005
R8295 VDD.n2770 VDD.n2769 25.6005
R8296 VDD.n2897 VDD.n2896 25.6005
R8297 VDD.n2896 VDD.n2895 25.6005
R8298 VDD.n2895 VDD.n2776 25.6005
R8299 VDD.n2889 VDD.n2776 25.6005
R8300 VDD.n2889 VDD.n2888 25.6005
R8301 VDD.n2888 VDD.n2887 25.6005
R8302 VDD.n2851 VDD.n2850 25.6005
R8303 VDD.n2853 VDD.n2851 25.6005
R8304 VDD.n2854 VDD.n2853 25.6005
R8305 VDD.n2856 VDD.n2854 25.6005
R8306 VDD.n2857 VDD.n2856 25.6005
R8307 VDD.n2859 VDD.n2857 25.6005
R8308 VDD.n2860 VDD.n2859 25.6005
R8309 VDD.n2862 VDD.n2860 25.6005
R8310 VDD.n2863 VDD.n2862 25.6005
R8311 VDD.n2865 VDD.n2863 25.6005
R8312 VDD.n2866 VDD.n2865 25.6005
R8313 VDD.n2868 VDD.n2866 25.6005
R8314 VDD.n2869 VDD.n2868 25.6005
R8315 VDD.n2871 VDD.n2869 25.6005
R8316 VDD.n2872 VDD.n2871 25.6005
R8317 VDD.n2874 VDD.n2872 25.6005
R8318 VDD.n2875 VDD.n2874 25.6005
R8319 VDD.n2877 VDD.n2875 25.6005
R8320 VDD.n2878 VDD.n2877 25.6005
R8321 VDD.n2880 VDD.n2878 25.6005
R8322 VDD.n2881 VDD.n2880 25.6005
R8323 VDD.n2883 VDD.n2881 25.6005
R8324 VDD.n2884 VDD.n2883 25.6005
R8325 VDD.n2837 VDD.n2836 25.6005
R8326 VDD.n2837 VDD.n2780 25.6005
R8327 VDD.n2843 VDD.n2780 25.6005
R8328 VDD.n2844 VDD.n2843 25.6005
R8329 VDD.n2845 VDD.n2844 25.6005
R8330 VDD.n2845 VDD.n2778 25.6005
R8331 VDD.n2831 VDD.n2830 25.6005
R8332 VDD.n4433 VDD.n4136 25.6005
R8333 VDD.n4434 VDD.n4433 25.6005
R8334 VDD.n4436 VDD.n4434 25.6005
R8335 VDD.n4436 VDD.n4435 25.6005
R8336 VDD.n4435 VDD.n4108 25.6005
R8337 VDD.n4480 VDD.n4108 25.6005
R8338 VDD.n4481 VDD.n4480 25.6005
R8339 VDD.n4482 VDD.n4481 25.6005
R8340 VDD.n4482 VDD.n4100 25.6005
R8341 VDD.n4421 VDD.n4420 25.6005
R8342 VDD.n4420 VDD.n4419 25.6005
R8343 VDD.n4419 VDD.n4416 25.6005
R8344 VDD.n4416 VDD.n4415 25.6005
R8345 VDD.n4415 VDD.n4412 25.6005
R8346 VDD.n4412 VDD.n4411 25.6005
R8347 VDD.n4411 VDD.n4408 25.6005
R8348 VDD.n4408 VDD.n4407 25.6005
R8349 VDD.n4407 VDD.n4404 25.6005
R8350 VDD.n4404 VDD.n4403 25.6005
R8351 VDD.n4403 VDD.n4400 25.6005
R8352 VDD.n4400 VDD.n4399 25.6005
R8353 VDD.n4399 VDD.n4396 25.6005
R8354 VDD.n4396 VDD.n4395 25.6005
R8355 VDD.n4395 VDD.n4392 25.6005
R8356 VDD.n4392 VDD.n4391 25.6005
R8357 VDD.n4389 VDD.n4119 25.6005
R8358 VDD.n4467 VDD.n4119 25.6005
R8359 VDD.n4468 VDD.n4467 25.6005
R8360 VDD.n4470 VDD.n4468 25.6005
R8361 VDD.n4470 VDD.n4469 25.6005
R8362 VDD.n4469 VDD.n4092 25.6005
R8363 VDD.n4501 VDD.n4092 25.6005
R8364 VDD.n4502 VDD.n4501 25.6005
R8365 VDD.n4504 VDD.n4502 25.6005
R8366 VDD.n4504 VDD.n4503 25.6005
R8367 VDD.n4503 VDD.n4069 25.6005
R8368 VDD.n4534 VDD.n4069 25.6005
R8369 VDD.n4669 VDD.n4668 25.6005
R8370 VDD.n5112 VDD.n5111 25.6005
R8371 VDD.n5111 VDD.n5110 25.6005
R8372 VDD.n5110 VDD.n3824 25.6005
R8373 VDD.n3863 VDD.n3824 25.6005
R8374 VDD.n3864 VDD.n3863 25.6005
R8375 VDD.n5089 VDD.n3864 25.6005
R8376 VDD.n5089 VDD.n5088 25.6005
R8377 VDD.n5088 VDD.n5087 25.6005
R8378 VDD.n5087 VDD.n3865 25.6005
R8379 VDD.n5077 VDD.n3865 25.6005
R8380 VDD.n5077 VDD.n5076 25.6005
R8381 VDD.n5076 VDD.n5075 25.6005
R8382 VDD.n5063 VDD.n3884 25.6005
R8383 VDD.n5063 VDD.n5062 25.6005
R8384 VDD.n5062 VDD.n5061 25.6005
R8385 VDD.n5061 VDD.n5059 25.6005
R8386 VDD.n5059 VDD.n5056 25.6005
R8387 VDD.n5056 VDD.n5055 25.6005
R8388 VDD.n5055 VDD.n5052 25.6005
R8389 VDD.n5052 VDD.n5051 25.6005
R8390 VDD.n5051 VDD.n5048 25.6005
R8391 VDD.n5048 VDD.n5047 25.6005
R8392 VDD.n5047 VDD.n5044 25.6005
R8393 VDD.n5044 VDD.n5043 25.6005
R8394 VDD.n5043 VDD.n5040 25.6005
R8395 VDD.n5040 VDD.n5039 25.6005
R8396 VDD.n5039 VDD.n5036 25.6005
R8397 VDD.n5036 VDD.n5035 25.6005
R8398 VDD.n3872 VDD.n3832 25.6005
R8399 VDD.n3875 VDD.n3872 25.6005
R8400 VDD.n3876 VDD.n3875 25.6005
R8401 VDD.n3877 VDD.n3876 25.6005
R8402 VDD.n5083 VDD.n3877 25.6005
R8403 VDD.n5083 VDD.n5082 25.6005
R8404 VDD.n5082 VDD.n5081 25.6005
R8405 VDD.n5081 VDD.n3878 25.6005
R8406 VDD.n5071 VDD.n3878 25.6005
R8407 VDD.n5104 VDD.n3833 25.6005
R8408 VDD.n3915 VDD.n3833 25.6005
R8409 VDD.n3916 VDD.n3915 25.6005
R8410 VDD.n4992 VDD.n3916 25.6005
R8411 VDD.n4993 VDD.n4992 25.6005
R8412 VDD.n4994 VDD.n4993 25.6005
R8413 VDD.n4994 VDD.n3910 25.6005
R8414 VDD.n5032 VDD.n3910 25.6005
R8415 VDD.n5033 VDD.n5032 25.6005
R8416 VDD.n4584 VDD.n4583 25.6005
R8417 VDD.n4583 VDD.n4582 25.6005
R8418 VDD.n4582 VDD.n4011 25.6005
R8419 VDD.n4650 VDD.n4011 25.6005
R8420 VDD.n4650 VDD.n4649 25.6005
R8421 VDD.n4649 VDD.n4648 25.6005
R8422 VDD.n4648 VDD.n4647 25.6005
R8423 VDD.n4647 VDD.n4015 25.6005
R8424 VDD.n4015 VDD.n4014 25.6005
R8425 VDD.n4014 VDD.n4013 25.6005
R8426 VDD.n4013 VDD.n3931 25.6005
R8427 VDD.n4727 VDD.n3931 25.6005
R8428 VDD.n4728 VDD.n4727 25.6005
R8429 VDD.n4054 VDD.n4053 25.6005
R8430 VDD.n4053 VDD.n4021 25.6005
R8431 VDD.n4626 VDD.n4021 25.6005
R8432 VDD.n4627 VDD.n4626 25.6005
R8433 VDD.n4637 VDD.n4627 25.6005
R8434 VDD.n4637 VDD.n4636 25.6005
R8435 VDD.n4636 VDD.n4635 25.6005
R8436 VDD.n4635 VDD.n4634 25.6005
R8437 VDD.n4634 VDD.n4632 25.6005
R8438 VDD.n4632 VDD.n4631 25.6005
R8439 VDD.n4631 VDD.n4629 25.6005
R8440 VDD.n4629 VDD.n4628 25.6005
R8441 VDD.n4628 VDD.n3930 25.6005
R8442 VDD.n4384 VDD.n4126 25.6005
R8443 VDD.n4463 VDD.n4126 25.6005
R8444 VDD.n4463 VDD.n4462 25.6005
R8445 VDD.n4462 VDD.n4461 25.6005
R8446 VDD.n4461 VDD.n4460 25.6005
R8447 VDD.n4460 VDD.n4099 25.6005
R8448 VDD.n4497 VDD.n4099 25.6005
R8449 VDD.n4497 VDD.n4496 25.6005
R8450 VDD.n4496 VDD.n4495 25.6005
R8451 VDD.n4383 VDD.n4382 25.6005
R8452 VDD.n4382 VDD.n4380 25.6005
R8453 VDD.n4380 VDD.n4377 25.6005
R8454 VDD.n4377 VDD.n4376 25.6005
R8455 VDD.n4376 VDD.n4373 25.6005
R8456 VDD.n4373 VDD.n4372 25.6005
R8457 VDD.n4372 VDD.n4369 25.6005
R8458 VDD.n4369 VDD.n4368 25.6005
R8459 VDD.n4368 VDD.n4365 25.6005
R8460 VDD.n4365 VDD.n4364 25.6005
R8461 VDD.n4364 VDD.n4361 25.6005
R8462 VDD.n4361 VDD.n4360 25.6005
R8463 VDD.n4360 VDD.n4357 25.6005
R8464 VDD.n4357 VDD.n4356 25.6005
R8465 VDD.n4356 VDD.n4140 25.6005
R8466 VDD.n4426 VDD.n4140 25.6005
R8467 VDD.n4429 VDD.n4427 25.6005
R8468 VDD.n4429 VDD.n4428 25.6005
R8469 VDD.n4428 VDD.n4112 25.6005
R8470 VDD.n4474 VDD.n4112 25.6005
R8471 VDD.n4475 VDD.n4474 25.6005
R8472 VDD.n4476 VDD.n4475 25.6005
R8473 VDD.n4476 VDD.n4106 25.6005
R8474 VDD.n4486 VDD.n4106 25.6005
R8475 VDD.n4487 VDD.n4486 25.6005
R8476 VDD.n4489 VDD.n4487 25.6005
R8477 VDD.n4489 VDD.n4488 25.6005
R8478 VDD.n4488 VDD.n4061 25.6005
R8479 VDD.n4541 VDD.n4061 25.6005
R8480 VDD.n4542 VDD.n4541 25.6005
R8481 VDD.n4543 VDD.n4542 25.6005
R8482 VDD.n4545 VDD.n4543 25.6005
R8483 VDD.n4545 VDD.n4544 25.6005
R8484 VDD.n4544 VDD.n4025 25.6005
R8485 VDD.n4621 VDD.n4025 25.6005
R8486 VDD.n4622 VDD.n4621 25.6005
R8487 VDD.n4623 VDD.n4622 25.6005
R8488 VDD.n4623 VDD.n4019 25.6005
R8489 VDD.n4641 VDD.n4019 25.6005
R8490 VDD.n4642 VDD.n4641 25.6005
R8491 VDD.n4643 VDD.n4642 25.6005
R8492 VDD.n4643 VDD.n3962 25.6005
R8493 VDD.n4700 VDD.n3962 25.6005
R8494 VDD.n4701 VDD.n4700 25.6005
R8495 VDD.n4703 VDD.n4701 25.6005
R8496 VDD.n4703 VDD.n4702 25.6005
R8497 VDD.n4702 VDD.n3925 25.6005
R8498 VDD.n4735 VDD.n3925 25.6005
R8499 VDD.n4736 VDD.n4735 25.6005
R8500 VDD.n4737 VDD.n4736 25.6005
R8501 VDD.n4737 VDD.n3918 25.6005
R8502 VDD.n4749 VDD.n3918 25.6005
R8503 VDD.n4750 VDD.n4749 25.6005
R8504 VDD.n4980 VDD.n4750 25.6005
R8505 VDD.n4981 VDD.n4980 25.6005
R8506 VDD.n4982 VDD.n4981 25.6005
R8507 VDD.n4983 VDD.n4982 25.6005
R8508 VDD.n4986 VDD.n4983 25.6005
R8509 VDD.n4987 VDD.n4986 25.6005
R8510 VDD.n4988 VDD.n4987 25.6005
R8511 VDD.n4988 VDD.n3912 25.6005
R8512 VDD.n4998 VDD.n3912 25.6005
R8513 VDD.n4999 VDD.n4998 25.6005
R8514 VDD.n5028 VDD.n4999 25.6005
R8515 VDD.n5028 VDD.n5027 25.6005
R8516 VDD.n5070 VDD.n5069 25.6005
R8517 VDD.n5069 VDD.n3891 25.6005
R8518 VDD.n5000 VDD.n3891 25.6005
R8519 VDD.n5003 VDD.n5000 25.6005
R8520 VDD.n5004 VDD.n5003 25.6005
R8521 VDD.n5007 VDD.n5004 25.6005
R8522 VDD.n5008 VDD.n5007 25.6005
R8523 VDD.n5011 VDD.n5008 25.6005
R8524 VDD.n5012 VDD.n5011 25.6005
R8525 VDD.n5015 VDD.n5012 25.6005
R8526 VDD.n5016 VDD.n5015 25.6005
R8527 VDD.n5019 VDD.n5016 25.6005
R8528 VDD.n5020 VDD.n5019 25.6005
R8529 VDD.n5023 VDD.n5020 25.6005
R8530 VDD.n5025 VDD.n5023 25.6005
R8531 VDD.n5026 VDD.n5025 25.6005
R8532 VDD.n4244 VDD.n4202 25.6005
R8533 VDD.n4213 VDD.n4202 25.6005
R8534 VDD.n4214 VDD.n4213 25.6005
R8535 VDD.n4217 VDD.n4214 25.6005
R8536 VDD.n4218 VDD.n4217 25.6005
R8537 VDD.n4221 VDD.n4218 25.6005
R8538 VDD.n4222 VDD.n4221 25.6005
R8539 VDD.n4225 VDD.n4222 25.6005
R8540 VDD.n4226 VDD.n4225 25.6005
R8541 VDD.n4229 VDD.n4226 25.6005
R8542 VDD.n4230 VDD.n4229 25.6005
R8543 VDD.n4233 VDD.n4230 25.6005
R8544 VDD.n4234 VDD.n4233 25.6005
R8545 VDD.n4237 VDD.n4234 25.6005
R8546 VDD.n4238 VDD.n4237 25.6005
R8547 VDD.n4239 VDD.n4238 25.6005
R8548 VDD.n4246 VDD.n4245 25.6005
R8549 VDD.n4246 VDD.n4194 25.6005
R8550 VDD.n4256 VDD.n4194 25.6005
R8551 VDD.n4257 VDD.n4256 25.6005
R8552 VDD.n4258 VDD.n4257 25.6005
R8553 VDD.n4258 VDD.n4186 25.6005
R8554 VDD.n4269 VDD.n4186 25.6005
R8555 VDD.n4270 VDD.n4269 25.6005
R8556 VDD.n4271 VDD.n4270 25.6005
R8557 VDD.n4271 VDD.n4179 25.6005
R8558 VDD.n4282 VDD.n4179 25.6005
R8559 VDD.n4283 VDD.n4282 25.6005
R8560 VDD.n4284 VDD.n4283 25.6005
R8561 VDD.n4284 VDD.n4172 25.6005
R8562 VDD.n4294 VDD.n4172 25.6005
R8563 VDD.n4295 VDD.n4294 25.6005
R8564 VDD.n4297 VDD.n4295 25.6005
R8565 VDD.n4297 VDD.n4296 25.6005
R8566 VDD.n4296 VDD.n4163 25.6005
R8567 VDD.n4347 VDD.n4163 25.6005
R8568 VDD.n4348 VDD.n4347 25.6005
R8569 VDD.n4352 VDD.n4348 25.6005
R8570 VDD.n4352 VDD.n4351 25.6005
R8571 VDD.n5145 VDD.n5144 25.6005
R8572 VDD.n5136 VDD.n3793 25.6005
R8573 VDD.n4799 VDD.n4784 25.6005
R8574 VDD.n4803 VDD.n4784 25.6005
R8575 VDD.n4804 VDD.n4803 25.6005
R8576 VDD.n4940 VDD.n4804 25.6005
R8577 VDD.n4940 VDD.n4939 25.6005
R8578 VDD.n4939 VDD.n4938 25.6005
R8579 VDD.n4938 VDD.n4805 25.6005
R8580 VDD.n4932 VDD.n4805 25.6005
R8581 VDD.n4932 VDD.n4931 25.6005
R8582 VDD.n4931 VDD.n4930 25.6005
R8583 VDD.n4930 VDD.n4812 25.6005
R8584 VDD.n4924 VDD.n4812 25.6005
R8585 VDD.n4924 VDD.n4923 25.6005
R8586 VDD.n4923 VDD.n4922 25.6005
R8587 VDD.n4922 VDD.n4818 25.6005
R8588 VDD.n4916 VDD.n4818 25.6005
R8589 VDD.n4916 VDD.n4915 25.6005
R8590 VDD.n4915 VDD.n4914 25.6005
R8591 VDD.n4914 VDD.n4826 25.6005
R8592 VDD.n4908 VDD.n4826 25.6005
R8593 VDD.n4908 VDD.n4907 25.6005
R8594 VDD.n4907 VDD.n4906 25.6005
R8595 VDD.n4906 VDD.n4833 25.6005
R8596 VDD.n4899 VDD.n4898 25.6005
R8597 VDD.n4898 VDD.n4897 25.6005
R8598 VDD.n4897 VDD.n4896 25.6005
R8599 VDD.n4896 VDD.n4894 25.6005
R8600 VDD.n4894 VDD.n4891 25.6005
R8601 VDD.n4891 VDD.n4890 25.6005
R8602 VDD.n4890 VDD.n4887 25.6005
R8603 VDD.n4887 VDD.n4886 25.6005
R8604 VDD.n4886 VDD.n4883 25.6005
R8605 VDD.n4883 VDD.n4882 25.6005
R8606 VDD.n4882 VDD.n4879 25.6005
R8607 VDD.n4879 VDD.n4878 25.6005
R8608 VDD.n4878 VDD.n4875 25.6005
R8609 VDD.n4875 VDD.n4874 25.6005
R8610 VDD.n4874 VDD.n4871 25.6005
R8611 VDD.n4871 VDD.n4870 25.6005
R8612 VDD.n4250 VDD.n4198 25.6005
R8613 VDD.n4251 VDD.n4250 25.6005
R8614 VDD.n4252 VDD.n4251 25.6005
R8615 VDD.n4252 VDD.n4190 25.6005
R8616 VDD.n4262 VDD.n4190 25.6005
R8617 VDD.n4263 VDD.n4262 25.6005
R8618 VDD.n4264 VDD.n4263 25.6005
R8619 VDD.n4264 VDD.n4182 25.6005
R8620 VDD.n4275 VDD.n4182 25.6005
R8621 VDD.n4276 VDD.n4275 25.6005
R8622 VDD.n4277 VDD.n4276 25.6005
R8623 VDD.n4277 VDD.n4176 25.6005
R8624 VDD.n4288 VDD.n4176 25.6005
R8625 VDD.n4289 VDD.n4288 25.6005
R8626 VDD.n4290 VDD.n4289 25.6005
R8627 VDD.n4290 VDD.n4168 25.6005
R8628 VDD.n4301 VDD.n4168 25.6005
R8629 VDD.n4302 VDD.n4301 25.6005
R8630 VDD.n4342 VDD.n4302 25.6005
R8631 VDD.n4342 VDD.n4341 25.6005
R8632 VDD.n4341 VDD.n4340 25.6005
R8633 VDD.n4340 VDD.n4338 25.6005
R8634 VDD.n4338 VDD.n4337 25.6005
R8635 VDD.n5149 VDD.n3449 25.6005
R8636 VDD.n3947 VDD.n3806 25.6005
R8637 VDD.n4948 VDD.n4947 25.6005
R8638 VDD.n4947 VDD.n4946 25.6005
R8639 VDD.n4946 VDD.n4778 25.6005
R8640 VDD.n4780 VDD.n4778 25.6005
R8641 VDD.n4846 VDD.n4780 25.6005
R8642 VDD.n4847 VDD.n4846 25.6005
R8643 VDD.n4848 VDD.n4847 25.6005
R8644 VDD.n4849 VDD.n4848 25.6005
R8645 VDD.n4851 VDD.n4849 25.6005
R8646 VDD.n4852 VDD.n4851 25.6005
R8647 VDD.n4853 VDD.n4852 25.6005
R8648 VDD.n4854 VDD.n4853 25.6005
R8649 VDD.n4856 VDD.n4854 25.6005
R8650 VDD.n4857 VDD.n4856 25.6005
R8651 VDD.n4858 VDD.n4857 25.6005
R8652 VDD.n4859 VDD.n4858 25.6005
R8653 VDD.n4861 VDD.n4859 25.6005
R8654 VDD.n4862 VDD.n4861 25.6005
R8655 VDD.n4863 VDD.n4862 25.6005
R8656 VDD.n4864 VDD.n4863 25.6005
R8657 VDD.n4866 VDD.n4864 25.6005
R8658 VDD.n4867 VDD.n4866 25.6005
R8659 VDD.n4868 VDD.n4867 25.6005
R8660 VDD.n157 VDD.n152 25.6005
R8661 VDD.n79 VDD.n78 25.6005
R8662 VDD.n80 VDD.n79 25.6005
R8663 VDD.n480 VDD.n80 25.6005
R8664 VDD.n480 VDD.n479 25.6005
R8665 VDD.n479 VDD.n478 25.6005
R8666 VDD.n478 VDD.n81 25.6005
R8667 VDD.n468 VDD.n81 25.6005
R8668 VDD.n468 VDD.n467 25.6005
R8669 VDD.n467 VDD.n466 25.6005
R8670 VDD.n466 VDD.n93 25.6005
R8671 VDD.n456 VDD.n93 25.6005
R8672 VDD.n456 VDD.n455 25.6005
R8673 VDD.n455 VDD.n454 25.6005
R8674 VDD.n454 VDD.n105 25.6005
R8675 VDD.n444 VDD.n105 25.6005
R8676 VDD.n444 VDD.n443 25.6005
R8677 VDD.n443 VDD.n442 25.6005
R8678 VDD.n442 VDD.n117 25.6005
R8679 VDD.n432 VDD.n117 25.6005
R8680 VDD.n432 VDD.n431 25.6005
R8681 VDD.n431 VDD.n430 25.6005
R8682 VDD.n430 VDD.n129 25.6005
R8683 VDD.n420 VDD.n129 25.6005
R8684 VDD.n53 VDD.n52 25.6005
R8685 VDD.n72 VDD.n53 25.6005
R8686 VDD.n72 VDD.n71 25.6005
R8687 VDD.n71 VDD.n70 25.6005
R8688 VDD.n70 VDD.n55 25.6005
R8689 VDD.n65 VDD.n55 25.6005
R8690 VDD.n504 VDD.n29 25.6005
R8691 VDD.n499 VDD.n29 25.6005
R8692 VDD.n499 VDD.n498 25.6005
R8693 VDD.n498 VDD.n497 25.6005
R8694 VDD.n497 VDD.n33 25.6005
R8695 VDD.n492 VDD.n33 25.6005
R8696 VDD.n491 VDD.n490 25.6005
R8697 VDD.n490 VDD.n36 25.6005
R8698 VDD.n352 VDD.n36 25.6005
R8699 VDD.n354 VDD.n352 25.6005
R8700 VDD.n355 VDD.n354 25.6005
R8701 VDD.n357 VDD.n355 25.6005
R8702 VDD.n358 VDD.n357 25.6005
R8703 VDD.n360 VDD.n358 25.6005
R8704 VDD.n361 VDD.n360 25.6005
R8705 VDD.n363 VDD.n361 25.6005
R8706 VDD.n364 VDD.n363 25.6005
R8707 VDD.n366 VDD.n364 25.6005
R8708 VDD.n367 VDD.n366 25.6005
R8709 VDD.n369 VDD.n367 25.6005
R8710 VDD.n370 VDD.n369 25.6005
R8711 VDD.n372 VDD.n370 25.6005
R8712 VDD.n373 VDD.n372 25.6005
R8713 VDD.n375 VDD.n373 25.6005
R8714 VDD.n376 VDD.n375 25.6005
R8715 VDD.n378 VDD.n376 25.6005
R8716 VDD.n379 VDD.n378 25.6005
R8717 VDD.n381 VDD.n379 25.6005
R8718 VDD.n382 VDD.n381 25.6005
R8719 VDD.n395 VDD.n394 25.6005
R8720 VDD.n394 VDD.n350 25.6005
R8721 VDD.n389 VDD.n350 25.6005
R8722 VDD.n389 VDD.n388 25.6005
R8723 VDD.n388 VDD.n387 25.6005
R8724 VDD.n387 VDD.n383 25.6005
R8725 VDD.n419 VDD.n418 25.6005
R8726 VDD.n418 VDD.n141 25.6005
R8727 VDD.n412 VDD.n141 25.6005
R8728 VDD.n412 VDD.n411 25.6005
R8729 VDD.n411 VDD.n410 25.6005
R8730 VDD.n410 VDD.n143 25.6005
R8731 VDD.n208 VDD.n207 25.6005
R8732 VDD.n214 VDD.n207 25.6005
R8733 VDD.n215 VDD.n214 25.6005
R8734 VDD.n216 VDD.n215 25.6005
R8735 VDD.n216 VDD.n205 25.6005
R8736 VDD.n205 VDD.n204 25.6005
R8737 VDD.n486 VDD.n44 25.6005
R8738 VDD.n486 VDD.n485 25.6005
R8739 VDD.n485 VDD.n484 25.6005
R8740 VDD.n484 VDD.n45 25.6005
R8741 VDD.n474 VDD.n45 25.6005
R8742 VDD.n474 VDD.n473 25.6005
R8743 VDD.n473 VDD.n472 25.6005
R8744 VDD.n472 VDD.n86 25.6005
R8745 VDD.n462 VDD.n86 25.6005
R8746 VDD.n462 VDD.n461 25.6005
R8747 VDD.n461 VDD.n460 25.6005
R8748 VDD.n460 VDD.n98 25.6005
R8749 VDD.n450 VDD.n98 25.6005
R8750 VDD.n450 VDD.n449 25.6005
R8751 VDD.n449 VDD.n448 25.6005
R8752 VDD.n448 VDD.n110 25.6005
R8753 VDD.n438 VDD.n110 25.6005
R8754 VDD.n438 VDD.n437 25.6005
R8755 VDD.n437 VDD.n436 25.6005
R8756 VDD.n436 VDD.n122 25.6005
R8757 VDD.n426 VDD.n122 25.6005
R8758 VDD.n426 VDD.n425 25.6005
R8759 VDD.n425 VDD.n424 25.6005
R8760 VDD.n167 VDD.n135 25.6005
R8761 VDD.n168 VDD.n167 25.6005
R8762 VDD.n169 VDD.n168 25.6005
R8763 VDD.n169 VDD.n163 25.6005
R8764 VDD.n175 VDD.n163 25.6005
R8765 VDD.n176 VDD.n175 25.6005
R8766 VDD.n303 VDD.n302 25.6005
R8767 VDD.n302 VDD.n301 25.6005
R8768 VDD.n301 VDD.n182 25.6005
R8769 VDD.n295 VDD.n182 25.6005
R8770 VDD.n295 VDD.n294 25.6005
R8771 VDD.n294 VDD.n293 25.6005
R8772 VDD.n257 VDD.n256 25.6005
R8773 VDD.n259 VDD.n257 25.6005
R8774 VDD.n260 VDD.n259 25.6005
R8775 VDD.n262 VDD.n260 25.6005
R8776 VDD.n263 VDD.n262 25.6005
R8777 VDD.n265 VDD.n263 25.6005
R8778 VDD.n266 VDD.n265 25.6005
R8779 VDD.n268 VDD.n266 25.6005
R8780 VDD.n269 VDD.n268 25.6005
R8781 VDD.n271 VDD.n269 25.6005
R8782 VDD.n272 VDD.n271 25.6005
R8783 VDD.n274 VDD.n272 25.6005
R8784 VDD.n275 VDD.n274 25.6005
R8785 VDD.n277 VDD.n275 25.6005
R8786 VDD.n278 VDD.n277 25.6005
R8787 VDD.n280 VDD.n278 25.6005
R8788 VDD.n281 VDD.n280 25.6005
R8789 VDD.n283 VDD.n281 25.6005
R8790 VDD.n284 VDD.n283 25.6005
R8791 VDD.n286 VDD.n284 25.6005
R8792 VDD.n287 VDD.n286 25.6005
R8793 VDD.n289 VDD.n287 25.6005
R8794 VDD.n290 VDD.n289 25.6005
R8795 VDD.n243 VDD.n242 25.6005
R8796 VDD.n243 VDD.n186 25.6005
R8797 VDD.n249 VDD.n186 25.6005
R8798 VDD.n250 VDD.n249 25.6005
R8799 VDD.n251 VDD.n250 25.6005
R8800 VDD.n251 VDD.n184 25.6005
R8801 VDD.n237 VDD.n236 25.6005
R8802 VDD.n1839 VDD.n1542 25.6005
R8803 VDD.n1840 VDD.n1839 25.6005
R8804 VDD.n1842 VDD.n1840 25.6005
R8805 VDD.n1842 VDD.n1841 25.6005
R8806 VDD.n1841 VDD.n1514 25.6005
R8807 VDD.n1886 VDD.n1514 25.6005
R8808 VDD.n1887 VDD.n1886 25.6005
R8809 VDD.n1888 VDD.n1887 25.6005
R8810 VDD.n1888 VDD.n1506 25.6005
R8811 VDD.n1827 VDD.n1826 25.6005
R8812 VDD.n1826 VDD.n1825 25.6005
R8813 VDD.n1825 VDD.n1822 25.6005
R8814 VDD.n1822 VDD.n1821 25.6005
R8815 VDD.n1821 VDD.n1818 25.6005
R8816 VDD.n1818 VDD.n1817 25.6005
R8817 VDD.n1817 VDD.n1814 25.6005
R8818 VDD.n1814 VDD.n1813 25.6005
R8819 VDD.n1813 VDD.n1810 25.6005
R8820 VDD.n1810 VDD.n1809 25.6005
R8821 VDD.n1809 VDD.n1806 25.6005
R8822 VDD.n1806 VDD.n1805 25.6005
R8823 VDD.n1805 VDD.n1802 25.6005
R8824 VDD.n1802 VDD.n1801 25.6005
R8825 VDD.n1801 VDD.n1798 25.6005
R8826 VDD.n1798 VDD.n1797 25.6005
R8827 VDD.n1795 VDD.n1525 25.6005
R8828 VDD.n1873 VDD.n1525 25.6005
R8829 VDD.n1874 VDD.n1873 25.6005
R8830 VDD.n1876 VDD.n1874 25.6005
R8831 VDD.n1876 VDD.n1875 25.6005
R8832 VDD.n1875 VDD.n1498 25.6005
R8833 VDD.n1907 VDD.n1498 25.6005
R8834 VDD.n1908 VDD.n1907 25.6005
R8835 VDD.n1910 VDD.n1908 25.6005
R8836 VDD.n1910 VDD.n1909 25.6005
R8837 VDD.n1909 VDD.n1475 25.6005
R8838 VDD.n1940 VDD.n1475 25.6005
R8839 VDD.n2075 VDD.n2074 25.6005
R8840 VDD.n2518 VDD.n2517 25.6005
R8841 VDD.n2517 VDD.n2516 25.6005
R8842 VDD.n2516 VDD.n1230 25.6005
R8843 VDD.n1269 VDD.n1230 25.6005
R8844 VDD.n1270 VDD.n1269 25.6005
R8845 VDD.n2495 VDD.n1270 25.6005
R8846 VDD.n2495 VDD.n2494 25.6005
R8847 VDD.n2494 VDD.n2493 25.6005
R8848 VDD.n2493 VDD.n1271 25.6005
R8849 VDD.n2483 VDD.n1271 25.6005
R8850 VDD.n2483 VDD.n2482 25.6005
R8851 VDD.n2482 VDD.n2481 25.6005
R8852 VDD.n2469 VDD.n1290 25.6005
R8853 VDD.n2469 VDD.n2468 25.6005
R8854 VDD.n2468 VDD.n2467 25.6005
R8855 VDD.n2467 VDD.n2465 25.6005
R8856 VDD.n2465 VDD.n2462 25.6005
R8857 VDD.n2462 VDD.n2461 25.6005
R8858 VDD.n2461 VDD.n2458 25.6005
R8859 VDD.n2458 VDD.n2457 25.6005
R8860 VDD.n2457 VDD.n2454 25.6005
R8861 VDD.n2454 VDD.n2453 25.6005
R8862 VDD.n2453 VDD.n2450 25.6005
R8863 VDD.n2450 VDD.n2449 25.6005
R8864 VDD.n2449 VDD.n2446 25.6005
R8865 VDD.n2446 VDD.n2445 25.6005
R8866 VDD.n2445 VDD.n2442 25.6005
R8867 VDD.n2442 VDD.n2441 25.6005
R8868 VDD.n1278 VDD.n1238 25.6005
R8869 VDD.n1281 VDD.n1278 25.6005
R8870 VDD.n1282 VDD.n1281 25.6005
R8871 VDD.n1283 VDD.n1282 25.6005
R8872 VDD.n2489 VDD.n1283 25.6005
R8873 VDD.n2489 VDD.n2488 25.6005
R8874 VDD.n2488 VDD.n2487 25.6005
R8875 VDD.n2487 VDD.n1284 25.6005
R8876 VDD.n2477 VDD.n1284 25.6005
R8877 VDD.n2510 VDD.n1239 25.6005
R8878 VDD.n1321 VDD.n1239 25.6005
R8879 VDD.n1322 VDD.n1321 25.6005
R8880 VDD.n2398 VDD.n1322 25.6005
R8881 VDD.n2399 VDD.n2398 25.6005
R8882 VDD.n2400 VDD.n2399 25.6005
R8883 VDD.n2400 VDD.n1316 25.6005
R8884 VDD.n2438 VDD.n1316 25.6005
R8885 VDD.n2439 VDD.n2438 25.6005
R8886 VDD.n1990 VDD.n1989 25.6005
R8887 VDD.n1989 VDD.n1988 25.6005
R8888 VDD.n1988 VDD.n1417 25.6005
R8889 VDD.n2056 VDD.n1417 25.6005
R8890 VDD.n2056 VDD.n2055 25.6005
R8891 VDD.n2055 VDD.n2054 25.6005
R8892 VDD.n2054 VDD.n2053 25.6005
R8893 VDD.n2053 VDD.n1421 25.6005
R8894 VDD.n1421 VDD.n1420 25.6005
R8895 VDD.n1420 VDD.n1419 25.6005
R8896 VDD.n1419 VDD.n1337 25.6005
R8897 VDD.n2133 VDD.n1337 25.6005
R8898 VDD.n2134 VDD.n2133 25.6005
R8899 VDD.n1460 VDD.n1459 25.6005
R8900 VDD.n1459 VDD.n1427 25.6005
R8901 VDD.n2032 VDD.n1427 25.6005
R8902 VDD.n2033 VDD.n2032 25.6005
R8903 VDD.n2043 VDD.n2033 25.6005
R8904 VDD.n2043 VDD.n2042 25.6005
R8905 VDD.n2042 VDD.n2041 25.6005
R8906 VDD.n2041 VDD.n2040 25.6005
R8907 VDD.n2040 VDD.n2038 25.6005
R8908 VDD.n2038 VDD.n2037 25.6005
R8909 VDD.n2037 VDD.n2035 25.6005
R8910 VDD.n2035 VDD.n2034 25.6005
R8911 VDD.n2034 VDD.n1336 25.6005
R8912 VDD.n1790 VDD.n1532 25.6005
R8913 VDD.n1869 VDD.n1532 25.6005
R8914 VDD.n1869 VDD.n1868 25.6005
R8915 VDD.n1868 VDD.n1867 25.6005
R8916 VDD.n1867 VDD.n1866 25.6005
R8917 VDD.n1866 VDD.n1505 25.6005
R8918 VDD.n1903 VDD.n1505 25.6005
R8919 VDD.n1903 VDD.n1902 25.6005
R8920 VDD.n1902 VDD.n1901 25.6005
R8921 VDD.n1789 VDD.n1788 25.6005
R8922 VDD.n1788 VDD.n1786 25.6005
R8923 VDD.n1786 VDD.n1783 25.6005
R8924 VDD.n1783 VDD.n1782 25.6005
R8925 VDD.n1782 VDD.n1779 25.6005
R8926 VDD.n1779 VDD.n1778 25.6005
R8927 VDD.n1778 VDD.n1775 25.6005
R8928 VDD.n1775 VDD.n1774 25.6005
R8929 VDD.n1774 VDD.n1771 25.6005
R8930 VDD.n1771 VDD.n1770 25.6005
R8931 VDD.n1770 VDD.n1767 25.6005
R8932 VDD.n1767 VDD.n1766 25.6005
R8933 VDD.n1766 VDD.n1763 25.6005
R8934 VDD.n1763 VDD.n1762 25.6005
R8935 VDD.n1762 VDD.n1546 25.6005
R8936 VDD.n1832 VDD.n1546 25.6005
R8937 VDD.n1835 VDD.n1833 25.6005
R8938 VDD.n1835 VDD.n1834 25.6005
R8939 VDD.n1834 VDD.n1518 25.6005
R8940 VDD.n1880 VDD.n1518 25.6005
R8941 VDD.n1881 VDD.n1880 25.6005
R8942 VDD.n1882 VDD.n1881 25.6005
R8943 VDD.n1882 VDD.n1512 25.6005
R8944 VDD.n1892 VDD.n1512 25.6005
R8945 VDD.n1893 VDD.n1892 25.6005
R8946 VDD.n1895 VDD.n1893 25.6005
R8947 VDD.n1895 VDD.n1894 25.6005
R8948 VDD.n1894 VDD.n1467 25.6005
R8949 VDD.n1947 VDD.n1467 25.6005
R8950 VDD.n1948 VDD.n1947 25.6005
R8951 VDD.n1949 VDD.n1948 25.6005
R8952 VDD.n1951 VDD.n1949 25.6005
R8953 VDD.n1951 VDD.n1950 25.6005
R8954 VDD.n1950 VDD.n1431 25.6005
R8955 VDD.n2027 VDD.n1431 25.6005
R8956 VDD.n2028 VDD.n2027 25.6005
R8957 VDD.n2029 VDD.n2028 25.6005
R8958 VDD.n2029 VDD.n1425 25.6005
R8959 VDD.n2047 VDD.n1425 25.6005
R8960 VDD.n2048 VDD.n2047 25.6005
R8961 VDD.n2049 VDD.n2048 25.6005
R8962 VDD.n2049 VDD.n1368 25.6005
R8963 VDD.n2106 VDD.n1368 25.6005
R8964 VDD.n2107 VDD.n2106 25.6005
R8965 VDD.n2109 VDD.n2107 25.6005
R8966 VDD.n2109 VDD.n2108 25.6005
R8967 VDD.n2108 VDD.n1331 25.6005
R8968 VDD.n2141 VDD.n1331 25.6005
R8969 VDD.n2142 VDD.n2141 25.6005
R8970 VDD.n2143 VDD.n2142 25.6005
R8971 VDD.n2143 VDD.n1324 25.6005
R8972 VDD.n2155 VDD.n1324 25.6005
R8973 VDD.n2156 VDD.n2155 25.6005
R8974 VDD.n2386 VDD.n2156 25.6005
R8975 VDD.n2387 VDD.n2386 25.6005
R8976 VDD.n2388 VDD.n2387 25.6005
R8977 VDD.n2389 VDD.n2388 25.6005
R8978 VDD.n2392 VDD.n2389 25.6005
R8979 VDD.n2393 VDD.n2392 25.6005
R8980 VDD.n2394 VDD.n2393 25.6005
R8981 VDD.n2394 VDD.n1318 25.6005
R8982 VDD.n2404 VDD.n1318 25.6005
R8983 VDD.n2405 VDD.n2404 25.6005
R8984 VDD.n2434 VDD.n2405 25.6005
R8985 VDD.n2434 VDD.n2433 25.6005
R8986 VDD.n2476 VDD.n2475 25.6005
R8987 VDD.n2475 VDD.n1297 25.6005
R8988 VDD.n2406 VDD.n1297 25.6005
R8989 VDD.n2409 VDD.n2406 25.6005
R8990 VDD.n2410 VDD.n2409 25.6005
R8991 VDD.n2413 VDD.n2410 25.6005
R8992 VDD.n2414 VDD.n2413 25.6005
R8993 VDD.n2417 VDD.n2414 25.6005
R8994 VDD.n2418 VDD.n2417 25.6005
R8995 VDD.n2421 VDD.n2418 25.6005
R8996 VDD.n2422 VDD.n2421 25.6005
R8997 VDD.n2425 VDD.n2422 25.6005
R8998 VDD.n2426 VDD.n2425 25.6005
R8999 VDD.n2429 VDD.n2426 25.6005
R9000 VDD.n2431 VDD.n2429 25.6005
R9001 VDD.n2432 VDD.n2431 25.6005
R9002 VDD.n1650 VDD.n1608 25.6005
R9003 VDD.n1619 VDD.n1608 25.6005
R9004 VDD.n1620 VDD.n1619 25.6005
R9005 VDD.n1623 VDD.n1620 25.6005
R9006 VDD.n1624 VDD.n1623 25.6005
R9007 VDD.n1627 VDD.n1624 25.6005
R9008 VDD.n1628 VDD.n1627 25.6005
R9009 VDD.n1631 VDD.n1628 25.6005
R9010 VDD.n1632 VDD.n1631 25.6005
R9011 VDD.n1635 VDD.n1632 25.6005
R9012 VDD.n1636 VDD.n1635 25.6005
R9013 VDD.n1639 VDD.n1636 25.6005
R9014 VDD.n1640 VDD.n1639 25.6005
R9015 VDD.n1643 VDD.n1640 25.6005
R9016 VDD.n1644 VDD.n1643 25.6005
R9017 VDD.n1645 VDD.n1644 25.6005
R9018 VDD.n1652 VDD.n1651 25.6005
R9019 VDD.n1652 VDD.n1600 25.6005
R9020 VDD.n1662 VDD.n1600 25.6005
R9021 VDD.n1663 VDD.n1662 25.6005
R9022 VDD.n1664 VDD.n1663 25.6005
R9023 VDD.n1664 VDD.n1592 25.6005
R9024 VDD.n1675 VDD.n1592 25.6005
R9025 VDD.n1676 VDD.n1675 25.6005
R9026 VDD.n1677 VDD.n1676 25.6005
R9027 VDD.n1677 VDD.n1585 25.6005
R9028 VDD.n1688 VDD.n1585 25.6005
R9029 VDD.n1689 VDD.n1688 25.6005
R9030 VDD.n1690 VDD.n1689 25.6005
R9031 VDD.n1690 VDD.n1578 25.6005
R9032 VDD.n1700 VDD.n1578 25.6005
R9033 VDD.n1701 VDD.n1700 25.6005
R9034 VDD.n1703 VDD.n1701 25.6005
R9035 VDD.n1703 VDD.n1702 25.6005
R9036 VDD.n1702 VDD.n1569 25.6005
R9037 VDD.n1753 VDD.n1569 25.6005
R9038 VDD.n1754 VDD.n1753 25.6005
R9039 VDD.n1758 VDD.n1754 25.6005
R9040 VDD.n1758 VDD.n1757 25.6005
R9041 VDD.n2551 VDD.n2550 25.6005
R9042 VDD.n2542 VDD.n1199 25.6005
R9043 VDD.n2205 VDD.n2190 25.6005
R9044 VDD.n2209 VDD.n2190 25.6005
R9045 VDD.n2210 VDD.n2209 25.6005
R9046 VDD.n2346 VDD.n2210 25.6005
R9047 VDD.n2346 VDD.n2345 25.6005
R9048 VDD.n2345 VDD.n2344 25.6005
R9049 VDD.n2344 VDD.n2211 25.6005
R9050 VDD.n2338 VDD.n2211 25.6005
R9051 VDD.n2338 VDD.n2337 25.6005
R9052 VDD.n2337 VDD.n2336 25.6005
R9053 VDD.n2336 VDD.n2218 25.6005
R9054 VDD.n2330 VDD.n2218 25.6005
R9055 VDD.n2330 VDD.n2329 25.6005
R9056 VDD.n2329 VDD.n2328 25.6005
R9057 VDD.n2328 VDD.n2224 25.6005
R9058 VDD.n2322 VDD.n2224 25.6005
R9059 VDD.n2322 VDD.n2321 25.6005
R9060 VDD.n2321 VDD.n2320 25.6005
R9061 VDD.n2320 VDD.n2232 25.6005
R9062 VDD.n2314 VDD.n2232 25.6005
R9063 VDD.n2314 VDD.n2313 25.6005
R9064 VDD.n2313 VDD.n2312 25.6005
R9065 VDD.n2312 VDD.n2239 25.6005
R9066 VDD.n2305 VDD.n2304 25.6005
R9067 VDD.n2304 VDD.n2303 25.6005
R9068 VDD.n2303 VDD.n2302 25.6005
R9069 VDD.n2302 VDD.n2300 25.6005
R9070 VDD.n2300 VDD.n2297 25.6005
R9071 VDD.n2297 VDD.n2296 25.6005
R9072 VDD.n2296 VDD.n2293 25.6005
R9073 VDD.n2293 VDD.n2292 25.6005
R9074 VDD.n2292 VDD.n2289 25.6005
R9075 VDD.n2289 VDD.n2288 25.6005
R9076 VDD.n2288 VDD.n2285 25.6005
R9077 VDD.n2285 VDD.n2284 25.6005
R9078 VDD.n2284 VDD.n2281 25.6005
R9079 VDD.n2281 VDD.n2280 25.6005
R9080 VDD.n2280 VDD.n2277 25.6005
R9081 VDD.n2277 VDD.n2276 25.6005
R9082 VDD.n1656 VDD.n1604 25.6005
R9083 VDD.n1657 VDD.n1656 25.6005
R9084 VDD.n1658 VDD.n1657 25.6005
R9085 VDD.n1658 VDD.n1596 25.6005
R9086 VDD.n1668 VDD.n1596 25.6005
R9087 VDD.n1669 VDD.n1668 25.6005
R9088 VDD.n1670 VDD.n1669 25.6005
R9089 VDD.n1670 VDD.n1588 25.6005
R9090 VDD.n1681 VDD.n1588 25.6005
R9091 VDD.n1682 VDD.n1681 25.6005
R9092 VDD.n1683 VDD.n1682 25.6005
R9093 VDD.n1683 VDD.n1582 25.6005
R9094 VDD.n1694 VDD.n1582 25.6005
R9095 VDD.n1695 VDD.n1694 25.6005
R9096 VDD.n1696 VDD.n1695 25.6005
R9097 VDD.n1696 VDD.n1574 25.6005
R9098 VDD.n1707 VDD.n1574 25.6005
R9099 VDD.n1708 VDD.n1707 25.6005
R9100 VDD.n1748 VDD.n1708 25.6005
R9101 VDD.n1748 VDD.n1747 25.6005
R9102 VDD.n1747 VDD.n1746 25.6005
R9103 VDD.n1746 VDD.n1744 25.6005
R9104 VDD.n1744 VDD.n1743 25.6005
R9105 VDD.n2555 VDD.n855 25.6005
R9106 VDD.n1353 VDD.n1212 25.6005
R9107 VDD.n2354 VDD.n2353 25.6005
R9108 VDD.n2353 VDD.n2352 25.6005
R9109 VDD.n2352 VDD.n2184 25.6005
R9110 VDD.n2186 VDD.n2184 25.6005
R9111 VDD.n2252 VDD.n2186 25.6005
R9112 VDD.n2253 VDD.n2252 25.6005
R9113 VDD.n2254 VDD.n2253 25.6005
R9114 VDD.n2255 VDD.n2254 25.6005
R9115 VDD.n2257 VDD.n2255 25.6005
R9116 VDD.n2258 VDD.n2257 25.6005
R9117 VDD.n2259 VDD.n2258 25.6005
R9118 VDD.n2260 VDD.n2259 25.6005
R9119 VDD.n2262 VDD.n2260 25.6005
R9120 VDD.n2263 VDD.n2262 25.6005
R9121 VDD.n2264 VDD.n2263 25.6005
R9122 VDD.n2265 VDD.n2264 25.6005
R9123 VDD.n2267 VDD.n2265 25.6005
R9124 VDD.n2268 VDD.n2267 25.6005
R9125 VDD.n2269 VDD.n2268 25.6005
R9126 VDD.n2270 VDD.n2269 25.6005
R9127 VDD.n2272 VDD.n2270 25.6005
R9128 VDD.n2273 VDD.n2272 25.6005
R9129 VDD.n2274 VDD.n2273 25.6005
R9130 VDD.n5720 VDD.n5715 25.6005
R9131 VDD.n5642 VDD.n5641 25.6005
R9132 VDD.n5643 VDD.n5642 25.6005
R9133 VDD.n6043 VDD.n5643 25.6005
R9134 VDD.n6043 VDD.n6042 25.6005
R9135 VDD.n6042 VDD.n6041 25.6005
R9136 VDD.n6041 VDD.n5644 25.6005
R9137 VDD.n6031 VDD.n5644 25.6005
R9138 VDD.n6031 VDD.n6030 25.6005
R9139 VDD.n6030 VDD.n6029 25.6005
R9140 VDD.n6029 VDD.n5656 25.6005
R9141 VDD.n6019 VDD.n5656 25.6005
R9142 VDD.n6019 VDD.n6018 25.6005
R9143 VDD.n6018 VDD.n6017 25.6005
R9144 VDD.n6017 VDD.n5668 25.6005
R9145 VDD.n6007 VDD.n5668 25.6005
R9146 VDD.n6007 VDD.n6006 25.6005
R9147 VDD.n6006 VDD.n6005 25.6005
R9148 VDD.n6005 VDD.n5680 25.6005
R9149 VDD.n5995 VDD.n5680 25.6005
R9150 VDD.n5995 VDD.n5994 25.6005
R9151 VDD.n5994 VDD.n5993 25.6005
R9152 VDD.n5993 VDD.n5692 25.6005
R9153 VDD.n5983 VDD.n5692 25.6005
R9154 VDD.n5616 VDD.n5615 25.6005
R9155 VDD.n5635 VDD.n5616 25.6005
R9156 VDD.n5635 VDD.n5634 25.6005
R9157 VDD.n5634 VDD.n5633 25.6005
R9158 VDD.n5633 VDD.n5618 25.6005
R9159 VDD.n5628 VDD.n5618 25.6005
R9160 VDD.n6067 VDD.n5592 25.6005
R9161 VDD.n6062 VDD.n5592 25.6005
R9162 VDD.n6062 VDD.n6061 25.6005
R9163 VDD.n6061 VDD.n6060 25.6005
R9164 VDD.n6060 VDD.n5596 25.6005
R9165 VDD.n6055 VDD.n5596 25.6005
R9166 VDD.n6054 VDD.n6053 25.6005
R9167 VDD.n6053 VDD.n5599 25.6005
R9168 VDD.n5915 VDD.n5599 25.6005
R9169 VDD.n5917 VDD.n5915 25.6005
R9170 VDD.n5918 VDD.n5917 25.6005
R9171 VDD.n5920 VDD.n5918 25.6005
R9172 VDD.n5921 VDD.n5920 25.6005
R9173 VDD.n5923 VDD.n5921 25.6005
R9174 VDD.n5924 VDD.n5923 25.6005
R9175 VDD.n5926 VDD.n5924 25.6005
R9176 VDD.n5927 VDD.n5926 25.6005
R9177 VDD.n5929 VDD.n5927 25.6005
R9178 VDD.n5930 VDD.n5929 25.6005
R9179 VDD.n5932 VDD.n5930 25.6005
R9180 VDD.n5933 VDD.n5932 25.6005
R9181 VDD.n5935 VDD.n5933 25.6005
R9182 VDD.n5936 VDD.n5935 25.6005
R9183 VDD.n5938 VDD.n5936 25.6005
R9184 VDD.n5939 VDD.n5938 25.6005
R9185 VDD.n5941 VDD.n5939 25.6005
R9186 VDD.n5942 VDD.n5941 25.6005
R9187 VDD.n5944 VDD.n5942 25.6005
R9188 VDD.n5945 VDD.n5944 25.6005
R9189 VDD.n5958 VDD.n5957 25.6005
R9190 VDD.n5957 VDD.n5913 25.6005
R9191 VDD.n5952 VDD.n5913 25.6005
R9192 VDD.n5952 VDD.n5951 25.6005
R9193 VDD.n5951 VDD.n5950 25.6005
R9194 VDD.n5950 VDD.n5946 25.6005
R9195 VDD.n5982 VDD.n5981 25.6005
R9196 VDD.n5981 VDD.n5704 25.6005
R9197 VDD.n5975 VDD.n5704 25.6005
R9198 VDD.n5975 VDD.n5974 25.6005
R9199 VDD.n5974 VDD.n5973 25.6005
R9200 VDD.n5973 VDD.n5706 25.6005
R9201 VDD.n5771 VDD.n5770 25.6005
R9202 VDD.n5777 VDD.n5770 25.6005
R9203 VDD.n5778 VDD.n5777 25.6005
R9204 VDD.n5779 VDD.n5778 25.6005
R9205 VDD.n5779 VDD.n5768 25.6005
R9206 VDD.n5768 VDD.n5767 25.6005
R9207 VDD.n6049 VDD.n5607 25.6005
R9208 VDD.n6049 VDD.n6048 25.6005
R9209 VDD.n6048 VDD.n6047 25.6005
R9210 VDD.n6047 VDD.n5608 25.6005
R9211 VDD.n6037 VDD.n5608 25.6005
R9212 VDD.n6037 VDD.n6036 25.6005
R9213 VDD.n6036 VDD.n6035 25.6005
R9214 VDD.n6035 VDD.n5649 25.6005
R9215 VDD.n6025 VDD.n5649 25.6005
R9216 VDD.n6025 VDD.n6024 25.6005
R9217 VDD.n6024 VDD.n6023 25.6005
R9218 VDD.n6023 VDD.n5661 25.6005
R9219 VDD.n6013 VDD.n5661 25.6005
R9220 VDD.n6013 VDD.n6012 25.6005
R9221 VDD.n6012 VDD.n6011 25.6005
R9222 VDD.n6011 VDD.n5673 25.6005
R9223 VDD.n6001 VDD.n5673 25.6005
R9224 VDD.n6001 VDD.n6000 25.6005
R9225 VDD.n6000 VDD.n5999 25.6005
R9226 VDD.n5999 VDD.n5685 25.6005
R9227 VDD.n5989 VDD.n5685 25.6005
R9228 VDD.n5989 VDD.n5988 25.6005
R9229 VDD.n5988 VDD.n5987 25.6005
R9230 VDD.n5730 VDD.n5698 25.6005
R9231 VDD.n5731 VDD.n5730 25.6005
R9232 VDD.n5732 VDD.n5731 25.6005
R9233 VDD.n5732 VDD.n5726 25.6005
R9234 VDD.n5738 VDD.n5726 25.6005
R9235 VDD.n5739 VDD.n5738 25.6005
R9236 VDD.n5866 VDD.n5865 25.6005
R9237 VDD.n5865 VDD.n5864 25.6005
R9238 VDD.n5864 VDD.n5745 25.6005
R9239 VDD.n5858 VDD.n5745 25.6005
R9240 VDD.n5858 VDD.n5857 25.6005
R9241 VDD.n5857 VDD.n5856 25.6005
R9242 VDD.n5820 VDD.n5819 25.6005
R9243 VDD.n5822 VDD.n5820 25.6005
R9244 VDD.n5823 VDD.n5822 25.6005
R9245 VDD.n5825 VDD.n5823 25.6005
R9246 VDD.n5826 VDD.n5825 25.6005
R9247 VDD.n5828 VDD.n5826 25.6005
R9248 VDD.n5829 VDD.n5828 25.6005
R9249 VDD.n5831 VDD.n5829 25.6005
R9250 VDD.n5832 VDD.n5831 25.6005
R9251 VDD.n5834 VDD.n5832 25.6005
R9252 VDD.n5835 VDD.n5834 25.6005
R9253 VDD.n5837 VDD.n5835 25.6005
R9254 VDD.n5838 VDD.n5837 25.6005
R9255 VDD.n5840 VDD.n5838 25.6005
R9256 VDD.n5841 VDD.n5840 25.6005
R9257 VDD.n5843 VDD.n5841 25.6005
R9258 VDD.n5844 VDD.n5843 25.6005
R9259 VDD.n5846 VDD.n5844 25.6005
R9260 VDD.n5847 VDD.n5846 25.6005
R9261 VDD.n5849 VDD.n5847 25.6005
R9262 VDD.n5850 VDD.n5849 25.6005
R9263 VDD.n5852 VDD.n5850 25.6005
R9264 VDD.n5853 VDD.n5852 25.6005
R9265 VDD.n5806 VDD.n5805 25.6005
R9266 VDD.n5806 VDD.n5749 25.6005
R9267 VDD.n5812 VDD.n5749 25.6005
R9268 VDD.n5813 VDD.n5812 25.6005
R9269 VDD.n5814 VDD.n5813 25.6005
R9270 VDD.n5814 VDD.n5747 25.6005
R9271 VDD.n5800 VDD.n5799 25.6005
R9272 VDD.n7402 VDD.n7105 25.6005
R9273 VDD.n7403 VDD.n7402 25.6005
R9274 VDD.n7405 VDD.n7403 25.6005
R9275 VDD.n7405 VDD.n7404 25.6005
R9276 VDD.n7404 VDD.n7077 25.6005
R9277 VDD.n7449 VDD.n7077 25.6005
R9278 VDD.n7450 VDD.n7449 25.6005
R9279 VDD.n7451 VDD.n7450 25.6005
R9280 VDD.n7451 VDD.n7069 25.6005
R9281 VDD.n7390 VDD.n7389 25.6005
R9282 VDD.n7389 VDD.n7388 25.6005
R9283 VDD.n7388 VDD.n7385 25.6005
R9284 VDD.n7385 VDD.n7384 25.6005
R9285 VDD.n7384 VDD.n7381 25.6005
R9286 VDD.n7381 VDD.n7380 25.6005
R9287 VDD.n7380 VDD.n7377 25.6005
R9288 VDD.n7377 VDD.n7376 25.6005
R9289 VDD.n7376 VDD.n7373 25.6005
R9290 VDD.n7373 VDD.n7372 25.6005
R9291 VDD.n7372 VDD.n7369 25.6005
R9292 VDD.n7369 VDD.n7368 25.6005
R9293 VDD.n7368 VDD.n7365 25.6005
R9294 VDD.n7365 VDD.n7364 25.6005
R9295 VDD.n7364 VDD.n7361 25.6005
R9296 VDD.n7361 VDD.n7360 25.6005
R9297 VDD.n7358 VDD.n7088 25.6005
R9298 VDD.n7436 VDD.n7088 25.6005
R9299 VDD.n7437 VDD.n7436 25.6005
R9300 VDD.n7439 VDD.n7437 25.6005
R9301 VDD.n7439 VDD.n7438 25.6005
R9302 VDD.n7438 VDD.n7061 25.6005
R9303 VDD.n7470 VDD.n7061 25.6005
R9304 VDD.n7471 VDD.n7470 25.6005
R9305 VDD.n7473 VDD.n7471 25.6005
R9306 VDD.n7473 VDD.n7472 25.6005
R9307 VDD.n7472 VDD.n7038 25.6005
R9308 VDD.n7503 VDD.n7038 25.6005
R9309 VDD.n7638 VDD.n7637 25.6005
R9310 VDD.n8081 VDD.n8080 25.6005
R9311 VDD.n8080 VDD.n8079 25.6005
R9312 VDD.n8079 VDD.n6793 25.6005
R9313 VDD.n6832 VDD.n6793 25.6005
R9314 VDD.n6833 VDD.n6832 25.6005
R9315 VDD.n8058 VDD.n6833 25.6005
R9316 VDD.n8058 VDD.n8057 25.6005
R9317 VDD.n8057 VDD.n8056 25.6005
R9318 VDD.n8056 VDD.n6834 25.6005
R9319 VDD.n8046 VDD.n6834 25.6005
R9320 VDD.n8046 VDD.n8045 25.6005
R9321 VDD.n8045 VDD.n8044 25.6005
R9322 VDD.n8032 VDD.n6853 25.6005
R9323 VDD.n8032 VDD.n8031 25.6005
R9324 VDD.n8031 VDD.n8030 25.6005
R9325 VDD.n8030 VDD.n8028 25.6005
R9326 VDD.n8028 VDD.n8025 25.6005
R9327 VDD.n8025 VDD.n8024 25.6005
R9328 VDD.n8024 VDD.n8021 25.6005
R9329 VDD.n8021 VDD.n8020 25.6005
R9330 VDD.n8020 VDD.n8017 25.6005
R9331 VDD.n8017 VDD.n8016 25.6005
R9332 VDD.n8016 VDD.n8013 25.6005
R9333 VDD.n8013 VDD.n8012 25.6005
R9334 VDD.n8012 VDD.n8009 25.6005
R9335 VDD.n8009 VDD.n8008 25.6005
R9336 VDD.n8008 VDD.n8005 25.6005
R9337 VDD.n8005 VDD.n8004 25.6005
R9338 VDD.n6841 VDD.n6801 25.6005
R9339 VDD.n6844 VDD.n6841 25.6005
R9340 VDD.n6845 VDD.n6844 25.6005
R9341 VDD.n6846 VDD.n6845 25.6005
R9342 VDD.n8052 VDD.n6846 25.6005
R9343 VDD.n8052 VDD.n8051 25.6005
R9344 VDD.n8051 VDD.n8050 25.6005
R9345 VDD.n8050 VDD.n6847 25.6005
R9346 VDD.n8040 VDD.n6847 25.6005
R9347 VDD.n8073 VDD.n6802 25.6005
R9348 VDD.n6884 VDD.n6802 25.6005
R9349 VDD.n6885 VDD.n6884 25.6005
R9350 VDD.n7961 VDD.n6885 25.6005
R9351 VDD.n7962 VDD.n7961 25.6005
R9352 VDD.n7963 VDD.n7962 25.6005
R9353 VDD.n7963 VDD.n6879 25.6005
R9354 VDD.n8001 VDD.n6879 25.6005
R9355 VDD.n8002 VDD.n8001 25.6005
R9356 VDD.n7553 VDD.n7552 25.6005
R9357 VDD.n7552 VDD.n7551 25.6005
R9358 VDD.n7551 VDD.n6980 25.6005
R9359 VDD.n7619 VDD.n6980 25.6005
R9360 VDD.n7619 VDD.n7618 25.6005
R9361 VDD.n7618 VDD.n7617 25.6005
R9362 VDD.n7617 VDD.n7616 25.6005
R9363 VDD.n7616 VDD.n6984 25.6005
R9364 VDD.n6984 VDD.n6983 25.6005
R9365 VDD.n6983 VDD.n6982 25.6005
R9366 VDD.n6982 VDD.n6900 25.6005
R9367 VDD.n7696 VDD.n6900 25.6005
R9368 VDD.n7697 VDD.n7696 25.6005
R9369 VDD.n7023 VDD.n7022 25.6005
R9370 VDD.n7022 VDD.n6990 25.6005
R9371 VDD.n7595 VDD.n6990 25.6005
R9372 VDD.n7596 VDD.n7595 25.6005
R9373 VDD.n7606 VDD.n7596 25.6005
R9374 VDD.n7606 VDD.n7605 25.6005
R9375 VDD.n7605 VDD.n7604 25.6005
R9376 VDD.n7604 VDD.n7603 25.6005
R9377 VDD.n7603 VDD.n7601 25.6005
R9378 VDD.n7601 VDD.n7600 25.6005
R9379 VDD.n7600 VDD.n7598 25.6005
R9380 VDD.n7598 VDD.n7597 25.6005
R9381 VDD.n7597 VDD.n6899 25.6005
R9382 VDD.n7353 VDD.n7095 25.6005
R9383 VDD.n7432 VDD.n7095 25.6005
R9384 VDD.n7432 VDD.n7431 25.6005
R9385 VDD.n7431 VDD.n7430 25.6005
R9386 VDD.n7430 VDD.n7429 25.6005
R9387 VDD.n7429 VDD.n7068 25.6005
R9388 VDD.n7466 VDD.n7068 25.6005
R9389 VDD.n7466 VDD.n7465 25.6005
R9390 VDD.n7465 VDD.n7464 25.6005
R9391 VDD.n7352 VDD.n7351 25.6005
R9392 VDD.n7351 VDD.n7349 25.6005
R9393 VDD.n7349 VDD.n7346 25.6005
R9394 VDD.n7346 VDD.n7345 25.6005
R9395 VDD.n7345 VDD.n7342 25.6005
R9396 VDD.n7342 VDD.n7341 25.6005
R9397 VDD.n7341 VDD.n7338 25.6005
R9398 VDD.n7338 VDD.n7337 25.6005
R9399 VDD.n7337 VDD.n7334 25.6005
R9400 VDD.n7334 VDD.n7333 25.6005
R9401 VDD.n7333 VDD.n7330 25.6005
R9402 VDD.n7330 VDD.n7329 25.6005
R9403 VDD.n7329 VDD.n7326 25.6005
R9404 VDD.n7326 VDD.n7325 25.6005
R9405 VDD.n7325 VDD.n7109 25.6005
R9406 VDD.n7395 VDD.n7109 25.6005
R9407 VDD.n7398 VDD.n7396 25.6005
R9408 VDD.n7398 VDD.n7397 25.6005
R9409 VDD.n7397 VDD.n7081 25.6005
R9410 VDD.n7443 VDD.n7081 25.6005
R9411 VDD.n7444 VDD.n7443 25.6005
R9412 VDD.n7445 VDD.n7444 25.6005
R9413 VDD.n7445 VDD.n7075 25.6005
R9414 VDD.n7455 VDD.n7075 25.6005
R9415 VDD.n7456 VDD.n7455 25.6005
R9416 VDD.n7458 VDD.n7456 25.6005
R9417 VDD.n7458 VDD.n7457 25.6005
R9418 VDD.n7457 VDD.n7030 25.6005
R9419 VDD.n7510 VDD.n7030 25.6005
R9420 VDD.n7511 VDD.n7510 25.6005
R9421 VDD.n7512 VDD.n7511 25.6005
R9422 VDD.n7514 VDD.n7512 25.6005
R9423 VDD.n7514 VDD.n7513 25.6005
R9424 VDD.n7513 VDD.n6994 25.6005
R9425 VDD.n7590 VDD.n6994 25.6005
R9426 VDD.n7591 VDD.n7590 25.6005
R9427 VDD.n7592 VDD.n7591 25.6005
R9428 VDD.n7592 VDD.n6988 25.6005
R9429 VDD.n7610 VDD.n6988 25.6005
R9430 VDD.n7611 VDD.n7610 25.6005
R9431 VDD.n7612 VDD.n7611 25.6005
R9432 VDD.n7612 VDD.n6931 25.6005
R9433 VDD.n7669 VDD.n6931 25.6005
R9434 VDD.n7670 VDD.n7669 25.6005
R9435 VDD.n7672 VDD.n7670 25.6005
R9436 VDD.n7672 VDD.n7671 25.6005
R9437 VDD.n7671 VDD.n6894 25.6005
R9438 VDD.n7704 VDD.n6894 25.6005
R9439 VDD.n7705 VDD.n7704 25.6005
R9440 VDD.n7706 VDD.n7705 25.6005
R9441 VDD.n7706 VDD.n6887 25.6005
R9442 VDD.n7718 VDD.n6887 25.6005
R9443 VDD.n7719 VDD.n7718 25.6005
R9444 VDD.n7949 VDD.n7719 25.6005
R9445 VDD.n7950 VDD.n7949 25.6005
R9446 VDD.n7951 VDD.n7950 25.6005
R9447 VDD.n7952 VDD.n7951 25.6005
R9448 VDD.n7955 VDD.n7952 25.6005
R9449 VDD.n7956 VDD.n7955 25.6005
R9450 VDD.n7957 VDD.n7956 25.6005
R9451 VDD.n7957 VDD.n6881 25.6005
R9452 VDD.n7967 VDD.n6881 25.6005
R9453 VDD.n7968 VDD.n7967 25.6005
R9454 VDD.n7997 VDD.n7968 25.6005
R9455 VDD.n7997 VDD.n7996 25.6005
R9456 VDD.n8039 VDD.n8038 25.6005
R9457 VDD.n8038 VDD.n6860 25.6005
R9458 VDD.n7969 VDD.n6860 25.6005
R9459 VDD.n7972 VDD.n7969 25.6005
R9460 VDD.n7973 VDD.n7972 25.6005
R9461 VDD.n7976 VDD.n7973 25.6005
R9462 VDD.n7977 VDD.n7976 25.6005
R9463 VDD.n7980 VDD.n7977 25.6005
R9464 VDD.n7981 VDD.n7980 25.6005
R9465 VDD.n7984 VDD.n7981 25.6005
R9466 VDD.n7985 VDD.n7984 25.6005
R9467 VDD.n7988 VDD.n7985 25.6005
R9468 VDD.n7989 VDD.n7988 25.6005
R9469 VDD.n7992 VDD.n7989 25.6005
R9470 VDD.n7994 VDD.n7992 25.6005
R9471 VDD.n7995 VDD.n7994 25.6005
R9472 VDD.n7213 VDD.n7171 25.6005
R9473 VDD.n7182 VDD.n7171 25.6005
R9474 VDD.n7183 VDD.n7182 25.6005
R9475 VDD.n7186 VDD.n7183 25.6005
R9476 VDD.n7187 VDD.n7186 25.6005
R9477 VDD.n7190 VDD.n7187 25.6005
R9478 VDD.n7191 VDD.n7190 25.6005
R9479 VDD.n7194 VDD.n7191 25.6005
R9480 VDD.n7195 VDD.n7194 25.6005
R9481 VDD.n7198 VDD.n7195 25.6005
R9482 VDD.n7199 VDD.n7198 25.6005
R9483 VDD.n7202 VDD.n7199 25.6005
R9484 VDD.n7203 VDD.n7202 25.6005
R9485 VDD.n7206 VDD.n7203 25.6005
R9486 VDD.n7207 VDD.n7206 25.6005
R9487 VDD.n7208 VDD.n7207 25.6005
R9488 VDD.n7215 VDD.n7214 25.6005
R9489 VDD.n7215 VDD.n7163 25.6005
R9490 VDD.n7225 VDD.n7163 25.6005
R9491 VDD.n7226 VDD.n7225 25.6005
R9492 VDD.n7227 VDD.n7226 25.6005
R9493 VDD.n7227 VDD.n7155 25.6005
R9494 VDD.n7238 VDD.n7155 25.6005
R9495 VDD.n7239 VDD.n7238 25.6005
R9496 VDD.n7240 VDD.n7239 25.6005
R9497 VDD.n7240 VDD.n7148 25.6005
R9498 VDD.n7251 VDD.n7148 25.6005
R9499 VDD.n7252 VDD.n7251 25.6005
R9500 VDD.n7253 VDD.n7252 25.6005
R9501 VDD.n7253 VDD.n7141 25.6005
R9502 VDD.n7263 VDD.n7141 25.6005
R9503 VDD.n7264 VDD.n7263 25.6005
R9504 VDD.n7266 VDD.n7264 25.6005
R9505 VDD.n7266 VDD.n7265 25.6005
R9506 VDD.n7265 VDD.n7132 25.6005
R9507 VDD.n7316 VDD.n7132 25.6005
R9508 VDD.n7317 VDD.n7316 25.6005
R9509 VDD.n7321 VDD.n7317 25.6005
R9510 VDD.n7321 VDD.n7320 25.6005
R9511 VDD.n8114 VDD.n8113 25.6005
R9512 VDD.n8105 VDD.n6762 25.6005
R9513 VDD.n7768 VDD.n7753 25.6005
R9514 VDD.n7772 VDD.n7753 25.6005
R9515 VDD.n7773 VDD.n7772 25.6005
R9516 VDD.n7909 VDD.n7773 25.6005
R9517 VDD.n7909 VDD.n7908 25.6005
R9518 VDD.n7908 VDD.n7907 25.6005
R9519 VDD.n7907 VDD.n7774 25.6005
R9520 VDD.n7901 VDD.n7774 25.6005
R9521 VDD.n7901 VDD.n7900 25.6005
R9522 VDD.n7900 VDD.n7899 25.6005
R9523 VDD.n7899 VDD.n7781 25.6005
R9524 VDD.n7893 VDD.n7781 25.6005
R9525 VDD.n7893 VDD.n7892 25.6005
R9526 VDD.n7892 VDD.n7891 25.6005
R9527 VDD.n7891 VDD.n7787 25.6005
R9528 VDD.n7885 VDD.n7787 25.6005
R9529 VDD.n7885 VDD.n7884 25.6005
R9530 VDD.n7884 VDD.n7883 25.6005
R9531 VDD.n7883 VDD.n7795 25.6005
R9532 VDD.n7877 VDD.n7795 25.6005
R9533 VDD.n7877 VDD.n7876 25.6005
R9534 VDD.n7876 VDD.n7875 25.6005
R9535 VDD.n7875 VDD.n7802 25.6005
R9536 VDD.n7868 VDD.n7867 25.6005
R9537 VDD.n7867 VDD.n7866 25.6005
R9538 VDD.n7866 VDD.n7865 25.6005
R9539 VDD.n7865 VDD.n7863 25.6005
R9540 VDD.n7863 VDD.n7860 25.6005
R9541 VDD.n7860 VDD.n7859 25.6005
R9542 VDD.n7859 VDD.n7856 25.6005
R9543 VDD.n7856 VDD.n7855 25.6005
R9544 VDD.n7855 VDD.n7852 25.6005
R9545 VDD.n7852 VDD.n7851 25.6005
R9546 VDD.n7851 VDD.n7848 25.6005
R9547 VDD.n7848 VDD.n7847 25.6005
R9548 VDD.n7847 VDD.n7844 25.6005
R9549 VDD.n7844 VDD.n7843 25.6005
R9550 VDD.n7843 VDD.n7840 25.6005
R9551 VDD.n7840 VDD.n7839 25.6005
R9552 VDD.n7219 VDD.n7167 25.6005
R9553 VDD.n7220 VDD.n7219 25.6005
R9554 VDD.n7221 VDD.n7220 25.6005
R9555 VDD.n7221 VDD.n7159 25.6005
R9556 VDD.n7231 VDD.n7159 25.6005
R9557 VDD.n7232 VDD.n7231 25.6005
R9558 VDD.n7233 VDD.n7232 25.6005
R9559 VDD.n7233 VDD.n7151 25.6005
R9560 VDD.n7244 VDD.n7151 25.6005
R9561 VDD.n7245 VDD.n7244 25.6005
R9562 VDD.n7246 VDD.n7245 25.6005
R9563 VDD.n7246 VDD.n7145 25.6005
R9564 VDD.n7257 VDD.n7145 25.6005
R9565 VDD.n7258 VDD.n7257 25.6005
R9566 VDD.n7259 VDD.n7258 25.6005
R9567 VDD.n7259 VDD.n7137 25.6005
R9568 VDD.n7270 VDD.n7137 25.6005
R9569 VDD.n7271 VDD.n7270 25.6005
R9570 VDD.n7311 VDD.n7271 25.6005
R9571 VDD.n7311 VDD.n7310 25.6005
R9572 VDD.n7310 VDD.n7309 25.6005
R9573 VDD.n7309 VDD.n7307 25.6005
R9574 VDD.n7307 VDD.n7306 25.6005
R9575 VDD.n8118 VDD.n6418 25.6005
R9576 VDD.n6916 VDD.n6775 25.6005
R9577 VDD.n7917 VDD.n7916 25.6005
R9578 VDD.n7916 VDD.n7915 25.6005
R9579 VDD.n7915 VDD.n7747 25.6005
R9580 VDD.n7749 VDD.n7747 25.6005
R9581 VDD.n7815 VDD.n7749 25.6005
R9582 VDD.n7816 VDD.n7815 25.6005
R9583 VDD.n7817 VDD.n7816 25.6005
R9584 VDD.n7818 VDD.n7817 25.6005
R9585 VDD.n7820 VDD.n7818 25.6005
R9586 VDD.n7821 VDD.n7820 25.6005
R9587 VDD.n7822 VDD.n7821 25.6005
R9588 VDD.n7823 VDD.n7822 25.6005
R9589 VDD.n7825 VDD.n7823 25.6005
R9590 VDD.n7826 VDD.n7825 25.6005
R9591 VDD.n7827 VDD.n7826 25.6005
R9592 VDD.n7828 VDD.n7827 25.6005
R9593 VDD.n7830 VDD.n7828 25.6005
R9594 VDD.n7831 VDD.n7830 25.6005
R9595 VDD.n7832 VDD.n7831 25.6005
R9596 VDD.n7833 VDD.n7832 25.6005
R9597 VDD.n7835 VDD.n7833 25.6005
R9598 VDD.n7836 VDD.n7835 25.6005
R9599 VDD.n7837 VDD.n7836 25.6005
R9600 VDD.n2608 VDD.n2604 24.8476
R9601 VDD.n2927 VDD.n2923 24.8476
R9602 VDD.n2906 VDD.n2905 24.8476
R9603 VDD.n2827 VDD.n2785 24.8476
R9604 VDD.n3141 VDD.n3140 24.8476
R9605 VDD.n4655 VDD.n3998 24.8476
R9606 VDD.n4667 VDD.n3999 24.8476
R9607 VDD.n4515 VDD.n3455 24.8476
R9608 VDD.n5143 VDD.n3456 24.8476
R9609 VDD.n5137 VDD.n3792 24.8476
R9610 VDD.n5122 VDD.n3812 24.8476
R9611 VDD.n5150 VDD.n3448 24.8476
R9612 VDD.n4566 VDD.n4564 24.8476
R9613 VDD.n3949 VDD.n3948 24.8476
R9614 VDD.n5127 VDD.n5126 24.8476
R9615 VDD.n3192 VDD.n3186 24.8476
R9616 VDD.n3613 VDD.n3607 24.8476
R9617 VDD.n3473 VDD.n3467 24.8476
R9618 VDD.n14 VDD.n10 24.8476
R9619 VDD.n333 VDD.n329 24.8476
R9620 VDD.n312 VDD.n311 24.8476
R9621 VDD.n233 VDD.n191 24.8476
R9622 VDD.n547 VDD.n546 24.8476
R9623 VDD.n2061 VDD.n1404 24.8476
R9624 VDD.n2073 VDD.n1405 24.8476
R9625 VDD.n1921 VDD.n861 24.8476
R9626 VDD.n2549 VDD.n862 24.8476
R9627 VDD.n2543 VDD.n1198 24.8476
R9628 VDD.n2528 VDD.n1218 24.8476
R9629 VDD.n2556 VDD.n854 24.8476
R9630 VDD.n1972 VDD.n1970 24.8476
R9631 VDD.n1355 VDD.n1354 24.8476
R9632 VDD.n2533 VDD.n2532 24.8476
R9633 VDD.n598 VDD.n592 24.8476
R9634 VDD.n1019 VDD.n1013 24.8476
R9635 VDD.n879 VDD.n873 24.8476
R9636 VDD.n5577 VDD.n5573 24.8476
R9637 VDD.n5896 VDD.n5892 24.8476
R9638 VDD.n5875 VDD.n5874 24.8476
R9639 VDD.n5796 VDD.n5754 24.8476
R9640 VDD.n5553 VDD.n5552 24.8476
R9641 VDD.n5530 VDD.n5529 24.8476
R9642 VDD.n5493 VDD.n5484 24.8476
R9643 VDD.n5437 VDD.n5313 24.8476
R9644 VDD.n5397 VDD.n5324 24.8476
R9645 VDD.n5371 VDD.n5333 24.8476
R9646 VDD.n5355 VDD.n5343 24.8476
R9647 VDD.n6110 VDD.n6109 24.8476
R9648 VDD.n7624 VDD.n6967 24.8476
R9649 VDD.n7636 VDD.n6968 24.8476
R9650 VDD.n7484 VDD.n6424 24.8476
R9651 VDD.n8112 VDD.n6425 24.8476
R9652 VDD.n8106 VDD.n6761 24.8476
R9653 VDD.n8091 VDD.n6781 24.8476
R9654 VDD.n8119 VDD.n6417 24.8476
R9655 VDD.n7535 VDD.n7533 24.8476
R9656 VDD.n6918 VDD.n6917 24.8476
R9657 VDD.n8096 VDD.n8095 24.8476
R9658 VDD.n6161 VDD.n6155 24.8476
R9659 VDD.n6582 VDD.n6576 24.8476
R9660 VDD.n6442 VDD.n6436 24.8476
R9661 VDD.n5431 VDD.n5430 24.4711
R9662 VDD.n5381 VDD.n5380 24.4711
R9663 VDD.n5413 VDD.n5411 24.0946
R9664 VDD.n2659 VDD.n2658 23.737
R9665 VDD.n2998 VDD.n2737 23.737
R9666 VDD.n65 VDD.n64 23.737
R9667 VDD.n404 VDD.n143 23.737
R9668 VDD.n5628 VDD.n5627 23.737
R9669 VDD.n5967 VDD.n5706 23.737
R9670 VDD.n2612 VDD.n2611 23.3417
R9671 VDD.n2931 VDD.n2930 23.3417
R9672 VDD.n2909 VDD.n2744 23.3417
R9673 VDD.n2826 VDD.n2787 23.3417
R9674 VDD.n3144 VDD.n3124 23.3417
R9675 VDD.n4656 VDD.n4654 23.3417
R9676 VDD.n4696 VDD.n3969 23.3417
R9677 VDD.n4518 VDD.n4516 23.3417
R9678 VDD.n4589 VDD.n4048 23.3417
R9679 VDD.n4714 VDD.n4713 23.3417
R9680 VDD.n5121 VDD.n3813 23.3417
R9681 VDD.n4529 VDD.n4074 23.3417
R9682 VDD.n4568 VDD.n4567 23.3417
R9683 VDD.n4718 VDD.n3945 23.3417
R9684 VDD.n4761 VDD.n3807 23.3417
R9685 VDD.n3193 VDD.n3184 23.3417
R9686 VDD.n3614 VDD.n3605 23.3417
R9687 VDD.n3474 VDD.n3465 23.3417
R9688 VDD.n18 VDD.n17 23.3417
R9689 VDD.n337 VDD.n336 23.3417
R9690 VDD.n315 VDD.n150 23.3417
R9691 VDD.n232 VDD.n193 23.3417
R9692 VDD.n550 VDD.n530 23.3417
R9693 VDD.n2062 VDD.n2060 23.3417
R9694 VDD.n2102 VDD.n1375 23.3417
R9695 VDD.n1924 VDD.n1922 23.3417
R9696 VDD.n1995 VDD.n1454 23.3417
R9697 VDD.n2120 VDD.n2119 23.3417
R9698 VDD.n2527 VDD.n1219 23.3417
R9699 VDD.n1935 VDD.n1480 23.3417
R9700 VDD.n1974 VDD.n1973 23.3417
R9701 VDD.n2124 VDD.n1351 23.3417
R9702 VDD.n2167 VDD.n1213 23.3417
R9703 VDD.n599 VDD.n590 23.3417
R9704 VDD.n1020 VDD.n1011 23.3417
R9705 VDD.n880 VDD.n871 23.3417
R9706 VDD.n5581 VDD.n5580 23.3417
R9707 VDD.n5900 VDD.n5899 23.3417
R9708 VDD.n5878 VDD.n5713 23.3417
R9709 VDD.n5795 VDD.n5756 23.3417
R9710 VDD.n6113 VDD.n6093 23.3417
R9711 VDD.n7625 VDD.n7623 23.3417
R9712 VDD.n7665 VDD.n6938 23.3417
R9713 VDD.n7487 VDD.n7485 23.3417
R9714 VDD.n7558 VDD.n7017 23.3417
R9715 VDD.n7683 VDD.n7682 23.3417
R9716 VDD.n8090 VDD.n6782 23.3417
R9717 VDD.n7498 VDD.n7043 23.3417
R9718 VDD.n7537 VDD.n7536 23.3417
R9719 VDD.n7687 VDD.n6914 23.3417
R9720 VDD.n7730 VDD.n6776 23.3417
R9721 VDD.n6162 VDD.n6153 23.3417
R9722 VDD.n6583 VDD.n6574 23.3417
R9723 VDD.n6443 VDD.n6434 23.3417
R9724 VDD.n2823 VDD.n2798 23.1723
R9725 VDD.n2771 VDD.n2770 23.1723
R9726 VDD.n229 VDD.n204 23.1723
R9727 VDD.n177 VDD.n176 23.1723
R9728 VDD.n5792 VDD.n5767 23.1723
R9729 VDD.n5740 VDD.n5739 23.1723
R9730 VDD.n5461 VDD.n5444 22.7713
R9731 VDD.n5489 VDD.n5488 22.4624
R9732 VDD.n5346 VDD.n5345 22.4624
R9733 VDD.n4241 VDD.n4200 22.4005
R9734 VDD.n4903 VDD.n4902 22.4005
R9735 VDD.n1647 VDD.n1606 22.4005
R9736 VDD.n2309 VDD.n2308 22.4005
R9737 VDD.n7210 VDD.n7169 22.4005
R9738 VDD.n7872 VDD.n7871 22.4005
R9739 VDD.n5456 VDD.n5446 22.2123
R9740 VDD.n5451 VDD.n5450 22.2123
R9741 VDD.n5494 VDD.n5491 22.2123
R9742 VDD.n5425 VDD.n5315 22.2123
R9743 VDD.n5385 VDD.n5332 22.2123
R9744 VDD.n5390 VDD.n5389 22.2123
R9745 VDD.n3082 VDD.n2632 21.9733
R9746 VDD.n3082 VDD.n2634 21.9733
R9747 VDD.n3076 VDD.n2643 21.9733
R9748 VDD.n3070 VDD.n2643 21.9733
R9749 VDD.n3064 VDD.n2682 21.9733
R9750 VDD.n3064 VDD.n2685 21.9733
R9751 VDD.n3058 VDD.n2685 21.9733
R9752 VDD.n3052 VDD.n2694 21.9733
R9753 VDD.n3052 VDD.n2697 21.9733
R9754 VDD.n3046 VDD.n2697 21.9733
R9755 VDD.n3040 VDD.n2706 21.9733
R9756 VDD.n3040 VDD.n2709 21.9733
R9757 VDD.n3034 VDD.n2709 21.9733
R9758 VDD.n3028 VDD.n2718 21.9733
R9759 VDD.n3028 VDD.n2721 21.9733
R9760 VDD.n3022 VDD.n2727 21.9733
R9761 VDD.n3016 VDD.n2727 21.9733
R9762 VDD.n488 VDD.n38 21.9733
R9763 VDD.n488 VDD.n40 21.9733
R9764 VDD.n482 VDD.n49 21.9733
R9765 VDD.n476 VDD.n49 21.9733
R9766 VDD.n470 VDD.n88 21.9733
R9767 VDD.n470 VDD.n91 21.9733
R9768 VDD.n464 VDD.n91 21.9733
R9769 VDD.n458 VDD.n100 21.9733
R9770 VDD.n458 VDD.n103 21.9733
R9771 VDD.n452 VDD.n103 21.9733
R9772 VDD.n446 VDD.n112 21.9733
R9773 VDD.n446 VDD.n115 21.9733
R9774 VDD.n440 VDD.n115 21.9733
R9775 VDD.n434 VDD.n124 21.9733
R9776 VDD.n434 VDD.n127 21.9733
R9777 VDD.n428 VDD.n133 21.9733
R9778 VDD.n422 VDD.n133 21.9733
R9779 VDD.n6051 VDD.n5601 21.9733
R9780 VDD.n6051 VDD.n5603 21.9733
R9781 VDD.n6045 VDD.n5612 21.9733
R9782 VDD.n6039 VDD.n5612 21.9733
R9783 VDD.n6033 VDD.n5651 21.9733
R9784 VDD.n6033 VDD.n5654 21.9733
R9785 VDD.n6027 VDD.n5654 21.9733
R9786 VDD.n6021 VDD.n5663 21.9733
R9787 VDD.n6021 VDD.n5666 21.9733
R9788 VDD.n6015 VDD.n5666 21.9733
R9789 VDD.n6009 VDD.n5675 21.9733
R9790 VDD.n6009 VDD.n5678 21.9733
R9791 VDD.n6003 VDD.n5678 21.9733
R9792 VDD.n5997 VDD.n5687 21.9733
R9793 VDD.n5997 VDD.n5690 21.9733
R9794 VDD.n5991 VDD.n5696 21.9733
R9795 VDD.n5985 VDD.n5696 21.9733
R9796 VDD.n2615 VDD.n2602 21.8358
R9797 VDD.n2934 VDD.n2921 21.8358
R9798 VDD.n3145 VDD.n3123 21.8358
R9799 VDD.n4035 VDD.n4004 21.8358
R9800 VDD.n4695 VDD.n3970 21.8358
R9801 VDD.n4519 VDD.n4082 21.8358
R9802 VDD.n4591 VDD.n4590 21.8358
R9803 VDD.n4712 VDD.n3954 21.8358
R9804 VDD.n5118 VDD.n5117 21.8358
R9805 VDD.n4530 VDD.n4073 21.8358
R9806 VDD.n4571 VDD.n4570 21.8358
R9807 VDD.n4719 VDD.n3944 21.8358
R9808 VDD.n4763 VDD.n4762 21.8358
R9809 VDD.n3197 VDD.n3196 21.8358
R9810 VDD.n3618 VDD.n3617 21.8358
R9811 VDD.n3478 VDD.n3477 21.8358
R9812 VDD.n21 VDD.n8 21.8358
R9813 VDD.n340 VDD.n327 21.8358
R9814 VDD.n551 VDD.n529 21.8358
R9815 VDD.n1441 VDD.n1410 21.8358
R9816 VDD.n2101 VDD.n1376 21.8358
R9817 VDD.n1925 VDD.n1488 21.8358
R9818 VDD.n1997 VDD.n1996 21.8358
R9819 VDD.n2118 VDD.n1360 21.8358
R9820 VDD.n2524 VDD.n2523 21.8358
R9821 VDD.n1936 VDD.n1479 21.8358
R9822 VDD.n1977 VDD.n1976 21.8358
R9823 VDD.n2125 VDD.n1350 21.8358
R9824 VDD.n2169 VDD.n2168 21.8358
R9825 VDD.n603 VDD.n602 21.8358
R9826 VDD.n1024 VDD.n1023 21.8358
R9827 VDD.n884 VDD.n883 21.8358
R9828 VDD.n5584 VDD.n5571 21.8358
R9829 VDD.n5903 VDD.n5890 21.8358
R9830 VDD.n6114 VDD.n6092 21.8358
R9831 VDD.n7004 VDD.n6973 21.8358
R9832 VDD.n7664 VDD.n6939 21.8358
R9833 VDD.n7488 VDD.n7051 21.8358
R9834 VDD.n7560 VDD.n7559 21.8358
R9835 VDD.n7681 VDD.n6923 21.8358
R9836 VDD.n8087 VDD.n8086 21.8358
R9837 VDD.n7499 VDD.n7042 21.8358
R9838 VDD.n7540 VDD.n7539 21.8358
R9839 VDD.n7688 VDD.n6913 21.8358
R9840 VDD.n7732 VDD.n7731 21.8358
R9841 VDD.n6166 VDD.n6165 21.8358
R9842 VDD.n6587 VDD.n6586 21.8358
R9843 VDD.n6447 VDD.n6446 21.8358
R9844 VDD.n5501 VDD.n5500 21.7826
R9845 VDD.n2771 VDD.n2749 21.7605
R9846 VDD.n2823 VDD.n2822 21.7605
R9847 VDD.n177 VDD.n155 21.7605
R9848 VDD.n229 VDD.n228 21.7605
R9849 VDD.n5740 VDD.n5718 21.7605
R9850 VDD.n5792 VDD.n5791 21.7605
R9851 VDD.n3076 VDD.t75 21.6502
R9852 VDD.t73 VDD.n2721 21.6502
R9853 VDD.n482 VDD.t121 21.6502
R9854 VDD.t123 VDD.n127 21.6502
R9855 VDD.n6045 VDD.t161 21.6502
R9856 VDD.t198 VDD.n5690 21.6502
R9857 VDD.n5376 VDD.n5332 20.7064
R9858 VDD.n2902 VDD.n2901 20.4805
R9859 VDD.n2817 VDD.n2782 20.4805
R9860 VDD.n308 VDD.n307 20.4805
R9861 VDD.n223 VDD.n188 20.4805
R9862 VDD.n5871 VDD.n5870 20.4805
R9863 VDD.n5786 VDD.n5751 20.4805
R9864 VDD.n3133 VDD.n3132 20.3299
R9865 VDD.n3158 VDD.n3157 20.3299
R9866 VDD.n3391 VDD.n3390 20.3299
R9867 VDD.n3404 VDD.n3403 20.3299
R9868 VDD.n3417 VDD.n3416 20.3299
R9869 VDD.n3430 VDD.n3429 20.3299
R9870 VDD.n3374 VDD.n3373 20.3299
R9871 VDD.n3360 VDD.n3359 20.3299
R9872 VDD.n3346 VDD.n3345 20.3299
R9873 VDD.n3114 VDD.n3113 20.3299
R9874 VDD.n5171 VDD.n5170 20.3299
R9875 VDD.n4036 VDD.n4033 20.3299
R9876 VDD.n3973 VDD.n3972 20.3299
R9877 VDD.n4350 VDD.n4349 20.3299
R9878 VDD.n4523 VDD.n4522 20.3299
R9879 VDD.n4603 VDD.n4046 20.3299
R9880 VDD.n4709 VDD.n4708 20.3299
R9881 VDD.n3844 VDD.n3815 20.3299
R9882 VDD.n4798 VDD.n4786 20.3299
R9883 VDD.n4334 VDD.n4303 20.3299
R9884 VDD.n4077 VDD.n4076 20.3299
R9885 VDD.n4569 VDD.n4038 20.3299
R9886 VDD.n3977 VDD.n3976 20.3299
R9887 VDD.n4974 VDD.n4752 20.3299
R9888 VDD.n4951 VDD.n4776 20.3299
R9889 VDD.n3200 VDD.n3199 20.3299
R9890 VDD.n3214 VDD.n3213 20.3299
R9891 VDD.n3288 VDD.n3287 20.3299
R9892 VDD.n3301 VDD.n3300 20.3299
R9893 VDD.n3314 VDD.n3313 20.3299
R9894 VDD.n3327 VDD.n3326 20.3299
R9895 VDD.n3271 VDD.n3270 20.3299
R9896 VDD.n3257 VDD.n3256 20.3299
R9897 VDD.n3243 VDD.n3242 20.3299
R9898 VDD.n3229 VDD.n3228 20.3299
R9899 VDD.n3170 VDD.n3169 20.3299
R9900 VDD.n3621 VDD.n3620 20.3299
R9901 VDD.n3635 VDD.n3634 20.3299
R9902 VDD.n3649 VDD.n3648 20.3299
R9903 VDD.n3662 VDD.n3661 20.3299
R9904 VDD.n3675 VDD.n3674 20.3299
R9905 VDD.n3688 VDD.n3687 20.3299
R9906 VDD.n3701 VDD.n3700 20.3299
R9907 VDD.n3714 VDD.n3713 20.3299
R9908 VDD.n3728 VDD.n3727 20.3299
R9909 VDD.n3741 VDD.n3740 20.3299
R9910 VDD.n3754 VDD.n3753 20.3299
R9911 VDD.n3767 VDD.n3766 20.3299
R9912 VDD.n3780 VDD.n3779 20.3299
R9913 VDD.n3581 VDD.n3580 20.3299
R9914 VDD.n3567 VDD.n3566 20.3299
R9915 VDD.n3553 VDD.n3552 20.3299
R9916 VDD.n3539 VDD.n3538 20.3299
R9917 VDD.n3525 VDD.n3524 20.3299
R9918 VDD.n3511 VDD.n3510 20.3299
R9919 VDD.n3496 VDD.n3495 20.3299
R9920 VDD.n3481 VDD.n3480 20.3299
R9921 VDD.n539 VDD.n538 20.3299
R9922 VDD.n564 VDD.n563 20.3299
R9923 VDD.n797 VDD.n796 20.3299
R9924 VDD.n810 VDD.n809 20.3299
R9925 VDD.n823 VDD.n822 20.3299
R9926 VDD.n836 VDD.n835 20.3299
R9927 VDD.n780 VDD.n779 20.3299
R9928 VDD.n766 VDD.n765 20.3299
R9929 VDD.n752 VDD.n751 20.3299
R9930 VDD.n520 VDD.n519 20.3299
R9931 VDD.n2577 VDD.n2576 20.3299
R9932 VDD.n1442 VDD.n1439 20.3299
R9933 VDD.n1379 VDD.n1378 20.3299
R9934 VDD.n1756 VDD.n1755 20.3299
R9935 VDD.n1929 VDD.n1928 20.3299
R9936 VDD.n2009 VDD.n1452 20.3299
R9937 VDD.n2115 VDD.n2114 20.3299
R9938 VDD.n1250 VDD.n1221 20.3299
R9939 VDD.n2204 VDD.n2192 20.3299
R9940 VDD.n1740 VDD.n1709 20.3299
R9941 VDD.n1483 VDD.n1482 20.3299
R9942 VDD.n1975 VDD.n1444 20.3299
R9943 VDD.n1383 VDD.n1382 20.3299
R9944 VDD.n2380 VDD.n2158 20.3299
R9945 VDD.n2357 VDD.n2182 20.3299
R9946 VDD.n606 VDD.n605 20.3299
R9947 VDD.n620 VDD.n619 20.3299
R9948 VDD.n694 VDD.n693 20.3299
R9949 VDD.n707 VDD.n706 20.3299
R9950 VDD.n720 VDD.n719 20.3299
R9951 VDD.n733 VDD.n732 20.3299
R9952 VDD.n677 VDD.n676 20.3299
R9953 VDD.n663 VDD.n662 20.3299
R9954 VDD.n649 VDD.n648 20.3299
R9955 VDD.n635 VDD.n634 20.3299
R9956 VDD.n576 VDD.n575 20.3299
R9957 VDD.n1027 VDD.n1026 20.3299
R9958 VDD.n1041 VDD.n1040 20.3299
R9959 VDD.n1055 VDD.n1054 20.3299
R9960 VDD.n1068 VDD.n1067 20.3299
R9961 VDD.n1081 VDD.n1080 20.3299
R9962 VDD.n1094 VDD.n1093 20.3299
R9963 VDD.n1107 VDD.n1106 20.3299
R9964 VDD.n1120 VDD.n1119 20.3299
R9965 VDD.n1134 VDD.n1133 20.3299
R9966 VDD.n1147 VDD.n1146 20.3299
R9967 VDD.n1160 VDD.n1159 20.3299
R9968 VDD.n1173 VDD.n1172 20.3299
R9969 VDD.n1186 VDD.n1185 20.3299
R9970 VDD.n987 VDD.n986 20.3299
R9971 VDD.n973 VDD.n972 20.3299
R9972 VDD.n959 VDD.n958 20.3299
R9973 VDD.n945 VDD.n944 20.3299
R9974 VDD.n931 VDD.n930 20.3299
R9975 VDD.n917 VDD.n916 20.3299
R9976 VDD.n902 VDD.n901 20.3299
R9977 VDD.n887 VDD.n886 20.3299
R9978 VDD.n6102 VDD.n6101 20.3299
R9979 VDD.n6127 VDD.n6126 20.3299
R9980 VDD.n6360 VDD.n6359 20.3299
R9981 VDD.n6373 VDD.n6372 20.3299
R9982 VDD.n6386 VDD.n6385 20.3299
R9983 VDD.n6399 VDD.n6398 20.3299
R9984 VDD.n6343 VDD.n6342 20.3299
R9985 VDD.n6329 VDD.n6328 20.3299
R9986 VDD.n6315 VDD.n6314 20.3299
R9987 VDD.n6083 VDD.n6082 20.3299
R9988 VDD.n8140 VDD.n8139 20.3299
R9989 VDD.n7005 VDD.n7002 20.3299
R9990 VDD.n6942 VDD.n6941 20.3299
R9991 VDD.n7319 VDD.n7318 20.3299
R9992 VDD.n7492 VDD.n7491 20.3299
R9993 VDD.n7572 VDD.n7015 20.3299
R9994 VDD.n7678 VDD.n7677 20.3299
R9995 VDD.n6813 VDD.n6784 20.3299
R9996 VDD.n7767 VDD.n7755 20.3299
R9997 VDD.n7303 VDD.n7272 20.3299
R9998 VDD.n7046 VDD.n7045 20.3299
R9999 VDD.n7538 VDD.n7007 20.3299
R10000 VDD.n6946 VDD.n6945 20.3299
R10001 VDD.n7943 VDD.n7721 20.3299
R10002 VDD.n7920 VDD.n7745 20.3299
R10003 VDD.n6169 VDD.n6168 20.3299
R10004 VDD.n6183 VDD.n6182 20.3299
R10005 VDD.n6257 VDD.n6256 20.3299
R10006 VDD.n6270 VDD.n6269 20.3299
R10007 VDD.n6283 VDD.n6282 20.3299
R10008 VDD.n6296 VDD.n6295 20.3299
R10009 VDD.n6240 VDD.n6239 20.3299
R10010 VDD.n6226 VDD.n6225 20.3299
R10011 VDD.n6212 VDD.n6211 20.3299
R10012 VDD.n6198 VDD.n6197 20.3299
R10013 VDD.n6139 VDD.n6138 20.3299
R10014 VDD.n6590 VDD.n6589 20.3299
R10015 VDD.n6604 VDD.n6603 20.3299
R10016 VDD.n6618 VDD.n6617 20.3299
R10017 VDD.n6631 VDD.n6630 20.3299
R10018 VDD.n6644 VDD.n6643 20.3299
R10019 VDD.n6657 VDD.n6656 20.3299
R10020 VDD.n6670 VDD.n6669 20.3299
R10021 VDD.n6683 VDD.n6682 20.3299
R10022 VDD.n6697 VDD.n6696 20.3299
R10023 VDD.n6710 VDD.n6709 20.3299
R10024 VDD.n6723 VDD.n6722 20.3299
R10025 VDD.n6736 VDD.n6735 20.3299
R10026 VDD.n6749 VDD.n6748 20.3299
R10027 VDD.n6550 VDD.n6549 20.3299
R10028 VDD.n6536 VDD.n6535 20.3299
R10029 VDD.n6522 VDD.n6521 20.3299
R10030 VDD.n6508 VDD.n6507 20.3299
R10031 VDD.n6494 VDD.n6493 20.3299
R10032 VDD.n6480 VDD.n6479 20.3299
R10033 VDD.n6465 VDD.n6464 20.3299
R10034 VDD.n6450 VDD.n6449 20.3299
R10035 VDD.n2897 VDD.n2755 20.1605
R10036 VDD.n2836 VDD.n2835 20.1605
R10037 VDD.n303 VDD.n161 20.1605
R10038 VDD.n242 VDD.n241 20.1605
R10039 VDD.n5866 VDD.n5724 20.1605
R10040 VDD.n5805 VDD.n5804 20.1605
R10041 VDD.n5515 VDD.n5477 19.3108
R10042 VDD.n3127 VDD.n3120 19.1835
R10043 VDD.n3152 VDD.n3119 19.1835
R10044 VDD.n3385 VDD.n3381 19.1835
R10045 VDD.n3398 VDD.n3380 19.1835
R10046 VDD.n3411 VDD.n3379 19.1835
R10047 VDD.n3424 VDD.n3378 19.1835
R10048 VDD.n3368 VDD.n3364 19.1835
R10049 VDD.n3354 VDD.n3350 19.1835
R10050 VDD.n3340 VDD.n3336 19.1835
R10051 VDD.n3108 VDD.n3104 19.1835
R10052 VDD.n5165 VDD.n3103 19.1835
R10053 VDD.n533 VDD.n526 19.1835
R10054 VDD.n558 VDD.n525 19.1835
R10055 VDD.n791 VDD.n787 19.1835
R10056 VDD.n804 VDD.n786 19.1835
R10057 VDD.n817 VDD.n785 19.1835
R10058 VDD.n830 VDD.n784 19.1835
R10059 VDD.n774 VDD.n770 19.1835
R10060 VDD.n760 VDD.n756 19.1835
R10061 VDD.n746 VDD.n742 19.1835
R10062 VDD.n514 VDD.n510 19.1835
R10063 VDD.n2571 VDD.n509 19.1835
R10064 VDD.n6096 VDD.n6089 19.1835
R10065 VDD.n6121 VDD.n6088 19.1835
R10066 VDD.n6354 VDD.n6350 19.1835
R10067 VDD.n6367 VDD.n6349 19.1835
R10068 VDD.n6380 VDD.n6348 19.1835
R10069 VDD.n6393 VDD.n6347 19.1835
R10070 VDD.n6337 VDD.n6333 19.1835
R10071 VDD.n6323 VDD.n6319 19.1835
R10072 VDD.n6309 VDD.n6305 19.1835
R10073 VDD.n6077 VDD.n6073 19.1835
R10074 VDD.n8134 VDD.n6072 19.1835
R10075 VDD.n3206 VDD.n3180 19.1564
R10076 VDD.n3219 VDD.n3208 19.1564
R10077 VDD.n3293 VDD.n3282 19.1564
R10078 VDD.n3306 VDD.n3295 19.1564
R10079 VDD.n3319 VDD.n3308 19.1564
R10080 VDD.n3332 VDD.n3321 19.1564
R10081 VDD.n3276 VDD.n3265 19.1564
R10082 VDD.n3262 VDD.n3251 19.1564
R10083 VDD.n3248 VDD.n3237 19.1564
R10084 VDD.n3234 VDD.n3223 19.1564
R10085 VDD.n3175 VDD.n3164 19.1564
R10086 VDD.n3627 VDD.n3601 19.1564
R10087 VDD.n3640 VDD.n3629 19.1564
R10088 VDD.n3654 VDD.n3643 19.1564
R10089 VDD.n3667 VDD.n3656 19.1564
R10090 VDD.n3680 VDD.n3669 19.1564
R10091 VDD.n3693 VDD.n3682 19.1564
R10092 VDD.n3706 VDD.n3695 19.1564
R10093 VDD.n3719 VDD.n3708 19.1564
R10094 VDD.n3733 VDD.n3722 19.1564
R10095 VDD.n3746 VDD.n3735 19.1564
R10096 VDD.n3759 VDD.n3748 19.1564
R10097 VDD.n3772 VDD.n3761 19.1564
R10098 VDD.n3785 VDD.n3774 19.1564
R10099 VDD.n3586 VDD.n3575 19.1564
R10100 VDD.n3572 VDD.n3561 19.1564
R10101 VDD.n3558 VDD.n3547 19.1564
R10102 VDD.n3544 VDD.n3533 19.1564
R10103 VDD.n3530 VDD.n3519 19.1564
R10104 VDD.n3516 VDD.n3505 19.1564
R10105 VDD.n3501 VDD.n3490 19.1564
R10106 VDD.n3487 VDD.n3461 19.1564
R10107 VDD.n612 VDD.n586 19.1564
R10108 VDD.n625 VDD.n614 19.1564
R10109 VDD.n699 VDD.n688 19.1564
R10110 VDD.n712 VDD.n701 19.1564
R10111 VDD.n725 VDD.n714 19.1564
R10112 VDD.n738 VDD.n727 19.1564
R10113 VDD.n682 VDD.n671 19.1564
R10114 VDD.n668 VDD.n657 19.1564
R10115 VDD.n654 VDD.n643 19.1564
R10116 VDD.n640 VDD.n629 19.1564
R10117 VDD.n581 VDD.n570 19.1564
R10118 VDD.n1033 VDD.n1007 19.1564
R10119 VDD.n1046 VDD.n1035 19.1564
R10120 VDD.n1060 VDD.n1049 19.1564
R10121 VDD.n1073 VDD.n1062 19.1564
R10122 VDD.n1086 VDD.n1075 19.1564
R10123 VDD.n1099 VDD.n1088 19.1564
R10124 VDD.n1112 VDD.n1101 19.1564
R10125 VDD.n1125 VDD.n1114 19.1564
R10126 VDD.n1139 VDD.n1128 19.1564
R10127 VDD.n1152 VDD.n1141 19.1564
R10128 VDD.n1165 VDD.n1154 19.1564
R10129 VDD.n1178 VDD.n1167 19.1564
R10130 VDD.n1191 VDD.n1180 19.1564
R10131 VDD.n992 VDD.n981 19.1564
R10132 VDD.n978 VDD.n967 19.1564
R10133 VDD.n964 VDD.n953 19.1564
R10134 VDD.n950 VDD.n939 19.1564
R10135 VDD.n936 VDD.n925 19.1564
R10136 VDD.n922 VDD.n911 19.1564
R10137 VDD.n907 VDD.n896 19.1564
R10138 VDD.n893 VDD.n867 19.1564
R10139 VDD.n6175 VDD.n6149 19.1564
R10140 VDD.n6188 VDD.n6177 19.1564
R10141 VDD.n6262 VDD.n6251 19.1564
R10142 VDD.n6275 VDD.n6264 19.1564
R10143 VDD.n6288 VDD.n6277 19.1564
R10144 VDD.n6301 VDD.n6290 19.1564
R10145 VDD.n6245 VDD.n6234 19.1564
R10146 VDD.n6231 VDD.n6220 19.1564
R10147 VDD.n6217 VDD.n6206 19.1564
R10148 VDD.n6203 VDD.n6192 19.1564
R10149 VDD.n6144 VDD.n6133 19.1564
R10150 VDD.n6596 VDD.n6570 19.1564
R10151 VDD.n6609 VDD.n6598 19.1564
R10152 VDD.n6623 VDD.n6612 19.1564
R10153 VDD.n6636 VDD.n6625 19.1564
R10154 VDD.n6649 VDD.n6638 19.1564
R10155 VDD.n6662 VDD.n6651 19.1564
R10156 VDD.n6675 VDD.n6664 19.1564
R10157 VDD.n6688 VDD.n6677 19.1564
R10158 VDD.n6702 VDD.n6691 19.1564
R10159 VDD.n6715 VDD.n6704 19.1564
R10160 VDD.n6728 VDD.n6717 19.1564
R10161 VDD.n6741 VDD.n6730 19.1564
R10162 VDD.n6754 VDD.n6743 19.1564
R10163 VDD.n6555 VDD.n6544 19.1564
R10164 VDD.n6541 VDD.n6530 19.1564
R10165 VDD.n6527 VDD.n6516 19.1564
R10166 VDD.n6513 VDD.n6502 19.1564
R10167 VDD.n6499 VDD.n6488 19.1564
R10168 VDD.n6485 VDD.n6474 19.1564
R10169 VDD.n6470 VDD.n6459 19.1564
R10170 VDD.n6456 VDD.n6430 19.1564
R10171 VDD.n3131 VDD.n3126 18.824
R10172 VDD.n3156 VDD.n3151 18.824
R10173 VDD.n3389 VDD.n3384 18.824
R10174 VDD.n3402 VDD.n3397 18.824
R10175 VDD.n3415 VDD.n3410 18.824
R10176 VDD.n3428 VDD.n3423 18.824
R10177 VDD.n3372 VDD.n3367 18.824
R10178 VDD.n3358 VDD.n3353 18.824
R10179 VDD.n3344 VDD.n3339 18.824
R10180 VDD.n3112 VDD.n3107 18.824
R10181 VDD.n5169 VDD.n5164 18.824
R10182 VDD.n4617 VDD.n4616 18.824
R10183 VDD.n4723 VDD.n3938 18.824
R10184 VDD.n4441 VDD.n4133 18.824
R10185 VDD.n4510 VDD.n4081 18.824
R10186 VDD.n4602 VDD.n4047 18.824
R10187 VDD.n4679 VDD.n3956 18.824
R10188 VDD.n3847 VDD.n3845 18.824
R10189 VDD.n4796 VDD.n4795 18.824
R10190 VDD.n4333 VDD.n4304 18.824
R10191 VDD.n4313 VDD.n4312 18.824
R10192 VDD.n4613 VDD.n4612 18.824
R10193 VDD.n4691 VDD.n3980 18.824
R10194 VDD.n4973 VDD.n4753 18.824
R10195 VDD.n4952 VDD.n4774 18.824
R10196 VDD.n3203 VDD.n3182 18.824
R10197 VDD.n3216 VDD.n3210 18.824
R10198 VDD.n3290 VDD.n3284 18.824
R10199 VDD.n3303 VDD.n3297 18.824
R10200 VDD.n3316 VDD.n3310 18.824
R10201 VDD.n3329 VDD.n3323 18.824
R10202 VDD.n3273 VDD.n3267 18.824
R10203 VDD.n3259 VDD.n3253 18.824
R10204 VDD.n3245 VDD.n3239 18.824
R10205 VDD.n3231 VDD.n3225 18.824
R10206 VDD.n3172 VDD.n3166 18.824
R10207 VDD.n3624 VDD.n3603 18.824
R10208 VDD.n3637 VDD.n3631 18.824
R10209 VDD.n3651 VDD.n3645 18.824
R10210 VDD.n3664 VDD.n3658 18.824
R10211 VDD.n3677 VDD.n3671 18.824
R10212 VDD.n3690 VDD.n3684 18.824
R10213 VDD.n3703 VDD.n3697 18.824
R10214 VDD.n3716 VDD.n3710 18.824
R10215 VDD.n3730 VDD.n3724 18.824
R10216 VDD.n3743 VDD.n3737 18.824
R10217 VDD.n3756 VDD.n3750 18.824
R10218 VDD.n3769 VDD.n3763 18.824
R10219 VDD.n3782 VDD.n3776 18.824
R10220 VDD.n3583 VDD.n3577 18.824
R10221 VDD.n3569 VDD.n3563 18.824
R10222 VDD.n3555 VDD.n3549 18.824
R10223 VDD.n3541 VDD.n3535 18.824
R10224 VDD.n3527 VDD.n3521 18.824
R10225 VDD.n3513 VDD.n3507 18.824
R10226 VDD.n3498 VDD.n3492 18.824
R10227 VDD.n3484 VDD.n3463 18.824
R10228 VDD.n537 VDD.n532 18.824
R10229 VDD.n562 VDD.n557 18.824
R10230 VDD.n795 VDD.n790 18.824
R10231 VDD.n808 VDD.n803 18.824
R10232 VDD.n821 VDD.n816 18.824
R10233 VDD.n834 VDD.n829 18.824
R10234 VDD.n778 VDD.n773 18.824
R10235 VDD.n764 VDD.n759 18.824
R10236 VDD.n750 VDD.n745 18.824
R10237 VDD.n518 VDD.n513 18.824
R10238 VDD.n2575 VDD.n2570 18.824
R10239 VDD.n2023 VDD.n2022 18.824
R10240 VDD.n2129 VDD.n1344 18.824
R10241 VDD.n1847 VDD.n1539 18.824
R10242 VDD.n1916 VDD.n1487 18.824
R10243 VDD.n2008 VDD.n1453 18.824
R10244 VDD.n2085 VDD.n1362 18.824
R10245 VDD.n1253 VDD.n1251 18.824
R10246 VDD.n2202 VDD.n2201 18.824
R10247 VDD.n1739 VDD.n1710 18.824
R10248 VDD.n1719 VDD.n1718 18.824
R10249 VDD.n2019 VDD.n2018 18.824
R10250 VDD.n2097 VDD.n1386 18.824
R10251 VDD.n2379 VDD.n2159 18.824
R10252 VDD.n2358 VDD.n2180 18.824
R10253 VDD.n609 VDD.n588 18.824
R10254 VDD.n622 VDD.n616 18.824
R10255 VDD.n696 VDD.n690 18.824
R10256 VDD.n709 VDD.n703 18.824
R10257 VDD.n722 VDD.n716 18.824
R10258 VDD.n735 VDD.n729 18.824
R10259 VDD.n679 VDD.n673 18.824
R10260 VDD.n665 VDD.n659 18.824
R10261 VDD.n651 VDD.n645 18.824
R10262 VDD.n637 VDD.n631 18.824
R10263 VDD.n578 VDD.n572 18.824
R10264 VDD.n1030 VDD.n1009 18.824
R10265 VDD.n1043 VDD.n1037 18.824
R10266 VDD.n1057 VDD.n1051 18.824
R10267 VDD.n1070 VDD.n1064 18.824
R10268 VDD.n1083 VDD.n1077 18.824
R10269 VDD.n1096 VDD.n1090 18.824
R10270 VDD.n1109 VDD.n1103 18.824
R10271 VDD.n1122 VDD.n1116 18.824
R10272 VDD.n1136 VDD.n1130 18.824
R10273 VDD.n1149 VDD.n1143 18.824
R10274 VDD.n1162 VDD.n1156 18.824
R10275 VDD.n1175 VDD.n1169 18.824
R10276 VDD.n1188 VDD.n1182 18.824
R10277 VDD.n989 VDD.n983 18.824
R10278 VDD.n975 VDD.n969 18.824
R10279 VDD.n961 VDD.n955 18.824
R10280 VDD.n947 VDD.n941 18.824
R10281 VDD.n933 VDD.n927 18.824
R10282 VDD.n919 VDD.n913 18.824
R10283 VDD.n904 VDD.n898 18.824
R10284 VDD.n890 VDD.n869 18.824
R10285 VDD.n5505 VDD.n5477 18.824
R10286 VDD.n5490 VDD.n5489 18.824
R10287 VDD.n5399 VDD.n5327 18.824
R10288 VDD.n5369 VDD.n5368 18.824
R10289 VDD.n5345 VDD.n5341 18.824
R10290 VDD.n6100 VDD.n6095 18.824
R10291 VDD.n6125 VDD.n6120 18.824
R10292 VDD.n6358 VDD.n6353 18.824
R10293 VDD.n6371 VDD.n6366 18.824
R10294 VDD.n6384 VDD.n6379 18.824
R10295 VDD.n6397 VDD.n6392 18.824
R10296 VDD.n6341 VDD.n6336 18.824
R10297 VDD.n6327 VDD.n6322 18.824
R10298 VDD.n6313 VDD.n6308 18.824
R10299 VDD.n6081 VDD.n6076 18.824
R10300 VDD.n8138 VDD.n8133 18.824
R10301 VDD.n7586 VDD.n7585 18.824
R10302 VDD.n7692 VDD.n6907 18.824
R10303 VDD.n7410 VDD.n7102 18.824
R10304 VDD.n7479 VDD.n7050 18.824
R10305 VDD.n7571 VDD.n7016 18.824
R10306 VDD.n7648 VDD.n6925 18.824
R10307 VDD.n6816 VDD.n6814 18.824
R10308 VDD.n7765 VDD.n7764 18.824
R10309 VDD.n7302 VDD.n7273 18.824
R10310 VDD.n7282 VDD.n7281 18.824
R10311 VDD.n7582 VDD.n7581 18.824
R10312 VDD.n7660 VDD.n6949 18.824
R10313 VDD.n7942 VDD.n7722 18.824
R10314 VDD.n7921 VDD.n7743 18.824
R10315 VDD.n6172 VDD.n6151 18.824
R10316 VDD.n6185 VDD.n6179 18.824
R10317 VDD.n6259 VDD.n6253 18.824
R10318 VDD.n6272 VDD.n6266 18.824
R10319 VDD.n6285 VDD.n6279 18.824
R10320 VDD.n6298 VDD.n6292 18.824
R10321 VDD.n6242 VDD.n6236 18.824
R10322 VDD.n6228 VDD.n6222 18.824
R10323 VDD.n6214 VDD.n6208 18.824
R10324 VDD.n6200 VDD.n6194 18.824
R10325 VDD.n6141 VDD.n6135 18.824
R10326 VDD.n6593 VDD.n6572 18.824
R10327 VDD.n6606 VDD.n6600 18.824
R10328 VDD.n6620 VDD.n6614 18.824
R10329 VDD.n6633 VDD.n6627 18.824
R10330 VDD.n6646 VDD.n6640 18.824
R10331 VDD.n6659 VDD.n6653 18.824
R10332 VDD.n6672 VDD.n6666 18.824
R10333 VDD.n6685 VDD.n6679 18.824
R10334 VDD.n6699 VDD.n6693 18.824
R10335 VDD.n6712 VDD.n6706 18.824
R10336 VDD.n6725 VDD.n6719 18.824
R10337 VDD.n6738 VDD.n6732 18.824
R10338 VDD.n6751 VDD.n6745 18.824
R10339 VDD.n6552 VDD.n6546 18.824
R10340 VDD.n6538 VDD.n6532 18.824
R10341 VDD.n6524 VDD.n6518 18.824
R10342 VDD.n6510 VDD.n6504 18.824
R10343 VDD.n6496 VDD.n6490 18.824
R10344 VDD.n6482 VDD.n6476 18.824
R10345 VDD.n6467 VDD.n6461 18.824
R10346 VDD.n6453 VDD.n6432 18.824
R10347 VDD.n2657 VDD.n2656 18.5605
R10348 VDD.n2997 VDD.n2739 18.5605
R10349 VDD.n63 VDD.n62 18.5605
R10350 VDD.n403 VDD.n145 18.5605
R10351 VDD.n5626 VDD.n5625 18.5605
R10352 VDD.n5966 VDD.n5708 18.5605
R10353 VDD.n3070 VDD.t67 17.7726
R10354 VDD.n2718 VDD.t63 17.7726
R10355 VDD.n476 VDD.t105 17.7726
R10356 VDD.n124 VDD.t343 17.7726
R10357 VDD.n6039 VDD.t163 17.7726
R10358 VDD.n5687 VDD.t212 17.7726
R10359 VDD.n3128 VDD.n3127 17.3181
R10360 VDD.n3153 VDD.n3152 17.3181
R10361 VDD.n3386 VDD.n3385 17.3181
R10362 VDD.n3399 VDD.n3398 17.3181
R10363 VDD.n3412 VDD.n3411 17.3181
R10364 VDD.n3425 VDD.n3424 17.3181
R10365 VDD.n3369 VDD.n3368 17.3181
R10366 VDD.n3355 VDD.n3354 17.3181
R10367 VDD.n3341 VDD.n3340 17.3181
R10368 VDD.n3109 VDD.n3108 17.3181
R10369 VDD.n5166 VDD.n5165 17.3181
R10370 VDD.n4533 VDD.n4070 17.3181
R10371 VDD.n4554 VDD.n4032 17.3181
R10372 VDD.n4722 VDD.n3939 17.3181
R10373 VDD.n4758 VDD.n3823 17.3181
R10374 VDD.n4443 VDD.n4442 17.3181
R10375 VDD.n4511 VDD.n4509 17.3181
R10376 VDD.n4599 VDD.n4598 17.3181
R10377 VDD.n4680 VDD.n3988 17.3181
R10378 VDD.n3849 VDD.n3848 17.3181
R10379 VDD.n4792 VDD.n4788 17.3181
R10380 VDD.n4330 VDD.n4329 17.3181
R10381 VDD.n4314 VDD.n4310 17.3181
R10382 VDD.n4609 VDD.n4041 17.3181
R10383 VDD.n4692 VDD.n3975 17.3181
R10384 VDD.n4970 VDD.n4969 17.3181
R10385 VDD.n4956 VDD.n4955 17.3181
R10386 VDD.n3204 VDD.n3180 17.3181
R10387 VDD.n3217 VDD.n3208 17.3181
R10388 VDD.n3291 VDD.n3282 17.3181
R10389 VDD.n3304 VDD.n3295 17.3181
R10390 VDD.n3317 VDD.n3308 17.3181
R10391 VDD.n3330 VDD.n3321 17.3181
R10392 VDD.n3274 VDD.n3265 17.3181
R10393 VDD.n3260 VDD.n3251 17.3181
R10394 VDD.n3246 VDD.n3237 17.3181
R10395 VDD.n3232 VDD.n3223 17.3181
R10396 VDD.n3173 VDD.n3164 17.3181
R10397 VDD.n3625 VDD.n3601 17.3181
R10398 VDD.n3638 VDD.n3629 17.3181
R10399 VDD.n3652 VDD.n3643 17.3181
R10400 VDD.n3665 VDD.n3656 17.3181
R10401 VDD.n3678 VDD.n3669 17.3181
R10402 VDD.n3691 VDD.n3682 17.3181
R10403 VDD.n3704 VDD.n3695 17.3181
R10404 VDD.n3717 VDD.n3708 17.3181
R10405 VDD.n3731 VDD.n3722 17.3181
R10406 VDD.n3744 VDD.n3735 17.3181
R10407 VDD.n3757 VDD.n3748 17.3181
R10408 VDD.n3770 VDD.n3761 17.3181
R10409 VDD.n3783 VDD.n3774 17.3181
R10410 VDD.n3584 VDD.n3575 17.3181
R10411 VDD.n3570 VDD.n3561 17.3181
R10412 VDD.n3556 VDD.n3547 17.3181
R10413 VDD.n3542 VDD.n3533 17.3181
R10414 VDD.n3528 VDD.n3519 17.3181
R10415 VDD.n3514 VDD.n3505 17.3181
R10416 VDD.n3499 VDD.n3490 17.3181
R10417 VDD.n3485 VDD.n3461 17.3181
R10418 VDD.n534 VDD.n533 17.3181
R10419 VDD.n559 VDD.n558 17.3181
R10420 VDD.n792 VDD.n791 17.3181
R10421 VDD.n805 VDD.n804 17.3181
R10422 VDD.n818 VDD.n817 17.3181
R10423 VDD.n831 VDD.n830 17.3181
R10424 VDD.n775 VDD.n774 17.3181
R10425 VDD.n761 VDD.n760 17.3181
R10426 VDD.n747 VDD.n746 17.3181
R10427 VDD.n515 VDD.n514 17.3181
R10428 VDD.n2572 VDD.n2571 17.3181
R10429 VDD.n1939 VDD.n1476 17.3181
R10430 VDD.n1960 VDD.n1438 17.3181
R10431 VDD.n2128 VDD.n1345 17.3181
R10432 VDD.n2164 VDD.n1229 17.3181
R10433 VDD.n1849 VDD.n1848 17.3181
R10434 VDD.n1917 VDD.n1915 17.3181
R10435 VDD.n2005 VDD.n2004 17.3181
R10436 VDD.n2086 VDD.n1394 17.3181
R10437 VDD.n1255 VDD.n1254 17.3181
R10438 VDD.n2198 VDD.n2194 17.3181
R10439 VDD.n1736 VDD.n1735 17.3181
R10440 VDD.n1720 VDD.n1716 17.3181
R10441 VDD.n2015 VDD.n1447 17.3181
R10442 VDD.n2098 VDD.n1381 17.3181
R10443 VDD.n2376 VDD.n2375 17.3181
R10444 VDD.n2362 VDD.n2361 17.3181
R10445 VDD.n610 VDD.n586 17.3181
R10446 VDD.n623 VDD.n614 17.3181
R10447 VDD.n697 VDD.n688 17.3181
R10448 VDD.n710 VDD.n701 17.3181
R10449 VDD.n723 VDD.n714 17.3181
R10450 VDD.n736 VDD.n727 17.3181
R10451 VDD.n680 VDD.n671 17.3181
R10452 VDD.n666 VDD.n657 17.3181
R10453 VDD.n652 VDD.n643 17.3181
R10454 VDD.n638 VDD.n629 17.3181
R10455 VDD.n579 VDD.n570 17.3181
R10456 VDD.n1031 VDD.n1007 17.3181
R10457 VDD.n1044 VDD.n1035 17.3181
R10458 VDD.n1058 VDD.n1049 17.3181
R10459 VDD.n1071 VDD.n1062 17.3181
R10460 VDD.n1084 VDD.n1075 17.3181
R10461 VDD.n1097 VDD.n1088 17.3181
R10462 VDD.n1110 VDD.n1101 17.3181
R10463 VDD.n1123 VDD.n1114 17.3181
R10464 VDD.n1137 VDD.n1128 17.3181
R10465 VDD.n1150 VDD.n1141 17.3181
R10466 VDD.n1163 VDD.n1154 17.3181
R10467 VDD.n1176 VDD.n1167 17.3181
R10468 VDD.n1189 VDD.n1180 17.3181
R10469 VDD.n990 VDD.n981 17.3181
R10470 VDD.n976 VDD.n967 17.3181
R10471 VDD.n962 VDD.n953 17.3181
R10472 VDD.n948 VDD.n939 17.3181
R10473 VDD.n934 VDD.n925 17.3181
R10474 VDD.n920 VDD.n911 17.3181
R10475 VDD.n905 VDD.n896 17.3181
R10476 VDD.n891 VDD.n867 17.3181
R10477 VDD.n6097 VDD.n6096 17.3181
R10478 VDD.n6122 VDD.n6121 17.3181
R10479 VDD.n6355 VDD.n6354 17.3181
R10480 VDD.n6368 VDD.n6367 17.3181
R10481 VDD.n6381 VDD.n6380 17.3181
R10482 VDD.n6394 VDD.n6393 17.3181
R10483 VDD.n6338 VDD.n6337 17.3181
R10484 VDD.n6324 VDD.n6323 17.3181
R10485 VDD.n6310 VDD.n6309 17.3181
R10486 VDD.n6078 VDD.n6077 17.3181
R10487 VDD.n8135 VDD.n8134 17.3181
R10488 VDD.n7502 VDD.n7039 17.3181
R10489 VDD.n7523 VDD.n7001 17.3181
R10490 VDD.n7691 VDD.n6908 17.3181
R10491 VDD.n7727 VDD.n6792 17.3181
R10492 VDD.n7412 VDD.n7411 17.3181
R10493 VDD.n7480 VDD.n7478 17.3181
R10494 VDD.n7568 VDD.n7567 17.3181
R10495 VDD.n7649 VDD.n6957 17.3181
R10496 VDD.n6818 VDD.n6817 17.3181
R10497 VDD.n7761 VDD.n7757 17.3181
R10498 VDD.n7299 VDD.n7298 17.3181
R10499 VDD.n7283 VDD.n7279 17.3181
R10500 VDD.n7578 VDD.n7010 17.3181
R10501 VDD.n7661 VDD.n6944 17.3181
R10502 VDD.n7939 VDD.n7938 17.3181
R10503 VDD.n7925 VDD.n7924 17.3181
R10504 VDD.n6173 VDD.n6149 17.3181
R10505 VDD.n6186 VDD.n6177 17.3181
R10506 VDD.n6260 VDD.n6251 17.3181
R10507 VDD.n6273 VDD.n6264 17.3181
R10508 VDD.n6286 VDD.n6277 17.3181
R10509 VDD.n6299 VDD.n6290 17.3181
R10510 VDD.n6243 VDD.n6234 17.3181
R10511 VDD.n6229 VDD.n6220 17.3181
R10512 VDD.n6215 VDD.n6206 17.3181
R10513 VDD.n6201 VDD.n6192 17.3181
R10514 VDD.n6142 VDD.n6133 17.3181
R10515 VDD.n6594 VDD.n6570 17.3181
R10516 VDD.n6607 VDD.n6598 17.3181
R10517 VDD.n6621 VDD.n6612 17.3181
R10518 VDD.n6634 VDD.n6625 17.3181
R10519 VDD.n6647 VDD.n6638 17.3181
R10520 VDD.n6660 VDD.n6651 17.3181
R10521 VDD.n6673 VDD.n6664 17.3181
R10522 VDD.n6686 VDD.n6677 17.3181
R10523 VDD.n6700 VDD.n6691 17.3181
R10524 VDD.n6713 VDD.n6704 17.3181
R10525 VDD.n6726 VDD.n6717 17.3181
R10526 VDD.n6739 VDD.n6730 17.3181
R10527 VDD.n6752 VDD.n6743 17.3181
R10528 VDD.n6553 VDD.n6544 17.3181
R10529 VDD.n6539 VDD.n6530 17.3181
R10530 VDD.n6525 VDD.n6516 17.3181
R10531 VDD.n6511 VDD.n6502 17.3181
R10532 VDD.n6497 VDD.n6488 17.3181
R10533 VDD.n6483 VDD.n6474 17.3181
R10534 VDD.n6468 VDD.n6459 17.3181
R10535 VDD.n6454 VDD.n6430 17.3181
R10536 VDD.n2652 VDD.n2622 17.2805
R10537 VDD.n2994 VDD.n2993 17.2805
R10538 VDD.n58 VDD.n28 17.2805
R10539 VDD.n400 VDD.n399 17.2805
R10540 VDD.n5621 VDD.n5591 17.2805
R10541 VDD.n5963 VDD.n5962 17.2805
R10542 VDD.n5410 VDD.n5322 17.208
R10543 VDD.n5406 VDD.n5324 16.9784
R10544 VDD.n3099 VDD.n3098 16.3958
R10545 VDD.n2989 VDD.n2942 16.3958
R10546 VDD.n505 VDD.n504 16.3958
R10547 VDD.n395 VDD.n348 16.3958
R10548 VDD.n6068 VDD.n6067 16.3958
R10549 VDD.n5958 VDD.n5911 16.3958
R10550 VDD.n5512 VDD 16.2995
R10551 VDD.n5154 VDD.n3444 15.8123
R10552 VDD.n4575 VDD.n4574 15.8123
R10553 VDD.n3942 VDD.n3941 15.8123
R10554 VDD.n4759 VDD.n4757 15.8123
R10555 VDD.n4455 VDD.n4130 15.8123
R10556 VDD.n4447 VDD.n4084 15.8123
R10557 VDD.n4596 VDD.n4595 15.8123
R10558 VDD.n4684 VDD.n4683 15.8123
R10559 VDD.n5099 VDD.n3841 15.8123
R10560 VDD.n4791 VDD.n4789 15.8123
R10561 VDD.n4327 VDD.n4326 15.8123
R10562 VDD.n4318 VDD.n4317 15.8123
R10563 VDD.n4608 VDD.n4002 15.8123
R10564 VDD.n3983 VDD.n3982 15.8123
R10565 VDD.n4967 VDD.n4966 15.8123
R10566 VDD.n4959 VDD.n4772 15.8123
R10567 VDD.n2560 VDD.n850 15.8123
R10568 VDD.n1981 VDD.n1980 15.8123
R10569 VDD.n1348 VDD.n1347 15.8123
R10570 VDD.n2165 VDD.n2163 15.8123
R10571 VDD.n1861 VDD.n1536 15.8123
R10572 VDD.n1853 VDD.n1490 15.8123
R10573 VDD.n2002 VDD.n2001 15.8123
R10574 VDD.n2090 VDD.n2089 15.8123
R10575 VDD.n2505 VDD.n1247 15.8123
R10576 VDD.n2197 VDD.n2195 15.8123
R10577 VDD.n1733 VDD.n1732 15.8123
R10578 VDD.n1724 VDD.n1723 15.8123
R10579 VDD.n2014 VDD.n1408 15.8123
R10580 VDD.n1389 VDD.n1388 15.8123
R10581 VDD.n2373 VDD.n2372 15.8123
R10582 VDD.n2365 VDD.n2178 15.8123
R10583 VDD.n5506 VDD.n5505 15.8123
R10584 VDD.n5402 VDD.n5327 15.8123
R10585 VDD.n5368 VDD.n5367 15.8123
R10586 VDD.n8123 VDD.n6413 15.8123
R10587 VDD.n7544 VDD.n7543 15.8123
R10588 VDD.n6911 VDD.n6910 15.8123
R10589 VDD.n7728 VDD.n7726 15.8123
R10590 VDD.n7424 VDD.n7099 15.8123
R10591 VDD.n7416 VDD.n7053 15.8123
R10592 VDD.n7565 VDD.n7564 15.8123
R10593 VDD.n7653 VDD.n7652 15.8123
R10594 VDD.n8068 VDD.n6810 15.8123
R10595 VDD.n7760 VDD.n7758 15.8123
R10596 VDD.n7296 VDD.n7295 15.8123
R10597 VDD.n7287 VDD.n7286 15.8123
R10598 VDD.n7577 VDD.n6971 15.8123
R10599 VDD.n6952 VDD.n6951 15.8123
R10600 VDD.n7936 VDD.n7935 15.8123
R10601 VDD.n7928 VDD.n7741 15.8123
R10602 VDD.n5363 VDD.n5339 15.7204
R10603 VDD.n5403 VDD.n5402 15.4725
R10604 VDD.n5418 VDD.n5319 14.4166
R10605 VDD.n5153 VDD.n3445 14.3064
R10606 VDD.n4553 VDD.n4552 14.3064
R10607 VDD.n5131 VDD.n3802 14.3064
R10608 VDD.n4755 VDD.n3803 14.3064
R10609 VDD.n5105 VDD.n3832 14.3064
R10610 VDD.n5105 VDD.n5104 14.3064
R10611 VDD.n4454 VDD.n4131 14.3064
R10612 VDD.n4450 VDD.n4448 14.3064
R10613 VDD.n4674 VDD.n3990 14.3064
R10614 VDD.n4675 VDD.n3987 14.3064
R10615 VDD.n5098 VDD.n3842 14.3064
R10616 VDD.n5094 VDD.n3853 14.3064
R10617 VDD.n4325 VDD.n4306 14.3064
R10618 VDD.n4321 VDD.n4308 14.3064
R10619 VDD.n4661 VDD.n4660 14.3064
R10620 VDD.n4664 VDD.n4663 14.3064
R10621 VDD.n4965 VDD.n4770 14.3064
R10622 VDD.n4961 VDD.n4960 14.3064
R10623 VDD.n2559 VDD.n851 14.3064
R10624 VDD.n1959 VDD.n1958 14.3064
R10625 VDD.n2537 VDD.n1208 14.3064
R10626 VDD.n2161 VDD.n1209 14.3064
R10627 VDD.n2511 VDD.n1238 14.3064
R10628 VDD.n2511 VDD.n2510 14.3064
R10629 VDD.n1860 VDD.n1537 14.3064
R10630 VDD.n1856 VDD.n1854 14.3064
R10631 VDD.n2080 VDD.n1396 14.3064
R10632 VDD.n2081 VDD.n1393 14.3064
R10633 VDD.n2504 VDD.n1248 14.3064
R10634 VDD.n2500 VDD.n1259 14.3064
R10635 VDD.n1731 VDD.n1712 14.3064
R10636 VDD.n1727 VDD.n1714 14.3064
R10637 VDD.n2067 VDD.n2066 14.3064
R10638 VDD.n2070 VDD.n2069 14.3064
R10639 VDD.n2371 VDD.n2176 14.3064
R10640 VDD.n2367 VDD.n2366 14.3064
R10641 VDD.n8122 VDD.n6414 14.3064
R10642 VDD.n7522 VDD.n7521 14.3064
R10643 VDD.n8100 VDD.n6771 14.3064
R10644 VDD.n7724 VDD.n6772 14.3064
R10645 VDD.n8074 VDD.n6801 14.3064
R10646 VDD.n8074 VDD.n8073 14.3064
R10647 VDD.n7423 VDD.n7100 14.3064
R10648 VDD.n7419 VDD.n7417 14.3064
R10649 VDD.n7643 VDD.n6959 14.3064
R10650 VDD.n7644 VDD.n6956 14.3064
R10651 VDD.n8067 VDD.n6811 14.3064
R10652 VDD.n8063 VDD.n6822 14.3064
R10653 VDD.n7294 VDD.n7275 14.3064
R10654 VDD.n7290 VDD.n7277 14.3064
R10655 VDD.n7630 VDD.n7629 14.3064
R10656 VDD.n7633 VDD.n7632 14.3064
R10657 VDD.n7934 VDD.n7739 14.3064
R10658 VDD.n7930 VDD.n7929 14.3064
R10659 VDD.n4248 VDD.n4200 13.6005
R10660 VDD.n4254 VDD.n4196 13.6005
R10661 VDD.n4260 VDD.n4192 13.6005
R10662 VDD.n4267 VDD.n4188 13.6005
R10663 VDD.n4267 VDD.n4266 13.6005
R10664 VDD.n4273 VDD.n4184 13.6005
R10665 VDD.n4280 VDD.n4279 13.6005
R10666 VDD.n4286 VDD.n4174 13.6005
R10667 VDD.n4292 VDD.n4174 13.6005
R10668 VDD.n4299 VDD.n4170 13.6005
R10669 VDD.n4344 VDD.n4165 13.6005
R10670 VDD.n4354 VDD.n4151 13.6005
R10671 VDD.n4942 VDD.n4781 13.6005
R10672 VDD.n4936 VDD.n4935 13.6005
R10673 VDD.n4934 VDD.n4810 13.6005
R10674 VDD.n4928 VDD.n4810 13.6005
R10675 VDD.n4927 VDD.n4926 13.6005
R10676 VDD.n4920 VDD.n4820 13.6005
R10677 VDD.n4919 VDD.n4918 13.6005
R10678 VDD.n4918 VDD.n4824 13.6005
R10679 VDD.n4912 VDD.n4911 13.6005
R10680 VDD.n4910 VDD.n4831 13.6005
R10681 VDD.n4904 VDD.n4903 13.6005
R10682 VDD.n1654 VDD.n1606 13.6005
R10683 VDD.n1660 VDD.n1602 13.6005
R10684 VDD.n1666 VDD.n1598 13.6005
R10685 VDD.n1673 VDD.n1594 13.6005
R10686 VDD.n1673 VDD.n1672 13.6005
R10687 VDD.n1679 VDD.n1590 13.6005
R10688 VDD.n1686 VDD.n1685 13.6005
R10689 VDD.n1692 VDD.n1580 13.6005
R10690 VDD.n1698 VDD.n1580 13.6005
R10691 VDD.n1705 VDD.n1576 13.6005
R10692 VDD.n1750 VDD.n1571 13.6005
R10693 VDD.n1760 VDD.n1557 13.6005
R10694 VDD.n2348 VDD.n2187 13.6005
R10695 VDD.n2342 VDD.n2341 13.6005
R10696 VDD.n2340 VDD.n2216 13.6005
R10697 VDD.n2334 VDD.n2216 13.6005
R10698 VDD.n2333 VDD.n2332 13.6005
R10699 VDD.n2326 VDD.n2226 13.6005
R10700 VDD.n2325 VDD.n2324 13.6005
R10701 VDD.n2324 VDD.n2230 13.6005
R10702 VDD.n2318 VDD.n2317 13.6005
R10703 VDD.n2316 VDD.n2237 13.6005
R10704 VDD.n2310 VDD.n2309 13.6005
R10705 VDD.n7217 VDD.n7169 13.6005
R10706 VDD.n7223 VDD.n7165 13.6005
R10707 VDD.n7229 VDD.n7161 13.6005
R10708 VDD.n7236 VDD.n7157 13.6005
R10709 VDD.n7236 VDD.n7235 13.6005
R10710 VDD.n7242 VDD.n7153 13.6005
R10711 VDD.n7249 VDD.n7248 13.6005
R10712 VDD.n7255 VDD.n7143 13.6005
R10713 VDD.n7261 VDD.n7143 13.6005
R10714 VDD.n7268 VDD.n7139 13.6005
R10715 VDD.n7313 VDD.n7134 13.6005
R10716 VDD.n7323 VDD.n7120 13.6005
R10717 VDD.n7911 VDD.n7750 13.6005
R10718 VDD.n7905 VDD.n7904 13.6005
R10719 VDD.n7903 VDD.n7779 13.6005
R10720 VDD.n7897 VDD.n7779 13.6005
R10721 VDD.n7896 VDD.n7895 13.6005
R10722 VDD.n7889 VDD.n7789 13.6005
R10723 VDD.n7888 VDD.n7887 13.6005
R10724 VDD.n7887 VDD.n7793 13.6005
R10725 VDD.n7881 VDD.n7880 13.6005
R10726 VDD.n7879 VDD.n7800 13.6005
R10727 VDD.n7873 VDD.n7872 13.6005
R10728 VDD.n5538 VDD.n5469 13.4622
R10729 VDD.n4478 VDD.n4094 13.4005
R10730 VDD.n4539 VDD.n3440 13.4005
R10731 VDD.n4043 VDD.n4023 13.4005
R10732 VDD.t629 VDD.n4006 13.4005
R10733 VDD.n4706 VDD.n3958 13.4005
R10734 VDD.n3920 VDD.n3810 13.4005
R10735 VDD.n5092 VDD.n3855 13.4005
R10736 VDD.n5073 VDD.n3889 13.4005
R10737 VDD.n1884 VDD.n1500 13.4005
R10738 VDD.n1945 VDD.n846 13.4005
R10739 VDD.n1449 VDD.n1429 13.4005
R10740 VDD.t10 VDD.n1412 13.4005
R10741 VDD.n2112 VDD.n1364 13.4005
R10742 VDD.n1326 VDD.n1216 13.4005
R10743 VDD.n2498 VDD.n1261 13.4005
R10744 VDD.n2479 VDD.n1295 13.4005
R10745 VDD.n7447 VDD.n7063 13.4005
R10746 VDD.n7508 VDD.n6409 13.4005
R10747 VDD.n7012 VDD.n6992 13.4005
R10748 VDD.t316 VDD.n6975 13.4005
R10749 VDD.n7675 VDD.n6927 13.4005
R10750 VDD.n6889 VDD.n6779 13.4005
R10751 VDD.n8061 VDD.n6824 13.4005
R10752 VDD.n8042 VDD.n6858 13.4005
R10753 VDD.n3058 VDD.t503 13.2488
R10754 VDD.n2706 VDD.t505 13.2488
R10755 VDD.n464 VDD.t31 13.2488
R10756 VDD.n112 VDD.t29 13.2488
R10757 VDD.n6027 VDD.t200 13.2488
R10758 VDD.n5675 VDD.t210 13.2488
R10759 VDD.n5422 VDD.n5317 13.2137
R10760 VDD.n4698 VDD.t597 13.2005
R10761 VDD.n2104 VDD.t12 13.2005
R10762 VDD.n7667 VDD.t183 13.2005
R10763 VDD.n5432 VDD.n5431 13.177
R10764 VDD.n5392 VDD.n5391 13.0943
R10765 VDD.n5147 VDD.t589 13.0005
R10766 VDD.n2553 VDD.t701 13.0005
R10767 VDD.n8116 VDD.t176 13.0005
R10768 VDD.n4551 VDD.n3445 12.8005
R10769 VDD.n4552 VDD.n4551 12.8005
R10770 VDD.n5131 VDD.n5130 12.8005
R10771 VDD.n5130 VDD.n3803 12.8005
R10772 VDD.n4739 VDD.t619 12.8005
R10773 VDD.n4451 VDD.n4131 12.8005
R10774 VDD.n4451 VDD.n4450 12.8005
R10775 VDD.n4676 VDD.n4674 12.8005
R10776 VDD.n4676 VDD.n4675 12.8005
R10777 VDD.n5095 VDD.n3842 12.8005
R10778 VDD.n5095 VDD.n5094 12.8005
R10779 VDD.n4322 VDD.n4306 12.8005
R10780 VDD.n4322 VDD.n4321 12.8005
R10781 VDD.n4662 VDD.n4661 12.8005
R10782 VDD.n4663 VDD.n4662 12.8005
R10783 VDD.n4962 VDD.n4770 12.8005
R10784 VDD.n4962 VDD.n4961 12.8005
R10785 VDD.n1957 VDD.n851 12.8005
R10786 VDD.n1958 VDD.n1957 12.8005
R10787 VDD.n2537 VDD.n2536 12.8005
R10788 VDD.n2536 VDD.n1209 12.8005
R10789 VDD.n2145 VDD.t324 12.8005
R10790 VDD.n1857 VDD.n1537 12.8005
R10791 VDD.n1857 VDD.n1856 12.8005
R10792 VDD.n2082 VDD.n2080 12.8005
R10793 VDD.n2082 VDD.n2081 12.8005
R10794 VDD.n2501 VDD.n1248 12.8005
R10795 VDD.n2501 VDD.n2500 12.8005
R10796 VDD.n1728 VDD.n1712 12.8005
R10797 VDD.n1728 VDD.n1727 12.8005
R10798 VDD.n2068 VDD.n2067 12.8005
R10799 VDD.n2069 VDD.n2068 12.8005
R10800 VDD.n2368 VDD.n2176 12.8005
R10801 VDD.n2368 VDD.n2367 12.8005
R10802 VDD.n7520 VDD.n6414 12.8005
R10803 VDD.n7521 VDD.n7520 12.8005
R10804 VDD.n8100 VDD.n8099 12.8005
R10805 VDD.n8099 VDD.n6772 12.8005
R10806 VDD.n7708 VDD.t370 12.8005
R10807 VDD.n7420 VDD.n7100 12.8005
R10808 VDD.n7420 VDD.n7419 12.8005
R10809 VDD.n7645 VDD.n7643 12.8005
R10810 VDD.n7645 VDD.n7644 12.8005
R10811 VDD.n8064 VDD.n6811 12.8005
R10812 VDD.n8064 VDD.n8063 12.8005
R10813 VDD.n7291 VDD.n7275 12.8005
R10814 VDD.n7291 VDD.n7290 12.8005
R10815 VDD.n7631 VDD.n7630 12.8005
R10816 VDD.n7632 VDD.n7631 12.8005
R10817 VDD.n7931 VDD.n7739 12.8005
R10818 VDD.n7931 VDD.n7930 12.8005
R10819 VDD.n4107 VDD.t603 12.6005
R10820 VDD.n1513 VDD.t498 12.6005
R10821 VDD.n7076 VDD.t561 12.6005
R10822 VDD.n5491 VDD.n5490 12.424
R10823 VDD.n4458 VDD.t429 12.4005
R10824 VDD.t615 VDD.n3838 12.4005
R10825 VDD.n1864 VDD.t99 12.4005
R10826 VDD.t454 VDD.n1244 12.4005
R10827 VDD.n7427 VDD.t38 12.4005
R10828 VDD.t181 VDD.n6807 12.4005
R10829 VDD.t653 VDD.n4138 12.2005
R10830 VDD.n3917 VDD.t424 12.2005
R10831 VDD.t452 VDD.n1544 12.2005
R10832 VDD.n1323 VDD.t146 12.2005
R10833 VDD.t373 VDD.n7107 12.2005
R10834 VDD.n6886 VDD.t22 12.2005
R10835 VDD.n4536 VDD.t413 12.0005
R10836 VDD.n5030 VDD.t635 12.0005
R10837 VDD.n1942 VDD.t334 12.0005
R10838 VDD.n2436 VDD.t189 12.0005
R10839 VDD.n7505 VDD.t2 12.0005
R10840 VDD.n7999 VDD.t341 12.0005
R10841 VDD.t631 VDD.n4170 11.8005
R10842 VDD.n5115 VDD.t427 11.8005
R10843 VDD.n4935 VDD.t633 11.8005
R10844 VDD.t97 VDD.n1576 11.8005
R10845 VDD.n2521 VDD.t195 11.8005
R10846 VDD.n2341 VDD.t501 11.8005
R10847 VDD.t156 VDD.n7139 11.8005
R10848 VDD.n8084 VDD.t216 11.8005
R10849 VDD.n7904 VDD.t268 11.8005
R10850 VDD.n4619 VDD.t398 11.6005
R10851 VDD.n2025 VDD.t81 11.6005
R10852 VDD.n7588 VDD.t230 11.6005
R10853 VDD.n4260 VDD.t621 11.4005
R10854 VDD.n4273 VDD.t609 11.4005
R10855 VDD.t410 VDD.n3933 11.4005
R10856 VDD.n4920 VDD.t661 11.4005
R10857 VDD.n4912 VDD.t641 11.4005
R10858 VDD.n1666 VDD.t6 11.4005
R10859 VDD.n1679 VDD.t174 11.4005
R10860 VDD.t52 VDD.n1339 11.4005
R10861 VDD.n2326 VDD.t221 11.4005
R10862 VDD.n2318 VDD.t36 11.4005
R10863 VDD.n7229 VDD.t158 11.4005
R10864 VDD.n7242 VDD.t8 11.4005
R10865 VDD.t579 VDD.n6902 11.4005
R10866 VDD.n7889 VDD.t509 11.4005
R10867 VDD.n7881 VDD.t283 11.4005
R10868 VDD.n5542 VDD.n5467 11.3631
R10869 VDD.n4494 VDD.n4100 11.2946
R10870 VDD.n5154 VDD.n5153 11.2946
R10871 VDD.n4575 VDD.n4553 11.2946
R10872 VDD.n3941 VDD.n3802 11.2946
R10873 VDD.n4757 VDD.n4755 11.2946
R10874 VDD.n4495 VDD.n4494 11.2946
R10875 VDD.n4455 VDD.n4454 11.2946
R10876 VDD.n4448 VDD.n4447 11.2946
R10877 VDD.n4595 VDD.n3990 11.2946
R10878 VDD.n4684 VDD.n3987 11.2946
R10879 VDD.n5099 VDD.n5098 11.2946
R10880 VDD.n4789 VDD.n3853 11.2946
R10881 VDD.n4326 VDD.n4325 11.2946
R10882 VDD.n4318 VDD.n4308 11.2946
R10883 VDD.n4660 VDD.n4002 11.2946
R10884 VDD.n4664 VDD.n3983 11.2946
R10885 VDD.n4966 VDD.n4965 11.2946
R10886 VDD.n4960 VDD.n4959 11.2946
R10887 VDD.n1900 VDD.n1506 11.2946
R10888 VDD.n2560 VDD.n2559 11.2946
R10889 VDD.n1981 VDD.n1959 11.2946
R10890 VDD.n1347 VDD.n1208 11.2946
R10891 VDD.n2163 VDD.n2161 11.2946
R10892 VDD.n1901 VDD.n1900 11.2946
R10893 VDD.n1861 VDD.n1860 11.2946
R10894 VDD.n1854 VDD.n1853 11.2946
R10895 VDD.n2001 VDD.n1396 11.2946
R10896 VDD.n2090 VDD.n1393 11.2946
R10897 VDD.n2505 VDD.n2504 11.2946
R10898 VDD.n2195 VDD.n1259 11.2946
R10899 VDD.n1732 VDD.n1731 11.2946
R10900 VDD.n1724 VDD.n1714 11.2946
R10901 VDD.n2066 VDD.n1408 11.2946
R10902 VDD.n2070 VDD.n1389 11.2946
R10903 VDD.n2372 VDD.n2371 11.2946
R10904 VDD.n2366 VDD.n2365 11.2946
R10905 VDD.n7463 VDD.n7069 11.2946
R10906 VDD.n8123 VDD.n8122 11.2946
R10907 VDD.n7544 VDD.n7522 11.2946
R10908 VDD.n6910 VDD.n6771 11.2946
R10909 VDD.n7726 VDD.n7724 11.2946
R10910 VDD.n7464 VDD.n7463 11.2946
R10911 VDD.n7424 VDD.n7423 11.2946
R10912 VDD.n7417 VDD.n7416 11.2946
R10913 VDD.n7564 VDD.n6959 11.2946
R10914 VDD.n7653 VDD.n6956 11.2946
R10915 VDD.n8068 VDD.n8067 11.2946
R10916 VDD.n7758 VDD.n6822 11.2946
R10917 VDD.n7295 VDD.n7294 11.2946
R10918 VDD.n7287 VDD.n7277 11.2946
R10919 VDD.n7629 VDD.n6971 11.2946
R10920 VDD.n7633 VDD.n6952 11.2946
R10921 VDD.n7935 VDD.n7934 11.2946
R10922 VDD.n7929 VDD.n7928 11.2946
R10923 VDD.n3984 VDD.t419 11.2005
R10924 VDD.n1390 VDD.t148 11.2005
R10925 VDD.n6953 VDD.t141 11.2005
R10926 VDD.t645 VDD.n4196 11.0005
R10927 VDD.n4279 VDD.t649 11.0005
R10928 VDD.n4020 VDD.t431 11.0005
R10929 VDD.t595 VDD.n4927 11.0005
R10930 VDD.t623 VDD.n4831 11.0005
R10931 VDD.t79 VDD.n1602 11.0005
R10932 VDD.n1685 VDD.t4 11.0005
R10933 VDD.n1426 VDD.t193 11.0005
R10934 VDD.t357 VDD.n2333 11.0005
R10935 VDD.t516 VDD.n2237 11.0005
R10936 VDD.t255 VDD.n7165 11.0005
R10937 VDD.n7248 VDD.t264 11.0005
R10938 VDD.n6989 VDD.t48 11.0005
R10939 VDD.t322 VDD.n7896 11.0005
R10940 VDD.t179 VDD.n7800 11.0005
R10941 VDD.n5237 VDD.n5193 10.8829
R10942 VDD.n5192 VDD.n5190 10.8829
R10943 VDD.n5231 VDD.n5192 10.8829
R10944 VDD.n5229 VDD.n5228 10.8829
R10945 VDD.n5230 VDD.n5229 10.8829
R10946 VDD.n5226 VDD.n5225 10.8829
R10947 VDD.n5213 VDD.n5212 10.8829
R10948 VDD.n5210 VDD.n5209 10.8829
R10949 VDD.n5299 VDD.n5298 10.8829
R10950 VDD.n5296 VDD.n5295 10.8829
R10951 VDD.n5297 VDD.n5296 10.8829
R10952 VDD.n5286 VDD.n5285 10.8829
R10953 VDD.n5285 VDD.n5253 10.8829
R10954 VDD.n5283 VDD.n5282 10.8829
R10955 VDD.n5273 VDD.n5272 10.8829
R10956 VDD.n5270 VDD.n5269 10.8829
R10957 VDD.n5133 VDD.t394 10.8005
R10958 VDD.n2539 VDD.t89 10.8005
R10959 VDD.n8102 VDD.t165 10.8005
R10960 VDD.n4344 VDD.t605 10.6005
R10961 VDD.n4059 VDD.t405 10.6005
R10962 VDD.n4942 VDD.t613 10.6005
R10963 VDD.n1750 VDD.t348 10.6005
R10964 VDD.n1465 VDD.t91 10.6005
R10965 VDD.n2348 VDD.t336 10.6005
R10966 VDD.n7313 VDD.t207 10.6005
R10967 VDD.n7028 VDD.t0 10.6005
R10968 VDD.n7911 VDD.t318 10.6005
R10969 VDD.n5102 VDD.t437 10.4005
R10970 VDD.n2508 VDD.t360 10.4005
R10971 VDD.n8071 VDD.t61 10.4005
R10972 VDD.n4507 VDD.t421 10.2005
R10973 VDD.t599 VDD.n3867 10.2005
R10974 VDD.n1913 VDD.t95 10.2005
R10975 VDD.t346 VDD.n1273 10.2005
R10976 VDD.n7476 VDD.t43 10.2005
R10977 VDD.t40 VDD.n6836 10.2005
R10978 VDD.n5381 VDD.n5333 10.1652
R10979 VDD.n4472 VDD.t625 10.0005
R10980 VDD.n5079 VDD.t402 10.0005
R10981 VDD.n1878 VDD.t468 10.0005
R10982 VDD.n2485 VDD.t228 10.0005
R10983 VDD.n7441 VDD.t167 10.0005
R10984 VDD.n8048 VDD.t152 10.0005
R10985 VDD.t400 VDD.n4121 9.8005
R10986 VDD.n4976 VDD.t601 9.8005
R10987 VDD.t50 VDD.n1527 9.8005
R10988 VDD.n2382 VDD.t246 9.8005
R10989 VDD.t297 VDD.n7090 9.8005
R10990 VDD.n7945 VDD.t559 9.8005
R10991 VDD.n4070 VDD.n3444 9.78874
R10992 VDD.n4574 VDD.n4554 9.78874
R10993 VDD.n3942 VDD.n3939 9.78874
R10994 VDD.n4759 VDD.n4758 9.78874
R10995 VDD.n4442 VDD.n4130 9.78874
R10996 VDD.n4509 VDD.n4084 9.78874
R10997 VDD.n4598 VDD.n4596 9.78874
R10998 VDD.n4683 VDD.n3988 9.78874
R10999 VDD.n3848 VDD.n3841 9.78874
R11000 VDD.n4792 VDD.n4791 9.78874
R11001 VDD.n4329 VDD.n4327 9.78874
R11002 VDD.n4317 VDD.n4310 9.78874
R11003 VDD.n4609 VDD.n4608 9.78874
R11004 VDD.n3982 VDD.n3975 9.78874
R11005 VDD.n4969 VDD.n4967 9.78874
R11006 VDD.n4956 VDD.n4772 9.78874
R11007 VDD.n1476 VDD.n850 9.78874
R11008 VDD.n1980 VDD.n1960 9.78874
R11009 VDD.n1348 VDD.n1345 9.78874
R11010 VDD.n2165 VDD.n2164 9.78874
R11011 VDD.n1848 VDD.n1536 9.78874
R11012 VDD.n1915 VDD.n1490 9.78874
R11013 VDD.n2004 VDD.n2002 9.78874
R11014 VDD.n2089 VDD.n1394 9.78874
R11015 VDD.n1254 VDD.n1247 9.78874
R11016 VDD.n2198 VDD.n2197 9.78874
R11017 VDD.n1735 VDD.n1733 9.78874
R11018 VDD.n1723 VDD.n1716 9.78874
R11019 VDD.n2015 VDD.n2014 9.78874
R11020 VDD.n1388 VDD.n1381 9.78874
R11021 VDD.n2375 VDD.n2373 9.78874
R11022 VDD.n2362 VDD.n2178 9.78874
R11023 VDD.n5552 VDD.n5442 9.78874
R11024 VDD.n5529 VDD.n5469 9.78874
R11025 VDD.n5494 VDD.n5493 9.78874
R11026 VDD.n5417 VDD.n5313 9.78874
R11027 VDD.n5398 VDD.n5397 9.78874
R11028 VDD.n5372 VDD.n5371 9.78874
R11029 VDD.n5358 VDD.n5343 9.78874
R11030 VDD.n7039 VDD.n6413 9.78874
R11031 VDD.n7543 VDD.n7523 9.78874
R11032 VDD.n6911 VDD.n6908 9.78874
R11033 VDD.n7728 VDD.n7727 9.78874
R11034 VDD.n7411 VDD.n7099 9.78874
R11035 VDD.n7478 VDD.n7053 9.78874
R11036 VDD.n7567 VDD.n7565 9.78874
R11037 VDD.n7652 VDD.n6957 9.78874
R11038 VDD.n6817 VDD.n6810 9.78874
R11039 VDD.n7761 VDD.n7760 9.78874
R11040 VDD.n7298 VDD.n7296 9.78874
R11041 VDD.n7286 VDD.n7279 9.78874
R11042 VDD.n7578 VDD.n7577 9.78874
R11043 VDD.n6951 VDD.n6944 9.78874
R11044 VDD.n7938 VDD.n7936 9.78874
R11045 VDD.n7925 VDD.n7741 9.78874
R11046 VDD.n5567 VDD.n5566 9.6955
R11047 VDD.n4078 VDD.t593 9.6005
R11048 VDD.n1484 VDD.t534 9.6005
R11049 VDD.n7047 VDD.t27 9.6005
R11050 VDD.n5479 VDD.n5475 9.52254
R11051 VDD.n4953 VDD.n4776 9.49615
R11052 VDD.n4798 VDD.n4797 9.49615
R11053 VDD.n4350 VDD.n4132 9.49615
R11054 VDD.n4332 VDD.n4303 9.49615
R11055 VDD.n2359 VDD.n2182 9.49615
R11056 VDD.n2204 VDD.n2203 9.49615
R11057 VDD.n1756 VDD.n1538 9.49615
R11058 VDD.n1738 VDD.n1709 9.49615
R11059 VDD.n7922 VDD.n7745 9.49615
R11060 VDD.n7767 VDD.n7766 9.49615
R11061 VDD.n7319 VDD.n7101 9.49615
R11062 VDD.n7301 VDD.n7272 9.49615
R11063 VDD.n5457 VDD.n5445 9.41227
R11064 VDD.n5546 VDD.n5544 9.41227
R11065 VDD.n5413 VDD.n5412 9.41227
R11066 VDD.n4716 VDD.t591 9.4005
R11067 VDD.n2122 VDD.t240 9.4005
R11068 VDD.n7685 VDD.t225 9.4005
R11069 VDD.n5208 VDD.n5207 9.338
R11070 VDD.n5268 VDD.n5267 9.338
R11071 VDD.n2942 VDD.n2941 9.30448
R11072 VDD.n3100 VDD.n3099 9.30448
R11073 VDD.n348 VDD.n347 9.30448
R11074 VDD.n506 VDD.n505 9.30448
R11075 VDD.n5911 VDD.n5910 9.30448
R11076 VDD.n6069 VDD.n6068 9.30448
R11077 VDD.n5198 VDD.n5197 9.30104
R11078 VDD.n2609 VDD.n2608 9.3005
R11079 VDD.n2611 VDD.n2610 9.3005
R11080 VDD.n2602 VDD.n2601 9.3005
R11081 VDD.n2617 VDD.n2616 9.3005
R11082 VDD.n2928 VDD.n2927 9.3005
R11083 VDD.n2930 VDD.n2929 9.3005
R11084 VDD.n2921 VDD.n2920 9.3005
R11085 VDD.n2936 VDD.n2935 9.3005
R11086 VDD.n2911 VDD.n2910 9.3005
R11087 VDD.n2905 VDD.n2904 9.3005
R11088 VDD.n2744 VDD.n2743 9.3005
R11089 VDD.n2752 VDD.n2748 9.3005
R11090 VDD.n2657 VDD.n2620 9.3005
R11091 VDD.n2652 VDD.n2621 9.3005
R11092 VDD.n2995 VDD.n2994 9.3005
R11093 VDD.n2997 VDD.n2996 9.3005
R11094 VDD.n2903 VDD.n2902 9.3005
R11095 VDD.n2771 VDD.n2747 9.3005
R11096 VDD.n2755 VDD.n2754 9.3005
R11097 VDD.n2797 VDD.n2785 9.3005
R11098 VDD.n2824 VDD.n2823 9.3005
R11099 VDD.n2817 VDD.n2816 9.3005
R11100 VDD.n2835 VDD.n2834 9.3005
R11101 VDD.n2826 VDD.n2825 9.3005
R11102 VDD.n2832 VDD.n2783 9.3005
R11103 VDD.n2796 VDD.n2795 9.3005
R11104 VDD.n3140 VDD.n3139 9.3005
R11105 VDD.n3124 VDD.n3122 9.3005
R11106 VDD.n3146 VDD.n3145 9.3005
R11107 VDD.n3132 VDD.n3121 9.3005
R11108 VDD.n3131 VDD.n3130 9.3005
R11109 VDD.n3129 VDD.n3128 9.3005
R11110 VDD.n3158 VDD.n3149 9.3005
R11111 VDD.n3156 VDD.n3155 9.3005
R11112 VDD.n3154 VDD.n3153 9.3005
R11113 VDD.n3391 VDD.n3382 9.3005
R11114 VDD.n3389 VDD.n3388 9.3005
R11115 VDD.n3387 VDD.n3386 9.3005
R11116 VDD.n3404 VDD.n3395 9.3005
R11117 VDD.n3402 VDD.n3401 9.3005
R11118 VDD.n3400 VDD.n3399 9.3005
R11119 VDD.n3417 VDD.n3408 9.3005
R11120 VDD.n3415 VDD.n3414 9.3005
R11121 VDD.n3413 VDD.n3412 9.3005
R11122 VDD.n3430 VDD.n3421 9.3005
R11123 VDD.n3428 VDD.n3427 9.3005
R11124 VDD.n3426 VDD.n3425 9.3005
R11125 VDD.n3374 VDD.n3365 9.3005
R11126 VDD.n3372 VDD.n3371 9.3005
R11127 VDD.n3370 VDD.n3369 9.3005
R11128 VDD.n3360 VDD.n3351 9.3005
R11129 VDD.n3358 VDD.n3357 9.3005
R11130 VDD.n3356 VDD.n3355 9.3005
R11131 VDD.n3346 VDD.n3337 9.3005
R11132 VDD.n3344 VDD.n3343 9.3005
R11133 VDD.n3342 VDD.n3341 9.3005
R11134 VDD.n3114 VDD.n3105 9.3005
R11135 VDD.n3112 VDD.n3111 9.3005
R11136 VDD.n3110 VDD.n3109 9.3005
R11137 VDD.n5171 VDD.n5162 9.3005
R11138 VDD.n5169 VDD.n5168 9.3005
R11139 VDD.n5167 VDD.n5166 9.3005
R11140 VDD.n4452 VDD.n4451 9.3005
R11141 VDD.n4448 VDD.n4446 9.3005
R11142 VDD.n4084 VDD.n4083 9.3005
R11143 VDD.n4512 VDD.n4511 9.3005
R11144 VDD.n4513 VDD.n4081 9.3005
R11145 VDD.n4522 VDD.n4521 9.3005
R11146 VDD.n4520 VDD.n4519 9.3005
R11147 VDD.n4516 VDD.n4514 9.3005
R11148 VDD.n3457 VDD.n3455 9.3005
R11149 VDD.n4677 VDD.n4676 9.3005
R11150 VDD.n4678 VDD.n3987 9.3005
R11151 VDD.n4683 VDD.n4682 9.3005
R11152 VDD.n4681 VDD.n4680 9.3005
R11153 VDD.n3956 VDD.n3955 9.3005
R11154 VDD.n4710 VDD.n4709 9.3005
R11155 VDD.n4712 VDD.n4711 9.3005
R11156 VDD.n4713 VDD.n3790 9.3005
R11157 VDD.n5138 VDD.n5137 9.3005
R11158 VDD.n5096 VDD.n5095 9.3005
R11159 VDD.n3853 VDD.n3852 9.3005
R11160 VDD.n4791 VDD.n4790 9.3005
R11161 VDD.n4788 VDD.n4787 9.3005
R11162 VDD.n4797 VDD.n4796 9.3005
R11163 VDD.n4133 VDD.n4132 9.3005
R11164 VDD.n4444 VDD.n4443 9.3005
R11165 VDD.n4445 VDD.n4130 9.3005
R11166 VDD.n4454 VDD.n4453 9.3005
R11167 VDD.n5143 VDD.n5142 9.3005
R11168 VDD.n4048 VDD.n3458 9.3005
R11169 VDD.n4592 VDD.n4591 9.3005
R11170 VDD.n4593 VDD.n4046 9.3005
R11171 VDD.n4602 VDD.n4601 9.3005
R11172 VDD.n4600 VDD.n4599 9.3005
R11173 VDD.n4596 VDD.n4594 9.3005
R11174 VDD.n3990 VDD.n3989 9.3005
R11175 VDD.n3812 VDD.n3791 9.3005
R11176 VDD.n5121 VDD.n5120 9.3005
R11177 VDD.n5119 VDD.n5118 9.3005
R11178 VDD.n3815 VDD.n3814 9.3005
R11179 VDD.n3845 VDD.n3843 9.3005
R11180 VDD.n3850 VDD.n3849 9.3005
R11181 VDD.n3851 VDD.n3841 9.3005
R11182 VDD.n5098 VDD.n5097 9.3005
R11183 VDD.n4963 VDD.n4962 9.3005
R11184 VDD.n4960 VDD.n4771 9.3005
R11185 VDD.n4775 VDD.n4772 9.3005
R11186 VDD.n4955 VDD.n4954 9.3005
R11187 VDD.n4953 VDD.n4952 9.3005
R11188 VDD.n4965 VDD.n4964 9.3005
R11189 VDD.n4967 VDD.n4767 9.3005
R11190 VDD.n4971 VDD.n4970 9.3005
R11191 VDD.n4973 VDD.n4972 9.3005
R11192 VDD.n4323 VDD.n4322 9.3005
R11193 VDD.n4308 VDD.n4307 9.3005
R11194 VDD.n4317 VDD.n4316 9.3005
R11195 VDD.n4315 VDD.n4314 9.3005
R11196 VDD.n4312 VDD.n4311 9.3005
R11197 VDD.n4325 VDD.n4324 9.3005
R11198 VDD.n4327 VDD.n4305 9.3005
R11199 VDD.n4331 VDD.n4330 9.3005
R11200 VDD.n4333 VDD.n4332 9.3005
R11201 VDD.n4551 VDD.n3447 9.3005
R11202 VDD.n4562 VDD.n4553 9.3005
R11203 VDD.n4574 VDD.n4573 9.3005
R11204 VDD.n4556 VDD.n4032 9.3005
R11205 VDD.n4616 VDD.n4615 9.3005
R11206 VDD.n4037 VDD.n4036 9.3005
R11207 VDD.n4039 VDD.n4004 9.3005
R11208 VDD.n4657 VDD.n4656 9.3005
R11209 VDD.n4658 VDD.n3998 9.3005
R11210 VDD.n5130 VDD.n5129 9.3005
R11211 VDD.n4755 VDD.n3805 9.3005
R11212 VDD.n4760 VDD.n4759 9.3005
R11213 VDD.n4765 VDD.n3823 9.3005
R11214 VDD.n4076 VDD.n4071 9.3005
R11215 VDD.n4531 VDD.n4530 9.3005
R11216 VDD.n4074 VDD.n3446 9.3005
R11217 VDD.n5151 VDD.n5150 9.3005
R11218 VDD.n4662 VDD.n4000 9.3005
R11219 VDD.n4665 VDD.n4664 9.3005
R11220 VDD.n3982 VDD.n3971 9.3005
R11221 VDD.n4693 VDD.n4692 9.3005
R11222 VDD.n3980 VDD.n3979 9.3005
R11223 VDD.n3976 VDD.n3940 9.3005
R11224 VDD.n4720 VDD.n4719 9.3005
R11225 VDD.n4557 VDD.n3945 9.3005
R11226 VDD.n3948 VDD.n3804 9.3005
R11227 VDD.n4533 VDD.n4532 9.3005
R11228 VDD.n4072 VDD.n3444 9.3005
R11229 VDD.n5153 VDD.n5152 9.3005
R11230 VDD.n4667 VDD.n4666 9.3005
R11231 VDD.n4001 VDD.n3969 9.3005
R11232 VDD.n4695 VDD.n4694 9.3005
R11233 VDD.n3974 VDD.n3973 9.3005
R11234 VDD.n3978 VDD.n3938 9.3005
R11235 VDD.n4722 VDD.n4721 9.3005
R11236 VDD.n3943 VDD.n3942 9.3005
R11237 VDD.n4558 VDD.n3802 9.3005
R11238 VDD.n4766 VDD.n4752 9.3005
R11239 VDD.n4764 VDD.n4763 9.3005
R11240 VDD.n4754 VDD.n3807 9.3005
R11241 VDD.n5128 VDD.n5127 9.3005
R11242 VDD.n4660 VDD.n4659 9.3005
R11243 VDD.n4608 VDD.n4003 9.3005
R11244 VDD.n4041 VDD.n4040 9.3005
R11245 VDD.n4614 VDD.n4613 9.3005
R11246 VDD.n4569 VDD.n4034 9.3005
R11247 VDD.n4572 VDD.n4571 9.3005
R11248 VDD.n4567 VDD.n4555 9.3005
R11249 VDD.n4564 VDD.n4563 9.3005
R11250 VDD.n3199 VDD.n3198 9.3005
R11251 VDD.n3182 VDD.n3181 9.3005
R11252 VDD.n3205 VDD.n3204 9.3005
R11253 VDD.n3186 VDD.n3185 9.3005
R11254 VDD.n3194 VDD.n3193 9.3005
R11255 VDD.n3196 VDD.n3195 9.3005
R11256 VDD.n3213 VDD.n3212 9.3005
R11257 VDD.n3210 VDD.n3209 9.3005
R11258 VDD.n3218 VDD.n3217 9.3005
R11259 VDD.n3287 VDD.n3286 9.3005
R11260 VDD.n3284 VDD.n3283 9.3005
R11261 VDD.n3292 VDD.n3291 9.3005
R11262 VDD.n3300 VDD.n3299 9.3005
R11263 VDD.n3297 VDD.n3296 9.3005
R11264 VDD.n3305 VDD.n3304 9.3005
R11265 VDD.n3313 VDD.n3312 9.3005
R11266 VDD.n3310 VDD.n3309 9.3005
R11267 VDD.n3318 VDD.n3317 9.3005
R11268 VDD.n3326 VDD.n3325 9.3005
R11269 VDD.n3323 VDD.n3322 9.3005
R11270 VDD.n3331 VDD.n3330 9.3005
R11271 VDD.n3270 VDD.n3269 9.3005
R11272 VDD.n3267 VDD.n3266 9.3005
R11273 VDD.n3275 VDD.n3274 9.3005
R11274 VDD.n3256 VDD.n3255 9.3005
R11275 VDD.n3253 VDD.n3252 9.3005
R11276 VDD.n3261 VDD.n3260 9.3005
R11277 VDD.n3242 VDD.n3241 9.3005
R11278 VDD.n3239 VDD.n3238 9.3005
R11279 VDD.n3247 VDD.n3246 9.3005
R11280 VDD.n3228 VDD.n3227 9.3005
R11281 VDD.n3225 VDD.n3224 9.3005
R11282 VDD.n3233 VDD.n3232 9.3005
R11283 VDD.n3169 VDD.n3168 9.3005
R11284 VDD.n3166 VDD.n3165 9.3005
R11285 VDD.n3174 VDD.n3173 9.3005
R11286 VDD.n3620 VDD.n3619 9.3005
R11287 VDD.n3603 VDD.n3602 9.3005
R11288 VDD.n3626 VDD.n3625 9.3005
R11289 VDD.n3607 VDD.n3606 9.3005
R11290 VDD.n3615 VDD.n3614 9.3005
R11291 VDD.n3617 VDD.n3616 9.3005
R11292 VDD.n3634 VDD.n3633 9.3005
R11293 VDD.n3631 VDD.n3630 9.3005
R11294 VDD.n3639 VDD.n3638 9.3005
R11295 VDD.n3648 VDD.n3647 9.3005
R11296 VDD.n3645 VDD.n3644 9.3005
R11297 VDD.n3653 VDD.n3652 9.3005
R11298 VDD.n3661 VDD.n3660 9.3005
R11299 VDD.n3658 VDD.n3657 9.3005
R11300 VDD.n3666 VDD.n3665 9.3005
R11301 VDD.n3674 VDD.n3673 9.3005
R11302 VDD.n3671 VDD.n3670 9.3005
R11303 VDD.n3679 VDD.n3678 9.3005
R11304 VDD.n3687 VDD.n3686 9.3005
R11305 VDD.n3684 VDD.n3683 9.3005
R11306 VDD.n3692 VDD.n3691 9.3005
R11307 VDD.n3700 VDD.n3699 9.3005
R11308 VDD.n3697 VDD.n3696 9.3005
R11309 VDD.n3705 VDD.n3704 9.3005
R11310 VDD.n3713 VDD.n3712 9.3005
R11311 VDD.n3710 VDD.n3709 9.3005
R11312 VDD.n3718 VDD.n3717 9.3005
R11313 VDD.n3727 VDD.n3726 9.3005
R11314 VDD.n3724 VDD.n3723 9.3005
R11315 VDD.n3732 VDD.n3731 9.3005
R11316 VDD.n3740 VDD.n3739 9.3005
R11317 VDD.n3737 VDD.n3736 9.3005
R11318 VDD.n3745 VDD.n3744 9.3005
R11319 VDD.n3753 VDD.n3752 9.3005
R11320 VDD.n3750 VDD.n3749 9.3005
R11321 VDD.n3758 VDD.n3757 9.3005
R11322 VDD.n3766 VDD.n3765 9.3005
R11323 VDD.n3763 VDD.n3762 9.3005
R11324 VDD.n3771 VDD.n3770 9.3005
R11325 VDD.n3779 VDD.n3778 9.3005
R11326 VDD.n3776 VDD.n3775 9.3005
R11327 VDD.n3784 VDD.n3783 9.3005
R11328 VDD.n3580 VDD.n3579 9.3005
R11329 VDD.n3577 VDD.n3576 9.3005
R11330 VDD.n3585 VDD.n3584 9.3005
R11331 VDD.n3566 VDD.n3565 9.3005
R11332 VDD.n3563 VDD.n3562 9.3005
R11333 VDD.n3571 VDD.n3570 9.3005
R11334 VDD.n3552 VDD.n3551 9.3005
R11335 VDD.n3549 VDD.n3548 9.3005
R11336 VDD.n3557 VDD.n3556 9.3005
R11337 VDD.n3538 VDD.n3537 9.3005
R11338 VDD.n3535 VDD.n3534 9.3005
R11339 VDD.n3543 VDD.n3542 9.3005
R11340 VDD.n3524 VDD.n3523 9.3005
R11341 VDD.n3521 VDD.n3520 9.3005
R11342 VDD.n3529 VDD.n3528 9.3005
R11343 VDD.n3510 VDD.n3509 9.3005
R11344 VDD.n3507 VDD.n3506 9.3005
R11345 VDD.n3515 VDD.n3514 9.3005
R11346 VDD.n3495 VDD.n3494 9.3005
R11347 VDD.n3492 VDD.n3491 9.3005
R11348 VDD.n3500 VDD.n3499 9.3005
R11349 VDD.n3480 VDD.n3479 9.3005
R11350 VDD.n3463 VDD.n3462 9.3005
R11351 VDD.n3486 VDD.n3485 9.3005
R11352 VDD.n3467 VDD.n3466 9.3005
R11353 VDD.n3475 VDD.n3474 9.3005
R11354 VDD.n3477 VDD.n3476 9.3005
R11355 VDD.n15 VDD.n14 9.3005
R11356 VDD.n17 VDD.n16 9.3005
R11357 VDD.n8 VDD.n7 9.3005
R11358 VDD.n23 VDD.n22 9.3005
R11359 VDD.n334 VDD.n333 9.3005
R11360 VDD.n336 VDD.n335 9.3005
R11361 VDD.n327 VDD.n326 9.3005
R11362 VDD.n342 VDD.n341 9.3005
R11363 VDD.n317 VDD.n316 9.3005
R11364 VDD.n311 VDD.n310 9.3005
R11365 VDD.n150 VDD.n149 9.3005
R11366 VDD.n158 VDD.n154 9.3005
R11367 VDD.n63 VDD.n26 9.3005
R11368 VDD.n58 VDD.n27 9.3005
R11369 VDD.n401 VDD.n400 9.3005
R11370 VDD.n403 VDD.n402 9.3005
R11371 VDD.n309 VDD.n308 9.3005
R11372 VDD.n177 VDD.n153 9.3005
R11373 VDD.n161 VDD.n160 9.3005
R11374 VDD.n203 VDD.n191 9.3005
R11375 VDD.n230 VDD.n229 9.3005
R11376 VDD.n223 VDD.n222 9.3005
R11377 VDD.n241 VDD.n240 9.3005
R11378 VDD.n232 VDD.n231 9.3005
R11379 VDD.n238 VDD.n189 9.3005
R11380 VDD.n202 VDD.n201 9.3005
R11381 VDD.n546 VDD.n545 9.3005
R11382 VDD.n530 VDD.n528 9.3005
R11383 VDD.n552 VDD.n551 9.3005
R11384 VDD.n538 VDD.n527 9.3005
R11385 VDD.n537 VDD.n536 9.3005
R11386 VDD.n535 VDD.n534 9.3005
R11387 VDD.n564 VDD.n555 9.3005
R11388 VDD.n562 VDD.n561 9.3005
R11389 VDD.n560 VDD.n559 9.3005
R11390 VDD.n797 VDD.n788 9.3005
R11391 VDD.n795 VDD.n794 9.3005
R11392 VDD.n793 VDD.n792 9.3005
R11393 VDD.n810 VDD.n801 9.3005
R11394 VDD.n808 VDD.n807 9.3005
R11395 VDD.n806 VDD.n805 9.3005
R11396 VDD.n823 VDD.n814 9.3005
R11397 VDD.n821 VDD.n820 9.3005
R11398 VDD.n819 VDD.n818 9.3005
R11399 VDD.n836 VDD.n827 9.3005
R11400 VDD.n834 VDD.n833 9.3005
R11401 VDD.n832 VDD.n831 9.3005
R11402 VDD.n780 VDD.n771 9.3005
R11403 VDD.n778 VDD.n777 9.3005
R11404 VDD.n776 VDD.n775 9.3005
R11405 VDD.n766 VDD.n757 9.3005
R11406 VDD.n764 VDD.n763 9.3005
R11407 VDD.n762 VDD.n761 9.3005
R11408 VDD.n752 VDD.n743 9.3005
R11409 VDD.n750 VDD.n749 9.3005
R11410 VDD.n748 VDD.n747 9.3005
R11411 VDD.n520 VDD.n511 9.3005
R11412 VDD.n518 VDD.n517 9.3005
R11413 VDD.n516 VDD.n515 9.3005
R11414 VDD.n2577 VDD.n2568 9.3005
R11415 VDD.n2575 VDD.n2574 9.3005
R11416 VDD.n2573 VDD.n2572 9.3005
R11417 VDD.n1858 VDD.n1857 9.3005
R11418 VDD.n1854 VDD.n1852 9.3005
R11419 VDD.n1490 VDD.n1489 9.3005
R11420 VDD.n1918 VDD.n1917 9.3005
R11421 VDD.n1919 VDD.n1487 9.3005
R11422 VDD.n1928 VDD.n1927 9.3005
R11423 VDD.n1926 VDD.n1925 9.3005
R11424 VDD.n1922 VDD.n1920 9.3005
R11425 VDD.n863 VDD.n861 9.3005
R11426 VDD.n2083 VDD.n2082 9.3005
R11427 VDD.n2084 VDD.n1393 9.3005
R11428 VDD.n2089 VDD.n2088 9.3005
R11429 VDD.n2087 VDD.n2086 9.3005
R11430 VDD.n1362 VDD.n1361 9.3005
R11431 VDD.n2116 VDD.n2115 9.3005
R11432 VDD.n2118 VDD.n2117 9.3005
R11433 VDD.n2119 VDD.n1196 9.3005
R11434 VDD.n2544 VDD.n2543 9.3005
R11435 VDD.n2502 VDD.n2501 9.3005
R11436 VDD.n1259 VDD.n1258 9.3005
R11437 VDD.n2197 VDD.n2196 9.3005
R11438 VDD.n2194 VDD.n2193 9.3005
R11439 VDD.n2203 VDD.n2202 9.3005
R11440 VDD.n1539 VDD.n1538 9.3005
R11441 VDD.n1850 VDD.n1849 9.3005
R11442 VDD.n1851 VDD.n1536 9.3005
R11443 VDD.n1860 VDD.n1859 9.3005
R11444 VDD.n2549 VDD.n2548 9.3005
R11445 VDD.n1454 VDD.n864 9.3005
R11446 VDD.n1998 VDD.n1997 9.3005
R11447 VDD.n1999 VDD.n1452 9.3005
R11448 VDD.n2008 VDD.n2007 9.3005
R11449 VDD.n2006 VDD.n2005 9.3005
R11450 VDD.n2002 VDD.n2000 9.3005
R11451 VDD.n1396 VDD.n1395 9.3005
R11452 VDD.n1218 VDD.n1197 9.3005
R11453 VDD.n2527 VDD.n2526 9.3005
R11454 VDD.n2525 VDD.n2524 9.3005
R11455 VDD.n1221 VDD.n1220 9.3005
R11456 VDD.n1251 VDD.n1249 9.3005
R11457 VDD.n1256 VDD.n1255 9.3005
R11458 VDD.n1257 VDD.n1247 9.3005
R11459 VDD.n2504 VDD.n2503 9.3005
R11460 VDD.n2369 VDD.n2368 9.3005
R11461 VDD.n2366 VDD.n2177 9.3005
R11462 VDD.n2181 VDD.n2178 9.3005
R11463 VDD.n2361 VDD.n2360 9.3005
R11464 VDD.n2359 VDD.n2358 9.3005
R11465 VDD.n2371 VDD.n2370 9.3005
R11466 VDD.n2373 VDD.n2173 9.3005
R11467 VDD.n2377 VDD.n2376 9.3005
R11468 VDD.n2379 VDD.n2378 9.3005
R11469 VDD.n1729 VDD.n1728 9.3005
R11470 VDD.n1714 VDD.n1713 9.3005
R11471 VDD.n1723 VDD.n1722 9.3005
R11472 VDD.n1721 VDD.n1720 9.3005
R11473 VDD.n1718 VDD.n1717 9.3005
R11474 VDD.n1731 VDD.n1730 9.3005
R11475 VDD.n1733 VDD.n1711 9.3005
R11476 VDD.n1737 VDD.n1736 9.3005
R11477 VDD.n1739 VDD.n1738 9.3005
R11478 VDD.n1957 VDD.n853 9.3005
R11479 VDD.n1968 VDD.n1959 9.3005
R11480 VDD.n1980 VDD.n1979 9.3005
R11481 VDD.n1962 VDD.n1438 9.3005
R11482 VDD.n2022 VDD.n2021 9.3005
R11483 VDD.n1443 VDD.n1442 9.3005
R11484 VDD.n1445 VDD.n1410 9.3005
R11485 VDD.n2063 VDD.n2062 9.3005
R11486 VDD.n2064 VDD.n1404 9.3005
R11487 VDD.n2536 VDD.n2535 9.3005
R11488 VDD.n2161 VDD.n1211 9.3005
R11489 VDD.n2166 VDD.n2165 9.3005
R11490 VDD.n2171 VDD.n1229 9.3005
R11491 VDD.n1482 VDD.n1477 9.3005
R11492 VDD.n1937 VDD.n1936 9.3005
R11493 VDD.n1480 VDD.n852 9.3005
R11494 VDD.n2557 VDD.n2556 9.3005
R11495 VDD.n2068 VDD.n1406 9.3005
R11496 VDD.n2071 VDD.n2070 9.3005
R11497 VDD.n1388 VDD.n1377 9.3005
R11498 VDD.n2099 VDD.n2098 9.3005
R11499 VDD.n1386 VDD.n1385 9.3005
R11500 VDD.n1382 VDD.n1346 9.3005
R11501 VDD.n2126 VDD.n2125 9.3005
R11502 VDD.n1963 VDD.n1351 9.3005
R11503 VDD.n1354 VDD.n1210 9.3005
R11504 VDD.n1939 VDD.n1938 9.3005
R11505 VDD.n1478 VDD.n850 9.3005
R11506 VDD.n2559 VDD.n2558 9.3005
R11507 VDD.n2073 VDD.n2072 9.3005
R11508 VDD.n1407 VDD.n1375 9.3005
R11509 VDD.n2101 VDD.n2100 9.3005
R11510 VDD.n1380 VDD.n1379 9.3005
R11511 VDD.n1384 VDD.n1344 9.3005
R11512 VDD.n2128 VDD.n2127 9.3005
R11513 VDD.n1349 VDD.n1348 9.3005
R11514 VDD.n1964 VDD.n1208 9.3005
R11515 VDD.n2172 VDD.n2158 9.3005
R11516 VDD.n2170 VDD.n2169 9.3005
R11517 VDD.n2160 VDD.n1213 9.3005
R11518 VDD.n2534 VDD.n2533 9.3005
R11519 VDD.n2066 VDD.n2065 9.3005
R11520 VDD.n2014 VDD.n1409 9.3005
R11521 VDD.n1447 VDD.n1446 9.3005
R11522 VDD.n2020 VDD.n2019 9.3005
R11523 VDD.n1975 VDD.n1440 9.3005
R11524 VDD.n1978 VDD.n1977 9.3005
R11525 VDD.n1973 VDD.n1961 9.3005
R11526 VDD.n1970 VDD.n1969 9.3005
R11527 VDD.n605 VDD.n604 9.3005
R11528 VDD.n588 VDD.n587 9.3005
R11529 VDD.n611 VDD.n610 9.3005
R11530 VDD.n592 VDD.n591 9.3005
R11531 VDD.n600 VDD.n599 9.3005
R11532 VDD.n602 VDD.n601 9.3005
R11533 VDD.n619 VDD.n618 9.3005
R11534 VDD.n616 VDD.n615 9.3005
R11535 VDD.n624 VDD.n623 9.3005
R11536 VDD.n693 VDD.n692 9.3005
R11537 VDD.n690 VDD.n689 9.3005
R11538 VDD.n698 VDD.n697 9.3005
R11539 VDD.n706 VDD.n705 9.3005
R11540 VDD.n703 VDD.n702 9.3005
R11541 VDD.n711 VDD.n710 9.3005
R11542 VDD.n719 VDD.n718 9.3005
R11543 VDD.n716 VDD.n715 9.3005
R11544 VDD.n724 VDD.n723 9.3005
R11545 VDD.n732 VDD.n731 9.3005
R11546 VDD.n729 VDD.n728 9.3005
R11547 VDD.n737 VDD.n736 9.3005
R11548 VDD.n676 VDD.n675 9.3005
R11549 VDD.n673 VDD.n672 9.3005
R11550 VDD.n681 VDD.n680 9.3005
R11551 VDD.n662 VDD.n661 9.3005
R11552 VDD.n659 VDD.n658 9.3005
R11553 VDD.n667 VDD.n666 9.3005
R11554 VDD.n648 VDD.n647 9.3005
R11555 VDD.n645 VDD.n644 9.3005
R11556 VDD.n653 VDD.n652 9.3005
R11557 VDD.n634 VDD.n633 9.3005
R11558 VDD.n631 VDD.n630 9.3005
R11559 VDD.n639 VDD.n638 9.3005
R11560 VDD.n575 VDD.n574 9.3005
R11561 VDD.n572 VDD.n571 9.3005
R11562 VDD.n580 VDD.n579 9.3005
R11563 VDD.n1026 VDD.n1025 9.3005
R11564 VDD.n1009 VDD.n1008 9.3005
R11565 VDD.n1032 VDD.n1031 9.3005
R11566 VDD.n1013 VDD.n1012 9.3005
R11567 VDD.n1021 VDD.n1020 9.3005
R11568 VDD.n1023 VDD.n1022 9.3005
R11569 VDD.n1040 VDD.n1039 9.3005
R11570 VDD.n1037 VDD.n1036 9.3005
R11571 VDD.n1045 VDD.n1044 9.3005
R11572 VDD.n1054 VDD.n1053 9.3005
R11573 VDD.n1051 VDD.n1050 9.3005
R11574 VDD.n1059 VDD.n1058 9.3005
R11575 VDD.n1067 VDD.n1066 9.3005
R11576 VDD.n1064 VDD.n1063 9.3005
R11577 VDD.n1072 VDD.n1071 9.3005
R11578 VDD.n1080 VDD.n1079 9.3005
R11579 VDD.n1077 VDD.n1076 9.3005
R11580 VDD.n1085 VDD.n1084 9.3005
R11581 VDD.n1093 VDD.n1092 9.3005
R11582 VDD.n1090 VDD.n1089 9.3005
R11583 VDD.n1098 VDD.n1097 9.3005
R11584 VDD.n1106 VDD.n1105 9.3005
R11585 VDD.n1103 VDD.n1102 9.3005
R11586 VDD.n1111 VDD.n1110 9.3005
R11587 VDD.n1119 VDD.n1118 9.3005
R11588 VDD.n1116 VDD.n1115 9.3005
R11589 VDD.n1124 VDD.n1123 9.3005
R11590 VDD.n1133 VDD.n1132 9.3005
R11591 VDD.n1130 VDD.n1129 9.3005
R11592 VDD.n1138 VDD.n1137 9.3005
R11593 VDD.n1146 VDD.n1145 9.3005
R11594 VDD.n1143 VDD.n1142 9.3005
R11595 VDD.n1151 VDD.n1150 9.3005
R11596 VDD.n1159 VDD.n1158 9.3005
R11597 VDD.n1156 VDD.n1155 9.3005
R11598 VDD.n1164 VDD.n1163 9.3005
R11599 VDD.n1172 VDD.n1171 9.3005
R11600 VDD.n1169 VDD.n1168 9.3005
R11601 VDD.n1177 VDD.n1176 9.3005
R11602 VDD.n1185 VDD.n1184 9.3005
R11603 VDD.n1182 VDD.n1181 9.3005
R11604 VDD.n1190 VDD.n1189 9.3005
R11605 VDD.n986 VDD.n985 9.3005
R11606 VDD.n983 VDD.n982 9.3005
R11607 VDD.n991 VDD.n990 9.3005
R11608 VDD.n972 VDD.n971 9.3005
R11609 VDD.n969 VDD.n968 9.3005
R11610 VDD.n977 VDD.n976 9.3005
R11611 VDD.n958 VDD.n957 9.3005
R11612 VDD.n955 VDD.n954 9.3005
R11613 VDD.n963 VDD.n962 9.3005
R11614 VDD.n944 VDD.n943 9.3005
R11615 VDD.n941 VDD.n940 9.3005
R11616 VDD.n949 VDD.n948 9.3005
R11617 VDD.n930 VDD.n929 9.3005
R11618 VDD.n927 VDD.n926 9.3005
R11619 VDD.n935 VDD.n934 9.3005
R11620 VDD.n916 VDD.n915 9.3005
R11621 VDD.n913 VDD.n912 9.3005
R11622 VDD.n921 VDD.n920 9.3005
R11623 VDD.n901 VDD.n900 9.3005
R11624 VDD.n898 VDD.n897 9.3005
R11625 VDD.n906 VDD.n905 9.3005
R11626 VDD.n886 VDD.n885 9.3005
R11627 VDD.n869 VDD.n868 9.3005
R11628 VDD.n892 VDD.n891 9.3005
R11629 VDD.n873 VDD.n872 9.3005
R11630 VDD.n881 VDD.n880 9.3005
R11631 VDD.n883 VDD.n882 9.3005
R11632 VDD.n5578 VDD.n5577 9.3005
R11633 VDD.n5580 VDD.n5579 9.3005
R11634 VDD.n5571 VDD.n5570 9.3005
R11635 VDD.n5586 VDD.n5585 9.3005
R11636 VDD.n5897 VDD.n5896 9.3005
R11637 VDD.n5899 VDD.n5898 9.3005
R11638 VDD.n5890 VDD.n5889 9.3005
R11639 VDD.n5905 VDD.n5904 9.3005
R11640 VDD.n5880 VDD.n5879 9.3005
R11641 VDD.n5874 VDD.n5873 9.3005
R11642 VDD.n5713 VDD.n5712 9.3005
R11643 VDD.n5721 VDD.n5717 9.3005
R11644 VDD.n5626 VDD.n5589 9.3005
R11645 VDD.n5621 VDD.n5590 9.3005
R11646 VDD.n5964 VDD.n5963 9.3005
R11647 VDD.n5966 VDD.n5965 9.3005
R11648 VDD.n5872 VDD.n5871 9.3005
R11649 VDD.n5740 VDD.n5716 9.3005
R11650 VDD.n5724 VDD.n5723 9.3005
R11651 VDD.n5766 VDD.n5754 9.3005
R11652 VDD.n5793 VDD.n5792 9.3005
R11653 VDD.n5786 VDD.n5785 9.3005
R11654 VDD.n5804 VDD.n5803 9.3005
R11655 VDD.n5795 VDD.n5794 9.3005
R11656 VDD.n5801 VDD.n5752 9.3005
R11657 VDD.n5765 VDD.n5764 9.3005
R11658 VDD.n5450 VDD.n5449 9.3005
R11659 VDD.n5451 VDD.n5447 9.3005
R11660 VDD.n5453 VDD.n5452 9.3005
R11661 VDD.n5454 VDD.n5446 9.3005
R11662 VDD.n5456 VDD.n5455 9.3005
R11663 VDD.n5458 VDD.n5457 9.3005
R11664 VDD.n5459 VDD.n5444 9.3005
R11665 VDD.n5461 VDD.n5460 9.3005
R11666 VDD.n5490 VDD.n5485 9.3005
R11667 VDD.n5495 VDD.n5494 9.3005
R11668 VDD.n5496 VDD.n5484 9.3005
R11669 VDD.n5498 VDD.n5497 9.3005
R11670 VDD.n5500 VDD.n5482 9.3005
R11671 VDD.n5502 VDD.n5501 9.3005
R11672 VDD.n5510 VDD.n5509 9.3005
R11673 VDD.n5508 VDD.n5507 9.3005
R11674 VDD.n5506 VDD.n5503 9.3005
R11675 VDD.n5477 VDD.n5476 9.3005
R11676 VDD.n5516 VDD.n5515 9.3005
R11677 VDD.n5517 VDD.n5475 9.3005
R11678 VDD.n5519 VDD.n5518 9.3005
R11679 VDD.n5521 VDD.n5473 9.3005
R11680 VDD.n5525 VDD.n5524 9.3005
R11681 VDD.n5526 VDD.n5470 9.3005
R11682 VDD.n5534 VDD.n5533 9.3005
R11683 VDD.n5532 VDD.n5531 9.3005
R11684 VDD.n5530 VDD.n5527 9.3005
R11685 VDD.n5469 VDD.n5468 9.3005
R11686 VDD.n5540 VDD.n5539 9.3005
R11687 VDD.n5542 VDD.n5541 9.3005
R11688 VDD.n5543 VDD.n5465 9.3005
R11689 VDD.n5547 VDD.n5546 9.3005
R11690 VDD.n5548 VDD.n5462 9.3005
R11691 VDD.n5557 VDD.n5556 9.3005
R11692 VDD.n5555 VDD.n5554 9.3005
R11693 VDD.n5553 VDD.n5550 9.3005
R11694 VDD.n5549 VDD.n5442 9.3005
R11695 VDD.n5564 VDD.n5563 9.3005
R11696 VDD.n5428 VDD.n5427 9.3005
R11697 VDD.n5430 VDD.n5429 9.3005
R11698 VDD.n5431 VDD.n5426 9.3005
R11699 VDD.n5432 VDD.n5316 9.3005
R11700 VDD.n5436 VDD.n5435 9.3005
R11701 VDD.n5434 VDD.n5433 9.3005
R11702 VDD.n5347 VDD.n5341 9.3005
R11703 VDD.n5358 VDD.n5357 9.3005
R11704 VDD.n5356 VDD.n5355 9.3005
R11705 VDD.n5354 VDD.n5348 9.3005
R11706 VDD.n5352 VDD.n5351 9.3005
R11707 VDD.n5350 VDD.n5339 9.3005
R11708 VDD.n5364 VDD.n5363 9.3005
R11709 VDD.n5365 VDD.n5338 9.3005
R11710 VDD.n5367 VDD.n5366 9.3005
R11711 VDD.n5369 VDD.n5336 9.3005
R11712 VDD.n5373 VDD.n5372 9.3005
R11713 VDD.n5374 VDD.n5333 9.3005
R11714 VDD.n5380 VDD.n5379 9.3005
R11715 VDD.n5378 VDD.n5377 9.3005
R11716 VDD.n5376 VDD.n5375 9.3005
R11717 VDD.n5332 VDD.n5331 9.3005
R11718 VDD.n5386 VDD.n5385 9.3005
R11719 VDD.n5387 VDD.n5330 9.3005
R11720 VDD.n5389 VDD.n5388 9.3005
R11721 VDD.n5390 VDD.n5328 9.3005
R11722 VDD.n5393 VDD.n5392 9.3005
R11723 VDD.n5394 VDD.n5325 9.3005
R11724 VDD.n5402 VDD.n5401 9.3005
R11725 VDD.n5400 VDD.n5399 9.3005
R11726 VDD.n5398 VDD.n5395 9.3005
R11727 VDD.n5324 VDD.n5323 9.3005
R11728 VDD.n5408 VDD.n5407 9.3005
R11729 VDD.n5410 VDD.n5409 9.3005
R11730 VDD.n5411 VDD.n5320 9.3005
R11731 VDD.n5414 VDD.n5413 9.3005
R11732 VDD.n5415 VDD.n5317 9.3005
R11733 VDD.n5421 VDD.n5420 9.3005
R11734 VDD.n5419 VDD.n5418 9.3005
R11735 VDD.n5417 VDD.n5416 9.3005
R11736 VDD.n5438 VDD.n5437 9.3005
R11737 VDD.n6109 VDD.n6108 9.3005
R11738 VDD.n6093 VDD.n6091 9.3005
R11739 VDD.n6115 VDD.n6114 9.3005
R11740 VDD.n6101 VDD.n6090 9.3005
R11741 VDD.n6100 VDD.n6099 9.3005
R11742 VDD.n6098 VDD.n6097 9.3005
R11743 VDD.n6127 VDD.n6118 9.3005
R11744 VDD.n6125 VDD.n6124 9.3005
R11745 VDD.n6123 VDD.n6122 9.3005
R11746 VDD.n6360 VDD.n6351 9.3005
R11747 VDD.n6358 VDD.n6357 9.3005
R11748 VDD.n6356 VDD.n6355 9.3005
R11749 VDD.n6373 VDD.n6364 9.3005
R11750 VDD.n6371 VDD.n6370 9.3005
R11751 VDD.n6369 VDD.n6368 9.3005
R11752 VDD.n6386 VDD.n6377 9.3005
R11753 VDD.n6384 VDD.n6383 9.3005
R11754 VDD.n6382 VDD.n6381 9.3005
R11755 VDD.n6399 VDD.n6390 9.3005
R11756 VDD.n6397 VDD.n6396 9.3005
R11757 VDD.n6395 VDD.n6394 9.3005
R11758 VDD.n6343 VDD.n6334 9.3005
R11759 VDD.n6341 VDD.n6340 9.3005
R11760 VDD.n6339 VDD.n6338 9.3005
R11761 VDD.n6329 VDD.n6320 9.3005
R11762 VDD.n6327 VDD.n6326 9.3005
R11763 VDD.n6325 VDD.n6324 9.3005
R11764 VDD.n6315 VDD.n6306 9.3005
R11765 VDD.n6313 VDD.n6312 9.3005
R11766 VDD.n6311 VDD.n6310 9.3005
R11767 VDD.n6083 VDD.n6074 9.3005
R11768 VDD.n6081 VDD.n6080 9.3005
R11769 VDD.n6079 VDD.n6078 9.3005
R11770 VDD.n8140 VDD.n8131 9.3005
R11771 VDD.n8138 VDD.n8137 9.3005
R11772 VDD.n8136 VDD.n8135 9.3005
R11773 VDD.n7421 VDD.n7420 9.3005
R11774 VDD.n7417 VDD.n7415 9.3005
R11775 VDD.n7053 VDD.n7052 9.3005
R11776 VDD.n7481 VDD.n7480 9.3005
R11777 VDD.n7482 VDD.n7050 9.3005
R11778 VDD.n7491 VDD.n7490 9.3005
R11779 VDD.n7489 VDD.n7488 9.3005
R11780 VDD.n7485 VDD.n7483 9.3005
R11781 VDD.n6426 VDD.n6424 9.3005
R11782 VDD.n7646 VDD.n7645 9.3005
R11783 VDD.n7647 VDD.n6956 9.3005
R11784 VDD.n7652 VDD.n7651 9.3005
R11785 VDD.n7650 VDD.n7649 9.3005
R11786 VDD.n6925 VDD.n6924 9.3005
R11787 VDD.n7679 VDD.n7678 9.3005
R11788 VDD.n7681 VDD.n7680 9.3005
R11789 VDD.n7682 VDD.n6759 9.3005
R11790 VDD.n8107 VDD.n8106 9.3005
R11791 VDD.n8065 VDD.n8064 9.3005
R11792 VDD.n6822 VDD.n6821 9.3005
R11793 VDD.n7760 VDD.n7759 9.3005
R11794 VDD.n7757 VDD.n7756 9.3005
R11795 VDD.n7766 VDD.n7765 9.3005
R11796 VDD.n7102 VDD.n7101 9.3005
R11797 VDD.n7413 VDD.n7412 9.3005
R11798 VDD.n7414 VDD.n7099 9.3005
R11799 VDD.n7423 VDD.n7422 9.3005
R11800 VDD.n8112 VDD.n8111 9.3005
R11801 VDD.n7017 VDD.n6427 9.3005
R11802 VDD.n7561 VDD.n7560 9.3005
R11803 VDD.n7562 VDD.n7015 9.3005
R11804 VDD.n7571 VDD.n7570 9.3005
R11805 VDD.n7569 VDD.n7568 9.3005
R11806 VDD.n7565 VDD.n7563 9.3005
R11807 VDD.n6959 VDD.n6958 9.3005
R11808 VDD.n6781 VDD.n6760 9.3005
R11809 VDD.n8090 VDD.n8089 9.3005
R11810 VDD.n8088 VDD.n8087 9.3005
R11811 VDD.n6784 VDD.n6783 9.3005
R11812 VDD.n6814 VDD.n6812 9.3005
R11813 VDD.n6819 VDD.n6818 9.3005
R11814 VDD.n6820 VDD.n6810 9.3005
R11815 VDD.n8067 VDD.n8066 9.3005
R11816 VDD.n7932 VDD.n7931 9.3005
R11817 VDD.n7929 VDD.n7740 9.3005
R11818 VDD.n7744 VDD.n7741 9.3005
R11819 VDD.n7924 VDD.n7923 9.3005
R11820 VDD.n7922 VDD.n7921 9.3005
R11821 VDD.n7934 VDD.n7933 9.3005
R11822 VDD.n7936 VDD.n7736 9.3005
R11823 VDD.n7940 VDD.n7939 9.3005
R11824 VDD.n7942 VDD.n7941 9.3005
R11825 VDD.n7292 VDD.n7291 9.3005
R11826 VDD.n7277 VDD.n7276 9.3005
R11827 VDD.n7286 VDD.n7285 9.3005
R11828 VDD.n7284 VDD.n7283 9.3005
R11829 VDD.n7281 VDD.n7280 9.3005
R11830 VDD.n7294 VDD.n7293 9.3005
R11831 VDD.n7296 VDD.n7274 9.3005
R11832 VDD.n7300 VDD.n7299 9.3005
R11833 VDD.n7302 VDD.n7301 9.3005
R11834 VDD.n7520 VDD.n6416 9.3005
R11835 VDD.n7531 VDD.n7522 9.3005
R11836 VDD.n7543 VDD.n7542 9.3005
R11837 VDD.n7525 VDD.n7001 9.3005
R11838 VDD.n7585 VDD.n7584 9.3005
R11839 VDD.n7006 VDD.n7005 9.3005
R11840 VDD.n7008 VDD.n6973 9.3005
R11841 VDD.n7626 VDD.n7625 9.3005
R11842 VDD.n7627 VDD.n6967 9.3005
R11843 VDD.n8099 VDD.n8098 9.3005
R11844 VDD.n7724 VDD.n6774 9.3005
R11845 VDD.n7729 VDD.n7728 9.3005
R11846 VDD.n7734 VDD.n6792 9.3005
R11847 VDD.n7045 VDD.n7040 9.3005
R11848 VDD.n7500 VDD.n7499 9.3005
R11849 VDD.n7043 VDD.n6415 9.3005
R11850 VDD.n8120 VDD.n8119 9.3005
R11851 VDD.n7631 VDD.n6969 9.3005
R11852 VDD.n7634 VDD.n7633 9.3005
R11853 VDD.n6951 VDD.n6940 9.3005
R11854 VDD.n7662 VDD.n7661 9.3005
R11855 VDD.n6949 VDD.n6948 9.3005
R11856 VDD.n6945 VDD.n6909 9.3005
R11857 VDD.n7689 VDD.n7688 9.3005
R11858 VDD.n7526 VDD.n6914 9.3005
R11859 VDD.n6917 VDD.n6773 9.3005
R11860 VDD.n7502 VDD.n7501 9.3005
R11861 VDD.n7041 VDD.n6413 9.3005
R11862 VDD.n8122 VDD.n8121 9.3005
R11863 VDD.n7636 VDD.n7635 9.3005
R11864 VDD.n6970 VDD.n6938 9.3005
R11865 VDD.n7664 VDD.n7663 9.3005
R11866 VDD.n6943 VDD.n6942 9.3005
R11867 VDD.n6947 VDD.n6907 9.3005
R11868 VDD.n7691 VDD.n7690 9.3005
R11869 VDD.n6912 VDD.n6911 9.3005
R11870 VDD.n7527 VDD.n6771 9.3005
R11871 VDD.n7735 VDD.n7721 9.3005
R11872 VDD.n7733 VDD.n7732 9.3005
R11873 VDD.n7723 VDD.n6776 9.3005
R11874 VDD.n8097 VDD.n8096 9.3005
R11875 VDD.n7629 VDD.n7628 9.3005
R11876 VDD.n7577 VDD.n6972 9.3005
R11877 VDD.n7010 VDD.n7009 9.3005
R11878 VDD.n7583 VDD.n7582 9.3005
R11879 VDD.n7538 VDD.n7003 9.3005
R11880 VDD.n7541 VDD.n7540 9.3005
R11881 VDD.n7536 VDD.n7524 9.3005
R11882 VDD.n7533 VDD.n7532 9.3005
R11883 VDD.n6168 VDD.n6167 9.3005
R11884 VDD.n6151 VDD.n6150 9.3005
R11885 VDD.n6174 VDD.n6173 9.3005
R11886 VDD.n6155 VDD.n6154 9.3005
R11887 VDD.n6163 VDD.n6162 9.3005
R11888 VDD.n6165 VDD.n6164 9.3005
R11889 VDD.n6182 VDD.n6181 9.3005
R11890 VDD.n6179 VDD.n6178 9.3005
R11891 VDD.n6187 VDD.n6186 9.3005
R11892 VDD.n6256 VDD.n6255 9.3005
R11893 VDD.n6253 VDD.n6252 9.3005
R11894 VDD.n6261 VDD.n6260 9.3005
R11895 VDD.n6269 VDD.n6268 9.3005
R11896 VDD.n6266 VDD.n6265 9.3005
R11897 VDD.n6274 VDD.n6273 9.3005
R11898 VDD.n6282 VDD.n6281 9.3005
R11899 VDD.n6279 VDD.n6278 9.3005
R11900 VDD.n6287 VDD.n6286 9.3005
R11901 VDD.n6295 VDD.n6294 9.3005
R11902 VDD.n6292 VDD.n6291 9.3005
R11903 VDD.n6300 VDD.n6299 9.3005
R11904 VDD.n6239 VDD.n6238 9.3005
R11905 VDD.n6236 VDD.n6235 9.3005
R11906 VDD.n6244 VDD.n6243 9.3005
R11907 VDD.n6225 VDD.n6224 9.3005
R11908 VDD.n6222 VDD.n6221 9.3005
R11909 VDD.n6230 VDD.n6229 9.3005
R11910 VDD.n6211 VDD.n6210 9.3005
R11911 VDD.n6208 VDD.n6207 9.3005
R11912 VDD.n6216 VDD.n6215 9.3005
R11913 VDD.n6197 VDD.n6196 9.3005
R11914 VDD.n6194 VDD.n6193 9.3005
R11915 VDD.n6202 VDD.n6201 9.3005
R11916 VDD.n6138 VDD.n6137 9.3005
R11917 VDD.n6135 VDD.n6134 9.3005
R11918 VDD.n6143 VDD.n6142 9.3005
R11919 VDD.n6589 VDD.n6588 9.3005
R11920 VDD.n6572 VDD.n6571 9.3005
R11921 VDD.n6595 VDD.n6594 9.3005
R11922 VDD.n6576 VDD.n6575 9.3005
R11923 VDD.n6584 VDD.n6583 9.3005
R11924 VDD.n6586 VDD.n6585 9.3005
R11925 VDD.n6603 VDD.n6602 9.3005
R11926 VDD.n6600 VDD.n6599 9.3005
R11927 VDD.n6608 VDD.n6607 9.3005
R11928 VDD.n6617 VDD.n6616 9.3005
R11929 VDD.n6614 VDD.n6613 9.3005
R11930 VDD.n6622 VDD.n6621 9.3005
R11931 VDD.n6630 VDD.n6629 9.3005
R11932 VDD.n6627 VDD.n6626 9.3005
R11933 VDD.n6635 VDD.n6634 9.3005
R11934 VDD.n6643 VDD.n6642 9.3005
R11935 VDD.n6640 VDD.n6639 9.3005
R11936 VDD.n6648 VDD.n6647 9.3005
R11937 VDD.n6656 VDD.n6655 9.3005
R11938 VDD.n6653 VDD.n6652 9.3005
R11939 VDD.n6661 VDD.n6660 9.3005
R11940 VDD.n6669 VDD.n6668 9.3005
R11941 VDD.n6666 VDD.n6665 9.3005
R11942 VDD.n6674 VDD.n6673 9.3005
R11943 VDD.n6682 VDD.n6681 9.3005
R11944 VDD.n6679 VDD.n6678 9.3005
R11945 VDD.n6687 VDD.n6686 9.3005
R11946 VDD.n6696 VDD.n6695 9.3005
R11947 VDD.n6693 VDD.n6692 9.3005
R11948 VDD.n6701 VDD.n6700 9.3005
R11949 VDD.n6709 VDD.n6708 9.3005
R11950 VDD.n6706 VDD.n6705 9.3005
R11951 VDD.n6714 VDD.n6713 9.3005
R11952 VDD.n6722 VDD.n6721 9.3005
R11953 VDD.n6719 VDD.n6718 9.3005
R11954 VDD.n6727 VDD.n6726 9.3005
R11955 VDD.n6735 VDD.n6734 9.3005
R11956 VDD.n6732 VDD.n6731 9.3005
R11957 VDD.n6740 VDD.n6739 9.3005
R11958 VDD.n6748 VDD.n6747 9.3005
R11959 VDD.n6745 VDD.n6744 9.3005
R11960 VDD.n6753 VDD.n6752 9.3005
R11961 VDD.n6549 VDD.n6548 9.3005
R11962 VDD.n6546 VDD.n6545 9.3005
R11963 VDD.n6554 VDD.n6553 9.3005
R11964 VDD.n6535 VDD.n6534 9.3005
R11965 VDD.n6532 VDD.n6531 9.3005
R11966 VDD.n6540 VDD.n6539 9.3005
R11967 VDD.n6521 VDD.n6520 9.3005
R11968 VDD.n6518 VDD.n6517 9.3005
R11969 VDD.n6526 VDD.n6525 9.3005
R11970 VDD.n6507 VDD.n6506 9.3005
R11971 VDD.n6504 VDD.n6503 9.3005
R11972 VDD.n6512 VDD.n6511 9.3005
R11973 VDD.n6493 VDD.n6492 9.3005
R11974 VDD.n6490 VDD.n6489 9.3005
R11975 VDD.n6498 VDD.n6497 9.3005
R11976 VDD.n6479 VDD.n6478 9.3005
R11977 VDD.n6476 VDD.n6475 9.3005
R11978 VDD.n6484 VDD.n6483 9.3005
R11979 VDD.n6464 VDD.n6463 9.3005
R11980 VDD.n6461 VDD.n6460 9.3005
R11981 VDD.n6469 VDD.n6468 9.3005
R11982 VDD.n6449 VDD.n6448 9.3005
R11983 VDD.n6432 VDD.n6431 9.3005
R11984 VDD.n6455 VDD.n6454 9.3005
R11985 VDD.n6436 VDD.n6435 9.3005
R11986 VDD.n6444 VDD.n6443 9.3005
R11987 VDD.n6446 VDD.n6445 9.3005
R11988 VDD.n5236 VDD.n5235 9.3005
R11989 VDD.n5234 VDD.n5232 9.3005
R11990 VDD.n5233 VDD.n5191 9.3005
R11991 VDD.n5242 VDD.n5189 9.3005
R11992 VDD.n5244 VDD.n5243 9.3005
R11993 VDD.n5215 VDD.n5214 9.3005
R11994 VDD.n5224 VDD.n5223 9.3005
R11995 VDD.n5222 VDD.n5199 9.3005
R11996 VDD.n5221 VDD.n5220 9.3005
R11997 VDD.n5218 VDD.n5217 9.3005
R11998 VDD.n5275 VDD.n5274 9.3005
R11999 VDD.n5281 VDD.n5280 9.3005
R12000 VDD.n5279 VDD.n5259 9.3005
R12001 VDD.n5278 VDD.n5277 9.3005
R12002 VDD.n5256 VDD.n5255 9.3005
R12003 VDD.n5288 VDD.n5287 9.3005
R12004 VDD.n5294 VDD.n5293 9.3005
R12005 VDD.n5292 VDD.n5254 9.3005
R12006 VDD.n5291 VDD.n5290 9.3005
R12007 VDD.n5249 VDD.n5248 9.3005
R12008 VDD.n5301 VDD.n5300 9.3005
R12009 VDD.n4586 VDD.t647 9.2005
R12010 VDD.n1992 VDD.t350 9.2005
R12011 VDD.n7555 VDD.t703 9.2005
R12012 VDD.n4672 VDD.t617 9.0005
R12013 VDD.n2078 VDD.t384 9.0005
R12014 VDD.n7641 VDD.t363 9.0005
R12015 VDD.n5511 VDD.n5510 8.92171
R12016 VDD.n4645 VDD.t607 8.8005
R12017 VDD.n2051 VDD.t292 8.8005
R12018 VDD.n7614 VDD.t326 8.8005
R12019 VDD.n2694 VDD.t503 8.72499
R12020 VDD.n3046 VDD.t505 8.72499
R12021 VDD.n100 VDD.t31 8.72499
R12022 VDD.n452 VDD.t29 8.72499
R12023 VDD.n5663 VDD.t200 8.72499
R12024 VDD.n6015 VDD.t210 8.72499
R12025 VDD.n5433 VDD.n5425 8.65932
R12026 VDD.t657 VDD.n4057 8.6005
R12027 VDD.t273 VDD.n1463 8.6005
R12028 VDD.t154 VDD.n7026 8.6005
R12029 VDD.n4733 VDD.t663 8.4005
R12030 VDD.n2139 VDD.t34 8.4005
R12031 VDD.n7702 VDD.t128 8.4005
R12032 VDD.n3128 VDD.n3126 8.28285
R12033 VDD.n3153 VDD.n3151 8.28285
R12034 VDD.n3386 VDD.n3384 8.28285
R12035 VDD.n3399 VDD.n3397 8.28285
R12036 VDD.n3412 VDD.n3410 8.28285
R12037 VDD.n3425 VDD.n3423 8.28285
R12038 VDD.n3369 VDD.n3367 8.28285
R12039 VDD.n3355 VDD.n3353 8.28285
R12040 VDD.n3341 VDD.n3339 8.28285
R12041 VDD.n3109 VDD.n3107 8.28285
R12042 VDD.n5166 VDD.n5164 8.28285
R12043 VDD.n4534 VDD.n4533 8.28285
R12044 VDD.n4617 VDD.n4032 8.28285
R12045 VDD.n4723 VDD.n4722 8.28285
R12046 VDD.n5112 VDD.n3823 8.28285
R12047 VDD.n4443 VDD.n4441 8.28285
R12048 VDD.n4511 VDD.n4510 8.28285
R12049 VDD.n4599 VDD.n4047 8.28285
R12050 VDD.n4680 VDD.n4679 8.28285
R12051 VDD.n3849 VDD.n3847 8.28285
R12052 VDD.n4795 VDD.n4788 8.28285
R12053 VDD.n4330 VDD.n4304 8.28285
R12054 VDD.n4314 VDD.n4313 8.28285
R12055 VDD.n4612 VDD.n4041 8.28285
R12056 VDD.n4692 VDD.n4691 8.28285
R12057 VDD.n4970 VDD.n4753 8.28285
R12058 VDD.n4955 VDD.n4774 8.28285
R12059 VDD.n3204 VDD.n3203 8.28285
R12060 VDD.n3217 VDD.n3216 8.28285
R12061 VDD.n3291 VDD.n3290 8.28285
R12062 VDD.n3304 VDD.n3303 8.28285
R12063 VDD.n3317 VDD.n3316 8.28285
R12064 VDD.n3330 VDD.n3329 8.28285
R12065 VDD.n3274 VDD.n3273 8.28285
R12066 VDD.n3260 VDD.n3259 8.28285
R12067 VDD.n3246 VDD.n3245 8.28285
R12068 VDD.n3232 VDD.n3231 8.28285
R12069 VDD.n3173 VDD.n3172 8.28285
R12070 VDD.n3625 VDD.n3624 8.28285
R12071 VDD.n3638 VDD.n3637 8.28285
R12072 VDD.n3652 VDD.n3651 8.28285
R12073 VDD.n3665 VDD.n3664 8.28285
R12074 VDD.n3678 VDD.n3677 8.28285
R12075 VDD.n3691 VDD.n3690 8.28285
R12076 VDD.n3704 VDD.n3703 8.28285
R12077 VDD.n3717 VDD.n3716 8.28285
R12078 VDD.n3731 VDD.n3730 8.28285
R12079 VDD.n3744 VDD.n3743 8.28285
R12080 VDD.n3757 VDD.n3756 8.28285
R12081 VDD.n3770 VDD.n3769 8.28285
R12082 VDD.n3783 VDD.n3782 8.28285
R12083 VDD.n3584 VDD.n3583 8.28285
R12084 VDD.n3570 VDD.n3569 8.28285
R12085 VDD.n3556 VDD.n3555 8.28285
R12086 VDD.n3542 VDD.n3541 8.28285
R12087 VDD.n3528 VDD.n3527 8.28285
R12088 VDD.n3514 VDD.n3513 8.28285
R12089 VDD.n3499 VDD.n3498 8.28285
R12090 VDD.n3485 VDD.n3484 8.28285
R12091 VDD.n534 VDD.n532 8.28285
R12092 VDD.n559 VDD.n557 8.28285
R12093 VDD.n792 VDD.n790 8.28285
R12094 VDD.n805 VDD.n803 8.28285
R12095 VDD.n818 VDD.n816 8.28285
R12096 VDD.n831 VDD.n829 8.28285
R12097 VDD.n775 VDD.n773 8.28285
R12098 VDD.n761 VDD.n759 8.28285
R12099 VDD.n747 VDD.n745 8.28285
R12100 VDD.n515 VDD.n513 8.28285
R12101 VDD.n2572 VDD.n2570 8.28285
R12102 VDD.n1940 VDD.n1939 8.28285
R12103 VDD.n2023 VDD.n1438 8.28285
R12104 VDD.n2129 VDD.n2128 8.28285
R12105 VDD.n2518 VDD.n1229 8.28285
R12106 VDD.n1849 VDD.n1847 8.28285
R12107 VDD.n1917 VDD.n1916 8.28285
R12108 VDD.n2005 VDD.n1453 8.28285
R12109 VDD.n2086 VDD.n2085 8.28285
R12110 VDD.n1255 VDD.n1253 8.28285
R12111 VDD.n2201 VDD.n2194 8.28285
R12112 VDD.n1736 VDD.n1710 8.28285
R12113 VDD.n1720 VDD.n1719 8.28285
R12114 VDD.n2018 VDD.n1447 8.28285
R12115 VDD.n2098 VDD.n2097 8.28285
R12116 VDD.n2376 VDD.n2159 8.28285
R12117 VDD.n2361 VDD.n2180 8.28285
R12118 VDD.n610 VDD.n609 8.28285
R12119 VDD.n623 VDD.n622 8.28285
R12120 VDD.n697 VDD.n696 8.28285
R12121 VDD.n710 VDD.n709 8.28285
R12122 VDD.n723 VDD.n722 8.28285
R12123 VDD.n736 VDD.n735 8.28285
R12124 VDD.n680 VDD.n679 8.28285
R12125 VDD.n666 VDD.n665 8.28285
R12126 VDD.n652 VDD.n651 8.28285
R12127 VDD.n638 VDD.n637 8.28285
R12128 VDD.n579 VDD.n578 8.28285
R12129 VDD.n1031 VDD.n1030 8.28285
R12130 VDD.n1044 VDD.n1043 8.28285
R12131 VDD.n1058 VDD.n1057 8.28285
R12132 VDD.n1071 VDD.n1070 8.28285
R12133 VDD.n1084 VDD.n1083 8.28285
R12134 VDD.n1097 VDD.n1096 8.28285
R12135 VDD.n1110 VDD.n1109 8.28285
R12136 VDD.n1123 VDD.n1122 8.28285
R12137 VDD.n1137 VDD.n1136 8.28285
R12138 VDD.n1150 VDD.n1149 8.28285
R12139 VDD.n1163 VDD.n1162 8.28285
R12140 VDD.n1176 VDD.n1175 8.28285
R12141 VDD.n1189 VDD.n1188 8.28285
R12142 VDD.n990 VDD.n989 8.28285
R12143 VDD.n976 VDD.n975 8.28285
R12144 VDD.n962 VDD.n961 8.28285
R12145 VDD.n948 VDD.n947 8.28285
R12146 VDD.n934 VDD.n933 8.28285
R12147 VDD.n920 VDD.n919 8.28285
R12148 VDD.n905 VDD.n904 8.28285
R12149 VDD.n891 VDD.n890 8.28285
R12150 VDD.n6097 VDD.n6095 8.28285
R12151 VDD.n6122 VDD.n6120 8.28285
R12152 VDD.n6355 VDD.n6353 8.28285
R12153 VDD.n6368 VDD.n6366 8.28285
R12154 VDD.n6381 VDD.n6379 8.28285
R12155 VDD.n6394 VDD.n6392 8.28285
R12156 VDD.n6338 VDD.n6336 8.28285
R12157 VDD.n6324 VDD.n6322 8.28285
R12158 VDD.n6310 VDD.n6308 8.28285
R12159 VDD.n6078 VDD.n6076 8.28285
R12160 VDD.n8135 VDD.n8133 8.28285
R12161 VDD.n7503 VDD.n7502 8.28285
R12162 VDD.n7586 VDD.n7001 8.28285
R12163 VDD.n7692 VDD.n7691 8.28285
R12164 VDD.n8081 VDD.n6792 8.28285
R12165 VDD.n7412 VDD.n7410 8.28285
R12166 VDD.n7480 VDD.n7479 8.28285
R12167 VDD.n7568 VDD.n7016 8.28285
R12168 VDD.n7649 VDD.n7648 8.28285
R12169 VDD.n6818 VDD.n6816 8.28285
R12170 VDD.n7764 VDD.n7757 8.28285
R12171 VDD.n7299 VDD.n7273 8.28285
R12172 VDD.n7283 VDD.n7282 8.28285
R12173 VDD.n7581 VDD.n7010 8.28285
R12174 VDD.n7661 VDD.n7660 8.28285
R12175 VDD.n7939 VDD.n7722 8.28285
R12176 VDD.n7924 VDD.n7743 8.28285
R12177 VDD.n6173 VDD.n6172 8.28285
R12178 VDD.n6186 VDD.n6185 8.28285
R12179 VDD.n6260 VDD.n6259 8.28285
R12180 VDD.n6273 VDD.n6272 8.28285
R12181 VDD.n6286 VDD.n6285 8.28285
R12182 VDD.n6299 VDD.n6298 8.28285
R12183 VDD.n6243 VDD.n6242 8.28285
R12184 VDD.n6229 VDD.n6228 8.28285
R12185 VDD.n6215 VDD.n6214 8.28285
R12186 VDD.n6201 VDD.n6200 8.28285
R12187 VDD.n6142 VDD.n6141 8.28285
R12188 VDD.n6594 VDD.n6593 8.28285
R12189 VDD.n6607 VDD.n6606 8.28285
R12190 VDD.n6621 VDD.n6620 8.28285
R12191 VDD.n6634 VDD.n6633 8.28285
R12192 VDD.n6647 VDD.n6646 8.28285
R12193 VDD.n6660 VDD.n6659 8.28285
R12194 VDD.n6673 VDD.n6672 8.28285
R12195 VDD.n6686 VDD.n6685 8.28285
R12196 VDD.n6700 VDD.n6699 8.28285
R12197 VDD.n6713 VDD.n6712 8.28285
R12198 VDD.n6726 VDD.n6725 8.28285
R12199 VDD.n6739 VDD.n6738 8.28285
R12200 VDD.n6752 VDD.n6751 8.28285
R12201 VDD.n6553 VDD.n6552 8.28285
R12202 VDD.n6539 VDD.n6538 8.28285
R12203 VDD.n6525 VDD.n6524 8.28285
R12204 VDD.n6511 VDD.n6510 8.28285
R12205 VDD.n6497 VDD.n6496 8.28285
R12206 VDD.n6483 VDD.n6482 8.28285
R12207 VDD.n6468 VDD.n6467 8.28285
R12208 VDD.n6454 VDD.n6453 8.28285
R12209 VDD.n4104 VDD.t637 8.2005
R12210 VDD.n1510 VDD.t242 8.2005
R12211 VDD.n7073 VDD.t85 8.2005
R12212 VDD.n2618 VDD.n2600 8.16726
R12213 VDD.n2937 VDD.n2919 8.16726
R12214 VDD.n24 VDD.n6 8.16726
R12215 VDD.n343 VDD.n325 8.16726
R12216 VDD.n5587 VDD.n5569 8.16726
R12217 VDD.n5906 VDD.n5888 8.16726
R12218 VDD.n4438 VDD.t392 8.0005
R12219 VDD.n5108 VDD.t627 8.0005
R12220 VDD.n5066 VDD.n3889 8.0005
R12221 VDD.n1844 VDD.t83 8.0005
R12222 VDD.n2514 VDD.t250 8.0005
R12223 VDD.n2472 VDD.n1295 8.0005
R12224 VDD.n7407 VDD.t20 8.0005
R12225 VDD.n8077 VDD.t329 8.0005
R12226 VDD.n8035 VDD.n6858 8.0005
R12227 VDD.n5247 VDD.n5187 7.9575
R12228 VDD.n2996 VDD.n2940 7.93978
R12229 VDD.n402 VDD.n346 7.93978
R12230 VDD.n5965 VDD.n5909 7.93978
R12231 VDD.n2941 VDD.n2940 7.93832
R12232 VDD.n347 VDD.n346 7.93832
R12233 VDD.n5910 VDD.n5909 7.93832
R12234 VDD.n5510 VDD.n5481 7.9292
R12235 VDD.n3101 VDD.n2620 7.9122
R12236 VDD.n507 VDD.n26 7.9122
R12237 VDD.n6070 VDD.n5589 7.9122
R12238 VDD.n2619 VDD.n2618 7.9105
R12239 VDD.n2938 VDD.n2937 7.9105
R12240 VDD.n2793 VDD.n2792 7.9105
R12241 VDD.n2913 VDD.n2912 7.9105
R12242 VDD.n3101 VDD.n3100 7.9105
R12243 VDD.n3148 VDD.n3120 7.9105
R12244 VDD.n3161 VDD.n3119 7.9105
R12245 VDD.n3394 VDD.n3381 7.9105
R12246 VDD.n3407 VDD.n3380 7.9105
R12247 VDD.n3420 VDD.n3379 7.9105
R12248 VDD.n3433 VDD.n3378 7.9105
R12249 VDD.n3377 VDD.n3364 7.9105
R12250 VDD.n3363 VDD.n3350 7.9105
R12251 VDD.n3349 VDD.n3336 7.9105
R12252 VDD.n3117 VDD.n3104 7.9105
R12253 VDD.n5174 VDD.n3103 7.9105
R12254 VDD.n3207 VDD.n3179 7.9105
R12255 VDD.n3220 VDD.n3178 7.9105
R12256 VDD.n3294 VDD.n3281 7.9105
R12257 VDD.n3307 VDD.n3280 7.9105
R12258 VDD.n3320 VDD.n3279 7.9105
R12259 VDD.n3333 VDD.n3278 7.9105
R12260 VDD.n3277 VDD.n3264 7.9105
R12261 VDD.n3263 VDD.n3250 7.9105
R12262 VDD.n3249 VDD.n3236 7.9105
R12263 VDD.n3235 VDD.n3222 7.9105
R12264 VDD.n3176 VDD.n3163 7.9105
R12265 VDD.n3176 VDD.n3175 7.9105
R12266 VDD.n3235 VDD.n3234 7.9105
R12267 VDD.n3249 VDD.n3248 7.9105
R12268 VDD.n3263 VDD.n3262 7.9105
R12269 VDD.n3277 VDD.n3276 7.9105
R12270 VDD.n3333 VDD.n3332 7.9105
R12271 VDD.n3320 VDD.n3319 7.9105
R12272 VDD.n3307 VDD.n3306 7.9105
R12273 VDD.n3294 VDD.n3293 7.9105
R12274 VDD.n3220 VDD.n3219 7.9105
R12275 VDD.n3207 VDD.n3206 7.9105
R12276 VDD.n3628 VDD.n3600 7.9105
R12277 VDD.n3641 VDD.n3599 7.9105
R12278 VDD.n3655 VDD.n3598 7.9105
R12279 VDD.n3668 VDD.n3597 7.9105
R12280 VDD.n3681 VDD.n3596 7.9105
R12281 VDD.n3694 VDD.n3595 7.9105
R12282 VDD.n3707 VDD.n3594 7.9105
R12283 VDD.n3720 VDD.n3593 7.9105
R12284 VDD.n3734 VDD.n3592 7.9105
R12285 VDD.n3747 VDD.n3591 7.9105
R12286 VDD.n3760 VDD.n3590 7.9105
R12287 VDD.n3773 VDD.n3589 7.9105
R12288 VDD.n3786 VDD.n3588 7.9105
R12289 VDD.n3587 VDD.n3574 7.9105
R12290 VDD.n3573 VDD.n3560 7.9105
R12291 VDD.n3559 VDD.n3546 7.9105
R12292 VDD.n3545 VDD.n3532 7.9105
R12293 VDD.n3531 VDD.n3518 7.9105
R12294 VDD.n3517 VDD.n3504 7.9105
R12295 VDD.n3502 VDD.n3489 7.9105
R12296 VDD.n3488 VDD.n3460 7.9105
R12297 VDD.n3488 VDD.n3487 7.9105
R12298 VDD.n3502 VDD.n3501 7.9105
R12299 VDD.n3517 VDD.n3516 7.9105
R12300 VDD.n3531 VDD.n3530 7.9105
R12301 VDD.n3545 VDD.n3544 7.9105
R12302 VDD.n3559 VDD.n3558 7.9105
R12303 VDD.n3573 VDD.n3572 7.9105
R12304 VDD.n3587 VDD.n3586 7.9105
R12305 VDD.n3786 VDD.n3785 7.9105
R12306 VDD.n3773 VDD.n3772 7.9105
R12307 VDD.n3760 VDD.n3759 7.9105
R12308 VDD.n3747 VDD.n3746 7.9105
R12309 VDD.n3734 VDD.n3733 7.9105
R12310 VDD.n3720 VDD.n3719 7.9105
R12311 VDD.n3707 VDD.n3706 7.9105
R12312 VDD.n3694 VDD.n3693 7.9105
R12313 VDD.n3681 VDD.n3680 7.9105
R12314 VDD.n3668 VDD.n3667 7.9105
R12315 VDD.n3655 VDD.n3654 7.9105
R12316 VDD.n3641 VDD.n3640 7.9105
R12317 VDD.n3628 VDD.n3627 7.9105
R12318 VDD.n5174 VDD.n5173 7.9105
R12319 VDD.n3117 VDD.n3116 7.9105
R12320 VDD.n3349 VDD.n3348 7.9105
R12321 VDD.n3363 VDD.n3362 7.9105
R12322 VDD.n3377 VDD.n3376 7.9105
R12323 VDD.n3433 VDD.n3432 7.9105
R12324 VDD.n3420 VDD.n3419 7.9105
R12325 VDD.n3407 VDD.n3406 7.9105
R12326 VDD.n3394 VDD.n3393 7.9105
R12327 VDD.n3161 VDD.n3160 7.9105
R12328 VDD.n3148 VDD.n3147 7.9105
R12329 VDD.n25 VDD.n24 7.9105
R12330 VDD.n344 VDD.n343 7.9105
R12331 VDD.n199 VDD.n198 7.9105
R12332 VDD.n319 VDD.n318 7.9105
R12333 VDD.n507 VDD.n506 7.9105
R12334 VDD.n554 VDD.n526 7.9105
R12335 VDD.n567 VDD.n525 7.9105
R12336 VDD.n800 VDD.n787 7.9105
R12337 VDD.n813 VDD.n786 7.9105
R12338 VDD.n826 VDD.n785 7.9105
R12339 VDD.n839 VDD.n784 7.9105
R12340 VDD.n783 VDD.n770 7.9105
R12341 VDD.n769 VDD.n756 7.9105
R12342 VDD.n755 VDD.n742 7.9105
R12343 VDD.n523 VDD.n510 7.9105
R12344 VDD.n2580 VDD.n509 7.9105
R12345 VDD.n613 VDD.n585 7.9105
R12346 VDD.n626 VDD.n584 7.9105
R12347 VDD.n700 VDD.n687 7.9105
R12348 VDD.n713 VDD.n686 7.9105
R12349 VDD.n726 VDD.n685 7.9105
R12350 VDD.n739 VDD.n684 7.9105
R12351 VDD.n683 VDD.n670 7.9105
R12352 VDD.n669 VDD.n656 7.9105
R12353 VDD.n655 VDD.n642 7.9105
R12354 VDD.n641 VDD.n628 7.9105
R12355 VDD.n582 VDD.n569 7.9105
R12356 VDD.n582 VDD.n581 7.9105
R12357 VDD.n641 VDD.n640 7.9105
R12358 VDD.n655 VDD.n654 7.9105
R12359 VDD.n669 VDD.n668 7.9105
R12360 VDD.n683 VDD.n682 7.9105
R12361 VDD.n739 VDD.n738 7.9105
R12362 VDD.n726 VDD.n725 7.9105
R12363 VDD.n713 VDD.n712 7.9105
R12364 VDD.n700 VDD.n699 7.9105
R12365 VDD.n626 VDD.n625 7.9105
R12366 VDD.n613 VDD.n612 7.9105
R12367 VDD.n1034 VDD.n1006 7.9105
R12368 VDD.n1047 VDD.n1005 7.9105
R12369 VDD.n1061 VDD.n1004 7.9105
R12370 VDD.n1074 VDD.n1003 7.9105
R12371 VDD.n1087 VDD.n1002 7.9105
R12372 VDD.n1100 VDD.n1001 7.9105
R12373 VDD.n1113 VDD.n1000 7.9105
R12374 VDD.n1126 VDD.n999 7.9105
R12375 VDD.n1140 VDD.n998 7.9105
R12376 VDD.n1153 VDD.n997 7.9105
R12377 VDD.n1166 VDD.n996 7.9105
R12378 VDD.n1179 VDD.n995 7.9105
R12379 VDD.n1192 VDD.n994 7.9105
R12380 VDD.n993 VDD.n980 7.9105
R12381 VDD.n979 VDD.n966 7.9105
R12382 VDD.n965 VDD.n952 7.9105
R12383 VDD.n951 VDD.n938 7.9105
R12384 VDD.n937 VDD.n924 7.9105
R12385 VDD.n923 VDD.n910 7.9105
R12386 VDD.n908 VDD.n895 7.9105
R12387 VDD.n894 VDD.n866 7.9105
R12388 VDD.n894 VDD.n893 7.9105
R12389 VDD.n908 VDD.n907 7.9105
R12390 VDD.n923 VDD.n922 7.9105
R12391 VDD.n937 VDD.n936 7.9105
R12392 VDD.n951 VDD.n950 7.9105
R12393 VDD.n965 VDD.n964 7.9105
R12394 VDD.n979 VDD.n978 7.9105
R12395 VDD.n993 VDD.n992 7.9105
R12396 VDD.n1192 VDD.n1191 7.9105
R12397 VDD.n1179 VDD.n1178 7.9105
R12398 VDD.n1166 VDD.n1165 7.9105
R12399 VDD.n1153 VDD.n1152 7.9105
R12400 VDD.n1140 VDD.n1139 7.9105
R12401 VDD.n1126 VDD.n1125 7.9105
R12402 VDD.n1113 VDD.n1112 7.9105
R12403 VDD.n1100 VDD.n1099 7.9105
R12404 VDD.n1087 VDD.n1086 7.9105
R12405 VDD.n1074 VDD.n1073 7.9105
R12406 VDD.n1061 VDD.n1060 7.9105
R12407 VDD.n1047 VDD.n1046 7.9105
R12408 VDD.n1034 VDD.n1033 7.9105
R12409 VDD.n2580 VDD.n2579 7.9105
R12410 VDD.n523 VDD.n522 7.9105
R12411 VDD.n755 VDD.n754 7.9105
R12412 VDD.n769 VDD.n768 7.9105
R12413 VDD.n783 VDD.n782 7.9105
R12414 VDD.n839 VDD.n838 7.9105
R12415 VDD.n826 VDD.n825 7.9105
R12416 VDD.n813 VDD.n812 7.9105
R12417 VDD.n800 VDD.n799 7.9105
R12418 VDD.n567 VDD.n566 7.9105
R12419 VDD.n554 VDD.n553 7.9105
R12420 VDD.n5588 VDD.n5587 7.9105
R12421 VDD.n5907 VDD.n5906 7.9105
R12422 VDD.n5762 VDD.n5761 7.9105
R12423 VDD.n5882 VDD.n5881 7.9105
R12424 VDD.n6070 VDD.n6069 7.9105
R12425 VDD.n6117 VDD.n6089 7.9105
R12426 VDD.n6130 VDD.n6088 7.9105
R12427 VDD.n6363 VDD.n6350 7.9105
R12428 VDD.n6376 VDD.n6349 7.9105
R12429 VDD.n6389 VDD.n6348 7.9105
R12430 VDD.n6402 VDD.n6347 7.9105
R12431 VDD.n6346 VDD.n6333 7.9105
R12432 VDD.n6332 VDD.n6319 7.9105
R12433 VDD.n6318 VDD.n6305 7.9105
R12434 VDD.n6086 VDD.n6073 7.9105
R12435 VDD.n8143 VDD.n6072 7.9105
R12436 VDD.n6176 VDD.n6148 7.9105
R12437 VDD.n6189 VDD.n6147 7.9105
R12438 VDD.n6263 VDD.n6250 7.9105
R12439 VDD.n6276 VDD.n6249 7.9105
R12440 VDD.n6289 VDD.n6248 7.9105
R12441 VDD.n6302 VDD.n6247 7.9105
R12442 VDD.n6246 VDD.n6233 7.9105
R12443 VDD.n6232 VDD.n6219 7.9105
R12444 VDD.n6218 VDD.n6205 7.9105
R12445 VDD.n6204 VDD.n6191 7.9105
R12446 VDD.n6145 VDD.n6132 7.9105
R12447 VDD.n6145 VDD.n6144 7.9105
R12448 VDD.n6204 VDD.n6203 7.9105
R12449 VDD.n6218 VDD.n6217 7.9105
R12450 VDD.n6232 VDD.n6231 7.9105
R12451 VDD.n6246 VDD.n6245 7.9105
R12452 VDD.n6302 VDD.n6301 7.9105
R12453 VDD.n6289 VDD.n6288 7.9105
R12454 VDD.n6276 VDD.n6275 7.9105
R12455 VDD.n6263 VDD.n6262 7.9105
R12456 VDD.n6189 VDD.n6188 7.9105
R12457 VDD.n6176 VDD.n6175 7.9105
R12458 VDD.n6597 VDD.n6569 7.9105
R12459 VDD.n6610 VDD.n6568 7.9105
R12460 VDD.n6624 VDD.n6567 7.9105
R12461 VDD.n6637 VDD.n6566 7.9105
R12462 VDD.n6650 VDD.n6565 7.9105
R12463 VDD.n6663 VDD.n6564 7.9105
R12464 VDD.n6676 VDD.n6563 7.9105
R12465 VDD.n6689 VDD.n6562 7.9105
R12466 VDD.n6703 VDD.n6561 7.9105
R12467 VDD.n6716 VDD.n6560 7.9105
R12468 VDD.n6729 VDD.n6559 7.9105
R12469 VDD.n6742 VDD.n6558 7.9105
R12470 VDD.n6755 VDD.n6557 7.9105
R12471 VDD.n6556 VDD.n6543 7.9105
R12472 VDD.n6542 VDD.n6529 7.9105
R12473 VDD.n6528 VDD.n6515 7.9105
R12474 VDD.n6514 VDD.n6501 7.9105
R12475 VDD.n6500 VDD.n6487 7.9105
R12476 VDD.n6486 VDD.n6473 7.9105
R12477 VDD.n6471 VDD.n6458 7.9105
R12478 VDD.n6457 VDD.n6429 7.9105
R12479 VDD.n6457 VDD.n6456 7.9105
R12480 VDD.n6471 VDD.n6470 7.9105
R12481 VDD.n6486 VDD.n6485 7.9105
R12482 VDD.n6500 VDD.n6499 7.9105
R12483 VDD.n6514 VDD.n6513 7.9105
R12484 VDD.n6528 VDD.n6527 7.9105
R12485 VDD.n6542 VDD.n6541 7.9105
R12486 VDD.n6556 VDD.n6555 7.9105
R12487 VDD.n6755 VDD.n6754 7.9105
R12488 VDD.n6742 VDD.n6741 7.9105
R12489 VDD.n6729 VDD.n6728 7.9105
R12490 VDD.n6716 VDD.n6715 7.9105
R12491 VDD.n6703 VDD.n6702 7.9105
R12492 VDD.n6689 VDD.n6688 7.9105
R12493 VDD.n6676 VDD.n6675 7.9105
R12494 VDD.n6663 VDD.n6662 7.9105
R12495 VDD.n6650 VDD.n6649 7.9105
R12496 VDD.n6637 VDD.n6636 7.9105
R12497 VDD.n6624 VDD.n6623 7.9105
R12498 VDD.n6610 VDD.n6609 7.9105
R12499 VDD.n6597 VDD.n6596 7.9105
R12500 VDD.n8143 VDD.n8142 7.9105
R12501 VDD.n6086 VDD.n6085 7.9105
R12502 VDD.n6318 VDD.n6317 7.9105
R12503 VDD.n6332 VDD.n6331 7.9105
R12504 VDD.n6346 VDD.n6345 7.9105
R12505 VDD.n6402 VDD.n6401 7.9105
R12506 VDD.n6389 VDD.n6388 7.9105
R12507 VDD.n6376 VDD.n6375 7.9105
R12508 VDD.n6363 VDD.n6362 7.9105
R12509 VDD.n6130 VDD.n6129 7.9105
R12510 VDD.n6117 VDD.n6116 7.9105
R12511 VDD.n5247 VDD.n5246 7.9105
R12512 VDD.n4439 VDD.t643 7.8005
R12513 VDD.n3913 VDD.t415 7.8005
R12514 VDD.n1845 VDD.t470 7.8005
R12515 VDD.n1319 VDD.t16 7.8005
R12516 VDD.n7408 VDD.t375 7.8005
R12517 VDD.n6882 VDD.t314 7.8005
R12518 VDD.n4423 VDD.n4151 7.6005
R12519 VDD.n4491 VDD.t390 7.6005
R12520 VDD.n4996 VDD.t655 7.6005
R12521 VDD.n1829 VDD.n1557 7.6005
R12522 VDD.n1897 VDD.t87 7.6005
R12523 VDD.n2402 VDD.t271 7.6005
R12524 VDD.n7392 VDD.n7120 7.6005
R12525 VDD.n7460 VDD.t144 7.6005
R12526 VDD.n7965 VDD.t214 7.6005
R12527 VDD.t611 VDD.n4165 7.4005
R12528 VDD.t396 VDD.n3826 7.4005
R12529 VDD.t651 VDD.n4781 7.4005
R12530 VDD.t542 VDD.n1571 7.4005
R12531 VDD.t111 VDD.n1232 7.4005
R12532 VDD.t248 VDD.n2187 7.4005
R12533 VDD.t138 VDD.n7134 7.4005
R12534 VDD.t46 VDD.n6795 7.4005
R12535 VDD.t507 VDD.n7750 7.4005
R12536 VDD.n4577 VDD.t388 7.2005
R12537 VDD.n1983 VDD.t93 7.2005
R12538 VDD.n7546 VDD.t262 7.2005
R12539 VDD.n5302 VDD 7.04882
R12540 VDD.n4254 VDD.t639 7.0005
R12541 VDD.n4280 VDD.t659 7.0005
R12542 VDD.t408 VDD.n3927 7.0005
R12543 VDD.n4926 VDD.t667 7.0005
R12544 VDD.t665 VDD.n4910 7.0005
R12545 VDD.n1660 VDD.t295 7.0005
R12546 VDD.n1686 VDD.t77 7.0005
R12547 VDD.t464 VDD.n1333 7.0005
R12548 VDD.n2332 VDD.t538 7.0005
R12549 VDD.t126 VDD.n2316 7.0005
R12550 VDD.n7223 VDD.t202 7.0005
R12551 VDD.n7249 VDD.t557 7.0005
R12552 VDD.t24 VDD.n6896 7.0005
R12553 VDD.n7895 VDD.t130 7.0005
R12554 VDD.t169 VDD.n7879 7.0005
R12555 VDD.n2912 VDD.n2742 6.83883
R12556 VDD.n2794 VDD.n2793 6.83883
R12557 VDD.n318 VDD.n148 6.83883
R12558 VDD.n200 VDD.n199 6.83883
R12559 VDD.n5881 VDD.n5711 6.83883
R12560 VDD.n5763 VDD.n5762 6.83883
R12561 VDD.n4671 VDD.t433 6.8005
R12562 VDD.n2077 VDD.t266 6.8005
R12563 VDD.n7640 VDD.t18 6.8005
R12564 VDD.n3133 VDD.n3131 6.77697
R12565 VDD.n3157 VDD.n3156 6.77697
R12566 VDD.n3390 VDD.n3389 6.77697
R12567 VDD.n3403 VDD.n3402 6.77697
R12568 VDD.n3416 VDD.n3415 6.77697
R12569 VDD.n3429 VDD.n3428 6.77697
R12570 VDD.n3373 VDD.n3372 6.77697
R12571 VDD.n3359 VDD.n3358 6.77697
R12572 VDD.n3345 VDD.n3344 6.77697
R12573 VDD.n3113 VDD.n3112 6.77697
R12574 VDD.n5170 VDD.n5169 6.77697
R12575 VDD.n4616 VDD.n4033 6.77697
R12576 VDD.n3972 VDD.n3938 6.77697
R12577 VDD.n4349 VDD.n4133 6.77697
R12578 VDD.n4523 VDD.n4081 6.77697
R12579 VDD.n4603 VDD.n4602 6.77697
R12580 VDD.n4708 VDD.n3956 6.77697
R12581 VDD.n3845 VDD.n3844 6.77697
R12582 VDD.n4796 VDD.n4786 6.77697
R12583 VDD.n4334 VDD.n4333 6.77697
R12584 VDD.n4312 VDD.n4077 6.77697
R12585 VDD.n4613 VDD.n4038 6.77697
R12586 VDD.n3980 VDD.n3977 6.77697
R12587 VDD.n4974 VDD.n4973 6.77697
R12588 VDD.n4952 VDD.n4951 6.77697
R12589 VDD.n3200 VDD.n3182 6.77697
R12590 VDD.n3214 VDD.n3210 6.77697
R12591 VDD.n3288 VDD.n3284 6.77697
R12592 VDD.n3301 VDD.n3297 6.77697
R12593 VDD.n3314 VDD.n3310 6.77697
R12594 VDD.n3327 VDD.n3323 6.77697
R12595 VDD.n3271 VDD.n3267 6.77697
R12596 VDD.n3257 VDD.n3253 6.77697
R12597 VDD.n3243 VDD.n3239 6.77697
R12598 VDD.n3229 VDD.n3225 6.77697
R12599 VDD.n3170 VDD.n3166 6.77697
R12600 VDD.n3621 VDD.n3603 6.77697
R12601 VDD.n3635 VDD.n3631 6.77697
R12602 VDD.n3649 VDD.n3645 6.77697
R12603 VDD.n3662 VDD.n3658 6.77697
R12604 VDD.n3675 VDD.n3671 6.77697
R12605 VDD.n3688 VDD.n3684 6.77697
R12606 VDD.n3701 VDD.n3697 6.77697
R12607 VDD.n3714 VDD.n3710 6.77697
R12608 VDD.n3728 VDD.n3724 6.77697
R12609 VDD.n3741 VDD.n3737 6.77697
R12610 VDD.n3754 VDD.n3750 6.77697
R12611 VDD.n3767 VDD.n3763 6.77697
R12612 VDD.n3780 VDD.n3776 6.77697
R12613 VDD.n3581 VDD.n3577 6.77697
R12614 VDD.n3567 VDD.n3563 6.77697
R12615 VDD.n3553 VDD.n3549 6.77697
R12616 VDD.n3539 VDD.n3535 6.77697
R12617 VDD.n3525 VDD.n3521 6.77697
R12618 VDD.n3511 VDD.n3507 6.77697
R12619 VDD.n3496 VDD.n3492 6.77697
R12620 VDD.n3481 VDD.n3463 6.77697
R12621 VDD.n539 VDD.n537 6.77697
R12622 VDD.n563 VDD.n562 6.77697
R12623 VDD.n796 VDD.n795 6.77697
R12624 VDD.n809 VDD.n808 6.77697
R12625 VDD.n822 VDD.n821 6.77697
R12626 VDD.n835 VDD.n834 6.77697
R12627 VDD.n779 VDD.n778 6.77697
R12628 VDD.n765 VDD.n764 6.77697
R12629 VDD.n751 VDD.n750 6.77697
R12630 VDD.n519 VDD.n518 6.77697
R12631 VDD.n2576 VDD.n2575 6.77697
R12632 VDD.n2022 VDD.n1439 6.77697
R12633 VDD.n1378 VDD.n1344 6.77697
R12634 VDD.n1755 VDD.n1539 6.77697
R12635 VDD.n1929 VDD.n1487 6.77697
R12636 VDD.n2009 VDD.n2008 6.77697
R12637 VDD.n2114 VDD.n1362 6.77697
R12638 VDD.n1251 VDD.n1250 6.77697
R12639 VDD.n2202 VDD.n2192 6.77697
R12640 VDD.n1740 VDD.n1739 6.77697
R12641 VDD.n1718 VDD.n1483 6.77697
R12642 VDD.n2019 VDD.n1444 6.77697
R12643 VDD.n1386 VDD.n1383 6.77697
R12644 VDD.n2380 VDD.n2379 6.77697
R12645 VDD.n2358 VDD.n2357 6.77697
R12646 VDD.n606 VDD.n588 6.77697
R12647 VDD.n620 VDD.n616 6.77697
R12648 VDD.n694 VDD.n690 6.77697
R12649 VDD.n707 VDD.n703 6.77697
R12650 VDD.n720 VDD.n716 6.77697
R12651 VDD.n733 VDD.n729 6.77697
R12652 VDD.n677 VDD.n673 6.77697
R12653 VDD.n663 VDD.n659 6.77697
R12654 VDD.n649 VDD.n645 6.77697
R12655 VDD.n635 VDD.n631 6.77697
R12656 VDD.n576 VDD.n572 6.77697
R12657 VDD.n1027 VDD.n1009 6.77697
R12658 VDD.n1041 VDD.n1037 6.77697
R12659 VDD.n1055 VDD.n1051 6.77697
R12660 VDD.n1068 VDD.n1064 6.77697
R12661 VDD.n1081 VDD.n1077 6.77697
R12662 VDD.n1094 VDD.n1090 6.77697
R12663 VDD.n1107 VDD.n1103 6.77697
R12664 VDD.n1120 VDD.n1116 6.77697
R12665 VDD.n1134 VDD.n1130 6.77697
R12666 VDD.n1147 VDD.n1143 6.77697
R12667 VDD.n1160 VDD.n1156 6.77697
R12668 VDD.n1173 VDD.n1169 6.77697
R12669 VDD.n1186 VDD.n1182 6.77697
R12670 VDD.n987 VDD.n983 6.77697
R12671 VDD.n973 VDD.n969 6.77697
R12672 VDD.n959 VDD.n955 6.77697
R12673 VDD.n945 VDD.n941 6.77697
R12674 VDD.n931 VDD.n927 6.77697
R12675 VDD.n917 VDD.n913 6.77697
R12676 VDD.n902 VDD.n898 6.77697
R12677 VDD.n887 VDD.n869 6.77697
R12678 VDD.n6102 VDD.n6100 6.77697
R12679 VDD.n6126 VDD.n6125 6.77697
R12680 VDD.n6359 VDD.n6358 6.77697
R12681 VDD.n6372 VDD.n6371 6.77697
R12682 VDD.n6385 VDD.n6384 6.77697
R12683 VDD.n6398 VDD.n6397 6.77697
R12684 VDD.n6342 VDD.n6341 6.77697
R12685 VDD.n6328 VDD.n6327 6.77697
R12686 VDD.n6314 VDD.n6313 6.77697
R12687 VDD.n6082 VDD.n6081 6.77697
R12688 VDD.n8139 VDD.n8138 6.77697
R12689 VDD.n7585 VDD.n7002 6.77697
R12690 VDD.n6941 VDD.n6907 6.77697
R12691 VDD.n7318 VDD.n7102 6.77697
R12692 VDD.n7492 VDD.n7050 6.77697
R12693 VDD.n7572 VDD.n7571 6.77697
R12694 VDD.n7677 VDD.n6925 6.77697
R12695 VDD.n6814 VDD.n6813 6.77697
R12696 VDD.n7765 VDD.n7755 6.77697
R12697 VDD.n7303 VDD.n7302 6.77697
R12698 VDD.n7281 VDD.n7046 6.77697
R12699 VDD.n7582 VDD.n7007 6.77697
R12700 VDD.n6949 VDD.n6946 6.77697
R12701 VDD.n7943 VDD.n7942 6.77697
R12702 VDD.n7921 VDD.n7920 6.77697
R12703 VDD.n6169 VDD.n6151 6.77697
R12704 VDD.n6183 VDD.n6179 6.77697
R12705 VDD.n6257 VDD.n6253 6.77697
R12706 VDD.n6270 VDD.n6266 6.77697
R12707 VDD.n6283 VDD.n6279 6.77697
R12708 VDD.n6296 VDD.n6292 6.77697
R12709 VDD.n6240 VDD.n6236 6.77697
R12710 VDD.n6226 VDD.n6222 6.77697
R12711 VDD.n6212 VDD.n6208 6.77697
R12712 VDD.n6198 VDD.n6194 6.77697
R12713 VDD.n6139 VDD.n6135 6.77697
R12714 VDD.n6590 VDD.n6572 6.77697
R12715 VDD.n6604 VDD.n6600 6.77697
R12716 VDD.n6618 VDD.n6614 6.77697
R12717 VDD.n6631 VDD.n6627 6.77697
R12718 VDD.n6644 VDD.n6640 6.77697
R12719 VDD.n6657 VDD.n6653 6.77697
R12720 VDD.n6670 VDD.n6666 6.77697
R12721 VDD.n6683 VDD.n6679 6.77697
R12722 VDD.n6697 VDD.n6693 6.77697
R12723 VDD.n6710 VDD.n6706 6.77697
R12724 VDD.n6723 VDD.n6719 6.77697
R12725 VDD.n6736 VDD.n6732 6.77697
R12726 VDD.n6749 VDD.n6745 6.77697
R12727 VDD.n6550 VDD.n6546 6.77697
R12728 VDD.n6536 VDD.n6532 6.77697
R12729 VDD.n6522 VDD.n6518 6.77697
R12730 VDD.n6508 VDD.n6504 6.77697
R12731 VDD.n6494 VDD.n6490 6.77697
R12732 VDD.n6480 VDD.n6476 6.77697
R12733 VDD.n6465 VDD.n6461 6.77697
R12734 VDD.n6450 VDD.n6432 6.77697
R12735 VDD.n5239 VDD.n5238 6.60764
R12736 VDD.t26 VDD.n5239 6.60764
R12737 VDD.n5241 VDD.n5240 6.60764
R12738 VDD.n5240 VDD.t26 6.60764
R12739 VDD.n5219 VDD.n5194 6.60764
R12740 VDD.t380 VDD.n5194 6.60764
R12741 VDD.n5227 VDD.n5195 6.60764
R12742 VDD.t380 VDD.n5195 6.60764
R12743 VDD.n5252 VDD.n5250 6.60764
R12744 VDD.t483 VDD.n5252 6.60764
R12745 VDD.n5289 VDD.n5251 6.60764
R12746 VDD.t483 VDD.n5251 6.60764
R12747 VDD.n5276 VDD.n5258 6.60764
R12748 VDD.t355 VDD.n5258 6.60764
R12749 VDD.n5284 VDD.n5257 6.60764
R12750 VDD.n5284 VDD.t355 6.60764
R12751 VDD.t639 VDD.n4192 6.6005
R12752 VDD.n4184 VDD.t659 6.6005
R12753 VDD.n4017 VDD.t433 6.6005
R12754 VDD.n4820 VDD.t667 6.6005
R12755 VDD.n4911 VDD.t665 6.6005
R12756 VDD.t295 VDD.n1598 6.6005
R12757 VDD.n1590 VDD.t77 6.6005
R12758 VDD.n1423 VDD.t266 6.6005
R12759 VDD.n2226 VDD.t538 6.6005
R12760 VDD.n2317 VDD.t126 6.6005
R12761 VDD.t202 VDD.n7161 6.6005
R12762 VDD.n7153 VDD.t557 6.6005
R12763 VDD.n6986 VDD.t18 6.6005
R12764 VDD.n7789 VDD.t130 6.6005
R12765 VDD.n7880 VDD.t169 6.6005
R12766 VDD.n5421 VDD.n5319 6.5566
R12767 VDD.n5391 VDD.n5325 6.5566
R12768 VDD.n5340 VDD.n5338 6.5566
R12769 VDD.n5205 VDD.t485 6.5015
R12770 VDD.n5205 VDD.t714 6.5015
R12771 VDD.n5265 VDD.t554 6.5015
R12772 VDD.n5265 VDD.t718 6.5015
R12773 VDD.n5563 VDD.n5562 6.46515
R12774 VDD.n5539 VDD.n5467 6.46515
R12775 VDD.n3952 VDD.t408 6.4005
R12776 VDD.n1358 VDD.t464 6.4005
R12777 VDD.n5445 VDD.n5444 6.4005
R12778 VDD.n5558 VDD.n5557 6.4005
R12779 VDD.n5544 VDD.n5543 6.4005
R12780 VDD.n5507 VDD.n5481 6.4005
R12781 VDD.n5412 VDD.n5317 6.4005
R12782 VDD.n5385 VDD.n5384 6.4005
R12783 VDD.n6921 VDD.t24 6.4005
R12784 VDD.n4299 VDD.t611 6.2005
R12785 VDD.n4587 VDD.t388 6.2005
R12786 VDD.n4936 VDD.t651 6.2005
R12787 VDD.n1705 VDD.t542 6.2005
R12788 VDD.n1993 VDD.t93 6.2005
R12789 VDD.n2342 VDD.t248 6.2005
R12790 VDD.n7268 VDD.t138 6.2005
R12791 VDD.n7556 VDD.t262 6.2005
R12792 VDD.n7905 VDD.t507 6.2005
R12793 VDD.n4423 VDD.n4142 6.0005
R12794 VDD.n4978 VDD.t396 6.0005
R12795 VDD.n1829 VDD.n1548 6.0005
R12796 VDD.n2384 VDD.t111 6.0005
R12797 VDD.n7392 VDD.n7111 6.0005
R12798 VDD.n7947 VDD.t46 6.0005
R12799 VDD.n5566 VDD.n5439 5.938
R12800 VDD.n4525 VDD.t390 5.8005
R12801 VDD.t655 VDD.n3880 5.8005
R12802 VDD.n1931 VDD.t87 5.8005
R12803 VDD.t271 VDD.n1286 5.8005
R12804 VDD.n7494 VDD.t144 5.8005
R12805 VDD.t214 VDD.n6849 5.8005
R12806 VDD.n5363 VDD.n5362 5.77611
R12807 VDD.n3099 VDD.n2622 5.7605
R12808 VDD.n2993 VDD.n2942 5.7605
R12809 VDD.n505 VDD.n28 5.7605
R12810 VDD.n399 VDD.n348 5.7605
R12811 VDD.n6068 VDD.n5591 5.7605
R12812 VDD.n5962 VDD.n5911 5.7605
R12813 VDD.n2917 VDD.t544 5.7135
R12814 VDD.n2917 VDD.t64 5.7135
R12815 VDD.n2915 VDD.t549 5.7135
R12816 VDD.n2915 VDD.t715 5.7135
R12817 VDD.n2740 VDD.t506 5.7135
R12818 VDD.n2740 VDD.t69 5.7135
R12819 VDD.n2788 VDD.t68 5.7135
R12820 VDD.n2788 VDD.t504 5.7135
R12821 VDD.n3150 VDD.t425 5.7135
R12822 VDD.n3150 VDD.t416 5.7135
R12823 VDD.n3383 VDD.t444 5.7135
R12824 VDD.n3383 VDD.t438 5.7135
R12825 VDD.n3396 VDD.t395 5.7135
R12826 VDD.n3396 VDD.t428 5.7135
R12827 VDD.n3409 VDD.t411 5.7135
R12828 VDD.n3409 VDD.t409 5.7135
R12829 VDD.n3422 VDD.t434 5.7135
R12830 VDD.n3422 VDD.t420 5.7135
R12831 VDD.n3366 VDD.t445 5.7135
R12832 VDD.n3366 VDD.t432 5.7135
R12833 VDD.n3352 VDD.t406 5.7135
R12834 VDD.n3352 VDD.t389 5.7135
R12835 VDD.n3338 VDD.t440 5.7135
R12836 VDD.n3338 VDD.t414 5.7135
R12837 VDD.n3106 VDD.t430 5.7135
R12838 VDD.n3106 VDD.t422 5.7135
R12839 VDD.n5163 VDD.t448 5.7135
R12840 VDD.n5163 VDD.t442 5.7135
R12841 VDD.n3215 VDD.t439 5.7135
R12842 VDD.n3215 VDD.t426 5.7135
R12843 VDD.n3289 VDD.t397 5.7135
R12844 VDD.n3289 VDD.t450 5.7135
R12845 VDD.n3302 VDD.t407 5.7135
R12846 VDD.n3302 VDD.t441 5.7135
R12847 VDD.n3315 VDD.t418 5.7135
R12848 VDD.n3315 VDD.t417 5.7135
R12849 VDD.n3328 VDD.t447 5.7135
R12850 VDD.n3328 VDD.t435 5.7135
R12851 VDD.n3272 VDD.t399 5.7135
R12852 VDD.n3272 VDD.t446 5.7135
R12853 VDD.n3258 VDD.t412 5.7135
R12854 VDD.n3258 VDD.t404 5.7135
R12855 VDD.n3244 VDD.t391 5.7135
R12856 VDD.n3244 VDD.t423 5.7135
R12857 VDD.n3230 VDD.t443 5.7135
R12858 VDD.n3230 VDD.t436 5.7135
R12859 VDD.n3171 VDD.t401 5.7135
R12860 VDD.n3171 VDD.t393 5.7135
R12861 VDD.n3636 VDD.t642 5.7135
R12862 VDD.n3636 VDD.t666 5.7135
R12863 VDD.n3650 VDD.t668 5.7135
R12864 VDD.n3650 VDD.t662 5.7135
R12865 VDD.n3663 VDD.t634 5.7135
R12866 VDD.n3663 VDD.t596 5.7135
R12867 VDD.n3676 VDD.t614 5.7135
R12868 VDD.n3676 VDD.t652 5.7135
R12869 VDD.n3689 VDD.t656 5.7135
R12870 VDD.n3689 VDD.t636 5.7135
R12871 VDD.n3702 VDD.t616 5.7135
R12872 VDD.n3702 VDD.t600 5.7135
R12873 VDD.n3715 VDD.t602 5.7135
R12874 VDD.n3715 VDD.t628 5.7135
R12875 VDD.n3729 VDD.t664 5.7135
R12876 VDD.n3729 VDD.t620 5.7135
R12877 VDD.n3742 VDD.t598 5.7135
R12878 VDD.n3742 VDD.t592 5.7135
R12879 VDD.n3755 VDD.t618 5.7135
R12880 VDD.n3755 VDD.t608 5.7135
R12881 VDD.n3768 VDD.t648 5.7135
R12882 VDD.n3768 VDD.t630 5.7135
R12883 VDD.n3781 VDD.t590 5.7135
R12884 VDD.n3781 VDD.t658 5.7135
R12885 VDD.n3582 VDD.t638 5.7135
R12886 VDD.n3582 VDD.t594 5.7135
R12887 VDD.n3568 VDD.t626 5.7135
R12888 VDD.n3568 VDD.t604 5.7135
R12889 VDD.n3554 VDD.t654 5.7135
R12890 VDD.n3554 VDD.t644 5.7135
R12891 VDD.n3540 VDD.t612 5.7135
R12892 VDD.n3540 VDD.t606 5.7135
R12893 VDD.n3526 VDD.t650 5.7135
R12894 VDD.n3526 VDD.t632 5.7135
R12895 VDD.n3512 VDD.t610 5.7135
R12896 VDD.n3512 VDD.t660 5.7135
R12897 VDD.n3497 VDD.t640 5.7135
R12898 VDD.n3497 VDD.t622 5.7135
R12899 VDD.n323 VDD.t30 5.7135
R12900 VDD.n323 VDD.t344 5.7135
R12901 VDD.n321 VDD.t106 5.7135
R12902 VDD.n321 VDD.t32 5.7135
R12903 VDD.n146 VDD.t705 5.7135
R12904 VDD.n146 VDD.t706 5.7135
R12905 VDD.n194 VDD.t253 5.7135
R12906 VDD.n194 VDD.t254 5.7135
R12907 VDD.n556 VDD.t378 5.7135
R12908 VDD.n556 VDD.t17 5.7135
R12909 VDD.n789 VDD.t112 5.7135
R12910 VDD.n789 VDD.t519 5.7135
R12911 VDD.n802 VDD.t90 5.7135
R12912 VDD.n802 VDD.t466 5.7135
R12913 VDD.n815 VDD.t332 5.7135
R12914 VDD.n815 VDD.t465 5.7135
R12915 VDD.n828 VDD.t267 5.7135
R12916 VDD.n828 VDD.t259 5.7135
R12917 VDD.n772 VDD.t178 5.7135
R12918 VDD.n772 VDD.t227 5.7135
R12919 VDD.n758 VDD.t92 5.7135
R12920 VDD.n758 VDD.t94 5.7135
R12921 VDD.n744 VDD.t88 5.7135
R12922 VDD.n744 VDD.t335 5.7135
R12923 VDD.n512 VDD.t160 5.7135
R12924 VDD.n512 VDD.t96 5.7135
R12925 VDD.n2569 VDD.t333 5.7135
R12926 VDD.n2569 VDD.t377 5.7135
R12927 VDD.n621 VDD.t147 5.7135
R12928 VDD.n621 VDD.t110 5.7135
R12929 VDD.n695 VDD.t309 5.7135
R12930 VDD.n695 VDD.t361 5.7135
R12931 VDD.n708 VDD.t197 5.7135
R12932 VDD.n708 VDD.t196 5.7135
R12933 VDD.n721 VDD.t53 5.7135
R12934 VDD.n721 VDD.t512 5.7135
R12935 VDD.n734 VDD.t285 5.7135
R12936 VDD.n734 VDD.t149 5.7135
R12937 VDD.n678 VDD.t82 5.7135
R12938 VDD.n678 VDD.t194 5.7135
R12939 VDD.n664 VDD.t286 5.7135
R12940 VDD.n664 VDD.t109 5.7135
R12941 VDD.n650 VDD.t513 5.7135
R12942 VDD.n650 VDD.t359 5.7135
R12943 VDD.n636 VDD.t100 5.7135
R12944 VDD.n636 VDD.t101 5.7135
R12945 VDD.n577 VDD.t51 5.7135
R12946 VDD.n577 VDD.t84 5.7135
R12947 VDD.n1042 VDD.t37 5.7135
R12948 VDD.n1042 VDD.t127 5.7135
R12949 VDD.n1056 VDD.t539 5.7135
R12950 VDD.n1056 VDD.t222 5.7135
R12951 VDD.n1069 VDD.t502 5.7135
R12952 VDD.n1069 VDD.t358 5.7135
R12953 VDD.n1082 VDD.t337 5.7135
R12954 VDD.n1082 VDD.t249 5.7135
R12955 VDD.n1095 VDD.t272 5.7135
R12956 VDD.n1095 VDD.t190 5.7135
R12957 VDD.n1108 VDD.t455 5.7135
R12958 VDD.n1108 VDD.t347 5.7135
R12959 VDD.n1121 VDD.t247 5.7135
R12960 VDD.n1121 VDD.t251 5.7135
R12961 VDD.n1135 VDD.t35 5.7135
R12962 VDD.n1135 VDD.t325 5.7135
R12963 VDD.n1148 VDD.t13 5.7135
R12964 VDD.n1148 VDD.t241 5.7135
R12965 VDD.n1161 VDD.t385 5.7135
R12966 VDD.n1161 VDD.t293 5.7135
R12967 VDD.n1174 VDD.t351 5.7135
R12968 VDD.n1174 VDD.t11 5.7135
R12969 VDD.n1187 VDD.t702 5.7135
R12970 VDD.n1187 VDD.t274 5.7135
R12971 VDD.n988 VDD.t243 5.7135
R12972 VDD.n988 VDD.t535 5.7135
R12973 VDD.n974 VDD.t469 5.7135
R12974 VDD.n974 VDD.t499 5.7135
R12975 VDD.n960 VDD.t453 5.7135
R12976 VDD.n960 VDD.t471 5.7135
R12977 VDD.n946 VDD.t543 5.7135
R12978 VDD.n946 VDD.t349 5.7135
R12979 VDD.n932 VDD.t5 5.7135
R12980 VDD.n932 VDD.t98 5.7135
R12981 VDD.n918 VDD.t175 5.7135
R12982 VDD.n918 VDD.t78 5.7135
R12983 VDD.n903 VDD.t296 5.7135
R12984 VDD.n903 VDD.t7 5.7135
R12985 VDD.n5886 VDD.t278 5.7135
R12986 VDD.n5886 VDD.t362 5.7135
R12987 VDD.n5884 VDD.t356 5.7135
R12988 VDD.n5884 VDD.t473 5.7135
R12989 VDD.n5709 VDD.t211 5.7135
R12990 VDD.n5709 VDD.t213 5.7135
R12991 VDD.n5757 VDD.t164 5.7135
R12992 VDD.n5757 VDD.t201 5.7135
R12993 VDD.n6119 VDD.t260 5.7135
R12994 VDD.n6119 VDD.t315 5.7135
R12995 VDD.n6352 VDD.t523 5.7135
R12996 VDD.n6352 VDD.t62 5.7135
R12997 VDD.n6365 VDD.t536 5.7135
R12998 VDD.n6365 VDD.t218 5.7135
R12999 VDD.n6378 VDD.t580 5.7135
R13000 VDD.n6378 VDD.t25 5.7135
R13001 VDD.n6391 VDD.t19 5.7135
R13002 VDD.n6391 VDD.t142 5.7135
R13003 VDD.n6335 VDD.t537 5.7135
R13004 VDD.n6335 VDD.t282 5.7135
R13005 VDD.n6321 VDD.t1 5.7135
R13006 VDD.n6321 VDD.t678 5.7135
R13007 VDD.n6307 VDD.t145 5.7135
R13008 VDD.n6307 VDD.t3 5.7135
R13009 VDD.n6075 VDD.t279 5.7135
R13010 VDD.n6075 VDD.t489 5.7135
R13011 VDD.n8132 VDD.t298 5.7135
R13012 VDD.n8132 VDD.t21 5.7135
R13013 VDD.n6184 VDD.t23 5.7135
R13014 VDD.n6184 VDD.t479 5.7135
R13015 VDD.n6258 VDD.t47 5.7135
R13016 VDD.n6258 VDD.t313 5.7135
R13017 VDD.n6271 VDD.t166 5.7135
R13018 VDD.n6271 VDD.t217 5.7135
R13019 VDD.n6284 VDD.t679 5.7135
R13020 VDD.n6284 VDD.t511 5.7135
R13021 VDD.n6297 VDD.t275 5.7135
R13022 VDD.n6297 VDD.t677 5.7135
R13023 VDD.n6241 VDD.t231 5.7135
R13024 VDD.n6241 VDD.t49 5.7135
R13025 VDD.n6227 VDD.t45 5.7135
R13026 VDD.n6227 VDD.t263 5.7135
R13027 VDD.n6213 VDD.t340 5.7135
R13028 VDD.n6213 VDD.t143 5.7135
R13029 VDD.n6199 VDD.t39 5.7135
R13030 VDD.n6199 VDD.t44 5.7135
R13031 VDD.n6140 VDD.t331 5.7135
R13032 VDD.n6140 VDD.t261 5.7135
R13033 VDD.n6605 VDD.t284 5.7135
R13034 VDD.n6605 VDD.t170 5.7135
R13035 VDD.n6619 VDD.t131 5.7135
R13036 VDD.n6619 VDD.t510 5.7135
R13037 VDD.n6632 VDD.t269 5.7135
R13038 VDD.n6632 VDD.t323 5.7135
R13039 VDD.n6645 VDD.t319 5.7135
R13040 VDD.n6645 VDD.t508 5.7135
R13041 VDD.n6658 VDD.t215 5.7135
R13042 VDD.n6658 VDD.t342 5.7135
R13043 VDD.n6671 VDD.t182 5.7135
R13044 VDD.n6671 VDD.t41 5.7135
R13045 VDD.n6684 VDD.t560 5.7135
R13046 VDD.n6684 VDD.t330 5.7135
R13047 VDD.n6698 VDD.t129 5.7135
R13048 VDD.n6698 VDD.t371 5.7135
R13049 VDD.n6711 VDD.t184 5.7135
R13050 VDD.n6711 VDD.t226 5.7135
R13051 VDD.n6724 VDD.t364 5.7135
R13052 VDD.n6724 VDD.t327 5.7135
R13053 VDD.n6737 VDD.t704 5.7135
R13054 VDD.n6737 VDD.t317 5.7135
R13055 VDD.n6750 VDD.t177 5.7135
R13056 VDD.n6750 VDD.t155 5.7135
R13057 VDD.n6551 VDD.t86 5.7135
R13058 VDD.n6551 VDD.t28 5.7135
R13059 VDD.n6537 VDD.t168 5.7135
R13060 VDD.n6537 VDD.t562 5.7135
R13061 VDD.n6523 VDD.t374 5.7135
R13062 VDD.n6523 VDD.t376 5.7135
R13063 VDD.n6509 VDD.t139 5.7135
R13064 VDD.n6509 VDD.t208 5.7135
R13065 VDD.n6495 VDD.t265 5.7135
R13066 VDD.n6495 VDD.t157 5.7135
R13067 VDD.n6481 VDD.t9 5.7135
R13068 VDD.n6481 VDD.t558 5.7135
R13069 VDD.n6466 VDD.t203 5.7135
R13070 VDD.n6466 VDD.t159 5.7135
R13071 VDD.n4465 VDD.t643 5.6005
R13072 VDD.n5085 VDD.t415 5.6005
R13073 VDD.n5066 VDD.n3908 5.6005
R13074 VDD.n1871 VDD.t470 5.6005
R13075 VDD.n2491 VDD.t16 5.6005
R13076 VDD.n2472 VDD.n1314 5.6005
R13077 VDD.n7434 VDD.t375 5.6005
R13078 VDD.n8054 VDD.t314 5.6005
R13079 VDD.n8035 VDD.n6877 5.6005
R13080 VDD.t392 VDD.n4114 5.4005
R13081 VDD.n3835 VDD.t627 5.4005
R13082 VDD.t83 VDD.n1520 5.4005
R13083 VDD.n1241 VDD.t250 5.4005
R13084 VDD.t20 VDD.n7083 5.4005
R13085 VDD.n6804 VDD.t329 5.4005
R13086 VDD.n2616 VDD.n2615 5.27109
R13087 VDD.n2935 VDD.n2934 5.27109
R13088 VDD.n3132 VDD.n3123 5.27109
R13089 VDD.n4036 VDD.n4035 5.27109
R13090 VDD.n3973 VDD.n3970 5.27109
R13091 VDD.n4351 VDD.n4350 5.27109
R13092 VDD.n4522 VDD.n4082 5.27109
R13093 VDD.n4590 VDD.n4046 5.27109
R13094 VDD.n4709 VDD.n3954 5.27109
R13095 VDD.n5117 VDD.n3815 5.27109
R13096 VDD.n4799 VDD.n4798 5.27109
R13097 VDD.n4337 VDD.n4303 5.27109
R13098 VDD.n4076 VDD.n4073 5.27109
R13099 VDD.n4570 VDD.n4569 5.27109
R13100 VDD.n3976 VDD.n3944 5.27109
R13101 VDD.n4762 VDD.n4752 5.27109
R13102 VDD.n4948 VDD.n4776 5.27109
R13103 VDD.n3199 VDD.n3197 5.27109
R13104 VDD.n3620 VDD.n3618 5.27109
R13105 VDD.n3480 VDD.n3478 5.27109
R13106 VDD.n22 VDD.n21 5.27109
R13107 VDD.n341 VDD.n340 5.27109
R13108 VDD.n538 VDD.n529 5.27109
R13109 VDD.n1442 VDD.n1441 5.27109
R13110 VDD.n1379 VDD.n1376 5.27109
R13111 VDD.n1757 VDD.n1756 5.27109
R13112 VDD.n1928 VDD.n1488 5.27109
R13113 VDD.n1996 VDD.n1452 5.27109
R13114 VDD.n2115 VDD.n1360 5.27109
R13115 VDD.n2523 VDD.n1221 5.27109
R13116 VDD.n2205 VDD.n2204 5.27109
R13117 VDD.n1743 VDD.n1709 5.27109
R13118 VDD.n1482 VDD.n1479 5.27109
R13119 VDD.n1976 VDD.n1975 5.27109
R13120 VDD.n1382 VDD.n1350 5.27109
R13121 VDD.n2168 VDD.n2158 5.27109
R13122 VDD.n2354 VDD.n2182 5.27109
R13123 VDD.n605 VDD.n603 5.27109
R13124 VDD.n1026 VDD.n1024 5.27109
R13125 VDD.n886 VDD.n884 5.27109
R13126 VDD.n5585 VDD.n5584 5.27109
R13127 VDD.n5904 VDD.n5903 5.27109
R13128 VDD.n6101 VDD.n6092 5.27109
R13129 VDD.n7005 VDD.n7004 5.27109
R13130 VDD.n6942 VDD.n6939 5.27109
R13131 VDD.n7320 VDD.n7319 5.27109
R13132 VDD.n7491 VDD.n7051 5.27109
R13133 VDD.n7559 VDD.n7015 5.27109
R13134 VDD.n7678 VDD.n6923 5.27109
R13135 VDD.n8086 VDD.n6784 5.27109
R13136 VDD.n7768 VDD.n7767 5.27109
R13137 VDD.n7306 VDD.n7272 5.27109
R13138 VDD.n7045 VDD.n7042 5.27109
R13139 VDD.n7539 VDD.n7538 5.27109
R13140 VDD.n6945 VDD.n6913 5.27109
R13141 VDD.n7731 VDD.n7721 5.27109
R13142 VDD.n7917 VDD.n7745 5.27109
R13143 VDD.n6168 VDD.n6166 5.27109
R13144 VDD.n6589 VDD.n6587 5.27109
R13145 VDD.n6449 VDD.n6447 5.27109
R13146 VDD.n4506 VDD.t637 5.2005
R13147 VDD.n1912 VDD.t242 5.2005
R13148 VDD.n7475 VDD.t85 5.2005
R13149 VDD.n2754 VDD.n2753 5.12506
R13150 VDD.n2834 VDD.n2833 5.12506
R13151 VDD.n160 VDD.n159 5.12506
R13152 VDD.n240 VDD.n239 5.12506
R13153 VDD.n5723 VDD.n5722 5.12506
R13154 VDD.n5803 VDD.n5802 5.12506
R13155 VDD.n5134 VDD.t663 5.0005
R13156 VDD.n2540 VDD.t34 5.0005
R13157 VDD.n8103 VDD.t128 5.0005
R13158 VDD.n4549 VDD.t657 4.8005
R13159 VDD.n1955 VDD.t273 4.8005
R13160 VDD.n7518 VDD.t154 4.8005
R13161 VDD.n4686 VDD.t607 4.6005
R13162 VDD.n2092 VDD.t292 4.6005
R13163 VDD.n7655 VDD.t326 4.6005
R13164 VDD.n2609 VDD.n2605 4.51911
R13165 VDD.n2928 VDD.n2924 4.51911
R13166 VDD.n3139 VDD.n3138 4.51911
R13167 VDD.n3188 VDD.n3185 4.51911
R13168 VDD.n3609 VDD.n3606 4.51911
R13169 VDD.n3469 VDD.n3466 4.51911
R13170 VDD.n15 VDD.n11 4.51911
R13171 VDD.n334 VDD.n330 4.51911
R13172 VDD.n545 VDD.n544 4.51911
R13173 VDD.n594 VDD.n591 4.51911
R13174 VDD.n1015 VDD.n1012 4.51911
R13175 VDD.n875 VDD.n872 4.51911
R13176 VDD.n5578 VDD.n5574 4.51911
R13177 VDD.n5897 VDD.n5893 4.51911
R13178 VDD.n6108 VDD.n6107 4.51911
R13179 VDD.n6157 VDD.n6154 4.51911
R13180 VDD.n6578 VDD.n6575 4.51911
R13181 VDD.n6438 VDD.n6435 4.51911
R13182 VDD.n4584 VDD.n4580 4.51815
R13183 VDD.n4580 VDD.n4054 4.51815
R13184 VDD.n1990 VDD.n1986 4.51815
R13185 VDD.n1986 VDD.n1460 4.51815
R13186 VDD.n7553 VDD.n7549 4.51815
R13187 VDD.n7549 VDD.n7023 4.51815
R13188 VDD.n5566 VDD.n5565 4.5005
R13189 VDD.n2656 VDD.n2652 4.4805
R13190 VDD.n2994 VDD.n2739 4.4805
R13191 VDD.n62 VDD.n58 4.4805
R13192 VDD.n400 VDD.n145 4.4805
R13193 VDD.n5625 VDD.n5621 4.4805
R13194 VDD.n5963 VDD.n5708 4.4805
R13195 VDD.n4639 VDD.t617 4.4005
R13196 VDD.n2045 VDD.t384 4.4005
R13197 VDD.n7608 VDD.t363 4.4005
R13198 VDD.n2682 VDD.t67 4.20118
R13199 VDD.n3034 VDD.t63 4.20118
R13200 VDD.n88 VDD.t105 4.20118
R13201 VDD.n440 VDD.t343 4.20118
R13202 VDD.n5651 VDD.t163 4.20118
R13203 VDD.n6003 VDD.t212 4.20118
R13204 VDD.t647 VDD.n4027 4.2005
R13205 VDD.t350 VDD.n1433 4.2005
R13206 VDD.t703 VDD.n6996 4.2005
R13207 VDD.n5359 VDD.n5341 4.14168
R13208 VDD.n4725 VDD.t591 4.0005
R13209 VDD.n2131 VDD.t240 4.0005
R13210 VDD.n7694 VDD.t225 4.0005
R13211 VDD.n5302 VDD.n5247 3.81358
R13212 VDD.t593 VDD.n4066 3.8005
R13213 VDD.t534 VDD.n1472 3.8005
R13214 VDD.t27 VDD.n7035 3.8005
R13215 VDD.n2791 VDD.n2790 3.7905
R13216 VDD.n2789 VDD.n2741 3.7905
R13217 VDD.n197 VDD.n196 3.7905
R13218 VDD.n195 VDD.n147 3.7905
R13219 VDD.n5760 VDD.n5759 3.7905
R13220 VDD.n5758 VDD.n5710 3.7905
R13221 VDD.n2612 VDD.n2602 3.76521
R13222 VDD.n2931 VDD.n2921 3.76521
R13223 VDD.n2910 VDD.n2909 3.76521
R13224 VDD.n2795 VDD.n2787 3.76521
R13225 VDD.n3145 VDD.n3144 3.76521
R13226 VDD.n4654 VDD.n4004 3.76521
R13227 VDD.n4696 VDD.n4695 3.76521
R13228 VDD.n4519 VDD.n4518 3.76521
R13229 VDD.n4591 VDD.n4589 3.76521
R13230 VDD.n4714 VDD.n4712 3.76521
R13231 VDD.n5118 VDD.n3813 3.76521
R13232 VDD.n4530 VDD.n4529 3.76521
R13233 VDD.n4571 VDD.n4568 3.76521
R13234 VDD.n4719 VDD.n4718 3.76521
R13235 VDD.n4763 VDD.n4761 3.76521
R13236 VDD.n3196 VDD.n3184 3.76521
R13237 VDD.n3617 VDD.n3605 3.76521
R13238 VDD.n3477 VDD.n3465 3.76521
R13239 VDD.n18 VDD.n8 3.76521
R13240 VDD.n337 VDD.n327 3.76521
R13241 VDD.n316 VDD.n315 3.76521
R13242 VDD.n201 VDD.n193 3.76521
R13243 VDD.n551 VDD.n550 3.76521
R13244 VDD.n2060 VDD.n1410 3.76521
R13245 VDD.n2102 VDD.n2101 3.76521
R13246 VDD.n1925 VDD.n1924 3.76521
R13247 VDD.n1997 VDD.n1995 3.76521
R13248 VDD.n2120 VDD.n2118 3.76521
R13249 VDD.n2524 VDD.n1219 3.76521
R13250 VDD.n1936 VDD.n1935 3.76521
R13251 VDD.n1977 VDD.n1974 3.76521
R13252 VDD.n2125 VDD.n2124 3.76521
R13253 VDD.n2169 VDD.n2167 3.76521
R13254 VDD.n602 VDD.n590 3.76521
R13255 VDD.n1023 VDD.n1011 3.76521
R13256 VDD.n883 VDD.n871 3.76521
R13257 VDD.n5581 VDD.n5571 3.76521
R13258 VDD.n5900 VDD.n5890 3.76521
R13259 VDD.n5879 VDD.n5878 3.76521
R13260 VDD.n5764 VDD.n5756 3.76521
R13261 VDD.n5554 VDD.n5464 3.76521
R13262 VDD.n5531 VDD.n5472 3.76521
R13263 VDD.n5520 VDD.n5519 3.76521
R13264 VDD.n5499 VDD.n5498 3.76521
R13265 VDD.n5436 VDD.n5315 3.76521
R13266 VDD.n5380 VDD.n5335 3.76521
R13267 VDD.n5354 VDD.n5353 3.76521
R13268 VDD.n6114 VDD.n6113 3.76521
R13269 VDD.n7623 VDD.n6973 3.76521
R13270 VDD.n7665 VDD.n7664 3.76521
R13271 VDD.n7488 VDD.n7487 3.76521
R13272 VDD.n7560 VDD.n7558 3.76521
R13273 VDD.n7683 VDD.n7681 3.76521
R13274 VDD.n8087 VDD.n6782 3.76521
R13275 VDD.n7499 VDD.n7498 3.76521
R13276 VDD.n7540 VDD.n7537 3.76521
R13277 VDD.n7688 VDD.n7687 3.76521
R13278 VDD.n7732 VDD.n7730 3.76521
R13279 VDD.n6165 VDD.n6153 3.76521
R13280 VDD.n6586 VDD.n6574 3.76521
R13281 VDD.n6446 VDD.n6434 3.76521
R13282 VDD.n4431 VDD.t400 3.6005
R13283 VDD.n5114 VDD.t601 3.6005
R13284 VDD.n1837 VDD.t50 3.6005
R13285 VDD.n2520 VDD.t246 3.6005
R13286 VDD.n7400 VDD.t297 3.6005
R13287 VDD.n8083 VDD.t559 3.6005
R13288 VDD.n4731 VDD.n4730 3.59719
R13289 VDD.n4730 VDD.n3923 3.59719
R13290 VDD.n4742 VDD.n3923 3.59719
R13291 VDD.n4745 VDD.n4744 3.59719
R13292 VDD.n4744 VDD.n3831 3.59719
R13293 VDD.n5106 VDD.n3831 3.59719
R13294 VDD.n4493 VDD.n4102 3.59719
R13295 VDD.n4102 VDD.n4065 3.59719
R13296 VDD.n4065 VDD.n3435 3.59719
R13297 VDD.n5158 VDD.n3437 3.59719
R13298 VDD.n4055 VDD.n3437 3.59719
R13299 VDD.n4579 VDD.n4055 3.59719
R13300 VDD.n2137 VDD.n2136 3.59719
R13301 VDD.n2136 VDD.n1329 3.59719
R13302 VDD.n2148 VDD.n1329 3.59719
R13303 VDD.n2151 VDD.n2150 3.59719
R13304 VDD.n2150 VDD.n1237 3.59719
R13305 VDD.n2512 VDD.n1237 3.59719
R13306 VDD.n1899 VDD.n1508 3.59719
R13307 VDD.n1508 VDD.n1471 3.59719
R13308 VDD.n1471 VDD.n841 3.59719
R13309 VDD.n2564 VDD.n843 3.59719
R13310 VDD.n1461 VDD.n843 3.59719
R13311 VDD.n1985 VDD.n1461 3.59719
R13312 VDD.n7700 VDD.n7699 3.59719
R13313 VDD.n7699 VDD.n6892 3.59719
R13314 VDD.n7711 VDD.n6892 3.59719
R13315 VDD.n7714 VDD.n7713 3.59719
R13316 VDD.n7713 VDD.n6800 3.59719
R13317 VDD.n8075 VDD.n6800 3.59719
R13318 VDD.n7462 VDD.n7071 3.59719
R13319 VDD.n7071 VDD.n7034 3.59719
R13320 VDD.n7034 VDD.n6404 3.59719
R13321 VDD.n8127 VDD.n6406 3.59719
R13322 VDD.n7024 VDD.n6406 3.59719
R13323 VDD.n7548 VDD.n7024 3.59719
R13324 VDD.n2939 VDD.n2938 3.49275
R13325 VDD.n345 VDD.n344 3.49275
R13326 VDD.n5908 VDD.n5907 3.49275
R13327 VDD.n5561 VDD.n5461 3.49141
R13328 VDD.n3211 VDD.n3178 3.44003
R13329 VDD.n3285 VDD.n3281 3.44003
R13330 VDD.n3298 VDD.n3280 3.44003
R13331 VDD.n3311 VDD.n3279 3.44003
R13332 VDD.n3324 VDD.n3278 3.44003
R13333 VDD.n3268 VDD.n3264 3.44003
R13334 VDD.n3254 VDD.n3250 3.44003
R13335 VDD.n3240 VDD.n3236 3.44003
R13336 VDD.n3226 VDD.n3222 3.44003
R13337 VDD.n3167 VDD.n3163 3.44003
R13338 VDD.n617 VDD.n584 3.44003
R13339 VDD.n691 VDD.n687 3.44003
R13340 VDD.n704 VDD.n686 3.44003
R13341 VDD.n717 VDD.n685 3.44003
R13342 VDD.n730 VDD.n684 3.44003
R13343 VDD.n674 VDD.n670 3.44003
R13344 VDD.n660 VDD.n656 3.44003
R13345 VDD.n646 VDD.n642 3.44003
R13346 VDD.n632 VDD.n628 3.44003
R13347 VDD.n573 VDD.n569 3.44003
R13348 VDD.n6180 VDD.n6147 3.44003
R13349 VDD.n6254 VDD.n6250 3.44003
R13350 VDD.n6267 VDD.n6249 3.44003
R13351 VDD.n6280 VDD.n6248 3.44003
R13352 VDD.n6293 VDD.n6247 3.44003
R13353 VDD.n6237 VDD.n6233 3.44003
R13354 VDD.n6223 VDD.n6219 3.44003
R13355 VDD.n6209 VDD.n6205 3.44003
R13356 VDD.n6195 VDD.n6191 3.44003
R13357 VDD.n6136 VDD.n6132 3.44003
R13358 VDD.n3160 VDD.n3159 3.42232
R13359 VDD.n3393 VDD.n3392 3.42232
R13360 VDD.n3406 VDD.n3405 3.42232
R13361 VDD.n3419 VDD.n3418 3.42232
R13362 VDD.n3432 VDD.n3431 3.42232
R13363 VDD.n3376 VDD.n3375 3.42232
R13364 VDD.n3362 VDD.n3361 3.42232
R13365 VDD.n3348 VDD.n3347 3.42232
R13366 VDD.n3116 VDD.n3115 3.42232
R13367 VDD.n5173 VDD.n5172 3.42232
R13368 VDD.n566 VDD.n565 3.42232
R13369 VDD.n799 VDD.n798 3.42232
R13370 VDD.n812 VDD.n811 3.42232
R13371 VDD.n825 VDD.n824 3.42232
R13372 VDD.n838 VDD.n837 3.42232
R13373 VDD.n782 VDD.n781 3.42232
R13374 VDD.n768 VDD.n767 3.42232
R13375 VDD.n754 VDD.n753 3.42232
R13376 VDD.n522 VDD.n521 3.42232
R13377 VDD.n2579 VDD.n2578 3.42232
R13378 VDD.n6129 VDD.n6128 3.42232
R13379 VDD.n6362 VDD.n6361 3.42232
R13380 VDD.n6375 VDD.n6374 3.42232
R13381 VDD.n6388 VDD.n6387 3.42232
R13382 VDD.n6401 VDD.n6400 3.42232
R13383 VDD.n6345 VDD.n6344 3.42232
R13384 VDD.n6331 VDD.n6330 3.42232
R13385 VDD.n6317 VDD.n6316 3.42232
R13386 VDD.n6085 VDD.n6084 3.42232
R13387 VDD.n8142 VDD.n8141 3.42232
R13388 VDD.n2914 VDD.n2913 3.41442
R13389 VDD.n320 VDD.n319 3.41442
R13390 VDD.n5883 VDD.n5882 3.41442
R13391 VDD.n2792 VDD.n2599 3.4105
R13392 VDD.n198 VDD.n5 3.4105
R13393 VDD.n5761 VDD.n5568 3.4105
R13394 VDD.n4457 VDD.t625 3.4005
R13395 VDD.n3911 VDD.t402 3.4005
R13396 VDD.n1863 VDD.t468 3.4005
R13397 VDD.n1317 VDD.t228 3.4005
R13398 VDD.n7426 VDD.t167 3.4005
R13399 VDD.n6880 VDD.t152 3.4005
R13400 VDD.n3632 VDD.n3599 3.389
R13401 VDD.n3646 VDD.n3598 3.389
R13402 VDD.n3659 VDD.n3597 3.389
R13403 VDD.n3672 VDD.n3596 3.389
R13404 VDD.n3685 VDD.n3595 3.389
R13405 VDD.n3698 VDD.n3594 3.389
R13406 VDD.n3711 VDD.n3593 3.389
R13407 VDD.n3725 VDD.n3592 3.389
R13408 VDD.n3738 VDD.n3591 3.389
R13409 VDD.n3751 VDD.n3590 3.389
R13410 VDD.n3764 VDD.n3589 3.389
R13411 VDD.n3777 VDD.n3588 3.389
R13412 VDD.n3578 VDD.n3574 3.389
R13413 VDD.n3564 VDD.n3560 3.389
R13414 VDD.n3550 VDD.n3546 3.389
R13415 VDD.n3536 VDD.n3532 3.389
R13416 VDD.n3522 VDD.n3518 3.389
R13417 VDD.n3508 VDD.n3504 3.389
R13418 VDD.n3493 VDD.n3489 3.389
R13419 VDD.n1038 VDD.n1005 3.389
R13420 VDD.n1052 VDD.n1004 3.389
R13421 VDD.n1065 VDD.n1003 3.389
R13422 VDD.n1078 VDD.n1002 3.389
R13423 VDD.n1091 VDD.n1001 3.389
R13424 VDD.n1104 VDD.n1000 3.389
R13425 VDD.n1117 VDD.n999 3.389
R13426 VDD.n1131 VDD.n998 3.389
R13427 VDD.n1144 VDD.n997 3.389
R13428 VDD.n1157 VDD.n996 3.389
R13429 VDD.n1170 VDD.n995 3.389
R13430 VDD.n1183 VDD.n994 3.389
R13431 VDD.n984 VDD.n980 3.389
R13432 VDD.n970 VDD.n966 3.389
R13433 VDD.n956 VDD.n952 3.389
R13434 VDD.n942 VDD.n938 3.389
R13435 VDD.n928 VDD.n924 3.389
R13436 VDD.n914 VDD.n910 3.389
R13437 VDD.n899 VDD.n895 3.389
R13438 VDD.n6601 VDD.n6568 3.389
R13439 VDD.n6615 VDD.n6567 3.389
R13440 VDD.n6628 VDD.n6566 3.389
R13441 VDD.n6641 VDD.n6565 3.389
R13442 VDD.n6654 VDD.n6564 3.389
R13443 VDD.n6667 VDD.n6563 3.389
R13444 VDD.n6680 VDD.n6562 3.389
R13445 VDD.n6694 VDD.n6561 3.389
R13446 VDD.n6707 VDD.n6560 3.389
R13447 VDD.n6720 VDD.n6559 3.389
R13448 VDD.n6733 VDD.n6558 3.389
R13449 VDD.n6746 VDD.n6557 3.389
R13450 VDD.n6547 VDD.n6543 3.389
R13451 VDD.n6533 VDD.n6529 3.389
R13452 VDD.n6519 VDD.n6515 3.389
R13453 VDD.n6505 VDD.n6501 3.389
R13454 VDD.n6491 VDD.n6487 3.389
R13455 VDD.n6477 VDD.n6473 3.389
R13456 VDD.n6462 VDD.n6458 3.389
R13457 VDD.n4731 VDD.n4729 3.38562
R13458 VDD.n2137 VDD.n2135 3.38562
R13459 VDD.n7700 VDD.n7698 3.38562
R13460 VDD.n5216 VDD 3.38175
R13461 VDD.n2658 VDD.n2657 3.2005
R13462 VDD.n2998 VDD.n2997 3.2005
R13463 VDD.n4484 VDD.t421 3.2005
R13464 VDD.n4990 VDD.t599 3.2005
R13465 VDD.n64 VDD.n63 3.2005
R13466 VDD.n404 VDD.n403 3.2005
R13467 VDD.n1890 VDD.t95 3.2005
R13468 VDD.n2396 VDD.t346 3.2005
R13469 VDD.n5627 VDD.n5626 3.2005
R13470 VDD.n5967 VDD.n5966 3.2005
R13471 VDD.n7453 VDD.t43 3.2005
R13472 VDD.n7959 VDD.t40 3.2005
R13473 VDD.n5188 VDD 3.13175
R13474 VDD.t605 VDD.n4142 3.0005
R13475 VDD.t437 VDD.n5101 3.0005
R13476 VDD.t613 VDD.n3908 3.0005
R13477 VDD.t348 VDD.n1548 3.0005
R13478 VDD.t360 VDD.n2507 3.0005
R13479 VDD.t336 VDD.n1314 3.0005
R13480 VDD.t207 VDD.n7111 3.0005
R13481 VDD.t61 VDD.n8070 3.0005
R13482 VDD.t318 VDD.n6877 3.0005
R13483 VDD.n4580 VDD.n4579 2.96248
R13484 VDD.n1986 VDD.n1985 2.96248
R13485 VDD.n7549 VDD.n7548 2.96248
R13486 VDD.t405 VDD.n3452 2.8005
R13487 VDD.t91 VDD.n858 2.8005
R13488 VDD.t0 VDD.n6421 2.8005
R13489 VDD.n4745 VDD.n3118 2.69802
R13490 VDD.n2151 VDD.n524 2.69802
R13491 VDD.n7714 VDD.n6087 2.69802
R13492 VDD.n5196 VDD 2.69321
R13493 VDD.n4248 VDD.t645 2.6005
R13494 VDD.n4286 VDD.t649 2.6005
R13495 VDD.n3924 VDD.t394 2.6005
R13496 VDD.n4928 VDD.t595 2.6005
R13497 VDD.n4904 VDD.t623 2.6005
R13498 VDD.n1654 VDD.t79 2.6005
R13499 VDD.n1692 VDD.t4 2.6005
R13500 VDD.n1330 VDD.t89 2.6005
R13501 VDD.n2334 VDD.t357 2.6005
R13502 VDD.n2310 VDD.t516 2.6005
R13503 VDD.n7217 VDD.t255 2.6005
R13504 VDD.n7255 VDD.t264 2.6005
R13505 VDD.n6893 VDD.t165 2.6005
R13506 VDD.n7897 VDD.t322 2.6005
R13507 VDD.n7873 VDD.t179 2.6005
R13508 VDD.n5511 VDD.n5480 2.58636
R13509 VDD.n2901 VDD.n2755 2.5605
R13510 VDD.n2835 VDD.n2782 2.5605
R13511 VDD.n307 VDD.n161 2.5605
R13512 VDD.n241 VDD.n188 2.5605
R13513 VDD.n5870 VDD.n5724 2.5605
R13514 VDD.n5804 VDD.n5751 2.5605
R13515 VDD.n5245 VDD 2.48488
R13516 VDD.n4652 VDD.t431 2.4005
R13517 VDD.n2058 VDD.t193 2.4005
R13518 VDD.n7621 VDD.t48 2.4005
R13519 VDD.n5159 VDD.n3435 2.27488
R13520 VDD.n2565 VDD.n841 2.27488
R13521 VDD.n8128 VDD.n6404 2.27488
R13522 VDD.n2611 VDD.n2604 2.25932
R13523 VDD.n2930 VDD.n2923 2.25932
R13524 VDD.n2906 VDD.n2744 2.25932
R13525 VDD.n2827 VDD.n2826 2.25932
R13526 VDD.n3141 VDD.n3124 2.25932
R13527 VDD.n4656 VDD.n4655 2.25932
R13528 VDD.n3999 VDD.n3969 2.25932
R13529 VDD.n4516 VDD.n4515 2.25932
R13530 VDD.n4048 VDD.n3456 2.25932
R13531 VDD.n4713 VDD.n3792 2.25932
R13532 VDD.n5122 VDD.n5121 2.25932
R13533 VDD.n4074 VDD.n3448 2.25932
R13534 VDD.n4567 VDD.n4566 2.25932
R13535 VDD.n3949 VDD.n3945 2.25932
R13536 VDD.n5126 VDD.n3807 2.25932
R13537 VDD.n3193 VDD.n3192 2.25932
R13538 VDD.n3614 VDD.n3613 2.25932
R13539 VDD.n3474 VDD.n3473 2.25932
R13540 VDD.n17 VDD.n10 2.25932
R13541 VDD.n336 VDD.n329 2.25932
R13542 VDD.n312 VDD.n150 2.25932
R13543 VDD.n233 VDD.n232 2.25932
R13544 VDD.n547 VDD.n530 2.25932
R13545 VDD.n2062 VDD.n2061 2.25932
R13546 VDD.n1405 VDD.n1375 2.25932
R13547 VDD.n1922 VDD.n1921 2.25932
R13548 VDD.n1454 VDD.n862 2.25932
R13549 VDD.n2119 VDD.n1198 2.25932
R13550 VDD.n2528 VDD.n2527 2.25932
R13551 VDD.n1480 VDD.n854 2.25932
R13552 VDD.n1973 VDD.n1972 2.25932
R13553 VDD.n1355 VDD.n1351 2.25932
R13554 VDD.n2532 VDD.n1213 2.25932
R13555 VDD.n599 VDD.n598 2.25932
R13556 VDD.n1020 VDD.n1019 2.25932
R13557 VDD.n880 VDD.n879 2.25932
R13558 VDD.n5580 VDD.n5573 2.25932
R13559 VDD.n5899 VDD.n5892 2.25932
R13560 VDD.n5875 VDD.n5713 2.25932
R13561 VDD.n5796 VDD.n5795 2.25932
R13562 VDD.n6110 VDD.n6093 2.25932
R13563 VDD.n7625 VDD.n7624 2.25932
R13564 VDD.n6968 VDD.n6938 2.25932
R13565 VDD.n7485 VDD.n7484 2.25932
R13566 VDD.n7017 VDD.n6425 2.25932
R13567 VDD.n7682 VDD.n6761 2.25932
R13568 VDD.n8091 VDD.n8090 2.25932
R13569 VDD.n7043 VDD.n6417 2.25932
R13570 VDD.n7536 VDD.n7535 2.25932
R13571 VDD.n6918 VDD.n6914 2.25932
R13572 VDD.n8095 VDD.n6776 2.25932
R13573 VDD.n6162 VDD.n6161 2.25932
R13574 VDD.n6583 VDD.n6582 2.25932
R13575 VDD.n6443 VDD.n6442 2.25932
R13576 VDD.t621 VDD.n4188 2.2005
R13577 VDD.n4266 VDD.t609 2.2005
R13578 VDD.t419 VDD.n3964 2.2005
R13579 VDD.t661 VDD.n4919 2.2005
R13580 VDD.t641 VDD.n4824 2.2005
R13581 VDD.t6 VDD.n1594 2.2005
R13582 VDD.n1672 VDD.t174 2.2005
R13583 VDD.t148 VDD.n1370 2.2005
R13584 VDD.t221 VDD.n2325 2.2005
R13585 VDD.t36 VDD.n2230 2.2005
R13586 VDD.t158 VDD.n7157 2.2005
R13587 VDD.n7235 VDD.t8 2.2005
R13588 VDD.t141 VDD.n6933 2.2005
R13589 VDD.t509 VDD.n7888 2.2005
R13590 VDD.t283 VDD.n7793 2.2005
R13591 VDD.t528 VDD.n5404 2.11161
R13592 VDD.n5422 VDD.n5421 2.02977
R13593 VDD.n5362 VDD.n5340 2.02977
R13594 VDD.n4494 VDD.n4493 2.01042
R13595 VDD.n1900 VDD.n1899 2.01042
R13596 VDD.n7463 VDD.n7462 2.01042
R13597 VDD.n4705 VDD.t410 2.0005
R13598 VDD.n2111 VDD.t52 2.0005
R13599 VDD.n7674 VDD.t579 2.0005
R13600 VDD.n5562 VDD.n5561 1.93989
R13601 VDD.n5160 VDD.n5159 1.846
R13602 VDD.n2566 VDD.n2565 1.846
R13603 VDD.n8129 VDD.n8128 1.846
R13604 VDD.n5160 VDD.n3118 1.84324
R13605 VDD.n2566 VDD.n524 1.84324
R13606 VDD.n8129 VDD.n6087 1.84324
R13607 VDD.n4292 VDD.t631 1.8005
R13608 VDD.n4605 VDD.t398 1.8005
R13609 VDD.t633 VDD.n4934 1.8005
R13610 VDD.n1698 VDD.t97 1.8005
R13611 VDD.n2011 VDD.t81 1.8005
R13612 VDD.t501 VDD.n2340 1.8005
R13613 VDD.n7261 VDD.t156 1.8005
R13614 VDD.n7574 VDD.t230 1.8005
R13615 VDD.t268 VDD.n7903 1.8005
R13616 VDD.n2940 VDD.n2939 1.74685
R13617 VDD.n346 VDD.n345 1.74685
R13618 VDD.n5909 VDD.n5908 1.74685
R13619 VDD.n5515 VDD.n5514 1.68131
R13620 VDD.n5514 VDD.n5479 1.68131
R13621 VDD.n4747 VDD.t427 1.6005
R13622 VDD.n2153 VDD.t195 1.6005
R13623 VDD.n7716 VDD.t216 1.6005
R13624 VDD.n5106 VDD.n5105 1.58728
R13625 VDD.n2512 VDD.n2511 1.58728
R13626 VDD.n8075 VDD.n8074 1.58728
R13627 VDD.n5407 VDD.n5322 1.56148
R13628 VDD.n4729 VDD.n4728 1.50638
R13629 VDD.n4729 VDD.n3930 1.50638
R13630 VDD.n2135 VDD.n2134 1.50638
R13631 VDD.n2135 VDD.n1336 1.50638
R13632 VDD.n7698 VDD.n7697 1.50638
R13633 VDD.n7698 VDD.n6899 1.50638
R13634 VDD.n3101 VDD.n2599 1.48637
R13635 VDD.n507 VDD.n5 1.48637
R13636 VDD.n6070 VDD.n5568 1.48637
R13637 VDD.n4561 VDD.n4560 1.41953
R13638 VDD.n4560 VDD.n4559 1.41953
R13639 VDD.n5141 VDD.n5140 1.41953
R13640 VDD.n5140 VDD.n5139 1.41953
R13641 VDD.n1967 VDD.n1966 1.41953
R13642 VDD.n1966 VDD.n1965 1.41953
R13643 VDD.n2547 VDD.n2546 1.41953
R13644 VDD.n2546 VDD.n2545 1.41953
R13645 VDD.n7530 VDD.n7529 1.41953
R13646 VDD.n7529 VDD.n7528 1.41953
R13647 VDD.n8110 VDD.n8109 1.41953
R13648 VDD.n8109 VDD.n8108 1.41953
R13649 VDD.t413 VDD.n4063 1.4005
R13650 VDD.t635 VDD.n3886 1.4005
R13651 VDD.t334 VDD.n1469 1.4005
R13652 VDD.t189 VDD.n1292 1.4005
R13653 VDD.t2 VDD.n7032 1.4005
R13654 VDD.t341 VDD.n6855 1.4005
R13655 VDD.n5159 VDD.n5158 1.32281
R13656 VDD.n2565 VDD.n2564 1.32281
R13657 VDD.n8128 VDD.n8127 1.32281
R13658 VDD.n2902 VDD.n2749 1.2805
R13659 VDD.n2822 VDD.n2817 1.2805
R13660 VDD.n308 VDD.n155 1.2805
R13661 VDD.n228 VDD.n223 1.2805
R13662 VDD.n5871 VDD.n5718 1.2805
R13663 VDD.n5791 VDD.n5786 1.2805
R13664 VDD.n4386 VDD.t653 1.2005
R13665 VDD.n5091 VDD.t424 1.2005
R13666 VDD.n1792 VDD.t452 1.2005
R13667 VDD.n2497 VDD.t146 1.2005
R13668 VDD.n7355 VDD.t373 1.2005
R13669 VDD.n8060 VDD.t22 1.2005
R13670 VDD.n5524 VDD.n5523 1.12991
R13671 VDD.n5535 VDD.n5470 1.12991
R13672 VDD.n5403 VDD.n5325 1.09318
R13673 VDD.n5488 VDD.n5485 1.07033
R13674 VDD.n5347 VDD.n5346 1.07033
R13675 VDD.t429 VDD.n4110 1.0005
R13676 VDD.n4768 VDD.t615 1.0005
R13677 VDD.t99 VDD.n1516 1.0005
R13678 VDD.n2174 VDD.t454 1.0005
R13679 VDD.t38 VDD.n7079 1.0005
R13680 VDD.n7737 VDD.t181 1.0005
R13681 VDD.n5293 VDD.n5288 1.0005
R13682 VDD.n3642 VDD.n3459 0.926359
R13683 VDD.n3788 VDD.n3503 0.926359
R13684 VDD.n1048 VDD.n865 0.926359
R13685 VDD.n1194 VDD.n909 0.926359
R13686 VDD.n6611 VDD.n6428 0.926359
R13687 VDD.n6757 VDD.n6472 0.926359
R13688 VDD.n5539 VDD.n5538 0.90555
R13689 VDD.n4742 VDD.n3118 0.899674
R13690 VDD.n2148 VDD.n524 0.899674
R13691 VDD.n7711 VDD.n6087 0.899674
R13692 VDD.n5161 VDD.n5160 0.83012
R13693 VDD.n2567 VDD.n2566 0.83012
R13694 VDD.n8130 VDD.n8129 0.83012
R13695 VDD.n3335 VDD.n3177 0.817389
R13696 VDD.n741 VDD.n583 0.817389
R13697 VDD.n6304 VDD.n6146 0.817389
R13698 VDD.n5160 VDD.n3162 0.813764
R13699 VDD.n2566 VDD.n568 0.813764
R13700 VDD.n8129 VDD.n6131 0.813764
R13701 VDD.n3335 VDD.n3221 0.805608
R13702 VDD.n741 VDD.n627 0.805608
R13703 VDD.n6304 VDD.n6190 0.805608
R13704 VDD.n4499 VDD.t603 0.8005
R13705 VDD.n1905 VDD.t498 0.8005
R13706 VDD.n7468 VDD.t561 0.8005
R13707 VDD.n5245 VDD.n5244 0.78925
R13708 VDD.n5160 VDD.n3434 0.764222
R13709 VDD.n2566 VDD.n840 0.764222
R13710 VDD.n8129 VDD.n6403 0.764222
R13711 VDD.n3721 VDD.n3459 0.759389
R13712 VDD.n3788 VDD.n3787 0.759389
R13713 VDD.n3335 VDD.n3334 0.759389
R13714 VDD.n1127 VDD.n865 0.759389
R13715 VDD.n1194 VDD.n1193 0.759389
R13716 VDD.n741 VDD.n740 0.759389
R13717 VDD.n6690 VDD.n6428 0.759389
R13718 VDD.n6757 VDD.n6756 0.759389
R13719 VDD.n6304 VDD.n6303 0.759389
R13720 VDD.n2608 VDD.n2607 0.753441
R13721 VDD.n2927 VDD.n2926 0.753441
R13722 VDD.n2905 VDD.n2746 0.753441
R13723 VDD.n2752 VDD.n2751 0.753441
R13724 VDD.n2830 VDD.n2785 0.753441
R13725 VDD.n2832 VDD.n2831 0.753441
R13726 VDD.n3140 VDD.n3137 0.753441
R13727 VDD.n4669 VDD.n3998 0.753441
R13728 VDD.n4668 VDD.n4667 0.753441
R13729 VDD.n5145 VDD.n3455 0.753441
R13730 VDD.n5144 VDD.n5143 0.753441
R13731 VDD.n5137 VDD.n5136 0.753441
R13732 VDD.n3812 VDD.n3793 0.753441
R13733 VDD.n5150 VDD.n5149 0.753441
R13734 VDD.n4564 VDD.n3449 0.753441
R13735 VDD.n3948 VDD.n3947 0.753441
R13736 VDD.n5127 VDD.n3806 0.753441
R13737 VDD.n3189 VDD.n3186 0.753441
R13738 VDD.n3610 VDD.n3607 0.753441
R13739 VDD.n3470 VDD.n3467 0.753441
R13740 VDD.n14 VDD.n13 0.753441
R13741 VDD.n333 VDD.n332 0.753441
R13742 VDD.n311 VDD.n152 0.753441
R13743 VDD.n158 VDD.n157 0.753441
R13744 VDD.n236 VDD.n191 0.753441
R13745 VDD.n238 VDD.n237 0.753441
R13746 VDD.n546 VDD.n543 0.753441
R13747 VDD.n2075 VDD.n1404 0.753441
R13748 VDD.n2074 VDD.n2073 0.753441
R13749 VDD.n2551 VDD.n861 0.753441
R13750 VDD.n2550 VDD.n2549 0.753441
R13751 VDD.n2543 VDD.n2542 0.753441
R13752 VDD.n1218 VDD.n1199 0.753441
R13753 VDD.n2556 VDD.n2555 0.753441
R13754 VDD.n1970 VDD.n855 0.753441
R13755 VDD.n1354 VDD.n1353 0.753441
R13756 VDD.n2533 VDD.n1212 0.753441
R13757 VDD.n595 VDD.n592 0.753441
R13758 VDD.n1016 VDD.n1013 0.753441
R13759 VDD.n876 VDD.n873 0.753441
R13760 VDD.n5577 VDD.n5576 0.753441
R13761 VDD.n5896 VDD.n5895 0.753441
R13762 VDD.n5874 VDD.n5715 0.753441
R13763 VDD.n5721 VDD.n5720 0.753441
R13764 VDD.n5799 VDD.n5754 0.753441
R13765 VDD.n5801 VDD.n5800 0.753441
R13766 VDD.n5545 VDD.n5462 0.753441
R13767 VDD.n5522 VDD.n5470 0.753441
R13768 VDD.n6109 VDD.n6106 0.753441
R13769 VDD.n7638 VDD.n6967 0.753441
R13770 VDD.n7637 VDD.n7636 0.753441
R13771 VDD.n8114 VDD.n6424 0.753441
R13772 VDD.n8113 VDD.n8112 0.753441
R13773 VDD.n8106 VDD.n8105 0.753441
R13774 VDD.n6781 VDD.n6762 0.753441
R13775 VDD.n8119 VDD.n8118 0.753441
R13776 VDD.n7533 VDD.n6418 0.753441
R13777 VDD.n6917 VDD.n6916 0.753441
R13778 VDD.n8096 VDD.n6775 0.753441
R13779 VDD.n6158 VDD.n6155 0.753441
R13780 VDD.n6579 VDD.n6576 0.753441
R13781 VDD.n6439 VDD.n6436 0.753441
R13782 VDD.n5223 VDD.n5215 0.708
R13783 VDD.n5280 VDD.n5275 0.708
R13784 VDD.n5124 VDD.t619 0.6005
R13785 VDD.n2530 VDD.t324 0.6005
R13786 VDD.n8093 VDD.t370 0.6005
R13787 VDD.n5310 VDD 0.516125
R13788 VDD.n5440 VDD 0.505708
R13789 VDD.n5244 VDD.n5189 0.5005
R13790 VDD.n5233 VDD.n5189 0.5005
R13791 VDD.n5234 VDD.n5233 0.5005
R13792 VDD.n5223 VDD.n5222 0.5005
R13793 VDD.n5222 VDD.n5221 0.5005
R13794 VDD.n5221 VDD.n5217 0.5005
R13795 VDD.n5280 VDD.n5279 0.5005
R13796 VDD.n5279 VDD.n5278 0.5005
R13797 VDD.n5278 VDD.n5255 0.5005
R13798 VDD.n5288 VDD.n5255 0.5005
R13799 VDD.n5293 VDD.n5292 0.5005
R13800 VDD.n5292 VDD.n5291 0.5005
R13801 VDD.n5291 VDD.n5248 0.5005
R13802 VDD.n5407 VDD.n5406 0.468793
R13803 VDD.n5235 VDD.n5234 0.44925
R13804 VDD.n5301 VDD.n5248 0.44925
R13805 VDD.n2790 VDD.n2599 0.404062
R13806 VDD.n196 VDD.n5 0.404062
R13807 VDD.n5759 VDD.n5568 0.404062
R13808 VDD.n5156 VDD.t589 0.4005
R13809 VDD.n2562 VDD.t701 0.4005
R13810 VDD.n8125 VDD.t176 0.4005
R13811 VDD.n3102 VDD.n3101 0.39283
R13812 VDD.n508 VDD.n507 0.39283
R13813 VDD.n6071 VDD.n6070 0.39283
R13814 VDD.n2914 VDD 0.390922
R13815 VDD.n320 VDD 0.390922
R13816 VDD.n5883 VDD 0.390922
R13817 VDD.n5501 VDD.n5480 0.388379
R13818 VDD.n5175 VDD.n5174 0.385322
R13819 VDD.n2581 VDD.n2580 0.385322
R13820 VDD.n8144 VDD.n8143 0.385322
R13821 VDD.n5309 VDD.n5303 0.3805
R13822 VDD.n5309 VDD.n5304 0.3805
R13823 VDD.n5309 VDD.n5308 0.3805
R13824 VDD.n5308 VDD.n5307 0.3805
R13825 VDD.n8151 VDD.n8150 0.3805
R13826 VDD.n8151 VDD.n5180 0.3805
R13827 VDD.n8146 VDD.n5180 0.3805
R13828 VDD.n8148 VDD.n8147 0.3805
R13829 VDD.n8147 VDD.n8146 0.3805
R13830 VDD.n8148 VDD.n5183 0.3805
R13831 VDD.n8146 VDD.n5183 0.3805
R13832 VDD.n8146 VDD.n8145 0.3805
R13833 VDD.n8155 VDD.n8154 0.3805
R13834 VDD.n8155 VDD.n2585 0.3805
R13835 VDD.n8152 VDD.n2585 0.3805
R13836 VDD.n8157 VDD.n3 0.3805
R13837 VDD.n8152 VDD.n3 0.3805
R13838 VDD.n8157 VDD.n1 0.3805
R13839 VDD.n8152 VDD.n1 0.3805
R13840 VDD.n8152 VDD.n2582 0.3805
R13841 VDD.n2597 VDD.n2596 0.3805
R13842 VDD.n2597 VDD.n2587 0.3805
R13843 VDD.n5177 VDD.n2587 0.3805
R13844 VDD.n2593 VDD.n2589 0.3805
R13845 VDD.n5177 VDD.n2589 0.3805
R13846 VDD.n2593 VDD.n2586 0.3805
R13847 VDD.n5177 VDD.n2586 0.3805
R13848 VDD.n5177 VDD.n5176 0.3805
R13849 VDD.n2939 VDD.n2914 0.323981
R13850 VDD.n345 VDD.n320 0.323981
R13851 VDD.n5908 VDD.n5883 0.323981
R13852 VDD.t75 VDD.n2634 0.323629
R13853 VDD.n3022 VDD.t73 0.323629
R13854 VDD.t121 VDD.n40 0.323629
R13855 VDD.n428 VDD.t123 0.323629
R13856 VDD.t161 VDD.n5603 0.323629
R13857 VDD.n5991 VDD.t198 0.323629
R13858 VDD.n5217 VDD.n5216 0.31175
R13859 VDD.n5311 VDD 0.285624
R13860 VDD.n5303 VDD.n5302 0.280336
R13861 VDD VDD.n5309 0.260645
R13862 VDD.n5235 VDD 0.24425
R13863 VDD VDD.n5301 0.24425
R13864 VDD.n5207 VDD.n5206 0.238
R13865 VDD.n5206 VDD.n5200 0.238
R13866 VDD.n5267 VDD.n5266 0.238
R13867 VDD.n5266 VDD.n5260 0.238
R13868 VDD.n5441 VDD 0.2305
R13869 VDD.n8155 VDD.n5177 0.21365
R13870 VDD.n8152 VDD.n8151 0.21075
R13871 VDD.n2792 VDD.n2791 0.204167
R13872 VDD.n2791 VDD.n2741 0.204167
R13873 VDD.n2918 VDD.n2916 0.204167
R13874 VDD.n198 VDD.n197 0.204167
R13875 VDD.n197 VDD.n147 0.204167
R13876 VDD.n324 VDD.n322 0.204167
R13877 VDD.n5761 VDD.n5760 0.204167
R13878 VDD.n5760 VDD.n5710 0.204167
R13879 VDD.n5887 VDD.n5885 0.204167
R13880 VDD.n4386 VDD.n4354 0.2005
R13881 VDD.n4431 VDD.n4138 0.2005
R13882 VDD.n4465 VDD.n4121 0.2005
R13883 VDD.n4439 VDD.n4438 0.2005
R13884 VDD.n4472 VDD.n4114 0.2005
R13885 VDD.n4458 VDD.n4457 0.2005
R13886 VDD.n4478 VDD.n4110 0.2005
R13887 VDD.n4499 VDD.n4094 0.2005
R13888 VDD.n4484 VDD.n4107 0.2005
R13889 VDD.n4507 VDD.n4506 0.2005
R13890 VDD.n4491 VDD.n4104 0.2005
R13891 VDD.n4525 VDD.n4078 0.2005
R13892 VDD.n4536 VDD.n4066 0.2005
R13893 VDD.n4539 VDD.n4063 0.2005
R13894 VDD.n5156 VDD.n3440 0.2005
R13895 VDD.n5147 VDD.n3452 0.2005
R13896 VDD.n4549 VDD.n4059 0.2005
R13897 VDD.n4577 VDD.n4057 0.2005
R13898 VDD.n4587 VDD.n4586 0.2005
R13899 VDD.n4619 VDD.n4027 0.2005
R13900 VDD.n4605 VDD.n4043 0.2005
R13901 VDD.t629 VDD.n4023 0.2005
R13902 VDD.n4652 VDD.n4006 0.2005
R13903 VDD.n4639 VDD.n4020 0.2005
R13904 VDD.n4672 VDD.n4671 0.2005
R13905 VDD.n4645 VDD.n4017 0.2005
R13906 VDD.n4686 VDD.n3984 0.2005
R13907 VDD.n4698 VDD.n3964 0.2005
R13908 VDD.n4689 VDD.t597 0.2005
R13909 VDD.n4689 VDD.n3958 0.2005
R13910 VDD.n4706 VDD.n4705 0.2005
R13911 VDD.n4725 VDD.n3933 0.2005
R13912 VDD.n4716 VDD.n3952 0.2005
R13913 VDD.n4733 VDD.n3927 0.2005
R13914 VDD.n5134 VDD.n5133 0.2005
R13915 VDD.n4739 VDD.n3924 0.2005
R13916 VDD.n5124 VDD.n3810 0.2005
R13917 VDD.n4747 VDD.n3920 0.2005
R13918 VDD.n5115 VDD.n5114 0.2005
R13919 VDD.n4978 VDD.n4976 0.2005
R13920 VDD.n5108 VDD.n3826 0.2005
R13921 VDD.n5102 VDD.n3835 0.2005
R13922 VDD.n5101 VDD.n3838 0.2005
R13923 VDD.n4768 VDD.n3855 0.2005
R13924 VDD.n5092 VDD.n5091 0.2005
R13925 VDD.n4990 VDD.n3917 0.2005
R13926 VDD.n5085 VDD.n3867 0.2005
R13927 VDD.n4996 VDD.n3913 0.2005
R13928 VDD.n5079 VDD.n3880 0.2005
R13929 VDD.n5030 VDD.n3911 0.2005
R13930 VDD.n5073 VDD.n3886 0.2005
R13931 VDD.n1792 VDD.n1760 0.2005
R13932 VDD.n1837 VDD.n1544 0.2005
R13933 VDD.n1871 VDD.n1527 0.2005
R13934 VDD.n1845 VDD.n1844 0.2005
R13935 VDD.n1878 VDD.n1520 0.2005
R13936 VDD.n1864 VDD.n1863 0.2005
R13937 VDD.n1884 VDD.n1516 0.2005
R13938 VDD.n1905 VDD.n1500 0.2005
R13939 VDD.n1890 VDD.n1513 0.2005
R13940 VDD.n1913 VDD.n1912 0.2005
R13941 VDD.n1897 VDD.n1510 0.2005
R13942 VDD.n1931 VDD.n1484 0.2005
R13943 VDD.n1942 VDD.n1472 0.2005
R13944 VDD.n1945 VDD.n1469 0.2005
R13945 VDD.n2562 VDD.n846 0.2005
R13946 VDD.n2553 VDD.n858 0.2005
R13947 VDD.n1955 VDD.n1465 0.2005
R13948 VDD.n1983 VDD.n1463 0.2005
R13949 VDD.n1993 VDD.n1992 0.2005
R13950 VDD.n2025 VDD.n1433 0.2005
R13951 VDD.n2011 VDD.n1449 0.2005
R13952 VDD.t10 VDD.n1429 0.2005
R13953 VDD.n2058 VDD.n1412 0.2005
R13954 VDD.n2045 VDD.n1426 0.2005
R13955 VDD.n2078 VDD.n2077 0.2005
R13956 VDD.n2051 VDD.n1423 0.2005
R13957 VDD.n2092 VDD.n1390 0.2005
R13958 VDD.n2104 VDD.n1370 0.2005
R13959 VDD.n2095 VDD.t12 0.2005
R13960 VDD.n2095 VDD.n1364 0.2005
R13961 VDD.n2112 VDD.n2111 0.2005
R13962 VDD.n2131 VDD.n1339 0.2005
R13963 VDD.n2122 VDD.n1358 0.2005
R13964 VDD.n2139 VDD.n1333 0.2005
R13965 VDD.n2540 VDD.n2539 0.2005
R13966 VDD.n2145 VDD.n1330 0.2005
R13967 VDD.n2530 VDD.n1216 0.2005
R13968 VDD.n2153 VDD.n1326 0.2005
R13969 VDD.n2521 VDD.n2520 0.2005
R13970 VDD.n2384 VDD.n2382 0.2005
R13971 VDD.n2514 VDD.n1232 0.2005
R13972 VDD.n2508 VDD.n1241 0.2005
R13973 VDD.n2507 VDD.n1244 0.2005
R13974 VDD.n2174 VDD.n1261 0.2005
R13975 VDD.n2498 VDD.n2497 0.2005
R13976 VDD.n2396 VDD.n1323 0.2005
R13977 VDD.n2491 VDD.n1273 0.2005
R13978 VDD.n2402 VDD.n1319 0.2005
R13979 VDD.n2485 VDD.n1286 0.2005
R13980 VDD.n2436 VDD.n1317 0.2005
R13981 VDD.n2479 VDD.n1292 0.2005
R13982 VDD.n7355 VDD.n7323 0.2005
R13983 VDD.n7400 VDD.n7107 0.2005
R13984 VDD.n7434 VDD.n7090 0.2005
R13985 VDD.n7408 VDD.n7407 0.2005
R13986 VDD.n7441 VDD.n7083 0.2005
R13987 VDD.n7427 VDD.n7426 0.2005
R13988 VDD.n7447 VDD.n7079 0.2005
R13989 VDD.n7468 VDD.n7063 0.2005
R13990 VDD.n7453 VDD.n7076 0.2005
R13991 VDD.n7476 VDD.n7475 0.2005
R13992 VDD.n7460 VDD.n7073 0.2005
R13993 VDD.n7494 VDD.n7047 0.2005
R13994 VDD.n7505 VDD.n7035 0.2005
R13995 VDD.n7508 VDD.n7032 0.2005
R13996 VDD.n8125 VDD.n6409 0.2005
R13997 VDD.n8116 VDD.n6421 0.2005
R13998 VDD.n7518 VDD.n7028 0.2005
R13999 VDD.n7546 VDD.n7026 0.2005
R14000 VDD.n7556 VDD.n7555 0.2005
R14001 VDD.n7588 VDD.n6996 0.2005
R14002 VDD.n7574 VDD.n7012 0.2005
R14003 VDD.t316 VDD.n6992 0.2005
R14004 VDD.n7621 VDD.n6975 0.2005
R14005 VDD.n7608 VDD.n6989 0.2005
R14006 VDD.n7641 VDD.n7640 0.2005
R14007 VDD.n7614 VDD.n6986 0.2005
R14008 VDD.n7655 VDD.n6953 0.2005
R14009 VDD.n7667 VDD.n6933 0.2005
R14010 VDD.n7658 VDD.t183 0.2005
R14011 VDD.n7658 VDD.n6927 0.2005
R14012 VDD.n7675 VDD.n7674 0.2005
R14013 VDD.n7694 VDD.n6902 0.2005
R14014 VDD.n7685 VDD.n6921 0.2005
R14015 VDD.n7702 VDD.n6896 0.2005
R14016 VDD.n8103 VDD.n8102 0.2005
R14017 VDD.n7708 VDD.n6893 0.2005
R14018 VDD.n8093 VDD.n6779 0.2005
R14019 VDD.n7716 VDD.n6889 0.2005
R14020 VDD.n8084 VDD.n8083 0.2005
R14021 VDD.n7947 VDD.n7945 0.2005
R14022 VDD.n8077 VDD.n6795 0.2005
R14023 VDD.n8071 VDD.n6804 0.2005
R14024 VDD.n8070 VDD.n6807 0.2005
R14025 VDD.n7737 VDD.n6824 0.2005
R14026 VDD.n8061 VDD.n8060 0.2005
R14027 VDD.n7959 VDD.n6886 0.2005
R14028 VDD.n8054 VDD.n6836 0.2005
R14029 VDD.n7965 VDD.n6882 0.2005
R14030 VDD.n8048 VDD.n6849 0.2005
R14031 VDD.n7999 VDD.n6880 0.2005
R14032 VDD.n8042 VDD.n6855 0.2005
R14033 VDD.n2913 VDD.n2741 0.20025
R14034 VDD.n2938 VDD.n2918 0.20025
R14035 VDD.n319 VDD.n147 0.20025
R14036 VDD.n344 VDD.n324 0.20025
R14037 VDD.n5882 VDD.n5710 0.20025
R14038 VDD.n5907 VDD.n5887 0.20025
R14039 VDD.n2610 VDD.n2601 0.196152
R14040 VDD.n2610 VDD.n2609 0.196152
R14041 VDD.n2929 VDD.n2920 0.196152
R14042 VDD.n2929 VDD.n2928 0.196152
R14043 VDD.n3139 VDD.n3122 0.196152
R14044 VDD.n3130 VDD.n3121 0.196152
R14045 VDD.n3155 VDD.n3149 0.196152
R14046 VDD.n3388 VDD.n3382 0.196152
R14047 VDD.n3401 VDD.n3395 0.196152
R14048 VDD.n3414 VDD.n3408 0.196152
R14049 VDD.n3427 VDD.n3421 0.196152
R14050 VDD.n3371 VDD.n3365 0.196152
R14051 VDD.n3357 VDD.n3351 0.196152
R14052 VDD.n3343 VDD.n3337 0.196152
R14053 VDD.n3111 VDD.n3105 0.196152
R14054 VDD.n5168 VDD.n5162 0.196152
R14055 VDD.n4972 VDD.n4971 0.196152
R14056 VDD.n4971 VDD.n4767 0.196152
R14057 VDD.n4964 VDD.n4767 0.196152
R14058 VDD.n4964 VDD.n4963 0.196152
R14059 VDD.n4963 VDD.n4771 0.196152
R14060 VDD.n4775 VDD.n4771 0.196152
R14061 VDD.n4954 VDD.n4775 0.196152
R14062 VDD.n4954 VDD.n4953 0.196152
R14063 VDD.n5120 VDD.n5119 0.196152
R14064 VDD.n5119 VDD.n3814 0.196152
R14065 VDD.n3843 VDD.n3814 0.196152
R14066 VDD.n3850 VDD.n3843 0.196152
R14067 VDD.n3851 VDD.n3850 0.196152
R14068 VDD.n5097 VDD.n3851 0.196152
R14069 VDD.n5097 VDD.n5096 0.196152
R14070 VDD.n5096 VDD.n3852 0.196152
R14071 VDD.n4790 VDD.n3852 0.196152
R14072 VDD.n4790 VDD.n4787 0.196152
R14073 VDD.n4797 VDD.n4787 0.196152
R14074 VDD.n4444 VDD.n4132 0.196152
R14075 VDD.n4445 VDD.n4444 0.196152
R14076 VDD.n4453 VDD.n4445 0.196152
R14077 VDD.n4453 VDD.n4452 0.196152
R14078 VDD.n4452 VDD.n4446 0.196152
R14079 VDD.n4446 VDD.n4083 0.196152
R14080 VDD.n4512 VDD.n4083 0.196152
R14081 VDD.n4513 VDD.n4512 0.196152
R14082 VDD.n4521 VDD.n4513 0.196152
R14083 VDD.n4521 VDD.n4520 0.196152
R14084 VDD.n4520 VDD.n4514 0.196152
R14085 VDD.n4332 VDD.n4331 0.196152
R14086 VDD.n4331 VDD.n4305 0.196152
R14087 VDD.n4324 VDD.n4305 0.196152
R14088 VDD.n4324 VDD.n4323 0.196152
R14089 VDD.n4323 VDD.n4307 0.196152
R14090 VDD.n4316 VDD.n4307 0.196152
R14091 VDD.n4316 VDD.n4315 0.196152
R14092 VDD.n4315 VDD.n4311 0.196152
R14093 VDD.n3198 VDD.n3181 0.196152
R14094 VDD.n3195 VDD.n3194 0.196152
R14095 VDD.n3194 VDD.n3185 0.196152
R14096 VDD.n3212 VDD.n3209 0.196152
R14097 VDD.n3286 VDD.n3283 0.196152
R14098 VDD.n3299 VDD.n3296 0.196152
R14099 VDD.n3312 VDD.n3309 0.196152
R14100 VDD.n3325 VDD.n3322 0.196152
R14101 VDD.n3269 VDD.n3266 0.196152
R14102 VDD.n3255 VDD.n3252 0.196152
R14103 VDD.n3241 VDD.n3238 0.196152
R14104 VDD.n3227 VDD.n3224 0.196152
R14105 VDD.n3168 VDD.n3165 0.196152
R14106 VDD.n3619 VDD.n3602 0.196152
R14107 VDD.n3615 VDD.n3606 0.196152
R14108 VDD.n3633 VDD.n3630 0.196152
R14109 VDD.n3647 VDD.n3644 0.196152
R14110 VDD.n3660 VDD.n3657 0.196152
R14111 VDD.n3673 VDD.n3670 0.196152
R14112 VDD.n3686 VDD.n3683 0.196152
R14113 VDD.n3699 VDD.n3696 0.196152
R14114 VDD.n3712 VDD.n3709 0.196152
R14115 VDD.n3726 VDD.n3723 0.196152
R14116 VDD.n3739 VDD.n3736 0.196152
R14117 VDD.n3752 VDD.n3749 0.196152
R14118 VDD.n3765 VDD.n3762 0.196152
R14119 VDD.n3778 VDD.n3775 0.196152
R14120 VDD.n3579 VDD.n3576 0.196152
R14121 VDD.n3565 VDD.n3562 0.196152
R14122 VDD.n3551 VDD.n3548 0.196152
R14123 VDD.n3537 VDD.n3534 0.196152
R14124 VDD.n3523 VDD.n3520 0.196152
R14125 VDD.n3509 VDD.n3506 0.196152
R14126 VDD.n3494 VDD.n3491 0.196152
R14127 VDD.n3479 VDD.n3462 0.196152
R14128 VDD.n3475 VDD.n3466 0.196152
R14129 VDD.n16 VDD.n7 0.196152
R14130 VDD.n16 VDD.n15 0.196152
R14131 VDD.n335 VDD.n326 0.196152
R14132 VDD.n335 VDD.n334 0.196152
R14133 VDD.n545 VDD.n528 0.196152
R14134 VDD.n536 VDD.n527 0.196152
R14135 VDD.n561 VDD.n555 0.196152
R14136 VDD.n794 VDD.n788 0.196152
R14137 VDD.n807 VDD.n801 0.196152
R14138 VDD.n820 VDD.n814 0.196152
R14139 VDD.n833 VDD.n827 0.196152
R14140 VDD.n777 VDD.n771 0.196152
R14141 VDD.n763 VDD.n757 0.196152
R14142 VDD.n749 VDD.n743 0.196152
R14143 VDD.n517 VDD.n511 0.196152
R14144 VDD.n2574 VDD.n2568 0.196152
R14145 VDD.n2378 VDD.n2377 0.196152
R14146 VDD.n2377 VDD.n2173 0.196152
R14147 VDD.n2370 VDD.n2173 0.196152
R14148 VDD.n2370 VDD.n2369 0.196152
R14149 VDD.n2369 VDD.n2177 0.196152
R14150 VDD.n2181 VDD.n2177 0.196152
R14151 VDD.n2360 VDD.n2181 0.196152
R14152 VDD.n2360 VDD.n2359 0.196152
R14153 VDD.n2526 VDD.n2525 0.196152
R14154 VDD.n2525 VDD.n1220 0.196152
R14155 VDD.n1249 VDD.n1220 0.196152
R14156 VDD.n1256 VDD.n1249 0.196152
R14157 VDD.n1257 VDD.n1256 0.196152
R14158 VDD.n2503 VDD.n1257 0.196152
R14159 VDD.n2503 VDD.n2502 0.196152
R14160 VDD.n2502 VDD.n1258 0.196152
R14161 VDD.n2196 VDD.n1258 0.196152
R14162 VDD.n2196 VDD.n2193 0.196152
R14163 VDD.n2203 VDD.n2193 0.196152
R14164 VDD.n1850 VDD.n1538 0.196152
R14165 VDD.n1851 VDD.n1850 0.196152
R14166 VDD.n1859 VDD.n1851 0.196152
R14167 VDD.n1859 VDD.n1858 0.196152
R14168 VDD.n1858 VDD.n1852 0.196152
R14169 VDD.n1852 VDD.n1489 0.196152
R14170 VDD.n1918 VDD.n1489 0.196152
R14171 VDD.n1919 VDD.n1918 0.196152
R14172 VDD.n1927 VDD.n1919 0.196152
R14173 VDD.n1927 VDD.n1926 0.196152
R14174 VDD.n1926 VDD.n1920 0.196152
R14175 VDD.n1738 VDD.n1737 0.196152
R14176 VDD.n1737 VDD.n1711 0.196152
R14177 VDD.n1730 VDD.n1711 0.196152
R14178 VDD.n1730 VDD.n1729 0.196152
R14179 VDD.n1729 VDD.n1713 0.196152
R14180 VDD.n1722 VDD.n1713 0.196152
R14181 VDD.n1722 VDD.n1721 0.196152
R14182 VDD.n1721 VDD.n1717 0.196152
R14183 VDD.n604 VDD.n587 0.196152
R14184 VDD.n601 VDD.n600 0.196152
R14185 VDD.n600 VDD.n591 0.196152
R14186 VDD.n618 VDD.n615 0.196152
R14187 VDD.n692 VDD.n689 0.196152
R14188 VDD.n705 VDD.n702 0.196152
R14189 VDD.n718 VDD.n715 0.196152
R14190 VDD.n731 VDD.n728 0.196152
R14191 VDD.n675 VDD.n672 0.196152
R14192 VDD.n661 VDD.n658 0.196152
R14193 VDD.n647 VDD.n644 0.196152
R14194 VDD.n633 VDD.n630 0.196152
R14195 VDD.n574 VDD.n571 0.196152
R14196 VDD.n1025 VDD.n1008 0.196152
R14197 VDD.n1021 VDD.n1012 0.196152
R14198 VDD.n1039 VDD.n1036 0.196152
R14199 VDD.n1053 VDD.n1050 0.196152
R14200 VDD.n1066 VDD.n1063 0.196152
R14201 VDD.n1079 VDD.n1076 0.196152
R14202 VDD.n1092 VDD.n1089 0.196152
R14203 VDD.n1105 VDD.n1102 0.196152
R14204 VDD.n1118 VDD.n1115 0.196152
R14205 VDD.n1132 VDD.n1129 0.196152
R14206 VDD.n1145 VDD.n1142 0.196152
R14207 VDD.n1158 VDD.n1155 0.196152
R14208 VDD.n1171 VDD.n1168 0.196152
R14209 VDD.n1184 VDD.n1181 0.196152
R14210 VDD.n985 VDD.n982 0.196152
R14211 VDD.n971 VDD.n968 0.196152
R14212 VDD.n957 VDD.n954 0.196152
R14213 VDD.n943 VDD.n940 0.196152
R14214 VDD.n929 VDD.n926 0.196152
R14215 VDD.n915 VDD.n912 0.196152
R14216 VDD.n900 VDD.n897 0.196152
R14217 VDD.n885 VDD.n868 0.196152
R14218 VDD.n881 VDD.n872 0.196152
R14219 VDD.n5579 VDD.n5570 0.196152
R14220 VDD.n5579 VDD.n5578 0.196152
R14221 VDD.n5898 VDD.n5889 0.196152
R14222 VDD.n5898 VDD.n5897 0.196152
R14223 VDD.n6108 VDD.n6091 0.196152
R14224 VDD.n6099 VDD.n6090 0.196152
R14225 VDD.n6124 VDD.n6118 0.196152
R14226 VDD.n6357 VDD.n6351 0.196152
R14227 VDD.n6370 VDD.n6364 0.196152
R14228 VDD.n6383 VDD.n6377 0.196152
R14229 VDD.n6396 VDD.n6390 0.196152
R14230 VDD.n6340 VDD.n6334 0.196152
R14231 VDD.n6326 VDD.n6320 0.196152
R14232 VDD.n6312 VDD.n6306 0.196152
R14233 VDD.n6080 VDD.n6074 0.196152
R14234 VDD.n8137 VDD.n8131 0.196152
R14235 VDD.n7941 VDD.n7940 0.196152
R14236 VDD.n7940 VDD.n7736 0.196152
R14237 VDD.n7933 VDD.n7736 0.196152
R14238 VDD.n7933 VDD.n7932 0.196152
R14239 VDD.n7932 VDD.n7740 0.196152
R14240 VDD.n7744 VDD.n7740 0.196152
R14241 VDD.n7923 VDD.n7744 0.196152
R14242 VDD.n7923 VDD.n7922 0.196152
R14243 VDD.n8089 VDD.n8088 0.196152
R14244 VDD.n8088 VDD.n6783 0.196152
R14245 VDD.n6812 VDD.n6783 0.196152
R14246 VDD.n6819 VDD.n6812 0.196152
R14247 VDD.n6820 VDD.n6819 0.196152
R14248 VDD.n8066 VDD.n6820 0.196152
R14249 VDD.n8066 VDD.n8065 0.196152
R14250 VDD.n8065 VDD.n6821 0.196152
R14251 VDD.n7759 VDD.n6821 0.196152
R14252 VDD.n7759 VDD.n7756 0.196152
R14253 VDD.n7766 VDD.n7756 0.196152
R14254 VDD.n7413 VDD.n7101 0.196152
R14255 VDD.n7414 VDD.n7413 0.196152
R14256 VDD.n7422 VDD.n7414 0.196152
R14257 VDD.n7422 VDD.n7421 0.196152
R14258 VDD.n7421 VDD.n7415 0.196152
R14259 VDD.n7415 VDD.n7052 0.196152
R14260 VDD.n7481 VDD.n7052 0.196152
R14261 VDD.n7482 VDD.n7481 0.196152
R14262 VDD.n7490 VDD.n7482 0.196152
R14263 VDD.n7490 VDD.n7489 0.196152
R14264 VDD.n7489 VDD.n7483 0.196152
R14265 VDD.n7301 VDD.n7300 0.196152
R14266 VDD.n7300 VDD.n7274 0.196152
R14267 VDD.n7293 VDD.n7274 0.196152
R14268 VDD.n7293 VDD.n7292 0.196152
R14269 VDD.n7292 VDD.n7276 0.196152
R14270 VDD.n7285 VDD.n7276 0.196152
R14271 VDD.n7285 VDD.n7284 0.196152
R14272 VDD.n7284 VDD.n7280 0.196152
R14273 VDD.n6167 VDD.n6150 0.196152
R14274 VDD.n6164 VDD.n6163 0.196152
R14275 VDD.n6163 VDD.n6154 0.196152
R14276 VDD.n6181 VDD.n6178 0.196152
R14277 VDD.n6255 VDD.n6252 0.196152
R14278 VDD.n6268 VDD.n6265 0.196152
R14279 VDD.n6281 VDD.n6278 0.196152
R14280 VDD.n6294 VDD.n6291 0.196152
R14281 VDD.n6238 VDD.n6235 0.196152
R14282 VDD.n6224 VDD.n6221 0.196152
R14283 VDD.n6210 VDD.n6207 0.196152
R14284 VDD.n6196 VDD.n6193 0.196152
R14285 VDD.n6137 VDD.n6134 0.196152
R14286 VDD.n6588 VDD.n6571 0.196152
R14287 VDD.n6584 VDD.n6575 0.196152
R14288 VDD.n6602 VDD.n6599 0.196152
R14289 VDD.n6616 VDD.n6613 0.196152
R14290 VDD.n6629 VDD.n6626 0.196152
R14291 VDD.n6642 VDD.n6639 0.196152
R14292 VDD.n6655 VDD.n6652 0.196152
R14293 VDD.n6668 VDD.n6665 0.196152
R14294 VDD.n6681 VDD.n6678 0.196152
R14295 VDD.n6695 VDD.n6692 0.196152
R14296 VDD.n6708 VDD.n6705 0.196152
R14297 VDD.n6721 VDD.n6718 0.196152
R14298 VDD.n6734 VDD.n6731 0.196152
R14299 VDD.n6747 VDD.n6744 0.196152
R14300 VDD.n6548 VDD.n6545 0.196152
R14301 VDD.n6534 VDD.n6531 0.196152
R14302 VDD.n6520 VDD.n6517 0.196152
R14303 VDD.n6506 VDD.n6503 0.196152
R14304 VDD.n6492 VDD.n6489 0.196152
R14305 VDD.n6478 VDD.n6475 0.196152
R14306 VDD.n6463 VDD.n6460 0.196152
R14307 VDD.n6448 VDD.n6431 0.196152
R14308 VDD.n6444 VDD.n6435 0.196152
R14309 VDD.n2916 VDD.n2619 0.193827
R14310 VDD.n322 VDD.n25 0.193827
R14311 VDD.n5885 VDD.n5588 0.193827
R14312 VDD.n8150 VDD.n5181 0.189561
R14313 VDD.n8145 VDD.n5178 0.189561
R14314 VDD.n8154 VDD.n8153 0.189561
R14315 VDD.n8156 VDD.n2582 0.189561
R14316 VDD.n2596 VDD.n2588 0.189561
R14317 VDD.n5176 VDD.n2598 0.189561
R14318 VDD.n3205 VDD.n3181 0.18951
R14319 VDD.n3218 VDD.n3209 0.18951
R14320 VDD.n3292 VDD.n3283 0.18951
R14321 VDD.n3305 VDD.n3296 0.18951
R14322 VDD.n3318 VDD.n3309 0.18951
R14323 VDD.n3331 VDD.n3322 0.18951
R14324 VDD.n3275 VDD.n3266 0.18951
R14325 VDD.n3261 VDD.n3252 0.18951
R14326 VDD.n3247 VDD.n3238 0.18951
R14327 VDD.n3233 VDD.n3224 0.18951
R14328 VDD.n3174 VDD.n3165 0.18951
R14329 VDD.n3626 VDD.n3602 0.18951
R14330 VDD.n3639 VDD.n3630 0.18951
R14331 VDD.n3653 VDD.n3644 0.18951
R14332 VDD.n3666 VDD.n3657 0.18951
R14333 VDD.n3679 VDD.n3670 0.18951
R14334 VDD.n3692 VDD.n3683 0.18951
R14335 VDD.n3705 VDD.n3696 0.18951
R14336 VDD.n3718 VDD.n3709 0.18951
R14337 VDD.n3732 VDD.n3723 0.18951
R14338 VDD.n3745 VDD.n3736 0.18951
R14339 VDD.n3758 VDD.n3749 0.18951
R14340 VDD.n3771 VDD.n3762 0.18951
R14341 VDD.n3784 VDD.n3775 0.18951
R14342 VDD.n3585 VDD.n3576 0.18951
R14343 VDD.n3571 VDD.n3562 0.18951
R14344 VDD.n3557 VDD.n3548 0.18951
R14345 VDD.n3543 VDD.n3534 0.18951
R14346 VDD.n3529 VDD.n3520 0.18951
R14347 VDD.n3515 VDD.n3506 0.18951
R14348 VDD.n3500 VDD.n3491 0.18951
R14349 VDD.n3486 VDD.n3462 0.18951
R14350 VDD.n611 VDD.n587 0.18951
R14351 VDD.n624 VDD.n615 0.18951
R14352 VDD.n698 VDD.n689 0.18951
R14353 VDD.n711 VDD.n702 0.18951
R14354 VDD.n724 VDD.n715 0.18951
R14355 VDD.n737 VDD.n728 0.18951
R14356 VDD.n681 VDD.n672 0.18951
R14357 VDD.n667 VDD.n658 0.18951
R14358 VDD.n653 VDD.n644 0.18951
R14359 VDD.n639 VDD.n630 0.18951
R14360 VDD.n580 VDD.n571 0.18951
R14361 VDD.n1032 VDD.n1008 0.18951
R14362 VDD.n1045 VDD.n1036 0.18951
R14363 VDD.n1059 VDD.n1050 0.18951
R14364 VDD.n1072 VDD.n1063 0.18951
R14365 VDD.n1085 VDD.n1076 0.18951
R14366 VDD.n1098 VDD.n1089 0.18951
R14367 VDD.n1111 VDD.n1102 0.18951
R14368 VDD.n1124 VDD.n1115 0.18951
R14369 VDD.n1138 VDD.n1129 0.18951
R14370 VDD.n1151 VDD.n1142 0.18951
R14371 VDD.n1164 VDD.n1155 0.18951
R14372 VDD.n1177 VDD.n1168 0.18951
R14373 VDD.n1190 VDD.n1181 0.18951
R14374 VDD.n991 VDD.n982 0.18951
R14375 VDD.n977 VDD.n968 0.18951
R14376 VDD.n963 VDD.n954 0.18951
R14377 VDD.n949 VDD.n940 0.18951
R14378 VDD.n935 VDD.n926 0.18951
R14379 VDD.n921 VDD.n912 0.18951
R14380 VDD.n906 VDD.n897 0.18951
R14381 VDD.n892 VDD.n868 0.18951
R14382 VDD.n6174 VDD.n6150 0.18951
R14383 VDD.n6187 VDD.n6178 0.18951
R14384 VDD.n6261 VDD.n6252 0.18951
R14385 VDD.n6274 VDD.n6265 0.18951
R14386 VDD.n6287 VDD.n6278 0.18951
R14387 VDD.n6300 VDD.n6291 0.18951
R14388 VDD.n6244 VDD.n6235 0.18951
R14389 VDD.n6230 VDD.n6221 0.18951
R14390 VDD.n6216 VDD.n6207 0.18951
R14391 VDD.n6202 VDD.n6193 0.18951
R14392 VDD.n6143 VDD.n6134 0.18951
R14393 VDD.n6595 VDD.n6571 0.18951
R14394 VDD.n6608 VDD.n6599 0.18951
R14395 VDD.n6622 VDD.n6613 0.18951
R14396 VDD.n6635 VDD.n6626 0.18951
R14397 VDD.n6648 VDD.n6639 0.18951
R14398 VDD.n6661 VDD.n6652 0.18951
R14399 VDD.n6674 VDD.n6665 0.18951
R14400 VDD.n6687 VDD.n6678 0.18951
R14401 VDD.n6701 VDD.n6692 0.18951
R14402 VDD.n6714 VDD.n6705 0.18951
R14403 VDD.n6727 VDD.n6718 0.18951
R14404 VDD.n6740 VDD.n6731 0.18951
R14405 VDD.n6753 VDD.n6744 0.18951
R14406 VDD.n6554 VDD.n6545 0.18951
R14407 VDD.n6540 VDD.n6531 0.18951
R14408 VDD.n6526 VDD.n6517 0.18951
R14409 VDD.n6512 VDD.n6503 0.18951
R14410 VDD.n6498 VDD.n6489 0.18951
R14411 VDD.n6484 VDD.n6475 0.18951
R14412 VDD.n6469 VDD.n6460 0.18951
R14413 VDD.n6455 VDD.n6431 0.18951
R14414 VDD.n5307 VDD.n5306 0.188144
R14415 VDD.n8149 VDD.n8148 0.188107
R14416 VDD.n5184 VDD.n5182 0.188107
R14417 VDD.n8151 VDD.n5179 0.188107
R14418 VDD.n5185 VDD.n5182 0.188107
R14419 VDD.n8157 VDD.n2 0.188107
R14420 VDD.n2584 VDD.n0 0.188107
R14421 VDD.n8155 VDD.n2583 0.188107
R14422 VDD.n4 VDD.n0 0.188107
R14423 VDD.n2595 VDD.n2593 0.188107
R14424 VDD.n2592 VDD.n2591 0.188107
R14425 VDD.n2597 VDD.n2594 0.188107
R14426 VDD.n2592 VDD.n2590 0.188107
R14427 VDD.n5305 VDD.n5186 0.187918
R14428 VDD.n3146 VDD.n3122 0.184196
R14429 VDD.n552 VDD.n528 0.184196
R14430 VDD.n6115 VDD.n6091 0.184196
R14431 VDD.n2617 VDD.n2601 0.180011
R14432 VDD.n2936 VDD.n2920 0.180011
R14433 VDD.n23 VDD.n7 0.180011
R14434 VDD.n342 VDD.n326 0.180011
R14435 VDD.n5586 VDD.n5570 0.180011
R14436 VDD.n5905 VDD.n5889 0.180011
R14437 VDD.n3130 VDD.n3129 0.176225
R14438 VDD.n3155 VDD.n3154 0.176225
R14439 VDD.n3388 VDD.n3387 0.176225
R14440 VDD.n3401 VDD.n3400 0.176225
R14441 VDD.n3414 VDD.n3413 0.176225
R14442 VDD.n3427 VDD.n3426 0.176225
R14443 VDD.n3371 VDD.n3370 0.176225
R14444 VDD.n3357 VDD.n3356 0.176225
R14445 VDD.n3343 VDD.n3342 0.176225
R14446 VDD.n3111 VDD.n3110 0.176225
R14447 VDD.n5168 VDD.n5167 0.176225
R14448 VDD.n536 VDD.n535 0.176225
R14449 VDD.n561 VDD.n560 0.176225
R14450 VDD.n794 VDD.n793 0.176225
R14451 VDD.n807 VDD.n806 0.176225
R14452 VDD.n820 VDD.n819 0.176225
R14453 VDD.n833 VDD.n832 0.176225
R14454 VDD.n777 VDD.n776 0.176225
R14455 VDD.n763 VDD.n762 0.176225
R14456 VDD.n749 VDD.n748 0.176225
R14457 VDD.n517 VDD.n516 0.176225
R14458 VDD.n2574 VDD.n2573 0.176225
R14459 VDD.n6099 VDD.n6098 0.176225
R14460 VDD.n6124 VDD.n6123 0.176225
R14461 VDD.n6357 VDD.n6356 0.176225
R14462 VDD.n6370 VDD.n6369 0.176225
R14463 VDD.n6383 VDD.n6382 0.176225
R14464 VDD.n6396 VDD.n6395 0.176225
R14465 VDD.n6340 VDD.n6339 0.176225
R14466 VDD.n6326 VDD.n6325 0.176225
R14467 VDD.n6312 VDD.n6311 0.176225
R14468 VDD.n6080 VDD.n6079 0.176225
R14469 VDD.n8137 VDD.n8136 0.176225
R14470 VDD.n3616 VDD.n3615 0.157626
R14471 VDD.n3476 VDD.n3475 0.157626
R14472 VDD.n1022 VDD.n1021 0.157626
R14473 VDD.n882 VDD.n881 0.157626
R14474 VDD.n6585 VDD.n6584 0.157626
R14475 VDD.n6445 VDD.n6444 0.157626
R14476 VDD.n2911 VDD.n2743 0.150564
R14477 VDD.n2825 VDD.n2796 0.150564
R14478 VDD.n317 VDD.n149 0.150564
R14479 VDD.n231 VDD.n202 0.150564
R14480 VDD.n5880 VDD.n5712 0.150564
R14481 VDD.n5794 VDD.n5765 0.150564
R14482 VDD.n3619 VDD.n3600 0.13335
R14483 VDD.n3633 VDD.n3599 0.13335
R14484 VDD.n3647 VDD.n3598 0.13335
R14485 VDD.n3660 VDD.n3597 0.13335
R14486 VDD.n3673 VDD.n3596 0.13335
R14487 VDD.n3686 VDD.n3595 0.13335
R14488 VDD.n3699 VDD.n3594 0.13335
R14489 VDD.n3712 VDD.n3593 0.13335
R14490 VDD.n3726 VDD.n3592 0.13335
R14491 VDD.n3739 VDD.n3591 0.13335
R14492 VDD.n3752 VDD.n3590 0.13335
R14493 VDD.n3765 VDD.n3589 0.13335
R14494 VDD.n3778 VDD.n3588 0.13335
R14495 VDD.n3579 VDD.n3574 0.13335
R14496 VDD.n3565 VDD.n3560 0.13335
R14497 VDD.n3551 VDD.n3546 0.13335
R14498 VDD.n3537 VDD.n3532 0.13335
R14499 VDD.n3523 VDD.n3518 0.13335
R14500 VDD.n3509 VDD.n3504 0.13335
R14501 VDD.n3494 VDD.n3489 0.13335
R14502 VDD.n3479 VDD.n3460 0.13335
R14503 VDD.n1025 VDD.n1006 0.13335
R14504 VDD.n1039 VDD.n1005 0.13335
R14505 VDD.n1053 VDD.n1004 0.13335
R14506 VDD.n1066 VDD.n1003 0.13335
R14507 VDD.n1079 VDD.n1002 0.13335
R14508 VDD.n1092 VDD.n1001 0.13335
R14509 VDD.n1105 VDD.n1000 0.13335
R14510 VDD.n1118 VDD.n999 0.13335
R14511 VDD.n1132 VDD.n998 0.13335
R14512 VDD.n1145 VDD.n997 0.13335
R14513 VDD.n1158 VDD.n996 0.13335
R14514 VDD.n1171 VDD.n995 0.13335
R14515 VDD.n1184 VDD.n994 0.13335
R14516 VDD.n985 VDD.n980 0.13335
R14517 VDD.n971 VDD.n966 0.13335
R14518 VDD.n957 VDD.n952 0.13335
R14519 VDD.n943 VDD.n938 0.13335
R14520 VDD.n929 VDD.n924 0.13335
R14521 VDD.n915 VDD.n910 0.13335
R14522 VDD.n900 VDD.n895 0.13335
R14523 VDD.n885 VDD.n866 0.13335
R14524 VDD.n6588 VDD.n6569 0.13335
R14525 VDD.n6602 VDD.n6568 0.13335
R14526 VDD.n6616 VDD.n6567 0.13335
R14527 VDD.n6629 VDD.n6566 0.13335
R14528 VDD.n6642 VDD.n6565 0.13335
R14529 VDD.n6655 VDD.n6564 0.13335
R14530 VDD.n6668 VDD.n6563 0.13335
R14531 VDD.n6681 VDD.n6562 0.13335
R14532 VDD.n6695 VDD.n6561 0.13335
R14533 VDD.n6708 VDD.n6560 0.13335
R14534 VDD.n6721 VDD.n6559 0.13335
R14535 VDD.n6734 VDD.n6558 0.13335
R14536 VDD.n6747 VDD.n6557 0.13335
R14537 VDD.n6548 VDD.n6543 0.13335
R14538 VDD.n6534 VDD.n6529 0.13335
R14539 VDD.n6520 VDD.n6515 0.13335
R14540 VDD.n6506 VDD.n6501 0.13335
R14541 VDD.n6492 VDD.n6487 0.13335
R14542 VDD.n6478 VDD.n6473 0.13335
R14543 VDD.n6463 VDD.n6458 0.13335
R14544 VDD.n6448 VDD.n6429 0.13335
R14545 VDD.n5120 VDD.n3791 0.127764
R14546 VDD.n2526 VDD.n1197 0.127764
R14547 VDD.n8089 VDD.n6760 0.127764
R14548 VDD.n4311 VDD.n4071 0.126643
R14549 VDD.n1717 VDD.n1477 0.126643
R14550 VDD.n7280 VDD.n7040 0.126643
R14551 VDD.n5460 VDD.n5459 0.120292
R14552 VDD.n5459 VDD.n5458 0.120292
R14553 VDD.n5455 VDD.n5454 0.120292
R14554 VDD.n5454 VDD.n5453 0.120292
R14555 VDD.n5453 VDD.n5447 0.120292
R14556 VDD.n5449 VDD.n5447 0.120292
R14557 VDD.n5495 VDD.n5485 0.120292
R14558 VDD.n5496 VDD.n5495 0.120292
R14559 VDD.n5497 VDD.n5496 0.120292
R14560 VDD.n5497 VDD.n5482 0.120292
R14561 VDD.n5502 VDD.n5482 0.120292
R14562 VDD.n5509 VDD.n5508 0.120292
R14563 VDD.n5508 VDD.n5503 0.120292
R14564 VDD.n5503 VDD.n5476 0.120292
R14565 VDD.n5516 VDD.n5476 0.120292
R14566 VDD.n5517 VDD.n5516 0.120292
R14567 VDD.n5518 VDD.n5517 0.120292
R14568 VDD.n5518 VDD.n5473 0.120292
R14569 VDD.n5525 VDD.n5473 0.120292
R14570 VDD.n5533 VDD.n5532 0.120292
R14571 VDD.n5532 VDD.n5527 0.120292
R14572 VDD.n5527 VDD.n5468 0.120292
R14573 VDD.n5540 VDD.n5468 0.120292
R14574 VDD.n5541 VDD.n5540 0.120292
R14575 VDD.n5541 VDD.n5465 0.120292
R14576 VDD.n5547 VDD.n5465 0.120292
R14577 VDD.n5556 VDD.n5555 0.120292
R14578 VDD.n5555 VDD.n5550 0.120292
R14579 VDD.n5550 VDD.n5549 0.120292
R14580 VDD.n5435 VDD.n5434 0.120292
R14581 VDD.n5434 VDD.n5316 0.120292
R14582 VDD.n5429 VDD.n5426 0.120292
R14583 VDD.n5429 VDD.n5428 0.120292
R14584 VDD.n5357 VDD.n5347 0.120292
R14585 VDD.n5357 VDD.n5356 0.120292
R14586 VDD.n5356 VDD.n5348 0.120292
R14587 VDD.n5351 VDD.n5348 0.120292
R14588 VDD.n5351 VDD.n5350 0.120292
R14589 VDD.n5365 VDD.n5364 0.120292
R14590 VDD.n5366 VDD.n5365 0.120292
R14591 VDD.n5366 VDD.n5336 0.120292
R14592 VDD.n5373 VDD.n5336 0.120292
R14593 VDD.n5374 VDD.n5373 0.120292
R14594 VDD.n5379 VDD.n5374 0.120292
R14595 VDD.n5379 VDD.n5378 0.120292
R14596 VDD.n5378 VDD.n5375 0.120292
R14597 VDD.n5386 VDD.n5331 0.120292
R14598 VDD.n5387 VDD.n5386 0.120292
R14599 VDD.n5388 VDD.n5387 0.120292
R14600 VDD.n5388 VDD.n5328 0.120292
R14601 VDD.n5394 VDD.n5393 0.120292
R14602 VDD.n5401 VDD.n5394 0.120292
R14603 VDD.n5401 VDD.n5400 0.120292
R14604 VDD.n5400 VDD.n5395 0.120292
R14605 VDD.n5395 VDD.n5323 0.120292
R14606 VDD.n5408 VDD.n5323 0.120292
R14607 VDD.n5409 VDD.n5408 0.120292
R14608 VDD.n5409 VDD.n5320 0.120292
R14609 VDD.n5415 VDD.n5414 0.120292
R14610 VDD.n5420 VDD.n5415 0.120292
R14611 VDD.n5420 VDD.n5419 0.120292
R14612 VDD.n5419 VDD.n5416 0.120292
R14613 VDD.n4972 VDD.n4766 0.117055
R14614 VDD.n2378 VDD.n2172 0.117055
R14615 VDD.n7941 VDD.n7735 0.117055
R14616 VDD.n5175 VDD.n3102 0.11095
R14617 VDD.n2581 VDD.n508 0.11095
R14618 VDD.n8144 VDD.n6071 0.11095
R14619 VDD.n2912 VDD.n2911 0.107565
R14620 VDD.n2796 VDD.n2793 0.107565
R14621 VDD.n318 VDD.n317 0.107565
R14622 VDD.n202 VDD.n199 0.107565
R14623 VDD.n5881 VDD.n5880 0.107565
R14624 VDD.n5765 VDD.n5762 0.107565
R14625 VDD.n5533 VDD 0.0968542
R14626 VDD.n5556 VDD 0.0968542
R14627 VDD.n8145 VDD.n8144 0.0937167
R14628 VDD.n5176 VDD.n5175 0.09356
R14629 VDD.n2582 VDD.n2581 0.09356
R14630 VDD.n3147 VDD.n3121 0.0790024
R14631 VDD.n3160 VDD.n3149 0.0790024
R14632 VDD.n3393 VDD.n3382 0.0790024
R14633 VDD.n3406 VDD.n3395 0.0790024
R14634 VDD.n3419 VDD.n3408 0.0790024
R14635 VDD.n3432 VDD.n3421 0.0790024
R14636 VDD.n3376 VDD.n3365 0.0790024
R14637 VDD.n3362 VDD.n3351 0.0790024
R14638 VDD.n3348 VDD.n3337 0.0790024
R14639 VDD.n3116 VDD.n3105 0.0790024
R14640 VDD.n5173 VDD.n5162 0.0790024
R14641 VDD.n553 VDD.n527 0.0790024
R14642 VDD.n566 VDD.n555 0.0790024
R14643 VDD.n799 VDD.n788 0.0790024
R14644 VDD.n812 VDD.n801 0.0790024
R14645 VDD.n825 VDD.n814 0.0790024
R14646 VDD.n838 VDD.n827 0.0790024
R14647 VDD.n782 VDD.n771 0.0790024
R14648 VDD.n768 VDD.n757 0.0790024
R14649 VDD.n754 VDD.n743 0.0790024
R14650 VDD.n522 VDD.n511 0.0790024
R14651 VDD.n2579 VDD.n2568 0.0790024
R14652 VDD.n6116 VDD.n6090 0.0790024
R14653 VDD.n6129 VDD.n6118 0.0790024
R14654 VDD.n6362 VDD.n6351 0.0790024
R14655 VDD.n6375 VDD.n6364 0.0790024
R14656 VDD.n6388 VDD.n6377 0.0790024
R14657 VDD.n6401 VDD.n6390 0.0790024
R14658 VDD.n6345 VDD.n6334 0.0790024
R14659 VDD.n6331 VDD.n6320 0.0790024
R14660 VDD.n6317 VDD.n6306 0.0790024
R14661 VDD.n6085 VDD.n6074 0.0790024
R14662 VDD.n8142 VDD.n8131 0.0790024
R14663 VDD.n4514 VDD.n3457 0.0664514
R14664 VDD.n1920 VDD.n863 0.0664514
R14665 VDD.n7483 VDD.n6426 0.0664514
R14666 VDD.n5246 VDD.n5188 0.063
R14667 VDD.n5246 VDD.n5245 0.063
R14668 VDD.n5216 VDD.n5187 0.063
R14669 VDD.n5196 VDD.n5187 0.063
R14670 VDD.n5439 VDD.n5310 0.0624835
R14671 VDD.n5197 VDD.n5188 0.0622084
R14672 VDD.n5460 VDD.n5441 0.0603958
R14673 VDD.n5458 VDD 0.0603958
R14674 VDD.n5455 VDD 0.0603958
R14675 VDD.n5509 VDD 0.0603958
R14676 VDD.n5526 VDD 0.0603958
R14677 VDD VDD.n5547 0.0603958
R14678 VDD.n5548 VDD 0.0603958
R14679 VDD.n5435 VDD.n5311 0.0603958
R14680 VDD.n5426 VDD 0.0603958
R14681 VDD.n5364 VDD 0.0603958
R14682 VDD VDD.n5331 0.0603958
R14683 VDD.n5393 VDD 0.0603958
R14684 VDD.n5414 VDD 0.0603958
R14685 VDD.n3198 VDD.n3179 0.0518285
R14686 VDD.n3195 VDD.n3179 0.0518285
R14687 VDD.n3212 VDD.n3178 0.0518285
R14688 VDD.n3286 VDD.n3281 0.0518285
R14689 VDD.n3299 VDD.n3280 0.0518285
R14690 VDD.n3312 VDD.n3279 0.0518285
R14691 VDD.n3325 VDD.n3278 0.0518285
R14692 VDD.n3269 VDD.n3264 0.0518285
R14693 VDD.n3255 VDD.n3250 0.0518285
R14694 VDD.n3241 VDD.n3236 0.0518285
R14695 VDD.n3227 VDD.n3222 0.0518285
R14696 VDD.n3168 VDD.n3163 0.0518285
R14697 VDD.n604 VDD.n585 0.0518285
R14698 VDD.n601 VDD.n585 0.0518285
R14699 VDD.n618 VDD.n584 0.0518285
R14700 VDD.n692 VDD.n687 0.0518285
R14701 VDD.n705 VDD.n686 0.0518285
R14702 VDD.n718 VDD.n685 0.0518285
R14703 VDD.n731 VDD.n684 0.0518285
R14704 VDD.n675 VDD.n670 0.0518285
R14705 VDD.n661 VDD.n656 0.0518285
R14706 VDD.n647 VDD.n642 0.0518285
R14707 VDD.n633 VDD.n628 0.0518285
R14708 VDD.n574 VDD.n569 0.0518285
R14709 VDD.n6167 VDD.n6148 0.0518285
R14710 VDD.n6164 VDD.n6148 0.0518285
R14711 VDD.n6181 VDD.n6147 0.0518285
R14712 VDD.n6255 VDD.n6250 0.0518285
R14713 VDD.n6268 VDD.n6249 0.0518285
R14714 VDD.n6281 VDD.n6248 0.0518285
R14715 VDD.n6294 VDD.n6247 0.0518285
R14716 VDD.n6238 VDD.n6233 0.0518285
R14717 VDD.n6224 VDD.n6219 0.0518285
R14718 VDD.n6210 VDD.n6205 0.0518285
R14719 VDD.n6196 VDD.n6191 0.0518285
R14720 VDD.n6137 VDD.n6132 0.0518285
R14721 VDD.n3249 VDD.n3235 0.0506333
R14722 VDD.n3277 VDD.n3263 0.0506333
R14723 VDD.n3320 VDD.n3307 0.0506333
R14724 VDD.n3307 VDD.n3294 0.0506333
R14725 VDD.n3220 VDD.n3207 0.0506333
R14726 VDD.n3349 VDD.n3117 0.0506333
R14727 VDD.n3363 VDD.n3349 0.0506333
R14728 VDD.n3420 VDD.n3407 0.0506333
R14729 VDD.n3407 VDD.n3394 0.0506333
R14730 VDD.n3161 VDD.n3148 0.0506333
R14731 VDD.n655 VDD.n641 0.0506333
R14732 VDD.n683 VDD.n669 0.0506333
R14733 VDD.n726 VDD.n713 0.0506333
R14734 VDD.n713 VDD.n700 0.0506333
R14735 VDD.n626 VDD.n613 0.0506333
R14736 VDD.n755 VDD.n523 0.0506333
R14737 VDD.n769 VDD.n755 0.0506333
R14738 VDD.n826 VDD.n813 0.0506333
R14739 VDD.n813 VDD.n800 0.0506333
R14740 VDD.n567 VDD.n554 0.0506333
R14741 VDD.n6218 VDD.n6204 0.0506333
R14742 VDD.n6246 VDD.n6232 0.0506333
R14743 VDD.n6289 VDD.n6276 0.0506333
R14744 VDD.n6276 VDD.n6263 0.0506333
R14745 VDD.n6189 VDD.n6176 0.0506333
R14746 VDD.n6318 VDD.n6086 0.0506333
R14747 VDD.n6332 VDD.n6318 0.0506333
R14748 VDD.n6389 VDD.n6376 0.0506333
R14749 VDD.n6376 VDD.n6363 0.0506333
R14750 VDD.n6130 VDD.n6117 0.0506333
R14751 VDD.n3263 VDD.n3249 0.0490667
R14752 VDD.n3333 VDD.n3320 0.0490667
R14753 VDD.n3377 VDD.n3363 0.0490667
R14754 VDD.n3433 VDD.n3420 0.0490667
R14755 VDD.n669 VDD.n655 0.0490667
R14756 VDD.n739 VDD.n726 0.0490667
R14757 VDD.n783 VDD.n769 0.0490667
R14758 VDD.n839 VDD.n826 0.0490667
R14759 VDD.n6232 VDD.n6218 0.0490667
R14760 VDD.n6302 VDD.n6289 0.0490667
R14761 VDD.n6346 VDD.n6332 0.0490667
R14762 VDD.n6402 VDD.n6389 0.0490667
R14763 VDD.n5438 VDD.n5311 0.0480207
R14764 VDD.n5565 VDD.n5440 0.0471667
R14765 VDD.n3531 VDD.n3517 0.0460758
R14766 VDD.n3559 VDD.n3545 0.0460758
R14767 VDD.n3587 VDD.n3573 0.0460758
R14768 VDD.n3773 VDD.n3760 0.0460758
R14769 VDD.n3747 VDD.n3734 0.0460758
R14770 VDD.n3707 VDD.n3694 0.0460758
R14771 VDD.n3694 VDD.n3681 0.0460758
R14772 VDD.n3668 VDD.n3655 0.0460758
R14773 VDD.n3641 VDD.n3628 0.0460758
R14774 VDD.n937 VDD.n923 0.0460758
R14775 VDD.n965 VDD.n951 0.0460758
R14776 VDD.n993 VDD.n979 0.0460758
R14777 VDD.n1179 VDD.n1166 0.0460758
R14778 VDD.n1153 VDD.n1140 0.0460758
R14779 VDD.n1113 VDD.n1100 0.0460758
R14780 VDD.n1100 VDD.n1087 0.0460758
R14781 VDD.n1074 VDD.n1061 0.0460758
R14782 VDD.n1047 VDD.n1034 0.0460758
R14783 VDD.n6500 VDD.n6486 0.0460758
R14784 VDD.n6528 VDD.n6514 0.0460758
R14785 VDD.n6556 VDD.n6542 0.0460758
R14786 VDD.n6742 VDD.n6729 0.0460758
R14787 VDD.n6716 VDD.n6703 0.0460758
R14788 VDD.n6676 VDD.n6663 0.0460758
R14789 VDD.n6663 VDD.n6650 0.0460758
R14790 VDD.n6637 VDD.n6624 0.0460758
R14791 VDD.n6610 VDD.n6597 0.0460758
R14792 VDD.n3502 VDD.n3488 0.0446515
R14793 VDD.n3545 VDD.n3531 0.0446515
R14794 VDD.n3573 VDD.n3559 0.0446515
R14795 VDD.n3786 VDD.n3773 0.0446515
R14796 VDD.n3760 VDD.n3747 0.0446515
R14797 VDD.n3720 VDD.n3707 0.0446515
R14798 VDD.n3681 VDD.n3668 0.0446515
R14799 VDD.n908 VDD.n894 0.0446515
R14800 VDD.n951 VDD.n937 0.0446515
R14801 VDD.n979 VDD.n965 0.0446515
R14802 VDD.n1192 VDD.n1179 0.0446515
R14803 VDD.n1166 VDD.n1153 0.0446515
R14804 VDD.n1126 VDD.n1113 0.0446515
R14805 VDD.n1087 VDD.n1074 0.0446515
R14806 VDD.n6471 VDD.n6457 0.0446515
R14807 VDD.n6514 VDD.n6500 0.0446515
R14808 VDD.n6542 VDD.n6528 0.0446515
R14809 VDD.n6755 VDD.n6742 0.0446515
R14810 VDD.n6729 VDD.n6716 0.0446515
R14811 VDD.n6689 VDD.n6676 0.0446515
R14812 VDD.n6650 VDD.n6637 0.0446515
R14813 VDD.n3206 VDD.n3205 0.0421667
R14814 VDD.n3219 VDD.n3218 0.0421667
R14815 VDD.n3293 VDD.n3292 0.0421667
R14816 VDD.n3306 VDD.n3305 0.0421667
R14817 VDD.n3319 VDD.n3318 0.0421667
R14818 VDD.n3332 VDD.n3331 0.0421667
R14819 VDD.n3276 VDD.n3275 0.0421667
R14820 VDD.n3262 VDD.n3261 0.0421667
R14821 VDD.n3248 VDD.n3247 0.0421667
R14822 VDD.n3234 VDD.n3233 0.0421667
R14823 VDD.n3175 VDD.n3174 0.0421667
R14824 VDD.n3627 VDD.n3626 0.0421667
R14825 VDD.n3640 VDD.n3639 0.0421667
R14826 VDD.n3654 VDD.n3653 0.0421667
R14827 VDD.n3667 VDD.n3666 0.0421667
R14828 VDD.n3680 VDD.n3679 0.0421667
R14829 VDD.n3693 VDD.n3692 0.0421667
R14830 VDD.n3706 VDD.n3705 0.0421667
R14831 VDD.n3719 VDD.n3718 0.0421667
R14832 VDD.n3733 VDD.n3732 0.0421667
R14833 VDD.n3746 VDD.n3745 0.0421667
R14834 VDD.n3759 VDD.n3758 0.0421667
R14835 VDD.n3772 VDD.n3771 0.0421667
R14836 VDD.n3785 VDD.n3784 0.0421667
R14837 VDD.n3586 VDD.n3585 0.0421667
R14838 VDD.n3572 VDD.n3571 0.0421667
R14839 VDD.n3558 VDD.n3557 0.0421667
R14840 VDD.n3544 VDD.n3543 0.0421667
R14841 VDD.n3530 VDD.n3529 0.0421667
R14842 VDD.n3516 VDD.n3515 0.0421667
R14843 VDD.n3501 VDD.n3500 0.0421667
R14844 VDD.n3487 VDD.n3486 0.0421667
R14845 VDD.n612 VDD.n611 0.0421667
R14846 VDD.n625 VDD.n624 0.0421667
R14847 VDD.n699 VDD.n698 0.0421667
R14848 VDD.n712 VDD.n711 0.0421667
R14849 VDD.n725 VDD.n724 0.0421667
R14850 VDD.n738 VDD.n737 0.0421667
R14851 VDD.n682 VDD.n681 0.0421667
R14852 VDD.n668 VDD.n667 0.0421667
R14853 VDD.n654 VDD.n653 0.0421667
R14854 VDD.n640 VDD.n639 0.0421667
R14855 VDD.n581 VDD.n580 0.0421667
R14856 VDD.n1033 VDD.n1032 0.0421667
R14857 VDD.n1046 VDD.n1045 0.0421667
R14858 VDD.n1060 VDD.n1059 0.0421667
R14859 VDD.n1073 VDD.n1072 0.0421667
R14860 VDD.n1086 VDD.n1085 0.0421667
R14861 VDD.n1099 VDD.n1098 0.0421667
R14862 VDD.n1112 VDD.n1111 0.0421667
R14863 VDD.n1125 VDD.n1124 0.0421667
R14864 VDD.n1139 VDD.n1138 0.0421667
R14865 VDD.n1152 VDD.n1151 0.0421667
R14866 VDD.n1165 VDD.n1164 0.0421667
R14867 VDD.n1178 VDD.n1177 0.0421667
R14868 VDD.n1191 VDD.n1190 0.0421667
R14869 VDD.n992 VDD.n991 0.0421667
R14870 VDD.n978 VDD.n977 0.0421667
R14871 VDD.n964 VDD.n963 0.0421667
R14872 VDD.n950 VDD.n949 0.0421667
R14873 VDD.n936 VDD.n935 0.0421667
R14874 VDD.n922 VDD.n921 0.0421667
R14875 VDD.n907 VDD.n906 0.0421667
R14876 VDD.n893 VDD.n892 0.0421667
R14877 VDD.n6175 VDD.n6174 0.0421667
R14878 VDD.n6188 VDD.n6187 0.0421667
R14879 VDD.n6262 VDD.n6261 0.0421667
R14880 VDD.n6275 VDD.n6274 0.0421667
R14881 VDD.n6288 VDD.n6287 0.0421667
R14882 VDD.n6301 VDD.n6300 0.0421667
R14883 VDD.n6245 VDD.n6244 0.0421667
R14884 VDD.n6231 VDD.n6230 0.0421667
R14885 VDD.n6217 VDD.n6216 0.0421667
R14886 VDD.n6203 VDD.n6202 0.0421667
R14887 VDD.n6144 VDD.n6143 0.0421667
R14888 VDD.n6596 VDD.n6595 0.0421667
R14889 VDD.n6609 VDD.n6608 0.0421667
R14890 VDD.n6623 VDD.n6622 0.0421667
R14891 VDD.n6636 VDD.n6635 0.0421667
R14892 VDD.n6649 VDD.n6648 0.0421667
R14893 VDD.n6662 VDD.n6661 0.0421667
R14894 VDD.n6675 VDD.n6674 0.0421667
R14895 VDD.n6688 VDD.n6687 0.0421667
R14896 VDD.n6702 VDD.n6701 0.0421667
R14897 VDD.n6715 VDD.n6714 0.0421667
R14898 VDD.n6728 VDD.n6727 0.0421667
R14899 VDD.n6741 VDD.n6740 0.0421667
R14900 VDD.n6754 VDD.n6753 0.0421667
R14901 VDD.n6555 VDD.n6554 0.0421667
R14902 VDD.n6541 VDD.n6540 0.0421667
R14903 VDD.n6527 VDD.n6526 0.0421667
R14904 VDD.n6513 VDD.n6512 0.0421667
R14905 VDD.n6499 VDD.n6498 0.0421667
R14906 VDD.n6485 VDD.n6484 0.0421667
R14907 VDD.n6470 VDD.n6469 0.0421667
R14908 VDD.n6456 VDD.n6455 0.0421667
R14909 VDD.n2996 VDD.n2995 0.0414091
R14910 VDD.n2621 VDD.n2620 0.0414091
R14911 VDD.n402 VDD.n401 0.0414091
R14912 VDD.n27 VDD.n26 0.0414091
R14913 VDD.n5965 VDD.n5964 0.0414091
R14914 VDD.n5590 VDD.n5589 0.0414091
R14915 VDD.n5564 VDD.n5441 0.0388333
R14916 VDD.n5197 VDD.n5196 0.0384591
R14917 VDD.n5215 VDD.n5200 0.038
R14918 VDD.n5275 VDD.n5260 0.038
R14919 VDD.n2995 VDD.n2941 0.0374318
R14920 VDD.n3100 VDD.n2621 0.0374318
R14921 VDD.n401 VDD.n347 0.0374318
R14922 VDD.n506 VDD.n27 0.0374318
R14923 VDD.n5964 VDD.n5910 0.0374318
R14924 VDD.n6069 VDD.n5590 0.0374318
R14925 VDD.n2618 VDD.n2617 0.03675
R14926 VDD.n2937 VDD.n2936 0.03675
R14927 VDD.n24 VDD.n23 0.03675
R14928 VDD.n343 VDD.n342 0.03675
R14929 VDD.n5587 VDD.n5586 0.03675
R14930 VDD.n5906 VDD.n5905 0.03675
R14931 VDD.n3147 VDD.n3146 0.0366111
R14932 VDD.n553 VDD.n552 0.0366111
R14933 VDD.n6116 VDD.n6115 0.0366111
R14934 VDD.n5549 VDD.n5440 0.0343542
R14935 VDD.n2747 VDD.n2743 0.0299118
R14936 VDD.n2904 VDD.n2903 0.0299118
R14937 VDD.n2754 VDD.n2748 0.0299118
R14938 VDD.n2825 VDD.n2824 0.0299118
R14939 VDD.n2816 VDD.n2797 0.0299118
R14940 VDD.n2834 VDD.n2783 0.0299118
R14941 VDD.n153 VDD.n149 0.0299118
R14942 VDD.n310 VDD.n309 0.0299118
R14943 VDD.n160 VDD.n154 0.0299118
R14944 VDD.n231 VDD.n230 0.0299118
R14945 VDD.n222 VDD.n203 0.0299118
R14946 VDD.n240 VDD.n189 0.0299118
R14947 VDD.n5716 VDD.n5712 0.0299118
R14948 VDD.n5873 VDD.n5872 0.0299118
R14949 VDD.n5723 VDD.n5717 0.0299118
R14950 VDD.n5794 VDD.n5793 0.0299118
R14951 VDD.n5785 VDD.n5766 0.0299118
R14952 VDD.n5803 VDD.n5752 0.0299118
R14953 VDD.n3129 VDD.n3120 0.0282778
R14954 VDD.n3154 VDD.n3119 0.0282778
R14955 VDD.n3387 VDD.n3381 0.0282778
R14956 VDD.n3400 VDD.n3380 0.0282778
R14957 VDD.n3413 VDD.n3379 0.0282778
R14958 VDD.n3426 VDD.n3378 0.0282778
R14959 VDD.n3370 VDD.n3364 0.0282778
R14960 VDD.n3356 VDD.n3350 0.0282778
R14961 VDD.n3342 VDD.n3336 0.0282778
R14962 VDD.n3110 VDD.n3104 0.0282778
R14963 VDD.n5167 VDD.n3103 0.0282778
R14964 VDD.n535 VDD.n526 0.0282778
R14965 VDD.n560 VDD.n525 0.0282778
R14966 VDD.n793 VDD.n787 0.0282778
R14967 VDD.n806 VDD.n786 0.0282778
R14968 VDD.n819 VDD.n785 0.0282778
R14969 VDD.n832 VDD.n784 0.0282778
R14970 VDD.n776 VDD.n770 0.0282778
R14971 VDD.n762 VDD.n756 0.0282778
R14972 VDD.n748 VDD.n742 0.0282778
R14973 VDD.n516 VDD.n510 0.0282778
R14974 VDD.n2573 VDD.n509 0.0282778
R14975 VDD.n6098 VDD.n6089 0.0282778
R14976 VDD.n6123 VDD.n6088 0.0282778
R14977 VDD.n6356 VDD.n6350 0.0282778
R14978 VDD.n6369 VDD.n6349 0.0282778
R14979 VDD.n6382 VDD.n6348 0.0282778
R14980 VDD.n6395 VDD.n6347 0.0282778
R14981 VDD.n6339 VDD.n6333 0.0282778
R14982 VDD.n6325 VDD.n6319 0.0282778
R14983 VDD.n6311 VDD.n6305 0.0282778
R14984 VDD.n6079 VDD.n6073 0.0282778
R14985 VDD.n8136 VDD.n6072 0.0282778
R14986 VDD.n5160 VDD.n3335 0.0282391
R14987 VDD.n2566 VDD.n741 0.0282391
R14988 VDD.n8129 VDD.n6304 0.0282391
R14989 VDD.n5142 VDD.n3457 0.0263621
R14990 VDD.n4592 VDD.n3458 0.0263621
R14991 VDD.n4593 VDD.n4592 0.0263621
R14992 VDD.n4601 VDD.n4593 0.0263621
R14993 VDD.n4601 VDD.n4600 0.0263621
R14994 VDD.n4600 VDD.n4594 0.0263621
R14995 VDD.n4594 VDD.n3989 0.0263621
R14996 VDD.n4677 VDD.n3989 0.0263621
R14997 VDD.n4678 VDD.n4677 0.0263621
R14998 VDD.n4682 VDD.n4678 0.0263621
R14999 VDD.n4682 VDD.n4681 0.0263621
R15000 VDD.n4681 VDD.n3955 0.0263621
R15001 VDD.n4710 VDD.n3955 0.0263621
R15002 VDD.n4711 VDD.n4710 0.0263621
R15003 VDD.n4711 VDD.n3790 0.0263621
R15004 VDD.n5138 VDD.n3791 0.0263621
R15005 VDD.n2548 VDD.n863 0.0263621
R15006 VDD.n1998 VDD.n864 0.0263621
R15007 VDD.n1999 VDD.n1998 0.0263621
R15008 VDD.n2007 VDD.n1999 0.0263621
R15009 VDD.n2007 VDD.n2006 0.0263621
R15010 VDD.n2006 VDD.n2000 0.0263621
R15011 VDD.n2000 VDD.n1395 0.0263621
R15012 VDD.n2083 VDD.n1395 0.0263621
R15013 VDD.n2084 VDD.n2083 0.0263621
R15014 VDD.n2088 VDD.n2084 0.0263621
R15015 VDD.n2088 VDD.n2087 0.0263621
R15016 VDD.n2087 VDD.n1361 0.0263621
R15017 VDD.n2116 VDD.n1361 0.0263621
R15018 VDD.n2117 VDD.n2116 0.0263621
R15019 VDD.n2117 VDD.n1196 0.0263621
R15020 VDD.n2544 VDD.n1197 0.0263621
R15021 VDD.n8111 VDD.n6426 0.0263621
R15022 VDD.n7561 VDD.n6427 0.0263621
R15023 VDD.n7562 VDD.n7561 0.0263621
R15024 VDD.n7570 VDD.n7562 0.0263621
R15025 VDD.n7570 VDD.n7569 0.0263621
R15026 VDD.n7569 VDD.n7563 0.0263621
R15027 VDD.n7563 VDD.n6958 0.0263621
R15028 VDD.n7646 VDD.n6958 0.0263621
R15029 VDD.n7647 VDD.n7646 0.0263621
R15030 VDD.n7651 VDD.n7647 0.0263621
R15031 VDD.n7651 VDD.n7650 0.0263621
R15032 VDD.n7650 VDD.n6924 0.0263621
R15033 VDD.n7679 VDD.n6924 0.0263621
R15034 VDD.n7680 VDD.n7679 0.0263621
R15035 VDD.n7680 VDD.n6759 0.0263621
R15036 VDD.n8107 VDD.n6760 0.0263621
R15037 VDD.n3334 VDD.n3333 0.02635
R15038 VDD.n3434 VDD.n3433 0.02635
R15039 VDD.n740 VDD.n739 0.02635
R15040 VDD.n840 VDD.n839 0.02635
R15041 VDD.n6303 VDD.n6302 0.02635
R15042 VDD.n6403 VDD.n6402 0.02635
R15043 VDD.n3102 VDD 0.025175
R15044 VDD.n508 VDD 0.025175
R15045 VDD.n3177 VDD.n3176 0.0247833
R15046 VDD.n3235 VDD.n3177 0.0247833
R15047 VDD.n3334 VDD.n3277 0.0247833
R15048 VDD.n3294 VDD.n3221 0.0247833
R15049 VDD.n3221 VDD.n3220 0.0247833
R15050 VDD.n5174 VDD.n5161 0.0247833
R15051 VDD.n5161 VDD.n3117 0.0247833
R15052 VDD.n3434 VDD.n3377 0.0247833
R15053 VDD.n3394 VDD.n3162 0.0247833
R15054 VDD.n3162 VDD.n3161 0.0247833
R15055 VDD.n583 VDD.n582 0.0247833
R15056 VDD.n641 VDD.n583 0.0247833
R15057 VDD.n740 VDD.n683 0.0247833
R15058 VDD.n700 VDD.n627 0.0247833
R15059 VDD.n627 VDD.n626 0.0247833
R15060 VDD.n2580 VDD.n2567 0.0247833
R15061 VDD.n2567 VDD.n523 0.0247833
R15062 VDD.n840 VDD.n783 0.0247833
R15063 VDD.n800 VDD.n568 0.0247833
R15064 VDD.n568 VDD.n567 0.0247833
R15065 VDD.n6146 VDD.n6145 0.0247833
R15066 VDD.n6204 VDD.n6146 0.0247833
R15067 VDD.n6303 VDD.n6246 0.0247833
R15068 VDD.n6263 VDD.n6190 0.0247833
R15069 VDD.n6190 VDD.n6189 0.0247833
R15070 VDD.n8143 VDD.n8130 0.0247833
R15071 VDD.n8130 VDD.n6086 0.0247833
R15072 VDD.n6403 VDD.n6346 0.0247833
R15073 VDD.n6363 VDD.n6131 0.0247833
R15074 VDD.n6131 VDD.n6130 0.0247833
R15075 VDD.n4560 VDD.n3789 0.0244565
R15076 VDD.n1966 VDD.n1195 0.0244565
R15077 VDD.n7529 VDD.n6758 0.0244565
R15078 VDD.n2790 VDD.n2789 0.0240625
R15079 VDD.n196 VDD.n195 0.0240625
R15080 VDD.n5759 VDD.n5758 0.0240625
R15081 VDD.n2904 VDD.n2747 0.0240294
R15082 VDD.n2903 VDD.n2748 0.0240294
R15083 VDD.n2824 VDD.n2797 0.0240294
R15084 VDD.n2816 VDD.n2783 0.0240294
R15085 VDD.n310 VDD.n153 0.0240294
R15086 VDD.n309 VDD.n154 0.0240294
R15087 VDD.n230 VDD.n203 0.0240294
R15088 VDD.n222 VDD.n189 0.0240294
R15089 VDD.n5873 VDD.n5716 0.0240294
R15090 VDD.n5872 VDD.n5717 0.0240294
R15091 VDD.n5793 VDD.n5766 0.0240294
R15092 VDD.n5785 VDD.n5752 0.0240294
R15093 VDD VDD.n5526 0.0239375
R15094 VDD VDD.n5548 0.0239375
R15095 VDD.n5416 VDD.n5310 0.0239375
R15096 VDD.n5139 VDD.n5138 0.0234885
R15097 VDD.n2545 VDD.n2544 0.0234885
R15098 VDD.n8108 VDD.n8107 0.0234885
R15099 VDD.n3503 VDD.n3502 0.0232879
R15100 VDD.n3517 VDD.n3503 0.0232879
R15101 VDD.n3787 VDD.n3587 0.0232879
R15102 VDD.n3787 VDD.n3786 0.0232879
R15103 VDD.n3734 VDD.n3721 0.0232879
R15104 VDD.n3721 VDD.n3720 0.0232879
R15105 VDD.n3655 VDD.n3642 0.0232879
R15106 VDD.n909 VDD.n908 0.0232879
R15107 VDD.n923 VDD.n909 0.0232879
R15108 VDD.n1193 VDD.n993 0.0232879
R15109 VDD.n1193 VDD.n1192 0.0232879
R15110 VDD.n1140 VDD.n1127 0.0232879
R15111 VDD.n1127 VDD.n1126 0.0232879
R15112 VDD.n1061 VDD.n1048 0.0232879
R15113 VDD.n6472 VDD.n6471 0.0232879
R15114 VDD.n6486 VDD.n6472 0.0232879
R15115 VDD.n6756 VDD.n6556 0.0232879
R15116 VDD.n6756 VDD.n6755 0.0232879
R15117 VDD.n6703 VDD.n6690 0.0232879
R15118 VDD.n6690 VDD.n6689 0.0232879
R15119 VDD.n6624 VDD.n6611 0.0232879
R15120 VDD.n5449 VDD 0.0226354
R15121 VDD.n5428 VDD 0.0226354
R15122 VDD.n5328 VDD 0.0226354
R15123 VDD.n3642 VDD.n3641 0.0218636
R15124 VDD.n1048 VDD.n1047 0.0218636
R15125 VDD.n6611 VDD.n6610 0.0218636
R15126 VDD.n6071 VDD.n5567 0.02165
R15127 VDD VDD.n5502 0.0213333
R15128 VDD VDD.n5525 0.0213333
R15129 VDD VDD.n5316 0.0213333
R15130 VDD.n5350 VDD 0.0213333
R15131 VDD.n5375 VDD 0.0213333
R15132 VDD.n5320 VDD 0.0213333
R15133 VDD.n5439 VDD.n5438 0.0149628
R15134 VDD.n5142 VDD.n5141 0.0141494
R15135 VDD.n2548 VDD.n2547 0.0141494
R15136 VDD.n8111 VDD.n8110 0.0141494
R15137 VDD.n2789 VDD 0.0136406
R15138 VDD.n195 VDD 0.0136406
R15139 VDD.n5758 VDD 0.0136406
R15140 VDD.n5141 VDD.n3458 0.0127126
R15141 VDD.n2547 VDD.n864 0.0127126
R15142 VDD.n8110 VDD.n6427 0.0127126
R15143 VDD.n4532 VDD.n4071 0.012359
R15144 VDD.n4531 VDD.n4072 0.012359
R15145 VDD.n5152 VDD.n3446 0.012359
R15146 VDD.n5151 VDD.n3447 0.012359
R15147 VDD.n4563 VDD.n4562 0.012359
R15148 VDD.n4573 VDD.n4555 0.012359
R15149 VDD.n4572 VDD.n4556 0.012359
R15150 VDD.n4615 VDD.n4034 0.012359
R15151 VDD.n4614 VDD.n4037 0.012359
R15152 VDD.n4040 VDD.n4039 0.012359
R15153 VDD.n4657 VDD.n4003 0.012359
R15154 VDD.n4659 VDD.n4658 0.012359
R15155 VDD.n4666 VDD.n4000 0.012359
R15156 VDD.n4665 VDD.n4001 0.012359
R15157 VDD.n4694 VDD.n3971 0.012359
R15158 VDD.n4693 VDD.n3974 0.012359
R15159 VDD.n3979 VDD.n3978 0.012359
R15160 VDD.n4721 VDD.n3940 0.012359
R15161 VDD.n4720 VDD.n3943 0.012359
R15162 VDD.n5129 VDD.n3804 0.012359
R15163 VDD.n5128 VDD.n3805 0.012359
R15164 VDD.n4760 VDD.n4754 0.012359
R15165 VDD.n4765 VDD.n4764 0.012359
R15166 VDD.n1938 VDD.n1477 0.012359
R15167 VDD.n1937 VDD.n1478 0.012359
R15168 VDD.n2558 VDD.n852 0.012359
R15169 VDD.n2557 VDD.n853 0.012359
R15170 VDD.n1969 VDD.n1968 0.012359
R15171 VDD.n1979 VDD.n1961 0.012359
R15172 VDD.n1978 VDD.n1962 0.012359
R15173 VDD.n2021 VDD.n1440 0.012359
R15174 VDD.n2020 VDD.n1443 0.012359
R15175 VDD.n1446 VDD.n1445 0.012359
R15176 VDD.n2063 VDD.n1409 0.012359
R15177 VDD.n2065 VDD.n2064 0.012359
R15178 VDD.n2072 VDD.n1406 0.012359
R15179 VDD.n2071 VDD.n1407 0.012359
R15180 VDD.n2100 VDD.n1377 0.012359
R15181 VDD.n2099 VDD.n1380 0.012359
R15182 VDD.n1385 VDD.n1384 0.012359
R15183 VDD.n2127 VDD.n1346 0.012359
R15184 VDD.n2126 VDD.n1349 0.012359
R15185 VDD.n2535 VDD.n1210 0.012359
R15186 VDD.n2534 VDD.n1211 0.012359
R15187 VDD.n2166 VDD.n2160 0.012359
R15188 VDD.n2171 VDD.n2170 0.012359
R15189 VDD.n7501 VDD.n7040 0.012359
R15190 VDD.n7500 VDD.n7041 0.012359
R15191 VDD.n8121 VDD.n6415 0.012359
R15192 VDD.n8120 VDD.n6416 0.012359
R15193 VDD.n7532 VDD.n7531 0.012359
R15194 VDD.n7542 VDD.n7524 0.012359
R15195 VDD.n7541 VDD.n7525 0.012359
R15196 VDD.n7584 VDD.n7003 0.012359
R15197 VDD.n7583 VDD.n7006 0.012359
R15198 VDD.n7009 VDD.n7008 0.012359
R15199 VDD.n7626 VDD.n6972 0.012359
R15200 VDD.n7628 VDD.n7627 0.012359
R15201 VDD.n7635 VDD.n6969 0.012359
R15202 VDD.n7634 VDD.n6970 0.012359
R15203 VDD.n7663 VDD.n6940 0.012359
R15204 VDD.n7662 VDD.n6943 0.012359
R15205 VDD.n6948 VDD.n6947 0.012359
R15206 VDD.n7690 VDD.n6909 0.012359
R15207 VDD.n7689 VDD.n6912 0.012359
R15208 VDD.n8098 VDD.n6773 0.012359
R15209 VDD.n8097 VDD.n6774 0.012359
R15210 VDD.n7729 VDD.n7723 0.012359
R15211 VDD.n7734 VDD.n7733 0.012359
R15212 VDD.n5308 VDD.n5305 0.0121
R15213 VDD.n5305 VDD.n5304 0.0121
R15214 VDD.n4532 VDD.n4531 0.0117179
R15215 VDD.n4072 VDD.n3446 0.0117179
R15216 VDD.n5152 VDD.n5151 0.0117179
R15217 VDD.n4563 VDD.n3447 0.0117179
R15218 VDD.n4573 VDD.n4572 0.0117179
R15219 VDD.n4556 VDD.n4034 0.0117179
R15220 VDD.n4615 VDD.n4614 0.0117179
R15221 VDD.n4040 VDD.n4037 0.0117179
R15222 VDD.n4039 VDD.n4003 0.0117179
R15223 VDD.n4659 VDD.n4657 0.0117179
R15224 VDD.n4658 VDD.n4000 0.0117179
R15225 VDD.n4666 VDD.n4665 0.0117179
R15226 VDD.n4001 VDD.n3971 0.0117179
R15227 VDD.n4694 VDD.n4693 0.0117179
R15228 VDD.n3979 VDD.n3974 0.0117179
R15229 VDD.n3978 VDD.n3940 0.0117179
R15230 VDD.n4721 VDD.n4720 0.0117179
R15231 VDD.n4557 VDD.n3943 0.0117179
R15232 VDD.n4558 VDD.n3804 0.0117179
R15233 VDD.n5129 VDD.n5128 0.0117179
R15234 VDD.n4754 VDD.n3805 0.0117179
R15235 VDD.n4764 VDD.n4760 0.0117179
R15236 VDD.n4766 VDD.n4765 0.0117179
R15237 VDD.n1938 VDD.n1937 0.0117179
R15238 VDD.n1478 VDD.n852 0.0117179
R15239 VDD.n2558 VDD.n2557 0.0117179
R15240 VDD.n1969 VDD.n853 0.0117179
R15241 VDD.n1979 VDD.n1978 0.0117179
R15242 VDD.n1962 VDD.n1440 0.0117179
R15243 VDD.n2021 VDD.n2020 0.0117179
R15244 VDD.n1446 VDD.n1443 0.0117179
R15245 VDD.n1445 VDD.n1409 0.0117179
R15246 VDD.n2065 VDD.n2063 0.0117179
R15247 VDD.n2064 VDD.n1406 0.0117179
R15248 VDD.n2072 VDD.n2071 0.0117179
R15249 VDD.n1407 VDD.n1377 0.0117179
R15250 VDD.n2100 VDD.n2099 0.0117179
R15251 VDD.n1385 VDD.n1380 0.0117179
R15252 VDD.n1384 VDD.n1346 0.0117179
R15253 VDD.n2127 VDD.n2126 0.0117179
R15254 VDD.n1963 VDD.n1349 0.0117179
R15255 VDD.n1964 VDD.n1210 0.0117179
R15256 VDD.n2535 VDD.n2534 0.0117179
R15257 VDD.n2160 VDD.n1211 0.0117179
R15258 VDD.n2170 VDD.n2166 0.0117179
R15259 VDD.n2172 VDD.n2171 0.0117179
R15260 VDD.n7501 VDD.n7500 0.0117179
R15261 VDD.n7041 VDD.n6415 0.0117179
R15262 VDD.n8121 VDD.n8120 0.0117179
R15263 VDD.n7532 VDD.n6416 0.0117179
R15264 VDD.n7542 VDD.n7541 0.0117179
R15265 VDD.n7525 VDD.n7003 0.0117179
R15266 VDD.n7584 VDD.n7583 0.0117179
R15267 VDD.n7009 VDD.n7006 0.0117179
R15268 VDD.n7008 VDD.n6972 0.0117179
R15269 VDD.n7628 VDD.n7626 0.0117179
R15270 VDD.n7627 VDD.n6969 0.0117179
R15271 VDD.n7635 VDD.n7634 0.0117179
R15272 VDD.n6970 VDD.n6940 0.0117179
R15273 VDD.n7663 VDD.n7662 0.0117179
R15274 VDD.n6948 VDD.n6943 0.0117179
R15275 VDD.n6947 VDD.n6909 0.0117179
R15276 VDD.n7690 VDD.n7689 0.0117179
R15277 VDD.n7526 VDD.n6912 0.0117179
R15278 VDD.n7527 VDD.n6773 0.0117179
R15279 VDD.n8098 VDD.n8097 0.0117179
R15280 VDD.n7723 VDD.n6774 0.0117179
R15281 VDD.n7733 VDD.n7729 0.0117179
R15282 VDD.n7735 VDD.n7734 0.0117179
R15283 VDD.n4561 VDD.n4555 0.0113974
R15284 VDD.n1967 VDD.n1961 0.0113974
R15285 VDD.n7530 VDD.n7524 0.0113974
R15286 VDD.n4560 VDD.n3335 0.0113225
R15287 VDD.n1966 VDD.n741 0.0113225
R15288 VDD.n7529 VDD.n6304 0.0113225
R15289 VDD.n5140 VDD.n3789 0.0110072
R15290 VDD.n2546 VDD.n1195 0.0110072
R15291 VDD.n8109 VDD.n6758 0.0110072
R15292 VDD.n3789 VDD.n3459 0.0106061
R15293 VDD.n1195 VDD.n865 0.0106061
R15294 VDD.n6758 VDD.n6428 0.0106061
R15295 VDD.n3101 VDD.n2619 0.0099
R15296 VDD.n507 VDD.n25 0.0099
R15297 VDD.n6070 VDD.n5588 0.0099
R15298 VDD.n4559 VDD.n4558 0.00979487
R15299 VDD.n1965 VDD.n1964 0.00979487
R15300 VDD.n7528 VDD.n7527 0.00979487
R15301 VDD.n3616 VDD.n3600 0.00883333
R15302 VDD.n3476 VDD.n3460 0.00883333
R15303 VDD.n1022 VDD.n1006 0.00883333
R15304 VDD.n882 VDD.n866 0.00883333
R15305 VDD.n5565 VDD.n5564 0.00883333
R15306 VDD.n6585 VDD.n6569 0.00883333
R15307 VDD.n6445 VDD.n6429 0.00883333
R15308 VDD.n3789 VDD.n3788 0.0079697
R15309 VDD.n1195 VDD.n1194 0.0079697
R15310 VDD.n6758 VDD.n6757 0.0079697
R15311 VDD.n5307 VDD.n5186 0.007165
R15312 VDD.n5309 VDD.n5186 0.007165
R15313 VDD.n2595 VDD.n2587 0.00678555
R15314 VDD.n2591 VDD.n2589 0.00678555
R15315 VDD.n2594 VDD.n2586 0.00678555
R15316 VDD.n5176 VDD.n2590 0.00678555
R15317 VDD.n2585 VDD.n2 0.00678555
R15318 VDD.n2584 VDD.n3 0.00678555
R15319 VDD.n2583 VDD.n1 0.00678555
R15320 VDD.n2582 VDD.n4 0.00678555
R15321 VDD.n8149 VDD.n5180 0.00678555
R15322 VDD.n8147 VDD.n5184 0.00678555
R15323 VDD.n5183 VDD.n5179 0.00678555
R15324 VDD.n8145 VDD.n5185 0.00678555
R15325 VDD.n8150 VDD.n8149 0.00678555
R15326 VDD.n5184 VDD.n5180 0.00678555
R15327 VDD.n8147 VDD.n5179 0.00678555
R15328 VDD.n5185 VDD.n5183 0.00678555
R15329 VDD.n8154 VDD.n2 0.00678555
R15330 VDD.n2585 VDD.n2584 0.00678555
R15331 VDD.n2583 VDD.n3 0.00678555
R15332 VDD.n4 VDD.n1 0.00678555
R15333 VDD.n2596 VDD.n2595 0.00678555
R15334 VDD.n2591 VDD.n2587 0.00678555
R15335 VDD.n2594 VDD.n2589 0.00678555
R15336 VDD.n2590 VDD.n2586 0.00678555
R15337 VDD.n5306 VDD.n5303 0.0067128
R15338 VDD.n5306 VDD.n5304 0.0067128
R15339 VDD.n8148 VDD.n5182 0.0063
R15340 VDD.n2593 VDD.n2592 0.0063
R15341 VDD VDD.n0 0.00485
R15342 VDD.n8146 VDD.n5181 0.00387804
R15343 VDD.n8151 VDD.n5178 0.00387804
R15344 VDD.n8153 VDD.n8152 0.00387804
R15345 VDD.n8156 VDD.n8155 0.00387804
R15346 VDD.n5177 VDD.n2588 0.00387804
R15347 VDD.n2598 VDD.n2597 0.00387804
R15348 VDD.n5182 VDD.n5181 0.00387804
R15349 VDD.n8148 VDD.n5178 0.00387804
R15350 VDD.n8153 VDD.n0 0.00387804
R15351 VDD.n8157 VDD.n8156 0.00387804
R15352 VDD.n2592 VDD.n2588 0.00387804
R15353 VDD.n2598 VDD.n2593 0.00387804
R15354 VDD.n2597 VDD 0.0034
R15355 VDD.n5139 VDD.n3790 0.00337356
R15356 VDD.n2545 VDD.n1196 0.00337356
R15357 VDD.n8108 VDD.n6759 0.00337356
R15358 VDD.n4559 VDD.n4557 0.0030641
R15359 VDD.n1965 VDD.n1963 0.0030641
R15360 VDD.n7528 VDD.n7526 0.0030641
R15361 VDD.n5567 VDD 0.00285
R15362 VDD VDD.n8157 0.00195
R15363 VDD.n4562 VDD.n4561 0.000820513
R15364 VDD.n1968 VDD.n1967 0.000820513
R15365 VDD.n7531 VDD.n7530 0.000820513
R15366 a_216625_n11375.n178 a_216625_n11375.n177 815.966
R15367 a_216625_n11375.n317 a_216625_n11375.n311 585
R15368 a_216625_n11375.n317 a_216625_n11375.n310 585
R15369 a_216625_n11375.n318 a_216625_n11375.n317 585
R15370 a_216625_n11375.n303 a_216625_n11375.n297 585
R15371 a_216625_n11375.n303 a_216625_n11375.n296 585
R15372 a_216625_n11375.n304 a_216625_n11375.n303 585
R15373 a_216625_n11375.n289 a_216625_n11375.n283 585
R15374 a_216625_n11375.n289 a_216625_n11375.n282 585
R15375 a_216625_n11375.n290 a_216625_n11375.n289 585
R15376 a_216625_n11375.n275 a_216625_n11375.n269 585
R15377 a_216625_n11375.n275 a_216625_n11375.n268 585
R15378 a_216625_n11375.n276 a_216625_n11375.n275 585
R15379 a_216625_n11375.n261 a_216625_n11375.n255 585
R15380 a_216625_n11375.n261 a_216625_n11375.n254 585
R15381 a_216625_n11375.n262 a_216625_n11375.n261 585
R15382 a_216625_n11375.n247 a_216625_n11375.n241 585
R15383 a_216625_n11375.n247 a_216625_n11375.n240 585
R15384 a_216625_n11375.n248 a_216625_n11375.n247 585
R15385 a_216625_n11375.n233 a_216625_n11375.n227 585
R15386 a_216625_n11375.n233 a_216625_n11375.n226 585
R15387 a_216625_n11375.n234 a_216625_n11375.n233 585
R15388 a_216625_n11375.n219 a_216625_n11375.n213 585
R15389 a_216625_n11375.n219 a_216625_n11375.n212 585
R15390 a_216625_n11375.n220 a_216625_n11375.n219 585
R15391 a_216625_n11375.n205 a_216625_n11375.n199 585
R15392 a_216625_n11375.n205 a_216625_n11375.n198 585
R15393 a_216625_n11375.n206 a_216625_n11375.n205 585
R15394 a_216625_n11375.n191 a_216625_n11375.n185 585
R15395 a_216625_n11375.n191 a_216625_n11375.n184 585
R15396 a_216625_n11375.n192 a_216625_n11375.n191 585
R15397 a_216625_n11375.n162 a_216625_n11375.n161 585
R15398 a_216625_n11375.n159 a_216625_n11375.n158 585
R15399 a_216625_n11375.n169 a_216625_n11375.n168 585
R15400 a_216625_n11375.n171 a_216625_n11375.n170 585
R15401 a_216625_n11375.n156 a_216625_n11375.n155 585
R15402 a_216625_n11375.n177 a_216625_n11375.n176 585
R15403 a_216625_n11375.n102 a_216625_n11375.t66 433.149
R15404 a_216625_n11375.t66 a_216625_n11375.n86 433.149
R15405 a_216625_n11375.n101 a_216625_n11375.t50 433.149
R15406 a_216625_n11375.t50 a_216625_n11375.n100 433.149
R15407 a_216625_n11375.t45 a_216625_n11375.n88 433.149
R15408 a_216625_n11375.n99 a_216625_n11375.t45 433.149
R15409 a_216625_n11375.t37 a_216625_n11375.n97 433.149
R15410 a_216625_n11375.n98 a_216625_n11375.t37 433.149
R15411 a_216625_n11375.n96 a_216625_n11375.t32 433.149
R15412 a_216625_n11375.t32 a_216625_n11375.n89 433.149
R15413 a_216625_n11375.n95 a_216625_n11375.t44 433.149
R15414 a_216625_n11375.t44 a_216625_n11375.n94 433.149
R15415 a_216625_n11375.t62 a_216625_n11375.n90 433.149
R15416 a_216625_n11375.n93 a_216625_n11375.t62 433.149
R15417 a_216625_n11375.t38 a_216625_n11375.n148 433.149
R15418 a_216625_n11375.n149 a_216625_n11375.t38 433.149
R15419 a_216625_n11375.t35 a_216625_n11375.n4 433.149
R15420 a_216625_n11375.n5 a_216625_n11375.t35 433.149
R15421 a_216625_n11375.t52 a_216625_n11375.n113 433.149
R15422 a_216625_n11375.n114 a_216625_n11375.t52 433.149
R15423 a_216625_n11375.n116 a_216625_n11375.t47 433.149
R15424 a_216625_n11375.t47 a_216625_n11375.n115 433.149
R15425 a_216625_n11375.n117 a_216625_n11375.t43 433.149
R15426 a_216625_n11375.t43 a_216625_n11375.n112 433.149
R15427 a_216625_n11375.t34 a_216625_n11375.n118 433.149
R15428 a_216625_n11375.n119 a_216625_n11375.t34 433.149
R15429 a_216625_n11375.t70 a_216625_n11375.n111 433.149
R15430 a_216625_n11375.n120 a_216625_n11375.t70 433.149
R15431 a_216625_n11375.n122 a_216625_n11375.t49 433.149
R15432 a_216625_n11375.t49 a_216625_n11375.n121 433.149
R15433 a_216625_n11375.n123 a_216625_n11375.t48 433.149
R15434 a_216625_n11375.t48 a_216625_n11375.n110 433.149
R15435 a_216625_n11375.t40 a_216625_n11375.n124 433.149
R15436 a_216625_n11375.n125 a_216625_n11375.t40 433.149
R15437 a_216625_n11375.t68 a_216625_n11375.n109 433.149
R15438 a_216625_n11375.n126 a_216625_n11375.t68 433.149
R15439 a_216625_n11375.n128 a_216625_n11375.t64 433.149
R15440 a_216625_n11375.t64 a_216625_n11375.n127 433.149
R15441 a_216625_n11375.n129 a_216625_n11375.t60 433.149
R15442 a_216625_n11375.t60 a_216625_n11375.n108 433.149
R15443 a_216625_n11375.t57 a_216625_n11375.n130 433.149
R15444 a_216625_n11375.n131 a_216625_n11375.t57 433.149
R15445 a_216625_n11375.t51 a_216625_n11375.n107 433.149
R15446 a_216625_n11375.n132 a_216625_n11375.t51 433.149
R15447 a_216625_n11375.n134 a_216625_n11375.t46 433.149
R15448 a_216625_n11375.t46 a_216625_n11375.n133 433.149
R15449 a_216625_n11375.n135 a_216625_n11375.t42 433.149
R15450 a_216625_n11375.t42 a_216625_n11375.n106 433.149
R15451 a_216625_n11375.t56 a_216625_n11375.n136 433.149
R15452 a_216625_n11375.n137 a_216625_n11375.t56 433.149
R15453 a_216625_n11375.t55 a_216625_n11375.n105 433.149
R15454 a_216625_n11375.n138 a_216625_n11375.t55 433.149
R15455 a_216625_n11375.n140 a_216625_n11375.t63 433.149
R15456 a_216625_n11375.t63 a_216625_n11375.n139 433.149
R15457 a_216625_n11375.n141 a_216625_n11375.t59 433.149
R15458 a_216625_n11375.t59 a_216625_n11375.n104 433.149
R15459 a_216625_n11375.t53 a_216625_n11375.n142 433.149
R15460 a_216625_n11375.n143 a_216625_n11375.t53 433.149
R15461 a_216625_n11375.t33 a_216625_n11375.n103 433.149
R15462 a_216625_n11375.n144 a_216625_n11375.t33 433.149
R15463 a_216625_n11375.n146 a_216625_n11375.t67 433.149
R15464 a_216625_n11375.t67 a_216625_n11375.n145 433.149
R15465 a_216625_n11375.n147 a_216625_n11375.t58 433.149
R15466 a_216625_n11375.t58 a_216625_n11375.n87 433.149
R15467 a_216625_n11375.n324 a_216625_n11375.t39 433.149
R15468 a_216625_n11375.t39 a_216625_n11375.n323 433.149
R15469 a_216625_n11375.t36 a_216625_n11375.n0 433.149
R15470 a_216625_n11375.n334 a_216625_n11375.t36 433.149
R15471 a_216625_n11375.t71 a_216625_n11375.n332 433.149
R15472 a_216625_n11375.n333 a_216625_n11375.t71 433.149
R15473 a_216625_n11375.n331 a_216625_n11375.t61 433.149
R15474 a_216625_n11375.t61 a_216625_n11375.n1 433.149
R15475 a_216625_n11375.n330 a_216625_n11375.t54 433.149
R15476 a_216625_n11375.t54 a_216625_n11375.n329 433.149
R15477 a_216625_n11375.t41 a_216625_n11375.n2 433.149
R15478 a_216625_n11375.n328 a_216625_n11375.t41 433.149
R15479 a_216625_n11375.t69 a_216625_n11375.n326 433.149
R15480 a_216625_n11375.n327 a_216625_n11375.t69 433.149
R15481 a_216625_n11375.n325 a_216625_n11375.t65 433.149
R15482 a_216625_n11375.t65 a_216625_n11375.n3 433.149
R15483 a_216625_n11375.t20 a_216625_n11375.n160 384.339
R15484 a_216625_n11375.n16 a_216625_n11375.n15 325.69
R15485 a_216625_n11375.n161 a_216625_n11375.n158 230.966
R15486 a_216625_n11375.n169 a_216625_n11375.n158 230.966
R15487 a_216625_n11375.n170 a_216625_n11375.n169 230.966
R15488 a_216625_n11375.n170 a_216625_n11375.n155 230.966
R15489 a_216625_n11375.n177 a_216625_n11375.n155 230.966
R15490 a_216625_n11375.n17 a_216625_n11375.n16 185
R15491 a_216625_n11375.n12 a_216625_n11375.n11 185
R15492 a_216625_n11375.n24 a_216625_n11375.n23 185
R15493 a_216625_n11375.n25 a_216625_n11375.n9 185
R15494 a_216625_n11375.n30 a_216625_n11375.n29 185
R15495 a_216625_n11375.n28 a_216625_n11375.n27 185
R15496 a_216625_n11375.n42 a_216625_n11375.n39 185
R15497 a_216625_n11375.n44 a_216625_n11375.n39 185
R15498 a_216625_n11375.n40 a_216625_n11375.n39 185
R15499 a_216625_n11375.n49 a_216625_n11375.n39 185
R15500 a_216625_n11375.n58 a_216625_n11375.n55 185
R15501 a_216625_n11375.n60 a_216625_n11375.n55 185
R15502 a_216625_n11375.n56 a_216625_n11375.n55 185
R15503 a_216625_n11375.n65 a_216625_n11375.n55 185
R15504 a_216625_n11375.n74 a_216625_n11375.n71 185
R15505 a_216625_n11375.n76 a_216625_n11375.n71 185
R15506 a_216625_n11375.n72 a_216625_n11375.n71 185
R15507 a_216625_n11375.n81 a_216625_n11375.n71 185
R15508 a_216625_n11375.n26 a_216625_n11375.t7 174.857
R15509 a_216625_n11375.n16 a_216625_n11375.n11 140.69
R15510 a_216625_n11375.n24 a_216625_n11375.n11 140.69
R15511 a_216625_n11375.n25 a_216625_n11375.n24 140.69
R15512 a_216625_n11375.n29 a_216625_n11375.n25 140.69
R15513 a_216625_n11375.n29 a_216625_n11375.n28 140.69
R15514 a_216625_n11375.n161 a_216625_n11375.t20 115.484
R15515 a_216625_n11375.n28 a_216625_n11375.t7 70.3453
R15516 a_216625_n11375.n317 a_216625_n11375.n316 51.6891
R15517 a_216625_n11375.n303 a_216625_n11375.n302 51.6891
R15518 a_216625_n11375.n289 a_216625_n11375.n288 51.6891
R15519 a_216625_n11375.n275 a_216625_n11375.n274 51.6891
R15520 a_216625_n11375.n261 a_216625_n11375.n260 51.6891
R15521 a_216625_n11375.n247 a_216625_n11375.n246 51.6891
R15522 a_216625_n11375.n233 a_216625_n11375.n232 51.6891
R15523 a_216625_n11375.n219 a_216625_n11375.n218 51.6891
R15524 a_216625_n11375.n205 a_216625_n11375.n204 51.6891
R15525 a_216625_n11375.n191 a_216625_n11375.n190 51.6891
R15526 a_216625_n11375.n316 a_216625_n11375.n315 29.8062
R15527 a_216625_n11375.n302 a_216625_n11375.n301 29.8062
R15528 a_216625_n11375.n288 a_216625_n11375.n287 29.8062
R15529 a_216625_n11375.n274 a_216625_n11375.n273 29.8062
R15530 a_216625_n11375.n260 a_216625_n11375.n259 29.8062
R15531 a_216625_n11375.n246 a_216625_n11375.n245 29.8062
R15532 a_216625_n11375.n232 a_216625_n11375.n231 29.8062
R15533 a_216625_n11375.n218 a_216625_n11375.n217 29.8062
R15534 a_216625_n11375.n204 a_216625_n11375.n203 29.8062
R15535 a_216625_n11375.n190 a_216625_n11375.n189 29.8062
R15536 a_216625_n11375.n162 a_216625_n11375.n160 29.3167
R15537 a_216625_n11375.n27 a_216625_n11375.n26 28.4333
R15538 a_216625_n11375.n51 a_216625_n11375.n50 26.8428
R15539 a_216625_n11375.n67 a_216625_n11375.n66 26.8428
R15540 a_216625_n11375.n83 a_216625_n11375.n82 26.8428
R15541 a_216625_n11375.n163 a_216625_n11375.n159 24.8476
R15542 a_216625_n11375.n30 a_216625_n11375.n10 24.8476
R15543 a_216625_n11375.n168 a_216625_n11375.n167 23.3417
R15544 a_216625_n11375.n31 a_216625_n11375.n9 23.3417
R15545 a_216625_n11375.n171 a_216625_n11375.n157 21.8358
R15546 a_216625_n11375.n23 a_216625_n11375.n22 21.8358
R15547 a_216625_n11375.n50 a_216625_n11375.n49 21.8358
R15548 a_216625_n11375.n66 a_216625_n11375.n65 21.8358
R15549 a_216625_n11375.n82 a_216625_n11375.n81 21.8358
R15550 a_216625_n11375.n315 a_216625_n11375.n311 20.3299
R15551 a_216625_n11375.n301 a_216625_n11375.n297 20.3299
R15552 a_216625_n11375.n287 a_216625_n11375.n283 20.3299
R15553 a_216625_n11375.n273 a_216625_n11375.n269 20.3299
R15554 a_216625_n11375.n259 a_216625_n11375.n255 20.3299
R15555 a_216625_n11375.n245 a_216625_n11375.n241 20.3299
R15556 a_216625_n11375.n231 a_216625_n11375.n227 20.3299
R15557 a_216625_n11375.n217 a_216625_n11375.n213 20.3299
R15558 a_216625_n11375.n203 a_216625_n11375.n199 20.3299
R15559 a_216625_n11375.n189 a_216625_n11375.n185 20.3299
R15560 a_216625_n11375.n172 a_216625_n11375.n156 20.3299
R15561 a_216625_n11375.n21 a_216625_n11375.n12 20.3299
R15562 a_216625_n11375.n48 a_216625_n11375.n40 20.3299
R15563 a_216625_n11375.n64 a_216625_n11375.n56 20.3299
R15564 a_216625_n11375.n80 a_216625_n11375.n72 20.3299
R15565 a_216625_n11375.n319 a_216625_n11375.n318 19.1618
R15566 a_216625_n11375.n305 a_216625_n11375.n304 19.1618
R15567 a_216625_n11375.n291 a_216625_n11375.n290 19.1618
R15568 a_216625_n11375.n277 a_216625_n11375.n276 19.1618
R15569 a_216625_n11375.n263 a_216625_n11375.n262 19.1618
R15570 a_216625_n11375.n249 a_216625_n11375.n248 19.1618
R15571 a_216625_n11375.n235 a_216625_n11375.n234 19.1618
R15572 a_216625_n11375.n221 a_216625_n11375.n220 19.1618
R15573 a_216625_n11375.n207 a_216625_n11375.n206 19.1618
R15574 a_216625_n11375.n193 a_216625_n11375.n192 19.1618
R15575 a_216625_n11375.n179 a_216625_n11375.n178 19.1618
R15576 a_216625_n11375.n15 a_216625_n11375.n6 19.1618
R15577 a_216625_n11375.n42 a_216625_n11375.n37 19.1618
R15578 a_216625_n11375.n58 a_216625_n11375.n36 19.1618
R15579 a_216625_n11375.n74 a_216625_n11375.n35 19.1618
R15580 a_216625_n11375.n312 a_216625_n11375.n310 18.824
R15581 a_216625_n11375.n298 a_216625_n11375.n296 18.824
R15582 a_216625_n11375.n284 a_216625_n11375.n282 18.824
R15583 a_216625_n11375.n270 a_216625_n11375.n268 18.824
R15584 a_216625_n11375.n256 a_216625_n11375.n254 18.824
R15585 a_216625_n11375.n242 a_216625_n11375.n240 18.824
R15586 a_216625_n11375.n228 a_216625_n11375.n226 18.824
R15587 a_216625_n11375.n214 a_216625_n11375.n212 18.824
R15588 a_216625_n11375.n200 a_216625_n11375.n198 18.824
R15589 a_216625_n11375.n186 a_216625_n11375.n184 18.824
R15590 a_216625_n11375.n176 a_216625_n11375.n175 18.824
R15591 a_216625_n11375.n18 a_216625_n11375.n17 18.824
R15592 a_216625_n11375.n45 a_216625_n11375.n44 18.824
R15593 a_216625_n11375.n61 a_216625_n11375.n60 18.824
R15594 a_216625_n11375.n77 a_216625_n11375.n76 18.824
R15595 a_216625_n11375.n318 a_216625_n11375.n309 17.3181
R15596 a_216625_n11375.n304 a_216625_n11375.n295 17.3181
R15597 a_216625_n11375.n290 a_216625_n11375.n281 17.3181
R15598 a_216625_n11375.n276 a_216625_n11375.n267 17.3181
R15599 a_216625_n11375.n262 a_216625_n11375.n253 17.3181
R15600 a_216625_n11375.n248 a_216625_n11375.n239 17.3181
R15601 a_216625_n11375.n234 a_216625_n11375.n225 17.3181
R15602 a_216625_n11375.n220 a_216625_n11375.n211 17.3181
R15603 a_216625_n11375.n206 a_216625_n11375.n197 17.3181
R15604 a_216625_n11375.n192 a_216625_n11375.n183 17.3181
R15605 a_216625_n11375.n178 a_216625_n11375.n154 17.3181
R15606 a_216625_n11375.n15 a_216625_n11375.n14 17.3181
R15607 a_216625_n11375.n43 a_216625_n11375.n42 17.3181
R15608 a_216625_n11375.n59 a_216625_n11375.n58 17.3181
R15609 a_216625_n11375.n75 a_216625_n11375.n74 17.3181
R15610 a_216625_n11375.n51 a_216625_n11375.n39 16.7801
R15611 a_216625_n11375.n67 a_216625_n11375.n55 16.7801
R15612 a_216625_n11375.n83 a_216625_n11375.n71 16.7801
R15613 a_216625_n11375.n309 a_216625_n11375.n308 9.3005
R15614 a_216625_n11375.n315 a_216625_n11375.n314 9.3005
R15615 a_216625_n11375.n313 a_216625_n11375.n312 9.3005
R15616 a_216625_n11375.n295 a_216625_n11375.n294 9.3005
R15617 a_216625_n11375.n301 a_216625_n11375.n300 9.3005
R15618 a_216625_n11375.n299 a_216625_n11375.n298 9.3005
R15619 a_216625_n11375.n281 a_216625_n11375.n280 9.3005
R15620 a_216625_n11375.n287 a_216625_n11375.n286 9.3005
R15621 a_216625_n11375.n285 a_216625_n11375.n284 9.3005
R15622 a_216625_n11375.n267 a_216625_n11375.n266 9.3005
R15623 a_216625_n11375.n273 a_216625_n11375.n272 9.3005
R15624 a_216625_n11375.n271 a_216625_n11375.n270 9.3005
R15625 a_216625_n11375.n253 a_216625_n11375.n252 9.3005
R15626 a_216625_n11375.n259 a_216625_n11375.n258 9.3005
R15627 a_216625_n11375.n257 a_216625_n11375.n256 9.3005
R15628 a_216625_n11375.n239 a_216625_n11375.n238 9.3005
R15629 a_216625_n11375.n245 a_216625_n11375.n244 9.3005
R15630 a_216625_n11375.n243 a_216625_n11375.n242 9.3005
R15631 a_216625_n11375.n225 a_216625_n11375.n224 9.3005
R15632 a_216625_n11375.n231 a_216625_n11375.n230 9.3005
R15633 a_216625_n11375.n229 a_216625_n11375.n228 9.3005
R15634 a_216625_n11375.n211 a_216625_n11375.n210 9.3005
R15635 a_216625_n11375.n217 a_216625_n11375.n216 9.3005
R15636 a_216625_n11375.n215 a_216625_n11375.n214 9.3005
R15637 a_216625_n11375.n197 a_216625_n11375.n196 9.3005
R15638 a_216625_n11375.n203 a_216625_n11375.n202 9.3005
R15639 a_216625_n11375.n201 a_216625_n11375.n200 9.3005
R15640 a_216625_n11375.n183 a_216625_n11375.n182 9.3005
R15641 a_216625_n11375.n189 a_216625_n11375.n188 9.3005
R15642 a_216625_n11375.n187 a_216625_n11375.n186 9.3005
R15643 a_216625_n11375.n164 a_216625_n11375.n163 9.3005
R15644 a_216625_n11375.n167 a_216625_n11375.n166 9.3005
R15645 a_216625_n11375.n154 a_216625_n11375.n153 9.3005
R15646 a_216625_n11375.n173 a_216625_n11375.n172 9.3005
R15647 a_216625_n11375.n175 a_216625_n11375.n174 9.3005
R15648 a_216625_n11375.n165 a_216625_n11375.n157 9.3005
R15649 a_216625_n11375.n10 a_216625_n11375.n8 9.3005
R15650 a_216625_n11375.n32 a_216625_n11375.n31 9.3005
R15651 a_216625_n11375.n22 a_216625_n11375.n7 9.3005
R15652 a_216625_n11375.n21 a_216625_n11375.n20 9.3005
R15653 a_216625_n11375.n19 a_216625_n11375.n18 9.3005
R15654 a_216625_n11375.n14 a_216625_n11375.n13 9.3005
R15655 a_216625_n11375.n50 a_216625_n11375.n38 9.3005
R15656 a_216625_n11375.n48 a_216625_n11375.n47 9.3005
R15657 a_216625_n11375.n46 a_216625_n11375.n45 9.3005
R15658 a_216625_n11375.n43 a_216625_n11375.n41 9.3005
R15659 a_216625_n11375.n66 a_216625_n11375.n54 9.3005
R15660 a_216625_n11375.n64 a_216625_n11375.n63 9.3005
R15661 a_216625_n11375.n62 a_216625_n11375.n61 9.3005
R15662 a_216625_n11375.n59 a_216625_n11375.n57 9.3005
R15663 a_216625_n11375.n82 a_216625_n11375.n70 9.3005
R15664 a_216625_n11375.n80 a_216625_n11375.n79 9.3005
R15665 a_216625_n11375.n78 a_216625_n11375.n77 9.3005
R15666 a_216625_n11375.n75 a_216625_n11375.n73 9.3005
R15667 a_216625_n11375.n310 a_216625_n11375.n309 8.28285
R15668 a_216625_n11375.n296 a_216625_n11375.n295 8.28285
R15669 a_216625_n11375.n282 a_216625_n11375.n281 8.28285
R15670 a_216625_n11375.n268 a_216625_n11375.n267 8.28285
R15671 a_216625_n11375.n254 a_216625_n11375.n253 8.28285
R15672 a_216625_n11375.n240 a_216625_n11375.n239 8.28285
R15673 a_216625_n11375.n226 a_216625_n11375.n225 8.28285
R15674 a_216625_n11375.n212 a_216625_n11375.n211 8.28285
R15675 a_216625_n11375.n198 a_216625_n11375.n197 8.28285
R15676 a_216625_n11375.n184 a_216625_n11375.n183 8.28285
R15677 a_216625_n11375.n176 a_216625_n11375.n154 8.28285
R15678 a_216625_n11375.n17 a_216625_n11375.n14 8.28285
R15679 a_216625_n11375.n44 a_216625_n11375.n43 8.28285
R15680 a_216625_n11375.n60 a_216625_n11375.n59 8.28285
R15681 a_216625_n11375.n76 a_216625_n11375.n75 8.28285
R15682 a_216625_n11375.n320 a_216625_n11375.n307 7.9105
R15683 a_216625_n11375.n306 a_216625_n11375.n293 7.9105
R15684 a_216625_n11375.n292 a_216625_n11375.n279 7.9105
R15685 a_216625_n11375.n278 a_216625_n11375.n265 7.9105
R15686 a_216625_n11375.n264 a_216625_n11375.n251 7.9105
R15687 a_216625_n11375.n250 a_216625_n11375.n237 7.9105
R15688 a_216625_n11375.n236 a_216625_n11375.n223 7.9105
R15689 a_216625_n11375.n222 a_216625_n11375.n209 7.9105
R15690 a_216625_n11375.n208 a_216625_n11375.n195 7.9105
R15691 a_216625_n11375.n194 a_216625_n11375.n181 7.9105
R15692 a_216625_n11375.n180 a_216625_n11375.n152 7.9105
R15693 a_216625_n11375.n34 a_216625_n11375.n6 7.9105
R15694 a_216625_n11375.n53 a_216625_n11375.n37 7.9105
R15695 a_216625_n11375.n69 a_216625_n11375.n36 7.9105
R15696 a_216625_n11375.n85 a_216625_n11375.n35 7.9105
R15697 a_216625_n11375.n85 a_216625_n11375.n84 7.9105
R15698 a_216625_n11375.n69 a_216625_n11375.n68 7.9105
R15699 a_216625_n11375.n53 a_216625_n11375.n52 7.9105
R15700 a_216625_n11375.n34 a_216625_n11375.n33 7.9105
R15701 a_216625_n11375.n180 a_216625_n11375.n179 7.9105
R15702 a_216625_n11375.n194 a_216625_n11375.n193 7.9105
R15703 a_216625_n11375.n208 a_216625_n11375.n207 7.9105
R15704 a_216625_n11375.n222 a_216625_n11375.n221 7.9105
R15705 a_216625_n11375.n236 a_216625_n11375.n235 7.9105
R15706 a_216625_n11375.n250 a_216625_n11375.n249 7.9105
R15707 a_216625_n11375.n264 a_216625_n11375.n263 7.9105
R15708 a_216625_n11375.n278 a_216625_n11375.n277 7.9105
R15709 a_216625_n11375.n292 a_216625_n11375.n291 7.9105
R15710 a_216625_n11375.n306 a_216625_n11375.n305 7.9105
R15711 a_216625_n11375.n320 a_216625_n11375.n319 7.9105
R15712 a_216625_n11375.n312 a_216625_n11375.n311 6.77697
R15713 a_216625_n11375.n298 a_216625_n11375.n297 6.77697
R15714 a_216625_n11375.n284 a_216625_n11375.n283 6.77697
R15715 a_216625_n11375.n270 a_216625_n11375.n269 6.77697
R15716 a_216625_n11375.n256 a_216625_n11375.n255 6.77697
R15717 a_216625_n11375.n242 a_216625_n11375.n241 6.77697
R15718 a_216625_n11375.n228 a_216625_n11375.n227 6.77697
R15719 a_216625_n11375.n214 a_216625_n11375.n213 6.77697
R15720 a_216625_n11375.n200 a_216625_n11375.n199 6.77697
R15721 a_216625_n11375.n186 a_216625_n11375.n185 6.77697
R15722 a_216625_n11375.n175 a_216625_n11375.n156 6.77697
R15723 a_216625_n11375.n18 a_216625_n11375.n12 6.77697
R15724 a_216625_n11375.n45 a_216625_n11375.n40 6.77697
R15725 a_216625_n11375.n61 a_216625_n11375.n56 6.77697
R15726 a_216625_n11375.n77 a_216625_n11375.n72 6.77697
R15727 a_216625_n11375.n317 a_216625_n11375.t25 5.7135
R15728 a_216625_n11375.n317 a_216625_n11375.t30 5.7135
R15729 a_216625_n11375.n303 a_216625_n11375.t19 5.7135
R15730 a_216625_n11375.n303 a_216625_n11375.t1 5.7135
R15731 a_216625_n11375.n289 a_216625_n11375.t14 5.7135
R15732 a_216625_n11375.n289 a_216625_n11375.t5 5.7135
R15733 a_216625_n11375.n275 a_216625_n11375.t27 5.7135
R15734 a_216625_n11375.n275 a_216625_n11375.t11 5.7135
R15735 a_216625_n11375.n261 a_216625_n11375.t28 5.7135
R15736 a_216625_n11375.n261 a_216625_n11375.t29 5.7135
R15737 a_216625_n11375.n247 a_216625_n11375.t6 5.7135
R15738 a_216625_n11375.n247 a_216625_n11375.t18 5.7135
R15739 a_216625_n11375.n233 a_216625_n11375.t17 5.7135
R15740 a_216625_n11375.n233 a_216625_n11375.t15 5.7135
R15741 a_216625_n11375.n219 a_216625_n11375.t9 5.7135
R15742 a_216625_n11375.n219 a_216625_n11375.t4 5.7135
R15743 a_216625_n11375.n205 a_216625_n11375.t3 5.7135
R15744 a_216625_n11375.n205 a_216625_n11375.t21 5.7135
R15745 a_216625_n11375.n191 a_216625_n11375.t16 5.7135
R15746 a_216625_n11375.n191 a_216625_n11375.t2 5.7135
R15747 a_216625_n11375.n151 a_216625_n11375.n150 5.58552
R15748 a_216625_n11375.n322 a_216625_n11375.n321 5.58552
R15749 a_216625_n11375.n26 a_216625_n11375.n8 5.33935
R15750 a_216625_n11375.n172 a_216625_n11375.n171 5.27109
R15751 a_216625_n11375.n23 a_216625_n11375.n21 5.27109
R15752 a_216625_n11375.n49 a_216625_n11375.n48 5.27109
R15753 a_216625_n11375.n65 a_216625_n11375.n64 5.27109
R15754 a_216625_n11375.n81 a_216625_n11375.n80 5.27109
R15755 a_216625_n11375.n164 a_216625_n11375.n160 4.51911
R15756 a_216625_n11375.n151 a_216625_n11375.n85 3.82472
R15757 a_216625_n11375.n321 a_216625_n11375.n34 3.80493
R15758 a_216625_n11375.n168 a_216625_n11375.n157 3.76521
R15759 a_216625_n11375.n22 a_216625_n11375.n9 3.76521
R15760 a_216625_n11375.n52 a_216625_n11375.n51 3.75827
R15761 a_216625_n11375.n68 a_216625_n11375.n67 3.75827
R15762 a_216625_n11375.n84 a_216625_n11375.n83 3.75827
R15763 a_216625_n11375.n39 a_216625_n11375.t8 3.4805
R15764 a_216625_n11375.n39 a_216625_n11375.t13 3.4805
R15765 a_216625_n11375.n55 a_216625_n11375.t26 3.4805
R15766 a_216625_n11375.n55 a_216625_n11375.t23 3.4805
R15767 a_216625_n11375.n71 a_216625_n11375.t24 3.4805
R15768 a_216625_n11375.n71 a_216625_n11375.t22 3.4805
R15769 a_216625_n11375.n316 a_216625_n11375.n307 3.43565
R15770 a_216625_n11375.n302 a_216625_n11375.n293 3.43565
R15771 a_216625_n11375.n288 a_216625_n11375.n279 3.43565
R15772 a_216625_n11375.n274 a_216625_n11375.n265 3.43565
R15773 a_216625_n11375.n260 a_216625_n11375.n251 3.43565
R15774 a_216625_n11375.n246 a_216625_n11375.n237 3.43565
R15775 a_216625_n11375.n232 a_216625_n11375.n223 3.43565
R15776 a_216625_n11375.n218 a_216625_n11375.n209 3.43565
R15777 a_216625_n11375.n204 a_216625_n11375.n195 3.43565
R15778 a_216625_n11375.n190 a_216625_n11375.n181 3.43565
R15779 a_216625_n11375.n91 a_216625_n11375.t31 2.84983
R15780 a_216625_n11375.t0 a_216625_n11375.n336 2.83411
R15781 a_216625_n11375.n91 a_216625_n11375.t10 2.7853
R15782 a_216625_n11375.n336 a_216625_n11375.t12 2.77004
R15783 a_216625_n11375.n167 a_216625_n11375.n159 2.25932
R15784 a_216625_n11375.n31 a_216625_n11375.n30 2.25932
R15785 a_216625_n11375.n321 a_216625_n11375.n320 1.75537
R15786 a_216625_n11375.n180 a_216625_n11375.n151 1.72874
R15787 a_216625_n11375.n93 a_216625_n11375.n92 1.11019
R15788 a_216625_n11375.n335 a_216625_n11375.n334 1.09519
R15789 a_216625_n11375.n92 a_216625_n11375.n90 1.06331
R15790 a_216625_n11375.n335 a_216625_n11375.n0 1.04831
R15791 a_216625_n11375.n163 a_216625_n11375.n162 0.753441
R15792 a_216625_n11375.n27 a_216625_n11375.n10 0.753441
R15793 a_216625_n11375.n327 a_216625_n11375.n3 0.3955
R15794 a_216625_n11375.n328 a_216625_n11375.n327 0.3955
R15795 a_216625_n11375.n329 a_216625_n11375.n328 0.3955
R15796 a_216625_n11375.n329 a_216625_n11375.n1 0.3955
R15797 a_216625_n11375.n333 a_216625_n11375.n1 0.3955
R15798 a_216625_n11375.n334 a_216625_n11375.n333 0.3955
R15799 a_216625_n11375.n145 a_216625_n11375.n87 0.3955
R15800 a_216625_n11375.n145 a_216625_n11375.n144 0.3955
R15801 a_216625_n11375.n144 a_216625_n11375.n143 0.3955
R15802 a_216625_n11375.n143 a_216625_n11375.n104 0.3955
R15803 a_216625_n11375.n139 a_216625_n11375.n104 0.3955
R15804 a_216625_n11375.n139 a_216625_n11375.n138 0.3955
R15805 a_216625_n11375.n138 a_216625_n11375.n137 0.3955
R15806 a_216625_n11375.n137 a_216625_n11375.n106 0.3955
R15807 a_216625_n11375.n133 a_216625_n11375.n106 0.3955
R15808 a_216625_n11375.n133 a_216625_n11375.n132 0.3955
R15809 a_216625_n11375.n132 a_216625_n11375.n131 0.3955
R15810 a_216625_n11375.n131 a_216625_n11375.n108 0.3955
R15811 a_216625_n11375.n127 a_216625_n11375.n108 0.3955
R15812 a_216625_n11375.n127 a_216625_n11375.n126 0.3955
R15813 a_216625_n11375.n126 a_216625_n11375.n125 0.3955
R15814 a_216625_n11375.n125 a_216625_n11375.n110 0.3955
R15815 a_216625_n11375.n121 a_216625_n11375.n110 0.3955
R15816 a_216625_n11375.n121 a_216625_n11375.n120 0.3955
R15817 a_216625_n11375.n120 a_216625_n11375.n119 0.3955
R15818 a_216625_n11375.n119 a_216625_n11375.n112 0.3955
R15819 a_216625_n11375.n115 a_216625_n11375.n112 0.3955
R15820 a_216625_n11375.n115 a_216625_n11375.n114 0.3955
R15821 a_216625_n11375.n114 a_216625_n11375.n5 0.3955
R15822 a_216625_n11375.n94 a_216625_n11375.n93 0.3955
R15823 a_216625_n11375.n94 a_216625_n11375.n89 0.3955
R15824 a_216625_n11375.n98 a_216625_n11375.n89 0.3955
R15825 a_216625_n11375.n99 a_216625_n11375.n98 0.3955
R15826 a_216625_n11375.n100 a_216625_n11375.n99 0.3955
R15827 a_216625_n11375.n100 a_216625_n11375.n86 0.3955
R15828 a_216625_n11375.n95 a_216625_n11375.n90 0.3955
R15829 a_216625_n11375.n96 a_216625_n11375.n95 0.3955
R15830 a_216625_n11375.n97 a_216625_n11375.n96 0.3955
R15831 a_216625_n11375.n97 a_216625_n11375.n88 0.3955
R15832 a_216625_n11375.n101 a_216625_n11375.n88 0.3955
R15833 a_216625_n11375.n102 a_216625_n11375.n101 0.3955
R15834 a_216625_n11375.n148 a_216625_n11375.n102 0.3955
R15835 a_216625_n11375.n148 a_216625_n11375.n147 0.3955
R15836 a_216625_n11375.n147 a_216625_n11375.n146 0.3955
R15837 a_216625_n11375.n146 a_216625_n11375.n103 0.3955
R15838 a_216625_n11375.n142 a_216625_n11375.n103 0.3955
R15839 a_216625_n11375.n142 a_216625_n11375.n141 0.3955
R15840 a_216625_n11375.n141 a_216625_n11375.n140 0.3955
R15841 a_216625_n11375.n140 a_216625_n11375.n105 0.3955
R15842 a_216625_n11375.n136 a_216625_n11375.n105 0.3955
R15843 a_216625_n11375.n136 a_216625_n11375.n135 0.3955
R15844 a_216625_n11375.n135 a_216625_n11375.n134 0.3955
R15845 a_216625_n11375.n134 a_216625_n11375.n107 0.3955
R15846 a_216625_n11375.n130 a_216625_n11375.n107 0.3955
R15847 a_216625_n11375.n130 a_216625_n11375.n129 0.3955
R15848 a_216625_n11375.n129 a_216625_n11375.n128 0.3955
R15849 a_216625_n11375.n128 a_216625_n11375.n109 0.3955
R15850 a_216625_n11375.n124 a_216625_n11375.n109 0.3955
R15851 a_216625_n11375.n124 a_216625_n11375.n123 0.3955
R15852 a_216625_n11375.n123 a_216625_n11375.n122 0.3955
R15853 a_216625_n11375.n122 a_216625_n11375.n111 0.3955
R15854 a_216625_n11375.n118 a_216625_n11375.n111 0.3955
R15855 a_216625_n11375.n118 a_216625_n11375.n117 0.3955
R15856 a_216625_n11375.n117 a_216625_n11375.n116 0.3955
R15857 a_216625_n11375.n116 a_216625_n11375.n113 0.3955
R15858 a_216625_n11375.n113 a_216625_n11375.n4 0.3955
R15859 a_216625_n11375.n324 a_216625_n11375.n4 0.3955
R15860 a_216625_n11375.n325 a_216625_n11375.n324 0.3955
R15861 a_216625_n11375.n326 a_216625_n11375.n325 0.3955
R15862 a_216625_n11375.n326 a_216625_n11375.n2 0.3955
R15863 a_216625_n11375.n330 a_216625_n11375.n2 0.3955
R15864 a_216625_n11375.n331 a_216625_n11375.n330 0.3955
R15865 a_216625_n11375.n332 a_216625_n11375.n331 0.3955
R15866 a_216625_n11375.n332 a_216625_n11375.n0 0.3955
R15867 a_216625_n11375.n323 a_216625_n11375.n5 0.370955
R15868 a_216625_n11375.n149 a_216625_n11375.n87 0.351864
R15869 a_216625_n11375.n92 a_216625_n11375.n91 0.349638
R15870 a_216625_n11375.n336 a_216625_n11375.n335 0.349638
R15871 a_216625_n11375.n314 a_216625_n11375.n313 0.196152
R15872 a_216625_n11375.n300 a_216625_n11375.n299 0.196152
R15873 a_216625_n11375.n286 a_216625_n11375.n285 0.196152
R15874 a_216625_n11375.n272 a_216625_n11375.n271 0.196152
R15875 a_216625_n11375.n258 a_216625_n11375.n257 0.196152
R15876 a_216625_n11375.n244 a_216625_n11375.n243 0.196152
R15877 a_216625_n11375.n230 a_216625_n11375.n229 0.196152
R15878 a_216625_n11375.n216 a_216625_n11375.n215 0.196152
R15879 a_216625_n11375.n202 a_216625_n11375.n201 0.196152
R15880 a_216625_n11375.n188 a_216625_n11375.n187 0.196152
R15881 a_216625_n11375.n166 a_216625_n11375.n164 0.196152
R15882 a_216625_n11375.n174 a_216625_n11375.n173 0.196152
R15883 a_216625_n11375.n20 a_216625_n11375.n19 0.196152
R15884 a_216625_n11375.n20 a_216625_n11375.n7 0.196152
R15885 a_216625_n11375.n47 a_216625_n11375.n46 0.196152
R15886 a_216625_n11375.n47 a_216625_n11375.n38 0.196152
R15887 a_216625_n11375.n63 a_216625_n11375.n62 0.196152
R15888 a_216625_n11375.n63 a_216625_n11375.n54 0.196152
R15889 a_216625_n11375.n79 a_216625_n11375.n78 0.196152
R15890 a_216625_n11375.n79 a_216625_n11375.n70 0.196152
R15891 a_216625_n11375.n166 a_216625_n11375.n165 0.194824
R15892 a_216625_n11375.n313 a_216625_n11375.n308 0.186853
R15893 a_216625_n11375.n299 a_216625_n11375.n294 0.186853
R15894 a_216625_n11375.n285 a_216625_n11375.n280 0.186853
R15895 a_216625_n11375.n271 a_216625_n11375.n266 0.186853
R15896 a_216625_n11375.n257 a_216625_n11375.n252 0.186853
R15897 a_216625_n11375.n243 a_216625_n11375.n238 0.186853
R15898 a_216625_n11375.n229 a_216625_n11375.n224 0.186853
R15899 a_216625_n11375.n215 a_216625_n11375.n210 0.186853
R15900 a_216625_n11375.n201 a_216625_n11375.n196 0.186853
R15901 a_216625_n11375.n187 a_216625_n11375.n182 0.186853
R15902 a_216625_n11375.n174 a_216625_n11375.n153 0.186853
R15903 a_216625_n11375.n19 a_216625_n11375.n13 0.186853
R15904 a_216625_n11375.n46 a_216625_n11375.n41 0.186853
R15905 a_216625_n11375.n62 a_216625_n11375.n57 0.186853
R15906 a_216625_n11375.n78 a_216625_n11375.n73 0.186853
R15907 a_216625_n11375.n32 a_216625_n11375.n8 0.184196
R15908 a_216625_n11375.n150 a_216625_n11375.n86 0.166409
R15909 a_216625_n11375.n322 a_216625_n11375.n3 0.131409
R15910 a_216625_n11375.n33 a_216625_n11375.n7 0.0790024
R15911 a_216625_n11375.n52 a_216625_n11375.n38 0.0790024
R15912 a_216625_n11375.n68 a_216625_n11375.n54 0.0790024
R15913 a_216625_n11375.n84 a_216625_n11375.n70 0.0790024
R15914 a_216625_n11375.n323 a_216625_n11375.n322 0.0709545
R15915 a_216625_n11375.n314 a_216625_n11375.n307 0.0572633
R15916 a_216625_n11375.n300 a_216625_n11375.n293 0.0572633
R15917 a_216625_n11375.n286 a_216625_n11375.n279 0.0572633
R15918 a_216625_n11375.n272 a_216625_n11375.n265 0.0572633
R15919 a_216625_n11375.n258 a_216625_n11375.n251 0.0572633
R15920 a_216625_n11375.n244 a_216625_n11375.n237 0.0572633
R15921 a_216625_n11375.n230 a_216625_n11375.n223 0.0572633
R15922 a_216625_n11375.n216 a_216625_n11375.n209 0.0572633
R15923 a_216625_n11375.n202 a_216625_n11375.n195 0.0572633
R15924 a_216625_n11375.n188 a_216625_n11375.n181 0.0572633
R15925 a_216625_n11375.n173 a_216625_n11375.n152 0.0572633
R15926 a_216625_n11375.n150 a_216625_n11375.n149 0.0550455
R15927 a_216625_n11375.n208 a_216625_n11375.n194 0.0506333
R15928 a_216625_n11375.n222 a_216625_n11375.n208 0.0506333
R15929 a_216625_n11375.n250 a_216625_n11375.n236 0.0506333
R15930 a_216625_n11375.n278 a_216625_n11375.n264 0.0506333
R15931 a_216625_n11375.n292 a_216625_n11375.n278 0.0506333
R15932 a_216625_n11375.n320 a_216625_n11375.n306 0.0506333
R15933 a_216625_n11375.n194 a_216625_n11375.n180 0.0490667
R15934 a_216625_n11375.n236 a_216625_n11375.n222 0.0490667
R15935 a_216625_n11375.n264 a_216625_n11375.n250 0.0490667
R15936 a_216625_n11375.n306 a_216625_n11375.n292 0.0490667
R15937 a_216625_n11375.n165 a_216625_n11375.n152 0.0477222
R15938 a_216625_n11375.n85 a_216625_n11375.n69 0.0400789
R15939 a_216625_n11375.n53 a_216625_n11375.n34 0.0400789
R15940 a_216625_n11375.n319 a_216625_n11375.n308 0.0393889
R15941 a_216625_n11375.n305 a_216625_n11375.n294 0.0393889
R15942 a_216625_n11375.n291 a_216625_n11375.n280 0.0393889
R15943 a_216625_n11375.n277 a_216625_n11375.n266 0.0393889
R15944 a_216625_n11375.n263 a_216625_n11375.n252 0.0393889
R15945 a_216625_n11375.n249 a_216625_n11375.n238 0.0393889
R15946 a_216625_n11375.n235 a_216625_n11375.n224 0.0393889
R15947 a_216625_n11375.n221 a_216625_n11375.n210 0.0393889
R15948 a_216625_n11375.n207 a_216625_n11375.n196 0.0393889
R15949 a_216625_n11375.n193 a_216625_n11375.n182 0.0393889
R15950 a_216625_n11375.n179 a_216625_n11375.n153 0.0393889
R15951 a_216625_n11375.n13 a_216625_n11375.n6 0.0393889
R15952 a_216625_n11375.n41 a_216625_n11375.n37 0.0393889
R15953 a_216625_n11375.n57 a_216625_n11375.n36 0.0393889
R15954 a_216625_n11375.n73 a_216625_n11375.n35 0.0393889
R15955 a_216625_n11375.n69 a_216625_n11375.n53 0.0388421
R15956 a_216625_n11375.n33 a_216625_n11375.n32 0.0366111
R15957 a_219526_n14006.n368 a_219526_n14006.n367 585
R15958 a_219526_n14006.n368 a_219526_n14006.n95 585
R15959 a_219526_n14006.n368 a_219526_n14006.n94 585
R15960 a_219526_n14006.n368 a_219526_n14006.n93 585
R15961 a_219526_n14006.n368 a_219526_n14006.n92 585
R15962 a_219526_n14006.n368 a_219526_n14006.n91 585
R15963 a_219526_n14006.n368 a_219526_n14006.n89 585
R15964 a_219526_n14006.n368 a_219526_n14006.n88 585
R15965 a_219526_n14006.n368 a_219526_n14006.n87 585
R15966 a_219526_n14006.n368 a_219526_n14006.n82 585
R15967 a_219526_n14006.n368 a_219526_n14006.n81 585
R15968 a_219526_n14006.n369 a_219526_n14006.n368 585
R15969 a_219526_n14006.n306 a_219526_n14006.n305 585
R15970 a_219526_n14006.n306 a_219526_n14006.n118 585
R15971 a_219526_n14006.n306 a_219526_n14006.n117 585
R15972 a_219526_n14006.n306 a_219526_n14006.n116 585
R15973 a_219526_n14006.n306 a_219526_n14006.n115 585
R15974 a_219526_n14006.n306 a_219526_n14006.n114 585
R15975 a_219526_n14006.n306 a_219526_n14006.n112 585
R15976 a_219526_n14006.n306 a_219526_n14006.n111 585
R15977 a_219526_n14006.n306 a_219526_n14006.n110 585
R15978 a_219526_n14006.n306 a_219526_n14006.n109 585
R15979 a_219526_n14006.n306 a_219526_n14006.n108 585
R15980 a_219526_n14006.n307 a_219526_n14006.n306 585
R15981 a_219526_n14006.n380 a_219526_n14006.n374 585
R15982 a_219526_n14006.n380 a_219526_n14006.n17 291.382
R15983 a_219526_n14006.n66 a_219526_n14006.n60 585
R15984 a_219526_n14006.n66 a_219526_n14006.n20 291.382
R15985 a_219526_n14006.n197 a_219526_n14006.n191 585
R15986 a_219526_n14006.n197 a_219526_n14006.n22 291.382
R15987 a_219526_n14006.n205 a_219526_n14006.n199 585
R15988 a_219526_n14006.n205 a_219526_n14006.n24 291.382
R15989 a_219526_n14006.n213 a_219526_n14006.n207 585
R15990 a_219526_n14006.n213 a_219526_n14006.n26 291.382
R15991 a_219526_n14006.n221 a_219526_n14006.n215 585
R15992 a_219526_n14006.n221 a_219526_n14006.n28 291.382
R15993 a_219526_n14006.n173 a_219526_n14006.n172 585
R15994 a_219526_n14006.n170 a_219526_n14006.n169 585
R15995 a_219526_n14006.n179 a_219526_n14006.n178 585
R15996 a_219526_n14006.n181 a_219526_n14006.n180 585
R15997 a_219526_n14006.n168 a_219526_n14006.n167 585
R15998 a_219526_n14006.n281 a_219526_n14006.n280 585
R15999 a_219526_n14006.n281 a_219526_n14006.n236 585
R16000 a_219526_n14006.n281 a_219526_n14006.n235 585
R16001 a_219526_n14006.n281 a_219526_n14006.n234 585
R16002 a_219526_n14006.n281 a_219526_n14006.n233 585
R16003 a_219526_n14006.n281 a_219526_n14006.n232 585
R16004 a_219526_n14006.n281 a_219526_n14006.n230 585
R16005 a_219526_n14006.n281 a_219526_n14006.n229 585
R16006 a_219526_n14006.n281 a_219526_n14006.n223 585
R16007 a_219526_n14006.n282 a_219526_n14006.n281 585
R16008 a_219526_n14006.n281 a_219526_n14006.n227 585
R16009 a_219526_n14006.n281 a_219526_n14006.n225 585
R16010 a_219526_n14006.n408 a_219526_n14006.n45 585
R16011 a_219526_n14006.n408 a_219526_n14006.n46 585
R16012 a_219526_n14006.n408 a_219526_n14006.n44 585
R16013 a_219526_n14006.n408 a_219526_n14006.n47 585
R16014 a_219526_n14006.n408 a_219526_n14006.n43 585
R16015 a_219526_n14006.n408 a_219526_n14006.n48 585
R16016 a_219526_n14006.n408 a_219526_n14006.n41 585
R16017 a_219526_n14006.n408 a_219526_n14006.n49 585
R16018 a_219526_n14006.n408 a_219526_n14006.n40 585
R16019 a_219526_n14006.n408 a_219526_n14006.n50 585
R16020 a_219526_n14006.n408 a_219526_n14006.n39 585
R16021 a_219526_n14006.n408 a_219526_n14006.n407 585
R16022 a_219526_n14006.n310 a_219526_n14006.t20 433.543
R16023 a_219526_n14006.n343 a_219526_n14006.t2 433.543
R16024 a_219526_n14006.n312 a_219526_n14006.t20 433.351
R16025 a_219526_n14006.n249 a_219526_n14006.t34 433.149
R16026 a_219526_n14006.t24 a_219526_n14006.n346 433.149
R16027 a_219526_n14006.n347 a_219526_n14006.t24 433.149
R16028 a_219526_n14006.t40 a_219526_n14006.n51 433.149
R16029 a_219526_n14006.n54 a_219526_n14006.t40 433.149
R16030 a_219526_n14006.n314 a_219526_n14006.t61 433.149
R16031 a_219526_n14006.t61 a_219526_n14006.n313 433.149
R16032 a_219526_n14006.n311 a_219526_n14006.t16 433.149
R16033 a_219526_n14006.t16 a_219526_n14006.n310 433.149
R16034 a_219526_n14006.t30 a_219526_n14006.n260 433.149
R16035 a_219526_n14006.n261 a_219526_n14006.t30 433.149
R16036 a_219526_n14006.t36 a_219526_n14006.n107 433.149
R16037 a_219526_n14006.n238 a_219526_n14006.t36 433.149
R16038 a_219526_n14006.n251 a_219526_n14006.t38 433.149
R16039 a_219526_n14006.t38 a_219526_n14006.n250 433.149
R16040 a_219526_n14006.n252 a_219526_n14006.t4 433.149
R16041 a_219526_n14006.t4 a_219526_n14006.n241 433.149
R16042 a_219526_n14006.t10 a_219526_n14006.n253 433.149
R16043 a_219526_n14006.n254 a_219526_n14006.t10 433.149
R16044 a_219526_n14006.t28 a_219526_n14006.n240 433.149
R16045 a_219526_n14006.n255 a_219526_n14006.t28 433.149
R16046 a_219526_n14006.n257 a_219526_n14006.t32 433.149
R16047 a_219526_n14006.t32 a_219526_n14006.n256 433.149
R16048 a_219526_n14006.n258 a_219526_n14006.t26 433.149
R16049 a_219526_n14006.t26 a_219526_n14006.n237 433.149
R16050 a_219526_n14006.n404 a_219526_n14006.t6 433.149
R16051 a_219526_n14006.t6 a_219526_n14006.n403 433.149
R16052 a_219526_n14006.t12 a_219526_n14006.n52 433.149
R16053 a_219526_n14006.n53 a_219526_n14006.t12 433.149
R16054 a_219526_n14006.n245 a_219526_n14006.t18 433.149
R16055 a_219526_n14006.t18 a_219526_n14006.n244 433.149
R16056 a_219526_n14006.n246 a_219526_n14006.t22 433.149
R16057 a_219526_n14006.t22 a_219526_n14006.n243 433.149
R16058 a_219526_n14006.t0 a_219526_n14006.n247 433.149
R16059 a_219526_n14006.n248 a_219526_n14006.t0 433.149
R16060 a_219526_n14006.n327 a_219526_n14006.t52 433.149
R16061 a_219526_n14006.t52 a_219526_n14006.n100 433.149
R16062 a_219526_n14006.n339 a_219526_n14006.t62 433.149
R16063 a_219526_n14006.t62 a_219526_n14006.n96 433.149
R16064 a_219526_n14006.n338 a_219526_n14006.t57 433.149
R16065 a_219526_n14006.t57 a_219526_n14006.n337 433.149
R16066 a_219526_n14006.t49 a_219526_n14006.n97 433.149
R16067 a_219526_n14006.n336 a_219526_n14006.t49 433.149
R16068 a_219526_n14006.t66 a_219526_n14006.n334 433.149
R16069 a_219526_n14006.n335 a_219526_n14006.t66 433.149
R16070 a_219526_n14006.n333 a_219526_n14006.t63 433.149
R16071 a_219526_n14006.t63 a_219526_n14006.n98 433.149
R16072 a_219526_n14006.n332 a_219526_n14006.t60 433.149
R16073 a_219526_n14006.t60 a_219526_n14006.n331 433.149
R16074 a_219526_n14006.t58 a_219526_n14006.n99 433.149
R16075 a_219526_n14006.n330 a_219526_n14006.t58 433.149
R16076 a_219526_n14006.t69 a_219526_n14006.n328 433.149
R16077 a_219526_n14006.n329 a_219526_n14006.t69 433.149
R16078 a_219526_n14006.n326 a_219526_n14006.t50 433.149
R16079 a_219526_n14006.t50 a_219526_n14006.n325 433.149
R16080 a_219526_n14006.t67 a_219526_n14006.n101 433.149
R16081 a_219526_n14006.n324 a_219526_n14006.t67 433.149
R16082 a_219526_n14006.t64 a_219526_n14006.n322 433.149
R16083 a_219526_n14006.n323 a_219526_n14006.t64 433.149
R16084 a_219526_n14006.n321 a_219526_n14006.t55 433.149
R16085 a_219526_n14006.t55 a_219526_n14006.n102 433.149
R16086 a_219526_n14006.n320 a_219526_n14006.t53 433.149
R16087 a_219526_n14006.t53 a_219526_n14006.n319 433.149
R16088 a_219526_n14006.t56 a_219526_n14006.n103 433.149
R16089 a_219526_n14006.n318 a_219526_n14006.t56 433.149
R16090 a_219526_n14006.t54 a_219526_n14006.n316 433.149
R16091 a_219526_n14006.n317 a_219526_n14006.t54 433.149
R16092 a_219526_n14006.n315 a_219526_n14006.t51 433.149
R16093 a_219526_n14006.t51 a_219526_n14006.n104 433.149
R16094 a_219526_n14006.t34 a_219526_n14006.n242 433.149
R16095 a_219526_n14006.n340 a_219526_n14006.t65 433.149
R16096 a_219526_n14006.n342 a_219526_n14006.t65 433.149
R16097 a_219526_n14006.n38 a_219526_n14006.t2 433.149
R16098 a_219526_n14006.n345 a_219526_n14006.t14 433.149
R16099 a_219526_n14006.t14 a_219526_n14006.n344 433.149
R16100 a_219526_n14006.n343 a_219526_n14006.t8 433.149
R16101 a_219526_n14006.t8 a_219526_n14006.n38 433.149
R16102 a_219526_n14006.t21 a_219526_n14006.n171 384.339
R16103 a_219526_n14006.n368 a_219526_n14006.n90 286.238
R16104 a_219526_n14006.n306 a_219526_n14006.n113 286.238
R16105 a_219526_n14006.n281 a_219526_n14006.n231 286.238
R16106 a_219526_n14006.n408 a_219526_n14006.n42 286.238
R16107 a_219526_n14006.n172 a_219526_n14006.n169 230.966
R16108 a_219526_n14006.n179 a_219526_n14006.n169 230.966
R16109 a_219526_n14006.n180 a_219526_n14006.n179 230.966
R16110 a_219526_n14006.n180 a_219526_n14006.n167 230.966
R16111 a_219526_n14006.n30 a_219526_n14006.n167 570.105
R16112 a_219526_n14006.n105 a_219526_n14006.t59 215.964
R16113 a_219526_n14006.n341 a_219526_n14006.t68 215.963
R16114 a_219526_n14006.n78 a_219526_n14006.n70 185
R16115 a_219526_n14006.n78 a_219526_n14006.n69 185
R16116 a_219526_n14006.n78 a_219526_n14006.n7 91.4184
R16117 a_219526_n14006.n135 a_219526_n14006.n127 185
R16118 a_219526_n14006.n135 a_219526_n14006.n126 185
R16119 a_219526_n14006.n135 a_219526_n14006.n9 91.4184
R16120 a_219526_n14006.n145 a_219526_n14006.n137 185
R16121 a_219526_n14006.n145 a_219526_n14006.n136 185
R16122 a_219526_n14006.n145 a_219526_n14006.n11 91.4184
R16123 a_219526_n14006.n154 a_219526_n14006.n153 185
R16124 a_219526_n14006.n151 a_219526_n14006.n150 185
R16125 a_219526_n14006.n159 a_219526_n14006.n158 185
R16126 a_219526_n14006.n161 a_219526_n14006.n160 185
R16127 a_219526_n14006.n147 a_219526_n14006.n146 185
R16128 a_219526_n14006.t47 a_219526_n14006.n152 174.857
R16129 a_219526_n14006.n153 a_219526_n14006.n150 140.69
R16130 a_219526_n14006.n159 a_219526_n14006.n150 140.69
R16131 a_219526_n14006.n160 a_219526_n14006.n159 140.69
R16132 a_219526_n14006.n160 a_219526_n14006.n146 140.69
R16133 a_219526_n14006.n13 a_219526_n14006.n146 256.962
R16134 a_219526_n14006.n172 a_219526_n14006.t21 115.484
R16135 a_219526_n14006.n153 a_219526_n14006.t47 70.3453
R16136 a_219526_n14006.n380 a_219526_n14006.n379 51.6891
R16137 a_219526_n14006.n66 a_219526_n14006.n65 51.6891
R16138 a_219526_n14006.n197 a_219526_n14006.n196 51.6891
R16139 a_219526_n14006.n205 a_219526_n14006.n204 51.6891
R16140 a_219526_n14006.n213 a_219526_n14006.n212 51.6891
R16141 a_219526_n14006.n221 a_219526_n14006.n220 51.6891
R16142 a_219526_n14006.n379 a_219526_n14006.n378 29.8062
R16143 a_219526_n14006.n65 a_219526_n14006.n64 29.8062
R16144 a_219526_n14006.n196 a_219526_n14006.n195 29.8062
R16145 a_219526_n14006.n204 a_219526_n14006.n203 29.8062
R16146 a_219526_n14006.n212 a_219526_n14006.n211 29.8062
R16147 a_219526_n14006.n220 a_219526_n14006.n219 29.8062
R16148 a_219526_n14006.n173 a_219526_n14006.n171 29.3167
R16149 a_219526_n14006.n154 a_219526_n14006.n152 28.4333
R16150 a_219526_n14006.n77 a_219526_n14006.n76 26.8423
R16151 a_219526_n14006.n134 a_219526_n14006.n133 26.8423
R16152 a_219526_n14006.n144 a_219526_n14006.n143 26.8423
R16153 a_219526_n14006.n355 a_219526_n14006.n91 24.8476
R16154 a_219526_n14006.n353 a_219526_n14006.n89 24.8476
R16155 a_219526_n14006.n293 a_219526_n14006.n114 24.8476
R16156 a_219526_n14006.n291 a_219526_n14006.n112 24.8476
R16157 a_219526_n14006.n155 a_219526_n14006.n151 24.8476
R16158 a_219526_n14006.n174 a_219526_n14006.n170 24.8476
R16159 a_219526_n14006.n268 a_219526_n14006.n232 24.8476
R16160 a_219526_n14006.n266 a_219526_n14006.n230 24.8476
R16161 a_219526_n14006.n389 a_219526_n14006.n48 24.8476
R16162 a_219526_n14006.n387 a_219526_n14006.n41 24.8476
R16163 a_219526_n14006.n357 a_219526_n14006.n92 23.3417
R16164 a_219526_n14006.n351 a_219526_n14006.n88 23.3417
R16165 a_219526_n14006.n295 a_219526_n14006.n115 23.3417
R16166 a_219526_n14006.n289 a_219526_n14006.n111 23.3417
R16167 a_219526_n14006.n158 a_219526_n14006.n157 23.3417
R16168 a_219526_n14006.n178 a_219526_n14006.n177 23.3417
R16169 a_219526_n14006.n270 a_219526_n14006.n233 23.3417
R16170 a_219526_n14006.n264 a_219526_n14006.n229 23.3417
R16171 a_219526_n14006.n391 a_219526_n14006.n43 23.3417
R16172 a_219526_n14006.n385 a_219526_n14006.n49 23.3417
R16173 a_219526_n14006.n359 a_219526_n14006.n93 21.8358
R16174 a_219526_n14006.n350 a_219526_n14006.n87 21.8358
R16175 a_219526_n14006.n297 a_219526_n14006.n116 21.8358
R16176 a_219526_n14006.n288 a_219526_n14006.n110 21.8358
R16177 a_219526_n14006.n76 a_219526_n14006.n70 21.8358
R16178 a_219526_n14006.n133 a_219526_n14006.n127 21.8358
R16179 a_219526_n14006.n143 a_219526_n14006.n137 21.8358
R16180 a_219526_n14006.n161 a_219526_n14006.n149 21.8358
R16181 a_219526_n14006.n181 a_219526_n14006.n0 21.8358
R16182 a_219526_n14006.n272 a_219526_n14006.n234 21.8358
R16183 a_219526_n14006.n228 a_219526_n14006.n223 21.8358
R16184 a_219526_n14006.n393 a_219526_n14006.n47 21.8358
R16185 a_219526_n14006.n384 a_219526_n14006.n40 21.8358
R16186 a_219526_n14006.n361 a_219526_n14006.n94 20.3299
R16187 a_219526_n14006.n86 a_219526_n14006.n82 20.3299
R16188 a_219526_n14006.n299 a_219526_n14006.n117 20.3299
R16189 a_219526_n14006.n122 a_219526_n14006.n109 20.3299
R16190 a_219526_n14006.n378 a_219526_n14006.n374 20.3299
R16191 a_219526_n14006.n73 a_219526_n14006.n69 20.3299
R16192 a_219526_n14006.n130 a_219526_n14006.n126 20.3299
R16193 a_219526_n14006.n140 a_219526_n14006.n136 20.3299
R16194 a_219526_n14006.n162 a_219526_n14006.n147 20.3299
R16195 a_219526_n14006.n64 a_219526_n14006.n60 20.3299
R16196 a_219526_n14006.n195 a_219526_n14006.n191 20.3299
R16197 a_219526_n14006.n203 a_219526_n14006.n199 20.3299
R16198 a_219526_n14006.n211 a_219526_n14006.n207 20.3299
R16199 a_219526_n14006.n219 a_219526_n14006.n215 20.3299
R16200 a_219526_n14006.n182 a_219526_n14006.n168 20.3299
R16201 a_219526_n14006.n274 a_219526_n14006.n235 20.3299
R16202 a_219526_n14006.n283 a_219526_n14006.n282 20.3299
R16203 a_219526_n14006.n395 a_219526_n14006.n44 20.3299
R16204 a_219526_n14006.n57 a_219526_n14006.n50 20.3299
R16205 a_219526_n14006.n367 a_219526_n14006.n349 19.0887
R16206 a_219526_n14006.n370 a_219526_n14006.n369 19.0887
R16207 a_219526_n14006.n305 a_219526_n14006.n119 19.0887
R16208 a_219526_n14006.n308 a_219526_n14006.n307 19.0887
R16209 a_219526_n14006.n280 a_219526_n14006.n263 19.0887
R16210 a_219526_n14006.n239 a_219526_n14006.n225 19.0887
R16211 a_219526_n14006.n401 a_219526_n14006.n45 19.0887
R16212 a_219526_n14006.n407 a_219526_n14006.n406 19.0887
R16213 a_219526_n14006.n363 a_219526_n14006.n95 18.824
R16214 a_219526_n14006.n83 a_219526_n14006.n81 18.824
R16215 a_219526_n14006.n301 a_219526_n14006.n118 18.824
R16216 a_219526_n14006.n120 a_219526_n14006.n108 18.824
R16217 a_219526_n14006.n375 a_219526_n14006.n17 24.6305
R16218 a_219526_n14006.n71 a_219526_n14006.n7 24.4363
R16219 a_219526_n14006.n128 a_219526_n14006.n9 24.4363
R16220 a_219526_n14006.n138 a_219526_n14006.n11 24.4363
R16221 a_219526_n14006.n13 a_219526_n14006.n165 22.9459
R16222 a_219526_n14006.n61 a_219526_n14006.n20 24.6305
R16223 a_219526_n14006.n192 a_219526_n14006.n22 24.6305
R16224 a_219526_n14006.n200 a_219526_n14006.n24 24.6305
R16225 a_219526_n14006.n208 a_219526_n14006.n26 24.6305
R16226 a_219526_n14006.n216 a_219526_n14006.n28 24.6305
R16227 a_219526_n14006.n30 a_219526_n14006.n185 23.6861
R16228 a_219526_n14006.n276 a_219526_n14006.n236 18.824
R16229 a_219526_n14006.n227 a_219526_n14006.n224 18.824
R16230 a_219526_n14006.n397 a_219526_n14006.n46 18.824
R16231 a_219526_n14006.n55 a_219526_n14006.n39 18.824
R16232 a_219526_n14006.n367 a_219526_n14006.n366 17.3181
R16233 a_219526_n14006.n369 a_219526_n14006.n80 17.3181
R16234 a_219526_n14006.n305 a_219526_n14006.n304 17.3181
R16235 a_219526_n14006.n307 a_219526_n14006.n33 17.3181
R16236 a_219526_n14006.n17 a_219526_n14006.n16 9.772
R16237 a_219526_n14006.n7 a_219526_n14006.n6 9.72509
R16238 a_219526_n14006.n9 a_219526_n14006.n8 9.72509
R16239 a_219526_n14006.n11 a_219526_n14006.n10 9.72509
R16240 a_219526_n14006.n13 a_219526_n14006.n12 11.3106
R16241 a_219526_n14006.n20 a_219526_n14006.n19 9.772
R16242 a_219526_n14006.n22 a_219526_n14006.n21 9.772
R16243 a_219526_n14006.n24 a_219526_n14006.n23 9.772
R16244 a_219526_n14006.n26 a_219526_n14006.n25 9.772
R16245 a_219526_n14006.n28 a_219526_n14006.n27 9.772
R16246 a_219526_n14006.n30 a_219526_n14006.n29 10.7354
R16247 a_219526_n14006.n280 a_219526_n14006.n279 17.3181
R16248 a_219526_n14006.n226 a_219526_n14006.n225 17.3181
R16249 a_219526_n14006.n399 a_219526_n14006.n45 17.3181
R16250 a_219526_n14006.n407 a_219526_n14006.n36 17.3181
R16251 a_219526_n14006.n78 a_219526_n14006.n77 16.7813
R16252 a_219526_n14006.n135 a_219526_n14006.n134 16.7813
R16253 a_219526_n14006.n145 a_219526_n14006.n144 16.7813
R16254 a_219526_n14006.n355 a_219526_n14006.n90 13.2799
R16255 a_219526_n14006.n353 a_219526_n14006.n90 13.2799
R16256 a_219526_n14006.n293 a_219526_n14006.n113 13.2799
R16257 a_219526_n14006.n291 a_219526_n14006.n113 13.2799
R16258 a_219526_n14006.n268 a_219526_n14006.n231 13.2799
R16259 a_219526_n14006.n266 a_219526_n14006.n231 13.2799
R16260 a_219526_n14006.n389 a_219526_n14006.n42 13.2799
R16261 a_219526_n14006.n387 a_219526_n14006.n42 13.2799
R16262 a_219526_n14006.n378 a_219526_n14006.n377 9.3005
R16263 a_219526_n14006.n376 a_219526_n14006.n375 9.3005
R16264 a_219526_n14006.n76 a_219526_n14006.n75 9.3005
R16265 a_219526_n14006.n74 a_219526_n14006.n73 9.3005
R16266 a_219526_n14006.n72 a_219526_n14006.n71 9.3005
R16267 a_219526_n14006.n133 a_219526_n14006.n132 9.3005
R16268 a_219526_n14006.n131 a_219526_n14006.n130 9.3005
R16269 a_219526_n14006.n129 a_219526_n14006.n128 9.3005
R16270 a_219526_n14006.n143 a_219526_n14006.n142 9.3005
R16271 a_219526_n14006.n141 a_219526_n14006.n140 9.3005
R16272 a_219526_n14006.n139 a_219526_n14006.n138 9.3005
R16273 a_219526_n14006.n156 a_219526_n14006.n155 9.3005
R16274 a_219526_n14006.n149 a_219526_n14006.n148 9.3005
R16275 a_219526_n14006.n163 a_219526_n14006.n162 9.3005
R16276 a_219526_n14006.n165 a_219526_n14006.n164 9.3005
R16277 a_219526_n14006.n157 a_219526_n14006.n18 9.3005
R16278 a_219526_n14006.n64 a_219526_n14006.n63 9.3005
R16279 a_219526_n14006.n62 a_219526_n14006.n61 9.3005
R16280 a_219526_n14006.n195 a_219526_n14006.n194 9.3005
R16281 a_219526_n14006.n193 a_219526_n14006.n192 9.3005
R16282 a_219526_n14006.n203 a_219526_n14006.n202 9.3005
R16283 a_219526_n14006.n201 a_219526_n14006.n200 9.3005
R16284 a_219526_n14006.n211 a_219526_n14006.n210 9.3005
R16285 a_219526_n14006.n209 a_219526_n14006.n208 9.3005
R16286 a_219526_n14006.n219 a_219526_n14006.n218 9.3005
R16287 a_219526_n14006.n217 a_219526_n14006.n216 9.3005
R16288 a_219526_n14006.n175 a_219526_n14006.n174 9.3005
R16289 a_219526_n14006.n177 a_219526_n14006.n176 9.3005
R16290 a_219526_n14006.n183 a_219526_n14006.n182 9.3005
R16291 a_219526_n14006.n185 a_219526_n14006.n184 9.3005
R16292 a_219526_n14006.n1 a_219526_n14006.n0 9.3005
R16293 a_219526_n14006.n269 a_219526_n14006.n268 9.3005
R16294 a_219526_n14006.n271 a_219526_n14006.n270 9.3005
R16295 a_219526_n14006.n273 a_219526_n14006.n272 9.3005
R16296 a_219526_n14006.n275 a_219526_n14006.n274 9.3005
R16297 a_219526_n14006.n277 a_219526_n14006.n276 9.3005
R16298 a_219526_n14006.n279 a_219526_n14006.n278 9.3005
R16299 a_219526_n14006.n267 a_219526_n14006.n266 9.3005
R16300 a_219526_n14006.n265 a_219526_n14006.n264 9.3005
R16301 a_219526_n14006.n228 a_219526_n14006.n2 9.3005
R16302 a_219526_n14006.n284 a_219526_n14006.n283 9.3005
R16303 a_219526_n14006.n224 a_219526_n14006.n31 9.3005
R16304 a_219526_n14006.n226 a_219526_n14006.n32 9.3005
R16305 a_219526_n14006.n34 a_219526_n14006.n33 9.3005
R16306 a_219526_n14006.n123 a_219526_n14006.n122 9.3005
R16307 a_219526_n14006.n121 a_219526_n14006.n120 9.3005
R16308 a_219526_n14006.n3 a_219526_n14006.n288 9.3005
R16309 a_219526_n14006.n294 a_219526_n14006.n293 9.3005
R16310 a_219526_n14006.n296 a_219526_n14006.n295 9.3005
R16311 a_219526_n14006.n298 a_219526_n14006.n297 9.3005
R16312 a_219526_n14006.n300 a_219526_n14006.n299 9.3005
R16313 a_219526_n14006.n302 a_219526_n14006.n301 9.3005
R16314 a_219526_n14006.n304 a_219526_n14006.n303 9.3005
R16315 a_219526_n14006.n292 a_219526_n14006.n291 9.3005
R16316 a_219526_n14006.n290 a_219526_n14006.n289 9.3005
R16317 a_219526_n14006.n356 a_219526_n14006.n355 9.3005
R16318 a_219526_n14006.n358 a_219526_n14006.n357 9.3005
R16319 a_219526_n14006.n360 a_219526_n14006.n359 9.3005
R16320 a_219526_n14006.n362 a_219526_n14006.n361 9.3005
R16321 a_219526_n14006.n364 a_219526_n14006.n363 9.3005
R16322 a_219526_n14006.n366 a_219526_n14006.n365 9.3005
R16323 a_219526_n14006.n354 a_219526_n14006.n353 9.3005
R16324 a_219526_n14006.n352 a_219526_n14006.n351 9.3005
R16325 a_219526_n14006.n4 a_219526_n14006.n350 9.3005
R16326 a_219526_n14006.n86 a_219526_n14006.n85 9.3005
R16327 a_219526_n14006.n84 a_219526_n14006.n83 9.3005
R16328 a_219526_n14006.n80 a_219526_n14006.n35 9.3005
R16329 a_219526_n14006.n390 a_219526_n14006.n389 9.3005
R16330 a_219526_n14006.n392 a_219526_n14006.n391 9.3005
R16331 a_219526_n14006.n394 a_219526_n14006.n393 9.3005
R16332 a_219526_n14006.n396 a_219526_n14006.n395 9.3005
R16333 a_219526_n14006.n398 a_219526_n14006.n397 9.3005
R16334 a_219526_n14006.n400 a_219526_n14006.n399 9.3005
R16335 a_219526_n14006.n388 a_219526_n14006.n387 9.3005
R16336 a_219526_n14006.n386 a_219526_n14006.n385 9.3005
R16337 a_219526_n14006.n5 a_219526_n14006.n384 9.3005
R16338 a_219526_n14006.n58 a_219526_n14006.n57 9.3005
R16339 a_219526_n14006.n56 a_219526_n14006.n55 9.3005
R16340 a_219526_n14006.n37 a_219526_n14006.n36 9.3005
R16341 a_219526_n14006.n366 a_219526_n14006.n95 8.28285
R16342 a_219526_n14006.n81 a_219526_n14006.n80 8.28285
R16343 a_219526_n14006.n304 a_219526_n14006.n118 8.28285
R16344 a_219526_n14006.n108 a_219526_n14006.n33 8.28285
R16345 a_219526_n14006.n279 a_219526_n14006.n236 8.28285
R16346 a_219526_n14006.n227 a_219526_n14006.n226 8.28285
R16347 a_219526_n14006.n399 a_219526_n14006.n46 8.28285
R16348 a_219526_n14006.n36 a_219526_n14006.n39 8.28285
R16349 a_219526_n14006.n381 a_219526_n14006.n373 7.9105
R16350 a_219526_n14006.n14 a_219526_n14006.n68 7.9105
R16351 a_219526_n14006.n14 a_219526_n14006.n125 7.9105
R16352 a_219526_n14006.n15 a_219526_n14006.n124 7.9105
R16353 a_219526_n14006.n15 a_219526_n14006.n18 7.9105
R16354 a_219526_n14006.n15 a_219526_n14006.n12 7.9105
R16355 a_219526_n14006.n15 a_219526_n14006.n10 7.9105
R16356 a_219526_n14006.n14 a_219526_n14006.n8 7.9105
R16357 a_219526_n14006.n14 a_219526_n14006.n6 7.9105
R16358 a_219526_n14006.n67 a_219526_n14006.n59 7.9105
R16359 a_219526_n14006.n198 a_219526_n14006.n190 7.9105
R16360 a_219526_n14006.n206 a_219526_n14006.n189 7.9105
R16361 a_219526_n14006.n214 a_219526_n14006.n188 7.9105
R16362 a_219526_n14006.n222 a_219526_n14006.n187 7.9105
R16363 a_219526_n14006.n186 a_219526_n14006.n1 7.9105
R16364 a_219526_n14006.n186 a_219526_n14006.n29 7.9105
R16365 a_219526_n14006.n222 a_219526_n14006.n27 7.9105
R16366 a_219526_n14006.n214 a_219526_n14006.n25 7.9105
R16367 a_219526_n14006.n206 a_219526_n14006.n23 7.9105
R16368 a_219526_n14006.n198 a_219526_n14006.n21 7.9105
R16369 a_219526_n14006.n67 a_219526_n14006.n19 7.9105
R16370 a_219526_n14006.n381 a_219526_n14006.n16 7.9105
R16371 a_219526_n14006.n285 a_219526_n14006.n2 7.9105
R16372 a_219526_n14006.n285 a_219526_n14006.n32 7.9105
R16373 a_219526_n14006.n383 a_219526_n14006.n37 7.9105
R16374 a_219526_n14006.n5 a_219526_n14006.n383 7.9105
R16375 a_219526_n14006.n363 a_219526_n14006.n94 6.77697
R16376 a_219526_n14006.n83 a_219526_n14006.n82 6.77697
R16377 a_219526_n14006.n301 a_219526_n14006.n117 6.77697
R16378 a_219526_n14006.n120 a_219526_n14006.n109 6.77697
R16379 a_219526_n14006.n375 a_219526_n14006.n374 6.77697
R16380 a_219526_n14006.n71 a_219526_n14006.n69 6.77697
R16381 a_219526_n14006.n128 a_219526_n14006.n126 6.77697
R16382 a_219526_n14006.n138 a_219526_n14006.n136 6.77697
R16383 a_219526_n14006.n165 a_219526_n14006.n147 6.77697
R16384 a_219526_n14006.n61 a_219526_n14006.n60 6.77697
R16385 a_219526_n14006.n192 a_219526_n14006.n191 6.77697
R16386 a_219526_n14006.n200 a_219526_n14006.n199 6.77697
R16387 a_219526_n14006.n208 a_219526_n14006.n207 6.77697
R16388 a_219526_n14006.n216 a_219526_n14006.n215 6.77697
R16389 a_219526_n14006.n185 a_219526_n14006.n168 6.77697
R16390 a_219526_n14006.n276 a_219526_n14006.n235 6.77697
R16391 a_219526_n14006.n282 a_219526_n14006.n224 6.77697
R16392 a_219526_n14006.n397 a_219526_n14006.n44 6.77697
R16393 a_219526_n14006.n55 a_219526_n14006.n50 6.77697
R16394 a_219526_n14006.n368 a_219526_n14006.t25 5.7135
R16395 a_219526_n14006.n368 a_219526_n14006.t15 5.7135
R16396 a_219526_n14006.n306 a_219526_n14006.t17 5.7135
R16397 a_219526_n14006.n306 a_219526_n14006.t37 5.7135
R16398 a_219526_n14006.n380 a_219526_n14006.t9 5.7135
R16399 a_219526_n14006.n380 a_219526_n14006.t3 5.7135
R16400 a_219526_n14006.n66 a_219526_n14006.t19 5.7135
R16401 a_219526_n14006.n66 a_219526_n14006.t13 5.7135
R16402 a_219526_n14006.n197 a_219526_n14006.t1 5.7135
R16403 a_219526_n14006.n197 a_219526_n14006.t23 5.7135
R16404 a_219526_n14006.n205 a_219526_n14006.t39 5.7135
R16405 a_219526_n14006.n205 a_219526_n14006.t35 5.7135
R16406 a_219526_n14006.n213 a_219526_n14006.t11 5.7135
R16407 a_219526_n14006.n213 a_219526_n14006.t5 5.7135
R16408 a_219526_n14006.n221 a_219526_n14006.t33 5.7135
R16409 a_219526_n14006.n221 a_219526_n14006.t29 5.7135
R16410 a_219526_n14006.n281 a_219526_n14006.t31 5.7135
R16411 a_219526_n14006.n281 a_219526_n14006.t27 5.7135
R16412 a_219526_n14006.n408 a_219526_n14006.t7 5.7135
R16413 a_219526_n14006.t41 a_219526_n14006.n408 5.7135
R16414 a_219526_n14006.n156 a_219526_n14006.n152 5.33935
R16415 a_219526_n14006.n361 a_219526_n14006.n93 5.27109
R16416 a_219526_n14006.n87 a_219526_n14006.n86 5.27109
R16417 a_219526_n14006.n299 a_219526_n14006.n116 5.27109
R16418 a_219526_n14006.n122 a_219526_n14006.n110 5.27109
R16419 a_219526_n14006.n73 a_219526_n14006.n70 5.27109
R16420 a_219526_n14006.n130 a_219526_n14006.n127 5.27109
R16421 a_219526_n14006.n140 a_219526_n14006.n137 5.27109
R16422 a_219526_n14006.n162 a_219526_n14006.n161 5.27109
R16423 a_219526_n14006.n182 a_219526_n14006.n181 5.27109
R16424 a_219526_n14006.n274 a_219526_n14006.n234 5.27109
R16425 a_219526_n14006.n283 a_219526_n14006.n223 5.27109
R16426 a_219526_n14006.n395 a_219526_n14006.n47 5.27109
R16427 a_219526_n14006.n57 a_219526_n14006.n40 5.27109
R16428 a_219526_n14006.n372 a_219526_n14006.n4 4.59906
R16429 a_219526_n14006.n3 a_219526_n14006.n287 4.59906
R16430 a_219526_n14006.n166 a_219526_n14006.n15 4.5738
R16431 a_219526_n14006.n371 a_219526_n14006.n14 4.57256
R16432 a_219526_n14006.n175 a_219526_n14006.n171 4.51911
R16433 a_219526_n14006.n166 a_219526_n14006.n34 4.5005
R16434 a_219526_n14006.n371 a_219526_n14006.n35 4.5005
R16435 a_219526_n14006.n359 a_219526_n14006.n92 3.76521
R16436 a_219526_n14006.n350 a_219526_n14006.n88 3.76521
R16437 a_219526_n14006.n297 a_219526_n14006.n115 3.76521
R16438 a_219526_n14006.n288 a_219526_n14006.n111 3.76521
R16439 a_219526_n14006.n158 a_219526_n14006.n149 3.76521
R16440 a_219526_n14006.n178 a_219526_n14006.n0 3.76521
R16441 a_219526_n14006.n272 a_219526_n14006.n233 3.76521
R16442 a_219526_n14006.n229 a_219526_n14006.n228 3.76521
R16443 a_219526_n14006.n393 a_219526_n14006.n43 3.76521
R16444 a_219526_n14006.n384 a_219526_n14006.n49 3.76521
R16445 a_219526_n14006.n77 a_219526_n14006.n68 3.76174
R16446 a_219526_n14006.n134 a_219526_n14006.n125 3.76174
R16447 a_219526_n14006.n144 a_219526_n14006.n124 3.76174
R16448 a_219526_n14006.n78 a_219526_n14006.t43 3.4805
R16449 a_219526_n14006.n78 a_219526_n14006.t48 3.4805
R16450 a_219526_n14006.n135 a_219526_n14006.t42 3.4805
R16451 a_219526_n14006.n135 a_219526_n14006.t44 3.4805
R16452 a_219526_n14006.n145 a_219526_n14006.t46 3.4805
R16453 a_219526_n14006.n145 a_219526_n14006.t45 3.4805
R16454 a_219526_n14006.n379 a_219526_n14006.n373 3.43565
R16455 a_219526_n14006.n65 a_219526_n14006.n59 3.43565
R16456 a_219526_n14006.n196 a_219526_n14006.n190 3.43565
R16457 a_219526_n14006.n204 a_219526_n14006.n189 3.43565
R16458 a_219526_n14006.n212 a_219526_n14006.n188 3.43565
R16459 a_219526_n14006.n220 a_219526_n14006.n187 3.43565
R16460 a_219526_n14006.n357 a_219526_n14006.n91 2.25932
R16461 a_219526_n14006.n351 a_219526_n14006.n89 2.25932
R16462 a_219526_n14006.n295 a_219526_n14006.n114 2.25932
R16463 a_219526_n14006.n289 a_219526_n14006.n112 2.25932
R16464 a_219526_n14006.n157 a_219526_n14006.n151 2.25932
R16465 a_219526_n14006.n177 a_219526_n14006.n170 2.25932
R16466 a_219526_n14006.n270 a_219526_n14006.n232 2.25932
R16467 a_219526_n14006.n264 a_219526_n14006.n230 2.25932
R16468 a_219526_n14006.n391 a_219526_n14006.n48 2.25932
R16469 a_219526_n14006.n385 a_219526_n14006.n41 2.25932
R16470 a_219526_n14006.n287 a_219526_n14006.n286 1.65697
R16471 a_219526_n14006.n382 a_219526_n14006.n372 1.65697
R16472 a_219526_n14006.n341 a_219526_n14006.n340 1.62034
R16473 a_219526_n14006.n314 a_219526_n14006.n105 1.61786
R16474 a_219526_n14006.n342 a_219526_n14006.n341 1.22534
R16475 a_219526_n14006.n313 a_219526_n14006.n105 1.22286
R16476 a_219526_n14006.n155 a_219526_n14006.n154 0.753441
R16477 a_219526_n14006.n174 a_219526_n14006.n173 0.753441
R16478 a_219526_n14006.n248 a_219526_n14006.n243 0.3955
R16479 a_219526_n14006.n244 a_219526_n14006.n243 0.3955
R16480 a_219526_n14006.n244 a_219526_n14006.n53 0.3955
R16481 a_219526_n14006.n403 a_219526_n14006.n53 0.3955
R16482 a_219526_n14006.n317 a_219526_n14006.n104 0.3955
R16483 a_219526_n14006.n318 a_219526_n14006.n317 0.3955
R16484 a_219526_n14006.n319 a_219526_n14006.n318 0.3955
R16485 a_219526_n14006.n319 a_219526_n14006.n102 0.3955
R16486 a_219526_n14006.n323 a_219526_n14006.n102 0.3955
R16487 a_219526_n14006.n324 a_219526_n14006.n323 0.3955
R16488 a_219526_n14006.n325 a_219526_n14006.n324 0.3955
R16489 a_219526_n14006.n330 a_219526_n14006.n329 0.3955
R16490 a_219526_n14006.n331 a_219526_n14006.n330 0.3955
R16491 a_219526_n14006.n331 a_219526_n14006.n98 0.3955
R16492 a_219526_n14006.n335 a_219526_n14006.n98 0.3955
R16493 a_219526_n14006.n336 a_219526_n14006.n335 0.3955
R16494 a_219526_n14006.n337 a_219526_n14006.n336 0.3955
R16495 a_219526_n14006.n337 a_219526_n14006.n96 0.3955
R16496 a_219526_n14006.n256 a_219526_n14006.n237 0.3955
R16497 a_219526_n14006.n256 a_219526_n14006.n255 0.3955
R16498 a_219526_n14006.n255 a_219526_n14006.n254 0.3955
R16499 a_219526_n14006.n254 a_219526_n14006.n241 0.3955
R16500 a_219526_n14006.n250 a_219526_n14006.n241 0.3955
R16501 a_219526_n14006.n261 a_219526_n14006.n238 0.3955
R16502 a_219526_n14006.n260 a_219526_n14006.n107 0.3955
R16503 a_219526_n14006.n315 a_219526_n14006.n314 0.3955
R16504 a_219526_n14006.n316 a_219526_n14006.n315 0.3955
R16505 a_219526_n14006.n316 a_219526_n14006.n103 0.3955
R16506 a_219526_n14006.n320 a_219526_n14006.n103 0.3955
R16507 a_219526_n14006.n321 a_219526_n14006.n320 0.3955
R16508 a_219526_n14006.n322 a_219526_n14006.n321 0.3955
R16509 a_219526_n14006.n322 a_219526_n14006.n101 0.3955
R16510 a_219526_n14006.n326 a_219526_n14006.n101 0.3955
R16511 a_219526_n14006.n327 a_219526_n14006.n326 0.3955
R16512 a_219526_n14006.n328 a_219526_n14006.n327 0.3955
R16513 a_219526_n14006.n328 a_219526_n14006.n99 0.3955
R16514 a_219526_n14006.n332 a_219526_n14006.n99 0.3955
R16515 a_219526_n14006.n333 a_219526_n14006.n332 0.3955
R16516 a_219526_n14006.n334 a_219526_n14006.n333 0.3955
R16517 a_219526_n14006.n334 a_219526_n14006.n97 0.3955
R16518 a_219526_n14006.n338 a_219526_n14006.n97 0.3955
R16519 a_219526_n14006.n339 a_219526_n14006.n338 0.3955
R16520 a_219526_n14006.n340 a_219526_n14006.n339 0.3955
R16521 a_219526_n14006.n344 a_219526_n14006.n343 0.3955
R16522 a_219526_n14006.n347 a_219526_n14006.n54 0.3955
R16523 a_219526_n14006.n346 a_219526_n14006.n51 0.3955
R16524 a_219526_n14006.n258 a_219526_n14006.n257 0.3955
R16525 a_219526_n14006.n257 a_219526_n14006.n240 0.3955
R16526 a_219526_n14006.n253 a_219526_n14006.n240 0.3955
R16527 a_219526_n14006.n253 a_219526_n14006.n252 0.3955
R16528 a_219526_n14006.n252 a_219526_n14006.n251 0.3955
R16529 a_219526_n14006.n251 a_219526_n14006.n242 0.3955
R16530 a_219526_n14006.n247 a_219526_n14006.n242 0.3955
R16531 a_219526_n14006.n247 a_219526_n14006.n246 0.3955
R16532 a_219526_n14006.n246 a_219526_n14006.n245 0.3955
R16533 a_219526_n14006.n245 a_219526_n14006.n52 0.3955
R16534 a_219526_n14006.n404 a_219526_n14006.n52 0.3955
R16535 a_219526_n14006.n342 a_219526_n14006.n96 0.2555
R16536 a_219526_n14006.n345 a_219526_n14006.n38 0.2555
R16537 a_219526_n14006.n313 a_219526_n14006.n104 0.2505
R16538 a_219526_n14006.n164 a_219526_n14006.n12 0.231176
R16539 a_219526_n14006.n139 a_219526_n14006.n10 0.231176
R16540 a_219526_n14006.n129 a_219526_n14006.n8 0.231176
R16541 a_219526_n14006.n72 a_219526_n14006.n6 0.231176
R16542 a_219526_n14006.n184 a_219526_n14006.n29 0.225742
R16543 a_219526_n14006.n217 a_219526_n14006.n27 0.225742
R16544 a_219526_n14006.n209 a_219526_n14006.n25 0.225742
R16545 a_219526_n14006.n201 a_219526_n14006.n23 0.225742
R16546 a_219526_n14006.n193 a_219526_n14006.n21 0.225742
R16547 a_219526_n14006.n62 a_219526_n14006.n19 0.225742
R16548 a_219526_n14006.n376 a_219526_n14006.n16 0.225742
R16549 a_219526_n14006.n263 a_219526_n14006.n262 0.204667
R16550 a_219526_n14006.n349 a_219526_n14006.n348 0.204667
R16551 a_219526_n14006.n402 a_219526_n14006.n401 0.204667
R16552 a_219526_n14006.n238 a_219526_n14006.n106 0.2005
R16553 a_219526_n14006.n259 a_219526_n14006.n239 0.2005
R16554 a_219526_n14006.n309 a_219526_n14006.n308 0.2005
R16555 a_219526_n14006.n370 a_219526_n14006.n79 0.2005
R16556 a_219526_n14006.n406 a_219526_n14006.n405 0.2005
R16557 a_219526_n14006.n377 a_219526_n14006.n376 0.196152
R16558 a_219526_n14006.n75 a_219526_n14006.n74 0.196152
R16559 a_219526_n14006.n74 a_219526_n14006.n72 0.196152
R16560 a_219526_n14006.n132 a_219526_n14006.n131 0.196152
R16561 a_219526_n14006.n131 a_219526_n14006.n129 0.196152
R16562 a_219526_n14006.n142 a_219526_n14006.n141 0.196152
R16563 a_219526_n14006.n141 a_219526_n14006.n139 0.196152
R16564 a_219526_n14006.n163 a_219526_n14006.n148 0.196152
R16565 a_219526_n14006.n164 a_219526_n14006.n163 0.196152
R16566 a_219526_n14006.n63 a_219526_n14006.n62 0.196152
R16567 a_219526_n14006.n194 a_219526_n14006.n193 0.196152
R16568 a_219526_n14006.n202 a_219526_n14006.n201 0.196152
R16569 a_219526_n14006.n210 a_219526_n14006.n209 0.196152
R16570 a_219526_n14006.n218 a_219526_n14006.n217 0.196152
R16571 a_219526_n14006.n176 a_219526_n14006.n175 0.196152
R16572 a_219526_n14006.n184 a_219526_n14006.n183 0.196152
R16573 a_219526_n14006.n311 a_219526_n14006.n106 0.1955
R16574 a_219526_n14006.n176 a_219526_n14006.n1 0.194824
R16575 a_219526_n14006.n312 a_219526_n14006.n311 0.193
R16576 a_219526_n14006.n38 a_219526_n14006.n342 0.191241
R16577 a_219526_n14006.n249 a_219526_n14006.n100 0.190315
R16578 a_219526_n14006.n18 a_219526_n14006.n156 0.186853
R16579 a_219526_n14006.n313 a_219526_n14006.n312 0.178741
R16580 a_219526_n14006.n119 a_219526_n14006.n106 0.152583
R16581 a_219526_n14006.n278 a_219526_n14006.n263 0.1505
R16582 a_219526_n14006.n278 a_219526_n14006.n277 0.1505
R16583 a_219526_n14006.n277 a_219526_n14006.n275 0.1505
R16584 a_219526_n14006.n275 a_219526_n14006.n273 0.1505
R16585 a_219526_n14006.n273 a_219526_n14006.n271 0.1505
R16586 a_219526_n14006.n271 a_219526_n14006.n269 0.1505
R16587 a_219526_n14006.n269 a_219526_n14006.n267 0.1505
R16588 a_219526_n14006.n267 a_219526_n14006.n265 0.1505
R16589 a_219526_n14006.n284 a_219526_n14006.n31 0.1505
R16590 a_219526_n14006.n123 a_219526_n14006.n121 0.1505
R16591 a_219526_n14006.n303 a_219526_n14006.n119 0.1505
R16592 a_219526_n14006.n303 a_219526_n14006.n302 0.1505
R16593 a_219526_n14006.n302 a_219526_n14006.n300 0.1505
R16594 a_219526_n14006.n300 a_219526_n14006.n298 0.1505
R16595 a_219526_n14006.n298 a_219526_n14006.n296 0.1505
R16596 a_219526_n14006.n296 a_219526_n14006.n294 0.1505
R16597 a_219526_n14006.n294 a_219526_n14006.n292 0.1505
R16598 a_219526_n14006.n292 a_219526_n14006.n290 0.1505
R16599 a_219526_n14006.n365 a_219526_n14006.n349 0.1505
R16600 a_219526_n14006.n365 a_219526_n14006.n364 0.1505
R16601 a_219526_n14006.n364 a_219526_n14006.n362 0.1505
R16602 a_219526_n14006.n362 a_219526_n14006.n360 0.1505
R16603 a_219526_n14006.n360 a_219526_n14006.n358 0.1505
R16604 a_219526_n14006.n358 a_219526_n14006.n356 0.1505
R16605 a_219526_n14006.n356 a_219526_n14006.n354 0.1505
R16606 a_219526_n14006.n354 a_219526_n14006.n352 0.1505
R16607 a_219526_n14006.n85 a_219526_n14006.n84 0.1505
R16608 a_219526_n14006.n58 a_219526_n14006.n56 0.1505
R16609 a_219526_n14006.n401 a_219526_n14006.n400 0.1505
R16610 a_219526_n14006.n400 a_219526_n14006.n398 0.1505
R16611 a_219526_n14006.n398 a_219526_n14006.n396 0.1505
R16612 a_219526_n14006.n396 a_219526_n14006.n394 0.1505
R16613 a_219526_n14006.n394 a_219526_n14006.n392 0.1505
R16614 a_219526_n14006.n392 a_219526_n14006.n390 0.1505
R16615 a_219526_n14006.n390 a_219526_n14006.n388 0.1505
R16616 a_219526_n14006.n388 a_219526_n14006.n386 0.1505
R16617 a_219526_n14006.n265 a_219526_n14006.n2 0.149806
R16618 a_219526_n14006.n290 a_219526_n14006.n3 0.149806
R16619 a_219526_n14006.n352 a_219526_n14006.n4 0.149806
R16620 a_219526_n14006.n386 a_219526_n14006.n5 0.149806
R16621 a_219526_n14006.n32 a_219526_n14006.n31 0.145639
R16622 a_219526_n14006.n121 a_219526_n14006.n34 0.145639
R16623 a_219526_n14006.n84 a_219526_n14006.n35 0.145639
R16624 a_219526_n14006.n56 a_219526_n14006.n37 0.145639
R16625 a_219526_n14006.n262 a_219526_n14006.n261 0.1305
R16626 a_219526_n14006.n260 a_219526_n14006.n259 0.1305
R16627 a_219526_n14006.n402 a_219526_n14006.n54 0.1305
R16628 a_219526_n14006.n405 a_219526_n14006.n51 0.1305
R16629 a_219526_n14006.n309 a_219526_n14006.n107 0.1255
R16630 a_219526_n14006.n348 a_219526_n14006.n347 0.1255
R16631 a_219526_n14006.n346 a_219526_n14006.n79 0.1255
R16632 a_219526_n14006.n310 a_219526_n14006.n309 0.1205
R16633 a_219526_n14006.n344 a_219526_n14006.n79 0.1205
R16634 a_219526_n14006.n348 a_219526_n14006.n345 0.1205
R16635 a_219526_n14006.n15 a_219526_n14006.n14 0.118
R16636 a_219526_n14006.n403 a_219526_n14006.n402 0.1155
R16637 a_219526_n14006.n262 a_219526_n14006.n237 0.1155
R16638 a_219526_n14006.n259 a_219526_n14006.n258 0.1155
R16639 a_219526_n14006.n405 a_219526_n14006.n404 0.1155
R16640 a_219526_n14006.n148 a_219526_n14006.n18 0.112457
R16641 a_219526_n14006.n406 a_219526_n14006.n37 0.10675
R16642 a_219526_n14006.n35 a_219526_n14006.n370 0.10675
R16643 a_219526_n14006.n308 a_219526_n14006.n34 0.10675
R16644 a_219526_n14006.n239 a_219526_n14006.n32 0.10675
R16645 a_219526_n14006.n183 a_219526_n14006.n1 0.104486
R16646 a_219526_n14006.n5 a_219526_n14006.n58 0.102583
R16647 a_219526_n14006.n85 a_219526_n14006.n4 0.102583
R16648 a_219526_n14006.n3 a_219526_n14006.n123 0.102583
R16649 a_219526_n14006.n2 a_219526_n14006.n284 0.102583
R16650 a_219526_n14006.n287 a_219526_n14006.n166 0.0990583
R16651 a_219526_n14006.n372 a_219526_n14006.n371 0.0990583
R16652 a_219526_n14006.n75 a_219526_n14006.n68 0.0735676
R16653 a_219526_n14006.n132 a_219526_n14006.n125 0.0735676
R16654 a_219526_n14006.n142 a_219526_n14006.n124 0.0735676
R16655 a_219526_n14006.n325 a_219526_n14006.n100 0.0605
R16656 a_219526_n14006.n250 a_219526_n14006.n249 0.0605
R16657 a_219526_n14006.n377 a_219526_n14006.n373 0.0572633
R16658 a_219526_n14006.n63 a_219526_n14006.n59 0.0572633
R16659 a_219526_n14006.n194 a_219526_n14006.n190 0.0572633
R16660 a_219526_n14006.n202 a_219526_n14006.n189 0.0572633
R16661 a_219526_n14006.n210 a_219526_n14006.n188 0.0572633
R16662 a_219526_n14006.n218 a_219526_n14006.n187 0.0572633
R16663 a_219526_n14006.n249 a_219526_n14006.n248 0.0555
R16664 a_219526_n14006.n329 a_219526_n14006.n100 0.0555
R16665 a_219526_n14006.n286 a_219526_n14006.n186 0.0506333
R16666 a_219526_n14006.n285 a_219526_n14006.n222 0.0506333
R16667 a_219526_n14006.n214 a_219526_n14006.n206 0.0506333
R16668 a_219526_n14006.n206 a_219526_n14006.n198 0.0506333
R16669 a_219526_n14006.n383 a_219526_n14006.n67 0.0506333
R16670 a_219526_n14006.n382 a_219526_n14006.n381 0.0506333
R16671 a_219526_n14006.n286 a_219526_n14006.n285 0.0490667
R16672 a_219526_n14006.n222 a_219526_n14006.n214 0.0490667
R16673 a_219526_n14006.n198 a_219526_n14006.n67 0.0490667
R16674 a_219526_n14006.n383 a_219526_n14006.n382 0.0490667
R16675 1Bit_Clk_ADC_0.x14.Y 1Bit_Clk_ADC_0.x14.Y.n20 305.704
R16676 1Bit_Clk_ADC_0.x14.Y 1Bit_Clk_ADC_0.x14.Y.t1 239.244
R16677 1Bit_Clk_ADC_0.x14.Y.n9 1Bit_Clk_ADC_0.x14.Y.t8 212.081
R16678 1Bit_Clk_ADC_0.x14.Y.n8 1Bit_Clk_ADC_0.x14.Y.t17 212.081
R16679 1Bit_Clk_ADC_0.x14.Y.n12 1Bit_Clk_ADC_0.x14.Y.t6 212.081
R16680 1Bit_Clk_ADC_0.x14.Y.n14 1Bit_Clk_ADC_0.x14.Y.t15 212.081
R16681 1Bit_Clk_ADC_0.x14.Y.n1 1Bit_Clk_ADC_0.x14.Y.t10 212.081
R16682 1Bit_Clk_ADC_0.x14.Y.n3 1Bit_Clk_ADC_0.x14.Y.t16 212.081
R16683 1Bit_Clk_ADC_0.x14.Y.n5 1Bit_Clk_ADC_0.x14.Y.t14 212.081
R16684 1Bit_Clk_ADC_0.x14.Y.n4 1Bit_Clk_ADC_0.x14.Y.t9 212.081
R16685 1Bit_Clk_ADC_0.x14.Y.n14 1Bit_Clk_ADC_0.x14.Y.n13 180.482
R16686 1Bit_Clk_ADC_0.x14.Y 1Bit_Clk_ADC_0.x14.Y.n6 158.656
R16687 1Bit_Clk_ADC_0.x14.Y 1Bit_Clk_ADC_0.x14.Y.n10 152
R16688 1Bit_Clk_ADC_0.x14.Y.n11 1Bit_Clk_ADC_0.x14.Y 152
R16689 1Bit_Clk_ADC_0.x14.Y.n16 1Bit_Clk_ADC_0.x14.Y.n15 152
R16690 1Bit_Clk_ADC_0.x14.Y.n2 1Bit_Clk_ADC_0.x14.Y.n0 152
R16691 1Bit_Clk_ADC_0.x14.Y.n9 1Bit_Clk_ADC_0.x14.Y.t4 139.78
R16692 1Bit_Clk_ADC_0.x14.Y.n8 1Bit_Clk_ADC_0.x14.Y.t13 139.78
R16693 1Bit_Clk_ADC_0.x14.Y.n12 1Bit_Clk_ADC_0.x14.Y.t18 139.78
R16694 1Bit_Clk_ADC_0.x14.Y.n14 1Bit_Clk_ADC_0.x14.Y.t11 139.78
R16695 1Bit_Clk_ADC_0.x14.Y.n1 1Bit_Clk_ADC_0.x14.Y.t5 139.78
R16696 1Bit_Clk_ADC_0.x14.Y.n3 1Bit_Clk_ADC_0.x14.Y.t12 139.78
R16697 1Bit_Clk_ADC_0.x14.Y.n5 1Bit_Clk_ADC_0.x14.Y.t7 139.78
R16698 1Bit_Clk_ADC_0.x14.Y.n4 1Bit_Clk_ADC_0.x14.Y.t3 139.78
R16699 1Bit_Clk_ADC_0.x14.Y.n5 1Bit_Clk_ADC_0.x14.Y.n4 61.346
R16700 1Bit_Clk_ADC_0.x14.Y.n20 1Bit_Clk_ADC_0.x14.Y.t0 31.6612
R16701 1Bit_Clk_ADC_0.x14.Y.n20 1Bit_Clk_ADC_0.x14.Y.t2 31.6612
R16702 1Bit_Clk_ADC_0.x14.Y.n10 1Bit_Clk_ADC_0.x14.Y.n9 30.6732
R16703 1Bit_Clk_ADC_0.x14.Y.n10 1Bit_Clk_ADC_0.x14.Y.n8 30.6732
R16704 1Bit_Clk_ADC_0.x14.Y.n11 1Bit_Clk_ADC_0.x14.Y.n8 30.6732
R16705 1Bit_Clk_ADC_0.x14.Y.n12 1Bit_Clk_ADC_0.x14.Y.n11 30.6732
R16706 1Bit_Clk_ADC_0.x14.Y.n15 1Bit_Clk_ADC_0.x14.Y.n12 30.6732
R16707 1Bit_Clk_ADC_0.x14.Y.n15 1Bit_Clk_ADC_0.x14.Y.n14 30.6732
R16708 1Bit_Clk_ADC_0.x14.Y.n2 1Bit_Clk_ADC_0.x14.Y.n1 30.6732
R16709 1Bit_Clk_ADC_0.x14.Y.n3 1Bit_Clk_ADC_0.x14.Y.n2 30.6732
R16710 1Bit_Clk_ADC_0.x14.Y.n6 1Bit_Clk_ADC_0.x14.Y.n3 30.6732
R16711 1Bit_Clk_ADC_0.x14.Y.n6 1Bit_Clk_ADC_0.x14.Y.n5 30.6732
R16712 1Bit_Clk_ADC_0.x14.Y.n19 1Bit_Clk_ADC_0.x14.Y.n18 18.9312
R16713 1Bit_Clk_ADC_0.x14.Y.n18 1Bit_Clk_ADC_0.x14.Y.n17 18.556
R16714 1Bit_Clk_ADC_0.x14.Y.n18 1Bit_Clk_ADC_0.x14.Y.n7 18.0371
R16715 1Bit_Clk_ADC_0.x14.Y.n13 1Bit_Clk_ADC_0.x14.Y 17.1525
R16716 1Bit_Clk_ADC_0.x14.Y.n17 1Bit_Clk_ADC_0.x14.Y.n16 16.6405
R16717 1Bit_Clk_ADC_0.x14.Y.n7 1Bit_Clk_ADC_0.x14.Y 9.7285
R16718 1Bit_Clk_ADC_0.x14.Y.n0 1Bit_Clk_ADC_0.x14.Y 8.7045
R16719 1Bit_Clk_ADC_0.x14.Y.n13 1Bit_Clk_ADC_0.x14.Y 6.4005
R16720 1Bit_Clk_ADC_0.x14.Y.n7 1Bit_Clk_ADC_0.x14.Y.n0 5.1205
R16721 1Bit_Clk_ADC_0.x14.Y.n17 1Bit_Clk_ADC_0.x14.Y 4.8645
R16722 1Bit_Clk_ADC_0.x14.Y.n16 1Bit_Clk_ADC_0.x14.Y 3.5845
R16723 1Bit_Clk_ADC_0.x14.Y 1Bit_Clk_ADC_0.x14.Y.n19 3.11845
R16724 1Bit_Clk_ADC_0.x14.Y.n19 1Bit_Clk_ADC_0.x14.Y 2.46204
R16725 GND.n3110 GND.n3109 150626
R16726 GND.n7690 GND.n2312 132052
R16727 GND.n7746 GND.n7736 54534.2
R16728 GND.n7741 GND.n7736 54534.2
R16729 GND.n7746 GND.n7737 54534.2
R16730 GND.n7741 GND.n7737 54534.2
R16731 GND.n9816 GND.n18 54534.2
R16732 GND.n9816 GND.n19 54534.2
R16733 GND.n9810 GND.n18 54534.2
R16734 GND.n9810 GND.n19 54534.2
R16735 GND.n9783 GND.n52 54534.2
R16736 GND.n9783 GND.n53 54534.2
R16737 GND.n9793 GND.n53 54534.2
R16738 GND.n9793 GND.n52 54534.2
R16739 GND.n8430 GND.n1800 54534.2
R16740 GND.n8430 GND.n1801 54534.2
R16741 GND.n1805 GND.n1801 54534.2
R16742 GND.n1805 GND.n1800 54534.2
R16743 GND.n9819 GND.n9818 22436.9
R16744 GND.n7703 GND.n2307 22436.9
R16745 GND.n7716 GND.n2273 10309.9
R16746 GND.n8031 GND.n8030 7076.19
R16747 GND.n5984 GND.n5983 6944.74
R16748 GND.n7720 GND.n2300 6871.82
R16749 GND.n7720 GND.n2301 6871.82
R16750 GND.n7721 GND.n2300 6871.82
R16751 GND.n7721 GND.n2301 6871.82
R16752 GND.n7705 GND.n2302 6871.82
R16753 GND.n7713 GND.n2302 6871.82
R16754 GND.n7705 GND.n2303 6871.82
R16755 GND.n7713 GND.n2303 6871.82
R16756 GND.n9453 GND.n9433 6871.82
R16757 GND.n9461 GND.n9433 6871.82
R16758 GND.n9453 GND.n9434 6871.82
R16759 GND.n9461 GND.n9434 6871.82
R16760 GND.n9442 GND.n9438 6871.82
R16761 GND.n9450 GND.n9438 6871.82
R16762 GND.n9442 GND.n9439 6871.82
R16763 GND.n9450 GND.n9439 6871.82
R16764 GND.n3113 GND.n3112 6475.12
R16765 GND.n8728 GND.n1653 5640.12
R16766 GND.n2934 GND.n2312 5503.96
R16767 GND.n5983 GND.n3696 5364.7
R16768 GND.n7693 GND.n2308 4925
R16769 GND.n7701 GND.n2308 4925
R16770 GND.n7693 GND.n2309 4925
R16771 GND.n7701 GND.n2309 4925
R16772 GND.n2118 GND.n13 4925
R16773 GND.n9821 GND.n13 4925
R16774 GND.n2118 GND.n14 4925
R16775 GND.n9821 GND.n14 4925
R16776 GND.n3112 GND.n3110 4039.17
R16777 GND.n7745 GND.n7744 3543.34
R16778 GND.n7745 GND.n7738 3543.34
R16779 GND.n9811 GND.n20 3543.34
R16780 GND.n9815 GND.n20 3543.34
R16781 GND.n9784 GND.n54 3543.34
R16782 GND.n9792 GND.n54 3543.34
R16783 GND.n8429 GND.n1802 3543.34
R16784 GND.n1806 GND.n1802 3543.34
R16785 GND.n7692 GND.n7690 3543.24
R16786 GND.n9797 GND.n50 3320.29
R16787 GND.n8499 GND.t20 3221.5
R16788 GND.n9792 GND.n9791 2581.08
R16789 GND.n8424 GND.n1806 2543.44
R16790 GND.n8429 GND.n8428 2458.22
R16791 GND.n9785 GND.n9784 2420.57
R16792 GND.n3111 GND.n2720 2316.25
R16793 GND GND.t385 2243.48
R16794 GND.n3399 GND.t105 2083.62
R16795 GND.n7740 GND.n7738 1722.85
R16796 GND.n9815 GND.n9814 1722.85
R16797 GND.n7744 GND.n7743 1673.07
R16798 GND.n9812 GND.n9811 1673.07
R16799 GND.n8030 GND.n2119 1509.34
R16800 GND.n9795 GND.n51 1389.5
R16801 GND.n504 GND.n229 1268.91
R16802 GND.n9343 GND.n294 1268.91
R16803 GND.n790 GND.n753 1268.91
R16804 GND.n9312 GND.n9311 1268.91
R16805 GND.n793 GND.n792 1268.91
R16806 GND.n9347 GND.n298 1268.91
R16807 GND.n322 GND.n316 1268.91
R16808 GND.n855 GND.n522 1268.91
R16809 GND.n4358 GND.n1921 1268.91
R16810 GND.n8237 GND.n1986 1268.91
R16811 GND.n4402 GND.n4265 1268.91
R16812 GND.n8206 GND.n8205 1268.91
R16813 GND.n4447 GND.n4267 1268.91
R16814 GND.n8241 GND.n1990 1268.91
R16815 GND.n2014 GND.n2008 1268.91
R16816 GND.n4439 GND.n4266 1268.91
R16817 GND.n7139 GND.n6677 1268.91
R16818 GND.n2577 GND.n2524 1268.91
R16819 GND.n7083 GND.n6673 1268.91
R16820 GND.n2610 GND.n2609 1268.91
R16821 GND.n6694 GND.n6676 1268.91
R16822 GND.n7363 GND.n2529 1268.91
R16823 GND.n7115 GND.n6674 1268.91
R16824 GND.n7332 GND.n7331 1268.91
R16825 GND.n7735 GND.n7734 1268.46
R16826 GND.n6802 GND.n2313 1252.97
R16827 GND.n7638 GND.n2340 1245.74
R16828 GND.n5620 GND.n2395 1245.74
R16829 GND.n5546 GND.n2338 1245.74
R16830 GND.n5616 GND.n5559 1245.74
R16831 GND.n7833 GND.n2258 1245.74
R16832 GND.n7984 GND.n2143 1245.74
R16833 GND.n7824 GND.n2256 1245.74
R16834 GND.n2194 GND.n2140 1245.74
R16835 GND.n9555 GND.n172 1245.74
R16836 GND.n9694 GND.n123 1245.74
R16837 GND.n9546 GND.n170 1245.74
R16838 GND.n9615 GND.n120 1245.74
R16839 GND.n9204 GND.n9139 1239.94
R16840 GND.n9171 GND.n9138 1239.94
R16841 GND.n617 GND.n574 1239.94
R16842 GND.n614 GND.n572 1239.94
R16843 GND.n8098 GND.n8033 1239.94
R16844 GND.n8065 GND.n2111 1239.94
R16845 GND.n8363 GND.n8362 1239.94
R16846 GND.n8395 GND.n1825 1239.94
R16847 GND.n6845 GND.n6804 1239.94
R16848 GND.n7495 GND.n7452 1239.94
R16849 GND.n7464 GND.n7450 1239.94
R16850 GND.n6847 GND.n6801 1239.94
R16851 GND.n6092 GND.n5986 1205.18
R16852 GND.n6094 GND.n3116 1205.18
R16853 GND.n6175 GND.n2865 1205.18
R16854 GND.n6185 GND.n2859 1205.18
R16855 GND.n6262 GND.n2768 1205.18
R16856 GND.n2813 GND.n2766 1205.18
R16857 GND.n6387 GND.n2737 1205.18
R16858 GND.n6390 GND.n6389 1205.18
R16859 GND.n5980 GND.n3720 1205.18
R16860 GND.n5897 GND.n5896 1205.18
R16861 GND.n5844 GND.n3811 1205.18
R16862 GND.n3982 GND.n3981 1205.18
R16863 GND.n5893 GND.n3726 1205.18
R16864 GND.n5276 GND.n3724 1205.18
R16865 GND.n5847 GND.n3786 1205.18
R16866 GND.n5311 GND.n3788 1205.18
R16867 GND.n5807 GND.n3840 1205.18
R16868 GND.n4080 GND.n4078 1205.18
R16869 GND.n4981 GND.n3896 1205.18
R16870 GND.n4112 GND.n4111 1205.18
R16871 GND.n5097 GND.n3847 1205.18
R16872 GND.n5369 GND.n5368 1205.18
R16873 GND.n5730 GND.n3902 1205.18
R16874 GND.n5402 GND.n5401 1205.18
R16875 GND.n1651 GND.n1093 1205.18
R16876 GND.n1527 GND.n1288 1205.18
R16877 GND.n1184 GND.n1089 1205.18
R16878 GND.n1351 GND.n1290 1205.18
R16879 GND.n1370 GND.n1092 1205.18
R16880 GND.n1525 GND.n1353 1205.18
R16881 GND.n1404 GND.n1090 1205.18
R16882 GND.n1489 GND.n1352 1205.18
R16883 GND.n8442 GND.n1794 1205.18
R16884 GND.n8730 GND.n1060 1205.18
R16885 GND.n8497 GND.n8441 1205.18
R16886 GND.n8696 GND.n1070 1205.18
R16887 GND.n3694 GND.n3139 1205.18
R16888 GND.n3570 GND.n3334 1205.18
R16889 GND.n3230 GND.n3135 1205.18
R16890 GND.n3344 GND.n3335 1205.18
R16891 GND.n8590 GND.n1798 1205.18
R16892 GND.n1721 GND.n1056 1205.18
R16893 GND.n8560 GND.n8559 1205.18
R16894 GND.n1687 GND.n1686 1205.18
R16895 GND.n3417 GND.n3138 1205.18
R16896 GND.n3568 GND.n3400 1205.18
R16897 GND.n3451 GND.n3136 1205.18
R16898 GND.n3532 GND.n3336 1205.18
R16899 GND.n3109 GND.n3108 1199.12
R16900 GND.n2935 GND.n2934 1174.88
R16901 GND.n7682 GND.n2325 1170.41
R16902 GND.n7588 GND.n2408 1170.41
R16903 GND.n7650 GND.n7649 1170.41
R16904 GND.n5590 GND.n2407 1170.41
R16905 GND.n7788 GND.n2267 1170.41
R16906 GND.n8027 GND.n2129 1170.41
R16907 GND.n7791 GND.n2270 1170.41
R16908 GND.n7996 GND.n7995 1170.41
R16909 GND.n9506 GND.n186 1170.41
R16910 GND.n9682 GND.n9620 1170.41
R16911 GND.n9475 GND.n9474 1170.41
R16912 GND.n9648 GND.n9621 1170.41
R16913 GND.n2998 GND.n2997 1170
R16914 GND.n3000 GND.n2999 1170
R16915 GND.n3079 GND.n3078 1170
R16916 GND.n3081 GND.n3080 1170
R16917 GND.n3112 GND.n3111 1152.21
R16918 GND.n9133 GND.n408 1124.06
R16919 GND.n9102 GND.n9101 1124.06
R16920 GND.n648 GND.n558 1124.06
R16921 GND.n679 GND.n561 1124.06
R16922 GND.n4568 GND.n2098 1124.06
R16923 GND.n4601 GND.n4600 1124.06
R16924 GND.n4314 GND.n1837 1124.06
R16925 GND.n8352 GND.n1839 1124.06
R16926 GND.n6914 GND.n6789 1124.06
R16927 GND.n6874 GND.n6791 1124.06
R16928 GND.n7550 GND.n2464 1124.06
R16929 GND.n7519 GND.n7518 1124.06
R16930 GND.n7624 GND.n2360 1077.71
R16931 GND.n5476 GND.n5471 1077.71
R16932 GND.n5517 GND.n2358 1077.71
R16933 GND.n5643 GND.n5464 1077.71
R16934 GND.n2232 GND.n2231 1077.71
R16935 GND.n7953 GND.n2165 1077.71
R16936 GND.n7863 GND.n2227 1077.71
R16937 GND.n7932 GND.n2179 1077.71
R16938 GND.n141 GND.n77 1077.71
R16939 GND.n9732 GND.n81 1077.71
R16940 GND.n9591 GND.n9590 1077.71
R16941 GND.n9711 GND.n95 1077.71
R16942 GND.n9818 GND.n9817 1030.62
R16943 GND.n3109 GND.n2892 1008.7
R16944 GND GND.t334 939.736
R16945 GND.n9463 GND.n9462 926.02
R16946 GND.n9798 GND.n9797 905.774
R16947 GND.t69 GND.n1815 887.173
R16948 GND.n9819 GND.n15 886.197
R16949 GND.n7704 GND.n7703 886.197
R16950 GND.n3110 GND.n2313 765.915
R16951 GND.n9809 GND.n9808 656.13
R16952 GND.n3110 GND.n2312 645.995
R16953 GND.t339 GND.t129 611.92
R16954 GND.t129 GND.t133 611.92
R16955 GND.t360 GND.t90 611.92
R16956 GND.t84 GND.t416 611.92
R16957 GND.t383 GND.t389 611.92
R16958 GND.n9809 GND.n25 587.528
R16959 GND.n9343 GND.n9342 585
R16960 GND.n9341 GND.n319 585
R16961 GND.n9340 GND.n318 585
R16962 GND.n9345 GND.n318 585
R16963 GND.n9339 GND.n9338 585
R16964 GND.n9337 GND.n9336 585
R16965 GND.n9335 GND.n9334 585
R16966 GND.n9333 GND.n9332 585
R16967 GND.n9331 GND.n9330 585
R16968 GND.n9329 GND.n9328 585
R16969 GND.n9327 GND.n9326 585
R16970 GND.n9325 GND.n9324 585
R16971 GND.n9323 GND.n9322 585
R16972 GND.n9321 GND.n9320 585
R16973 GND.n9319 GND.n9318 585
R16974 GND.n9317 GND.n9316 585
R16975 GND.n9315 GND.n9314 585
R16976 GND.n9313 GND.n9312 585
R16977 GND.n9311 GND.n320 585
R16978 GND.n9311 GND.n9310 585
R16979 GND.n966 GND.n295 585
R16980 GND.n9352 GND.n295 585
R16981 GND.n967 GND.n348 585
R16982 GND.n9280 GND.n348 585
R16983 GND.n968 GND.n287 585
R16984 GND.n9358 GND.n287 585
R16985 GND.n971 GND.n970 585
R16986 GND.n970 GND.n358 585
R16987 GND.n973 GND.n276 585
R16988 GND.n9366 GND.n276 585
R16989 GND.n965 GND.n447 585
R16990 GND.n9046 GND.n447 585
R16991 GND.n962 GND.n267 585
R16992 GND.n9375 GND.n267 585
R16993 GND.n961 GND.n960 585
R16994 GND.n960 GND.t39 585
R16995 GND.n959 GND.n257 585
R16996 GND.n9381 GND.n257 585
R16997 GND.n472 GND.n464 585
R16998 GND.n8975 GND.n464 585
R16999 GND.n953 GND.n245 585
R17000 GND.n9390 GND.n245 585
R17001 GND.n951 GND.n950 585
R17002 GND.n950 GND.n949 585
R17003 GND.n786 GND.n235 585
R17004 GND.n9398 GND.n235 585
R17005 GND.n787 GND.n491 585
R17006 GND.n926 GND.n491 585
R17007 GND.n788 GND.n226 585
R17008 GND.n9404 GND.n226 585
R17009 GND.n790 GND.n789 585
R17010 GND.n791 GND.n790 585
R17011 GND.n785 GND.n753 585
R17012 GND.n784 GND.n783 585
R17013 GND.n782 GND.n781 585
R17014 GND.n780 GND.n779 585
R17015 GND.n778 GND.n777 585
R17016 GND.n776 GND.n775 585
R17017 GND.n774 GND.n773 585
R17018 GND.n772 GND.n771 585
R17019 GND.n770 GND.n769 585
R17020 GND.n768 GND.n767 585
R17021 GND.n766 GND.n765 585
R17022 GND.n764 GND.n763 585
R17023 GND.n762 GND.n761 585
R17024 GND.n760 GND.n759 585
R17025 GND.n758 GND.n757 585
R17026 GND.n756 GND.n755 585
R17027 GND.n754 GND.n504 585
R17028 GND.n856 GND.n504 585
R17029 GND.n231 GND.n229 585
R17030 GND.n791 GND.n229 585
R17031 GND.n9403 GND.n9402 585
R17032 GND.n9404 GND.n9403 585
R17033 GND.n9401 GND.n230 585
R17034 GND.n926 GND.n230 585
R17035 GND.n9400 GND.n9399 585
R17036 GND.n9399 GND.n9398 585
R17037 GND.n249 GND.n233 585
R17038 GND.n949 GND.n233 585
R17039 GND.n9389 GND.n9388 585
R17040 GND.n9390 GND.n9389 585
R17041 GND.n251 GND.n248 585
R17042 GND.n8975 GND.n248 585
R17043 GND.n9383 GND.n9382 585
R17044 GND.n9382 GND.n9381 585
R17045 GND.n255 GND.n254 585
R17046 GND.t39 GND.n255 585
R17047 GND.n9374 GND.n9373 585
R17048 GND.n9375 GND.n9374 585
R17049 GND.n271 GND.n270 585
R17050 GND.n9046 GND.n270 585
R17051 GND.n9368 GND.n9367 585
R17052 GND.n9367 GND.n9366 585
R17053 GND.n291 GND.n274 585
R17054 GND.n358 GND.n274 585
R17055 GND.n9357 GND.n9356 585
R17056 GND.n9358 GND.n9357 585
R17057 GND.n9355 GND.n290 585
R17058 GND.n9280 GND.n290 585
R17059 GND.n9354 GND.n9353 585
R17060 GND.n9353 GND.n9352 585
R17061 GND.n294 GND.n293 585
R17062 GND.n9310 GND.n294 585
R17063 GND.n855 GND.n854 585
R17064 GND.n856 GND.n855 585
R17065 GND.n823 GND.n521 585
R17066 GND.n822 GND.n821 585
R17067 GND.n820 GND.n819 585
R17068 GND.n818 GND.n817 585
R17069 GND.n816 GND.n815 585
R17070 GND.n814 GND.n813 585
R17071 GND.n812 GND.n811 585
R17072 GND.n810 GND.n809 585
R17073 GND.n808 GND.n807 585
R17074 GND.n806 GND.n805 585
R17075 GND.n804 GND.n803 585
R17076 GND.n802 GND.n801 585
R17077 GND.n800 GND.n799 585
R17078 GND.n798 GND.n797 585
R17079 GND.n796 GND.n795 585
R17080 GND.n794 GND.n793 585
R17081 GND.n792 GND.n524 585
R17082 GND.n792 GND.n791 585
R17083 GND.n523 GND.n228 585
R17084 GND.n9404 GND.n228 585
R17085 GND.n239 GND.n237 585
R17086 GND.n926 GND.n237 585
R17087 GND.n9397 GND.n9396 585
R17088 GND.n9398 GND.n9397 585
R17089 GND.n240 GND.n238 585
R17090 GND.n949 GND.n238 585
R17091 GND.n9392 GND.n9391 585
R17092 GND.n9391 GND.n9390 585
R17093 GND.n261 GND.n243 585
R17094 GND.n8975 GND.n243 585
R17095 GND.n9380 GND.n9379 585
R17096 GND.n9381 GND.n9380 585
R17097 GND.n9378 GND.n260 585
R17098 GND.t39 GND.n260 585
R17099 GND.n9377 GND.n9376 585
R17100 GND.n9376 GND.n9375 585
R17101 GND.n280 GND.n265 585
R17102 GND.n9046 GND.n265 585
R17103 GND.n9365 GND.n9364 585
R17104 GND.n9366 GND.n9365 585
R17105 GND.n282 GND.n279 585
R17106 GND.n358 GND.n279 585
R17107 GND.n9360 GND.n9359 585
R17108 GND.n9359 GND.n9358 585
R17109 GND.n285 GND.n284 585
R17110 GND.n9280 GND.n285 585
R17111 GND.n9351 GND.n9350 585
R17112 GND.n9352 GND.n9351 585
R17113 GND.n9349 GND.n298 585
R17114 GND.n9310 GND.n298 585
R17115 GND.n9348 GND.n9347 585
R17116 GND.n300 GND.n299 585
R17117 GND.n8984 GND.n8983 585
R17118 GND.n8986 GND.n8985 585
R17119 GND.n8988 GND.n8987 585
R17120 GND.n8990 GND.n8989 585
R17121 GND.n8992 GND.n8991 585
R17122 GND.n8994 GND.n8993 585
R17123 GND.n8996 GND.n8995 585
R17124 GND.n8998 GND.n8997 585
R17125 GND.n9000 GND.n8999 585
R17126 GND.n9002 GND.n9001 585
R17127 GND.n9004 GND.n9003 585
R17128 GND.n9006 GND.n9005 585
R17129 GND.n9008 GND.n9007 585
R17130 GND.n9010 GND.n9009 585
R17131 GND.n9011 GND.n316 585
R17132 GND.n9345 GND.n316 585
R17133 GND.n9012 GND.n322 585
R17134 GND.n9310 GND.n322 585
R17135 GND.n9013 GND.n296 585
R17136 GND.n9352 GND.n296 585
R17137 GND.n9014 GND.n349 585
R17138 GND.n9280 GND.n349 585
R17139 GND.n9015 GND.n288 585
R17140 GND.n9358 GND.n288 585
R17141 GND.n8982 GND.n8981 585
R17142 GND.n8981 GND.n358 585
R17143 GND.n9019 GND.n277 585
R17144 GND.n9366 GND.n277 585
R17145 GND.n9021 GND.n448 585
R17146 GND.n9046 GND.n448 585
R17147 GND.n9023 GND.n268 585
R17148 GND.n9375 GND.n268 585
R17149 GND.n9024 GND.n8980 585
R17150 GND.n8980 GND.t39 585
R17151 GND.n8979 GND.n258 585
R17152 GND.n9381 GND.n258 585
R17153 GND.n8977 GND.n8976 585
R17154 GND.n8976 GND.n8975 585
R17155 GND.n846 GND.n246 585
R17156 GND.n9390 GND.n246 585
R17157 GND.n824 GND.n476 585
R17158 GND.n949 GND.n476 585
R17159 GND.n850 GND.n236 585
R17160 GND.n9398 GND.n236 585
R17161 GND.n851 GND.n492 585
R17162 GND.n926 GND.n492 585
R17163 GND.n852 GND.n227 585
R17164 GND.n9404 GND.n227 585
R17165 GND.n853 GND.n522 585
R17166 GND.n791 GND.n522 585
R17167 GND.n9428 GND.n193 585
R17168 GND.n735 GND.n193 585
R17169 GND.n9427 GND.n9426 585
R17170 GND.n9426 GND.n9425 585
R17171 GND.n216 GND.n196 585
R17172 GND.n200 GND.n196 585
R17173 GND.n217 GND.n212 585
R17174 GND.n857 GND.n212 585
R17175 GND.n9413 GND.n9412 585
R17176 GND.n9414 GND.n9413 585
R17177 GND.n215 GND.n213 585
R17178 GND.n752 GND.n213 585
R17179 GND.n9407 GND.n9406 585
R17180 GND.n9406 GND.n9405 585
R17181 GND.n831 GND.n223 585
R17182 GND.n927 GND.n223 585
R17183 GND.n830 GND.n829 585
R17184 GND.n829 GND.n234 585
R17185 GND.n838 GND.n837 585
R17186 GND.n838 GND.n475 585
R17187 GND.n839 GND.n827 585
R17188 GND.n839 GND.n244 585
R17189 GND.n841 GND.n840 585
R17190 GND.n840 GND.n463 585
R17191 GND.n458 GND.n457 585
R17192 GND.n457 GND.n256 585
R17193 GND.n9029 GND.n9028 585
R17194 GND.n9030 GND.n9029 585
R17195 GND.n9027 GND.n445 585
R17196 GND.n445 GND.n266 585
R17197 GND.n9049 GND.n9048 585
R17198 GND.n9048 GND.n9047 585
R17199 GND.n9050 GND.n439 585
R17200 GND.n439 GND.n275 585
R17201 GND.n9058 GND.n9057 585
R17202 GND.n9059 GND.n9058 585
R17203 GND.n441 GND.n346 585
R17204 GND.n346 GND.n286 585
R17205 GND.n9283 GND.n9282 585
R17206 GND.n9282 GND.n9281 585
R17207 GND.n343 GND.n342 585
R17208 GND.n351 GND.n342 585
R17209 GND.n9289 GND.n9288 585
R17210 GND.n9289 GND.n321 585
R17211 GND.n9291 GND.n9290 585
R17212 GND.n9290 GND.n324 585
R17213 GND.n9292 GND.n336 585
R17214 GND.n336 GND.n317 585
R17215 GND.n9298 GND.n9297 585
R17216 GND.n9299 GND.n9298 585
R17217 GND.n339 GND.n337 585
R17218 GND.n371 GND.n337 585
R17219 GND.n387 GND.n386 585
R17220 GND.n386 GND.n372 585
R17221 GND.n9083 GND.n427 585
R17222 GND.n9083 GND.n372 585
R17223 GND.n9082 GND.n9081 585
R17224 GND.n9082 GND.n371 585
R17225 GND.n428 GND.n334 585
R17226 GND.n9299 GND.n334 585
R17227 GND.n9077 GND.n9076 585
R17228 GND.n9076 GND.n317 585
R17229 GND.n9075 GND.n9074 585
R17230 GND.n9075 GND.n324 585
R17231 GND.n432 GND.n431 585
R17232 GND.n431 GND.n321 585
R17233 GND.n9069 GND.n9068 585
R17234 GND.n9068 GND.n351 585
R17235 GND.n9066 GND.n347 585
R17236 GND.n9281 GND.n347 585
R17237 GND.n438 GND.n434 585
R17238 GND.n438 GND.n286 585
R17239 GND.n9061 GND.n9060 585
R17240 GND.n9060 GND.n9059 585
R17241 GND.n9034 GND.n437 585
R17242 GND.n437 GND.n275 585
R17243 GND.n9036 GND.n446 585
R17244 GND.n9047 GND.n446 585
R17245 GND.n9033 GND.n9032 585
R17246 GND.n9032 GND.n266 585
R17247 GND.n9031 GND.n455 585
R17248 GND.n9031 GND.n9030 585
R17249 GND.n484 GND.n456 585
R17250 GND.n456 GND.n256 585
R17251 GND.n939 GND.n938 585
R17252 GND.n938 GND.n463 585
R17253 GND.n937 GND.n483 585
R17254 GND.n937 GND.n244 585
R17255 GND.n936 GND.n935 585
R17256 GND.n936 GND.n475 585
R17257 GND.n487 GND.n486 585
R17258 GND.n486 GND.n234 585
R17259 GND.n929 GND.n928 585
R17260 GND.n928 GND.n927 585
R17261 GND.n526 GND.n225 585
R17262 GND.n9405 GND.n225 585
R17263 GND.n751 GND.n750 585
R17264 GND.n752 GND.n751 585
R17265 GND.n744 GND.n210 585
R17266 GND.n9414 GND.n210 585
R17267 GND.n743 GND.n503 585
R17268 GND.n857 GND.n503 585
R17269 GND.n741 GND.n740 585
R17270 GND.n740 GND.n200 585
R17271 GND.n738 GND.n198 585
R17272 GND.n9425 GND.n198 585
R17273 GND.n737 GND.n736 585
R17274 GND.n736 GND.n735 585
R17275 GND.n726 GND.n725 585
R17276 GND.n725 GND.n724 585
R17277 GND.n535 GND.n201 585
R17278 GND.n201 GND.n197 585
R17279 GND.n9423 GND.n9422 585
R17280 GND.n9424 GND.n9423 585
R17281 GND.n204 GND.n202 585
R17282 GND.n858 GND.n202 585
R17283 GND.n9417 GND.n9416 585
R17284 GND.n9416 GND.n9415 585
R17285 GND.n913 GND.n208 585
R17286 GND.n211 GND.n208 585
R17287 GND.n916 GND.n915 585
R17288 GND.n915 GND.n224 585
R17289 GND.n917 GND.n909 585
R17290 GND.n909 GND.n490 585
R17291 GND.n924 GND.n923 585
R17292 GND.n925 GND.n924 585
R17293 GND.n911 GND.n478 585
R17294 GND.n494 GND.n478 585
R17295 GND.n947 GND.n946 585
R17296 GND.n948 GND.n947 585
R17297 GND.n480 GND.n466 585
R17298 GND.n466 GND.n247 585
R17299 GND.n8973 GND.n8972 585
R17300 GND.n8974 GND.n8973 585
R17301 GND.n469 GND.n467 585
R17302 GND.n467 GND.n259 585
R17303 GND.n890 GND.n889 585
R17304 GND.n891 GND.n890 585
R17305 GND.n887 GND.n450 585
R17306 GND.n450 GND.n269 585
R17307 GND.n9044 GND.n9043 585
R17308 GND.n9045 GND.n9044 585
R17309 GND.n452 GND.n357 585
R17310 GND.n357 GND.n278 585
R17311 GND.n9270 GND.n9269 585
R17312 GND.n9269 GND.n9268 585
R17313 GND.n9271 GND.n352 585
R17314 GND.n352 GND.n289 585
R17315 GND.n9278 GND.n9277 585
R17316 GND.n9279 GND.n9278 585
R17317 GND.n354 GND.n325 585
R17318 GND.n325 GND.n297 585
R17319 GND.n9308 GND.n9307 585
R17320 GND.n9309 GND.n9308 585
R17321 GND.n328 GND.n326 585
R17322 GND.n326 GND.n301 585
R17323 GND.n9302 GND.n9301 585
R17324 GND.n9301 GND.n9300 585
R17325 GND.n374 GND.n332 585
R17326 GND.n335 GND.n332 585
R17327 GND.n9242 GND.n9241 585
R17328 GND.n9243 GND.n9242 585
R17329 GND.n9238 GND.n373 585
R17330 GND.n378 GND.n373 585
R17331 GND.n9148 GND.n370 585
R17332 GND.n378 GND.n370 585
R17333 GND.n9245 GND.n9244 585
R17334 GND.n9244 GND.n9243 585
R17335 GND.n369 GND.n367 585
R17336 GND.n369 GND.n335 585
R17337 GND.n9250 GND.n333 585
R17338 GND.n9300 GND.n333 585
R17339 GND.n9253 GND.n9252 585
R17340 GND.n9252 GND.n301 585
R17341 GND.n365 GND.n323 585
R17342 GND.n9309 GND.n323 585
R17343 GND.n9259 GND.n9258 585
R17344 GND.n9258 GND.n297 585
R17345 GND.n9261 GND.n350 585
R17346 GND.n9279 GND.n350 585
R17347 GND.n362 GND.n360 585
R17348 GND.n360 GND.n289 585
R17349 GND.n9267 GND.n9266 585
R17350 GND.n9268 GND.n9267 585
R17351 GND.n880 GND.n359 585
R17352 GND.n359 GND.n278 585
R17353 GND.n878 GND.n449 585
R17354 GND.n9045 GND.n449 585
R17355 GND.n886 GND.n885 585
R17356 GND.n886 GND.n269 585
R17357 GND.n892 GND.n876 585
R17358 GND.n892 GND.n891 585
R17359 GND.n894 GND.n893 585
R17360 GND.n893 GND.n259 585
R17361 GND.n874 GND.n465 585
R17362 GND.n8974 GND.n465 585
R17363 GND.n900 GND.n899 585
R17364 GND.n899 GND.n247 585
R17365 GND.n902 GND.n477 585
R17366 GND.n948 GND.n477 585
R17367 GND.n497 GND.n495 585
R17368 GND.n495 GND.n494 585
R17369 GND.n908 GND.n907 585
R17370 GND.n925 GND.n908 585
R17371 GND.n869 GND.n493 585
R17372 GND.n493 GND.n490 585
R17373 GND.n868 GND.n867 585
R17374 GND.n867 GND.n224 585
R17375 GND.n866 GND.n865 585
R17376 GND.n866 GND.n211 585
R17377 GND.n500 GND.n209 585
R17378 GND.n9415 GND.n209 585
R17379 GND.n860 GND.n859 585
R17380 GND.n859 GND.n858 585
R17381 GND.n718 GND.n199 585
R17382 GND.n9424 GND.n199 585
R17383 GND.n717 GND.n538 585
R17384 GND.n538 GND.n197 585
R17385 GND.n723 GND.n722 585
R17386 GND.n724 GND.n723 585
R17387 GND.n8237 GND.n8236 585
R17388 GND.n8235 GND.n2011 585
R17389 GND.n8234 GND.n2010 585
R17390 GND.n8239 GND.n2010 585
R17391 GND.n8233 GND.n8232 585
R17392 GND.n8231 GND.n8230 585
R17393 GND.n8229 GND.n8228 585
R17394 GND.n8227 GND.n8226 585
R17395 GND.n8225 GND.n8224 585
R17396 GND.n8223 GND.n8222 585
R17397 GND.n8221 GND.n8220 585
R17398 GND.n8219 GND.n8218 585
R17399 GND.n8217 GND.n8216 585
R17400 GND.n8215 GND.n8214 585
R17401 GND.n8213 GND.n8212 585
R17402 GND.n8211 GND.n8210 585
R17403 GND.n8209 GND.n8208 585
R17404 GND.n8207 GND.n8206 585
R17405 GND.n8205 GND.n2012 585
R17406 GND.n8205 GND.n8204 585
R17407 GND.n4698 GND.n1987 585
R17408 GND.n8246 GND.n1987 585
R17409 GND.n4699 GND.n2040 585
R17410 GND.n8174 GND.n2040 585
R17411 GND.n4700 GND.n1979 585
R17412 GND.n8252 GND.n1979 585
R17413 GND.n4703 GND.n4702 585
R17414 GND.n4702 GND.n2050 585
R17415 GND.n4705 GND.n1968 585
R17416 GND.n8260 GND.n1968 585
R17417 GND.n4695 GND.n4694 585
R17418 GND.n4694 GND.n4196 585
R17419 GND.n4711 GND.n1959 585
R17420 GND.n8269 GND.n1959 585
R17421 GND.n4713 GND.n4712 585
R17422 GND.t40 GND.n4713 585
R17423 GND.n4693 GND.n1949 585
R17424 GND.n8275 GND.n1949 585
R17425 GND.n4491 GND.n4211 585
R17426 GND.n4492 GND.n4491 585
R17427 GND.n4687 GND.n1937 585
R17428 GND.n8284 GND.n1937 585
R17429 GND.n4685 GND.n4684 585
R17430 GND.n4684 GND.n4683 585
R17431 GND.n4397 GND.n1927 585
R17432 GND.n8292 GND.n1927 585
R17433 GND.n4398 GND.n4253 585
R17434 GND.n4503 GND.n4253 585
R17435 GND.n4399 GND.n1918 585
R17436 GND.n8298 GND.n1918 585
R17437 GND.n4400 GND.n4265 585
R17438 GND.n4448 GND.n4265 585
R17439 GND.n4402 GND.n4401 585
R17440 GND.n4396 GND.n4366 585
R17441 GND.n4395 GND.n4394 585
R17442 GND.n4393 GND.n4392 585
R17443 GND.n4391 GND.n4390 585
R17444 GND.n4389 GND.n4388 585
R17445 GND.n4387 GND.n4386 585
R17446 GND.n4385 GND.n4384 585
R17447 GND.n4383 GND.n4382 585
R17448 GND.n4381 GND.n4380 585
R17449 GND.n4379 GND.n4378 585
R17450 GND.n4377 GND.n4376 585
R17451 GND.n4375 GND.n4374 585
R17452 GND.n4373 GND.n4372 585
R17453 GND.n4371 GND.n4370 585
R17454 GND.n4369 GND.n4368 585
R17455 GND.n4367 GND.n4358 585
R17456 GND.n4440 GND.n4358 585
R17457 GND.n1923 GND.n1921 585
R17458 GND.n4448 GND.n1921 585
R17459 GND.n8297 GND.n8296 585
R17460 GND.n8298 GND.n8297 585
R17461 GND.n8295 GND.n1922 585
R17462 GND.n4503 GND.n1922 585
R17463 GND.n8294 GND.n8293 585
R17464 GND.n8293 GND.n8292 585
R17465 GND.n1941 GND.n1925 585
R17466 GND.n4683 GND.n1925 585
R17467 GND.n8283 GND.n8282 585
R17468 GND.n8284 GND.n8283 585
R17469 GND.n1943 GND.n1940 585
R17470 GND.n4492 GND.n1940 585
R17471 GND.n8277 GND.n8276 585
R17472 GND.n8276 GND.n8275 585
R17473 GND.n1947 GND.n1946 585
R17474 GND.t40 GND.n1947 585
R17475 GND.n8268 GND.n8267 585
R17476 GND.n8269 GND.n8268 585
R17477 GND.n1963 GND.n1962 585
R17478 GND.n4196 GND.n1962 585
R17479 GND.n8262 GND.n8261 585
R17480 GND.n8261 GND.n8260 585
R17481 GND.n1983 GND.n1966 585
R17482 GND.n2050 GND.n1966 585
R17483 GND.n8251 GND.n8250 585
R17484 GND.n8252 GND.n8251 585
R17485 GND.n8249 GND.n1982 585
R17486 GND.n8174 GND.n1982 585
R17487 GND.n8248 GND.n8247 585
R17488 GND.n8247 GND.n8246 585
R17489 GND.n1986 GND.n1985 585
R17490 GND.n8204 GND.n1986 585
R17491 GND.n4439 GND.n4438 585
R17492 GND.n4440 GND.n4439 585
R17493 GND.n4436 GND.n4411 585
R17494 GND.n4435 GND.n4434 585
R17495 GND.n4433 GND.n4432 585
R17496 GND.n4431 GND.n4430 585
R17497 GND.n4429 GND.n4428 585
R17498 GND.n4427 GND.n4426 585
R17499 GND.n4425 GND.n4424 585
R17500 GND.n4423 GND.n4422 585
R17501 GND.n4421 GND.n4420 585
R17502 GND.n4419 GND.n4418 585
R17503 GND.n4417 GND.n4416 585
R17504 GND.n4415 GND.n4414 585
R17505 GND.n4413 GND.n4412 585
R17506 GND.n4269 GND.n4268 585
R17507 GND.n4443 GND.n4442 585
R17508 GND.n4444 GND.n4267 585
R17509 GND.n4447 GND.n4446 585
R17510 GND.n4448 GND.n4447 585
R17511 GND.n4445 GND.n1920 585
R17512 GND.n8298 GND.n1920 585
R17513 GND.n1931 GND.n1929 585
R17514 GND.n4503 GND.n1929 585
R17515 GND.n8291 GND.n8290 585
R17516 GND.n8292 GND.n8291 585
R17517 GND.n1932 GND.n1930 585
R17518 GND.n4683 GND.n1930 585
R17519 GND.n8286 GND.n8285 585
R17520 GND.n8285 GND.n8284 585
R17521 GND.n1953 GND.n1935 585
R17522 GND.n4492 GND.n1935 585
R17523 GND.n8274 GND.n8273 585
R17524 GND.n8275 GND.n8274 585
R17525 GND.n8272 GND.n1952 585
R17526 GND.t40 GND.n1952 585
R17527 GND.n8271 GND.n8270 585
R17528 GND.n8270 GND.n8269 585
R17529 GND.n1972 GND.n1957 585
R17530 GND.n4196 GND.n1957 585
R17531 GND.n8259 GND.n8258 585
R17532 GND.n8260 GND.n8259 585
R17533 GND.n1974 GND.n1971 585
R17534 GND.n2050 GND.n1971 585
R17535 GND.n8254 GND.n8253 585
R17536 GND.n8253 GND.n8252 585
R17537 GND.n1977 GND.n1976 585
R17538 GND.n8174 GND.n1977 585
R17539 GND.n8245 GND.n8244 585
R17540 GND.n8246 GND.n8245 585
R17541 GND.n8243 GND.n1990 585
R17542 GND.n8204 GND.n1990 585
R17543 GND.n8242 GND.n8241 585
R17544 GND.n1992 GND.n1991 585
R17545 GND.n4727 GND.n4726 585
R17546 GND.n4729 GND.n4728 585
R17547 GND.n4731 GND.n4730 585
R17548 GND.n4733 GND.n4732 585
R17549 GND.n4735 GND.n4734 585
R17550 GND.n4737 GND.n4736 585
R17551 GND.n4739 GND.n4738 585
R17552 GND.n4741 GND.n4740 585
R17553 GND.n4743 GND.n4742 585
R17554 GND.n4745 GND.n4744 585
R17555 GND.n4747 GND.n4746 585
R17556 GND.n4749 GND.n4748 585
R17557 GND.n4751 GND.n4750 585
R17558 GND.n4753 GND.n4752 585
R17559 GND.n4754 GND.n2008 585
R17560 GND.n8239 GND.n2008 585
R17561 GND.n4755 GND.n2014 585
R17562 GND.n8204 GND.n2014 585
R17563 GND.n4756 GND.n1988 585
R17564 GND.n8246 GND.n1988 585
R17565 GND.n4757 GND.n2041 585
R17566 GND.n8174 GND.n2041 585
R17567 GND.n4758 GND.n1980 585
R17568 GND.n8252 GND.n1980 585
R17569 GND.n4761 GND.n4760 585
R17570 GND.n4760 GND.n2050 585
R17571 GND.n4763 GND.n1969 585
R17572 GND.n8260 GND.n1969 585
R17573 GND.n4725 GND.n4724 585
R17574 GND.n4724 GND.n4196 585
R17575 GND.n4722 GND.n1960 585
R17576 GND.n8269 GND.n1960 585
R17577 GND.n4721 GND.n4205 585
R17578 GND.t40 GND.n4205 585
R17579 GND.n4204 GND.n1950 585
R17580 GND.n8275 GND.n1950 585
R17581 GND.n4494 GND.n4493 585
R17582 GND.n4493 GND.n4492 585
R17583 GND.n4496 GND.n1938 585
R17584 GND.n8284 GND.n1938 585
R17585 GND.n4255 GND.n4215 585
R17586 GND.n4683 GND.n4215 585
R17587 GND.n4500 GND.n1928 585
R17588 GND.n8292 GND.n1928 585
R17589 GND.n4502 GND.n4501 585
R17590 GND.n4503 GND.n4502 585
R17591 GND.n4254 GND.n1919 585
R17592 GND.n8298 GND.n1919 585
R17593 GND.n4437 GND.n4266 585
R17594 GND.n4448 GND.n4266 585
R17595 GND.n4345 GND.n4344 585
R17596 GND.n4346 GND.n4345 585
R17597 GND.n4343 GND.n4335 585
R17598 GND.n4335 GND.n1895 585
R17599 GND.n4338 GND.n4337 585
R17600 GND.n4337 GND.n1896 585
R17601 GND.n4339 GND.n1908 585
R17602 GND.n4357 GND.n1908 585
R17603 GND.n8307 GND.n8306 585
R17604 GND.n8308 GND.n8307 585
R17605 GND.n1911 GND.n1909 585
R17606 GND.n4449 GND.n1909 585
R17607 GND.n8301 GND.n8300 585
R17608 GND.n8300 GND.n8299 585
R17609 GND.n4474 GND.n1915 585
R17610 GND.n4504 GND.n1915 585
R17611 GND.n4478 GND.n4477 585
R17612 GND.n4478 GND.n1926 585
R17613 GND.n4480 GND.n4479 585
R17614 GND.n4479 GND.n4214 585
R17615 GND.n4481 GND.n4470 585
R17616 GND.n4470 GND.n1936 585
R17617 GND.n4489 GND.n4488 585
R17618 GND.n4490 GND.n4489 585
R17619 GND.n4209 GND.n4207 585
R17620 GND.n4209 GND.n1948 585
R17621 GND.n4716 GND.n4715 585
R17622 GND.n4715 GND.n4714 585
R17623 GND.n4208 GND.n4197 585
R17624 GND.n4197 GND.n1958 585
R17625 GND.n4770 GND.n4769 585
R17626 GND.n4771 GND.n4770 585
R17627 GND.n4200 GND.n4198 585
R17628 GND.n4198 GND.n1967 585
R17629 GND.n4646 GND.n4645 585
R17630 GND.n4647 GND.n4646 585
R17631 GND.n4642 GND.n2038 585
R17632 GND.n2038 GND.n1978 585
R17633 GND.n8177 GND.n8176 585
R17634 GND.n8176 GND.n8175 585
R17635 GND.n2035 GND.n2034 585
R17636 GND.n2043 GND.n2034 585
R17637 GND.n8183 GND.n8182 585
R17638 GND.n8183 GND.n2013 585
R17639 GND.n8185 GND.n8184 585
R17640 GND.n8184 GND.n2016 585
R17641 GND.n8186 GND.n2028 585
R17642 GND.n2028 GND.n2009 585
R17643 GND.n8192 GND.n8191 585
R17644 GND.n8193 GND.n8192 585
R17645 GND.n2031 GND.n2029 585
R17646 GND.n2063 GND.n2029 585
R17647 GND.n2077 GND.n2076 585
R17648 GND.n2076 GND.n2064 585
R17649 GND.n4619 GND.n4558 585
R17650 GND.n4619 GND.n2064 585
R17651 GND.n4621 GND.n4620 585
R17652 GND.n4620 GND.n2063 585
R17653 GND.n4623 GND.n2026 585
R17654 GND.n8193 GND.n2026 585
R17655 GND.n4626 GND.n4625 585
R17656 GND.n4625 GND.n2009 585
R17657 GND.n4556 GND.n4555 585
R17658 GND.n4555 GND.n2016 585
R17659 GND.n4632 GND.n4631 585
R17660 GND.n4632 GND.n2013 585
R17661 GND.n4634 GND.n4633 585
R17662 GND.n4633 GND.n2043 585
R17663 GND.n4551 GND.n2039 585
R17664 GND.n8175 GND.n2039 585
R17665 GND.n4640 GND.n4639 585
R17666 GND.n4640 GND.n1978 585
R17667 GND.n4649 GND.n4648 585
R17668 GND.n4648 GND.n4647 585
R17669 GND.n4651 GND.n4194 585
R17670 GND.n4194 GND.n1967 585
R17671 GND.n4772 GND.n4195 585
R17672 GND.n4772 GND.n4771 585
R17673 GND.n4774 GND.n4773 585
R17674 GND.n4773 GND.n1958 585
R17675 GND.n4775 GND.n4192 585
R17676 GND.n4714 GND.n4192 585
R17677 GND.n4259 GND.n4191 585
R17678 GND.n4259 GND.n1948 585
R17679 GND.n4469 GND.n4468 585
R17680 GND.n4490 GND.n4469 585
R17681 GND.n4465 GND.n4258 585
R17682 GND.n4258 GND.n1936 585
R17683 GND.n4458 GND.n4260 585
R17684 GND.n4458 GND.n4214 585
R17685 GND.n4460 GND.n4459 585
R17686 GND.n4459 GND.n1926 585
R17687 GND.n4456 GND.n4252 585
R17688 GND.n4504 GND.n4252 585
R17689 GND.n4262 GND.n1917 585
R17690 GND.n8299 GND.n1917 585
R17691 GND.n4451 GND.n4450 585
R17692 GND.n4450 GND.n4449 585
R17693 GND.n4273 GND.n1906 585
R17694 GND.n8308 GND.n1906 585
R17695 GND.n4356 GND.n4355 585
R17696 GND.n4357 GND.n4356 585
R17697 GND.n4350 GND.n4271 585
R17698 GND.n4271 GND.n1896 585
R17699 GND.n4349 GND.n4348 585
R17700 GND.n4348 GND.n1895 585
R17701 GND.n4347 GND.n4274 585
R17702 GND.n4347 GND.n4346 585
R17703 GND.n8328 GND.n8327 585
R17704 GND.n8327 GND.n8326 585
R17705 GND.n1898 GND.n1870 585
R17706 GND.n4333 GND.n1870 585
R17707 GND.n8317 GND.n8316 585
R17708 GND.n8318 GND.n8317 585
R17709 GND.n1900 GND.n1897 585
R17710 GND.n4270 GND.n1897 585
R17711 GND.n8311 GND.n8310 585
R17712 GND.n8310 GND.n8309 585
R17713 GND.n4510 GND.n1904 585
R17714 GND.n1907 GND.n1904 585
R17715 GND.n4513 GND.n4512 585
R17716 GND.n4512 GND.n1916 585
R17717 GND.n4514 GND.n4506 585
R17718 GND.n4506 GND.n4505 585
R17719 GND.n4521 GND.n4520 585
R17720 GND.n4522 GND.n4521 585
R17721 GND.n4508 GND.n4217 585
R17722 GND.n4524 GND.n4217 585
R17723 GND.n4681 GND.n4680 585
R17724 GND.n4682 GND.n4681 585
R17725 GND.n4220 GND.n4218 585
R17726 GND.n4218 GND.n1939 585
R17727 GND.n4674 GND.n4673 585
R17728 GND.n4673 GND.n4672 585
R17729 GND.n4542 GND.n4225 585
R17730 GND.n4225 GND.n1951 585
R17731 GND.n4544 GND.n4543 585
R17732 GND.n4543 GND.n4210 585
R17733 GND.n4546 GND.n4541 585
R17734 GND.n4541 GND.n1961 585
R17735 GND.n4660 GND.n4659 585
R17736 GND.n4661 GND.n4660 585
R17737 GND.n4548 GND.n2049 585
R17738 GND.n2049 GND.n1970 585
R17739 GND.n8164 GND.n8163 585
R17740 GND.n8163 GND.n8162 585
R17741 GND.n8165 GND.n2044 585
R17742 GND.n2044 GND.n1981 585
R17743 GND.n8172 GND.n8171 585
R17744 GND.n8173 GND.n8172 585
R17745 GND.n2046 GND.n2017 585
R17746 GND.n2017 GND.n1989 585
R17747 GND.n8202 GND.n8201 585
R17748 GND.n8203 GND.n8202 585
R17749 GND.n2020 GND.n2018 585
R17750 GND.n2018 GND.n1993 585
R17751 GND.n8196 GND.n8195 585
R17752 GND.n8195 GND.n8194 585
R17753 GND.n2066 GND.n2024 585
R17754 GND.n2027 GND.n2024 585
R17755 GND.n8136 GND.n8135 585
R17756 GND.n8137 GND.n8136 585
R17757 GND.n8132 GND.n2065 585
R17758 GND.n2112 GND.n2065 585
R17759 GND.n8042 GND.n2062 585
R17760 GND.n2112 GND.n2062 585
R17761 GND.n8139 GND.n8138 585
R17762 GND.n8138 GND.n8137 585
R17763 GND.n2061 GND.n2059 585
R17764 GND.n2061 GND.n2027 585
R17765 GND.n8144 GND.n2025 585
R17766 GND.n8194 GND.n2025 585
R17767 GND.n8147 GND.n8146 585
R17768 GND.n8146 GND.n1993 585
R17769 GND.n2057 GND.n2015 585
R17770 GND.n8203 GND.n2015 585
R17771 GND.n8153 GND.n8152 585
R17772 GND.n8152 GND.n1989 585
R17773 GND.n8155 GND.n2042 585
R17774 GND.n8173 GND.n2042 585
R17775 GND.n2054 GND.n2052 585
R17776 GND.n2052 GND.n1981 585
R17777 GND.n8161 GND.n8160 585
R17778 GND.n8162 GND.n8161 585
R17779 GND.n4537 GND.n2051 585
R17780 GND.n2051 GND.n1970 585
R17781 GND.n4662 GND.n4540 585
R17782 GND.n4662 GND.n4661 585
R17783 GND.n4664 GND.n4663 585
R17784 GND.n4663 GND.n1961 585
R17785 GND.n4536 GND.n4534 585
R17786 GND.n4536 GND.n4210 585
R17787 GND.n4229 GND.n4227 585
R17788 GND.n4227 GND.n1951 585
R17789 GND.n4671 GND.n4670 585
R17790 GND.n4672 GND.n4671 585
R17791 GND.n4529 GND.n4226 585
R17792 GND.n4226 GND.n1939 585
R17793 GND.n4528 GND.n4216 585
R17794 GND.n4682 GND.n4216 585
R17795 GND.n4526 GND.n4525 585
R17796 GND.n4525 GND.n4524 585
R17797 GND.n4523 GND.n4251 585
R17798 GND.n4523 GND.n4522 585
R17799 GND.n4233 GND.n4232 585
R17800 GND.n4505 GND.n4232 585
R17801 GND.n4245 GND.n4244 585
R17802 GND.n4244 GND.n1916 585
R17803 GND.n4243 GND.n4242 585
R17804 GND.n4243 GND.n1907 585
R17805 GND.n4236 GND.n1905 585
R17806 GND.n8309 GND.n1905 585
R17807 GND.n4237 GND.n1894 585
R17808 GND.n4270 GND.n1894 585
R17809 GND.n8320 GND.n8319 585
R17810 GND.n8319 GND.n8318 585
R17811 GND.n1891 GND.n1873 585
R17812 GND.n4333 GND.n1873 585
R17813 GND.n8325 GND.n8324 585
R17814 GND.n8326 GND.n8325 585
R17815 GND.n3566 GND.n3400 585
R17816 GND.n3565 GND.n3564 585
R17817 GND.n3562 GND.n3401 585
R17818 GND.n3560 GND.n3559 585
R17819 GND.n3558 GND.n3402 585
R17820 GND.n3557 GND.n3556 585
R17821 GND.n3554 GND.n3403 585
R17822 GND.n3552 GND.n3551 585
R17823 GND.n3550 GND.n3404 585
R17824 GND.n3549 GND.n3548 585
R17825 GND.n3546 GND.n3405 585
R17826 GND.n3544 GND.n3543 585
R17827 GND.n3542 GND.n3406 585
R17828 GND.n3541 GND.n3540 585
R17829 GND.n3538 GND.n3407 585
R17830 GND.n3536 GND.n3535 585
R17831 GND.n3534 GND.n3408 585
R17832 GND.n3533 GND.n3532 585
R17833 GND.n3530 GND.n3336 585
R17834 GND.n3569 GND.n3336 585
R17835 GND.n3529 GND.n3528 585
R17836 GND.n3528 GND.n3331 585
R17837 GND.n3527 GND.n3330 585
R17838 GND.n3575 GND.n3330 585
R17839 GND.n3526 GND.n3525 585
R17840 GND.n3525 GND.n3325 585
R17841 GND.n3524 GND.n3324 585
R17842 GND.n3581 GND.n3324 585
R17843 GND.n3523 GND.n3522 585
R17844 GND.n3522 GND.n3319 585
R17845 GND.n3521 GND.n3318 585
R17846 GND.n3587 GND.n3318 585
R17847 GND.n3520 GND.n3519 585
R17848 GND.n3519 GND.n3313 585
R17849 GND.n3518 GND.n3312 585
R17850 GND.n3593 GND.n3312 585
R17851 GND.n3517 GND.n3516 585
R17852 GND.n3516 GND.n3307 585
R17853 GND.n3515 GND.n3306 585
R17854 GND.n3599 GND.n3306 585
R17855 GND.n3514 GND.n3513 585
R17856 GND.n3513 GND.n3298 585
R17857 GND.n3512 GND.n3297 585
R17858 GND.n3605 GND.n3297 585
R17859 GND.n3511 GND.n3510 585
R17860 GND.n3510 GND.n3291 585
R17861 GND.n3509 GND.n3290 585
R17862 GND.n3611 GND.n3290 585
R17863 GND.n3508 GND.n3507 585
R17864 GND.n3507 GND.n3283 585
R17865 GND.n3409 GND.n3282 585
R17866 GND.n3617 GND.n3282 585
R17867 GND.n3489 GND.n3488 585
R17868 GND.n3488 GND.n3276 585
R17869 GND.n3492 GND.n3275 585
R17870 GND.n3623 GND.n3275 585
R17871 GND.n3494 GND.n3493 585
R17872 GND.n3493 GND.n3269 585
R17873 GND.n3495 GND.n3268 585
R17874 GND.n3629 GND.n3268 585
R17875 GND.n3497 GND.n3496 585
R17876 GND.n3496 GND.t151 585
R17877 GND.n3486 GND.n3262 585
R17878 GND.n3635 GND.n3262 585
R17879 GND.n3484 GND.n3483 585
R17880 GND.n3483 GND.n3196 585
R17881 GND.n3480 GND.n3195 585
R17882 GND.n3641 GND.n3195 585
R17883 GND.n3479 GND.n3478 585
R17884 GND.n3478 GND.n3190 585
R17885 GND.n3477 GND.n3189 585
R17886 GND.n3647 GND.n3189 585
R17887 GND.n3476 GND.n3475 585
R17888 GND.n3475 GND.n3184 585
R17889 GND.n3474 GND.n3183 585
R17890 GND.n3653 GND.n3183 585
R17891 GND.n3473 GND.n3472 585
R17892 GND.n3472 GND.n3178 585
R17893 GND.n3471 GND.n3177 585
R17894 GND.n3659 GND.n3177 585
R17895 GND.n3470 GND.n3469 585
R17896 GND.n3469 GND.n3172 585
R17897 GND.n3468 GND.n3171 585
R17898 GND.n3665 GND.n3171 585
R17899 GND.n3467 GND.n3466 585
R17900 GND.n3466 GND.n3166 585
R17901 GND.n3465 GND.n3165 585
R17902 GND.n3671 GND.n3165 585
R17903 GND.n3464 GND.n3463 585
R17904 GND.n3463 GND.n3160 585
R17905 GND.n3462 GND.n3159 585
R17906 GND.n3677 GND.n3159 585
R17907 GND.n3461 GND.n3460 585
R17908 GND.n3460 GND.n3154 585
R17909 GND.n3459 GND.n3153 585
R17910 GND.n3683 GND.n3153 585
R17911 GND.n3458 GND.n3457 585
R17912 GND.n3457 GND.n3146 585
R17913 GND.n3456 GND.n3145 585
R17914 GND.n3689 GND.n3145 585
R17915 GND.n3455 GND.n3454 585
R17916 GND.n3454 GND.n3137 585
R17917 GND.n3453 GND.n3136 585
R17918 GND.n3695 GND.n3136 585
R17919 GND.n3452 GND.n3451 585
R17920 GND.n3450 GND.n3449 585
R17921 GND.n3448 GND.n3447 585
R17922 GND.n3446 GND.n3445 585
R17923 GND.n3444 GND.n3443 585
R17924 GND.n3442 GND.n3441 585
R17925 GND.n3440 GND.n3439 585
R17926 GND.n3438 GND.n3437 585
R17927 GND.n3436 GND.n3435 585
R17928 GND.n3434 GND.n3433 585
R17929 GND.n3432 GND.n3431 585
R17930 GND.n3430 GND.n3429 585
R17931 GND.n3428 GND.n3427 585
R17932 GND.n3426 GND.n3425 585
R17933 GND.n3424 GND.n3423 585
R17934 GND.n3422 GND.n3421 585
R17935 GND.n3420 GND.n3419 585
R17936 GND.n3418 GND.n3417 585
R17937 GND.n3416 GND.n3138 585
R17938 GND.n3695 GND.n3138 585
R17939 GND.n3149 GND.n3147 585
R17940 GND.n3147 GND.n3137 585
R17941 GND.n3688 GND.n3687 585
R17942 GND.n3689 GND.n3688 585
R17943 GND.n3686 GND.n3148 585
R17944 GND.n3148 GND.n3146 585
R17945 GND.n3685 GND.n3684 585
R17946 GND.n3684 GND.n3683 585
R17947 GND.n3151 GND.n3150 585
R17948 GND.n3154 GND.n3151 585
R17949 GND.n3676 GND.n3675 585
R17950 GND.n3677 GND.n3676 585
R17951 GND.n3674 GND.n3161 585
R17952 GND.n3161 GND.n3160 585
R17953 GND.n3673 GND.n3672 585
R17954 GND.n3672 GND.n3671 585
R17955 GND.n3163 GND.n3162 585
R17956 GND.n3166 GND.n3163 585
R17957 GND.n3664 GND.n3663 585
R17958 GND.n3665 GND.n3664 585
R17959 GND.n3662 GND.n3173 585
R17960 GND.n3173 GND.n3172 585
R17961 GND.n3661 GND.n3660 585
R17962 GND.n3660 GND.n3659 585
R17963 GND.n3175 GND.n3174 585
R17964 GND.n3178 GND.n3175 585
R17965 GND.n3652 GND.n3651 585
R17966 GND.n3653 GND.n3652 585
R17967 GND.n3650 GND.n3185 585
R17968 GND.n3185 GND.n3184 585
R17969 GND.n3649 GND.n3648 585
R17970 GND.n3648 GND.n3647 585
R17971 GND.n3187 GND.n3186 585
R17972 GND.n3190 GND.n3187 585
R17973 GND.n3640 GND.n3639 585
R17974 GND.n3641 GND.n3640 585
R17975 GND.n3638 GND.n3197 585
R17976 GND.n3197 GND.n3196 585
R17977 GND.n3263 GND.n3260 585
R17978 GND.n3635 GND.n3263 585
R17979 GND.n3272 GND.n3270 585
R17980 GND.n3270 GND.t151 585
R17981 GND.n3628 GND.n3627 585
R17982 GND.n3629 GND.n3628 585
R17983 GND.n3626 GND.n3271 585
R17984 GND.n3271 GND.n3269 585
R17985 GND.n3277 GND.n3273 585
R17986 GND.n3623 GND.n3277 585
R17987 GND.n3286 GND.n3284 585
R17988 GND.n3284 GND.n3276 585
R17989 GND.n3616 GND.n3615 585
R17990 GND.n3617 GND.n3616 585
R17991 GND.n3614 GND.n3285 585
R17992 GND.n3285 GND.n3283 585
R17993 GND.n3301 GND.n3292 585
R17994 GND.n3611 GND.n3292 585
R17995 GND.n3302 GND.n3299 585
R17996 GND.n3299 GND.n3291 585
R17997 GND.n3604 GND.n3603 585
R17998 GND.n3605 GND.n3604 585
R17999 GND.n3602 GND.n3300 585
R18000 GND.n3300 GND.n3298 585
R18001 GND.n3601 GND.n3600 585
R18002 GND.n3600 GND.n3599 585
R18003 GND.n3304 GND.n3303 585
R18004 GND.n3307 GND.n3304 585
R18005 GND.n3592 GND.n3591 585
R18006 GND.n3593 GND.n3592 585
R18007 GND.n3590 GND.n3314 585
R18008 GND.n3314 GND.n3313 585
R18009 GND.n3589 GND.n3588 585
R18010 GND.n3588 GND.n3587 585
R18011 GND.n3316 GND.n3315 585
R18012 GND.n3319 GND.n3316 585
R18013 GND.n3580 GND.n3579 585
R18014 GND.n3581 GND.n3580 585
R18015 GND.n3578 GND.n3326 585
R18016 GND.n3326 GND.n3325 585
R18017 GND.n3577 GND.n3576 585
R18018 GND.n3576 GND.n3575 585
R18019 GND.n3328 GND.n3327 585
R18020 GND.n3331 GND.n3328 585
R18021 GND.n3568 GND.n3567 585
R18022 GND.n3569 GND.n3568 585
R18023 GND.n1721 GND.n1720 585
R18024 GND.n1719 GND.n1662 585
R18025 GND.n1718 GND.n1717 585
R18026 GND.n1716 GND.n1715 585
R18027 GND.n1714 GND.n1713 585
R18028 GND.n1712 GND.n1711 585
R18029 GND.n1710 GND.n1709 585
R18030 GND.n1708 GND.n1707 585
R18031 GND.n1706 GND.n1705 585
R18032 GND.n1704 GND.n1703 585
R18033 GND.n1702 GND.n1701 585
R18034 GND.n1700 GND.n1699 585
R18035 GND.n1698 GND.n1697 585
R18036 GND.n1696 GND.n1695 585
R18037 GND.n1694 GND.n1693 585
R18038 GND.n1692 GND.n1691 585
R18039 GND.n1690 GND.n1689 585
R18040 GND.n1688 GND.n1687 585
R18041 GND.n1686 GND.n1685 585
R18042 GND.n1686 GND.n1059 585
R18043 GND.n1684 GND.n1058 585
R18044 GND.n8735 GND.n1058 585
R18045 GND.n1683 GND.n1682 585
R18046 GND.n1682 GND.n1053 585
R18047 GND.n1681 GND.n1052 585
R18048 GND.n8741 GND.n1052 585
R18049 GND.n1680 GND.n1679 585
R18050 GND.n1679 GND.n1047 585
R18051 GND.n1678 GND.n1046 585
R18052 GND.n8747 GND.n1046 585
R18053 GND.n1677 GND.n1676 585
R18054 GND.n1676 GND.n1041 585
R18055 GND.n1675 GND.n1040 585
R18056 GND.n8753 GND.n1040 585
R18057 GND.n1674 GND.n1673 585
R18058 GND.n1673 GND.n1035 585
R18059 GND.n1672 GND.n1034 585
R18060 GND.n8759 GND.n1034 585
R18061 GND.n1671 GND.n1670 585
R18062 GND.n1670 GND.n1029 585
R18063 GND.n1669 GND.n1028 585
R18064 GND.n8765 GND.n1028 585
R18065 GND.n1668 GND.n1667 585
R18066 GND.n1667 GND.n1023 585
R18067 GND.n1666 GND.n1022 585
R18068 GND.n8771 GND.n1022 585
R18069 GND.n1665 GND.n1664 585
R18070 GND.n1664 GND.n1015 585
R18071 GND.n1663 GND.n1014 585
R18072 GND.n8777 GND.n1014 585
R18073 GND.n1003 GND.n1001 585
R18074 GND.n1006 GND.n1003 585
R18075 GND.n8785 GND.n8784 585
R18076 GND.n8784 GND.n8783 585
R18077 GND.n1002 GND.n1000 585
R18078 GND.n1004 GND.n1002 585
R18079 GND.n8517 GND.n1728 585
R18080 GND.n8666 GND.n1728 585
R18081 GND.n8521 GND.n8520 585
R18082 GND.n8520 GND.n1727 585
R18083 GND.n8522 GND.n1735 585
R18084 GND.t6 GND.n1735 585
R18085 GND.n8524 GND.n8523 585
R18086 GND.n8523 GND.n1733 585
R18087 GND.n8525 GND.n1741 585
R18088 GND.n8653 GND.n1741 585
R18089 GND.n8515 GND.n8514 585
R18090 GND.n8514 GND.n1739 585
R18091 GND.n8511 GND.n1747 585
R18092 GND.n8647 GND.n1747 585
R18093 GND.n8534 GND.n8533 585
R18094 GND.n8533 GND.n1745 585
R18095 GND.n8535 GND.n1753 585
R18096 GND.n8639 GND.n1753 585
R18097 GND.n8537 GND.n8536 585
R18098 GND.n8536 GND.n1752 585
R18099 GND.n8538 GND.n1760 585
R18100 GND.n8633 GND.n1760 585
R18101 GND.n8540 GND.n8539 585
R18102 GND.n8539 GND.n1758 585
R18103 GND.n8541 GND.n1767 585
R18104 GND.n8625 GND.n1767 585
R18105 GND.n8543 GND.n8542 585
R18106 GND.n8542 GND.n1765 585
R18107 GND.n8544 GND.n1773 585
R18108 GND.n8619 GND.n1773 585
R18109 GND.n8546 GND.n8545 585
R18110 GND.n8545 GND.n1771 585
R18111 GND.n8547 GND.n1779 585
R18112 GND.n8613 GND.n1779 585
R18113 GND.n8549 GND.n8548 585
R18114 GND.n8548 GND.n1777 585
R18115 GND.n8550 GND.n1785 585
R18116 GND.n8607 GND.n1785 585
R18117 GND.n8552 GND.n8551 585
R18118 GND.n8551 GND.n1783 585
R18119 GND.n8553 GND.n1791 585
R18120 GND.n8601 GND.n1791 585
R18121 GND.n8555 GND.n8554 585
R18122 GND.n8554 GND.n1789 585
R18123 GND.n8556 GND.n1797 585
R18124 GND.n8595 GND.n1797 585
R18125 GND.n8559 GND.n8557 585
R18126 GND.n8559 GND.n1795 585
R18127 GND.n8561 GND.n8560 585
R18128 GND.n8562 GND.n8510 585
R18129 GND.n8564 GND.n8563 585
R18130 GND.n8566 GND.n8508 585
R18131 GND.n8568 GND.n8567 585
R18132 GND.n8569 GND.n8507 585
R18133 GND.n8571 GND.n8570 585
R18134 GND.n8573 GND.n8505 585
R18135 GND.n8575 GND.n8574 585
R18136 GND.n8576 GND.n8504 585
R18137 GND.n8578 GND.n8577 585
R18138 GND.n8580 GND.n8502 585
R18139 GND.n8582 GND.n8581 585
R18140 GND.n8583 GND.n8501 585
R18141 GND.n8585 GND.n8584 585
R18142 GND.n8587 GND.n8500 585
R18143 GND.n8588 GND.n1799 585
R18144 GND.n8591 GND.n8590 585
R18145 GND.n8592 GND.n1798 585
R18146 GND.n1798 GND.n1795 585
R18147 GND.n8594 GND.n8593 585
R18148 GND.n8595 GND.n8594 585
R18149 GND.n1788 GND.n1787 585
R18150 GND.n1789 GND.n1788 585
R18151 GND.n8603 GND.n8602 585
R18152 GND.n8602 GND.n8601 585
R18153 GND.n8604 GND.n1786 585
R18154 GND.n1786 GND.n1783 585
R18155 GND.n8606 GND.n8605 585
R18156 GND.n8607 GND.n8606 585
R18157 GND.n1776 GND.n1775 585
R18158 GND.n1777 GND.n1776 585
R18159 GND.n8615 GND.n8614 585
R18160 GND.n8614 GND.n8613 585
R18161 GND.n8616 GND.n1774 585
R18162 GND.n1774 GND.n1771 585
R18163 GND.n8618 GND.n8617 585
R18164 GND.n8619 GND.n8618 585
R18165 GND.n1764 GND.n1763 585
R18166 GND.n1765 GND.n1764 585
R18167 GND.n8627 GND.n8626 585
R18168 GND.n8626 GND.n8625 585
R18169 GND.n8628 GND.n1761 585
R18170 GND.n1761 GND.n1758 585
R18171 GND.n8632 GND.n8631 585
R18172 GND.n8633 GND.n8632 585
R18173 GND.n8630 GND.n1762 585
R18174 GND.n1762 GND.n1752 585
R18175 GND.n8629 GND.n1754 585
R18176 GND.n8639 GND.n1754 585
R18177 GND.n8642 GND.n1748 585
R18178 GND.n1748 GND.n1745 585
R18179 GND.n8646 GND.n8645 585
R18180 GND.n8647 GND.n8646 585
R18181 GND.n8644 GND.n1738 585
R18182 GND.n1739 GND.n1738 585
R18183 GND.n8654 GND.n1737 585
R18184 GND.n8654 GND.n8653 585
R18185 GND.n8656 GND.n8655 585
R18186 GND.n8655 GND.n1733 585
R18187 GND.n8659 GND.n1734 585
R18188 GND.t6 GND.n1734 585
R18189 GND.n8658 GND.n8657 585
R18190 GND.n8657 GND.n1727 585
R18191 GND.n1729 GND.n1724 585
R18192 GND.n8666 GND.n1729 585
R18193 GND.n8669 GND.n1725 585
R18194 GND.n1725 GND.n1004 585
R18195 GND.n8670 GND.n1007 585
R18196 GND.n8783 GND.n1007 585
R18197 GND.n1018 GND.n1016 585
R18198 GND.n1016 GND.n1006 585
R18199 GND.n8776 GND.n8775 585
R18200 GND.n8777 GND.n8776 585
R18201 GND.n8774 GND.n1017 585
R18202 GND.n1017 GND.n1015 585
R18203 GND.n8773 GND.n8772 585
R18204 GND.n8772 GND.n8771 585
R18205 GND.n1020 GND.n1019 585
R18206 GND.n1023 GND.n1020 585
R18207 GND.n8764 GND.n8763 585
R18208 GND.n8765 GND.n8764 585
R18209 GND.n8762 GND.n1030 585
R18210 GND.n1030 GND.n1029 585
R18211 GND.n8761 GND.n8760 585
R18212 GND.n8760 GND.n8759 585
R18213 GND.n1032 GND.n1031 585
R18214 GND.n1035 GND.n1032 585
R18215 GND.n8752 GND.n8751 585
R18216 GND.n8753 GND.n8752 585
R18217 GND.n8750 GND.n1042 585
R18218 GND.n1042 GND.n1041 585
R18219 GND.n8749 GND.n8748 585
R18220 GND.n8748 GND.n8747 585
R18221 GND.n1044 GND.n1043 585
R18222 GND.n1047 GND.n1044 585
R18223 GND.n8740 GND.n8739 585
R18224 GND.n8741 GND.n8740 585
R18225 GND.n8738 GND.n1054 585
R18226 GND.n1054 GND.n1053 585
R18227 GND.n8737 GND.n8736 585
R18228 GND.n8736 GND.n8735 585
R18229 GND.n1056 GND.n1055 585
R18230 GND.n1059 GND.n1056 585
R18231 GND.n3334 GND.n3333 585
R18232 GND.n3397 GND.n3396 585
R18233 GND.n3395 GND.n3345 585
R18234 GND.n3399 GND.n3345 585
R18235 GND.n3394 GND.n3393 585
R18236 GND.n3392 GND.n3391 585
R18237 GND.n3390 GND.n3389 585
R18238 GND.n3388 GND.n3387 585
R18239 GND.n3386 GND.n3385 585
R18240 GND.n3384 GND.n3383 585
R18241 GND.n3382 GND.n3381 585
R18242 GND.n3380 GND.n3379 585
R18243 GND.n3378 GND.n3377 585
R18244 GND.n3376 GND.n3375 585
R18245 GND.n3374 GND.n3373 585
R18246 GND.n3372 GND.n3371 585
R18247 GND.n3370 GND.n3369 585
R18248 GND.n3368 GND.n3367 585
R18249 GND.n3366 GND.n3344 585
R18250 GND.n3399 GND.n3344 585
R18251 GND.n3365 GND.n3335 585
R18252 GND.n3569 GND.n3335 585
R18253 GND.n3364 GND.n3363 585
R18254 GND.n3363 GND.n3331 585
R18255 GND.n3362 GND.n3329 585
R18256 GND.n3575 GND.n3329 585
R18257 GND.n3361 GND.n3360 585
R18258 GND.n3360 GND.n3325 585
R18259 GND.n3359 GND.n3323 585
R18260 GND.n3581 GND.n3323 585
R18261 GND.n3358 GND.n3357 585
R18262 GND.n3357 GND.n3319 585
R18263 GND.n3356 GND.n3317 585
R18264 GND.n3587 GND.n3317 585
R18265 GND.n3355 GND.n3354 585
R18266 GND.n3354 GND.n3313 585
R18267 GND.n3353 GND.n3311 585
R18268 GND.n3593 GND.n3311 585
R18269 GND.n3352 GND.n3351 585
R18270 GND.n3351 GND.n3307 585
R18271 GND.n3350 GND.n3305 585
R18272 GND.n3599 GND.n3305 585
R18273 GND.n3349 GND.n3348 585
R18274 GND.n3348 GND.n3298 585
R18275 GND.n3347 GND.n3296 585
R18276 GND.n3605 GND.n3296 585
R18277 GND.n3346 GND.n3288 585
R18278 GND.n3291 GND.n3288 585
R18279 GND.n3612 GND.n3289 585
R18280 GND.n3612 GND.n3611 585
R18281 GND.n3614 GND.n3613 585
R18282 GND.n3613 GND.n3283 585
R18283 GND.n3615 GND.n3281 585
R18284 GND.n3617 GND.n3281 585
R18285 GND.n3286 GND.n3274 585
R18286 GND.n3276 GND.n3274 585
R18287 GND.n3624 GND.n3273 585
R18288 GND.n3624 GND.n3623 585
R18289 GND.n3626 GND.n3625 585
R18290 GND.n3625 GND.n3269 585
R18291 GND.n3627 GND.n3267 585
R18292 GND.n3629 GND.n3267 585
R18293 GND.n3272 GND.n3261 585
R18294 GND.t151 GND.n3261 585
R18295 GND.n3636 GND.n3260 585
R18296 GND.n3636 GND.n3635 585
R18297 GND.n3638 GND.n3637 585
R18298 GND.n3637 GND.n3196 585
R18299 GND.n3639 GND.n3194 585
R18300 GND.n3641 GND.n3194 585
R18301 GND.n3258 GND.n3257 585
R18302 GND.n3257 GND.n3190 585
R18303 GND.n3256 GND.n3188 585
R18304 GND.n3647 GND.n3188 585
R18305 GND.n3255 GND.n3254 585
R18306 GND.n3254 GND.n3184 585
R18307 GND.n3253 GND.n3182 585
R18308 GND.n3653 GND.n3182 585
R18309 GND.n3252 GND.n3251 585
R18310 GND.n3251 GND.n3178 585
R18311 GND.n3250 GND.n3176 585
R18312 GND.n3659 GND.n3176 585
R18313 GND.n3249 GND.n3248 585
R18314 GND.n3248 GND.n3172 585
R18315 GND.n3247 GND.n3170 585
R18316 GND.n3665 GND.n3170 585
R18317 GND.n3246 GND.n3245 585
R18318 GND.n3245 GND.n3166 585
R18319 GND.n3244 GND.n3164 585
R18320 GND.n3671 GND.n3164 585
R18321 GND.n3243 GND.n3242 585
R18322 GND.n3242 GND.n3160 585
R18323 GND.n3241 GND.n3158 585
R18324 GND.n3677 GND.n3158 585
R18325 GND.n3240 GND.n3239 585
R18326 GND.n3239 GND.n3154 585
R18327 GND.n3238 GND.n3152 585
R18328 GND.n3683 GND.n3152 585
R18329 GND.n3237 GND.n3236 585
R18330 GND.n3236 GND.n3146 585
R18331 GND.n3235 GND.n3144 585
R18332 GND.n3689 GND.n3144 585
R18333 GND.n3234 GND.n3233 585
R18334 GND.n3233 GND.n3137 585
R18335 GND.n3232 GND.n3135 585
R18336 GND.n3695 GND.n3135 585
R18337 GND.n3231 GND.n3230 585
R18338 GND.n3229 GND.n3228 585
R18339 GND.n3227 GND.n3226 585
R18340 GND.n3225 GND.n3224 585
R18341 GND.n3223 GND.n3222 585
R18342 GND.n3221 GND.n3220 585
R18343 GND.n3219 GND.n3218 585
R18344 GND.n3217 GND.n3216 585
R18345 GND.n3215 GND.n3214 585
R18346 GND.n3213 GND.n3212 585
R18347 GND.n3211 GND.n3210 585
R18348 GND.n3209 GND.n3208 585
R18349 GND.n3207 GND.n3206 585
R18350 GND.n3205 GND.n3204 585
R18351 GND.n3203 GND.n3202 585
R18352 GND.n3201 GND.n3200 585
R18353 GND.n3199 GND.n3198 585
R18354 GND.n3141 GND.n3139 585
R18355 GND.n3694 GND.n3693 585
R18356 GND.n3695 GND.n3694 585
R18357 GND.n3692 GND.n3140 585
R18358 GND.n3140 GND.n3137 585
R18359 GND.n3691 GND.n3690 585
R18360 GND.n3690 GND.n3689 585
R18361 GND.n3143 GND.n3142 585
R18362 GND.n3146 GND.n3143 585
R18363 GND.n3682 GND.n3681 585
R18364 GND.n3683 GND.n3682 585
R18365 GND.n3680 GND.n3155 585
R18366 GND.n3155 GND.n3154 585
R18367 GND.n3679 GND.n3678 585
R18368 GND.n3678 GND.n3677 585
R18369 GND.n3157 GND.n3156 585
R18370 GND.n3160 GND.n3157 585
R18371 GND.n3670 GND.n3669 585
R18372 GND.n3671 GND.n3670 585
R18373 GND.n3668 GND.n3167 585
R18374 GND.n3167 GND.n3166 585
R18375 GND.n3667 GND.n3666 585
R18376 GND.n3666 GND.n3665 585
R18377 GND.n3169 GND.n3168 585
R18378 GND.n3172 GND.n3169 585
R18379 GND.n3658 GND.n3657 585
R18380 GND.n3659 GND.n3658 585
R18381 GND.n3656 GND.n3179 585
R18382 GND.n3179 GND.n3178 585
R18383 GND.n3655 GND.n3654 585
R18384 GND.n3654 GND.n3653 585
R18385 GND.n3181 GND.n3180 585
R18386 GND.n3184 GND.n3181 585
R18387 GND.n3646 GND.n3645 585
R18388 GND.n3647 GND.n3646 585
R18389 GND.n3644 GND.n3191 585
R18390 GND.n3191 GND.n3190 585
R18391 GND.n3643 GND.n3642 585
R18392 GND.n3642 GND.n3641 585
R18393 GND.n3193 GND.n3192 585
R18394 GND.n3196 GND.n3193 585
R18395 GND.n3634 GND.n3633 585
R18396 GND.n3635 GND.n3634 585
R18397 GND.n3632 GND.n3264 585
R18398 GND.n3264 GND.t151 585
R18399 GND.n3631 GND.n3630 585
R18400 GND.n3630 GND.n3629 585
R18401 GND.n3266 GND.n3265 585
R18402 GND.n3269 GND.n3266 585
R18403 GND.n3622 GND.n3621 585
R18404 GND.n3623 GND.n3622 585
R18405 GND.n3620 GND.n3278 585
R18406 GND.n3278 GND.n3276 585
R18407 GND.n3619 GND.n3618 585
R18408 GND.n3618 GND.n3617 585
R18409 GND.n3280 GND.n3279 585
R18410 GND.n3283 GND.n3280 585
R18411 GND.n3610 GND.n3609 585
R18412 GND.n3611 GND.n3610 585
R18413 GND.n3608 GND.n3293 585
R18414 GND.n3293 GND.n3291 585
R18415 GND.n3607 GND.n3606 585
R18416 GND.n3606 GND.n3605 585
R18417 GND.n3295 GND.n3294 585
R18418 GND.n3298 GND.n3295 585
R18419 GND.n3598 GND.n3597 585
R18420 GND.n3599 GND.n3598 585
R18421 GND.n3596 GND.n3308 585
R18422 GND.n3308 GND.n3307 585
R18423 GND.n3595 GND.n3594 585
R18424 GND.n3594 GND.n3593 585
R18425 GND.n3310 GND.n3309 585
R18426 GND.n3313 GND.n3310 585
R18427 GND.n3586 GND.n3585 585
R18428 GND.n3587 GND.n3586 585
R18429 GND.n3584 GND.n3320 585
R18430 GND.n3320 GND.n3319 585
R18431 GND.n3583 GND.n3582 585
R18432 GND.n3582 GND.n3581 585
R18433 GND.n3322 GND.n3321 585
R18434 GND.n3325 GND.n3322 585
R18435 GND.n3574 GND.n3573 585
R18436 GND.n3575 GND.n3574 585
R18437 GND.n3572 GND.n3332 585
R18438 GND.n3332 GND.n3331 585
R18439 GND.n3571 GND.n3570 585
R18440 GND.n3570 GND.n3569 585
R18441 GND.n8731 GND.n8730 585
R18442 GND.n1062 GND.n1061 585
R18443 GND.n8727 GND.n8726 585
R18444 GND.n8728 GND.n8727 585
R18445 GND.n8725 GND.n1723 585
R18446 GND.n8724 GND.n8723 585
R18447 GND.n8722 GND.n8721 585
R18448 GND.n8720 GND.n8719 585
R18449 GND.n8718 GND.n8717 585
R18450 GND.n8716 GND.n8715 585
R18451 GND.n8714 GND.n8713 585
R18452 GND.n8712 GND.n8711 585
R18453 GND.n8710 GND.n8709 585
R18454 GND.n8708 GND.n8707 585
R18455 GND.n8706 GND.n8705 585
R18456 GND.n8704 GND.n8703 585
R18457 GND.n8702 GND.n8701 585
R18458 GND.n8700 GND.n8699 585
R18459 GND.n8698 GND.n1070 585
R18460 GND.n8728 GND.n1070 585
R18461 GND.n8697 GND.n8696 585
R18462 GND.n8696 GND.n1059 585
R18463 GND.n8695 GND.n1057 585
R18464 GND.n8735 GND.n1057 585
R18465 GND.n8694 GND.n8693 585
R18466 GND.n8693 GND.n1053 585
R18467 GND.n8692 GND.n1051 585
R18468 GND.n8741 GND.n1051 585
R18469 GND.n8691 GND.n8690 585
R18470 GND.n8690 GND.n1047 585
R18471 GND.n8689 GND.n1045 585
R18472 GND.n8747 GND.n1045 585
R18473 GND.n8688 GND.n8687 585
R18474 GND.n8687 GND.n1041 585
R18475 GND.n8686 GND.n1039 585
R18476 GND.n8753 GND.n1039 585
R18477 GND.n8685 GND.n8684 585
R18478 GND.n8684 GND.n1035 585
R18479 GND.n8683 GND.n1033 585
R18480 GND.n8759 GND.n1033 585
R18481 GND.n8682 GND.n8681 585
R18482 GND.n8681 GND.n1029 585
R18483 GND.n8680 GND.n1027 585
R18484 GND.n8765 GND.n1027 585
R18485 GND.n8679 GND.n8678 585
R18486 GND.n8678 GND.n1023 585
R18487 GND.n8677 GND.n1021 585
R18488 GND.n8771 GND.n1021 585
R18489 GND.n8676 GND.n8675 585
R18490 GND.n8675 GND.n1015 585
R18491 GND.n8674 GND.n1013 585
R18492 GND.n8777 GND.n1013 585
R18493 GND.n8673 GND.n8672 585
R18494 GND.n8672 GND.n1006 585
R18495 GND.n8670 GND.n1005 585
R18496 GND.n8783 GND.n1005 585
R18497 GND.n8669 GND.n8668 585
R18498 GND.n8668 GND.n1004 585
R18499 GND.n8667 GND.n1724 585
R18500 GND.n8667 GND.n8666 585
R18501 GND.n8658 GND.n1726 585
R18502 GND.n1727 GND.n1726 585
R18503 GND.n8660 GND.n8659 585
R18504 GND.t6 GND.n8660 585
R18505 GND.n8656 GND.n1736 585
R18506 GND.n1736 GND.n1733 585
R18507 GND.n1740 GND.n1737 585
R18508 GND.n8653 GND.n1740 585
R18509 GND.n8644 GND.n8643 585
R18510 GND.n8643 GND.n1739 585
R18511 GND.n8645 GND.n1746 585
R18512 GND.n8647 GND.n1746 585
R18513 GND.n8642 GND.n8641 585
R18514 GND.n8641 GND.n1745 585
R18515 GND.n8640 GND.n1751 585
R18516 GND.n8640 GND.n8639 585
R18517 GND.n8475 GND.n1750 585
R18518 GND.n1752 GND.n1750 585
R18519 GND.n8476 GND.n1759 585
R18520 GND.n8633 GND.n1759 585
R18521 GND.n8478 GND.n8477 585
R18522 GND.n8477 GND.n1758 585
R18523 GND.n8479 GND.n1766 585
R18524 GND.n8625 GND.n1766 585
R18525 GND.n8481 GND.n8480 585
R18526 GND.n8480 GND.n1765 585
R18527 GND.n8482 GND.n1772 585
R18528 GND.n8619 GND.n1772 585
R18529 GND.n8484 GND.n8483 585
R18530 GND.n8483 GND.n1771 585
R18531 GND.n8485 GND.n1778 585
R18532 GND.n8613 GND.n1778 585
R18533 GND.n8487 GND.n8486 585
R18534 GND.n8486 GND.n1777 585
R18535 GND.n8488 GND.n1784 585
R18536 GND.n8607 GND.n1784 585
R18537 GND.n8490 GND.n8489 585
R18538 GND.n8489 GND.n1783 585
R18539 GND.n8491 GND.n1790 585
R18540 GND.n8601 GND.n1790 585
R18541 GND.n8493 GND.n8492 585
R18542 GND.n8492 GND.n1789 585
R18543 GND.n8494 GND.n1796 585
R18544 GND.n8595 GND.n1796 585
R18545 GND.n8495 GND.n8441 585
R18546 GND.n8441 GND.n1795 585
R18547 GND.n8497 GND.n8496 585
R18548 GND.n8474 GND.n8440 585
R18549 GND.n8473 GND.n8472 585
R18550 GND.n8471 GND.n8470 585
R18551 GND.n8469 GND.n8468 585
R18552 GND.n8467 GND.n8466 585
R18553 GND.n8465 GND.n8464 585
R18554 GND.n8463 GND.n8462 585
R18555 GND.n8461 GND.n8460 585
R18556 GND.n8459 GND.n8458 585
R18557 GND.n8457 GND.n8456 585
R18558 GND.n8455 GND.n8454 585
R18559 GND.n8453 GND.n8452 585
R18560 GND.n8451 GND.n8450 585
R18561 GND.n8449 GND.n8448 585
R18562 GND.n8447 GND.n8446 585
R18563 GND.n8445 GND.n8444 585
R18564 GND.n8443 GND.n8442 585
R18565 GND.n1794 GND.n1793 585
R18566 GND.n1795 GND.n1794 585
R18567 GND.n8597 GND.n8596 585
R18568 GND.n8596 GND.n8595 585
R18569 GND.n8598 GND.n1792 585
R18570 GND.n1792 GND.n1789 585
R18571 GND.n8600 GND.n8599 585
R18572 GND.n8601 GND.n8600 585
R18573 GND.n1782 GND.n1781 585
R18574 GND.n1783 GND.n1782 585
R18575 GND.n8609 GND.n8608 585
R18576 GND.n8608 GND.n8607 585
R18577 GND.n8610 GND.n1780 585
R18578 GND.n1780 GND.n1777 585
R18579 GND.n8612 GND.n8611 585
R18580 GND.n8613 GND.n8612 585
R18581 GND.n1770 GND.n1769 585
R18582 GND.n1771 GND.n1770 585
R18583 GND.n8621 GND.n8620 585
R18584 GND.n8620 GND.n8619 585
R18585 GND.n8622 GND.n1768 585
R18586 GND.n1768 GND.n1765 585
R18587 GND.n8624 GND.n8623 585
R18588 GND.n8625 GND.n8624 585
R18589 GND.n1757 GND.n1756 585
R18590 GND.n1758 GND.n1757 585
R18591 GND.n8635 GND.n8634 585
R18592 GND.n8634 GND.n8633 585
R18593 GND.n8636 GND.n1755 585
R18594 GND.n1755 GND.n1752 585
R18595 GND.n8638 GND.n8637 585
R18596 GND.n8639 GND.n8638 585
R18597 GND.n1744 GND.n1743 585
R18598 GND.n1745 GND.n1744 585
R18599 GND.n8649 GND.n8648 585
R18600 GND.n8648 GND.n8647 585
R18601 GND.n8650 GND.n1742 585
R18602 GND.n1742 GND.n1739 585
R18603 GND.n8652 GND.n8651 585
R18604 GND.n8653 GND.n8652 585
R18605 GND.n1732 GND.n1731 585
R18606 GND.n1733 GND.n1732 585
R18607 GND.n8662 GND.n8661 585
R18608 GND.n8661 GND.t6 585
R18609 GND.n8663 GND.n1730 585
R18610 GND.n1730 GND.n1727 585
R18611 GND.n8665 GND.n8664 585
R18612 GND.n8666 GND.n8665 585
R18613 GND.n1010 GND.n1008 585
R18614 GND.n1008 GND.n1004 585
R18615 GND.n8782 GND.n8781 585
R18616 GND.n8783 GND.n8782 585
R18617 GND.n8780 GND.n1009 585
R18618 GND.n1009 GND.n1006 585
R18619 GND.n8779 GND.n8778 585
R18620 GND.n8778 GND.n8777 585
R18621 GND.n1012 GND.n1011 585
R18622 GND.n1015 GND.n1012 585
R18623 GND.n8770 GND.n8769 585
R18624 GND.n8771 GND.n8770 585
R18625 GND.n8768 GND.n1024 585
R18626 GND.n1024 GND.n1023 585
R18627 GND.n8767 GND.n8766 585
R18628 GND.n8766 GND.n8765 585
R18629 GND.n1026 GND.n1025 585
R18630 GND.n1029 GND.n1026 585
R18631 GND.n8758 GND.n8757 585
R18632 GND.n8759 GND.n8758 585
R18633 GND.n8756 GND.n1036 585
R18634 GND.n1036 GND.n1035 585
R18635 GND.n8755 GND.n8754 585
R18636 GND.n8754 GND.n8753 585
R18637 GND.n1038 GND.n1037 585
R18638 GND.n1041 GND.n1038 585
R18639 GND.n8746 GND.n8745 585
R18640 GND.n8747 GND.n8746 585
R18641 GND.n8744 GND.n1048 585
R18642 GND.n1048 GND.n1047 585
R18643 GND.n8743 GND.n8742 585
R18644 GND.n8742 GND.n8741 585
R18645 GND.n1050 GND.n1049 585
R18646 GND.n1053 GND.n1050 585
R18647 GND.n8734 GND.n8733 585
R18648 GND.n8735 GND.n8734 585
R18649 GND.n8732 GND.n1060 585
R18650 GND.n1060 GND.n1059 585
R18651 GND.n1523 GND.n1353 585
R18652 GND.n1522 GND.n1521 585
R18653 GND.n1519 GND.n1354 585
R18654 GND.n1517 GND.n1516 585
R18655 GND.n1515 GND.n1355 585
R18656 GND.n1514 GND.n1513 585
R18657 GND.n1511 GND.n1356 585
R18658 GND.n1509 GND.n1508 585
R18659 GND.n1507 GND.n1357 585
R18660 GND.n1506 GND.n1505 585
R18661 GND.n1503 GND.n1358 585
R18662 GND.n1501 GND.n1500 585
R18663 GND.n1499 GND.n1359 585
R18664 GND.n1498 GND.n1497 585
R18665 GND.n1495 GND.n1360 585
R18666 GND.n1493 GND.n1492 585
R18667 GND.n1491 GND.n1361 585
R18668 GND.n1490 GND.n1489 585
R18669 GND.n1487 GND.n1352 585
R18670 GND.n1526 GND.n1352 585
R18671 GND.n1486 GND.n1485 585
R18672 GND.n1485 GND.n1285 585
R18673 GND.n1484 GND.n1284 585
R18674 GND.n1532 GND.n1284 585
R18675 GND.n1483 GND.n1482 585
R18676 GND.n1482 GND.n1279 585
R18677 GND.n1481 GND.n1278 585
R18678 GND.n1538 GND.n1278 585
R18679 GND.n1480 GND.n1479 585
R18680 GND.n1479 GND.n1273 585
R18681 GND.n1478 GND.n1272 585
R18682 GND.n1544 GND.n1272 585
R18683 GND.n1477 GND.n1476 585
R18684 GND.n1476 GND.n1267 585
R18685 GND.n1475 GND.n1266 585
R18686 GND.n1550 GND.n1266 585
R18687 GND.n1474 GND.n1473 585
R18688 GND.n1473 GND.n1261 585
R18689 GND.n1472 GND.n1260 585
R18690 GND.n1556 GND.n1260 585
R18691 GND.n1471 GND.n1470 585
R18692 GND.n1470 GND.n1252 585
R18693 GND.n1469 GND.n1251 585
R18694 GND.n1562 GND.n1251 585
R18695 GND.n1468 GND.n1467 585
R18696 GND.n1467 GND.n1245 585
R18697 GND.n1466 GND.n1244 585
R18698 GND.n1568 GND.n1244 585
R18699 GND.n1465 GND.n1464 585
R18700 GND.n1464 GND.n1237 585
R18701 GND.n1362 GND.n1236 585
R18702 GND.n1574 GND.n1236 585
R18703 GND.n1442 GND.n1441 585
R18704 GND.n1441 GND.n1230 585
R18705 GND.n1445 GND.n1229 585
R18706 GND.n1580 GND.n1229 585
R18707 GND.n1447 GND.n1446 585
R18708 GND.n1446 GND.n1223 585
R18709 GND.n1448 GND.n1222 585
R18710 GND.n1586 GND.n1222 585
R18711 GND.n1450 GND.n1449 585
R18712 GND.n1449 GND.t310 585
R18713 GND.n1439 GND.n1216 585
R18714 GND.n1592 GND.n1216 585
R18715 GND.n1437 GND.n1436 585
R18716 GND.n1436 GND.n1150 585
R18717 GND.n1433 GND.n1149 585
R18718 GND.n1598 GND.n1149 585
R18719 GND.n1432 GND.n1431 585
R18720 GND.n1431 GND.n1144 585
R18721 GND.n1430 GND.n1143 585
R18722 GND.n1604 GND.n1143 585
R18723 GND.n1429 GND.n1428 585
R18724 GND.n1428 GND.n1138 585
R18725 GND.n1427 GND.n1137 585
R18726 GND.n1610 GND.n1137 585
R18727 GND.n1426 GND.n1425 585
R18728 GND.n1425 GND.n1132 585
R18729 GND.n1424 GND.n1131 585
R18730 GND.n1616 GND.n1131 585
R18731 GND.n1423 GND.n1422 585
R18732 GND.n1422 GND.n1126 585
R18733 GND.n1421 GND.n1125 585
R18734 GND.n1622 GND.n1125 585
R18735 GND.n1420 GND.n1419 585
R18736 GND.n1419 GND.n1120 585
R18737 GND.n1418 GND.n1119 585
R18738 GND.n1628 GND.n1119 585
R18739 GND.n1417 GND.n1416 585
R18740 GND.n1416 GND.n1114 585
R18741 GND.n1415 GND.n1113 585
R18742 GND.n1634 GND.n1113 585
R18743 GND.n1414 GND.n1413 585
R18744 GND.n1413 GND.n1108 585
R18745 GND.n1412 GND.n1107 585
R18746 GND.n1640 GND.n1107 585
R18747 GND.n1411 GND.n1410 585
R18748 GND.n1410 GND.n1100 585
R18749 GND.n1409 GND.n1099 585
R18750 GND.n1646 GND.n1099 585
R18751 GND.n1408 GND.n1407 585
R18752 GND.n1407 GND.n1091 585
R18753 GND.n1406 GND.n1090 585
R18754 GND.n1652 GND.n1090 585
R18755 GND.n1405 GND.n1404 585
R18756 GND.n1403 GND.n1402 585
R18757 GND.n1401 GND.n1400 585
R18758 GND.n1399 GND.n1398 585
R18759 GND.n1397 GND.n1396 585
R18760 GND.n1395 GND.n1394 585
R18761 GND.n1393 GND.n1392 585
R18762 GND.n1391 GND.n1390 585
R18763 GND.n1389 GND.n1388 585
R18764 GND.n1387 GND.n1386 585
R18765 GND.n1385 GND.n1384 585
R18766 GND.n1383 GND.n1382 585
R18767 GND.n1381 GND.n1380 585
R18768 GND.n1379 GND.n1378 585
R18769 GND.n1377 GND.n1376 585
R18770 GND.n1375 GND.n1374 585
R18771 GND.n1373 GND.n1372 585
R18772 GND.n1371 GND.n1370 585
R18773 GND.n1369 GND.n1092 585
R18774 GND.n1652 GND.n1092 585
R18775 GND.n1103 GND.n1101 585
R18776 GND.n1101 GND.n1091 585
R18777 GND.n1645 GND.n1644 585
R18778 GND.n1646 GND.n1645 585
R18779 GND.n1643 GND.n1102 585
R18780 GND.n1102 GND.n1100 585
R18781 GND.n1642 GND.n1641 585
R18782 GND.n1641 GND.n1640 585
R18783 GND.n1105 GND.n1104 585
R18784 GND.n1108 GND.n1105 585
R18785 GND.n1633 GND.n1632 585
R18786 GND.n1634 GND.n1633 585
R18787 GND.n1631 GND.n1115 585
R18788 GND.n1115 GND.n1114 585
R18789 GND.n1630 GND.n1629 585
R18790 GND.n1629 GND.n1628 585
R18791 GND.n1117 GND.n1116 585
R18792 GND.n1120 GND.n1117 585
R18793 GND.n1621 GND.n1620 585
R18794 GND.n1622 GND.n1621 585
R18795 GND.n1619 GND.n1127 585
R18796 GND.n1127 GND.n1126 585
R18797 GND.n1618 GND.n1617 585
R18798 GND.n1617 GND.n1616 585
R18799 GND.n1129 GND.n1128 585
R18800 GND.n1132 GND.n1129 585
R18801 GND.n1609 GND.n1608 585
R18802 GND.n1610 GND.n1609 585
R18803 GND.n1607 GND.n1139 585
R18804 GND.n1139 GND.n1138 585
R18805 GND.n1606 GND.n1605 585
R18806 GND.n1605 GND.n1604 585
R18807 GND.n1141 GND.n1140 585
R18808 GND.n1144 GND.n1141 585
R18809 GND.n1597 GND.n1596 585
R18810 GND.n1598 GND.n1597 585
R18811 GND.n1595 GND.n1151 585
R18812 GND.n1151 GND.n1150 585
R18813 GND.n1217 GND.n1214 585
R18814 GND.n1592 GND.n1217 585
R18815 GND.n1226 GND.n1224 585
R18816 GND.n1224 GND.t310 585
R18817 GND.n1585 GND.n1584 585
R18818 GND.n1586 GND.n1585 585
R18819 GND.n1583 GND.n1225 585
R18820 GND.n1225 GND.n1223 585
R18821 GND.n1231 GND.n1227 585
R18822 GND.n1580 GND.n1231 585
R18823 GND.n1240 GND.n1238 585
R18824 GND.n1238 GND.n1230 585
R18825 GND.n1573 GND.n1572 585
R18826 GND.n1574 GND.n1573 585
R18827 GND.n1571 GND.n1239 585
R18828 GND.n1239 GND.n1237 585
R18829 GND.n1255 GND.n1246 585
R18830 GND.n1568 GND.n1246 585
R18831 GND.n1256 GND.n1253 585
R18832 GND.n1253 GND.n1245 585
R18833 GND.n1561 GND.n1560 585
R18834 GND.n1562 GND.n1561 585
R18835 GND.n1559 GND.n1254 585
R18836 GND.n1254 GND.n1252 585
R18837 GND.n1558 GND.n1557 585
R18838 GND.n1557 GND.n1556 585
R18839 GND.n1258 GND.n1257 585
R18840 GND.n1261 GND.n1258 585
R18841 GND.n1549 GND.n1548 585
R18842 GND.n1550 GND.n1549 585
R18843 GND.n1547 GND.n1268 585
R18844 GND.n1268 GND.n1267 585
R18845 GND.n1546 GND.n1545 585
R18846 GND.n1545 GND.n1544 585
R18847 GND.n1270 GND.n1269 585
R18848 GND.n1273 GND.n1270 585
R18849 GND.n1537 GND.n1536 585
R18850 GND.n1538 GND.n1537 585
R18851 GND.n1535 GND.n1280 585
R18852 GND.n1280 GND.n1279 585
R18853 GND.n1534 GND.n1533 585
R18854 GND.n1533 GND.n1532 585
R18855 GND.n1282 GND.n1281 585
R18856 GND.n1285 GND.n1282 585
R18857 GND.n1525 GND.n1524 585
R18858 GND.n1526 GND.n1525 585
R18859 GND.n1288 GND.n1287 585
R18860 GND.n1319 GND.n1317 585
R18861 GND.n1320 GND.n1316 585
R18862 GND.n1320 GND.n51 585
R18863 GND.n1323 GND.n1322 585
R18864 GND.n1324 GND.n1315 585
R18865 GND.n1326 GND.n1325 585
R18866 GND.n1328 GND.n1314 585
R18867 GND.n1331 GND.n1330 585
R18868 GND.n1332 GND.n1313 585
R18869 GND.n1334 GND.n1333 585
R18870 GND.n1336 GND.n1312 585
R18871 GND.n1339 GND.n1338 585
R18872 GND.n1340 GND.n1311 585
R18873 GND.n1342 GND.n1341 585
R18874 GND.n1344 GND.n1310 585
R18875 GND.n1345 GND.n1309 585
R18876 GND.n1348 GND.n1347 585
R18877 GND.n1349 GND.n1290 585
R18878 GND.n1290 GND.n51 585
R18879 GND.n1351 GND.n1350 585
R18880 GND.n1526 GND.n1351 585
R18881 GND.n1308 GND.n1289 585
R18882 GND.n1289 GND.n1285 585
R18883 GND.n1307 GND.n1283 585
R18884 GND.n1532 GND.n1283 585
R18885 GND.n1306 GND.n1305 585
R18886 GND.n1305 GND.n1279 585
R18887 GND.n1304 GND.n1277 585
R18888 GND.n1538 GND.n1277 585
R18889 GND.n1303 GND.n1302 585
R18890 GND.n1302 GND.n1273 585
R18891 GND.n1301 GND.n1271 585
R18892 GND.n1544 GND.n1271 585
R18893 GND.n1300 GND.n1299 585
R18894 GND.n1299 GND.n1267 585
R18895 GND.n1298 GND.n1265 585
R18896 GND.n1550 GND.n1265 585
R18897 GND.n1297 GND.n1296 585
R18898 GND.n1296 GND.n1261 585
R18899 GND.n1295 GND.n1259 585
R18900 GND.n1556 GND.n1259 585
R18901 GND.n1294 GND.n1293 585
R18902 GND.n1293 GND.n1252 585
R18903 GND.n1292 GND.n1250 585
R18904 GND.n1562 GND.n1250 585
R18905 GND.n1291 GND.n1242 585
R18906 GND.n1245 GND.n1242 585
R18907 GND.n1569 GND.n1243 585
R18908 GND.n1569 GND.n1568 585
R18909 GND.n1571 GND.n1570 585
R18910 GND.n1570 GND.n1237 585
R18911 GND.n1572 GND.n1235 585
R18912 GND.n1574 GND.n1235 585
R18913 GND.n1240 GND.n1228 585
R18914 GND.n1230 GND.n1228 585
R18915 GND.n1581 GND.n1227 585
R18916 GND.n1581 GND.n1580 585
R18917 GND.n1583 GND.n1582 585
R18918 GND.n1582 GND.n1223 585
R18919 GND.n1584 GND.n1221 585
R18920 GND.n1586 GND.n1221 585
R18921 GND.n1226 GND.n1215 585
R18922 GND.t310 GND.n1215 585
R18923 GND.n1593 GND.n1214 585
R18924 GND.n1593 GND.n1592 585
R18925 GND.n1595 GND.n1594 585
R18926 GND.n1594 GND.n1150 585
R18927 GND.n1596 GND.n1148 585
R18928 GND.n1598 GND.n1148 585
R18929 GND.n1212 GND.n1211 585
R18930 GND.n1211 GND.n1144 585
R18931 GND.n1210 GND.n1142 585
R18932 GND.n1604 GND.n1142 585
R18933 GND.n1209 GND.n1208 585
R18934 GND.n1208 GND.n1138 585
R18935 GND.n1207 GND.n1136 585
R18936 GND.n1610 GND.n1136 585
R18937 GND.n1206 GND.n1205 585
R18938 GND.n1205 GND.n1132 585
R18939 GND.n1204 GND.n1130 585
R18940 GND.n1616 GND.n1130 585
R18941 GND.n1203 GND.n1202 585
R18942 GND.n1202 GND.n1126 585
R18943 GND.n1201 GND.n1124 585
R18944 GND.n1622 GND.n1124 585
R18945 GND.n1200 GND.n1199 585
R18946 GND.n1199 GND.n1120 585
R18947 GND.n1198 GND.n1118 585
R18948 GND.n1628 GND.n1118 585
R18949 GND.n1197 GND.n1196 585
R18950 GND.n1196 GND.n1114 585
R18951 GND.n1195 GND.n1112 585
R18952 GND.n1634 GND.n1112 585
R18953 GND.n1194 GND.n1193 585
R18954 GND.n1193 GND.n1108 585
R18955 GND.n1192 GND.n1106 585
R18956 GND.n1640 GND.n1106 585
R18957 GND.n1191 GND.n1190 585
R18958 GND.n1190 GND.n1100 585
R18959 GND.n1189 GND.n1098 585
R18960 GND.n1646 GND.n1098 585
R18961 GND.n1188 GND.n1187 585
R18962 GND.n1187 GND.n1091 585
R18963 GND.n1186 GND.n1089 585
R18964 GND.n1652 GND.n1089 585
R18965 GND.n1185 GND.n1184 585
R18966 GND.n1183 GND.n1182 585
R18967 GND.n1181 GND.n1180 585
R18968 GND.n1179 GND.n1178 585
R18969 GND.n1177 GND.n1176 585
R18970 GND.n1175 GND.n1174 585
R18971 GND.n1173 GND.n1172 585
R18972 GND.n1171 GND.n1170 585
R18973 GND.n1169 GND.n1168 585
R18974 GND.n1167 GND.n1166 585
R18975 GND.n1165 GND.n1164 585
R18976 GND.n1163 GND.n1162 585
R18977 GND.n1161 GND.n1160 585
R18978 GND.n1159 GND.n1158 585
R18979 GND.n1157 GND.n1156 585
R18980 GND.n1155 GND.n1154 585
R18981 GND.n1153 GND.n1152 585
R18982 GND.n1095 GND.n1093 585
R18983 GND.n1651 GND.n1650 585
R18984 GND.n1652 GND.n1651 585
R18985 GND.n1649 GND.n1094 585
R18986 GND.n1094 GND.n1091 585
R18987 GND.n1648 GND.n1647 585
R18988 GND.n1647 GND.n1646 585
R18989 GND.n1097 GND.n1096 585
R18990 GND.n1100 GND.n1097 585
R18991 GND.n1639 GND.n1638 585
R18992 GND.n1640 GND.n1639 585
R18993 GND.n1637 GND.n1109 585
R18994 GND.n1109 GND.n1108 585
R18995 GND.n1636 GND.n1635 585
R18996 GND.n1635 GND.n1634 585
R18997 GND.n1111 GND.n1110 585
R18998 GND.n1114 GND.n1111 585
R18999 GND.n1627 GND.n1626 585
R19000 GND.n1628 GND.n1627 585
R19001 GND.n1625 GND.n1121 585
R19002 GND.n1121 GND.n1120 585
R19003 GND.n1624 GND.n1623 585
R19004 GND.n1623 GND.n1622 585
R19005 GND.n1123 GND.n1122 585
R19006 GND.n1126 GND.n1123 585
R19007 GND.n1615 GND.n1614 585
R19008 GND.n1616 GND.n1615 585
R19009 GND.n1613 GND.n1133 585
R19010 GND.n1133 GND.n1132 585
R19011 GND.n1612 GND.n1611 585
R19012 GND.n1611 GND.n1610 585
R19013 GND.n1135 GND.n1134 585
R19014 GND.n1138 GND.n1135 585
R19015 GND.n1603 GND.n1602 585
R19016 GND.n1604 GND.n1603 585
R19017 GND.n1601 GND.n1145 585
R19018 GND.n1145 GND.n1144 585
R19019 GND.n1600 GND.n1599 585
R19020 GND.n1599 GND.n1598 585
R19021 GND.n1147 GND.n1146 585
R19022 GND.n1150 GND.n1147 585
R19023 GND.n1591 GND.n1590 585
R19024 GND.n1592 GND.n1591 585
R19025 GND.n1589 GND.n1218 585
R19026 GND.n1218 GND.t310 585
R19027 GND.n1588 GND.n1587 585
R19028 GND.n1587 GND.n1586 585
R19029 GND.n1220 GND.n1219 585
R19030 GND.n1223 GND.n1220 585
R19031 GND.n1579 GND.n1578 585
R19032 GND.n1580 GND.n1579 585
R19033 GND.n1577 GND.n1232 585
R19034 GND.n1232 GND.n1230 585
R19035 GND.n1576 GND.n1575 585
R19036 GND.n1575 GND.n1574 585
R19037 GND.n1234 GND.n1233 585
R19038 GND.n1237 GND.n1234 585
R19039 GND.n1567 GND.n1566 585
R19040 GND.n1568 GND.n1567 585
R19041 GND.n1565 GND.n1247 585
R19042 GND.n1247 GND.n1245 585
R19043 GND.n1564 GND.n1563 585
R19044 GND.n1563 GND.n1562 585
R19045 GND.n1249 GND.n1248 585
R19046 GND.n1252 GND.n1249 585
R19047 GND.n1555 GND.n1554 585
R19048 GND.n1556 GND.n1555 585
R19049 GND.n1553 GND.n1262 585
R19050 GND.n1262 GND.n1261 585
R19051 GND.n1552 GND.n1551 585
R19052 GND.n1551 GND.n1550 585
R19053 GND.n1264 GND.n1263 585
R19054 GND.n1267 GND.n1264 585
R19055 GND.n1543 GND.n1542 585
R19056 GND.n1544 GND.n1543 585
R19057 GND.n1541 GND.n1274 585
R19058 GND.n1274 GND.n1273 585
R19059 GND.n1540 GND.n1539 585
R19060 GND.n1539 GND.n1538 585
R19061 GND.n1276 GND.n1275 585
R19062 GND.n1279 GND.n1276 585
R19063 GND.n1531 GND.n1530 585
R19064 GND.n1532 GND.n1531 585
R19065 GND.n1529 GND.n1286 585
R19066 GND.n1286 GND.n1285 585
R19067 GND.n1528 GND.n1527 585
R19068 GND.n1527 GND.n1526 585
R19069 GND.n9202 GND.n9139 585
R19070 GND.n9201 GND.n9200 585
R19071 GND.n9198 GND.n9140 585
R19072 GND.n9198 GND.n50 585
R19073 GND.n9197 GND.n9196 585
R19074 GND.n9195 GND.n9194 585
R19075 GND.n9193 GND.n9142 585
R19076 GND.n9191 GND.n9190 585
R19077 GND.n9189 GND.n9143 585
R19078 GND.n9188 GND.n9187 585
R19079 GND.n9185 GND.n9144 585
R19080 GND.n9183 GND.n9182 585
R19081 GND.n9181 GND.n9145 585
R19082 GND.n9180 GND.n9179 585
R19083 GND.n9177 GND.n9146 585
R19084 GND.n9175 GND.n9174 585
R19085 GND.n9173 GND.n9147 585
R19086 GND.n9172 GND.n9171 585
R19087 GND.n9169 GND.n9138 585
R19088 GND.n9205 GND.n9138 585
R19089 GND.n9168 GND.n9137 585
R19090 GND.n9206 GND.n9137 585
R19091 GND.n9167 GND.n9136 585
R19092 GND.n9207 GND.n9136 585
R19093 GND.n9166 GND.n9165 585
R19094 GND.n9165 GND.n9164 585
R19095 GND.n9163 GND.n411 585
R19096 GND.n9213 GND.n411 585
R19097 GND.n9162 GND.n9161 585
R19098 GND.n9161 GND.n409 585
R19099 GND.n9160 GND.n9159 585
R19100 GND.n9160 GND.n403 585
R19101 GND.n9158 GND.n401 585
R19102 GND.n9221 GND.n401 585
R19103 GND.n9157 GND.n9156 585
R19104 GND.n9156 GND.n9155 585
R19105 GND.n9154 GND.n393 585
R19106 GND.n9227 GND.n393 585
R19107 GND.n9153 GND.n9152 585
R19108 GND.n9152 GND.n391 585
R19109 GND.n9151 GND.n9150 585
R19110 GND.n9151 GND.n383 585
R19111 GND.n9149 GND.n381 585
R19112 GND.n9235 GND.n381 585
R19113 GND.n9237 GND.n9236 585
R19114 GND.n9236 GND.n9235 585
R19115 GND.n377 GND.n376 585
R19116 GND.n383 GND.n377 585
R19117 GND.n397 GND.n395 585
R19118 GND.n395 GND.n391 585
R19119 GND.n9226 GND.n9225 585
R19120 GND.n9227 GND.n9226 585
R19121 GND.n9224 GND.n396 585
R19122 GND.n9155 GND.n396 585
R19123 GND.n9223 GND.n9222 585
R19124 GND.n9222 GND.n9221 585
R19125 GND.n399 GND.n398 585
R19126 GND.n403 GND.n399 585
R19127 GND.n415 GND.n413 585
R19128 GND.n413 GND.n409 585
R19129 GND.n9212 GND.n9211 585
R19130 GND.n9213 GND.n9212 585
R19131 GND.n9210 GND.n414 585
R19132 GND.n9164 GND.n414 585
R19133 GND.n9209 GND.n9208 585
R19134 GND.n9208 GND.n9207 585
R19135 GND.n417 GND.n416 585
R19136 GND.n9206 GND.n417 585
R19137 GND.n9204 GND.n9203 585
R19138 GND.n9205 GND.n9204 585
R19139 GND.n9133 GND.n9132 585
R19140 GND.n9131 GND.n426 585
R19141 GND.n9130 GND.n425 585
R19142 GND.n9135 GND.n425 585
R19143 GND.n9129 GND.n9128 585
R19144 GND.n9127 GND.n9126 585
R19145 GND.n9125 GND.n9124 585
R19146 GND.n9123 GND.n9122 585
R19147 GND.n9121 GND.n9120 585
R19148 GND.n9119 GND.n9118 585
R19149 GND.n9117 GND.n9116 585
R19150 GND.n9115 GND.n9114 585
R19151 GND.n9113 GND.n9112 585
R19152 GND.n9111 GND.n9110 585
R19153 GND.n9109 GND.n9108 585
R19154 GND.n9107 GND.n9106 585
R19155 GND.n9105 GND.n9104 585
R19156 GND.n9103 GND.n9102 585
R19157 GND.n9101 GND.n9100 585
R19158 GND.n9101 GND.n412 585
R19159 GND.n9099 GND.n410 585
R19160 GND.n9214 GND.n410 585
R19161 GND.n9098 GND.n9097 585
R19162 GND.n9097 GND.n9096 585
R19163 GND.n9095 GND.n402 585
R19164 GND.n9220 GND.n402 585
R19165 GND.n9094 GND.n9093 585
R19166 GND.n9093 GND.n400 585
R19167 GND.n9092 GND.n9091 585
R19168 GND.n9092 GND.n394 585
R19169 GND.n9090 GND.n392 585
R19170 GND.n9228 GND.n392 585
R19171 GND.n9089 GND.n9088 585
R19172 GND.n9088 GND.n9087 585
R19173 GND.n9086 GND.n382 585
R19174 GND.n9234 GND.n382 585
R19175 GND.n9085 GND.n9084 585
R19176 GND.n9084 GND.n380 585
R19177 GND.n388 GND.n384 585
R19178 GND.n384 GND.n380 585
R19179 GND.n9233 GND.n9232 585
R19180 GND.n9234 GND.n9233 585
R19181 GND.n9231 GND.n385 585
R19182 GND.n9087 GND.n385 585
R19183 GND.n9230 GND.n9229 585
R19184 GND.n9229 GND.n9228 585
R19185 GND.n390 GND.n389 585
R19186 GND.n394 GND.n390 585
R19187 GND.n406 GND.n404 585
R19188 GND.n404 GND.n400 585
R19189 GND.n9219 GND.n9218 585
R19190 GND.n9220 GND.n9219 585
R19191 GND.n9217 GND.n405 585
R19192 GND.n9096 GND.n405 585
R19193 GND.n9216 GND.n9215 585
R19194 GND.n9215 GND.n9214 585
R19195 GND.n408 GND.n407 585
R19196 GND.n412 GND.n408 585
R19197 GND.n9620 GND.n9619 585
R19198 GND.n9678 GND.n9677 585
R19199 GND.n9676 GND.n9629 585
R19200 GND.n9680 GND.n9629 585
R19201 GND.n9675 GND.n9674 585
R19202 GND.n9673 GND.n9672 585
R19203 GND.n9671 GND.n9670 585
R19204 GND.n9669 GND.n9668 585
R19205 GND.n9667 GND.n9666 585
R19206 GND.n9665 GND.n9664 585
R19207 GND.n9663 GND.n9662 585
R19208 GND.n9661 GND.n9660 585
R19209 GND.n9659 GND.n9658 585
R19210 GND.n9657 GND.n9656 585
R19211 GND.n9655 GND.n9654 585
R19212 GND.n9653 GND.n9652 585
R19213 GND.n9651 GND.n9650 585
R19214 GND.n9649 GND.n9648 585
R19215 GND.n9647 GND.n9621 585
R19216 GND.n9681 GND.n9621 585
R19217 GND.n9646 GND.n9645 585
R19218 GND.n9645 GND.n9617 585
R19219 GND.n9644 GND.n9616 585
R19220 GND.n9687 GND.n9616 585
R19221 GND.n9643 GND.n9642 585
R19222 GND.n9642 GND.n121 585
R19223 GND.n9641 GND.n119 585
R19224 GND.n9696 GND.n119 585
R19225 GND.n9640 GND.n9639 585
R19226 GND.n9639 GND.n9638 585
R19227 GND.n9637 GND.n107 585
R19228 GND.n9702 GND.n107 585
R19229 GND.n9636 GND.n9635 585
R19230 GND.n9635 GND.n96 585
R19231 GND.n9634 GND.n9630 585
R19232 GND.n9634 GND.n90 585
R19233 GND.n9633 GND.n9632 585
R19234 GND.n9633 GND.n103 585
R19235 GND.n9631 GND.n64 585
R19236 GND.n82 GND.n64 585
R19237 GND.n9761 GND.n9760 585
R19238 GND.n9760 GND.n9759 585
R19239 GND.n63 GND.n62 585
R19240 GND.n153 GND.n63 585
R19241 GND.n9519 GND.n74 585
R19242 GND.n9750 GND.n74 585
R19243 GND.n9521 GND.n9520 585
R19244 GND.n9521 GND.n160 585
R19245 GND.n9528 GND.n9527 585
R19246 GND.n9527 GND.n9526 585
R19247 GND.n9529 GND.n183 585
R19248 GND.n183 GND.n166 585
R19249 GND.n9531 GND.n9530 585
R19250 GND.n9533 GND.n9531 585
R19251 GND.n9518 GND.n182 585
R19252 GND.n182 GND.n171 585
R19253 GND.n9517 GND.n9516 585
R19254 GND.n9516 GND.n176 585
R19255 GND.n9515 GND.n174 585
R19256 GND.n9540 GND.n174 585
R19257 GND.n9514 GND.n9513 585
R19258 GND.n9513 GND.n9512 585
R19259 GND.n185 GND.n184 585
R19260 GND.n9511 GND.n185 585
R19261 GND.n9474 GND.n9473 585
R19262 GND.n9474 GND.n9464 585
R19263 GND.n9476 GND.n9475 585
R19264 GND.n9478 GND.n9477 585
R19265 GND.n9480 GND.n9479 585
R19266 GND.n9482 GND.n9481 585
R19267 GND.n9484 GND.n9483 585
R19268 GND.n9486 GND.n9485 585
R19269 GND.n9488 GND.n9487 585
R19270 GND.n9490 GND.n9489 585
R19271 GND.n9492 GND.n9491 585
R19272 GND.n9494 GND.n9493 585
R19273 GND.n9496 GND.n9495 585
R19274 GND.n9498 GND.n9497 585
R19275 GND.n9500 GND.n9499 585
R19276 GND.n9501 GND.n9472 585
R19277 GND.n9503 GND.n9502 585
R19278 GND.n188 GND.n187 585
R19279 GND.n9507 GND.n9506 585
R19280 GND.n9506 GND.n9505 585
R19281 GND.n9508 GND.n186 585
R19282 GND.n9464 GND.n186 585
R19283 GND.n9510 GND.n9509 585
R19284 GND.n9511 GND.n9510 585
R19285 GND.n179 GND.n177 585
R19286 GND.n9512 GND.n177 585
R19287 GND.n9539 GND.n9538 585
R19288 GND.n9540 GND.n9539 585
R19289 GND.n9537 GND.n178 585
R19290 GND.n178 GND.n176 585
R19291 GND.n9536 GND.n9535 585
R19292 GND.n9535 GND.n171 585
R19293 GND.n9534 GND.n180 585
R19294 GND.n9534 GND.n9533 585
R19295 GND.n9523 GND.n181 585
R19296 GND.n181 GND.n166 585
R19297 GND.n9525 GND.n9524 585
R19298 GND.n9526 GND.n9525 585
R19299 GND.n73 GND.n72 585
R19300 GND.n160 GND.n73 585
R19301 GND.n9752 GND.n9751 585
R19302 GND.n9751 GND.n9750 585
R19303 GND.n9753 GND.n67 585
R19304 GND.n153 GND.n67 585
R19305 GND.n9758 GND.n9757 585
R19306 GND.n9759 GND.n9758 585
R19307 GND.n70 GND.n68 585
R19308 GND.n82 GND.n68 585
R19309 GND.n112 GND.n111 585
R19310 GND.n112 GND.n103 585
R19311 GND.n114 GND.n113 585
R19312 GND.n113 GND.n90 585
R19313 GND.n115 GND.n109 585
R19314 GND.n109 GND.n96 585
R19315 GND.n9701 GND.n9700 585
R19316 GND.n9702 GND.n9701 585
R19317 GND.n9699 GND.n110 585
R19318 GND.n9638 GND.n110 585
R19319 GND.n9698 GND.n9697 585
R19320 GND.n9697 GND.n9696 585
R19321 GND.n117 GND.n116 585
R19322 GND.n121 GND.n117 585
R19323 GND.n9686 GND.n9685 585
R19324 GND.n9687 GND.n9686 585
R19325 GND.n9684 GND.n9618 585
R19326 GND.n9618 GND.n9617 585
R19327 GND.n9683 GND.n9682 585
R19328 GND.n9682 GND.n9681 585
R19329 GND.n9692 GND.n123 585
R19330 GND.n9691 GND.n9690 585
R19331 GND.n128 GND.n127 585
R19332 GND.n9688 GND.n128 585
R19333 GND.n9609 GND.n9608 585
R19334 GND.n9610 GND.n130 585
R19335 GND.n9615 GND.n9614 585
R19336 GND.n9688 GND.n9615 585
R19337 GND.n9613 GND.n120 585
R19338 GND.n9695 GND.n120 585
R19339 GND.n9612 GND.n9611 585
R19340 GND.n9611 GND.n118 585
R19341 GND.n106 GND.n105 585
R19342 GND.n108 GND.n106 585
R19343 GND.n9705 GND.n9704 585
R19344 GND.n9704 GND.n9703 585
R19345 GND.n9706 GND.n91 585
R19346 GND.n9735 GND.n91 585
R19347 GND.n9708 GND.n9707 585
R19348 GND.n9709 GND.n9708 585
R19349 GND.n104 GND.n84 585
R19350 GND.n9741 GND.n84 585
R19351 GND.n9567 GND.n9566 585
R19352 GND.n9566 GND.n9565 585
R19353 GND.n9572 GND.n9571 585
R19354 GND.n9572 GND.n65 585
R19355 GND.n9574 GND.n9573 585
R19356 GND.n9573 GND.n76 585
R19357 GND.n9575 GND.n161 585
R19358 GND.n9588 GND.n161 585
R19359 GND.n9576 GND.n168 585
R19360 GND.n9522 GND.n168 585
R19361 GND.n9578 GND.n9577 585
R19362 GND.n9579 GND.n9578 585
R19363 GND.n9563 GND.n167 585
R19364 GND.n9532 GND.n167 585
R19365 GND.n9562 GND.n9561 585
R19366 GND.n9561 GND.n9560 585
R19367 GND.n170 GND.n169 585
R19368 GND.n175 GND.n170 585
R19369 GND.n9547 GND.n9546 585
R19370 GND.n9548 GND.n9543 585
R19371 GND.n9550 GND.n9549 585
R19372 GND.n9552 GND.n9542 585
R19373 GND.n9553 GND.n173 585
R19374 GND.n9556 GND.n9555 585
R19375 GND.n9557 GND.n172 585
R19376 GND.n175 GND.n172 585
R19377 GND.n9559 GND.n9558 585
R19378 GND.n9560 GND.n9559 585
R19379 GND.n165 GND.n164 585
R19380 GND.n9532 GND.n165 585
R19381 GND.n9581 GND.n9580 585
R19382 GND.n9580 GND.n9579 585
R19383 GND.n9582 GND.n162 585
R19384 GND.n9522 GND.n162 585
R19385 GND.n9587 GND.n9586 585
R19386 GND.n9588 GND.n9587 585
R19387 GND.n9585 GND.n163 585
R19388 GND.n163 GND.n76 585
R19389 GND.n9584 GND.n9583 585
R19390 GND.n9583 GND.n65 585
R19391 GND.n87 GND.n85 585
R19392 GND.n9565 GND.n85 585
R19393 GND.n9740 GND.n9739 585
R19394 GND.n9741 GND.n9740 585
R19395 GND.n9738 GND.n86 585
R19396 GND.n9709 GND.n86 585
R19397 GND.n9737 GND.n9736 585
R19398 GND.n9736 GND.n9735 585
R19399 GND.n89 GND.n88 585
R19400 GND.n9703 GND.n89 585
R19401 GND.n125 GND.n124 585
R19402 GND.n124 GND.n108 585
R19403 GND.n126 GND.n122 585
R19404 GND.n122 GND.n118 585
R19405 GND.n9694 GND.n9693 585
R19406 GND.n9695 GND.n9694 585
R19407 GND.n9732 GND.n9731 585
R19408 GND.n9730 GND.n98 585
R19409 GND.n9729 GND.n97 585
R19410 GND.n9734 GND.n97 585
R19411 GND.n9728 GND.n9727 585
R19412 GND.n9721 GND.n100 585
R19413 GND.n9723 GND.n9722 585
R19414 GND.n9719 GND.n9718 585
R19415 GND.n9717 GND.n9716 585
R19416 GND.n9715 GND.n9714 585
R19417 GND.n9713 GND.n95 585
R19418 GND.n9734 GND.n95 585
R19419 GND.n9712 GND.n9711 585
R19420 GND.n9711 GND.n9710 585
R19421 GND.n102 GND.n83 585
R19422 GND.n9742 GND.n83 585
R19423 GND.n152 GND.n151 585
R19424 GND.n152 GND.n66 585
R19425 GND.n156 GND.n155 585
R19426 GND.n155 GND.n154 585
R19427 GND.n157 GND.n75 585
R19428 GND.n9749 GND.n75 585
R19429 GND.n9590 GND.n158 585
R19430 GND.n9590 GND.n9589 585
R19431 GND.n9592 GND.n9591 585
R19432 GND.n9593 GND.n150 585
R19433 GND.n9595 GND.n9594 585
R19434 GND.n9597 GND.n137 585
R19435 GND.n9599 GND.n9598 585
R19436 GND.n140 GND.n135 585
R19437 GND.n147 GND.n146 585
R19438 GND.n145 GND.n139 585
R19439 GND.n144 GND.n143 585
R19440 GND.n142 GND.n141 585
R19441 GND.n79 GND.n77 585
R19442 GND.n9589 GND.n77 585
R19443 GND.n9748 GND.n9747 585
R19444 GND.n9749 GND.n9748 585
R19445 GND.n9746 GND.n78 585
R19446 GND.n154 GND.n78 585
R19447 GND.n9745 GND.n9744 585
R19448 GND.n9744 GND.n66 585
R19449 GND.n9743 GND.n80 585
R19450 GND.n9743 GND.n9742 585
R19451 GND.n99 GND.n81 585
R19452 GND.n9710 GND.n81 585
R19453 GND.n8096 GND.n8033 585
R19454 GND.n8095 GND.n8094 585
R19455 GND.n8092 GND.n8034 585
R19456 GND.n8092 GND.n8032 585
R19457 GND.n8091 GND.n8090 585
R19458 GND.n8089 GND.n8088 585
R19459 GND.n8087 GND.n8036 585
R19460 GND.n8085 GND.n8084 585
R19461 GND.n8083 GND.n8037 585
R19462 GND.n8082 GND.n8081 585
R19463 GND.n8079 GND.n8038 585
R19464 GND.n8077 GND.n8076 585
R19465 GND.n8075 GND.n8039 585
R19466 GND.n8074 GND.n8073 585
R19467 GND.n8071 GND.n8040 585
R19468 GND.n8069 GND.n8068 585
R19469 GND.n8067 GND.n8041 585
R19470 GND.n8066 GND.n8065 585
R19471 GND.n8063 GND.n2111 585
R19472 GND.n8099 GND.n2111 585
R19473 GND.n8062 GND.n2110 585
R19474 GND.n8100 GND.n2110 585
R19475 GND.n8061 GND.n2109 585
R19476 GND.n8101 GND.n2109 585
R19477 GND.n8060 GND.n8059 585
R19478 GND.n8059 GND.n8058 585
R19479 GND.n8057 GND.n2101 585
R19480 GND.n8107 GND.n2101 585
R19481 GND.n8056 GND.n8055 585
R19482 GND.n8055 GND.n2099 585
R19483 GND.n8054 GND.n8053 585
R19484 GND.n8054 GND.n2093 585
R19485 GND.n8052 GND.n2091 585
R19486 GND.n8115 GND.n2091 585
R19487 GND.n8051 GND.n8050 585
R19488 GND.n8050 GND.n8049 585
R19489 GND.n8048 GND.n2083 585
R19490 GND.n8121 GND.n2083 585
R19491 GND.n8047 GND.n8046 585
R19492 GND.n8046 GND.n2081 585
R19493 GND.n8045 GND.n8044 585
R19494 GND.n8045 GND.n2073 585
R19495 GND.n8043 GND.n2071 585
R19496 GND.n8129 GND.n2071 585
R19497 GND.n8131 GND.n8130 585
R19498 GND.n8130 GND.n8129 585
R19499 GND.n2069 GND.n2068 585
R19500 GND.n2073 GND.n2069 585
R19501 GND.n2087 GND.n2085 585
R19502 GND.n2085 GND.n2081 585
R19503 GND.n8120 GND.n8119 585
R19504 GND.n8121 GND.n8120 585
R19505 GND.n8118 GND.n2086 585
R19506 GND.n8049 GND.n2086 585
R19507 GND.n8117 GND.n8116 585
R19508 GND.n8116 GND.n8115 585
R19509 GND.n2089 GND.n2088 585
R19510 GND.n2093 GND.n2089 585
R19511 GND.n2105 GND.n2103 585
R19512 GND.n2103 GND.n2099 585
R19513 GND.n8106 GND.n8105 585
R19514 GND.n8107 GND.n8106 585
R19515 GND.n8104 GND.n2104 585
R19516 GND.n8058 GND.n2104 585
R19517 GND.n8103 GND.n8102 585
R19518 GND.n8102 GND.n8101 585
R19519 GND.n2107 GND.n2106 585
R19520 GND.n8100 GND.n2107 585
R19521 GND.n8098 GND.n8097 585
R19522 GND.n8099 GND.n8098 585
R19523 GND.n4568 GND.n4567 585
R19524 GND.n4571 GND.n4570 585
R19525 GND.n4572 GND.n4566 585
R19526 GND.n4566 GND.n2108 585
R19527 GND.n4574 GND.n4573 585
R19528 GND.n4576 GND.n4565 585
R19529 GND.n4579 GND.n4578 585
R19530 GND.n4580 GND.n4564 585
R19531 GND.n4582 GND.n4581 585
R19532 GND.n4584 GND.n4563 585
R19533 GND.n4587 GND.n4586 585
R19534 GND.n4588 GND.n4562 585
R19535 GND.n4590 GND.n4589 585
R19536 GND.n4592 GND.n4561 585
R19537 GND.n4595 GND.n4594 585
R19538 GND.n4596 GND.n4560 585
R19539 GND.n4598 GND.n4597 585
R19540 GND.n4600 GND.n4559 585
R19541 GND.n4602 GND.n4601 585
R19542 GND.n4601 GND.n2102 585
R19543 GND.n4603 GND.n2100 585
R19544 GND.n8108 GND.n2100 585
R19545 GND.n4606 GND.n4605 585
R19546 GND.n4605 GND.n4604 585
R19547 GND.n4607 GND.n2092 585
R19548 GND.n8114 GND.n2092 585
R19549 GND.n4609 GND.n4608 585
R19550 GND.n4609 GND.n2090 585
R19551 GND.n4611 GND.n4610 585
R19552 GND.n4610 GND.n2084 585
R19553 GND.n4612 GND.n2082 585
R19554 GND.n8122 GND.n2082 585
R19555 GND.n4615 GND.n4614 585
R19556 GND.n4614 GND.n4613 585
R19557 GND.n4616 GND.n2072 585
R19558 GND.n8128 GND.n2072 585
R19559 GND.n4618 GND.n4617 585
R19560 GND.n4618 GND.n2070 585
R19561 GND.n2078 GND.n2074 585
R19562 GND.n2074 GND.n2070 585
R19563 GND.n8127 GND.n8126 585
R19564 GND.n8128 GND.n8127 585
R19565 GND.n8125 GND.n2075 585
R19566 GND.n4613 GND.n2075 585
R19567 GND.n8124 GND.n8123 585
R19568 GND.n8123 GND.n8122 585
R19569 GND.n2080 GND.n2079 585
R19570 GND.n2084 GND.n2080 585
R19571 GND.n2096 GND.n2094 585
R19572 GND.n2094 GND.n2090 585
R19573 GND.n8113 GND.n8112 585
R19574 GND.n8114 GND.n8113 585
R19575 GND.n8111 GND.n2095 585
R19576 GND.n4604 GND.n2095 585
R19577 GND.n8110 GND.n8109 585
R19578 GND.n8109 GND.n8108 585
R19579 GND.n2098 GND.n2097 585
R19580 GND.n2102 GND.n2098 585
R19581 GND.n716 GND.n537 585
R19582 GND.n537 GND.n190 585
R19583 GND.n715 GND.n531 585
R19584 GND.n730 GND.n531 585
R19585 GND.n714 GND.n713 585
R19586 GND.n713 GND.n712 585
R19587 GND.n540 GND.n539 585
R19588 GND.n551 GND.n540 585
R19589 GND.n620 GND.n548 585
R19590 GND.n703 GND.n548 585
R19591 GND.n622 GND.n621 585
R19592 GND.n621 GND.n546 585
R19593 GND.n623 GND.n555 585
R19594 GND.n696 GND.n555 585
R19595 GND.n625 GND.n624 585
R19596 GND.n625 GND.n560 585
R19597 GND.n627 GND.n626 585
R19598 GND.n626 GND.n559 585
R19599 GND.n628 GND.n567 585
R19600 GND.n639 GND.n567 585
R19601 GND.n629 GND.n575 585
R19602 GND.n575 GND.n566 585
R19603 GND.n631 GND.n630 585
R19604 GND.n632 GND.n631 585
R19605 GND.n619 GND.n574 585
R19606 GND.n574 GND.n573 585
R19607 GND.n618 GND.n617 585
R19608 GND.n577 GND.n576 585
R19609 GND.n587 GND.n586 585
R19610 GND.n589 GND.n588 585
R19611 GND.n591 GND.n590 585
R19612 GND.n593 GND.n592 585
R19613 GND.n595 GND.n594 585
R19614 GND.n597 GND.n596 585
R19615 GND.n599 GND.n598 585
R19616 GND.n601 GND.n600 585
R19617 GND.n603 GND.n602 585
R19618 GND.n605 GND.n604 585
R19619 GND.n607 GND.n606 585
R19620 GND.n609 GND.n608 585
R19621 GND.n611 GND.n610 585
R19622 GND.n612 GND.n585 585
R19623 GND.n614 GND.n613 585
R19624 GND.n615 GND.n614 585
R19625 GND.n572 GND.n571 585
R19626 GND.n573 GND.n572 585
R19627 GND.n634 GND.n633 585
R19628 GND.n633 GND.n632 585
R19629 GND.n635 GND.n569 585
R19630 GND.n569 GND.n566 585
R19631 GND.n638 GND.n637 585
R19632 GND.n639 GND.n638 585
R19633 GND.n636 GND.n570 585
R19634 GND.n570 GND.n559 585
R19635 GND.n554 GND.n553 585
R19636 GND.n560 GND.n554 585
R19637 GND.n698 GND.n697 585
R19638 GND.n697 GND.n696 585
R19639 GND.n699 GND.n550 585
R19640 GND.n550 GND.n546 585
R19641 GND.n702 GND.n701 585
R19642 GND.n703 GND.n702 585
R19643 GND.n700 GND.n552 585
R19644 GND.n552 GND.n551 585
R19645 GND.n534 GND.n532 585
R19646 GND.n712 GND.n532 585
R19647 GND.n729 GND.n728 585
R19648 GND.n730 GND.n729 585
R19649 GND.n727 GND.n533 585
R19650 GND.n533 GND.n190 585
R19651 GND.n734 GND.n191 585
R19652 GND.n9431 GND.n191 585
R19653 GND.n733 GND.n732 585
R19654 GND.n732 GND.n731 585
R19655 GND.n529 GND.n528 585
R19656 GND.n530 GND.n529 585
R19657 GND.n689 GND.n541 585
R19658 GND.n711 GND.n541 585
R19659 GND.n691 GND.n690 585
R19660 GND.n690 GND.n549 585
R19661 GND.n692 GND.n547 585
R19662 GND.n704 GND.n547 585
R19663 GND.n694 GND.n693 585
R19664 GND.n695 GND.n694 585
R19665 GND.n688 GND.n556 585
R19666 GND.n562 GND.n556 585
R19667 GND.n687 GND.n686 585
R19668 GND.n686 GND.n685 585
R19669 GND.n558 GND.n557 585
R19670 GND.n568 GND.n558 585
R19671 GND.n649 GND.n648 585
R19672 GND.n651 GND.n650 585
R19673 GND.n653 GND.n652 585
R19674 GND.n655 GND.n654 585
R19675 GND.n657 GND.n656 585
R19676 GND.n659 GND.n658 585
R19677 GND.n661 GND.n660 585
R19678 GND.n663 GND.n662 585
R19679 GND.n665 GND.n664 585
R19680 GND.n667 GND.n666 585
R19681 GND.n669 GND.n668 585
R19682 GND.n671 GND.n670 585
R19683 GND.n673 GND.n672 585
R19684 GND.n674 GND.n647 585
R19685 GND.n676 GND.n675 585
R19686 GND.n565 GND.n564 585
R19687 GND.n680 GND.n679 585
R19688 GND.n679 GND.n678 585
R19689 GND.n681 GND.n561 585
R19690 GND.n568 GND.n561 585
R19691 GND.n684 GND.n683 585
R19692 GND.n685 GND.n684 585
R19693 GND.n682 GND.n563 585
R19694 GND.n563 GND.n562 585
R19695 GND.n545 GND.n544 585
R19696 GND.n695 GND.n545 585
R19697 GND.n706 GND.n705 585
R19698 GND.n705 GND.n704 585
R19699 GND.n707 GND.n542 585
R19700 GND.n549 GND.n542 585
R19701 GND.n710 GND.n709 585
R19702 GND.n711 GND.n710 585
R19703 GND.n708 GND.n543 585
R19704 GND.n543 GND.n530 585
R19705 GND.n194 GND.n192 585
R19706 GND.n731 GND.n192 585
R19707 GND.n9430 GND.n9429 585
R19708 GND.n9431 GND.n9430 585
R19709 GND.n8027 GND.n8026 585
R19710 GND.n8025 GND.n2128 585
R19711 GND.n8024 GND.n2127 585
R19712 GND.n8029 GND.n2127 585
R19713 GND.n8023 GND.n8022 585
R19714 GND.n8021 GND.n8020 585
R19715 GND.n8019 GND.n8018 585
R19716 GND.n8017 GND.n8016 585
R19717 GND.n8015 GND.n8014 585
R19718 GND.n8013 GND.n8012 585
R19719 GND.n8011 GND.n8010 585
R19720 GND.n8009 GND.n8008 585
R19721 GND.n8007 GND.n8006 585
R19722 GND.n8005 GND.n8004 585
R19723 GND.n8003 GND.n8002 585
R19724 GND.n8001 GND.n8000 585
R19725 GND.n7999 GND.n7998 585
R19726 GND.n7997 GND.n7996 585
R19727 GND.n7995 GND.n2131 585
R19728 GND.n7995 GND.n7994 585
R19729 GND.n7899 GND.n2132 585
R19730 GND.n7993 GND.n2132 585
R19731 GND.n7901 GND.n7900 585
R19732 GND.n7900 GND.n2133 585
R19733 GND.n7902 GND.n2138 585
R19734 GND.n7987 GND.n2138 585
R19735 GND.n7904 GND.n7903 585
R19736 GND.n7905 GND.n7904 585
R19737 GND.n7898 GND.n2193 585
R19738 GND.n7911 GND.n2193 585
R19739 GND.n7897 GND.n2190 585
R19740 GND.n7923 GND.n2190 585
R19741 GND.n7896 GND.n7895 585
R19742 GND.n7895 GND.n2180 585
R19743 GND.n7894 GND.n2201 585
R19744 GND.n7894 GND.n2174 585
R19745 GND.n7893 GND.n7892 585
R19746 GND.n7893 GND.n2186 585
R19747 GND.n7891 GND.n2202 585
R19748 GND.n2202 GND.n2166 585
R19749 GND.n2252 GND.n2203 585
R19750 GND.n2253 GND.n2252 585
R19751 GND.n7887 GND.n2158 585
R19752 GND.n7970 GND.n2158 585
R19753 GND.n7885 GND.n7884 585
R19754 GND.n7884 GND.n7883 585
R19755 GND.n2206 GND.n2205 585
R19756 GND.n7873 GND.n2206 585
R19757 GND.n7796 GND.n7795 585
R19758 GND.n7795 GND.n2213 585
R19759 GND.n7797 GND.n2220 585
R19760 GND.n7867 GND.n2220 585
R19761 GND.n7800 GND.n7798 585
R19762 GND.n7800 GND.n7799 585
R19763 GND.n7801 GND.n7794 585
R19764 GND.n7801 GND.n2257 585
R19765 GND.n7803 GND.n7802 585
R19766 GND.n7802 GND.n2263 585
R19767 GND.n7804 GND.n2261 585
R19768 GND.n7817 GND.n2261 585
R19769 GND.n7806 GND.n7805 585
R19770 GND.n7807 GND.n7806 585
R19771 GND.n7793 GND.n2268 585
R19772 GND.n7808 GND.n2268 585
R19773 GND.n7792 GND.n7791 585
R19774 GND.n7791 GND.n7790 585
R19775 GND.n2270 GND.n2269 585
R19776 GND.n7759 GND.n7758 585
R19777 GND.n7761 GND.n7760 585
R19778 GND.n7763 GND.n7762 585
R19779 GND.n7765 GND.n7764 585
R19780 GND.n7767 GND.n7766 585
R19781 GND.n7769 GND.n7768 585
R19782 GND.n7771 GND.n7770 585
R19783 GND.n7773 GND.n7772 585
R19784 GND.n7775 GND.n7774 585
R19785 GND.n7777 GND.n7776 585
R19786 GND.n7779 GND.n7778 585
R19787 GND.n7781 GND.n7780 585
R19788 GND.n7783 GND.n7782 585
R19789 GND.n7785 GND.n7784 585
R19790 GND.n7786 GND.n7757 585
R19791 GND.n7788 GND.n7787 585
R19792 GND.n7789 GND.n7788 585
R19793 GND.n2267 GND.n2266 585
R19794 GND.n7790 GND.n2267 585
R19795 GND.n7810 GND.n7809 585
R19796 GND.n7809 GND.n7808 585
R19797 GND.n7811 GND.n2264 585
R19798 GND.n7807 GND.n2264 585
R19799 GND.n7816 GND.n7815 585
R19800 GND.n7817 GND.n7816 585
R19801 GND.n7814 GND.n2265 585
R19802 GND.n2265 GND.n2263 585
R19803 GND.n7813 GND.n7812 585
R19804 GND.n7812 GND.n2257 585
R19805 GND.n2218 GND.n2217 585
R19806 GND.n7799 GND.n2218 585
R19807 GND.n7869 GND.n7868 585
R19808 GND.n7868 GND.n7867 585
R19809 GND.n7870 GND.n2216 585
R19810 GND.n2216 GND.n2213 585
R19811 GND.n7872 GND.n7871 585
R19812 GND.n7873 GND.n7872 585
R19813 GND.n2155 GND.n2154 585
R19814 GND.n7883 GND.n2155 585
R19815 GND.n7972 GND.n7971 585
R19816 GND.n7971 GND.n7970 585
R19817 GND.n2157 GND.n2156 585
R19818 GND.n2253 GND.n2157 585
R19819 GND.n7915 GND.n7914 585
R19820 GND.n7915 GND.n2166 585
R19821 GND.n7916 GND.n7913 585
R19822 GND.n7916 GND.n2186 585
R19823 GND.n7918 GND.n7917 585
R19824 GND.n7917 GND.n2174 585
R19825 GND.n7919 GND.n2192 585
R19826 GND.n2192 GND.n2180 585
R19827 GND.n7922 GND.n7921 585
R19828 GND.n7923 GND.n7922 585
R19829 GND.n7920 GND.n7912 585
R19830 GND.n7912 GND.n7911 585
R19831 GND.n2136 GND.n2135 585
R19832 GND.n7905 GND.n2136 585
R19833 GND.n7989 GND.n7988 585
R19834 GND.n7988 GND.n7987 585
R19835 GND.n7990 GND.n2134 585
R19836 GND.n2134 GND.n2133 585
R19837 GND.n7992 GND.n7991 585
R19838 GND.n7993 GND.n7992 585
R19839 GND.n2130 GND.n2129 585
R19840 GND.n7994 GND.n2129 585
R19841 GND.n7984 GND.n7983 585
R19842 GND.n7982 GND.n2142 585
R19843 GND.n7981 GND.n2141 585
R19844 GND.n7986 GND.n2141 585
R19845 GND.n2146 GND.n2145 585
R19846 GND.n2196 GND.n2195 585
R19847 GND.n2197 GND.n2140 585
R19848 GND.n7986 GND.n2140 585
R19849 GND.n2198 GND.n2194 585
R19850 GND.n2194 GND.n2137 585
R19851 GND.n2200 GND.n2199 585
R19852 GND.n7910 GND.n2200 585
R19853 GND.n2189 GND.n2188 585
R19854 GND.n2191 GND.n2189 585
R19855 GND.n7926 GND.n7925 585
R19856 GND.n7925 GND.n7924 585
R19857 GND.n7927 GND.n2175 585
R19858 GND.n7956 GND.n2175 585
R19859 GND.n7929 GND.n7928 585
R19860 GND.n7930 GND.n7929 585
R19861 GND.n2187 GND.n2168 585
R19862 GND.n7962 GND.n2168 585
R19863 GND.n7854 GND.n7853 585
R19864 GND.n7855 GND.n7854 585
R19865 GND.n7850 GND.n2254 585
R19866 GND.n2254 GND.n2160 585
R19867 GND.n7848 GND.n2208 585
R19868 GND.n7881 GND.n2208 585
R19869 GND.n7847 GND.n7846 585
R19870 GND.n7846 GND.n7845 585
R19871 GND.n7844 GND.n2214 585
R19872 GND.n7874 GND.n2214 585
R19873 GND.n7843 GND.n2221 585
R19874 GND.n7866 GND.n2221 585
R19875 GND.n7842 GND.n7841 585
R19876 GND.n7841 GND.n2219 585
R19877 GND.n7840 GND.n2255 585
R19878 GND.n7840 GND.n7839 585
R19879 GND.n7822 GND.n2256 585
R19880 GND.n2262 GND.n2256 585
R19881 GND.n7825 GND.n7824 585
R19882 GND.n7826 GND.n7820 585
R19883 GND.n7828 GND.n7827 585
R19884 GND.n7830 GND.n7819 585
R19885 GND.n7831 GND.n2260 585
R19886 GND.n7834 GND.n7833 585
R19887 GND.n7835 GND.n2258 585
R19888 GND.n2262 GND.n2258 585
R19889 GND.n7838 GND.n7837 585
R19890 GND.n7839 GND.n7838 585
R19891 GND.n7836 GND.n2259 585
R19892 GND.n2259 GND.n2219 585
R19893 GND.n2212 GND.n2211 585
R19894 GND.n7866 GND.n2212 585
R19895 GND.n7876 GND.n7875 585
R19896 GND.n7875 GND.n7874 585
R19897 GND.n7877 GND.n2209 585
R19898 GND.n7845 GND.n2209 585
R19899 GND.n7880 GND.n7879 585
R19900 GND.n7881 GND.n7880 585
R19901 GND.n7878 GND.n2210 585
R19902 GND.n2210 GND.n2160 585
R19903 GND.n2171 GND.n2169 585
R19904 GND.n7855 GND.n2169 585
R19905 GND.n7961 GND.n7960 585
R19906 GND.n7962 GND.n7961 585
R19907 GND.n7959 GND.n2170 585
R19908 GND.n7930 GND.n2170 585
R19909 GND.n7958 GND.n7957 585
R19910 GND.n7957 GND.n7956 585
R19911 GND.n2173 GND.n2172 585
R19912 GND.n7924 GND.n2173 585
R19913 GND.n7907 GND.n7906 585
R19914 GND.n7906 GND.n2191 585
R19915 GND.n7909 GND.n7908 585
R19916 GND.n7910 GND.n7909 585
R19917 GND.n2144 GND.n2143 585
R19918 GND.n2143 GND.n2137 585
R19919 GND.n7953 GND.n7952 585
R19920 GND.n7951 GND.n2182 585
R19921 GND.n7950 GND.n2181 585
R19922 GND.n7955 GND.n2181 585
R19923 GND.n7949 GND.n7948 585
R19924 GND.n7942 GND.n2183 585
R19925 GND.n7944 GND.n7943 585
R19926 GND.n7940 GND.n7939 585
R19927 GND.n7938 GND.n7937 585
R19928 GND.n7936 GND.n7935 585
R19929 GND.n7934 GND.n2179 585
R19930 GND.n7955 GND.n2179 585
R19931 GND.n7933 GND.n7932 585
R19932 GND.n7932 GND.n7931 585
R19933 GND.n2185 GND.n2167 585
R19934 GND.n7963 GND.n2167 585
R19935 GND.n7858 GND.n7857 585
R19936 GND.n7857 GND.n7856 585
R19937 GND.n7859 GND.n2159 585
R19938 GND.n7969 GND.n2159 585
R19939 GND.n7860 GND.n2207 585
R19940 GND.n7882 GND.n2207 585
R19941 GND.n7861 GND.n2227 585
R19942 GND.n2227 GND.n2215 585
R19943 GND.n7863 GND.n7862 585
R19944 GND.n2251 GND.n2226 585
R19945 GND.n2250 GND.n2249 585
R19946 GND.n2248 GND.n2247 585
R19947 GND.n2246 GND.n2245 585
R19948 GND.n2238 GND.n2229 585
R19949 GND.n2240 GND.n2239 585
R19950 GND.n2237 GND.n2236 585
R19951 GND.n2235 GND.n2234 585
R19952 GND.n2233 GND.n2232 585
R19953 GND.n2231 GND.n2230 585
R19954 GND.n2231 GND.n2215 585
R19955 GND.n2163 GND.n2161 585
R19956 GND.n7882 GND.n2161 585
R19957 GND.n7968 GND.n7967 585
R19958 GND.n7969 GND.n7968 585
R19959 GND.n7966 GND.n2162 585
R19960 GND.n7856 GND.n2162 585
R19961 GND.n7965 GND.n7964 585
R19962 GND.n7964 GND.n7963 585
R19963 GND.n2165 GND.n2164 585
R19964 GND.n7931 GND.n2165 585
R19965 GND.n2659 GND.n2658 585
R19966 GND.n2658 GND.n2657 585
R19967 GND.n2660 GND.n2480 585
R19968 GND.n7428 GND.n2480 585
R19969 GND.n2663 GND.n2662 585
R19970 GND.n2662 GND.n2478 585
R19971 GND.n2647 GND.n2488 585
R19972 GND.n7420 GND.n2488 585
R19973 GND.n2669 GND.n2668 585
R19974 GND.n2669 GND.n2496 585
R19975 GND.n2672 GND.n2671 585
R19976 GND.n2671 GND.n2670 585
R19977 GND.n2644 GND.n2507 585
R19978 GND.n7389 GND.n2507 585
R19979 GND.n2679 GND.n2678 585
R19980 GND.n2678 GND.n2677 585
R19981 GND.n2681 GND.n2515 585
R19982 GND.n7375 GND.n2515 585
R19983 GND.n2641 GND.n2640 585
R19984 GND.n2640 GND.n2617 585
R19985 GND.n2687 GND.n2686 585
R19986 GND.n2687 GND.n2545 585
R19987 GND.n7246 GND.n7245 585
R19988 GND.n7245 GND.n7244 585
R19989 GND.n2639 GND.n2637 585
R19990 GND.n2639 GND.n2555 585
R19991 GND.n7192 GND.n6635 585
R19992 GND.n7192 GND.n7191 585
R19993 GND.n7194 GND.n7193 585
R19994 GND.n7193 GND.n6609 585
R19995 GND.n6636 GND.n6634 585
R19996 GND.n6636 GND.n6629 585
R19997 GND.n7164 GND.n7163 585
R19998 GND.n7163 GND.n6618 585
R19999 GND.n7161 GND.n6649 585
R20000 GND.n7174 GND.n6649 585
R20001 GND.n6662 GND.n6658 585
R20002 GND.n6683 GND.n6662 585
R20003 GND.n7156 GND.n7155 585
R20004 GND.n7155 GND.n7154 585
R20005 GND.n6928 GND.n6661 585
R20006 GND.n6688 GND.n6661 585
R20007 GND.n6927 GND.n6672 585
R20008 GND.n7141 GND.n6672 585
R20009 GND.n6935 GND.n6933 585
R20010 GND.n6935 GND.n6934 585
R20011 GND.n6937 GND.n6936 585
R20012 GND.n6936 GND.n6693 585
R20013 GND.n6924 GND.n6750 585
R20014 GND.n7012 GND.n6750 585
R20015 GND.n6942 GND.n6941 585
R20016 GND.n6941 GND.n6757 585
R20017 GND.n6943 GND.n6755 585
R20018 GND.n6999 GND.n6755 585
R20019 GND.n7001 GND.n7000 585
R20020 GND.n7000 GND.n6999 585
R20021 GND.n7002 GND.n6751 585
R20022 GND.n6757 GND.n6751 585
R20023 GND.n7011 GND.n7010 585
R20024 GND.n7012 GND.n7011 585
R20025 GND.n7004 GND.n6752 585
R20026 GND.n6752 GND.n6693 585
R20027 GND.n7005 GND.n6670 585
R20028 GND.n6934 GND.n6670 585
R20029 GND.n7143 GND.n7142 585
R20030 GND.n7142 GND.n7141 585
R20031 GND.n7144 GND.n6665 585
R20032 GND.n6688 GND.n6665 585
R20033 GND.n7153 GND.n7152 585
R20034 GND.n7154 GND.n7153 585
R20035 GND.n6667 GND.n6645 585
R20036 GND.n6683 GND.n6645 585
R20037 GND.n7175 GND.n6647 585
R20038 GND.n7175 GND.n7174 585
R20039 GND.n7176 GND.n6643 585
R20040 GND.n7176 GND.n6618 585
R20041 GND.n7178 GND.n7177 585
R20042 GND.n7177 GND.n6629 585
R20043 GND.n6638 GND.n6637 585
R20044 GND.n6637 GND.n6609 585
R20045 GND.n7190 GND.n7189 585
R20046 GND.n7191 GND.n7190 585
R20047 GND.n7188 GND.n2690 585
R20048 GND.n2690 GND.n2555 585
R20049 GND.n7243 GND.n7242 585
R20050 GND.n7244 GND.n7243 585
R20051 GND.n2693 GND.n2691 585
R20052 GND.n2691 GND.n2545 585
R20053 GND.n7236 GND.n2514 585
R20054 GND.n2617 GND.n2514 585
R20055 GND.n7377 GND.n7376 585
R20056 GND.n7376 GND.n7375 585
R20057 GND.n7378 GND.n2508 585
R20058 GND.n2677 GND.n2508 585
R20059 GND.n7388 GND.n7387 585
R20060 GND.n7389 GND.n7388 585
R20061 GND.n2511 GND.n2509 585
R20062 GND.n2670 GND.n2509 585
R20063 GND.n7382 GND.n2486 585
R20064 GND.n2496 GND.n2486 585
R20065 GND.n7422 GND.n7421 585
R20066 GND.n7421 GND.n7420 585
R20067 GND.n2483 GND.n2482 585
R20068 GND.n2482 GND.n2478 585
R20069 GND.n7427 GND.n7426 585
R20070 GND.n7428 GND.n7427 585
R20071 GND.n2423 GND.n2421 585
R20072 GND.n2657 GND.n2421 585
R20073 GND.n7364 GND.n7363 585
R20074 GND.n7361 GND.n2531 585
R20075 GND.n7360 GND.n7359 585
R20076 GND.n7358 GND.n7357 585
R20077 GND.n7356 GND.n2533 585
R20078 GND.n7354 GND.n7353 585
R20079 GND.n7352 GND.n2534 585
R20080 GND.n7351 GND.n7350 585
R20081 GND.n7348 GND.n2535 585
R20082 GND.n7346 GND.n7345 585
R20083 GND.n7344 GND.n2536 585
R20084 GND.n7343 GND.n7342 585
R20085 GND.n7340 GND.n2537 585
R20086 GND.n7338 GND.n7337 585
R20087 GND.n7336 GND.n2538 585
R20088 GND.n7335 GND.n7334 585
R20089 GND.n7332 GND.n2539 585
R20090 GND.n7332 GND.n2487 585
R20091 GND.n7331 GND.n7330 585
R20092 GND.n7331 GND.n2495 585
R20093 GND.n7329 GND.n2526 585
R20094 GND.n7368 GND.n2526 585
R20095 GND.n7328 GND.n7327 585
R20096 GND.n7327 GND.n2505 585
R20097 GND.n7326 GND.n2517 585
R20098 GND.n7374 GND.n2517 585
R20099 GND.n2544 GND.n2540 585
R20100 GND.n7297 GND.n2544 585
R20101 GND.n7322 GND.n7321 585
R20102 GND.n7321 GND.n7320 585
R20103 GND.n7233 GND.n2543 585
R20104 GND.n2689 GND.n2543 585
R20105 GND.n7232 GND.n2557 585
R20106 GND.n7309 GND.n2557 585
R20107 GND.n7231 GND.n7230 585
R20108 GND.n7230 GND.t238 585
R20109 GND.n7229 GND.n2695 585
R20110 GND.n7229 GND.n7228 585
R20111 GND.n7184 GND.n6608 585
R20112 GND.n7202 GND.n6608 585
R20113 GND.n6640 GND.n6620 585
R20114 GND.n7219 GND.n6620 585
R20115 GND.n7119 GND.n6651 585
R20116 GND.n7173 GND.n6651 585
R20117 GND.n7121 GND.n6685 585
R20118 GND.n7133 GND.n6685 585
R20119 GND.n7122 GND.n6690 585
R20120 GND.n6690 GND.n6664 585
R20121 GND.n7124 GND.n7123 585
R20122 GND.n7125 GND.n7124 585
R20123 GND.n7117 GND.n6674 585
R20124 GND.n7140 GND.n6674 585
R20125 GND.n7116 GND.n7115 585
R20126 GND.n6692 GND.n6691 585
R20127 GND.n6729 GND.n6728 585
R20128 GND.n6727 GND.n6701 585
R20129 GND.n6726 GND.n6725 585
R20130 GND.n6724 GND.n6723 585
R20131 GND.n6722 GND.n6721 585
R20132 GND.n6720 GND.n6719 585
R20133 GND.n6718 GND.n6717 585
R20134 GND.n6716 GND.n6715 585
R20135 GND.n6714 GND.n6713 585
R20136 GND.n6712 GND.n6711 585
R20137 GND.n6710 GND.n6709 585
R20138 GND.n6708 GND.n6707 585
R20139 GND.n6706 GND.n6705 585
R20140 GND.n6704 GND.n6703 585
R20141 GND.n6702 GND.n6694 585
R20142 GND.n7113 GND.n6694 585
R20143 GND.n6687 GND.n6676 585
R20144 GND.n7140 GND.n6676 585
R20145 GND.n7127 GND.n7126 585
R20146 GND.n7126 GND.n7125 585
R20147 GND.n7128 GND.n6686 585
R20148 GND.n6686 GND.n6664 585
R20149 GND.n7132 GND.n7131 585
R20150 GND.n7133 GND.n7132 585
R20151 GND.n7129 GND.n6622 585
R20152 GND.n7173 GND.n6622 585
R20153 GND.n7218 GND.n7217 585
R20154 GND.n7219 GND.n7218 585
R20155 GND.n6625 GND.n6623 585
R20156 GND.n7202 GND.n6623 585
R20157 GND.n7211 GND.n6612 585
R20158 GND.n7228 GND.n6612 585
R20159 GND.n2561 GND.n2559 585
R20160 GND.t238 GND.n2559 585
R20161 GND.n7308 GND.n7307 585
R20162 GND.n7309 GND.n7308 585
R20163 GND.n2562 GND.n2560 585
R20164 GND.n2689 GND.n2560 585
R20165 GND.n7290 GND.n2548 585
R20166 GND.n7320 GND.n2548 585
R20167 GND.n7296 GND.n7295 585
R20168 GND.n7297 GND.n7296 585
R20169 GND.n7292 GND.n2519 585
R20170 GND.n7374 GND.n2519 585
R20171 GND.n2530 GND.n2528 585
R20172 GND.n2528 GND.n2505 585
R20173 GND.n7367 GND.n7366 585
R20174 GND.n7368 GND.n7367 585
R20175 GND.n7365 GND.n2529 585
R20176 GND.n2529 GND.n2495 585
R20177 GND.n2577 GND.n2576 585
R20178 GND.n2580 GND.n2579 585
R20179 GND.n2581 GND.n2575 585
R20180 GND.n2575 GND.n2487 585
R20181 GND.n2583 GND.n2582 585
R20182 GND.n2585 GND.n2574 585
R20183 GND.n2588 GND.n2587 585
R20184 GND.n2589 GND.n2573 585
R20185 GND.n2591 GND.n2590 585
R20186 GND.n2593 GND.n2572 585
R20187 GND.n2596 GND.n2595 585
R20188 GND.n2597 GND.n2571 585
R20189 GND.n2599 GND.n2598 585
R20190 GND.n2601 GND.n2570 585
R20191 GND.n2604 GND.n2603 585
R20192 GND.n2605 GND.n2569 585
R20193 GND.n2607 GND.n2606 585
R20194 GND.n2609 GND.n2568 585
R20195 GND.n2611 GND.n2610 585
R20196 GND.n2610 GND.n2495 585
R20197 GND.n2612 GND.n2525 585
R20198 GND.n7368 GND.n2525 585
R20199 GND.n2614 GND.n2613 585
R20200 GND.n2613 GND.n2505 585
R20201 GND.n2615 GND.n2516 585
R20202 GND.n7374 GND.n2516 585
R20203 GND.n7299 GND.n7298 585
R20204 GND.n7298 GND.n7297 585
R20205 GND.n7301 GND.n2546 585
R20206 GND.n7320 GND.n2546 585
R20207 GND.n2688 GND.n2567 585
R20208 GND.n2689 GND.n2688 585
R20209 GND.n7207 GND.n2556 585
R20210 GND.n7309 GND.n2556 585
R20211 GND.n7209 GND.n7208 585
R20212 GND.n7208 GND.t238 585
R20213 GND.n7206 GND.n6610 585
R20214 GND.n7228 GND.n6610 585
R20215 GND.n7204 GND.n7203 585
R20216 GND.n7203 GND.n7202 585
R20217 GND.n7074 GND.n6619 585
R20218 GND.n7219 GND.n6619 585
R20219 GND.n7073 GND.n6650 585
R20220 GND.n7173 GND.n6650 585
R20221 GND.n7078 GND.n6684 585
R20222 GND.n7133 GND.n6684 585
R20223 GND.n7080 GND.n7079 585
R20224 GND.n7079 GND.n6664 585
R20225 GND.n7081 GND.n6689 585
R20226 GND.n7125 GND.n6689 585
R20227 GND.n7082 GND.n6673 585
R20228 GND.n7140 GND.n6673 585
R20229 GND.n7084 GND.n7083 585
R20230 GND.n7086 GND.n7085 585
R20231 GND.n7088 GND.n7087 585
R20232 GND.n7090 GND.n7089 585
R20233 GND.n7092 GND.n7091 585
R20234 GND.n7094 GND.n7093 585
R20235 GND.n7096 GND.n7095 585
R20236 GND.n7098 GND.n7097 585
R20237 GND.n7100 GND.n7099 585
R20238 GND.n7102 GND.n7101 585
R20239 GND.n7104 GND.n7103 585
R20240 GND.n7106 GND.n7105 585
R20241 GND.n7108 GND.n7107 585
R20242 GND.n7109 GND.n7071 585
R20243 GND.n7111 GND.n7110 585
R20244 GND.n7072 GND.n7070 585
R20245 GND.n6679 GND.n6677 585
R20246 GND.n7113 GND.n6677 585
R20247 GND.n7139 GND.n7138 585
R20248 GND.n7140 GND.n7139 585
R20249 GND.n7137 GND.n6678 585
R20250 GND.n7125 GND.n6678 585
R20251 GND.n7136 GND.n7135 585
R20252 GND.n7135 GND.n6664 585
R20253 GND.n7134 GND.n6682 585
R20254 GND.n7134 GND.n7133 585
R20255 GND.n6680 GND.n6617 585
R20256 GND.n7173 GND.n6617 585
R20257 GND.n7221 GND.n7220 585
R20258 GND.n7220 GND.n7219 585
R20259 GND.n6614 GND.n6613 585
R20260 GND.n7202 GND.n6613 585
R20261 GND.n7227 GND.n7226 585
R20262 GND.n7228 GND.n7227 585
R20263 GND.n2554 GND.n2553 585
R20264 GND.t238 GND.n2554 585
R20265 GND.n7311 GND.n7310 585
R20266 GND.n7310 GND.n7309 585
R20267 GND.n7312 GND.n2549 585
R20268 GND.n2689 GND.n2549 585
R20269 GND.n7319 GND.n7318 585
R20270 GND.n7320 GND.n7319 585
R20271 GND.n2551 GND.n2520 585
R20272 GND.n7297 GND.n2520 585
R20273 GND.n7373 GND.n7372 585
R20274 GND.n7374 GND.n7373 585
R20275 GND.n7371 GND.n2521 585
R20276 GND.n2521 GND.n2505 585
R20277 GND.n7370 GND.n7369 585
R20278 GND.n7369 GND.n7368 585
R20279 GND.n2524 GND.n2523 585
R20280 GND.n2524 GND.n2495 585
R20281 GND.n7550 GND.n7549 585
R20282 GND.n7548 GND.n2463 585
R20283 GND.n7547 GND.n2462 585
R20284 GND.n7552 GND.n2462 585
R20285 GND.n7546 GND.n7545 585
R20286 GND.n7544 GND.n7543 585
R20287 GND.n7542 GND.n7541 585
R20288 GND.n7540 GND.n7539 585
R20289 GND.n7538 GND.n7537 585
R20290 GND.n7536 GND.n7535 585
R20291 GND.n7534 GND.n7533 585
R20292 GND.n7532 GND.n7531 585
R20293 GND.n7530 GND.n7529 585
R20294 GND.n7528 GND.n7527 585
R20295 GND.n7526 GND.n7525 585
R20296 GND.n7524 GND.n7523 585
R20297 GND.n7522 GND.n7521 585
R20298 GND.n7520 GND.n7519 585
R20299 GND.n7518 GND.n2466 585
R20300 GND.n7518 GND.n2452 585
R20301 GND.n7517 GND.n7516 585
R20302 GND.n7517 GND.n2446 585
R20303 GND.n7515 GND.n2444 585
R20304 GND.n7560 GND.n2444 585
R20305 GND.n7514 GND.n7513 585
R20306 GND.n7513 GND.n7512 585
R20307 GND.n2467 GND.n2437 585
R20308 GND.n7566 GND.n2437 585
R20309 GND.n2649 GND.n2648 585
R20310 GND.n2649 GND.n2435 585
R20311 GND.n2651 GND.n2650 585
R20312 GND.n2650 GND.n2429 585
R20313 GND.n2652 GND.n2427 585
R20314 GND.n7574 GND.n2427 585
R20315 GND.n2655 GND.n2654 585
R20316 GND.n2654 GND.n2653 585
R20317 GND.n2656 GND.n2419 585
R20318 GND.n7580 GND.n2419 585
R20319 GND.n7579 GND.n7578 585
R20320 GND.n7580 GND.n7579 585
R20321 GND.n7577 GND.n2422 585
R20322 GND.n2653 GND.n2422 585
R20323 GND.n7576 GND.n7575 585
R20324 GND.n7575 GND.n7574 585
R20325 GND.n2425 GND.n2424 585
R20326 GND.n2429 GND.n2425 585
R20327 GND.n2441 GND.n2439 585
R20328 GND.n2439 GND.n2435 585
R20329 GND.n7565 GND.n7564 585
R20330 GND.n7566 GND.n7565 585
R20331 GND.n7563 GND.n2440 585
R20332 GND.n7512 GND.n2440 585
R20333 GND.n7562 GND.n7561 585
R20334 GND.n7561 GND.n7560 585
R20335 GND.n2443 GND.n2442 585
R20336 GND.n2446 GND.n2443 585
R20337 GND.n2465 GND.n2464 585
R20338 GND.n2464 GND.n2452 585
R20339 GND.n1890 GND.n1872 585
R20340 GND.n2271 GND.n1872 585
R20341 GND.n1889 GND.n1864 585
R20342 GND.n8332 GND.n1864 585
R20343 GND.n1888 GND.n1887 585
R20344 GND.n1887 GND.n1862 585
R20345 GND.n1886 GND.n1885 585
R20346 GND.n1886 GND.n1856 585
R20347 GND.n1884 GND.n1854 585
R20348 GND.n8340 GND.n1854 585
R20349 GND.n1883 GND.n1882 585
R20350 GND.n1882 GND.n1881 585
R20351 GND.n1880 GND.n1846 585
R20352 GND.n8346 GND.n1846 585
R20353 GND.n1879 GND.n1878 585
R20354 GND.n1878 GND.n1844 585
R20355 GND.n1877 GND.n1876 585
R20356 GND.n1877 GND.n1838 585
R20357 GND.n1875 GND.n1836 585
R20358 GND.n8354 GND.n1836 585
R20359 GND.n1874 GND.n1829 585
R20360 GND.n1834 GND.n1829 585
R20361 GND.n8361 GND.n1830 585
R20362 GND.n8361 GND.n8360 585
R20363 GND.n8362 GND.n1828 585
R20364 GND.n8362 GND.n1816 585
R20365 GND.n8364 GND.n8363 585
R20366 GND.n8366 GND.n8365 585
R20367 GND.n8368 GND.n8367 585
R20368 GND.n8370 GND.n8369 585
R20369 GND.n8372 GND.n8371 585
R20370 GND.n8374 GND.n8373 585
R20371 GND.n8376 GND.n8375 585
R20372 GND.n8378 GND.n8377 585
R20373 GND.n8380 GND.n8379 585
R20374 GND.n8382 GND.n8381 585
R20375 GND.n8384 GND.n8383 585
R20376 GND.n8386 GND.n8385 585
R20377 GND.n8388 GND.n8387 585
R20378 GND.n8390 GND.n8389 585
R20379 GND.n8392 GND.n8391 585
R20380 GND.n8393 GND.n1826 585
R20381 GND.n8395 GND.n8394 585
R20382 GND.n8396 GND.n8395 585
R20383 GND.n1827 GND.n1825 585
R20384 GND.n1825 GND.n1816 585
R20385 GND.n8359 GND.n8358 585
R20386 GND.n8360 GND.n8359 585
R20387 GND.n8357 GND.n1831 585
R20388 GND.n1834 GND.n1831 585
R20389 GND.n8356 GND.n8355 585
R20390 GND.n8355 GND.n8354 585
R20391 GND.n1833 GND.n1832 585
R20392 GND.n1838 GND.n1833 585
R20393 GND.n1850 GND.n1848 585
R20394 GND.n1848 GND.n1844 585
R20395 GND.n8345 GND.n8344 585
R20396 GND.n8346 GND.n8345 585
R20397 GND.n8343 GND.n1849 585
R20398 GND.n1881 GND.n1849 585
R20399 GND.n8342 GND.n8341 585
R20400 GND.n8341 GND.n8340 585
R20401 GND.n1852 GND.n1851 585
R20402 GND.n1856 GND.n1852 585
R20403 GND.n1868 GND.n1866 585
R20404 GND.n1866 GND.n1862 585
R20405 GND.n8331 GND.n8330 585
R20406 GND.n8332 GND.n8331 585
R20407 GND.n8329 GND.n1867 585
R20408 GND.n2271 GND.n1867 585
R20409 GND.n4332 GND.n4331 585
R20410 GND.n4332 GND.n2272 585
R20411 GND.n4330 GND.n4275 585
R20412 GND.n4275 GND.n1865 585
R20413 GND.n4329 GND.n1863 585
R20414 GND.n8333 GND.n1863 585
R20415 GND.n4328 GND.n4327 585
R20416 GND.n4327 GND.n4326 585
R20417 GND.n4325 GND.n1855 585
R20418 GND.n8339 GND.n1855 585
R20419 GND.n4324 GND.n4323 585
R20420 GND.n4323 GND.n1853 585
R20421 GND.n4322 GND.n4321 585
R20422 GND.n4322 GND.n1847 585
R20423 GND.n4320 GND.n1845 585
R20424 GND.n8347 GND.n1845 585
R20425 GND.n4319 GND.n4318 585
R20426 GND.n4318 GND.n4317 585
R20427 GND.n4316 GND.n1837 585
R20428 GND.n8353 GND.n1837 585
R20429 GND.n4315 GND.n4314 585
R20430 GND.n4312 GND.n4276 585
R20431 GND.n4311 GND.n4310 585
R20432 GND.n4309 GND.n4308 585
R20433 GND.n4307 GND.n4278 585
R20434 GND.n4305 GND.n4304 585
R20435 GND.n4303 GND.n4279 585
R20436 GND.n4302 GND.n4301 585
R20437 GND.n4299 GND.n4280 585
R20438 GND.n4297 GND.n4296 585
R20439 GND.n4295 GND.n4281 585
R20440 GND.n4294 GND.n4293 585
R20441 GND.n4291 GND.n4282 585
R20442 GND.n4289 GND.n4288 585
R20443 GND.n4287 GND.n4283 585
R20444 GND.n4286 GND.n4285 585
R20445 GND.n1841 GND.n1839 585
R20446 GND.n1839 GND.n1835 585
R20447 GND.n8352 GND.n8351 585
R20448 GND.n8353 GND.n8352 585
R20449 GND.n8350 GND.n1840 585
R20450 GND.n4317 GND.n1840 585
R20451 GND.n8349 GND.n8348 585
R20452 GND.n8348 GND.n8347 585
R20453 GND.n1843 GND.n1842 585
R20454 GND.n1847 GND.n1843 585
R20455 GND.n1859 GND.n1857 585
R20456 GND.n1857 GND.n1853 585
R20457 GND.n8338 GND.n8337 585
R20458 GND.n8339 GND.n8338 585
R20459 GND.n8336 GND.n1858 585
R20460 GND.n4326 GND.n1858 585
R20461 GND.n8335 GND.n8334 585
R20462 GND.n8334 GND.n8333 585
R20463 GND.n1861 GND.n1860 585
R20464 GND.n1865 GND.n1861 585
R20465 GND.n4336 GND.n4334 585
R20466 GND.n4334 GND.n2272 585
R20467 GND.n5370 GND.n5369 585
R20468 GND.n5369 GND.n3843 585
R20469 GND.n5371 GND.n3845 585
R20470 GND.n5777 GND.n3845 585
R20471 GND.n5374 GND.n5373 585
R20472 GND.n5373 GND.n5372 585
R20473 GND.n5375 GND.n3853 585
R20474 GND.n5771 GND.n3853 585
R20475 GND.n5377 GND.n5376 585
R20476 GND.n5377 GND.n3855 585
R20477 GND.n5379 GND.n5378 585
R20478 GND.n5378 GND.n3861 585
R20479 GND.n5380 GND.n3863 585
R20480 GND.n5763 GND.n3863 585
R20481 GND.n5383 GND.n5382 585
R20482 GND.n5382 GND.n5381 585
R20483 GND.n5384 GND.n3871 585
R20484 GND.n5757 GND.n3871 585
R20485 GND.n5386 GND.n5385 585
R20486 GND.n5386 GND.n3873 585
R20487 GND.n5388 GND.n5387 585
R20488 GND.n5387 GND.n3879 585
R20489 GND.n5389 GND.n3881 585
R20490 GND.n5749 GND.n3881 585
R20491 GND.n5392 GND.n5391 585
R20492 GND.n5391 GND.n5390 585
R20493 GND.n5393 GND.n3889 585
R20494 GND.n5743 GND.n3889 585
R20495 GND.n5395 GND.n5394 585
R20496 GND.n5395 GND.n3891 585
R20497 GND.n5397 GND.n5396 585
R20498 GND.n5396 GND.n3897 585
R20499 GND.n5398 GND.n3899 585
R20500 GND.n5735 GND.n3899 585
R20501 GND.n5401 GND.n5399 585
R20502 GND.n5401 GND.n5400 585
R20503 GND.n5403 GND.n5402 585
R20504 GND.n5405 GND.n5404 585
R20505 GND.n5407 GND.n5406 585
R20506 GND.n5409 GND.n5408 585
R20507 GND.n5411 GND.n5410 585
R20508 GND.n5413 GND.n5412 585
R20509 GND.n5415 GND.n5414 585
R20510 GND.n5417 GND.n5416 585
R20511 GND.n5419 GND.n5418 585
R20512 GND.n5421 GND.n5420 585
R20513 GND.n5423 GND.n5422 585
R20514 GND.n5425 GND.n5424 585
R20515 GND.n5427 GND.n5426 585
R20516 GND.n5429 GND.n5428 585
R20517 GND.n5431 GND.n5430 585
R20518 GND.n5434 GND.n5433 585
R20519 GND.n5432 GND.n5027 585
R20520 GND.n5025 GND.n5024 585
R20521 GND.n5023 GND.n5022 585
R20522 GND.n5021 GND.n5020 585
R20523 GND.n5019 GND.n5018 585
R20524 GND.n5017 GND.n5016 585
R20525 GND.n5015 GND.n5005 585
R20526 GND.n5694 GND.n5693 585
R20527 GND.n5696 GND.n5695 585
R20528 GND.n5698 GND.n5697 585
R20529 GND.n5700 GND.n5699 585
R20530 GND.n5702 GND.n5701 585
R20531 GND.n5704 GND.n5703 585
R20532 GND.n5706 GND.n5705 585
R20533 GND.n5708 GND.n5707 585
R20534 GND.n5710 GND.n5709 585
R20535 GND.n5712 GND.n5711 585
R20536 GND.n5714 GND.n5713 585
R20537 GND.n5716 GND.n5715 585
R20538 GND.n5718 GND.n5717 585
R20539 GND.n5720 GND.n5719 585
R20540 GND.n5722 GND.n5721 585
R20541 GND.n5724 GND.n5723 585
R20542 GND.n5725 GND.n5003 585
R20543 GND.n5727 GND.n5726 585
R20544 GND.n3905 GND.n3904 585
R20545 GND.n5731 GND.n5730 585
R20546 GND.n5730 GND.n5729 585
R20547 GND.n5732 GND.n3902 585
R20548 GND.n5400 GND.n3902 585
R20549 GND.n5734 GND.n5733 585
R20550 GND.n5735 GND.n5734 585
R20551 GND.n3903 GND.n3901 585
R20552 GND.n3901 GND.n3897 585
R20553 GND.n3887 GND.n3886 585
R20554 GND.n3891 GND.n3887 585
R20555 GND.n5745 GND.n5744 585
R20556 GND.n5744 GND.n5743 585
R20557 GND.n5746 GND.n3884 585
R20558 GND.n5390 GND.n3884 585
R20559 GND.n5748 GND.n5747 585
R20560 GND.n5749 GND.n5748 585
R20561 GND.n3885 GND.n3883 585
R20562 GND.n3883 GND.n3879 585
R20563 GND.n3869 GND.n3868 585
R20564 GND.n3873 GND.n3869 585
R20565 GND.n5759 GND.n5758 585
R20566 GND.n5758 GND.n5757 585
R20567 GND.n5760 GND.n3866 585
R20568 GND.n5381 GND.n3866 585
R20569 GND.n5762 GND.n5761 585
R20570 GND.n5763 GND.n5762 585
R20571 GND.n3867 GND.n3865 585
R20572 GND.n3865 GND.n3861 585
R20573 GND.n3851 GND.n3850 585
R20574 GND.n3855 GND.n3851 585
R20575 GND.n5773 GND.n5772 585
R20576 GND.n5772 GND.n5771 585
R20577 GND.n5774 GND.n3848 585
R20578 GND.n5372 GND.n3848 585
R20579 GND.n5776 GND.n5775 585
R20580 GND.n5777 GND.n5776 585
R20581 GND.n3849 GND.n3847 585
R20582 GND.n3847 GND.n3843 585
R20583 GND.n5097 GND.n5096 585
R20584 GND.n5100 GND.n5099 585
R20585 GND.n5101 GND.n5095 585
R20586 GND.n5095 GND.n3837 585
R20587 GND.n5103 GND.n5102 585
R20588 GND.n5105 GND.n5094 585
R20589 GND.n5108 GND.n5107 585
R20590 GND.n5109 GND.n5093 585
R20591 GND.n5111 GND.n5110 585
R20592 GND.n5113 GND.n5092 585
R20593 GND.n5116 GND.n5115 585
R20594 GND.n5117 GND.n5091 585
R20595 GND.n5119 GND.n5118 585
R20596 GND.n5121 GND.n5090 585
R20597 GND.n5124 GND.n5123 585
R20598 GND.n5125 GND.n5089 585
R20599 GND.n5127 GND.n5126 585
R20600 GND.n5129 GND.n5088 585
R20601 GND.n5132 GND.n5131 585
R20602 GND.n5047 GND.n5046 585
R20603 GND.n5141 GND.n5140 585
R20604 GND.n5143 GND.n5045 585
R20605 GND.n5146 GND.n5145 585
R20606 GND.n5043 GND.n5042 585
R20607 GND.n5153 GND.n5152 585
R20608 GND.n5155 GND.n5041 585
R20609 GND.n5159 GND.n5158 585
R20610 GND.n5156 GND.n5037 585
R20611 GND.n5338 GND.n5039 585
R20612 GND.n5340 GND.n5035 585
R20613 GND.n5342 GND.n5341 585
R20614 GND.n5344 GND.n5034 585
R20615 GND.n5347 GND.n5346 585
R20616 GND.n5348 GND.n5033 585
R20617 GND.n5350 GND.n5349 585
R20618 GND.n5352 GND.n5032 585
R20619 GND.n5355 GND.n5354 585
R20620 GND.n5356 GND.n5031 585
R20621 GND.n5358 GND.n5357 585
R20622 GND.n5360 GND.n5030 585
R20623 GND.n5363 GND.n5362 585
R20624 GND.n5364 GND.n5029 585
R20625 GND.n5366 GND.n5365 585
R20626 GND.n5368 GND.n5028 585
R20627 GND.n4081 GND.n4080 585
R20628 GND.n4080 GND.n4079 585
R20629 GND.n4082 GND.n3844 585
R20630 GND.n5778 GND.n3844 585
R20631 GND.n4084 GND.n4083 585
R20632 GND.n4084 GND.n3846 585
R20633 GND.n4086 GND.n4085 585
R20634 GND.n4085 GND.n3852 585
R20635 GND.n4087 GND.n3854 585
R20636 GND.n5770 GND.n3854 585
R20637 GND.n4090 GND.n4089 585
R20638 GND.n4089 GND.n4088 585
R20639 GND.n4091 GND.n3862 585
R20640 GND.n5764 GND.n3862 585
R20641 GND.n4093 GND.n4092 585
R20642 GND.n4093 GND.n3864 585
R20643 GND.n4095 GND.n4094 585
R20644 GND.n4094 GND.n3870 585
R20645 GND.n4096 GND.n3872 585
R20646 GND.n5756 GND.n3872 585
R20647 GND.n4099 GND.n4098 585
R20648 GND.n4098 GND.n4097 585
R20649 GND.n4100 GND.n3880 585
R20650 GND.n5750 GND.n3880 585
R20651 GND.n4102 GND.n4101 585
R20652 GND.n4102 GND.n3882 585
R20653 GND.n4104 GND.n4103 585
R20654 GND.n4103 GND.n3888 585
R20655 GND.n4105 GND.n3890 585
R20656 GND.n5742 GND.n3890 585
R20657 GND.n4108 GND.n4107 585
R20658 GND.n4107 GND.n4106 585
R20659 GND.n4109 GND.n3898 585
R20660 GND.n5736 GND.n3898 585
R20661 GND.n4111 GND.n4110 585
R20662 GND.n4111 GND.n3900 585
R20663 GND.n4113 GND.n4112 585
R20664 GND.n4115 GND.n4114 585
R20665 GND.n4117 GND.n4116 585
R20666 GND.n4119 GND.n4118 585
R20667 GND.n4121 GND.n4120 585
R20668 GND.n4123 GND.n4122 585
R20669 GND.n4125 GND.n4124 585
R20670 GND.n4127 GND.n4126 585
R20671 GND.n4129 GND.n4128 585
R20672 GND.n4131 GND.n4130 585
R20673 GND.n4133 GND.n4132 585
R20674 GND.n4135 GND.n4134 585
R20675 GND.n4137 GND.n4136 585
R20676 GND.n4139 GND.n4138 585
R20677 GND.n4141 GND.n4140 585
R20678 GND.n4143 GND.n4142 585
R20679 GND.n4145 GND.n4144 585
R20680 GND.n4148 GND.n4147 585
R20681 GND.n4146 GND.n3951 585
R20682 GND.n3949 GND.n3948 585
R20683 GND.n3947 GND.n3946 585
R20684 GND.n3945 GND.n3944 585
R20685 GND.n3943 GND.n3942 585
R20686 GND.n3941 GND.n3940 585
R20687 GND.n3939 GND.n3929 585
R20688 GND.n4948 GND.n4947 585
R20689 GND.n4950 GND.n4949 585
R20690 GND.n4952 GND.n4951 585
R20691 GND.n4954 GND.n4953 585
R20692 GND.n4956 GND.n4955 585
R20693 GND.n4958 GND.n4957 585
R20694 GND.n4960 GND.n4959 585
R20695 GND.n4962 GND.n4961 585
R20696 GND.n4964 GND.n4963 585
R20697 GND.n4966 GND.n4965 585
R20698 GND.n4968 GND.n4967 585
R20699 GND.n4970 GND.n4969 585
R20700 GND.n4972 GND.n4971 585
R20701 GND.n4974 GND.n4973 585
R20702 GND.n4976 GND.n4975 585
R20703 GND.n4978 GND.n4977 585
R20704 GND.n4979 GND.n3927 585
R20705 GND.n4981 GND.n4980 585
R20706 GND.n4982 GND.n4981 585
R20707 GND.n3896 GND.n3895 585
R20708 GND.n3900 GND.n3896 585
R20709 GND.n5738 GND.n5737 585
R20710 GND.n5737 GND.n5736 585
R20711 GND.n5739 GND.n3893 585
R20712 GND.n4106 GND.n3893 585
R20713 GND.n5741 GND.n5740 585
R20714 GND.n5742 GND.n5741 585
R20715 GND.n3894 GND.n3892 585
R20716 GND.n3892 GND.n3888 585
R20717 GND.n3878 GND.n3877 585
R20718 GND.n3882 GND.n3878 585
R20719 GND.n5752 GND.n5751 585
R20720 GND.n5751 GND.n5750 585
R20721 GND.n5753 GND.n3875 585
R20722 GND.n4097 GND.n3875 585
R20723 GND.n5755 GND.n5754 585
R20724 GND.n5756 GND.n5755 585
R20725 GND.n3876 GND.n3874 585
R20726 GND.n3874 GND.n3870 585
R20727 GND.n3860 GND.n3859 585
R20728 GND.n3864 GND.n3860 585
R20729 GND.n5766 GND.n5765 585
R20730 GND.n5765 GND.n5764 585
R20731 GND.n5767 GND.n3857 585
R20732 GND.n4088 GND.n3857 585
R20733 GND.n5769 GND.n5768 585
R20734 GND.n5770 GND.n5769 585
R20735 GND.n3858 GND.n3856 585
R20736 GND.n3856 GND.n3852 585
R20737 GND.n3842 GND.n3841 585
R20738 GND.n3846 GND.n3842 585
R20739 GND.n5780 GND.n5779 585
R20740 GND.n5779 GND.n5778 585
R20741 GND.n5781 GND.n3840 585
R20742 GND.n4079 GND.n3840 585
R20743 GND.n5807 GND.n5806 585
R20744 GND.n5805 GND.n3839 585
R20745 GND.n5804 GND.n3838 585
R20746 GND.n5809 GND.n3838 585
R20747 GND.n5803 GND.n5802 585
R20748 GND.n5801 GND.n5800 585
R20749 GND.n5799 GND.n5798 585
R20750 GND.n5797 GND.n5796 585
R20751 GND.n5795 GND.n5794 585
R20752 GND.n5793 GND.n5792 585
R20753 GND.n5791 GND.n5790 585
R20754 GND.n5789 GND.n5788 585
R20755 GND.n5787 GND.n5786 585
R20756 GND.n5785 GND.n5784 585
R20757 GND.n5783 GND.n5782 585
R20758 GND.n3816 GND.n3815 585
R20759 GND.n5812 GND.n5811 585
R20760 GND.n3817 GND.n3814 585
R20761 GND.n4019 GND.n4016 585
R20762 GND.n4021 GND.n4020 585
R20763 GND.n4025 GND.n4022 585
R20764 GND.n4027 GND.n4026 585
R20765 GND.n4031 GND.n4028 585
R20766 GND.n4033 GND.n4032 585
R20767 GND.n4037 GND.n4034 585
R20768 GND.n4039 GND.n4038 585
R20769 GND.n4043 GND.n4040 585
R20770 GND.n4046 GND.n4045 585
R20771 GND.n4048 GND.n4047 585
R20772 GND.n4050 GND.n4049 585
R20773 GND.n4052 GND.n4051 585
R20774 GND.n4054 GND.n4053 585
R20775 GND.n4056 GND.n4055 585
R20776 GND.n4058 GND.n4057 585
R20777 GND.n4060 GND.n4059 585
R20778 GND.n4062 GND.n4061 585
R20779 GND.n4064 GND.n4063 585
R20780 GND.n4066 GND.n4065 585
R20781 GND.n4068 GND.n4067 585
R20782 GND.n4070 GND.n4069 585
R20783 GND.n4072 GND.n4071 585
R20784 GND.n4074 GND.n4073 585
R20785 GND.n4076 GND.n4075 585
R20786 GND.n4078 GND.n4077 585
R20787 GND.n5278 GND.n3724 585
R20788 GND.n5894 GND.n3724 585
R20789 GND.n5281 GND.n5280 585
R20790 GND.n5280 GND.n5279 585
R20791 GND.n5282 GND.n3732 585
R20792 GND.n5888 GND.n3732 585
R20793 GND.n5284 GND.n5283 585
R20794 GND.n5284 GND.n3734 585
R20795 GND.n5286 GND.n5285 585
R20796 GND.n5285 GND.n3742 585
R20797 GND.n5287 GND.n3744 585
R20798 GND.n5880 GND.n3744 585
R20799 GND.n5290 GND.n5289 585
R20800 GND.n5289 GND.n5288 585
R20801 GND.n5291 GND.n3752 585
R20802 GND.n5874 GND.n3752 585
R20803 GND.n5293 GND.n5292 585
R20804 GND.n5293 GND.n3754 585
R20805 GND.n5295 GND.n5294 585
R20806 GND.n5294 GND.n3760 585
R20807 GND.n5296 GND.n3762 585
R20808 GND.n5866 GND.n3762 585
R20809 GND.n5299 GND.n5298 585
R20810 GND.n5298 GND.n5297 585
R20811 GND.n5300 GND.n3770 585
R20812 GND.n5860 GND.n3770 585
R20813 GND.n5302 GND.n5301 585
R20814 GND.n5302 GND.n3772 585
R20815 GND.n5304 GND.n5303 585
R20816 GND.n5303 GND.n3778 585
R20817 GND.n5305 GND.n3780 585
R20818 GND.n5852 GND.n3780 585
R20819 GND.n5308 GND.n5307 585
R20820 GND.n5307 GND.n5306 585
R20821 GND.n5309 GND.n3788 585
R20822 GND.n5846 GND.n3788 585
R20823 GND.n5311 GND.n5310 585
R20824 GND.n5313 GND.n5171 585
R20825 GND.n5315 GND.n5314 585
R20826 GND.n5316 GND.n5170 585
R20827 GND.n5318 GND.n5317 585
R20828 GND.n5320 GND.n5168 585
R20829 GND.n5322 GND.n5321 585
R20830 GND.n5323 GND.n5167 585
R20831 GND.n5325 GND.n5324 585
R20832 GND.n5327 GND.n5165 585
R20833 GND.n5329 GND.n5328 585
R20834 GND.n5330 GND.n5164 585
R20835 GND.n5332 GND.n5331 585
R20836 GND.n5334 GND.n5163 585
R20837 GND.n5335 GND.n5036 585
R20838 GND.n5338 GND.n5337 585
R20839 GND.n5162 GND.n5037 585
R20840 GND.n5160 GND.n5159 585
R20841 GND.n5041 GND.n5040 585
R20842 GND.n5152 GND.n5151 585
R20843 GND.n5149 GND.n5043 585
R20844 GND.n5147 GND.n5146 585
R20845 GND.n5045 GND.n5044 585
R20846 GND.n5140 GND.n5139 585
R20847 GND.n5137 GND.n5047 585
R20848 GND.n5135 GND.n5134 585
R20849 GND.n5087 GND.n5048 585
R20850 GND.n5086 GND.n5085 585
R20851 GND.n5083 GND.n5049 585
R20852 GND.n5081 GND.n5080 585
R20853 GND.n5079 GND.n5050 585
R20854 GND.n5078 GND.n5077 585
R20855 GND.n5075 GND.n5051 585
R20856 GND.n5073 GND.n5072 585
R20857 GND.n5071 GND.n5052 585
R20858 GND.n5070 GND.n5069 585
R20859 GND.n5067 GND.n5053 585
R20860 GND.n5065 GND.n5064 585
R20861 GND.n5063 GND.n5054 585
R20862 GND.n5062 GND.n5061 585
R20863 GND.n5059 GND.n5055 585
R20864 GND.n5057 GND.n5056 585
R20865 GND.n3786 GND.n3785 585
R20866 GND.n3789 GND.n3786 585
R20867 GND.n5848 GND.n5847 585
R20868 GND.n5847 GND.n5846 585
R20869 GND.n5849 GND.n3783 585
R20870 GND.n5306 GND.n3783 585
R20871 GND.n5851 GND.n5850 585
R20872 GND.n5852 GND.n5851 585
R20873 GND.n3784 GND.n3782 585
R20874 GND.n3782 GND.n3778 585
R20875 GND.n3768 GND.n3767 585
R20876 GND.n3772 GND.n3768 585
R20877 GND.n5862 GND.n5861 585
R20878 GND.n5861 GND.n5860 585
R20879 GND.n5863 GND.n3765 585
R20880 GND.n5297 GND.n3765 585
R20881 GND.n5865 GND.n5864 585
R20882 GND.n5866 GND.n5865 585
R20883 GND.n3766 GND.n3764 585
R20884 GND.n3764 GND.n3760 585
R20885 GND.n3750 GND.n3749 585
R20886 GND.n3754 GND.n3750 585
R20887 GND.n5876 GND.n5875 585
R20888 GND.n5875 GND.n5874 585
R20889 GND.n5877 GND.n3747 585
R20890 GND.n5288 GND.n3747 585
R20891 GND.n5879 GND.n5878 585
R20892 GND.n5880 GND.n5879 585
R20893 GND.n3748 GND.n3746 585
R20894 GND.n3746 GND.n3742 585
R20895 GND.n3730 GND.n3729 585
R20896 GND.n3734 GND.n3730 585
R20897 GND.n5890 GND.n5889 585
R20898 GND.n5889 GND.n5888 585
R20899 GND.n5891 GND.n3727 585
R20900 GND.n5279 GND.n3727 585
R20901 GND.n5893 GND.n5892 585
R20902 GND.n5894 GND.n5893 585
R20903 GND.n3728 GND.n3726 585
R20904 GND.n5196 GND.n5195 585
R20905 GND.n5197 GND.n5193 585
R20906 GND.n5193 GND.n3717 585
R20907 GND.n5199 GND.n5198 585
R20908 GND.n5201 GND.n5192 585
R20909 GND.n5204 GND.n5203 585
R20910 GND.n5205 GND.n5191 585
R20911 GND.n5207 GND.n5206 585
R20912 GND.n5209 GND.n5190 585
R20913 GND.n5212 GND.n5211 585
R20914 GND.n5213 GND.n5189 585
R20915 GND.n5215 GND.n5214 585
R20916 GND.n5217 GND.n5188 585
R20917 GND.n5220 GND.n5219 585
R20918 GND.n5221 GND.n5187 585
R20919 GND.n5223 GND.n5222 585
R20920 GND.n5225 GND.n5186 585
R20921 GND.n5228 GND.n5227 585
R20922 GND.n5229 GND.n5185 585
R20923 GND.n5231 GND.n5230 585
R20924 GND.n5233 GND.n5184 585
R20925 GND.n5236 GND.n5235 585
R20926 GND.n5237 GND.n5183 585
R20927 GND.n5239 GND.n5238 585
R20928 GND.n5241 GND.n5182 585
R20929 GND.n5244 GND.n5243 585
R20930 GND.n5245 GND.n5181 585
R20931 GND.n5247 GND.n5246 585
R20932 GND.n5249 GND.n5180 585
R20933 GND.n5252 GND.n5251 585
R20934 GND.n5253 GND.n5179 585
R20935 GND.n5255 GND.n5254 585
R20936 GND.n5257 GND.n5178 585
R20937 GND.n5260 GND.n5259 585
R20938 GND.n5261 GND.n5177 585
R20939 GND.n5263 GND.n5262 585
R20940 GND.n5265 GND.n5176 585
R20941 GND.n5268 GND.n5267 585
R20942 GND.n5269 GND.n5175 585
R20943 GND.n5271 GND.n5270 585
R20944 GND.n5273 GND.n5174 585
R20945 GND.n5274 GND.n5173 585
R20946 GND.n5277 GND.n5276 585
R20947 GND.n5896 GND.n3722 585
R20948 GND.n5896 GND.n5895 585
R20949 GND.n3953 GND.n3723 585
R20950 GND.n3725 GND.n3723 585
R20951 GND.n3955 GND.n3954 585
R20952 GND.n3954 GND.n3731 585
R20953 GND.n3956 GND.n3733 585
R20954 GND.n5887 GND.n3733 585
R20955 GND.n3959 GND.n3958 585
R20956 GND.n3958 GND.n3957 585
R20957 GND.n3960 GND.n3743 585
R20958 GND.n5881 GND.n3743 585
R20959 GND.n3962 GND.n3961 585
R20960 GND.n3962 GND.n3745 585
R20961 GND.n3964 GND.n3963 585
R20962 GND.n3963 GND.n3751 585
R20963 GND.n3965 GND.n3753 585
R20964 GND.n5873 GND.n3753 585
R20965 GND.n3968 GND.n3967 585
R20966 GND.n3967 GND.n3966 585
R20967 GND.n3969 GND.n3761 585
R20968 GND.n5867 GND.n3761 585
R20969 GND.n3971 GND.n3970 585
R20970 GND.n3971 GND.n3763 585
R20971 GND.n3973 GND.n3972 585
R20972 GND.n3972 GND.n3769 585
R20973 GND.n3974 GND.n3771 585
R20974 GND.n5859 GND.n3771 585
R20975 GND.n3977 GND.n3976 585
R20976 GND.n3976 GND.n3975 585
R20977 GND.n3978 GND.n3779 585
R20978 GND.n5853 GND.n3779 585
R20979 GND.n3980 GND.n3979 585
R20980 GND.n3980 GND.n3781 585
R20981 GND.n3981 GND.n3952 585
R20982 GND.n3981 GND.n3787 585
R20983 GND.n3983 GND.n3982 585
R20984 GND.n3985 GND.n3984 585
R20985 GND.n3987 GND.n3986 585
R20986 GND.n3989 GND.n3988 585
R20987 GND.n3991 GND.n3990 585
R20988 GND.n3993 GND.n3992 585
R20989 GND.n3995 GND.n3994 585
R20990 GND.n3997 GND.n3996 585
R20991 GND.n3999 GND.n3998 585
R20992 GND.n4001 GND.n4000 585
R20993 GND.n4003 GND.n4002 585
R20994 GND.n4005 GND.n4004 585
R20995 GND.n4007 GND.n4006 585
R20996 GND.n4009 GND.n4008 585
R20997 GND.n4011 GND.n4010 585
R20998 GND.n4013 GND.n4012 585
R20999 GND.n4015 GND.n4014 585
R21000 GND.n4043 GND.n4042 585
R21001 GND.n4041 GND.n4038 585
R21002 GND.n4037 GND.n4036 585
R21003 GND.n4035 GND.n4032 585
R21004 GND.n4031 GND.n4030 585
R21005 GND.n4029 GND.n4026 585
R21006 GND.n4025 GND.n4024 585
R21007 GND.n4023 GND.n4020 585
R21008 GND.n4019 GND.n4018 585
R21009 GND.n4017 GND.n3814 585
R21010 GND.n5815 GND.n5814 585
R21011 GND.n5817 GND.n5816 585
R21012 GND.n5819 GND.n5818 585
R21013 GND.n5821 GND.n5820 585
R21014 GND.n5823 GND.n5822 585
R21015 GND.n5825 GND.n5824 585
R21016 GND.n5827 GND.n5826 585
R21017 GND.n5829 GND.n5828 585
R21018 GND.n5831 GND.n5830 585
R21019 GND.n5833 GND.n5832 585
R21020 GND.n5835 GND.n5834 585
R21021 GND.n5837 GND.n5836 585
R21022 GND.n5839 GND.n5838 585
R21023 GND.n5841 GND.n5840 585
R21024 GND.n5842 GND.n3812 585
R21025 GND.n5844 GND.n5843 585
R21026 GND.n5845 GND.n5844 585
R21027 GND.n3813 GND.n3811 585
R21028 GND.n3811 GND.n3787 585
R21029 GND.n3777 GND.n3776 585
R21030 GND.n3781 GND.n3777 585
R21031 GND.n5855 GND.n5854 585
R21032 GND.n5854 GND.n5853 585
R21033 GND.n5856 GND.n3774 585
R21034 GND.n3975 GND.n3774 585
R21035 GND.n5858 GND.n5857 585
R21036 GND.n5859 GND.n5858 585
R21037 GND.n3775 GND.n3773 585
R21038 GND.n3773 GND.n3769 585
R21039 GND.n3759 GND.n3758 585
R21040 GND.n3763 GND.n3759 585
R21041 GND.n5869 GND.n5868 585
R21042 GND.n5868 GND.n5867 585
R21043 GND.n5870 GND.n3756 585
R21044 GND.n3966 GND.n3756 585
R21045 GND.n5872 GND.n5871 585
R21046 GND.n5873 GND.n5872 585
R21047 GND.n3757 GND.n3755 585
R21048 GND.n3755 GND.n3751 585
R21049 GND.n3741 GND.n3740 585
R21050 GND.n3745 GND.n3741 585
R21051 GND.n5883 GND.n5882 585
R21052 GND.n5882 GND.n5881 585
R21053 GND.n5884 GND.n3736 585
R21054 GND.n3957 GND.n3736 585
R21055 GND.n5886 GND.n5885 585
R21056 GND.n5887 GND.n5886 585
R21057 GND.n3739 GND.n3735 585
R21058 GND.n3735 GND.n3731 585
R21059 GND.n3738 GND.n3737 585
R21060 GND.n3737 GND.n3725 585
R21061 GND.n3721 GND.n3720 585
R21062 GND.n5895 GND.n3720 585
R21063 GND.n5980 GND.n5979 585
R21064 GND.n5978 GND.n3719 585
R21065 GND.n5977 GND.n3718 585
R21066 GND.n5982 GND.n3718 585
R21067 GND.n5976 GND.n5975 585
R21068 GND.n5974 GND.n5973 585
R21069 GND.n5972 GND.n5971 585
R21070 GND.n5970 GND.n5969 585
R21071 GND.n5968 GND.n5967 585
R21072 GND.n5966 GND.n5965 585
R21073 GND.n5964 GND.n5963 585
R21074 GND.n5962 GND.n5961 585
R21075 GND.n5960 GND.n5959 585
R21076 GND.n5958 GND.n5957 585
R21077 GND.n5956 GND.n5955 585
R21078 GND.n5954 GND.n5953 585
R21079 GND.n5952 GND.n5951 585
R21080 GND.n5950 GND.n5949 585
R21081 GND.n5948 GND.n5947 585
R21082 GND.n5946 GND.n5945 585
R21083 GND.n5944 GND.n5943 585
R21084 GND.n5942 GND.n5941 585
R21085 GND.n5940 GND.n5939 585
R21086 GND.n5938 GND.n5937 585
R21087 GND.n5936 GND.n5935 585
R21088 GND.n5934 GND.n5933 585
R21089 GND.n5932 GND.n5931 585
R21090 GND.n5930 GND.n5929 585
R21091 GND.n5928 GND.n5927 585
R21092 GND.n5926 GND.n5925 585
R21093 GND.n5924 GND.n5923 585
R21094 GND.n5922 GND.n5921 585
R21095 GND.n5920 GND.n5919 585
R21096 GND.n5918 GND.n5917 585
R21097 GND.n5916 GND.n5915 585
R21098 GND.n5914 GND.n5913 585
R21099 GND.n5912 GND.n5911 585
R21100 GND.n5910 GND.n5909 585
R21101 GND.n5908 GND.n5907 585
R21102 GND.n5906 GND.n5905 585
R21103 GND.n5904 GND.n5903 585
R21104 GND.n5902 GND.n5901 585
R21105 GND.n5900 GND.n5899 585
R21106 GND.n5898 GND.n5897 585
R21107 GND.n2766 GND.n2765 585
R21108 GND.n2767 GND.n2766 585
R21109 GND.n6269 GND.n6268 585
R21110 GND.n6268 GND.n6267 585
R21111 GND.n6270 GND.n2764 585
R21112 GND.n2764 GND.n2763 585
R21113 GND.n6272 GND.n6271 585
R21114 GND.n6273 GND.n6272 585
R21115 GND.n2758 GND.n2757 585
R21116 GND.n2759 GND.n2758 585
R21117 GND.n6281 GND.n6280 585
R21118 GND.n6280 GND.n6279 585
R21119 GND.n6282 GND.n2756 585
R21120 GND.n2756 GND.n2755 585
R21121 GND.n6284 GND.n6283 585
R21122 GND.n6286 GND.n6284 585
R21123 GND.n2751 GND.n2750 585
R21124 GND.n6285 GND.n2751 585
R21125 GND.n6294 GND.n6293 585
R21126 GND.n6293 GND.n6292 585
R21127 GND.n6295 GND.n2749 585
R21128 GND.n2749 GND.n2748 585
R21129 GND.n6297 GND.n6296 585
R21130 GND.n6298 GND.n6297 585
R21131 GND.n2743 GND.n2742 585
R21132 GND.n2744 GND.n2743 585
R21133 GND.n6306 GND.n6305 585
R21134 GND.n6305 GND.n6304 585
R21135 GND.n6307 GND.n2741 585
R21136 GND.n2741 GND.n2740 585
R21137 GND.n6310 GND.n6309 585
R21138 GND.n6311 GND.n6310 585
R21139 GND.n6308 GND.n2734 585
R21140 GND.n2735 GND.n2734 585
R21141 GND.n6389 GND.n2732 585
R21142 GND.n6389 GND.n6388 585
R21143 GND.n6391 GND.n6390 585
R21144 GND.n6392 GND.n2731 585
R21145 GND.n6394 GND.n6393 585
R21146 GND.n6396 GND.n2729 585
R21147 GND.n6398 GND.n6397 585
R21148 GND.n6399 GND.n2728 585
R21149 GND.n6401 GND.n6400 585
R21150 GND.n6403 GND.n2726 585
R21151 GND.n6405 GND.n6404 585
R21152 GND.n6406 GND.n2725 585
R21153 GND.n6408 GND.n6407 585
R21154 GND.n6410 GND.n2723 585
R21155 GND.n6412 GND.n6411 585
R21156 GND.n6413 GND.n2722 585
R21157 GND.n6415 GND.n6414 585
R21158 GND.n6417 GND.n2721 585
R21159 GND.n6418 GND.n2718 585
R21160 GND.n6421 GND.n6420 585
R21161 GND.n2719 GND.n2717 585
R21162 GND.n6338 GND.n6336 585
R21163 GND.n6342 GND.n6341 585
R21164 GND.n6344 GND.n6334 585
R21165 GND.n6345 GND.n6331 585
R21166 GND.n6348 GND.n6347 585
R21167 GND.n6333 GND.n6330 585
R21168 GND.n6327 GND.n6326 585
R21169 GND.n6357 GND.n6356 585
R21170 GND.n6359 GND.n6324 585
R21171 GND.n6361 GND.n6360 585
R21172 GND.n6362 GND.n6323 585
R21173 GND.n6364 GND.n6363 585
R21174 GND.n6366 GND.n6321 585
R21175 GND.n6368 GND.n6367 585
R21176 GND.n6369 GND.n6320 585
R21177 GND.n6371 GND.n6370 585
R21178 GND.n6373 GND.n6318 585
R21179 GND.n6375 GND.n6374 585
R21180 GND.n6376 GND.n6317 585
R21181 GND.n6378 GND.n6377 585
R21182 GND.n6380 GND.n6316 585
R21183 GND.n6381 GND.n6315 585
R21184 GND.n6384 GND.n6383 585
R21185 GND.n6385 GND.n2737 585
R21186 GND.n2737 GND.n2720 585
R21187 GND.n6387 GND.n6386 585
R21188 GND.n6388 GND.n6387 585
R21189 GND.n6314 GND.n2736 585
R21190 GND.n2736 GND.n2735 585
R21191 GND.n6313 GND.n6312 585
R21192 GND.n6312 GND.n6311 585
R21193 GND.n2739 GND.n2738 585
R21194 GND.n2740 GND.n2739 585
R21195 GND.n6303 GND.n6302 585
R21196 GND.n6304 GND.n6303 585
R21197 GND.n6301 GND.n2745 585
R21198 GND.n2745 GND.n2744 585
R21199 GND.n6300 GND.n6299 585
R21200 GND.n6299 GND.n6298 585
R21201 GND.n2747 GND.n2746 585
R21202 GND.n2748 GND.n2747 585
R21203 GND.n6291 GND.n6290 585
R21204 GND.n6292 GND.n6291 585
R21205 GND.n6289 GND.n2752 585
R21206 GND.n6285 GND.n2752 585
R21207 GND.n6288 GND.n6287 585
R21208 GND.n6287 GND.n6286 585
R21209 GND.n2754 GND.n2753 585
R21210 GND.n2755 GND.n2754 585
R21211 GND.n6278 GND.n6277 585
R21212 GND.n6279 GND.n6278 585
R21213 GND.n6276 GND.n2760 585
R21214 GND.n2760 GND.n2759 585
R21215 GND.n6275 GND.n6274 585
R21216 GND.n6274 GND.n6273 585
R21217 GND.n2762 GND.n2761 585
R21218 GND.n2763 GND.n2762 585
R21219 GND.n6266 GND.n6265 585
R21220 GND.n6267 GND.n6266 585
R21221 GND.n6264 GND.n2768 585
R21222 GND.n2768 GND.n2767 585
R21223 GND.n6263 GND.n6262 585
R21224 GND.n2770 GND.n2769 585
R21225 GND.n6259 GND.n6258 585
R21226 GND.n6260 GND.n6259 585
R21227 GND.n6257 GND.n2792 585
R21228 GND.n6256 GND.n6255 585
R21229 GND.n6254 GND.n6253 585
R21230 GND.n6252 GND.n6251 585
R21231 GND.n6250 GND.n6249 585
R21232 GND.n6248 GND.n6247 585
R21233 GND.n6246 GND.n6245 585
R21234 GND.n6244 GND.n6243 585
R21235 GND.n6242 GND.n6241 585
R21236 GND.n6240 GND.n6239 585
R21237 GND.n6238 GND.n6237 585
R21238 GND.n6236 GND.n6235 585
R21239 GND.n6234 GND.n6233 585
R21240 GND.n6231 GND.n2794 585
R21241 GND.n2796 GND.n2795 585
R21242 GND.n6226 GND.n2799 585
R21243 GND.n6225 GND.n2800 585
R21244 GND.n6224 GND.n2801 585
R21245 GND.n2803 GND.n2802 585
R21246 GND.n6219 GND.n2806 585
R21247 GND.n6218 GND.n2807 585
R21248 GND.n6217 GND.n2808 585
R21249 GND.n2810 GND.n2809 585
R21250 GND.n2846 GND.n2845 585
R21251 GND.n2844 GND.n2843 585
R21252 GND.n2842 GND.n2841 585
R21253 GND.n2840 GND.n2839 585
R21254 GND.n2838 GND.n2837 585
R21255 GND.n2836 GND.n2835 585
R21256 GND.n2834 GND.n2833 585
R21257 GND.n2832 GND.n2831 585
R21258 GND.n2830 GND.n2829 585
R21259 GND.n2828 GND.n2827 585
R21260 GND.n2826 GND.n2825 585
R21261 GND.n2824 GND.n2823 585
R21262 GND.n2822 GND.n2821 585
R21263 GND.n2820 GND.n2819 585
R21264 GND.n2818 GND.n2817 585
R21265 GND.n2816 GND.n2815 585
R21266 GND.n2814 GND.n2813 585
R21267 GND.n6095 GND.n6094 585
R21268 GND.n6094 GND.n6093 585
R21269 GND.n6096 GND.n3114 585
R21270 GND.n5985 GND.n3114 585
R21271 GND.n6098 GND.n6097 585
R21272 GND.n6099 GND.n6098 585
R21273 GND.n2887 GND.n2886 585
R21274 GND.n2888 GND.n2887 585
R21275 GND.n6107 GND.n6106 585
R21276 GND.n6106 GND.n6105 585
R21277 GND.n6108 GND.n2885 585
R21278 GND.n2885 GND.n2884 585
R21279 GND.n6110 GND.n6109 585
R21280 GND.n6111 GND.n6110 585
R21281 GND.n2879 GND.n2878 585
R21282 GND.n2880 GND.n2879 585
R21283 GND.n6119 GND.n6118 585
R21284 GND.n6118 GND.n6117 585
R21285 GND.n6120 GND.n2877 585
R21286 GND.n2877 GND.n2876 585
R21287 GND.n6122 GND.n6121 585
R21288 GND.n6123 GND.n6122 585
R21289 GND.n2871 GND.n2870 585
R21290 GND.n2872 GND.n2871 585
R21291 GND.n6131 GND.n6130 585
R21292 GND.n6130 GND.n6129 585
R21293 GND.n6132 GND.n2869 585
R21294 GND.n2869 GND.n2868 585
R21295 GND.n6134 GND.n6133 585
R21296 GND.n6135 GND.n6134 585
R21297 GND.n2861 GND.n2860 585
R21298 GND.n2862 GND.n2861 585
R21299 GND.n6182 GND.n6181 585
R21300 GND.n6181 GND.n6180 585
R21301 GND.n6183 GND.n2859 585
R21302 GND.n2863 GND.n2859 585
R21303 GND.n6185 GND.n6184 585
R21304 GND.n6187 GND.n2857 585
R21305 GND.n6189 GND.n6188 585
R21306 GND.n6190 GND.n2856 585
R21307 GND.n6192 GND.n6191 585
R21308 GND.n6194 GND.n2854 585
R21309 GND.n6196 GND.n6195 585
R21310 GND.n6197 GND.n2853 585
R21311 GND.n6199 GND.n6198 585
R21312 GND.n6201 GND.n2851 585
R21313 GND.n6203 GND.n6202 585
R21314 GND.n6204 GND.n2850 585
R21315 GND.n6206 GND.n6205 585
R21316 GND.n6208 GND.n2848 585
R21317 GND.n6210 GND.n6209 585
R21318 GND.n6211 GND.n2812 585
R21319 GND.n6213 GND.n6212 585
R21320 GND.n6215 GND.n2810 585
R21321 GND.n6217 GND.n6216 585
R21322 GND.n6218 GND.n2805 585
R21323 GND.n6220 GND.n6219 585
R21324 GND.n6222 GND.n2803 585
R21325 GND.n6224 GND.n6223 585
R21326 GND.n6225 GND.n2798 585
R21327 GND.n6227 GND.n6226 585
R21328 GND.n6229 GND.n2796 585
R21329 GND.n6231 GND.n6230 585
R21330 GND.n6149 GND.n2793 585
R21331 GND.n6151 GND.n6150 585
R21332 GND.n6153 GND.n6147 585
R21333 GND.n6155 GND.n6154 585
R21334 GND.n6156 GND.n6146 585
R21335 GND.n6158 GND.n6157 585
R21336 GND.n6160 GND.n6144 585
R21337 GND.n6162 GND.n6161 585
R21338 GND.n6163 GND.n6143 585
R21339 GND.n6165 GND.n6164 585
R21340 GND.n6167 GND.n6141 585
R21341 GND.n6169 GND.n6168 585
R21342 GND.n6170 GND.n6140 585
R21343 GND.n6172 GND.n6171 585
R21344 GND.n6174 GND.n6139 585
R21345 GND.n6176 GND.n6175 585
R21346 GND.n6175 GND.n2771 585
R21347 GND.n6177 GND.n2865 585
R21348 GND.n2865 GND.n2863 585
R21349 GND.n6179 GND.n6178 585
R21350 GND.n6180 GND.n6179 585
R21351 GND.n6138 GND.n2864 585
R21352 GND.n2864 GND.n2862 585
R21353 GND.n6137 GND.n6136 585
R21354 GND.n6136 GND.n6135 585
R21355 GND.n2867 GND.n2866 585
R21356 GND.n2868 GND.n2867 585
R21357 GND.n6128 GND.n6127 585
R21358 GND.n6129 GND.n6128 585
R21359 GND.n6126 GND.n2873 585
R21360 GND.n2873 GND.n2872 585
R21361 GND.n6125 GND.n6124 585
R21362 GND.n6124 GND.n6123 585
R21363 GND.n2875 GND.n2874 585
R21364 GND.n2876 GND.n2875 585
R21365 GND.n6116 GND.n6115 585
R21366 GND.n6117 GND.n6116 585
R21367 GND.n6114 GND.n2881 585
R21368 GND.n2881 GND.n2880 585
R21369 GND.n6113 GND.n6112 585
R21370 GND.n6112 GND.n6111 585
R21371 GND.n2883 GND.n2882 585
R21372 GND.n2884 GND.n2883 585
R21373 GND.n6104 GND.n6103 585
R21374 GND.n6105 GND.n6104 585
R21375 GND.n6102 GND.n2889 585
R21376 GND.n2889 GND.n2888 585
R21377 GND.n6101 GND.n6100 585
R21378 GND.n6100 GND.n6099 585
R21379 GND.n2891 GND.n2890 585
R21380 GND.n5985 GND.n2891 585
R21381 GND.n6092 GND.n6091 585
R21382 GND.n6093 GND.n6092 585
R21383 GND.n6090 GND.n5986 585
R21384 GND.n6089 GND.n6088 585
R21385 GND.n6086 GND.n5987 585
R21386 GND.n6086 GND.n5984 585
R21387 GND.n6085 GND.n6084 585
R21388 GND.n6083 GND.n6082 585
R21389 GND.n6081 GND.n5989 585
R21390 GND.n6079 GND.n6078 585
R21391 GND.n6077 GND.n5990 585
R21392 GND.n6076 GND.n6075 585
R21393 GND.n6073 GND.n5991 585
R21394 GND.n6071 GND.n6070 585
R21395 GND.n6069 GND.n5992 585
R21396 GND.n6068 GND.n6067 585
R21397 GND.n6065 GND.n5993 585
R21398 GND.n6063 GND.n6062 585
R21399 GND.n6061 GND.n5994 585
R21400 GND.n6060 GND.n6059 585
R21401 GND.n6057 GND.n5995 585
R21402 GND.n6055 GND.n6054 585
R21403 GND.n6053 GND.n5996 585
R21404 GND.n6052 GND.n6051 585
R21405 GND.n6049 GND.n5997 585
R21406 GND.n6047 GND.n6046 585
R21407 GND.n6045 GND.n5998 585
R21408 GND.n6044 GND.n6043 585
R21409 GND.n6041 GND.n5999 585
R21410 GND.n6039 GND.n6038 585
R21411 GND.n6037 GND.n6000 585
R21412 GND.n6036 GND.n6035 585
R21413 GND.n6033 GND.n6001 585
R21414 GND.n6031 GND.n6030 585
R21415 GND.n6029 GND.n6002 585
R21416 GND.n6028 GND.n6027 585
R21417 GND.n6025 GND.n6003 585
R21418 GND.n6023 GND.n6022 585
R21419 GND.n6021 GND.n6004 585
R21420 GND.n6020 GND.n6019 585
R21421 GND.n6017 GND.n6005 585
R21422 GND.n6015 GND.n6014 585
R21423 GND.n6013 GND.n6006 585
R21424 GND.n6012 GND.n6011 585
R21425 GND.n6009 GND.n6007 585
R21426 GND.n3116 GND.n3115 585
R21427 GND.n7586 GND.n2408 585
R21428 GND.n7585 GND.n7584 585
R21429 GND.n2410 GND.n2409 585
R21430 GND.n7582 GND.n2410 585
R21431 GND.n5565 GND.n5564 585
R21432 GND.n5567 GND.n5566 585
R21433 GND.n5569 GND.n5568 585
R21434 GND.n5571 GND.n5570 585
R21435 GND.n5573 GND.n5572 585
R21436 GND.n5575 GND.n5574 585
R21437 GND.n5577 GND.n5576 585
R21438 GND.n5579 GND.n5578 585
R21439 GND.n5581 GND.n5580 585
R21440 GND.n5583 GND.n5582 585
R21441 GND.n5585 GND.n5584 585
R21442 GND.n5587 GND.n5586 585
R21443 GND.n5589 GND.n5588 585
R21444 GND.n5591 GND.n5590 585
R21445 GND.n5592 GND.n2407 585
R21446 GND.n7589 GND.n2407 585
R21447 GND.n5593 GND.n2406 585
R21448 GND.n7590 GND.n2406 585
R21449 GND.n5594 GND.n2405 585
R21450 GND.n7591 GND.n2405 585
R21451 GND.n5596 GND.n5595 585
R21452 GND.n5595 GND.n5558 585
R21453 GND.n5597 GND.n2398 585
R21454 GND.n7597 GND.n2398 585
R21455 GND.n5599 GND.n5598 585
R21456 GND.n5599 GND.n2396 585
R21457 GND.n5601 GND.n5600 585
R21458 GND.n5600 GND.n2390 585
R21459 GND.n5602 GND.n2388 585
R21460 GND.n7605 GND.n2388 585
R21461 GND.n5604 GND.n5603 585
R21462 GND.n5605 GND.n5604 585
R21463 GND.n5563 GND.n2380 585
R21464 GND.n7611 GND.n2380 585
R21465 GND.n5662 GND.n5446 585
R21466 GND.n5662 GND.n5661 585
R21467 GND.n5664 GND.n5663 585
R21468 GND.n5663 GND.n2368 585
R21469 GND.n5445 GND.n5444 585
R21470 GND.n5445 GND.n2365 585
R21471 GND.n5509 GND.n5508 585
R21472 GND.n5508 GND.n5461 585
R21473 GND.n5510 GND.n2357 585
R21474 GND.n7626 GND.n2357 585
R21475 GND.n5512 GND.n5511 585
R21476 GND.n5513 GND.n5512 585
R21477 GND.n5507 GND.n2347 585
R21478 GND.n7632 GND.n2347 585
R21479 GND.n5506 GND.n5505 585
R21480 GND.n5505 GND.n2345 585
R21481 GND.n5504 GND.n5503 585
R21482 GND.n5504 GND.n2339 585
R21483 GND.n5502 GND.n2337 585
R21484 GND.n7640 GND.n2337 585
R21485 GND.n5501 GND.n2336 585
R21486 GND.n7641 GND.n2336 585
R21487 GND.n5500 GND.n2329 585
R21488 GND.n2331 GND.n2329 585
R21489 GND.n7648 GND.n2330 585
R21490 GND.n7648 GND.n7647 585
R21491 GND.n7649 GND.n2328 585
R21492 GND.n7649 GND.n2316 585
R21493 GND.n7651 GND.n7650 585
R21494 GND.n7653 GND.n7652 585
R21495 GND.n7655 GND.n7654 585
R21496 GND.n7657 GND.n7656 585
R21497 GND.n7659 GND.n7658 585
R21498 GND.n7661 GND.n7660 585
R21499 GND.n7663 GND.n7662 585
R21500 GND.n7665 GND.n7664 585
R21501 GND.n7667 GND.n7666 585
R21502 GND.n7669 GND.n7668 585
R21503 GND.n7671 GND.n7670 585
R21504 GND.n7673 GND.n7672 585
R21505 GND.n7675 GND.n7674 585
R21506 GND.n7677 GND.n7676 585
R21507 GND.n7679 GND.n7678 585
R21508 GND.n7680 GND.n2326 585
R21509 GND.n7682 GND.n7681 585
R21510 GND.n7683 GND.n7682 585
R21511 GND.n2327 GND.n2325 585
R21512 GND.n2325 GND.n2316 585
R21513 GND.n7646 GND.n7645 585
R21514 GND.n7647 GND.n7646 585
R21515 GND.n7644 GND.n2332 585
R21516 GND.n2332 GND.n2331 585
R21517 GND.n7643 GND.n7642 585
R21518 GND.n7642 GND.n7641 585
R21519 GND.n2334 GND.n2333 585
R21520 GND.n7640 GND.n2334 585
R21521 GND.n2352 GND.n2351 585
R21522 GND.n2351 GND.n2339 585
R21523 GND.n2353 GND.n2349 585
R21524 GND.n2349 GND.n2345 585
R21525 GND.n7631 GND.n7630 585
R21526 GND.n7632 GND.n7631 585
R21527 GND.n7629 GND.n2350 585
R21528 GND.n5513 GND.n2350 585
R21529 GND.n7628 GND.n7627 585
R21530 GND.n7627 GND.n7626 585
R21531 GND.n2355 GND.n2354 585
R21532 GND.n5461 GND.n2355 585
R21533 GND.n5455 GND.n5454 585
R21534 GND.n5454 GND.n2365 585
R21535 GND.n5453 GND.n5452 585
R21536 GND.n5453 GND.n2368 585
R21537 GND.n2384 GND.n2382 585
R21538 GND.n5661 GND.n2382 585
R21539 GND.n7610 GND.n7609 585
R21540 GND.n7611 GND.n7610 585
R21541 GND.n7608 GND.n2383 585
R21542 GND.n5605 GND.n2383 585
R21543 GND.n7607 GND.n7606 585
R21544 GND.n7606 GND.n7605 585
R21545 GND.n2386 GND.n2385 585
R21546 GND.n2390 GND.n2386 585
R21547 GND.n2402 GND.n2400 585
R21548 GND.n2400 GND.n2396 585
R21549 GND.n7596 GND.n7595 585
R21550 GND.n7597 GND.n7596 585
R21551 GND.n7594 GND.n2401 585
R21552 GND.n5558 GND.n2401 585
R21553 GND.n7593 GND.n7592 585
R21554 GND.n7592 GND.n7591 585
R21555 GND.n2404 GND.n2403 585
R21556 GND.n7590 GND.n2404 585
R21557 GND.n7588 GND.n7587 585
R21558 GND.n7589 GND.n7588 585
R21559 GND.n5620 GND.n5619 585
R21560 GND.n5618 GND.n5617 585
R21561 GND.n5556 GND.n5554 585
R21562 GND.n5622 GND.n5556 585
R21563 GND.n5625 GND.n5624 585
R21564 GND.n5557 GND.n5555 585
R21565 GND.n5616 GND.n5615 585
R21566 GND.n5622 GND.n5616 585
R21567 GND.n5614 GND.n5559 585
R21568 GND.n5559 GND.n2399 585
R21569 GND.n5613 GND.n2397 585
R21570 GND.n7598 GND.n2397 585
R21571 GND.n5612 GND.n5611 585
R21572 GND.n5611 GND.n5610 585
R21573 GND.n5609 GND.n2389 585
R21574 GND.n7604 GND.n2389 585
R21575 GND.n5608 GND.n5607 585
R21576 GND.n5607 GND.n5606 585
R21577 GND.n5561 GND.n5560 585
R21578 GND.n5562 GND.n5561 585
R21579 GND.n5449 GND.n2379 585
R21580 GND.n7612 GND.n2379 585
R21581 GND.n5659 GND.n5658 585
R21582 GND.n5660 GND.n5659 585
R21583 GND.n5654 GND.n2367 585
R21584 GND.n7618 GND.n2367 585
R21585 GND.n5653 GND.n5652 585
R21586 GND.n5652 GND.n5651 585
R21587 GND.n5460 GND.n5459 585
R21588 GND.n5460 GND.n2359 585
R21589 GND.n5537 GND.n5536 585
R21590 GND.n5537 GND.n2356 585
R21591 GND.n5539 GND.n5538 585
R21592 GND.n5538 GND.n2348 585
R21593 GND.n5540 GND.n2346 585
R21594 GND.n7633 GND.n2346 585
R21595 GND.n5543 GND.n5542 585
R21596 GND.n5542 GND.n5541 585
R21597 GND.n5544 GND.n2338 585
R21598 GND.n7639 GND.n2338 585
R21599 GND.n5546 GND.n5545 585
R21600 GND.n5548 GND.n5530 585
R21601 GND.n5550 GND.n5549 585
R21602 GND.n5534 GND.n5529 585
R21603 GND.n5533 GND.n5532 585
R21604 GND.n2342 GND.n2340 585
R21605 GND.n7638 GND.n7637 585
R21606 GND.n7639 GND.n7638 585
R21607 GND.n7636 GND.n2341 585
R21608 GND.n5541 GND.n2341 585
R21609 GND.n7635 GND.n7634 585
R21610 GND.n7634 GND.n7633 585
R21611 GND.n2344 GND.n2343 585
R21612 GND.n2348 GND.n2344 585
R21613 GND.n2372 GND.n2371 585
R21614 GND.n2372 GND.n2356 585
R21615 GND.n2374 GND.n2373 585
R21616 GND.n2373 GND.n2359 585
R21617 GND.n2375 GND.n2369 585
R21618 GND.n5651 GND.n2369 585
R21619 GND.n7617 GND.n7616 585
R21620 GND.n7618 GND.n7617 585
R21621 GND.n7615 GND.n2370 585
R21622 GND.n5660 GND.n2370 585
R21623 GND.n7614 GND.n7613 585
R21624 GND.n7613 GND.n7612 585
R21625 GND.n2377 GND.n2376 585
R21626 GND.n5562 GND.n2377 585
R21627 GND.n2393 GND.n2391 585
R21628 GND.n5606 GND.n2391 585
R21629 GND.n7603 GND.n7602 585
R21630 GND.n7604 GND.n7603 585
R21631 GND.n7601 GND.n2392 585
R21632 GND.n5610 GND.n2392 585
R21633 GND.n7600 GND.n7599 585
R21634 GND.n7599 GND.n7598 585
R21635 GND.n2395 GND.n2394 585
R21636 GND.n2399 GND.n2395 585
R21637 GND.n5476 GND.n5475 585
R21638 GND.n5478 GND.n5470 585
R21639 GND.n5479 GND.n5469 585
R21640 GND.n5479 GND.n2387 585
R21641 GND.n5482 GND.n5481 585
R21642 GND.n5483 GND.n5467 585
R21643 GND.n5634 GND.n5633 585
R21644 GND.n5636 GND.n5466 585
R21645 GND.n5637 GND.n5465 585
R21646 GND.n5640 GND.n5639 585
R21647 GND.n5641 GND.n5464 585
R21648 GND.n5464 GND.n2387 585
R21649 GND.n5643 GND.n5642 585
R21650 GND.n5643 GND.n2381 585
R21651 GND.n5644 GND.n5463 585
R21652 GND.n5644 GND.n2378 585
R21653 GND.n5646 GND.n5645 585
R21654 GND.n5645 GND.n5447 585
R21655 GND.n5647 GND.n2366 585
R21656 GND.n7619 GND.n2366 585
R21657 GND.n5649 GND.n5648 585
R21658 GND.n5650 GND.n5649 585
R21659 GND.n5462 GND.n2358 585
R21660 GND.n7625 GND.n2358 585
R21661 GND.n5518 GND.n5517 585
R21662 GND.n5519 GND.n5515 585
R21663 GND.n5521 GND.n5520 585
R21664 GND.n5523 GND.n5490 585
R21665 GND.n5525 GND.n5524 585
R21666 GND.n5493 GND.n5488 585
R21667 GND.n5498 GND.n5497 585
R21668 GND.n5496 GND.n5492 585
R21669 GND.n5495 GND.n5494 585
R21670 GND.n2362 GND.n2360 585
R21671 GND.n7624 GND.n7623 585
R21672 GND.n7625 GND.n7624 585
R21673 GND.n7622 GND.n2361 585
R21674 GND.n5650 GND.n2361 585
R21675 GND.n7621 GND.n7620 585
R21676 GND.n7620 GND.n7619 585
R21677 GND.n2364 GND.n2363 585
R21678 GND.n5447 GND.n2364 585
R21679 GND.n5473 GND.n5472 585
R21680 GND.n5472 GND.n2378 585
R21681 GND.n5474 GND.n5471 585
R21682 GND.n5471 GND.n2381 585
R21683 GND.n6944 GND.n6764 585
R21684 GND.n6984 GND.n6764 585
R21685 GND.n6946 GND.n6945 585
R21686 GND.n6945 GND.n6762 585
R21687 GND.n6947 GND.n6768 585
R21688 GND.n6970 GND.n6768 585
R21689 GND.n6950 GND.n6949 585
R21690 GND.n6949 GND.n6948 585
R21691 GND.n6951 GND.n6774 585
R21692 GND.n6963 GND.n6774 585
R21693 GND.n6953 GND.n6952 585
R21694 GND.n6954 GND.n6953 585
R21695 GND.n6923 GND.n6782 585
R21696 GND.n6782 GND.n6780 585
R21697 GND.n6922 GND.n6921 585
R21698 GND.n6921 GND.n6920 585
R21699 GND.n6784 GND.n6783 585
R21700 GND.n6793 GND.n6784 585
R21701 GND.n6873 GND.n6791 585
R21702 GND.n6913 GND.n6791 585
R21703 GND.n6875 GND.n6874 585
R21704 GND.n6877 GND.n6876 585
R21705 GND.n6879 GND.n6878 585
R21706 GND.n6881 GND.n6880 585
R21707 GND.n6883 GND.n6882 585
R21708 GND.n6885 GND.n6884 585
R21709 GND.n6887 GND.n6886 585
R21710 GND.n6889 GND.n6888 585
R21711 GND.n6891 GND.n6890 585
R21712 GND.n6893 GND.n6892 585
R21713 GND.n6895 GND.n6894 585
R21714 GND.n6897 GND.n6896 585
R21715 GND.n6899 GND.n6898 585
R21716 GND.n6900 GND.n6871 585
R21717 GND.n6902 GND.n6901 585
R21718 GND.n6872 GND.n6870 585
R21719 GND.n6789 GND.n6788 585
R21720 GND.n6904 GND.n6789 585
R21721 GND.n6915 GND.n6914 585
R21722 GND.n6914 GND.n6913 585
R21723 GND.n6916 GND.n6786 585
R21724 GND.n6793 GND.n6786 585
R21725 GND.n6919 GND.n6918 585
R21726 GND.n6920 GND.n6919 585
R21727 GND.n6917 GND.n6787 585
R21728 GND.n6787 GND.n6780 585
R21729 GND.n6772 GND.n6771 585
R21730 GND.n6954 GND.n6772 585
R21731 GND.n6965 GND.n6964 585
R21732 GND.n6964 GND.n6963 585
R21733 GND.n6966 GND.n6769 585
R21734 GND.n6948 GND.n6769 585
R21735 GND.n6969 GND.n6968 585
R21736 GND.n6970 GND.n6969 585
R21737 GND.n6967 GND.n6770 585
R21738 GND.n6770 GND.n6762 585
R21739 GND.n6754 GND.n6753 585
R21740 GND.n6984 GND.n6754 585
R21741 GND.n6801 GND.n6800 585
R21742 GND.n6802 GND.n6801 585
R21743 GND.n6813 GND.n6812 585
R21744 GND.n6815 GND.n6811 585
R21745 GND.n6818 GND.n6817 585
R21746 GND.n6819 GND.n6810 585
R21747 GND.n6821 GND.n6820 585
R21748 GND.n6823 GND.n6809 585
R21749 GND.n6826 GND.n6825 585
R21750 GND.n6827 GND.n6808 585
R21751 GND.n6829 GND.n6828 585
R21752 GND.n6831 GND.n6807 585
R21753 GND.n6834 GND.n6833 585
R21754 GND.n6835 GND.n6806 585
R21755 GND.n6837 GND.n6836 585
R21756 GND.n6839 GND.n6805 585
R21757 GND.n6842 GND.n6841 585
R21758 GND.n6843 GND.n6804 585
R21759 GND.n6845 GND.n6844 585
R21760 GND.n6846 GND.n6845 585
R21761 GND.n6797 GND.n6796 585
R21762 GND.n6803 GND.n6797 585
R21763 GND.n6907 GND.n6906 585
R21764 GND.n6906 GND.n6905 585
R21765 GND.n6908 GND.n6794 585
R21766 GND.n6794 GND.n6790 585
R21767 GND.n6911 GND.n6910 585
R21768 GND.n6912 GND.n6911 585
R21769 GND.n6909 GND.n6795 585
R21770 GND.n6795 GND.n6785 585
R21771 GND.n6779 GND.n6778 585
R21772 GND.n6855 GND.n6779 585
R21773 GND.n6957 GND.n6956 585
R21774 GND.n6956 GND.n6955 585
R21775 GND.n6958 GND.n6776 585
R21776 GND.n6776 GND.n6773 585
R21777 GND.n6961 GND.n6960 585
R21778 GND.n6962 GND.n6961 585
R21779 GND.n6959 GND.n6777 585
R21780 GND.n6777 GND.n6767 585
R21781 GND.n6761 GND.n6760 585
R21782 GND.n6971 GND.n6761 585
R21783 GND.n6987 GND.n6986 585
R21784 GND.n6986 GND.n6985 585
R21785 GND.n6988 GND.n6758 585
R21786 GND.n6982 GND.n6758 585
R21787 GND.n6997 GND.n6996 585
R21788 GND.n6998 GND.n6997 585
R21789 GND.n6990 GND.n6759 585
R21790 GND.n6759 GND.n6749 585
R21791 GND.n6991 GND.n6732 585
R21792 GND.n7013 GND.n6732 585
R21793 GND.n7061 GND.n7060 585
R21794 GND.n7062 GND.n7061 585
R21795 GND.n6735 GND.n6733 585
R21796 GND.n6733 GND.n6671 585
R21797 GND.n7055 GND.n7054 585
R21798 GND.n7054 GND.n6675 585
R21799 GND.n7053 GND.n7052 585
R21800 GND.n7053 GND.n6663 585
R21801 GND.n7046 GND.n7045 585
R21802 GND.n7045 GND.n7044 585
R21803 GND.n7047 GND.n6653 585
R21804 GND.n6653 GND.n6648 585
R21805 GND.n7171 GND.n7170 585
R21806 GND.n7172 GND.n7171 585
R21807 GND.n6655 GND.n6631 585
R21808 GND.n6631 GND.n6621 585
R21809 GND.n7200 GND.n7199 585
R21810 GND.n7201 GND.n7200 585
R21811 GND.n2633 GND.n2632 585
R21812 GND.n6611 GND.n2632 585
R21813 GND.n7252 GND.n7251 585
R21814 GND.n7253 GND.n7252 585
R21815 GND.n2634 GND.n2624 585
R21816 GND.n2624 GND.n2558 585
R21817 GND.n7279 GND.n7278 585
R21818 GND.n7278 GND.n7277 585
R21819 GND.n7280 GND.n2619 585
R21820 GND.n2619 GND.n2547 585
R21821 GND.n7287 GND.n7286 585
R21822 GND.n7288 GND.n7287 585
R21823 GND.n2621 GND.n2504 585
R21824 GND.n2518 GND.n2504 585
R21825 GND.n7392 GND.n7391 585
R21826 GND.n7391 GND.n7390 585
R21827 GND.n7393 GND.n2497 585
R21828 GND.n2527 GND.n2497 585
R21829 GND.n7403 GND.n7402 585
R21830 GND.n7404 GND.n7403 585
R21831 GND.n2501 GND.n2499 585
R21832 GND.n2499 GND.n2498 585
R21833 GND.n7397 GND.n2477 585
R21834 GND.n7419 GND.n2477 585
R21835 GND.n7431 GND.n7430 585
R21836 GND.n7430 GND.n7429 585
R21837 GND.n2474 GND.n2472 585
R21838 GND.n2481 GND.n2472 585
R21839 GND.n7437 GND.n7436 585
R21840 GND.n7438 GND.n7437 585
R21841 GND.n7435 GND.n2473 585
R21842 GND.n2473 GND.n2420 585
R21843 GND.n2432 GND.n2430 585
R21844 GND.n2430 GND.n2426 585
R21845 GND.n7572 GND.n7571 585
R21846 GND.n7573 GND.n7572 585
R21847 GND.n7570 GND.n2431 585
R21848 GND.n7444 GND.n2431 585
R21849 GND.n7569 GND.n7568 585
R21850 GND.n7568 GND.n7567 585
R21851 GND.n2434 GND.n2433 585
R21852 GND.n2438 GND.n2434 585
R21853 GND.n2449 GND.n2447 585
R21854 GND.n7511 GND.n2447 585
R21855 GND.n7558 GND.n7557 585
R21856 GND.n7559 GND.n7558 585
R21857 GND.n7556 GND.n2448 585
R21858 GND.n7505 GND.n2448 585
R21859 GND.n7555 GND.n7554 585
R21860 GND.n7554 GND.n7553 585
R21861 GND.n2451 GND.n2450 585
R21862 GND.n2461 GND.n2451 585
R21863 GND.n7499 GND.n7498 585
R21864 GND.n7500 GND.n7499 585
R21865 GND.n7497 GND.n7452 585
R21866 GND.n7452 GND.n7451 585
R21867 GND.n7496 GND.n7495 585
R21868 GND.n7454 GND.n7453 585
R21869 GND.n7492 GND.n7491 585
R21870 GND.n7493 GND.n7492 585
R21871 GND.n7490 GND.n7462 585
R21872 GND.n7489 GND.n7488 585
R21873 GND.n7487 GND.n7486 585
R21874 GND.n7485 GND.n7484 585
R21875 GND.n7483 GND.n7482 585
R21876 GND.n7481 GND.n7480 585
R21877 GND.n7479 GND.n7478 585
R21878 GND.n7477 GND.n7476 585
R21879 GND.n7475 GND.n7474 585
R21880 GND.n7473 GND.n7472 585
R21881 GND.n7471 GND.n7470 585
R21882 GND.n7469 GND.n7468 585
R21883 GND.n7467 GND.n7466 585
R21884 GND.n7465 GND.n7464 585
R21885 GND.n7463 GND.n7450 585
R21886 GND.n7451 GND.n7450 585
R21887 GND.n7501 GND.n7449 585
R21888 GND.n7501 GND.n7500 585
R21889 GND.n7503 GND.n7502 585
R21890 GND.n7502 GND.n2461 585
R21891 GND.n7504 GND.n2453 585
R21892 GND.n7553 GND.n2453 585
R21893 GND.n7507 GND.n7506 585
R21894 GND.n7506 GND.n7505 585
R21895 GND.n7508 GND.n2445 585
R21896 GND.n7559 GND.n2445 585
R21897 GND.n7510 GND.n7509 585
R21898 GND.n7511 GND.n7510 585
R21899 GND.n7448 GND.n2468 585
R21900 GND.n2468 GND.n2438 585
R21901 GND.n7447 GND.n2436 585
R21902 GND.n7567 GND.n2436 585
R21903 GND.n7446 GND.n7445 585
R21904 GND.n7445 GND.n7444 585
R21905 GND.n7443 GND.n2428 585
R21906 GND.n7573 GND.n2428 585
R21907 GND.n7442 GND.n7441 585
R21908 GND.n7441 GND.n2426 585
R21909 GND.n7440 GND.n2469 585
R21910 GND.n7440 GND.n2420 585
R21911 GND.n7439 GND.n2471 585
R21912 GND.n7439 GND.n7438 585
R21913 GND.n7412 GND.n2470 585
R21914 GND.n2481 GND.n2470 585
R21915 GND.n2491 GND.n2479 585
R21916 GND.n7429 GND.n2479 585
R21917 GND.n7418 GND.n7417 585
R21918 GND.n7419 GND.n7418 585
R21919 GND.n7407 GND.n2489 585
R21920 GND.n2498 GND.n2489 585
R21921 GND.n7406 GND.n7405 585
R21922 GND.n7405 GND.n7404 585
R21923 GND.n7262 GND.n2494 585
R21924 GND.n2527 GND.n2494 585
R21925 GND.n7261 GND.n2506 585
R21926 GND.n7390 GND.n2506 585
R21927 GND.n7268 GND.n7267 585
R21928 GND.n7267 GND.n2518 585
R21929 GND.n7270 GND.n2618 585
R21930 GND.n7288 GND.n2618 585
R21931 GND.n2628 GND.n2626 585
R21932 GND.n2626 GND.n2547 585
R21933 GND.n7276 GND.n7275 585
R21934 GND.n7277 GND.n7276 585
R21935 GND.n7256 GND.n2625 585
R21936 GND.n2625 GND.n2558 585
R21937 GND.n7255 GND.n7254 585
R21938 GND.n7254 GND.n7253 585
R21939 GND.n2631 GND.n2630 585
R21940 GND.n6611 GND.n2631 585
R21941 GND.n7029 GND.n6630 585
R21942 GND.n7201 GND.n6630 585
R21943 GND.n7035 GND.n7034 585
R21944 GND.n7034 GND.n6621 585
R21945 GND.n7037 GND.n6652 585
R21946 GND.n7172 GND.n6652 585
R21947 GND.n6742 GND.n6740 585
R21948 GND.n6740 GND.n6648 585
R21949 GND.n7043 GND.n7042 585
R21950 GND.n7044 GND.n7043 585
R21951 GND.n7024 GND.n6739 585
R21952 GND.n6739 GND.n6663 585
R21953 GND.n7023 GND.n7022 585
R21954 GND.n7022 GND.n6675 585
R21955 GND.n7021 GND.n7020 585
R21956 GND.n7021 GND.n6671 585
R21957 GND.n6745 GND.n6731 585
R21958 GND.n7062 GND.n6731 585
R21959 GND.n7015 GND.n7014 585
R21960 GND.n7014 GND.n7013 585
R21961 GND.n6976 GND.n6748 585
R21962 GND.n6749 GND.n6748 585
R21963 GND.n6975 GND.n6756 585
R21964 GND.n6998 GND.n6756 585
R21965 GND.n6981 GND.n6980 585
R21966 GND.n6982 GND.n6981 585
R21967 GND.n6974 GND.n6763 585
R21968 GND.n6985 GND.n6763 585
R21969 GND.n6973 GND.n6972 585
R21970 GND.n6972 GND.n6971 585
R21971 GND.n6766 GND.n6765 585
R21972 GND.n6767 GND.n6766 585
R21973 GND.n6850 GND.n6775 585
R21974 GND.n6962 GND.n6775 585
R21975 GND.n6852 GND.n6851 585
R21976 GND.n6851 GND.n6773 585
R21977 GND.n6853 GND.n6781 585
R21978 GND.n6955 GND.n6781 585
R21979 GND.n6856 GND.n6854 585
R21980 GND.n6856 GND.n6855 585
R21981 GND.n6858 GND.n6857 585
R21982 GND.n6857 GND.n6785 585
R21983 GND.n6859 GND.n6792 585
R21984 GND.n6912 GND.n6792 585
R21985 GND.n6860 GND.n6799 585
R21986 GND.n6799 GND.n6790 585
R21987 GND.n6862 GND.n6861 585
R21988 GND.n6905 GND.n6862 585
R21989 GND.n6849 GND.n6798 585
R21990 GND.n6803 GND.n6798 585
R21991 GND.n6848 GND.n6847 585
R21992 GND.n6847 GND.n6846 585
R21993 GND.n2892 GND 573.913
R21994 GND.t14 GND.t372 568.212
R21995 GND.t139 GND.t63 568.212
R21996 GND.t137 GND.t45 568.212
R21997 GND.n3111 GND.n2313 544.87
R21998 GND.n2999 GND.t146 509.935
R21999 GND.n7735 GND.n2274 483.204
R22000 GND.n5729 GND.n2274 471.378
R22001 GND.t142 GND 466.226
R22002 GND GND.t294 466.226
R22003 GND.t391 GND 466.226
R22004 GND.t389 GND 458.94
R22005 GND.n8397 GND.n1815 457.69
R22006 GND.n7719 GND.n7718 446.495
R22007 GND.n7719 GND.n7717 446.495
R22008 GND.n7712 GND.n2304 446.495
R22009 GND.n7706 GND.n2304 446.495
R22010 GND.n9460 GND.n9435 446.495
R22011 GND.n9454 GND.n9435 446.495
R22012 GND.n9449 GND.n9440 446.495
R22013 GND.n9443 GND.n9440 446.495
R22014 GND GND.t360 407.947
R22015 GND.t416 GND 407.947
R22016 GND.t372 GND 407.947
R22017 GND.t112 GND.t317 407.947
R22018 GND.t272 GND.t318 407.947
R22019 GND.t110 GND.t315 407.947
R22020 GND.t199 GND.t316 407.947
R22021 GND.t368 GND.t292 407.947
R22022 GND.t369 GND.t296 407.947
R22023 GND.t298 GND.t366 407.947
R22024 GND.t294 GND.t367 407.947
R22025 GND.t269 GND.t332 407.947
R22026 GND.t397 GND.t8 407.947
R22027 GND.t346 GND.t37 407.947
R22028 GND.t347 GND.t344 407.947
R22029 GND.t387 GND.t364 407.947
R22030 GND.t393 GND.t362 407.947
R22031 GND.t363 GND.t381 407.947
R22032 GND.t365 GND.t391 407.947
R22033 GND.n7624 GND.n2361 394
R22034 GND.n7620 GND.n2361 394
R22035 GND.n7620 GND.n2364 394
R22036 GND.n5472 GND.n2364 394
R22037 GND.n5472 GND.n5471 394
R22038 GND.n5494 GND.n5492 394
R22039 GND.n5498 GND.n5493 394
R22040 GND.n5524 GND.n5523 394
R22041 GND.n5521 GND.n5515 394
R22042 GND.n5649 GND.n2358 394
R22043 GND.n5649 GND.n2366 394
R22044 GND.n5645 GND.n2366 394
R22045 GND.n5645 GND.n5644 394
R22046 GND.n5644 GND.n5643 394
R22047 GND.n5479 GND.n5478 394
R22048 GND.n5481 GND.n5479 394
R22049 GND.n5634 GND.n5467 394
R22050 GND.n5637 GND.n5636 394
R22051 GND.n5639 GND.n5464 394
R22052 GND.n7638 GND.n2341 394
R22053 GND.n7634 GND.n2341 394
R22054 GND.n7634 GND.n2344 394
R22055 GND.n2372 GND.n2344 394
R22056 GND.n2373 GND.n2372 394
R22057 GND.n2373 GND.n2369 394
R22058 GND.n7617 GND.n2369 394
R22059 GND.n7617 GND.n2370 394
R22060 GND.n7613 GND.n2370 394
R22061 GND.n7613 GND.n2377 394
R22062 GND.n2391 GND.n2377 394
R22063 GND.n7603 GND.n2391 394
R22064 GND.n7603 GND.n2392 394
R22065 GND.n7599 GND.n2392 394
R22066 GND.n7599 GND.n2395 394
R22067 GND.n5534 GND.n5533 394
R22068 GND.n5549 GND.n5548 394
R22069 GND.n5542 GND.n2338 394
R22070 GND.n5542 GND.n2346 394
R22071 GND.n5538 GND.n2346 394
R22072 GND.n5538 GND.n5537 394
R22073 GND.n5537 GND.n5460 394
R22074 GND.n5652 GND.n5460 394
R22075 GND.n5652 GND.n2367 394
R22076 GND.n5659 GND.n2367 394
R22077 GND.n5659 GND.n2379 394
R22078 GND.n5561 GND.n2379 394
R22079 GND.n5607 GND.n5561 394
R22080 GND.n5607 GND.n2389 394
R22081 GND.n5611 GND.n2389 394
R22082 GND.n5611 GND.n2397 394
R22083 GND.n5559 GND.n2397 394
R22084 GND.n5617 GND.n5556 394
R22085 GND.n5624 GND.n5556 394
R22086 GND.n5616 GND.n5557 394
R22087 GND.n7646 GND.n2325 394
R22088 GND.n7646 GND.n2332 394
R22089 GND.n7642 GND.n2332 394
R22090 GND.n7642 GND.n2334 394
R22091 GND.n2351 GND.n2334 394
R22092 GND.n2351 GND.n2349 394
R22093 GND.n7631 GND.n2349 394
R22094 GND.n7631 GND.n2350 394
R22095 GND.n7627 GND.n2350 394
R22096 GND.n7627 GND.n2355 394
R22097 GND.n5454 GND.n2355 394
R22098 GND.n5454 GND.n5453 394
R22099 GND.n5453 GND.n2382 394
R22100 GND.n7610 GND.n2382 394
R22101 GND.n7610 GND.n2383 394
R22102 GND.n7606 GND.n2383 394
R22103 GND.n7606 GND.n2386 394
R22104 GND.n2400 GND.n2386 394
R22105 GND.n7596 GND.n2400 394
R22106 GND.n7596 GND.n2401 394
R22107 GND.n7592 GND.n2401 394
R22108 GND.n7592 GND.n2404 394
R22109 GND.n7588 GND.n2404 394
R22110 GND.n7682 GND.n2326 394
R22111 GND.n7678 GND.n7677 394
R22112 GND.n7674 GND.n7673 394
R22113 GND.n7670 GND.n7669 394
R22114 GND.n7666 GND.n7665 394
R22115 GND.n7662 GND.n7661 394
R22116 GND.n7658 GND.n7657 394
R22117 GND.n7654 GND.n7653 394
R22118 GND.n7649 GND.n7648 394
R22119 GND.n7648 GND.n2329 394
R22120 GND.n2336 GND.n2329 394
R22121 GND.n2337 GND.n2336 394
R22122 GND.n5504 GND.n2337 394
R22123 GND.n5505 GND.n5504 394
R22124 GND.n5505 GND.n2347 394
R22125 GND.n5512 GND.n2347 394
R22126 GND.n5512 GND.n2357 394
R22127 GND.n5508 GND.n2357 394
R22128 GND.n5508 GND.n5445 394
R22129 GND.n5663 GND.n5445 394
R22130 GND.n5663 GND.n5662 394
R22131 GND.n5662 GND.n2380 394
R22132 GND.n5604 GND.n2380 394
R22133 GND.n5604 GND.n2388 394
R22134 GND.n5600 GND.n2388 394
R22135 GND.n5600 GND.n5599 394
R22136 GND.n5599 GND.n2398 394
R22137 GND.n5595 GND.n2398 394
R22138 GND.n5595 GND.n2405 394
R22139 GND.n2406 GND.n2405 394
R22140 GND.n2407 GND.n2406 394
R22141 GND.n7584 GND.n2410 394
R22142 GND.n5564 GND.n2410 394
R22143 GND.n5568 GND.n5567 394
R22144 GND.n5572 GND.n5571 394
R22145 GND.n5576 GND.n5575 394
R22146 GND.n5580 GND.n5579 394
R22147 GND.n5584 GND.n5583 394
R22148 GND.n5588 GND.n5587 394
R22149 GND.n6088 GND.n6086 394
R22150 GND.n6086 GND.n6085 394
R22151 GND.n6082 GND.n6081 394
R22152 GND.n6079 GND.n5990 394
R22153 GND.n6075 GND.n6073 394
R22154 GND.n6071 GND.n5992 394
R22155 GND.n6067 GND.n6065 394
R22156 GND.n6063 GND.n5994 394
R22157 GND.n6059 GND.n6057 394
R22158 GND.n6055 GND.n5996 394
R22159 GND.n6051 GND.n6049 394
R22160 GND.n6047 GND.n5998 394
R22161 GND.n6043 GND.n6041 394
R22162 GND.n6039 GND.n6000 394
R22163 GND.n6035 GND.n6033 394
R22164 GND.n6031 GND.n6002 394
R22165 GND.n6027 GND.n6025 394
R22166 GND.n6023 GND.n6004 394
R22167 GND.n6019 GND.n6017 394
R22168 GND.n6015 GND.n6006 394
R22169 GND.n6011 GND.n6009 394
R22170 GND.n6092 GND.n2891 394
R22171 GND.n6100 GND.n2891 394
R22172 GND.n6100 GND.n2889 394
R22173 GND.n6104 GND.n2889 394
R22174 GND.n6104 GND.n2883 394
R22175 GND.n6112 GND.n2883 394
R22176 GND.n6112 GND.n2881 394
R22177 GND.n6116 GND.n2881 394
R22178 GND.n6116 GND.n2875 394
R22179 GND.n6124 GND.n2875 394
R22180 GND.n6124 GND.n2873 394
R22181 GND.n6128 GND.n2873 394
R22182 GND.n6128 GND.n2867 394
R22183 GND.n6136 GND.n2867 394
R22184 GND.n6136 GND.n2864 394
R22185 GND.n6179 GND.n2864 394
R22186 GND.n6179 GND.n2865 394
R22187 GND.n6175 GND.n6174 394
R22188 GND.n6172 GND.n6140 394
R22189 GND.n6168 GND.n6167 394
R22190 GND.n6165 GND.n6143 394
R22191 GND.n6161 GND.n6160 394
R22192 GND.n6158 GND.n6146 394
R22193 GND.n6154 GND.n6153 394
R22194 GND.n6151 GND.n6149 394
R22195 GND.n6230 GND.n6229 394
R22196 GND.n6227 GND.n2798 394
R22197 GND.n6223 GND.n6222 394
R22198 GND.n6220 GND.n2805 394
R22199 GND.n6216 GND.n6215 394
R22200 GND.n6213 GND.n2812 394
R22201 GND.n6209 GND.n6208 394
R22202 GND.n6206 GND.n2850 394
R22203 GND.n6202 GND.n6201 394
R22204 GND.n6199 GND.n2853 394
R22205 GND.n6195 GND.n6194 394
R22206 GND.n6192 GND.n2856 394
R22207 GND.n6188 GND.n6187 394
R22208 GND.n6094 GND.n3114 394
R22209 GND.n6098 GND.n3114 394
R22210 GND.n6098 GND.n2887 394
R22211 GND.n6106 GND.n2887 394
R22212 GND.n6106 GND.n2885 394
R22213 GND.n6110 GND.n2885 394
R22214 GND.n6110 GND.n2879 394
R22215 GND.n6118 GND.n2879 394
R22216 GND.n6118 GND.n2877 394
R22217 GND.n6122 GND.n2877 394
R22218 GND.n6122 GND.n2871 394
R22219 GND.n6130 GND.n2871 394
R22220 GND.n6130 GND.n2869 394
R22221 GND.n6134 GND.n2869 394
R22222 GND.n6134 GND.n2861 394
R22223 GND.n6181 GND.n2861 394
R22224 GND.n6181 GND.n2859 394
R22225 GND.n6259 GND.n2770 394
R22226 GND.n6259 GND.n2792 394
R22227 GND.n6255 GND.n6254 394
R22228 GND.n6251 GND.n6250 394
R22229 GND.n6247 GND.n6246 394
R22230 GND.n6243 GND.n6242 394
R22231 GND.n6239 GND.n6238 394
R22232 GND.n6235 GND.n6234 394
R22233 GND.n2795 GND.n2794 394
R22234 GND.n2800 GND.n2799 394
R22235 GND.n2802 GND.n2801 394
R22236 GND.n2807 GND.n2806 394
R22237 GND.n2809 GND.n2808 394
R22238 GND.n2845 GND.n2844 394
R22239 GND.n2841 GND.n2840 394
R22240 GND.n2837 GND.n2836 394
R22241 GND.n2833 GND.n2832 394
R22242 GND.n2829 GND.n2828 394
R22243 GND.n2825 GND.n2824 394
R22244 GND.n2821 GND.n2820 394
R22245 GND.n2817 GND.n2816 394
R22246 GND.n6266 GND.n2768 394
R22247 GND.n6266 GND.n2762 394
R22248 GND.n6274 GND.n2762 394
R22249 GND.n6274 GND.n2760 394
R22250 GND.n6278 GND.n2760 394
R22251 GND.n6278 GND.n2754 394
R22252 GND.n6287 GND.n2754 394
R22253 GND.n6287 GND.n2752 394
R22254 GND.n6291 GND.n2752 394
R22255 GND.n6291 GND.n2747 394
R22256 GND.n6299 GND.n2747 394
R22257 GND.n6299 GND.n2745 394
R22258 GND.n6303 GND.n2745 394
R22259 GND.n6303 GND.n2739 394
R22260 GND.n6312 GND.n2739 394
R22261 GND.n6312 GND.n2736 394
R22262 GND.n6387 GND.n2736 394
R22263 GND.n6383 GND.n2737 394
R22264 GND.n6381 GND.n6380 394
R22265 GND.n6378 GND.n6317 394
R22266 GND.n6374 GND.n6373 394
R22267 GND.n6371 GND.n6320 394
R22268 GND.n6367 GND.n6366 394
R22269 GND.n6364 GND.n6323 394
R22270 GND.n6360 GND.n6359 394
R22271 GND.n6357 GND.n6326 394
R22272 GND.n6347 GND.n6333 394
R22273 GND.n6345 GND.n6344 394
R22274 GND.n6342 GND.n6336 394
R22275 GND.n6420 GND.n2719 394
R22276 GND.n6418 GND.n6417 394
R22277 GND.n6415 GND.n2722 394
R22278 GND.n6411 GND.n6410 394
R22279 GND.n6408 GND.n2725 394
R22280 GND.n6404 GND.n6403 394
R22281 GND.n6401 GND.n2728 394
R22282 GND.n6397 GND.n6396 394
R22283 GND.n6394 GND.n2731 394
R22284 GND.n6268 GND.n2766 394
R22285 GND.n6268 GND.n2764 394
R22286 GND.n6272 GND.n2764 394
R22287 GND.n6272 GND.n2758 394
R22288 GND.n6280 GND.n2758 394
R22289 GND.n6280 GND.n2756 394
R22290 GND.n6284 GND.n2756 394
R22291 GND.n6284 GND.n2751 394
R22292 GND.n6293 GND.n2751 394
R22293 GND.n6293 GND.n2749 394
R22294 GND.n6297 GND.n2749 394
R22295 GND.n6297 GND.n2743 394
R22296 GND.n6305 GND.n2743 394
R22297 GND.n6305 GND.n2741 394
R22298 GND.n6310 GND.n2741 394
R22299 GND.n6310 GND.n2734 394
R22300 GND.n6389 GND.n2734 394
R22301 GND.n3719 GND.n3718 394
R22302 GND.n5975 GND.n3718 394
R22303 GND.n5973 GND.n5972 394
R22304 GND.n5969 GND.n5968 394
R22305 GND.n5965 GND.n5964 394
R22306 GND.n5961 GND.n5960 394
R22307 GND.n5957 GND.n5956 394
R22308 GND.n5953 GND.n5952 394
R22309 GND.n5949 GND.n5948 394
R22310 GND.n5945 GND.n5944 394
R22311 GND.n5941 GND.n5940 394
R22312 GND.n5937 GND.n5936 394
R22313 GND.n5933 GND.n5932 394
R22314 GND.n5929 GND.n5928 394
R22315 GND.n5925 GND.n5924 394
R22316 GND.n5921 GND.n5920 394
R22317 GND.n5917 GND.n5916 394
R22318 GND.n5913 GND.n5912 394
R22319 GND.n5909 GND.n5908 394
R22320 GND.n5905 GND.n5904 394
R22321 GND.n5901 GND.n5900 394
R22322 GND.n3737 GND.n3720 394
R22323 GND.n3737 GND.n3735 394
R22324 GND.n5886 GND.n3735 394
R22325 GND.n5886 GND.n3736 394
R22326 GND.n5882 GND.n3736 394
R22327 GND.n5882 GND.n3741 394
R22328 GND.n3755 GND.n3741 394
R22329 GND.n5872 GND.n3755 394
R22330 GND.n5872 GND.n3756 394
R22331 GND.n5868 GND.n3756 394
R22332 GND.n5868 GND.n3759 394
R22333 GND.n3773 GND.n3759 394
R22334 GND.n5858 GND.n3773 394
R22335 GND.n5858 GND.n3774 394
R22336 GND.n5854 GND.n3774 394
R22337 GND.n5854 GND.n3777 394
R22338 GND.n3811 GND.n3777 394
R22339 GND.n5844 GND.n3812 394
R22340 GND.n5840 GND.n5839 394
R22341 GND.n5836 GND.n5835 394
R22342 GND.n5832 GND.n5831 394
R22343 GND.n5828 GND.n5827 394
R22344 GND.n5824 GND.n5823 394
R22345 GND.n5820 GND.n5819 394
R22346 GND.n5816 GND.n5815 394
R22347 GND.n4018 GND.n4017 394
R22348 GND.n4024 GND.n4023 394
R22349 GND.n4030 GND.n4029 394
R22350 GND.n4036 GND.n4035 394
R22351 GND.n4042 GND.n4041 394
R22352 GND.n4014 GND.n4013 394
R22353 GND.n4010 GND.n4009 394
R22354 GND.n4006 GND.n4005 394
R22355 GND.n4002 GND.n4001 394
R22356 GND.n3998 GND.n3997 394
R22357 GND.n3994 GND.n3993 394
R22358 GND.n3990 GND.n3989 394
R22359 GND.n3986 GND.n3985 394
R22360 GND.n5896 GND.n3723 394
R22361 GND.n3954 GND.n3723 394
R22362 GND.n3954 GND.n3733 394
R22363 GND.n3958 GND.n3733 394
R22364 GND.n3958 GND.n3743 394
R22365 GND.n3962 GND.n3743 394
R22366 GND.n3963 GND.n3962 394
R22367 GND.n3963 GND.n3753 394
R22368 GND.n3967 GND.n3753 394
R22369 GND.n3967 GND.n3761 394
R22370 GND.n3971 GND.n3761 394
R22371 GND.n3972 GND.n3971 394
R22372 GND.n3972 GND.n3771 394
R22373 GND.n3976 GND.n3771 394
R22374 GND.n3976 GND.n3779 394
R22375 GND.n3980 GND.n3779 394
R22376 GND.n3981 GND.n3980 394
R22377 GND.n5195 GND.n5193 394
R22378 GND.n5199 GND.n5193 394
R22379 GND.n5203 GND.n5201 394
R22380 GND.n5207 GND.n5191 394
R22381 GND.n5211 GND.n5209 394
R22382 GND.n5215 GND.n5189 394
R22383 GND.n5219 GND.n5217 394
R22384 GND.n5223 GND.n5187 394
R22385 GND.n5227 GND.n5225 394
R22386 GND.n5231 GND.n5185 394
R22387 GND.n5235 GND.n5233 394
R22388 GND.n5239 GND.n5183 394
R22389 GND.n5243 GND.n5241 394
R22390 GND.n5247 GND.n5181 394
R22391 GND.n5251 GND.n5249 394
R22392 GND.n5255 GND.n5179 394
R22393 GND.n5259 GND.n5257 394
R22394 GND.n5263 GND.n5177 394
R22395 GND.n5267 GND.n5265 394
R22396 GND.n5271 GND.n5175 394
R22397 GND.n5274 GND.n5273 394
R22398 GND.n5893 GND.n3727 394
R22399 GND.n5889 GND.n3727 394
R22400 GND.n5889 GND.n3730 394
R22401 GND.n3746 GND.n3730 394
R22402 GND.n5879 GND.n3746 394
R22403 GND.n5879 GND.n3747 394
R22404 GND.n5875 GND.n3747 394
R22405 GND.n5875 GND.n3750 394
R22406 GND.n3764 GND.n3750 394
R22407 GND.n5865 GND.n3764 394
R22408 GND.n5865 GND.n3765 394
R22409 GND.n5861 GND.n3765 394
R22410 GND.n5861 GND.n3768 394
R22411 GND.n3782 GND.n3768 394
R22412 GND.n5851 GND.n3782 394
R22413 GND.n5851 GND.n3783 394
R22414 GND.n5847 GND.n3783 394
R22415 GND.n5057 GND.n3786 394
R22416 GND.n5061 GND.n5059 394
R22417 GND.n5065 GND.n5054 394
R22418 GND.n5069 GND.n5067 394
R22419 GND.n5073 GND.n5052 394
R22420 GND.n5077 GND.n5075 394
R22421 GND.n5081 GND.n5050 394
R22422 GND.n5085 GND.n5083 394
R22423 GND.n5135 GND.n5048 394
R22424 GND.n5139 GND.n5137 394
R22425 GND.n5147 GND.n5044 394
R22426 GND.n5151 GND.n5149 394
R22427 GND.n5160 GND.n5040 394
R22428 GND.n5337 GND.n5162 394
R22429 GND.n5335 GND.n5334 394
R22430 GND.n5332 GND.n5164 394
R22431 GND.n5328 GND.n5327 394
R22432 GND.n5325 GND.n5167 394
R22433 GND.n5321 GND.n5320 394
R22434 GND.n5318 GND.n5170 394
R22435 GND.n5314 GND.n5313 394
R22436 GND.n5280 GND.n3724 394
R22437 GND.n5280 GND.n3732 394
R22438 GND.n5284 GND.n3732 394
R22439 GND.n5285 GND.n5284 394
R22440 GND.n5285 GND.n3744 394
R22441 GND.n5289 GND.n3744 394
R22442 GND.n5289 GND.n3752 394
R22443 GND.n5293 GND.n3752 394
R22444 GND.n5294 GND.n5293 394
R22445 GND.n5294 GND.n3762 394
R22446 GND.n5298 GND.n3762 394
R22447 GND.n5298 GND.n3770 394
R22448 GND.n5302 GND.n3770 394
R22449 GND.n5303 GND.n5302 394
R22450 GND.n5303 GND.n3780 394
R22451 GND.n5307 GND.n3780 394
R22452 GND.n5307 GND.n3788 394
R22453 GND.n3839 GND.n3838 394
R22454 GND.n5802 GND.n3838 394
R22455 GND.n5800 GND.n5799 394
R22456 GND.n5796 GND.n5795 394
R22457 GND.n5792 GND.n5791 394
R22458 GND.n5788 GND.n5787 394
R22459 GND.n5784 GND.n5783 394
R22460 GND.n5811 GND.n3816 394
R22461 GND.n4016 GND.n3817 394
R22462 GND.n4022 GND.n4021 394
R22463 GND.n4028 GND.n4027 394
R22464 GND.n4034 GND.n4033 394
R22465 GND.n4040 GND.n4039 394
R22466 GND.n4047 GND.n4046 394
R22467 GND.n4051 GND.n4050 394
R22468 GND.n4055 GND.n4054 394
R22469 GND.n4059 GND.n4058 394
R22470 GND.n4063 GND.n4062 394
R22471 GND.n4067 GND.n4066 394
R22472 GND.n4071 GND.n4070 394
R22473 GND.n4075 GND.n4074 394
R22474 GND.n5779 GND.n3840 394
R22475 GND.n5779 GND.n3842 394
R22476 GND.n3856 GND.n3842 394
R22477 GND.n5769 GND.n3856 394
R22478 GND.n5769 GND.n3857 394
R22479 GND.n5765 GND.n3857 394
R22480 GND.n5765 GND.n3860 394
R22481 GND.n3874 GND.n3860 394
R22482 GND.n5755 GND.n3874 394
R22483 GND.n5755 GND.n3875 394
R22484 GND.n5751 GND.n3875 394
R22485 GND.n5751 GND.n3878 394
R22486 GND.n3892 GND.n3878 394
R22487 GND.n5741 GND.n3892 394
R22488 GND.n5741 GND.n3893 394
R22489 GND.n5737 GND.n3893 394
R22490 GND.n5737 GND.n3896 394
R22491 GND.n4981 GND.n3927 394
R22492 GND.n4977 GND.n4976 394
R22493 GND.n4973 GND.n4972 394
R22494 GND.n4969 GND.n4968 394
R22495 GND.n4965 GND.n4964 394
R22496 GND.n4961 GND.n4960 394
R22497 GND.n4957 GND.n4956 394
R22498 GND.n4953 GND.n4952 394
R22499 GND.n4949 GND.n4948 394
R22500 GND.n3940 GND.n3939 394
R22501 GND.n3944 GND.n3943 394
R22502 GND.n3948 GND.n3947 394
R22503 GND.n4147 GND.n4146 394
R22504 GND.n4144 GND.n4143 394
R22505 GND.n4140 GND.n4139 394
R22506 GND.n4136 GND.n4135 394
R22507 GND.n4132 GND.n4131 394
R22508 GND.n4128 GND.n4127 394
R22509 GND.n4124 GND.n4123 394
R22510 GND.n4120 GND.n4119 394
R22511 GND.n4116 GND.n4115 394
R22512 GND.n4080 GND.n3844 394
R22513 GND.n4084 GND.n3844 394
R22514 GND.n4085 GND.n4084 394
R22515 GND.n4085 GND.n3854 394
R22516 GND.n4089 GND.n3854 394
R22517 GND.n4089 GND.n3862 394
R22518 GND.n4093 GND.n3862 394
R22519 GND.n4094 GND.n4093 394
R22520 GND.n4094 GND.n3872 394
R22521 GND.n4098 GND.n3872 394
R22522 GND.n4098 GND.n3880 394
R22523 GND.n4102 GND.n3880 394
R22524 GND.n4103 GND.n4102 394
R22525 GND.n4103 GND.n3890 394
R22526 GND.n4107 GND.n3890 394
R22527 GND.n4107 GND.n3898 394
R22528 GND.n4111 GND.n3898 394
R22529 GND.n5099 GND.n5095 394
R22530 GND.n5103 GND.n5095 394
R22531 GND.n5107 GND.n5105 394
R22532 GND.n5111 GND.n5093 394
R22533 GND.n5115 GND.n5113 394
R22534 GND.n5119 GND.n5091 394
R22535 GND.n5123 GND.n5121 394
R22536 GND.n5127 GND.n5089 394
R22537 GND.n5131 GND.n5129 394
R22538 GND.n5141 GND.n5046 394
R22539 GND.n5145 GND.n5143 394
R22540 GND.n5153 GND.n5042 394
R22541 GND.n5158 GND.n5155 394
R22542 GND.n5156 GND.n5039 394
R22543 GND.n5342 GND.n5035 394
R22544 GND.n5346 GND.n5344 394
R22545 GND.n5350 GND.n5033 394
R22546 GND.n5354 GND.n5352 394
R22547 GND.n5358 GND.n5031 394
R22548 GND.n5362 GND.n5360 394
R22549 GND.n5366 GND.n5029 394
R22550 GND.n5776 GND.n3847 394
R22551 GND.n5776 GND.n3848 394
R22552 GND.n5772 GND.n3848 394
R22553 GND.n5772 GND.n3851 394
R22554 GND.n3865 GND.n3851 394
R22555 GND.n5762 GND.n3865 394
R22556 GND.n5762 GND.n3866 394
R22557 GND.n5758 GND.n3866 394
R22558 GND.n5758 GND.n3869 394
R22559 GND.n3883 GND.n3869 394
R22560 GND.n5748 GND.n3883 394
R22561 GND.n5748 GND.n3884 394
R22562 GND.n5744 GND.n3884 394
R22563 GND.n5744 GND.n3887 394
R22564 GND.n3901 GND.n3887 394
R22565 GND.n5734 GND.n3901 394
R22566 GND.n5734 GND.n3902 394
R22567 GND.n5730 GND.n3905 394
R22568 GND.n5727 GND.n5003 394
R22569 GND.n5723 GND.n5722 394
R22570 GND.n5719 GND.n5718 394
R22571 GND.n5715 GND.n5714 394
R22572 GND.n5711 GND.n5710 394
R22573 GND.n5707 GND.n5706 394
R22574 GND.n5703 GND.n5702 394
R22575 GND.n5699 GND.n5698 394
R22576 GND.n5695 GND.n5694 394
R22577 GND.n5016 GND.n5015 394
R22578 GND.n5020 GND.n5019 394
R22579 GND.n5024 GND.n5023 394
R22580 GND.n5433 GND.n5432 394
R22581 GND.n5430 GND.n5429 394
R22582 GND.n5426 GND.n5425 394
R22583 GND.n5422 GND.n5421 394
R22584 GND.n5418 GND.n5417 394
R22585 GND.n5414 GND.n5413 394
R22586 GND.n5410 GND.n5409 394
R22587 GND.n5406 GND.n5405 394
R22588 GND.n5369 GND.n3845 394
R22589 GND.n5373 GND.n3845 394
R22590 GND.n5373 GND.n3853 394
R22591 GND.n5377 GND.n3853 394
R22592 GND.n5378 GND.n5377 394
R22593 GND.n5378 GND.n3863 394
R22594 GND.n5382 GND.n3863 394
R22595 GND.n5382 GND.n3871 394
R22596 GND.n5386 GND.n3871 394
R22597 GND.n5387 GND.n5386 394
R22598 GND.n5387 GND.n3881 394
R22599 GND.n5391 GND.n3881 394
R22600 GND.n5391 GND.n3889 394
R22601 GND.n5395 GND.n3889 394
R22602 GND.n5396 GND.n5395 394
R22603 GND.n5396 GND.n3899 394
R22604 GND.n5401 GND.n3899 394
R22605 GND.n2231 GND.n2161 394
R22606 GND.n7968 GND.n2161 394
R22607 GND.n7968 GND.n2162 394
R22608 GND.n7964 GND.n2162 394
R22609 GND.n7964 GND.n2165 394
R22610 GND.n2236 GND.n2235 394
R22611 GND.n2239 GND.n2238 394
R22612 GND.n2247 GND.n2246 394
R22613 GND.n2249 GND.n2226 394
R22614 GND.n2227 GND.n2207 394
R22615 GND.n2207 GND.n2159 394
R22616 GND.n7857 GND.n2159 394
R22617 GND.n7857 GND.n2167 394
R22618 GND.n7932 GND.n2167 394
R22619 GND.n2182 GND.n2181 394
R22620 GND.n7948 GND.n2181 394
R22621 GND.n7943 GND.n7942 394
R22622 GND.n7939 GND.n7938 394
R22623 GND.n7935 GND.n2179 394
R22624 GND.n7838 GND.n2258 394
R22625 GND.n7838 GND.n2259 394
R22626 GND.n2259 GND.n2212 394
R22627 GND.n7875 GND.n2212 394
R22628 GND.n7875 GND.n2209 394
R22629 GND.n7880 GND.n2209 394
R22630 GND.n7880 GND.n2210 394
R22631 GND.n2210 GND.n2169 394
R22632 GND.n7961 GND.n2169 394
R22633 GND.n7961 GND.n2170 394
R22634 GND.n7957 GND.n2170 394
R22635 GND.n7957 GND.n2173 394
R22636 GND.n7906 GND.n2173 394
R22637 GND.n7909 GND.n7906 394
R22638 GND.n7909 GND.n2143 394
R22639 GND.n7831 GND.n7830 394
R22640 GND.n7828 GND.n7820 394
R22641 GND.n7840 GND.n2256 394
R22642 GND.n7841 GND.n7840 394
R22643 GND.n7841 GND.n2221 394
R22644 GND.n2221 GND.n2214 394
R22645 GND.n7846 GND.n2214 394
R22646 GND.n7846 GND.n2208 394
R22647 GND.n2254 GND.n2208 394
R22648 GND.n7854 GND.n2254 394
R22649 GND.n7854 GND.n2168 394
R22650 GND.n7929 GND.n2168 394
R22651 GND.n7929 GND.n2175 394
R22652 GND.n7925 GND.n2175 394
R22653 GND.n7925 GND.n2189 394
R22654 GND.n2200 GND.n2189 394
R22655 GND.n2200 GND.n2194 394
R22656 GND.n2142 GND.n2141 394
R22657 GND.n2145 GND.n2141 394
R22658 GND.n2195 GND.n2140 394
R22659 GND.n7809 GND.n2267 394
R22660 GND.n7809 GND.n2264 394
R22661 GND.n7816 GND.n2264 394
R22662 GND.n7816 GND.n2265 394
R22663 GND.n7812 GND.n2265 394
R22664 GND.n7812 GND.n2218 394
R22665 GND.n7868 GND.n2218 394
R22666 GND.n7868 GND.n2216 394
R22667 GND.n7872 GND.n2216 394
R22668 GND.n7872 GND.n2155 394
R22669 GND.n7971 GND.n2155 394
R22670 GND.n7971 GND.n2157 394
R22671 GND.n7915 GND.n2157 394
R22672 GND.n7916 GND.n7915 394
R22673 GND.n7917 GND.n7916 394
R22674 GND.n7917 GND.n2192 394
R22675 GND.n7922 GND.n2192 394
R22676 GND.n7922 GND.n7912 394
R22677 GND.n7912 GND.n2136 394
R22678 GND.n7988 GND.n2136 394
R22679 GND.n7988 GND.n2134 394
R22680 GND.n7992 GND.n2134 394
R22681 GND.n7992 GND.n2129 394
R22682 GND.n7788 GND.n7757 394
R22683 GND.n7784 GND.n7783 394
R22684 GND.n7780 GND.n7779 394
R22685 GND.n7776 GND.n7775 394
R22686 GND.n7772 GND.n7771 394
R22687 GND.n7768 GND.n7767 394
R22688 GND.n7764 GND.n7763 394
R22689 GND.n7760 GND.n7759 394
R22690 GND.n7791 GND.n2268 394
R22691 GND.n7806 GND.n2268 394
R22692 GND.n7806 GND.n2261 394
R22693 GND.n7802 GND.n2261 394
R22694 GND.n7802 GND.n7801 394
R22695 GND.n7801 GND.n7800 394
R22696 GND.n7800 GND.n2220 394
R22697 GND.n7795 GND.n2220 394
R22698 GND.n7795 GND.n2206 394
R22699 GND.n7884 GND.n2206 394
R22700 GND.n7884 GND.n2158 394
R22701 GND.n2252 GND.n2158 394
R22702 GND.n2252 GND.n2202 394
R22703 GND.n7893 GND.n2202 394
R22704 GND.n7894 GND.n7893 394
R22705 GND.n7895 GND.n7894 394
R22706 GND.n7895 GND.n2190 394
R22707 GND.n2193 GND.n2190 394
R22708 GND.n7904 GND.n2193 394
R22709 GND.n7904 GND.n2138 394
R22710 GND.n7900 GND.n2138 394
R22711 GND.n7900 GND.n2132 394
R22712 GND.n7995 GND.n2132 394
R22713 GND.n2128 GND.n2127 394
R22714 GND.n8022 GND.n2127 394
R22715 GND.n8020 GND.n8019 394
R22716 GND.n8016 GND.n8015 394
R22717 GND.n8012 GND.n8011 394
R22718 GND.n8008 GND.n8007 394
R22719 GND.n8004 GND.n8003 394
R22720 GND.n8000 GND.n7999 394
R22721 GND.n9748 GND.n77 394
R22722 GND.n9748 GND.n78 394
R22723 GND.n9744 GND.n78 394
R22724 GND.n9744 GND.n9743 394
R22725 GND.n9743 GND.n81 394
R22726 GND.n143 GND.n139 394
R22727 GND.n147 GND.n140 394
R22728 GND.n9598 GND.n9597 394
R22729 GND.n9595 GND.n150 394
R22730 GND.n9590 GND.n75 394
R22731 GND.n155 GND.n75 394
R22732 GND.n155 GND.n152 394
R22733 GND.n152 GND.n83 394
R22734 GND.n9711 GND.n83 394
R22735 GND.n98 GND.n97 394
R22736 GND.n9727 GND.n97 394
R22737 GND.n9722 GND.n9721 394
R22738 GND.n9718 GND.n9717 394
R22739 GND.n9714 GND.n95 394
R22740 GND.n9559 GND.n172 394
R22741 GND.n9559 GND.n165 394
R22742 GND.n9580 GND.n165 394
R22743 GND.n9580 GND.n162 394
R22744 GND.n9587 GND.n162 394
R22745 GND.n9587 GND.n163 394
R22746 GND.n9583 GND.n163 394
R22747 GND.n9583 GND.n85 394
R22748 GND.n9740 GND.n85 394
R22749 GND.n9740 GND.n86 394
R22750 GND.n9736 GND.n86 394
R22751 GND.n9736 GND.n89 394
R22752 GND.n124 GND.n89 394
R22753 GND.n124 GND.n122 394
R22754 GND.n9694 GND.n122 394
R22755 GND.n9553 GND.n9552 394
R22756 GND.n9550 GND.n9543 394
R22757 GND.n9561 GND.n170 394
R22758 GND.n9561 GND.n167 394
R22759 GND.n9578 GND.n167 394
R22760 GND.n9578 GND.n168 394
R22761 GND.n168 GND.n161 394
R22762 GND.n9573 GND.n161 394
R22763 GND.n9573 GND.n9572 394
R22764 GND.n9572 GND.n9566 394
R22765 GND.n9566 GND.n84 394
R22766 GND.n9708 GND.n84 394
R22767 GND.n9708 GND.n91 394
R22768 GND.n9704 GND.n91 394
R22769 GND.n9704 GND.n106 394
R22770 GND.n9611 GND.n106 394
R22771 GND.n9611 GND.n120 394
R22772 GND.n9690 GND.n128 394
R22773 GND.n9608 GND.n128 394
R22774 GND.n9615 GND.n130 394
R22775 GND.n9510 GND.n186 394
R22776 GND.n9510 GND.n177 394
R22777 GND.n9539 GND.n177 394
R22778 GND.n9539 GND.n178 394
R22779 GND.n9535 GND.n178 394
R22780 GND.n9535 GND.n9534 394
R22781 GND.n9534 GND.n181 394
R22782 GND.n9525 GND.n181 394
R22783 GND.n9525 GND.n73 394
R22784 GND.n9751 GND.n73 394
R22785 GND.n9751 GND.n67 394
R22786 GND.n9758 GND.n67 394
R22787 GND.n9758 GND.n68 394
R22788 GND.n112 GND.n68 394
R22789 GND.n113 GND.n112 394
R22790 GND.n113 GND.n109 394
R22791 GND.n9701 GND.n109 394
R22792 GND.n9701 GND.n110 394
R22793 GND.n9697 GND.n110 394
R22794 GND.n9697 GND.n117 394
R22795 GND.n9686 GND.n117 394
R22796 GND.n9686 GND.n9618 394
R22797 GND.n9682 GND.n9618 394
R22798 GND.n9506 GND.n188 394
R22799 GND.n9503 GND.n9472 394
R22800 GND.n9499 GND.n9498 394
R22801 GND.n9495 GND.n9494 394
R22802 GND.n9491 GND.n9490 394
R22803 GND.n9487 GND.n9486 394
R22804 GND.n9483 GND.n9482 394
R22805 GND.n9479 GND.n9478 394
R22806 GND.n9474 GND.n185 394
R22807 GND.n9513 GND.n185 394
R22808 GND.n9513 GND.n174 394
R22809 GND.n9516 GND.n174 394
R22810 GND.n9516 GND.n182 394
R22811 GND.n9531 GND.n182 394
R22812 GND.n9531 GND.n183 394
R22813 GND.n9527 GND.n183 394
R22814 GND.n9527 GND.n9521 394
R22815 GND.n9521 GND.n74 394
R22816 GND.n74 GND.n63 394
R22817 GND.n9760 GND.n63 394
R22818 GND.n9760 GND.n64 394
R22819 GND.n9633 GND.n64 394
R22820 GND.n9634 GND.n9633 394
R22821 GND.n9635 GND.n9634 394
R22822 GND.n9635 GND.n107 394
R22823 GND.n9639 GND.n107 394
R22824 GND.n9639 GND.n119 394
R22825 GND.n9642 GND.n119 394
R22826 GND.n9642 GND.n9616 394
R22827 GND.n9645 GND.n9616 394
R22828 GND.n9645 GND.n9621 394
R22829 GND.n9678 GND.n9629 394
R22830 GND.n9674 GND.n9629 394
R22831 GND.n9672 GND.n9671 394
R22832 GND.n9668 GND.n9667 394
R22833 GND.n9664 GND.n9663 394
R22834 GND.n9660 GND.n9659 394
R22835 GND.n9656 GND.n9655 394
R22836 GND.n9652 GND.n9651 394
R22837 GND.n1651 GND.n1094 394
R22838 GND.n1647 GND.n1094 394
R22839 GND.n1647 GND.n1097 394
R22840 GND.n1639 GND.n1097 394
R22841 GND.n1639 GND.n1109 394
R22842 GND.n1635 GND.n1109 394
R22843 GND.n1635 GND.n1111 394
R22844 GND.n1627 GND.n1111 394
R22845 GND.n1627 GND.n1121 394
R22846 GND.n1623 GND.n1121 394
R22847 GND.n1623 GND.n1123 394
R22848 GND.n1615 GND.n1123 394
R22849 GND.n1615 GND.n1133 394
R22850 GND.n1611 GND.n1133 394
R22851 GND.n1611 GND.n1135 394
R22852 GND.n1603 GND.n1135 394
R22853 GND.n1603 GND.n1145 394
R22854 GND.n1599 GND.n1145 394
R22855 GND.n1599 GND.n1147 394
R22856 GND.n1591 GND.n1147 394
R22857 GND.n1591 GND.n1218 394
R22858 GND.n1587 GND.n1218 394
R22859 GND.n1587 GND.n1220 394
R22860 GND.n1579 GND.n1220 394
R22861 GND.n1579 GND.n1232 394
R22862 GND.n1575 GND.n1232 394
R22863 GND.n1575 GND.n1234 394
R22864 GND.n1567 GND.n1234 394
R22865 GND.n1567 GND.n1247 394
R22866 GND.n1563 GND.n1247 394
R22867 GND.n1563 GND.n1249 394
R22868 GND.n1555 GND.n1249 394
R22869 GND.n1555 GND.n1262 394
R22870 GND.n1551 GND.n1262 394
R22871 GND.n1551 GND.n1264 394
R22872 GND.n1543 GND.n1264 394
R22873 GND.n1543 GND.n1274 394
R22874 GND.n1539 GND.n1274 394
R22875 GND.n1539 GND.n1276 394
R22876 GND.n1531 GND.n1276 394
R22877 GND.n1531 GND.n1286 394
R22878 GND.n1527 GND.n1286 394
R22879 GND.n1154 GND.n1153 394
R22880 GND.n1158 GND.n1157 394
R22881 GND.n1162 GND.n1161 394
R22882 GND.n1166 GND.n1165 394
R22883 GND.n1170 GND.n1169 394
R22884 GND.n1174 GND.n1173 394
R22885 GND.n1178 GND.n1177 394
R22886 GND.n1182 GND.n1181 394
R22887 GND.n1187 GND.n1089 394
R22888 GND.n1187 GND.n1098 394
R22889 GND.n1190 GND.n1098 394
R22890 GND.n1190 GND.n1106 394
R22891 GND.n1193 GND.n1106 394
R22892 GND.n1193 GND.n1112 394
R22893 GND.n1196 GND.n1112 394
R22894 GND.n1196 GND.n1118 394
R22895 GND.n1199 GND.n1118 394
R22896 GND.n1199 GND.n1124 394
R22897 GND.n1202 GND.n1124 394
R22898 GND.n1202 GND.n1130 394
R22899 GND.n1205 GND.n1130 394
R22900 GND.n1205 GND.n1136 394
R22901 GND.n1208 GND.n1136 394
R22902 GND.n1208 GND.n1142 394
R22903 GND.n1211 GND.n1142 394
R22904 GND.n1211 GND.n1148 394
R22905 GND.n1594 GND.n1148 394
R22906 GND.n1594 GND.n1593 394
R22907 GND.n1593 GND.n1215 394
R22908 GND.n1221 GND.n1215 394
R22909 GND.n1582 GND.n1221 394
R22910 GND.n1582 GND.n1581 394
R22911 GND.n1581 GND.n1228 394
R22912 GND.n1235 GND.n1228 394
R22913 GND.n1570 GND.n1235 394
R22914 GND.n1570 GND.n1569 394
R22915 GND.n1569 GND.n1242 394
R22916 GND.n1250 GND.n1242 394
R22917 GND.n1293 GND.n1250 394
R22918 GND.n1293 GND.n1259 394
R22919 GND.n1296 GND.n1259 394
R22920 GND.n1296 GND.n1265 394
R22921 GND.n1299 GND.n1265 394
R22922 GND.n1299 GND.n1271 394
R22923 GND.n1302 GND.n1271 394
R22924 GND.n1302 GND.n1277 394
R22925 GND.n1305 GND.n1277 394
R22926 GND.n1305 GND.n1283 394
R22927 GND.n1289 GND.n1283 394
R22928 GND.n1351 GND.n1289 394
R22929 GND.n1320 GND.n1319 394
R22930 GND.n1322 GND.n1320 394
R22931 GND.n1326 GND.n1315 394
R22932 GND.n1330 GND.n1328 394
R22933 GND.n1334 GND.n1313 394
R22934 GND.n1338 GND.n1336 394
R22935 GND.n1342 GND.n1311 394
R22936 GND.n1345 GND.n1344 394
R22937 GND.n1347 GND.n1290 394
R22938 GND.n1101 GND.n1092 394
R22939 GND.n1645 GND.n1101 394
R22940 GND.n1645 GND.n1102 394
R22941 GND.n1641 GND.n1102 394
R22942 GND.n1641 GND.n1105 394
R22943 GND.n1633 GND.n1105 394
R22944 GND.n1633 GND.n1115 394
R22945 GND.n1629 GND.n1115 394
R22946 GND.n1629 GND.n1117 394
R22947 GND.n1621 GND.n1117 394
R22948 GND.n1621 GND.n1127 394
R22949 GND.n1617 GND.n1127 394
R22950 GND.n1617 GND.n1129 394
R22951 GND.n1609 GND.n1129 394
R22952 GND.n1609 GND.n1139 394
R22953 GND.n1605 GND.n1139 394
R22954 GND.n1605 GND.n1141 394
R22955 GND.n1597 GND.n1141 394
R22956 GND.n1597 GND.n1151 394
R22957 GND.n1217 GND.n1151 394
R22958 GND.n1224 GND.n1217 394
R22959 GND.n1585 GND.n1224 394
R22960 GND.n1585 GND.n1225 394
R22961 GND.n1231 GND.n1225 394
R22962 GND.n1238 GND.n1231 394
R22963 GND.n1573 GND.n1238 394
R22964 GND.n1573 GND.n1239 394
R22965 GND.n1246 GND.n1239 394
R22966 GND.n1253 GND.n1246 394
R22967 GND.n1561 GND.n1253 394
R22968 GND.n1561 GND.n1254 394
R22969 GND.n1557 GND.n1254 394
R22970 GND.n1557 GND.n1258 394
R22971 GND.n1549 GND.n1258 394
R22972 GND.n1549 GND.n1268 394
R22973 GND.n1545 GND.n1268 394
R22974 GND.n1545 GND.n1270 394
R22975 GND.n1537 GND.n1270 394
R22976 GND.n1537 GND.n1280 394
R22977 GND.n1533 GND.n1280 394
R22978 GND.n1533 GND.n1282 394
R22979 GND.n1525 GND.n1282 394
R22980 GND.n1374 GND.n1373 394
R22981 GND.n1378 GND.n1377 394
R22982 GND.n1382 GND.n1381 394
R22983 GND.n1386 GND.n1385 394
R22984 GND.n1390 GND.n1389 394
R22985 GND.n1394 GND.n1393 394
R22986 GND.n1398 GND.n1397 394
R22987 GND.n1402 GND.n1401 394
R22988 GND.n1407 GND.n1090 394
R22989 GND.n1407 GND.n1099 394
R22990 GND.n1410 GND.n1099 394
R22991 GND.n1410 GND.n1107 394
R22992 GND.n1413 GND.n1107 394
R22993 GND.n1413 GND.n1113 394
R22994 GND.n1416 GND.n1113 394
R22995 GND.n1416 GND.n1119 394
R22996 GND.n1419 GND.n1119 394
R22997 GND.n1419 GND.n1125 394
R22998 GND.n1422 GND.n1125 394
R22999 GND.n1422 GND.n1131 394
R23000 GND.n1425 GND.n1131 394
R23001 GND.n1425 GND.n1137 394
R23002 GND.n1428 GND.n1137 394
R23003 GND.n1428 GND.n1143 394
R23004 GND.n1431 GND.n1143 394
R23005 GND.n1431 GND.n1149 394
R23006 GND.n1436 GND.n1149 394
R23007 GND.n1436 GND.n1216 394
R23008 GND.n1449 GND.n1216 394
R23009 GND.n1449 GND.n1222 394
R23010 GND.n1446 GND.n1222 394
R23011 GND.n1446 GND.n1229 394
R23012 GND.n1441 GND.n1229 394
R23013 GND.n1441 GND.n1236 394
R23014 GND.n1464 GND.n1236 394
R23015 GND.n1464 GND.n1244 394
R23016 GND.n1467 GND.n1244 394
R23017 GND.n1467 GND.n1251 394
R23018 GND.n1470 GND.n1251 394
R23019 GND.n1470 GND.n1260 394
R23020 GND.n1473 GND.n1260 394
R23021 GND.n1473 GND.n1266 394
R23022 GND.n1476 GND.n1266 394
R23023 GND.n1476 GND.n1272 394
R23024 GND.n1479 GND.n1272 394
R23025 GND.n1479 GND.n1278 394
R23026 GND.n1482 GND.n1278 394
R23027 GND.n1482 GND.n1284 394
R23028 GND.n1485 GND.n1284 394
R23029 GND.n1485 GND.n1352 394
R23030 GND.n1521 GND.n1519 394
R23031 GND.n1517 GND.n1355 394
R23032 GND.n1513 GND.n1511 394
R23033 GND.n1509 GND.n1357 394
R23034 GND.n1505 GND.n1503 394
R23035 GND.n1501 GND.n1359 394
R23036 GND.n1497 GND.n1495 394
R23037 GND.n1493 GND.n1361 394
R23038 GND.n8596 GND.n1794 394
R23039 GND.n8596 GND.n1792 394
R23040 GND.n8600 GND.n1792 394
R23041 GND.n8600 GND.n1782 394
R23042 GND.n8608 GND.n1782 394
R23043 GND.n8608 GND.n1780 394
R23044 GND.n8612 GND.n1780 394
R23045 GND.n8612 GND.n1770 394
R23046 GND.n8620 GND.n1770 394
R23047 GND.n8620 GND.n1768 394
R23048 GND.n8624 GND.n1768 394
R23049 GND.n8624 GND.n1757 394
R23050 GND.n8634 GND.n1757 394
R23051 GND.n8634 GND.n1755 394
R23052 GND.n8638 GND.n1755 394
R23053 GND.n8638 GND.n1744 394
R23054 GND.n8648 GND.n1744 394
R23055 GND.n8648 GND.n1742 394
R23056 GND.n8652 GND.n1742 394
R23057 GND.n8652 GND.n1732 394
R23058 GND.n8661 GND.n1732 394
R23059 GND.n8661 GND.n1730 394
R23060 GND.n8665 GND.n1730 394
R23061 GND.n8665 GND.n1008 394
R23062 GND.n8782 GND.n1008 394
R23063 GND.n8782 GND.n1009 394
R23064 GND.n8778 GND.n1009 394
R23065 GND.n8778 GND.n1012 394
R23066 GND.n8770 GND.n1012 394
R23067 GND.n8770 GND.n1024 394
R23068 GND.n8766 GND.n1024 394
R23069 GND.n8766 GND.n1026 394
R23070 GND.n8758 GND.n1026 394
R23071 GND.n8758 GND.n1036 394
R23072 GND.n8754 GND.n1036 394
R23073 GND.n8754 GND.n1038 394
R23074 GND.n8746 GND.n1038 394
R23075 GND.n8746 GND.n1048 394
R23076 GND.n8742 GND.n1048 394
R23077 GND.n8742 GND.n1050 394
R23078 GND.n8734 GND.n1050 394
R23079 GND.n8734 GND.n1060 394
R23080 GND.n8446 GND.n8445 394
R23081 GND.n8450 GND.n8449 394
R23082 GND.n8454 GND.n8453 394
R23083 GND.n8458 GND.n8457 394
R23084 GND.n8462 GND.n8461 394
R23085 GND.n8466 GND.n8465 394
R23086 GND.n8470 GND.n8469 394
R23087 GND.n8472 GND.n8440 394
R23088 GND.n8441 GND.n1796 394
R23089 GND.n8492 GND.n1796 394
R23090 GND.n8492 GND.n1790 394
R23091 GND.n8489 GND.n1790 394
R23092 GND.n8489 GND.n1784 394
R23093 GND.n8486 GND.n1784 394
R23094 GND.n8486 GND.n1778 394
R23095 GND.n8483 GND.n1778 394
R23096 GND.n8483 GND.n1772 394
R23097 GND.n8480 GND.n1772 394
R23098 GND.n8480 GND.n1766 394
R23099 GND.n8477 GND.n1766 394
R23100 GND.n8477 GND.n1759 394
R23101 GND.n1759 GND.n1750 394
R23102 GND.n8640 GND.n1750 394
R23103 GND.n8641 GND.n8640 394
R23104 GND.n8641 GND.n1746 394
R23105 GND.n8643 GND.n1746 394
R23106 GND.n8643 GND.n1740 394
R23107 GND.n1740 GND.n1736 394
R23108 GND.n8660 GND.n1736 394
R23109 GND.n8660 GND.n1726 394
R23110 GND.n8667 GND.n1726 394
R23111 GND.n8668 GND.n8667 394
R23112 GND.n8668 GND.n1005 394
R23113 GND.n8672 GND.n1005 394
R23114 GND.n8672 GND.n1013 394
R23115 GND.n8675 GND.n1013 394
R23116 GND.n8675 GND.n1021 394
R23117 GND.n8678 GND.n1021 394
R23118 GND.n8678 GND.n1027 394
R23119 GND.n8681 GND.n1027 394
R23120 GND.n8681 GND.n1033 394
R23121 GND.n8684 GND.n1033 394
R23122 GND.n8684 GND.n1039 394
R23123 GND.n8687 GND.n1039 394
R23124 GND.n8687 GND.n1045 394
R23125 GND.n8690 GND.n1045 394
R23126 GND.n8690 GND.n1051 394
R23127 GND.n8693 GND.n1051 394
R23128 GND.n8693 GND.n1057 394
R23129 GND.n8696 GND.n1057 394
R23130 GND.n8727 GND.n1062 394
R23131 GND.n8727 GND.n1723 394
R23132 GND.n8723 GND.n8722 394
R23133 GND.n8719 GND.n8718 394
R23134 GND.n8715 GND.n8714 394
R23135 GND.n8711 GND.n8710 394
R23136 GND.n8707 GND.n8706 394
R23137 GND.n8703 GND.n8702 394
R23138 GND.n8699 GND.n1070 394
R23139 GND.n3694 GND.n3140 394
R23140 GND.n3690 GND.n3140 394
R23141 GND.n3690 GND.n3143 394
R23142 GND.n3682 GND.n3143 394
R23143 GND.n3682 GND.n3155 394
R23144 GND.n3678 GND.n3155 394
R23145 GND.n3678 GND.n3157 394
R23146 GND.n3670 GND.n3157 394
R23147 GND.n3670 GND.n3167 394
R23148 GND.n3666 GND.n3167 394
R23149 GND.n3666 GND.n3169 394
R23150 GND.n3658 GND.n3169 394
R23151 GND.n3658 GND.n3179 394
R23152 GND.n3654 GND.n3179 394
R23153 GND.n3654 GND.n3181 394
R23154 GND.n3646 GND.n3181 394
R23155 GND.n3646 GND.n3191 394
R23156 GND.n3642 GND.n3191 394
R23157 GND.n3642 GND.n3193 394
R23158 GND.n3634 GND.n3193 394
R23159 GND.n3634 GND.n3264 394
R23160 GND.n3630 GND.n3264 394
R23161 GND.n3630 GND.n3266 394
R23162 GND.n3622 GND.n3266 394
R23163 GND.n3622 GND.n3278 394
R23164 GND.n3618 GND.n3278 394
R23165 GND.n3618 GND.n3280 394
R23166 GND.n3610 GND.n3280 394
R23167 GND.n3610 GND.n3293 394
R23168 GND.n3606 GND.n3293 394
R23169 GND.n3606 GND.n3295 394
R23170 GND.n3598 GND.n3295 394
R23171 GND.n3598 GND.n3308 394
R23172 GND.n3594 GND.n3308 394
R23173 GND.n3594 GND.n3310 394
R23174 GND.n3586 GND.n3310 394
R23175 GND.n3586 GND.n3320 394
R23176 GND.n3582 GND.n3320 394
R23177 GND.n3582 GND.n3322 394
R23178 GND.n3574 GND.n3322 394
R23179 GND.n3574 GND.n3332 394
R23180 GND.n3570 GND.n3332 394
R23181 GND.n3200 GND.n3199 394
R23182 GND.n3204 GND.n3203 394
R23183 GND.n3208 GND.n3207 394
R23184 GND.n3212 GND.n3211 394
R23185 GND.n3216 GND.n3215 394
R23186 GND.n3220 GND.n3219 394
R23187 GND.n3224 GND.n3223 394
R23188 GND.n3228 GND.n3227 394
R23189 GND.n3233 GND.n3135 394
R23190 GND.n3233 GND.n3144 394
R23191 GND.n3236 GND.n3144 394
R23192 GND.n3236 GND.n3152 394
R23193 GND.n3239 GND.n3152 394
R23194 GND.n3239 GND.n3158 394
R23195 GND.n3242 GND.n3158 394
R23196 GND.n3242 GND.n3164 394
R23197 GND.n3245 GND.n3164 394
R23198 GND.n3245 GND.n3170 394
R23199 GND.n3248 GND.n3170 394
R23200 GND.n3248 GND.n3176 394
R23201 GND.n3251 GND.n3176 394
R23202 GND.n3251 GND.n3182 394
R23203 GND.n3254 GND.n3182 394
R23204 GND.n3254 GND.n3188 394
R23205 GND.n3257 GND.n3188 394
R23206 GND.n3257 GND.n3194 394
R23207 GND.n3637 GND.n3194 394
R23208 GND.n3637 GND.n3636 394
R23209 GND.n3636 GND.n3261 394
R23210 GND.n3267 GND.n3261 394
R23211 GND.n3625 GND.n3267 394
R23212 GND.n3625 GND.n3624 394
R23213 GND.n3624 GND.n3274 394
R23214 GND.n3281 GND.n3274 394
R23215 GND.n3613 GND.n3281 394
R23216 GND.n3613 GND.n3612 394
R23217 GND.n3612 GND.n3288 394
R23218 GND.n3296 GND.n3288 394
R23219 GND.n3348 GND.n3296 394
R23220 GND.n3348 GND.n3305 394
R23221 GND.n3351 GND.n3305 394
R23222 GND.n3351 GND.n3311 394
R23223 GND.n3354 GND.n3311 394
R23224 GND.n3354 GND.n3317 394
R23225 GND.n3357 GND.n3317 394
R23226 GND.n3357 GND.n3323 394
R23227 GND.n3360 GND.n3323 394
R23228 GND.n3360 GND.n3329 394
R23229 GND.n3363 GND.n3329 394
R23230 GND.n3363 GND.n3335 394
R23231 GND.n3397 GND.n3345 394
R23232 GND.n3393 GND.n3345 394
R23233 GND.n3391 GND.n3390 394
R23234 GND.n3387 GND.n3386 394
R23235 GND.n3383 GND.n3382 394
R23236 GND.n3379 GND.n3378 394
R23237 GND.n3375 GND.n3374 394
R23238 GND.n3371 GND.n3370 394
R23239 GND.n3367 GND.n3344 394
R23240 GND.n8594 GND.n1798 394
R23241 GND.n8594 GND.n1788 394
R23242 GND.n8602 GND.n1788 394
R23243 GND.n8602 GND.n1786 394
R23244 GND.n8606 GND.n1786 394
R23245 GND.n8606 GND.n1776 394
R23246 GND.n8614 GND.n1776 394
R23247 GND.n8614 GND.n1774 394
R23248 GND.n8618 GND.n1774 394
R23249 GND.n8618 GND.n1764 394
R23250 GND.n8626 GND.n1764 394
R23251 GND.n8626 GND.n1761 394
R23252 GND.n8632 GND.n1761 394
R23253 GND.n8632 GND.n1762 394
R23254 GND.n1762 GND.n1754 394
R23255 GND.n1754 GND.n1748 394
R23256 GND.n8646 GND.n1748 394
R23257 GND.n8646 GND.n1738 394
R23258 GND.n8654 GND.n1738 394
R23259 GND.n8655 GND.n8654 394
R23260 GND.n8655 GND.n1734 394
R23261 GND.n8657 GND.n1734 394
R23262 GND.n8657 GND.n1729 394
R23263 GND.n1729 GND.n1725 394
R23264 GND.n1725 GND.n1007 394
R23265 GND.n1016 GND.n1007 394
R23266 GND.n8776 GND.n1016 394
R23267 GND.n8776 GND.n1017 394
R23268 GND.n8772 GND.n1017 394
R23269 GND.n8772 GND.n1020 394
R23270 GND.n8764 GND.n1020 394
R23271 GND.n8764 GND.n1030 394
R23272 GND.n8760 GND.n1030 394
R23273 GND.n8760 GND.n1032 394
R23274 GND.n8752 GND.n1032 394
R23275 GND.n8752 GND.n1042 394
R23276 GND.n8748 GND.n1042 394
R23277 GND.n8748 GND.n1044 394
R23278 GND.n8740 GND.n1044 394
R23279 GND.n8740 GND.n1054 394
R23280 GND.n8736 GND.n1054 394
R23281 GND.n8736 GND.n1056 394
R23282 GND.n8588 GND.n8587 394
R23283 GND.n8585 GND.n8501 394
R23284 GND.n8581 GND.n8580 394
R23285 GND.n8578 GND.n8504 394
R23286 GND.n8574 GND.n8573 394
R23287 GND.n8571 GND.n8507 394
R23288 GND.n8567 GND.n8566 394
R23289 GND.n8564 GND.n8510 394
R23290 GND.n8559 GND.n1797 394
R23291 GND.n8554 GND.n1797 394
R23292 GND.n8554 GND.n1791 394
R23293 GND.n8551 GND.n1791 394
R23294 GND.n8551 GND.n1785 394
R23295 GND.n8548 GND.n1785 394
R23296 GND.n8548 GND.n1779 394
R23297 GND.n8545 GND.n1779 394
R23298 GND.n8545 GND.n1773 394
R23299 GND.n8542 GND.n1773 394
R23300 GND.n8542 GND.n1767 394
R23301 GND.n8539 GND.n1767 394
R23302 GND.n8539 GND.n1760 394
R23303 GND.n8536 GND.n1760 394
R23304 GND.n8536 GND.n1753 394
R23305 GND.n8533 GND.n1753 394
R23306 GND.n8533 GND.n1747 394
R23307 GND.n8514 GND.n1747 394
R23308 GND.n8514 GND.n1741 394
R23309 GND.n8523 GND.n1741 394
R23310 GND.n8523 GND.n1735 394
R23311 GND.n8520 GND.n1735 394
R23312 GND.n8520 GND.n1728 394
R23313 GND.n1728 GND.n1002 394
R23314 GND.n8784 GND.n1002 394
R23315 GND.n8784 GND.n1003 394
R23316 GND.n1014 GND.n1003 394
R23317 GND.n1664 GND.n1014 394
R23318 GND.n1664 GND.n1022 394
R23319 GND.n1667 GND.n1022 394
R23320 GND.n1667 GND.n1028 394
R23321 GND.n1670 GND.n1028 394
R23322 GND.n1670 GND.n1034 394
R23323 GND.n1673 GND.n1034 394
R23324 GND.n1673 GND.n1040 394
R23325 GND.n1676 GND.n1040 394
R23326 GND.n1676 GND.n1046 394
R23327 GND.n1679 GND.n1046 394
R23328 GND.n1679 GND.n1052 394
R23329 GND.n1682 GND.n1052 394
R23330 GND.n1682 GND.n1058 394
R23331 GND.n1686 GND.n1058 394
R23332 GND.n1717 GND.n1662 394
R23333 GND.n1715 GND.n1714 394
R23334 GND.n1711 GND.n1710 394
R23335 GND.n1707 GND.n1706 394
R23336 GND.n1703 GND.n1702 394
R23337 GND.n1699 GND.n1698 394
R23338 GND.n1695 GND.n1694 394
R23339 GND.n1691 GND.n1690 394
R23340 GND.n9200 GND.n9198 394
R23341 GND.n9198 GND.n9197 394
R23342 GND.n9194 GND.n9193 394
R23343 GND.n9191 GND.n9143 394
R23344 GND.n9187 GND.n9185 394
R23345 GND.n9183 GND.n9145 394
R23346 GND.n9179 GND.n9177 394
R23347 GND.n9175 GND.n9147 394
R23348 GND.n631 GND.n574 394
R23349 GND.n631 GND.n575 394
R23350 GND.n575 GND.n567 394
R23351 GND.n626 GND.n567 394
R23352 GND.n626 GND.n625 394
R23353 GND.n625 GND.n555 394
R23354 GND.n621 GND.n555 394
R23355 GND.n621 GND.n548 394
R23356 GND.n548 GND.n540 394
R23357 GND.n713 GND.n540 394
R23358 GND.n713 GND.n531 394
R23359 GND.n537 GND.n531 394
R23360 GND.n723 GND.n537 394
R23361 GND.n723 GND.n538 394
R23362 GND.n538 GND.n199 394
R23363 GND.n859 GND.n199 394
R23364 GND.n859 GND.n209 394
R23365 GND.n866 GND.n209 394
R23366 GND.n867 GND.n866 394
R23367 GND.n867 GND.n493 394
R23368 GND.n908 GND.n493 394
R23369 GND.n908 GND.n495 394
R23370 GND.n495 GND.n477 394
R23371 GND.n899 GND.n477 394
R23372 GND.n899 GND.n465 394
R23373 GND.n893 GND.n465 394
R23374 GND.n893 GND.n892 394
R23375 GND.n892 GND.n886 394
R23376 GND.n886 GND.n449 394
R23377 GND.n449 GND.n359 394
R23378 GND.n9267 GND.n359 394
R23379 GND.n9267 GND.n360 394
R23380 GND.n360 GND.n350 394
R23381 GND.n9258 GND.n350 394
R23382 GND.n9258 GND.n323 394
R23383 GND.n9252 GND.n323 394
R23384 GND.n9252 GND.n333 394
R23385 GND.n369 GND.n333 394
R23386 GND.n9244 GND.n369 394
R23387 GND.n9244 GND.n370 394
R23388 GND.n381 GND.n370 394
R23389 GND.n9151 GND.n381 394
R23390 GND.n9152 GND.n9151 394
R23391 GND.n9152 GND.n393 394
R23392 GND.n9156 GND.n393 394
R23393 GND.n9156 GND.n401 394
R23394 GND.n9160 GND.n401 394
R23395 GND.n9161 GND.n9160 394
R23396 GND.n9161 GND.n411 394
R23397 GND.n9165 GND.n411 394
R23398 GND.n9165 GND.n9136 394
R23399 GND.n9137 GND.n9136 394
R23400 GND.n9138 GND.n9137 394
R23401 GND.n614 GND.n585 394
R23402 GND.n610 GND.n609 394
R23403 GND.n606 GND.n605 394
R23404 GND.n602 GND.n601 394
R23405 GND.n598 GND.n597 394
R23406 GND.n594 GND.n593 394
R23407 GND.n590 GND.n589 394
R23408 GND.n586 GND.n577 394
R23409 GND.n633 GND.n572 394
R23410 GND.n633 GND.n569 394
R23411 GND.n638 GND.n569 394
R23412 GND.n638 GND.n570 394
R23413 GND.n570 GND.n554 394
R23414 GND.n697 GND.n554 394
R23415 GND.n697 GND.n550 394
R23416 GND.n702 GND.n550 394
R23417 GND.n702 GND.n552 394
R23418 GND.n552 GND.n532 394
R23419 GND.n729 GND.n532 394
R23420 GND.n729 GND.n533 394
R23421 GND.n725 GND.n533 394
R23422 GND.n725 GND.n201 394
R23423 GND.n9423 GND.n201 394
R23424 GND.n9423 GND.n202 394
R23425 GND.n9416 GND.n202 394
R23426 GND.n9416 GND.n208 394
R23427 GND.n915 GND.n208 394
R23428 GND.n915 GND.n909 394
R23429 GND.n924 GND.n909 394
R23430 GND.n924 GND.n478 394
R23431 GND.n947 GND.n478 394
R23432 GND.n947 GND.n466 394
R23433 GND.n8973 GND.n466 394
R23434 GND.n8973 GND.n467 394
R23435 GND.n890 GND.n467 394
R23436 GND.n890 GND.n450 394
R23437 GND.n9044 GND.n450 394
R23438 GND.n9044 GND.n357 394
R23439 GND.n9269 GND.n357 394
R23440 GND.n9269 GND.n352 394
R23441 GND.n9278 GND.n352 394
R23442 GND.n9278 GND.n325 394
R23443 GND.n9308 GND.n325 394
R23444 GND.n9308 GND.n326 394
R23445 GND.n9301 GND.n326 394
R23446 GND.n9301 GND.n332 394
R23447 GND.n9242 GND.n332 394
R23448 GND.n9242 GND.n373 394
R23449 GND.n9236 GND.n373 394
R23450 GND.n9236 GND.n377 394
R23451 GND.n395 GND.n377 394
R23452 GND.n9226 GND.n395 394
R23453 GND.n9226 GND.n396 394
R23454 GND.n9222 GND.n396 394
R23455 GND.n9222 GND.n399 394
R23456 GND.n413 GND.n399 394
R23457 GND.n9212 GND.n413 394
R23458 GND.n9212 GND.n414 394
R23459 GND.n9208 GND.n414 394
R23460 GND.n9208 GND.n417 394
R23461 GND.n9204 GND.n417 394
R23462 GND.n426 GND.n425 394
R23463 GND.n9128 GND.n425 394
R23464 GND.n9126 GND.n9125 394
R23465 GND.n9122 GND.n9121 394
R23466 GND.n9118 GND.n9117 394
R23467 GND.n9114 GND.n9113 394
R23468 GND.n9110 GND.n9109 394
R23469 GND.n9106 GND.n9105 394
R23470 GND.n686 GND.n558 394
R23471 GND.n686 GND.n556 394
R23472 GND.n694 GND.n556 394
R23473 GND.n694 GND.n547 394
R23474 GND.n690 GND.n547 394
R23475 GND.n690 GND.n541 394
R23476 GND.n541 GND.n529 394
R23477 GND.n732 GND.n529 394
R23478 GND.n732 GND.n191 394
R23479 GND.n736 GND.n191 394
R23480 GND.n736 GND.n198 394
R23481 GND.n740 GND.n198 394
R23482 GND.n740 GND.n503 394
R23483 GND.n503 GND.n210 394
R23484 GND.n751 GND.n210 394
R23485 GND.n751 GND.n225 394
R23486 GND.n928 GND.n225 394
R23487 GND.n928 GND.n486 394
R23488 GND.n936 GND.n486 394
R23489 GND.n937 GND.n936 394
R23490 GND.n938 GND.n937 394
R23491 GND.n938 GND.n456 394
R23492 GND.n9031 GND.n456 394
R23493 GND.n9032 GND.n9031 394
R23494 GND.n9032 GND.n446 394
R23495 GND.n446 GND.n437 394
R23496 GND.n9060 GND.n437 394
R23497 GND.n9060 GND.n438 394
R23498 GND.n438 GND.n347 394
R23499 GND.n9068 GND.n347 394
R23500 GND.n9068 GND.n431 394
R23501 GND.n9075 GND.n431 394
R23502 GND.n9076 GND.n9075 394
R23503 GND.n9076 GND.n334 394
R23504 GND.n9082 GND.n334 394
R23505 GND.n9083 GND.n9082 394
R23506 GND.n9084 GND.n9083 394
R23507 GND.n9084 GND.n382 394
R23508 GND.n9088 GND.n382 394
R23509 GND.n9088 GND.n392 394
R23510 GND.n9092 GND.n392 394
R23511 GND.n9093 GND.n9092 394
R23512 GND.n9093 GND.n402 394
R23513 GND.n9097 GND.n402 394
R23514 GND.n9097 GND.n410 394
R23515 GND.n9101 GND.n410 394
R23516 GND.n679 GND.n565 394
R23517 GND.n676 GND.n647 394
R23518 GND.n672 GND.n671 394
R23519 GND.n668 GND.n667 394
R23520 GND.n664 GND.n663 394
R23521 GND.n660 GND.n659 394
R23522 GND.n656 GND.n655 394
R23523 GND.n652 GND.n651 394
R23524 GND.n684 GND.n561 394
R23525 GND.n684 GND.n563 394
R23526 GND.n563 GND.n545 394
R23527 GND.n705 GND.n545 394
R23528 GND.n705 GND.n542 394
R23529 GND.n710 GND.n542 394
R23530 GND.n710 GND.n543 394
R23531 GND.n543 GND.n192 394
R23532 GND.n9430 GND.n192 394
R23533 GND.n9430 GND.n193 394
R23534 GND.n9426 GND.n193 394
R23535 GND.n9426 GND.n196 394
R23536 GND.n212 GND.n196 394
R23537 GND.n9413 GND.n212 394
R23538 GND.n9413 GND.n213 394
R23539 GND.n9406 GND.n213 394
R23540 GND.n9406 GND.n223 394
R23541 GND.n829 GND.n223 394
R23542 GND.n838 GND.n829 394
R23543 GND.n839 GND.n838 394
R23544 GND.n840 GND.n839 394
R23545 GND.n840 GND.n457 394
R23546 GND.n9029 GND.n457 394
R23547 GND.n9029 GND.n445 394
R23548 GND.n9048 GND.n445 394
R23549 GND.n9048 GND.n439 394
R23550 GND.n9058 GND.n439 394
R23551 GND.n9058 GND.n346 394
R23552 GND.n9282 GND.n346 394
R23553 GND.n9282 GND.n342 394
R23554 GND.n9289 GND.n342 394
R23555 GND.n9290 GND.n9289 394
R23556 GND.n9290 GND.n336 394
R23557 GND.n9298 GND.n336 394
R23558 GND.n9298 GND.n337 394
R23559 GND.n386 GND.n337 394
R23560 GND.n386 GND.n384 394
R23561 GND.n9233 GND.n384 394
R23562 GND.n9233 GND.n385 394
R23563 GND.n9229 GND.n385 394
R23564 GND.n9229 GND.n390 394
R23565 GND.n404 GND.n390 394
R23566 GND.n9219 GND.n404 394
R23567 GND.n9219 GND.n405 394
R23568 GND.n9215 GND.n405 394
R23569 GND.n9215 GND.n408 394
R23570 GND.n9403 GND.n229 394
R23571 GND.n9403 GND.n230 394
R23572 GND.n9399 GND.n230 394
R23573 GND.n9399 GND.n233 394
R23574 GND.n9389 GND.n233 394
R23575 GND.n9389 GND.n248 394
R23576 GND.n9382 GND.n248 394
R23577 GND.n9382 GND.n255 394
R23578 GND.n9374 GND.n255 394
R23579 GND.n9374 GND.n270 394
R23580 GND.n9367 GND.n270 394
R23581 GND.n9367 GND.n274 394
R23582 GND.n9357 GND.n274 394
R23583 GND.n9357 GND.n290 394
R23584 GND.n9353 GND.n290 394
R23585 GND.n9353 GND.n294 394
R23586 GND.n755 GND.n504 394
R23587 GND.n759 GND.n758 394
R23588 GND.n763 GND.n762 394
R23589 GND.n767 GND.n766 394
R23590 GND.n771 GND.n770 394
R23591 GND.n775 GND.n774 394
R23592 GND.n779 GND.n778 394
R23593 GND.n783 GND.n782 394
R23594 GND.n790 GND.n226 394
R23595 GND.n491 GND.n226 394
R23596 GND.n491 GND.n235 394
R23597 GND.n950 GND.n235 394
R23598 GND.n950 GND.n245 394
R23599 GND.n464 GND.n245 394
R23600 GND.n464 GND.n257 394
R23601 GND.n960 GND.n257 394
R23602 GND.n960 GND.n267 394
R23603 GND.n447 GND.n267 394
R23604 GND.n447 GND.n276 394
R23605 GND.n970 GND.n276 394
R23606 GND.n970 GND.n287 394
R23607 GND.n348 GND.n287 394
R23608 GND.n348 GND.n295 394
R23609 GND.n9311 GND.n295 394
R23610 GND.n319 GND.n318 394
R23611 GND.n9338 GND.n318 394
R23612 GND.n9336 GND.n9335 394
R23613 GND.n9332 GND.n9331 394
R23614 GND.n9328 GND.n9327 394
R23615 GND.n9324 GND.n9323 394
R23616 GND.n9320 GND.n9319 394
R23617 GND.n9316 GND.n9315 394
R23618 GND.n792 GND.n228 394
R23619 GND.n237 GND.n228 394
R23620 GND.n9397 GND.n237 394
R23621 GND.n9397 GND.n238 394
R23622 GND.n9391 GND.n238 394
R23623 GND.n9391 GND.n243 394
R23624 GND.n9380 GND.n243 394
R23625 GND.n9380 GND.n260 394
R23626 GND.n9376 GND.n260 394
R23627 GND.n9376 GND.n265 394
R23628 GND.n9365 GND.n265 394
R23629 GND.n9365 GND.n279 394
R23630 GND.n9359 GND.n279 394
R23631 GND.n9359 GND.n285 394
R23632 GND.n9351 GND.n285 394
R23633 GND.n9351 GND.n298 394
R23634 GND.n8983 GND.n300 394
R23635 GND.n8987 GND.n8986 394
R23636 GND.n8991 GND.n8990 394
R23637 GND.n8995 GND.n8994 394
R23638 GND.n8999 GND.n8998 394
R23639 GND.n9003 GND.n9002 394
R23640 GND.n9007 GND.n9006 394
R23641 GND.n9009 GND.n316 394
R23642 GND.n522 GND.n227 394
R23643 GND.n492 GND.n227 394
R23644 GND.n492 GND.n236 394
R23645 GND.n476 GND.n236 394
R23646 GND.n476 GND.n246 394
R23647 GND.n8976 GND.n246 394
R23648 GND.n8976 GND.n258 394
R23649 GND.n8980 GND.n258 394
R23650 GND.n8980 GND.n268 394
R23651 GND.n448 GND.n268 394
R23652 GND.n448 GND.n277 394
R23653 GND.n8981 GND.n277 394
R23654 GND.n8981 GND.n288 394
R23655 GND.n349 GND.n288 394
R23656 GND.n349 GND.n296 394
R23657 GND.n322 GND.n296 394
R23658 GND.n797 GND.n796 394
R23659 GND.n801 GND.n800 394
R23660 GND.n805 GND.n804 394
R23661 GND.n809 GND.n808 394
R23662 GND.n813 GND.n812 394
R23663 GND.n817 GND.n816 394
R23664 GND.n821 GND.n820 394
R23665 GND.n855 GND.n521 394
R23666 GND.n3147 GND.n3138 394
R23667 GND.n3688 GND.n3147 394
R23668 GND.n3688 GND.n3148 394
R23669 GND.n3684 GND.n3148 394
R23670 GND.n3684 GND.n3151 394
R23671 GND.n3676 GND.n3151 394
R23672 GND.n3676 GND.n3161 394
R23673 GND.n3672 GND.n3161 394
R23674 GND.n3672 GND.n3163 394
R23675 GND.n3664 GND.n3163 394
R23676 GND.n3664 GND.n3173 394
R23677 GND.n3660 GND.n3173 394
R23678 GND.n3660 GND.n3175 394
R23679 GND.n3652 GND.n3175 394
R23680 GND.n3652 GND.n3185 394
R23681 GND.n3648 GND.n3185 394
R23682 GND.n3648 GND.n3187 394
R23683 GND.n3640 GND.n3187 394
R23684 GND.n3640 GND.n3197 394
R23685 GND.n3263 GND.n3197 394
R23686 GND.n3270 GND.n3263 394
R23687 GND.n3628 GND.n3270 394
R23688 GND.n3628 GND.n3271 394
R23689 GND.n3277 GND.n3271 394
R23690 GND.n3284 GND.n3277 394
R23691 GND.n3616 GND.n3284 394
R23692 GND.n3616 GND.n3285 394
R23693 GND.n3292 GND.n3285 394
R23694 GND.n3299 GND.n3292 394
R23695 GND.n3604 GND.n3299 394
R23696 GND.n3604 GND.n3300 394
R23697 GND.n3600 GND.n3300 394
R23698 GND.n3600 GND.n3304 394
R23699 GND.n3592 GND.n3304 394
R23700 GND.n3592 GND.n3314 394
R23701 GND.n3588 GND.n3314 394
R23702 GND.n3588 GND.n3316 394
R23703 GND.n3580 GND.n3316 394
R23704 GND.n3580 GND.n3326 394
R23705 GND.n3576 GND.n3326 394
R23706 GND.n3576 GND.n3328 394
R23707 GND.n3568 GND.n3328 394
R23708 GND.n3421 GND.n3420 394
R23709 GND.n3425 GND.n3424 394
R23710 GND.n3429 GND.n3428 394
R23711 GND.n3433 GND.n3432 394
R23712 GND.n3437 GND.n3436 394
R23713 GND.n3441 GND.n3440 394
R23714 GND.n3445 GND.n3444 394
R23715 GND.n3449 GND.n3448 394
R23716 GND.n3454 GND.n3136 394
R23717 GND.n3454 GND.n3145 394
R23718 GND.n3457 GND.n3145 394
R23719 GND.n3457 GND.n3153 394
R23720 GND.n3460 GND.n3153 394
R23721 GND.n3460 GND.n3159 394
R23722 GND.n3463 GND.n3159 394
R23723 GND.n3463 GND.n3165 394
R23724 GND.n3466 GND.n3165 394
R23725 GND.n3466 GND.n3171 394
R23726 GND.n3469 GND.n3171 394
R23727 GND.n3469 GND.n3177 394
R23728 GND.n3472 GND.n3177 394
R23729 GND.n3472 GND.n3183 394
R23730 GND.n3475 GND.n3183 394
R23731 GND.n3475 GND.n3189 394
R23732 GND.n3478 GND.n3189 394
R23733 GND.n3478 GND.n3195 394
R23734 GND.n3483 GND.n3195 394
R23735 GND.n3483 GND.n3262 394
R23736 GND.n3496 GND.n3262 394
R23737 GND.n3496 GND.n3268 394
R23738 GND.n3493 GND.n3268 394
R23739 GND.n3493 GND.n3275 394
R23740 GND.n3488 GND.n3275 394
R23741 GND.n3488 GND.n3282 394
R23742 GND.n3507 GND.n3282 394
R23743 GND.n3507 GND.n3290 394
R23744 GND.n3510 GND.n3290 394
R23745 GND.n3510 GND.n3297 394
R23746 GND.n3513 GND.n3297 394
R23747 GND.n3513 GND.n3306 394
R23748 GND.n3516 GND.n3306 394
R23749 GND.n3516 GND.n3312 394
R23750 GND.n3519 GND.n3312 394
R23751 GND.n3519 GND.n3318 394
R23752 GND.n3522 GND.n3318 394
R23753 GND.n3522 GND.n3324 394
R23754 GND.n3525 GND.n3324 394
R23755 GND.n3525 GND.n3330 394
R23756 GND.n3528 GND.n3330 394
R23757 GND.n3528 GND.n3336 394
R23758 GND.n3564 GND.n3562 394
R23759 GND.n3560 GND.n3402 394
R23760 GND.n3556 GND.n3554 394
R23761 GND.n3552 GND.n3404 394
R23762 GND.n3548 GND.n3546 394
R23763 GND.n3544 GND.n3406 394
R23764 GND.n3540 GND.n3538 394
R23765 GND.n3536 GND.n3408 394
R23766 GND.n8094 GND.n8092 394
R23767 GND.n8092 GND.n8091 394
R23768 GND.n8088 GND.n8087 394
R23769 GND.n8085 GND.n8037 394
R23770 GND.n8081 GND.n8079 394
R23771 GND.n8077 GND.n8039 394
R23772 GND.n8073 GND.n8071 394
R23773 GND.n8069 GND.n8041 394
R23774 GND.n8362 GND.n8361 394
R23775 GND.n8361 GND.n1829 394
R23776 GND.n1836 GND.n1829 394
R23777 GND.n1877 GND.n1836 394
R23778 GND.n1878 GND.n1877 394
R23779 GND.n1878 GND.n1846 394
R23780 GND.n1882 GND.n1846 394
R23781 GND.n1882 GND.n1854 394
R23782 GND.n1886 GND.n1854 394
R23783 GND.n1887 GND.n1886 394
R23784 GND.n1887 GND.n1864 394
R23785 GND.n1872 GND.n1864 394
R23786 GND.n8325 GND.n1872 394
R23787 GND.n8325 GND.n1873 394
R23788 GND.n8319 GND.n1873 394
R23789 GND.n8319 GND.n1894 394
R23790 GND.n1905 GND.n1894 394
R23791 GND.n4243 GND.n1905 394
R23792 GND.n4244 GND.n4243 394
R23793 GND.n4244 GND.n4232 394
R23794 GND.n4523 GND.n4232 394
R23795 GND.n4525 GND.n4523 394
R23796 GND.n4525 GND.n4216 394
R23797 GND.n4226 GND.n4216 394
R23798 GND.n4671 GND.n4226 394
R23799 GND.n4671 GND.n4227 394
R23800 GND.n4536 GND.n4227 394
R23801 GND.n4663 GND.n4536 394
R23802 GND.n4663 GND.n4662 394
R23803 GND.n4662 GND.n2051 394
R23804 GND.n8161 GND.n2051 394
R23805 GND.n8161 GND.n2052 394
R23806 GND.n2052 GND.n2042 394
R23807 GND.n8152 GND.n2042 394
R23808 GND.n8152 GND.n2015 394
R23809 GND.n8146 GND.n2015 394
R23810 GND.n8146 GND.n2025 394
R23811 GND.n2061 GND.n2025 394
R23812 GND.n8138 GND.n2061 394
R23813 GND.n8138 GND.n2062 394
R23814 GND.n2071 GND.n2062 394
R23815 GND.n8045 GND.n2071 394
R23816 GND.n8046 GND.n8045 394
R23817 GND.n8046 GND.n2083 394
R23818 GND.n8050 GND.n2083 394
R23819 GND.n8050 GND.n2091 394
R23820 GND.n8054 GND.n2091 394
R23821 GND.n8055 GND.n8054 394
R23822 GND.n8055 GND.n2101 394
R23823 GND.n8059 GND.n2101 394
R23824 GND.n8059 GND.n2109 394
R23825 GND.n2110 GND.n2109 394
R23826 GND.n2111 GND.n2110 394
R23827 GND.n8395 GND.n1826 394
R23828 GND.n8391 GND.n8390 394
R23829 GND.n8387 GND.n8386 394
R23830 GND.n8383 GND.n8382 394
R23831 GND.n8379 GND.n8378 394
R23832 GND.n8375 GND.n8374 394
R23833 GND.n8371 GND.n8370 394
R23834 GND.n8367 GND.n8366 394
R23835 GND.n8359 GND.n1825 394
R23836 GND.n8359 GND.n1831 394
R23837 GND.n8355 GND.n1831 394
R23838 GND.n8355 GND.n1833 394
R23839 GND.n1848 GND.n1833 394
R23840 GND.n8345 GND.n1848 394
R23841 GND.n8345 GND.n1849 394
R23842 GND.n8341 GND.n1849 394
R23843 GND.n8341 GND.n1852 394
R23844 GND.n1866 GND.n1852 394
R23845 GND.n8331 GND.n1866 394
R23846 GND.n8331 GND.n1867 394
R23847 GND.n8327 GND.n1867 394
R23848 GND.n8327 GND.n1870 394
R23849 GND.n8317 GND.n1870 394
R23850 GND.n8317 GND.n1897 394
R23851 GND.n8310 GND.n1897 394
R23852 GND.n8310 GND.n1904 394
R23853 GND.n4512 GND.n1904 394
R23854 GND.n4512 GND.n4506 394
R23855 GND.n4521 GND.n4506 394
R23856 GND.n4521 GND.n4217 394
R23857 GND.n4681 GND.n4217 394
R23858 GND.n4681 GND.n4218 394
R23859 GND.n4673 GND.n4218 394
R23860 GND.n4673 GND.n4225 394
R23861 GND.n4543 GND.n4225 394
R23862 GND.n4543 GND.n4541 394
R23863 GND.n4660 GND.n4541 394
R23864 GND.n4660 GND.n2049 394
R23865 GND.n8163 GND.n2049 394
R23866 GND.n8163 GND.n2044 394
R23867 GND.n8172 GND.n2044 394
R23868 GND.n8172 GND.n2017 394
R23869 GND.n8202 GND.n2017 394
R23870 GND.n8202 GND.n2018 394
R23871 GND.n8195 GND.n2018 394
R23872 GND.n8195 GND.n2024 394
R23873 GND.n8136 GND.n2024 394
R23874 GND.n8136 GND.n2065 394
R23875 GND.n8130 GND.n2065 394
R23876 GND.n8130 GND.n2069 394
R23877 GND.n2085 GND.n2069 394
R23878 GND.n8120 GND.n2085 394
R23879 GND.n8120 GND.n2086 394
R23880 GND.n8116 GND.n2086 394
R23881 GND.n8116 GND.n2089 394
R23882 GND.n2103 GND.n2089 394
R23883 GND.n8106 GND.n2103 394
R23884 GND.n8106 GND.n2104 394
R23885 GND.n8102 GND.n2104 394
R23886 GND.n8102 GND.n2107 394
R23887 GND.n8098 GND.n2107 394
R23888 GND.n4570 GND.n4566 394
R23889 GND.n4574 GND.n4566 394
R23890 GND.n4578 GND.n4576 394
R23891 GND.n4582 GND.n4564 394
R23892 GND.n4586 GND.n4584 394
R23893 GND.n4590 GND.n4562 394
R23894 GND.n4594 GND.n4592 394
R23895 GND.n4598 GND.n4560 394
R23896 GND.n4318 GND.n1837 394
R23897 GND.n4318 GND.n1845 394
R23898 GND.n4322 GND.n1845 394
R23899 GND.n4323 GND.n4322 394
R23900 GND.n4323 GND.n1855 394
R23901 GND.n4327 GND.n1855 394
R23902 GND.n4327 GND.n1863 394
R23903 GND.n4275 GND.n1863 394
R23904 GND.n4332 GND.n4275 394
R23905 GND.n4347 GND.n4332 394
R23906 GND.n4348 GND.n4347 394
R23907 GND.n4348 GND.n4271 394
R23908 GND.n4356 GND.n4271 394
R23909 GND.n4356 GND.n1906 394
R23910 GND.n4450 GND.n1906 394
R23911 GND.n4450 GND.n1917 394
R23912 GND.n4252 GND.n1917 394
R23913 GND.n4459 GND.n4252 394
R23914 GND.n4459 GND.n4458 394
R23915 GND.n4458 GND.n4258 394
R23916 GND.n4469 GND.n4258 394
R23917 GND.n4469 GND.n4259 394
R23918 GND.n4259 GND.n4192 394
R23919 GND.n4773 GND.n4192 394
R23920 GND.n4773 GND.n4772 394
R23921 GND.n4772 GND.n4194 394
R23922 GND.n4648 GND.n4194 394
R23923 GND.n4648 GND.n4640 394
R23924 GND.n4640 GND.n2039 394
R23925 GND.n4633 GND.n2039 394
R23926 GND.n4633 GND.n4632 394
R23927 GND.n4632 GND.n4555 394
R23928 GND.n4625 GND.n4555 394
R23929 GND.n4625 GND.n2026 394
R23930 GND.n4620 GND.n2026 394
R23931 GND.n4620 GND.n4619 394
R23932 GND.n4619 GND.n4618 394
R23933 GND.n4618 GND.n2072 394
R23934 GND.n4614 GND.n2072 394
R23935 GND.n4614 GND.n2082 394
R23936 GND.n4610 GND.n2082 394
R23937 GND.n4610 GND.n4609 394
R23938 GND.n4609 GND.n2092 394
R23939 GND.n4605 GND.n2092 394
R23940 GND.n4605 GND.n2100 394
R23941 GND.n4601 GND.n2100 394
R23942 GND.n4285 GND.n1839 394
R23943 GND.n4289 GND.n4283 394
R23944 GND.n4293 GND.n4291 394
R23945 GND.n4297 GND.n4281 394
R23946 GND.n4301 GND.n4299 394
R23947 GND.n4305 GND.n4279 394
R23948 GND.n4308 GND.n4307 394
R23949 GND.n4312 GND.n4311 394
R23950 GND.n8352 GND.n1840 394
R23951 GND.n8348 GND.n1840 394
R23952 GND.n8348 GND.n1843 394
R23953 GND.n1857 GND.n1843 394
R23954 GND.n8338 GND.n1857 394
R23955 GND.n8338 GND.n1858 394
R23956 GND.n8334 GND.n1858 394
R23957 GND.n8334 GND.n1861 394
R23958 GND.n4334 GND.n1861 394
R23959 GND.n4345 GND.n4334 394
R23960 GND.n4345 GND.n4335 394
R23961 GND.n4337 GND.n4335 394
R23962 GND.n4337 GND.n1908 394
R23963 GND.n8307 GND.n1908 394
R23964 GND.n8307 GND.n1909 394
R23965 GND.n8300 GND.n1909 394
R23966 GND.n8300 GND.n1915 394
R23967 GND.n4478 GND.n1915 394
R23968 GND.n4479 GND.n4478 394
R23969 GND.n4479 GND.n4470 394
R23970 GND.n4489 GND.n4470 394
R23971 GND.n4489 GND.n4209 394
R23972 GND.n4715 GND.n4209 394
R23973 GND.n4715 GND.n4197 394
R23974 GND.n4770 GND.n4197 394
R23975 GND.n4770 GND.n4198 394
R23976 GND.n4646 GND.n4198 394
R23977 GND.n4646 GND.n2038 394
R23978 GND.n8176 GND.n2038 394
R23979 GND.n8176 GND.n2034 394
R23980 GND.n8183 GND.n2034 394
R23981 GND.n8184 GND.n8183 394
R23982 GND.n8184 GND.n2028 394
R23983 GND.n8192 GND.n2028 394
R23984 GND.n8192 GND.n2029 394
R23985 GND.n2076 GND.n2029 394
R23986 GND.n2076 GND.n2074 394
R23987 GND.n8127 GND.n2074 394
R23988 GND.n8127 GND.n2075 394
R23989 GND.n8123 GND.n2075 394
R23990 GND.n8123 GND.n2080 394
R23991 GND.n2094 GND.n2080 394
R23992 GND.n8113 GND.n2094 394
R23993 GND.n8113 GND.n2095 394
R23994 GND.n8109 GND.n2095 394
R23995 GND.n8109 GND.n2098 394
R23996 GND.n8297 GND.n1921 394
R23997 GND.n8297 GND.n1922 394
R23998 GND.n8293 GND.n1922 394
R23999 GND.n8293 GND.n1925 394
R24000 GND.n8283 GND.n1925 394
R24001 GND.n8283 GND.n1940 394
R24002 GND.n8276 GND.n1940 394
R24003 GND.n8276 GND.n1947 394
R24004 GND.n8268 GND.n1947 394
R24005 GND.n8268 GND.n1962 394
R24006 GND.n8261 GND.n1962 394
R24007 GND.n8261 GND.n1966 394
R24008 GND.n8251 GND.n1966 394
R24009 GND.n8251 GND.n1982 394
R24010 GND.n8247 GND.n1982 394
R24011 GND.n8247 GND.n1986 394
R24012 GND.n4368 GND.n4358 394
R24013 GND.n4372 GND.n4371 394
R24014 GND.n4376 GND.n4375 394
R24015 GND.n4380 GND.n4379 394
R24016 GND.n4384 GND.n4383 394
R24017 GND.n4388 GND.n4387 394
R24018 GND.n4392 GND.n4391 394
R24019 GND.n4394 GND.n4366 394
R24020 GND.n4265 GND.n1918 394
R24021 GND.n4253 GND.n1918 394
R24022 GND.n4253 GND.n1927 394
R24023 GND.n4684 GND.n1927 394
R24024 GND.n4684 GND.n1937 394
R24025 GND.n4491 GND.n1937 394
R24026 GND.n4491 GND.n1949 394
R24027 GND.n4713 GND.n1949 394
R24028 GND.n4713 GND.n1959 394
R24029 GND.n4694 GND.n1959 394
R24030 GND.n4694 GND.n1968 394
R24031 GND.n4702 GND.n1968 394
R24032 GND.n4702 GND.n1979 394
R24033 GND.n2040 GND.n1979 394
R24034 GND.n2040 GND.n1987 394
R24035 GND.n8205 GND.n1987 394
R24036 GND.n2011 GND.n2010 394
R24037 GND.n8232 GND.n2010 394
R24038 GND.n8230 GND.n8229 394
R24039 GND.n8226 GND.n8225 394
R24040 GND.n8222 GND.n8221 394
R24041 GND.n8218 GND.n8217 394
R24042 GND.n8214 GND.n8213 394
R24043 GND.n8210 GND.n8209 394
R24044 GND.n4447 GND.n1920 394
R24045 GND.n1929 GND.n1920 394
R24046 GND.n8291 GND.n1929 394
R24047 GND.n8291 GND.n1930 394
R24048 GND.n8285 GND.n1930 394
R24049 GND.n8285 GND.n1935 394
R24050 GND.n8274 GND.n1935 394
R24051 GND.n8274 GND.n1952 394
R24052 GND.n8270 GND.n1952 394
R24053 GND.n8270 GND.n1957 394
R24054 GND.n8259 GND.n1957 394
R24055 GND.n8259 GND.n1971 394
R24056 GND.n8253 GND.n1971 394
R24057 GND.n8253 GND.n1977 394
R24058 GND.n8245 GND.n1977 394
R24059 GND.n8245 GND.n1990 394
R24060 GND.n4726 GND.n1992 394
R24061 GND.n4730 GND.n4729 394
R24062 GND.n4734 GND.n4733 394
R24063 GND.n4738 GND.n4737 394
R24064 GND.n4742 GND.n4741 394
R24065 GND.n4746 GND.n4745 394
R24066 GND.n4750 GND.n4749 394
R24067 GND.n4752 GND.n2008 394
R24068 GND.n4266 GND.n1919 394
R24069 GND.n4502 GND.n1919 394
R24070 GND.n4502 GND.n1928 394
R24071 GND.n4215 GND.n1928 394
R24072 GND.n4215 GND.n1938 394
R24073 GND.n4493 GND.n1938 394
R24074 GND.n4493 GND.n1950 394
R24075 GND.n4205 GND.n1950 394
R24076 GND.n4205 GND.n1960 394
R24077 GND.n4724 GND.n1960 394
R24078 GND.n4724 GND.n1969 394
R24079 GND.n4760 GND.n1969 394
R24080 GND.n4760 GND.n1980 394
R24081 GND.n2041 GND.n1980 394
R24082 GND.n2041 GND.n1988 394
R24083 GND.n2014 GND.n1988 394
R24084 GND.n4442 GND.n4269 394
R24085 GND.n4414 GND.n4413 394
R24086 GND.n4418 GND.n4417 394
R24087 GND.n4422 GND.n4421 394
R24088 GND.n4426 GND.n4425 394
R24089 GND.n4430 GND.n4429 394
R24090 GND.n4434 GND.n4433 394
R24091 GND.n4439 GND.n4411 394
R24092 GND.n7139 GND.n6678 394
R24093 GND.n7135 GND.n6678 394
R24094 GND.n7135 GND.n7134 394
R24095 GND.n7134 GND.n6617 394
R24096 GND.n7220 GND.n6617 394
R24097 GND.n7220 GND.n6613 394
R24098 GND.n7227 GND.n6613 394
R24099 GND.n7227 GND.n2554 394
R24100 GND.n7310 GND.n2554 394
R24101 GND.n7310 GND.n2549 394
R24102 GND.n7319 GND.n2549 394
R24103 GND.n7319 GND.n2520 394
R24104 GND.n7373 GND.n2520 394
R24105 GND.n7373 GND.n2521 394
R24106 GND.n7369 GND.n2521 394
R24107 GND.n7369 GND.n2524 394
R24108 GND.n7070 GND.n6677 394
R24109 GND.n7111 GND.n7071 394
R24110 GND.n7107 GND.n7106 394
R24111 GND.n7103 GND.n7102 394
R24112 GND.n7099 GND.n7098 394
R24113 GND.n7095 GND.n7094 394
R24114 GND.n7091 GND.n7090 394
R24115 GND.n7087 GND.n7086 394
R24116 GND.n6689 GND.n6673 394
R24117 GND.n7079 GND.n6689 394
R24118 GND.n7079 GND.n6684 394
R24119 GND.n6684 GND.n6650 394
R24120 GND.n6650 GND.n6619 394
R24121 GND.n7203 GND.n6619 394
R24122 GND.n7203 GND.n6610 394
R24123 GND.n7208 GND.n6610 394
R24124 GND.n7208 GND.n2556 394
R24125 GND.n2688 GND.n2556 394
R24126 GND.n2688 GND.n2546 394
R24127 GND.n7298 GND.n2546 394
R24128 GND.n7298 GND.n2516 394
R24129 GND.n2613 GND.n2516 394
R24130 GND.n2613 GND.n2525 394
R24131 GND.n2610 GND.n2525 394
R24132 GND.n2579 GND.n2575 394
R24133 GND.n2583 GND.n2575 394
R24134 GND.n2587 GND.n2585 394
R24135 GND.n2591 GND.n2573 394
R24136 GND.n2595 GND.n2593 394
R24137 GND.n2599 GND.n2571 394
R24138 GND.n2603 GND.n2601 394
R24139 GND.n2607 GND.n2569 394
R24140 GND.n7126 GND.n6676 394
R24141 GND.n7126 GND.n6686 394
R24142 GND.n7132 GND.n6686 394
R24143 GND.n7132 GND.n6622 394
R24144 GND.n7218 GND.n6622 394
R24145 GND.n7218 GND.n6623 394
R24146 GND.n6623 GND.n6612 394
R24147 GND.n6612 GND.n2559 394
R24148 GND.n7308 GND.n2559 394
R24149 GND.n7308 GND.n2560 394
R24150 GND.n2560 GND.n2548 394
R24151 GND.n7296 GND.n2548 394
R24152 GND.n7296 GND.n2519 394
R24153 GND.n2528 GND.n2519 394
R24154 GND.n7367 GND.n2528 394
R24155 GND.n7367 GND.n2529 394
R24156 GND.n6703 GND.n6694 394
R24157 GND.n6707 GND.n6706 394
R24158 GND.n6711 GND.n6710 394
R24159 GND.n6715 GND.n6714 394
R24160 GND.n6719 GND.n6718 394
R24161 GND.n6723 GND.n6722 394
R24162 GND.n6725 GND.n6701 394
R24163 GND.n6729 GND.n6692 394
R24164 GND.n7124 GND.n6674 394
R24165 GND.n7124 GND.n6690 394
R24166 GND.n6690 GND.n6685 394
R24167 GND.n6685 GND.n6651 394
R24168 GND.n6651 GND.n6620 394
R24169 GND.n6620 GND.n6608 394
R24170 GND.n7229 GND.n6608 394
R24171 GND.n7230 GND.n7229 394
R24172 GND.n7230 GND.n2557 394
R24173 GND.n2557 GND.n2543 394
R24174 GND.n7321 GND.n2543 394
R24175 GND.n7321 GND.n2544 394
R24176 GND.n2544 GND.n2517 394
R24177 GND.n7327 GND.n2517 394
R24178 GND.n7327 GND.n2526 394
R24179 GND.n7331 GND.n2526 394
R24180 GND.n7361 GND.n7360 394
R24181 GND.n7357 GND.n7356 394
R24182 GND.n7354 GND.n2534 394
R24183 GND.n7350 GND.n7348 394
R24184 GND.n7346 GND.n2536 394
R24185 GND.n7342 GND.n7340 394
R24186 GND.n7338 GND.n2538 394
R24187 GND.n7334 GND.n7332 394
R24188 GND.n6870 GND.n6789 394
R24189 GND.n6902 GND.n6871 394
R24190 GND.n6898 GND.n6897 394
R24191 GND.n6894 GND.n6893 394
R24192 GND.n6890 GND.n6889 394
R24193 GND.n6886 GND.n6885 394
R24194 GND.n6882 GND.n6881 394
R24195 GND.n6878 GND.n6877 394
R24196 GND.n6914 GND.n6786 394
R24197 GND.n6919 GND.n6786 394
R24198 GND.n6919 GND.n6787 394
R24199 GND.n6787 GND.n6772 394
R24200 GND.n6964 GND.n6772 394
R24201 GND.n6964 GND.n6769 394
R24202 GND.n6969 GND.n6769 394
R24203 GND.n6969 GND.n6770 394
R24204 GND.n6770 GND.n6754 394
R24205 GND.n7000 GND.n6754 394
R24206 GND.n7000 GND.n6751 394
R24207 GND.n7011 GND.n6751 394
R24208 GND.n7011 GND.n6752 394
R24209 GND.n6752 GND.n6670 394
R24210 GND.n7142 GND.n6670 394
R24211 GND.n7142 GND.n6665 394
R24212 GND.n7153 GND.n6665 394
R24213 GND.n7153 GND.n6645 394
R24214 GND.n7175 GND.n6645 394
R24215 GND.n7176 GND.n7175 394
R24216 GND.n7177 GND.n7176 394
R24217 GND.n7177 GND.n6637 394
R24218 GND.n7190 GND.n6637 394
R24219 GND.n7190 GND.n2690 394
R24220 GND.n7243 GND.n2690 394
R24221 GND.n7243 GND.n2691 394
R24222 GND.n2691 GND.n2514 394
R24223 GND.n7376 GND.n2514 394
R24224 GND.n7376 GND.n2508 394
R24225 GND.n7388 GND.n2508 394
R24226 GND.n7388 GND.n2509 394
R24227 GND.n2509 GND.n2486 394
R24228 GND.n7421 GND.n2486 394
R24229 GND.n7421 GND.n2482 394
R24230 GND.n7427 GND.n2482 394
R24231 GND.n7427 GND.n2421 394
R24232 GND.n7579 GND.n2421 394
R24233 GND.n7579 GND.n2422 394
R24234 GND.n7575 GND.n2422 394
R24235 GND.n7575 GND.n2425 394
R24236 GND.n2439 GND.n2425 394
R24237 GND.n7565 GND.n2439 394
R24238 GND.n7565 GND.n2440 394
R24239 GND.n7561 GND.n2440 394
R24240 GND.n7561 GND.n2443 394
R24241 GND.n2464 GND.n2443 394
R24242 GND.n2463 GND.n2462 394
R24243 GND.n7545 GND.n2462 394
R24244 GND.n7543 GND.n7542 394
R24245 GND.n7539 GND.n7538 394
R24246 GND.n7535 GND.n7534 394
R24247 GND.n7531 GND.n7530 394
R24248 GND.n7527 GND.n7526 394
R24249 GND.n7523 GND.n7522 394
R24250 GND.n6791 GND.n6784 394
R24251 GND.n6921 GND.n6784 394
R24252 GND.n6921 GND.n6782 394
R24253 GND.n6953 GND.n6782 394
R24254 GND.n6953 GND.n6774 394
R24255 GND.n6949 GND.n6774 394
R24256 GND.n6949 GND.n6768 394
R24257 GND.n6945 GND.n6768 394
R24258 GND.n6945 GND.n6764 394
R24259 GND.n6764 GND.n6755 394
R24260 GND.n6941 GND.n6755 394
R24261 GND.n6941 GND.n6750 394
R24262 GND.n6936 GND.n6750 394
R24263 GND.n6936 GND.n6935 394
R24264 GND.n6935 GND.n6672 394
R24265 GND.n6672 GND.n6661 394
R24266 GND.n7155 GND.n6661 394
R24267 GND.n7155 GND.n6662 394
R24268 GND.n6662 GND.n6649 394
R24269 GND.n7163 GND.n6649 394
R24270 GND.n7163 GND.n6636 394
R24271 GND.n7193 GND.n6636 394
R24272 GND.n7193 GND.n7192 394
R24273 GND.n7192 GND.n2639 394
R24274 GND.n7245 GND.n2639 394
R24275 GND.n7245 GND.n2687 394
R24276 GND.n2687 GND.n2640 394
R24277 GND.n2640 GND.n2515 394
R24278 GND.n2678 GND.n2515 394
R24279 GND.n2678 GND.n2507 394
R24280 GND.n2671 GND.n2507 394
R24281 GND.n2671 GND.n2669 394
R24282 GND.n2669 GND.n2488 394
R24283 GND.n2662 GND.n2488 394
R24284 GND.n2662 GND.n2480 394
R24285 GND.n2658 GND.n2480 394
R24286 GND.n2658 GND.n2419 394
R24287 GND.n2654 GND.n2419 394
R24288 GND.n2654 GND.n2427 394
R24289 GND.n2650 GND.n2427 394
R24290 GND.n2650 GND.n2649 394
R24291 GND.n2649 GND.n2437 394
R24292 GND.n7513 GND.n2437 394
R24293 GND.n7513 GND.n2444 394
R24294 GND.n7517 GND.n2444 394
R24295 GND.n7518 GND.n7517 394
R24296 GND.n6845 GND.n6797 394
R24297 GND.n6906 GND.n6797 394
R24298 GND.n6906 GND.n6794 394
R24299 GND.n6911 GND.n6794 394
R24300 GND.n6911 GND.n6795 394
R24301 GND.n6795 GND.n6779 394
R24302 GND.n6956 GND.n6779 394
R24303 GND.n6956 GND.n6776 394
R24304 GND.n6961 GND.n6776 394
R24305 GND.n6961 GND.n6777 394
R24306 GND.n6777 GND.n6761 394
R24307 GND.n6986 GND.n6761 394
R24308 GND.n6986 GND.n6758 394
R24309 GND.n6997 GND.n6758 394
R24310 GND.n6997 GND.n6759 394
R24311 GND.n6759 GND.n6732 394
R24312 GND.n7061 GND.n6732 394
R24313 GND.n7061 GND.n6733 394
R24314 GND.n7054 GND.n6733 394
R24315 GND.n7054 GND.n7053 394
R24316 GND.n7053 GND.n7045 394
R24317 GND.n7045 GND.n6653 394
R24318 GND.n7171 GND.n6653 394
R24319 GND.n7171 GND.n6631 394
R24320 GND.n7200 GND.n6631 394
R24321 GND.n7200 GND.n2632 394
R24322 GND.n7252 GND.n2632 394
R24323 GND.n7252 GND.n2624 394
R24324 GND.n7278 GND.n2624 394
R24325 GND.n7278 GND.n2619 394
R24326 GND.n7287 GND.n2619 394
R24327 GND.n7287 GND.n2504 394
R24328 GND.n7391 GND.n2504 394
R24329 GND.n7391 GND.n2497 394
R24330 GND.n7403 GND.n2497 394
R24331 GND.n7403 GND.n2499 394
R24332 GND.n2499 GND.n2477 394
R24333 GND.n7430 GND.n2477 394
R24334 GND.n7430 GND.n2472 394
R24335 GND.n7437 GND.n2472 394
R24336 GND.n7437 GND.n2473 394
R24337 GND.n2473 GND.n2430 394
R24338 GND.n7572 GND.n2430 394
R24339 GND.n7572 GND.n2431 394
R24340 GND.n7568 GND.n2431 394
R24341 GND.n7568 GND.n2434 394
R24342 GND.n2447 GND.n2434 394
R24343 GND.n7558 GND.n2447 394
R24344 GND.n7558 GND.n2448 394
R24345 GND.n7554 GND.n2448 394
R24346 GND.n7554 GND.n2451 394
R24347 GND.n7499 GND.n2451 394
R24348 GND.n7499 GND.n7452 394
R24349 GND.n7492 GND.n7454 394
R24350 GND.n7492 GND.n7462 394
R24351 GND.n7488 GND.n7487 394
R24352 GND.n7484 GND.n7483 394
R24353 GND.n7480 GND.n7479 394
R24354 GND.n7476 GND.n7475 394
R24355 GND.n7472 GND.n7471 394
R24356 GND.n7468 GND.n7467 394
R24357 GND.n6847 GND.n6798 394
R24358 GND.n6862 GND.n6798 394
R24359 GND.n6862 GND.n6799 394
R24360 GND.n6799 GND.n6792 394
R24361 GND.n6857 GND.n6792 394
R24362 GND.n6857 GND.n6856 394
R24363 GND.n6856 GND.n6781 394
R24364 GND.n6851 GND.n6781 394
R24365 GND.n6851 GND.n6775 394
R24366 GND.n6775 GND.n6766 394
R24367 GND.n6972 GND.n6766 394
R24368 GND.n6972 GND.n6763 394
R24369 GND.n6981 GND.n6763 394
R24370 GND.n6981 GND.n6756 394
R24371 GND.n6756 GND.n6748 394
R24372 GND.n7014 GND.n6748 394
R24373 GND.n7014 GND.n6731 394
R24374 GND.n7021 GND.n6731 394
R24375 GND.n7022 GND.n7021 394
R24376 GND.n7022 GND.n6739 394
R24377 GND.n7043 GND.n6739 394
R24378 GND.n7043 GND.n6740 394
R24379 GND.n6740 GND.n6652 394
R24380 GND.n7034 GND.n6652 394
R24381 GND.n7034 GND.n6630 394
R24382 GND.n6630 GND.n2631 394
R24383 GND.n7254 GND.n2631 394
R24384 GND.n7254 GND.n2625 394
R24385 GND.n7276 GND.n2625 394
R24386 GND.n7276 GND.n2626 394
R24387 GND.n2626 GND.n2618 394
R24388 GND.n7267 GND.n2618 394
R24389 GND.n7267 GND.n2506 394
R24390 GND.n2506 GND.n2494 394
R24391 GND.n7405 GND.n2494 394
R24392 GND.n7405 GND.n2489 394
R24393 GND.n7418 GND.n2489 394
R24394 GND.n7418 GND.n2479 394
R24395 GND.n2479 GND.n2470 394
R24396 GND.n7439 GND.n2470 394
R24397 GND.n7440 GND.n7439 394
R24398 GND.n7441 GND.n7440 394
R24399 GND.n7441 GND.n2428 394
R24400 GND.n7445 GND.n2428 394
R24401 GND.n7445 GND.n2436 394
R24402 GND.n2468 GND.n2436 394
R24403 GND.n7510 GND.n2468 394
R24404 GND.n7510 GND.n2445 394
R24405 GND.n7506 GND.n2445 394
R24406 GND.n7506 GND.n2453 394
R24407 GND.n7502 GND.n2453 394
R24408 GND.n7502 GND.n7501 394
R24409 GND.n7501 GND.n7450 394
R24410 GND.n6841 GND.n6839 394
R24411 GND.n6837 GND.n6806 394
R24412 GND.n6833 GND.n6831 394
R24413 GND.n6829 GND.n6808 394
R24414 GND.n6825 GND.n6823 394
R24415 GND.n6821 GND.n6810 394
R24416 GND.n6817 GND.n6815 394
R24417 GND.n6813 GND.n6801 394
R24418 GND.n9791 GND.n55 389.272
R24419 GND.n9787 GND.n55 389.272
R24420 GND.n8426 GND.n8425 389.272
R24421 GND.n8425 GND.n8424 389.272
R24422 GND.n5983 GND.n5982 379.416
R24423 GND.t430 GND.t47 365.217
R24424 GND.t47 GND.t149 365.217
R24425 GND.t359 GND.t135 349.67
R24426 GND.t361 GND.t131 349.67
R24427 GND.t94 GND.t141 349.67
R24428 GND.t88 GND.t144 349.67
R24429 GND.t96 GND.t373 349.67
R24430 GND.t278 GND.t374 349.67
R24431 GND.n7747 GND.n2274 349.257
R24432 GND.t149 GND.t339 345.717
R24433 GND.t395 GND.n2892 335.099
R24434 GND.n7718 GND.n2299 325.753
R24435 GND.n7712 GND.n7711 325.753
R24436 GND.n9460 GND.n9459 325.753
R24437 GND.n9449 GND.n9448 325.753
R24438 GND.n7694 GND.n2310 320
R24439 GND.n7700 GND.n2310 320
R24440 GND.n9822 GND.n12 320
R24441 GND.n2117 GND.n12 320
R24442 GND.n9783 GND.t152 316.002
R24443 GND.n9794 GND.t357 312.788
R24444 GND.n9795 GND.n9794 306.404
R24445 GND.t377 GND.n7683 290.356
R24446 GND.n9786 GND.n9785 289.163
R24447 GND.n2915 GND.t46 286.433
R24448 GND.n2971 GND.t15 285.481
R24449 GND.n3095 GND.t384 285.481
R24450 GND.n3107 GND.t386 282.327
R24451 GND.n8431 GND.n25 277.108
R24452 GND.t133 GND.t359 262.252
R24453 GND.t135 GND.t361 262.252
R24454 GND.t131 GND.t358 262.252
R24455 GND.t90 GND.t145 262.252
R24456 GND.t92 GND.n2998 262.252
R24457 GND.t141 GND.t92 262.252
R24458 GND.t144 GND.t94 262.252
R24459 GND.t148 GND.t88 262.252
R24460 GND.t373 GND.t84 262.252
R24461 GND.t374 GND.t96 262.252
R24462 GND.t371 GND.t278 262.252
R24463 GND.n9820 GND.n9819 260.283
R24464 GND.n7703 GND.n7702 260.283
R24465 GND.n7717 GND.n2298 257.236
R24466 GND.n7707 GND.n7706 257.236
R24467 GND.n9455 GND.n9454 257.236
R24468 GND.n9444 GND.n9443 257.236
R24469 GND.n7700 GND.n7699 255.087
R24470 GND.n9823 GND.n9822 255.087
R24471 GND.n7695 GND.n7694 252.827
R24472 GND.n2117 GND.n2116 252.827
R24473 GND.n8428 GND.n1803 251.516
R24474 GND.n7743 GND.n7742 247.38
R24475 GND.n9812 GND.n21 247.38
R24476 GND.t153 GND.t81 244.084
R24477 GND.n2895 GND.t335 242.66
R24478 GND.n9680 GND.t124 224.244
R24479 GND.n7689 GND.t377 223.273
R24480 GND.n9345 GND.n9344 218.815
R24481 GND.n9345 GND.n302 218.815
R24482 GND.n9345 GND.n303 218.815
R24483 GND.n9345 GND.n304 218.815
R24484 GND.n9345 GND.n305 218.815
R24485 GND.n9345 GND.n306 218.815
R24486 GND.n9345 GND.n307 218.815
R24487 GND.n9345 GND.n308 218.815
R24488 GND.n856 GND.n512 218.815
R24489 GND.n856 GND.n511 218.815
R24490 GND.n856 GND.n510 218.815
R24491 GND.n856 GND.n509 218.815
R24492 GND.n856 GND.n508 218.815
R24493 GND.n856 GND.n507 218.815
R24494 GND.n856 GND.n506 218.815
R24495 GND.n856 GND.n505 218.815
R24496 GND.n856 GND.n520 218.815
R24497 GND.n856 GND.n519 218.815
R24498 GND.n856 GND.n518 218.815
R24499 GND.n856 GND.n517 218.815
R24500 GND.n856 GND.n516 218.815
R24501 GND.n856 GND.n515 218.815
R24502 GND.n856 GND.n514 218.815
R24503 GND.n856 GND.n513 218.815
R24504 GND.n9346 GND.n9345 218.815
R24505 GND.n9345 GND.n309 218.815
R24506 GND.n9345 GND.n310 218.815
R24507 GND.n9345 GND.n311 218.815
R24508 GND.n9345 GND.n312 218.815
R24509 GND.n9345 GND.n313 218.815
R24510 GND.n9345 GND.n314 218.815
R24511 GND.n9345 GND.n315 218.815
R24512 GND.n8239 GND.n8238 218.815
R24513 GND.n8239 GND.n1994 218.815
R24514 GND.n8239 GND.n1995 218.815
R24515 GND.n8239 GND.n1996 218.815
R24516 GND.n8239 GND.n1997 218.815
R24517 GND.n8239 GND.n1998 218.815
R24518 GND.n8239 GND.n1999 218.815
R24519 GND.n8239 GND.n2000 218.815
R24520 GND.n4440 GND.n4403 218.815
R24521 GND.n4440 GND.n4365 218.815
R24522 GND.n4440 GND.n4364 218.815
R24523 GND.n4440 GND.n4363 218.815
R24524 GND.n4440 GND.n4362 218.815
R24525 GND.n4440 GND.n4361 218.815
R24526 GND.n4440 GND.n4360 218.815
R24527 GND.n4440 GND.n4359 218.815
R24528 GND.n4440 GND.n4410 218.815
R24529 GND.n4440 GND.n4409 218.815
R24530 GND.n4440 GND.n4408 218.815
R24531 GND.n4440 GND.n4407 218.815
R24532 GND.n4440 GND.n4406 218.815
R24533 GND.n4440 GND.n4405 218.815
R24534 GND.n4440 GND.n4404 218.815
R24535 GND.n4441 GND.n4440 218.815
R24536 GND.n8240 GND.n8239 218.815
R24537 GND.n8239 GND.n2001 218.815
R24538 GND.n8239 GND.n2002 218.815
R24539 GND.n8239 GND.n2003 218.815
R24540 GND.n8239 GND.n2004 218.815
R24541 GND.n8239 GND.n2005 218.815
R24542 GND.n8239 GND.n2006 218.815
R24543 GND.n8239 GND.n2007 218.815
R24544 GND.n3563 GND.n3399 218.815
R24545 GND.n3561 GND.n3399 218.815
R24546 GND.n3555 GND.n3399 218.815
R24547 GND.n3553 GND.n3399 218.815
R24548 GND.n3547 GND.n3399 218.815
R24549 GND.n3545 GND.n3399 218.815
R24550 GND.n3539 GND.n3399 218.815
R24551 GND.n3537 GND.n3399 218.815
R24552 GND.n3531 GND.n3399 218.815
R24553 GND.n3696 GND.n3134 218.815
R24554 GND.n3696 GND.n3133 218.815
R24555 GND.n3696 GND.n3132 218.815
R24556 GND.n3696 GND.n3131 218.815
R24557 GND.n3696 GND.n3130 218.815
R24558 GND.n3696 GND.n3129 218.815
R24559 GND.n3696 GND.n3128 218.815
R24560 GND.n3696 GND.n3127 218.815
R24561 GND.n3696 GND.n3126 218.815
R24562 GND.n8728 GND.n1722 218.815
R24563 GND.n8728 GND.n1661 218.815
R24564 GND.n8728 GND.n1660 218.815
R24565 GND.n8728 GND.n1659 218.815
R24566 GND.n8728 GND.n1658 218.815
R24567 GND.n8728 GND.n1657 218.815
R24568 GND.n8728 GND.n1656 218.815
R24569 GND.n8728 GND.n1655 218.815
R24570 GND.n8728 GND.n1654 218.815
R24571 GND.n8558 GND.n8499 218.815
R24572 GND.n8565 GND.n8499 218.815
R24573 GND.n8509 GND.n8499 218.815
R24574 GND.n8572 GND.n8499 218.815
R24575 GND.n8506 GND.n8499 218.815
R24576 GND.n8579 GND.n8499 218.815
R24577 GND.n8503 GND.n8499 218.815
R24578 GND.n8586 GND.n8499 218.815
R24579 GND.n8589 GND.n8499 218.815
R24580 GND.n3399 GND.n3398 218.815
R24581 GND.n3399 GND.n3337 218.815
R24582 GND.n3399 GND.n3338 218.815
R24583 GND.n3399 GND.n3339 218.815
R24584 GND.n3399 GND.n3340 218.815
R24585 GND.n3399 GND.n3341 218.815
R24586 GND.n3399 GND.n3342 218.815
R24587 GND.n3399 GND.n3343 218.815
R24588 GND.n3696 GND.n3125 218.815
R24589 GND.n3696 GND.n3124 218.815
R24590 GND.n3696 GND.n3123 218.815
R24591 GND.n3696 GND.n3122 218.815
R24592 GND.n3696 GND.n3121 218.815
R24593 GND.n3696 GND.n3120 218.815
R24594 GND.n3696 GND.n3119 218.815
R24595 GND.n3696 GND.n3118 218.815
R24596 GND.n3696 GND.n3117 218.815
R24597 GND.n8729 GND.n8728 218.815
R24598 GND.n8728 GND.n1063 218.815
R24599 GND.n8728 GND.n1064 218.815
R24600 GND.n8728 GND.n1065 218.815
R24601 GND.n8728 GND.n1066 218.815
R24602 GND.n8728 GND.n1067 218.815
R24603 GND.n8728 GND.n1068 218.815
R24604 GND.n8728 GND.n1069 218.815
R24605 GND.n8499 GND.n8498 218.815
R24606 GND.n8499 GND.n8439 218.815
R24607 GND.n8499 GND.n8438 218.815
R24608 GND.n8499 GND.n8437 218.815
R24609 GND.n8499 GND.n8436 218.815
R24610 GND.n8499 GND.n8435 218.815
R24611 GND.n8499 GND.n8434 218.815
R24612 GND.n8499 GND.n8433 218.815
R24613 GND.n8499 GND.n8432 218.815
R24614 GND.n1520 GND.n51 218.815
R24615 GND.n1518 GND.n51 218.815
R24616 GND.n1512 GND.n51 218.815
R24617 GND.n1510 GND.n51 218.815
R24618 GND.n1504 GND.n51 218.815
R24619 GND.n1502 GND.n51 218.815
R24620 GND.n1496 GND.n51 218.815
R24621 GND.n1494 GND.n51 218.815
R24622 GND.n1488 GND.n51 218.815
R24623 GND.n1653 GND.n1088 218.815
R24624 GND.n1653 GND.n1087 218.815
R24625 GND.n1653 GND.n1086 218.815
R24626 GND.n1653 GND.n1085 218.815
R24627 GND.n1653 GND.n1084 218.815
R24628 GND.n1653 GND.n1083 218.815
R24629 GND.n1653 GND.n1082 218.815
R24630 GND.n1653 GND.n1081 218.815
R24631 GND.n1653 GND.n1080 218.815
R24632 GND.n1318 GND.n51 218.815
R24633 GND.n1321 GND.n51 218.815
R24634 GND.n1327 GND.n51 218.815
R24635 GND.n1329 GND.n51 218.815
R24636 GND.n1335 GND.n51 218.815
R24637 GND.n1337 GND.n51 218.815
R24638 GND.n1343 GND.n51 218.815
R24639 GND.n1346 GND.n51 218.815
R24640 GND.n1653 GND.n1079 218.815
R24641 GND.n1653 GND.n1078 218.815
R24642 GND.n1653 GND.n1077 218.815
R24643 GND.n1653 GND.n1076 218.815
R24644 GND.n1653 GND.n1075 218.815
R24645 GND.n1653 GND.n1074 218.815
R24646 GND.n1653 GND.n1073 218.815
R24647 GND.n1653 GND.n1072 218.815
R24648 GND.n1653 GND.n1071 218.815
R24649 GND.n9199 GND.n50 218.815
R24650 GND.n9141 GND.n50 218.815
R24651 GND.n9192 GND.n50 218.815
R24652 GND.n9186 GND.n50 218.815
R24653 GND.n9184 GND.n50 218.815
R24654 GND.n9178 GND.n50 218.815
R24655 GND.n9176 GND.n50 218.815
R24656 GND.n9170 GND.n50 218.815
R24657 GND.n9135 GND.n9134 218.815
R24658 GND.n9135 GND.n418 218.815
R24659 GND.n9135 GND.n419 218.815
R24660 GND.n9135 GND.n420 218.815
R24661 GND.n9135 GND.n421 218.815
R24662 GND.n9135 GND.n422 218.815
R24663 GND.n9135 GND.n423 218.815
R24664 GND.n9135 GND.n424 218.815
R24665 GND.n9680 GND.n9679 218.815
R24666 GND.n9680 GND.n9622 218.815
R24667 GND.n9680 GND.n9623 218.815
R24668 GND.n9680 GND.n9624 218.815
R24669 GND.n9680 GND.n9625 218.815
R24670 GND.n9680 GND.n9626 218.815
R24671 GND.n9680 GND.n9627 218.815
R24672 GND.n9680 GND.n9628 218.815
R24673 GND.n9505 GND.n9465 218.815
R24674 GND.n9505 GND.n9466 218.815
R24675 GND.n9505 GND.n9467 218.815
R24676 GND.n9505 GND.n9468 218.815
R24677 GND.n9505 GND.n9469 218.815
R24678 GND.n9505 GND.n9470 218.815
R24679 GND.n9505 GND.n9471 218.815
R24680 GND.n9505 GND.n9504 218.815
R24681 GND.n9689 GND.n9688 218.815
R24682 GND.n9688 GND.n129 218.815
R24683 GND.n9545 GND.n9541 218.815
R24684 GND.n9551 GND.n9541 218.815
R24685 GND.n9554 GND.n9541 218.815
R24686 GND.n9734 GND.n9733 218.815
R24687 GND.n9734 GND.n92 218.815
R24688 GND.n9734 GND.n93 218.815
R24689 GND.n9734 GND.n94 218.815
R24690 GND.n159 GND.n149 218.815
R24691 GND.n9596 GND.n149 218.815
R24692 GND.n149 GND.n136 218.815
R24693 GND.n149 GND.n148 218.815
R24694 GND.n149 GND.n138 218.815
R24695 GND.n8093 GND.n8032 218.815
R24696 GND.n8035 GND.n8032 218.815
R24697 GND.n8086 GND.n8032 218.815
R24698 GND.n8080 GND.n8032 218.815
R24699 GND.n8078 GND.n8032 218.815
R24700 GND.n8072 GND.n8032 218.815
R24701 GND.n8070 GND.n8032 218.815
R24702 GND.n8064 GND.n8032 218.815
R24703 GND.n4569 GND.n2108 218.815
R24704 GND.n4575 GND.n2108 218.815
R24705 GND.n4577 GND.n2108 218.815
R24706 GND.n4583 GND.n2108 218.815
R24707 GND.n4585 GND.n2108 218.815
R24708 GND.n4591 GND.n2108 218.815
R24709 GND.n4593 GND.n2108 218.815
R24710 GND.n4599 GND.n2108 218.815
R24711 GND.n616 GND.n615 218.815
R24712 GND.n615 GND.n578 218.815
R24713 GND.n615 GND.n579 218.815
R24714 GND.n615 GND.n580 218.815
R24715 GND.n615 GND.n581 218.815
R24716 GND.n615 GND.n582 218.815
R24717 GND.n615 GND.n583 218.815
R24718 GND.n615 GND.n584 218.815
R24719 GND.n678 GND.n640 218.815
R24720 GND.n678 GND.n641 218.815
R24721 GND.n678 GND.n642 218.815
R24722 GND.n678 GND.n643 218.815
R24723 GND.n678 GND.n644 218.815
R24724 GND.n678 GND.n645 218.815
R24725 GND.n678 GND.n646 218.815
R24726 GND.n678 GND.n677 218.815
R24727 GND.n8029 GND.n8028 218.815
R24728 GND.n8029 GND.n2120 218.815
R24729 GND.n8029 GND.n2121 218.815
R24730 GND.n8029 GND.n2122 218.815
R24731 GND.n8029 GND.n2123 218.815
R24732 GND.n8029 GND.n2124 218.815
R24733 GND.n8029 GND.n2125 218.815
R24734 GND.n8029 GND.n2126 218.815
R24735 GND.n7789 GND.n7749 218.815
R24736 GND.n7789 GND.n7750 218.815
R24737 GND.n7789 GND.n7751 218.815
R24738 GND.n7789 GND.n7752 218.815
R24739 GND.n7789 GND.n7753 218.815
R24740 GND.n7789 GND.n7754 218.815
R24741 GND.n7789 GND.n7755 218.815
R24742 GND.n7789 GND.n7756 218.815
R24743 GND.n7986 GND.n7985 218.815
R24744 GND.n7986 GND.n2139 218.815
R24745 GND.n7823 GND.n7818 218.815
R24746 GND.n7829 GND.n7818 218.815
R24747 GND.n7832 GND.n7818 218.815
R24748 GND.n7955 GND.n7954 218.815
R24749 GND.n7955 GND.n2176 218.815
R24750 GND.n7955 GND.n2177 218.815
R24751 GND.n7955 GND.n2178 218.815
R24752 GND.n7865 GND.n7864 218.815
R24753 GND.n7865 GND.n2225 218.815
R24754 GND.n7865 GND.n2224 218.815
R24755 GND.n7865 GND.n2223 218.815
R24756 GND.n7865 GND.n2222 218.815
R24757 GND.n7362 GND.n2487 218.815
R24758 GND.n2532 GND.n2487 218.815
R24759 GND.n7355 GND.n2487 218.815
R24760 GND.n7349 GND.n2487 218.815
R24761 GND.n7347 GND.n2487 218.815
R24762 GND.n7341 GND.n2487 218.815
R24763 GND.n7339 GND.n2487 218.815
R24764 GND.n7333 GND.n2487 218.815
R24765 GND.n7114 GND.n7113 218.815
R24766 GND.n7113 GND.n6730 218.815
R24767 GND.n7113 GND.n6700 218.815
R24768 GND.n7113 GND.n6699 218.815
R24769 GND.n7113 GND.n6698 218.815
R24770 GND.n7113 GND.n6697 218.815
R24771 GND.n7113 GND.n6696 218.815
R24772 GND.n7113 GND.n6695 218.815
R24773 GND.n2578 GND.n2487 218.815
R24774 GND.n2584 GND.n2487 218.815
R24775 GND.n2586 GND.n2487 218.815
R24776 GND.n2592 GND.n2487 218.815
R24777 GND.n2594 GND.n2487 218.815
R24778 GND.n2600 GND.n2487 218.815
R24779 GND.n2602 GND.n2487 218.815
R24780 GND.n2608 GND.n2487 218.815
R24781 GND.n7113 GND.n7063 218.815
R24782 GND.n7113 GND.n7064 218.815
R24783 GND.n7113 GND.n7065 218.815
R24784 GND.n7113 GND.n7066 218.815
R24785 GND.n7113 GND.n7067 218.815
R24786 GND.n7113 GND.n7068 218.815
R24787 GND.n7113 GND.n7069 218.815
R24788 GND.n7113 GND.n7112 218.815
R24789 GND.n7552 GND.n7551 218.815
R24790 GND.n7552 GND.n2454 218.815
R24791 GND.n7552 GND.n2455 218.815
R24792 GND.n7552 GND.n2456 218.815
R24793 GND.n7552 GND.n2457 218.815
R24794 GND.n7552 GND.n2458 218.815
R24795 GND.n7552 GND.n2459 218.815
R24796 GND.n7552 GND.n2460 218.815
R24797 GND.n8396 GND.n1817 218.815
R24798 GND.n8396 GND.n1818 218.815
R24799 GND.n8396 GND.n1819 218.815
R24800 GND.n8396 GND.n1820 218.815
R24801 GND.n8396 GND.n1821 218.815
R24802 GND.n8396 GND.n1822 218.815
R24803 GND.n8396 GND.n1823 218.815
R24804 GND.n8396 GND.n1824 218.815
R24805 GND.n4313 GND.n1835 218.815
R24806 GND.n4277 GND.n1835 218.815
R24807 GND.n4306 GND.n1835 218.815
R24808 GND.n4300 GND.n1835 218.815
R24809 GND.n4298 GND.n1835 218.815
R24810 GND.n4292 GND.n1835 218.815
R24811 GND.n4290 GND.n1835 218.815
R24812 GND.n4284 GND.n1835 218.815
R24813 GND.n5729 GND.n4983 218.815
R24814 GND.n5729 GND.n4984 218.815
R24815 GND.n5729 GND.n4985 218.815
R24816 GND.n5729 GND.n4986 218.815
R24817 GND.n5729 GND.n4987 218.815
R24818 GND.n5729 GND.n4988 218.815
R24819 GND.n5729 GND.n4989 218.815
R24820 GND.n5729 GND.n4990 218.815
R24821 GND.n5729 GND.n4991 218.815
R24822 GND.n5729 GND.n4992 218.815
R24823 GND.n5729 GND.n4993 218.815
R24824 GND.n5729 GND.n4994 218.815
R24825 GND.n5729 GND.n4995 218.815
R24826 GND.n5729 GND.n4996 218.815
R24827 GND.n5729 GND.n4997 218.815
R24828 GND.n5729 GND.n4998 218.815
R24829 GND.n5729 GND.n4999 218.815
R24830 GND.n5729 GND.n5000 218.815
R24831 GND.n5729 GND.n5001 218.815
R24832 GND.n5729 GND.n5002 218.815
R24833 GND.n5729 GND.n5728 218.815
R24834 GND.n5098 GND.n3837 218.815
R24835 GND.n5104 GND.n3837 218.815
R24836 GND.n5106 GND.n3837 218.815
R24837 GND.n5112 GND.n3837 218.815
R24838 GND.n5114 GND.n3837 218.815
R24839 GND.n5120 GND.n3837 218.815
R24840 GND.n5122 GND.n3837 218.815
R24841 GND.n5128 GND.n3837 218.815
R24842 GND.n5130 GND.n3837 218.815
R24843 GND.n5142 GND.n3837 218.815
R24844 GND.n5144 GND.n3837 218.815
R24845 GND.n5154 GND.n3837 218.815
R24846 GND.n5157 GND.n3837 218.815
R24847 GND.n5038 GND.n3837 218.815
R24848 GND.n5343 GND.n3837 218.815
R24849 GND.n5345 GND.n3837 218.815
R24850 GND.n5351 GND.n3837 218.815
R24851 GND.n5353 GND.n3837 218.815
R24852 GND.n5359 GND.n3837 218.815
R24853 GND.n5361 GND.n3837 218.815
R24854 GND.n5367 GND.n3837 218.815
R24855 GND.n4982 GND.n3906 218.815
R24856 GND.n4982 GND.n3907 218.815
R24857 GND.n4982 GND.n3908 218.815
R24858 GND.n4982 GND.n3909 218.815
R24859 GND.n4982 GND.n3910 218.815
R24860 GND.n4982 GND.n3911 218.815
R24861 GND.n4982 GND.n3912 218.815
R24862 GND.n4982 GND.n3913 218.815
R24863 GND.n4982 GND.n3914 218.815
R24864 GND.n4982 GND.n3915 218.815
R24865 GND.n4982 GND.n3916 218.815
R24866 GND.n4982 GND.n3917 218.815
R24867 GND.n4982 GND.n3918 218.815
R24868 GND.n4982 GND.n3919 218.815
R24869 GND.n4982 GND.n3920 218.815
R24870 GND.n4982 GND.n3921 218.815
R24871 GND.n4982 GND.n3922 218.815
R24872 GND.n4982 GND.n3923 218.815
R24873 GND.n4982 GND.n3924 218.815
R24874 GND.n4982 GND.n3925 218.815
R24875 GND.n4982 GND.n3926 218.815
R24876 GND.n5809 GND.n5808 218.815
R24877 GND.n5809 GND.n3818 218.815
R24878 GND.n5809 GND.n3819 218.815
R24879 GND.n5809 GND.n3820 218.815
R24880 GND.n5809 GND.n3821 218.815
R24881 GND.n5809 GND.n3822 218.815
R24882 GND.n5809 GND.n3823 218.815
R24883 GND.n5810 GND.n5809 218.815
R24884 GND.n5809 GND.n3824 218.815
R24885 GND.n5809 GND.n3825 218.815
R24886 GND.n5809 GND.n3826 218.815
R24887 GND.n5809 GND.n3827 218.815
R24888 GND.n5809 GND.n3828 218.815
R24889 GND.n5809 GND.n3829 218.815
R24890 GND.n5809 GND.n3830 218.815
R24891 GND.n5809 GND.n3831 218.815
R24892 GND.n5809 GND.n3832 218.815
R24893 GND.n5809 GND.n3833 218.815
R24894 GND.n5809 GND.n3834 218.815
R24895 GND.n5809 GND.n3835 218.815
R24896 GND.n5809 GND.n3836 218.815
R24897 GND.n5312 GND.n3789 218.815
R24898 GND.n5172 GND.n3789 218.815
R24899 GND.n5319 GND.n3789 218.815
R24900 GND.n5169 GND.n3789 218.815
R24901 GND.n5326 GND.n3789 218.815
R24902 GND.n5166 GND.n3789 218.815
R24903 GND.n5333 GND.n3789 218.815
R24904 GND.n5336 GND.n3789 218.815
R24905 GND.n5161 GND.n3789 218.815
R24906 GND.n5150 GND.n3789 218.815
R24907 GND.n5148 GND.n3789 218.815
R24908 GND.n5138 GND.n3789 218.815
R24909 GND.n5136 GND.n3789 218.815
R24910 GND.n5084 GND.n3789 218.815
R24911 GND.n5082 GND.n3789 218.815
R24912 GND.n5076 GND.n3789 218.815
R24913 GND.n5074 GND.n3789 218.815
R24914 GND.n5068 GND.n3789 218.815
R24915 GND.n5066 GND.n3789 218.815
R24916 GND.n5060 GND.n3789 218.815
R24917 GND.n5058 GND.n3789 218.815
R24918 GND.n5194 GND.n3717 218.815
R24919 GND.n5200 GND.n3717 218.815
R24920 GND.n5202 GND.n3717 218.815
R24921 GND.n5208 GND.n3717 218.815
R24922 GND.n5210 GND.n3717 218.815
R24923 GND.n5216 GND.n3717 218.815
R24924 GND.n5218 GND.n3717 218.815
R24925 GND.n5224 GND.n3717 218.815
R24926 GND.n5226 GND.n3717 218.815
R24927 GND.n5232 GND.n3717 218.815
R24928 GND.n5234 GND.n3717 218.815
R24929 GND.n5240 GND.n3717 218.815
R24930 GND.n5242 GND.n3717 218.815
R24931 GND.n5248 GND.n3717 218.815
R24932 GND.n5250 GND.n3717 218.815
R24933 GND.n5256 GND.n3717 218.815
R24934 GND.n5258 GND.n3717 218.815
R24935 GND.n5264 GND.n3717 218.815
R24936 GND.n5266 GND.n3717 218.815
R24937 GND.n5272 GND.n3717 218.815
R24938 GND.n5275 GND.n3717 218.815
R24939 GND.n5845 GND.n3790 218.815
R24940 GND.n5845 GND.n3791 218.815
R24941 GND.n5845 GND.n3792 218.815
R24942 GND.n5845 GND.n3793 218.815
R24943 GND.n5845 GND.n3794 218.815
R24944 GND.n5845 GND.n3795 218.815
R24945 GND.n5845 GND.n3796 218.815
R24946 GND.n5845 GND.n3797 218.815
R24947 GND.n5845 GND.n3798 218.815
R24948 GND.n5845 GND.n3799 218.815
R24949 GND.n5845 GND.n3800 218.815
R24950 GND.n5845 GND.n3801 218.815
R24951 GND.n5845 GND.n3802 218.815
R24952 GND.n5845 GND.n3803 218.815
R24953 GND.n5845 GND.n3804 218.815
R24954 GND.n5845 GND.n3805 218.815
R24955 GND.n5845 GND.n3806 218.815
R24956 GND.n5845 GND.n3807 218.815
R24957 GND.n5845 GND.n3808 218.815
R24958 GND.n5845 GND.n3809 218.815
R24959 GND.n5845 GND.n3810 218.815
R24960 GND.n5982 GND.n5981 218.815
R24961 GND.n5982 GND.n3697 218.815
R24962 GND.n5982 GND.n3698 218.815
R24963 GND.n5982 GND.n3699 218.815
R24964 GND.n5982 GND.n3700 218.815
R24965 GND.n5982 GND.n3701 218.815
R24966 GND.n5982 GND.n3702 218.815
R24967 GND.n5982 GND.n3703 218.815
R24968 GND.n5982 GND.n3704 218.815
R24969 GND.n5982 GND.n3705 218.815
R24970 GND.n5982 GND.n3706 218.815
R24971 GND.n5982 GND.n3707 218.815
R24972 GND.n5982 GND.n3708 218.815
R24973 GND.n5982 GND.n3709 218.815
R24974 GND.n5982 GND.n3710 218.815
R24975 GND.n5982 GND.n3711 218.815
R24976 GND.n5982 GND.n3712 218.815
R24977 GND.n5982 GND.n3713 218.815
R24978 GND.n5982 GND.n3714 218.815
R24979 GND.n5982 GND.n3715 218.815
R24980 GND.n5982 GND.n3716 218.815
R24981 GND.n2733 GND.n2720 218.815
R24982 GND.n6395 GND.n2720 218.815
R24983 GND.n2730 GND.n2720 218.815
R24984 GND.n6402 GND.n2720 218.815
R24985 GND.n2727 GND.n2720 218.815
R24986 GND.n6409 GND.n2720 218.815
R24987 GND.n2724 GND.n2720 218.815
R24988 GND.n6416 GND.n2720 218.815
R24989 GND.n6419 GND.n2720 218.815
R24990 GND.n6335 GND.n2720 218.815
R24991 GND.n6343 GND.n2720 218.815
R24992 GND.n6346 GND.n2720 218.815
R24993 GND.n6332 GND.n2720 218.815
R24994 GND.n6358 GND.n2720 218.815
R24995 GND.n6325 GND.n2720 218.815
R24996 GND.n6365 GND.n2720 218.815
R24997 GND.n6322 GND.n2720 218.815
R24998 GND.n6372 GND.n2720 218.815
R24999 GND.n6319 GND.n2720 218.815
R25000 GND.n6379 GND.n2720 218.815
R25001 GND.n6382 GND.n2720 218.815
R25002 GND.n6261 GND.n6260 218.815
R25003 GND.n6260 GND.n2772 218.815
R25004 GND.n6260 GND.n2773 218.815
R25005 GND.n6260 GND.n2774 218.815
R25006 GND.n6260 GND.n2775 218.815
R25007 GND.n6260 GND.n2776 218.815
R25008 GND.n6260 GND.n2777 218.815
R25009 GND.n6260 GND.n2778 218.815
R25010 GND.n6260 GND.n2779 218.815
R25011 GND.n6260 GND.n2780 218.815
R25012 GND.n6260 GND.n2781 218.815
R25013 GND.n6260 GND.n2782 218.815
R25014 GND.n6260 GND.n2783 218.815
R25015 GND.n6260 GND.n2784 218.815
R25016 GND.n6260 GND.n2785 218.815
R25017 GND.n6260 GND.n2786 218.815
R25018 GND.n6260 GND.n2787 218.815
R25019 GND.n6260 GND.n2788 218.815
R25020 GND.n6260 GND.n2789 218.815
R25021 GND.n6260 GND.n2790 218.815
R25022 GND.n6260 GND.n2791 218.815
R25023 GND.n6186 GND.n2771 218.815
R25024 GND.n2858 GND.n2771 218.815
R25025 GND.n6193 GND.n2771 218.815
R25026 GND.n2855 GND.n2771 218.815
R25027 GND.n6200 GND.n2771 218.815
R25028 GND.n2852 GND.n2771 218.815
R25029 GND.n6207 GND.n2771 218.815
R25030 GND.n2849 GND.n2771 218.815
R25031 GND.n6214 GND.n2771 218.815
R25032 GND.n2811 GND.n2771 218.815
R25033 GND.n6221 GND.n2771 218.815
R25034 GND.n2804 GND.n2771 218.815
R25035 GND.n6228 GND.n2771 218.815
R25036 GND.n2797 GND.n2771 218.815
R25037 GND.n6152 GND.n2771 218.815
R25038 GND.n6148 GND.n2771 218.815
R25039 GND.n6159 GND.n2771 218.815
R25040 GND.n6145 GND.n2771 218.815
R25041 GND.n6166 GND.n2771 218.815
R25042 GND.n6142 GND.n2771 218.815
R25043 GND.n6173 GND.n2771 218.815
R25044 GND.n6087 GND.n5984 218.815
R25045 GND.n5988 GND.n5984 218.815
R25046 GND.n6080 GND.n5984 218.815
R25047 GND.n6074 GND.n5984 218.815
R25048 GND.n6072 GND.n5984 218.815
R25049 GND.n6066 GND.n5984 218.815
R25050 GND.n6064 GND.n5984 218.815
R25051 GND.n6058 GND.n5984 218.815
R25052 GND.n6056 GND.n5984 218.815
R25053 GND.n6050 GND.n5984 218.815
R25054 GND.n6048 GND.n5984 218.815
R25055 GND.n6042 GND.n5984 218.815
R25056 GND.n6040 GND.n5984 218.815
R25057 GND.n6034 GND.n5984 218.815
R25058 GND.n6032 GND.n5984 218.815
R25059 GND.n6026 GND.n5984 218.815
R25060 GND.n6024 GND.n5984 218.815
R25061 GND.n6018 GND.n5984 218.815
R25062 GND.n6016 GND.n5984 218.815
R25063 GND.n6010 GND.n5984 218.815
R25064 GND.n6008 GND.n5984 218.815
R25065 GND.n7583 GND.n7582 218.815
R25066 GND.n7582 GND.n2411 218.815
R25067 GND.n7582 GND.n2412 218.815
R25068 GND.n7582 GND.n2413 218.815
R25069 GND.n7582 GND.n2414 218.815
R25070 GND.n7582 GND.n2415 218.815
R25071 GND.n7582 GND.n2416 218.815
R25072 GND.n7582 GND.n2417 218.815
R25073 GND.n7683 GND.n2317 218.815
R25074 GND.n7683 GND.n2318 218.815
R25075 GND.n7683 GND.n2319 218.815
R25076 GND.n7683 GND.n2320 218.815
R25077 GND.n7683 GND.n2321 218.815
R25078 GND.n7683 GND.n2322 218.815
R25079 GND.n7683 GND.n2323 218.815
R25080 GND.n7683 GND.n2324 218.815
R25081 GND.n5622 GND.n5621 218.815
R25082 GND.n5623 GND.n5622 218.815
R25083 GND.n5547 GND.n2335 218.815
R25084 GND.n5535 GND.n2335 218.815
R25085 GND.n5531 GND.n2335 218.815
R25086 GND.n5477 GND.n2387 218.815
R25087 GND.n5480 GND.n2387 218.815
R25088 GND.n5635 GND.n2387 218.815
R25089 GND.n5638 GND.n2387 218.815
R25090 GND.n5516 GND.n5514 218.815
R25091 GND.n5522 GND.n5514 218.815
R25092 GND.n5514 GND.n5489 218.815
R25093 GND.n5514 GND.n5499 218.815
R25094 GND.n5514 GND.n5491 218.815
R25095 GND.n6904 GND.n6863 218.815
R25096 GND.n6904 GND.n6864 218.815
R25097 GND.n6904 GND.n6865 218.815
R25098 GND.n6904 GND.n6866 218.815
R25099 GND.n6904 GND.n6867 218.815
R25100 GND.n6904 GND.n6868 218.815
R25101 GND.n6904 GND.n6869 218.815
R25102 GND.n6904 GND.n6903 218.815
R25103 GND.n6814 GND.n6802 218.815
R25104 GND.n6816 GND.n6802 218.815
R25105 GND.n6822 GND.n6802 218.815
R25106 GND.n6824 GND.n6802 218.815
R25107 GND.n6830 GND.n6802 218.815
R25108 GND.n6832 GND.n6802 218.815
R25109 GND.n6838 GND.n6802 218.815
R25110 GND.n6840 GND.n6802 218.815
R25111 GND.n7494 GND.n7493 218.815
R25112 GND.n7493 GND.n7455 218.815
R25113 GND.n7493 GND.n7456 218.815
R25114 GND.n7493 GND.n7457 218.815
R25115 GND.n7493 GND.n7458 218.815
R25116 GND.n7493 GND.n7459 218.815
R25117 GND.n7493 GND.n7460 218.815
R25118 GND.n7493 GND.n7461 218.815
R25119 GND GND.t112 218.543
R25120 GND.t332 GND 218.543
R25121 GND.n3097 GND.n3096 207.213
R25122 GND.n3006 GND.n2919 207.213
R25123 GND.n3041 GND.n3039 207.213
R25124 GND.n2978 GND.n2970 207.213
R25125 GND.n2964 GND.n2963 207.213
R25126 GND.n2942 GND.n2941 207.213
R25127 GND.n2940 GND.n2933 207.213
R25128 GND.n2925 GND.n2924 207.213
R25129 GND.n2991 GND.n2960 207.213
R25130 GND.n3001 GND.n2923 207.213
R25131 GND.n2917 GND.n2916 207.213
R25132 GND.n3015 GND.n3014 207.213
R25133 GND.n3025 GND.n2912 207.213
R25134 GND.n2906 GND.n2905 207.213
R25135 GND.n3046 GND.n3045 207.213
R25136 GND.n3048 GND.n3047 207.213
R25137 GND.n2904 GND.n2903 207.213
R25138 GND.n9796 GND.n9795 205.056
R25139 GND.t358 GND 203.975
R25140 GND GND.t148 203.975
R25141 GND GND.t371 203.975
R25142 GND.t317 GND.t272 203.975
R25143 GND.t318 GND.t110 203.975
R25144 GND.t315 GND.t199 203.975
R25145 GND.t316 GND.t368 203.975
R25146 GND.t292 GND.t369 203.975
R25147 GND.t367 GND.t298 203.975
R25148 GND.t8 GND.t269 203.975
R25149 GND.t37 GND.t397 203.975
R25150 GND.t344 GND.t346 203.975
R25151 GND.t364 GND.t347 203.975
R25152 GND.t362 GND.t387 203.975
R25153 GND.t381 GND.t365 203.975
R25154 GND.n9463 GND.n9432 194.953
R25155 GND.n3090 GND.n3089 194.788
R25156 GND.n3080 GND.t393 189.405
R25157 GND.n6598 GND.n6592 185
R25158 GND.n6598 GND.n6591 185
R25159 GND.n6599 GND.n6598 185
R25160 GND.n6584 GND.n6578 185
R25161 GND.n6584 GND.n6577 185
R25162 GND.n6585 GND.n6584 185
R25163 GND.n6570 GND.n6564 185
R25164 GND.n6570 GND.n6563 185
R25165 GND.n6571 GND.n6570 185
R25166 GND.n6556 GND.n6550 185
R25167 GND.n6556 GND.n6549 185
R25168 GND.n6557 GND.n6556 185
R25169 GND.n6542 GND.n6536 185
R25170 GND.n6542 GND.n6535 185
R25171 GND.n6543 GND.n6542 185
R25172 GND.n2708 GND.n2702 185
R25173 GND.n2708 GND.n2701 185
R25174 GND.n2709 GND.n2708 185
R25175 GND.n6457 GND.n6451 185
R25176 GND.n6457 GND.n6450 185
R25177 GND.n6458 GND.n6457 185
R25178 GND.n6471 GND.n6465 185
R25179 GND.n6471 GND.n6464 185
R25180 GND.n6472 GND.n6471 185
R25181 GND.n6484 GND.n6478 185
R25182 GND.n6484 GND.n6477 185
R25183 GND.n6485 GND.n6484 185
R25184 GND.n6497 GND.n6491 185
R25185 GND.n6497 GND.n6490 185
R25186 GND.n6498 GND.n6497 185
R25187 GND.n6510 GND.n6504 185
R25188 GND.n6510 GND.n6503 185
R25189 GND.n6511 GND.n6510 185
R25190 GND.n6523 GND.n6517 185
R25191 GND.n6523 GND.n6516 185
R25192 GND.n6524 GND.n6523 185
R25193 GND.n6438 GND.n6432 185
R25194 GND.n6438 GND.n6431 185
R25195 GND.n6439 GND.n6438 185
R25196 GND.n8961 GND.n8955 185
R25197 GND.n8961 GND.n8954 185
R25198 GND.n8962 GND.n8961 185
R25199 GND.n8947 GND.n8941 185
R25200 GND.n8947 GND.n8940 185
R25201 GND.n8948 GND.n8947 185
R25202 GND.n8933 GND.n8927 185
R25203 GND.n8933 GND.n8926 185
R25204 GND.n8934 GND.n8933 185
R25205 GND.n8919 GND.n8913 185
R25206 GND.n8919 GND.n8912 185
R25207 GND.n8920 GND.n8919 185
R25208 GND.n8905 GND.n8899 185
R25209 GND.n8905 GND.n8898 185
R25210 GND.n8906 GND.n8905 185
R25211 GND.n991 GND.n985 185
R25212 GND.n991 GND.n984 185
R25213 GND.n992 GND.n991 185
R25214 GND.n8821 GND.n8815 185
R25215 GND.n8821 GND.n8814 185
R25216 GND.n8822 GND.n8821 185
R25217 GND.n8835 GND.n8829 185
R25218 GND.n8835 GND.n8828 185
R25219 GND.n8836 GND.n8835 185
R25220 GND.n8848 GND.n8842 185
R25221 GND.n8848 GND.n8841 185
R25222 GND.n8849 GND.n8848 185
R25223 GND.n8861 GND.n8855 185
R25224 GND.n8861 GND.n8854 185
R25225 GND.n8862 GND.n8861 185
R25226 GND.n8874 GND.n8868 185
R25227 GND.n8874 GND.n8867 185
R25228 GND.n8875 GND.n8874 185
R25229 GND.n8887 GND.n8881 185
R25230 GND.n8887 GND.n8880 185
R25231 GND.n8888 GND.n8887 185
R25232 GND.n8802 GND.n8796 185
R25233 GND.n8802 GND.n8795 185
R25234 GND.n8803 GND.n8802 185
R25235 GND.n4860 GND.n4854 185
R25236 GND.n4860 GND.n4853 185
R25237 GND.n4861 GND.n4860 185
R25238 GND.n4846 GND.n4840 185
R25239 GND.n4846 GND.n4839 185
R25240 GND.n4847 GND.n4846 185
R25241 GND.n4832 GND.n4826 185
R25242 GND.n4832 GND.n4825 185
R25243 GND.n4833 GND.n4832 185
R25244 GND.n4818 GND.n4812 185
R25245 GND.n4818 GND.n4811 185
R25246 GND.n4819 GND.n4818 185
R25247 GND.n4804 GND.n4798 185
R25248 GND.n4804 GND.n4797 185
R25249 GND.n4805 GND.n4804 185
R25250 GND.n4789 GND.n4783 185
R25251 GND.n4789 GND.n4782 185
R25252 GND.n4790 GND.n4789 185
R25253 GND.n4183 GND.n4177 185
R25254 GND.n4183 GND.n4176 185
R25255 GND.n4184 GND.n4183 185
R25256 GND.n4877 GND.n4871 185
R25257 GND.n4877 GND.n4870 185
R25258 GND.n4878 GND.n4877 185
R25259 GND.n4890 GND.n4884 185
R25260 GND.n4890 GND.n4883 185
R25261 GND.n4891 GND.n4890 185
R25262 GND.n4903 GND.n4897 185
R25263 GND.n4903 GND.n4896 185
R25264 GND.n4904 GND.n4903 185
R25265 GND.n4916 GND.n4910 185
R25266 GND.n4916 GND.n4909 185
R25267 GND.n4917 GND.n4916 185
R25268 GND.n4929 GND.n4923 185
R25269 GND.n4929 GND.n4922 185
R25270 GND.n4930 GND.n4929 185
R25271 GND.n4164 GND.n4158 185
R25272 GND.n4164 GND.n4157 185
R25273 GND.n4165 GND.n4164 185
R25274 GND.t366 GND.n3079 174.834
R25275 GND.n7742 GND.n7740 160.037
R25276 GND.n9814 GND.n21 160.037
R25277 GND.n7690 GND.n2313 154.131
R25278 GND.n9808 GND.t379 153.792
R25279 GND.n8397 GND.t407 153.792
R25280 GND GND.t395 152.981
R25281 GND.n9798 GND.t124 150.475
R25282 GND.n9796 GND.t357 148.613
R25283 GND.n5494 GND.n5491 147.374
R25284 GND.n5499 GND.n5498 147.374
R25285 GND.n5524 GND.n5489 147.374
R25286 GND.n5522 GND.n5521 147.374
R25287 GND.n5517 GND.n5516 147.374
R25288 GND.n5477 GND.n5476 147.374
R25289 GND.n5481 GND.n5480 147.374
R25290 GND.n5635 GND.n5634 147.374
R25291 GND.n5638 GND.n5637 147.374
R25292 GND.n5533 GND.n5531 147.374
R25293 GND.n5549 GND.n5535 147.374
R25294 GND.n5547 GND.n5546 147.374
R25295 GND.n5621 GND.n5620 147.374
R25296 GND.n5624 GND.n5623 147.374
R25297 GND.n7678 GND.n2324 147.374
R25298 GND.n7674 GND.n2323 147.374
R25299 GND.n7670 GND.n2322 147.374
R25300 GND.n7666 GND.n2321 147.374
R25301 GND.n7662 GND.n2320 147.374
R25302 GND.n7658 GND.n2319 147.374
R25303 GND.n7654 GND.n2318 147.374
R25304 GND.n7650 GND.n2317 147.374
R25305 GND.n7583 GND.n2408 147.374
R25306 GND.n5564 GND.n2411 147.374
R25307 GND.n5568 GND.n2412 147.374
R25308 GND.n5572 GND.n2413 147.374
R25309 GND.n5576 GND.n2414 147.374
R25310 GND.n5580 GND.n2415 147.374
R25311 GND.n5584 GND.n2416 147.374
R25312 GND.n5588 GND.n2417 147.374
R25313 GND.n6087 GND.n5986 147.374
R25314 GND.n6085 GND.n5988 147.374
R25315 GND.n6081 GND.n6080 147.374
R25316 GND.n6074 GND.n5990 147.374
R25317 GND.n6073 GND.n6072 147.374
R25318 GND.n6066 GND.n5992 147.374
R25319 GND.n6065 GND.n6064 147.374
R25320 GND.n6058 GND.n5994 147.374
R25321 GND.n6057 GND.n6056 147.374
R25322 GND.n6050 GND.n5996 147.374
R25323 GND.n6049 GND.n6048 147.374
R25324 GND.n6042 GND.n5998 147.374
R25325 GND.n6041 GND.n6040 147.374
R25326 GND.n6034 GND.n6000 147.374
R25327 GND.n6033 GND.n6032 147.374
R25328 GND.n6026 GND.n6002 147.374
R25329 GND.n6025 GND.n6024 147.374
R25330 GND.n6018 GND.n6004 147.374
R25331 GND.n6017 GND.n6016 147.374
R25332 GND.n6010 GND.n6006 147.374
R25333 GND.n6009 GND.n6008 147.374
R25334 GND.n6173 GND.n6172 147.374
R25335 GND.n6168 GND.n6142 147.374
R25336 GND.n6166 GND.n6165 147.374
R25337 GND.n6161 GND.n6145 147.374
R25338 GND.n6159 GND.n6158 147.374
R25339 GND.n6154 GND.n6148 147.374
R25340 GND.n6152 GND.n6151 147.374
R25341 GND.n6230 GND.n2797 147.374
R25342 GND.n6228 GND.n6227 147.374
R25343 GND.n6223 GND.n2804 147.374
R25344 GND.n6221 GND.n6220 147.374
R25345 GND.n6216 GND.n2811 147.374
R25346 GND.n6214 GND.n6213 147.374
R25347 GND.n6209 GND.n2849 147.374
R25348 GND.n6207 GND.n6206 147.374
R25349 GND.n6202 GND.n2852 147.374
R25350 GND.n6200 GND.n6199 147.374
R25351 GND.n6195 GND.n2855 147.374
R25352 GND.n6193 GND.n6192 147.374
R25353 GND.n6188 GND.n2858 147.374
R25354 GND.n6186 GND.n6185 147.374
R25355 GND.n6262 GND.n6261 147.374
R25356 GND.n2792 GND.n2772 147.374
R25357 GND.n6254 GND.n2773 147.374
R25358 GND.n6250 GND.n2774 147.374
R25359 GND.n6246 GND.n2775 147.374
R25360 GND.n6242 GND.n2776 147.374
R25361 GND.n6238 GND.n2777 147.374
R25362 GND.n6234 GND.n2778 147.374
R25363 GND.n2795 GND.n2779 147.374
R25364 GND.n2800 GND.n2780 147.374
R25365 GND.n2802 GND.n2781 147.374
R25366 GND.n2807 GND.n2782 147.374
R25367 GND.n2809 GND.n2783 147.374
R25368 GND.n2844 GND.n2784 147.374
R25369 GND.n2840 GND.n2785 147.374
R25370 GND.n2836 GND.n2786 147.374
R25371 GND.n2832 GND.n2787 147.374
R25372 GND.n2828 GND.n2788 147.374
R25373 GND.n2824 GND.n2789 147.374
R25374 GND.n2820 GND.n2790 147.374
R25375 GND.n2816 GND.n2791 147.374
R25376 GND.n6382 GND.n6381 147.374
R25377 GND.n6379 GND.n6378 147.374
R25378 GND.n6374 GND.n6319 147.374
R25379 GND.n6372 GND.n6371 147.374
R25380 GND.n6367 GND.n6322 147.374
R25381 GND.n6365 GND.n6364 147.374
R25382 GND.n6360 GND.n6325 147.374
R25383 GND.n6358 GND.n6357 147.374
R25384 GND.n6333 GND.n6332 147.374
R25385 GND.n6346 GND.n6345 147.374
R25386 GND.n6343 GND.n6342 147.374
R25387 GND.n6335 GND.n2719 147.374
R25388 GND.n6419 GND.n6418 147.374
R25389 GND.n6416 GND.n6415 147.374
R25390 GND.n6411 GND.n2724 147.374
R25391 GND.n6409 GND.n6408 147.374
R25392 GND.n6404 GND.n2727 147.374
R25393 GND.n6402 GND.n6401 147.374
R25394 GND.n6397 GND.n2730 147.374
R25395 GND.n6395 GND.n6394 147.374
R25396 GND.n6390 GND.n2733 147.374
R25397 GND.n5981 GND.n5980 147.374
R25398 GND.n5975 GND.n3697 147.374
R25399 GND.n5972 GND.n3698 147.374
R25400 GND.n5968 GND.n3699 147.374
R25401 GND.n5964 GND.n3700 147.374
R25402 GND.n5960 GND.n3701 147.374
R25403 GND.n5956 GND.n3702 147.374
R25404 GND.n5952 GND.n3703 147.374
R25405 GND.n5948 GND.n3704 147.374
R25406 GND.n5944 GND.n3705 147.374
R25407 GND.n5940 GND.n3706 147.374
R25408 GND.n5936 GND.n3707 147.374
R25409 GND.n5932 GND.n3708 147.374
R25410 GND.n5928 GND.n3709 147.374
R25411 GND.n5924 GND.n3710 147.374
R25412 GND.n5920 GND.n3711 147.374
R25413 GND.n5916 GND.n3712 147.374
R25414 GND.n5912 GND.n3713 147.374
R25415 GND.n5908 GND.n3714 147.374
R25416 GND.n5904 GND.n3715 147.374
R25417 GND.n5900 GND.n3716 147.374
R25418 GND.n5840 GND.n3810 147.374
R25419 GND.n5836 GND.n3809 147.374
R25420 GND.n5832 GND.n3808 147.374
R25421 GND.n5828 GND.n3807 147.374
R25422 GND.n5824 GND.n3806 147.374
R25423 GND.n5820 GND.n3805 147.374
R25424 GND.n5816 GND.n3804 147.374
R25425 GND.n4017 GND.n3803 147.374
R25426 GND.n4023 GND.n3802 147.374
R25427 GND.n4029 GND.n3801 147.374
R25428 GND.n4035 GND.n3800 147.374
R25429 GND.n4041 GND.n3799 147.374
R25430 GND.n4014 GND.n3798 147.374
R25431 GND.n4010 GND.n3797 147.374
R25432 GND.n4006 GND.n3796 147.374
R25433 GND.n4002 GND.n3795 147.374
R25434 GND.n3998 GND.n3794 147.374
R25435 GND.n3994 GND.n3793 147.374
R25436 GND.n3990 GND.n3792 147.374
R25437 GND.n3986 GND.n3791 147.374
R25438 GND.n3982 GND.n3790 147.374
R25439 GND.n5194 GND.n3726 147.374
R25440 GND.n5200 GND.n5199 147.374
R25441 GND.n5203 GND.n5202 147.374
R25442 GND.n5208 GND.n5207 147.374
R25443 GND.n5211 GND.n5210 147.374
R25444 GND.n5216 GND.n5215 147.374
R25445 GND.n5219 GND.n5218 147.374
R25446 GND.n5224 GND.n5223 147.374
R25447 GND.n5227 GND.n5226 147.374
R25448 GND.n5232 GND.n5231 147.374
R25449 GND.n5235 GND.n5234 147.374
R25450 GND.n5240 GND.n5239 147.374
R25451 GND.n5243 GND.n5242 147.374
R25452 GND.n5248 GND.n5247 147.374
R25453 GND.n5251 GND.n5250 147.374
R25454 GND.n5256 GND.n5255 147.374
R25455 GND.n5259 GND.n5258 147.374
R25456 GND.n5264 GND.n5263 147.374
R25457 GND.n5267 GND.n5266 147.374
R25458 GND.n5272 GND.n5271 147.374
R25459 GND.n5275 GND.n5274 147.374
R25460 GND.n5059 GND.n5058 147.374
R25461 GND.n5060 GND.n5054 147.374
R25462 GND.n5067 GND.n5066 147.374
R25463 GND.n5068 GND.n5052 147.374
R25464 GND.n5075 GND.n5074 147.374
R25465 GND.n5076 GND.n5050 147.374
R25466 GND.n5083 GND.n5082 147.374
R25467 GND.n5084 GND.n5048 147.374
R25468 GND.n5137 GND.n5136 147.374
R25469 GND.n5138 GND.n5044 147.374
R25470 GND.n5149 GND.n5148 147.374
R25471 GND.n5150 GND.n5040 147.374
R25472 GND.n5162 GND.n5161 147.374
R25473 GND.n5336 GND.n5335 147.374
R25474 GND.n5333 GND.n5332 147.374
R25475 GND.n5328 GND.n5166 147.374
R25476 GND.n5326 GND.n5325 147.374
R25477 GND.n5321 GND.n5169 147.374
R25478 GND.n5319 GND.n5318 147.374
R25479 GND.n5314 GND.n5172 147.374
R25480 GND.n5312 GND.n5311 147.374
R25481 GND.n5808 GND.n5807 147.374
R25482 GND.n5802 GND.n3818 147.374
R25483 GND.n5799 GND.n3819 147.374
R25484 GND.n5795 GND.n3820 147.374
R25485 GND.n5791 GND.n3821 147.374
R25486 GND.n5787 GND.n3822 147.374
R25487 GND.n5783 GND.n3823 147.374
R25488 GND.n5811 GND.n5810 147.374
R25489 GND.n4016 GND.n3824 147.374
R25490 GND.n4022 GND.n3825 147.374
R25491 GND.n4028 GND.n3826 147.374
R25492 GND.n4034 GND.n3827 147.374
R25493 GND.n4040 GND.n3828 147.374
R25494 GND.n4047 GND.n3829 147.374
R25495 GND.n4051 GND.n3830 147.374
R25496 GND.n4055 GND.n3831 147.374
R25497 GND.n4059 GND.n3832 147.374
R25498 GND.n4063 GND.n3833 147.374
R25499 GND.n4067 GND.n3834 147.374
R25500 GND.n4071 GND.n3835 147.374
R25501 GND.n4075 GND.n3836 147.374
R25502 GND.n4977 GND.n3926 147.374
R25503 GND.n4973 GND.n3925 147.374
R25504 GND.n4969 GND.n3924 147.374
R25505 GND.n4965 GND.n3923 147.374
R25506 GND.n4961 GND.n3922 147.374
R25507 GND.n4957 GND.n3921 147.374
R25508 GND.n4953 GND.n3920 147.374
R25509 GND.n4949 GND.n3919 147.374
R25510 GND.n3939 GND.n3918 147.374
R25511 GND.n3943 GND.n3917 147.374
R25512 GND.n3947 GND.n3916 147.374
R25513 GND.n4146 GND.n3915 147.374
R25514 GND.n4144 GND.n3914 147.374
R25515 GND.n4140 GND.n3913 147.374
R25516 GND.n4136 GND.n3912 147.374
R25517 GND.n4132 GND.n3911 147.374
R25518 GND.n4128 GND.n3910 147.374
R25519 GND.n4124 GND.n3909 147.374
R25520 GND.n4120 GND.n3908 147.374
R25521 GND.n4116 GND.n3907 147.374
R25522 GND.n4112 GND.n3906 147.374
R25523 GND.n5098 GND.n5097 147.374
R25524 GND.n5104 GND.n5103 147.374
R25525 GND.n5107 GND.n5106 147.374
R25526 GND.n5112 GND.n5111 147.374
R25527 GND.n5115 GND.n5114 147.374
R25528 GND.n5120 GND.n5119 147.374
R25529 GND.n5123 GND.n5122 147.374
R25530 GND.n5128 GND.n5127 147.374
R25531 GND.n5131 GND.n5130 147.374
R25532 GND.n5142 GND.n5141 147.374
R25533 GND.n5145 GND.n5144 147.374
R25534 GND.n5154 GND.n5153 147.374
R25535 GND.n5158 GND.n5157 147.374
R25536 GND.n5039 GND.n5038 147.374
R25537 GND.n5343 GND.n5342 147.374
R25538 GND.n5346 GND.n5345 147.374
R25539 GND.n5351 GND.n5350 147.374
R25540 GND.n5354 GND.n5353 147.374
R25541 GND.n5359 GND.n5358 147.374
R25542 GND.n5362 GND.n5361 147.374
R25543 GND.n5367 GND.n5366 147.374
R25544 GND.n5728 GND.n5727 147.374
R25545 GND.n5723 GND.n5002 147.374
R25546 GND.n5719 GND.n5001 147.374
R25547 GND.n5715 GND.n5000 147.374
R25548 GND.n5711 GND.n4999 147.374
R25549 GND.n5707 GND.n4998 147.374
R25550 GND.n5703 GND.n4997 147.374
R25551 GND.n5699 GND.n4996 147.374
R25552 GND.n5695 GND.n4995 147.374
R25553 GND.n5015 GND.n4994 147.374
R25554 GND.n5019 GND.n4993 147.374
R25555 GND.n5023 GND.n4992 147.374
R25556 GND.n5432 GND.n4991 147.374
R25557 GND.n5430 GND.n4990 147.374
R25558 GND.n5426 GND.n4989 147.374
R25559 GND.n5422 GND.n4988 147.374
R25560 GND.n5418 GND.n4987 147.374
R25561 GND.n5414 GND.n4986 147.374
R25562 GND.n5410 GND.n4985 147.374
R25563 GND.n5406 GND.n4984 147.374
R25564 GND.n5402 GND.n4983 147.374
R25565 GND.n2235 GND.n2222 147.374
R25566 GND.n2239 GND.n2223 147.374
R25567 GND.n2246 GND.n2224 147.374
R25568 GND.n2249 GND.n2225 147.374
R25569 GND.n7864 GND.n7863 147.374
R25570 GND.n7954 GND.n7953 147.374
R25571 GND.n7948 GND.n2176 147.374
R25572 GND.n7943 GND.n2177 147.374
R25573 GND.n7938 GND.n2178 147.374
R25574 GND.n7832 GND.n7831 147.374
R25575 GND.n7829 GND.n7828 147.374
R25576 GND.n7824 GND.n7823 147.374
R25577 GND.n7985 GND.n7984 147.374
R25578 GND.n2145 GND.n2139 147.374
R25579 GND.n7784 GND.n7756 147.374
R25580 GND.n7780 GND.n7755 147.374
R25581 GND.n7776 GND.n7754 147.374
R25582 GND.n7772 GND.n7753 147.374
R25583 GND.n7768 GND.n7752 147.374
R25584 GND.n7764 GND.n7751 147.374
R25585 GND.n7760 GND.n7750 147.374
R25586 GND.n7749 GND.n2270 147.374
R25587 GND.n8028 GND.n8027 147.374
R25588 GND.n8022 GND.n2120 147.374
R25589 GND.n8019 GND.n2121 147.374
R25590 GND.n8015 GND.n2122 147.374
R25591 GND.n8011 GND.n2123 147.374
R25592 GND.n8007 GND.n2124 147.374
R25593 GND.n8003 GND.n2125 147.374
R25594 GND.n7999 GND.n2126 147.374
R25595 GND.n143 GND.n138 147.374
R25596 GND.n148 GND.n147 147.374
R25597 GND.n9598 GND.n136 147.374
R25598 GND.n9596 GND.n9595 147.374
R25599 GND.n9591 GND.n159 147.374
R25600 GND.n9733 GND.n9732 147.374
R25601 GND.n9727 GND.n92 147.374
R25602 GND.n9722 GND.n93 147.374
R25603 GND.n9717 GND.n94 147.374
R25604 GND.n9554 GND.n9553 147.374
R25605 GND.n9551 GND.n9550 147.374
R25606 GND.n9546 GND.n9545 147.374
R25607 GND.n9689 GND.n123 147.374
R25608 GND.n9608 GND.n129 147.374
R25609 GND.n9504 GND.n9503 147.374
R25610 GND.n9499 GND.n9471 147.374
R25611 GND.n9495 GND.n9470 147.374
R25612 GND.n9491 GND.n9469 147.374
R25613 GND.n9487 GND.n9468 147.374
R25614 GND.n9483 GND.n9467 147.374
R25615 GND.n9479 GND.n9466 147.374
R25616 GND.n9475 GND.n9465 147.374
R25617 GND.n9679 GND.n9620 147.374
R25618 GND.n9674 GND.n9622 147.374
R25619 GND.n9671 GND.n9623 147.374
R25620 GND.n9667 GND.n9624 147.374
R25621 GND.n9663 GND.n9625 147.374
R25622 GND.n9659 GND.n9626 147.374
R25623 GND.n9655 GND.n9627 147.374
R25624 GND.n9651 GND.n9628 147.374
R25625 GND.n1153 GND.n1071 147.374
R25626 GND.n1157 GND.n1072 147.374
R25627 GND.n1161 GND.n1073 147.374
R25628 GND.n1165 GND.n1074 147.374
R25629 GND.n1169 GND.n1075 147.374
R25630 GND.n1173 GND.n1076 147.374
R25631 GND.n1177 GND.n1077 147.374
R25632 GND.n1181 GND.n1078 147.374
R25633 GND.n1184 GND.n1079 147.374
R25634 GND.n1318 GND.n1288 147.374
R25635 GND.n1322 GND.n1321 147.374
R25636 GND.n1327 GND.n1326 147.374
R25637 GND.n1330 GND.n1329 147.374
R25638 GND.n1335 GND.n1334 147.374
R25639 GND.n1338 GND.n1337 147.374
R25640 GND.n1343 GND.n1342 147.374
R25641 GND.n1346 GND.n1345 147.374
R25642 GND.n1373 GND.n1080 147.374
R25643 GND.n1377 GND.n1081 147.374
R25644 GND.n1381 GND.n1082 147.374
R25645 GND.n1385 GND.n1083 147.374
R25646 GND.n1389 GND.n1084 147.374
R25647 GND.n1393 GND.n1085 147.374
R25648 GND.n1397 GND.n1086 147.374
R25649 GND.n1401 GND.n1087 147.374
R25650 GND.n1404 GND.n1088 147.374
R25651 GND.n1520 GND.n1353 147.374
R25652 GND.n1519 GND.n1518 147.374
R25653 GND.n1512 GND.n1355 147.374
R25654 GND.n1511 GND.n1510 147.374
R25655 GND.n1504 GND.n1357 147.374
R25656 GND.n1503 GND.n1502 147.374
R25657 GND.n1496 GND.n1359 147.374
R25658 GND.n1495 GND.n1494 147.374
R25659 GND.n1488 GND.n1361 147.374
R25660 GND.n8445 GND.n8432 147.374
R25661 GND.n8449 GND.n8433 147.374
R25662 GND.n8453 GND.n8434 147.374
R25663 GND.n8457 GND.n8435 147.374
R25664 GND.n8461 GND.n8436 147.374
R25665 GND.n8465 GND.n8437 147.374
R25666 GND.n8469 GND.n8438 147.374
R25667 GND.n8472 GND.n8439 147.374
R25668 GND.n8498 GND.n8497 147.374
R25669 GND.n8730 GND.n8729 147.374
R25670 GND.n1723 GND.n1063 147.374
R25671 GND.n8722 GND.n1064 147.374
R25672 GND.n8718 GND.n1065 147.374
R25673 GND.n8714 GND.n1066 147.374
R25674 GND.n8710 GND.n1067 147.374
R25675 GND.n8706 GND.n1068 147.374
R25676 GND.n8702 GND.n1069 147.374
R25677 GND.n3199 GND.n3117 147.374
R25678 GND.n3203 GND.n3118 147.374
R25679 GND.n3207 GND.n3119 147.374
R25680 GND.n3211 GND.n3120 147.374
R25681 GND.n3215 GND.n3121 147.374
R25682 GND.n3219 GND.n3122 147.374
R25683 GND.n3223 GND.n3123 147.374
R25684 GND.n3227 GND.n3124 147.374
R25685 GND.n3230 GND.n3125 147.374
R25686 GND.n3398 GND.n3334 147.374
R25687 GND.n3393 GND.n3337 147.374
R25688 GND.n3390 GND.n3338 147.374
R25689 GND.n3386 GND.n3339 147.374
R25690 GND.n3382 GND.n3340 147.374
R25691 GND.n3378 GND.n3341 147.374
R25692 GND.n3374 GND.n3342 147.374
R25693 GND.n3370 GND.n3343 147.374
R25694 GND.n8589 GND.n8588 147.374
R25695 GND.n8586 GND.n8585 147.374
R25696 GND.n8581 GND.n8503 147.374
R25697 GND.n8579 GND.n8578 147.374
R25698 GND.n8574 GND.n8506 147.374
R25699 GND.n8572 GND.n8571 147.374
R25700 GND.n8567 GND.n8509 147.374
R25701 GND.n8565 GND.n8564 147.374
R25702 GND.n8560 GND.n8558 147.374
R25703 GND.n1722 GND.n1721 147.374
R25704 GND.n1717 GND.n1661 147.374
R25705 GND.n1714 GND.n1660 147.374
R25706 GND.n1710 GND.n1659 147.374
R25707 GND.n1706 GND.n1658 147.374
R25708 GND.n1702 GND.n1657 147.374
R25709 GND.n1698 GND.n1656 147.374
R25710 GND.n1694 GND.n1655 147.374
R25711 GND.n1690 GND.n1654 147.374
R25712 GND.n9199 GND.n9139 147.374
R25713 GND.n9197 GND.n9141 147.374
R25714 GND.n9193 GND.n9192 147.374
R25715 GND.n9186 GND.n9143 147.374
R25716 GND.n9185 GND.n9184 147.374
R25717 GND.n9178 GND.n9145 147.374
R25718 GND.n9177 GND.n9176 147.374
R25719 GND.n9170 GND.n9147 147.374
R25720 GND.n610 GND.n584 147.374
R25721 GND.n606 GND.n583 147.374
R25722 GND.n602 GND.n582 147.374
R25723 GND.n598 GND.n581 147.374
R25724 GND.n594 GND.n580 147.374
R25725 GND.n590 GND.n579 147.374
R25726 GND.n586 GND.n578 147.374
R25727 GND.n617 GND.n616 147.374
R25728 GND.n9134 GND.n9133 147.374
R25729 GND.n9128 GND.n418 147.374
R25730 GND.n9125 GND.n419 147.374
R25731 GND.n9121 GND.n420 147.374
R25732 GND.n9117 GND.n421 147.374
R25733 GND.n9113 GND.n422 147.374
R25734 GND.n9109 GND.n423 147.374
R25735 GND.n9105 GND.n424 147.374
R25736 GND.n677 GND.n676 147.374
R25737 GND.n672 GND.n646 147.374
R25738 GND.n668 GND.n645 147.374
R25739 GND.n664 GND.n644 147.374
R25740 GND.n660 GND.n643 147.374
R25741 GND.n656 GND.n642 147.374
R25742 GND.n652 GND.n641 147.374
R25743 GND.n648 GND.n640 147.374
R25744 GND.n758 GND.n505 147.374
R25745 GND.n762 GND.n506 147.374
R25746 GND.n766 GND.n507 147.374
R25747 GND.n770 GND.n508 147.374
R25748 GND.n774 GND.n509 147.374
R25749 GND.n778 GND.n510 147.374
R25750 GND.n782 GND.n511 147.374
R25751 GND.n753 GND.n512 147.374
R25752 GND.n9344 GND.n9343 147.374
R25753 GND.n9338 GND.n302 147.374
R25754 GND.n9335 GND.n303 147.374
R25755 GND.n9331 GND.n304 147.374
R25756 GND.n9327 GND.n305 147.374
R25757 GND.n9323 GND.n306 147.374
R25758 GND.n9319 GND.n307 147.374
R25759 GND.n9315 GND.n308 147.374
R25760 GND.n9344 GND.n319 147.374
R25761 GND.n9336 GND.n302 147.374
R25762 GND.n9332 GND.n303 147.374
R25763 GND.n9328 GND.n304 147.374
R25764 GND.n9324 GND.n305 147.374
R25765 GND.n9320 GND.n306 147.374
R25766 GND.n9316 GND.n307 147.374
R25767 GND.n9312 GND.n308 147.374
R25768 GND.n783 GND.n512 147.374
R25769 GND.n779 GND.n511 147.374
R25770 GND.n775 GND.n510 147.374
R25771 GND.n771 GND.n509 147.374
R25772 GND.n767 GND.n508 147.374
R25773 GND.n763 GND.n507 147.374
R25774 GND.n759 GND.n506 147.374
R25775 GND.n755 GND.n505 147.374
R25776 GND.n9347 GND.n9346 147.374
R25777 GND.n8983 GND.n309 147.374
R25778 GND.n8987 GND.n310 147.374
R25779 GND.n8991 GND.n311 147.374
R25780 GND.n8995 GND.n312 147.374
R25781 GND.n8999 GND.n313 147.374
R25782 GND.n9003 GND.n314 147.374
R25783 GND.n9007 GND.n315 147.374
R25784 GND.n793 GND.n513 147.374
R25785 GND.n797 GND.n514 147.374
R25786 GND.n801 GND.n515 147.374
R25787 GND.n805 GND.n516 147.374
R25788 GND.n809 GND.n517 147.374
R25789 GND.n813 GND.n518 147.374
R25790 GND.n817 GND.n519 147.374
R25791 GND.n821 GND.n520 147.374
R25792 GND.n521 GND.n520 147.374
R25793 GND.n820 GND.n519 147.374
R25794 GND.n816 GND.n518 147.374
R25795 GND.n812 GND.n517 147.374
R25796 GND.n808 GND.n516 147.374
R25797 GND.n804 GND.n515 147.374
R25798 GND.n800 GND.n514 147.374
R25799 GND.n796 GND.n513 147.374
R25800 GND.n9346 GND.n300 147.374
R25801 GND.n8986 GND.n309 147.374
R25802 GND.n8990 GND.n310 147.374
R25803 GND.n8994 GND.n311 147.374
R25804 GND.n8998 GND.n312 147.374
R25805 GND.n9002 GND.n313 147.374
R25806 GND.n9006 GND.n314 147.374
R25807 GND.n9009 GND.n315 147.374
R25808 GND.n3420 GND.n3126 147.374
R25809 GND.n3424 GND.n3127 147.374
R25810 GND.n3428 GND.n3128 147.374
R25811 GND.n3432 GND.n3129 147.374
R25812 GND.n3436 GND.n3130 147.374
R25813 GND.n3440 GND.n3131 147.374
R25814 GND.n3444 GND.n3132 147.374
R25815 GND.n3448 GND.n3133 147.374
R25816 GND.n3451 GND.n3134 147.374
R25817 GND.n3563 GND.n3400 147.374
R25818 GND.n3562 GND.n3561 147.374
R25819 GND.n3555 GND.n3402 147.374
R25820 GND.n3554 GND.n3553 147.374
R25821 GND.n3547 GND.n3404 147.374
R25822 GND.n3546 GND.n3545 147.374
R25823 GND.n3539 GND.n3406 147.374
R25824 GND.n3538 GND.n3537 147.374
R25825 GND.n3531 GND.n3408 147.374
R25826 GND.n8093 GND.n8033 147.374
R25827 GND.n8091 GND.n8035 147.374
R25828 GND.n8087 GND.n8086 147.374
R25829 GND.n8080 GND.n8037 147.374
R25830 GND.n8079 GND.n8078 147.374
R25831 GND.n8072 GND.n8039 147.374
R25832 GND.n8071 GND.n8070 147.374
R25833 GND.n8064 GND.n8041 147.374
R25834 GND.n8391 GND.n1824 147.374
R25835 GND.n8387 GND.n1823 147.374
R25836 GND.n8383 GND.n1822 147.374
R25837 GND.n8379 GND.n1821 147.374
R25838 GND.n8375 GND.n1820 147.374
R25839 GND.n8371 GND.n1819 147.374
R25840 GND.n8367 GND.n1818 147.374
R25841 GND.n8363 GND.n1817 147.374
R25842 GND.n4569 GND.n4568 147.374
R25843 GND.n4575 GND.n4574 147.374
R25844 GND.n4578 GND.n4577 147.374
R25845 GND.n4583 GND.n4582 147.374
R25846 GND.n4586 GND.n4585 147.374
R25847 GND.n4591 GND.n4590 147.374
R25848 GND.n4594 GND.n4593 147.374
R25849 GND.n4599 GND.n4598 147.374
R25850 GND.n4284 GND.n4283 147.374
R25851 GND.n4291 GND.n4290 147.374
R25852 GND.n4292 GND.n4281 147.374
R25853 GND.n4299 GND.n4298 147.374
R25854 GND.n4300 GND.n4279 147.374
R25855 GND.n4307 GND.n4306 147.374
R25856 GND.n4311 GND.n4277 147.374
R25857 GND.n4314 GND.n4313 147.374
R25858 GND.n4371 GND.n4359 147.374
R25859 GND.n4375 GND.n4360 147.374
R25860 GND.n4379 GND.n4361 147.374
R25861 GND.n4383 GND.n4362 147.374
R25862 GND.n4387 GND.n4363 147.374
R25863 GND.n4391 GND.n4364 147.374
R25864 GND.n4394 GND.n4365 147.374
R25865 GND.n4403 GND.n4402 147.374
R25866 GND.n8238 GND.n8237 147.374
R25867 GND.n8232 GND.n1994 147.374
R25868 GND.n8229 GND.n1995 147.374
R25869 GND.n8225 GND.n1996 147.374
R25870 GND.n8221 GND.n1997 147.374
R25871 GND.n8217 GND.n1998 147.374
R25872 GND.n8213 GND.n1999 147.374
R25873 GND.n8209 GND.n2000 147.374
R25874 GND.n8238 GND.n2011 147.374
R25875 GND.n8230 GND.n1994 147.374
R25876 GND.n8226 GND.n1995 147.374
R25877 GND.n8222 GND.n1996 147.374
R25878 GND.n8218 GND.n1997 147.374
R25879 GND.n8214 GND.n1998 147.374
R25880 GND.n8210 GND.n1999 147.374
R25881 GND.n8206 GND.n2000 147.374
R25882 GND.n4403 GND.n4366 147.374
R25883 GND.n4392 GND.n4365 147.374
R25884 GND.n4388 GND.n4364 147.374
R25885 GND.n4384 GND.n4363 147.374
R25886 GND.n4380 GND.n4362 147.374
R25887 GND.n4376 GND.n4361 147.374
R25888 GND.n4372 GND.n4360 147.374
R25889 GND.n4368 GND.n4359 147.374
R25890 GND.n8241 GND.n8240 147.374
R25891 GND.n4726 GND.n2001 147.374
R25892 GND.n4730 GND.n2002 147.374
R25893 GND.n4734 GND.n2003 147.374
R25894 GND.n4738 GND.n2004 147.374
R25895 GND.n4742 GND.n2005 147.374
R25896 GND.n4746 GND.n2006 147.374
R25897 GND.n4750 GND.n2007 147.374
R25898 GND.n4441 GND.n4267 147.374
R25899 GND.n4404 GND.n4269 147.374
R25900 GND.n4414 GND.n4405 147.374
R25901 GND.n4418 GND.n4406 147.374
R25902 GND.n4422 GND.n4407 147.374
R25903 GND.n4426 GND.n4408 147.374
R25904 GND.n4430 GND.n4409 147.374
R25905 GND.n4434 GND.n4410 147.374
R25906 GND.n4411 GND.n4410 147.374
R25907 GND.n4433 GND.n4409 147.374
R25908 GND.n4429 GND.n4408 147.374
R25909 GND.n4425 GND.n4407 147.374
R25910 GND.n4421 GND.n4406 147.374
R25911 GND.n4417 GND.n4405 147.374
R25912 GND.n4413 GND.n4404 147.374
R25913 GND.n4442 GND.n4441 147.374
R25914 GND.n8240 GND.n1992 147.374
R25915 GND.n4729 GND.n2001 147.374
R25916 GND.n4733 GND.n2002 147.374
R25917 GND.n4737 GND.n2003 147.374
R25918 GND.n4741 GND.n2004 147.374
R25919 GND.n4745 GND.n2005 147.374
R25920 GND.n4749 GND.n2006 147.374
R25921 GND.n4752 GND.n2007 147.374
R25922 GND.n3564 GND.n3563 147.374
R25923 GND.n3561 GND.n3560 147.374
R25924 GND.n3556 GND.n3555 147.374
R25925 GND.n3553 GND.n3552 147.374
R25926 GND.n3548 GND.n3547 147.374
R25927 GND.n3545 GND.n3544 147.374
R25928 GND.n3540 GND.n3539 147.374
R25929 GND.n3537 GND.n3536 147.374
R25930 GND.n3532 GND.n3531 147.374
R25931 GND.n3449 GND.n3134 147.374
R25932 GND.n3445 GND.n3133 147.374
R25933 GND.n3441 GND.n3132 147.374
R25934 GND.n3437 GND.n3131 147.374
R25935 GND.n3433 GND.n3130 147.374
R25936 GND.n3429 GND.n3129 147.374
R25937 GND.n3425 GND.n3128 147.374
R25938 GND.n3421 GND.n3127 147.374
R25939 GND.n3417 GND.n3126 147.374
R25940 GND.n1722 GND.n1662 147.374
R25941 GND.n1715 GND.n1661 147.374
R25942 GND.n1711 GND.n1660 147.374
R25943 GND.n1707 GND.n1659 147.374
R25944 GND.n1703 GND.n1658 147.374
R25945 GND.n1699 GND.n1657 147.374
R25946 GND.n1695 GND.n1656 147.374
R25947 GND.n1691 GND.n1655 147.374
R25948 GND.n1687 GND.n1654 147.374
R25949 GND.n8558 GND.n8510 147.374
R25950 GND.n8566 GND.n8565 147.374
R25951 GND.n8509 GND.n8507 147.374
R25952 GND.n8573 GND.n8572 147.374
R25953 GND.n8506 GND.n8504 147.374
R25954 GND.n8580 GND.n8579 147.374
R25955 GND.n8503 GND.n8501 147.374
R25956 GND.n8587 GND.n8586 147.374
R25957 GND.n8590 GND.n8589 147.374
R25958 GND.n3398 GND.n3397 147.374
R25959 GND.n3391 GND.n3337 147.374
R25960 GND.n3387 GND.n3338 147.374
R25961 GND.n3383 GND.n3339 147.374
R25962 GND.n3379 GND.n3340 147.374
R25963 GND.n3375 GND.n3341 147.374
R25964 GND.n3371 GND.n3342 147.374
R25965 GND.n3367 GND.n3343 147.374
R25966 GND.n3228 GND.n3125 147.374
R25967 GND.n3224 GND.n3124 147.374
R25968 GND.n3220 GND.n3123 147.374
R25969 GND.n3216 GND.n3122 147.374
R25970 GND.n3212 GND.n3121 147.374
R25971 GND.n3208 GND.n3120 147.374
R25972 GND.n3204 GND.n3119 147.374
R25973 GND.n3200 GND.n3118 147.374
R25974 GND.n3139 GND.n3117 147.374
R25975 GND.n8729 GND.n1062 147.374
R25976 GND.n8723 GND.n1063 147.374
R25977 GND.n8719 GND.n1064 147.374
R25978 GND.n8715 GND.n1065 147.374
R25979 GND.n8711 GND.n1066 147.374
R25980 GND.n8707 GND.n1067 147.374
R25981 GND.n8703 GND.n1068 147.374
R25982 GND.n8699 GND.n1069 147.374
R25983 GND.n8498 GND.n8440 147.374
R25984 GND.n8470 GND.n8439 147.374
R25985 GND.n8466 GND.n8438 147.374
R25986 GND.n8462 GND.n8437 147.374
R25987 GND.n8458 GND.n8436 147.374
R25988 GND.n8454 GND.n8435 147.374
R25989 GND.n8450 GND.n8434 147.374
R25990 GND.n8446 GND.n8433 147.374
R25991 GND.n8442 GND.n8432 147.374
R25992 GND.n1521 GND.n1520 147.374
R25993 GND.n1518 GND.n1517 147.374
R25994 GND.n1513 GND.n1512 147.374
R25995 GND.n1510 GND.n1509 147.374
R25996 GND.n1505 GND.n1504 147.374
R25997 GND.n1502 GND.n1501 147.374
R25998 GND.n1497 GND.n1496 147.374
R25999 GND.n1494 GND.n1493 147.374
R26000 GND.n1489 GND.n1488 147.374
R26001 GND.n1402 GND.n1088 147.374
R26002 GND.n1398 GND.n1087 147.374
R26003 GND.n1394 GND.n1086 147.374
R26004 GND.n1390 GND.n1085 147.374
R26005 GND.n1386 GND.n1084 147.374
R26006 GND.n1382 GND.n1083 147.374
R26007 GND.n1378 GND.n1082 147.374
R26008 GND.n1374 GND.n1081 147.374
R26009 GND.n1370 GND.n1080 147.374
R26010 GND.n1319 GND.n1318 147.374
R26011 GND.n1321 GND.n1315 147.374
R26012 GND.n1328 GND.n1327 147.374
R26013 GND.n1329 GND.n1313 147.374
R26014 GND.n1336 GND.n1335 147.374
R26015 GND.n1337 GND.n1311 147.374
R26016 GND.n1344 GND.n1343 147.374
R26017 GND.n1347 GND.n1346 147.374
R26018 GND.n1182 GND.n1079 147.374
R26019 GND.n1178 GND.n1078 147.374
R26020 GND.n1174 GND.n1077 147.374
R26021 GND.n1170 GND.n1076 147.374
R26022 GND.n1166 GND.n1075 147.374
R26023 GND.n1162 GND.n1074 147.374
R26024 GND.n1158 GND.n1073 147.374
R26025 GND.n1154 GND.n1072 147.374
R26026 GND.n1093 GND.n1071 147.374
R26027 GND.n9200 GND.n9199 147.374
R26028 GND.n9194 GND.n9141 147.374
R26029 GND.n9192 GND.n9191 147.374
R26030 GND.n9187 GND.n9186 147.374
R26031 GND.n9184 GND.n9183 147.374
R26032 GND.n9179 GND.n9178 147.374
R26033 GND.n9176 GND.n9175 147.374
R26034 GND.n9171 GND.n9170 147.374
R26035 GND.n9134 GND.n426 147.374
R26036 GND.n9126 GND.n418 147.374
R26037 GND.n9122 GND.n419 147.374
R26038 GND.n9118 GND.n420 147.374
R26039 GND.n9114 GND.n421 147.374
R26040 GND.n9110 GND.n422 147.374
R26041 GND.n9106 GND.n423 147.374
R26042 GND.n9102 GND.n424 147.374
R26043 GND.n9679 GND.n9678 147.374
R26044 GND.n9672 GND.n9622 147.374
R26045 GND.n9668 GND.n9623 147.374
R26046 GND.n9664 GND.n9624 147.374
R26047 GND.n9660 GND.n9625 147.374
R26048 GND.n9656 GND.n9626 147.374
R26049 GND.n9652 GND.n9627 147.374
R26050 GND.n9648 GND.n9628 147.374
R26051 GND.n9478 GND.n9465 147.374
R26052 GND.n9482 GND.n9466 147.374
R26053 GND.n9486 GND.n9467 147.374
R26054 GND.n9490 GND.n9468 147.374
R26055 GND.n9494 GND.n9469 147.374
R26056 GND.n9498 GND.n9470 147.374
R26057 GND.n9472 GND.n9471 147.374
R26058 GND.n9504 GND.n188 147.374
R26059 GND.n9690 GND.n9689 147.374
R26060 GND.n130 GND.n129 147.374
R26061 GND.n9545 GND.n9543 147.374
R26062 GND.n9552 GND.n9551 147.374
R26063 GND.n9555 GND.n9554 147.374
R26064 GND.n9733 GND.n98 147.374
R26065 GND.n9721 GND.n92 147.374
R26066 GND.n9718 GND.n93 147.374
R26067 GND.n9714 GND.n94 147.374
R26068 GND.n159 GND.n150 147.374
R26069 GND.n9597 GND.n9596 147.374
R26070 GND.n140 GND.n136 147.374
R26071 GND.n148 GND.n139 147.374
R26072 GND.n141 GND.n138 147.374
R26073 GND.n8094 GND.n8093 147.374
R26074 GND.n8088 GND.n8035 147.374
R26075 GND.n8086 GND.n8085 147.374
R26076 GND.n8081 GND.n8080 147.374
R26077 GND.n8078 GND.n8077 147.374
R26078 GND.n8073 GND.n8072 147.374
R26079 GND.n8070 GND.n8069 147.374
R26080 GND.n8065 GND.n8064 147.374
R26081 GND.n4570 GND.n4569 147.374
R26082 GND.n4576 GND.n4575 147.374
R26083 GND.n4577 GND.n4564 147.374
R26084 GND.n4584 GND.n4583 147.374
R26085 GND.n4585 GND.n4562 147.374
R26086 GND.n4592 GND.n4591 147.374
R26087 GND.n4593 GND.n4560 147.374
R26088 GND.n4600 GND.n4599 147.374
R26089 GND.n616 GND.n577 147.374
R26090 GND.n589 GND.n578 147.374
R26091 GND.n593 GND.n579 147.374
R26092 GND.n597 GND.n580 147.374
R26093 GND.n601 GND.n581 147.374
R26094 GND.n605 GND.n582 147.374
R26095 GND.n609 GND.n583 147.374
R26096 GND.n585 GND.n584 147.374
R26097 GND.n651 GND.n640 147.374
R26098 GND.n655 GND.n641 147.374
R26099 GND.n659 GND.n642 147.374
R26100 GND.n663 GND.n643 147.374
R26101 GND.n667 GND.n644 147.374
R26102 GND.n671 GND.n645 147.374
R26103 GND.n647 GND.n646 147.374
R26104 GND.n677 GND.n565 147.374
R26105 GND.n8028 GND.n2128 147.374
R26106 GND.n8020 GND.n2120 147.374
R26107 GND.n8016 GND.n2121 147.374
R26108 GND.n8012 GND.n2122 147.374
R26109 GND.n8008 GND.n2123 147.374
R26110 GND.n8004 GND.n2124 147.374
R26111 GND.n8000 GND.n2125 147.374
R26112 GND.n7996 GND.n2126 147.374
R26113 GND.n7759 GND.n7749 147.374
R26114 GND.n7763 GND.n7750 147.374
R26115 GND.n7767 GND.n7751 147.374
R26116 GND.n7771 GND.n7752 147.374
R26117 GND.n7775 GND.n7753 147.374
R26118 GND.n7779 GND.n7754 147.374
R26119 GND.n7783 GND.n7755 147.374
R26120 GND.n7757 GND.n7756 147.374
R26121 GND.n7985 GND.n2142 147.374
R26122 GND.n2195 GND.n2139 147.374
R26123 GND.n7823 GND.n7820 147.374
R26124 GND.n7830 GND.n7829 147.374
R26125 GND.n7833 GND.n7832 147.374
R26126 GND.n7954 GND.n2182 147.374
R26127 GND.n7942 GND.n2176 147.374
R26128 GND.n7939 GND.n2177 147.374
R26129 GND.n7935 GND.n2178 147.374
R26130 GND.n7864 GND.n2226 147.374
R26131 GND.n2247 GND.n2225 147.374
R26132 GND.n2238 GND.n2224 147.374
R26133 GND.n2236 GND.n2223 147.374
R26134 GND.n2232 GND.n2222 147.374
R26135 GND.n7112 GND.n7111 147.374
R26136 GND.n7107 GND.n7069 147.374
R26137 GND.n7103 GND.n7068 147.374
R26138 GND.n7099 GND.n7067 147.374
R26139 GND.n7095 GND.n7066 147.374
R26140 GND.n7091 GND.n7065 147.374
R26141 GND.n7087 GND.n7064 147.374
R26142 GND.n7083 GND.n7063 147.374
R26143 GND.n2578 GND.n2577 147.374
R26144 GND.n2584 GND.n2583 147.374
R26145 GND.n2587 GND.n2586 147.374
R26146 GND.n2592 GND.n2591 147.374
R26147 GND.n2595 GND.n2594 147.374
R26148 GND.n2600 GND.n2599 147.374
R26149 GND.n2603 GND.n2602 147.374
R26150 GND.n2608 GND.n2607 147.374
R26151 GND.n6706 GND.n6695 147.374
R26152 GND.n6710 GND.n6696 147.374
R26153 GND.n6714 GND.n6697 147.374
R26154 GND.n6718 GND.n6698 147.374
R26155 GND.n6722 GND.n6699 147.374
R26156 GND.n6725 GND.n6700 147.374
R26157 GND.n6730 GND.n6729 147.374
R26158 GND.n7115 GND.n7114 147.374
R26159 GND.n7363 GND.n7362 147.374
R26160 GND.n7360 GND.n2532 147.374
R26161 GND.n7356 GND.n7355 147.374
R26162 GND.n7349 GND.n2534 147.374
R26163 GND.n7348 GND.n7347 147.374
R26164 GND.n7341 GND.n2536 147.374
R26165 GND.n7340 GND.n7339 147.374
R26166 GND.n7333 GND.n2538 147.374
R26167 GND.n6903 GND.n6902 147.374
R26168 GND.n6898 GND.n6869 147.374
R26169 GND.n6894 GND.n6868 147.374
R26170 GND.n6890 GND.n6867 147.374
R26171 GND.n6886 GND.n6866 147.374
R26172 GND.n6882 GND.n6865 147.374
R26173 GND.n6878 GND.n6864 147.374
R26174 GND.n6874 GND.n6863 147.374
R26175 GND.n7551 GND.n7550 147.374
R26176 GND.n7545 GND.n2454 147.374
R26177 GND.n7542 GND.n2455 147.374
R26178 GND.n7538 GND.n2456 147.374
R26179 GND.n7534 GND.n2457 147.374
R26180 GND.n7530 GND.n2458 147.374
R26181 GND.n7526 GND.n2459 147.374
R26182 GND.n7522 GND.n2460 147.374
R26183 GND.n7362 GND.n7361 147.374
R26184 GND.n7357 GND.n2532 147.374
R26185 GND.n7355 GND.n7354 147.374
R26186 GND.n7350 GND.n7349 147.374
R26187 GND.n7347 GND.n7346 147.374
R26188 GND.n7342 GND.n7341 147.374
R26189 GND.n7339 GND.n7338 147.374
R26190 GND.n7334 GND.n7333 147.374
R26191 GND.n7114 GND.n6692 147.374
R26192 GND.n6730 GND.n6701 147.374
R26193 GND.n6723 GND.n6700 147.374
R26194 GND.n6719 GND.n6699 147.374
R26195 GND.n6715 GND.n6698 147.374
R26196 GND.n6711 GND.n6697 147.374
R26197 GND.n6707 GND.n6696 147.374
R26198 GND.n6703 GND.n6695 147.374
R26199 GND.n2579 GND.n2578 147.374
R26200 GND.n2585 GND.n2584 147.374
R26201 GND.n2586 GND.n2573 147.374
R26202 GND.n2593 GND.n2592 147.374
R26203 GND.n2594 GND.n2571 147.374
R26204 GND.n2601 GND.n2600 147.374
R26205 GND.n2602 GND.n2569 147.374
R26206 GND.n2609 GND.n2608 147.374
R26207 GND.n7086 GND.n7063 147.374
R26208 GND.n7090 GND.n7064 147.374
R26209 GND.n7094 GND.n7065 147.374
R26210 GND.n7098 GND.n7066 147.374
R26211 GND.n7102 GND.n7067 147.374
R26212 GND.n7106 GND.n7068 147.374
R26213 GND.n7071 GND.n7069 147.374
R26214 GND.n7112 GND.n7070 147.374
R26215 GND.n7551 GND.n2463 147.374
R26216 GND.n7543 GND.n2454 147.374
R26217 GND.n7539 GND.n2455 147.374
R26218 GND.n7535 GND.n2456 147.374
R26219 GND.n7531 GND.n2457 147.374
R26220 GND.n7527 GND.n2458 147.374
R26221 GND.n7523 GND.n2459 147.374
R26222 GND.n7519 GND.n2460 147.374
R26223 GND.n8366 GND.n1817 147.374
R26224 GND.n8370 GND.n1818 147.374
R26225 GND.n8374 GND.n1819 147.374
R26226 GND.n8378 GND.n1820 147.374
R26227 GND.n8382 GND.n1821 147.374
R26228 GND.n8386 GND.n1822 147.374
R26229 GND.n8390 GND.n1823 147.374
R26230 GND.n1826 GND.n1824 147.374
R26231 GND.n4313 GND.n4312 147.374
R26232 GND.n4308 GND.n4277 147.374
R26233 GND.n4306 GND.n4305 147.374
R26234 GND.n4301 GND.n4300 147.374
R26235 GND.n4298 GND.n4297 147.374
R26236 GND.n4293 GND.n4292 147.374
R26237 GND.n4290 GND.n4289 147.374
R26238 GND.n4285 GND.n4284 147.374
R26239 GND.n5405 GND.n4983 147.374
R26240 GND.n5409 GND.n4984 147.374
R26241 GND.n5413 GND.n4985 147.374
R26242 GND.n5417 GND.n4986 147.374
R26243 GND.n5421 GND.n4987 147.374
R26244 GND.n5425 GND.n4988 147.374
R26245 GND.n5429 GND.n4989 147.374
R26246 GND.n5433 GND.n4990 147.374
R26247 GND.n5024 GND.n4991 147.374
R26248 GND.n5020 GND.n4992 147.374
R26249 GND.n5016 GND.n4993 147.374
R26250 GND.n5694 GND.n4994 147.374
R26251 GND.n5698 GND.n4995 147.374
R26252 GND.n5702 GND.n4996 147.374
R26253 GND.n5706 GND.n4997 147.374
R26254 GND.n5710 GND.n4998 147.374
R26255 GND.n5714 GND.n4999 147.374
R26256 GND.n5718 GND.n5000 147.374
R26257 GND.n5722 GND.n5001 147.374
R26258 GND.n5003 GND.n5002 147.374
R26259 GND.n5728 GND.n3905 147.374
R26260 GND.n5099 GND.n5098 147.374
R26261 GND.n5105 GND.n5104 147.374
R26262 GND.n5106 GND.n5093 147.374
R26263 GND.n5113 GND.n5112 147.374
R26264 GND.n5114 GND.n5091 147.374
R26265 GND.n5121 GND.n5120 147.374
R26266 GND.n5122 GND.n5089 147.374
R26267 GND.n5129 GND.n5128 147.374
R26268 GND.n5130 GND.n5046 147.374
R26269 GND.n5143 GND.n5142 147.374
R26270 GND.n5144 GND.n5042 147.374
R26271 GND.n5155 GND.n5154 147.374
R26272 GND.n5157 GND.n5156 147.374
R26273 GND.n5038 GND.n5035 147.374
R26274 GND.n5344 GND.n5343 147.374
R26275 GND.n5345 GND.n5033 147.374
R26276 GND.n5352 GND.n5351 147.374
R26277 GND.n5353 GND.n5031 147.374
R26278 GND.n5360 GND.n5359 147.374
R26279 GND.n5361 GND.n5029 147.374
R26280 GND.n5368 GND.n5367 147.374
R26281 GND.n4115 GND.n3906 147.374
R26282 GND.n4119 GND.n3907 147.374
R26283 GND.n4123 GND.n3908 147.374
R26284 GND.n4127 GND.n3909 147.374
R26285 GND.n4131 GND.n3910 147.374
R26286 GND.n4135 GND.n3911 147.374
R26287 GND.n4139 GND.n3912 147.374
R26288 GND.n4143 GND.n3913 147.374
R26289 GND.n4147 GND.n3914 147.374
R26290 GND.n3948 GND.n3915 147.374
R26291 GND.n3944 GND.n3916 147.374
R26292 GND.n3940 GND.n3917 147.374
R26293 GND.n4948 GND.n3918 147.374
R26294 GND.n4952 GND.n3919 147.374
R26295 GND.n4956 GND.n3920 147.374
R26296 GND.n4960 GND.n3921 147.374
R26297 GND.n4964 GND.n3922 147.374
R26298 GND.n4968 GND.n3923 147.374
R26299 GND.n4972 GND.n3924 147.374
R26300 GND.n4976 GND.n3925 147.374
R26301 GND.n3927 GND.n3926 147.374
R26302 GND.n5808 GND.n3839 147.374
R26303 GND.n5800 GND.n3818 147.374
R26304 GND.n5796 GND.n3819 147.374
R26305 GND.n5792 GND.n3820 147.374
R26306 GND.n5788 GND.n3821 147.374
R26307 GND.n5784 GND.n3822 147.374
R26308 GND.n3823 GND.n3816 147.374
R26309 GND.n5810 GND.n3817 147.374
R26310 GND.n4021 GND.n3824 147.374
R26311 GND.n4027 GND.n3825 147.374
R26312 GND.n4033 GND.n3826 147.374
R26313 GND.n4039 GND.n3827 147.374
R26314 GND.n4046 GND.n3828 147.374
R26315 GND.n4050 GND.n3829 147.374
R26316 GND.n4054 GND.n3830 147.374
R26317 GND.n4058 GND.n3831 147.374
R26318 GND.n4062 GND.n3832 147.374
R26319 GND.n4066 GND.n3833 147.374
R26320 GND.n4070 GND.n3834 147.374
R26321 GND.n4074 GND.n3835 147.374
R26322 GND.n4078 GND.n3836 147.374
R26323 GND.n5313 GND.n5312 147.374
R26324 GND.n5172 GND.n5170 147.374
R26325 GND.n5320 GND.n5319 147.374
R26326 GND.n5169 GND.n5167 147.374
R26327 GND.n5327 GND.n5326 147.374
R26328 GND.n5166 GND.n5164 147.374
R26329 GND.n5334 GND.n5333 147.374
R26330 GND.n5337 GND.n5336 147.374
R26331 GND.n5161 GND.n5160 147.374
R26332 GND.n5151 GND.n5150 147.374
R26333 GND.n5148 GND.n5147 147.374
R26334 GND.n5139 GND.n5138 147.374
R26335 GND.n5136 GND.n5135 147.374
R26336 GND.n5085 GND.n5084 147.374
R26337 GND.n5082 GND.n5081 147.374
R26338 GND.n5077 GND.n5076 147.374
R26339 GND.n5074 GND.n5073 147.374
R26340 GND.n5069 GND.n5068 147.374
R26341 GND.n5066 GND.n5065 147.374
R26342 GND.n5061 GND.n5060 147.374
R26343 GND.n5058 GND.n5057 147.374
R26344 GND.n5195 GND.n5194 147.374
R26345 GND.n5201 GND.n5200 147.374
R26346 GND.n5202 GND.n5191 147.374
R26347 GND.n5209 GND.n5208 147.374
R26348 GND.n5210 GND.n5189 147.374
R26349 GND.n5217 GND.n5216 147.374
R26350 GND.n5218 GND.n5187 147.374
R26351 GND.n5225 GND.n5224 147.374
R26352 GND.n5226 GND.n5185 147.374
R26353 GND.n5233 GND.n5232 147.374
R26354 GND.n5234 GND.n5183 147.374
R26355 GND.n5241 GND.n5240 147.374
R26356 GND.n5242 GND.n5181 147.374
R26357 GND.n5249 GND.n5248 147.374
R26358 GND.n5250 GND.n5179 147.374
R26359 GND.n5257 GND.n5256 147.374
R26360 GND.n5258 GND.n5177 147.374
R26361 GND.n5265 GND.n5264 147.374
R26362 GND.n5266 GND.n5175 147.374
R26363 GND.n5273 GND.n5272 147.374
R26364 GND.n5276 GND.n5275 147.374
R26365 GND.n3985 GND.n3790 147.374
R26366 GND.n3989 GND.n3791 147.374
R26367 GND.n3993 GND.n3792 147.374
R26368 GND.n3997 GND.n3793 147.374
R26369 GND.n4001 GND.n3794 147.374
R26370 GND.n4005 GND.n3795 147.374
R26371 GND.n4009 GND.n3796 147.374
R26372 GND.n4013 GND.n3797 147.374
R26373 GND.n4042 GND.n3798 147.374
R26374 GND.n4036 GND.n3799 147.374
R26375 GND.n4030 GND.n3800 147.374
R26376 GND.n4024 GND.n3801 147.374
R26377 GND.n4018 GND.n3802 147.374
R26378 GND.n5815 GND.n3803 147.374
R26379 GND.n5819 GND.n3804 147.374
R26380 GND.n5823 GND.n3805 147.374
R26381 GND.n5827 GND.n3806 147.374
R26382 GND.n5831 GND.n3807 147.374
R26383 GND.n5835 GND.n3808 147.374
R26384 GND.n5839 GND.n3809 147.374
R26385 GND.n3812 GND.n3810 147.374
R26386 GND.n5981 GND.n3719 147.374
R26387 GND.n5973 GND.n3697 147.374
R26388 GND.n5969 GND.n3698 147.374
R26389 GND.n5965 GND.n3699 147.374
R26390 GND.n5961 GND.n3700 147.374
R26391 GND.n5957 GND.n3701 147.374
R26392 GND.n5953 GND.n3702 147.374
R26393 GND.n5949 GND.n3703 147.374
R26394 GND.n5945 GND.n3704 147.374
R26395 GND.n5941 GND.n3705 147.374
R26396 GND.n5937 GND.n3706 147.374
R26397 GND.n5933 GND.n3707 147.374
R26398 GND.n5929 GND.n3708 147.374
R26399 GND.n5925 GND.n3709 147.374
R26400 GND.n5921 GND.n3710 147.374
R26401 GND.n5917 GND.n3711 147.374
R26402 GND.n5913 GND.n3712 147.374
R26403 GND.n5909 GND.n3713 147.374
R26404 GND.n5905 GND.n3714 147.374
R26405 GND.n5901 GND.n3715 147.374
R26406 GND.n5897 GND.n3716 147.374
R26407 GND.n2733 GND.n2731 147.374
R26408 GND.n6396 GND.n6395 147.374
R26409 GND.n2730 GND.n2728 147.374
R26410 GND.n6403 GND.n6402 147.374
R26411 GND.n2727 GND.n2725 147.374
R26412 GND.n6410 GND.n6409 147.374
R26413 GND.n2724 GND.n2722 147.374
R26414 GND.n6417 GND.n6416 147.374
R26415 GND.n6420 GND.n6419 147.374
R26416 GND.n6336 GND.n6335 147.374
R26417 GND.n6344 GND.n6343 147.374
R26418 GND.n6347 GND.n6346 147.374
R26419 GND.n6332 GND.n6326 147.374
R26420 GND.n6359 GND.n6358 147.374
R26421 GND.n6325 GND.n6323 147.374
R26422 GND.n6366 GND.n6365 147.374
R26423 GND.n6322 GND.n6320 147.374
R26424 GND.n6373 GND.n6372 147.374
R26425 GND.n6319 GND.n6317 147.374
R26426 GND.n6380 GND.n6379 147.374
R26427 GND.n6383 GND.n6382 147.374
R26428 GND.n6261 GND.n2770 147.374
R26429 GND.n6255 GND.n2772 147.374
R26430 GND.n6251 GND.n2773 147.374
R26431 GND.n6247 GND.n2774 147.374
R26432 GND.n6243 GND.n2775 147.374
R26433 GND.n6239 GND.n2776 147.374
R26434 GND.n6235 GND.n2777 147.374
R26435 GND.n2794 GND.n2778 147.374
R26436 GND.n2799 GND.n2779 147.374
R26437 GND.n2801 GND.n2780 147.374
R26438 GND.n2806 GND.n2781 147.374
R26439 GND.n2808 GND.n2782 147.374
R26440 GND.n2845 GND.n2783 147.374
R26441 GND.n2841 GND.n2784 147.374
R26442 GND.n2837 GND.n2785 147.374
R26443 GND.n2833 GND.n2786 147.374
R26444 GND.n2829 GND.n2787 147.374
R26445 GND.n2825 GND.n2788 147.374
R26446 GND.n2821 GND.n2789 147.374
R26447 GND.n2817 GND.n2790 147.374
R26448 GND.n2813 GND.n2791 147.374
R26449 GND.n6187 GND.n6186 147.374
R26450 GND.n2858 GND.n2856 147.374
R26451 GND.n6194 GND.n6193 147.374
R26452 GND.n2855 GND.n2853 147.374
R26453 GND.n6201 GND.n6200 147.374
R26454 GND.n2852 GND.n2850 147.374
R26455 GND.n6208 GND.n6207 147.374
R26456 GND.n2849 GND.n2812 147.374
R26457 GND.n6215 GND.n6214 147.374
R26458 GND.n2811 GND.n2805 147.374
R26459 GND.n6222 GND.n6221 147.374
R26460 GND.n2804 GND.n2798 147.374
R26461 GND.n6229 GND.n6228 147.374
R26462 GND.n6149 GND.n2797 147.374
R26463 GND.n6153 GND.n6152 147.374
R26464 GND.n6148 GND.n6146 147.374
R26465 GND.n6160 GND.n6159 147.374
R26466 GND.n6145 GND.n6143 147.374
R26467 GND.n6167 GND.n6166 147.374
R26468 GND.n6142 GND.n6140 147.374
R26469 GND.n6174 GND.n6173 147.374
R26470 GND.n6088 GND.n6087 147.374
R26471 GND.n6082 GND.n5988 147.374
R26472 GND.n6080 GND.n6079 147.374
R26473 GND.n6075 GND.n6074 147.374
R26474 GND.n6072 GND.n6071 147.374
R26475 GND.n6067 GND.n6066 147.374
R26476 GND.n6064 GND.n6063 147.374
R26477 GND.n6059 GND.n6058 147.374
R26478 GND.n6056 GND.n6055 147.374
R26479 GND.n6051 GND.n6050 147.374
R26480 GND.n6048 GND.n6047 147.374
R26481 GND.n6043 GND.n6042 147.374
R26482 GND.n6040 GND.n6039 147.374
R26483 GND.n6035 GND.n6034 147.374
R26484 GND.n6032 GND.n6031 147.374
R26485 GND.n6027 GND.n6026 147.374
R26486 GND.n6024 GND.n6023 147.374
R26487 GND.n6019 GND.n6018 147.374
R26488 GND.n6016 GND.n6015 147.374
R26489 GND.n6011 GND.n6010 147.374
R26490 GND.n6008 GND.n3116 147.374
R26491 GND.n7584 GND.n7583 147.374
R26492 GND.n5567 GND.n2411 147.374
R26493 GND.n5571 GND.n2412 147.374
R26494 GND.n5575 GND.n2413 147.374
R26495 GND.n5579 GND.n2414 147.374
R26496 GND.n5583 GND.n2415 147.374
R26497 GND.n5587 GND.n2416 147.374
R26498 GND.n5590 GND.n2417 147.374
R26499 GND.n7653 GND.n2317 147.374
R26500 GND.n7657 GND.n2318 147.374
R26501 GND.n7661 GND.n2319 147.374
R26502 GND.n7665 GND.n2320 147.374
R26503 GND.n7669 GND.n2321 147.374
R26504 GND.n7673 GND.n2322 147.374
R26505 GND.n7677 GND.n2323 147.374
R26506 GND.n2326 GND.n2324 147.374
R26507 GND.n5621 GND.n5617 147.374
R26508 GND.n5623 GND.n5557 147.374
R26509 GND.n5548 GND.n5547 147.374
R26510 GND.n5535 GND.n5534 147.374
R26511 GND.n5531 GND.n2340 147.374
R26512 GND.n5478 GND.n5477 147.374
R26513 GND.n5480 GND.n5467 147.374
R26514 GND.n5636 GND.n5635 147.374
R26515 GND.n5639 GND.n5638 147.374
R26516 GND.n5516 GND.n5515 147.374
R26517 GND.n5523 GND.n5522 147.374
R26518 GND.n5493 GND.n5489 147.374
R26519 GND.n5499 GND.n5492 147.374
R26520 GND.n5491 GND.n2360 147.374
R26521 GND.n6877 GND.n6863 147.374
R26522 GND.n6881 GND.n6864 147.374
R26523 GND.n6885 GND.n6865 147.374
R26524 GND.n6889 GND.n6866 147.374
R26525 GND.n6893 GND.n6867 147.374
R26526 GND.n6897 GND.n6868 147.374
R26527 GND.n6871 GND.n6869 147.374
R26528 GND.n6903 GND.n6870 147.374
R26529 GND.n7495 GND.n7494 147.374
R26530 GND.n7462 GND.n7455 147.374
R26531 GND.n7487 GND.n7456 147.374
R26532 GND.n7483 GND.n7457 147.374
R26533 GND.n7479 GND.n7458 147.374
R26534 GND.n7475 GND.n7459 147.374
R26535 GND.n7471 GND.n7460 147.374
R26536 GND.n7467 GND.n7461 147.374
R26537 GND.n6840 GND.n6804 147.374
R26538 GND.n6839 GND.n6838 147.374
R26539 GND.n6832 GND.n6806 147.374
R26540 GND.n6831 GND.n6830 147.374
R26541 GND.n6824 GND.n6808 147.374
R26542 GND.n6823 GND.n6822 147.374
R26543 GND.n6816 GND.n6810 147.374
R26544 GND.n6815 GND.n6814 147.374
R26545 GND.n6814 GND.n6813 147.374
R26546 GND.n6817 GND.n6816 147.374
R26547 GND.n6822 GND.n6821 147.374
R26548 GND.n6825 GND.n6824 147.374
R26549 GND.n6830 GND.n6829 147.374
R26550 GND.n6833 GND.n6832 147.374
R26551 GND.n6838 GND.n6837 147.374
R26552 GND.n6841 GND.n6840 147.374
R26553 GND.n7494 GND.n7454 147.374
R26554 GND.n7488 GND.n7455 147.374
R26555 GND.n7484 GND.n7456 147.374
R26556 GND.n7480 GND.n7457 147.374
R26557 GND.n7476 GND.n7458 147.374
R26558 GND.n7472 GND.n7459 147.374
R26559 GND.n7468 GND.n7460 147.374
R26560 GND.n7464 GND.n7461 147.374
R26561 GND.n8426 GND.n1803 146.825
R26562 GND.n14 GND.n11 146.25
R26563 GND.n2114 GND.n14 146.25
R26564 GND.n13 GND.n12 146.25
R26565 GND.n2114 GND.n13 146.25
R26566 GND.n2311 GND.n2309 146.25
R26567 GND.n7691 GND.n2309 146.25
R26568 GND.n2310 GND.n2308 146.25
R26569 GND.n7691 GND.n2308 146.25
R26570 GND.n9797 GND.n9796 141.834
R26571 GND.n7723 GND.n2298 141.766
R26572 GND.n7708 GND.n7707 141.766
R26573 GND.n9456 GND.n9455 141.766
R26574 GND.n9445 GND.n9444 141.766
R26575 GND.n7734 GND.t82 138.244
R26576 GND.t70 GND.n16 138.201
R26577 GND.n9432 GND.t153 134.816
R26578 GND.t418 GND.t427 131.518
R26579 GND.t105 GND.t57 131.518
R26580 GND.t57 GND.t418 131.518
R26581 GND.t20 GND.t427 131.518
R26582 GND.n7748 GND.n2273 126.046
R26583 GND.t81 GND.n25 125.581
R26584 GND.n2119 GND.t341 125.493
R26585 GND.n9820 GND.t290 125.493
R26586 GND.t311 GND.n15 125.493
R26587 GND.n9451 GND.t7 125.493
R26588 GND.n9452 GND.t17 125.493
R26589 GND.n9462 GND.t16 125.493
R26590 GND.n7692 GND.t286 125.493
R26591 GND.n7702 GND.t348 125.493
R26592 GND.n7704 GND.t288 125.493
R26593 GND.n7714 GND.t26 125.493
R26594 GND.t0 GND.n7715 125.493
R26595 GND.t314 GND.n7716 125.493
R26596 GND.t376 GND.n7747 114.344
R26597 GND.n7690 GND.n7689 113.591
R26598 GND.t409 GND.t104 112.284
R26599 GND.t163 GND.t357 112.284
R26600 GND.t104 GND.t163 112.284
R26601 GND.t152 GND.t409 112.284
R26602 GND.n7722 GND.n2299 111.918
R26603 GND.n7711 GND.n2305 111.918
R26604 GND.n9459 GND.n9436 111.918
R26605 GND.n9448 GND.n9441 111.918
R26606 GND.n9787 GND.n9786 109.177
R26607 GND.t105 GND.n17 97.2365
R26608 GND.n9818 GND.n16 96.6695
R26609 GND.n6093 GND.n5984 94.0436
R26610 GND.n2863 GND.n2771 94.0436
R26611 GND.n6260 GND.n2767 94.0436
R26612 GND.n6388 GND.n2720 94.0436
R26613 GND.n2998 GND.t145 87.4177
R26614 GND.n9452 GND.n9451 83.6625
R26615 GND.n7715 GND.n7714 83.6625
R26616 GND.n754 GND.n231 82.4476
R26617 GND.n9342 GND.n293 82.4476
R26618 GND.n789 GND.n785 82.4476
R26619 GND.n9313 GND.n320 82.4476
R26620 GND.n794 GND.n524 82.4476
R26621 GND.n854 GND.n853 82.4476
R26622 GND.n9349 GND.n9348 82.4476
R26623 GND.n9012 GND.n9011 82.4476
R26624 GND.n4367 GND.n1923 82.4476
R26625 GND.n8236 GND.n1985 82.4476
R26626 GND.n4401 GND.n4400 82.4476
R26627 GND.n8207 GND.n2012 82.4476
R26628 GND.n4446 GND.n4444 82.4476
R26629 GND.n4438 GND.n4437 82.4476
R26630 GND.n8243 GND.n8242 82.4476
R26631 GND.n4755 GND.n4754 82.4476
R26632 GND.n7138 GND.n6679 82.4476
R26633 GND.n7084 GND.n7082 82.4476
R26634 GND.n2576 GND.n2523 82.4476
R26635 GND.n2611 GND.n2568 82.4476
R26636 GND.n6702 GND.n6687 82.4476
R26637 GND.n7117 GND.n7116 82.4476
R26638 GND.n7365 GND.n7364 82.4476
R26639 GND.n7330 GND.n2539 82.4476
R26640 GND.n5615 GND.n5614 80.9417
R26641 GND.n5619 GND.n2394 80.9417
R26642 GND.n7637 GND.n2342 80.9417
R26643 GND.n5545 GND.n5544 80.9417
R26644 GND.n9614 GND.n9613 80.9417
R26645 GND.n9693 GND.n9692 80.9417
R26646 GND.n9557 GND.n9556 80.9417
R26647 GND.n9547 GND.n169 80.9417
R26648 GND.n2198 GND.n2197 80.9417
R26649 GND.n7983 GND.n2144 80.9417
R26650 GND.n7835 GND.n7834 80.9417
R26651 GND.n7825 GND.n7822 80.9417
R26652 GND.n613 GND.n571 80.5652
R26653 GND.n619 GND.n618 80.5652
R26654 GND.n9203 GND.n9202 80.5652
R26655 GND.n9172 GND.n9169 80.5652
R26656 GND.n8394 GND.n1827 80.5652
R26657 GND.n8364 GND.n1828 80.5652
R26658 GND.n8097 GND.n8096 80.5652
R26659 GND.n8066 GND.n8063 80.5652
R26660 GND.n6844 GND.n6843 80.5652
R26661 GND.n6848 GND.n6800 80.5652
R26662 GND.n7497 GND.n7496 80.5652
R26663 GND.n7465 GND.n7463 80.5652
R26664 GND.n5552 GND.t424 79.0275
R26665 GND.n131 GND.t331 79.0275
R26666 GND.n2147 GND.t304 79.0275
R26667 GND.n5627 GND.t402 79.027
R26668 GND.n9606 GND.t262 79.027
R26669 GND.n7979 GND.t282 79.027
R26670 GND.n5848 GND.n3785 78.3064
R26671 GND.n5892 GND.n3728 78.3064
R26672 GND.n5278 GND.n5277 78.3064
R26673 GND.n5310 GND.n5309 78.3064
R26674 GND.n5370 GND.n5028 78.3064
R26675 GND.n5096 GND.n3849 78.3064
R26676 GND.n5732 GND.n5731 78.3064
R26677 GND.n5403 GND.n5399 78.3064
R26678 GND.n6177 GND.n6176 78.3064
R26679 GND.n6091 GND.n6090 78.3064
R26680 GND.n6095 GND.n3115 78.3064
R26681 GND.n6184 GND.n6183 78.3064
R26682 GND.n6391 GND.n2732 78.3064
R26683 GND.n2814 GND.n2765 78.3064
R26684 GND.n6264 GND.n6263 78.3064
R26685 GND.n6386 GND.n6385 78.3064
R26686 GND.n1186 GND.n1185 78.3064
R26687 GND.n1650 GND.n1095 78.3064
R26688 GND.n1528 GND.n1287 78.3064
R26689 GND.n1350 GND.n1349 78.3064
R26690 GND.n1490 GND.n1487 78.3064
R26691 GND.n1524 GND.n1523 78.3064
R26692 GND.n1371 GND.n1369 78.3064
R26693 GND.n1406 GND.n1405 78.3064
R26694 GND.n8496 GND.n8495 78.3064
R26695 GND.n8443 GND.n1793 78.3064
R26696 GND.n8732 GND.n8731 78.3064
R26697 GND.n8698 GND.n8697 78.3064
R26698 GND.n1720 GND.n1055 78.3064
R26699 GND.n8592 GND.n8591 78.3064
R26700 GND.n8561 GND.n8557 78.3064
R26701 GND.n1688 GND.n1685 78.3064
R26702 GND.n3232 GND.n3231 78.3064
R26703 GND.n3693 GND.n3141 78.3064
R26704 GND.n3571 GND.n3333 78.3064
R26705 GND.n3366 GND.n3365 78.3064
R26706 GND.n3533 GND.n3530 78.3064
R26707 GND.n3567 GND.n3566 78.3064
R26708 GND.n3418 GND.n3416 78.3064
R26709 GND.n3453 GND.n3452 78.3064
R26710 GND.n5843 GND.n3813 78.3064
R26711 GND.n5979 GND.n3721 78.3064
R26712 GND.n5898 GND.n3722 78.3064
R26713 GND.n3983 GND.n3952 78.3064
R26714 GND.n4113 GND.n4110 78.3064
R26715 GND.n4081 GND.n4077 78.3064
R26716 GND.n5806 GND.n5781 78.3064
R26717 GND.n4980 GND.n3895 78.3064
R26718 GND.n6260 GND.n2771 76.6282
R26719 GND.n7587 GND.n7586 76.0476
R26720 GND.n5592 GND.n5591 76.0476
R26721 GND.n7651 GND.n2328 76.0476
R26722 GND.n7681 GND.n2327 76.0476
R26723 GND.n9683 GND.n9619 76.0476
R26724 GND.n9649 GND.n9647 76.0476
R26725 GND.n9476 GND.n9473 76.0476
R26726 GND.n9508 GND.n9507 76.0476
R26727 GND.n8026 GND.n2130 76.0476
R26728 GND.n7997 GND.n2131 76.0476
R26729 GND.n7792 GND.n2269 76.0476
R26730 GND.n7787 GND.n2266 76.0476
R26731 GND.t20 GND.t3 74.6993
R26732 GND.t352 GND.t311 74.3667
R26733 GND.t353 GND.t352 74.3667
R26734 GND.t12 GND.t353 74.3667
R26735 GND.t351 GND.t12 74.3667
R26736 GND.t351 GND.t31 74.3667
R26737 GND.t31 GND.t154 74.3667
R26738 GND.t154 GND.t53 74.3667
R26739 GND.t53 GND.t7 74.3667
R26740 GND.t17 GND.t150 74.3667
R26741 GND.t150 GND.t263 74.3667
R26742 GND.t263 GND.t49 74.3667
R26743 GND.t49 GND.t48 74.3667
R26744 GND.t48 GND.t340 74.3667
R26745 GND.t340 GND.t431 74.3667
R26746 GND.t431 GND.t343 74.3667
R26747 GND.t343 GND.t16 74.3667
R26748 GND.t288 GND.t223 74.3667
R26749 GND.t223 GND.t350 74.3667
R26750 GND.t350 GND.t27 74.3667
R26751 GND.t27 GND.t205 74.3667
R26752 GND.t205 GND.t28 74.3667
R26753 GND.t28 GND.t289 74.3667
R26754 GND.t289 GND.t204 74.3667
R26755 GND.t204 GND.t26 74.3667
R26756 GND.t336 GND.t0 74.3667
R26757 GND.t337 GND.t336 74.3667
R26758 GND.t166 GND.t337 74.3667
R26759 GND.t101 GND.t166 74.3667
R26760 GND.t101 GND.t42 74.3667
R26761 GND.t42 GND.t354 74.3667
R26762 GND.t354 GND.t159 74.3667
R26763 GND.t159 GND.t314 74.3667
R26764 GND.n681 GND.n680 73.0358
R26765 GND.n649 GND.n557 73.0358
R26766 GND.n9132 GND.n407 73.0358
R26767 GND.n9103 GND.n9100 73.0358
R26768 GND.n8351 GND.n1841 73.0358
R26769 GND.n4316 GND.n4315 73.0358
R26770 GND.n4567 GND.n2097 73.0358
R26771 GND.n4602 GND.n4559 73.0358
R26772 GND.n6915 GND.n6788 73.0358
R26773 GND.n6875 GND.n6873 73.0358
R26774 GND.n7549 GND.n2465 73.0358
R26775 GND.n7520 GND.n2466 73.0358
R26776 GND.n5628 GND.n5553 73.0311
R26777 GND.n9605 GND.n132 73.0311
R26778 GND.n7978 GND.n2148 73.0311
R26779 GND.n7623 GND.n2362 70.024
R26780 GND.n5475 GND.n5474 70.024
R26781 GND.n5642 GND.n5641 70.024
R26782 GND.n5518 GND.n5462 70.024
R26783 GND.n142 GND.n79 70.024
R26784 GND.n9731 GND.n99 70.024
R26785 GND.n9713 GND.n9712 70.024
R26786 GND.n9592 GND.n158 70.024
R26787 GND.n2233 GND.n2230 70.024
R26788 GND.n7952 GND.n2164 70.024
R26789 GND.n7934 GND.n7933 70.024
R26790 GND.n7862 GND.n7861 70.024
R26791 GND.n7493 GND.t82 62.1041
R26792 GND.t224 GND.n2273 61.3874
R26793 GND.n6093 GND.n5985 59.2128
R26794 GND.n6099 GND.n2888 59.2128
R26795 GND.n6105 GND.n2888 59.2128
R26796 GND.n6105 GND.n2884 59.2128
R26797 GND.n6111 GND.n2884 59.2128
R26798 GND.n6111 GND.n2880 59.2128
R26799 GND.n6117 GND.n2880 59.2128
R26800 GND.n6123 GND.n2876 59.2128
R26801 GND.n6123 GND.n2872 59.2128
R26802 GND.n6129 GND.n2872 59.2128
R26803 GND.n6129 GND.n2868 59.2128
R26804 GND.n6135 GND.n2868 59.2128
R26805 GND.n6135 GND.n2862 59.2128
R26806 GND.n6180 GND.n2862 59.2128
R26807 GND.n6180 GND.n2863 59.2128
R26808 GND.n6267 GND.n2767 59.2128
R26809 GND.n6267 GND.n2763 59.2128
R26810 GND.n6273 GND.n2763 59.2128
R26811 GND.n6273 GND.n2759 59.2128
R26812 GND.n6279 GND.n2759 59.2128
R26813 GND.n6279 GND.n2755 59.2128
R26814 GND.n6286 GND.n2755 59.2128
R26815 GND.n6286 GND.n6285 59.2128
R26816 GND.n6292 GND.n2748 59.2128
R26817 GND.n6298 GND.n2748 59.2128
R26818 GND.n6298 GND.n2744 59.2128
R26819 GND.n6304 GND.n2744 59.2128
R26820 GND.n6304 GND.n2740 59.2128
R26821 GND.n6311 GND.n2740 59.2128
R26822 GND.n6311 GND.n2735 59.2128
R26823 GND.n6388 GND.n2735 59.2128
R26824 GND.n2999 GND.t102 58.2786
R26825 GND.n7695 GND.n2311 55.5568
R26826 GND.n2116 GND.n11 55.5568
R26827 GND.n7747 GND.t69 54.7135
R26828 GND.n9205 GND.n50 53.8036
R26829 GND.n6846 GND.n6802 53.8036
R26830 GND.n7699 GND.n2311 53.298
R26831 GND.n9823 GND.n11 53.298
R26832 GND.n615 GND.t379 51.3116
R26833 GND.t407 GND.n8396 51.3116
R26834 GND.n3696 GND.n3695 48.9824
R26835 GND.n3569 GND.n3399 48.9824
R26836 GND.n8499 GND.n1795 48.9824
R26837 GND.n8728 GND.n1059 48.9824
R26838 GND.n1653 GND.n1652 48.9824
R26839 GND.n1526 GND.n51 48.9824
R26840 GND.n5985 GND.n3113 48.7636
R26841 GND.n2937 GND.n2931 43.9358
R26842 GND.n3102 GND.n3101 43.9358
R26843 GND.t146 GND.t14 43.7091
R26844 GND.t102 GND.t139 43.7091
R26845 GND.t63 GND.t137 43.7091
R26846 GND.t45 GND.t142 43.7091
R26847 GND.n8031 GND.t70 43.6575
R26848 GND.n2934 GND.t430 43.4788
R26849 GND.n2939 GND.n2935 42.1528
R26850 GND.n9441 GND.n9439 41.7862
R26851 GND.n9439 GND.t351 41.7862
R26852 GND.n9440 GND.n9438 41.7862
R26853 GND.t351 GND.n9438 41.7862
R26854 GND.n9436 GND.n9434 41.7862
R26855 GND.t48 GND.n9434 41.7862
R26856 GND.n9435 GND.n9433 41.7862
R26857 GND.t48 GND.n9433 41.7862
R26858 GND.n2305 GND.n2303 41.7862
R26859 GND.t205 GND.n2303 41.7862
R26860 GND.n2304 GND.n2302 41.7862
R26861 GND.t205 GND.n2302 41.7862
R26862 GND.n7722 GND.n7721 41.7862
R26863 GND.n7721 GND.t101 41.7862
R26864 GND.n7720 GND.n7719 41.7862
R26865 GND.t101 GND.n7720 41.7862
R26866 GND.t341 GND.n2114 37.1836
R26867 GND.n2114 GND.t290 37.1836
R26868 GND.t286 GND.n7691 37.1836
R26869 GND.n7691 GND.t348 37.1836
R26870 GND.n9798 GND.n48 37.1524
R26871 GND.n1810 GND.n16 37.1524
R26872 GND.n9808 GND.n27 37.1524
R26873 GND.n7734 GND.n2276 37.1524
R26874 GND.n8411 GND.n8397 37.1524
R26875 GND.n7689 GND.n2315 37.1524
R26876 GND.n2987 GND.n2962 34.6358
R26877 GND.n2987 GND.n2986 34.6358
R26878 GND.n2979 GND.n2969 34.6358
R26879 GND.n2947 GND.n2931 34.6358
R26880 GND.n2948 GND.n2947 34.6358
R26881 GND.n2948 GND.n2928 34.6358
R26882 GND.n2944 GND.n2943 34.6358
R26883 GND.n2953 GND.n2929 34.6358
R26884 GND.n2990 GND.n2961 34.6358
R26885 GND.n2983 GND.n2961 34.6358
R26886 GND.n2983 GND.n2982 34.6358
R26887 GND.n2982 GND.n2967 34.6358
R26888 GND.n2974 GND.n2967 34.6358
R26889 GND.n3016 GND.n3013 34.6358
R26890 GND.n3024 GND.n2913 34.6358
R26891 GND.n3026 GND.n2909 34.6358
R26892 GND.n3021 GND.n3019 34.6358
R26893 GND.n3021 GND.n3020 34.6358
R26894 GND.n3020 GND.n2910 34.6358
R26895 GND.n3031 GND.n2910 34.6358
R26896 GND.n3073 GND.n3072 34.6358
R26897 GND.n3072 GND.n3038 34.6358
R26898 GND.n3065 GND.n3064 34.6358
R26899 GND.n3057 GND.n3052 34.6358
R26900 GND.n3069 GND.n3068 34.6358
R26901 GND.n3068 GND.n3042 34.6358
R26902 GND.n3061 GND.n3042 34.6358
R26903 GND.n3061 GND.n3060 34.6358
R26904 GND.n3060 GND.n3050 34.6358
R26905 GND.n3091 GND.n3090 34.6358
R26906 GND.n3090 GND.n3088 34.6358
R26907 GND.n3098 GND.n3097 34.6358
R26908 GND.n3097 GND.n2893 34.6358
R26909 GND.n9822 GND.n9821 34.4123
R26910 GND.n9821 GND.n9820 34.4123
R26911 GND.n2118 GND.n2117 34.4123
R26912 GND.n2119 GND.n2118 34.4123
R26913 GND.n9450 GND.n9449 34.4123
R26914 GND.n9451 GND.n9450 34.4123
R26915 GND.n9443 GND.n9442 34.4123
R26916 GND.n9442 GND.n15 34.4123
R26917 GND.n9461 GND.n9460 34.4123
R26918 GND.n9462 GND.n9461 34.4123
R26919 GND.n9454 GND.n9453 34.4123
R26920 GND.n9453 GND.n9452 34.4123
R26921 GND.n7701 GND.n7700 34.4123
R26922 GND.n7702 GND.n7701 34.4123
R26923 GND.n7694 GND.n7693 34.4123
R26924 GND.n7693 GND.n7692 34.4123
R26925 GND.n7713 GND.n7712 34.4123
R26926 GND.n7714 GND.n7713 34.4123
R26927 GND.n7706 GND.n7705 34.4123
R26928 GND.n7705 GND.n7704 34.4123
R26929 GND.n7718 GND.n2301 34.4123
R26930 GND.n7716 GND.n2301 34.4123
R26931 GND.n7717 GND.n2300 34.4123
R26932 GND.n7715 GND.n2300 34.4123
R26933 GND.n2978 GND.n2977 33.8829
R26934 GND.n2942 GND.n2929 33.8829
R26935 GND.n2991 GND.n2990 33.8829
R26936 GND.n3013 GND.n2917 33.8829
R26937 GND.n3016 GND.n3015 33.8829
R26938 GND.n3046 GND.n3038 33.8829
R26939 GND.n3069 GND.n3041 33.8829
R26940 GND.n2899 GND.n2897 32.377
R26941 GND.n9206 GND.n9205 31.0057
R26942 GND.n6846 GND.n6803 31.0057
R26943 GND.n3057 GND.n3056 30.8711
R26944 GND.n3092 GND.n3091 30.4946
R26945 GND.n6904 GND.n6790 30.0938
R26946 GND.n7723 GND.n7722 29.8476
R26947 GND.n7708 GND.n2305 29.8476
R26948 GND.n9456 GND.n9436 29.8476
R26949 GND.n9445 GND.n9441 29.8476
R26950 GND.n6117 GND.t414 29.6067
R26951 GND.t414 GND.n2876 29.6067
R26952 GND.n6285 GND.t61 29.6067
R26953 GND.n6292 GND.t61 29.6067
R26954 GND.n3056 GND.n3050 29.3652
R26955 GND.n3079 GND.t296 29.1396
R26956 GND.n3695 GND.n3137 28.4686
R26957 GND.n3689 GND.n3137 28.4686
R26958 GND.n3689 GND.n3146 28.4686
R26959 GND.n3683 GND.n3146 28.4686
R26960 GND.n3683 GND.n3154 28.4686
R26961 GND.n3677 GND.n3154 28.4686
R26962 GND.n3677 GND.n3160 28.4686
R26963 GND.n3671 GND.n3160 28.4686
R26964 GND.n3671 GND.n3166 28.4686
R26965 GND.n3665 GND.n3166 28.4686
R26966 GND.n3665 GND.n3172 28.4686
R26967 GND.n3659 GND.n3172 28.4686
R26968 GND.n3659 GND.n3178 28.4686
R26969 GND.n3653 GND.n3178 28.4686
R26970 GND.n3653 GND.n3184 28.4686
R26971 GND.n3647 GND.n3184 28.4686
R26972 GND.n3647 GND.n3190 28.4686
R26973 GND.n3641 GND.n3190 28.4686
R26974 GND.n3641 GND.n3196 28.4686
R26975 GND.n3635 GND.n3196 28.4686
R26976 GND.n3635 GND.t151 28.4686
R26977 GND.n3629 GND.t151 28.4686
R26978 GND.n3629 GND.n3269 28.4686
R26979 GND.n3623 GND.n3269 28.4686
R26980 GND.n3623 GND.n3276 28.4686
R26981 GND.n3617 GND.n3276 28.4686
R26982 GND.n3617 GND.n3283 28.4686
R26983 GND.n3611 GND.n3283 28.4686
R26984 GND.n3611 GND.n3291 28.4686
R26985 GND.n3605 GND.n3291 28.4686
R26986 GND.n3605 GND.n3298 28.4686
R26987 GND.n3599 GND.n3298 28.4686
R26988 GND.n3599 GND.n3307 28.4686
R26989 GND.n3593 GND.n3307 28.4686
R26990 GND.n3593 GND.n3313 28.4686
R26991 GND.n3587 GND.n3313 28.4686
R26992 GND.n3587 GND.n3319 28.4686
R26993 GND.n3581 GND.n3319 28.4686
R26994 GND.n3581 GND.n3325 28.4686
R26995 GND.n3575 GND.n3325 28.4686
R26996 GND.n3575 GND.n3331 28.4686
R26997 GND.n3569 GND.n3331 28.4686
R26998 GND.n8595 GND.n1795 28.4686
R26999 GND.n8595 GND.n1789 28.4686
R27000 GND.n8601 GND.n1789 28.4686
R27001 GND.n8601 GND.n1783 28.4686
R27002 GND.n8607 GND.n1783 28.4686
R27003 GND.n8607 GND.n1777 28.4686
R27004 GND.n8613 GND.n1777 28.4686
R27005 GND.n8613 GND.n1771 28.4686
R27006 GND.n8619 GND.n1771 28.4686
R27007 GND.n8619 GND.n1765 28.4686
R27008 GND.n8625 GND.n1765 28.4686
R27009 GND.n8625 GND.n1758 28.4686
R27010 GND.n8633 GND.n1758 28.4686
R27011 GND.n8633 GND.n1752 28.4686
R27012 GND.n8639 GND.n1752 28.4686
R27013 GND.n8639 GND.n1745 28.4686
R27014 GND.n8647 GND.n1745 28.4686
R27015 GND.n8647 GND.n1739 28.4686
R27016 GND.n8653 GND.n1739 28.4686
R27017 GND.n8653 GND.n1733 28.4686
R27018 GND.t6 GND.n1733 28.4686
R27019 GND.t6 GND.n1727 28.4686
R27020 GND.n8666 GND.n1727 28.4686
R27021 GND.n8666 GND.n1004 28.4686
R27022 GND.n8783 GND.n1004 28.4686
R27023 GND.n8783 GND.n1006 28.4686
R27024 GND.n8777 GND.n1006 28.4686
R27025 GND.n8777 GND.n1015 28.4686
R27026 GND.n8771 GND.n1015 28.4686
R27027 GND.n8771 GND.n1023 28.4686
R27028 GND.n8765 GND.n1023 28.4686
R27029 GND.n8765 GND.n1029 28.4686
R27030 GND.n8759 GND.n1029 28.4686
R27031 GND.n8759 GND.n1035 28.4686
R27032 GND.n8753 GND.n1035 28.4686
R27033 GND.n8753 GND.n1041 28.4686
R27034 GND.n8747 GND.n1041 28.4686
R27035 GND.n8747 GND.n1047 28.4686
R27036 GND.n8741 GND.n1047 28.4686
R27037 GND.n8741 GND.n1053 28.4686
R27038 GND.n8735 GND.n1053 28.4686
R27039 GND.n8735 GND.n1059 28.4686
R27040 GND.n1652 GND.n1091 28.4686
R27041 GND.n1646 GND.n1091 28.4686
R27042 GND.n1646 GND.n1100 28.4686
R27043 GND.n1640 GND.n1100 28.4686
R27044 GND.n1640 GND.n1108 28.4686
R27045 GND.n1634 GND.n1108 28.4686
R27046 GND.n1634 GND.n1114 28.4686
R27047 GND.n1628 GND.n1114 28.4686
R27048 GND.n1628 GND.n1120 28.4686
R27049 GND.n1622 GND.n1120 28.4686
R27050 GND.n1622 GND.n1126 28.4686
R27051 GND.n1616 GND.n1126 28.4686
R27052 GND.n1616 GND.n1132 28.4686
R27053 GND.n1610 GND.n1132 28.4686
R27054 GND.n1610 GND.n1138 28.4686
R27055 GND.n1604 GND.n1138 28.4686
R27056 GND.n1604 GND.n1144 28.4686
R27057 GND.n1598 GND.n1144 28.4686
R27058 GND.n1598 GND.n1150 28.4686
R27059 GND.n1592 GND.n1150 28.4686
R27060 GND.n1592 GND.t310 28.4686
R27061 GND.n1586 GND.t310 28.4686
R27062 GND.n1586 GND.n1223 28.4686
R27063 GND.n1580 GND.n1223 28.4686
R27064 GND.n1580 GND.n1230 28.4686
R27065 GND.n1574 GND.n1230 28.4686
R27066 GND.n1574 GND.n1237 28.4686
R27067 GND.n1568 GND.n1237 28.4686
R27068 GND.n1568 GND.n1245 28.4686
R27069 GND.n1562 GND.n1245 28.4686
R27070 GND.n1562 GND.n1252 28.4686
R27071 GND.n1556 GND.n1252 28.4686
R27072 GND.n1556 GND.n1261 28.4686
R27073 GND.n1550 GND.n1261 28.4686
R27074 GND.n1550 GND.n1267 28.4686
R27075 GND.n1544 GND.n1267 28.4686
R27076 GND.n1544 GND.n1273 28.4686
R27077 GND.n1538 GND.n1273 28.4686
R27078 GND.n1538 GND.n1279 28.4686
R27079 GND.n1532 GND.n1279 28.4686
R27080 GND.n1532 GND.n1285 28.4686
R27081 GND.n1526 GND.n1285 28.4686
R27082 GND.n7697 GND.t349 28.3395
R27083 GND.n7696 GND.t287 28.3395
R27084 GND.n10 GND.t291 28.3395
R27085 GND.n2115 GND.t342 28.3395
R27086 GND.n9164 GND.n9135 28.2699
R27087 GND.n2977 GND.n2971 28.2358
R27088 GND.n3095 GND.n2897 28.2358
R27089 GND.n2969 GND.n2964 27.8593
R27090 GND.n2944 GND.n2940 27.8593
R27091 GND.n3025 GND.n3024 27.8593
R27092 GND.n3064 GND.n3048 27.8593
R27093 GND.n6597 GND.n6596 27.6063
R27094 GND.n6583 GND.n6582 27.6063
R27095 GND.n6569 GND.n6568 27.6063
R27096 GND.n6555 GND.n6554 27.6063
R27097 GND.n6541 GND.n6540 27.6063
R27098 GND.n2707 GND.n2706 27.6063
R27099 GND.n6456 GND.n6455 27.6063
R27100 GND.n6470 GND.n6469 27.6063
R27101 GND.n6483 GND.n6482 27.6063
R27102 GND.n6496 GND.n6495 27.6063
R27103 GND.n6509 GND.n6508 27.6063
R27104 GND.n6522 GND.n6521 27.6063
R27105 GND.n6437 GND.n6436 27.6063
R27106 GND.n8960 GND.n8959 27.6063
R27107 GND.n8946 GND.n8945 27.6063
R27108 GND.n8932 GND.n8931 27.6063
R27109 GND.n8918 GND.n8917 27.6063
R27110 GND.n8904 GND.n8903 27.6063
R27111 GND.n990 GND.n989 27.6063
R27112 GND.n8820 GND.n8819 27.6063
R27113 GND.n8834 GND.n8833 27.6063
R27114 GND.n8847 GND.n8846 27.6063
R27115 GND.n8860 GND.n8859 27.6063
R27116 GND.n8873 GND.n8872 27.6063
R27117 GND.n8886 GND.n8885 27.6063
R27118 GND.n8801 GND.n8800 27.6063
R27119 GND.n4859 GND.n4858 27.6063
R27120 GND.n4845 GND.n4844 27.6063
R27121 GND.n4831 GND.n4830 27.6063
R27122 GND.n4817 GND.n4816 27.6063
R27123 GND.n4803 GND.n4802 27.6063
R27124 GND.n4788 GND.n4787 27.6063
R27125 GND.n4182 GND.n4181 27.6063
R27126 GND.n4876 GND.n4875 27.6063
R27127 GND.n4889 GND.n4888 27.6063
R27128 GND.n4902 GND.n4901 27.6063
R27129 GND.n4915 GND.n4914 27.6063
R27130 GND.n4928 GND.n4927 27.6063
R27131 GND.n4163 GND.n4162 27.6063
R27132 GND.n3019 GND.n2915 27.1064
R27133 GND.t265 GND.n9206 25.9901
R27134 GND.n6803 GND.t215 25.9901
R27135 GND.n5056 GND.n3785 25.6005
R27136 GND.n5056 GND.n5055 25.6005
R27137 GND.n5062 GND.n5055 25.6005
R27138 GND.n5063 GND.n5062 25.6005
R27139 GND.n5064 GND.n5063 25.6005
R27140 GND.n5064 GND.n5053 25.6005
R27141 GND.n5070 GND.n5053 25.6005
R27142 GND.n5071 GND.n5070 25.6005
R27143 GND.n5072 GND.n5071 25.6005
R27144 GND.n5072 GND.n5051 25.6005
R27145 GND.n5078 GND.n5051 25.6005
R27146 GND.n5079 GND.n5078 25.6005
R27147 GND.n5080 GND.n5079 25.6005
R27148 GND.n5080 GND.n5049 25.6005
R27149 GND.n5086 GND.n5049 25.6005
R27150 GND.n5087 GND.n5086 25.6005
R27151 GND.n5134 GND.n5087 25.6005
R27152 GND.n5892 GND.n5891 25.6005
R27153 GND.n5891 GND.n5890 25.6005
R27154 GND.n5890 GND.n3729 25.6005
R27155 GND.n3748 GND.n3729 25.6005
R27156 GND.n5878 GND.n3748 25.6005
R27157 GND.n5878 GND.n5877 25.6005
R27158 GND.n5877 GND.n5876 25.6005
R27159 GND.n5876 GND.n3749 25.6005
R27160 GND.n3766 GND.n3749 25.6005
R27161 GND.n5864 GND.n3766 25.6005
R27162 GND.n5864 GND.n5863 25.6005
R27163 GND.n5863 GND.n5862 25.6005
R27164 GND.n5862 GND.n3767 25.6005
R27165 GND.n3784 GND.n3767 25.6005
R27166 GND.n5850 GND.n3784 25.6005
R27167 GND.n5850 GND.n5849 25.6005
R27168 GND.n5849 GND.n5848 25.6005
R27169 GND.n5196 GND.n3728 25.6005
R27170 GND.n5197 GND.n5196 25.6005
R27171 GND.n5198 GND.n5197 25.6005
R27172 GND.n5198 GND.n5192 25.6005
R27173 GND.n5204 GND.n5192 25.6005
R27174 GND.n5205 GND.n5204 25.6005
R27175 GND.n5206 GND.n5205 25.6005
R27176 GND.n5206 GND.n5190 25.6005
R27177 GND.n5212 GND.n5190 25.6005
R27178 GND.n5213 GND.n5212 25.6005
R27179 GND.n5214 GND.n5213 25.6005
R27180 GND.n5214 GND.n5188 25.6005
R27181 GND.n5220 GND.n5188 25.6005
R27182 GND.n5221 GND.n5220 25.6005
R27183 GND.n5222 GND.n5221 25.6005
R27184 GND.n5222 GND.n5186 25.6005
R27185 GND.n5228 GND.n5186 25.6005
R27186 GND.n5229 GND.n5228 25.6005
R27187 GND.n5230 GND.n5229 25.6005
R27188 GND.n5230 GND.n5184 25.6005
R27189 GND.n5236 GND.n5184 25.6005
R27190 GND.n5237 GND.n5236 25.6005
R27191 GND.n5238 GND.n5237 25.6005
R27192 GND.n5238 GND.n5182 25.6005
R27193 GND.n5244 GND.n5182 25.6005
R27194 GND.n5245 GND.n5244 25.6005
R27195 GND.n5246 GND.n5245 25.6005
R27196 GND.n5246 GND.n5180 25.6005
R27197 GND.n5252 GND.n5180 25.6005
R27198 GND.n5253 GND.n5252 25.6005
R27199 GND.n5254 GND.n5253 25.6005
R27200 GND.n5254 GND.n5178 25.6005
R27201 GND.n5260 GND.n5178 25.6005
R27202 GND.n5261 GND.n5260 25.6005
R27203 GND.n5262 GND.n5261 25.6005
R27204 GND.n5262 GND.n5176 25.6005
R27205 GND.n5268 GND.n5176 25.6005
R27206 GND.n5269 GND.n5268 25.6005
R27207 GND.n5270 GND.n5269 25.6005
R27208 GND.n5270 GND.n5174 25.6005
R27209 GND.n5174 GND.n5173 25.6005
R27210 GND.n5277 GND.n5173 25.6005
R27211 GND.n5281 GND.n5278 25.6005
R27212 GND.n5282 GND.n5281 25.6005
R27213 GND.n5283 GND.n5282 25.6005
R27214 GND.n5286 GND.n5283 25.6005
R27215 GND.n5287 GND.n5286 25.6005
R27216 GND.n5290 GND.n5287 25.6005
R27217 GND.n5291 GND.n5290 25.6005
R27218 GND.n5292 GND.n5291 25.6005
R27219 GND.n5295 GND.n5292 25.6005
R27220 GND.n5296 GND.n5295 25.6005
R27221 GND.n5299 GND.n5296 25.6005
R27222 GND.n5300 GND.n5299 25.6005
R27223 GND.n5301 GND.n5300 25.6005
R27224 GND.n5304 GND.n5301 25.6005
R27225 GND.n5305 GND.n5304 25.6005
R27226 GND.n5308 GND.n5305 25.6005
R27227 GND.n5309 GND.n5308 25.6005
R27228 GND.n5341 GND.n5340 25.6005
R27229 GND.n5341 GND.n5034 25.6005
R27230 GND.n5347 GND.n5034 25.6005
R27231 GND.n5348 GND.n5347 25.6005
R27232 GND.n5349 GND.n5348 25.6005
R27233 GND.n5349 GND.n5032 25.6005
R27234 GND.n5355 GND.n5032 25.6005
R27235 GND.n5356 GND.n5355 25.6005
R27236 GND.n5357 GND.n5356 25.6005
R27237 GND.n5357 GND.n5030 25.6005
R27238 GND.n5363 GND.n5030 25.6005
R27239 GND.n5364 GND.n5363 25.6005
R27240 GND.n5365 GND.n5364 25.6005
R27241 GND.n5365 GND.n5028 25.6005
R27242 GND.n5163 GND.n5036 25.6005
R27243 GND.n5331 GND.n5163 25.6005
R27244 GND.n5331 GND.n5330 25.6005
R27245 GND.n5330 GND.n5329 25.6005
R27246 GND.n5329 GND.n5165 25.6005
R27247 GND.n5324 GND.n5165 25.6005
R27248 GND.n5324 GND.n5323 25.6005
R27249 GND.n5323 GND.n5322 25.6005
R27250 GND.n5322 GND.n5168 25.6005
R27251 GND.n5317 GND.n5168 25.6005
R27252 GND.n5317 GND.n5316 25.6005
R27253 GND.n5316 GND.n5315 25.6005
R27254 GND.n5315 GND.n5171 25.6005
R27255 GND.n5310 GND.n5171 25.6005
R27256 GND.n5100 GND.n5096 25.6005
R27257 GND.n5101 GND.n5100 25.6005
R27258 GND.n5102 GND.n5101 25.6005
R27259 GND.n5102 GND.n5094 25.6005
R27260 GND.n5108 GND.n5094 25.6005
R27261 GND.n5109 GND.n5108 25.6005
R27262 GND.n5110 GND.n5109 25.6005
R27263 GND.n5110 GND.n5092 25.6005
R27264 GND.n5116 GND.n5092 25.6005
R27265 GND.n5117 GND.n5116 25.6005
R27266 GND.n5118 GND.n5117 25.6005
R27267 GND.n5118 GND.n5090 25.6005
R27268 GND.n5124 GND.n5090 25.6005
R27269 GND.n5125 GND.n5124 25.6005
R27270 GND.n5126 GND.n5125 25.6005
R27271 GND.n5126 GND.n5088 25.6005
R27272 GND.n5132 GND.n5088 25.6005
R27273 GND.n5775 GND.n3849 25.6005
R27274 GND.n5775 GND.n5774 25.6005
R27275 GND.n5774 GND.n5773 25.6005
R27276 GND.n5773 GND.n3850 25.6005
R27277 GND.n3867 GND.n3850 25.6005
R27278 GND.n5761 GND.n3867 25.6005
R27279 GND.n5761 GND.n5760 25.6005
R27280 GND.n5760 GND.n5759 25.6005
R27281 GND.n5759 GND.n3868 25.6005
R27282 GND.n3885 GND.n3868 25.6005
R27283 GND.n5747 GND.n3885 25.6005
R27284 GND.n5747 GND.n5746 25.6005
R27285 GND.n5746 GND.n5745 25.6005
R27286 GND.n5745 GND.n3886 25.6005
R27287 GND.n3903 GND.n3886 25.6005
R27288 GND.n5733 GND.n3903 25.6005
R27289 GND.n5733 GND.n5732 25.6005
R27290 GND.n5731 GND.n3904 25.6005
R27291 GND.n5726 GND.n3904 25.6005
R27292 GND.n5726 GND.n5725 25.6005
R27293 GND.n5725 GND.n5724 25.6005
R27294 GND.n5724 GND.n5721 25.6005
R27295 GND.n5721 GND.n5720 25.6005
R27296 GND.n5720 GND.n5717 25.6005
R27297 GND.n5717 GND.n5716 25.6005
R27298 GND.n5716 GND.n5713 25.6005
R27299 GND.n5713 GND.n5712 25.6005
R27300 GND.n5712 GND.n5709 25.6005
R27301 GND.n5709 GND.n5708 25.6005
R27302 GND.n5708 GND.n5705 25.6005
R27303 GND.n5705 GND.n5704 25.6005
R27304 GND.n5704 GND.n5701 25.6005
R27305 GND.n5701 GND.n5700 25.6005
R27306 GND.n5700 GND.n5697 25.6005
R27307 GND.n5697 GND.n5696 25.6005
R27308 GND.n5021 GND.n5018 25.6005
R27309 GND.n5022 GND.n5021 25.6005
R27310 GND.n5431 GND.n5428 25.6005
R27311 GND.n5428 GND.n5427 25.6005
R27312 GND.n5427 GND.n5424 25.6005
R27313 GND.n5424 GND.n5423 25.6005
R27314 GND.n5423 GND.n5420 25.6005
R27315 GND.n5420 GND.n5419 25.6005
R27316 GND.n5419 GND.n5416 25.6005
R27317 GND.n5416 GND.n5415 25.6005
R27318 GND.n5415 GND.n5412 25.6005
R27319 GND.n5412 GND.n5411 25.6005
R27320 GND.n5411 GND.n5408 25.6005
R27321 GND.n5408 GND.n5407 25.6005
R27322 GND.n5407 GND.n5404 25.6005
R27323 GND.n5404 GND.n5403 25.6005
R27324 GND.n5371 GND.n5370 25.6005
R27325 GND.n5374 GND.n5371 25.6005
R27326 GND.n5375 GND.n5374 25.6005
R27327 GND.n5376 GND.n5375 25.6005
R27328 GND.n5379 GND.n5376 25.6005
R27329 GND.n5380 GND.n5379 25.6005
R27330 GND.n5383 GND.n5380 25.6005
R27331 GND.n5384 GND.n5383 25.6005
R27332 GND.n5385 GND.n5384 25.6005
R27333 GND.n5388 GND.n5385 25.6005
R27334 GND.n5389 GND.n5388 25.6005
R27335 GND.n5392 GND.n5389 25.6005
R27336 GND.n5393 GND.n5392 25.6005
R27337 GND.n5394 GND.n5393 25.6005
R27338 GND.n5397 GND.n5394 25.6005
R27339 GND.n5398 GND.n5397 25.6005
R27340 GND.n5399 GND.n5398 25.6005
R27341 GND.n6176 GND.n6139 25.6005
R27342 GND.n6171 GND.n6139 25.6005
R27343 GND.n6171 GND.n6170 25.6005
R27344 GND.n6170 GND.n6169 25.6005
R27345 GND.n6169 GND.n6141 25.6005
R27346 GND.n6164 GND.n6141 25.6005
R27347 GND.n6164 GND.n6163 25.6005
R27348 GND.n6163 GND.n6162 25.6005
R27349 GND.n6162 GND.n6144 25.6005
R27350 GND.n6157 GND.n6144 25.6005
R27351 GND.n6157 GND.n6156 25.6005
R27352 GND.n6156 GND.n6155 25.6005
R27353 GND.n6155 GND.n6147 25.6005
R27354 GND.n6150 GND.n6147 25.6005
R27355 GND.n6150 GND.n2793 25.6005
R27356 GND.n6091 GND.n2890 25.6005
R27357 GND.n6101 GND.n2890 25.6005
R27358 GND.n6102 GND.n6101 25.6005
R27359 GND.n6103 GND.n6102 25.6005
R27360 GND.n6103 GND.n2882 25.6005
R27361 GND.n6113 GND.n2882 25.6005
R27362 GND.n6114 GND.n6113 25.6005
R27363 GND.n6115 GND.n6114 25.6005
R27364 GND.n6115 GND.n2874 25.6005
R27365 GND.n6125 GND.n2874 25.6005
R27366 GND.n6126 GND.n6125 25.6005
R27367 GND.n6127 GND.n6126 25.6005
R27368 GND.n6127 GND.n2866 25.6005
R27369 GND.n6137 GND.n2866 25.6005
R27370 GND.n6138 GND.n6137 25.6005
R27371 GND.n6178 GND.n6138 25.6005
R27372 GND.n6178 GND.n6177 25.6005
R27373 GND.n6090 GND.n6089 25.6005
R27374 GND.n6089 GND.n5987 25.6005
R27375 GND.n6084 GND.n5987 25.6005
R27376 GND.n6084 GND.n6083 25.6005
R27377 GND.n6083 GND.n5989 25.6005
R27378 GND.n6078 GND.n5989 25.6005
R27379 GND.n6078 GND.n6077 25.6005
R27380 GND.n6077 GND.n6076 25.6005
R27381 GND.n6076 GND.n5991 25.6005
R27382 GND.n6070 GND.n5991 25.6005
R27383 GND.n6070 GND.n6069 25.6005
R27384 GND.n6069 GND.n6068 25.6005
R27385 GND.n6068 GND.n5993 25.6005
R27386 GND.n6062 GND.n5993 25.6005
R27387 GND.n6062 GND.n6061 25.6005
R27388 GND.n6061 GND.n6060 25.6005
R27389 GND.n6060 GND.n5995 25.6005
R27390 GND.n6054 GND.n5995 25.6005
R27391 GND.n6054 GND.n6053 25.6005
R27392 GND.n6053 GND.n6052 25.6005
R27393 GND.n6052 GND.n5997 25.6005
R27394 GND.n6046 GND.n5997 25.6005
R27395 GND.n6046 GND.n6045 25.6005
R27396 GND.n6045 GND.n6044 25.6005
R27397 GND.n6044 GND.n5999 25.6005
R27398 GND.n6038 GND.n5999 25.6005
R27399 GND.n6038 GND.n6037 25.6005
R27400 GND.n6037 GND.n6036 25.6005
R27401 GND.n6036 GND.n6001 25.6005
R27402 GND.n6030 GND.n6001 25.6005
R27403 GND.n6030 GND.n6029 25.6005
R27404 GND.n6029 GND.n6028 25.6005
R27405 GND.n6028 GND.n6003 25.6005
R27406 GND.n6022 GND.n6003 25.6005
R27407 GND.n6022 GND.n6021 25.6005
R27408 GND.n6021 GND.n6020 25.6005
R27409 GND.n6020 GND.n6005 25.6005
R27410 GND.n6014 GND.n6005 25.6005
R27411 GND.n6014 GND.n6013 25.6005
R27412 GND.n6013 GND.n6012 25.6005
R27413 GND.n6012 GND.n6007 25.6005
R27414 GND.n6007 GND.n3115 25.6005
R27415 GND.n6096 GND.n6095 25.6005
R27416 GND.n6097 GND.n6096 25.6005
R27417 GND.n6097 GND.n2886 25.6005
R27418 GND.n6107 GND.n2886 25.6005
R27419 GND.n6108 GND.n6107 25.6005
R27420 GND.n6109 GND.n6108 25.6005
R27421 GND.n6109 GND.n2878 25.6005
R27422 GND.n6119 GND.n2878 25.6005
R27423 GND.n6120 GND.n6119 25.6005
R27424 GND.n6121 GND.n6120 25.6005
R27425 GND.n6121 GND.n2870 25.6005
R27426 GND.n6131 GND.n2870 25.6005
R27427 GND.n6132 GND.n6131 25.6005
R27428 GND.n6133 GND.n6132 25.6005
R27429 GND.n6133 GND.n2860 25.6005
R27430 GND.n6182 GND.n2860 25.6005
R27431 GND.n6183 GND.n6182 25.6005
R27432 GND.n6421 GND.n2718 25.6005
R27433 GND.n2721 GND.n2718 25.6005
R27434 GND.n6414 GND.n2721 25.6005
R27435 GND.n6414 GND.n6413 25.6005
R27436 GND.n6413 GND.n6412 25.6005
R27437 GND.n6412 GND.n2723 25.6005
R27438 GND.n6407 GND.n2723 25.6005
R27439 GND.n6407 GND.n6406 25.6005
R27440 GND.n6406 GND.n6405 25.6005
R27441 GND.n6405 GND.n2726 25.6005
R27442 GND.n6400 GND.n2726 25.6005
R27443 GND.n6400 GND.n6399 25.6005
R27444 GND.n6399 GND.n6398 25.6005
R27445 GND.n6398 GND.n2729 25.6005
R27446 GND.n6393 GND.n2729 25.6005
R27447 GND.n6393 GND.n6392 25.6005
R27448 GND.n6392 GND.n6391 25.6005
R27449 GND.n6269 GND.n2765 25.6005
R27450 GND.n6270 GND.n6269 25.6005
R27451 GND.n6271 GND.n6270 25.6005
R27452 GND.n6271 GND.n2757 25.6005
R27453 GND.n6281 GND.n2757 25.6005
R27454 GND.n6282 GND.n6281 25.6005
R27455 GND.n6283 GND.n6282 25.6005
R27456 GND.n6283 GND.n2750 25.6005
R27457 GND.n6294 GND.n2750 25.6005
R27458 GND.n6295 GND.n6294 25.6005
R27459 GND.n6296 GND.n6295 25.6005
R27460 GND.n6296 GND.n2742 25.6005
R27461 GND.n6306 GND.n2742 25.6005
R27462 GND.n6307 GND.n6306 25.6005
R27463 GND.n6309 GND.n6307 25.6005
R27464 GND.n6309 GND.n6308 25.6005
R27465 GND.n6308 GND.n2732 25.6005
R27466 GND.n2846 GND.n2843 25.6005
R27467 GND.n2843 GND.n2842 25.6005
R27468 GND.n2842 GND.n2839 25.6005
R27469 GND.n2839 GND.n2838 25.6005
R27470 GND.n2838 GND.n2835 25.6005
R27471 GND.n2835 GND.n2834 25.6005
R27472 GND.n2834 GND.n2831 25.6005
R27473 GND.n2831 GND.n2830 25.6005
R27474 GND.n2830 GND.n2827 25.6005
R27475 GND.n2827 GND.n2826 25.6005
R27476 GND.n2826 GND.n2823 25.6005
R27477 GND.n2823 GND.n2822 25.6005
R27478 GND.n2822 GND.n2819 25.6005
R27479 GND.n2819 GND.n2818 25.6005
R27480 GND.n2818 GND.n2815 25.6005
R27481 GND.n2815 GND.n2814 25.6005
R27482 GND.n6212 GND.n6211 25.6005
R27483 GND.n6211 GND.n6210 25.6005
R27484 GND.n6210 GND.n2848 25.6005
R27485 GND.n6205 GND.n2848 25.6005
R27486 GND.n6205 GND.n6204 25.6005
R27487 GND.n6204 GND.n6203 25.6005
R27488 GND.n6203 GND.n2851 25.6005
R27489 GND.n6198 GND.n2851 25.6005
R27490 GND.n6198 GND.n6197 25.6005
R27491 GND.n6197 GND.n6196 25.6005
R27492 GND.n6196 GND.n2854 25.6005
R27493 GND.n6191 GND.n2854 25.6005
R27494 GND.n6191 GND.n6190 25.6005
R27495 GND.n6190 GND.n6189 25.6005
R27496 GND.n6189 GND.n2857 25.6005
R27497 GND.n6184 GND.n2857 25.6005
R27498 GND.n6263 GND.n2769 25.6005
R27499 GND.n6258 GND.n2769 25.6005
R27500 GND.n6258 GND.n6257 25.6005
R27501 GND.n6257 GND.n6256 25.6005
R27502 GND.n6256 GND.n6253 25.6005
R27503 GND.n6253 GND.n6252 25.6005
R27504 GND.n6252 GND.n6249 25.6005
R27505 GND.n6249 GND.n6248 25.6005
R27506 GND.n6248 GND.n6245 25.6005
R27507 GND.n6245 GND.n6244 25.6005
R27508 GND.n6244 GND.n6241 25.6005
R27509 GND.n6241 GND.n6240 25.6005
R27510 GND.n6240 GND.n6237 25.6005
R27511 GND.n6237 GND.n6236 25.6005
R27512 GND.n6236 GND.n6233 25.6005
R27513 GND.n6265 GND.n6264 25.6005
R27514 GND.n6265 GND.n2761 25.6005
R27515 GND.n6275 GND.n2761 25.6005
R27516 GND.n6276 GND.n6275 25.6005
R27517 GND.n6277 GND.n6276 25.6005
R27518 GND.n6277 GND.n2753 25.6005
R27519 GND.n6288 GND.n2753 25.6005
R27520 GND.n6289 GND.n6288 25.6005
R27521 GND.n6290 GND.n6289 25.6005
R27522 GND.n6290 GND.n2746 25.6005
R27523 GND.n6300 GND.n2746 25.6005
R27524 GND.n6301 GND.n6300 25.6005
R27525 GND.n6302 GND.n6301 25.6005
R27526 GND.n6302 GND.n2738 25.6005
R27527 GND.n6313 GND.n2738 25.6005
R27528 GND.n6314 GND.n6313 25.6005
R27529 GND.n6386 GND.n6314 25.6005
R27530 GND.n6385 GND.n6384 25.6005
R27531 GND.n6384 GND.n6315 25.6005
R27532 GND.n6316 GND.n6315 25.6005
R27533 GND.n6377 GND.n6316 25.6005
R27534 GND.n6377 GND.n6376 25.6005
R27535 GND.n6376 GND.n6375 25.6005
R27536 GND.n6375 GND.n6318 25.6005
R27537 GND.n6370 GND.n6318 25.6005
R27538 GND.n6370 GND.n6369 25.6005
R27539 GND.n6369 GND.n6368 25.6005
R27540 GND.n6368 GND.n6321 25.6005
R27541 GND.n6363 GND.n6321 25.6005
R27542 GND.n6363 GND.n6362 25.6005
R27543 GND.n6362 GND.n6361 25.6005
R27544 GND.n6361 GND.n6324 25.6005
R27545 GND.n6348 GND.n6331 25.6005
R27546 GND.n6334 GND.n6331 25.6005
R27547 GND.n5608 GND.n5560 25.6005
R27548 GND.n5609 GND.n5608 25.6005
R27549 GND.n5612 GND.n5609 25.6005
R27550 GND.n5613 GND.n5612 25.6005
R27551 GND.n5614 GND.n5613 25.6005
R27552 GND.n5615 GND.n5555 25.6005
R27553 GND.n5619 GND.n5618 25.6005
R27554 GND.n7637 GND.n7636 25.6005
R27555 GND.n7636 GND.n7635 25.6005
R27556 GND.n7635 GND.n2343 25.6005
R27557 GND.n2371 GND.n2343 25.6005
R27558 GND.n2374 GND.n2371 25.6005
R27559 GND.n2375 GND.n2374 25.6005
R27560 GND.n7616 GND.n2375 25.6005
R27561 GND.n7616 GND.n7615 25.6005
R27562 GND.n7615 GND.n7614 25.6005
R27563 GND.n7614 GND.n2376 25.6005
R27564 GND.n2393 GND.n2376 25.6005
R27565 GND.n7602 GND.n2393 25.6005
R27566 GND.n7602 GND.n7601 25.6005
R27567 GND.n7601 GND.n7600 25.6005
R27568 GND.n7600 GND.n2394 25.6005
R27569 GND.n5532 GND.n2342 25.6005
R27570 GND.n5545 GND.n5530 25.6005
R27571 GND.n5544 GND.n5543 25.6005
R27572 GND.n5543 GND.n5540 25.6005
R27573 GND.n5540 GND.n5539 25.6005
R27574 GND.n5539 GND.n5536 25.6005
R27575 GND.n5536 GND.n5459 25.6005
R27576 GND.n7609 GND.n7608 25.6005
R27577 GND.n7608 GND.n7607 25.6005
R27578 GND.n7607 GND.n2385 25.6005
R27579 GND.n2402 GND.n2385 25.6005
R27580 GND.n7595 GND.n2402 25.6005
R27581 GND.n7595 GND.n7594 25.6005
R27582 GND.n7594 GND.n7593 25.6005
R27583 GND.n7593 GND.n2403 25.6005
R27584 GND.n7587 GND.n2403 25.6005
R27585 GND.n7586 GND.n7585 25.6005
R27586 GND.n7585 GND.n2409 25.6005
R27587 GND.n5565 GND.n2409 25.6005
R27588 GND.n5566 GND.n5565 25.6005
R27589 GND.n5569 GND.n5566 25.6005
R27590 GND.n5570 GND.n5569 25.6005
R27591 GND.n5573 GND.n5570 25.6005
R27592 GND.n5574 GND.n5573 25.6005
R27593 GND.n5577 GND.n5574 25.6005
R27594 GND.n5578 GND.n5577 25.6005
R27595 GND.n5581 GND.n5578 25.6005
R27596 GND.n5582 GND.n5581 25.6005
R27597 GND.n5585 GND.n5582 25.6005
R27598 GND.n5586 GND.n5585 25.6005
R27599 GND.n5589 GND.n5586 25.6005
R27600 GND.n5591 GND.n5589 25.6005
R27601 GND.n5603 GND.n5563 25.6005
R27602 GND.n5603 GND.n5602 25.6005
R27603 GND.n5602 GND.n5601 25.6005
R27604 GND.n5601 GND.n5598 25.6005
R27605 GND.n5598 GND.n5597 25.6005
R27606 GND.n5597 GND.n5596 25.6005
R27607 GND.n5596 GND.n5594 25.6005
R27608 GND.n5594 GND.n5593 25.6005
R27609 GND.n5593 GND.n5592 25.6005
R27610 GND.n2330 GND.n2328 25.6005
R27611 GND.n5500 GND.n2330 25.6005
R27612 GND.n5501 GND.n5500 25.6005
R27613 GND.n5502 GND.n5501 25.6005
R27614 GND.n5503 GND.n5502 25.6005
R27615 GND.n5506 GND.n5503 25.6005
R27616 GND.n5507 GND.n5506 25.6005
R27617 GND.n5511 GND.n5507 25.6005
R27618 GND.n5511 GND.n5510 25.6005
R27619 GND.n7681 GND.n7680 25.6005
R27620 GND.n7680 GND.n7679 25.6005
R27621 GND.n7679 GND.n7676 25.6005
R27622 GND.n7676 GND.n7675 25.6005
R27623 GND.n7675 GND.n7672 25.6005
R27624 GND.n7672 GND.n7671 25.6005
R27625 GND.n7671 GND.n7668 25.6005
R27626 GND.n7668 GND.n7667 25.6005
R27627 GND.n7667 GND.n7664 25.6005
R27628 GND.n7664 GND.n7663 25.6005
R27629 GND.n7663 GND.n7660 25.6005
R27630 GND.n7660 GND.n7659 25.6005
R27631 GND.n7659 GND.n7656 25.6005
R27632 GND.n7656 GND.n7655 25.6005
R27633 GND.n7655 GND.n7652 25.6005
R27634 GND.n7652 GND.n7651 25.6005
R27635 GND.n7645 GND.n2327 25.6005
R27636 GND.n7645 GND.n7644 25.6005
R27637 GND.n7644 GND.n7643 25.6005
R27638 GND.n7643 GND.n2333 25.6005
R27639 GND.n2352 GND.n2333 25.6005
R27640 GND.n2353 GND.n2352 25.6005
R27641 GND.n7630 GND.n2353 25.6005
R27642 GND.n7630 GND.n7629 25.6005
R27643 GND.n7629 GND.n7628 25.6005
R27644 GND.n5495 GND.n2362 25.6005
R27645 GND.n5496 GND.n5495 25.6005
R27646 GND.n7623 GND.n7622 25.6005
R27647 GND.n7622 GND.n7621 25.6005
R27648 GND.n7621 GND.n2363 25.6005
R27649 GND.n5473 GND.n2363 25.6005
R27650 GND.n5474 GND.n5473 25.6005
R27651 GND.n5475 GND.n5470 25.6005
R27652 GND.n5470 GND.n5469 25.6005
R27653 GND.n5640 GND.n5465 25.6005
R27654 GND.n5641 GND.n5640 25.6005
R27655 GND.n5648 GND.n5462 25.6005
R27656 GND.n5648 GND.n5647 25.6005
R27657 GND.n5647 GND.n5646 25.6005
R27658 GND.n5646 GND.n5463 25.6005
R27659 GND.n5642 GND.n5463 25.6005
R27660 GND.n5520 GND.n5519 25.6005
R27661 GND.n5519 GND.n5518 25.6005
R27662 GND.n1188 GND.n1186 25.6005
R27663 GND.n1189 GND.n1188 25.6005
R27664 GND.n1191 GND.n1189 25.6005
R27665 GND.n1192 GND.n1191 25.6005
R27666 GND.n1194 GND.n1192 25.6005
R27667 GND.n1195 GND.n1194 25.6005
R27668 GND.n1197 GND.n1195 25.6005
R27669 GND.n1198 GND.n1197 25.6005
R27670 GND.n1200 GND.n1198 25.6005
R27671 GND.n1201 GND.n1200 25.6005
R27672 GND.n1203 GND.n1201 25.6005
R27673 GND.n1204 GND.n1203 25.6005
R27674 GND.n1206 GND.n1204 25.6005
R27675 GND.n1207 GND.n1206 25.6005
R27676 GND.n1209 GND.n1207 25.6005
R27677 GND.n1210 GND.n1209 25.6005
R27678 GND.n1212 GND.n1210 25.6005
R27679 GND.n1152 GND.n1095 25.6005
R27680 GND.n1155 GND.n1152 25.6005
R27681 GND.n1156 GND.n1155 25.6005
R27682 GND.n1159 GND.n1156 25.6005
R27683 GND.n1160 GND.n1159 25.6005
R27684 GND.n1163 GND.n1160 25.6005
R27685 GND.n1164 GND.n1163 25.6005
R27686 GND.n1167 GND.n1164 25.6005
R27687 GND.n1168 GND.n1167 25.6005
R27688 GND.n1171 GND.n1168 25.6005
R27689 GND.n1172 GND.n1171 25.6005
R27690 GND.n1175 GND.n1172 25.6005
R27691 GND.n1176 GND.n1175 25.6005
R27692 GND.n1179 GND.n1176 25.6005
R27693 GND.n1180 GND.n1179 25.6005
R27694 GND.n1183 GND.n1180 25.6005
R27695 GND.n1185 GND.n1183 25.6005
R27696 GND.n1650 GND.n1649 25.6005
R27697 GND.n1649 GND.n1648 25.6005
R27698 GND.n1648 GND.n1096 25.6005
R27699 GND.n1638 GND.n1096 25.6005
R27700 GND.n1638 GND.n1637 25.6005
R27701 GND.n1637 GND.n1636 25.6005
R27702 GND.n1636 GND.n1110 25.6005
R27703 GND.n1626 GND.n1110 25.6005
R27704 GND.n1626 GND.n1625 25.6005
R27705 GND.n1625 GND.n1624 25.6005
R27706 GND.n1624 GND.n1122 25.6005
R27707 GND.n1614 GND.n1122 25.6005
R27708 GND.n1614 GND.n1613 25.6005
R27709 GND.n1613 GND.n1612 25.6005
R27710 GND.n1612 GND.n1134 25.6005
R27711 GND.n1602 GND.n1134 25.6005
R27712 GND.n1602 GND.n1601 25.6005
R27713 GND.n1601 GND.n1600 25.6005
R27714 GND.n1600 GND.n1146 25.6005
R27715 GND.n1590 GND.n1146 25.6005
R27716 GND.n1590 GND.n1589 25.6005
R27717 GND.n1589 GND.n1588 25.6005
R27718 GND.n1588 GND.n1219 25.6005
R27719 GND.n1578 GND.n1219 25.6005
R27720 GND.n1578 GND.n1577 25.6005
R27721 GND.n1577 GND.n1576 25.6005
R27722 GND.n1576 GND.n1233 25.6005
R27723 GND.n1566 GND.n1233 25.6005
R27724 GND.n1566 GND.n1565 25.6005
R27725 GND.n1565 GND.n1564 25.6005
R27726 GND.n1564 GND.n1248 25.6005
R27727 GND.n1554 GND.n1248 25.6005
R27728 GND.n1554 GND.n1553 25.6005
R27729 GND.n1553 GND.n1552 25.6005
R27730 GND.n1552 GND.n1263 25.6005
R27731 GND.n1542 GND.n1263 25.6005
R27732 GND.n1542 GND.n1541 25.6005
R27733 GND.n1541 GND.n1540 25.6005
R27734 GND.n1540 GND.n1275 25.6005
R27735 GND.n1530 GND.n1275 25.6005
R27736 GND.n1530 GND.n1529 25.6005
R27737 GND.n1529 GND.n1528 25.6005
R27738 GND.n1317 GND.n1287 25.6005
R27739 GND.n1317 GND.n1316 25.6005
R27740 GND.n1323 GND.n1316 25.6005
R27741 GND.n1324 GND.n1323 25.6005
R27742 GND.n1325 GND.n1324 25.6005
R27743 GND.n1325 GND.n1314 25.6005
R27744 GND.n1331 GND.n1314 25.6005
R27745 GND.n1332 GND.n1331 25.6005
R27746 GND.n1333 GND.n1332 25.6005
R27747 GND.n1333 GND.n1312 25.6005
R27748 GND.n1339 GND.n1312 25.6005
R27749 GND.n1340 GND.n1339 25.6005
R27750 GND.n1341 GND.n1340 25.6005
R27751 GND.n1341 GND.n1310 25.6005
R27752 GND.n1310 GND.n1309 25.6005
R27753 GND.n1348 GND.n1309 25.6005
R27754 GND.n1349 GND.n1348 25.6005
R27755 GND.n1448 GND.n1447 25.6005
R27756 GND.n1447 GND.n1445 25.6005
R27757 GND.n1468 GND.n1466 25.6005
R27758 GND.n1469 GND.n1468 25.6005
R27759 GND.n1471 GND.n1469 25.6005
R27760 GND.n1472 GND.n1471 25.6005
R27761 GND.n1474 GND.n1472 25.6005
R27762 GND.n1475 GND.n1474 25.6005
R27763 GND.n1477 GND.n1475 25.6005
R27764 GND.n1478 GND.n1477 25.6005
R27765 GND.n1480 GND.n1478 25.6005
R27766 GND.n1481 GND.n1480 25.6005
R27767 GND.n1483 GND.n1481 25.6005
R27768 GND.n1484 GND.n1483 25.6005
R27769 GND.n1486 GND.n1484 25.6005
R27770 GND.n1487 GND.n1486 25.6005
R27771 GND.n1523 GND.n1522 25.6005
R27772 GND.n1522 GND.n1354 25.6005
R27773 GND.n1516 GND.n1354 25.6005
R27774 GND.n1516 GND.n1515 25.6005
R27775 GND.n1515 GND.n1514 25.6005
R27776 GND.n1514 GND.n1356 25.6005
R27777 GND.n1508 GND.n1356 25.6005
R27778 GND.n1508 GND.n1507 25.6005
R27779 GND.n1507 GND.n1506 25.6005
R27780 GND.n1506 GND.n1358 25.6005
R27781 GND.n1500 GND.n1358 25.6005
R27782 GND.n1500 GND.n1499 25.6005
R27783 GND.n1499 GND.n1498 25.6005
R27784 GND.n1498 GND.n1360 25.6005
R27785 GND.n1492 GND.n1360 25.6005
R27786 GND.n1492 GND.n1491 25.6005
R27787 GND.n1491 GND.n1490 25.6005
R27788 GND.n1256 GND.n1255 25.6005
R27789 GND.n1560 GND.n1256 25.6005
R27790 GND.n1560 GND.n1559 25.6005
R27791 GND.n1559 GND.n1558 25.6005
R27792 GND.n1558 GND.n1257 25.6005
R27793 GND.n1548 GND.n1257 25.6005
R27794 GND.n1548 GND.n1547 25.6005
R27795 GND.n1547 GND.n1546 25.6005
R27796 GND.n1546 GND.n1269 25.6005
R27797 GND.n1536 GND.n1269 25.6005
R27798 GND.n1536 GND.n1535 25.6005
R27799 GND.n1535 GND.n1534 25.6005
R27800 GND.n1534 GND.n1281 25.6005
R27801 GND.n1524 GND.n1281 25.6005
R27802 GND.n1291 GND.n1243 25.6005
R27803 GND.n1292 GND.n1291 25.6005
R27804 GND.n1294 GND.n1292 25.6005
R27805 GND.n1295 GND.n1294 25.6005
R27806 GND.n1297 GND.n1295 25.6005
R27807 GND.n1298 GND.n1297 25.6005
R27808 GND.n1300 GND.n1298 25.6005
R27809 GND.n1301 GND.n1300 25.6005
R27810 GND.n1303 GND.n1301 25.6005
R27811 GND.n1304 GND.n1303 25.6005
R27812 GND.n1306 GND.n1304 25.6005
R27813 GND.n1307 GND.n1306 25.6005
R27814 GND.n1308 GND.n1307 25.6005
R27815 GND.n1350 GND.n1308 25.6005
R27816 GND.n1369 GND.n1103 25.6005
R27817 GND.n1644 GND.n1103 25.6005
R27818 GND.n1644 GND.n1643 25.6005
R27819 GND.n1643 GND.n1642 25.6005
R27820 GND.n1642 GND.n1104 25.6005
R27821 GND.n1632 GND.n1104 25.6005
R27822 GND.n1632 GND.n1631 25.6005
R27823 GND.n1631 GND.n1630 25.6005
R27824 GND.n1630 GND.n1116 25.6005
R27825 GND.n1620 GND.n1116 25.6005
R27826 GND.n1620 GND.n1619 25.6005
R27827 GND.n1619 GND.n1618 25.6005
R27828 GND.n1618 GND.n1128 25.6005
R27829 GND.n1608 GND.n1128 25.6005
R27830 GND.n1608 GND.n1607 25.6005
R27831 GND.n1607 GND.n1606 25.6005
R27832 GND.n1606 GND.n1140 25.6005
R27833 GND.n1372 GND.n1371 25.6005
R27834 GND.n1375 GND.n1372 25.6005
R27835 GND.n1376 GND.n1375 25.6005
R27836 GND.n1379 GND.n1376 25.6005
R27837 GND.n1380 GND.n1379 25.6005
R27838 GND.n1383 GND.n1380 25.6005
R27839 GND.n1384 GND.n1383 25.6005
R27840 GND.n1387 GND.n1384 25.6005
R27841 GND.n1388 GND.n1387 25.6005
R27842 GND.n1391 GND.n1388 25.6005
R27843 GND.n1392 GND.n1391 25.6005
R27844 GND.n1395 GND.n1392 25.6005
R27845 GND.n1396 GND.n1395 25.6005
R27846 GND.n1399 GND.n1396 25.6005
R27847 GND.n1400 GND.n1399 25.6005
R27848 GND.n1403 GND.n1400 25.6005
R27849 GND.n1405 GND.n1403 25.6005
R27850 GND.n1408 GND.n1406 25.6005
R27851 GND.n1409 GND.n1408 25.6005
R27852 GND.n1411 GND.n1409 25.6005
R27853 GND.n1412 GND.n1411 25.6005
R27854 GND.n1414 GND.n1412 25.6005
R27855 GND.n1415 GND.n1414 25.6005
R27856 GND.n1417 GND.n1415 25.6005
R27857 GND.n1418 GND.n1417 25.6005
R27858 GND.n1420 GND.n1418 25.6005
R27859 GND.n1421 GND.n1420 25.6005
R27860 GND.n1423 GND.n1421 25.6005
R27861 GND.n1424 GND.n1423 25.6005
R27862 GND.n1426 GND.n1424 25.6005
R27863 GND.n1427 GND.n1426 25.6005
R27864 GND.n1429 GND.n1427 25.6005
R27865 GND.n1430 GND.n1429 25.6005
R27866 GND.n1432 GND.n1430 25.6005
R27867 GND.n1433 GND.n1432 25.6005
R27868 GND.n9707 GND.n9706 25.6005
R27869 GND.n9706 GND.n9705 25.6005
R27870 GND.n9705 GND.n105 25.6005
R27871 GND.n9612 GND.n105 25.6005
R27872 GND.n9613 GND.n9612 25.6005
R27873 GND.n9614 GND.n9610 25.6005
R27874 GND.n9692 GND.n9691 25.6005
R27875 GND.n9558 GND.n9557 25.6005
R27876 GND.n9558 GND.n164 25.6005
R27877 GND.n9581 GND.n164 25.6005
R27878 GND.n9582 GND.n9581 25.6005
R27879 GND.n9586 GND.n9582 25.6005
R27880 GND.n9586 GND.n9585 25.6005
R27881 GND.n9585 GND.n9584 25.6005
R27882 GND.n9584 GND.n87 25.6005
R27883 GND.n9739 GND.n87 25.6005
R27884 GND.n9739 GND.n9738 25.6005
R27885 GND.n9738 GND.n9737 25.6005
R27886 GND.n9737 GND.n88 25.6005
R27887 GND.n125 GND.n88 25.6005
R27888 GND.n126 GND.n125 25.6005
R27889 GND.n9693 GND.n126 25.6005
R27890 GND.n9556 GND.n173 25.6005
R27891 GND.n9548 GND.n9547 25.6005
R27892 GND.n9562 GND.n169 25.6005
R27893 GND.n9563 GND.n9562 25.6005
R27894 GND.n9577 GND.n9563 25.6005
R27895 GND.n9577 GND.n9576 25.6005
R27896 GND.n9576 GND.n9575 25.6005
R27897 GND.n114 GND.n111 25.6005
R27898 GND.n115 GND.n114 25.6005
R27899 GND.n9700 GND.n115 25.6005
R27900 GND.n9700 GND.n9699 25.6005
R27901 GND.n9699 GND.n9698 25.6005
R27902 GND.n9698 GND.n116 25.6005
R27903 GND.n9685 GND.n116 25.6005
R27904 GND.n9685 GND.n9684 25.6005
R27905 GND.n9684 GND.n9683 25.6005
R27906 GND.n9677 GND.n9619 25.6005
R27907 GND.n9677 GND.n9676 25.6005
R27908 GND.n9676 GND.n9675 25.6005
R27909 GND.n9675 GND.n9673 25.6005
R27910 GND.n9673 GND.n9670 25.6005
R27911 GND.n9670 GND.n9669 25.6005
R27912 GND.n9669 GND.n9666 25.6005
R27913 GND.n9666 GND.n9665 25.6005
R27914 GND.n9665 GND.n9662 25.6005
R27915 GND.n9662 GND.n9661 25.6005
R27916 GND.n9661 GND.n9658 25.6005
R27917 GND.n9658 GND.n9657 25.6005
R27918 GND.n9657 GND.n9654 25.6005
R27919 GND.n9654 GND.n9653 25.6005
R27920 GND.n9653 GND.n9650 25.6005
R27921 GND.n9650 GND.n9649 25.6005
R27922 GND.n9632 GND.n9630 25.6005
R27923 GND.n9636 GND.n9630 25.6005
R27924 GND.n9637 GND.n9636 25.6005
R27925 GND.n9640 GND.n9637 25.6005
R27926 GND.n9641 GND.n9640 25.6005
R27927 GND.n9643 GND.n9641 25.6005
R27928 GND.n9644 GND.n9643 25.6005
R27929 GND.n9646 GND.n9644 25.6005
R27930 GND.n9647 GND.n9646 25.6005
R27931 GND.n9473 GND.n184 25.6005
R27932 GND.n9514 GND.n184 25.6005
R27933 GND.n9515 GND.n9514 25.6005
R27934 GND.n9517 GND.n9515 25.6005
R27935 GND.n9518 GND.n9517 25.6005
R27936 GND.n9530 GND.n9518 25.6005
R27937 GND.n9530 GND.n9529 25.6005
R27938 GND.n9529 GND.n9528 25.6005
R27939 GND.n9528 GND.n9520 25.6005
R27940 GND.n9507 GND.n187 25.6005
R27941 GND.n9502 GND.n187 25.6005
R27942 GND.n9502 GND.n9501 25.6005
R27943 GND.n9501 GND.n9500 25.6005
R27944 GND.n9500 GND.n9497 25.6005
R27945 GND.n9497 GND.n9496 25.6005
R27946 GND.n9496 GND.n9493 25.6005
R27947 GND.n9493 GND.n9492 25.6005
R27948 GND.n9492 GND.n9489 25.6005
R27949 GND.n9489 GND.n9488 25.6005
R27950 GND.n9488 GND.n9485 25.6005
R27951 GND.n9485 GND.n9484 25.6005
R27952 GND.n9484 GND.n9481 25.6005
R27953 GND.n9481 GND.n9480 25.6005
R27954 GND.n9480 GND.n9477 25.6005
R27955 GND.n9477 GND.n9476 25.6005
R27956 GND.n9509 GND.n9508 25.6005
R27957 GND.n9509 GND.n179 25.6005
R27958 GND.n9538 GND.n179 25.6005
R27959 GND.n9538 GND.n9537 25.6005
R27960 GND.n9537 GND.n9536 25.6005
R27961 GND.n9536 GND.n180 25.6005
R27962 GND.n9523 GND.n180 25.6005
R27963 GND.n9524 GND.n9523 25.6005
R27964 GND.n9524 GND.n72 25.6005
R27965 GND.n144 GND.n142 25.6005
R27966 GND.n145 GND.n144 25.6005
R27967 GND.n9747 GND.n79 25.6005
R27968 GND.n9747 GND.n9746 25.6005
R27969 GND.n9746 GND.n9745 25.6005
R27970 GND.n9745 GND.n80 25.6005
R27971 GND.n99 GND.n80 25.6005
R27972 GND.n9731 GND.n9730 25.6005
R27973 GND.n9730 GND.n9729 25.6005
R27974 GND.n9716 GND.n9715 25.6005
R27975 GND.n9715 GND.n9713 25.6005
R27976 GND.n158 GND.n157 25.6005
R27977 GND.n157 GND.n156 25.6005
R27978 GND.n156 GND.n151 25.6005
R27979 GND.n151 GND.n102 25.6005
R27980 GND.n9712 GND.n102 25.6005
R27981 GND.n9594 GND.n9593 25.6005
R27982 GND.n9593 GND.n9592 25.6005
R27983 GND.n9402 GND.n231 25.6005
R27984 GND.n9402 GND.n9401 25.6005
R27985 GND.n9401 GND.n9400 25.6005
R27986 GND.n9383 GND.n254 25.6005
R27987 GND.n9373 GND.n254 25.6005
R27988 GND.n9356 GND.n9355 25.6005
R27989 GND.n9355 GND.n9354 25.6005
R27990 GND.n9354 GND.n293 25.6005
R27991 GND.n756 GND.n754 25.6005
R27992 GND.n757 GND.n756 25.6005
R27993 GND.n760 GND.n757 25.6005
R27994 GND.n761 GND.n760 25.6005
R27995 GND.n764 GND.n761 25.6005
R27996 GND.n765 GND.n764 25.6005
R27997 GND.n768 GND.n765 25.6005
R27998 GND.n769 GND.n768 25.6005
R27999 GND.n772 GND.n769 25.6005
R28000 GND.n773 GND.n772 25.6005
R28001 GND.n776 GND.n773 25.6005
R28002 GND.n777 GND.n776 25.6005
R28003 GND.n780 GND.n777 25.6005
R28004 GND.n781 GND.n780 25.6005
R28005 GND.n784 GND.n781 25.6005
R28006 GND.n785 GND.n784 25.6005
R28007 GND.n789 GND.n788 25.6005
R28008 GND.n788 GND.n787 25.6005
R28009 GND.n787 GND.n786 25.6005
R28010 GND.n961 GND.n959 25.6005
R28011 GND.n962 GND.n961 25.6005
R28012 GND.n968 GND.n967 25.6005
R28013 GND.n967 GND.n966 25.6005
R28014 GND.n966 GND.n320 25.6005
R28015 GND.n9342 GND.n9341 25.6005
R28016 GND.n9341 GND.n9340 25.6005
R28017 GND.n9340 GND.n9339 25.6005
R28018 GND.n9339 GND.n9337 25.6005
R28019 GND.n9337 GND.n9334 25.6005
R28020 GND.n9334 GND.n9333 25.6005
R28021 GND.n9333 GND.n9330 25.6005
R28022 GND.n9330 GND.n9329 25.6005
R28023 GND.n9329 GND.n9326 25.6005
R28024 GND.n9326 GND.n9325 25.6005
R28025 GND.n9325 GND.n9322 25.6005
R28026 GND.n9322 GND.n9321 25.6005
R28027 GND.n9321 GND.n9318 25.6005
R28028 GND.n9318 GND.n9317 25.6005
R28029 GND.n9317 GND.n9314 25.6005
R28030 GND.n9314 GND.n9313 25.6005
R28031 GND.n795 GND.n794 25.6005
R28032 GND.n798 GND.n795 25.6005
R28033 GND.n799 GND.n798 25.6005
R28034 GND.n802 GND.n799 25.6005
R28035 GND.n803 GND.n802 25.6005
R28036 GND.n806 GND.n803 25.6005
R28037 GND.n807 GND.n806 25.6005
R28038 GND.n810 GND.n807 25.6005
R28039 GND.n811 GND.n810 25.6005
R28040 GND.n814 GND.n811 25.6005
R28041 GND.n815 GND.n814 25.6005
R28042 GND.n818 GND.n815 25.6005
R28043 GND.n819 GND.n818 25.6005
R28044 GND.n822 GND.n819 25.6005
R28045 GND.n823 GND.n822 25.6005
R28046 GND.n854 GND.n823 25.6005
R28047 GND.n524 GND.n523 25.6005
R28048 GND.n523 GND.n239 25.6005
R28049 GND.n9396 GND.n239 25.6005
R28050 GND.n9379 GND.n9378 25.6005
R28051 GND.n9378 GND.n9377 25.6005
R28052 GND.n9360 GND.n284 25.6005
R28053 GND.n9350 GND.n284 25.6005
R28054 GND.n9350 GND.n9349 25.6005
R28055 GND.n9348 GND.n299 25.6005
R28056 GND.n8984 GND.n299 25.6005
R28057 GND.n8985 GND.n8984 25.6005
R28058 GND.n8988 GND.n8985 25.6005
R28059 GND.n8989 GND.n8988 25.6005
R28060 GND.n8992 GND.n8989 25.6005
R28061 GND.n8993 GND.n8992 25.6005
R28062 GND.n8996 GND.n8993 25.6005
R28063 GND.n8997 GND.n8996 25.6005
R28064 GND.n9000 GND.n8997 25.6005
R28065 GND.n9001 GND.n9000 25.6005
R28066 GND.n9004 GND.n9001 25.6005
R28067 GND.n9005 GND.n9004 25.6005
R28068 GND.n9008 GND.n9005 25.6005
R28069 GND.n9010 GND.n9008 25.6005
R28070 GND.n9011 GND.n9010 25.6005
R28071 GND.n853 GND.n852 25.6005
R28072 GND.n852 GND.n851 25.6005
R28073 GND.n851 GND.n850 25.6005
R28074 GND.n9024 GND.n8979 25.6005
R28075 GND.n9024 GND.n9023 25.6005
R28076 GND.n9015 GND.n9014 25.6005
R28077 GND.n9014 GND.n9013 25.6005
R28078 GND.n9013 GND.n9012 25.6005
R28079 GND.n680 GND.n564 25.6005
R28080 GND.n675 GND.n564 25.6005
R28081 GND.n675 GND.n674 25.6005
R28082 GND.n674 GND.n673 25.6005
R28083 GND.n673 GND.n670 25.6005
R28084 GND.n670 GND.n669 25.6005
R28085 GND.n669 GND.n666 25.6005
R28086 GND.n666 GND.n665 25.6005
R28087 GND.n665 GND.n662 25.6005
R28088 GND.n662 GND.n661 25.6005
R28089 GND.n661 GND.n658 25.6005
R28090 GND.n658 GND.n657 25.6005
R28091 GND.n657 GND.n654 25.6005
R28092 GND.n654 GND.n653 25.6005
R28093 GND.n653 GND.n650 25.6005
R28094 GND.n650 GND.n649 25.6005
R28095 GND.n683 GND.n681 25.6005
R28096 GND.n683 GND.n682 25.6005
R28097 GND.n682 GND.n544 25.6005
R28098 GND.n706 GND.n544 25.6005
R28099 GND.n707 GND.n706 25.6005
R28100 GND.n709 GND.n707 25.6005
R28101 GND.n709 GND.n708 25.6005
R28102 GND.n708 GND.n194 25.6005
R28103 GND.n9429 GND.n194 25.6005
R28104 GND.n9429 GND.n9428 25.6005
R28105 GND.n9428 GND.n9427 25.6005
R28106 GND.n9028 GND.n458 25.6005
R28107 GND.n9028 GND.n9027 25.6005
R28108 GND.n387 GND.n339 25.6005
R28109 GND.n388 GND.n387 25.6005
R28110 GND.n9232 GND.n388 25.6005
R28111 GND.n9232 GND.n9231 25.6005
R28112 GND.n9231 GND.n9230 25.6005
R28113 GND.n9230 GND.n389 25.6005
R28114 GND.n406 GND.n389 25.6005
R28115 GND.n9218 GND.n406 25.6005
R28116 GND.n9218 GND.n9217 25.6005
R28117 GND.n9217 GND.n9216 25.6005
R28118 GND.n9216 GND.n407 25.6005
R28119 GND.n9132 GND.n9131 25.6005
R28120 GND.n9131 GND.n9130 25.6005
R28121 GND.n9130 GND.n9129 25.6005
R28122 GND.n9129 GND.n9127 25.6005
R28123 GND.n9127 GND.n9124 25.6005
R28124 GND.n9124 GND.n9123 25.6005
R28125 GND.n9123 GND.n9120 25.6005
R28126 GND.n9120 GND.n9119 25.6005
R28127 GND.n9119 GND.n9116 25.6005
R28128 GND.n9116 GND.n9115 25.6005
R28129 GND.n9115 GND.n9112 25.6005
R28130 GND.n9112 GND.n9111 25.6005
R28131 GND.n9111 GND.n9108 25.6005
R28132 GND.n9108 GND.n9107 25.6005
R28133 GND.n9107 GND.n9104 25.6005
R28134 GND.n9104 GND.n9103 25.6005
R28135 GND.n687 GND.n557 25.6005
R28136 GND.n688 GND.n687 25.6005
R28137 GND.n693 GND.n688 25.6005
R28138 GND.n693 GND.n692 25.6005
R28139 GND.n692 GND.n691 25.6005
R28140 GND.n691 GND.n689 25.6005
R28141 GND.n689 GND.n528 25.6005
R28142 GND.n733 GND.n528 25.6005
R28143 GND.n734 GND.n733 25.6005
R28144 GND.n737 GND.n734 25.6005
R28145 GND.n738 GND.n737 25.6005
R28146 GND.n484 GND.n455 25.6005
R28147 GND.n9033 GND.n455 25.6005
R28148 GND.n9081 GND.n427 25.6005
R28149 GND.n9085 GND.n427 25.6005
R28150 GND.n9086 GND.n9085 25.6005
R28151 GND.n9089 GND.n9086 25.6005
R28152 GND.n9090 GND.n9089 25.6005
R28153 GND.n9091 GND.n9090 25.6005
R28154 GND.n9094 GND.n9091 25.6005
R28155 GND.n9095 GND.n9094 25.6005
R28156 GND.n9098 GND.n9095 25.6005
R28157 GND.n9099 GND.n9098 25.6005
R28158 GND.n9100 GND.n9099 25.6005
R28159 GND.n613 GND.n612 25.6005
R28160 GND.n612 GND.n611 25.6005
R28161 GND.n611 GND.n608 25.6005
R28162 GND.n608 GND.n607 25.6005
R28163 GND.n607 GND.n604 25.6005
R28164 GND.n604 GND.n603 25.6005
R28165 GND.n603 GND.n600 25.6005
R28166 GND.n600 GND.n599 25.6005
R28167 GND.n599 GND.n596 25.6005
R28168 GND.n596 GND.n595 25.6005
R28169 GND.n595 GND.n592 25.6005
R28170 GND.n592 GND.n591 25.6005
R28171 GND.n591 GND.n588 25.6005
R28172 GND.n588 GND.n587 25.6005
R28173 GND.n587 GND.n576 25.6005
R28174 GND.n618 GND.n576 25.6005
R28175 GND.n634 GND.n571 25.6005
R28176 GND.n635 GND.n634 25.6005
R28177 GND.n637 GND.n635 25.6005
R28178 GND.n637 GND.n636 25.6005
R28179 GND.n636 GND.n553 25.6005
R28180 GND.n698 GND.n553 25.6005
R28181 GND.n699 GND.n698 25.6005
R28182 GND.n701 GND.n699 25.6005
R28183 GND.n701 GND.n700 25.6005
R28184 GND.n700 GND.n534 25.6005
R28185 GND.n728 GND.n534 25.6005
R28186 GND.n728 GND.n727 25.6005
R28187 GND.n727 GND.n726 25.6005
R28188 GND.n889 GND.n469 25.6005
R28189 GND.n9238 GND.n9237 25.6005
R28190 GND.n9237 GND.n376 25.6005
R28191 GND.n397 GND.n376 25.6005
R28192 GND.n9225 GND.n397 25.6005
R28193 GND.n9225 GND.n9224 25.6005
R28194 GND.n9224 GND.n9223 25.6005
R28195 GND.n9223 GND.n398 25.6005
R28196 GND.n415 GND.n398 25.6005
R28197 GND.n9211 GND.n415 25.6005
R28198 GND.n9211 GND.n9210 25.6005
R28199 GND.n9210 GND.n9209 25.6005
R28200 GND.n9209 GND.n416 25.6005
R28201 GND.n9203 GND.n416 25.6005
R28202 GND.n9202 GND.n9201 25.6005
R28203 GND.n9201 GND.n9140 25.6005
R28204 GND.n9196 GND.n9140 25.6005
R28205 GND.n9196 GND.n9195 25.6005
R28206 GND.n9195 GND.n9142 25.6005
R28207 GND.n9190 GND.n9142 25.6005
R28208 GND.n9190 GND.n9189 25.6005
R28209 GND.n9189 GND.n9188 25.6005
R28210 GND.n9188 GND.n9144 25.6005
R28211 GND.n9182 GND.n9144 25.6005
R28212 GND.n9182 GND.n9181 25.6005
R28213 GND.n9181 GND.n9180 25.6005
R28214 GND.n9180 GND.n9146 25.6005
R28215 GND.n9174 GND.n9146 25.6005
R28216 GND.n9174 GND.n9173 25.6005
R28217 GND.n9173 GND.n9172 25.6005
R28218 GND.n630 GND.n619 25.6005
R28219 GND.n630 GND.n629 25.6005
R28220 GND.n629 GND.n628 25.6005
R28221 GND.n628 GND.n627 25.6005
R28222 GND.n627 GND.n624 25.6005
R28223 GND.n624 GND.n623 25.6005
R28224 GND.n623 GND.n622 25.6005
R28225 GND.n622 GND.n620 25.6005
R28226 GND.n620 GND.n539 25.6005
R28227 GND.n714 GND.n539 25.6005
R28228 GND.n715 GND.n714 25.6005
R28229 GND.n716 GND.n715 25.6005
R28230 GND.n722 GND.n716 25.6005
R28231 GND.n894 GND.n876 25.6005
R28232 GND.n9149 GND.n9148 25.6005
R28233 GND.n9150 GND.n9149 25.6005
R28234 GND.n9153 GND.n9150 25.6005
R28235 GND.n9154 GND.n9153 25.6005
R28236 GND.n9157 GND.n9154 25.6005
R28237 GND.n9158 GND.n9157 25.6005
R28238 GND.n9159 GND.n9158 25.6005
R28239 GND.n9162 GND.n9159 25.6005
R28240 GND.n9163 GND.n9162 25.6005
R28241 GND.n9166 GND.n9163 25.6005
R28242 GND.n9167 GND.n9166 25.6005
R28243 GND.n9168 GND.n9167 25.6005
R28244 GND.n9169 GND.n9168 25.6005
R28245 GND.n8495 GND.n8494 25.6005
R28246 GND.n8494 GND.n8493 25.6005
R28247 GND.n8493 GND.n8491 25.6005
R28248 GND.n8491 GND.n8490 25.6005
R28249 GND.n8490 GND.n8488 25.6005
R28250 GND.n8488 GND.n8487 25.6005
R28251 GND.n8487 GND.n8485 25.6005
R28252 GND.n8485 GND.n8484 25.6005
R28253 GND.n8484 GND.n8482 25.6005
R28254 GND.n8482 GND.n8481 25.6005
R28255 GND.n8481 GND.n8479 25.6005
R28256 GND.n8479 GND.n8478 25.6005
R28257 GND.n8478 GND.n8476 25.6005
R28258 GND.n8476 GND.n8475 25.6005
R28259 GND.n8475 GND.n1751 25.6005
R28260 GND.n8444 GND.n8443 25.6005
R28261 GND.n8447 GND.n8444 25.6005
R28262 GND.n8448 GND.n8447 25.6005
R28263 GND.n8451 GND.n8448 25.6005
R28264 GND.n8452 GND.n8451 25.6005
R28265 GND.n8455 GND.n8452 25.6005
R28266 GND.n8456 GND.n8455 25.6005
R28267 GND.n8459 GND.n8456 25.6005
R28268 GND.n8460 GND.n8459 25.6005
R28269 GND.n8463 GND.n8460 25.6005
R28270 GND.n8464 GND.n8463 25.6005
R28271 GND.n8467 GND.n8464 25.6005
R28272 GND.n8468 GND.n8467 25.6005
R28273 GND.n8471 GND.n8468 25.6005
R28274 GND.n8473 GND.n8471 25.6005
R28275 GND.n8474 GND.n8473 25.6005
R28276 GND.n8496 GND.n8474 25.6005
R28277 GND.n8597 GND.n1793 25.6005
R28278 GND.n8598 GND.n8597 25.6005
R28279 GND.n8599 GND.n8598 25.6005
R28280 GND.n8599 GND.n1781 25.6005
R28281 GND.n8609 GND.n1781 25.6005
R28282 GND.n8610 GND.n8609 25.6005
R28283 GND.n8611 GND.n8610 25.6005
R28284 GND.n8611 GND.n1769 25.6005
R28285 GND.n8621 GND.n1769 25.6005
R28286 GND.n8622 GND.n8621 25.6005
R28287 GND.n8623 GND.n8622 25.6005
R28288 GND.n8623 GND.n1756 25.6005
R28289 GND.n8635 GND.n1756 25.6005
R28290 GND.n8636 GND.n8635 25.6005
R28291 GND.n8637 GND.n8636 25.6005
R28292 GND.n8637 GND.n1743 25.6005
R28293 GND.n8649 GND.n1743 25.6005
R28294 GND.n8650 GND.n8649 25.6005
R28295 GND.n8651 GND.n8650 25.6005
R28296 GND.n8651 GND.n1731 25.6005
R28297 GND.n8662 GND.n1731 25.6005
R28298 GND.n8663 GND.n8662 25.6005
R28299 GND.n8664 GND.n8663 25.6005
R28300 GND.n8664 GND.n1010 25.6005
R28301 GND.n8781 GND.n1010 25.6005
R28302 GND.n8781 GND.n8780 25.6005
R28303 GND.n8780 GND.n8779 25.6005
R28304 GND.n8779 GND.n1011 25.6005
R28305 GND.n8769 GND.n1011 25.6005
R28306 GND.n8769 GND.n8768 25.6005
R28307 GND.n8768 GND.n8767 25.6005
R28308 GND.n8767 GND.n1025 25.6005
R28309 GND.n8757 GND.n1025 25.6005
R28310 GND.n8757 GND.n8756 25.6005
R28311 GND.n8756 GND.n8755 25.6005
R28312 GND.n8755 GND.n1037 25.6005
R28313 GND.n8745 GND.n1037 25.6005
R28314 GND.n8745 GND.n8744 25.6005
R28315 GND.n8744 GND.n8743 25.6005
R28316 GND.n8743 GND.n1049 25.6005
R28317 GND.n8733 GND.n1049 25.6005
R28318 GND.n8733 GND.n8732 25.6005
R28319 GND.n8731 GND.n1061 25.6005
R28320 GND.n8726 GND.n1061 25.6005
R28321 GND.n8726 GND.n8725 25.6005
R28322 GND.n8725 GND.n8724 25.6005
R28323 GND.n8724 GND.n8721 25.6005
R28324 GND.n8721 GND.n8720 25.6005
R28325 GND.n8720 GND.n8717 25.6005
R28326 GND.n8717 GND.n8716 25.6005
R28327 GND.n8716 GND.n8713 25.6005
R28328 GND.n8713 GND.n8712 25.6005
R28329 GND.n8712 GND.n8709 25.6005
R28330 GND.n8709 GND.n8708 25.6005
R28331 GND.n8708 GND.n8705 25.6005
R28332 GND.n8705 GND.n8704 25.6005
R28333 GND.n8704 GND.n8701 25.6005
R28334 GND.n8701 GND.n8700 25.6005
R28335 GND.n8700 GND.n8698 25.6005
R28336 GND.n8775 GND.n1018 25.6005
R28337 GND.n8775 GND.n8774 25.6005
R28338 GND.n8774 GND.n8773 25.6005
R28339 GND.n8773 GND.n1019 25.6005
R28340 GND.n8763 GND.n1019 25.6005
R28341 GND.n8763 GND.n8762 25.6005
R28342 GND.n8762 GND.n8761 25.6005
R28343 GND.n8761 GND.n1031 25.6005
R28344 GND.n8751 GND.n1031 25.6005
R28345 GND.n8751 GND.n8750 25.6005
R28346 GND.n8750 GND.n8749 25.6005
R28347 GND.n8749 GND.n1043 25.6005
R28348 GND.n8739 GND.n1043 25.6005
R28349 GND.n8739 GND.n8738 25.6005
R28350 GND.n8738 GND.n8737 25.6005
R28351 GND.n8737 GND.n1055 25.6005
R28352 GND.n8674 GND.n8673 25.6005
R28353 GND.n8676 GND.n8674 25.6005
R28354 GND.n8677 GND.n8676 25.6005
R28355 GND.n8679 GND.n8677 25.6005
R28356 GND.n8680 GND.n8679 25.6005
R28357 GND.n8682 GND.n8680 25.6005
R28358 GND.n8683 GND.n8682 25.6005
R28359 GND.n8685 GND.n8683 25.6005
R28360 GND.n8686 GND.n8685 25.6005
R28361 GND.n8688 GND.n8686 25.6005
R28362 GND.n8689 GND.n8688 25.6005
R28363 GND.n8691 GND.n8689 25.6005
R28364 GND.n8692 GND.n8691 25.6005
R28365 GND.n8694 GND.n8692 25.6005
R28366 GND.n8695 GND.n8694 25.6005
R28367 GND.n8697 GND.n8695 25.6005
R28368 GND.n8593 GND.n8592 25.6005
R28369 GND.n8593 GND.n1787 25.6005
R28370 GND.n8603 GND.n1787 25.6005
R28371 GND.n8604 GND.n8603 25.6005
R28372 GND.n8605 GND.n8604 25.6005
R28373 GND.n8605 GND.n1775 25.6005
R28374 GND.n8615 GND.n1775 25.6005
R28375 GND.n8616 GND.n8615 25.6005
R28376 GND.n8617 GND.n8616 25.6005
R28377 GND.n8617 GND.n1763 25.6005
R28378 GND.n8627 GND.n1763 25.6005
R28379 GND.n8628 GND.n8627 25.6005
R28380 GND.n8631 GND.n8628 25.6005
R28381 GND.n8631 GND.n8630 25.6005
R28382 GND.n8630 GND.n8629 25.6005
R28383 GND.n8591 GND.n1799 25.6005
R28384 GND.n8500 GND.n1799 25.6005
R28385 GND.n8584 GND.n8500 25.6005
R28386 GND.n8584 GND.n8583 25.6005
R28387 GND.n8583 GND.n8582 25.6005
R28388 GND.n8582 GND.n8502 25.6005
R28389 GND.n8577 GND.n8502 25.6005
R28390 GND.n8577 GND.n8576 25.6005
R28391 GND.n8576 GND.n8575 25.6005
R28392 GND.n8575 GND.n8505 25.6005
R28393 GND.n8570 GND.n8505 25.6005
R28394 GND.n8570 GND.n8569 25.6005
R28395 GND.n8569 GND.n8568 25.6005
R28396 GND.n8568 GND.n8508 25.6005
R28397 GND.n8563 GND.n8508 25.6005
R28398 GND.n8563 GND.n8562 25.6005
R28399 GND.n8562 GND.n8561 25.6005
R28400 GND.n8557 GND.n8556 25.6005
R28401 GND.n8556 GND.n8555 25.6005
R28402 GND.n8555 GND.n8553 25.6005
R28403 GND.n8553 GND.n8552 25.6005
R28404 GND.n8552 GND.n8550 25.6005
R28405 GND.n8550 GND.n8549 25.6005
R28406 GND.n8549 GND.n8547 25.6005
R28407 GND.n8547 GND.n8546 25.6005
R28408 GND.n8546 GND.n8544 25.6005
R28409 GND.n8544 GND.n8543 25.6005
R28410 GND.n8543 GND.n8541 25.6005
R28411 GND.n8541 GND.n8540 25.6005
R28412 GND.n8540 GND.n8538 25.6005
R28413 GND.n8538 GND.n8537 25.6005
R28414 GND.n8537 GND.n8535 25.6005
R28415 GND.n8525 GND.n8524 25.6005
R28416 GND.n8524 GND.n8522 25.6005
R28417 GND.n8785 GND.n1001 25.6005
R28418 GND.n1663 GND.n1001 25.6005
R28419 GND.n1665 GND.n1663 25.6005
R28420 GND.n1666 GND.n1665 25.6005
R28421 GND.n1668 GND.n1666 25.6005
R28422 GND.n1669 GND.n1668 25.6005
R28423 GND.n1671 GND.n1669 25.6005
R28424 GND.n1672 GND.n1671 25.6005
R28425 GND.n1674 GND.n1672 25.6005
R28426 GND.n1675 GND.n1674 25.6005
R28427 GND.n1677 GND.n1675 25.6005
R28428 GND.n1678 GND.n1677 25.6005
R28429 GND.n1680 GND.n1678 25.6005
R28430 GND.n1681 GND.n1680 25.6005
R28431 GND.n1683 GND.n1681 25.6005
R28432 GND.n1684 GND.n1683 25.6005
R28433 GND.n1685 GND.n1684 25.6005
R28434 GND.n1720 GND.n1719 25.6005
R28435 GND.n1719 GND.n1718 25.6005
R28436 GND.n1718 GND.n1716 25.6005
R28437 GND.n1716 GND.n1713 25.6005
R28438 GND.n1713 GND.n1712 25.6005
R28439 GND.n1712 GND.n1709 25.6005
R28440 GND.n1709 GND.n1708 25.6005
R28441 GND.n1708 GND.n1705 25.6005
R28442 GND.n1705 GND.n1704 25.6005
R28443 GND.n1704 GND.n1701 25.6005
R28444 GND.n1701 GND.n1700 25.6005
R28445 GND.n1700 GND.n1697 25.6005
R28446 GND.n1697 GND.n1696 25.6005
R28447 GND.n1696 GND.n1693 25.6005
R28448 GND.n1693 GND.n1692 25.6005
R28449 GND.n1692 GND.n1689 25.6005
R28450 GND.n1689 GND.n1688 25.6005
R28451 GND.n3234 GND.n3232 25.6005
R28452 GND.n3235 GND.n3234 25.6005
R28453 GND.n3237 GND.n3235 25.6005
R28454 GND.n3238 GND.n3237 25.6005
R28455 GND.n3240 GND.n3238 25.6005
R28456 GND.n3241 GND.n3240 25.6005
R28457 GND.n3243 GND.n3241 25.6005
R28458 GND.n3244 GND.n3243 25.6005
R28459 GND.n3246 GND.n3244 25.6005
R28460 GND.n3247 GND.n3246 25.6005
R28461 GND.n3249 GND.n3247 25.6005
R28462 GND.n3250 GND.n3249 25.6005
R28463 GND.n3252 GND.n3250 25.6005
R28464 GND.n3253 GND.n3252 25.6005
R28465 GND.n3255 GND.n3253 25.6005
R28466 GND.n3256 GND.n3255 25.6005
R28467 GND.n3258 GND.n3256 25.6005
R28468 GND.n3198 GND.n3141 25.6005
R28469 GND.n3201 GND.n3198 25.6005
R28470 GND.n3202 GND.n3201 25.6005
R28471 GND.n3205 GND.n3202 25.6005
R28472 GND.n3206 GND.n3205 25.6005
R28473 GND.n3209 GND.n3206 25.6005
R28474 GND.n3210 GND.n3209 25.6005
R28475 GND.n3213 GND.n3210 25.6005
R28476 GND.n3214 GND.n3213 25.6005
R28477 GND.n3217 GND.n3214 25.6005
R28478 GND.n3218 GND.n3217 25.6005
R28479 GND.n3221 GND.n3218 25.6005
R28480 GND.n3222 GND.n3221 25.6005
R28481 GND.n3225 GND.n3222 25.6005
R28482 GND.n3226 GND.n3225 25.6005
R28483 GND.n3229 GND.n3226 25.6005
R28484 GND.n3231 GND.n3229 25.6005
R28485 GND.n3693 GND.n3692 25.6005
R28486 GND.n3692 GND.n3691 25.6005
R28487 GND.n3691 GND.n3142 25.6005
R28488 GND.n3681 GND.n3142 25.6005
R28489 GND.n3681 GND.n3680 25.6005
R28490 GND.n3680 GND.n3679 25.6005
R28491 GND.n3679 GND.n3156 25.6005
R28492 GND.n3669 GND.n3156 25.6005
R28493 GND.n3669 GND.n3668 25.6005
R28494 GND.n3668 GND.n3667 25.6005
R28495 GND.n3667 GND.n3168 25.6005
R28496 GND.n3657 GND.n3168 25.6005
R28497 GND.n3657 GND.n3656 25.6005
R28498 GND.n3656 GND.n3655 25.6005
R28499 GND.n3655 GND.n3180 25.6005
R28500 GND.n3645 GND.n3180 25.6005
R28501 GND.n3645 GND.n3644 25.6005
R28502 GND.n3644 GND.n3643 25.6005
R28503 GND.n3643 GND.n3192 25.6005
R28504 GND.n3633 GND.n3192 25.6005
R28505 GND.n3633 GND.n3632 25.6005
R28506 GND.n3632 GND.n3631 25.6005
R28507 GND.n3631 GND.n3265 25.6005
R28508 GND.n3621 GND.n3265 25.6005
R28509 GND.n3621 GND.n3620 25.6005
R28510 GND.n3620 GND.n3619 25.6005
R28511 GND.n3619 GND.n3279 25.6005
R28512 GND.n3609 GND.n3279 25.6005
R28513 GND.n3609 GND.n3608 25.6005
R28514 GND.n3608 GND.n3607 25.6005
R28515 GND.n3607 GND.n3294 25.6005
R28516 GND.n3597 GND.n3294 25.6005
R28517 GND.n3597 GND.n3596 25.6005
R28518 GND.n3596 GND.n3595 25.6005
R28519 GND.n3595 GND.n3309 25.6005
R28520 GND.n3585 GND.n3309 25.6005
R28521 GND.n3585 GND.n3584 25.6005
R28522 GND.n3584 GND.n3583 25.6005
R28523 GND.n3583 GND.n3321 25.6005
R28524 GND.n3573 GND.n3321 25.6005
R28525 GND.n3573 GND.n3572 25.6005
R28526 GND.n3572 GND.n3571 25.6005
R28527 GND.n3396 GND.n3333 25.6005
R28528 GND.n3396 GND.n3395 25.6005
R28529 GND.n3395 GND.n3394 25.6005
R28530 GND.n3394 GND.n3392 25.6005
R28531 GND.n3392 GND.n3389 25.6005
R28532 GND.n3389 GND.n3388 25.6005
R28533 GND.n3388 GND.n3385 25.6005
R28534 GND.n3385 GND.n3384 25.6005
R28535 GND.n3384 GND.n3381 25.6005
R28536 GND.n3381 GND.n3380 25.6005
R28537 GND.n3380 GND.n3377 25.6005
R28538 GND.n3377 GND.n3376 25.6005
R28539 GND.n3376 GND.n3373 25.6005
R28540 GND.n3373 GND.n3372 25.6005
R28541 GND.n3372 GND.n3369 25.6005
R28542 GND.n3369 GND.n3368 25.6005
R28543 GND.n3368 GND.n3366 25.6005
R28544 GND.n3495 GND.n3494 25.6005
R28545 GND.n3494 GND.n3492 25.6005
R28546 GND.n3511 GND.n3509 25.6005
R28547 GND.n3512 GND.n3511 25.6005
R28548 GND.n3514 GND.n3512 25.6005
R28549 GND.n3515 GND.n3514 25.6005
R28550 GND.n3517 GND.n3515 25.6005
R28551 GND.n3518 GND.n3517 25.6005
R28552 GND.n3520 GND.n3518 25.6005
R28553 GND.n3521 GND.n3520 25.6005
R28554 GND.n3523 GND.n3521 25.6005
R28555 GND.n3524 GND.n3523 25.6005
R28556 GND.n3526 GND.n3524 25.6005
R28557 GND.n3527 GND.n3526 25.6005
R28558 GND.n3529 GND.n3527 25.6005
R28559 GND.n3530 GND.n3529 25.6005
R28560 GND.n3566 GND.n3565 25.6005
R28561 GND.n3565 GND.n3401 25.6005
R28562 GND.n3559 GND.n3401 25.6005
R28563 GND.n3559 GND.n3558 25.6005
R28564 GND.n3558 GND.n3557 25.6005
R28565 GND.n3557 GND.n3403 25.6005
R28566 GND.n3551 GND.n3403 25.6005
R28567 GND.n3551 GND.n3550 25.6005
R28568 GND.n3550 GND.n3549 25.6005
R28569 GND.n3549 GND.n3405 25.6005
R28570 GND.n3543 GND.n3405 25.6005
R28571 GND.n3543 GND.n3542 25.6005
R28572 GND.n3542 GND.n3541 25.6005
R28573 GND.n3541 GND.n3407 25.6005
R28574 GND.n3535 GND.n3407 25.6005
R28575 GND.n3535 GND.n3534 25.6005
R28576 GND.n3534 GND.n3533 25.6005
R28577 GND.n3302 GND.n3301 25.6005
R28578 GND.n3603 GND.n3302 25.6005
R28579 GND.n3603 GND.n3602 25.6005
R28580 GND.n3602 GND.n3601 25.6005
R28581 GND.n3601 GND.n3303 25.6005
R28582 GND.n3591 GND.n3303 25.6005
R28583 GND.n3591 GND.n3590 25.6005
R28584 GND.n3590 GND.n3589 25.6005
R28585 GND.n3589 GND.n3315 25.6005
R28586 GND.n3579 GND.n3315 25.6005
R28587 GND.n3579 GND.n3578 25.6005
R28588 GND.n3578 GND.n3577 25.6005
R28589 GND.n3577 GND.n3327 25.6005
R28590 GND.n3567 GND.n3327 25.6005
R28591 GND.n3346 GND.n3289 25.6005
R28592 GND.n3347 GND.n3346 25.6005
R28593 GND.n3349 GND.n3347 25.6005
R28594 GND.n3350 GND.n3349 25.6005
R28595 GND.n3352 GND.n3350 25.6005
R28596 GND.n3353 GND.n3352 25.6005
R28597 GND.n3355 GND.n3353 25.6005
R28598 GND.n3356 GND.n3355 25.6005
R28599 GND.n3358 GND.n3356 25.6005
R28600 GND.n3359 GND.n3358 25.6005
R28601 GND.n3361 GND.n3359 25.6005
R28602 GND.n3362 GND.n3361 25.6005
R28603 GND.n3364 GND.n3362 25.6005
R28604 GND.n3365 GND.n3364 25.6005
R28605 GND.n3416 GND.n3149 25.6005
R28606 GND.n3687 GND.n3149 25.6005
R28607 GND.n3687 GND.n3686 25.6005
R28608 GND.n3686 GND.n3685 25.6005
R28609 GND.n3685 GND.n3150 25.6005
R28610 GND.n3675 GND.n3150 25.6005
R28611 GND.n3675 GND.n3674 25.6005
R28612 GND.n3674 GND.n3673 25.6005
R28613 GND.n3673 GND.n3162 25.6005
R28614 GND.n3663 GND.n3162 25.6005
R28615 GND.n3663 GND.n3662 25.6005
R28616 GND.n3662 GND.n3661 25.6005
R28617 GND.n3661 GND.n3174 25.6005
R28618 GND.n3651 GND.n3174 25.6005
R28619 GND.n3651 GND.n3650 25.6005
R28620 GND.n3650 GND.n3649 25.6005
R28621 GND.n3649 GND.n3186 25.6005
R28622 GND.n3419 GND.n3418 25.6005
R28623 GND.n3422 GND.n3419 25.6005
R28624 GND.n3423 GND.n3422 25.6005
R28625 GND.n3426 GND.n3423 25.6005
R28626 GND.n3427 GND.n3426 25.6005
R28627 GND.n3430 GND.n3427 25.6005
R28628 GND.n3431 GND.n3430 25.6005
R28629 GND.n3434 GND.n3431 25.6005
R28630 GND.n3435 GND.n3434 25.6005
R28631 GND.n3438 GND.n3435 25.6005
R28632 GND.n3439 GND.n3438 25.6005
R28633 GND.n3442 GND.n3439 25.6005
R28634 GND.n3443 GND.n3442 25.6005
R28635 GND.n3446 GND.n3443 25.6005
R28636 GND.n3447 GND.n3446 25.6005
R28637 GND.n3450 GND.n3447 25.6005
R28638 GND.n3452 GND.n3450 25.6005
R28639 GND.n3455 GND.n3453 25.6005
R28640 GND.n3456 GND.n3455 25.6005
R28641 GND.n3458 GND.n3456 25.6005
R28642 GND.n3459 GND.n3458 25.6005
R28643 GND.n3461 GND.n3459 25.6005
R28644 GND.n3462 GND.n3461 25.6005
R28645 GND.n3464 GND.n3462 25.6005
R28646 GND.n3465 GND.n3464 25.6005
R28647 GND.n3467 GND.n3465 25.6005
R28648 GND.n3468 GND.n3467 25.6005
R28649 GND.n3470 GND.n3468 25.6005
R28650 GND.n3471 GND.n3470 25.6005
R28651 GND.n3473 GND.n3471 25.6005
R28652 GND.n3474 GND.n3473 25.6005
R28653 GND.n3476 GND.n3474 25.6005
R28654 GND.n3477 GND.n3476 25.6005
R28655 GND.n3479 GND.n3477 25.6005
R28656 GND.n3480 GND.n3479 25.6005
R28657 GND.n5843 GND.n5842 25.6005
R28658 GND.n5842 GND.n5841 25.6005
R28659 GND.n5841 GND.n5838 25.6005
R28660 GND.n5838 GND.n5837 25.6005
R28661 GND.n5837 GND.n5834 25.6005
R28662 GND.n5834 GND.n5833 25.6005
R28663 GND.n5833 GND.n5830 25.6005
R28664 GND.n5830 GND.n5829 25.6005
R28665 GND.n5829 GND.n5826 25.6005
R28666 GND.n5826 GND.n5825 25.6005
R28667 GND.n5825 GND.n5822 25.6005
R28668 GND.n5822 GND.n5821 25.6005
R28669 GND.n5821 GND.n5818 25.6005
R28670 GND.n5818 GND.n5817 25.6005
R28671 GND.n5817 GND.n5814 25.6005
R28672 GND.n3738 GND.n3721 25.6005
R28673 GND.n3739 GND.n3738 25.6005
R28674 GND.n5885 GND.n3739 25.6005
R28675 GND.n5885 GND.n5884 25.6005
R28676 GND.n5884 GND.n5883 25.6005
R28677 GND.n5883 GND.n3740 25.6005
R28678 GND.n3757 GND.n3740 25.6005
R28679 GND.n5871 GND.n3757 25.6005
R28680 GND.n5871 GND.n5870 25.6005
R28681 GND.n5870 GND.n5869 25.6005
R28682 GND.n5869 GND.n3758 25.6005
R28683 GND.n3775 GND.n3758 25.6005
R28684 GND.n5857 GND.n3775 25.6005
R28685 GND.n5857 GND.n5856 25.6005
R28686 GND.n5856 GND.n5855 25.6005
R28687 GND.n5855 GND.n3776 25.6005
R28688 GND.n3813 GND.n3776 25.6005
R28689 GND.n5979 GND.n5978 25.6005
R28690 GND.n5978 GND.n5977 25.6005
R28691 GND.n5977 GND.n5976 25.6005
R28692 GND.n5976 GND.n5974 25.6005
R28693 GND.n5974 GND.n5971 25.6005
R28694 GND.n5971 GND.n5970 25.6005
R28695 GND.n5970 GND.n5967 25.6005
R28696 GND.n5967 GND.n5966 25.6005
R28697 GND.n5966 GND.n5963 25.6005
R28698 GND.n5963 GND.n5962 25.6005
R28699 GND.n5962 GND.n5959 25.6005
R28700 GND.n5959 GND.n5958 25.6005
R28701 GND.n5958 GND.n5955 25.6005
R28702 GND.n5955 GND.n5954 25.6005
R28703 GND.n5954 GND.n5951 25.6005
R28704 GND.n5951 GND.n5950 25.6005
R28705 GND.n5950 GND.n5947 25.6005
R28706 GND.n5947 GND.n5946 25.6005
R28707 GND.n5946 GND.n5943 25.6005
R28708 GND.n5943 GND.n5942 25.6005
R28709 GND.n5942 GND.n5939 25.6005
R28710 GND.n5939 GND.n5938 25.6005
R28711 GND.n5938 GND.n5935 25.6005
R28712 GND.n5935 GND.n5934 25.6005
R28713 GND.n5934 GND.n5931 25.6005
R28714 GND.n5931 GND.n5930 25.6005
R28715 GND.n5930 GND.n5927 25.6005
R28716 GND.n5927 GND.n5926 25.6005
R28717 GND.n5926 GND.n5923 25.6005
R28718 GND.n5923 GND.n5922 25.6005
R28719 GND.n5922 GND.n5919 25.6005
R28720 GND.n5919 GND.n5918 25.6005
R28721 GND.n5918 GND.n5915 25.6005
R28722 GND.n5915 GND.n5914 25.6005
R28723 GND.n5914 GND.n5911 25.6005
R28724 GND.n5911 GND.n5910 25.6005
R28725 GND.n5910 GND.n5907 25.6005
R28726 GND.n5907 GND.n5906 25.6005
R28727 GND.n5906 GND.n5903 25.6005
R28728 GND.n5903 GND.n5902 25.6005
R28729 GND.n5902 GND.n5899 25.6005
R28730 GND.n5899 GND.n5898 25.6005
R28731 GND.n3953 GND.n3722 25.6005
R28732 GND.n3955 GND.n3953 25.6005
R28733 GND.n3956 GND.n3955 25.6005
R28734 GND.n3959 GND.n3956 25.6005
R28735 GND.n3960 GND.n3959 25.6005
R28736 GND.n3961 GND.n3960 25.6005
R28737 GND.n3964 GND.n3961 25.6005
R28738 GND.n3965 GND.n3964 25.6005
R28739 GND.n3968 GND.n3965 25.6005
R28740 GND.n3969 GND.n3968 25.6005
R28741 GND.n3970 GND.n3969 25.6005
R28742 GND.n3973 GND.n3970 25.6005
R28743 GND.n3974 GND.n3973 25.6005
R28744 GND.n3977 GND.n3974 25.6005
R28745 GND.n3978 GND.n3977 25.6005
R28746 GND.n3979 GND.n3978 25.6005
R28747 GND.n3979 GND.n3952 25.6005
R28748 GND.n4148 GND.n4145 25.6005
R28749 GND.n4145 GND.n4142 25.6005
R28750 GND.n4142 GND.n4141 25.6005
R28751 GND.n4141 GND.n4138 25.6005
R28752 GND.n4138 GND.n4137 25.6005
R28753 GND.n4137 GND.n4134 25.6005
R28754 GND.n4134 GND.n4133 25.6005
R28755 GND.n4133 GND.n4130 25.6005
R28756 GND.n4130 GND.n4129 25.6005
R28757 GND.n4129 GND.n4126 25.6005
R28758 GND.n4126 GND.n4125 25.6005
R28759 GND.n4125 GND.n4122 25.6005
R28760 GND.n4122 GND.n4121 25.6005
R28761 GND.n4121 GND.n4118 25.6005
R28762 GND.n4118 GND.n4117 25.6005
R28763 GND.n4117 GND.n4114 25.6005
R28764 GND.n4114 GND.n4113 25.6005
R28765 GND.n4082 GND.n4081 25.6005
R28766 GND.n4083 GND.n4082 25.6005
R28767 GND.n4086 GND.n4083 25.6005
R28768 GND.n4087 GND.n4086 25.6005
R28769 GND.n4090 GND.n4087 25.6005
R28770 GND.n4091 GND.n4090 25.6005
R28771 GND.n4092 GND.n4091 25.6005
R28772 GND.n4095 GND.n4092 25.6005
R28773 GND.n4096 GND.n4095 25.6005
R28774 GND.n4099 GND.n4096 25.6005
R28775 GND.n4100 GND.n4099 25.6005
R28776 GND.n4101 GND.n4100 25.6005
R28777 GND.n4104 GND.n4101 25.6005
R28778 GND.n4105 GND.n4104 25.6005
R28779 GND.n4108 GND.n4105 25.6005
R28780 GND.n4109 GND.n4108 25.6005
R28781 GND.n4110 GND.n4109 25.6005
R28782 GND.n4048 GND.n4045 25.6005
R28783 GND.n4049 GND.n4048 25.6005
R28784 GND.n4052 GND.n4049 25.6005
R28785 GND.n4053 GND.n4052 25.6005
R28786 GND.n4056 GND.n4053 25.6005
R28787 GND.n4057 GND.n4056 25.6005
R28788 GND.n4060 GND.n4057 25.6005
R28789 GND.n4061 GND.n4060 25.6005
R28790 GND.n4064 GND.n4061 25.6005
R28791 GND.n4065 GND.n4064 25.6005
R28792 GND.n4068 GND.n4065 25.6005
R28793 GND.n4069 GND.n4068 25.6005
R28794 GND.n4072 GND.n4069 25.6005
R28795 GND.n4073 GND.n4072 25.6005
R28796 GND.n4076 GND.n4073 25.6005
R28797 GND.n4077 GND.n4076 25.6005
R28798 GND.n4015 GND.n4012 25.6005
R28799 GND.n4012 GND.n4011 25.6005
R28800 GND.n4011 GND.n4008 25.6005
R28801 GND.n4008 GND.n4007 25.6005
R28802 GND.n4007 GND.n4004 25.6005
R28803 GND.n4004 GND.n4003 25.6005
R28804 GND.n4003 GND.n4000 25.6005
R28805 GND.n4000 GND.n3999 25.6005
R28806 GND.n3999 GND.n3996 25.6005
R28807 GND.n3996 GND.n3995 25.6005
R28808 GND.n3995 GND.n3992 25.6005
R28809 GND.n3992 GND.n3991 25.6005
R28810 GND.n3991 GND.n3988 25.6005
R28811 GND.n3988 GND.n3987 25.6005
R28812 GND.n3987 GND.n3984 25.6005
R28813 GND.n3984 GND.n3983 25.6005
R28814 GND.n5806 GND.n5805 25.6005
R28815 GND.n5805 GND.n5804 25.6005
R28816 GND.n5804 GND.n5803 25.6005
R28817 GND.n5803 GND.n5801 25.6005
R28818 GND.n5801 GND.n5798 25.6005
R28819 GND.n5798 GND.n5797 25.6005
R28820 GND.n5797 GND.n5794 25.6005
R28821 GND.n5794 GND.n5793 25.6005
R28822 GND.n5793 GND.n5790 25.6005
R28823 GND.n5790 GND.n5789 25.6005
R28824 GND.n5789 GND.n5786 25.6005
R28825 GND.n5786 GND.n5785 25.6005
R28826 GND.n5785 GND.n5782 25.6005
R28827 GND.n5782 GND.n3815 25.6005
R28828 GND.n5812 GND.n3815 25.6005
R28829 GND.n5781 GND.n5780 25.6005
R28830 GND.n5780 GND.n3841 25.6005
R28831 GND.n3858 GND.n3841 25.6005
R28832 GND.n5768 GND.n3858 25.6005
R28833 GND.n5768 GND.n5767 25.6005
R28834 GND.n5767 GND.n5766 25.6005
R28835 GND.n5766 GND.n3859 25.6005
R28836 GND.n3876 GND.n3859 25.6005
R28837 GND.n5754 GND.n3876 25.6005
R28838 GND.n5754 GND.n5753 25.6005
R28839 GND.n5753 GND.n5752 25.6005
R28840 GND.n5752 GND.n3877 25.6005
R28841 GND.n3894 GND.n3877 25.6005
R28842 GND.n5740 GND.n3894 25.6005
R28843 GND.n5740 GND.n5739 25.6005
R28844 GND.n5739 GND.n5738 25.6005
R28845 GND.n5738 GND.n3895 25.6005
R28846 GND.n4980 GND.n4979 25.6005
R28847 GND.n4979 GND.n4978 25.6005
R28848 GND.n4978 GND.n4975 25.6005
R28849 GND.n4975 GND.n4974 25.6005
R28850 GND.n4974 GND.n4971 25.6005
R28851 GND.n4971 GND.n4970 25.6005
R28852 GND.n4970 GND.n4967 25.6005
R28853 GND.n4967 GND.n4966 25.6005
R28854 GND.n4966 GND.n4963 25.6005
R28855 GND.n4963 GND.n4962 25.6005
R28856 GND.n4962 GND.n4959 25.6005
R28857 GND.n4959 GND.n4958 25.6005
R28858 GND.n4958 GND.n4955 25.6005
R28859 GND.n4955 GND.n4954 25.6005
R28860 GND.n4954 GND.n4951 25.6005
R28861 GND.n3942 GND.n3941 25.6005
R28862 GND.n3945 GND.n3942 25.6005
R28863 GND.n7928 GND.n7927 25.6005
R28864 GND.n7927 GND.n7926 25.6005
R28865 GND.n7926 GND.n2188 25.6005
R28866 GND.n2199 GND.n2188 25.6005
R28867 GND.n2199 GND.n2198 25.6005
R28868 GND.n2197 GND.n2196 25.6005
R28869 GND.n7983 GND.n7982 25.6005
R28870 GND.n7837 GND.n7835 25.6005
R28871 GND.n7837 GND.n7836 25.6005
R28872 GND.n7836 GND.n2211 25.6005
R28873 GND.n7876 GND.n2211 25.6005
R28874 GND.n7877 GND.n7876 25.6005
R28875 GND.n7879 GND.n7877 25.6005
R28876 GND.n7879 GND.n7878 25.6005
R28877 GND.n7878 GND.n2171 25.6005
R28878 GND.n7960 GND.n2171 25.6005
R28879 GND.n7960 GND.n7959 25.6005
R28880 GND.n7959 GND.n7958 25.6005
R28881 GND.n7958 GND.n2172 25.6005
R28882 GND.n7907 GND.n2172 25.6005
R28883 GND.n7908 GND.n7907 25.6005
R28884 GND.n7908 GND.n2144 25.6005
R28885 GND.n7834 GND.n2260 25.6005
R28886 GND.n7826 GND.n7825 25.6005
R28887 GND.n7822 GND.n2255 25.6005
R28888 GND.n7842 GND.n2255 25.6005
R28889 GND.n7843 GND.n7842 25.6005
R28890 GND.n7844 GND.n7843 25.6005
R28891 GND.n7847 GND.n7844 25.6005
R28892 GND.n7918 GND.n7913 25.6005
R28893 GND.n7919 GND.n7918 25.6005
R28894 GND.n7921 GND.n7919 25.6005
R28895 GND.n7921 GND.n7920 25.6005
R28896 GND.n7920 GND.n2135 25.6005
R28897 GND.n7989 GND.n2135 25.6005
R28898 GND.n7990 GND.n7989 25.6005
R28899 GND.n7991 GND.n7990 25.6005
R28900 GND.n7991 GND.n2130 25.6005
R28901 GND.n8026 GND.n8025 25.6005
R28902 GND.n8025 GND.n8024 25.6005
R28903 GND.n8024 GND.n8023 25.6005
R28904 GND.n8023 GND.n8021 25.6005
R28905 GND.n8021 GND.n8018 25.6005
R28906 GND.n8018 GND.n8017 25.6005
R28907 GND.n8017 GND.n8014 25.6005
R28908 GND.n8014 GND.n8013 25.6005
R28909 GND.n8013 GND.n8010 25.6005
R28910 GND.n8010 GND.n8009 25.6005
R28911 GND.n8009 GND.n8006 25.6005
R28912 GND.n8006 GND.n8005 25.6005
R28913 GND.n8005 GND.n8002 25.6005
R28914 GND.n8002 GND.n8001 25.6005
R28915 GND.n8001 GND.n7998 25.6005
R28916 GND.n7998 GND.n7997 25.6005
R28917 GND.n7892 GND.n2201 25.6005
R28918 GND.n7896 GND.n2201 25.6005
R28919 GND.n7897 GND.n7896 25.6005
R28920 GND.n7898 GND.n7897 25.6005
R28921 GND.n7903 GND.n7898 25.6005
R28922 GND.n7903 GND.n7902 25.6005
R28923 GND.n7902 GND.n7901 25.6005
R28924 GND.n7901 GND.n7899 25.6005
R28925 GND.n7899 GND.n2131 25.6005
R28926 GND.n7793 GND.n7792 25.6005
R28927 GND.n7805 GND.n7793 25.6005
R28928 GND.n7805 GND.n7804 25.6005
R28929 GND.n7804 GND.n7803 25.6005
R28930 GND.n7803 GND.n7794 25.6005
R28931 GND.n7798 GND.n7794 25.6005
R28932 GND.n7798 GND.n7797 25.6005
R28933 GND.n7797 GND.n7796 25.6005
R28934 GND.n7796 GND.n2205 25.6005
R28935 GND.n7787 GND.n7786 25.6005
R28936 GND.n7786 GND.n7785 25.6005
R28937 GND.n7785 GND.n7782 25.6005
R28938 GND.n7782 GND.n7781 25.6005
R28939 GND.n7781 GND.n7778 25.6005
R28940 GND.n7778 GND.n7777 25.6005
R28941 GND.n7777 GND.n7774 25.6005
R28942 GND.n7774 GND.n7773 25.6005
R28943 GND.n7773 GND.n7770 25.6005
R28944 GND.n7770 GND.n7769 25.6005
R28945 GND.n7769 GND.n7766 25.6005
R28946 GND.n7766 GND.n7765 25.6005
R28947 GND.n7765 GND.n7762 25.6005
R28948 GND.n7762 GND.n7761 25.6005
R28949 GND.n7761 GND.n7758 25.6005
R28950 GND.n7758 GND.n2269 25.6005
R28951 GND.n7810 GND.n2266 25.6005
R28952 GND.n7811 GND.n7810 25.6005
R28953 GND.n7815 GND.n7811 25.6005
R28954 GND.n7815 GND.n7814 25.6005
R28955 GND.n7814 GND.n7813 25.6005
R28956 GND.n7813 GND.n2217 25.6005
R28957 GND.n7869 GND.n2217 25.6005
R28958 GND.n7870 GND.n7869 25.6005
R28959 GND.n7871 GND.n7870 25.6005
R28960 GND.n2234 GND.n2233 25.6005
R28961 GND.n2237 GND.n2234 25.6005
R28962 GND.n2230 GND.n2163 25.6005
R28963 GND.n7967 GND.n2163 25.6005
R28964 GND.n7967 GND.n7966 25.6005
R28965 GND.n7966 GND.n7965 25.6005
R28966 GND.n7965 GND.n2164 25.6005
R28967 GND.n7952 GND.n7951 25.6005
R28968 GND.n7951 GND.n7950 25.6005
R28969 GND.n7937 GND.n7936 25.6005
R28970 GND.n7936 GND.n7934 25.6005
R28971 GND.n7861 GND.n7860 25.6005
R28972 GND.n7860 GND.n7859 25.6005
R28973 GND.n7859 GND.n7858 25.6005
R28974 GND.n7858 GND.n2185 25.6005
R28975 GND.n7933 GND.n2185 25.6005
R28976 GND.n2251 GND.n2250 25.6005
R28977 GND.n7862 GND.n2251 25.6005
R28978 GND.n8296 GND.n1923 25.6005
R28979 GND.n8296 GND.n8295 25.6005
R28980 GND.n8295 GND.n8294 25.6005
R28981 GND.n8277 GND.n1946 25.6005
R28982 GND.n8267 GND.n1946 25.6005
R28983 GND.n8250 GND.n8249 25.6005
R28984 GND.n8249 GND.n8248 25.6005
R28985 GND.n8248 GND.n1985 25.6005
R28986 GND.n4369 GND.n4367 25.6005
R28987 GND.n4370 GND.n4369 25.6005
R28988 GND.n4373 GND.n4370 25.6005
R28989 GND.n4374 GND.n4373 25.6005
R28990 GND.n4377 GND.n4374 25.6005
R28991 GND.n4378 GND.n4377 25.6005
R28992 GND.n4381 GND.n4378 25.6005
R28993 GND.n4382 GND.n4381 25.6005
R28994 GND.n4385 GND.n4382 25.6005
R28995 GND.n4386 GND.n4385 25.6005
R28996 GND.n4389 GND.n4386 25.6005
R28997 GND.n4390 GND.n4389 25.6005
R28998 GND.n4393 GND.n4390 25.6005
R28999 GND.n4395 GND.n4393 25.6005
R29000 GND.n4396 GND.n4395 25.6005
R29001 GND.n4401 GND.n4396 25.6005
R29002 GND.n4400 GND.n4399 25.6005
R29003 GND.n4399 GND.n4398 25.6005
R29004 GND.n4398 GND.n4397 25.6005
R29005 GND.n4712 GND.n4693 25.6005
R29006 GND.n4712 GND.n4711 25.6005
R29007 GND.n4700 GND.n4699 25.6005
R29008 GND.n4699 GND.n4698 25.6005
R29009 GND.n4698 GND.n2012 25.6005
R29010 GND.n8236 GND.n8235 25.6005
R29011 GND.n8235 GND.n8234 25.6005
R29012 GND.n8234 GND.n8233 25.6005
R29013 GND.n8233 GND.n8231 25.6005
R29014 GND.n8231 GND.n8228 25.6005
R29015 GND.n8228 GND.n8227 25.6005
R29016 GND.n8227 GND.n8224 25.6005
R29017 GND.n8224 GND.n8223 25.6005
R29018 GND.n8223 GND.n8220 25.6005
R29019 GND.n8220 GND.n8219 25.6005
R29020 GND.n8219 GND.n8216 25.6005
R29021 GND.n8216 GND.n8215 25.6005
R29022 GND.n8215 GND.n8212 25.6005
R29023 GND.n8212 GND.n8211 25.6005
R29024 GND.n8211 GND.n8208 25.6005
R29025 GND.n8208 GND.n8207 25.6005
R29026 GND.n4444 GND.n4443 25.6005
R29027 GND.n4443 GND.n4268 25.6005
R29028 GND.n4412 GND.n4268 25.6005
R29029 GND.n4415 GND.n4412 25.6005
R29030 GND.n4416 GND.n4415 25.6005
R29031 GND.n4419 GND.n4416 25.6005
R29032 GND.n4420 GND.n4419 25.6005
R29033 GND.n4423 GND.n4420 25.6005
R29034 GND.n4424 GND.n4423 25.6005
R29035 GND.n4427 GND.n4424 25.6005
R29036 GND.n4428 GND.n4427 25.6005
R29037 GND.n4431 GND.n4428 25.6005
R29038 GND.n4432 GND.n4431 25.6005
R29039 GND.n4435 GND.n4432 25.6005
R29040 GND.n4436 GND.n4435 25.6005
R29041 GND.n4438 GND.n4436 25.6005
R29042 GND.n4446 GND.n4445 25.6005
R29043 GND.n4445 GND.n1931 25.6005
R29044 GND.n8290 GND.n1931 25.6005
R29045 GND.n8273 GND.n8272 25.6005
R29046 GND.n8272 GND.n8271 25.6005
R29047 GND.n8254 GND.n1976 25.6005
R29048 GND.n8244 GND.n1976 25.6005
R29049 GND.n8244 GND.n8243 25.6005
R29050 GND.n8242 GND.n1991 25.6005
R29051 GND.n4727 GND.n1991 25.6005
R29052 GND.n4728 GND.n4727 25.6005
R29053 GND.n4731 GND.n4728 25.6005
R29054 GND.n4732 GND.n4731 25.6005
R29055 GND.n4735 GND.n4732 25.6005
R29056 GND.n4736 GND.n4735 25.6005
R29057 GND.n4739 GND.n4736 25.6005
R29058 GND.n4740 GND.n4739 25.6005
R29059 GND.n4743 GND.n4740 25.6005
R29060 GND.n4744 GND.n4743 25.6005
R29061 GND.n4747 GND.n4744 25.6005
R29062 GND.n4748 GND.n4747 25.6005
R29063 GND.n4751 GND.n4748 25.6005
R29064 GND.n4753 GND.n4751 25.6005
R29065 GND.n4754 GND.n4753 25.6005
R29066 GND.n4437 GND.n4254 25.6005
R29067 GND.n4501 GND.n4254 25.6005
R29068 GND.n4501 GND.n4500 25.6005
R29069 GND.n4721 GND.n4204 25.6005
R29070 GND.n4722 GND.n4721 25.6005
R29071 GND.n4758 GND.n4757 25.6005
R29072 GND.n4757 GND.n4756 25.6005
R29073 GND.n4756 GND.n4755 25.6005
R29074 GND.n4286 GND.n1841 25.6005
R29075 GND.n4287 GND.n4286 25.6005
R29076 GND.n4288 GND.n4287 25.6005
R29077 GND.n4288 GND.n4282 25.6005
R29078 GND.n4294 GND.n4282 25.6005
R29079 GND.n4295 GND.n4294 25.6005
R29080 GND.n4296 GND.n4295 25.6005
R29081 GND.n4296 GND.n4280 25.6005
R29082 GND.n4302 GND.n4280 25.6005
R29083 GND.n4303 GND.n4302 25.6005
R29084 GND.n4304 GND.n4303 25.6005
R29085 GND.n4304 GND.n4278 25.6005
R29086 GND.n4309 GND.n4278 25.6005
R29087 GND.n4310 GND.n4309 25.6005
R29088 GND.n4310 GND.n4276 25.6005
R29089 GND.n4315 GND.n4276 25.6005
R29090 GND.n8351 GND.n8350 25.6005
R29091 GND.n8350 GND.n8349 25.6005
R29092 GND.n8349 GND.n1842 25.6005
R29093 GND.n1859 GND.n1842 25.6005
R29094 GND.n8337 GND.n1859 25.6005
R29095 GND.n8337 GND.n8336 25.6005
R29096 GND.n8336 GND.n8335 25.6005
R29097 GND.n8335 GND.n1860 25.6005
R29098 GND.n4336 GND.n1860 25.6005
R29099 GND.n4344 GND.n4336 25.6005
R29100 GND.n4344 GND.n4343 25.6005
R29101 GND.n4716 GND.n4207 25.6005
R29102 GND.n4716 GND.n4208 25.6005
R29103 GND.n2077 GND.n2031 25.6005
R29104 GND.n2078 GND.n2077 25.6005
R29105 GND.n8126 GND.n2078 25.6005
R29106 GND.n8126 GND.n8125 25.6005
R29107 GND.n8125 GND.n8124 25.6005
R29108 GND.n8124 GND.n2079 25.6005
R29109 GND.n2096 GND.n2079 25.6005
R29110 GND.n8112 GND.n2096 25.6005
R29111 GND.n8112 GND.n8111 25.6005
R29112 GND.n8111 GND.n8110 25.6005
R29113 GND.n8110 GND.n2097 25.6005
R29114 GND.n4571 GND.n4567 25.6005
R29115 GND.n4572 GND.n4571 25.6005
R29116 GND.n4573 GND.n4572 25.6005
R29117 GND.n4573 GND.n4565 25.6005
R29118 GND.n4579 GND.n4565 25.6005
R29119 GND.n4580 GND.n4579 25.6005
R29120 GND.n4581 GND.n4580 25.6005
R29121 GND.n4581 GND.n4563 25.6005
R29122 GND.n4587 GND.n4563 25.6005
R29123 GND.n4588 GND.n4587 25.6005
R29124 GND.n4589 GND.n4588 25.6005
R29125 GND.n4589 GND.n4561 25.6005
R29126 GND.n4595 GND.n4561 25.6005
R29127 GND.n4596 GND.n4595 25.6005
R29128 GND.n4597 GND.n4596 25.6005
R29129 GND.n4597 GND.n4559 25.6005
R29130 GND.n4319 GND.n4316 25.6005
R29131 GND.n4320 GND.n4319 25.6005
R29132 GND.n4321 GND.n4320 25.6005
R29133 GND.n4324 GND.n4321 25.6005
R29134 GND.n4325 GND.n4324 25.6005
R29135 GND.n4328 GND.n4325 25.6005
R29136 GND.n4329 GND.n4328 25.6005
R29137 GND.n4330 GND.n4329 25.6005
R29138 GND.n4331 GND.n4330 25.6005
R29139 GND.n4331 GND.n4274 25.6005
R29140 GND.n4349 GND.n4274 25.6005
R29141 GND.n4775 GND.n4191 25.6005
R29142 GND.n4775 GND.n4774 25.6005
R29143 GND.n4621 GND.n4558 25.6005
R29144 GND.n4617 GND.n4558 25.6005
R29145 GND.n4617 GND.n4616 25.6005
R29146 GND.n4616 GND.n4615 25.6005
R29147 GND.n4615 GND.n4612 25.6005
R29148 GND.n4612 GND.n4611 25.6005
R29149 GND.n4611 GND.n4608 25.6005
R29150 GND.n4608 GND.n4607 25.6005
R29151 GND.n4607 GND.n4606 25.6005
R29152 GND.n4606 GND.n4603 25.6005
R29153 GND.n4603 GND.n4602 25.6005
R29154 GND.n8394 GND.n8393 25.6005
R29155 GND.n8393 GND.n8392 25.6005
R29156 GND.n8392 GND.n8389 25.6005
R29157 GND.n8389 GND.n8388 25.6005
R29158 GND.n8388 GND.n8385 25.6005
R29159 GND.n8385 GND.n8384 25.6005
R29160 GND.n8384 GND.n8381 25.6005
R29161 GND.n8381 GND.n8380 25.6005
R29162 GND.n8380 GND.n8377 25.6005
R29163 GND.n8377 GND.n8376 25.6005
R29164 GND.n8376 GND.n8373 25.6005
R29165 GND.n8373 GND.n8372 25.6005
R29166 GND.n8372 GND.n8369 25.6005
R29167 GND.n8369 GND.n8368 25.6005
R29168 GND.n8368 GND.n8365 25.6005
R29169 GND.n8365 GND.n8364 25.6005
R29170 GND.n8358 GND.n1827 25.6005
R29171 GND.n8358 GND.n8357 25.6005
R29172 GND.n8357 GND.n8356 25.6005
R29173 GND.n8356 GND.n1832 25.6005
R29174 GND.n1850 GND.n1832 25.6005
R29175 GND.n8344 GND.n1850 25.6005
R29176 GND.n8344 GND.n8343 25.6005
R29177 GND.n8343 GND.n8342 25.6005
R29178 GND.n8342 GND.n1851 25.6005
R29179 GND.n1868 GND.n1851 25.6005
R29180 GND.n8330 GND.n1868 25.6005
R29181 GND.n8330 GND.n8329 25.6005
R29182 GND.n8329 GND.n8328 25.6005
R29183 GND.n4544 GND.n4542 25.6005
R29184 GND.n8132 GND.n8131 25.6005
R29185 GND.n8131 GND.n2068 25.6005
R29186 GND.n2087 GND.n2068 25.6005
R29187 GND.n8119 GND.n2087 25.6005
R29188 GND.n8119 GND.n8118 25.6005
R29189 GND.n8118 GND.n8117 25.6005
R29190 GND.n8117 GND.n2088 25.6005
R29191 GND.n2105 GND.n2088 25.6005
R29192 GND.n8105 GND.n2105 25.6005
R29193 GND.n8105 GND.n8104 25.6005
R29194 GND.n8104 GND.n8103 25.6005
R29195 GND.n8103 GND.n2106 25.6005
R29196 GND.n8097 GND.n2106 25.6005
R29197 GND.n8096 GND.n8095 25.6005
R29198 GND.n8095 GND.n8034 25.6005
R29199 GND.n8090 GND.n8034 25.6005
R29200 GND.n8090 GND.n8089 25.6005
R29201 GND.n8089 GND.n8036 25.6005
R29202 GND.n8084 GND.n8036 25.6005
R29203 GND.n8084 GND.n8083 25.6005
R29204 GND.n8083 GND.n8082 25.6005
R29205 GND.n8082 GND.n8038 25.6005
R29206 GND.n8076 GND.n8038 25.6005
R29207 GND.n8076 GND.n8075 25.6005
R29208 GND.n8075 GND.n8074 25.6005
R29209 GND.n8074 GND.n8040 25.6005
R29210 GND.n8068 GND.n8040 25.6005
R29211 GND.n8068 GND.n8067 25.6005
R29212 GND.n8067 GND.n8066 25.6005
R29213 GND.n1830 GND.n1828 25.6005
R29214 GND.n1874 GND.n1830 25.6005
R29215 GND.n1875 GND.n1874 25.6005
R29216 GND.n1876 GND.n1875 25.6005
R29217 GND.n1879 GND.n1876 25.6005
R29218 GND.n1880 GND.n1879 25.6005
R29219 GND.n1883 GND.n1880 25.6005
R29220 GND.n1884 GND.n1883 25.6005
R29221 GND.n1885 GND.n1884 25.6005
R29222 GND.n1888 GND.n1885 25.6005
R29223 GND.n1889 GND.n1888 25.6005
R29224 GND.n1890 GND.n1889 25.6005
R29225 GND.n8324 GND.n1890 25.6005
R29226 GND.n4534 GND.n4229 25.6005
R29227 GND.n8043 GND.n8042 25.6005
R29228 GND.n8044 GND.n8043 25.6005
R29229 GND.n8047 GND.n8044 25.6005
R29230 GND.n8048 GND.n8047 25.6005
R29231 GND.n8051 GND.n8048 25.6005
R29232 GND.n8052 GND.n8051 25.6005
R29233 GND.n8053 GND.n8052 25.6005
R29234 GND.n8056 GND.n8053 25.6005
R29235 GND.n8057 GND.n8056 25.6005
R29236 GND.n8060 GND.n8057 25.6005
R29237 GND.n8061 GND.n8060 25.6005
R29238 GND.n8062 GND.n8061 25.6005
R29239 GND.n8063 GND.n8062 25.6005
R29240 GND.n7072 GND.n6679 25.6005
R29241 GND.n7110 GND.n7072 25.6005
R29242 GND.n7110 GND.n7109 25.6005
R29243 GND.n7109 GND.n7108 25.6005
R29244 GND.n7108 GND.n7105 25.6005
R29245 GND.n7105 GND.n7104 25.6005
R29246 GND.n7104 GND.n7101 25.6005
R29247 GND.n7101 GND.n7100 25.6005
R29248 GND.n7100 GND.n7097 25.6005
R29249 GND.n7097 GND.n7096 25.6005
R29250 GND.n7096 GND.n7093 25.6005
R29251 GND.n7093 GND.n7092 25.6005
R29252 GND.n7092 GND.n7089 25.6005
R29253 GND.n7089 GND.n7088 25.6005
R29254 GND.n7088 GND.n7085 25.6005
R29255 GND.n7085 GND.n7084 25.6005
R29256 GND.n7138 GND.n7137 25.6005
R29257 GND.n7137 GND.n7136 25.6005
R29258 GND.n7136 GND.n6682 25.6005
R29259 GND.n7226 GND.n2553 25.6005
R29260 GND.n7311 GND.n2553 25.6005
R29261 GND.n7372 GND.n7371 25.6005
R29262 GND.n7371 GND.n7370 25.6005
R29263 GND.n7370 GND.n2523 25.6005
R29264 GND.n2580 GND.n2576 25.6005
R29265 GND.n2581 GND.n2580 25.6005
R29266 GND.n2582 GND.n2581 25.6005
R29267 GND.n2582 GND.n2574 25.6005
R29268 GND.n2588 GND.n2574 25.6005
R29269 GND.n2589 GND.n2588 25.6005
R29270 GND.n2590 GND.n2589 25.6005
R29271 GND.n2590 GND.n2572 25.6005
R29272 GND.n2596 GND.n2572 25.6005
R29273 GND.n2597 GND.n2596 25.6005
R29274 GND.n2598 GND.n2597 25.6005
R29275 GND.n2598 GND.n2570 25.6005
R29276 GND.n2604 GND.n2570 25.6005
R29277 GND.n2605 GND.n2604 25.6005
R29278 GND.n2606 GND.n2605 25.6005
R29279 GND.n2606 GND.n2568 25.6005
R29280 GND.n7082 GND.n7081 25.6005
R29281 GND.n7081 GND.n7080 25.6005
R29282 GND.n7080 GND.n7078 25.6005
R29283 GND.n7209 GND.n7206 25.6005
R29284 GND.n7209 GND.n7207 25.6005
R29285 GND.n2615 GND.n2614 25.6005
R29286 GND.n2614 GND.n2612 25.6005
R29287 GND.n2612 GND.n2611 25.6005
R29288 GND.n6704 GND.n6702 25.6005
R29289 GND.n6705 GND.n6704 25.6005
R29290 GND.n6708 GND.n6705 25.6005
R29291 GND.n6709 GND.n6708 25.6005
R29292 GND.n6712 GND.n6709 25.6005
R29293 GND.n6713 GND.n6712 25.6005
R29294 GND.n6716 GND.n6713 25.6005
R29295 GND.n6717 GND.n6716 25.6005
R29296 GND.n6720 GND.n6717 25.6005
R29297 GND.n6721 GND.n6720 25.6005
R29298 GND.n6724 GND.n6721 25.6005
R29299 GND.n6726 GND.n6724 25.6005
R29300 GND.n6727 GND.n6726 25.6005
R29301 GND.n6728 GND.n6727 25.6005
R29302 GND.n6728 GND.n6691 25.6005
R29303 GND.n7116 GND.n6691 25.6005
R29304 GND.n7127 GND.n6687 25.6005
R29305 GND.n7128 GND.n7127 25.6005
R29306 GND.n7131 GND.n7128 25.6005
R29307 GND.n7211 GND.n2561 25.6005
R29308 GND.n7307 GND.n2561 25.6005
R29309 GND.n7292 GND.n2530 25.6005
R29310 GND.n7366 GND.n2530 25.6005
R29311 GND.n7366 GND.n7365 25.6005
R29312 GND.n7364 GND.n2531 25.6005
R29313 GND.n7359 GND.n2531 25.6005
R29314 GND.n7359 GND.n7358 25.6005
R29315 GND.n7358 GND.n2533 25.6005
R29316 GND.n7353 GND.n2533 25.6005
R29317 GND.n7353 GND.n7352 25.6005
R29318 GND.n7352 GND.n7351 25.6005
R29319 GND.n7351 GND.n2535 25.6005
R29320 GND.n7345 GND.n2535 25.6005
R29321 GND.n7345 GND.n7344 25.6005
R29322 GND.n7344 GND.n7343 25.6005
R29323 GND.n7343 GND.n2537 25.6005
R29324 GND.n7337 GND.n2537 25.6005
R29325 GND.n7337 GND.n7336 25.6005
R29326 GND.n7336 GND.n7335 25.6005
R29327 GND.n7335 GND.n2539 25.6005
R29328 GND.n7123 GND.n7117 25.6005
R29329 GND.n7123 GND.n7122 25.6005
R29330 GND.n7122 GND.n7121 25.6005
R29331 GND.n7231 GND.n2695 25.6005
R29332 GND.n7232 GND.n7231 25.6005
R29333 GND.n7328 GND.n7326 25.6005
R29334 GND.n7329 GND.n7328 25.6005
R29335 GND.n7330 GND.n7329 25.6005
R29336 GND.n6872 GND.n6788 25.6005
R29337 GND.n6901 GND.n6872 25.6005
R29338 GND.n6901 GND.n6900 25.6005
R29339 GND.n6900 GND.n6899 25.6005
R29340 GND.n6899 GND.n6896 25.6005
R29341 GND.n6896 GND.n6895 25.6005
R29342 GND.n6895 GND.n6892 25.6005
R29343 GND.n6892 GND.n6891 25.6005
R29344 GND.n6891 GND.n6888 25.6005
R29345 GND.n6888 GND.n6887 25.6005
R29346 GND.n6887 GND.n6884 25.6005
R29347 GND.n6884 GND.n6883 25.6005
R29348 GND.n6883 GND.n6880 25.6005
R29349 GND.n6880 GND.n6879 25.6005
R29350 GND.n6879 GND.n6876 25.6005
R29351 GND.n6876 GND.n6875 25.6005
R29352 GND.n6916 GND.n6915 25.6005
R29353 GND.n6918 GND.n6916 25.6005
R29354 GND.n6918 GND.n6917 25.6005
R29355 GND.n6917 GND.n6771 25.6005
R29356 GND.n6965 GND.n6771 25.6005
R29357 GND.n6966 GND.n6965 25.6005
R29358 GND.n6968 GND.n6966 25.6005
R29359 GND.n6968 GND.n6967 25.6005
R29360 GND.n6967 GND.n6753 25.6005
R29361 GND.n7001 GND.n6753 25.6005
R29362 GND.n7002 GND.n7001 25.6005
R29363 GND.n7189 GND.n6638 25.6005
R29364 GND.n7189 GND.n7188 25.6005
R29365 GND.n7426 GND.n2423 25.6005
R29366 GND.n7578 GND.n2423 25.6005
R29367 GND.n7578 GND.n7577 25.6005
R29368 GND.n7577 GND.n7576 25.6005
R29369 GND.n7576 GND.n2424 25.6005
R29370 GND.n2441 GND.n2424 25.6005
R29371 GND.n7564 GND.n2441 25.6005
R29372 GND.n7564 GND.n7563 25.6005
R29373 GND.n7563 GND.n7562 25.6005
R29374 GND.n7562 GND.n2442 25.6005
R29375 GND.n2465 GND.n2442 25.6005
R29376 GND.n7549 GND.n7548 25.6005
R29377 GND.n7548 GND.n7547 25.6005
R29378 GND.n7547 GND.n7546 25.6005
R29379 GND.n7546 GND.n7544 25.6005
R29380 GND.n7544 GND.n7541 25.6005
R29381 GND.n7541 GND.n7540 25.6005
R29382 GND.n7540 GND.n7537 25.6005
R29383 GND.n7537 GND.n7536 25.6005
R29384 GND.n7536 GND.n7533 25.6005
R29385 GND.n7533 GND.n7532 25.6005
R29386 GND.n7532 GND.n7529 25.6005
R29387 GND.n7529 GND.n7528 25.6005
R29388 GND.n7528 GND.n7525 25.6005
R29389 GND.n7525 GND.n7524 25.6005
R29390 GND.n7524 GND.n7521 25.6005
R29391 GND.n7521 GND.n7520 25.6005
R29392 GND.n6873 GND.n6783 25.6005
R29393 GND.n6922 GND.n6783 25.6005
R29394 GND.n6923 GND.n6922 25.6005
R29395 GND.n6952 GND.n6923 25.6005
R29396 GND.n6952 GND.n6951 25.6005
R29397 GND.n6951 GND.n6950 25.6005
R29398 GND.n6950 GND.n6947 25.6005
R29399 GND.n6947 GND.n6946 25.6005
R29400 GND.n6946 GND.n6944 25.6005
R29401 GND.n6944 GND.n6943 25.6005
R29402 GND.n6943 GND.n6942 25.6005
R29403 GND.n7194 GND.n6635 25.6005
R29404 GND.n6635 GND.n2637 25.6005
R29405 GND.n2660 GND.n2659 25.6005
R29406 GND.n2659 GND.n2656 25.6005
R29407 GND.n2656 GND.n2655 25.6005
R29408 GND.n2655 GND.n2652 25.6005
R29409 GND.n2652 GND.n2651 25.6005
R29410 GND.n2651 GND.n2648 25.6005
R29411 GND.n2648 GND.n2467 25.6005
R29412 GND.n7514 GND.n2467 25.6005
R29413 GND.n7515 GND.n7514 25.6005
R29414 GND.n7516 GND.n7515 25.6005
R29415 GND.n7516 GND.n2466 25.6005
R29416 GND.n6843 GND.n6842 25.6005
R29417 GND.n6842 GND.n6805 25.6005
R29418 GND.n6836 GND.n6805 25.6005
R29419 GND.n6836 GND.n6835 25.6005
R29420 GND.n6835 GND.n6834 25.6005
R29421 GND.n6834 GND.n6807 25.6005
R29422 GND.n6828 GND.n6807 25.6005
R29423 GND.n6828 GND.n6827 25.6005
R29424 GND.n6827 GND.n6826 25.6005
R29425 GND.n6826 GND.n6809 25.6005
R29426 GND.n6820 GND.n6809 25.6005
R29427 GND.n6820 GND.n6819 25.6005
R29428 GND.n6819 GND.n6818 25.6005
R29429 GND.n6818 GND.n6811 25.6005
R29430 GND.n6812 GND.n6811 25.6005
R29431 GND.n6812 GND.n6800 25.6005
R29432 GND.n6844 GND.n6796 25.6005
R29433 GND.n6907 GND.n6796 25.6005
R29434 GND.n6908 GND.n6907 25.6005
R29435 GND.n6910 GND.n6908 25.6005
R29436 GND.n6910 GND.n6909 25.6005
R29437 GND.n6909 GND.n6778 25.6005
R29438 GND.n6957 GND.n6778 25.6005
R29439 GND.n6958 GND.n6957 25.6005
R29440 GND.n6960 GND.n6958 25.6005
R29441 GND.n6960 GND.n6959 25.6005
R29442 GND.n6959 GND.n6760 25.6005
R29443 GND.n6987 GND.n6760 25.6005
R29444 GND.n6988 GND.n6987 25.6005
R29445 GND.n7251 GND.n2633 25.6005
R29446 GND.n7436 GND.n7435 25.6005
R29447 GND.n7435 GND.n2432 25.6005
R29448 GND.n7571 GND.n2432 25.6005
R29449 GND.n7571 GND.n7570 25.6005
R29450 GND.n7570 GND.n7569 25.6005
R29451 GND.n7569 GND.n2433 25.6005
R29452 GND.n2449 GND.n2433 25.6005
R29453 GND.n7557 GND.n2449 25.6005
R29454 GND.n7557 GND.n7556 25.6005
R29455 GND.n7556 GND.n7555 25.6005
R29456 GND.n7555 GND.n2450 25.6005
R29457 GND.n7498 GND.n2450 25.6005
R29458 GND.n7498 GND.n7497 25.6005
R29459 GND.n7496 GND.n7453 25.6005
R29460 GND.n7491 GND.n7453 25.6005
R29461 GND.n7491 GND.n7490 25.6005
R29462 GND.n7490 GND.n7489 25.6005
R29463 GND.n7489 GND.n7486 25.6005
R29464 GND.n7486 GND.n7485 25.6005
R29465 GND.n7485 GND.n7482 25.6005
R29466 GND.n7482 GND.n7481 25.6005
R29467 GND.n7481 GND.n7478 25.6005
R29468 GND.n7478 GND.n7477 25.6005
R29469 GND.n7477 GND.n7474 25.6005
R29470 GND.n7474 GND.n7473 25.6005
R29471 GND.n7473 GND.n7470 25.6005
R29472 GND.n7470 GND.n7469 25.6005
R29473 GND.n7469 GND.n7466 25.6005
R29474 GND.n7466 GND.n7465 25.6005
R29475 GND.n6849 GND.n6848 25.6005
R29476 GND.n6861 GND.n6849 25.6005
R29477 GND.n6861 GND.n6860 25.6005
R29478 GND.n6860 GND.n6859 25.6005
R29479 GND.n6859 GND.n6858 25.6005
R29480 GND.n6858 GND.n6854 25.6005
R29481 GND.n6854 GND.n6853 25.6005
R29482 GND.n6853 GND.n6852 25.6005
R29483 GND.n6852 GND.n6850 25.6005
R29484 GND.n6850 GND.n6765 25.6005
R29485 GND.n6973 GND.n6765 25.6005
R29486 GND.n6974 GND.n6973 25.6005
R29487 GND.n6980 GND.n6974 25.6005
R29488 GND.n7255 GND.n2630 25.6005
R29489 GND.n2471 GND.n2469 25.6005
R29490 GND.n7442 GND.n2469 25.6005
R29491 GND.n7443 GND.n7442 25.6005
R29492 GND.n7446 GND.n7443 25.6005
R29493 GND.n7447 GND.n7446 25.6005
R29494 GND.n7448 GND.n7447 25.6005
R29495 GND.n7509 GND.n7448 25.6005
R29496 GND.n7509 GND.n7508 25.6005
R29497 GND.n7508 GND.n7507 25.6005
R29498 GND.n7507 GND.n7504 25.6005
R29499 GND.n7504 GND.n7503 25.6005
R29500 GND.n7503 GND.n7449 25.6005
R29501 GND.n7463 GND.n7449 25.6005
R29502 GND.n5510 GND.n5509 25.4876
R29503 GND.n7628 GND.n2354 25.4876
R29504 GND.n9520 GND.n9519 25.4876
R29505 GND.n9752 GND.n72 25.4876
R29506 GND.n7885 GND.n2205 25.4876
R29507 GND.n7871 GND.n2154 25.4876
R29508 GND.n5550 GND.n5530 25.384
R29509 GND.n9549 GND.n9548 25.384
R29510 GND.n7827 GND.n7826 25.384
R29511 GND.n5653 GND.n5459 25.3181
R29512 GND.n9575 GND.n9574 25.3181
R29513 GND.n7848 GND.n7847 25.3181
R29514 GND.n5134 GND.n5133 25.224
R29515 GND.n5133 GND.n5132 25.224
R29516 GND.n1213 GND.n1212 25.224
R29517 GND.n1213 GND.n1140 25.224
R29518 GND.n3259 GND.n3258 25.224
R29519 GND.n3259 GND.n3186 25.224
R29520 GND.n5466 GND.n5465 25.1487
R29521 GND.n5520 GND.n5490 25.1487
R29522 GND.n9719 GND.n9716 25.1487
R29523 GND.n9594 GND.n137 25.1487
R29524 GND.n7940 GND.n7937 25.1487
R29525 GND.n2250 GND.n2248 25.1487
R29526 GND.n3096 GND.t390 24.9236
R29527 GND.n3096 GND.t396 24.9236
R29528 GND.n2919 GND.t103 24.9236
R29529 GND.n2919 GND.t64 24.9236
R29530 GND.n3039 GND.t299 24.9236
R29531 GND.n3039 GND.t295 24.9236
R29532 GND.n2970 GND.t97 24.9236
R29533 GND.n2970 GND.t279 24.9236
R29534 GND.n2963 GND.t417 24.9236
R29535 GND.n2963 GND.t85 24.9236
R29536 GND.n2941 GND.t136 24.9236
R29537 GND.n2941 GND.t132 24.9236
R29538 GND.n2933 GND.t130 24.9236
R29539 GND.n2933 GND.t134 24.9236
R29540 GND.n2924 GND.t91 24.9236
R29541 GND.n2924 GND.t93 24.9236
R29542 GND.n2960 GND.t95 24.9236
R29543 GND.n2960 GND.t89 24.9236
R29544 GND.n2923 GND.t147 24.9236
R29545 GND.n2923 GND.t140 24.9236
R29546 GND.n2916 GND.t138 24.9236
R29547 GND.n2916 GND.t143 24.9236
R29548 GND.n3014 GND.t113 24.9236
R29549 GND.n3014 GND.t273 24.9236
R29550 GND.n2912 GND.t111 24.9236
R29551 GND.n2912 GND.t200 24.9236
R29552 GND.n2905 GND.t293 24.9236
R29553 GND.n2905 GND.t297 24.9236
R29554 GND.n3045 GND.t333 24.9236
R29555 GND.n3045 GND.t9 24.9236
R29556 GND.n3047 GND.t38 24.9236
R29557 GND.n3047 GND.t345 24.9236
R29558 GND.n3089 GND.t382 24.9236
R29559 GND.n3089 GND.t392 24.9236
R29560 GND.n2903 GND.t388 24.9236
R29561 GND.n2903 GND.t394 24.9236
R29562 GND.n6341 GND.n6334 24.8551
R29563 GND.n8522 GND.n8521 24.8551
R29564 GND.n3946 GND.n3945 24.8551
R29565 GND.n8972 GND.n8971 24.8476
R29566 GND.n888 GND.n887 24.8476
R29567 GND.n895 GND.n874 24.8476
R29568 GND.n885 GND.n877 24.8476
R29569 GND.n4674 GND.n4224 24.8476
R29570 GND.n4546 GND.n4545 24.8476
R29571 GND.n4670 GND.n4669 24.8476
R29572 GND.n4665 GND.n4664 24.8476
R29573 GND.n7199 GND.n7198 24.8476
R29574 GND.n7250 GND.n2634 24.8476
R29575 GND.n7030 GND.n7029 24.8476
R29576 GND.n7257 GND.n7256 24.8476
R29577 GND.n5497 GND.n5496 24.584
R29578 GND.n5482 GND.n5469 24.584
R29579 GND.n146 GND.n145 24.584
R29580 GND.n9729 GND.n9728 24.584
R29581 GND.n2240 GND.n2237 24.584
R29582 GND.n7950 GND.n7949 24.584
R29583 GND.n7734 GND.n7733 24.5614
R29584 GND.n9802 GND.n9798 24.5614
R29585 GND.n8406 GND.n16 24.5614
R29586 GND.n9808 GND.n9807 24.5614
R29587 GND.n8398 GND.n8397 24.5614
R29588 GND.n7689 GND.n7688 24.5614
R29589 GND.n2847 GND.n2846 24.4711
R29590 GND.n6212 GND.n2847 24.4711
R29591 GND.n8671 GND.n1018 24.4711
R29592 GND.n8673 GND.n8671 24.4711
R29593 GND.n4045 GND.n4044 24.4711
R29594 GND.n4044 GND.n4015 24.4711
R29595 GND.n5018 GND.n5017 24.3581
R29596 GND.n1450 GND.n1448 24.3581
R29597 GND.n3497 GND.n3495 24.3581
R29598 GND.t225 GND.t213 24.2386
R29599 GND.t72 GND.t425 24.2386
R29600 GND.n2962 GND.n2959 24.0946
R29601 GND.n3101 GND.n2895 24.0946
R29602 GND.n9384 GND.n251 24.0946
R29603 GND.n9372 GND.n271 24.0946
R29604 GND.n958 GND.n472 24.0946
R29605 GND.n965 GND.n963 24.0946
R29606 GND.n262 GND.n261 24.0946
R29607 GND.n280 GND.n264 24.0946
R29608 GND.n8978 GND.n8977 24.0946
R29609 GND.n9022 GND.n9021 24.0946
R29610 GND.n841 GND.n828 24.0946
R29611 GND.n9049 GND.n444 24.0946
R29612 GND.n939 GND.n485 24.0946
R29613 GND.n9037 GND.n9036 24.0946
R29614 GND.n8278 GND.n1943 24.0946
R29615 GND.n8266 GND.n1963 24.0946
R29616 GND.n4692 GND.n4211 24.0946
R29617 GND.n4710 GND.n4695 24.0946
R29618 GND.n1954 GND.n1953 24.0946
R29619 GND.n1972 GND.n1956 24.0946
R29620 GND.n4494 GND.n4257 24.0946
R29621 GND.n4725 GND.n4723 24.0946
R29622 GND.n4488 GND.n4487 24.0946
R29623 GND.n4769 GND.n4199 24.0946
R29624 GND.n4468 GND.n4467 24.0946
R29625 GND.n4195 GND.n4193 24.0946
R29626 GND.n7225 GND.n6614 24.0946
R29627 GND.n7313 GND.n7312 24.0946
R29628 GND.n7205 GND.n7204 24.0946
R29629 GND.n2567 GND.n2564 24.0946
R29630 GND.n7212 GND.n6625 24.0946
R29631 GND.n7306 GND.n2562 24.0946
R29632 GND.n7185 GND.n7184 24.0946
R29633 GND.n7234 GND.n7233 24.0946
R29634 GND.n7178 GND.n6644 24.0946
R29635 GND.n7242 GND.n2692 24.0946
R29636 GND.n7195 GND.n6634 24.0946
R29637 GND.n7247 GND.n7246 24.0946
R29638 GND.n5560 GND.n5449 23.8499
R29639 GND.n9707 GND.n104 23.8499
R29640 GND.n7928 GND.n2187 23.8499
R29641 GND.n3092 GND.n2895 23.7181
R29642 GND.n7609 GND.n2384 23.6805
R29643 GND.n5563 GND.n5446 23.6805
R29644 GND.n111 GND.n70 23.6805
R29645 GND.n9632 GND.n9631 23.6805
R29646 GND.n7914 GND.n7913 23.6805
R29647 GND.n7892 GND.n7891 23.6805
R29648 GND.n735 GND.n197 23.6071
R29649 GND.n9425 GND.n9424 23.6071
R29650 GND.n858 GND.n200 23.6071
R29651 GND.n9414 GND.n211 23.6071
R29652 GND.n9300 GND.n317 23.6071
R29653 GND.n9299 GND.n335 23.6071
R29654 GND.n9243 GND.n371 23.6071
R29655 GND.n4346 GND.n4333 23.6071
R29656 GND.n8318 GND.n1895 23.6071
R29657 GND.n4270 GND.n1896 23.6071
R29658 GND.n8308 GND.n1907 23.6071
R29659 GND.n8194 GND.n2009 23.6071
R29660 GND.n8193 GND.n2027 23.6071
R29661 GND.n8137 GND.n2063 23.6071
R29662 GND.n6999 GND.n6998 23.6071
R29663 GND.n6757 GND.n6749 23.6071
R29664 GND.n7013 GND.n7012 23.6071
R29665 GND.n6934 GND.n6671 23.6071
R29666 GND.n7420 GND.n7419 23.6071
R29667 GND.n7429 GND.n2478 23.6071
R29668 GND.n7428 GND.n2481 23.6071
R29669 GND.n480 GND.n468 23.3417
R29670 GND.n9043 GND.n451 23.3417
R29671 GND.n900 GND.n898 23.3417
R29672 GND.n884 GND.n878 23.3417
R29673 GND.n4675 GND.n4220 23.3417
R29674 GND.n4659 GND.n4547 23.3417
R29675 GND.n4529 GND.n4228 23.3417
R29676 GND.n4540 GND.n4535 23.3417
R29677 GND.n6655 GND.n6632 23.3417
R29678 GND.n7279 GND.n2623 23.3417
R29679 GND.n7035 GND.n7033 23.3417
R29680 GND.n7275 GND.n2627 23.3417
R29681 GND.n5532 GND.n5529 23.2193
R29682 GND.n9542 GND.n173 23.2193
R29683 GND.n7819 GND.n2260 23.2193
R29684 GND.n5625 GND.n5555 23.0238
R29685 GND.n5618 GND.n5554 23.0238
R29686 GND.n9610 GND.n9609 23.0238
R29687 GND.n9691 GND.n127 23.0238
R29688 GND.n2196 GND.n2146 23.0238
R29689 GND.n7982 GND.n7981 23.0238
R29690 GND.n2992 GND.n2959 22.5887
R29691 GND.n3032 GND.n2909 22.5887
R29692 GND.n9388 GND.n9387 22.5887
R29693 GND.n9369 GND.n9368 22.5887
R29694 GND.n954 GND.n953 22.5887
R29695 GND.n974 GND.n973 22.5887
R29696 GND.n9392 GND.n242 22.5887
R29697 GND.n9364 GND.n281 22.5887
R29698 GND.n846 GND.n462 22.5887
R29699 GND.n9020 GND.n9019 22.5887
R29700 GND.n842 GND.n827 22.5887
R29701 GND.n9051 GND.n9050 22.5887
R29702 GND.n940 GND.n483 22.5887
R29703 GND.n9035 GND.n9034 22.5887
R29704 GND.n8282 GND.n8281 22.5887
R29705 GND.n8263 GND.n8262 22.5887
R29706 GND.n4688 GND.n4687 22.5887
R29707 GND.n4706 GND.n4705 22.5887
R29708 GND.n8286 GND.n1934 22.5887
R29709 GND.n8258 GND.n1973 22.5887
R29710 GND.n4496 GND.n4495 22.5887
R29711 GND.n4764 GND.n4763 22.5887
R29712 GND.n4481 GND.n4471 22.5887
R29713 GND.n4768 GND.n4200 22.5887
R29714 GND.n4466 GND.n4465 22.5887
R29715 GND.n4652 GND.n4651 22.5887
R29716 GND.n7222 GND.n7221 22.5887
R29717 GND.n7318 GND.n2550 22.5887
R29718 GND.n7074 GND.n6628 22.5887
R29719 GND.n7302 GND.n7301 22.5887
R29720 GND.n7217 GND.n7216 22.5887
R29721 GND.n7290 GND.n7289 22.5887
R29722 GND.n7183 GND.n6640 22.5887
R29723 GND.n7322 GND.n2542 22.5887
R29724 GND.n7179 GND.n6643 22.5887
R29725 GND.n7241 GND.n2693 22.5887
R29726 GND.n7165 GND.n7164 22.5887
R29727 GND.n2686 GND.n2638 22.5887
R29728 GND.t3 GND.n8431 22.5377
R29729 GND.n3009 GND.n2915 22.2123
R29730 GND.n3098 GND.n3095 22.2123
R29731 GND.n6356 GND.n6324 21.8734
R29732 GND.n8535 GND.n8534 21.8734
R29733 GND.n4951 GND.n4950 21.8734
R29734 GND.n946 GND.n945 21.8358
R29735 GND.n9042 GND.n452 21.8358
R29736 GND.n902 GND.n901 21.8358
R29737 GND.n881 GND.n880 21.8358
R29738 GND.n4680 GND.n4679 21.8358
R29739 GND.n4658 GND.n4548 21.8358
R29740 GND.n4530 GND.n4528 21.8358
R29741 GND.n4539 GND.n4537 21.8358
R29742 GND.n7170 GND.n7169 21.8358
R29743 GND.n7281 GND.n7280 21.8358
R29744 GND.n7037 GND.n7036 21.8358
R29745 GND.n7274 GND.n2628 21.8358
R29746 GND.n7683 GND.n2316 21.8132
R29747 GND.n324 GND.t231 21.6398
R29748 GND.n2016 GND.t33 21.6398
R29749 GND.t116 GND.n2496 21.6398
R29750 GND.n5434 GND.n5431 21.3765
R29751 GND.n1466 GND.n1465 21.3765
R29752 GND.n3509 GND.n3508 21.3765
R29753 GND.n3032 GND.n3031 21.0829
R29754 GND.n3108 GND.n2893 21.0829
R29755 GND.n250 GND.n249 21.0829
R29756 GND.n291 GND.n273 21.0829
R29757 GND.n952 GND.n951 21.0829
R29758 GND.n972 GND.n971 21.0829
R29759 GND.n9393 GND.n240 21.0829
R29760 GND.n9363 GND.n282 21.0829
R29761 GND.n847 GND.n824 21.0829
R29762 GND.n9018 GND.n8982 21.0829
R29763 GND.n837 GND.n836 21.0829
R29764 GND.n9057 GND.n440 21.0829
R29765 GND.n935 GND.n934 21.0829
R29766 GND.n9061 GND.n436 21.0829
R29767 GND.n1942 GND.n1941 21.0829
R29768 GND.n1983 GND.n1965 21.0829
R29769 GND.n4686 GND.n4685 21.0829
R29770 GND.n4704 GND.n4703 21.0829
R29771 GND.n8287 GND.n1932 21.0829
R29772 GND.n8257 GND.n1974 21.0829
R29773 GND.n4497 GND.n4255 21.0829
R29774 GND.n4762 GND.n4761 21.0829
R29775 GND.n4482 GND.n4480 21.0829
R29776 GND.n4645 GND.n4641 21.0829
R29777 GND.n4464 GND.n4260 21.0829
R29778 GND.n4650 GND.n4649 21.0829
R29779 GND.n6680 GND.n6616 21.0829
R29780 GND.n7317 GND.n2551 21.0829
R29781 GND.n7075 GND.n7073 21.0829
R29782 GND.n7300 GND.n7299 21.0829
R29783 GND.n7129 GND.n6624 21.0829
R29784 GND.n7295 GND.n7291 21.0829
R29785 GND.n7119 GND.n7118 21.0829
R29786 GND.n7323 GND.n2540 21.0829
R29787 GND.n6647 GND.n6646 21.0829
R29788 GND.n7237 GND.n7236 21.0829
R29789 GND.n7162 GND.n7161 21.0829
R29790 GND.n2685 GND.n2641 21.0829
R29791 GND.n9425 GND.n197 20.9841
R29792 GND.n9424 GND.n200 20.9841
R29793 GND.n858 GND.n857 20.9841
R29794 GND.n752 GND.n211 20.9841
R29795 GND.n791 GND.n224 20.9841
R29796 GND.n9405 GND.n224 20.9841
R29797 GND.n927 GND.n490 20.9841
R29798 GND.n925 GND.n234 20.9841
R29799 GND.n494 GND.n475 20.9841
R29800 GND.n949 GND.n948 20.9841
R29801 GND.n948 GND.n244 20.9841
R29802 GND.n9390 GND.n247 20.9841
R29803 GND.n8974 GND.n256 20.9841
R29804 GND.n9381 GND.n259 20.9841
R29805 GND.n9030 GND.n259 20.9841
R29806 GND.n891 GND.t39 20.9841
R29807 GND.n891 GND.n266 20.9841
R29808 GND.n9375 GND.n269 20.9841
R29809 GND.n9045 GND.n275 20.9841
R29810 GND.n9366 GND.n278 20.9841
R29811 GND.n9059 GND.n278 20.9841
R29812 GND.n9268 GND.n358 20.9841
R29813 GND.n9358 GND.n289 20.9841
R29814 GND.n9280 GND.n9279 20.9841
R29815 GND.n9279 GND.n351 20.9841
R29816 GND.n9352 GND.n297 20.9841
R29817 GND.n321 GND.n297 20.9841
R29818 GND.n9310 GND.n9309 20.9841
R29819 GND.n9309 GND.n324 20.9841
R29820 GND.n9300 GND.n9299 20.9841
R29821 GND.n371 GND.n335 20.9841
R29822 GND.n9243 GND.n372 20.9841
R29823 GND.n4333 GND.n1895 20.9841
R29824 GND.n8318 GND.n1896 20.9841
R29825 GND.n4357 GND.n4270 20.9841
R29826 GND.n4449 GND.n1907 20.9841
R29827 GND.n4448 GND.n1916 20.9841
R29828 GND.n8299 GND.n1916 20.9841
R29829 GND.n4505 GND.n4504 20.9841
R29830 GND.n4522 GND.n1926 20.9841
R29831 GND.n4524 GND.n4214 20.9841
R29832 GND.n4683 GND.n4682 20.9841
R29833 GND.n4682 GND.n1936 20.9841
R29834 GND.n8284 GND.n1939 20.9841
R29835 GND.n4672 GND.n1948 20.9841
R29836 GND.n8275 GND.n1951 20.9841
R29837 GND.n4714 GND.n1951 20.9841
R29838 GND.t40 GND.n4210 20.9841
R29839 GND.n4210 GND.n1958 20.9841
R29840 GND.n8269 GND.n1961 20.9841
R29841 GND.n4661 GND.n1967 20.9841
R29842 GND.n8260 GND.n1970 20.9841
R29843 GND.n4647 GND.n1970 20.9841
R29844 GND.n8162 GND.n2050 20.9841
R29845 GND.n8252 GND.n1981 20.9841
R29846 GND.n8174 GND.n8173 20.9841
R29847 GND.n8173 GND.n2043 20.9841
R29848 GND.n8246 GND.n1989 20.9841
R29849 GND.n2013 GND.n1989 20.9841
R29850 GND.n8204 GND.n8203 20.9841
R29851 GND.n8203 GND.n2016 20.9841
R29852 GND.n8194 GND.n8193 20.9841
R29853 GND.n2063 GND.n2027 20.9841
R29854 GND.n8137 GND.n2064 20.9841
R29855 GND.n6998 GND.n6757 20.9841
R29856 GND.n7012 GND.n6749 20.9841
R29857 GND.n7013 GND.n6693 20.9841
R29858 GND.n7141 GND.n6671 20.9841
R29859 GND.n7140 GND.n6675 20.9841
R29860 GND.n6688 GND.n6675 20.9841
R29861 GND.n7154 GND.n6663 20.9841
R29862 GND.n7044 GND.n6683 20.9841
R29863 GND.n7174 GND.n6648 20.9841
R29864 GND.n7173 GND.n7172 20.9841
R29865 GND.n7172 GND.n6618 20.9841
R29866 GND.n7219 GND.n6621 20.9841
R29867 GND.n7201 GND.n6609 20.9841
R29868 GND.n7228 GND.n6611 20.9841
R29869 GND.n7191 GND.n6611 20.9841
R29870 GND.n7253 GND.t238 20.9841
R29871 GND.n7253 GND.n2555 20.9841
R29872 GND.n7309 GND.n2558 20.9841
R29873 GND.n7277 GND.n2545 20.9841
R29874 GND.n7320 GND.n2547 20.9841
R29875 GND.n2617 GND.n2547 20.9841
R29876 GND.n7297 GND.n7288 20.9841
R29877 GND.n7374 GND.n2518 20.9841
R29878 GND.n7390 GND.n2505 20.9841
R29879 GND.n7390 GND.n7389 20.9841
R29880 GND.n7368 GND.n2527 20.9841
R29881 GND.n2670 GND.n2527 20.9841
R29882 GND.n7404 GND.n2495 20.9841
R29883 GND.n7404 GND.n2496 20.9841
R29884 GND.n7419 GND.n2478 20.9841
R29885 GND.n7429 GND.n7428 20.9841
R29886 GND.n2657 GND.n2481 20.9841
R29887 GND.n6596 GND.n6592 20.3299
R29888 GND.n6582 GND.n6578 20.3299
R29889 GND.n6568 GND.n6564 20.3299
R29890 GND.n6554 GND.n6550 20.3299
R29891 GND.n6540 GND.n6536 20.3299
R29892 GND.n2706 GND.n2702 20.3299
R29893 GND.n6455 GND.n6451 20.3299
R29894 GND.n6469 GND.n6465 20.3299
R29895 GND.n6482 GND.n6478 20.3299
R29896 GND.n6495 GND.n6491 20.3299
R29897 GND.n6508 GND.n6504 20.3299
R29898 GND.n6521 GND.n6517 20.3299
R29899 GND.n6436 GND.n6432 20.3299
R29900 GND.n8959 GND.n8955 20.3299
R29901 GND.n8945 GND.n8941 20.3299
R29902 GND.n8931 GND.n8927 20.3299
R29903 GND.n8917 GND.n8913 20.3299
R29904 GND.n8903 GND.n8899 20.3299
R29905 GND.n989 GND.n985 20.3299
R29906 GND.n8819 GND.n8815 20.3299
R29907 GND.n8833 GND.n8829 20.3299
R29908 GND.n8846 GND.n8842 20.3299
R29909 GND.n8859 GND.n8855 20.3299
R29910 GND.n8872 GND.n8868 20.3299
R29911 GND.n8885 GND.n8881 20.3299
R29912 GND.n8800 GND.n8796 20.3299
R29913 GND.n911 GND.n479 20.3299
R29914 GND.n9270 GND.n356 20.3299
R29915 GND.n903 GND.n497 20.3299
R29916 GND.n9266 GND.n361 20.3299
R29917 GND.n4858 GND.n4854 20.3299
R29918 GND.n4844 GND.n4840 20.3299
R29919 GND.n4830 GND.n4826 20.3299
R29920 GND.n4816 GND.n4812 20.3299
R29921 GND.n4802 GND.n4798 20.3299
R29922 GND.n4787 GND.n4783 20.3299
R29923 GND.n4181 GND.n4177 20.3299
R29924 GND.n4875 GND.n4871 20.3299
R29925 GND.n4888 GND.n4884 20.3299
R29926 GND.n4901 GND.n4897 20.3299
R29927 GND.n4914 GND.n4910 20.3299
R29928 GND.n4927 GND.n4923 20.3299
R29929 GND.n4162 GND.n4158 20.3299
R29930 GND.n4508 GND.n4219 20.3299
R29931 GND.n8164 GND.n2048 20.3299
R29932 GND.n4527 GND.n4526 20.3299
R29933 GND.n8160 GND.n2053 20.3299
R29934 GND.n7047 GND.n6654 20.3299
R29935 GND.n7286 GND.n2620 20.3299
R29936 GND.n7038 GND.n6742 20.3299
R29937 GND.n7271 GND.n7270 20.3299
R29938 GND.t99 GND.n9414 20.3284
R29939 GND.t270 GND.n8308 20.3284
R29940 GND.n6934 GND.t421 20.3284
R29941 GND.n7582 GND.t192 19.9612
R29942 GND.n490 GND.t43 19.6726
R29943 GND.n4505 GND.t13 19.6726
R29944 GND.t239 GND.n6663 19.6726
R29945 GND.n9400 GND.n232 19.577
R29946 GND.n9356 GND.n292 19.577
R29947 GND.n786 GND.n474 19.577
R29948 GND.n969 GND.n968 19.577
R29949 GND.n9396 GND.n9395 19.577
R29950 GND.n9361 GND.n9360 19.577
R29951 GND.n850 GND.n849 19.577
R29952 GND.n9016 GND.n9015 19.577
R29953 GND.n835 GND.n830 19.577
R29954 GND.n9056 GND.n441 19.577
R29955 GND.n933 GND.n487 19.577
R29956 GND.n9062 GND.n434 19.577
R29957 GND.n8294 GND.n1924 19.577
R29958 GND.n8250 GND.n1984 19.577
R29959 GND.n4397 GND.n4213 19.577
R29960 GND.n4701 GND.n4700 19.577
R29961 GND.n8290 GND.n8289 19.577
R29962 GND.n8255 GND.n8254 19.577
R29963 GND.n4500 GND.n4499 19.577
R29964 GND.n4759 GND.n4758 19.577
R29965 GND.n4477 GND.n4473 19.577
R29966 GND.n4644 GND.n4642 19.577
R29967 GND.n4461 GND.n4460 19.577
R29968 GND.n4639 GND.n4550 19.577
R29969 GND.n6682 GND.n6681 19.577
R29970 GND.n7372 GND.n2522 19.577
R29971 GND.n7078 GND.n7077 19.577
R29972 GND.n2616 GND.n2615 19.577
R29973 GND.n7131 GND.n7130 19.577
R29974 GND.n7294 GND.n7292 19.577
R29975 GND.n7121 GND.n7120 19.577
R29976 GND.n7326 GND.n7325 19.577
R29977 GND.n7148 GND.n6667 19.577
R29978 GND.n7377 GND.n2513 19.577
R29979 GND.n7160 GND.n6658 19.577
R29980 GND.n2682 GND.n2681 19.577
R29981 GND.n6600 GND.n6599 19.1591
R29982 GND.n6586 GND.n6585 19.1591
R29983 GND.n6572 GND.n6571 19.1591
R29984 GND.n6558 GND.n6557 19.1591
R29985 GND.n6544 GND.n6543 19.1591
R29986 GND.n2710 GND.n2709 19.1591
R29987 GND.n6459 GND.n6458 19.1591
R29988 GND.n6473 GND.n6472 19.1591
R29989 GND.n6486 GND.n6485 19.1591
R29990 GND.n6499 GND.n6498 19.1591
R29991 GND.n6512 GND.n6511 19.1591
R29992 GND.n6525 GND.n6524 19.1591
R29993 GND.n6440 GND.n6439 19.1591
R29994 GND.n8963 GND.n8962 19.1591
R29995 GND.n8949 GND.n8948 19.1591
R29996 GND.n8935 GND.n8934 19.1591
R29997 GND.n8921 GND.n8920 19.1591
R29998 GND.n8907 GND.n8906 19.1591
R29999 GND.n993 GND.n992 19.1591
R30000 GND.n8823 GND.n8822 19.1591
R30001 GND.n8837 GND.n8836 19.1591
R30002 GND.n8850 GND.n8849 19.1591
R30003 GND.n8863 GND.n8862 19.1591
R30004 GND.n8876 GND.n8875 19.1591
R30005 GND.n8889 GND.n8888 19.1591
R30006 GND.n8804 GND.n8803 19.1591
R30007 GND.n4862 GND.n4861 19.1591
R30008 GND.n4848 GND.n4847 19.1591
R30009 GND.n4834 GND.n4833 19.1591
R30010 GND.n4820 GND.n4819 19.1591
R30011 GND.n4806 GND.n4805 19.1591
R30012 GND.n4791 GND.n4790 19.1591
R30013 GND.n4185 GND.n4184 19.1591
R30014 GND.n4879 GND.n4878 19.1591
R30015 GND.n4892 GND.n4891 19.1591
R30016 GND.n4905 GND.n4904 19.1591
R30017 GND.n4918 GND.n4917 19.1591
R30018 GND.n4931 GND.n4930 19.1591
R30019 GND.n4166 GND.n4165 19.1591
R30020 GND.n6593 GND.n6591 18.824
R30021 GND.n6579 GND.n6577 18.824
R30022 GND.n6565 GND.n6563 18.824
R30023 GND.n6551 GND.n6549 18.824
R30024 GND.n6537 GND.n6535 18.824
R30025 GND.n2703 GND.n2701 18.824
R30026 GND.n6452 GND.n6450 18.824
R30027 GND.n6466 GND.n6464 18.824
R30028 GND.n6479 GND.n6477 18.824
R30029 GND.n6492 GND.n6490 18.824
R30030 GND.n6505 GND.n6503 18.824
R30031 GND.n6518 GND.n6516 18.824
R30032 GND.n6433 GND.n6431 18.824
R30033 GND.n8956 GND.n8954 18.824
R30034 GND.n8942 GND.n8940 18.824
R30035 GND.n8928 GND.n8926 18.824
R30036 GND.n8914 GND.n8912 18.824
R30037 GND.n8900 GND.n8898 18.824
R30038 GND.n986 GND.n984 18.824
R30039 GND.n8816 GND.n8814 18.824
R30040 GND.n8830 GND.n8828 18.824
R30041 GND.n8843 GND.n8841 18.824
R30042 GND.n8856 GND.n8854 18.824
R30043 GND.n8869 GND.n8867 18.824
R30044 GND.n8882 GND.n8880 18.824
R30045 GND.n8797 GND.n8795 18.824
R30046 GND.n536 GND.n535 18.824
R30047 GND.n923 GND.n922 18.824
R30048 GND.n9272 GND.n9271 18.824
R30049 GND.n9241 GND.n9240 18.824
R30050 GND.n721 GND.n717 18.824
R30051 GND.n907 GND.n906 18.824
R30052 GND.n9265 GND.n362 18.824
R30053 GND.n9245 GND.n368 18.824
R30054 GND.n4855 GND.n4853 18.824
R30055 GND.n4841 GND.n4839 18.824
R30056 GND.n4827 GND.n4825 18.824
R30057 GND.n4813 GND.n4811 18.824
R30058 GND.n4799 GND.n4797 18.824
R30059 GND.n4784 GND.n4782 18.824
R30060 GND.n4178 GND.n4176 18.824
R30061 GND.n4872 GND.n4870 18.824
R30062 GND.n4885 GND.n4883 18.824
R30063 GND.n4898 GND.n4896 18.824
R30064 GND.n4911 GND.n4909 18.824
R30065 GND.n4924 GND.n4922 18.824
R30066 GND.n4159 GND.n4157 18.824
R30067 GND.n1898 GND.n1869 18.824
R30068 GND.n4520 GND.n4519 18.824
R30069 GND.n8166 GND.n8165 18.824
R30070 GND.n8135 GND.n8134 18.824
R30071 GND.n8323 GND.n1891 18.824
R30072 GND.n4251 GND.n4231 18.824
R30073 GND.n8159 GND.n2054 18.824
R30074 GND.n8139 GND.n2060 18.824
R30075 GND.n6996 GND.n6989 18.824
R30076 GND.n7048 GND.n7046 18.824
R30077 GND.n7285 GND.n2621 18.824
R30078 GND.n7434 GND.n2474 18.824
R30079 GND.n6979 GND.n6975 18.824
R30080 GND.n7042 GND.n7041 18.824
R30081 GND.n7269 GND.n7268 18.824
R30082 GND.n7412 GND.n7411 18.824
R30083 GND.n9798 GND.n49 18.7784
R30084 GND.n8419 GND.n16 18.7784
R30085 GND.n9808 GND.n26 18.7784
R30086 GND.n7734 GND.n2275 18.7784
R30087 GND.n8397 GND.n1814 18.7784
R30088 GND.n7689 GND.n2314 18.7784
R30089 GND.n8032 GND.n8031 18.4271
R30090 GND.n832 GND.n831 18.0711
R30091 GND.n9283 GND.n345 18.0711
R30092 GND.n930 GND.n929 18.0711
R30093 GND.n9066 GND.n9065 18.0711
R30094 GND.n4476 GND.n4474 18.0711
R30095 GND.n8177 GND.n2037 18.0711
R30096 GND.n4457 GND.n4456 18.0711
R30097 GND.n4638 GND.n4551 18.0711
R30098 GND.n7152 GND.n7151 18.0711
R30099 GND.n7379 GND.n7378 18.0711
R30100 GND.n7157 GND.n7156 18.0711
R30101 GND.n2680 GND.n2679 18.0711
R30102 GND.n5022 GND.n5014 17.7398
R30103 GND.n1445 GND.n1444 17.7398
R30104 GND.n3492 GND.n3491 17.7398
R30105 GND.t206 GND.n8974 17.7054
R30106 GND.n4672 GND.t183 17.7054
R30107 GND.t108 GND.n7201 17.7054
R30108 GND.n5895 GND.n3717 17.4326
R30109 GND.n5846 GND.n5845 17.4326
R30110 GND.n4079 GND.n3837 17.4326
R30111 GND.n5400 GND.n4982 17.4326
R30112 GND.n6599 GND.n6590 17.3181
R30113 GND.n6585 GND.n6576 17.3181
R30114 GND.n6571 GND.n6562 17.3181
R30115 GND.n6557 GND.n6548 17.3181
R30116 GND.n6543 GND.n6534 17.3181
R30117 GND.n2709 GND.n2700 17.3181
R30118 GND.n6458 GND.n6449 17.3181
R30119 GND.n6472 GND.n6463 17.3181
R30120 GND.n6485 GND.n6476 17.3181
R30121 GND.n6498 GND.n6489 17.3181
R30122 GND.n6511 GND.n6502 17.3181
R30123 GND.n6524 GND.n6515 17.3181
R30124 GND.n6439 GND.n6430 17.3181
R30125 GND.n8962 GND.n8953 17.3181
R30126 GND.n8948 GND.n8939 17.3181
R30127 GND.n8934 GND.n8925 17.3181
R30128 GND.n8920 GND.n8911 17.3181
R30129 GND.n8906 GND.n8897 17.3181
R30130 GND.n992 GND.n983 17.3181
R30131 GND.n8822 GND.n8813 17.3181
R30132 GND.n8836 GND.n8827 17.3181
R30133 GND.n8849 GND.n8840 17.3181
R30134 GND.n8862 GND.n8853 17.3181
R30135 GND.n8875 GND.n8866 17.3181
R30136 GND.n8888 GND.n8879 17.3181
R30137 GND.n8803 GND.n8794 17.3181
R30138 GND.n9422 GND.n203 17.3181
R30139 GND.n917 GND.n910 17.3181
R30140 GND.n9277 GND.n353 17.3181
R30141 GND.n375 GND.n374 17.3181
R30142 GND.n719 GND.n718 17.3181
R30143 GND.n869 GND.n496 17.3181
R30144 GND.n9262 GND.n9261 17.3181
R30145 GND.n9246 GND.n367 17.3181
R30146 GND.n4861 GND.n4852 17.3181
R30147 GND.n4847 GND.n4838 17.3181
R30148 GND.n4833 GND.n4824 17.3181
R30149 GND.n4819 GND.n4810 17.3181
R30150 GND.n4805 GND.n4796 17.3181
R30151 GND.n4790 GND.n4781 17.3181
R30152 GND.n4184 GND.n4175 17.3181
R30153 GND.n4878 GND.n4869 17.3181
R30154 GND.n4891 GND.n4882 17.3181
R30155 GND.n4904 GND.n4895 17.3181
R30156 GND.n4917 GND.n4908 17.3181
R30157 GND.n4930 GND.n4921 17.3181
R30158 GND.n4165 GND.n4156 17.3181
R30159 GND.n8316 GND.n1899 17.3181
R30160 GND.n4514 GND.n4507 17.3181
R30161 GND.n8171 GND.n2045 17.3181
R30162 GND.n2067 GND.n2066 17.3181
R30163 GND.n8321 GND.n8320 17.3181
R30164 GND.n4250 GND.n4233 17.3181
R30165 GND.n8156 GND.n8155 17.3181
R30166 GND.n8140 GND.n2059 17.3181
R30167 GND.n6995 GND.n6990 17.3181
R30168 GND.n7052 GND.n7051 17.3181
R30169 GND.n7392 GND.n2503 17.3181
R30170 GND.n7432 GND.n7431 17.3181
R30171 GND.n6977 GND.n6976 17.3181
R30172 GND.n7024 GND.n6741 17.3181
R30173 GND.n7266 GND.n7261 17.3181
R30174 GND.n7413 GND.n2491 17.3181
R30175 GND.n5664 GND.n5443 17.2805
R30176 GND.n5452 GND.n5451 17.2805
R30177 GND.n9761 GND.n61 17.2805
R30178 GND.n9757 GND.n9756 17.2805
R30179 GND.n7890 GND.n2203 17.2805
R30180 GND.n2156 GND.n2153 17.2805
R30181 GND.n6349 GND.n6348 16.9869
R30182 GND.n8526 GND.n8525 16.9869
R30183 GND.n3941 GND.n3932 16.9869
R30184 GND.n7493 GND.n7451 16.7316
R30185 GND.n8099 GND.n8032 16.7262
R30186 GND.n615 GND.n573 16.7262
R30187 GND.n8396 GND.n1816 16.7262
R30188 GND.n216 GND.n195 16.5652
R30189 GND.n9407 GND.n222 16.5652
R30190 GND.n9284 GND.n343 16.5652
R30191 GND.n9297 GND.n9296 16.5652
R30192 GND.n741 GND.n739 16.5652
R30193 GND.n526 GND.n489 16.5652
R30194 GND.n9069 GND.n9067 16.5652
R30195 GND.n9080 GND.n428 16.5652
R30196 GND.n4342 GND.n4338 16.5652
R30197 GND.n8301 GND.n1914 16.5652
R30198 GND.n8178 GND.n2035 16.5652
R30199 GND.n8191 GND.n8190 16.5652
R30200 GND.n4351 GND.n4350 16.5652
R30201 GND.n4455 GND.n4262 16.5652
R30202 GND.n4635 GND.n4634 16.5652
R30203 GND.n4623 GND.n4622 16.5652
R30204 GND.n7010 GND.n7003 16.5652
R30205 GND.n7144 GND.n6666 16.5652
R30206 GND.n7387 GND.n2510 16.5652
R30207 GND.n7425 GND.n2483 16.5652
R30208 GND.n6940 GND.n6924 16.5652
R30209 GND.n6928 GND.n6660 16.5652
R30210 GND.n2676 GND.n2644 16.5652
R30211 GND.n2663 GND.n2661 16.5652
R30212 GND.n9235 GND.n380 16.415
R30213 GND.n9234 GND.n383 16.415
R30214 GND.n9087 GND.n391 16.415
R30215 GND.n9155 GND.n394 16.415
R30216 GND.n9221 GND.n400 16.415
R30217 GND.n9220 GND.n403 16.415
R30218 GND.n9096 GND.n409 16.415
R30219 GND.n9214 GND.n9213 16.415
R30220 GND.n9164 GND.n412 16.415
R30221 GND.n6913 GND.n6912 16.415
R30222 GND.n6793 GND.n6785 16.415
R30223 GND.n6955 GND.n6780 16.415
R30224 GND.n6954 GND.n6773 16.415
R30225 GND.n6963 GND.n6962 16.415
R30226 GND.n6948 GND.n6767 16.415
R30227 GND.n6971 GND.n6970 16.415
R30228 GND.n6985 GND.n6762 16.415
R30229 GND.t325 GND.n269 16.3939
R30230 GND.t164 GND.n1961 16.3939
R30231 GND.t120 GND.n2558 16.3939
R30232 GND.n9505 GND.n9464 16.3597
R30233 GND.n7790 GND.n7789 16.3597
R30234 GND.n5658 GND.n5657 16.3205
R30235 GND.n9568 GND.n9567 16.3205
R30236 GND.n7853 GND.n7852 16.3205
R30237 GND.n5665 GND.n5444 16.0005
R30238 GND.n5455 GND.n5450 16.0005
R30239 GND.n9762 GND.n62 16.0005
R30240 GND.n9753 GND.n69 16.0005
R30241 GND.n7888 GND.n7887 16.0005
R30242 GND.n7972 GND.n2152 16.0005
R30243 GND.n3009 GND.n3008 15.8123
R30244 GND.n9421 GND.n204 15.8123
R30245 GND.n918 GND.n916 15.8123
R30246 GND.n9276 GND.n354 15.8123
R30247 GND.n9302 GND.n331 15.8123
R30248 GND.n860 GND.n502 15.8123
R30249 GND.n870 GND.n868 15.8123
R30250 GND.n9260 GND.n9259 15.8123
R30251 GND.n9250 GND.n9249 15.8123
R30252 GND.n8315 GND.n1900 15.8123
R30253 GND.n4515 GND.n4513 15.8123
R30254 GND.n8170 GND.n2046 15.8123
R30255 GND.n8196 GND.n2023 15.8123
R30256 GND.n4237 GND.n1893 15.8123
R30257 GND.n4246 GND.n4245 15.8123
R30258 GND.n8154 GND.n8153 15.8123
R30259 GND.n8144 GND.n8143 15.8123
R30260 GND.n6992 GND.n6991 15.8123
R30261 GND.n7055 GND.n6738 15.8123
R30262 GND.n7394 GND.n7393 15.8123
R30263 GND.n7397 GND.n2476 15.8123
R30264 GND.n7015 GND.n6747 15.8123
R30265 GND.n7025 GND.n7023 15.8123
R30266 GND.n7263 GND.n7262 15.8123
R30267 GND.n7417 GND.n7416 15.8123
R30268 GND.n9398 GND.t237 15.7382
R30269 GND.n8292 GND.t11 15.7382
R30270 GND.n7133 GND.t210 15.7382
R30271 GND.n6598 GND.n6597 15.4484
R30272 GND.n6584 GND.n6583 15.4484
R30273 GND.n6570 GND.n6569 15.4484
R30274 GND.n6556 GND.n6555 15.4484
R30275 GND.n6542 GND.n6541 15.4484
R30276 GND.n2708 GND.n2707 15.4484
R30277 GND.n6457 GND.n6456 15.4484
R30278 GND.n6471 GND.n6470 15.4484
R30279 GND.n6484 GND.n6483 15.4484
R30280 GND.n6497 GND.n6496 15.4484
R30281 GND.n6510 GND.n6509 15.4484
R30282 GND.n6523 GND.n6522 15.4484
R30283 GND.n6438 GND.n6437 15.4484
R30284 GND.n8961 GND.n8960 15.4484
R30285 GND.n8947 GND.n8946 15.4484
R30286 GND.n8933 GND.n8932 15.4484
R30287 GND.n8919 GND.n8918 15.4484
R30288 GND.n8905 GND.n8904 15.4484
R30289 GND.n991 GND.n990 15.4484
R30290 GND.n8821 GND.n8820 15.4484
R30291 GND.n8835 GND.n8834 15.4484
R30292 GND.n8848 GND.n8847 15.4484
R30293 GND.n8861 GND.n8860 15.4484
R30294 GND.n8874 GND.n8873 15.4484
R30295 GND.n8887 GND.n8886 15.4484
R30296 GND.n8802 GND.n8801 15.4484
R30297 GND.n4860 GND.n4859 15.4484
R30298 GND.n4846 GND.n4845 15.4484
R30299 GND.n4832 GND.n4831 15.4484
R30300 GND.n4818 GND.n4817 15.4484
R30301 GND.n4804 GND.n4803 15.4484
R30302 GND.n4789 GND.n4788 15.4484
R30303 GND.n4183 GND.n4182 15.4484
R30304 GND.n4877 GND.n4876 15.4484
R30305 GND.n4890 GND.n4889 15.4484
R30306 GND.n4903 GND.n4902 15.4484
R30307 GND.n4916 GND.n4915 15.4484
R30308 GND.n4929 GND.n4928 15.4484
R30309 GND.n4164 GND.n4163 15.4484
R30310 GND.n9345 GND.n301 15.0825
R30311 GND.n8239 GND.n1993 15.0825
R30312 GND.n2498 GND.n2487 15.0825
R30313 GND.n218 GND.n217 15.0593
R30314 GND.n9408 GND.n215 15.0593
R30315 GND.n9288 GND.n9287 15.0593
R30316 GND.n9292 GND.n338 15.0593
R30317 GND.n743 GND.n742 15.0593
R30318 GND.n750 GND.n749 15.0593
R30319 GND.n9070 GND.n432 15.0593
R30320 GND.n9078 GND.n9077 15.0593
R30321 GND.n4340 GND.n4339 15.0593
R30322 GND.n8302 GND.n1911 15.0593
R30323 GND.n8182 GND.n8181 15.0593
R30324 GND.n8186 GND.n2030 15.0593
R30325 GND.n4355 GND.n4272 15.0593
R30326 GND.n4452 GND.n4451 15.0593
R30327 GND.n4631 GND.n4554 15.0593
R30328 GND.n4626 GND.n4624 15.0593
R30329 GND.n7009 GND.n7004 15.0593
R30330 GND.n7145 GND.n7143 15.0593
R30331 GND.n7386 GND.n2511 15.0593
R30332 GND.n7423 GND.n7422 15.0593
R30333 GND.n6938 GND.n6937 15.0593
R30334 GND.n6929 GND.n6927 15.0593
R30335 GND.n2673 GND.n2672 15.0593
R30336 GND.n2664 GND.n2647 15.0593
R30337 GND.n5654 GND.n5448 15.0405
R30338 GND.n9571 GND.n9570 15.0405
R30339 GND.n7851 GND.n7850 15.0405
R30340 GND.t55 GND.n9680 14.9707
R30341 GND.n8029 GND.t167 14.9707
R30342 GND.n5509 GND.n5442 14.7205
R30343 GND.n5456 GND.n2354 14.7205
R30344 GND.n9519 GND.n60 14.7205
R30345 GND.n9754 GND.n9752 14.7205
R30346 GND.n7886 GND.n7885 14.7205
R30347 GND.n7973 GND.n2154 14.7205
R30348 GND.n9235 GND.n9234 14.5912
R30349 GND.n9087 GND.n383 14.5912
R30350 GND.n9228 GND.n391 14.5912
R30351 GND.n9227 GND.n394 14.5912
R30352 GND.n9155 GND.n400 14.5912
R30353 GND.n9221 GND.n9220 14.5912
R30354 GND.n9214 GND.n409 14.5912
R30355 GND.n9213 GND.n412 14.5912
R30356 GND.n6913 GND.n6790 14.5912
R30357 GND.n6912 GND.n6793 14.5912
R30358 GND.n6920 GND.n6785 14.5912
R30359 GND.n6855 GND.n6780 14.5912
R30360 GND.n6955 GND.n6954 14.5912
R30361 GND.n6963 GND.n6773 14.5912
R30362 GND.n6970 GND.n6767 14.5912
R30363 GND.n6971 GND.n6762 14.5912
R30364 GND.n6985 GND.n6984 14.5912
R30365 GND.n3080 GND.t363 14.57
R30366 GND.n9046 GND.t10 14.4267
R30367 GND.t5 GND.n4196 14.4267
R30368 GND.n2689 GND.t52 14.4267
R30369 GND.n7748 GND.t376 14.3158
R30370 GND.n2974 GND.n2973 14.3064
R30371 GND.n3008 GND.n3007 14.3064
R30372 GND.n9418 GND.n9417 14.3064
R30373 GND.n914 GND.n913 14.3064
R30374 GND.n9307 GND.n327 14.3064
R30375 GND.n9303 GND.n328 14.3064
R30376 GND.n861 GND.n500 14.3064
R30377 GND.n865 GND.n499 14.3064
R30378 GND.n9257 GND.n365 14.3064
R30379 GND.n9253 GND.n9251 14.3064
R30380 GND.n8312 GND.n8311 14.3064
R30381 GND.n4511 GND.n4510 14.3064
R30382 GND.n8201 GND.n2019 14.3064
R30383 GND.n8197 GND.n2020 14.3064
R30384 GND.n4238 GND.n4236 14.3064
R30385 GND.n4242 GND.n4235 14.3064
R30386 GND.n8151 GND.n2057 14.3064
R30387 GND.n8147 GND.n8145 14.3064
R30388 GND.n7060 GND.n6734 14.3064
R30389 GND.n7056 GND.n6735 14.3064
R30390 GND.n7402 GND.n2500 14.3064
R30391 GND.n7398 GND.n2501 14.3064
R30392 GND.n7016 GND.n6745 14.3064
R30393 GND.n7020 GND.n6744 14.3064
R30394 GND.n7406 GND.n2493 14.3064
R30395 GND.n7407 GND.n2490 14.3064
R30396 GND.n7647 GND.n2331 13.9936
R30397 GND.n7641 GND.n7640 13.9936
R30398 GND.n7591 GND.n7590 13.9936
R30399 GND.n7590 GND.n7589 13.9936
R30400 GND.n5553 GND.t80 13.9205
R30401 GND.n5553 GND.t191 13.9205
R30402 GND.n132 GND.t268 13.9205
R30403 GND.n132 GND.t313 13.9205
R30404 GND.n2148 GND.t356 13.9205
R30405 GND.n2148 GND.t176 13.9205
R30406 GND.n5809 GND.n3789 13.875
R30407 GND.n5655 GND.n5653 13.7605
R30408 GND.n5484 GND.n5483 13.7605
R30409 GND.n5488 GND.n5486 13.7605
R30410 GND.n9574 GND.n9564 13.7605
R30411 GND.n9726 GND.n100 13.7605
R30412 GND.n135 GND.n133 13.7605
R30413 GND.n7849 GND.n7848 13.7605
R30414 GND.n7947 GND.n2183 13.7605
R30415 GND.n2241 GND.n2229 13.7605
R30416 GND.n9412 GND.n214 13.5534
R30417 GND.n9412 GND.n9411 13.5534
R30418 GND.n9291 GND.n341 13.5534
R30419 GND.n9293 GND.n9291 13.5534
R30420 GND.n745 GND.n744 13.5534
R30421 GND.n744 GND.n525 13.5534
R30422 GND.n9074 GND.n9073 13.5534
R30423 GND.n9074 GND.n430 13.5534
R30424 GND.n8306 GND.n1910 13.5534
R30425 GND.n8306 GND.n8305 13.5534
R30426 GND.n8185 GND.n2033 13.5534
R30427 GND.n8187 GND.n8185 13.5534
R30428 GND.n4354 GND.n4273 13.5534
R30429 GND.n4273 GND.n4264 13.5534
R30430 GND.n4630 GND.n4556 13.5534
R30431 GND.n4627 GND.n4556 13.5534
R30432 GND.n7006 GND.n7005 13.5534
R30433 GND.n7005 GND.n6669 13.5534
R30434 GND.n7383 GND.n7382 13.5534
R30435 GND.n7382 GND.n2485 13.5534
R30436 GND.n6933 GND.n6926 13.5534
R30437 GND.n6933 GND.n6932 13.5534
R30438 GND.n2668 GND.n2646 13.5534
R30439 GND.n2668 GND.n2667 13.5534
R30440 GND.n7639 GND.n2339 13.3762
R30441 GND.n7633 GND.n7632 13.3762
R30442 GND.n7626 GND.n2356 13.3762
R30443 GND.n7618 GND.n2368 13.3762
R30444 GND.n5605 GND.n5562 13.3762
R30445 GND.n7604 GND.n2390 13.3762
R30446 GND.n7598 GND.n7597 13.3762
R30447 GND.n5558 GND.n2399 13.3762
R30448 GND.t235 GND.n9227 13.2233
R30449 GND.n5696 GND.n5004 13.2221
R30450 GND.n1435 GND.n1433 13.2221
R30451 GND.n3482 GND.n3480 13.2221
R30452 GND.t219 GND.t192 13.1869
R30453 GND.t167 GND.t301 13.1826
R30454 GND.t2 GND.n286 13.1153
R30455 GND.t415 GND.n1978 13.1153
R30456 GND.n7375 GND.t74 13.1153
R30457 GND.n9417 GND.n207 12.8005
R30458 GND.n913 GND.n207 12.8005
R30459 GND.n9307 GND.n9306 12.8005
R30460 GND.n9306 GND.n328 12.8005
R30461 GND.n864 GND.n500 12.8005
R30462 GND.n865 GND.n864 12.8005
R30463 GND.n9254 GND.n365 12.8005
R30464 GND.n9254 GND.n9253 12.8005
R30465 GND.n8311 GND.n1903 12.8005
R30466 GND.n4510 GND.n1903 12.8005
R30467 GND.n8201 GND.n8200 12.8005
R30468 GND.n8200 GND.n2020 12.8005
R30469 GND.n4241 GND.n4236 12.8005
R30470 GND.n4242 GND.n4241 12.8005
R30471 GND.n8148 GND.n2057 12.8005
R30472 GND.n8148 GND.n8147 12.8005
R30473 GND.n7060 GND.n7059 12.8005
R30474 GND.n7059 GND.n6735 12.8005
R30475 GND.n7402 GND.n7401 12.8005
R30476 GND.n7401 GND.n2501 12.8005
R30477 GND.n7019 GND.n6745 12.8005
R30478 GND.n7020 GND.n7019 12.8005
R30479 GND.n7408 GND.n7406 12.8005
R30480 GND.n7408 GND.n7407 12.8005
R30481 GND.n3103 GND.n2712 12.7044
R30482 GND.n5633 GND.n5468 12.4805
R30483 GND.n5526 GND.n5525 12.4805
R30484 GND.n9724 GND.n9723 12.4805
R30485 GND.n9600 GND.n9599 12.4805
R30486 GND.n7945 GND.n7944 12.4805
R30487 GND.n2245 GND.n2244 12.4805
R30488 GND.n6422 GND.n6421 12.4692
R30489 GND.n8786 GND.n8785 12.4692
R30490 GND.n4149 GND.n4148 12.4692
R30491 GND.n9281 GND.t244 12.4595
R30492 GND.t240 GND.n372 12.4595
R30493 GND.n8175 GND.t211 12.4595
R30494 GND.t301 GND.n2064 12.4595
R30495 GND.n2677 GND.t75 12.4595
R30496 GND.n2657 GND.t219 12.4595
R30497 GND.n6962 GND.t114 12.3114
R30498 GND.n217 GND.n214 12.0476
R30499 GND.n9411 GND.n215 12.0476
R30500 GND.n9288 GND.n341 12.0476
R30501 GND.n9293 GND.n9292 12.0476
R30502 GND.n745 GND.n743 12.0476
R30503 GND.n750 GND.n525 12.0476
R30504 GND.n9073 GND.n432 12.0476
R30505 GND.n9077 GND.n430 12.0476
R30506 GND.n4339 GND.n1910 12.0476
R30507 GND.n8305 GND.n1911 12.0476
R30508 GND.n8182 GND.n2033 12.0476
R30509 GND.n8187 GND.n8186 12.0476
R30510 GND.n4355 GND.n4354 12.0476
R30511 GND.n4451 GND.n4264 12.0476
R30512 GND.n4631 GND.n4630 12.0476
R30513 GND.n4627 GND.n4626 12.0476
R30514 GND.n7006 GND.n7004 12.0476
R30515 GND.n7143 GND.n6669 12.0476
R30516 GND.n7383 GND.n2511 12.0476
R30517 GND.n7422 GND.n2485 12.0476
R30518 GND.n6937 GND.n6926 12.0476
R30519 GND.n6932 GND.n6927 12.0476
R30520 GND.n2672 GND.n2646 12.0476
R30521 GND.n2667 GND.n2647 12.0476
R30522 GND.n856 GND.t255 11.8038
R30523 GND.n463 GND.t41 11.8038
R30524 GND.n4440 GND.t155 11.8038
R30525 GND.n4490 GND.t305 11.8038
R30526 GND.n7113 GND.t410 11.8038
R30527 GND.n6629 GND.t300 11.8038
R30528 GND.n9505 GND.n9463 11.7297
R30529 GND.n7789 GND.n7748 11.7297
R30530 GND.n3107 GND.n3106 11.5593
R30531 GND.n6855 GND.t284 11.3995
R30532 GND.n5458 GND.n5441 11.3205
R30533 GND.n5668 GND.n5667 11.3205
R30534 GND.n7726 GND.n7725 11.3205
R30535 GND.n7726 GND.n2295 11.3205
R30536 GND.n71 GND.n59 11.3205
R30537 GND.n9765 GND.n9764 11.3205
R30538 GND.n7976 GND.n7975 11.3205
R30539 GND.n2204 GND.n2150 11.3205
R30540 GND.n5622 GND.n5558 11.3184
R30541 GND.n3108 GND.n3107 11.2946
R30542 GND.n9418 GND.n204 11.2946
R30543 GND.n916 GND.n914 11.2946
R30544 GND.n354 GND.n327 11.2946
R30545 GND.n9303 GND.n9302 11.2946
R30546 GND.n861 GND.n860 11.2946
R30547 GND.n868 GND.n499 11.2946
R30548 GND.n9259 GND.n9257 11.2946
R30549 GND.n9251 GND.n9250 11.2946
R30550 GND.n8312 GND.n1900 11.2946
R30551 GND.n4513 GND.n4511 11.2946
R30552 GND.n2046 GND.n2019 11.2946
R30553 GND.n8197 GND.n8196 11.2946
R30554 GND.n4238 GND.n4237 11.2946
R30555 GND.n4245 GND.n4235 11.2946
R30556 GND.n8153 GND.n8151 11.2946
R30557 GND.n8145 GND.n8144 11.2946
R30558 GND.n6991 GND.n6734 11.2946
R30559 GND.n7056 GND.n7055 11.2946
R30560 GND.n7393 GND.n2500 11.2946
R30561 GND.n7398 GND.n7397 11.2946
R30562 GND.n7016 GND.n7015 11.2946
R30563 GND.n7023 GND.n6744 11.2946
R30564 GND.n7262 GND.n2493 11.2946
R30565 GND.n7417 GND.n2490 11.2946
R30566 GND.n5632 GND.n5466 11.2005
R30567 GND.n5490 GND.n5487 11.2005
R30568 GND.n9720 GND.n9719 11.2005
R30569 GND.n137 GND.n134 11.2005
R30570 GND.n7941 GND.n7940 11.2005
R30571 GND.n2248 GND.n2228 11.2005
R30572 GND.n735 GND.t225 11.148
R30573 GND.n857 GND.n856 11.148
R30574 GND.n926 GND.t257 11.148
R30575 GND.n4346 GND.t72 11.148
R30576 GND.n4440 GND.n4357 11.148
R30577 GND.n4503 GND.t428 11.148
R30578 GND.n6999 GND.t201 11.148
R30579 GND.n7113 GND.n6693 11.148
R30580 GND.t77 GND.n6664 11.148
R30581 GND.n9817 GND.n17 11.0565
R30582 GND.n6984 GND.n6983 10.9922
R30583 GND.n5541 GND.t400 10.7011
R30584 GND.t401 GND.n2396 10.7011
R30585 GND.n5633 GND.n5632 10.5605
R30586 GND.n5525 GND.n5487 10.5605
R30587 GND.n9723 GND.n9720 10.5605
R30588 GND.n9599 GND.n134 10.5605
R30589 GND.n7944 GND.n7941 10.5605
R30590 GND.n2245 GND.n2228 10.5605
R30591 GND.n218 GND.n216 10.5417
R30592 GND.n9408 GND.n9407 10.5417
R30593 GND.n9287 GND.n343 10.5417
R30594 GND.n9297 GND.n338 10.5417
R30595 GND.n742 GND.n741 10.5417
R30596 GND.n749 GND.n526 10.5417
R30597 GND.n9070 GND.n9069 10.5417
R30598 GND.n9078 GND.n428 10.5417
R30599 GND.n4340 GND.n4338 10.5417
R30600 GND.n8302 GND.n8301 10.5417
R30601 GND.n8181 GND.n2035 10.5417
R30602 GND.n8191 GND.n2030 10.5417
R30603 GND.n4350 GND.n4272 10.5417
R30604 GND.n4452 GND.n4262 10.5417
R30605 GND.n4634 GND.n4554 10.5417
R30606 GND.n4624 GND.n4623 10.5417
R30607 GND.n7010 GND.n7009 10.5417
R30608 GND.n7145 GND.n7144 10.5417
R30609 GND.n7387 GND.n7386 10.5417
R30610 GND.n7423 GND.n2483 10.5417
R30611 GND.n6938 GND.n6924 10.5417
R30612 GND.n6929 GND.n6928 10.5417
R30613 GND.n2673 GND.n2644 10.5417
R30614 GND.n2664 GND.n2663 10.5417
R30615 GND.n9512 GND.n9511 10.4951
R30616 GND.n9540 GND.n176 10.4951
R30617 GND.n9687 GND.n9617 10.4951
R30618 GND.n9681 GND.n9617 10.4951
R30619 GND.n7808 GND.n7807 10.4951
R30620 GND.n7817 GND.n2263 10.4951
R30621 GND.n7993 GND.n2133 10.4951
R30622 GND.n7994 GND.n7993 10.4951
R30623 GND.t259 GND.n403 10.4875
R30624 GND.n6099 GND.n3113 10.4497
R30625 GND.n5894 GND.n3725 10.3174
R30626 GND.n5279 GND.n3731 10.3174
R30627 GND.n5888 GND.n5887 10.3174
R30628 GND.n3957 GND.n3734 10.3174
R30629 GND.n5881 GND.n3742 10.3174
R30630 GND.n5880 GND.n3745 10.3174
R30631 GND.n5288 GND.n3751 10.3174
R30632 GND.n5874 GND.n5873 10.3174
R30633 GND.n5867 GND.n3760 10.3174
R30634 GND.n5866 GND.n3763 10.3174
R30635 GND.n5297 GND.n3769 10.3174
R30636 GND.n5860 GND.n5859 10.3174
R30637 GND.n3975 GND.n3772 10.3174
R30638 GND.n5853 GND.n3778 10.3174
R30639 GND.n5852 GND.n3781 10.3174
R30640 GND.n5306 GND.n3787 10.3174
R30641 GND.n5778 GND.n3843 10.3174
R30642 GND.n5777 GND.n3846 10.3174
R30643 GND.n5372 GND.n3852 10.3174
R30644 GND.n5771 GND.n5770 10.3174
R30645 GND.n4088 GND.n3855 10.3174
R30646 GND.n5764 GND.n3861 10.3174
R30647 GND.n5763 GND.n3864 10.3174
R30648 GND.n5381 GND.n3870 10.3174
R30649 GND.n4097 GND.n3873 10.3174
R30650 GND.n5750 GND.n3879 10.3174
R30651 GND.n5749 GND.n3882 10.3174
R30652 GND.n5390 GND.n3888 10.3174
R30653 GND.n5743 GND.n5742 10.3174
R30654 GND.n4106 GND.n3891 10.3174
R30655 GND.n5736 GND.n3897 10.3174
R30656 GND.n5735 GND.n3900 10.3174
R30657 GND.n7641 GND.n2335 10.0837
R30658 GND.n175 GND.n171 10.0321
R30659 GND.n9532 GND.n166 10.0321
R30660 GND.n9522 GND.n160 10.0321
R30661 GND.n9759 GND.n65 10.0321
R30662 GND.n9709 GND.n90 10.0321
R30663 GND.n9703 GND.n9702 10.0321
R30664 GND.n9696 GND.n118 10.0321
R30665 GND.n9695 GND.n121 10.0321
R30666 GND.n2262 GND.n2257 10.0321
R30667 GND.n7867 GND.n2219 10.0321
R30668 GND.n7874 GND.n7873 10.0321
R30669 GND.n2253 GND.n2160 10.0321
R30670 GND.n7930 GND.n2174 10.0321
R30671 GND.n7924 GND.n7923 10.0321
R30672 GND.n7910 GND.n7905 10.0321
R30673 GND.n7987 GND.n2137 10.0321
R30674 GND.n380 GND.n379 9.91643
R30675 GND.n9422 GND.n9421 9.78874
R30676 GND.n918 GND.n917 9.78874
R30677 GND.n9277 GND.n9276 9.78874
R30678 GND.n374 GND.n331 9.78874
R30679 GND.n718 GND.n502 9.78874
R30680 GND.n870 GND.n869 9.78874
R30681 GND.n9261 GND.n9260 9.78874
R30682 GND.n9249 GND.n367 9.78874
R30683 GND.n8316 GND.n8315 9.78874
R30684 GND.n4515 GND.n4514 9.78874
R30685 GND.n8171 GND.n8170 9.78874
R30686 GND.n2066 GND.n2023 9.78874
R30687 GND.n8320 GND.n1893 9.78874
R30688 GND.n4246 GND.n4233 9.78874
R30689 GND.n8155 GND.n8154 9.78874
R30690 GND.n8143 GND.n2059 9.78874
R30691 GND.n6992 GND.n6990 9.78874
R30692 GND.n7052 GND.n6738 9.78874
R30693 GND.n7394 GND.n7392 9.78874
R30694 GND.n7431 GND.n2476 9.78874
R30695 GND.n6976 GND.n6747 9.78874
R30696 GND.n7025 GND.n7024 9.78874
R30697 GND.n7263 GND.n7261 9.78874
R30698 GND.n7416 GND.n2491 9.78874
R30699 GND.n7500 GND.n7451 9.64216
R30700 GND.n8100 GND.n8099 9.63905
R30701 GND.n632 GND.n573 9.63905
R30702 GND.n8360 GND.n1816 9.63905
R30703 GND.n7414 GND.n7411 9.49615
R30704 GND.n9247 GND.n368 9.49615
R30705 GND.n739 GND.n527 9.49615
R30706 GND.n849 GND.n848 9.49615
R30707 GND.n9395 GND.n9394 9.49615
R30708 GND.n9362 GND.n9361 9.49615
R30709 GND.n969 GND.n964 9.49615
R30710 GND.n474 GND.n473 9.49615
R30711 GND.n252 GND.n232 9.49615
R30712 GND.n292 GND.n272 9.49615
R30713 GND.n9296 GND.n9295 9.49615
R30714 GND.n9017 GND.n9016 9.49615
R30715 GND.n219 GND.n195 9.49615
R30716 GND.n9240 GND.n9239 9.49615
R30717 GND.n9080 GND.n9079 9.49615
R30718 GND.n536 GND.n205 9.49615
R30719 GND.n721 GND.n720 9.49615
R30720 GND.n8141 GND.n2060 9.49615
R30721 GND.n4352 GND.n4351 9.49615
R30722 GND.n4499 GND.n4498 9.49615
R30723 GND.n8289 GND.n8288 9.49615
R30724 GND.n8256 GND.n8255 9.49615
R30725 GND.n4701 GND.n4697 9.49615
R30726 GND.n4213 GND.n4212 9.49615
R30727 GND.n1944 GND.n1924 9.49615
R30728 GND.n1984 GND.n1964 9.49615
R30729 GND.n8190 GND.n8189 9.49615
R30730 GND.n4759 GND.n4203 9.49615
R30731 GND.n4342 GND.n4341 9.49615
R30732 GND.n8134 GND.n8133 9.49615
R30733 GND.n4622 GND.n4557 9.49615
R30734 GND.n1901 GND.n1869 9.49615
R30735 GND.n8323 GND.n8322 9.49615
R30736 GND.n6994 GND.n6989 9.49615
R30737 GND.n7434 GND.n7433 9.49615
R30738 GND.n2665 GND.n2661 9.49615
R30739 GND.n6940 GND.n6939 9.49615
R30740 GND.n7120 GND.n6641 9.49615
R30741 GND.n7077 GND.n7076 9.49615
R30742 GND.n6681 GND.n6615 9.49615
R30743 GND.n7316 GND.n2522 9.49615
R30744 GND.n7294 GND.n7293 9.49615
R30745 GND.n2616 GND.n2566 9.49615
R30746 GND.n7130 GND.n6626 9.49615
R30747 GND.n7425 GND.n7424 9.49615
R30748 GND.n7325 GND.n7324 9.49615
R30749 GND.n7008 GND.n7003 9.49615
R30750 GND.n6979 GND.n6978 9.49615
R30751 GND.n5552 GND.n5551 9.43925
R30752 GND.n9544 GND.n131 9.43925
R30753 GND.n7821 GND.n2147 9.43925
R30754 GND.n5627 GND.n5626 9.4255
R30755 GND.n9607 GND.n9606 9.4255
R30756 GND.n7980 GND.n7979 9.4255
R30757 GND.n5485 GND.n5484 9.39047
R30758 GND.n5527 GND.n5487 9.39047
R30759 GND.n9726 GND.n9725 9.39047
R30760 GND.n9601 GND.n134 9.39047
R30761 GND.n7947 GND.n7946 9.39047
R30762 GND.n2243 GND.n2228 9.39047
R30763 GND.n5666 GND.n5443 9.3755
R30764 GND.n7696 GND.n7695 9.3755
R30765 GND.n9763 GND.n61 9.3755
R30766 GND.n7890 GND.n7889 9.3755
R30767 GND.n2116 GND.n2115 9.3755
R30768 GND.n5528 GND.n5486 9.3709
R30769 GND.n5632 GND.n5631 9.3709
R30770 GND.n9602 GND.n133 9.3709
R30771 GND.n9720 GND.n101 9.3709
R30772 GND.n2242 GND.n2241 9.3709
R30773 GND.n7941 GND.n2184 9.3709
R30774 GND.n5667 GND.n5442 9.37029
R30775 GND.n9764 GND.n60 9.37029
R30776 GND.n7886 GND.n2204 9.37029
R30777 GND.n678 GND.n639 9.35557
R30778 GND.n8354 GND.n1835 9.35557
R30779 GND.n5014 GND.n5013 9.30943
R30780 GND.n5436 GND.n5435 9.30943
R30781 GND.n5006 GND.n5004 9.30943
R30782 GND.n5690 GND.n5008 9.30943
R30783 GND.n6355 GND.n6354 9.30943
R30784 GND.n6350 GND.n6349 9.30943
R30785 GND.n6340 GND.n6339 9.30943
R30786 GND.n6423 GND.n6422 9.30943
R30787 GND.n8519 GND.n8518 9.30943
R30788 GND.n8787 GND.n8786 9.30943
R30789 GND.n1444 GND.n1443 9.30943
R30790 GND.n1463 GND.n1462 9.30943
R30791 GND.n1435 GND.n1434 9.30943
R30792 GND.n1452 GND.n1451 9.30943
R30793 GND.n8532 GND.n8531 9.30943
R30794 GND.n8527 GND.n8526 9.30943
R30795 GND.n3491 GND.n3490 9.30943
R30796 GND.n3506 GND.n3505 9.30943
R30797 GND.n3482 GND.n3481 9.30943
R30798 GND.n3499 GND.n3498 9.30943
R30799 GND.n3930 GND.n3928 9.30943
R30800 GND.n4944 GND.n3932 9.30943
R30801 GND.n3938 GND.n3937 9.30943
R30802 GND.n4150 GND.n4149 9.30943
R30803 GND.n6590 GND.n6589 9.3005
R30804 GND.n6594 GND.n6593 9.3005
R30805 GND.n6596 GND.n6595 9.3005
R30806 GND.n6576 GND.n6575 9.3005
R30807 GND.n6580 GND.n6579 9.3005
R30808 GND.n6582 GND.n6581 9.3005
R30809 GND.n6562 GND.n6561 9.3005
R30810 GND.n6566 GND.n6565 9.3005
R30811 GND.n6568 GND.n6567 9.3005
R30812 GND.n6548 GND.n6547 9.3005
R30813 GND.n6552 GND.n6551 9.3005
R30814 GND.n6554 GND.n6553 9.3005
R30815 GND.n6534 GND.n6533 9.3005
R30816 GND.n6538 GND.n6537 9.3005
R30817 GND.n6540 GND.n6539 9.3005
R30818 GND.n2700 GND.n2699 9.3005
R30819 GND.n2704 GND.n2703 9.3005
R30820 GND.n2706 GND.n2705 9.3005
R30821 GND.n6449 GND.n6448 9.3005
R30822 GND.n6453 GND.n6452 9.3005
R30823 GND.n6455 GND.n6454 9.3005
R30824 GND.n6463 GND.n6462 9.3005
R30825 GND.n6467 GND.n6466 9.3005
R30826 GND.n6469 GND.n6468 9.3005
R30827 GND.n6476 GND.n6475 9.3005
R30828 GND.n6480 GND.n6479 9.3005
R30829 GND.n6482 GND.n6481 9.3005
R30830 GND.n6489 GND.n6488 9.3005
R30831 GND.n6493 GND.n6492 9.3005
R30832 GND.n6495 GND.n6494 9.3005
R30833 GND.n6502 GND.n6501 9.3005
R30834 GND.n6506 GND.n6505 9.3005
R30835 GND.n6508 GND.n6507 9.3005
R30836 GND.n6515 GND.n6514 9.3005
R30837 GND.n6519 GND.n6518 9.3005
R30838 GND.n6521 GND.n6520 9.3005
R30839 GND.n6430 GND.n6429 9.3005
R30840 GND.n6434 GND.n6433 9.3005
R30841 GND.n6436 GND.n6435 9.3005
R30842 GND.n5692 GND.n5691 9.3005
R30843 GND.n5026 GND.n5012 9.3005
R30844 GND.n6329 GND.n6328 9.3005
R30845 GND.n6337 GND.n2716 9.3005
R30846 GND.n3104 GND.n2893 9.3005
R30847 GND.n3011 GND.n2915 9.3005
R30848 GND.n2896 GND.n2895 9.3005
R30849 GND.n3101 GND.n3100 9.3005
R30850 GND.n3093 GND.n3092 9.3005
R30851 GND.n3085 GND.n2901 9.3005
R30852 GND.n3084 GND.n2900 9.3005
R30853 GND.n3053 GND.n2902 9.3005
R30854 GND.n3051 GND.n3050 9.3005
R30855 GND.n3060 GND.n3059 9.3005
R30856 GND.n3062 GND.n3061 9.3005
R30857 GND.n3044 GND.n3042 9.3005
R30858 GND.n3068 GND.n3067 9.3005
R30859 GND.n3070 GND.n3069 9.3005
R30860 GND.n3040 GND.n3036 9.3005
R30861 GND.n3075 GND.n2907 9.3005
R30862 GND.n3035 GND.n3034 9.3005
R30863 GND.n3031 GND.n3030 9.3005
R30864 GND.n3028 GND.n2910 9.3005
R30865 GND.n3020 GND.n2911 9.3005
R30866 GND.n3022 GND.n3021 9.3005
R30867 GND.n3019 GND.n3018 9.3005
R30868 GND.n3010 GND.n3009 9.3005
R30869 GND.n3006 GND.n3005 9.3005
R30870 GND.n3003 GND.n3002 9.3005
R30871 GND.n2972 GND.n2971 9.3005
R30872 GND.n2977 GND.n2976 9.3005
R30873 GND.n2980 GND.n2979 9.3005
R30874 GND.n2969 GND.n2966 9.3005
R30875 GND.n2986 GND.n2985 9.3005
R30876 GND.n2988 GND.n2987 9.3005
R30877 GND.n2962 GND.n2958 9.3005
R30878 GND.n2994 GND.n2926 9.3005
R30879 GND.n2957 GND.n2956 9.3005
R30880 GND.n2939 GND.n2938 9.3005
R30881 GND.n2945 GND.n2944 9.3005
R30882 GND.n2943 GND.n2930 9.3005
R30883 GND.n2950 GND.n2929 9.3005
R30884 GND.n2953 GND.n2952 9.3005
R30885 GND.n2932 GND.n2931 9.3005
R30886 GND.n2947 GND.n2946 9.3005
R30887 GND.n2949 GND.n2948 9.3005
R30888 GND.n2951 GND.n2928 9.3005
R30889 GND.n2955 GND.n2927 9.3005
R30890 GND.n2996 GND.n2995 9.3005
R30891 GND.n2993 GND.n2992 9.3005
R30892 GND.n2990 GND.n2989 9.3005
R30893 GND.n2965 GND.n2961 9.3005
R30894 GND.n2984 GND.n2983 9.3005
R30895 GND.n2982 GND.n2981 9.3005
R30896 GND.n2968 GND.n2967 9.3005
R30897 GND.n2975 GND.n2974 9.3005
R30898 GND.n2922 GND.n2921 9.3005
R30899 GND.n3004 GND.n2920 9.3005
R30900 GND.n3007 GND.n2918 9.3005
R30901 GND.n3013 GND.n3012 9.3005
R30902 GND.n3017 GND.n3016 9.3005
R30903 GND.n2914 GND.n2913 9.3005
R30904 GND.n3024 GND.n3023 9.3005
R30905 GND.n3027 GND.n3026 9.3005
R30906 GND.n3029 GND.n2909 9.3005
R30907 GND.n3033 GND.n2908 9.3005
R30908 GND.n3077 GND.n3076 9.3005
R30909 GND.n3074 GND.n3073 9.3005
R30910 GND.n3072 GND.n3071 9.3005
R30911 GND.n3043 GND.n3038 9.3005
R30912 GND.n3066 GND.n3065 9.3005
R30913 GND.n3064 GND.n3063 9.3005
R30914 GND.n3052 GND.n3049 9.3005
R30915 GND.n3058 GND.n3057 9.3005
R30916 GND.n3055 GND.n3054 9.3005
R30917 GND.n3083 GND.n3082 9.3005
R30918 GND.n3087 GND.n3086 9.3005
R30919 GND.n2898 GND.n2897 9.3005
R30920 GND.n3095 GND.n3094 9.3005
R30921 GND.n3099 GND.n3098 9.3005
R30922 GND.n3097 GND.n2894 9.3005
R30923 GND.n5666 GND.n5665 9.3005
R30924 GND.n5457 GND.n5451 9.3005
R30925 GND.n5457 GND.n5450 9.3005
R30926 GND.n5457 GND.n5456 9.3005
R30927 GND.n5656 GND.n5655 9.3005
R30928 GND.n5656 GND.n5448 9.3005
R30929 GND.n5657 GND.n5656 9.3005
R30930 GND.n5485 GND.n5468 9.3005
R30931 GND.n5527 GND.n5526 9.3005
R30932 GND.n7709 GND.n7708 9.3005
R30933 GND.n7711 GND.n7710 9.3005
R30934 GND.n7707 GND.n2306 9.3005
R30935 GND.n7724 GND.n7723 9.3005
R30936 GND.n2299 GND.n2297 9.3005
R30937 GND.n2298 GND.n2296 9.3005
R30938 GND.n7699 GND.n7698 9.3005
R30939 GND.n8953 GND.n8952 9.3005
R30940 GND.n8957 GND.n8956 9.3005
R30941 GND.n8959 GND.n8958 9.3005
R30942 GND.n8939 GND.n8938 9.3005
R30943 GND.n8943 GND.n8942 9.3005
R30944 GND.n8945 GND.n8944 9.3005
R30945 GND.n8925 GND.n8924 9.3005
R30946 GND.n8929 GND.n8928 9.3005
R30947 GND.n8931 GND.n8930 9.3005
R30948 GND.n8911 GND.n8910 9.3005
R30949 GND.n8915 GND.n8914 9.3005
R30950 GND.n8917 GND.n8916 9.3005
R30951 GND.n8897 GND.n8896 9.3005
R30952 GND.n8901 GND.n8900 9.3005
R30953 GND.n8903 GND.n8902 9.3005
R30954 GND.n983 GND.n982 9.3005
R30955 GND.n987 GND.n986 9.3005
R30956 GND.n989 GND.n988 9.3005
R30957 GND.n8813 GND.n8812 9.3005
R30958 GND.n8817 GND.n8816 9.3005
R30959 GND.n8819 GND.n8818 9.3005
R30960 GND.n8827 GND.n8826 9.3005
R30961 GND.n8831 GND.n8830 9.3005
R30962 GND.n8833 GND.n8832 9.3005
R30963 GND.n8840 GND.n8839 9.3005
R30964 GND.n8844 GND.n8843 9.3005
R30965 GND.n8846 GND.n8845 9.3005
R30966 GND.n8853 GND.n8852 9.3005
R30967 GND.n8857 GND.n8856 9.3005
R30968 GND.n8859 GND.n8858 9.3005
R30969 GND.n8866 GND.n8865 9.3005
R30970 GND.n8870 GND.n8869 9.3005
R30971 GND.n8872 GND.n8871 9.3005
R30972 GND.n8879 GND.n8878 9.3005
R30973 GND.n8883 GND.n8882 9.3005
R30974 GND.n8885 GND.n8884 9.3005
R30975 GND.n8794 GND.n8793 9.3005
R30976 GND.n8798 GND.n8797 9.3005
R30977 GND.n8800 GND.n8799 9.3005
R30978 GND.n1440 GND.n1363 9.3005
R30979 GND.n1438 GND.n1368 9.3005
R30980 GND.n9791 GND.n9790 9.3005
R30981 GND.n9789 GND.n55 9.3005
R30982 GND.n9788 GND.n9787 9.3005
R30983 GND.n9763 GND.n9762 9.3005
R30984 GND.n9756 GND.n9755 9.3005
R30985 GND.n9755 GND.n69 9.3005
R30986 GND.n9755 GND.n9754 9.3005
R30987 GND.n9569 GND.n9564 9.3005
R30988 GND.n9570 GND.n9569 9.3005
R30989 GND.n9569 GND.n9568 9.3005
R30990 GND.n9725 GND.n9724 9.3005
R30991 GND.n9601 GND.n9600 9.3005
R30992 GND.n252 GND.n250 9.3005
R30993 GND.n9387 GND.n9386 9.3005
R30994 GND.n9385 GND.n9384 9.3005
R30995 GND.n254 GND.n253 9.3005
R30996 GND.n9372 GND.n9371 9.3005
R30997 GND.n9370 GND.n9369 9.3005
R30998 GND.n273 GND.n272 9.3005
R30999 GND.n952 GND.n473 9.3005
R31000 GND.n955 GND.n954 9.3005
R31001 GND.n958 GND.n957 9.3005
R31002 GND.n972 GND.n964 9.3005
R31003 GND.n975 GND.n974 9.3005
R31004 GND.n977 GND.n963 9.3005
R31005 GND.n961 GND.n263 9.3005
R31006 GND.n9394 GND.n9393 9.3005
R31007 GND.n242 GND.n241 9.3005
R31008 GND.n957 GND.n262 9.3005
R31009 GND.n9378 GND.n263 9.3005
R31010 GND.n977 GND.n264 9.3005
R31011 GND.n283 GND.n281 9.3005
R31012 GND.n9363 GND.n9362 9.3005
R31013 GND.n848 GND.n847 9.3005
R31014 GND.n845 GND.n462 9.3005
R31015 GND.n9018 GND.n9017 9.3005
R31016 GND.n9020 GND.n442 9.3005
R31017 GND.n8978 GND.n459 9.3005
R31018 GND.n9022 GND.n443 9.3005
R31019 GND.n9025 GND.n9024 9.3005
R31020 GND.n9411 GND.n9410 9.3005
R31021 GND.n9409 GND.n9408 9.3005
R31022 GND.n222 GND.n221 9.3005
R31023 GND.n833 GND.n832 9.3005
R31024 GND.n835 GND.n834 9.3005
R31025 GND.n836 GND.n826 9.3005
R31026 GND.n843 GND.n842 9.3005
R31027 GND.n828 GND.n825 9.3005
R31028 GND.n9294 GND.n9293 9.3005
R31029 GND.n9295 GND.n338 9.3005
R31030 GND.n219 GND.n218 9.3005
R31031 GND.n220 GND.n214 9.3005
R31032 GND.n9028 GND.n9026 9.3005
R31033 GND.n460 GND.n444 9.3005
R31034 GND.n9052 GND.n9051 9.3005
R31035 GND.n9054 GND.n440 9.3005
R31036 GND.n9056 GND.n9055 9.3005
R31037 GND.n345 GND.n344 9.3005
R31038 GND.n9285 GND.n9284 9.3005
R31039 GND.n9287 GND.n9286 9.3005
R31040 GND.n341 GND.n340 9.3005
R31041 GND.n747 GND.n525 9.3005
R31042 GND.n749 GND.n748 9.3005
R31043 GND.n489 GND.n488 9.3005
R31044 GND.n931 GND.n930 9.3005
R31045 GND.n933 GND.n932 9.3005
R31046 GND.n934 GND.n482 9.3005
R31047 GND.n941 GND.n940 9.3005
R31048 GND.n746 GND.n745 9.3005
R31049 GND.n742 GND.n527 9.3005
R31050 GND.n430 GND.n429 9.3005
R31051 GND.n9079 GND.n9078 9.3005
R31052 GND.n9073 GND.n9072 9.3005
R31053 GND.n9071 GND.n9070 9.3005
R31054 GND.n9067 GND.n433 9.3005
R31055 GND.n9065 GND.n9064 9.3005
R31056 GND.n9063 GND.n9062 9.3005
R31057 GND.n436 GND.n435 9.3005
R31058 GND.n9035 GND.n453 9.3005
R31059 GND.n485 GND.n470 9.3005
R31060 GND.n9038 GND.n9037 9.3005
R31061 GND.n8969 GND.n455 9.3005
R31062 GND.n207 GND.n206 9.3005
R31063 GND.n914 GND.n912 9.3005
R31064 GND.n919 GND.n918 9.3005
R31065 GND.n920 GND.n910 9.3005
R31066 GND.n922 GND.n921 9.3005
R31067 GND.n481 GND.n479 9.3005
R31068 GND.n945 GND.n944 9.3005
R31069 GND.n942 GND.n468 9.3005
R31070 GND.n8971 GND.n8970 9.3005
R31071 GND.n9306 GND.n9305 9.3005
R31072 GND.n9304 GND.n9303 9.3005
R31073 GND.n331 GND.n330 9.3005
R31074 GND.n9239 GND.n375 9.3005
R31075 GND.n205 GND.n203 9.3005
R31076 GND.n9421 GND.n9420 9.3005
R31077 GND.n9419 GND.n9418 9.3005
R31078 GND.n888 GND.n454 9.3005
R31079 GND.n9039 GND.n451 9.3005
R31080 GND.n9042 GND.n9041 9.3005
R31081 GND.n356 GND.n355 9.3005
R31082 GND.n9273 GND.n9272 9.3005
R31083 GND.n9274 GND.n353 9.3005
R31084 GND.n9276 GND.n9275 9.3005
R31085 GND.n329 GND.n327 9.3005
R31086 GND.n9255 GND.n9254 9.3005
R31087 GND.n9251 GND.n366 9.3005
R31088 GND.n9249 GND.n9248 9.3005
R31089 GND.n9247 GND.n9246 9.3005
R31090 GND.n9257 GND.n9256 9.3005
R31091 GND.n9260 GND.n364 9.3005
R31092 GND.n9263 GND.n9262 9.3005
R31093 GND.n9265 GND.n9264 9.3005
R31094 GND.n363 GND.n361 9.3005
R31095 GND.n882 GND.n881 9.3005
R31096 GND.n864 GND.n863 9.3005
R31097 GND.n499 GND.n498 9.3005
R31098 GND.n871 GND.n870 9.3005
R31099 GND.n872 GND.n496 9.3005
R31100 GND.n906 GND.n905 9.3005
R31101 GND.n904 GND.n903 9.3005
R31102 GND.n901 GND.n873 9.3005
R31103 GND.n862 GND.n861 9.3005
R31104 GND.n502 GND.n501 9.3005
R31105 GND.n720 GND.n719 9.3005
R31106 GND.n898 GND.n897 9.3005
R31107 GND.n896 GND.n895 9.3005
R31108 GND.n884 GND.n883 9.3005
R31109 GND.n879 GND.n877 9.3005
R31110 GND.n8513 GND.n8512 9.3005
R31111 GND.n8516 GND.n999 9.3005
R31112 GND.n3487 GND.n3410 9.3005
R31113 GND.n3485 GND.n3415 9.3005
R31114 GND.n4852 GND.n4851 9.3005
R31115 GND.n4856 GND.n4855 9.3005
R31116 GND.n4858 GND.n4857 9.3005
R31117 GND.n4838 GND.n4837 9.3005
R31118 GND.n4842 GND.n4841 9.3005
R31119 GND.n4844 GND.n4843 9.3005
R31120 GND.n4824 GND.n4823 9.3005
R31121 GND.n4828 GND.n4827 9.3005
R31122 GND.n4830 GND.n4829 9.3005
R31123 GND.n4810 GND.n4809 9.3005
R31124 GND.n4814 GND.n4813 9.3005
R31125 GND.n4816 GND.n4815 9.3005
R31126 GND.n4796 GND.n4795 9.3005
R31127 GND.n4800 GND.n4799 9.3005
R31128 GND.n4802 GND.n4801 9.3005
R31129 GND.n4781 GND.n4780 9.3005
R31130 GND.n4785 GND.n4784 9.3005
R31131 GND.n4787 GND.n4786 9.3005
R31132 GND.n4175 GND.n4174 9.3005
R31133 GND.n4179 GND.n4178 9.3005
R31134 GND.n4181 GND.n4180 9.3005
R31135 GND.n4869 GND.n4868 9.3005
R31136 GND.n4873 GND.n4872 9.3005
R31137 GND.n4875 GND.n4874 9.3005
R31138 GND.n4882 GND.n4881 9.3005
R31139 GND.n4886 GND.n4885 9.3005
R31140 GND.n4888 GND.n4887 9.3005
R31141 GND.n4895 GND.n4894 9.3005
R31142 GND.n4899 GND.n4898 9.3005
R31143 GND.n4901 GND.n4900 9.3005
R31144 GND.n4908 GND.n4907 9.3005
R31145 GND.n4912 GND.n4911 9.3005
R31146 GND.n4914 GND.n4913 9.3005
R31147 GND.n4921 GND.n4920 9.3005
R31148 GND.n4925 GND.n4924 9.3005
R31149 GND.n4927 GND.n4926 9.3005
R31150 GND.n4156 GND.n4155 9.3005
R31151 GND.n4160 GND.n4159 9.3005
R31152 GND.n4162 GND.n4161 9.3005
R31153 GND.n4946 GND.n4945 9.3005
R31154 GND.n3950 GND.n3936 9.3005
R31155 GND.n7889 GND.n7888 9.3005
R31156 GND.n7974 GND.n2153 9.3005
R31157 GND.n7974 GND.n2152 9.3005
R31158 GND.n7974 GND.n7973 9.3005
R31159 GND.n7849 GND.n2151 9.3005
R31160 GND.n7851 GND.n2151 9.3005
R31161 GND.n7852 GND.n2151 9.3005
R31162 GND.n7946 GND.n7945 9.3005
R31163 GND.n2244 GND.n2243 9.3005
R31164 GND.n1944 GND.n1942 9.3005
R31165 GND.n8281 GND.n8280 9.3005
R31166 GND.n8279 GND.n8278 9.3005
R31167 GND.n1946 GND.n1945 9.3005
R31168 GND.n8266 GND.n8265 9.3005
R31169 GND.n8264 GND.n8263 9.3005
R31170 GND.n1965 GND.n1964 9.3005
R31171 GND.n4686 GND.n4212 9.3005
R31172 GND.n4689 GND.n4688 9.3005
R31173 GND.n4692 GND.n4691 9.3005
R31174 GND.n4704 GND.n4697 9.3005
R31175 GND.n4707 GND.n4706 9.3005
R31176 GND.n4710 GND.n4709 9.3005
R31177 GND.n4712 GND.n1955 9.3005
R31178 GND.n8288 GND.n8287 9.3005
R31179 GND.n1934 GND.n1933 9.3005
R31180 GND.n4691 GND.n1954 9.3005
R31181 GND.n8272 GND.n1955 9.3005
R31182 GND.n4709 GND.n1956 9.3005
R31183 GND.n1975 GND.n1973 9.3005
R31184 GND.n8257 GND.n8256 9.3005
R31185 GND.n4498 GND.n4497 9.3005
R31186 GND.n4495 GND.n4256 9.3005
R31187 GND.n4762 GND.n4203 9.3005
R31188 GND.n4765 GND.n4764 9.3005
R31189 GND.n4257 GND.n4206 9.3005
R31190 GND.n4723 GND.n4201 9.3005
R31191 GND.n4721 GND.n4720 9.3005
R31192 GND.n8305 GND.n8304 9.3005
R31193 GND.n8303 GND.n8302 9.3005
R31194 GND.n1914 GND.n1913 9.3005
R31195 GND.n4476 GND.n4475 9.3005
R31196 GND.n4473 GND.n4472 9.3005
R31197 GND.n4483 GND.n4482 9.3005
R31198 GND.n4484 GND.n4471 9.3005
R31199 GND.n4487 GND.n4486 9.3005
R31200 GND.n8188 GND.n8187 9.3005
R31201 GND.n8189 GND.n2030 9.3005
R31202 GND.n4341 GND.n4340 9.3005
R31203 GND.n1912 GND.n1910 9.3005
R31204 GND.n4717 GND.n4716 9.3005
R31205 GND.n4718 GND.n4199 9.3005
R31206 GND.n4768 GND.n4767 9.3005
R31207 GND.n4641 GND.n4202 9.3005
R31208 GND.n4644 GND.n4643 9.3005
R31209 GND.n2037 GND.n2036 9.3005
R31210 GND.n8179 GND.n8178 9.3005
R31211 GND.n8181 GND.n8180 9.3005
R31212 GND.n2033 GND.n2032 9.3005
R31213 GND.n4264 GND.n4263 9.3005
R31214 GND.n4453 GND.n4452 9.3005
R31215 GND.n4455 GND.n4454 9.3005
R31216 GND.n4457 GND.n4261 9.3005
R31217 GND.n4462 GND.n4461 9.3005
R31218 GND.n4464 GND.n4463 9.3005
R31219 GND.n4466 GND.n4222 9.3005
R31220 GND.n4354 GND.n4353 9.3005
R31221 GND.n4352 GND.n4272 9.3005
R31222 GND.n4628 GND.n4627 9.3005
R31223 GND.n4624 GND.n4557 9.3005
R31224 GND.n4630 GND.n4629 9.3005
R31225 GND.n4554 GND.n4553 9.3005
R31226 GND.n4636 GND.n4635 9.3005
R31227 GND.n4638 GND.n4637 9.3005
R31228 GND.n4552 GND.n4550 9.3005
R31229 GND.n4650 GND.n4549 9.3005
R31230 GND.n4653 GND.n4652 9.3005
R31231 GND.n4467 GND.n4223 9.3005
R31232 GND.n4654 GND.n4193 9.3005
R31233 GND.n4776 GND.n4775 9.3005
R31234 GND.n1903 GND.n1902 9.3005
R31235 GND.n4511 GND.n4509 9.3005
R31236 GND.n4516 GND.n4515 9.3005
R31237 GND.n4517 GND.n4507 9.3005
R31238 GND.n4519 GND.n4518 9.3005
R31239 GND.n4221 GND.n4219 9.3005
R31240 GND.n4679 GND.n4678 9.3005
R31241 GND.n4676 GND.n4675 9.3005
R31242 GND.n4224 GND.n4189 9.3005
R31243 GND.n8200 GND.n8199 9.3005
R31244 GND.n8198 GND.n8197 9.3005
R31245 GND.n2023 GND.n2022 9.3005
R31246 GND.n8133 GND.n2067 9.3005
R31247 GND.n1901 GND.n1899 9.3005
R31248 GND.n8315 GND.n8314 9.3005
R31249 GND.n8313 GND.n8312 9.3005
R31250 GND.n4545 GND.n4190 9.3005
R31251 GND.n4655 GND.n4547 9.3005
R31252 GND.n4658 GND.n4657 9.3005
R31253 GND.n2048 GND.n2047 9.3005
R31254 GND.n8167 GND.n8166 9.3005
R31255 GND.n8168 GND.n2045 9.3005
R31256 GND.n8170 GND.n8169 9.3005
R31257 GND.n2021 GND.n2019 9.3005
R31258 GND.n8149 GND.n8148 9.3005
R31259 GND.n8145 GND.n2058 9.3005
R31260 GND.n8143 GND.n8142 9.3005
R31261 GND.n8141 GND.n8140 9.3005
R31262 GND.n8151 GND.n8150 9.3005
R31263 GND.n8154 GND.n2056 9.3005
R31264 GND.n8157 GND.n8156 9.3005
R31265 GND.n8159 GND.n8158 9.3005
R31266 GND.n2055 GND.n2053 9.3005
R31267 GND.n4539 GND.n4538 9.3005
R31268 GND.n4241 GND.n4240 9.3005
R31269 GND.n4235 GND.n4234 9.3005
R31270 GND.n4247 GND.n4246 9.3005
R31271 GND.n4250 GND.n4249 9.3005
R31272 GND.n4248 GND.n4231 9.3005
R31273 GND.n4527 GND.n4230 9.3005
R31274 GND.n4531 GND.n4530 9.3005
R31275 GND.n4239 GND.n4238 9.3005
R31276 GND.n1893 GND.n1892 9.3005
R31277 GND.n8322 GND.n8321 9.3005
R31278 GND.n4532 GND.n4228 9.3005
R31279 GND.n4669 GND.n4668 9.3005
R31280 GND.n4535 GND.n4533 9.3005
R31281 GND.n4666 GND.n4665 9.3005
R31282 GND.n9446 GND.n9445 9.3005
R31283 GND.n9448 GND.n9447 9.3005
R31284 GND.n9444 GND.n9 9.3005
R31285 GND.n9457 GND.n9456 9.3005
R31286 GND.n9459 GND.n9458 9.3005
R31287 GND.n9455 GND.n9437 9.3005
R31288 GND.n9824 GND.n9823 9.3005
R31289 GND.n8427 GND.n8426 9.3005
R31290 GND.n8425 GND.n1804 9.3005
R31291 GND.n8424 GND.n8423 9.3005
R31292 GND.n6616 GND.n6615 9.3005
R31293 GND.n7223 GND.n7222 9.3005
R31294 GND.n7225 GND.n7224 9.3005
R31295 GND.n2553 GND.n2552 9.3005
R31296 GND.n7314 GND.n7313 9.3005
R31297 GND.n7315 GND.n2550 9.3005
R31298 GND.n7317 GND.n7316 9.3005
R31299 GND.n7076 GND.n7075 9.3005
R31300 GND.n6628 GND.n6627 9.3005
R31301 GND.n7300 GND.n2566 9.3005
R31302 GND.n7303 GND.n7302 9.3005
R31303 GND.n7213 GND.n7205 9.3005
R31304 GND.n7305 GND.n2564 9.3005
R31305 GND.n7210 GND.n7209 9.3005
R31306 GND.n6626 GND.n6624 9.3005
R31307 GND.n7216 GND.n7215 9.3005
R31308 GND.n7213 GND.n7212 9.3005
R31309 GND.n7210 GND.n2561 9.3005
R31310 GND.n7306 GND.n7305 9.3005
R31311 GND.n7289 GND.n2565 9.3005
R31312 GND.n7293 GND.n7291 9.3005
R31313 GND.n7118 GND.n6641 9.3005
R31314 GND.n7183 GND.n7182 9.3005
R31315 GND.n7324 GND.n7323 9.3005
R31316 GND.n2542 GND.n2541 9.3005
R31317 GND.n7186 GND.n7185 9.3005
R31318 GND.n7235 GND.n7234 9.3005
R31319 GND.n7231 GND.n6607 9.3005
R31320 GND.n6669 GND.n6668 9.3005
R31321 GND.n7146 GND.n7145 9.3005
R31322 GND.n7147 GND.n6666 9.3005
R31323 GND.n7151 GND.n7150 9.3005
R31324 GND.n7149 GND.n7148 9.3005
R31325 GND.n6646 GND.n6642 9.3005
R31326 GND.n7180 GND.n7179 9.3005
R31327 GND.n6644 GND.n6639 9.3005
R31328 GND.n2485 GND.n2484 9.3005
R31329 GND.n7424 GND.n7423 9.3005
R31330 GND.n7009 GND.n7008 9.3005
R31331 GND.n7007 GND.n7006 9.3005
R31332 GND.n7189 GND.n7187 9.3005
R31333 GND.n2694 GND.n2692 9.3005
R31334 GND.n7241 GND.n7240 9.3005
R31335 GND.n7238 GND.n7237 9.3005
R31336 GND.n2513 GND.n2512 9.3005
R31337 GND.n7380 GND.n7379 9.3005
R31338 GND.n7381 GND.n2510 9.3005
R31339 GND.n7386 GND.n7385 9.3005
R31340 GND.n7384 GND.n7383 9.3005
R31341 GND.n6932 GND.n6931 9.3005
R31342 GND.n6930 GND.n6929 9.3005
R31343 GND.n6660 GND.n6659 9.3005
R31344 GND.n7158 GND.n7157 9.3005
R31345 GND.n7160 GND.n7159 9.3005
R31346 GND.n7162 GND.n6657 9.3005
R31347 GND.n7166 GND.n7165 9.3005
R31348 GND.n7196 GND.n7195 9.3005
R31349 GND.n2667 GND.n2666 9.3005
R31350 GND.n2665 GND.n2664 9.3005
R31351 GND.n2646 GND.n2645 9.3005
R31352 GND.n2674 GND.n2673 9.3005
R31353 GND.n2676 GND.n2675 9.3005
R31354 GND.n2680 GND.n2643 9.3005
R31355 GND.n2683 GND.n2682 9.3005
R31356 GND.n2685 GND.n2684 9.3005
R31357 GND.n2642 GND.n2638 9.3005
R31358 GND.n7248 GND.n7247 9.3005
R31359 GND.n6635 GND.n2635 9.3005
R31360 GND.n6926 GND.n6925 9.3005
R31361 GND.n6939 GND.n6938 9.3005
R31362 GND.n7059 GND.n7058 9.3005
R31363 GND.n7057 GND.n7056 9.3005
R31364 GND.n6738 GND.n6737 9.3005
R31365 GND.n7051 GND.n7050 9.3005
R31366 GND.n7049 GND.n7048 9.3005
R31367 GND.n6656 GND.n6654 9.3005
R31368 GND.n7169 GND.n7168 9.3005
R31369 GND.n6633 GND.n6632 9.3005
R31370 GND.n7198 GND.n7197 9.3005
R31371 GND.n7401 GND.n7400 9.3005
R31372 GND.n7399 GND.n7398 9.3005
R31373 GND.n2476 GND.n2475 9.3005
R31374 GND.n7433 GND.n7432 9.3005
R31375 GND.n6995 GND.n6994 9.3005
R31376 GND.n6993 GND.n6992 9.3005
R31377 GND.n6736 GND.n6734 9.3005
R31378 GND.n7250 GND.n7249 9.3005
R31379 GND.n2636 GND.n2623 9.3005
R31380 GND.n7282 GND.n7281 9.3005
R31381 GND.n7283 GND.n2620 9.3005
R31382 GND.n7285 GND.n7284 9.3005
R31383 GND.n2503 GND.n2502 9.3005
R31384 GND.n7395 GND.n7394 9.3005
R31385 GND.n7396 GND.n2500 9.3005
R31386 GND.n7409 GND.n7408 9.3005
R31387 GND.n7410 GND.n2490 9.3005
R31388 GND.n7416 GND.n7415 9.3005
R31389 GND.n7414 GND.n7413 9.3005
R31390 GND.n2493 GND.n2492 9.3005
R31391 GND.n7264 GND.n7263 9.3005
R31392 GND.n7266 GND.n7265 9.3005
R31393 GND.n7269 GND.n7260 9.3005
R31394 GND.n7272 GND.n7271 9.3005
R31395 GND.n7274 GND.n7273 9.3005
R31396 GND.n7019 GND.n7018 9.3005
R31397 GND.n6744 GND.n6743 9.3005
R31398 GND.n7026 GND.n7025 9.3005
R31399 GND.n7027 GND.n6741 9.3005
R31400 GND.n7041 GND.n7040 9.3005
R31401 GND.n7039 GND.n7038 9.3005
R31402 GND.n7036 GND.n7028 9.3005
R31403 GND.n7017 GND.n7016 9.3005
R31404 GND.n6747 GND.n6746 9.3005
R31405 GND.n6978 GND.n6977 9.3005
R31406 GND.n7033 GND.n7032 9.3005
R31407 GND.n7031 GND.n7030 9.3005
R31408 GND.n7259 GND.n2627 9.3005
R31409 GND.n7258 GND.n7257 9.3005
R31410 GND.n5483 GND.n5468 9.2805
R31411 GND.n5526 GND.n5488 9.2805
R31412 GND.n9724 GND.n100 9.2805
R31413 GND.n9600 GND.n135 9.2805
R31414 GND.n7945 GND.n2183 9.2805
R31415 GND.n2244 GND.n2229 9.2805
R31416 GND.t41 GND.n247 9.18083
R31417 GND.t305 GND.n1939 9.18083
R31418 GND.t300 GND.n6621 9.18083
R31419 GND.t87 GND.n2365 9.05485
R31420 GND.n9427 GND.n195 9.03579
R31421 GND.n831 GND.n222 9.03579
R31422 GND.n9284 GND.n9283 9.03579
R31423 GND.n9296 GND.n339 9.03579
R31424 GND.n739 GND.n738 9.03579
R31425 GND.n929 GND.n489 9.03579
R31426 GND.n9067 GND.n9066 9.03579
R31427 GND.n9081 GND.n9080 9.03579
R31428 GND.n4343 GND.n4342 9.03579
R31429 GND.n4474 GND.n1914 9.03579
R31430 GND.n8178 GND.n8177 9.03579
R31431 GND.n8190 GND.n2031 9.03579
R31432 GND.n4351 GND.n4349 9.03579
R31433 GND.n4456 GND.n4455 9.03579
R31434 GND.n4635 GND.n4551 9.03579
R31435 GND.n4622 GND.n4621 9.03579
R31436 GND.n7003 GND.n7002 9.03579
R31437 GND.n7152 GND.n6666 9.03579
R31438 GND.n7378 GND.n2510 9.03579
R31439 GND.n7426 GND.n7425 9.03579
R31440 GND.n6942 GND.n6940 9.03579
R31441 GND.n7156 GND.n6660 9.03579
R31442 GND.n2679 GND.n2676 9.03579
R31443 GND.n2661 GND.n2660 9.03579
R31444 GND.t160 GND.n5660 8.84906
R31445 GND.n3088 GND.n2900 8.8069
R31446 GND.n7553 GND.n7552 8.79143
R31447 GND.n8058 GND.n2108 8.78859
R31448 GND.n6232 GND.n2793 8.65932
R31449 GND.n6233 GND.n6232 8.65932
R31450 GND.n1751 GND.n1749 8.65932
R31451 GND.n8629 GND.n1749 8.65932
R31452 GND.n5814 GND.n5813 8.65932
R31453 GND.n5813 GND.n5812 8.65932
R31454 GND.n5435 GND.n5027 8.5765
R31455 GND.n1463 GND.n1362 8.5765
R31456 GND.n3506 GND.n3409 8.5765
R31457 GND.t306 GND.n925 8.52509
R31458 GND.n4522 GND.t35 8.52509
R31459 GND.n7044 GND.t118 8.52509
R31460 GND.n9688 GND.n121 8.48875
R31461 GND.n7987 GND.n7986 8.48875
R31462 GND.n6355 GND.n6327 8.3205
R31463 GND.n8532 GND.n8511 8.3205
R31464 GND.n4947 GND.n3928 8.3205
R31465 GND.n6591 GND.n6590 8.28285
R31466 GND.n6577 GND.n6576 8.28285
R31467 GND.n6563 GND.n6562 8.28285
R31468 GND.n6549 GND.n6548 8.28285
R31469 GND.n6535 GND.n6534 8.28285
R31470 GND.n2701 GND.n2700 8.28285
R31471 GND.n6450 GND.n6449 8.28285
R31472 GND.n6464 GND.n6463 8.28285
R31473 GND.n6477 GND.n6476 8.28285
R31474 GND.n6490 GND.n6489 8.28285
R31475 GND.n6503 GND.n6502 8.28285
R31476 GND.n6516 GND.n6515 8.28285
R31477 GND.n6431 GND.n6430 8.28285
R31478 GND.n8954 GND.n8953 8.28285
R31479 GND.n8940 GND.n8939 8.28285
R31480 GND.n8926 GND.n8925 8.28285
R31481 GND.n8912 GND.n8911 8.28285
R31482 GND.n8898 GND.n8897 8.28285
R31483 GND.n984 GND.n983 8.28285
R31484 GND.n8814 GND.n8813 8.28285
R31485 GND.n8828 GND.n8827 8.28285
R31486 GND.n8841 GND.n8840 8.28285
R31487 GND.n8854 GND.n8853 8.28285
R31488 GND.n8867 GND.n8866 8.28285
R31489 GND.n8880 GND.n8879 8.28285
R31490 GND.n8795 GND.n8794 8.28285
R31491 GND.n535 GND.n203 8.28285
R31492 GND.n923 GND.n910 8.28285
R31493 GND.n9271 GND.n353 8.28285
R31494 GND.n9241 GND.n375 8.28285
R31495 GND.n719 GND.n717 8.28285
R31496 GND.n907 GND.n496 8.28285
R31497 GND.n9262 GND.n362 8.28285
R31498 GND.n9246 GND.n9245 8.28285
R31499 GND.n4853 GND.n4852 8.28285
R31500 GND.n4839 GND.n4838 8.28285
R31501 GND.n4825 GND.n4824 8.28285
R31502 GND.n4811 GND.n4810 8.28285
R31503 GND.n4797 GND.n4796 8.28285
R31504 GND.n4782 GND.n4781 8.28285
R31505 GND.n4176 GND.n4175 8.28285
R31506 GND.n4870 GND.n4869 8.28285
R31507 GND.n4883 GND.n4882 8.28285
R31508 GND.n4896 GND.n4895 8.28285
R31509 GND.n4909 GND.n4908 8.28285
R31510 GND.n4922 GND.n4921 8.28285
R31511 GND.n4157 GND.n4156 8.28285
R31512 GND.n1899 GND.n1898 8.28285
R31513 GND.n4520 GND.n4507 8.28285
R31514 GND.n8165 GND.n2045 8.28285
R31515 GND.n8135 GND.n2067 8.28285
R31516 GND.n8321 GND.n1891 8.28285
R31517 GND.n4251 GND.n4250 8.28285
R31518 GND.n8156 GND.n2054 8.28285
R31519 GND.n8140 GND.n8139 8.28285
R31520 GND.n6996 GND.n6995 8.28285
R31521 GND.n7051 GND.n7046 8.28285
R31522 GND.n2621 GND.n2503 8.28285
R31523 GND.n7432 GND.n2474 8.28285
R31524 GND.n6977 GND.n6975 8.28285
R31525 GND.n7042 GND.n6741 8.28285
R31526 GND.n7268 GND.n7266 8.28285
R31527 GND.n7413 GND.n7412 8.28285
R31528 GND.n5628 GND.n5552 8.09988
R31529 GND.n9605 GND.n131 8.09988
R31530 GND.n7978 GND.n2147 8.09988
R31531 GND.n5628 GND.n5627 8.0985
R31532 GND.n9606 GND.n9605 8.0985
R31533 GND.n7979 GND.n7978 8.0985
R31534 GND.n7500 GND.t22 8.08248
R31535 GND.t194 GND.n8100 8.07988
R31536 GND.n632 GND.t250 8.07988
R31537 GND.n8360 GND.t276 8.07988
R31538 GND.n5026 GND.n5025 8.0645
R31539 GND.n1442 GND.n1440 8.0645
R31540 GND.n3489 GND.n3487 8.0645
R31541 GND.n9560 GND.t246 8.02575
R31542 GND.n9638 GND.t261 8.02575
R31543 GND.n7839 GND.t86 8.02575
R31544 GND.n7911 GND.t281 8.02575
R31545 GND.n5655 GND.n5654 8.0005
R31546 GND.n5484 GND.n5482 8.0005
R31547 GND.n5497 GND.n5486 8.0005
R31548 GND.n9571 GND.n9564 8.0005
R31549 GND.n9728 GND.n9726 8.0005
R31550 GND.n146 GND.n133 8.0005
R31551 GND.n7850 GND.n7849 8.0005
R31552 GND.n7949 GND.n7947 8.0005
R31553 GND.n2241 GND.n2240 8.0005
R31554 GND.n5630 GND.n5528 7.94599
R31555 GND.n9603 GND.n9602 7.94599
R31556 GND.n2242 GND.n2149 7.94599
R31557 GND.n5631 GND.n5630 7.9455
R31558 GND.n9603 GND.n101 7.9455
R31559 GND.n2184 GND.n2149 7.9455
R31560 GND.n6601 GND.n6588 7.9105
R31561 GND.n6587 GND.n6574 7.9105
R31562 GND.n6573 GND.n6560 7.9105
R31563 GND.n6559 GND.n6546 7.9105
R31564 GND.n6545 GND.n6532 7.9105
R31565 GND.n2711 GND.n2698 7.9105
R31566 GND.n2711 GND.n2710 7.9105
R31567 GND.n6545 GND.n6544 7.9105
R31568 GND.n6559 GND.n6558 7.9105
R31569 GND.n6573 GND.n6572 7.9105
R31570 GND.n6587 GND.n6586 7.9105
R31571 GND.n6601 GND.n6600 7.9105
R31572 GND.n6460 GND.n6447 7.9105
R31573 GND.n6474 GND.n6446 7.9105
R31574 GND.n6487 GND.n6445 7.9105
R31575 GND.n6500 GND.n6444 7.9105
R31576 GND.n6513 GND.n6443 7.9105
R31577 GND.n6526 GND.n6442 7.9105
R31578 GND.n6441 GND.n6428 7.9105
R31579 GND.n6441 GND.n6440 7.9105
R31580 GND.n6526 GND.n6525 7.9105
R31581 GND.n6513 GND.n6512 7.9105
R31582 GND.n6500 GND.n6499 7.9105
R31583 GND.n6487 GND.n6486 7.9105
R31584 GND.n6474 GND.n6473 7.9105
R31585 GND.n6460 GND.n6459 7.9105
R31586 GND.n8964 GND.n8951 7.9105
R31587 GND.n8950 GND.n8937 7.9105
R31588 GND.n8936 GND.n8923 7.9105
R31589 GND.n8922 GND.n8909 7.9105
R31590 GND.n8908 GND.n8895 7.9105
R31591 GND.n994 GND.n981 7.9105
R31592 GND.n994 GND.n993 7.9105
R31593 GND.n8908 GND.n8907 7.9105
R31594 GND.n8922 GND.n8921 7.9105
R31595 GND.n8936 GND.n8935 7.9105
R31596 GND.n8950 GND.n8949 7.9105
R31597 GND.n8964 GND.n8963 7.9105
R31598 GND.n8824 GND.n8811 7.9105
R31599 GND.n8838 GND.n8810 7.9105
R31600 GND.n8851 GND.n8809 7.9105
R31601 GND.n8864 GND.n8808 7.9105
R31602 GND.n8877 GND.n8807 7.9105
R31603 GND.n8890 GND.n8806 7.9105
R31604 GND.n8805 GND.n8792 7.9105
R31605 GND.n8805 GND.n8804 7.9105
R31606 GND.n8890 GND.n8889 7.9105
R31607 GND.n8877 GND.n8876 7.9105
R31608 GND.n8864 GND.n8863 7.9105
R31609 GND.n8851 GND.n8850 7.9105
R31610 GND.n8838 GND.n8837 7.9105
R31611 GND.n8824 GND.n8823 7.9105
R31612 GND.n4863 GND.n4850 7.9105
R31613 GND.n4849 GND.n4836 7.9105
R31614 GND.n4835 GND.n4822 7.9105
R31615 GND.n4821 GND.n4808 7.9105
R31616 GND.n4807 GND.n4794 7.9105
R31617 GND.n4792 GND.n4779 7.9105
R31618 GND.n4792 GND.n4791 7.9105
R31619 GND.n4807 GND.n4806 7.9105
R31620 GND.n4821 GND.n4820 7.9105
R31621 GND.n4835 GND.n4834 7.9105
R31622 GND.n4849 GND.n4848 7.9105
R31623 GND.n4863 GND.n4862 7.9105
R31624 GND.n4186 GND.n4173 7.9105
R31625 GND.n4880 GND.n4172 7.9105
R31626 GND.n4893 GND.n4171 7.9105
R31627 GND.n4906 GND.n4170 7.9105
R31628 GND.n4919 GND.n4169 7.9105
R31629 GND.n4932 GND.n4168 7.9105
R31630 GND.n4167 GND.n4154 7.9105
R31631 GND.n4167 GND.n4166 7.9105
R31632 GND.n4932 GND.n4931 7.9105
R31633 GND.n4919 GND.n4918 7.9105
R31634 GND.n4906 GND.n4905 7.9105
R31635 GND.n4893 GND.n4892 7.9105
R31636 GND.n4880 GND.n4879 7.9105
R31637 GND.n4186 GND.n4185 7.9105
R31638 GND.n5340 GND.n5339 7.90638
R31639 GND.n5339 GND.n5036 7.90638
R31640 GND.n1255 GND.n1241 7.90638
R31641 GND.n1243 GND.n1241 7.90638
R31642 GND.n3301 GND.n3287 7.90638
R31643 GND.n3289 GND.n3287 7.90638
R31644 GND.n9268 GND.t2 7.86935
R31645 GND.n8162 GND.t415 7.86935
R31646 GND.n7288 GND.t74 7.86935
R31647 GND.t126 GND.n2359 7.82016
R31648 GND.t190 GND.n7611 7.82016
R31649 GND.n7582 GND.n7581 7.82016
R31650 GND.n6330 GND.n6329 7.8085
R31651 GND.n8515 GND.n8513 7.8085
R31652 GND.n4946 GND.n3929 7.8085
R31653 GND.n2955 GND.n2954 7.7829
R31654 GND.n9541 GND.n9540 7.56276
R31655 GND.n7818 GND.n7817 7.56276
R31656 GND.n3040 GND.n3037 7.52991
R31657 GND.n832 GND.n830 7.52991
R31658 GND.n441 GND.n345 7.52991
R31659 GND.n930 GND.n487 7.52991
R31660 GND.n9065 GND.n434 7.52991
R31661 GND.n4477 GND.n4476 7.52991
R31662 GND.n4642 GND.n2037 7.52991
R31663 GND.n4460 GND.n4457 7.52991
R31664 GND.n4639 GND.n4638 7.52991
R31665 GND.n7151 GND.n6667 7.52991
R31666 GND.n7379 GND.n7377 7.52991
R31667 GND.n7157 GND.n6658 7.52991
R31668 GND.n2681 GND.n2680 7.52991
R31669 GND.n3037 GND.n2907 7.3733
R31670 GND.t334 GND.t383 7.28527
R31671 GND.t321 GND.n289 7.21361
R31672 GND.t177 GND.n1981 7.21361
R31673 GND.t217 GND.n2518 7.21361
R31674 GND.n7647 GND.t18 7.20282
R31675 GND.n5008 GND.n5005 7.0405
R31676 GND.n5444 GND.n5442 7.0405
R31677 GND.n5456 GND.n5455 7.0405
R31678 GND.n1451 GND.n1439 7.0405
R31679 GND.n62 GND.n60 7.0405
R31680 GND.n9754 GND.n9753 7.0405
R31681 GND.n3498 GND.n3486 7.0405
R31682 GND.n7887 GND.n7886 7.0405
R31683 GND.n7973 GND.n7972 7.0405
R31684 GND.n5140 GND.n5047 6.9637
R31685 GND.n5140 GND.n5045 6.9637
R31686 GND.n5146 GND.n5045 6.9637
R31687 GND.n5146 GND.n5043 6.9637
R31688 GND.n5152 GND.n5043 6.9637
R31689 GND.n5152 GND.n5041 6.9637
R31690 GND.n5159 GND.n5041 6.9637
R31691 GND.n5159 GND.n5037 6.9637
R31692 GND.n5338 GND.n5037 6.9637
R31693 GND.n6231 GND.n2796 6.9637
R31694 GND.n6226 GND.n2796 6.9637
R31695 GND.n6226 GND.n6225 6.9637
R31696 GND.n6225 GND.n6224 6.9637
R31697 GND.n6224 GND.n2803 6.9637
R31698 GND.n6219 GND.n2803 6.9637
R31699 GND.n6219 GND.n6218 6.9637
R31700 GND.n6218 GND.n6217 6.9637
R31701 GND.n6217 GND.n2810 6.9637
R31702 GND.n2997 GND.n2996 6.9637
R31703 GND.n3081 GND.n2904 6.9637
R31704 GND.n1596 GND.n1595 6.9637
R31705 GND.n1595 GND.n1214 6.9637
R31706 GND.n1226 GND.n1214 6.9637
R31707 GND.n1584 GND.n1226 6.9637
R31708 GND.n1584 GND.n1583 6.9637
R31709 GND.n1583 GND.n1227 6.9637
R31710 GND.n1240 GND.n1227 6.9637
R31711 GND.n1572 GND.n1240 6.9637
R31712 GND.n1572 GND.n1571 6.9637
R31713 GND.n8645 GND.n8642 6.9637
R31714 GND.n8645 GND.n8644 6.9637
R31715 GND.n8644 GND.n1737 6.9637
R31716 GND.n8656 GND.n1737 6.9637
R31717 GND.n8659 GND.n8656 6.9637
R31718 GND.n8659 GND.n8658 6.9637
R31719 GND.n8658 GND.n1724 6.9637
R31720 GND.n8669 GND.n1724 6.9637
R31721 GND.n8670 GND.n8669 6.9637
R31722 GND.n3639 GND.n3638 6.9637
R31723 GND.n3638 GND.n3260 6.9637
R31724 GND.n3272 GND.n3260 6.9637
R31725 GND.n3627 GND.n3272 6.9637
R31726 GND.n3627 GND.n3626 6.9637
R31727 GND.n3626 GND.n3273 6.9637
R31728 GND.n3286 GND.n3273 6.9637
R31729 GND.n3615 GND.n3286 6.9637
R31730 GND.n3615 GND.n3614 6.9637
R31731 GND.n4019 GND.n3814 6.9637
R31732 GND.n4020 GND.n4019 6.9637
R31733 GND.n4025 GND.n4020 6.9637
R31734 GND.n4026 GND.n4025 6.9637
R31735 GND.n4031 GND.n4026 6.9637
R31736 GND.n4032 GND.n4031 6.9637
R31737 GND.n4037 GND.n4032 6.9637
R31738 GND.n4038 GND.n4037 6.9637
R31739 GND.n4043 GND.n4038 6.9637
R31740 GND.t18 GND.n2316 6.79126
R31741 GND.n5514 GND.n5513 6.79126
R31742 GND.n7605 GND.n2387 6.79126
R31743 GND.n153 GND.t32 6.7911
R31744 GND.n7970 GND.t51 6.7911
R31745 GND.n6340 GND.n6338 6.7845
R31746 GND.n8519 GND.n8517 6.7845
R31747 GND.n3949 GND.n3938 6.7845
R31748 GND.n6593 GND.n6592 6.77697
R31749 GND.n6579 GND.n6578 6.77697
R31750 GND.n6565 GND.n6564 6.77697
R31751 GND.n6551 GND.n6550 6.77697
R31752 GND.n6537 GND.n6536 6.77697
R31753 GND.n2703 GND.n2702 6.77697
R31754 GND.n6452 GND.n6451 6.77697
R31755 GND.n6466 GND.n6465 6.77697
R31756 GND.n6479 GND.n6478 6.77697
R31757 GND.n6492 GND.n6491 6.77697
R31758 GND.n6505 GND.n6504 6.77697
R31759 GND.n6518 GND.n6517 6.77697
R31760 GND.n6433 GND.n6432 6.77697
R31761 GND.n2986 GND.n2964 6.77697
R31762 GND.n2940 GND.n2939 6.77697
R31763 GND.n3026 GND.n3025 6.77697
R31764 GND.n3052 GND.n3048 6.77697
R31765 GND.n8956 GND.n8955 6.77697
R31766 GND.n8942 GND.n8941 6.77697
R31767 GND.n8928 GND.n8927 6.77697
R31768 GND.n8914 GND.n8913 6.77697
R31769 GND.n8900 GND.n8899 6.77697
R31770 GND.n986 GND.n985 6.77697
R31771 GND.n8816 GND.n8815 6.77697
R31772 GND.n8830 GND.n8829 6.77697
R31773 GND.n8843 GND.n8842 6.77697
R31774 GND.n8856 GND.n8855 6.77697
R31775 GND.n8869 GND.n8868 6.77697
R31776 GND.n8882 GND.n8881 6.77697
R31777 GND.n8797 GND.n8796 6.77697
R31778 GND.n726 GND.n536 6.77697
R31779 GND.n922 GND.n911 6.77697
R31780 GND.n9272 GND.n9270 6.77697
R31781 GND.n9240 GND.n9238 6.77697
R31782 GND.n722 GND.n721 6.77697
R31783 GND.n906 GND.n497 6.77697
R31784 GND.n9266 GND.n9265 6.77697
R31785 GND.n9148 GND.n368 6.77697
R31786 GND.n4855 GND.n4854 6.77697
R31787 GND.n4841 GND.n4840 6.77697
R31788 GND.n4827 GND.n4826 6.77697
R31789 GND.n4813 GND.n4812 6.77697
R31790 GND.n4799 GND.n4798 6.77697
R31791 GND.n4784 GND.n4783 6.77697
R31792 GND.n4178 GND.n4177 6.77697
R31793 GND.n4872 GND.n4871 6.77697
R31794 GND.n4885 GND.n4884 6.77697
R31795 GND.n4898 GND.n4897 6.77697
R31796 GND.n4911 GND.n4910 6.77697
R31797 GND.n4924 GND.n4923 6.77697
R31798 GND.n4159 GND.n4158 6.77697
R31799 GND.n8328 GND.n1869 6.77697
R31800 GND.n4519 GND.n4508 6.77697
R31801 GND.n8166 GND.n8164 6.77697
R31802 GND.n8134 GND.n8132 6.77697
R31803 GND.n8324 GND.n8323 6.77697
R31804 GND.n4526 GND.n4231 6.77697
R31805 GND.n8160 GND.n8159 6.77697
R31806 GND.n8042 GND.n2060 6.77697
R31807 GND.n6989 GND.n6988 6.77697
R31808 GND.n7048 GND.n7047 6.77697
R31809 GND.n7286 GND.n7285 6.77697
R31810 GND.n7436 GND.n7434 6.77697
R31811 GND.n6980 GND.n6979 6.77697
R31812 GND.n7041 GND.n6742 6.77697
R31813 GND.n7270 GND.n7269 6.77697
R31814 GND.n7411 GND.n2471 6.77697
R31815 GND.n5658 GND.n5448 6.7205
R31816 GND.n9570 GND.n9567 6.7205
R31817 GND.n7853 GND.n7851 6.7205
R31818 GND.n9565 GND.t280 6.63677
R31819 GND.n7855 GND.t50 6.63677
R31820 GND.n5514 GND.n2348 6.58548
R31821 GND.n5606 GND.n2387 6.58548
R31822 GND.n9826 GND.n9825 6.56408
R31823 GND.t10 GND.n9045 6.55788
R31824 GND.n4661 GND.t5 6.55788
R31825 GND.n7277 GND.t52 6.55788
R31826 GND.n5693 GND.n5692 6.5285
R31827 GND.n1438 GND.n1437 6.5285
R31828 GND.n3485 GND.n3484 6.5285
R31829 GND.n1802 GND.n1800 6.42907
R31830 GND.t418 GND.n1800 6.42907
R31831 GND.n54 GND.n52 6.42907
R31832 GND.t104 GND.n52 6.42907
R31833 GND.n9786 GND.n53 6.42907
R31834 GND.t104 GND.n53 6.42907
R31835 GND.n9811 GND.n9810 6.42907
R31836 GND.n9810 GND.n9809 6.42907
R31837 GND.n9816 GND.n9815 6.42907
R31838 GND.n9817 GND.n9816 6.42907
R31839 GND.n1803 GND.n1801 6.42907
R31840 GND.t418 GND.n1801 6.42907
R31841 GND.n7744 GND.n7737 6.42907
R31842 GND.n7737 GND.n1815 6.42907
R31843 GND.n7738 GND.n7736 6.42907
R31844 GND.n7736 GND.n7735 6.42907
R31845 GND.n6337 GND.n2717 6.2725
R31846 GND.n8516 GND.n1000 6.2725
R31847 GND.n3951 GND.n3950 6.2725
R31848 GND.n5551 GND.n5550 6.2405
R31849 GND.n9549 GND.n9544 6.2405
R31850 GND.n7827 GND.n7821 6.2405
R31851 GND.n2954 GND.n2928 6.02403
R31852 GND.n3073 GND.n3037 6.02403
R31853 GND.n249 GND.n232 6.02403
R31854 GND.n292 GND.n291 6.02403
R31855 GND.n951 GND.n474 6.02403
R31856 GND.n971 GND.n969 6.02403
R31857 GND.n9395 GND.n240 6.02403
R31858 GND.n9361 GND.n282 6.02403
R31859 GND.n849 GND.n824 6.02403
R31860 GND.n9016 GND.n8982 6.02403
R31861 GND.n837 GND.n835 6.02403
R31862 GND.n9057 GND.n9056 6.02403
R31863 GND.n935 GND.n933 6.02403
R31864 GND.n9062 GND.n9061 6.02403
R31865 GND.n1941 GND.n1924 6.02403
R31866 GND.n1984 GND.n1983 6.02403
R31867 GND.n4685 GND.n4213 6.02403
R31868 GND.n4703 GND.n4701 6.02403
R31869 GND.n8289 GND.n1932 6.02403
R31870 GND.n8255 GND.n1974 6.02403
R31871 GND.n4499 GND.n4255 6.02403
R31872 GND.n4761 GND.n4759 6.02403
R31873 GND.n4480 GND.n4473 6.02403
R31874 GND.n4645 GND.n4644 6.02403
R31875 GND.n4461 GND.n4260 6.02403
R31876 GND.n4649 GND.n4550 6.02403
R31877 GND.n6681 GND.n6680 6.02403
R31878 GND.n2551 GND.n2522 6.02403
R31879 GND.n7077 GND.n7073 6.02403
R31880 GND.n7299 GND.n2616 6.02403
R31881 GND.n7130 GND.n7129 6.02403
R31882 GND.n7295 GND.n7294 6.02403
R31883 GND.n7120 GND.n7119 6.02403
R31884 GND.n7325 GND.n2540 6.02403
R31885 GND.n7148 GND.n6647 6.02403
R31886 GND.n7236 GND.n2513 6.02403
R31887 GND.n7161 GND.n7160 6.02403
R31888 GND.n2682 GND.n2641 6.02403
R31889 GND.n9345 GND.n317 5.90214
R31890 GND.n8239 GND.n2009 5.90214
R31891 GND.n7420 GND.n2487 5.90214
R31892 GND.n9588 GND.t252 5.86511
R31893 GND.n103 GND.t312 5.86511
R31894 GND.n7845 GND.t186 5.86511
R31895 GND.n2186 GND.t175 5.86511
R31896 GND.n8030 GND.n8029 5.86511
R31897 GND.n9790 GND.n9782 5.81173
R31898 GND.n5665 GND.n5664 5.7605
R31899 GND.n5452 GND.n5450 5.7605
R31900 GND.n9762 GND.n9761 5.7605
R31901 GND.n9757 GND.n69 5.7605
R31902 GND.n7888 GND.n2203 5.7605
R31903 GND.n2156 GND.n2152 5.7605
R31904 GND.n2973 GND.n2922 5.5301
R31905 GND.n5657 GND.n5449 5.4405
R31906 GND.n9568 GND.n104 5.4405
R31907 GND.n7852 GND.n2187 5.4405
R31908 GND.n9511 GND.t213 5.40211
R31909 GND.n7808 GND.t425 5.40211
R31910 GND.n946 GND.n479 5.27109
R31911 GND.n452 GND.n356 5.27109
R31912 GND.n903 GND.n902 5.27109
R31913 GND.n880 GND.n361 5.27109
R31914 GND.n4680 GND.n4219 5.27109
R31915 GND.n4548 GND.n2048 5.27109
R31916 GND.n4528 GND.n4527 5.27109
R31917 GND.n4537 GND.n2053 5.27109
R31918 GND.n7170 GND.n6654 5.27109
R31919 GND.n7280 GND.n2620 5.27109
R31920 GND.n7038 GND.n7037 5.27109
R31921 GND.n7271 GND.n2628 5.27109
R31922 GND.n494 GND.t237 5.2464
R31923 GND.n4524 GND.t11 5.2464
R31924 GND.t210 GND.n6648 5.2464
R31925 GND.n3008 GND.n3006 5.1205
R31926 GND.n7580 GND.n2420 5.10491
R31927 GND.n2653 GND.n2426 5.10491
R31928 GND.n7574 GND.n7573 5.10491
R31929 GND.n7567 GND.n2435 5.10491
R31930 GND.n7566 GND.n2438 5.10491
R31931 GND.n7512 GND.n7511 5.10491
R31932 GND.n7560 GND.n7559 5.10491
R31933 GND.n7505 GND.n2446 5.10491
R31934 GND.n7553 GND.n2452 5.10491
R31935 GND.n8129 GND.n2070 5.10326
R31936 GND.n8128 GND.n2073 5.10326
R31937 GND.n4613 GND.n2081 5.10326
R31938 GND.n8049 GND.n2084 5.10326
R31939 GND.n8115 GND.n2090 5.10326
R31940 GND.n8114 GND.n2093 5.10326
R31941 GND.n4604 GND.n2099 5.10326
R31942 GND.n8108 GND.n8107 5.10326
R31943 GND.n8058 GND.n2102 5.10326
R31944 GND.n568 GND.n559 5.10326
R31945 GND.n685 GND.n560 5.10326
R31946 GND.n695 GND.n546 5.10326
R31947 GND.n704 GND.n703 5.10326
R31948 GND.n551 GND.n549 5.10326
R31949 GND.n712 GND.n711 5.10326
R31950 GND.n730 GND.n530 5.10326
R31951 GND.n731 GND.n190 5.10326
R31952 GND.n8353 GND.n1838 5.10326
R31953 GND.n4317 GND.n1844 5.10326
R31954 GND.n1881 GND.n1847 5.10326
R31955 GND.n8340 GND.n1853 5.10326
R31956 GND.n8339 GND.n1856 5.10326
R31957 GND.n4326 GND.n1862 5.10326
R31958 GND.n8333 GND.n8332 5.10326
R31959 GND.n2271 GND.n1865 5.10326
R31960 GND.n9464 GND.t213 5.09345
R31961 GND.n9526 GND.n149 5.09345
R31962 GND.n9734 GND.n96 5.09345
R31963 GND.n7790 GND.t425 5.09345
R31964 GND.n7865 GND.n2213 5.09345
R31965 GND.n7955 GND.n2180 5.09345
R31966 GND.n2113 GND.n2112 5.05588
R31967 GND.n7438 GND.n2418 5.05559
R31968 GND.n9207 GND.t265 5.01604
R31969 GND.n6905 GND.t215 5.01604
R31970 GND.n5461 GND.t79 4.93923
R31971 GND.n7612 GND.t203 4.93923
R31972 GND.n9579 GND.n149 4.93912
R31973 GND.n9735 GND.n9734 4.93912
R31974 GND.n7866 GND.n7865 4.93912
R31975 GND.n7956 GND.n7955 4.93912
R31976 GND.n724 GND.n189 4.84085
R31977 GND.n8326 GND.n1871 4.84085
R31978 GND.n5626 GND.n5554 4.83606
R31979 GND.n5626 GND.n5625 4.83606
R31980 GND.n9607 GND.n127 4.83606
R31981 GND.n9609 GND.n9607 4.83606
R31982 GND.n7981 GND.n7980 4.83606
R31983 GND.n7980 GND.n2146 4.83606
R31984 GND.n5339 GND.n5338 4.8133
R31985 GND.n1571 GND.n1241 4.8133
R31986 GND.n3614 GND.n3287 4.8133
R31987 GND.n3000 GND.n2920 4.7109
R31988 GND.n3078 GND.n2906 4.7109
R31989 GND.n5551 GND.n5529 4.6405
R31990 GND.n9544 GND.n9542 4.6405
R31991 GND.n7821 GND.n7819 4.6405
R31992 GND.n6232 GND.n6231 4.6085
R31993 GND.n8642 GND.n1749 4.6085
R31994 GND.n5813 GND.n3814 4.6085
R31995 GND.n2653 GND.n2420 4.53775
R31996 GND.n7574 GND.n2426 4.53775
R31997 GND.n7573 GND.n2429 4.53775
R31998 GND.n7444 GND.n2435 4.53775
R31999 GND.n7567 GND.n7566 4.53775
R32000 GND.n7512 GND.n2438 4.53775
R32001 GND.n7559 GND.n2446 4.53775
R32002 GND.n7505 GND.n2452 4.53775
R32003 GND.n8129 GND.n8128 4.53629
R32004 GND.n4613 GND.n2073 4.53629
R32005 GND.n8122 GND.n2081 4.53629
R32006 GND.n8121 GND.n2084 4.53629
R32007 GND.n8049 GND.n2090 4.53629
R32008 GND.n8115 GND.n8114 4.53629
R32009 GND.n8108 GND.n2099 4.53629
R32010 GND.n8107 GND.n2102 4.53629
R32011 GND.n639 GND.n568 4.53629
R32012 GND.n685 GND.n559 4.53629
R32013 GND.n562 GND.n560 4.53629
R32014 GND.n696 GND.n695 4.53629
R32015 GND.n704 GND.n546 4.53629
R32016 GND.n703 GND.n549 4.53629
R32017 GND.n712 GND.n530 4.53629
R32018 GND.n731 GND.n730 4.53629
R32019 GND.n9431 GND.n190 4.53629
R32020 GND.n8354 GND.n8353 4.53629
R32021 GND.n4317 GND.n1838 4.53629
R32022 GND.n8347 GND.n1844 4.53629
R32023 GND.n8346 GND.n1847 4.53629
R32024 GND.n1881 GND.n1853 4.53629
R32025 GND.n8340 GND.n8339 4.53629
R32026 GND.n8333 GND.n1862 4.53629
R32027 GND.n8332 GND.n1865 4.53629
R32028 GND.n2272 GND.n2271 4.53629
R32029 GND.n5661 GND.t160 4.52767
R32030 GND.n5013 GND.n5010 4.5255
R32031 GND.n5437 GND.n5436 4.5255
R32032 GND.n5009 GND.n5006 4.5255
R32033 GND.n5690 GND.n5689 4.5255
R32034 GND.n6354 GND.n6353 4.5255
R32035 GND.n6351 GND.n6350 4.5255
R32036 GND.n6339 GND.n2714 4.5255
R32037 GND.n6424 GND.n6423 4.5255
R32038 GND.n8518 GND.n997 4.5255
R32039 GND.n8788 GND.n8787 4.5255
R32040 GND.n1443 GND.n1365 4.5255
R32041 GND.n1462 GND.n1461 4.5255
R32042 GND.n1434 GND.n1366 4.5255
R32043 GND.n1453 GND.n1452 4.5255
R32044 GND.n8531 GND.n8530 4.5255
R32045 GND.n8528 GND.n8527 4.5255
R32046 GND.n3490 GND.n3412 4.5255
R32047 GND.n3505 GND.n3504 4.5255
R32048 GND.n3481 GND.n3413 4.5255
R32049 GND.n3500 GND.n3499 4.5255
R32050 GND.n3933 GND.n3930 4.5255
R32051 GND.n4944 GND.n4943 4.5255
R32052 GND.n3937 GND.n3934 4.5255
R32053 GND.n4151 GND.n4150 4.5255
R32054 GND.n2954 GND.n2953 4.51815
R32055 GND.n9388 GND.n250 4.51815
R32056 GND.n9368 GND.n273 4.51815
R32057 GND.n953 GND.n952 4.51815
R32058 GND.n973 GND.n972 4.51815
R32059 GND.n9393 GND.n9392 4.51815
R32060 GND.n9364 GND.n9363 4.51815
R32061 GND.n847 GND.n846 4.51815
R32062 GND.n9019 GND.n9018 4.51815
R32063 GND.n836 GND.n827 4.51815
R32064 GND.n9050 GND.n440 4.51815
R32065 GND.n934 GND.n483 4.51815
R32066 GND.n9034 GND.n436 4.51815
R32067 GND.n8282 GND.n1942 4.51815
R32068 GND.n8262 GND.n1965 4.51815
R32069 GND.n4687 GND.n4686 4.51815
R32070 GND.n4705 GND.n4704 4.51815
R32071 GND.n8287 GND.n8286 4.51815
R32072 GND.n8258 GND.n8257 4.51815
R32073 GND.n4497 GND.n4496 4.51815
R32074 GND.n4763 GND.n4762 4.51815
R32075 GND.n4482 GND.n4481 4.51815
R32076 GND.n4641 GND.n4200 4.51815
R32077 GND.n4465 GND.n4464 4.51815
R32078 GND.n4651 GND.n4650 4.51815
R32079 GND.n7221 GND.n6616 4.51815
R32080 GND.n7318 GND.n7317 4.51815
R32081 GND.n7075 GND.n7074 4.51815
R32082 GND.n7301 GND.n7300 4.51815
R32083 GND.n7217 GND.n6624 4.51815
R32084 GND.n7291 GND.n7290 4.51815
R32085 GND.n7118 GND.n6640 4.51815
R32086 GND.n7323 GND.n7322 4.51815
R32087 GND.n6646 GND.n6643 4.51815
R32088 GND.n7237 GND.n2693 4.51815
R32089 GND.n7164 GND.n7162 4.51815
R32090 GND.n2686 GND.n2685 4.51815
R32091 GND.n5012 GND.n5011 4.5005
R32092 GND.n5691 GND.n5007 4.5005
R32093 GND.n6352 GND.n6328 4.5005
R32094 GND.n2716 GND.n2715 4.5005
R32095 GND.n999 GND.n998 4.5005
R32096 GND.n1364 GND.n1363 4.5005
R32097 GND.n1368 GND.n1367 4.5005
R32098 GND.n8529 GND.n8512 4.5005
R32099 GND.n3411 GND.n3410 4.5005
R32100 GND.n3415 GND.n3414 4.5005
R32101 GND.n4945 GND.n3931 4.5005
R32102 GND.n3936 GND.n3935 4.5005
R32103 GND.n5446 GND.n5443 4.4805
R32104 GND.n5451 GND.n2384 4.4805
R32105 GND.n9631 GND.n61 4.4805
R32106 GND.n9756 GND.n70 4.4805
R32107 GND.n7891 GND.n7890 4.4805
R32108 GND.n7914 GND.n2153 4.4805
R32109 GND.n5651 GND.t87 4.32189
R32110 GND.t375 GND.n3754 4.26958
R32111 GND.n3966 GND.t4 4.26958
R32112 GND.n5757 GND.t370 4.26958
R32113 GND.t62 GND.n5756 4.26958
R32114 GND.n7444 GND.t412 4.11238
R32115 GND.t171 GND.n8121 4.11106
R32116 GND.n6920 GND.t187 4.10413
R32117 GND.n379 GND.t323 4.03523
R32118 GND.n551 GND.t308 3.82757
R32119 GND.t197 GND.n1856 3.82757
R32120 GND.n945 GND.n480 3.76521
R32121 GND.n9043 GND.n9042 3.76521
R32122 GND.n901 GND.n900 3.76521
R32123 GND.n881 GND.n878 3.76521
R32124 GND.n4679 GND.n4220 3.76521
R32125 GND.n4659 GND.n4658 3.76521
R32126 GND.n4530 GND.n4529 3.76521
R32127 GND.n4540 GND.n4539 3.76521
R32128 GND.n7169 GND.n6655 3.76521
R32129 GND.n7281 GND.n7279 3.76521
R32130 GND.n7036 GND.n7035 3.76521
R32131 GND.n7275 GND.n7274 3.76521
R32132 GND.n2335 GND.t283 3.70455
R32133 GND.n9750 GND.t267 3.70446
R32134 GND.n9741 GND.t98 3.70446
R32135 GND.n7883 GND.t355 3.70446
R32136 GND.n7962 GND.t338 3.70446
R32137 GND.n379 GND.n378 3.62715
R32138 GND.n696 GND.t248 3.54409
R32139 GND.t122 GND.n8346 3.54409
R32140 GND.n6983 GND.t398 3.49733
R32141 GND.n6598 GND.t68 3.4805
R32142 GND.n6598 GND.t60 3.4805
R32143 GND.n6584 GND.t117 3.4805
R32144 GND.n6584 GND.t220 3.4805
R32145 GND.n6570 GND.t121 3.4805
R32146 GND.n6570 GND.t218 3.4805
R32147 GND.n6556 GND.t78 3.4805
R32148 GND.n6556 GND.t25 3.4805
R32149 GND.n6542 GND.t399 3.4805
R32150 GND.n6542 GND.t411 3.4805
R32151 GND.n2708 GND.t188 3.4805
R32152 GND.n2708 GND.t115 3.4805
R32153 GND.n6457 GND.t66 3.4805
R32154 GND.n6457 GND.t23 3.4805
R32155 GND.n6471 GND.t128 3.4805
R32156 GND.n6471 GND.t413 3.4805
R32157 GND.n6484 GND.t76 3.4805
R32158 GND.n6484 GND.t107 3.4805
R32159 GND.n6497 GND.t109 3.4805
R32160 GND.n6497 GND.t222 3.4805
R32161 GND.n6510 GND.t422 3.4805
R32162 GND.n6510 GND.t119 3.4805
R32163 GND.n6523 GND.t420 3.4805
R32164 GND.n6523 GND.t202 3.4805
R32165 GND.n6438 GND.t216 3.4805
R32166 GND.n6438 GND.t285 3.4805
R32167 GND.n8961 GND.t228 3.4805
R32168 GND.n8961 GND.t260 3.4805
R32169 GND.n8947 GND.t232 3.4805
R32170 GND.n8947 GND.t241 3.4805
R32171 GND.n8933 GND.t326 3.4805
R32172 GND.n8933 GND.t322 3.4805
R32173 GND.n8919 GND.t258 3.4805
R32174 GND.n8919 GND.t328 3.4805
R32175 GND.n8905 GND.t209 3.4805
R32176 GND.n8905 GND.t256 3.4805
R32177 GND.n991 GND.t320 3.4805
R32178 GND.n991 GND.t309 3.4805
R32179 GND.n8821 GND.t230 3.4805
R32180 GND.n8821 GND.t266 3.4805
R32181 GND.n8835 GND.t324 3.4805
R32182 GND.n8835 GND.t236 3.4805
R32183 GND.n8848 GND.t245 3.4805
R32184 GND.n8848 GND.t234 3.4805
R32185 GND.n8861 GND.t207 3.4805
R32186 GND.n8861 GND.t254 3.4805
R32187 GND.n8874 GND.t100 3.4805
R32188 GND.n8874 GND.t307 3.4805
R32189 GND.n8887 GND.t243 3.4805
R32190 GND.n8887 GND.t226 3.4805
R32191 GND.n8802 GND.t251 3.4805
R32192 GND.n8802 GND.t249 3.4805
R32193 GND.n4860 GND.t174 3.4805
R32194 GND.n4860 GND.t275 3.4805
R32195 GND.n4846 GND.t34 3.4805
R32196 GND.n4846 GND.t302 3.4805
R32197 GND.n4832 GND.t165 3.4805
R32198 GND.n4832 GND.t178 3.4805
R32199 GND.n4818 GND.t429 3.4805
R32200 GND.n4818 GND.t406 3.4805
R32201 GND.n4804 GND.t180 3.4805
R32202 GND.n4804 GND.t156 3.4805
R32203 GND.n4789 GND.t404 3.4805
R32204 GND.n4789 GND.t198 3.4805
R32205 GND.n4183 GND.t170 3.4805
R32206 GND.n4183 GND.t195 3.4805
R32207 GND.n4877 GND.t30 3.4805
R32208 GND.n4877 GND.t172 3.4805
R32209 GND.n4890 GND.t212 3.4805
R32210 GND.n4890 GND.t182 3.4805
R32211 GND.n4903 GND.t184 3.4805
R32212 GND.n4903 GND.t158 3.4805
R32213 GND.n4916 GND.t271 3.4805
R32214 GND.n4916 GND.t36 3.4805
R32215 GND.n4929 GND.t162 3.4805
R32216 GND.n4929 GND.t73 3.4805
R32217 GND.n4164 GND.t277 3.4805
R32218 GND.n4164 GND.t123 3.4805
R32219 GND.n6983 GND.n6982 3.47289
R32220 GND.n5438 GND.n5437 3.42801
R32221 GND.n5438 GND.n5010 3.42801
R32222 GND.n5689 GND.n5688 3.42801
R32223 GND.n5688 GND.n5009 3.42801
R32224 GND.n6351 GND.n2713 3.42801
R32225 GND.n6353 GND.n2713 3.42801
R32226 GND.n6425 GND.n6424 3.42801
R32227 GND.n6425 GND.n2714 3.42801
R32228 GND.n8789 GND.n8788 3.42801
R32229 GND.n8789 GND.n997 3.42801
R32230 GND.n1461 GND.n1460 3.42801
R32231 GND.n1460 GND.n1365 3.42801
R32232 GND.n1454 GND.n1453 3.42801
R32233 GND.n1454 GND.n1366 3.42801
R32234 GND.n8530 GND.n996 3.42801
R32235 GND.n8528 GND.n996 3.42801
R32236 GND.n3504 GND.n3503 3.42801
R32237 GND.n3503 GND.n3412 3.42801
R32238 GND.n3501 GND.n3500 3.42801
R32239 GND.n3501 GND.n3413 3.42801
R32240 GND.n4943 GND.n4942 3.42801
R32241 GND.n4942 GND.n3933 3.42801
R32242 GND.n4152 GND.n4151 3.42801
R32243 GND.n4152 GND.n3934 3.42801
R32244 GND.n5629 GND.n5628 3.4105
R32245 GND.n9605 GND.n9604 3.4105
R32246 GND.n7978 GND.n7977 3.4105
R32247 GND.t280 GND.n82 3.3958
R32248 GND.t50 GND.n2166 3.3958
R32249 GND.n3091 GND.n2899 3.38874
R32250 GND.n6597 GND.n6588 3.38531
R32251 GND.n6583 GND.n6574 3.38531
R32252 GND.n6569 GND.n6560 3.38531
R32253 GND.n6555 GND.n6546 3.38531
R32254 GND.n6541 GND.n6532 3.38531
R32255 GND.n2707 GND.n2698 3.38531
R32256 GND.n6456 GND.n6447 3.38531
R32257 GND.n6470 GND.n6446 3.38531
R32258 GND.n6483 GND.n6445 3.38531
R32259 GND.n6496 GND.n6444 3.38531
R32260 GND.n6509 GND.n6443 3.38531
R32261 GND.n6522 GND.n6442 3.38531
R32262 GND.n6437 GND.n6428 3.38531
R32263 GND.n8960 GND.n8951 3.38531
R32264 GND.n8946 GND.n8937 3.38531
R32265 GND.n8932 GND.n8923 3.38531
R32266 GND.n8918 GND.n8909 3.38531
R32267 GND.n8904 GND.n8895 3.38531
R32268 GND.n990 GND.n981 3.38531
R32269 GND.n8820 GND.n8811 3.38531
R32270 GND.n8834 GND.n8810 3.38531
R32271 GND.n8847 GND.n8809 3.38531
R32272 GND.n8860 GND.n8808 3.38531
R32273 GND.n8873 GND.n8807 3.38531
R32274 GND.n8886 GND.n8806 3.38531
R32275 GND.n8801 GND.n8792 3.38531
R32276 GND.n4859 GND.n4850 3.38531
R32277 GND.n4845 GND.n4836 3.38531
R32278 GND.n4831 GND.n4822 3.38531
R32279 GND.n4817 GND.n4808 3.38531
R32280 GND.n4803 GND.n4794 3.38531
R32281 GND.n4788 GND.n4779 3.38531
R32282 GND.n4182 GND.n4173 3.38531
R32283 GND.n4876 GND.n4172 3.38531
R32284 GND.n4889 GND.n4171 3.38531
R32285 GND.n4902 GND.n4170 3.38531
R32286 GND.n4915 GND.n4169 3.38531
R32287 GND.n4928 GND.n4168 3.38531
R32288 GND.n4163 GND.n4154 3.38531
R32289 GND.n9463 GND.n189 3.38095
R32290 GND.n7748 GND.n1871 3.38095
R32291 GND.n9047 GND.t253 3.27919
R32292 GND.n4771 GND.t157 3.27919
R32293 GND.n7244 GND.t221 3.27919
R32294 GND.n3033 GND.n3032 3.2773
R32295 GND.t274 GND.n2093 3.2606
R32296 GND.t32 GND.n76 3.24147
R32297 GND.n7881 GND.t51 3.24147
R32298 GND.n9784 GND.n9783 3.21479
R32299 GND.n9793 GND.n9792 3.21479
R32300 GND.n9794 GND.n9793 3.21479
R32301 GND.n21 GND.n19 3.21479
R32302 GND.n9432 GND.n19 3.21479
R32303 GND.n20 GND.n18 3.21479
R32304 GND.t3 GND.n18 3.21479
R32305 GND.n8430 GND.n8429 3.21479
R32306 GND.n8431 GND.n8430 3.21479
R32307 GND.n1806 GND.n1805 3.21479
R32308 GND.n1805 GND.n17 3.21479
R32309 GND.n7742 GND.n7741 3.21479
R32310 GND.n7741 GND.t224 3.21479
R32311 GND.n7746 GND.n7745 3.21479
R32312 GND.t69 GND.n7746 3.21479
R32313 GND.n8423 GND.n8422 3.20815
R32314 GND.n9096 GND.t229 3.19221
R32315 GND.n9387 GND.n251 3.01226
R32316 GND.n9369 GND.n271 3.01226
R32317 GND.n954 GND.n472 3.01226
R32318 GND.n974 GND.n965 3.01226
R32319 GND.n261 GND.n242 3.01226
R32320 GND.n281 GND.n280 3.01226
R32321 GND.n8977 GND.n462 3.01226
R32322 GND.n9021 GND.n9020 3.01226
R32323 GND.n842 GND.n841 3.01226
R32324 GND.n9051 GND.n9049 3.01226
R32325 GND.n940 GND.n939 3.01226
R32326 GND.n9036 GND.n9035 3.01226
R32327 GND.n8281 GND.n1943 3.01226
R32328 GND.n8263 GND.n1963 3.01226
R32329 GND.n4688 GND.n4211 3.01226
R32330 GND.n4706 GND.n4695 3.01226
R32331 GND.n1953 GND.n1934 3.01226
R32332 GND.n1973 GND.n1972 3.01226
R32333 GND.n4495 GND.n4494 3.01226
R32334 GND.n4764 GND.n4725 3.01226
R32335 GND.n4488 GND.n4471 3.01226
R32336 GND.n4769 GND.n4768 3.01226
R32337 GND.n4468 GND.n4466 3.01226
R32338 GND.n4652 GND.n4195 3.01226
R32339 GND.n7222 GND.n6614 3.01226
R32340 GND.n7312 GND.n2550 3.01226
R32341 GND.n7204 GND.n6628 3.01226
R32342 GND.n7302 GND.n2567 3.01226
R32343 GND.n7216 GND.n6625 3.01226
R32344 GND.n7289 GND.n2562 3.01226
R32345 GND.n7184 GND.n7183 3.01226
R32346 GND.n7233 GND.n2542 3.01226
R32347 GND.n7179 GND.n7178 3.01226
R32348 GND.n7242 GND.n7241 3.01226
R32349 GND.n7165 GND.n6634 3.01226
R32350 GND.n7246 GND.n2638 3.01226
R32351 GND.n6422 GND.n2717 2.9445
R32352 GND.n8786 GND.n1000 2.9445
R32353 GND.n4149 GND.n3951 2.9445
R32354 GND.n7581 GND.n2418 2.91552
R32355 GND.n8030 GND.n2113 2.91475
R32356 GND.n2959 GND.n2926 2.8677
R32357 GND.n3001 GND.n3000 2.8677
R32358 GND.n9541 GND.t247 2.77847
R32359 GND.n7818 GND.t196 2.77847
R32360 GND.n9207 GND.n9135 2.73625
R32361 GND.n5693 GND.n5004 2.6885
R32362 GND.n1437 GND.n1435 2.6885
R32363 GND.n3484 GND.n3482 2.6885
R32364 GND.n791 GND.n752 2.62345
R32365 GND.n9405 GND.n9404 2.62345
R32366 GND.n927 GND.n926 2.62345
R32367 GND.n9398 GND.n234 2.62345
R32368 GND.n949 GND.n475 2.62345
R32369 GND.n9390 GND.n244 2.62345
R32370 GND.n8975 GND.n463 2.62345
R32371 GND.n9381 GND.n256 2.62345
R32372 GND.n9030 GND.t39 2.62345
R32373 GND.n9375 GND.n266 2.62345
R32374 GND.n9047 GND.n9046 2.62345
R32375 GND.n9366 GND.n275 2.62345
R32376 GND.n9059 GND.n358 2.62345
R32377 GND.n9358 GND.n286 2.62345
R32378 GND.n9281 GND.n9280 2.62345
R32379 GND.n9310 GND.n321 2.62345
R32380 GND.n4449 GND.n4448 2.62345
R32381 GND.n8299 GND.n8298 2.62345
R32382 GND.n4504 GND.n4503 2.62345
R32383 GND.n8292 GND.n1926 2.62345
R32384 GND.n4683 GND.n4214 2.62345
R32385 GND.n8284 GND.n1936 2.62345
R32386 GND.n4492 GND.n4490 2.62345
R32387 GND.n8275 GND.n1948 2.62345
R32388 GND.n4714 GND.t40 2.62345
R32389 GND.n8269 GND.n1958 2.62345
R32390 GND.n4771 GND.n4196 2.62345
R32391 GND.n8260 GND.n1967 2.62345
R32392 GND.n4647 GND.n2050 2.62345
R32393 GND.n8252 GND.n1978 2.62345
R32394 GND.n8175 GND.n8174 2.62345
R32395 GND.n8204 GND.n2013 2.62345
R32396 GND.n7141 GND.n7140 2.62345
R32397 GND.n7125 GND.n6688 2.62345
R32398 GND.n7154 GND.n6664 2.62345
R32399 GND.n7133 GND.n6683 2.62345
R32400 GND.n7174 GND.n7173 2.62345
R32401 GND.n7219 GND.n6618 2.62345
R32402 GND.n7202 GND.n6629 2.62345
R32403 GND.n7228 GND.n6609 2.62345
R32404 GND.n7191 GND.t238 2.62345
R32405 GND.n7309 GND.n2555 2.62345
R32406 GND.n7244 GND.n2689 2.62345
R32407 GND.n7320 GND.n2545 2.62345
R32408 GND.n7297 GND.n2617 2.62345
R32409 GND.n7375 GND.n7374 2.62345
R32410 GND.n2677 GND.n2505 2.62345
R32411 GND.n2670 GND.n2495 2.62345
R32412 GND.n2277 GND.t83 2.60536
R32413 GND.n7684 GND.t193 2.60536
R32414 GND.n7685 GND.t19 2.60536
R32415 GND.n7686 GND.t378 2.60536
R32416 GND.n9801 GND.t125 2.60536
R32417 GND.n9800 GND.t56 2.60536
R32418 GND.n9799 GND.t214 2.60536
R32419 GND.n28 GND.t380 2.60536
R32420 GND.n8405 GND.t71 2.60536
R32421 GND.n8404 GND.t168 2.60536
R32422 GND.n8403 GND.t426 2.60536
R32423 GND.n8402 GND.t408 2.60536
R32424 GND.n5622 GND.t58 2.46987
R32425 GND.n3078 GND.n3077 2.4581
R32426 GND.n6338 GND.n6337 2.4325
R32427 GND.n8517 GND.n8516 2.4325
R32428 GND.n3950 GND.n3949 2.4325
R32429 GND.n7511 GND.n2307 2.41091
R32430 GND.n9228 GND.t227 2.28029
R32431 GND.n8972 GND.n468 2.25932
R32432 GND.n887 GND.n451 2.25932
R32433 GND.n898 GND.n874 2.25932
R32434 GND.n885 GND.n884 2.25932
R32435 GND.n4675 GND.n4674 2.25932
R32436 GND.n4547 GND.n4546 2.25932
R32437 GND.n4670 GND.n4228 2.25932
R32438 GND.n4664 GND.n4535 2.25932
R32439 GND.n7199 GND.n6632 2.25932
R32440 GND.n2634 GND.n2623 2.25932
R32441 GND.n7033 GND.n7029 2.25932
R32442 GND.n7256 GND.n2627 2.25932
R32443 GND.n5692 GND.n5005 2.1765
R32444 GND.n1439 GND.n1438 2.1765
R32445 GND.n3486 GND.n3485 2.1765
R32446 GND.t423 GND.n2345 2.05831
R32447 GND.n5610 GND.t189 2.05831
R32448 GND.n7698 GND.n2306 1.9855
R32449 GND.n8975 GND.t327 1.96771
R32450 GND.n4492 GND.t405 1.96771
R32451 GND.n7202 GND.t24 1.96771
R32452 GND.n6341 GND.n6340 1.9205
R32453 GND.n8521 GND.n8519 1.9205
R32454 GND.n3946 GND.n3938 1.9205
R32455 GND.n7589 GND.t192 1.85253
R32456 GND.n9688 GND.t264 1.85248
R32457 GND.n7986 GND.t185 1.85248
R32458 GND.n3034 GND.n2906 1.8437
R32459 GND.n3053 GND.n2904 1.8437
R32460 GND.n5982 GND.n3717 1.77928
R32461 GND.n5895 GND.n5894 1.77928
R32462 GND.n5279 GND.n3725 1.77928
R32463 GND.n5888 GND.n3731 1.77928
R32464 GND.n5887 GND.n3734 1.77928
R32465 GND.n3957 GND.n3742 1.77928
R32466 GND.n5881 GND.n5880 1.77928
R32467 GND.n5288 GND.n3745 1.77928
R32468 GND.n5874 GND.n3751 1.77928
R32469 GND.n5873 GND.n3754 1.77928
R32470 GND.t4 GND.t375 1.77928
R32471 GND.n3966 GND.n3760 1.77928
R32472 GND.n5867 GND.n5866 1.77928
R32473 GND.n5297 GND.n3763 1.77928
R32474 GND.n5860 GND.n3769 1.77928
R32475 GND.n5859 GND.n3772 1.77928
R32476 GND.n3975 GND.n3778 1.77928
R32477 GND.n5853 GND.n5852 1.77928
R32478 GND.n5306 GND.n3781 1.77928
R32479 GND.n5846 GND.n3787 1.77928
R32480 GND.n5845 GND.n3789 1.77928
R32481 GND.n5809 GND.n3837 1.77928
R32482 GND.n4079 GND.n3843 1.77928
R32483 GND.n5778 GND.n5777 1.77928
R32484 GND.n5372 GND.n3846 1.77928
R32485 GND.n5771 GND.n3852 1.77928
R32486 GND.n5770 GND.n3855 1.77928
R32487 GND.n4088 GND.n3861 1.77928
R32488 GND.n5764 GND.n5763 1.77928
R32489 GND.n5381 GND.n3864 1.77928
R32490 GND.n5757 GND.n3870 1.77928
R32491 GND.t370 GND.t62 1.77928
R32492 GND.n5756 GND.n3873 1.77928
R32493 GND.n4097 GND.n3879 1.77928
R32494 GND.n5750 GND.n5749 1.77928
R32495 GND.n5390 GND.n3882 1.77928
R32496 GND.n5743 GND.n3888 1.77928
R32497 GND.n5742 GND.n3891 1.77928
R32498 GND.n4106 GND.n3897 1.77928
R32499 GND.n5736 GND.n5735 1.77928
R32500 GND.n5400 GND.n3900 1.77928
R32501 GND.n5729 GND.n4982 1.77928
R32502 GND.t127 GND.n2418 1.74971
R32503 GND.t29 GND.n2113 1.74925
R32504 GND.n6426 GND.n6425 1.6975
R32505 GND.n6426 GND.n2713 1.6975
R32506 GND.n1459 GND.n1454 1.6975
R32507 GND.n1460 GND.n1459 1.6975
R32508 GND.n8790 GND.n8789 1.6975
R32509 GND.n8790 GND.n996 1.6975
R32510 GND.n4941 GND.n4152 1.6975
R32511 GND.n4942 GND.n4941 1.6975
R32512 GND.n3502 GND.n3501 1.6975
R32513 GND.n3503 GND.n3502 1.6975
R32514 GND.n5688 GND.n5687 1.6975
R32515 GND.n5687 GND.n5438 1.6975
R32516 GND.n7688 GND.n7686 1.68459
R32517 GND.n9807 GND.n28 1.68459
R32518 GND.n8402 GND.n8398 1.68459
R32519 GND.n5017 GND.n5008 1.6645
R32520 GND.n1451 GND.n1450 1.6645
R32521 GND.n3498 GND.n3497 1.6645
R32522 GND.n7733 GND.n2277 1.66167
R32523 GND.n9802 GND.n9801 1.66167
R32524 GND.n8406 GND.n8405 1.66167
R32525 GND.t22 GND.n2461 1.56018
R32526 GND.n8101 GND.t194 1.55968
R32527 GND.t250 GND.n566 1.55968
R32528 GND.n1834 GND.t276 1.55968
R32529 GND.n9533 GND.t330 1.54382
R32530 GND.t329 GND.n108 1.54382
R32531 GND.n7799 GND.t303 1.54382
R32532 GND.t21 GND.n2191 1.54382
R32533 GND.n7739 GND.n7 1.51986
R32534 GND.n9813 GND.n24 1.51986
R32535 GND.n979 GND.n978 1.51971
R32536 GND.n4696 GND.n4187 1.51971
R32537 GND.n6605 GND.n2563 1.51971
R32538 GND.t208 GND.n189 1.51615
R32539 GND.t179 GND.n1871 1.51615
R32540 GND.n9384 GND.n9383 1.50638
R32541 GND.n9373 GND.n9372 1.50638
R32542 GND.n959 GND.n958 1.50638
R32543 GND.n963 GND.n962 1.50638
R32544 GND.n9379 GND.n262 1.50638
R32545 GND.n9377 GND.n264 1.50638
R32546 GND.n8979 GND.n8978 1.50638
R32547 GND.n9023 GND.n9022 1.50638
R32548 GND.n828 GND.n458 1.50638
R32549 GND.n9027 GND.n444 1.50638
R32550 GND.n485 GND.n484 1.50638
R32551 GND.n9037 GND.n9033 1.50638
R32552 GND.n8278 GND.n8277 1.50638
R32553 GND.n8267 GND.n8266 1.50638
R32554 GND.n4693 GND.n4692 1.50638
R32555 GND.n4711 GND.n4710 1.50638
R32556 GND.n8273 GND.n1954 1.50638
R32557 GND.n8271 GND.n1956 1.50638
R32558 GND.n4257 GND.n4204 1.50638
R32559 GND.n4723 GND.n4722 1.50638
R32560 GND.n4487 GND.n4207 1.50638
R32561 GND.n4208 GND.n4199 1.50638
R32562 GND.n4467 GND.n4191 1.50638
R32563 GND.n4774 GND.n4193 1.50638
R32564 GND.n7226 GND.n7225 1.50638
R32565 GND.n7313 GND.n7311 1.50638
R32566 GND.n7206 GND.n7205 1.50638
R32567 GND.n7207 GND.n2564 1.50638
R32568 GND.n7212 GND.n7211 1.50638
R32569 GND.n7307 GND.n7306 1.50638
R32570 GND.n7185 GND.n2695 1.50638
R32571 GND.n7234 GND.n7232 1.50638
R32572 GND.n6644 GND.n6638 1.50638
R32573 GND.n7188 GND.n2692 1.50638
R32574 GND.n7195 GND.n7194 1.50638
R32575 GND.n7247 GND.n2637 1.50638
R32576 GND.n9825 GND.n9 1.43919
R32577 GND.n875 GND.n471 1.43699
R32578 GND.n4667 GND.n4188 1.43699
R32579 GND.n6529 GND.n2629 1.43699
R32580 GND.n2956 GND.n2925 1.4341
R32581 GND.n3002 GND.n3001 1.4341
R32582 GND.n979 GND.n461 1.41953
R32583 GND.n8969 GND.n8968 1.41953
R32584 GND.n4719 GND.n4187 1.41953
R32585 GND.n4777 GND.n4776 1.41953
R32586 GND.n6606 GND.n6605 1.41953
R32587 GND.n2696 GND.n2635 1.41953
R32588 GND.n6349 GND.n6330 1.4085
R32589 GND.n8526 GND.n8515 1.4085
R32590 GND.n3932 GND.n3929 1.4085
R32591 GND.n9681 GND.t55 1.38949
R32592 GND.n7994 GND.t167 1.38949
R32593 GND.n6948 GND.t419 1.36838
R32594 GND.n9404 GND.t43 1.31198
R32595 GND.t257 GND.t306 1.31198
R32596 GND.t327 GND.t206 1.31198
R32597 GND.t253 GND.t325 1.31198
R32598 GND.t244 GND.t321 1.31198
R32599 GND.n351 GND.t1 1.31198
R32600 GND.n9352 GND.t1 1.31198
R32601 GND.t231 GND.t233 1.31198
R32602 GND.n8298 GND.t13 1.31198
R32603 GND.t428 GND.t35 1.31198
R32604 GND.t405 GND.t183 1.31198
R32605 GND.t157 GND.t164 1.31198
R32606 GND.t211 GND.t177 1.31198
R32607 GND.n2043 GND.t54 1.31198
R32608 GND.n8246 GND.t54 1.31198
R32609 GND.t33 GND.t181 1.31198
R32610 GND.n7125 GND.t239 1.31198
R32611 GND.t118 GND.t77 1.31198
R32612 GND.t24 GND.t108 1.31198
R32613 GND.t221 GND.t120 1.31198
R32614 GND.t75 GND.t217 1.31198
R32615 GND.n7389 GND.t44 1.31198
R32616 GND.n7368 GND.t44 1.31198
R32617 GND.t106 GND.t116 1.31198
R32618 GND.n9780 GND.n49 1.30521
R32619 GND.n8420 GND.n8419 1.30521
R32620 GND.n995 GND.n26 1.30521
R32621 GND.n5684 GND.n2275 1.30521
R32622 GND.n4939 GND.n1814 1.30521
R32623 GND.n5439 GND.n2314 1.30521
R32624 GND.n562 GND.t319 1.27619
R32625 GND.n8347 GND.t403 1.27619
R32626 GND.n9770 GND.n49 1.2598
R32627 GND.n8419 GND.n8418 1.2598
R32628 GND.n9768 GND.n26 1.2598
R32629 GND.n5674 GND.n2275 1.2598
R32630 GND.n8412 GND.n1814 1.2598
R32631 GND.n5671 GND.n2314 1.2598
R32632 GND.n7687 GND.n2278 1.21056
R32633 GND.n9806 GND.n9805 1.2101
R32634 GND.n8410 GND.n8409 1.2101
R32635 GND.n5678 GND.n5671 1.20311
R32636 GND.n9774 GND.n9768 1.20311
R32637 GND.n8413 GND.n8412 1.20311
R32638 GND.n5025 GND.n5014 1.1525
R32639 GND.n1444 GND.n1442 1.1525
R32640 GND.n3491 GND.n3489 1.1525
R32641 GND.n5675 GND.n5674 1.13828
R32642 GND.n7732 GND.n7731 1.13828
R32643 GND.n9804 GND.n9803 1.13828
R32644 GND.n9771 GND.n9770 1.13828
R32645 GND.n8408 GND.n8407 1.13828
R32646 GND.n8418 GND.n8417 1.13828
R32647 GND.n7687 GND.n2315 1.1243
R32648 GND.n7732 GND.n2276 1.1243
R32649 GND.n9803 GND.n48 1.1243
R32650 GND.n9806 GND.n27 1.1243
R32651 GND.n8407 GND.n1810 1.1243
R32652 GND.n8411 GND.n8410 1.1243
R32653 GND.n4940 GND.n4939 1.03305
R32654 GND.n8791 GND.n995 1.03266
R32655 GND.n3056 GND.n3055 1.0245
R32656 GND.n7727 GND.n7726 1.01931
R32657 GND.n7581 GND.n7580 0.993024
R32658 GND.n7560 GND.t65 0.993024
R32659 GND.n8030 GND.n2070 0.992704
R32660 GND.n4604 GND.t169 0.992704
R32661 GND.n9463 GND.n9431 0.992704
R32662 GND.n7748 GND.n2272 0.992704
R32663 GND.t227 GND.t235 0.912417
R32664 GND.t229 GND.t259 0.912417
R32665 GND.n6905 GND.n6904 0.912417
R32666 GND.t284 GND.t187 0.912417
R32667 GND.t419 GND.t114 0.912417
R32668 GND.n6329 GND.n6327 0.8965
R32669 GND.n8513 GND.n8511 0.8965
R32670 GND.n4947 GND.n4946 0.8965
R32671 GND.t59 GND.n2307 0.851235
R32672 GND.n7552 GND.n2461 0.851235
R32673 GND.n8101 GND.n2108 0.850961
R32674 GND.n6531 GND.n6530 0.759389
R32675 GND.n6528 GND.n6527 0.759389
R32676 GND.n8894 GND.n8893 0.759389
R32677 GND.n8892 GND.n8891 0.759389
R32678 GND.n8825 GND.n980 0.759389
R32679 GND.n8966 GND.n8965 0.759389
R32680 GND.n4793 GND.n4153 0.759389
R32681 GND.n4934 GND.n4933 0.759389
R32682 GND.n4867 GND.n4866 0.759389
R32683 GND.n4865 GND.n4864 0.759389
R32684 GND.n6461 GND.n2697 0.759389
R32685 GND.n6603 GND.n6602 0.759389
R32686 GND.n2979 GND.n2978 0.753441
R32687 GND.n2943 GND.n2942 0.753441
R32688 GND.n2992 GND.n2991 0.753441
R32689 GND.n3007 GND.n2917 0.753441
R32690 GND.n3015 GND.n2913 0.753441
R32691 GND.n3065 GND.n3046 0.753441
R32692 GND.n3041 GND.n3040 0.753441
R32693 GND.n8971 GND.n469 0.753441
R32694 GND.n889 GND.n888 0.753441
R32695 GND.n895 GND.n894 0.753441
R32696 GND.n877 GND.n876 0.753441
R32697 GND.n4542 GND.n4224 0.753441
R32698 GND.n4545 GND.n4544 0.753441
R32699 GND.n4669 GND.n4229 0.753441
R32700 GND.n4665 GND.n4534 0.753441
R32701 GND.n7198 GND.n2633 0.753441
R32702 GND.n7251 GND.n7250 0.753441
R32703 GND.n7030 GND.n2630 0.753441
R32704 GND.n7257 GND.n7255 0.753441
R32705 GND.n9803 GND.n9802 0.726297
R32706 GND.n8407 GND.n8406 0.726297
R32707 GND.n9807 GND.n9806 0.726297
R32708 GND.n7733 GND.n7732 0.726297
R32709 GND.n8410 GND.n8398 0.726297
R32710 GND.n7688 GND.n7687 0.726297
R32711 GND.t67 GND.n2429 0.709446
R32712 GND.n9788 GND.n9785 0.709347
R32713 GND.n8428 GND.n8427 0.709347
R32714 GND.n8122 GND.t173 0.709217
R32715 GND.n9790 GND.n9789 0.688
R32716 GND.n9789 GND.n9788 0.688
R32717 GND.n8423 GND.n1804 0.688
R32718 GND.n8427 GND.n1804 0.688
R32719 GND.n9415 GND.t255 0.656238
R32720 GND.n9415 GND.t99 0.656238
R32721 GND.t233 GND.n301 0.656238
R32722 GND.n8309 GND.t155 0.656238
R32723 GND.n8309 GND.t270 0.656238
R32724 GND.t181 GND.n1993 0.656238
R32725 GND.t410 GND.n7062 0.656238
R32726 GND.n7062 GND.t421 0.656238
R32727 GND.n2498 GND.t106 0.656238
R32728 GND.n5027 GND.n5026 0.6405
R32729 GND.n1440 GND.n1362 0.6405
R32730 GND.n3487 GND.n3409 0.6405
R32731 GND.n7640 GND.n7639 0.617842
R32732 GND.n5541 GND.n2339 0.617842
R32733 GND.t400 GND.t423 0.617842
R32734 GND.n7633 GND.n2345 0.617842
R32735 GND.n7632 GND.n2348 0.617842
R32736 GND.n5513 GND.n2356 0.617842
R32737 GND.t79 GND.t126 0.617842
R32738 GND.t203 GND.t190 0.617842
R32739 GND.n5606 GND.n5605 0.617842
R32740 GND.n7605 GND.n7604 0.617842
R32741 GND.n5610 GND.n2390 0.617842
R32742 GND.t189 GND.t401 0.617842
R32743 GND.n7598 GND.n2396 0.617842
R32744 GND.n7597 GND.n2399 0.617842
R32745 GND.n2997 GND.n2925 0.6149
R32746 GND.n6427 GND.n2712 0.589937
R32747 GND.n4941 GND.n4940 0.548285
R32748 GND.n6427 GND.n6426 0.547165
R32749 GND.n8791 GND.n8790 0.547165
R32750 GND.n3502 GND.n1807 0.547165
R32751 GND.n5687 GND.n5686 0.547165
R32752 GND.n9825 GND.n9824 0.541695
R32753 GND.t323 GND.t240 0.538397
R32754 GND.t398 GND.t201 0.538397
R32755 GND.n1459 GND.n1458 0.535303
R32756 GND.n7709 GND.n2306 0.5005
R32757 GND.n7710 GND.n7709 0.5005
R32758 GND.n7724 GND.n2297 0.5005
R32759 GND.n9446 GND.n9 0.5005
R32760 GND.n9447 GND.n9446 0.5005
R32761 GND.n9447 GND.n9437 0.5005
R32762 GND.n9457 GND.n9437 0.5005
R32763 GND.n9458 GND.n9457 0.5005
R32764 GND.n7710 GND.n2295 0.49675
R32765 GND.n2936 GND 0.484875
R32766 GND.n176 GND.n175 0.463495
R32767 GND.n9560 GND.n171 0.463495
R32768 GND.t330 GND.t246 0.463495
R32769 GND.n9533 GND.n9532 0.463495
R32770 GND.n9579 GND.n166 0.463495
R32771 GND.n9526 GND.n9522 0.463495
R32772 GND.t252 GND.t267 0.463495
R32773 GND.t312 GND.t98 0.463495
R32774 GND.n9735 GND.n90 0.463495
R32775 GND.n9703 GND.n96 0.463495
R32776 GND.n9702 GND.n108 0.463495
R32777 GND.t261 GND.t329 0.463495
R32778 GND.n9638 GND.n118 0.463495
R32779 GND.n9696 GND.n9695 0.463495
R32780 GND.n2263 GND.n2262 0.463495
R32781 GND.n7839 GND.n2257 0.463495
R32782 GND.t303 GND.t86 0.463495
R32783 GND.n7799 GND.n2219 0.463495
R32784 GND.n7867 GND.n7866 0.463495
R32785 GND.n7874 GND.n2213 0.463495
R32786 GND.t186 GND.t355 0.463495
R32787 GND.t175 GND.t338 0.463495
R32788 GND.n7956 GND.n2174 0.463495
R32789 GND.n7924 GND.n2180 0.463495
R32790 GND.n7923 GND.n2191 0.463495
R32791 GND.t281 GND.t21 0.463495
R32792 GND.n7911 GND.n7910 0.463495
R32793 GND.n7905 GND.n2137 0.463495
R32794 GND.n5439 GND.n2712 0.443226
R32795 GND.n711 GND.t242 0.42573
R32796 GND.n4326 GND.t161 0.42573
R32797 GND.n7625 GND.n2359 0.412061
R32798 GND.n5651 GND.n5650 0.412061
R32799 GND.n7619 GND.n7618 0.412061
R32800 GND.n5660 GND.n5447 0.412061
R32801 GND.n7612 GND.n2378 0.412061
R32802 GND.n5562 GND.n2381 0.412061
R32803 GND.n2956 GND.n2955 0.4101
R32804 GND.n2996 GND.n2926 0.4101
R32805 GND.n3002 GND.n2922 0.4101
R32806 GND.n3006 GND.n2920 0.4101
R32807 GND.n3034 GND.n3033 0.4101
R32808 GND.n3077 GND.n2907 0.4101
R32809 GND.n3055 GND.n3053 0.4101
R32810 GND.n3082 GND.n2900 0.4101
R32811 GND.n3087 GND.n2901 0.4101
R32812 GND.n6356 GND.n6355 0.3845
R32813 GND.n8534 GND.n8532 0.3845
R32814 GND.n4950 GND.n3928 0.3845
R32815 GND.n5679 GND.n5678 0.3805
R32816 GND.n5678 GND.n5672 0.3805
R32817 GND.n5683 GND.n5669 0.3805
R32818 GND.n5680 GND.n5440 0.3805
R32819 GND.n9775 GND.n9774 0.3805
R32820 GND.n9774 GND.n9769 0.3805
R32821 GND.n9779 GND.n9766 0.3805
R32822 GND.n9776 GND.n58 0.3805
R32823 GND.n1458 GND.n1457 0.3805
R32824 GND.n1457 GND.n56 0.3805
R32825 GND.n8414 GND.n8413 0.3805
R32826 GND.n8413 GND.n1812 0.3805
R32827 GND.n4936 GND.n1809 0.3805
R32828 GND.n4938 GND.n1813 0.3805
R32829 GND.n2294 GND.n2293 0.3805
R32830 GND.n2293 GND.n2292 0.3805
R32831 GND.n2292 GND.n2291 0.3805
R32832 GND.n2287 GND.n2286 0.3805
R32833 GND.n2291 GND.n2286 0.3805
R32834 GND.n2287 GND.n2285 0.3805
R32835 GND.n2291 GND.n2285 0.3805
R32836 GND.n2291 GND.n2290 0.3805
R32837 GND.n9829 GND.n9828 0.3805
R32838 GND.n9832 GND.n2 0.3805
R32839 GND.n9829 GND.n2 0.3805
R32840 GND.n9832 GND.n5 0.3805
R32841 GND.n9829 GND.n5 0.3805
R32842 GND.n9832 GND.n1 0.3805
R32843 GND.n9829 GND.n1 0.3805
R32844 GND.n9832 GND.n9831 0.3805
R32845 GND.n44 GND.n43 0.3805
R32846 GND.n40 GND.n33 0.3805
R32847 GND.n43 GND.n33 0.3805
R32848 GND.n40 GND.n36 0.3805
R32849 GND.n43 GND.n36 0.3805
R32850 GND.n40 GND.n32 0.3805
R32851 GND.n43 GND.n32 0.3805
R32852 GND.n43 GND.n42 0.3805
R32853 GND.n2973 GND.n2971 0.376971
R32854 GND.n9770 GND.n48 0.356443
R32855 GND.n8418 GND.n1810 0.356443
R32856 GND.n9768 GND.n27 0.356443
R32857 GND.n5674 GND.n2276 0.356443
R32858 GND.n8412 GND.n8411 0.356443
R32859 GND.n5671 GND.n2315 0.356443
R32860 GND.n5686 GND.n5685 0.349946
R32861 GND.n7686 GND.n7685 0.323417
R32862 GND.n7684 GND.n2277 0.323417
R32863 GND.n9799 GND.n28 0.323417
R32864 GND.n9801 GND.n9800 0.323417
R32865 GND.n8403 GND.n8402 0.323417
R32866 GND.n8405 GND.n8404 0.323417
R32867 GND.n7685 GND.n7684 0.321333
R32868 GND.n9800 GND.n9799 0.321333
R32869 GND.n8404 GND.n8403 0.321333
R32870 GND.n9589 GND.n9588 0.309164
R32871 GND.n9749 GND.n76 0.309164
R32872 GND.n154 GND.n65 0.309164
R32873 GND.n9565 GND.n66 0.309164
R32874 GND.n9742 GND.n9741 0.309164
R32875 GND.n9710 GND.n9709 0.309164
R32876 GND.n7845 GND.n2215 0.309164
R32877 GND.n7882 GND.n7881 0.309164
R32878 GND.n7969 GND.n2160 0.309164
R32879 GND.n7856 GND.n7855 0.309164
R32880 GND.n7963 GND.n7962 0.309164
R32881 GND.n7931 GND.n7930 0.309164
R32882 GND.n2847 GND.n2810 0.3077
R32883 GND.n8671 GND.n8670 0.3077
R32884 GND.n4044 GND.n4043 0.3077
R32885 GND.n7743 GND.n7739 0.300787
R32886 GND.n9813 GND.n9812 0.300787
R32887 GND.n8 GND 0.288767
R32888 GND.t412 GND.t67 0.284078
R32889 GND.t65 GND.t59 0.284078
R32890 GND.t173 GND.t171 0.283987
R32891 GND.t169 GND.t274 0.283987
R32892 GND.n678 GND.n566 0.283987
R32893 GND.t319 GND.t248 0.283987
R32894 GND.t308 GND.t242 0.283987
R32895 GND.n1835 GND.n1834 0.283987
R32896 GND.t403 GND.t122 0.283987
R32897 GND.t161 GND.t197 0.283987
R32898 GND.n8422 GND.n1807 0.281502
R32899 GND.n9782 GND.n56 0.269106
R32900 GND.n7725 GND.n7724 0.25425
R32901 GND.n7697 GND.n7696 0.2505
R32902 GND.n2115 GND.n10 0.2505
R32903 GND.n7725 GND.n2296 0.24675
R32904 GND.n4866 GND.n1807 0.239239
R32905 GND.n5686 GND.n2697 0.239239
R32906 GND.n8892 GND.n8791 0.237409
R32907 GND.n6528 GND.n6427 0.237409
R32908 GND.n4940 GND.n4934 0.236355
R32909 GND.t219 GND.t127 0.233662
R32910 GND.t301 GND.t29 0.2336
R32911 GND.t225 GND.t208 0.2336
R32912 GND.t72 GND.t179 0.2336
R32913 GND.n7740 GND.n7739 0.233287
R32914 GND.n9814 GND.n9813 0.233287
R32915 GND.t283 GND.n2331 0.206281
R32916 GND.n7626 GND.n7625 0.206281
R32917 GND.n5650 GND.n5461 0.206281
R32918 GND.n7619 GND.n2365 0.206281
R32919 GND.n5447 GND.n2368 0.206281
R32920 GND.n5661 GND.n2378 0.206281
R32921 GND.n7611 GND.n2381 0.206281
R32922 GND.n7591 GND.t58 0.206281
R32923 GND.n3082 GND.n3081 0.2053
R32924 GND.n3088 GND.n3087 0.2053
R32925 GND.n2901 GND.n2899 0.2053
R32926 GND.n2297 GND 0.203
R32927 GND.n9458 GND 0.203
R32928 GND.n7273 GND.n7272 0.196152
R32929 GND.n7272 GND.n7260 0.196152
R32930 GND.n7265 GND.n7260 0.196152
R32931 GND.n7265 GND.n7264 0.196152
R32932 GND.n7264 GND.n2492 0.196152
R32933 GND.n7409 GND.n2492 0.196152
R32934 GND.n7410 GND.n7409 0.196152
R32935 GND.n7415 GND.n7410 0.196152
R32936 GND.n7415 GND.n7414 0.196152
R32937 GND.n882 GND.n363 0.196152
R32938 GND.n9264 GND.n363 0.196152
R32939 GND.n9264 GND.n9263 0.196152
R32940 GND.n9263 GND.n364 0.196152
R32941 GND.n9256 GND.n364 0.196152
R32942 GND.n9256 GND.n9255 0.196152
R32943 GND.n9255 GND.n366 0.196152
R32944 GND.n9248 GND.n366 0.196152
R32945 GND.n9248 GND.n9247 0.196152
R32946 GND.n746 GND.n527 0.196152
R32947 GND.n747 GND.n746 0.196152
R32948 GND.n748 GND.n747 0.196152
R32949 GND.n748 GND.n488 0.196152
R32950 GND.n931 GND.n488 0.196152
R32951 GND.n932 GND.n931 0.196152
R32952 GND.n932 GND.n482 0.196152
R32953 GND.n941 GND.n482 0.196152
R32954 GND.n848 GND.n845 0.196152
R32955 GND.n9394 GND.n241 0.196152
R32956 GND.n9362 GND.n283 0.196152
R32957 GND.n975 GND.n964 0.196152
R32958 GND.n955 GND.n473 0.196152
R32959 GND.n9386 GND.n252 0.196152
R32960 GND.n9386 GND.n9385 0.196152
R32961 GND.n9385 GND.n253 0.196152
R32962 GND.n9371 GND.n253 0.196152
R32963 GND.n9371 GND.n9370 0.196152
R32964 GND.n9370 GND.n272 0.196152
R32965 GND.n9055 GND.n9054 0.196152
R32966 GND.n9055 GND.n344 0.196152
R32967 GND.n9285 GND.n344 0.196152
R32968 GND.n9286 GND.n9285 0.196152
R32969 GND.n9286 GND.n340 0.196152
R32970 GND.n9294 GND.n340 0.196152
R32971 GND.n9295 GND.n9294 0.196152
R32972 GND.n9017 GND.n442 0.196152
R32973 GND.n220 GND.n219 0.196152
R32974 GND.n9410 GND.n220 0.196152
R32975 GND.n9410 GND.n9409 0.196152
R32976 GND.n9409 GND.n221 0.196152
R32977 GND.n833 GND.n221 0.196152
R32978 GND.n834 GND.n833 0.196152
R32979 GND.n834 GND.n826 0.196152
R32980 GND.n843 GND.n826 0.196152
R32981 GND.n9041 GND.n355 0.196152
R32982 GND.n9273 GND.n355 0.196152
R32983 GND.n9274 GND.n9273 0.196152
R32984 GND.n9275 GND.n9274 0.196152
R32985 GND.n9275 GND.n329 0.196152
R32986 GND.n9305 GND.n329 0.196152
R32987 GND.n9305 GND.n9304 0.196152
R32988 GND.n9304 GND.n330 0.196152
R32989 GND.n9239 GND.n330 0.196152
R32990 GND.n453 GND.n435 0.196152
R32991 GND.n9063 GND.n435 0.196152
R32992 GND.n9064 GND.n9063 0.196152
R32993 GND.n9064 GND.n433 0.196152
R32994 GND.n9071 GND.n433 0.196152
R32995 GND.n9072 GND.n9071 0.196152
R32996 GND.n9072 GND.n429 0.196152
R32997 GND.n9079 GND.n429 0.196152
R32998 GND.n9420 GND.n205 0.196152
R32999 GND.n9420 GND.n9419 0.196152
R33000 GND.n9419 GND.n206 0.196152
R33001 GND.n912 GND.n206 0.196152
R33002 GND.n919 GND.n912 0.196152
R33003 GND.n920 GND.n919 0.196152
R33004 GND.n921 GND.n920 0.196152
R33005 GND.n921 GND.n481 0.196152
R33006 GND.n944 GND.n481 0.196152
R33007 GND.n720 GND.n501 0.196152
R33008 GND.n862 GND.n501 0.196152
R33009 GND.n863 GND.n862 0.196152
R33010 GND.n863 GND.n498 0.196152
R33011 GND.n871 GND.n498 0.196152
R33012 GND.n872 GND.n871 0.196152
R33013 GND.n905 GND.n872 0.196152
R33014 GND.n905 GND.n904 0.196152
R33015 GND.n904 GND.n873 0.196152
R33016 GND.n4538 GND.n2055 0.196152
R33017 GND.n8158 GND.n2055 0.196152
R33018 GND.n8158 GND.n8157 0.196152
R33019 GND.n8157 GND.n2056 0.196152
R33020 GND.n8150 GND.n2056 0.196152
R33021 GND.n8150 GND.n8149 0.196152
R33022 GND.n8149 GND.n2058 0.196152
R33023 GND.n8142 GND.n2058 0.196152
R33024 GND.n8142 GND.n8141 0.196152
R33025 GND.n4353 GND.n4352 0.196152
R33026 GND.n4353 GND.n4263 0.196152
R33027 GND.n4453 GND.n4263 0.196152
R33028 GND.n4454 GND.n4453 0.196152
R33029 GND.n4454 GND.n4261 0.196152
R33030 GND.n4462 GND.n4261 0.196152
R33031 GND.n4463 GND.n4462 0.196152
R33032 GND.n4463 GND.n4222 0.196152
R33033 GND.n4498 GND.n4256 0.196152
R33034 GND.n8288 GND.n1933 0.196152
R33035 GND.n8256 GND.n1975 0.196152
R33036 GND.n4707 GND.n4697 0.196152
R33037 GND.n4689 GND.n4212 0.196152
R33038 GND.n8280 GND.n1944 0.196152
R33039 GND.n8280 GND.n8279 0.196152
R33040 GND.n8279 GND.n1945 0.196152
R33041 GND.n8265 GND.n1945 0.196152
R33042 GND.n8265 GND.n8264 0.196152
R33043 GND.n8264 GND.n1964 0.196152
R33044 GND.n4643 GND.n4202 0.196152
R33045 GND.n4643 GND.n2036 0.196152
R33046 GND.n8179 GND.n2036 0.196152
R33047 GND.n8180 GND.n8179 0.196152
R33048 GND.n8180 GND.n2032 0.196152
R33049 GND.n8188 GND.n2032 0.196152
R33050 GND.n8189 GND.n8188 0.196152
R33051 GND.n4765 GND.n4203 0.196152
R33052 GND.n4341 GND.n1912 0.196152
R33053 GND.n8304 GND.n1912 0.196152
R33054 GND.n8304 GND.n8303 0.196152
R33055 GND.n8303 GND.n1913 0.196152
R33056 GND.n4475 GND.n1913 0.196152
R33057 GND.n4475 GND.n4472 0.196152
R33058 GND.n4483 GND.n4472 0.196152
R33059 GND.n4484 GND.n4483 0.196152
R33060 GND.n4657 GND.n2047 0.196152
R33061 GND.n8167 GND.n2047 0.196152
R33062 GND.n8168 GND.n8167 0.196152
R33063 GND.n8169 GND.n8168 0.196152
R33064 GND.n8169 GND.n2021 0.196152
R33065 GND.n8199 GND.n2021 0.196152
R33066 GND.n8199 GND.n8198 0.196152
R33067 GND.n8198 GND.n2022 0.196152
R33068 GND.n8133 GND.n2022 0.196152
R33069 GND.n4653 GND.n4549 0.196152
R33070 GND.n4552 GND.n4549 0.196152
R33071 GND.n4637 GND.n4552 0.196152
R33072 GND.n4637 GND.n4636 0.196152
R33073 GND.n4636 GND.n4553 0.196152
R33074 GND.n4629 GND.n4553 0.196152
R33075 GND.n4629 GND.n4628 0.196152
R33076 GND.n4628 GND.n4557 0.196152
R33077 GND.n8314 GND.n1901 0.196152
R33078 GND.n8314 GND.n8313 0.196152
R33079 GND.n8313 GND.n1902 0.196152
R33080 GND.n4509 GND.n1902 0.196152
R33081 GND.n4516 GND.n4509 0.196152
R33082 GND.n4517 GND.n4516 0.196152
R33083 GND.n4518 GND.n4517 0.196152
R33084 GND.n4518 GND.n4221 0.196152
R33085 GND.n4678 GND.n4221 0.196152
R33086 GND.n8322 GND.n1892 0.196152
R33087 GND.n4239 GND.n1892 0.196152
R33088 GND.n4240 GND.n4239 0.196152
R33089 GND.n4240 GND.n4234 0.196152
R33090 GND.n4247 GND.n4234 0.196152
R33091 GND.n4249 GND.n4247 0.196152
R33092 GND.n4249 GND.n4248 0.196152
R33093 GND.n4248 GND.n4230 0.196152
R33094 GND.n4531 GND.n4230 0.196152
R33095 GND.n6994 GND.n6993 0.196152
R33096 GND.n6993 GND.n6736 0.196152
R33097 GND.n7058 GND.n6736 0.196152
R33098 GND.n7058 GND.n7057 0.196152
R33099 GND.n7057 GND.n6737 0.196152
R33100 GND.n7050 GND.n6737 0.196152
R33101 GND.n7050 GND.n7049 0.196152
R33102 GND.n7049 GND.n6656 0.196152
R33103 GND.n7168 GND.n6656 0.196152
R33104 GND.n7283 GND.n7282 0.196152
R33105 GND.n7284 GND.n7283 0.196152
R33106 GND.n7284 GND.n2502 0.196152
R33107 GND.n7395 GND.n2502 0.196152
R33108 GND.n7396 GND.n7395 0.196152
R33109 GND.n7400 GND.n7396 0.196152
R33110 GND.n7400 GND.n7399 0.196152
R33111 GND.n7399 GND.n2475 0.196152
R33112 GND.n7433 GND.n2475 0.196152
R33113 GND.n2684 GND.n2642 0.196152
R33114 GND.n2684 GND.n2683 0.196152
R33115 GND.n2683 GND.n2643 0.196152
R33116 GND.n2675 GND.n2643 0.196152
R33117 GND.n2675 GND.n2674 0.196152
R33118 GND.n2674 GND.n2645 0.196152
R33119 GND.n2666 GND.n2645 0.196152
R33120 GND.n2666 GND.n2665 0.196152
R33121 GND.n6939 GND.n6925 0.196152
R33122 GND.n6931 GND.n6925 0.196152
R33123 GND.n6931 GND.n6930 0.196152
R33124 GND.n6930 GND.n6659 0.196152
R33125 GND.n7158 GND.n6659 0.196152
R33126 GND.n7159 GND.n7158 0.196152
R33127 GND.n7159 GND.n6657 0.196152
R33128 GND.n7166 GND.n6657 0.196152
R33129 GND.n7182 GND.n6641 0.196152
R33130 GND.n7076 GND.n6627 0.196152
R33131 GND.n7223 GND.n6615 0.196152
R33132 GND.n7224 GND.n7223 0.196152
R33133 GND.n7224 GND.n2552 0.196152
R33134 GND.n7314 GND.n2552 0.196152
R33135 GND.n7315 GND.n7314 0.196152
R33136 GND.n7316 GND.n7315 0.196152
R33137 GND.n7293 GND.n2565 0.196152
R33138 GND.n7303 GND.n2566 0.196152
R33139 GND.n7215 GND.n6626 0.196152
R33140 GND.n7238 GND.n2512 0.196152
R33141 GND.n7380 GND.n2512 0.196152
R33142 GND.n7381 GND.n7380 0.196152
R33143 GND.n7385 GND.n7381 0.196152
R33144 GND.n7385 GND.n7384 0.196152
R33145 GND.n7384 GND.n2484 0.196152
R33146 GND.n7424 GND.n2484 0.196152
R33147 GND.n7324 GND.n2541 0.196152
R33148 GND.n7008 GND.n7007 0.196152
R33149 GND.n7007 GND.n6668 0.196152
R33150 GND.n7146 GND.n6668 0.196152
R33151 GND.n7147 GND.n7146 0.196152
R33152 GND.n7150 GND.n7147 0.196152
R33153 GND.n7150 GND.n7149 0.196152
R33154 GND.n7149 GND.n6642 0.196152
R33155 GND.n7180 GND.n6642 0.196152
R33156 GND.n6978 GND.n6746 0.196152
R33157 GND.n7017 GND.n6746 0.196152
R33158 GND.n7018 GND.n7017 0.196152
R33159 GND.n7018 GND.n6743 0.196152
R33160 GND.n7026 GND.n6743 0.196152
R33161 GND.n7027 GND.n7026 0.196152
R33162 GND.n7040 GND.n7027 0.196152
R33163 GND.n7040 GND.n7039 0.196152
R33164 GND.n7039 GND.n7028 0.196152
R33165 GND.n9054 GND.n9053 0.193435
R33166 GND.n4766 GND.n4202 0.193435
R33167 GND.n7239 GND.n7238 0.193435
R33168 GND.n45 GND 0.191049
R33169 GND.n5669 GND.n5668 0.189724
R33170 GND.n9766 GND.n9765 0.189724
R33171 GND.n4936 GND.n2150 0.189724
R33172 GND.n9805 GND.n29 0.189608
R33173 GND.n8409 GND.n8399 0.189608
R33174 GND.n2294 GND.n2280 0.189561
R33175 GND.n2290 GND.n2282 0.189561
R33176 GND.n9828 GND.n3 0.189561
R33177 GND.n9831 GND.n9830 0.189561
R33178 GND.n44 GND.n31 0.189561
R33179 GND.n42 GND.n41 0.189561
R33180 GND.n5673 GND.n2278 0.189282
R33181 GND.n2287 GND.n2281 0.189062
R33182 GND.n2288 GND.n2284 0.189062
R33183 GND.n2293 GND.n2283 0.189062
R33184 GND.n2289 GND.n2288 0.189062
R33185 GND.n9827 GND.n0 0.189062
R33186 GND.n23 GND.n22 0.189062
R33187 GND.n4 GND.n0 0.189062
R33188 GND.n23 GND.n6 0.189062
R33189 GND.n34 GND.n30 0.189062
R33190 GND.n38 GND.n37 0.189062
R33191 GND.n35 GND.n34 0.189062
R33192 GND.n39 GND.n38 0.189062
R33193 GND.n6594 GND.n6589 0.188181
R33194 GND.n6580 GND.n6575 0.188181
R33195 GND.n6566 GND.n6561 0.188181
R33196 GND.n6552 GND.n6547 0.188181
R33197 GND.n6538 GND.n6533 0.188181
R33198 GND.n2704 GND.n2699 0.188181
R33199 GND.n6453 GND.n6448 0.188181
R33200 GND.n6467 GND.n6462 0.188181
R33201 GND.n6480 GND.n6475 0.188181
R33202 GND.n6493 GND.n6488 0.188181
R33203 GND.n6506 GND.n6501 0.188181
R33204 GND.n6519 GND.n6514 0.188181
R33205 GND.n6434 GND.n6429 0.188181
R33206 GND.n8957 GND.n8952 0.188181
R33207 GND.n8943 GND.n8938 0.188181
R33208 GND.n8929 GND.n8924 0.188181
R33209 GND.n8915 GND.n8910 0.188181
R33210 GND.n8901 GND.n8896 0.188181
R33211 GND.n987 GND.n982 0.188181
R33212 GND.n8817 GND.n8812 0.188181
R33213 GND.n8831 GND.n8826 0.188181
R33214 GND.n8844 GND.n8839 0.188181
R33215 GND.n8857 GND.n8852 0.188181
R33216 GND.n8870 GND.n8865 0.188181
R33217 GND.n8883 GND.n8878 0.188181
R33218 GND.n8798 GND.n8793 0.188181
R33219 GND.n4856 GND.n4851 0.188181
R33220 GND.n4842 GND.n4837 0.188181
R33221 GND.n4828 GND.n4823 0.188181
R33222 GND.n4814 GND.n4809 0.188181
R33223 GND.n4800 GND.n4795 0.188181
R33224 GND.n4785 GND.n4780 0.188181
R33225 GND.n4179 GND.n4174 0.188181
R33226 GND.n4873 GND.n4868 0.188181
R33227 GND.n4886 GND.n4881 0.188181
R33228 GND.n4899 GND.n4894 0.188181
R33229 GND.n4912 GND.n4907 0.188181
R33230 GND.n4925 GND.n4920 0.188181
R33231 GND.n4160 GND.n4155 0.188181
R33232 GND.n5677 GND.n5673 0.188144
R33233 GND.n9773 GND.n29 0.188144
R33234 GND.n8399 GND.n1811 0.188144
R33235 GND.n5676 GND.n5670 0.185301
R33236 GND.n5681 GND.n5440 0.185301
R33237 GND.n5683 GND.n5682 0.185301
R33238 GND.n9772 GND.n9767 0.185301
R33239 GND.n9777 GND.n58 0.185301
R33240 GND.n9779 GND.n9778 0.185301
R33241 GND.n8416 GND.n8415 0.185301
R33242 GND.n4938 GND.n4937 0.185301
R33243 GND.n4935 GND.n1809 0.185301
R33244 GND.n1456 GND.n1455 0.185134
R33245 GND.n2936 GND.n2935 0.161919
R33246 GND.n6595 GND.n6594 0.158954
R33247 GND.n6581 GND.n6580 0.158954
R33248 GND.n6567 GND.n6566 0.158954
R33249 GND.n6553 GND.n6552 0.158954
R33250 GND.n6539 GND.n6538 0.158954
R33251 GND.n2705 GND.n2704 0.158954
R33252 GND.n6454 GND.n6453 0.158954
R33253 GND.n6468 GND.n6467 0.158954
R33254 GND.n6481 GND.n6480 0.158954
R33255 GND.n6494 GND.n6493 0.158954
R33256 GND.n6507 GND.n6506 0.158954
R33257 GND.n6520 GND.n6519 0.158954
R33258 GND.n6435 GND.n6434 0.158954
R33259 GND.n8958 GND.n8957 0.158954
R33260 GND.n8944 GND.n8943 0.158954
R33261 GND.n8930 GND.n8929 0.158954
R33262 GND.n8916 GND.n8915 0.158954
R33263 GND.n8902 GND.n8901 0.158954
R33264 GND.n988 GND.n987 0.158954
R33265 GND.n8818 GND.n8817 0.158954
R33266 GND.n8832 GND.n8831 0.158954
R33267 GND.n8845 GND.n8844 0.158954
R33268 GND.n8858 GND.n8857 0.158954
R33269 GND.n8871 GND.n8870 0.158954
R33270 GND.n8884 GND.n8883 0.158954
R33271 GND.n8799 GND.n8798 0.158954
R33272 GND.n4857 GND.n4856 0.158954
R33273 GND.n4843 GND.n4842 0.158954
R33274 GND.n4829 GND.n4828 0.158954
R33275 GND.n4815 GND.n4814 0.158954
R33276 GND.n4801 GND.n4800 0.158954
R33277 GND.n4786 GND.n4785 0.158954
R33278 GND.n4180 GND.n4179 0.158954
R33279 GND.n4874 GND.n4873 0.158954
R33280 GND.n4887 GND.n4886 0.158954
R33281 GND.n4900 GND.n4899 0.158954
R33282 GND.n4913 GND.n4912 0.158954
R33283 GND.n4926 GND.n4925 0.158954
R33284 GND.n4161 GND.n4160 0.158954
R33285 GND.n9512 GND.t247 0.154832
R33286 GND.n9589 GND.n160 0.154832
R33287 GND.n9750 GND.n9749 0.154832
R33288 GND.n154 GND.n153 0.154832
R33289 GND.n9759 GND.n66 0.154832
R33290 GND.n9742 GND.n82 0.154832
R33291 GND.n9710 GND.n103 0.154832
R33292 GND.t264 GND.n9687 0.154832
R33293 GND.n7807 GND.t196 0.154832
R33294 GND.n7873 GND.n2215 0.154832
R33295 GND.n7883 GND.n7882 0.154832
R33296 GND.n7970 GND.n7969 0.154832
R33297 GND.n7856 GND.n2253 0.154832
R33298 GND.n7963 GND.n2166 0.154832
R33299 GND.n7931 GND.n2186 0.154832
R33300 GND.t185 GND.n2133 0.154832
R33301 GND.n43 GND.n24 0.145891
R33302 GND.n1456 GND.n980 0.144344
R33303 GND.n7273 GND.n7259 0.140424
R33304 GND.n883 GND.n882 0.140424
R33305 GND.n4538 GND.n4533 0.140424
R33306 GND.n9829 GND.n7 0.135741
R33307 GND.n897 GND.n873 0.131508
R33308 GND.n4532 GND.n4531 0.131508
R33309 GND.n7032 GND.n7028 0.131508
R33310 GND.n5435 GND.n5434 0.1285
R33311 GND.n1465 GND.n1463 0.1285
R33312 GND.n3508 GND.n3506 0.1285
R33313 GND.n9041 GND.n9040 0.128217
R33314 GND.n4657 GND.n4656 0.128217
R33315 GND.n7282 GND.n2622 0.128217
R33316 GND.n944 GND.n943 0.117348
R33317 GND.n4678 GND.n4677 0.117348
R33318 GND.n7168 GND.n7167 0.117348
R33319 GND.n3106 GND.n3105 0.112479
R33320 GND.n5680 GND.n5679 0.110167
R33321 GND.n9776 GND.n9775 0.110167
R33322 GND.n8414 GND.n1813 0.110167
R33323 GND.n3105 GND 0.106269
R33324 GND.n5133 GND.n5047 0.1029
R33325 GND.n1596 GND.n1213 0.1029
R33326 GND.n3639 GND.n3259 0.1029
R33327 GND.n6573 GND.n6559 0.0910185
R33328 GND.n6587 GND.n6573 0.0910185
R33329 GND.n6526 GND.n6513 0.0910185
R33330 GND.n6500 GND.n6487 0.0910185
R33331 GND.n6487 GND.n6474 0.0910185
R33332 GND.n8936 GND.n8922 0.0910185
R33333 GND.n8950 GND.n8936 0.0910185
R33334 GND.n8890 GND.n8877 0.0910185
R33335 GND.n8864 GND.n8851 0.0910185
R33336 GND.n8851 GND.n8838 0.0910185
R33337 GND.n4835 GND.n4821 0.0910185
R33338 GND.n4849 GND.n4835 0.0910185
R33339 GND.n4932 GND.n4919 0.0910185
R33340 GND.n4906 GND.n4893 0.0910185
R33341 GND.n4893 GND.n4880 0.0910185
R33342 GND.n7731 GND.n7730 0.0900158
R33343 GND.n5675 GND.n2279 0.0900158
R33344 GND.n9804 GND.n47 0.0900158
R33345 GND.n9771 GND.n57 0.0900158
R33346 GND.n8408 GND.n8401 0.0900158
R33347 GND.n8417 GND.n1808 0.0900158
R33348 GND.n6559 GND.n6545 0.0892778
R33349 GND.n6513 GND.n6500 0.0892778
R33350 GND.n8922 GND.n8908 0.0892778
R33351 GND.n8877 GND.n8864 0.0892778
R33352 GND.n4821 GND.n4807 0.0892778
R33353 GND.n4919 GND.n4906 0.0892778
R33354 GND.n5685 GND.n5684 0.0863711
R33355 GND.n9781 GND.n9780 0.0863711
R33356 GND.n8421 GND.n8420 0.0863711
R33357 GND.n2293 GND.n7 0.0755085
R33358 GND.n7698 GND.n7697 0.0755
R33359 GND.n9824 GND.n10 0.0755
R33360 GND.n5013 GND.n5012 0.0719286
R33361 GND.n5436 GND.n5012 0.0719286
R33362 GND.n5691 GND.n5006 0.0719286
R33363 GND.n5691 GND.n5690 0.0719286
R33364 GND.n6354 GND.n6328 0.0719286
R33365 GND.n6350 GND.n6328 0.0719286
R33366 GND.n6339 GND.n2716 0.0719286
R33367 GND.n6423 GND.n2716 0.0719286
R33368 GND.n8518 GND.n999 0.0719286
R33369 GND.n8787 GND.n999 0.0719286
R33370 GND.n1443 GND.n1363 0.0719286
R33371 GND.n1462 GND.n1363 0.0719286
R33372 GND.n1434 GND.n1368 0.0719286
R33373 GND.n1452 GND.n1368 0.0719286
R33374 GND.n8531 GND.n8512 0.0719286
R33375 GND.n8527 GND.n8512 0.0719286
R33376 GND.n3490 GND.n3410 0.0719286
R33377 GND.n3505 GND.n3410 0.0719286
R33378 GND.n3481 GND.n3415 0.0719286
R33379 GND.n3499 GND.n3415 0.0719286
R33380 GND.n4945 GND.n3930 0.0719286
R33381 GND.n4945 GND.n4944 0.0719286
R33382 GND.n3937 GND.n3936 0.0719286
R33383 GND.n4150 GND.n3936 0.0719286
R33384 GND.n5668 GND.n5441 0.071
R33385 GND.n9765 GND.n59 0.071
R33386 GND.n7976 GND.n2150 0.071
R33387 GND.n7731 GND.n2278 0.0703691
R33388 GND.n9805 GND.n9804 0.0698941
R33389 GND.n8409 GND.n8408 0.0698941
R33390 GND.n9782 GND.n9781 0.0694333
R33391 GND.n8422 GND.n8421 0.0689437
R33392 GND.n24 GND.n23 0.0682585
R33393 GND.n8967 GND.n979 0.0617955
R33394 GND.n4778 GND.n4187 0.0617955
R33395 GND.n6605 GND.n6604 0.0617955
R33396 GND.n5440 GND.n5439 0.0610133
R33397 GND.n995 GND.n58 0.0610133
R33398 GND.n4939 GND.n4938 0.0610133
R33399 GND.n2938 GND.n2932 0.0593235
R33400 GND.n2946 GND.n2945 0.0593235
R33401 GND.n2949 GND.n2930 0.0593235
R33402 GND.n2952 GND.n2927 0.0593235
R33403 GND.n2995 GND.n2957 0.0593235
R33404 GND.n2994 GND.n2993 0.0593235
R33405 GND.n2989 GND.n2958 0.0593235
R33406 GND.n2985 GND.n2984 0.0593235
R33407 GND.n2981 GND.n2966 0.0593235
R33408 GND.n2980 GND.n2968 0.0593235
R33409 GND.n2972 GND.n2921 0.0593235
R33410 GND.n3004 GND.n3003 0.0593235
R33411 GND.n3005 GND.n2918 0.0593235
R33412 GND.n3012 GND.n3010 0.0593235
R33413 GND.n3023 GND.n3022 0.0593235
R33414 GND.n3027 GND.n2911 0.0593235
R33415 GND.n3029 GND.n3028 0.0593235
R33416 GND.n3030 GND.n2908 0.0593235
R33417 GND.n3076 GND.n3035 0.0593235
R33418 GND.n3075 GND.n3074 0.0593235
R33419 GND.n3071 GND.n3036 0.0593235
R33420 GND.n3063 GND.n3044 0.0593235
R33421 GND.n3062 GND.n3049 0.0593235
R33422 GND.n3059 GND.n3058 0.0593235
R33423 GND.n3054 GND.n3051 0.0593235
R33424 GND.n3083 GND.n2902 0.0593235
R33425 GND.n3086 GND.n3084 0.0593235
R33426 GND.n3085 GND.n2898 0.0593235
R33427 GND.n3099 GND.n2896 0.0593235
R33428 GND.n3100 GND.n2894 0.0593235
R33429 GND.n5684 GND.n5683 0.0586933
R33430 GND.n9780 GND.n9779 0.0586933
R33431 GND.n8420 GND.n1809 0.0586933
R33432 GND.n7728 GND 0.0541248
R33433 GND GND.n2914 0.0499652
R33434 GND GND.n3066 0.0499652
R33435 GND.n6531 GND.n2711 0.0457593
R33436 GND.n6545 GND.n6531 0.0457593
R33437 GND.n6602 GND.n6601 0.0457593
R33438 GND.n6527 GND.n6526 0.0457593
R33439 GND.n6461 GND.n6460 0.0457593
R33440 GND.n8894 GND.n994 0.0457593
R33441 GND.n8908 GND.n8894 0.0457593
R33442 GND.n8965 GND.n8964 0.0457593
R33443 GND.n8891 GND.n8890 0.0457593
R33444 GND.n8825 GND.n8824 0.0457593
R33445 GND.n4793 GND.n4792 0.0457593
R33446 GND.n4807 GND.n4793 0.0457593
R33447 GND.n4864 GND.n4863 0.0457593
R33448 GND.n4933 GND.n4932 0.0457593
R33449 GND.n4867 GND.n4186 0.0457593
R33450 GND.n6602 GND.n6587 0.0440185
R33451 GND.n6527 GND.n6441 0.0440185
R33452 GND.n6474 GND.n6461 0.0440185
R33453 GND.n8965 GND.n8950 0.0440185
R33454 GND.n8891 GND.n8805 0.0440185
R33455 GND.n8838 GND.n8825 0.0440185
R33456 GND.n4864 GND.n4849 0.0440185
R33457 GND.n4933 GND.n4167 0.0440185
R33458 GND.n4880 GND.n4867 0.0440185
R33459 GND.n5630 GND.n5629 0.0433385
R33460 GND.n9604 GND.n9603 0.0433385
R33461 GND.n7977 GND.n2149 0.0433385
R33462 GND GND.n5675 0.0430057
R33463 GND GND.n9771 0.0430057
R33464 GND.n8417 GND 0.0430057
R33465 GND.n5656 GND.n5458 0.0429107
R33466 GND.n9569 GND.n71 0.0429107
R33467 GND.n7975 GND.n2151 0.0429107
R33468 GND.n5011 GND.n5010 0.0421667
R33469 GND.n5437 GND.n5011 0.0421667
R33470 GND.n5009 GND.n5007 0.0421667
R33471 GND.n5689 GND.n5007 0.0421667
R33472 GND.n6353 GND.n6352 0.0421667
R33473 GND.n6352 GND.n6351 0.0421667
R33474 GND.n2715 GND.n2714 0.0421667
R33475 GND.n6424 GND.n2715 0.0421667
R33476 GND.n998 GND.n997 0.0421667
R33477 GND.n8788 GND.n998 0.0421667
R33478 GND.n1365 GND.n1364 0.0421667
R33479 GND.n1461 GND.n1364 0.0421667
R33480 GND.n1367 GND.n1366 0.0421667
R33481 GND.n1453 GND.n1367 0.0421667
R33482 GND.n8530 GND.n8529 0.0421667
R33483 GND.n8529 GND.n8528 0.0421667
R33484 GND.n3412 GND.n3411 0.0421667
R33485 GND.n3504 GND.n3411 0.0421667
R33486 GND.n3414 GND.n3413 0.0421667
R33487 GND.n3500 GND.n3414 0.0421667
R33488 GND.n3933 GND.n3931 0.0421667
R33489 GND.n4943 GND.n3931 0.0421667
R33490 GND.n3935 GND.n3934 0.0421667
R33491 GND.n4151 GND.n3935 0.0421667
R33492 GND.n6600 GND.n6589 0.0407778
R33493 GND.n6586 GND.n6575 0.0407778
R33494 GND.n6572 GND.n6561 0.0407778
R33495 GND.n6558 GND.n6547 0.0407778
R33496 GND.n6544 GND.n6533 0.0407778
R33497 GND.n2710 GND.n2699 0.0407778
R33498 GND.n6459 GND.n6448 0.0407778
R33499 GND.n6473 GND.n6462 0.0407778
R33500 GND.n6486 GND.n6475 0.0407778
R33501 GND.n6499 GND.n6488 0.0407778
R33502 GND.n6512 GND.n6501 0.0407778
R33503 GND.n6525 GND.n6514 0.0407778
R33504 GND.n6440 GND.n6429 0.0407778
R33505 GND.n8963 GND.n8952 0.0407778
R33506 GND.n8949 GND.n8938 0.0407778
R33507 GND.n8935 GND.n8924 0.0407778
R33508 GND.n8921 GND.n8910 0.0407778
R33509 GND.n8907 GND.n8896 0.0407778
R33510 GND.n993 GND.n982 0.0407778
R33511 GND.n8823 GND.n8812 0.0407778
R33512 GND.n8837 GND.n8826 0.0407778
R33513 GND.n8850 GND.n8839 0.0407778
R33514 GND.n8863 GND.n8852 0.0407778
R33515 GND.n8876 GND.n8865 0.0407778
R33516 GND.n8889 GND.n8878 0.0407778
R33517 GND.n8804 GND.n8793 0.0407778
R33518 GND.n4862 GND.n4851 0.0407778
R33519 GND.n4848 GND.n4837 0.0407778
R33520 GND.n4834 GND.n4823 0.0407778
R33521 GND.n4820 GND.n4809 0.0407778
R33522 GND.n4806 GND.n4795 0.0407778
R33523 GND.n4791 GND.n4780 0.0407778
R33524 GND.n4185 GND.n4174 0.0407778
R33525 GND.n4879 GND.n4868 0.0407778
R33526 GND.n4892 GND.n4881 0.0407778
R33527 GND.n4905 GND.n4894 0.0407778
R33528 GND.n4918 GND.n4907 0.0407778
R33529 GND.n4931 GND.n4920 0.0407778
R33530 GND.n4166 GND.n4155 0.0407778
R33531 GND.n5458 GND.n5457 0.0384464
R33532 GND.n9755 GND.n71 0.0384464
R33533 GND.n7975 GND.n7974 0.0384464
R33534 GND.n8401 GND.n8400 0.0358479
R33535 GND.n897 GND.n896 0.0356562
R33536 GND.n883 GND.n879 0.0356562
R33537 GND.n4668 GND.n4532 0.0356562
R33538 GND.n4666 GND.n4533 0.0356562
R33539 GND.n7032 GND.n7031 0.0356562
R33540 GND.n7259 GND.n7258 0.0356562
R33541 GND.n957 GND.n263 0.0351154
R33542 GND.n4691 GND.n1955 0.0351154
R33543 GND.n7213 GND.n7210 0.0351154
R33544 GND.n978 GND.n977 0.0346346
R33545 GND.n4709 GND.n4696 0.0346346
R33546 GND.n7305 GND.n2563 0.0346346
R33547 GND.n3104 GND 0.0341538
R33548 GND.n47 GND.n46 0.0338896
R33549 GND.n57 GND.n47 0.0337917
R33550 GND.n8401 GND.n1808 0.0337917
R33551 GND.n7730 GND.n2279 0.0337917
R33552 GND.n977 GND.n976 0.0336731
R33553 GND.n4709 GND.n4708 0.0336731
R33554 GND.n7305 GND.n7304 0.0336731
R33555 GND.n9026 GND.n459 0.0331923
R33556 GND.n9052 GND.n443 0.0331923
R33557 GND.n4717 GND.n4206 0.0331923
R33558 GND.n4767 GND.n4201 0.0331923
R33559 GND.n7187 GND.n7186 0.0331923
R33560 GND.n7240 GND.n7235 0.0331923
R33561 GND.n957 GND.n956 0.0327115
R33562 GND.n461 GND.n460 0.0327115
R33563 GND.n4691 GND.n4690 0.0327115
R33564 GND.n4719 GND.n4718 0.0327115
R33565 GND.n7214 GND.n7213 0.0327115
R33566 GND.n6606 GND.n2694 0.0327115
R33567 GND.n9781 GND.n57 0.0318333
R33568 GND.n8421 GND.n1808 0.0318333
R33569 GND.n5685 GND.n2279 0.0318333
R33570 GND.n2937 GND.n2936 0.0312487
R33571 GND.n2965 GND 0.0312487
R33572 GND.n844 GND.n825 0.0307885
R33573 GND.n4486 GND.n4485 0.0307885
R33574 GND.n7181 GND.n6639 0.0307885
R33575 GND.n2951 GND 0.0285749
R33576 GND GND.n2975 0.0285749
R33577 GND.n3017 GND 0.0285749
R33578 GND.n3043 GND 0.0285749
R33579 GND.n3094 GND 0.0285749
R33580 GND.n943 GND.n941 0.0249565
R33581 GND.n844 GND.n843 0.0249565
R33582 GND.n9040 GND.n453 0.0249565
R33583 GND.n4677 GND.n4222 0.0249565
R33584 GND.n4485 GND.n4484 0.0249565
R33585 GND.n4656 GND.n4653 0.0249565
R33586 GND.n2642 GND.n2622 0.0249565
R33587 GND.n7167 GND.n7166 0.0249565
R33588 GND.n7181 GND.n7180 0.0249565
R33589 GND.n5682 GND.n5681 0.0242951
R33590 GND.n9778 GND.n9777 0.0242951
R33591 GND.n4937 GND.n4935 0.0242951
R33592 GND.n5673 GND.n5672 0.024
R33593 GND.n9769 GND.n29 0.024
R33594 GND.n8399 GND.n1812 0.024
R33595 GND.n3106 GND 0.0226354
R33596 GND.n45 GND.n44 0.0221396
R33597 GND.n7729 GND 0.0210625
R33598 GND.n5676 GND 0.0203443
R33599 GND.n9772 GND 0.0203443
R33600 GND GND.n8416 0.0203443
R33601 GND.n5629 GND.n5441 0.0191042
R33602 GND.n9604 GND.n59 0.0191042
R33603 GND.n7977 GND.n7976 0.0191042
R33604 GND.n7730 GND.n7729 0.0191042
R33605 GND.n879 GND.n875 0.0190547
R33606 GND.n4667 GND.n4666 0.0190547
R33607 GND.n7258 GND.n2629 0.0190547
R33608 GND.n8970 GND.n470 0.0187692
R33609 GND.n8969 GND.n454 0.0187692
R33610 GND.n9039 GND.n9038 0.0187692
R33611 GND.n4223 GND.n4189 0.0187692
R33612 GND.n4776 GND.n4190 0.0187692
R33613 GND.n4655 GND.n4654 0.0187692
R33614 GND.n7197 GND.n7196 0.0187692
R33615 GND.n7249 GND.n2635 0.0187692
R33616 GND.n7248 GND.n2636 0.0187692
R33617 GND.n896 GND.n875 0.0171016
R33618 GND.n4668 GND.n4667 0.0171016
R33619 GND.n7031 GND.n2629 0.0171016
R33620 GND.n942 GND.n470 0.0168462
R33621 GND.n8970 GND.n8969 0.0168462
R33622 GND.n9038 GND.n454 0.0168462
R33623 GND.n4676 GND.n4223 0.0168462
R33624 GND.n4776 GND.n4189 0.0168462
R33625 GND.n4654 GND.n4190 0.0168462
R33626 GND.n7196 GND.n6633 0.0168462
R33627 GND.n7197 GND.n2635 0.0168462
R33628 GND.n7249 GND.n7248 0.0168462
R33629 GND.n1457 GND.n1456 0.0168125
R33630 GND.n8893 GND.n471 0.0165676
R33631 GND.n8967 GND.n8966 0.0165676
R33632 GND.n4188 GND.n4153 0.0165676
R33633 GND.n4865 GND.n4778 0.0165676
R33634 GND.n6530 GND.n6529 0.0165676
R33635 GND.n6604 GND.n6603 0.0165676
R33636 GND.n943 GND.n942 0.0144423
R33637 GND.n4677 GND.n4676 0.0144423
R33638 GND.n7167 GND.n6633 0.0144423
R33639 GND.n845 GND.n844 0.014087
R33640 GND.n956 GND.n241 0.014087
R33641 GND.n956 GND.n955 0.014087
R33642 GND.n4485 GND.n4256 0.014087
R33643 GND.n4690 GND.n1933 0.014087
R33644 GND.n4690 GND.n4689 0.014087
R33645 GND.n7182 GND.n7181 0.014087
R33646 GND.n7214 GND.n6627 0.014087
R33647 GND.n7215 GND.n7214 0.014087
R33648 GND.n1455 GND.n56 0.0127323
R33649 GND.n1458 GND.n1455 0.0127323
R33650 GND.n9040 GND.n9039 0.0125192
R33651 GND.n4656 GND.n4655 0.0125192
R33652 GND.n2636 GND.n2622 0.0125192
R33653 GND.n5682 GND.n5680 0.0123976
R33654 GND.n5672 GND.n5670 0.0123976
R33655 GND.n5679 GND.n5670 0.0123976
R33656 GND.n5681 GND.n5669 0.0123976
R33657 GND.n9778 GND.n9776 0.0123976
R33658 GND.n9769 GND.n9767 0.0123976
R33659 GND.n9775 GND.n9767 0.0123976
R33660 GND.n9777 GND.n9766 0.0123976
R33661 GND.n4935 GND.n1813 0.0123976
R33662 GND.n8415 GND.n1812 0.0123976
R33663 GND.n8415 GND.n8414 0.0123976
R33664 GND.n4937 GND.n4936 0.0123976
R33665 GND.n9826 GND.n8 0.0123479
R33666 GND.n7727 GND.n2294 0.01225
R33667 GND GND.n3102 0.0118636
R33668 GND.n3103 GND 0.0118636
R33669 GND.n5683 GND.n5440 0.0113267
R33670 GND.n9779 GND.n58 0.0113267
R33671 GND.n4938 GND.n1809 0.0113267
R33672 GND GND.n2950 0.0111952
R33673 GND.n2976 GND 0.0111952
R33674 GND.n3070 GND 0.0111952
R33675 GND GND.n3093 0.0111952
R33676 GND.n9828 GND.n9826 0.0102917
R33677 GND.n7728 GND.n7727 0.0102917
R33678 GND.n6595 GND.n6588 0.0102222
R33679 GND.n6581 GND.n6574 0.0102222
R33680 GND.n6567 GND.n6560 0.0102222
R33681 GND.n6553 GND.n6546 0.0102222
R33682 GND.n6539 GND.n6532 0.0102222
R33683 GND.n2705 GND.n2698 0.0102222
R33684 GND.n6454 GND.n6447 0.0102222
R33685 GND.n6468 GND.n6446 0.0102222
R33686 GND.n6481 GND.n6445 0.0102222
R33687 GND.n6494 GND.n6444 0.0102222
R33688 GND.n6507 GND.n6443 0.0102222
R33689 GND.n6520 GND.n6442 0.0102222
R33690 GND.n6435 GND.n6428 0.0102222
R33691 GND.n8958 GND.n8951 0.0102222
R33692 GND.n8944 GND.n8937 0.0102222
R33693 GND.n8930 GND.n8923 0.0102222
R33694 GND.n8916 GND.n8909 0.0102222
R33695 GND.n8902 GND.n8895 0.0102222
R33696 GND.n988 GND.n981 0.0102222
R33697 GND.n8818 GND.n8811 0.0102222
R33698 GND.n8832 GND.n8810 0.0102222
R33699 GND.n8845 GND.n8809 0.0102222
R33700 GND.n8858 GND.n8808 0.0102222
R33701 GND.n8871 GND.n8807 0.0102222
R33702 GND.n8884 GND.n8806 0.0102222
R33703 GND.n8799 GND.n8792 0.0102222
R33704 GND.n4857 GND.n4850 0.0102222
R33705 GND.n4843 GND.n4836 0.0102222
R33706 GND.n4829 GND.n4822 0.0102222
R33707 GND.n4815 GND.n4808 0.0102222
R33708 GND.n4801 GND.n4794 0.0102222
R33709 GND.n4786 GND.n4779 0.0102222
R33710 GND.n4180 GND.n4173 0.0102222
R33711 GND.n4874 GND.n4172 0.0102222
R33712 GND.n4887 GND.n4171 0.0102222
R33713 GND.n4900 GND.n4170 0.0102222
R33714 GND.n4913 GND.n4169 0.0102222
R33715 GND.n4926 GND.n4168 0.0102222
R33716 GND.n4161 GND.n4154 0.0102222
R33717 GND.n3018 GND 0.00985829
R33718 GND.n3067 GND 0.00985829
R33719 GND.n38 GND 0.0092
R33720 GND.n976 GND.n283 0.00865217
R33721 GND.n976 GND.n975 0.00865217
R33722 GND.n9053 GND.n442 0.00865217
R33723 GND.n4708 GND.n1975 0.00865217
R33724 GND.n4708 GND.n4707 0.00865217
R33725 GND.n4766 GND.n4765 0.00865217
R33726 GND.n7304 GND.n2565 0.00865217
R33727 GND.n7304 GND.n7303 0.00865217
R33728 GND.n7239 GND.n2541 0.00865217
R33729 GND.n2988 GND 0.00852139
R33730 GND.n3011 GND 0.00852139
R33731 GND GND.n3103 0.00852139
R33732 GND.n5677 GND.n5676 0.0067128
R33733 GND.n5678 GND.n5677 0.0067128
R33734 GND.n9773 GND.n9772 0.0067128
R33735 GND.n9774 GND.n9773 0.0067128
R33736 GND.n8416 GND.n1811 0.0067128
R33737 GND.n8413 GND.n1811 0.0067128
R33738 GND.n2288 GND.n2287 0.0063
R33739 GND.n43 GND.n34 0.0063
R33740 GND.n46 GND 0.00627708
R33741 GND.n5667 GND.n5666 0.00570833
R33742 GND.n9764 GND.n9763 0.00570833
R33743 GND.n7889 GND.n2204 0.00570833
R33744 GND.n3105 GND.n3104 0.00530769
R33745 GND.n5631 GND.n5485 0.00496429
R33746 GND.n5528 GND.n5527 0.00496429
R33747 GND.n9725 GND.n101 0.00496429
R33748 GND.n9602 GND.n9601 0.00496429
R33749 GND.n7946 GND.n2184 0.00496429
R33750 GND.n2243 GND.n2242 0.00496429
R33751 GND.n33 GND.n30 0.00487671
R33752 GND.n37 GND.n36 0.00487671
R33753 GND.n35 GND.n32 0.00487671
R33754 GND.n42 GND.n39 0.00487671
R33755 GND.n9827 GND.n2 0.00487671
R33756 GND.n22 GND.n5 0.00487671
R33757 GND.n4 GND.n1 0.00487671
R33758 GND.n9831 GND.n6 0.00487671
R33759 GND.n2292 GND.n2281 0.00487671
R33760 GND.n2286 GND.n2284 0.00487671
R33761 GND.n2285 GND.n2283 0.00487671
R33762 GND.n2290 GND.n2289 0.00487671
R33763 GND.n2294 GND.n2281 0.00487671
R33764 GND.n2292 GND.n2284 0.00487671
R33765 GND.n2286 GND.n2283 0.00487671
R33766 GND.n2289 GND.n2285 0.00487671
R33767 GND.n9828 GND.n9827 0.00487671
R33768 GND.n22 GND.n2 0.00487671
R33769 GND.n5 GND.n4 0.00487671
R33770 GND.n6 GND.n1 0.00487671
R33771 GND.n44 GND.n30 0.00487671
R33772 GND.n37 GND.n33 0.00487671
R33773 GND.n36 GND.n35 0.00487671
R33774 GND.n39 GND.n32 0.00487671
R33775 GND GND.n0 0.00485
R33776 GND.n8893 GND.n8892 0.00457568
R33777 GND.n8966 GND.n980 0.00457568
R33778 GND.n4934 GND.n4153 0.00457568
R33779 GND.n4866 GND.n4865 0.00457568
R33780 GND.n6530 GND.n6528 0.00457568
R33781 GND.n6603 GND.n2697 0.00457568
R33782 GND.n8400 GND 0.00431875
R33783 GND.n2296 GND.n2295 0.00425
R33784 GND.n2291 GND.n2280 0.00387804
R33785 GND.n2293 GND.n2282 0.00387804
R33786 GND.n9830 GND.n0 0.00387804
R33787 GND.n23 GND.n3 0.00387804
R33788 GND.n41 GND.n40 0.00387804
R33789 GND.n38 GND.n31 0.00387804
R33790 GND.n2288 GND.n2280 0.00387804
R33791 GND.n2287 GND.n2282 0.00387804
R33792 GND.n9832 GND.n3 0.00387804
R33793 GND.n9830 GND.n9829 0.00387804
R33794 GND.n40 GND.n31 0.00387804
R33795 GND.n41 GND.n34 0.00387804
R33796 GND.n2938 GND.n2937 0.0031738
R33797 GND.n2945 GND.n2932 0.0031738
R33798 GND.n2946 GND.n2930 0.0031738
R33799 GND.n2950 GND.n2949 0.0031738
R33800 GND.n2952 GND.n2951 0.0031738
R33801 GND.n2957 GND.n2927 0.0031738
R33802 GND.n2995 GND.n2994 0.0031738
R33803 GND.n2993 GND.n2958 0.0031738
R33804 GND.n2989 GND.n2988 0.0031738
R33805 GND.n2985 GND.n2965 0.0031738
R33806 GND.n2984 GND.n2966 0.0031738
R33807 GND.n2981 GND.n2980 0.0031738
R33808 GND.n2976 GND.n2968 0.0031738
R33809 GND.n2975 GND.n2972 0.0031738
R33810 GND.n3003 GND.n2921 0.0031738
R33811 GND.n3005 GND.n3004 0.0031738
R33812 GND.n3010 GND.n2918 0.0031738
R33813 GND.n3012 GND.n3011 0.0031738
R33814 GND.n3018 GND.n3017 0.0031738
R33815 GND.n3022 GND.n2914 0.0031738
R33816 GND.n3023 GND.n2911 0.0031738
R33817 GND.n3028 GND.n3027 0.0031738
R33818 GND.n3030 GND.n3029 0.0031738
R33819 GND.n3035 GND.n2908 0.0031738
R33820 GND.n3076 GND.n3075 0.0031738
R33821 GND.n3074 GND.n3036 0.0031738
R33822 GND.n3071 GND.n3070 0.0031738
R33823 GND.n3067 GND.n3043 0.0031738
R33824 GND.n3066 GND.n3044 0.0031738
R33825 GND.n3063 GND.n3062 0.0031738
R33826 GND.n3059 GND.n3049 0.0031738
R33827 GND.n3058 GND.n3051 0.0031738
R33828 GND.n3054 GND.n2902 0.0031738
R33829 GND.n3084 GND.n3083 0.0031738
R33830 GND.n3086 GND.n3085 0.0031738
R33831 GND.n3093 GND.n2898 0.0031738
R33832 GND.n3094 GND.n2896 0.0031738
R33833 GND.n3100 GND.n3099 0.0031738
R33834 GND.n3102 GND.n2894 0.0031738
R33835 GND.n825 GND.n459 0.00242308
R33836 GND.n9026 GND.n9025 0.00242308
R33837 GND.n460 GND.n443 0.00242308
R33838 GND.n4486 GND.n4206 0.00242308
R33839 GND.n4720 GND.n4717 0.00242308
R33840 GND.n4718 GND.n4201 0.00242308
R33841 GND.n7186 GND.n6639 0.00242308
R33842 GND.n7187 GND.n6607 0.00242308
R33843 GND.n7235 GND.n2694 0.00242308
R33844 GND GND.n9832 0.00195
R33845 GND.n8400 GND.n8 0.0014641
R33846 GND.n46 GND.n45 0.00113729
R33847 GND.n978 GND.n263 0.000980769
R33848 GND.n9025 GND.n461 0.000980769
R33849 GND.n9053 GND.n9052 0.000980769
R33850 GND.n4696 GND.n1955 0.000980769
R33851 GND.n4720 GND.n4719 0.000980769
R33852 GND.n4767 GND.n4766 0.000980769
R33853 GND.n7210 GND.n2563 0.000980769
R33854 GND.n6607 GND.n6606 0.000980769
R33855 GND.n7240 GND.n7239 0.000980769
R33856 GND.n7729 GND.n7728 0.000589524
R33857 GND.n8968 GND.n471 0.000578378
R33858 GND.n8968 GND.n8967 0.000578378
R33859 GND.n4777 GND.n4188 0.000578378
R33860 GND.n4778 GND.n4777 0.000578378
R33861 GND.n6529 GND.n2696 0.000578378
R33862 GND.n6604 GND.n2696 0.000578378
R33863 1Bit_Clk_ADC_0.x3.B.n41 1Bit_Clk_ADC_0.x3.B.n40 256.104
R33864 1Bit_Clk_ADC_0.x3.B.n45 1Bit_Clk_ADC_0.x3.B.n44 243.68
R33865 1Bit_Clk_ADC_0.x3.B.n3 1Bit_Clk_ADC_0.x3.B.n1 241.847
R33866 1Bit_Clk_ADC_0.x3.B.n4 1Bit_Clk_ADC_0.x3.B.t21 212.081
R33867 1Bit_Clk_ADC_0.x3.B.n11 1Bit_Clk_ADC_0.x3.B.t35 212.081
R33868 1Bit_Clk_ADC_0.x3.B.n5 1Bit_Clk_ADC_0.x3.B.t28 212.081
R33869 1Bit_Clk_ADC_0.x3.B.n6 1Bit_Clk_ADC_0.x3.B.t14 212.081
R33870 1Bit_Clk_ADC_0.x3.B.n25 1Bit_Clk_ADC_0.x3.B.t31 212.081
R33871 1Bit_Clk_ADC_0.x3.B.n24 1Bit_Clk_ADC_0.x3.B.t25 212.081
R33872 1Bit_Clk_ADC_0.x3.B.n30 1Bit_Clk_ADC_0.x3.B.t15 212.081
R33873 1Bit_Clk_ADC_0.x3.B.n32 1Bit_Clk_ADC_0.x3.B.t30 212.081
R33874 1Bit_Clk_ADC_0.x3.B.n16 1Bit_Clk_ADC_0.x3.B.t20 212.081
R33875 1Bit_Clk_ADC_0.x3.B.n18 1Bit_Clk_ADC_0.x3.B.t17 212.081
R33876 1Bit_Clk_ADC_0.x3.B.n15 1Bit_Clk_ADC_0.x3.B.t18 212.081
R33877 1Bit_Clk_ADC_0.x3.B.n23 1Bit_Clk_ADC_0.x3.B.t12 212.081
R33878 1Bit_Clk_ADC_0.x3.B.n45 1Bit_Clk_ADC_0.x3.B.n43 205.28
R33879 1Bit_Clk_ADC_0.x3.B.n41 1Bit_Clk_ADC_0.x3.B.n39 202.094
R33880 1Bit_Clk_ADC_0.x3.B.n0 1Bit_Clk_ADC_0.x3.B.n23 188.516
R33881 1Bit_Clk_ADC_0.x3.B.n3 1Bit_Clk_ADC_0.x3.B.n2 185
R33882 1Bit_Clk_ADC_0.x3.B.n4 1Bit_Clk_ADC_0.x3.B 182.786
R33883 1Bit_Clk_ADC_0.x3.B.n32 1Bit_Clk_ADC_0.x3.B.n31 180.482
R33884 1Bit_Clk_ADC_0.x3.B.n17 1Bit_Clk_ADC_0.x3.B 154.304
R33885 1Bit_Clk_ADC_0.x3.B.n13 1Bit_Clk_ADC_0.x3.B.n12 152
R33886 1Bit_Clk_ADC_0.x3.B.n10 1Bit_Clk_ADC_0.x3.B.n9 152
R33887 1Bit_Clk_ADC_0.x3.B.n8 1Bit_Clk_ADC_0.x3.B.n7 152
R33888 1Bit_Clk_ADC_0.x3.B.n34 1Bit_Clk_ADC_0.x3.B.n33 152
R33889 1Bit_Clk_ADC_0.x3.B.n29 1Bit_Clk_ADC_0.x3.B.n28 152
R33890 1Bit_Clk_ADC_0.x3.B.n27 1Bit_Clk_ADC_0.x3.B.n26 152
R33891 1Bit_Clk_ADC_0.x3.B.n22 1Bit_Clk_ADC_0.x3.B.n21 152
R33892 1Bit_Clk_ADC_0.x3.B.n20 1Bit_Clk_ADC_0.x3.B.n19 152
R33893 1Bit_Clk_ADC_0.x3.B.n4 1Bit_Clk_ADC_0.x3.B.t16 139.78
R33894 1Bit_Clk_ADC_0.x3.B.n11 1Bit_Clk_ADC_0.x3.B.t26 139.78
R33895 1Bit_Clk_ADC_0.x3.B.n5 1Bit_Clk_ADC_0.x3.B.t22 139.78
R33896 1Bit_Clk_ADC_0.x3.B.n6 1Bit_Clk_ADC_0.x3.B.t32 139.78
R33897 1Bit_Clk_ADC_0.x3.B.n25 1Bit_Clk_ADC_0.x3.B.t24 139.78
R33898 1Bit_Clk_ADC_0.x3.B.n24 1Bit_Clk_ADC_0.x3.B.t19 139.78
R33899 1Bit_Clk_ADC_0.x3.B.n30 1Bit_Clk_ADC_0.x3.B.t29 139.78
R33900 1Bit_Clk_ADC_0.x3.B.n32 1Bit_Clk_ADC_0.x3.B.t23 139.78
R33901 1Bit_Clk_ADC_0.x3.B.n16 1Bit_Clk_ADC_0.x3.B.t13 139.78
R33902 1Bit_Clk_ADC_0.x3.B.n18 1Bit_Clk_ADC_0.x3.B.t33 139.78
R33903 1Bit_Clk_ADC_0.x3.B.n15 1Bit_Clk_ADC_0.x3.B.t34 139.78
R33904 1Bit_Clk_ADC_0.x3.B.n23 1Bit_Clk_ADC_0.x3.B.t27 139.78
R33905 1Bit_Clk_ADC_0.x3.B.n12 1Bit_Clk_ADC_0.x3.B.n4 30.6732
R33906 1Bit_Clk_ADC_0.x3.B.n12 1Bit_Clk_ADC_0.x3.B.n11 30.6732
R33907 1Bit_Clk_ADC_0.x3.B.n11 1Bit_Clk_ADC_0.x3.B.n10 30.6732
R33908 1Bit_Clk_ADC_0.x3.B.n10 1Bit_Clk_ADC_0.x3.B.n5 30.6732
R33909 1Bit_Clk_ADC_0.x3.B.n7 1Bit_Clk_ADC_0.x3.B.n5 30.6732
R33910 1Bit_Clk_ADC_0.x3.B.n7 1Bit_Clk_ADC_0.x3.B.n6 30.6732
R33911 1Bit_Clk_ADC_0.x3.B.n26 1Bit_Clk_ADC_0.x3.B.n25 30.6732
R33912 1Bit_Clk_ADC_0.x3.B.n26 1Bit_Clk_ADC_0.x3.B.n24 30.6732
R33913 1Bit_Clk_ADC_0.x3.B.n29 1Bit_Clk_ADC_0.x3.B.n24 30.6732
R33914 1Bit_Clk_ADC_0.x3.B.n30 1Bit_Clk_ADC_0.x3.B.n29 30.6732
R33915 1Bit_Clk_ADC_0.x3.B.n33 1Bit_Clk_ADC_0.x3.B.n30 30.6732
R33916 1Bit_Clk_ADC_0.x3.B.n33 1Bit_Clk_ADC_0.x3.B.n32 30.6732
R33917 1Bit_Clk_ADC_0.x3.B.n17 1Bit_Clk_ADC_0.x3.B.n16 30.6732
R33918 1Bit_Clk_ADC_0.x3.B.n18 1Bit_Clk_ADC_0.x3.B.n17 30.6732
R33919 1Bit_Clk_ADC_0.x3.B.n19 1Bit_Clk_ADC_0.x3.B.n18 30.6732
R33920 1Bit_Clk_ADC_0.x3.B.n19 1Bit_Clk_ADC_0.x3.B.n15 30.6732
R33921 1Bit_Clk_ADC_0.x3.B.n22 1Bit_Clk_ADC_0.x3.B.n15 30.6732
R33922 1Bit_Clk_ADC_0.x3.B.n23 1Bit_Clk_ADC_0.x3.B.n22 30.6732
R33923 1Bit_Clk_ADC_0.x3.B.n39 1Bit_Clk_ADC_0.x3.B.t8 26.5955
R33924 1Bit_Clk_ADC_0.x3.B.n39 1Bit_Clk_ADC_0.x3.B.t9 26.5955
R33925 1Bit_Clk_ADC_0.x3.B.n40 1Bit_Clk_ADC_0.x3.B.t10 26.5955
R33926 1Bit_Clk_ADC_0.x3.B.n40 1Bit_Clk_ADC_0.x3.B.t11 26.5955
R33927 1Bit_Clk_ADC_0.x3.B.n43 1Bit_Clk_ADC_0.x3.B.t2 26.5955
R33928 1Bit_Clk_ADC_0.x3.B.n43 1Bit_Clk_ADC_0.x3.B.t0 26.5955
R33929 1Bit_Clk_ADC_0.x3.B.n44 1Bit_Clk_ADC_0.x3.B.t1 26.5955
R33930 1Bit_Clk_ADC_0.x3.B.n44 1Bit_Clk_ADC_0.x3.B.t3 26.5955
R33931 1Bit_Clk_ADC_0.x3.B.n2 1Bit_Clk_ADC_0.x3.B.t4 24.9236
R33932 1Bit_Clk_ADC_0.x3.B.n2 1Bit_Clk_ADC_0.x3.B.t5 24.9236
R33933 1Bit_Clk_ADC_0.x3.B.n1 1Bit_Clk_ADC_0.x3.B.t6 24.9236
R33934 1Bit_Clk_ADC_0.x3.B.n1 1Bit_Clk_ADC_0.x3.B.t7 24.9236
R33935 1Bit_Clk_ADC_0.x3.B 1Bit_Clk_ADC_0.x3.B.n45 22.9652
R33936 1Bit_Clk_ADC_0.x3.B.n28 1Bit_Clk_ADC_0.x3.B.n27 21.5045
R33937 1Bit_Clk_ADC_0.x3.B.n38 1Bit_Clk_ADC_0.x3.B.n3 21.4064
R33938 1Bit_Clk_ADC_0.x3.B.n37 1Bit_Clk_ADC_0.x3.B.n14 20.3538
R33939 1Bit_Clk_ADC_0.x3.B.n20 1Bit_Clk_ADC_0.x3.B 19.2005
R33940 1Bit_Clk_ADC_0.x3.B.n35 1Bit_Clk_ADC_0.x3.B 17.6645
R33941 1Bit_Clk_ADC_0.x3.B.n31 1Bit_Clk_ADC_0.x3.B 17.1525
R33942 1Bit_Clk_ADC_0.x3.B.n21 1Bit_Clk_ADC_0.x3.B 17.1525
R33943 1Bit_Clk_ADC_0.x3.B.n0 1Bit_Clk_ADC_0.x3.B 16.8965
R33944 1Bit_Clk_ADC_0.x3.B.n9 1Bit_Clk_ADC_0.x3.B 16.3845
R33945 1Bit_Clk_ADC_0.x3.B.n14 1Bit_Clk_ADC_0.x3.B 15.3605
R33946 1Bit_Clk_ADC_0.x3.B 1Bit_Clk_ADC_0.x3.B.n8 14.3365
R33947 1Bit_Clk_ADC_0.x3.B.n42 1Bit_Clk_ADC_0.x3.B.n41 13.9299
R33948 1Bit_Clk_ADC_0.x3.B 1Bit_Clk_ADC_0.x3.B.n42 13.9299
R33949 1Bit_Clk_ADC_0.x3.B.n36 1Bit_Clk_ADC_0.x3.B.n35 10.863
R33950 1Bit_Clk_ADC_0.x3.B.n36 1Bit_Clk_ADC_0.x3.B.n0 9.488
R33951 1Bit_Clk_ADC_0.x3.B.n38 1Bit_Clk_ADC_0.x3.B.n37 9.3005
R33952 1Bit_Clk_ADC_0.x3.B.n8 1Bit_Clk_ADC_0.x3.B 9.2165
R33953 1Bit_Clk_ADC_0.x3.B.n9 1Bit_Clk_ADC_0.x3.B 7.1685
R33954 1Bit_Clk_ADC_0.x3.B.n0 1Bit_Clk_ADC_0.x3.B 6.6565
R33955 1Bit_Clk_ADC_0.x3.B.n31 1Bit_Clk_ADC_0.x3.B 6.4005
R33956 1Bit_Clk_ADC_0.x3.B.n21 1Bit_Clk_ADC_0.x3.B 6.4005
R33957 1Bit_Clk_ADC_0.x3.B.n42 1Bit_Clk_ADC_0.x3.B 5.26405
R33958 1Bit_Clk_ADC_0.x3.B.n13 1Bit_Clk_ADC_0.x3.B 5.1205
R33959 1Bit_Clk_ADC_0.x3.B 1Bit_Clk_ADC_0.x3.B.n20 4.3525
R33960 1Bit_Clk_ADC_0.x3.B.n34 1Bit_Clk_ADC_0.x3.B 3.5845
R33961 1Bit_Clk_ADC_0.x3.B.n14 1Bit_Clk_ADC_0.x3.B.n13 3.0725
R33962 1Bit_Clk_ADC_0.x3.B.n42 1Bit_Clk_ADC_0.x3.B 2.87153
R33963 1Bit_Clk_ADC_0.x3.B.n35 1Bit_Clk_ADC_0.x3.B.n34 2.3045
R33964 1Bit_Clk_ADC_0.x3.B 1Bit_Clk_ADC_0.x3.B.n38 1.55564
R33965 1Bit_Clk_ADC_0.x3.B.n28 1Bit_Clk_ADC_0.x3.B 1.5365
R33966 1Bit_Clk_ADC_0.x3.B.n37 1Bit_Clk_ADC_0.x3.B.n36 1.29878
R33967 1Bit_Clk_ADC_0.x3.B.n27 1Bit_Clk_ADC_0.x3.B 0.5125
R33968 OUT.n68 OUT.t30 1038.79
R33969 OUT.n82 OUT.t16 1038.79
R33970 OUT.n59 OUT.t50 1038.78
R33971 OUT.n60 OUT.t35 1038.78
R33972 OUT.n68 OUT.t39 1038.55
R33973 OUT.n69 OUT.t41 1038.55
R33974 OUT.n70 OUT.t72 1038.55
R33975 OUT.n71 OUT.t28 1038.55
R33976 OUT.n72 OUT.t63 1038.55
R33977 OUT.n73 OUT.t70 1038.55
R33978 OUT.n74 OUT.t71 1038.55
R33979 OUT.n75 OUT.t27 1038.55
R33980 OUT.n76 OUT.t61 1038.55
R33981 OUT.n82 OUT.t87 1038.55
R33982 OUT.n35 OUT.t29 1038.55
R33983 OUT.n36 OUT.t38 1038.55
R33984 OUT.n37 OUT.t15 1038.55
R33985 OUT.n38 OUT.t21 1038.55
R33986 OUT.n39 OUT.t22 1038.55
R33987 OUT.n40 OUT.t54 1038.55
R33988 OUT.n41 OUT.t81 1038.55
R33989 OUT.n42 OUT.t42 1038.55
R33990 OUT.n43 OUT.t49 1038.55
R33991 OUT.n44 OUT.t78 1038.55
R33992 OUT.n45 OUT.t80 1038.55
R33993 OUT.n46 OUT.t40 1038.55
R33994 OUT.n59 OUT.t14 1038.54
R33995 OUT.n67 OUT.t32 1038.54
R33996 OUT.n66 OUT.t24 1038.54
R33997 OUT.n65 OUT.t68 1038.54
R33998 OUT.n64 OUT.t65 1038.54
R33999 OUT.n63 OUT.t33 1038.54
R34000 OUT.n62 OUT.t74 1038.54
R34001 OUT.n61 OUT.t69 1038.54
R34002 OUT.n60 OUT.t36 1038.54
R34003 OUT.n47 OUT.t85 1038.54
R34004 OUT.n48 OUT.t76 1038.54
R34005 OUT.n49 OUT.t75 1038.54
R34006 OUT.n50 OUT.t45 1038.54
R34007 OUT.n51 OUT.t86 1038.54
R34008 OUT.n52 OUT.t58 1038.54
R34009 OUT.n53 OUT.t53 1038.54
R34010 OUT.n54 OUT.t52 1038.54
R34011 OUT.n55 OUT.t17 1038.54
R34012 OUT.n56 OUT.t67 1038.54
R34013 OUT.n57 OUT.t34 1038.54
R34014 OUT OUT.t82 1029.08
R34015 OUT OUT.t25 1029.08
R34016 OUT.n33 OUT.t31 1028.97
R34017 OUT.n24 OUT.t59 1024.54
R34018 OUT.n85 OUT.t79 1024.51
R34019 OUT.n27 OUT.t56 1024.51
R34020 OUT.n89 OUT.t51 1024.08
R34021 OUT.n90 OUT.t44 1024.08
R34022 OUT.n91 OUT.t43 1024.08
R34023 OUT.n92 OUT.t84 1024.08
R34024 OUT.n93 OUT.t12 1024.08
R34025 OUT.n88 OUT.t77 1024.08
R34026 OUT.n87 OUT.t48 1024.08
R34027 OUT.n86 OUT.t47 1024.08
R34028 OUT.n85 OUT.t13 1024.08
R34029 OUT.n26 OUT.t26 1024.08
R34030 OUT.n25 OUT.t19 1024.08
R34031 OUT.n24 OUT.t62 1024.08
R34032 OUT.n30 OUT.t55 1024.08
R34033 OUT.n29 OUT.t23 1024.08
R34034 OUT.n28 OUT.t66 1024.08
R34035 OUT.n27 OUT.t64 1024.08
R34036 OUT.n2 OUT.n1 256.103
R34037 OUT.n5 OUT.n3 243.68
R34038 OUT.n9 OUT.n7 241.847
R34039 OUT.n11 OUT.t60 212.081
R34040 OUT.n14 OUT.t20 212.081
R34041 OUT.n16 OUT.t83 212.081
R34042 OUT.n15 OUT.t46 212.081
R34043 OUT.n5 OUT.n4 205.28
R34044 OUT.n2 OUT.n0 202.095
R34045 OUT.n9 OUT.n8 185
R34046 OUT.n18 OUT.n17 154.816
R34047 OUT.n13 OUT.n12 152
R34048 OUT.n11 OUT.t37 139.78
R34049 OUT.n14 OUT.t73 139.78
R34050 OUT.n16 OUT.t57 139.78
R34051 OUT.n15 OUT.t18 139.78
R34052 OUT.n16 OUT.n15 61.346
R34053 OUT.n13 OUT.n11 30.6732
R34054 OUT.n14 OUT.n13 30.6732
R34055 OUT.n17 OUT.n14 30.6732
R34056 OUT.n17 OUT.n16 30.6732
R34057 OUT.n0 OUT.t11 26.5955
R34058 OUT.n0 OUT.t9 26.5955
R34059 OUT.n3 OUT.t2 26.5955
R34060 OUT.n3 OUT.t3 26.5955
R34061 OUT.n4 OUT.t0 26.5955
R34062 OUT.n4 OUT.t1 26.5955
R34063 OUT.n1 OUT.t8 26.5955
R34064 OUT.n1 OUT.t10 26.5955
R34065 OUT.n8 OUT.t4 24.9236
R34066 OUT.n8 OUT.t6 24.9236
R34067 OUT.n7 OUT.t5 24.9236
R34068 OUT.n7 OUT.t7 24.9236
R34069 OUT OUT.n5 22.9652
R34070 OUT OUT.n9 18.8943
R34071 OUT.n19 OUT.n10 15.4113
R34072 OUT.n19 OUT.n18 14.9099
R34073 OUT.n12 OUT 14.8485
R34074 OUT.n6 OUT.n2 13.9299
R34075 OUT.n6 OUT 13.9299
R34076 OUT.n89 OUT.n88 11.077
R34077 OUT.n47 OUT.n46 11.038
R34078 OUT.n78 OUT.n77 9.27134
R34079 OUT.n32 OUT.n31 8.81565
R34080 OUT.n12 OUT 8.7045
R34081 OUT.n31 OUT.n26 5.79686
R34082 OUT.n77 OUT.n67 5.65425
R34083 OUT.n78 OUT.n59 5.63925
R34084 OUT.n10 OUT 5.62293
R34085 OUT.n31 OUT.n30 5.56709
R34086 OUT.n77 OUT.n76 5.40925
R34087 OUT.n94 OUT.n93 4.88925
R34088 OUT.n58 OUT.n57 4.82675
R34089 OUT.n83 OUT.n82 4.70675
R34090 OUT.n35 OUT.n34 4.70675
R34091 OUT OUT.n98 4.09615
R34092 OUT.n18 OUT 3.8405
R34093 OUT.n20 OUT.n19 3.4105
R34094 OUT.n98 OUT.n58 2.94106
R34095 OUT.n10 OUT 2.51265
R34096 OUT.n93 OUT.n92 2.3755
R34097 OUT.n98 OUT.n97 2.0245
R34098 OUT.n79 OUT 1.9755
R34099 OUT.n84 OUT 1.4755
R34100 OUT.n95 OUT 1.2005
R34101 OUT OUT.n6 1.19676
R34102 OUT.n34 OUT.n23 1.0255
R34103 OUT.n56 OUT.n55 1.0105
R34104 OUT.n37 OUT.n36 1.0105
R34105 OUT.n97 OUT.n80 0.853
R34106 OUT.n97 OUT.n96 0.853
R34107 OUT.n81 OUT 0.8505
R34108 OUT.n33 OUT.n32 0.7505
R34109 OUT.n23 OUT 0.678625
R34110 OUT.n32 OUT 0.6255
R34111 OUT.n95 OUT 0.6005
R34112 OUT.n25 OUT.n24 0.4605
R34113 OUT.n26 OUT.n25 0.4605
R34114 OUT.n86 OUT.n85 0.428449
R34115 OUT.n87 OUT.n86 0.428449
R34116 OUT.n88 OUT.n87 0.428449
R34117 OUT.n28 OUT.n27 0.428449
R34118 OUT.n29 OUT.n28 0.428449
R34119 OUT.n30 OUT.n29 0.428449
R34120 OUT.n79 OUT.n78 0.4005
R34121 OUT.n34 OUT.n33 0.313
R34122 OUT.n61 OUT.n60 0.2405
R34123 OUT.n62 OUT.n61 0.2405
R34124 OUT.n63 OUT.n62 0.2405
R34125 OUT.n64 OUT.n63 0.2405
R34126 OUT.n65 OUT.n64 0.2405
R34127 OUT.n66 OUT.n65 0.2405
R34128 OUT.n67 OUT.n66 0.2405
R34129 OUT.n69 OUT.n68 0.2405
R34130 OUT.n70 OUT.n69 0.2405
R34131 OUT.n71 OUT.n70 0.2405
R34132 OUT.n72 OUT.n71 0.2405
R34133 OUT.n73 OUT.n72 0.2405
R34134 OUT.n74 OUT.n73 0.2405
R34135 OUT.n75 OUT.n74 0.2405
R34136 OUT.n76 OUT.n75 0.2405
R34137 OUT.n92 OUT.n91 0.2405
R34138 OUT.n91 OUT.n90 0.2405
R34139 OUT.n90 OUT.n89 0.2405
R34140 OUT.n57 OUT.n56 0.2405
R34141 OUT.n55 OUT.n54 0.2405
R34142 OUT.n54 OUT.n53 0.2405
R34143 OUT.n53 OUT.n52 0.2405
R34144 OUT.n52 OUT.n51 0.2405
R34145 OUT.n51 OUT.n50 0.2405
R34146 OUT.n50 OUT.n49 0.2405
R34147 OUT.n49 OUT.n48 0.2405
R34148 OUT.n48 OUT.n47 0.2405
R34149 OUT.n36 OUT.n35 0.2405
R34150 OUT.n38 OUT.n37 0.2405
R34151 OUT.n39 OUT.n38 0.2405
R34152 OUT.n40 OUT.n39 0.2405
R34153 OUT.n41 OUT.n40 0.2405
R34154 OUT.n42 OUT.n41 0.2405
R34155 OUT.n43 OUT.n42 0.2405
R34156 OUT.n44 OUT.n43 0.2405
R34157 OUT.n45 OUT.n44 0.2405
R34158 OUT.n46 OUT.n45 0.2405
R34159 OUT.n84 OUT.n83 0.213
R34160 OUT.n58 OUT.n23 0.11925
R34161 OUT OUT.n22 0.109775
R34162 OUT.n96 OUT.n95 0.06925
R34163 OUT.n80 OUT.n79 0.06925
R34164 OUT.n81 OUT.n80 0.06925
R34165 OUT.n94 OUT.n84 0.0505
R34166 OUT.n22 OUT 0.04891
R34167 OUT.n21 OUT.n20 0.024
R34168 OUT.n20 OUT 0.024
R34169 OUT.n96 OUT.n94 0.01925
R34170 OUT.n83 OUT.n81 0.013
R34171 OUT.n21 OUT 0.00833333
R34172 OUT.n22 OUT.n21 0.000891667
R34173 a_216435_n47946.n19 a_216435_n47946.t13 1038.55
R34174 a_216435_n47946.n18 a_216435_n47946.t16 1038.55
R34175 a_216435_n47946.n17 a_216435_n47946.t17 1038.55
R34176 a_216435_n47946.n16 a_216435_n47946.t26 1038.55
R34177 a_216435_n47946.n15 a_216435_n47946.t10 1038.55
R34178 a_216435_n47946.n14 a_216435_n47946.t21 1038.55
R34179 a_216435_n47946.n13 a_216435_n47946.t23 1038.55
R34180 a_216435_n47946.n12 a_216435_n47946.t8 1038.55
R34181 a_216435_n47946.n11 a_216435_n47946.t9 1038.55
R34182 a_216435_n47946.n10 a_216435_n47946.t20 1038.55
R34183 a_216435_n47946.n9 a_216435_n47946.t11 1038.54
R34184 a_216435_n47946.n8 a_216435_n47946.t7 1038.54
R34185 a_216435_n47946.n7 a_216435_n47946.t6 1038.54
R34186 a_216435_n47946.n6 a_216435_n47946.t22 1038.54
R34187 a_216435_n47946.n5 a_216435_n47946.t12 1038.54
R34188 a_216435_n47946.n4 a_216435_n47946.t29 1038.54
R34189 a_216435_n47946.n3 a_216435_n47946.t25 1038.54
R34190 a_216435_n47946.n2 a_216435_n47946.t24 1038.54
R34191 a_216435_n47946.n1 a_216435_n47946.t14 1038.54
R34192 a_216435_n47946.n21 a_216435_n47946.t30 1024.54
R34193 a_216435_n47946.n24 a_216435_n47946.t28 1024.51
R34194 a_216435_n47946.n23 a_216435_n47946.t19 1024.08
R34195 a_216435_n47946.n22 a_216435_n47946.t15 1024.08
R34196 a_216435_n47946.n21 a_216435_n47946.t31 1024.08
R34197 a_216435_n47946.n27 a_216435_n47946.t27 1024.08
R34198 a_216435_n47946.n26 a_216435_n47946.t18 1024.08
R34199 a_216435_n47946.n25 a_216435_n47946.t33 1024.08
R34200 a_216435_n47946.n24 a_216435_n47946.t32 1024.08
R34201 a_216435_n47946.n31 a_216435_n47946.n30 52.1388
R34202 a_216435_n47946.n33 a_216435_n47946.n32 48.672
R34203 a_216435_n47946.n32 a_216435_n47946.n0 19.8859
R34204 a_216435_n47946.n10 a_216435_n47946.n9 11.038
R34205 a_216435_n47946.n29 a_216435_n47946.n28 9.2841
R34206 a_216435_n47946.n30 a_216435_n47946.t4 6.5015
R34207 a_216435_n47946.n30 a_216435_n47946.t3 6.5015
R34208 a_216435_n47946.n33 a_216435_n47946.t2 6.5015
R34209 a_216435_n47946.t5 a_216435_n47946.n33 6.5015
R34210 a_216435_n47946.n20 a_216435_n47946.n1 6.48538
R34211 a_216435_n47946.n28 a_216435_n47946.n23 5.79686
R34212 a_216435_n47946.n28 a_216435_n47946.n27 5.56709
R34213 a_216435_n47946.n20 a_216435_n47946.n19 4.86925
R34214 a_216435_n47946.n0 a_216435_n47946.t0 3.9605
R34215 a_216435_n47946.n0 a_216435_n47946.t1 3.9605
R34216 a_216435_n47946.n31 a_216435_n47946.n29 3.62905
R34217 a_216435_n47946.n32 a_216435_n47946.n31 3.48527
R34218 a_216435_n47946.n22 a_216435_n47946.n21 0.4605
R34219 a_216435_n47946.n23 a_216435_n47946.n22 0.4605
R34220 a_216435_n47946.n25 a_216435_n47946.n24 0.428449
R34221 a_216435_n47946.n26 a_216435_n47946.n25 0.428449
R34222 a_216435_n47946.n27 a_216435_n47946.n26 0.428449
R34223 a_216435_n47946.n19 a_216435_n47946.n18 0.2405
R34224 a_216435_n47946.n18 a_216435_n47946.n17 0.2405
R34225 a_216435_n47946.n17 a_216435_n47946.n16 0.2405
R34226 a_216435_n47946.n16 a_216435_n47946.n15 0.2405
R34227 a_216435_n47946.n15 a_216435_n47946.n14 0.2405
R34228 a_216435_n47946.n14 a_216435_n47946.n13 0.2405
R34229 a_216435_n47946.n13 a_216435_n47946.n12 0.2405
R34230 a_216435_n47946.n12 a_216435_n47946.n11 0.2405
R34231 a_216435_n47946.n11 a_216435_n47946.n10 0.2405
R34232 a_216435_n47946.n2 a_216435_n47946.n1 0.2405
R34233 a_216435_n47946.n3 a_216435_n47946.n2 0.2405
R34234 a_216435_n47946.n4 a_216435_n47946.n3 0.2405
R34235 a_216435_n47946.n5 a_216435_n47946.n4 0.2405
R34236 a_216435_n47946.n6 a_216435_n47946.n5 0.2405
R34237 a_216435_n47946.n7 a_216435_n47946.n6 0.2405
R34238 a_216435_n47946.n8 a_216435_n47946.n7 0.2405
R34239 a_216435_n47946.n9 a_216435_n47946.n8 0.2405
R34240 a_216435_n47946.n29 a_216435_n47946.n20 0.188
R34241 a_155026_n27776.n6 a_155026_n27776.n5 22.4024
R34242 a_155026_n27776.n7 a_155026_n27776.n2 18.9924
R34243 a_155026_n27776.n4 a_155026_n27776.n3 18.9924
R34244 a_155026_n27776.n7 a_155026_n27776.n6 3.716
R34245 a_155026_n27776.n6 a_155026_n27776.n4 3.71013
R34246 a_155026_n27776.n3 a_155026_n27776.t5 3.4805
R34247 a_155026_n27776.n3 a_155026_n27776.t4 3.4805
R34248 a_155026_n27776.n2 a_155026_n27776.t8 3.4805
R34249 a_155026_n27776.n2 a_155026_n27776.t7 3.4805
R34250 a_155026_n27776.n5 a_155026_n27776.t6 3.4805
R34251 a_155026_n27776.n5 a_155026_n27776.t1 3.4805
R34252 a_155026_n27776.n9 a_155026_n27776.t2 3.04088
R34253 a_155026_n27776.n0 a_155026_n27776.t9 3.03453
R34254 a_155026_n27776.t0 a_155026_n27776.n9 2.59519
R34255 a_155026_n27776.n0 a_155026_n27776.t3 2.59419
R34256 a_155026_n27776.n8 a_155026_n27776.n7 2.55108
R34257 a_155026_n27776.n4 a_155026_n27776.n1 2.55108
R34258 a_155026_n27776.n8 a_155026_n27776.n1 0.293114
R34259 a_155026_n27776.n9 a_155026_n27776.n8 0.078625
R34260 a_155026_n27776.n1 a_155026_n27776.n0 0.0672614
R34261 1Bit_DAC_0.OUT.n1 1Bit_DAC_0.OUT.t36 57.0195
R34262 1Bit_DAC_0.OUT.n54 1Bit_DAC_0.OUT.t11 56.9568
R34263 1Bit_DAC_0.OUT.n30 1Bit_DAC_0.OUT.n27 50.515
R34264 1Bit_DAC_0.OUT.n32 1Bit_DAC_0.OUT.n31 50.4558
R34265 1Bit_DAC_0.OUT.n34 1Bit_DAC_0.OUT.n33 50.4558
R34266 1Bit_DAC_0.OUT.n51 1Bit_DAC_0.OUT.n50 50.4558
R34267 1Bit_DAC_0.OUT.n11 1Bit_DAC_0.OUT.n10 50.4558
R34268 1Bit_DAC_0.OUT.n9 1Bit_DAC_0.OUT.n8 50.4558
R34269 1Bit_DAC_0.OUT.n36 1Bit_DAC_0.OUT.n35 50.438
R34270 1Bit_DAC_0.OUT.n47 1Bit_DAC_0.OUT.n46 50.438
R34271 1Bit_DAC_0.OUT.n17 1Bit_DAC_0.OUT.n16 50.438
R34272 1Bit_DAC_0.OUT.n13 1Bit_DAC_0.OUT.n12 50.438
R34273 1Bit_DAC_0.OUT.n7 1Bit_DAC_0.OUT.n6 50.438
R34274 1Bit_DAC_0.OUT.n5 1Bit_DAC_0.OUT.n4 50.438
R34275 1Bit_DAC_0.OUT.n1 1Bit_DAC_0.OUT.n0 50.438
R34276 1Bit_DAC_0.OUT.n29 1Bit_DAC_0.OUT.n28 50.4246
R34277 1Bit_DAC_0.OUT.n39 1Bit_DAC_0.OUT.n38 50.4246
R34278 1Bit_DAC_0.OUT.n43 1Bit_DAC_0.OUT.n42 50.4246
R34279 1Bit_DAC_0.OUT.n15 1Bit_DAC_0.OUT.n14 50.4246
R34280 1Bit_DAC_0.OUT.n3 1Bit_DAC_0.OUT.n2 50.4246
R34281 1Bit_DAC_0.OUT.n37 1Bit_DAC_0.OUT.t42 25.1211
R34282 1Bit_DAC_0.OUT.n25 1Bit_DAC_0.OUT.t6 25.1211
R34283 1Bit_DAC_0.OUT.n20 1Bit_DAC_0.OUT.n18 21.23
R34284 1Bit_DAC_0.OUT.n41 1Bit_DAC_0.OUT.n40 21.179
R34285 1Bit_DAC_0.OUT.n49 1Bit_DAC_0.OUT.n48 21.179
R34286 1Bit_DAC_0.OUT.n53 1Bit_DAC_0.OUT.n52 21.179
R34287 1Bit_DAC_0.OUT.n24 1Bit_DAC_0.OUT.n23 21.179
R34288 1Bit_DAC_0.OUT.n20 1Bit_DAC_0.OUT.n19 21.179
R34289 1Bit_DAC_0.OUT.n45 1Bit_DAC_0.OUT.n44 21.1611
R34290 1Bit_DAC_0.OUT.n22 1Bit_DAC_0.OUT.n21 21.1611
R34291 1Bit_DAC_0.OUT.n28 1Bit_DAC_0.OUT.t12 6.5015
R34292 1Bit_DAC_0.OUT.n28 1Bit_DAC_0.OUT.t8 6.5015
R34293 1Bit_DAC_0.OUT.n27 1Bit_DAC_0.OUT.t2 6.5015
R34294 1Bit_DAC_0.OUT.n27 1Bit_DAC_0.OUT.t0 6.5015
R34295 1Bit_DAC_0.OUT.n35 1Bit_DAC_0.OUT.t22 6.5015
R34296 1Bit_DAC_0.OUT.n35 1Bit_DAC_0.OUT.t16 6.5015
R34297 1Bit_DAC_0.OUT.n38 1Bit_DAC_0.OUT.t18 6.5015
R34298 1Bit_DAC_0.OUT.n38 1Bit_DAC_0.OUT.t10 6.5015
R34299 1Bit_DAC_0.OUT.n42 1Bit_DAC_0.OUT.t21 6.5015
R34300 1Bit_DAC_0.OUT.n42 1Bit_DAC_0.OUT.t15 6.5015
R34301 1Bit_DAC_0.OUT.n31 1Bit_DAC_0.OUT.t13 6.5015
R34302 1Bit_DAC_0.OUT.n31 1Bit_DAC_0.OUT.t19 6.5015
R34303 1Bit_DAC_0.OUT.n33 1Bit_DAC_0.OUT.t20 6.5015
R34304 1Bit_DAC_0.OUT.n33 1Bit_DAC_0.OUT.t27 6.5015
R34305 1Bit_DAC_0.OUT.n46 1Bit_DAC_0.OUT.t1 6.5015
R34306 1Bit_DAC_0.OUT.n46 1Bit_DAC_0.OUT.t24 6.5015
R34307 1Bit_DAC_0.OUT.n50 1Bit_DAC_0.OUT.t9 6.5015
R34308 1Bit_DAC_0.OUT.n50 1Bit_DAC_0.OUT.t14 6.5015
R34309 1Bit_DAC_0.OUT.n16 1Bit_DAC_0.OUT.t33 6.5015
R34310 1Bit_DAC_0.OUT.n16 1Bit_DAC_0.OUT.t43 6.5015
R34311 1Bit_DAC_0.OUT.n14 1Bit_DAC_0.OUT.t39 6.5015
R34312 1Bit_DAC_0.OUT.n14 1Bit_DAC_0.OUT.t31 6.5015
R34313 1Bit_DAC_0.OUT.n12 1Bit_DAC_0.OUT.t52 6.5015
R34314 1Bit_DAC_0.OUT.n12 1Bit_DAC_0.OUT.t30 6.5015
R34315 1Bit_DAC_0.OUT.n6 1Bit_DAC_0.OUT.t48 6.5015
R34316 1Bit_DAC_0.OUT.n6 1Bit_DAC_0.OUT.t45 6.5015
R34317 1Bit_DAC_0.OUT.n4 1Bit_DAC_0.OUT.t38 6.5015
R34318 1Bit_DAC_0.OUT.n4 1Bit_DAC_0.OUT.t50 6.5015
R34319 1Bit_DAC_0.OUT.n10 1Bit_DAC_0.OUT.t53 6.5015
R34320 1Bit_DAC_0.OUT.n10 1Bit_DAC_0.OUT.t51 6.5015
R34321 1Bit_DAC_0.OUT.n8 1Bit_DAC_0.OUT.t44 6.5015
R34322 1Bit_DAC_0.OUT.n8 1Bit_DAC_0.OUT.t41 6.5015
R34323 1Bit_DAC_0.OUT.n2 1Bit_DAC_0.OUT.t56 6.5015
R34324 1Bit_DAC_0.OUT.n2 1Bit_DAC_0.OUT.t40 6.5015
R34325 1Bit_DAC_0.OUT.n0 1Bit_DAC_0.OUT.t32 6.5015
R34326 1Bit_DAC_0.OUT.n0 1Bit_DAC_0.OUT.t37 6.5015
R34327 1Bit_DAC_0.OUT.n29 1Bit_DAC_0.OUT.t28 4.07308
R34328 1Bit_DAC_0.OUT.n40 1Bit_DAC_0.OUT.t34 3.9605
R34329 1Bit_DAC_0.OUT.n40 1Bit_DAC_0.OUT.t35 3.9605
R34330 1Bit_DAC_0.OUT.n44 1Bit_DAC_0.OUT.t47 3.9605
R34331 1Bit_DAC_0.OUT.n44 1Bit_DAC_0.OUT.t54 3.9605
R34332 1Bit_DAC_0.OUT.n48 1Bit_DAC_0.OUT.t55 3.9605
R34333 1Bit_DAC_0.OUT.n48 1Bit_DAC_0.OUT.t46 3.9605
R34334 1Bit_DAC_0.OUT.n52 1Bit_DAC_0.OUT.t29 3.9605
R34335 1Bit_DAC_0.OUT.n52 1Bit_DAC_0.OUT.t49 3.9605
R34336 1Bit_DAC_0.OUT.n23 1Bit_DAC_0.OUT.t3 3.9605
R34337 1Bit_DAC_0.OUT.n23 1Bit_DAC_0.OUT.t25 3.9605
R34338 1Bit_DAC_0.OUT.n21 1Bit_DAC_0.OUT.t23 3.9605
R34339 1Bit_DAC_0.OUT.n21 1Bit_DAC_0.OUT.t4 3.9605
R34340 1Bit_DAC_0.OUT.n19 1Bit_DAC_0.OUT.t5 3.9605
R34341 1Bit_DAC_0.OUT.n19 1Bit_DAC_0.OUT.t17 3.9605
R34342 1Bit_DAC_0.OUT.n18 1Bit_DAC_0.OUT.t26 3.9605
R34343 1Bit_DAC_0.OUT.n18 1Bit_DAC_0.OUT.t7 3.9605
R34344 1Bit_DAC_0.OUT.n26 1Bit_DAC_0.OUT.n17 0.0663
R34345 1Bit_DAC_0.OUT.n3 1Bit_DAC_0.OUT.n1 0.0631667
R34346 1Bit_DAC_0.OUT.n7 1Bit_DAC_0.OUT.n5 0.0631667
R34347 1Bit_DAC_0.OUT.n9 1Bit_DAC_0.OUT.n7 0.0631667
R34348 1Bit_DAC_0.OUT.n11 1Bit_DAC_0.OUT.n9 0.0631667
R34349 1Bit_DAC_0.OUT.n13 1Bit_DAC_0.OUT.n11 0.0631667
R34350 1Bit_DAC_0.OUT.n15 1Bit_DAC_0.OUT.n13 0.0631667
R34351 1Bit_DAC_0.OUT.n24 1Bit_DAC_0.OUT.n22 0.0631667
R34352 1Bit_DAC_0.OUT.n22 1Bit_DAC_0.OUT.n20 0.0569
R34353 1Bit_DAC_0.OUT.n25 1Bit_DAC_0.OUT.n24 0.0569
R34354 1Bit_DAC_0.OUT.n5 1Bit_DAC_0.OUT.n3 0.0506333
R34355 1Bit_DAC_0.OUT.n17 1Bit_DAC_0.OUT.n15 0.0443667
R34356 1Bit_DAC_0.OUT.n26 1Bit_DAC_0.OUT.n25 0.0349667
R34357 1Bit_DAC_0.OUT.n36 1Bit_DAC_0.OUT.n34 0.024
R34358 1Bit_DAC_0.OUT.n34 1Bit_DAC_0.OUT.n32 0.024
R34359 1Bit_DAC_0.OUT.n32 1Bit_DAC_0.OUT.n30 0.0205533
R34360 1Bit_DAC_0.OUT 1Bit_DAC_0.OUT.n26 0.0146
R34361 1Bit_DAC_0.OUT.n43 1Bit_DAC_0.OUT.n41 0.0146
R34362 1Bit_DAC_0.OUT.n39 1Bit_DAC_0.OUT.n37 0.0146
R34363 1Bit_DAC_0.OUT 1Bit_DAC_0.OUT.n54 0.013425
R34364 1Bit_DAC_0.OUT.n54 1Bit_DAC_0.OUT.n53 0.01225
R34365 1Bit_DAC_0.OUT.n53 1Bit_DAC_0.OUT.n51 0.01225
R34366 1Bit_DAC_0.OUT.n51 1Bit_DAC_0.OUT.n49 0.01225
R34367 1Bit_DAC_0.OUT.n49 1Bit_DAC_0.OUT.n47 0.01225
R34368 1Bit_DAC_0.OUT.n47 1Bit_DAC_0.OUT.n45 0.01225
R34369 1Bit_DAC_0.OUT.n41 1Bit_DAC_0.OUT.n39 0.0099
R34370 1Bit_DAC_0.OUT.n37 1Bit_DAC_0.OUT.n36 0.0099
R34371 1Bit_DAC_0.OUT.n30 1Bit_DAC_0.OUT.n29 0.008725
R34372 1Bit_DAC_0.OUT.n45 1Bit_DAC_0.OUT.n43 0.00755
R34373 VREFP.n1 VREFP.t44 57.5333
R34374 VREFP.n36 VREFP.t10 57.4858
R34375 VREFP.n49 VREFP.n36 51.9355
R34376 VREFP.n3 VREFP.n2 50.9572
R34377 VREFP.n9 VREFP.n8 50.9572
R34378 VREFP.n13 VREFP.n12 50.9572
R34379 VREFP.n40 VREFP.n39 50.9572
R34380 VREFP.n46 VREFP.n45 50.9572
R34381 VREFP.n51 VREFP.n50 50.9572
R34382 VREFP.n1 VREFP.n0 50.9468
R34383 VREFP.n5 VREFP.n4 50.9468
R34384 VREFP.n7 VREFP.n6 50.9468
R34385 VREFP.n11 VREFP.n10 50.9468
R34386 VREFP.n15 VREFP.n14 50.9468
R34387 VREFP.n17 VREFP.n16 50.9468
R34388 VREFP.n38 VREFP.n37 50.9468
R34389 VREFP.n42 VREFP.n41 50.9468
R34390 VREFP.n44 VREFP.n43 50.9468
R34391 VREFP.n48 VREFP.n47 50.9468
R34392 VREFP.n53 VREFP.n52 50.9468
R34393 VREFP.n55 VREFP.n54 50.9468
R34394 VREFP.n25 VREFP.t21 26.2585
R34395 VREFP.n35 VREFP.t33 26.2585
R34396 VREFP.n20 VREFP.n18 22.3849
R34397 VREFP.n30 VREFP.n28 22.3849
R34398 VREFP.n22 VREFP.n21 22.3124
R34399 VREFP.n32 VREFP.n31 22.3124
R34400 VREFP.n20 VREFP.n19 22.302
R34401 VREFP.n24 VREFP.n23 22.302
R34402 VREFP.n30 VREFP.n29 22.302
R34403 VREFP.n34 VREFP.n33 22.302
R34404 VREFP.n0 VREFP.t52 6.5015
R34405 VREFP.n0 VREFP.t50 6.5015
R34406 VREFP.n2 VREFP.t53 6.5015
R34407 VREFP.n2 VREFP.t54 6.5015
R34408 VREFP.n4 VREFP.t41 6.5015
R34409 VREFP.n4 VREFP.t55 6.5015
R34410 VREFP.n6 VREFP.t43 6.5015
R34411 VREFP.n6 VREFP.t42 6.5015
R34412 VREFP.n8 VREFP.t51 6.5015
R34413 VREFP.n8 VREFP.t49 6.5015
R34414 VREFP.n10 VREFP.t38 6.5015
R34415 VREFP.n10 VREFP.t37 6.5015
R34416 VREFP.n12 VREFP.t45 6.5015
R34417 VREFP.n12 VREFP.t39 6.5015
R34418 VREFP.n14 VREFP.t46 6.5015
R34419 VREFP.n14 VREFP.t40 6.5015
R34420 VREFP.n16 VREFP.t48 6.5015
R34421 VREFP.n16 VREFP.t47 6.5015
R34422 VREFP.n37 VREFP.t11 6.5015
R34423 VREFP.n37 VREFP.t19 6.5015
R34424 VREFP.n39 VREFP.t9 6.5015
R34425 VREFP.n39 VREFP.t18 6.5015
R34426 VREFP.n41 VREFP.t12 6.5015
R34427 VREFP.n41 VREFP.t5 6.5015
R34428 VREFP.n43 VREFP.t7 6.5015
R34429 VREFP.n43 VREFP.t13 6.5015
R34430 VREFP.n45 VREFP.t15 6.5015
R34431 VREFP.n45 VREFP.t30 6.5015
R34432 VREFP.n47 VREFP.t4 6.5015
R34433 VREFP.n47 VREFP.t17 6.5015
R34434 VREFP.n50 VREFP.t6 6.5015
R34435 VREFP.n50 VREFP.t16 6.5015
R34436 VREFP.n52 VREFP.t31 6.5015
R34437 VREFP.n52 VREFP.t8 6.5015
R34438 VREFP.n54 VREFP.t14 6.5015
R34439 VREFP.n54 VREFP.t29 6.5015
R34440 VREFP.n56 VREFP.n55 6.03712
R34441 VREFP.n26 VREFP.n17 6.03204
R34442 VREFP.n26 VREFP.n25 4.05675
R34443 VREFP.n18 VREFP.t23 3.9605
R34444 VREFP.n18 VREFP.t22 3.9605
R34445 VREFP.n19 VREFP.t26 3.9605
R34446 VREFP.n19 VREFP.t24 3.9605
R34447 VREFP.n21 VREFP.t27 3.9605
R34448 VREFP.n21 VREFP.t25 3.9605
R34449 VREFP.n23 VREFP.t20 3.9605
R34450 VREFP.n23 VREFP.t28 3.9605
R34451 VREFP.n28 VREFP.t3 3.9605
R34452 VREFP.n28 VREFP.t0 3.9605
R34453 VREFP.n29 VREFP.t2 3.9605
R34454 VREFP.n29 VREFP.t32 3.9605
R34455 VREFP.n31 VREFP.t1 3.9605
R34456 VREFP.n31 VREFP.t34 3.9605
R34457 VREFP.n33 VREFP.t35 3.9605
R34458 VREFP.n33 VREFP.t36 3.9605
R34459 VREFP.n57 VREFP.n56 3.4105
R34460 VREFP.n58 VREFP.n57 2.39545
R34461 VREFP.n57 VREFP.n35 0.64675
R34462 VREFP.n56 VREFP 0.438
R34463 VREFP VREFP.n58 0.382375
R34464 VREFP.n27 VREFP 0.2755
R34465 VREFP.n58 VREFP 0.226687
R34466 VREFP.n27 VREFP.n26 0.163
R34467 VREFP.n55 VREFP.n53 0.0954495
R34468 VREFP.n53 VREFP.n51 0.0954495
R34469 VREFP.n48 VREFP.n46 0.0954495
R34470 VREFP.n44 VREFP.n42 0.0954495
R34471 VREFP.n42 VREFP.n40 0.0954495
R34472 VREFP.n17 VREFP.n15 0.0945
R34473 VREFP.n15 VREFP.n13 0.0945
R34474 VREFP.n11 VREFP.n9 0.0945
R34475 VREFP.n7 VREFP.n5 0.0945
R34476 VREFP.n5 VREFP.n3 0.0945
R34477 VREFP.n25 VREFP.n24 0.0945
R34478 VREFP.n24 VREFP.n22 0.0945
R34479 VREFP.n35 VREFP.n34 0.0945
R34480 VREFP.n34 VREFP.n32 0.0945
R34481 VREFP.n46 VREFP.n44 0.0859545
R34482 VREFP.n40 VREFP.n38 0.0859545
R34483 VREFP.n13 VREFP.n11 0.0851
R34484 VREFP.n9 VREFP.n7 0.0851
R34485 VREFP.n3 VREFP.n1 0.0851
R34486 VREFP.n22 VREFP.n20 0.0851
R34487 VREFP.n32 VREFP.n30 0.0851
R34488 VREFP VREFP.n27 0.0652059
R34489 VREFP.n51 VREFP.n49 0.0650657
R34490 VREFP.n38 VREFP.n36 0.0484495
R34491 VREFP.n49 VREFP.n48 0.0213889
R34492 a_219318_n20038.n83 a_219318_n20038.n14 15.3734
R34493 a_219318_n20038.n83 a_219318_n20038.n78 185
R34494 a_219318_n20038.n83 a_219318_n20038.n22 91.4184
R34495 a_219318_n20038.n109 a_219318_n20038.n16 15.3734
R34496 a_219318_n20038.n109 a_219318_n20038.n104 185
R34497 a_219318_n20038.n109 a_219318_n20038.n24 91.4184
R34498 a_219318_n20038.n115 a_219318_n20038.n18 15.3734
R34499 a_219318_n20038.n115 a_219318_n20038.n110 185
R34500 a_219318_n20038.n115 a_219318_n20038.n26 91.4184
R34501 a_219318_n20038.n123 a_219318_n20038.n122 185
R34502 a_219318_n20038.n120 a_219318_n20038.n119 185
R34503 a_219318_n20038.n128 a_219318_n20038.n127 185
R34504 a_219318_n20038.n130 a_219318_n20038.n129 185
R34505 a_219318_n20038.n117 a_219318_n20038.n116 185
R34506 a_219318_n20038.n91 a_219318_n20038.n90 185
R34507 a_219318_n20038.n92 a_219318_n20038.n85 185
R34508 a_219318_n20038.n101 a_219318_n20038.n100 185
R34509 a_219318_n20038.n99 a_219318_n20038.n98 185
R34510 a_219318_n20038.n94 a_219318_n20038.n93 185
R34511 a_219318_n20038.n32 a_219318_n20038.n170 91.4185
R34512 a_219318_n20038.n56 a_219318_n20038.n170 14.3253
R34513 a_219318_n20038.n34 a_219318_n20038.n167 91.4185
R34514 a_219318_n20038.n58 a_219318_n20038.n167 14.3253
R34515 a_219318_n20038.n36 a_219318_n20038.n164 91.4185
R34516 a_219318_n20038.n60 a_219318_n20038.n164 14.3253
R34517 a_219318_n20038.n38 a_219318_n20038.n161 91.4185
R34518 a_219318_n20038.n62 a_219318_n20038.n161 14.3253
R34519 a_219318_n20038.n40 a_219318_n20038.n158 91.4185
R34520 a_219318_n20038.n64 a_219318_n20038.n158 14.3253
R34521 a_219318_n20038.n42 a_219318_n20038.n155 91.4185
R34522 a_219318_n20038.n66 a_219318_n20038.n155 14.3253
R34523 a_219318_n20038.n154 a_219318_n20038.n153 185
R34524 a_219318_n20038.n151 a_219318_n20038.n137 185
R34525 a_219318_n20038.n141 a_219318_n20038.n138 185
R34526 a_219318_n20038.n146 a_219318_n20038.n145 185
R34527 a_219318_n20038.n144 a_219318_n20038.n143 185
R34528 a_219318_n20038.n178 a_219318_n20038.n177 185
R34529 a_219318_n20038.n185 a_219318_n20038.n184 185
R34530 a_219318_n20038.n186 a_219318_n20038.n175 185
R34531 a_219318_n20038.n191 a_219318_n20038.n190 185
R34532 a_219318_n20038.n189 a_219318_n20038.n188 185
R34533 a_219318_n20038.n48 a_219318_n20038.n193 91.4187
R34534 a_219318_n20038.n194 a_219318_n20038.n193 185
R34535 a_219318_n20038.n8 a_219318_n20038.n193 15.371
R34536 a_219318_n20038.n50 a_219318_n20038.n72 91.4187
R34537 a_219318_n20038.n73 a_219318_n20038.n72 185
R34538 a_219318_n20038.n10 a_219318_n20038.n72 15.371
R34539 a_219318_n20038.n200 a_219318_n20038.n52 91.4187
R34540 a_219318_n20038.n200 a_219318_n20038.n69 185
R34541 a_219318_n20038.n200 a_219318_n20038.n12 15.371
R34542 a_219318_n20038.t15 a_219318_n20038.n121 174.857
R34543 a_219318_n20038.n95 a_219318_n20038.t0 174.857
R34544 a_219318_n20038.n142 a_219318_n20038.t12 174.857
R34545 a_219318_n20038.n187 a_219318_n20038.t23 174.857
R34546 a_219318_n20038.n122 a_219318_n20038.n119 140.69
R34547 a_219318_n20038.n128 a_219318_n20038.n119 140.69
R34548 a_219318_n20038.n129 a_219318_n20038.n128 140.69
R34549 a_219318_n20038.n129 a_219318_n20038.n116 140.69
R34550 a_219318_n20038.n28 a_219318_n20038.n116 256.962
R34551 a_219318_n20038.n91 a_219318_n20038.n30 256.962
R34552 a_219318_n20038.n92 a_219318_n20038.n91 140.69
R34553 a_219318_n20038.n100 a_219318_n20038.n92 140.69
R34554 a_219318_n20038.n100 a_219318_n20038.n99 140.69
R34555 a_219318_n20038.n99 a_219318_n20038.n93 140.69
R34556 a_219318_n20038.n43 a_219318_n20038.n154 256.962
R34557 a_219318_n20038.n154 a_219318_n20038.n137 140.69
R34558 a_219318_n20038.n141 a_219318_n20038.n137 140.69
R34559 a_219318_n20038.n145 a_219318_n20038.n141 140.69
R34560 a_219318_n20038.n145 a_219318_n20038.n144 140.69
R34561 a_219318_n20038.n46 a_219318_n20038.n177 256.962
R34562 a_219318_n20038.n185 a_219318_n20038.n177 140.69
R34563 a_219318_n20038.n186 a_219318_n20038.n185 140.69
R34564 a_219318_n20038.n190 a_219318_n20038.n186 140.69
R34565 a_219318_n20038.n190 a_219318_n20038.n189 140.69
R34566 a_219318_n20038.n122 a_219318_n20038.t15 70.3453
R34567 a_219318_n20038.t0 a_219318_n20038.n93 70.3453
R34568 a_219318_n20038.n144 a_219318_n20038.t12 70.3453
R34569 a_219318_n20038.n189 a_219318_n20038.t23 70.3453
R34570 a_219318_n20038.n123 a_219318_n20038.n121 28.4333
R34571 a_219318_n20038.n95 a_219318_n20038.n94 28.4333
R34572 a_219318_n20038.n143 a_219318_n20038.n142 28.4333
R34573 a_219318_n20038.n188 a_219318_n20038.n187 28.4333
R34574 a_219318_n20038.n14 a_219318_n20038.n13 3.21237
R34575 a_219318_n20038.n124 a_219318_n20038.n120 24.8476
R34576 a_219318_n20038.n98 a_219318_n20038.n97 24.8476
R34577 a_219318_n20038.n146 a_219318_n20038.n140 24.8476
R34578 a_219318_n20038.n191 a_219318_n20038.n176 24.8476
R34579 a_219318_n20038.n127 a_219318_n20038.n126 23.3417
R34580 a_219318_n20038.n101 a_219318_n20038.n86 23.3417
R34581 a_219318_n20038.n147 a_219318_n20038.n138 23.3417
R34582 a_219318_n20038.n192 a_219318_n20038.n175 23.3417
R34583 a_219318_n20038.n14 a_219318_n20038.n81 27.6334
R34584 a_219318_n20038.n16 a_219318_n20038.n107 27.6334
R34585 a_219318_n20038.n18 a_219318_n20038.n113 27.6334
R34586 a_219318_n20038.n130 a_219318_n20038.n118 21.8358
R34587 a_219318_n20038.n102 a_219318_n20038.n85 21.8358
R34588 a_219318_n20038.n151 a_219318_n20038.n150 21.8358
R34589 a_219318_n20038.n184 a_219318_n20038.n183 21.8358
R34590 a_219318_n20038.n81 a_219318_n20038.n78 20.3299
R34591 a_219318_n20038.n107 a_219318_n20038.n104 20.3299
R34592 a_219318_n20038.n113 a_219318_n20038.n110 20.3299
R34593 a_219318_n20038.n131 a_219318_n20038.n117 20.3299
R34594 a_219318_n20038.n90 a_219318_n20038.n89 20.3299
R34595 a_219318_n20038.n153 a_219318_n20038.n152 20.3299
R34596 a_219318_n20038.n182 a_219318_n20038.n178 20.3299
R34597 a_219318_n20038.n198 a_219318_n20038.n194 20.3299
R34598 a_219318_n20038.n77 a_219318_n20038.n73 20.3299
R34599 a_219318_n20038.n70 a_219318_n20038.n69 20.3299
R34600 a_219318_n20038.n79 a_219318_n20038.n22 24.4363
R34601 a_219318_n20038.n105 a_219318_n20038.n24 24.4363
R34602 a_219318_n20038.n111 a_219318_n20038.n26 24.4363
R34603 a_219318_n20038.n28 a_219318_n20038.n134 22.9459
R34604 a_219318_n20038.n22 a_219318_n20038.n21 9.72509
R34605 a_219318_n20038.n24 a_219318_n20038.n23 9.72509
R34606 a_219318_n20038.n26 a_219318_n20038.n25 9.72509
R34607 a_219318_n20038.n28 a_219318_n20038.n27 11.3106
R34608 a_219318_n20038.n29 a_219318_n20038.n30 11.3108
R34609 a_219318_n20038.n31 a_219318_n20038.n32 9.72532
R34610 a_219318_n20038.n33 a_219318_n20038.n34 9.72532
R34611 a_219318_n20038.n35 a_219318_n20038.n36 9.72532
R34612 a_219318_n20038.n37 a_219318_n20038.n38 9.72532
R34613 a_219318_n20038.n39 a_219318_n20038.n40 9.72532
R34614 a_219318_n20038.n41 a_219318_n20038.n42 9.72532
R34615 a_219318_n20038.n44 a_219318_n20038.n43 11.3108
R34616 a_219318_n20038.n46 a_219318_n20038.n45 11.3109
R34617 a_219318_n20038.n47 a_219318_n20038.n48 9.72555
R34618 a_219318_n20038.n49 a_219318_n20038.n50 9.72555
R34619 a_219318_n20038.n53 a_219318_n20038.n52 9.72555
R34620 a_219318_n20038.n16 a_219318_n20038.n15 3.21237
R34621 a_219318_n20038.n18 a_219318_n20038.n17 3.21237
R34622 a_219318_n20038.n7 a_219318_n20038.n8 3.21131
R34623 a_219318_n20038.n9 a_219318_n20038.n10 3.21131
R34624 a_219318_n20038.n12 a_219318_n20038.n11 3.21131
R34625 a_219318_n20038.n55 a_219318_n20038.n56 2.85029
R34626 a_219318_n20038.n57 a_219318_n20038.n58 2.85029
R34627 a_219318_n20038.n59 a_219318_n20038.n60 2.85029
R34628 a_219318_n20038.n61 a_219318_n20038.n62 2.85029
R34629 a_219318_n20038.n63 a_219318_n20038.n64 2.85029
R34630 a_219318_n20038.n65 a_219318_n20038.n66 2.85029
R34631 a_219318_n20038.n82 a_219318_n20038.n81 9.3005
R34632 a_219318_n20038.n80 a_219318_n20038.n79 9.3005
R34633 a_219318_n20038.n108 a_219318_n20038.n107 9.3005
R34634 a_219318_n20038.n106 a_219318_n20038.n105 9.3005
R34635 a_219318_n20038.n114 a_219318_n20038.n113 9.3005
R34636 a_219318_n20038.n112 a_219318_n20038.n111 9.3005
R34637 a_219318_n20038.n125 a_219318_n20038.n124 9.3005
R34638 a_219318_n20038.n118 a_219318_n20038.n3 9.3005
R34639 a_219318_n20038.n132 a_219318_n20038.n131 9.3005
R34640 a_219318_n20038.n134 a_219318_n20038.n133 9.3005
R34641 a_219318_n20038.n126 a_219318_n20038.n3 9.3005
R34642 a_219318_n20038.n97 a_219318_n20038.n96 9.3005
R34643 a_219318_n20038.n86 a_219318_n20038.n84 9.3005
R34644 a_219318_n20038.n103 a_219318_n20038.n102 9.3005
R34645 a_219318_n20038.n89 a_219318_n20038.n54 9.3005
R34646 a_219318_n20038.n88 a_219318_n20038.n87 9.3005
R34647 a_219318_n20038.n172 a_219318_n20038.n171 9.3005
R34648 a_219318_n20038.n169 a_219318_n20038.n168 9.3005
R34649 a_219318_n20038.n166 a_219318_n20038.n165 9.3005
R34650 a_219318_n20038.n163 a_219318_n20038.n162 9.3005
R34651 a_219318_n20038.n160 a_219318_n20038.n159 9.3005
R34652 a_219318_n20038.n157 a_219318_n20038.n156 9.3005
R34653 a_219318_n20038.n140 a_219318_n20038.n139 9.3005
R34654 a_219318_n20038.n148 a_219318_n20038.n147 9.3005
R34655 a_219318_n20038.n150 a_219318_n20038.n149 9.3005
R34656 a_219318_n20038.n152 a_219318_n20038.n68 9.3005
R34657 a_219318_n20038.n136 a_219318_n20038.n67 9.3005
R34658 a_219318_n20038.n176 a_219318_n20038.n174 9.3005
R34659 a_219318_n20038.n2 a_219318_n20038.n192 9.3005
R34660 a_219318_n20038.n183 a_219318_n20038.n2 9.3005
R34661 a_219318_n20038.n182 a_219318_n20038.n181 9.3005
R34662 a_219318_n20038.n180 a_219318_n20038.n179 9.3005
R34663 a_219318_n20038.n198 a_219318_n20038.n197 9.3005
R34664 a_219318_n20038.n196 a_219318_n20038.n195 9.3005
R34665 a_219318_n20038.n77 a_219318_n20038.n76 9.3005
R34666 a_219318_n20038.n75 a_219318_n20038.n74 9.3005
R34667 a_219318_n20038.n71 a_219318_n20038.n70 9.3005
R34668 a_219318_n20038.n199 a_219318_n20038.n51 9.3005
R34669 a_219318_n20038.n30 a_219318_n20038.n88 22.9458
R34670 a_219318_n20038.n32 a_219318_n20038.n172 24.4362
R34671 a_219318_n20038.n34 a_219318_n20038.n169 24.4362
R34672 a_219318_n20038.n36 a_219318_n20038.n166 24.4362
R34673 a_219318_n20038.n38 a_219318_n20038.n163 24.4362
R34674 a_219318_n20038.n40 a_219318_n20038.n160 24.4362
R34675 a_219318_n20038.n42 a_219318_n20038.n157 24.4362
R34676 a_219318_n20038.n43 a_219318_n20038.n136 22.9458
R34677 a_219318_n20038.n179 a_219318_n20038.n46 22.9457
R34678 a_219318_n20038.n195 a_219318_n20038.n48 24.4361
R34679 a_219318_n20038.n74 a_219318_n20038.n50 24.4361
R34680 a_219318_n20038.n52 a_219318_n20038.n51 24.4361
R34681 a_219318_n20038.n1 a_219318_n20038.n13 7.9105
R34682 a_219318_n20038.n1 a_219318_n20038.n15 7.9105
R34683 a_219318_n20038.n1 a_219318_n20038.n17 7.9105
R34684 a_219318_n20038.n1 a_219318_n20038.n3 7.9105
R34685 a_219318_n20038.n1 a_219318_n20038.n27 7.9105
R34686 a_219318_n20038.n1 a_219318_n20038.n25 7.9105
R34687 a_219318_n20038.n1 a_219318_n20038.n23 7.9105
R34688 a_219318_n20038.n1 a_219318_n20038.n21 7.9105
R34689 a_219318_n20038.n6 a_219318_n20038.n31 7.9105
R34690 a_219318_n20038.n6 a_219318_n20038.n33 7.9105
R34691 a_219318_n20038.n5 a_219318_n20038.n35 7.9105
R34692 a_219318_n20038.n5 a_219318_n20038.n37 7.9105
R34693 a_219318_n20038.n4 a_219318_n20038.n39 7.9105
R34694 a_219318_n20038.n4 a_219318_n20038.n41 7.9105
R34695 a_219318_n20038.n4 a_219318_n20038.n65 7.9105
R34696 a_219318_n20038.n4 a_219318_n20038.n63 7.9105
R34697 a_219318_n20038.n5 a_219318_n20038.n61 7.9105
R34698 a_219318_n20038.n5 a_219318_n20038.n59 7.9105
R34699 a_219318_n20038.n6 a_219318_n20038.n57 7.9105
R34700 a_219318_n20038.n6 a_219318_n20038.n55 7.9105
R34701 a_219318_n20038.n0 a_219318_n20038.n45 7.9105
R34702 a_219318_n20038.n0 a_219318_n20038.n47 7.9105
R34703 a_219318_n20038.n0 a_219318_n20038.n49 7.9105
R34704 a_219318_n20038.n0 a_219318_n20038.n9 7.9105
R34705 a_219318_n20038.n0 a_219318_n20038.n7 7.9105
R34706 a_219318_n20038.n0 a_219318_n20038.n2 7.9105
R34707 a_219318_n20038.n0 a_219318_n20038.n53 7.9105
R34708 a_219318_n20038.n11 a_219318_n20038.n0 7.9105
R34709 a_219318_n20038.n79 a_219318_n20038.n78 6.77697
R34710 a_219318_n20038.n105 a_219318_n20038.n104 6.77697
R34711 a_219318_n20038.n111 a_219318_n20038.n110 6.77697
R34712 a_219318_n20038.n134 a_219318_n20038.n117 6.77697
R34713 a_219318_n20038.n90 a_219318_n20038.n88 6.77697
R34714 a_219318_n20038.n56 a_219318_n20038.n172 28.3048
R34715 a_219318_n20038.n58 a_219318_n20038.n169 28.3048
R34716 a_219318_n20038.n60 a_219318_n20038.n166 28.3048
R34717 a_219318_n20038.n62 a_219318_n20038.n163 28.3048
R34718 a_219318_n20038.n64 a_219318_n20038.n160 28.3048
R34719 a_219318_n20038.n66 a_219318_n20038.n157 28.3048
R34720 a_219318_n20038.n153 a_219318_n20038.n136 6.77697
R34721 a_219318_n20038.n179 a_219318_n20038.n178 6.77697
R34722 a_219318_n20038.n195 a_219318_n20038.n194 6.77697
R34723 a_219318_n20038.n74 a_219318_n20038.n73 6.77697
R34724 a_219318_n20038.n51 a_219318_n20038.n69 6.77697
R34725 a_219318_n20038.n125 a_219318_n20038.n121 5.33935
R34726 a_219318_n20038.n96 a_219318_n20038.n95 5.33935
R34727 a_219318_n20038.n142 a_219318_n20038.n139 5.33935
R34728 a_219318_n20038.n187 a_219318_n20038.n174 5.33935
R34729 a_219318_n20038.n131 a_219318_n20038.n130 5.27109
R34730 a_219318_n20038.n89 a_219318_n20038.n85 5.27109
R34731 a_219318_n20038.n152 a_219318_n20038.n151 5.27109
R34732 a_219318_n20038.n184 a_219318_n20038.n182 5.27109
R34733 a_219318_n20038.n8 a_219318_n20038.n198 27.6341
R34734 a_219318_n20038.n10 a_219318_n20038.n77 27.6341
R34735 a_219318_n20038.n12 a_219318_n20038.n70 27.6341
R34736 a_219318_n20038.n19 a_219318_n20038.n54 4.56989
R34737 a_219318_n20038.n20 a_219318_n20038.n68 4.56989
R34738 a_219318_n20038.n19 a_219318_n20038.n29 4.5005
R34739 a_219318_n20038.n20 a_219318_n20038.n44 4.5005
R34740 a_219318_n20038.n127 a_219318_n20038.n118 3.76521
R34741 a_219318_n20038.n102 a_219318_n20038.n101 3.76521
R34742 a_219318_n20038.n150 a_219318_n20038.n138 3.76521
R34743 a_219318_n20038.n183 a_219318_n20038.n175 3.76521
R34744 a_219318_n20038.n83 a_219318_n20038.t4 3.4805
R34745 a_219318_n20038.n83 a_219318_n20038.t1 3.4805
R34746 a_219318_n20038.n109 a_219318_n20038.t14 3.4805
R34747 a_219318_n20038.n109 a_219318_n20038.t2 3.4805
R34748 a_219318_n20038.n115 a_219318_n20038.t11 3.4805
R34749 a_219318_n20038.n115 a_219318_n20038.t17 3.4805
R34750 a_219318_n20038.n170 a_219318_n20038.t25 3.4805
R34751 a_219318_n20038.n170 a_219318_n20038.t3 3.4805
R34752 a_219318_n20038.n167 a_219318_n20038.t6 3.4805
R34753 a_219318_n20038.n167 a_219318_n20038.t9 3.4805
R34754 a_219318_n20038.n164 a_219318_n20038.t13 3.4805
R34755 a_219318_n20038.n164 a_219318_n20038.t5 3.4805
R34756 a_219318_n20038.n161 a_219318_n20038.t8 3.4805
R34757 a_219318_n20038.n161 a_219318_n20038.t7 3.4805
R34758 a_219318_n20038.n158 a_219318_n20038.t10 3.4805
R34759 a_219318_n20038.n158 a_219318_n20038.t27 3.4805
R34760 a_219318_n20038.n155 a_219318_n20038.t16 3.4805
R34761 a_219318_n20038.n155 a_219318_n20038.t26 3.4805
R34762 a_219318_n20038.n193 a_219318_n20038.t19 3.4805
R34763 a_219318_n20038.n193 a_219318_n20038.t18 3.4805
R34764 a_219318_n20038.n72 a_219318_n20038.t22 3.4805
R34765 a_219318_n20038.n72 a_219318_n20038.t21 3.4805
R34766 a_219318_n20038.n200 a_219318_n20038.t20 3.4805
R34767 a_219318_n20038.t24 a_219318_n20038.n200 3.4805
R34768 a_219318_n20038.n135 a_219318_n20038.n1 2.68111
R34769 a_219318_n20038.n173 a_219318_n20038.n1 2.5834
R34770 a_219318_n20038.n173 a_219318_n20038.n19 2.26061
R34771 a_219318_n20038.n20 a_219318_n20038.n135 2.26061
R34772 a_219318_n20038.n126 a_219318_n20038.n120 2.25932
R34773 a_219318_n20038.n98 a_219318_n20038.n86 2.25932
R34774 a_219318_n20038.n147 a_219318_n20038.n146 2.25932
R34775 a_219318_n20038.n192 a_219318_n20038.n191 2.25932
R34776 a_219318_n20038.n0 a_219318_n20038.n173 1.93434
R34777 a_219318_n20038.n135 a_219318_n20038.n0 1.83663
R34778 a_219318_n20038.n19 a_219318_n20038.n6 1.83146
R34779 a_219318_n20038.n4 a_219318_n20038.n20 1.82972
R34780 a_219318_n20038.n124 a_219318_n20038.n123 0.753441
R34781 a_219318_n20038.n97 a_219318_n20038.n94 0.753441
R34782 a_219318_n20038.n143 a_219318_n20038.n140 0.753441
R34783 a_219318_n20038.n188 a_219318_n20038.n176 0.753441
R34784 a_219318_n20038.n3 a_219318_n20038.n125 0.298809
R34785 a_219318_n20038.n2 a_219318_n20038.n174 0.298809
R34786 a_219318_n20038.n11 a_219318_n20038.n71 0.274655
R34787 a_219318_n20038.n76 a_219318_n20038.n9 0.274655
R34788 a_219318_n20038.n197 a_219318_n20038.n7 0.274655
R34789 a_219318_n20038.n5 a_219318_n20038.n4 0.270315
R34790 a_219318_n20038.n17 a_219318_n20038.n114 0.26922
R34791 a_219318_n20038.n15 a_219318_n20038.n108 0.26922
R34792 a_219318_n20038.n13 a_219318_n20038.n82 0.26922
R34793 a_219318_n20038.n133 a_219318_n20038.n27 0.231176
R34794 a_219318_n20038.n112 a_219318_n20038.n25 0.231176
R34795 a_219318_n20038.n106 a_219318_n20038.n23 0.231176
R34796 a_219318_n20038.n80 a_219318_n20038.n21 0.231176
R34797 a_219318_n20038.n44 a_219318_n20038.n67 0.228459
R34798 a_219318_n20038.n156 a_219318_n20038.n41 0.228459
R34799 a_219318_n20038.n159 a_219318_n20038.n39 0.228459
R34800 a_219318_n20038.n162 a_219318_n20038.n37 0.228459
R34801 a_219318_n20038.n165 a_219318_n20038.n35 0.228459
R34802 a_219318_n20038.n168 a_219318_n20038.n33 0.228459
R34803 a_219318_n20038.n171 a_219318_n20038.n31 0.228459
R34804 a_219318_n20038.n87 a_219318_n20038.n29 0.228459
R34805 a_219318_n20038.n53 a_219318_n20038.n199 0.225742
R34806 a_219318_n20038.n75 a_219318_n20038.n49 0.225742
R34807 a_219318_n20038.n196 a_219318_n20038.n47 0.225742
R34808 a_219318_n20038.n180 a_219318_n20038.n45 0.225742
R34809 a_219318_n20038.n82 a_219318_n20038.n80 0.196152
R34810 a_219318_n20038.n108 a_219318_n20038.n106 0.196152
R34811 a_219318_n20038.n114 a_219318_n20038.n112 0.196152
R34812 a_219318_n20038.n132 a_219318_n20038.n3 0.196152
R34813 a_219318_n20038.n133 a_219318_n20038.n132 0.196152
R34814 a_219318_n20038.n103 a_219318_n20038.n84 0.196152
R34815 a_219318_n20038.n96 a_219318_n20038.n84 0.196152
R34816 a_219318_n20038.n149 a_219318_n20038.n148 0.196152
R34817 a_219318_n20038.n148 a_219318_n20038.n139 0.196152
R34818 a_219318_n20038.n181 a_219318_n20038.n180 0.196152
R34819 a_219318_n20038.n181 a_219318_n20038.n2 0.196152
R34820 a_219318_n20038.n197 a_219318_n20038.n196 0.196152
R34821 a_219318_n20038.n76 a_219318_n20038.n75 0.196152
R34822 a_219318_n20038.n199 a_219318_n20038.n71 0.196152
R34823 a_219318_n20038.n6 a_219318_n20038.n5 0.179796
R34824 a_219318_n20038.n156 a_219318_n20038.n65 0.168676
R34825 a_219318_n20038.n159 a_219318_n20038.n63 0.168676
R34826 a_219318_n20038.n162 a_219318_n20038.n61 0.168676
R34827 a_219318_n20038.n165 a_219318_n20038.n59 0.168676
R34828 a_219318_n20038.n168 a_219318_n20038.n57 0.168676
R34829 a_219318_n20038.n171 a_219318_n20038.n55 0.168676
R34830 a_219318_n20038.n87 a_219318_n20038.n54 0.158954
R34831 a_219318_n20038.n68 a_219318_n20038.n67 0.158954
R34832 a_219318_n20038.n149 a_219318_n20038.n68 0.140355
R34833 a_219318_n20038.n54 a_219318_n20038.n103 0.140355
R34834 a_188130_n13996.n66 a_188130_n13996.n60 585
R34835 a_188130_n13996.n66 a_188130_n13996.n17 291.382
R34836 a_188130_n13996.n349 a_188130_n13996.n348 585
R34837 a_188130_n13996.n348 a_188130_n13996.n347 585
R34838 a_188130_n13996.n348 a_188130_n13996.n99 585
R34839 a_188130_n13996.n348 a_188130_n13996.n98 585
R34840 a_188130_n13996.n348 a_188130_n13996.n97 585
R34841 a_188130_n13996.n348 a_188130_n13996.n96 585
R34842 a_188130_n13996.n348 a_188130_n13996.n94 585
R34843 a_188130_n13996.n348 a_188130_n13996.n93 585
R34844 a_188130_n13996.n348 a_188130_n13996.n92 585
R34845 a_188130_n13996.n348 a_188130_n13996.n91 585
R34846 a_188130_n13996.n348 a_188130_n13996.n90 585
R34847 a_188130_n13996.n348 a_188130_n13996.n89 585
R34848 a_188130_n13996.n273 a_188130_n13996.n272 585
R34849 a_188130_n13996.n273 a_188130_n13996.n118 585
R34850 a_188130_n13996.n273 a_188130_n13996.n117 585
R34851 a_188130_n13996.n273 a_188130_n13996.n116 585
R34852 a_188130_n13996.n273 a_188130_n13996.n115 585
R34853 a_188130_n13996.n273 a_188130_n13996.n114 585
R34854 a_188130_n13996.n273 a_188130_n13996.n112 585
R34855 a_188130_n13996.n273 a_188130_n13996.n111 585
R34856 a_188130_n13996.n273 a_188130_n13996.n110 585
R34857 a_188130_n13996.n273 a_188130_n13996.n109 585
R34858 a_188130_n13996.n273 a_188130_n13996.n108 585
R34859 a_188130_n13996.n274 a_188130_n13996.n273 585
R34860 a_188130_n13996.n179 a_188130_n13996.n178 585
R34861 a_188130_n13996.n178 a_188130_n13996.n177 585
R34862 a_188130_n13996.n178 a_188130_n13996.n134 585
R34863 a_188130_n13996.n178 a_188130_n13996.n133 585
R34864 a_188130_n13996.n178 a_188130_n13996.n132 585
R34865 a_188130_n13996.n178 a_188130_n13996.n131 585
R34866 a_188130_n13996.n178 a_188130_n13996.n129 585
R34867 a_188130_n13996.n178 a_188130_n13996.n128 585
R34868 a_188130_n13996.n178 a_188130_n13996.n127 585
R34869 a_188130_n13996.n178 a_188130_n13996.n126 585
R34870 a_188130_n13996.n178 a_188130_n13996.n125 585
R34871 a_188130_n13996.n178 a_188130_n13996.n124 585
R34872 a_188130_n13996.n378 a_188130_n13996.n377 585
R34873 a_188130_n13996.n378 a_188130_n13996.n82 585
R34874 a_188130_n13996.n378 a_188130_n13996.n81 585
R34875 a_188130_n13996.n378 a_188130_n13996.n80 585
R34876 a_188130_n13996.n378 a_188130_n13996.n79 585
R34877 a_188130_n13996.n378 a_188130_n13996.n78 585
R34878 a_188130_n13996.n378 a_188130_n13996.n76 585
R34879 a_188130_n13996.n378 a_188130_n13996.n75 585
R34880 a_188130_n13996.n378 a_188130_n13996.n69 585
R34881 a_188130_n13996.n379 a_188130_n13996.n378 585
R34882 a_188130_n13996.n378 a_188130_n13996.n73 585
R34883 a_188130_n13996.n378 a_188130_n13996.n71 585
R34884 a_188130_n13996.n389 a_188130_n13996.n383 585
R34885 a_188130_n13996.n389 a_188130_n13996.n26 291.382
R34886 a_188130_n13996.n397 a_188130_n13996.n391 585
R34887 a_188130_n13996.n397 a_188130_n13996.n28 291.382
R34888 a_188130_n13996.n405 a_188130_n13996.n399 585
R34889 a_188130_n13996.n405 a_188130_n13996.n30 291.382
R34890 a_188130_n13996.n49 a_188130_n13996.n43 585
R34891 a_188130_n13996.n49 a_188130_n13996.n32 291.382
R34892 a_188130_n13996.n143 a_188130_n13996.n142 585
R34893 a_188130_n13996.n140 a_188130_n13996.n139 585
R34894 a_188130_n13996.n149 a_188130_n13996.n148 585
R34895 a_188130_n13996.n151 a_188130_n13996.n150 585
R34896 a_188130_n13996.n138 a_188130_n13996.n137 585
R34897 a_188130_n13996.n408 a_188130_n13996.n41 585
R34898 a_188130_n13996.n408 a_188130_n13996.n36 291.382
R34899 a_188130_n13996.t6 a_188130_n13996.n190 433.543
R34900 a_188130_n13996.t30 a_188130_n13996.n211 433.543
R34901 a_188130_n13996.n191 a_188130_n13996.t6 433.351
R34902 a_188130_n13996.n235 a_188130_n13996.t22 433.149
R34903 a_188130_n13996.n353 a_188130_n13996.t24 433.149
R34904 a_188130_n13996.t24 a_188130_n13996.n352 433.149
R34905 a_188130_n13996.n354 a_188130_n13996.t28 433.149
R34906 a_188130_n13996.t28 a_188130_n13996.n83 433.149
R34907 a_188130_n13996.n194 a_188130_n13996.t66 433.149
R34908 a_188130_n13996.t66 a_188130_n13996.n192 433.149
R34909 a_188130_n13996.t42 a_188130_n13996.n119 433.149
R34910 a_188130_n13996.n190 a_188130_n13996.t42 433.149
R34911 a_188130_n13996.n246 a_188130_n13996.t12 433.149
R34912 a_188130_n13996.t12 a_188130_n13996.n120 433.149
R34913 a_188130_n13996.t14 a_188130_n13996.n247 433.149
R34914 a_188130_n13996.n248 a_188130_n13996.t14 433.149
R34915 a_188130_n13996.t36 a_188130_n13996.n183 433.149
R34916 a_188130_n13996.n236 a_188130_n13996.t36 433.149
R34917 a_188130_n13996.n238 a_188130_n13996.t44 433.149
R34918 a_188130_n13996.t44 a_188130_n13996.n237 433.149
R34919 a_188130_n13996.n239 a_188130_n13996.t10 433.149
R34920 a_188130_n13996.t10 a_188130_n13996.n182 433.149
R34921 a_188130_n13996.t20 a_188130_n13996.n240 433.149
R34922 a_188130_n13996.n241 a_188130_n13996.t20 433.149
R34923 a_188130_n13996.t26 a_188130_n13996.n121 433.149
R34924 a_188130_n13996.n242 a_188130_n13996.t26 433.149
R34925 a_188130_n13996.n244 a_188130_n13996.t38 433.149
R34926 a_188130_n13996.t38 a_188130_n13996.n243 433.149
R34927 a_188130_n13996.t34 a_188130_n13996.n357 433.149
R34928 a_188130_n13996.n358 a_188130_n13996.t34 433.149
R34929 a_188130_n13996.n85 a_188130_n13996.t32 433.149
R34930 a_188130_n13996.t32 a_188130_n13996.n84 433.149
R34931 a_188130_n13996.t40 a_188130_n13996.n229 433.149
R34932 a_188130_n13996.n230 a_188130_n13996.t40 433.149
R34933 a_188130_n13996.n232 a_188130_n13996.t4 433.149
R34934 a_188130_n13996.t4 a_188130_n13996.n231 433.149
R34935 a_188130_n13996.n233 a_188130_n13996.t16 433.149
R34936 a_188130_n13996.t16 a_188130_n13996.n184 433.149
R34937 a_188130_n13996.t55 a_188130_n13996.n227 433.149
R34938 a_188130_n13996.n228 a_188130_n13996.t55 433.149
R34939 a_188130_n13996.t57 a_188130_n13996.n215 433.149
R34940 a_188130_n13996.n216 a_188130_n13996.t57 433.149
R34941 a_188130_n13996.t54 a_188130_n13996.n209 433.149
R34942 a_188130_n13996.n217 a_188130_n13996.t54 433.149
R34943 a_188130_n13996.n219 a_188130_n13996.t52 433.149
R34944 a_188130_n13996.t52 a_188130_n13996.n218 433.149
R34945 a_188130_n13996.n220 a_188130_n13996.t49 433.149
R34946 a_188130_n13996.t49 a_188130_n13996.n208 433.149
R34947 a_188130_n13996.t50 a_188130_n13996.n221 433.149
R34948 a_188130_n13996.n222 a_188130_n13996.t50 433.149
R34949 a_188130_n13996.t67 a_188130_n13996.n207 433.149
R34950 a_188130_n13996.n223 a_188130_n13996.t67 433.149
R34951 a_188130_n13996.n225 a_188130_n13996.t64 433.149
R34952 a_188130_n13996.t64 a_188130_n13996.n224 433.149
R34953 a_188130_n13996.n226 a_188130_n13996.t58 433.149
R34954 a_188130_n13996.t58 a_188130_n13996.n186 433.149
R34955 a_188130_n13996.n206 a_188130_n13996.t69 433.149
R34956 a_188130_n13996.t69 a_188130_n13996.n185 433.149
R34957 a_188130_n13996.n205 a_188130_n13996.t65 433.149
R34958 a_188130_n13996.t65 a_188130_n13996.n204 433.149
R34959 a_188130_n13996.t61 a_188130_n13996.n187 433.149
R34960 a_188130_n13996.n203 a_188130_n13996.t61 433.149
R34961 a_188130_n13996.t56 a_188130_n13996.n201 433.149
R34962 a_188130_n13996.n202 a_188130_n13996.t56 433.149
R34963 a_188130_n13996.n200 a_188130_n13996.t53 433.149
R34964 a_188130_n13996.t53 a_188130_n13996.n188 433.149
R34965 a_188130_n13996.n199 a_188130_n13996.t68 433.149
R34966 a_188130_n13996.t68 a_188130_n13996.n198 433.149
R34967 a_188130_n13996.t60 a_188130_n13996.n189 433.149
R34968 a_188130_n13996.n197 a_188130_n13996.t60 433.149
R34969 a_188130_n13996.t59 a_188130_n13996.n195 433.149
R34970 a_188130_n13996.n196 a_188130_n13996.t59 433.149
R34971 a_188130_n13996.t22 a_188130_n13996.n234 433.149
R34972 a_188130_n13996.n214 a_188130_n13996.t62 433.149
R34973 a_188130_n13996.t62 a_188130_n13996.n212 433.149
R34974 a_188130_n13996.n39 a_188130_n13996.t30 433.149
R34975 a_188130_n13996.t18 a_188130_n13996.n38 433.149
R34976 a_188130_n13996.n210 a_188130_n13996.t18 433.149
R34977 a_188130_n13996.n211 a_188130_n13996.t8 433.149
R34978 a_188130_n13996.n39 a_188130_n13996.t8 433.149
R34979 a_188130_n13996.t7 a_188130_n13996.n141 384.339
R34980 a_188130_n13996.n348 a_188130_n13996.n95 286.238
R34981 a_188130_n13996.n273 a_188130_n13996.n113 286.238
R34982 a_188130_n13996.n178 a_188130_n13996.n130 286.238
R34983 a_188130_n13996.n378 a_188130_n13996.n77 286.238
R34984 a_188130_n13996.n142 a_188130_n13996.n139 230.966
R34985 a_188130_n13996.n149 a_188130_n13996.n139 230.966
R34986 a_188130_n13996.n150 a_188130_n13996.n149 230.966
R34987 a_188130_n13996.n150 a_188130_n13996.n137 230.966
R34988 a_188130_n13996.n34 a_188130_n13996.n137 570.105
R34989 a_188130_n13996.n193 a_188130_n13996.t63 215.964
R34990 a_188130_n13996.n213 a_188130_n13996.t51 215.963
R34991 a_188130_n13996.n329 a_188130_n13996.n321 185
R34992 a_188130_n13996.n329 a_188130_n13996.n320 185
R34993 a_188130_n13996.n329 a_188130_n13996.n8 91.4184
R34994 a_188130_n13996.n318 a_188130_n13996.n310 185
R34995 a_188130_n13996.n318 a_188130_n13996.n309 185
R34996 a_188130_n13996.n318 a_188130_n13996.n10 91.4184
R34997 a_188130_n13996.n307 a_188130_n13996.n299 185
R34998 a_188130_n13996.n307 a_188130_n13996.n298 185
R34999 a_188130_n13996.n307 a_188130_n13996.n12 91.4184
R35000 a_188130_n13996.n285 a_188130_n13996.n284 185
R35001 a_188130_n13996.n282 a_188130_n13996.n281 185
R35002 a_188130_n13996.n290 a_188130_n13996.n289 185
R35003 a_188130_n13996.n292 a_188130_n13996.n291 185
R35004 a_188130_n13996.n278 a_188130_n13996.n277 185
R35005 a_188130_n13996.t2 a_188130_n13996.n283 174.857
R35006 a_188130_n13996.n284 a_188130_n13996.n281 140.69
R35007 a_188130_n13996.n290 a_188130_n13996.n281 140.69
R35008 a_188130_n13996.n291 a_188130_n13996.n290 140.69
R35009 a_188130_n13996.n291 a_188130_n13996.n277 140.69
R35010 a_188130_n13996.n14 a_188130_n13996.n277 256.962
R35011 a_188130_n13996.n142 a_188130_n13996.t7 115.484
R35012 a_188130_n13996.n284 a_188130_n13996.t2 70.3453
R35013 a_188130_n13996.n408 a_188130_n13996.n40 51.6894
R35014 a_188130_n13996.n66 a_188130_n13996.n65 51.6891
R35015 a_188130_n13996.n389 a_188130_n13996.n388 51.6891
R35016 a_188130_n13996.n397 a_188130_n13996.n396 51.6891
R35017 a_188130_n13996.n405 a_188130_n13996.n404 51.6891
R35018 a_188130_n13996.n49 a_188130_n13996.n48 51.6891
R35019 a_188130_n13996.n65 a_188130_n13996.n64 29.8062
R35020 a_188130_n13996.n388 a_188130_n13996.n387 29.8062
R35021 a_188130_n13996.n396 a_188130_n13996.n395 29.8062
R35022 a_188130_n13996.n404 a_188130_n13996.n403 29.8062
R35023 a_188130_n13996.n48 a_188130_n13996.n47 29.8062
R35024 a_188130_n13996.n53 a_188130_n13996.n40 29.8061
R35025 a_188130_n13996.n143 a_188130_n13996.n141 29.3167
R35026 a_188130_n13996.n285 a_188130_n13996.n283 28.4333
R35027 a_188130_n13996.n328 a_188130_n13996.n327 26.8423
R35028 a_188130_n13996.n317 a_188130_n13996.n316 26.8423
R35029 a_188130_n13996.n306 a_188130_n13996.n305 26.8423
R35030 a_188130_n13996.n337 a_188130_n13996.n96 24.8476
R35031 a_188130_n13996.n335 a_188130_n13996.n94 24.8476
R35032 a_188130_n13996.n286 a_188130_n13996.n282 24.8476
R35033 a_188130_n13996.n260 a_188130_n13996.n114 24.8476
R35034 a_188130_n13996.n258 a_188130_n13996.n112 24.8476
R35035 a_188130_n13996.n167 a_188130_n13996.n131 24.8476
R35036 a_188130_n13996.n165 a_188130_n13996.n129 24.8476
R35037 a_188130_n13996.n365 a_188130_n13996.n78 24.8476
R35038 a_188130_n13996.n363 a_188130_n13996.n76 24.8476
R35039 a_188130_n13996.n144 a_188130_n13996.n140 24.8476
R35040 a_188130_n13996.n339 a_188130_n13996.n97 23.3417
R35041 a_188130_n13996.n333 a_188130_n13996.n93 23.3417
R35042 a_188130_n13996.n289 a_188130_n13996.n288 23.3417
R35043 a_188130_n13996.n262 a_188130_n13996.n115 23.3417
R35044 a_188130_n13996.n256 a_188130_n13996.n111 23.3417
R35045 a_188130_n13996.n169 a_188130_n13996.n132 23.3417
R35046 a_188130_n13996.n163 a_188130_n13996.n128 23.3417
R35047 a_188130_n13996.n367 a_188130_n13996.n79 23.3417
R35048 a_188130_n13996.n361 a_188130_n13996.n75 23.3417
R35049 a_188130_n13996.n148 a_188130_n13996.n147 23.3417
R35050 a_188130_n13996.n341 a_188130_n13996.n98 21.8358
R35051 a_188130_n13996.n332 a_188130_n13996.n92 21.8358
R35052 a_188130_n13996.n327 a_188130_n13996.n321 21.8358
R35053 a_188130_n13996.n316 a_188130_n13996.n310 21.8358
R35054 a_188130_n13996.n305 a_188130_n13996.n299 21.8358
R35055 a_188130_n13996.n292 a_188130_n13996.n280 21.8358
R35056 a_188130_n13996.n264 a_188130_n13996.n116 21.8358
R35057 a_188130_n13996.n255 a_188130_n13996.n110 21.8358
R35058 a_188130_n13996.n171 a_188130_n13996.n133 21.8358
R35059 a_188130_n13996.n162 a_188130_n13996.n127 21.8358
R35060 a_188130_n13996.n369 a_188130_n13996.n80 21.8358
R35061 a_188130_n13996.n74 a_188130_n13996.n69 21.8358
R35062 a_188130_n13996.n151 a_188130_n13996.n5 21.8358
R35063 a_188130_n13996.n64 a_188130_n13996.n60 20.3299
R35064 a_188130_n13996.n343 a_188130_n13996.n99 20.3299
R35065 a_188130_n13996.n100 a_188130_n13996.n91 20.3299
R35066 a_188130_n13996.n324 a_188130_n13996.n320 20.3299
R35067 a_188130_n13996.n313 a_188130_n13996.n309 20.3299
R35068 a_188130_n13996.n302 a_188130_n13996.n298 20.3299
R35069 a_188130_n13996.n293 a_188130_n13996.n278 20.3299
R35070 a_188130_n13996.n266 a_188130_n13996.n117 20.3299
R35071 a_188130_n13996.n253 a_188130_n13996.n109 20.3299
R35072 a_188130_n13996.n173 a_188130_n13996.n134 20.3299
R35073 a_188130_n13996.n135 a_188130_n13996.n126 20.3299
R35074 a_188130_n13996.n371 a_188130_n13996.n81 20.3299
R35075 a_188130_n13996.n380 a_188130_n13996.n379 20.3299
R35076 a_188130_n13996.n387 a_188130_n13996.n383 20.3299
R35077 a_188130_n13996.n395 a_188130_n13996.n391 20.3299
R35078 a_188130_n13996.n403 a_188130_n13996.n399 20.3299
R35079 a_188130_n13996.n47 a_188130_n13996.n43 20.3299
R35080 a_188130_n13996.n152 a_188130_n13996.n138 20.3299
R35081 a_188130_n13996.n53 a_188130_n13996.n41 20.3299
R35082 a_188130_n13996.n350 a_188130_n13996.n349 19.0887
R35083 a_188130_n13996.n105 a_188130_n13996.n89 19.0887
R35084 a_188130_n13996.n272 a_188130_n13996.n250 19.0887
R35085 a_188130_n13996.n275 a_188130_n13996.n274 19.0887
R35086 a_188130_n13996.n180 a_188130_n13996.n179 19.0887
R35087 a_188130_n13996.n124 a_188130_n13996.n19 19.0887
R35088 a_188130_n13996.n377 a_188130_n13996.n360 19.0887
R35089 a_188130_n13996.n355 a_188130_n13996.n71 19.0887
R35090 a_188130_n13996.n61 a_188130_n13996.n17 24.6305
R35091 a_188130_n13996.n347 a_188130_n13996.n346 18.824
R35092 a_188130_n13996.n102 a_188130_n13996.n90 18.824
R35093 a_188130_n13996.n322 a_188130_n13996.n8 24.4363
R35094 a_188130_n13996.n311 a_188130_n13996.n10 24.4363
R35095 a_188130_n13996.n300 a_188130_n13996.n12 24.4363
R35096 a_188130_n13996.n14 a_188130_n13996.n296 22.9459
R35097 a_188130_n13996.n268 a_188130_n13996.n118 18.824
R35098 a_188130_n13996.n251 a_188130_n13996.n108 18.824
R35099 a_188130_n13996.n177 a_188130_n13996.n176 18.824
R35100 a_188130_n13996.n158 a_188130_n13996.n125 18.824
R35101 a_188130_n13996.n373 a_188130_n13996.n82 18.824
R35102 a_188130_n13996.n73 a_188130_n13996.n70 18.824
R35103 a_188130_n13996.n384 a_188130_n13996.n26 24.6305
R35104 a_188130_n13996.n392 a_188130_n13996.n28 24.6305
R35105 a_188130_n13996.n400 a_188130_n13996.n30 24.6305
R35106 a_188130_n13996.n44 a_188130_n13996.n32 24.6305
R35107 a_188130_n13996.n34 a_188130_n13996.n155 23.6861
R35108 a_188130_n13996.n51 a_188130_n13996.n36 24.6305
R35109 a_188130_n13996.n17 a_188130_n13996.n16 9.772
R35110 a_188130_n13996.n349 a_188130_n13996.n88 17.3181
R35111 a_188130_n13996.n104 a_188130_n13996.n89 17.3181
R35112 a_188130_n13996.n8 a_188130_n13996.n7 9.72509
R35113 a_188130_n13996.n10 a_188130_n13996.n9 9.72509
R35114 a_188130_n13996.n12 a_188130_n13996.n11 9.72509
R35115 a_188130_n13996.n14 a_188130_n13996.n13 11.3106
R35116 a_188130_n13996.n272 a_188130_n13996.n271 17.3181
R35117 a_188130_n13996.n274 a_188130_n13996.n107 17.3181
R35118 a_188130_n13996.n179 a_188130_n13996.n123 17.3181
R35119 a_188130_n13996.n160 a_188130_n13996.n124 17.3181
R35120 a_188130_n13996.n377 a_188130_n13996.n376 17.3181
R35121 a_188130_n13996.n72 a_188130_n13996.n71 17.3181
R35122 a_188130_n13996.n26 a_188130_n13996.n25 9.772
R35123 a_188130_n13996.n28 a_188130_n13996.n27 9.772
R35124 a_188130_n13996.n30 a_188130_n13996.n29 9.772
R35125 a_188130_n13996.n32 a_188130_n13996.n31 9.772
R35126 a_188130_n13996.n34 a_188130_n13996.n33 10.7354
R35127 a_188130_n13996.n36 a_188130_n13996.n35 9.772
R35128 a_188130_n13996.n329 a_188130_n13996.n328 16.7813
R35129 a_188130_n13996.n318 a_188130_n13996.n317 16.7813
R35130 a_188130_n13996.n307 a_188130_n13996.n306 16.7813
R35131 a_188130_n13996.n337 a_188130_n13996.n95 13.2799
R35132 a_188130_n13996.n335 a_188130_n13996.n95 13.2799
R35133 a_188130_n13996.n260 a_188130_n13996.n113 13.2799
R35134 a_188130_n13996.n258 a_188130_n13996.n113 13.2799
R35135 a_188130_n13996.n167 a_188130_n13996.n130 13.2799
R35136 a_188130_n13996.n165 a_188130_n13996.n130 13.2799
R35137 a_188130_n13996.n365 a_188130_n13996.n77 13.2799
R35138 a_188130_n13996.n363 a_188130_n13996.n77 13.2799
R35139 a_188130_n13996.n64 a_188130_n13996.n63 9.3005
R35140 a_188130_n13996.n62 a_188130_n13996.n61 9.3005
R35141 a_188130_n13996.n327 a_188130_n13996.n326 9.3005
R35142 a_188130_n13996.n325 a_188130_n13996.n324 9.3005
R35143 a_188130_n13996.n323 a_188130_n13996.n322 9.3005
R35144 a_188130_n13996.n316 a_188130_n13996.n315 9.3005
R35145 a_188130_n13996.n314 a_188130_n13996.n313 9.3005
R35146 a_188130_n13996.n312 a_188130_n13996.n311 9.3005
R35147 a_188130_n13996.n305 a_188130_n13996.n304 9.3005
R35148 a_188130_n13996.n303 a_188130_n13996.n302 9.3005
R35149 a_188130_n13996.n301 a_188130_n13996.n300 9.3005
R35150 a_188130_n13996.n287 a_188130_n13996.n286 9.3005
R35151 a_188130_n13996.n280 a_188130_n13996.n279 9.3005
R35152 a_188130_n13996.n294 a_188130_n13996.n293 9.3005
R35153 a_188130_n13996.n296 a_188130_n13996.n295 9.3005
R35154 a_188130_n13996.n288 a_188130_n13996.n18 9.3005
R35155 a_188130_n13996.n381 a_188130_n13996.n380 9.3005
R35156 a_188130_n13996.n70 a_188130_n13996.n23 9.3005
R35157 a_188130_n13996.n74 a_188130_n13996.n0 9.3005
R35158 a_188130_n13996.n366 a_188130_n13996.n365 9.3005
R35159 a_188130_n13996.n368 a_188130_n13996.n367 9.3005
R35160 a_188130_n13996.n370 a_188130_n13996.n369 9.3005
R35161 a_188130_n13996.n372 a_188130_n13996.n371 9.3005
R35162 a_188130_n13996.n374 a_188130_n13996.n373 9.3005
R35163 a_188130_n13996.n376 a_188130_n13996.n375 9.3005
R35164 a_188130_n13996.n364 a_188130_n13996.n363 9.3005
R35165 a_188130_n13996.n362 a_188130_n13996.n361 9.3005
R35166 a_188130_n13996.n168 a_188130_n13996.n167 9.3005
R35167 a_188130_n13996.n170 a_188130_n13996.n169 9.3005
R35168 a_188130_n13996.n172 a_188130_n13996.n171 9.3005
R35169 a_188130_n13996.n174 a_188130_n13996.n173 9.3005
R35170 a_188130_n13996.n176 a_188130_n13996.n175 9.3005
R35171 a_188130_n13996.n123 a_188130_n13996.n122 9.3005
R35172 a_188130_n13996.n166 a_188130_n13996.n165 9.3005
R35173 a_188130_n13996.n164 a_188130_n13996.n163 9.3005
R35174 a_188130_n13996.n1 a_188130_n13996.n162 9.3005
R35175 a_188130_n13996.n136 a_188130_n13996.n135 9.3005
R35176 a_188130_n13996.n159 a_188130_n13996.n158 9.3005
R35177 a_188130_n13996.n20 a_188130_n13996.n160 9.3005
R35178 a_188130_n13996.n107 a_188130_n13996.n21 9.3005
R35179 a_188130_n13996.n254 a_188130_n13996.n253 9.3005
R35180 a_188130_n13996.n252 a_188130_n13996.n251 9.3005
R35181 a_188130_n13996.n3 a_188130_n13996.n255 9.3005
R35182 a_188130_n13996.n261 a_188130_n13996.n260 9.3005
R35183 a_188130_n13996.n263 a_188130_n13996.n262 9.3005
R35184 a_188130_n13996.n265 a_188130_n13996.n264 9.3005
R35185 a_188130_n13996.n267 a_188130_n13996.n266 9.3005
R35186 a_188130_n13996.n269 a_188130_n13996.n268 9.3005
R35187 a_188130_n13996.n271 a_188130_n13996.n270 9.3005
R35188 a_188130_n13996.n259 a_188130_n13996.n258 9.3005
R35189 a_188130_n13996.n257 a_188130_n13996.n256 9.3005
R35190 a_188130_n13996.n338 a_188130_n13996.n337 9.3005
R35191 a_188130_n13996.n340 a_188130_n13996.n339 9.3005
R35192 a_188130_n13996.n342 a_188130_n13996.n341 9.3005
R35193 a_188130_n13996.n344 a_188130_n13996.n343 9.3005
R35194 a_188130_n13996.n346 a_188130_n13996.n345 9.3005
R35195 a_188130_n13996.n88 a_188130_n13996.n87 9.3005
R35196 a_188130_n13996.n336 a_188130_n13996.n335 9.3005
R35197 a_188130_n13996.n334 a_188130_n13996.n333 9.3005
R35198 a_188130_n13996.n4 a_188130_n13996.n332 9.3005
R35199 a_188130_n13996.n101 a_188130_n13996.n100 9.3005
R35200 a_188130_n13996.n103 a_188130_n13996.n102 9.3005
R35201 a_188130_n13996.n22 a_188130_n13996.n104 9.3005
R35202 a_188130_n13996.n72 a_188130_n13996.n24 9.3005
R35203 a_188130_n13996.n387 a_188130_n13996.n386 9.3005
R35204 a_188130_n13996.n385 a_188130_n13996.n384 9.3005
R35205 a_188130_n13996.n395 a_188130_n13996.n394 9.3005
R35206 a_188130_n13996.n393 a_188130_n13996.n392 9.3005
R35207 a_188130_n13996.n403 a_188130_n13996.n402 9.3005
R35208 a_188130_n13996.n401 a_188130_n13996.n400 9.3005
R35209 a_188130_n13996.n47 a_188130_n13996.n46 9.3005
R35210 a_188130_n13996.n45 a_188130_n13996.n44 9.3005
R35211 a_188130_n13996.n145 a_188130_n13996.n144 9.3005
R35212 a_188130_n13996.n147 a_188130_n13996.n146 9.3005
R35213 a_188130_n13996.n153 a_188130_n13996.n152 9.3005
R35214 a_188130_n13996.n155 a_188130_n13996.n154 9.3005
R35215 a_188130_n13996.n6 a_188130_n13996.n5 9.3005
R35216 a_188130_n13996.n54 a_188130_n13996.n53 9.3005
R35217 a_188130_n13996.n52 a_188130_n13996.n51 9.3005
R35218 a_188130_n13996.n347 a_188130_n13996.n88 8.28285
R35219 a_188130_n13996.n104 a_188130_n13996.n90 8.28285
R35220 a_188130_n13996.n271 a_188130_n13996.n118 8.28285
R35221 a_188130_n13996.n108 a_188130_n13996.n107 8.28285
R35222 a_188130_n13996.n177 a_188130_n13996.n123 8.28285
R35223 a_188130_n13996.n160 a_188130_n13996.n125 8.28285
R35224 a_188130_n13996.n376 a_188130_n13996.n82 8.28285
R35225 a_188130_n13996.n73 a_188130_n13996.n72 8.28285
R35226 a_188130_n13996.n67 a_188130_n13996.n59 7.9105
R35227 a_188130_n13996.n37 a_188130_n13996.n319 7.9105
R35228 a_188130_n13996.n37 a_188130_n13996.n308 7.9105
R35229 a_188130_n13996.n15 a_188130_n13996.n297 7.9105
R35230 a_188130_n13996.n15 a_188130_n13996.n18 7.9105
R35231 a_188130_n13996.n15 a_188130_n13996.n13 7.9105
R35232 a_188130_n13996.n15 a_188130_n13996.n11 7.9105
R35233 a_188130_n13996.n37 a_188130_n13996.n9 7.9105
R35234 a_188130_n13996.n37 a_188130_n13996.n7 7.9105
R35235 a_188130_n13996.n382 a_188130_n13996.n24 7.9105
R35236 a_188130_n13996.n390 a_188130_n13996.n58 7.9105
R35237 a_188130_n13996.n398 a_188130_n13996.n57 7.9105
R35238 a_188130_n13996.n406 a_188130_n13996.n56 7.9105
R35239 a_188130_n13996.n50 a_188130_n13996.n42 7.9105
R35240 a_188130_n13996.n156 a_188130_n13996.n6 7.9105
R35241 a_188130_n13996.n156 a_188130_n13996.n33 7.9105
R35242 a_188130_n13996.n50 a_188130_n13996.n31 7.9105
R35243 a_188130_n13996.n406 a_188130_n13996.n29 7.9105
R35244 a_188130_n13996.n398 a_188130_n13996.n27 7.9105
R35245 a_188130_n13996.n390 a_188130_n13996.n25 7.9105
R35246 a_188130_n13996.n382 a_188130_n13996.n0 7.9105
R35247 a_188130_n13996.n1 a_188130_n13996.n161 7.9105
R35248 a_188130_n13996.n161 a_188130_n13996.n20 7.9105
R35249 a_188130_n13996.n67 a_188130_n13996.n16 7.9105
R35250 a_188130_n13996.n35 a_188130_n13996.n407 7.9105
R35251 a_188130_n13996.n407 a_188130_n13996.n55 7.9105
R35252 a_188130_n13996.n61 a_188130_n13996.n60 6.77697
R35253 a_188130_n13996.n346 a_188130_n13996.n99 6.77697
R35254 a_188130_n13996.n102 a_188130_n13996.n91 6.77697
R35255 a_188130_n13996.n322 a_188130_n13996.n320 6.77697
R35256 a_188130_n13996.n311 a_188130_n13996.n309 6.77697
R35257 a_188130_n13996.n300 a_188130_n13996.n298 6.77697
R35258 a_188130_n13996.n296 a_188130_n13996.n278 6.77697
R35259 a_188130_n13996.n268 a_188130_n13996.n117 6.77697
R35260 a_188130_n13996.n251 a_188130_n13996.n109 6.77697
R35261 a_188130_n13996.n176 a_188130_n13996.n134 6.77697
R35262 a_188130_n13996.n158 a_188130_n13996.n126 6.77697
R35263 a_188130_n13996.n373 a_188130_n13996.n81 6.77697
R35264 a_188130_n13996.n379 a_188130_n13996.n70 6.77697
R35265 a_188130_n13996.n384 a_188130_n13996.n383 6.77697
R35266 a_188130_n13996.n392 a_188130_n13996.n391 6.77697
R35267 a_188130_n13996.n400 a_188130_n13996.n399 6.77697
R35268 a_188130_n13996.n44 a_188130_n13996.n43 6.77697
R35269 a_188130_n13996.n155 a_188130_n13996.n138 6.77697
R35270 a_188130_n13996.n51 a_188130_n13996.n41 6.77697
R35271 a_188130_n13996.n66 a_188130_n13996.t9 5.7135
R35272 a_188130_n13996.n66 a_188130_n13996.t31 5.7135
R35273 a_188130_n13996.n348 a_188130_n13996.t25 5.7135
R35274 a_188130_n13996.n348 a_188130_n13996.t19 5.7135
R35275 a_188130_n13996.n273 a_188130_n13996.t43 5.7135
R35276 a_188130_n13996.n273 a_188130_n13996.t15 5.7135
R35277 a_188130_n13996.n178 a_188130_n13996.t13 5.7135
R35278 a_188130_n13996.n178 a_188130_n13996.t39 5.7135
R35279 a_188130_n13996.n378 a_188130_n13996.t35 5.7135
R35280 a_188130_n13996.n378 a_188130_n13996.t29 5.7135
R35281 a_188130_n13996.n389 a_188130_n13996.t41 5.7135
R35282 a_188130_n13996.n389 a_188130_n13996.t33 5.7135
R35283 a_188130_n13996.n397 a_188130_n13996.t17 5.7135
R35284 a_188130_n13996.n397 a_188130_n13996.t5 5.7135
R35285 a_188130_n13996.n405 a_188130_n13996.t37 5.7135
R35286 a_188130_n13996.n405 a_188130_n13996.t23 5.7135
R35287 a_188130_n13996.n49 a_188130_n13996.t27 5.7135
R35288 a_188130_n13996.n49 a_188130_n13996.t21 5.7135
R35289 a_188130_n13996.n408 a_188130_n13996.t11 5.7135
R35290 a_188130_n13996.t45 a_188130_n13996.n408 5.7135
R35291 a_188130_n13996.n287 a_188130_n13996.n283 5.33935
R35292 a_188130_n13996.n343 a_188130_n13996.n98 5.27109
R35293 a_188130_n13996.n100 a_188130_n13996.n92 5.27109
R35294 a_188130_n13996.n324 a_188130_n13996.n321 5.27109
R35295 a_188130_n13996.n313 a_188130_n13996.n310 5.27109
R35296 a_188130_n13996.n302 a_188130_n13996.n299 5.27109
R35297 a_188130_n13996.n293 a_188130_n13996.n292 5.27109
R35298 a_188130_n13996.n266 a_188130_n13996.n116 5.27109
R35299 a_188130_n13996.n253 a_188130_n13996.n110 5.27109
R35300 a_188130_n13996.n173 a_188130_n13996.n133 5.27109
R35301 a_188130_n13996.n135 a_188130_n13996.n127 5.27109
R35302 a_188130_n13996.n371 a_188130_n13996.n80 5.27109
R35303 a_188130_n13996.n380 a_188130_n13996.n69 5.27109
R35304 a_188130_n13996.n152 a_188130_n13996.n151 5.27109
R35305 a_188130_n13996.n3 a_188130_n13996.n2 4.59906
R35306 a_188130_n13996.n4 a_188130_n13996.n331 4.59906
R35307 a_188130_n13996.n15 a_188130_n13996.n276 4.5738
R35308 a_188130_n13996.n330 a_188130_n13996.n37 4.57256
R35309 a_188130_n13996.n145 a_188130_n13996.n141 4.51911
R35310 a_188130_n13996.n276 a_188130_n13996.n21 4.5005
R35311 a_188130_n13996.n330 a_188130_n13996.n22 4.5005
R35312 a_188130_n13996.n341 a_188130_n13996.n97 3.76521
R35313 a_188130_n13996.n332 a_188130_n13996.n93 3.76521
R35314 a_188130_n13996.n289 a_188130_n13996.n280 3.76521
R35315 a_188130_n13996.n264 a_188130_n13996.n115 3.76521
R35316 a_188130_n13996.n255 a_188130_n13996.n111 3.76521
R35317 a_188130_n13996.n171 a_188130_n13996.n132 3.76521
R35318 a_188130_n13996.n162 a_188130_n13996.n128 3.76521
R35319 a_188130_n13996.n369 a_188130_n13996.n79 3.76521
R35320 a_188130_n13996.n75 a_188130_n13996.n74 3.76521
R35321 a_188130_n13996.n148 a_188130_n13996.n5 3.76521
R35322 a_188130_n13996.n328 a_188130_n13996.n319 3.76174
R35323 a_188130_n13996.n317 a_188130_n13996.n308 3.76174
R35324 a_188130_n13996.n306 a_188130_n13996.n297 3.76174
R35325 a_188130_n13996.n329 a_188130_n13996.t48 3.4805
R35326 a_188130_n13996.n329 a_188130_n13996.t3 3.4805
R35327 a_188130_n13996.n318 a_188130_n13996.t46 3.4805
R35328 a_188130_n13996.n318 a_188130_n13996.t0 3.4805
R35329 a_188130_n13996.n307 a_188130_n13996.t1 3.4805
R35330 a_188130_n13996.n307 a_188130_n13996.t47 3.4805
R35331 a_188130_n13996.n55 a_188130_n13996.n40 3.43567
R35332 a_188130_n13996.n65 a_188130_n13996.n59 3.43565
R35333 a_188130_n13996.n388 a_188130_n13996.n58 3.43565
R35334 a_188130_n13996.n396 a_188130_n13996.n57 3.43565
R35335 a_188130_n13996.n404 a_188130_n13996.n56 3.43565
R35336 a_188130_n13996.n48 a_188130_n13996.n42 3.43565
R35337 a_188130_n13996.n339 a_188130_n13996.n96 2.25932
R35338 a_188130_n13996.n333 a_188130_n13996.n94 2.25932
R35339 a_188130_n13996.n288 a_188130_n13996.n282 2.25932
R35340 a_188130_n13996.n262 a_188130_n13996.n114 2.25932
R35341 a_188130_n13996.n256 a_188130_n13996.n112 2.25932
R35342 a_188130_n13996.n169 a_188130_n13996.n131 2.25932
R35343 a_188130_n13996.n163 a_188130_n13996.n129 2.25932
R35344 a_188130_n13996.n367 a_188130_n13996.n78 2.25932
R35345 a_188130_n13996.n361 a_188130_n13996.n76 2.25932
R35346 a_188130_n13996.n147 a_188130_n13996.n140 2.25932
R35347 a_188130_n13996.n157 a_188130_n13996.n2 1.65697
R35348 a_188130_n13996.n331 a_188130_n13996.n68 1.65697
R35349 a_188130_n13996.n214 a_188130_n13996.n213 1.62034
R35350 a_188130_n13996.n194 a_188130_n13996.n193 1.61786
R35351 a_188130_n13996.n213 a_188130_n13996.n212 1.22534
R35352 a_188130_n13996.n193 a_188130_n13996.n192 1.22286
R35353 a_188130_n13996.n286 a_188130_n13996.n285 0.753441
R35354 a_188130_n13996.n144 a_188130_n13996.n143 0.753441
R35355 a_188130_n13996.n231 a_188130_n13996.n184 0.3955
R35356 a_188130_n13996.n231 a_188130_n13996.n230 0.3955
R35357 a_188130_n13996.n230 a_188130_n13996.n84 0.3955
R35358 a_188130_n13996.n358 a_188130_n13996.n84 0.3955
R35359 a_188130_n13996.n197 a_188130_n13996.n196 0.3955
R35360 a_188130_n13996.n198 a_188130_n13996.n197 0.3955
R35361 a_188130_n13996.n198 a_188130_n13996.n188 0.3955
R35362 a_188130_n13996.n202 a_188130_n13996.n188 0.3955
R35363 a_188130_n13996.n203 a_188130_n13996.n202 0.3955
R35364 a_188130_n13996.n204 a_188130_n13996.n203 0.3955
R35365 a_188130_n13996.n204 a_188130_n13996.n185 0.3955
R35366 a_188130_n13996.n224 a_188130_n13996.n186 0.3955
R35367 a_188130_n13996.n224 a_188130_n13996.n223 0.3955
R35368 a_188130_n13996.n223 a_188130_n13996.n222 0.3955
R35369 a_188130_n13996.n222 a_188130_n13996.n208 0.3955
R35370 a_188130_n13996.n218 a_188130_n13996.n208 0.3955
R35371 a_188130_n13996.n218 a_188130_n13996.n217 0.3955
R35372 a_188130_n13996.n217 a_188130_n13996.n216 0.3955
R35373 a_188130_n13996.n243 a_188130_n13996.n242 0.3955
R35374 a_188130_n13996.n242 a_188130_n13996.n241 0.3955
R35375 a_188130_n13996.n241 a_188130_n13996.n182 0.3955
R35376 a_188130_n13996.n237 a_188130_n13996.n182 0.3955
R35377 a_188130_n13996.n237 a_188130_n13996.n236 0.3955
R35378 a_188130_n13996.n248 a_188130_n13996.n120 0.3955
R35379 a_188130_n13996.n247 a_188130_n13996.n246 0.3955
R35380 a_188130_n13996.n195 a_188130_n13996.n194 0.3955
R35381 a_188130_n13996.n195 a_188130_n13996.n189 0.3955
R35382 a_188130_n13996.n199 a_188130_n13996.n189 0.3955
R35383 a_188130_n13996.n200 a_188130_n13996.n199 0.3955
R35384 a_188130_n13996.n201 a_188130_n13996.n200 0.3955
R35385 a_188130_n13996.n201 a_188130_n13996.n187 0.3955
R35386 a_188130_n13996.n205 a_188130_n13996.n187 0.3955
R35387 a_188130_n13996.n206 a_188130_n13996.n205 0.3955
R35388 a_188130_n13996.n227 a_188130_n13996.n206 0.3955
R35389 a_188130_n13996.n227 a_188130_n13996.n226 0.3955
R35390 a_188130_n13996.n226 a_188130_n13996.n225 0.3955
R35391 a_188130_n13996.n225 a_188130_n13996.n207 0.3955
R35392 a_188130_n13996.n221 a_188130_n13996.n207 0.3955
R35393 a_188130_n13996.n221 a_188130_n13996.n220 0.3955
R35394 a_188130_n13996.n220 a_188130_n13996.n219 0.3955
R35395 a_188130_n13996.n219 a_188130_n13996.n209 0.3955
R35396 a_188130_n13996.n215 a_188130_n13996.n209 0.3955
R35397 a_188130_n13996.n215 a_188130_n13996.n214 0.3955
R35398 a_188130_n13996.n211 a_188130_n13996.n210 0.3955
R35399 a_188130_n13996.n352 a_188130_n13996.n83 0.3955
R35400 a_188130_n13996.n354 a_188130_n13996.n353 0.3955
R35401 a_188130_n13996.n244 a_188130_n13996.n121 0.3955
R35402 a_188130_n13996.n240 a_188130_n13996.n121 0.3955
R35403 a_188130_n13996.n240 a_188130_n13996.n239 0.3955
R35404 a_188130_n13996.n239 a_188130_n13996.n238 0.3955
R35405 a_188130_n13996.n238 a_188130_n13996.n183 0.3955
R35406 a_188130_n13996.n234 a_188130_n13996.n183 0.3955
R35407 a_188130_n13996.n234 a_188130_n13996.n233 0.3955
R35408 a_188130_n13996.n233 a_188130_n13996.n232 0.3955
R35409 a_188130_n13996.n232 a_188130_n13996.n229 0.3955
R35410 a_188130_n13996.n229 a_188130_n13996.n85 0.3955
R35411 a_188130_n13996.n357 a_188130_n13996.n85 0.3955
R35412 a_188130_n13996.n216 a_188130_n13996.n212 0.2555
R35413 a_188130_n13996.n39 a_188130_n13996.n38 0.2555
R35414 a_188130_n13996.n196 a_188130_n13996.n192 0.2505
R35415 a_188130_n13996.n295 a_188130_n13996.n13 0.231176
R35416 a_188130_n13996.n301 a_188130_n13996.n11 0.231176
R35417 a_188130_n13996.n312 a_188130_n13996.n9 0.231176
R35418 a_188130_n13996.n323 a_188130_n13996.n7 0.231176
R35419 a_188130_n13996.n52 a_188130_n13996.n35 0.225742
R35420 a_188130_n13996.n154 a_188130_n13996.n33 0.225742
R35421 a_188130_n13996.n45 a_188130_n13996.n31 0.225742
R35422 a_188130_n13996.n401 a_188130_n13996.n29 0.225742
R35423 a_188130_n13996.n393 a_188130_n13996.n27 0.225742
R35424 a_188130_n13996.n385 a_188130_n13996.n25 0.225742
R35425 a_188130_n13996.n62 a_188130_n13996.n16 0.225742
R35426 a_188130_n13996.n360 a_188130_n13996.n359 0.204667
R35427 a_188130_n13996.n181 a_188130_n13996.n180 0.204667
R35428 a_188130_n13996.n351 a_188130_n13996.n350 0.204667
R35429 a_188130_n13996.n249 a_188130_n13996.n248 0.2005
R35430 a_188130_n13996.n245 a_188130_n13996.n19 0.2005
R35431 a_188130_n13996.n275 a_188130_n13996.n106 0.2005
R35432 a_188130_n13996.n105 a_188130_n13996.n86 0.2005
R35433 a_188130_n13996.n356 a_188130_n13996.n355 0.2005
R35434 a_188130_n13996.n63 a_188130_n13996.n62 0.196152
R35435 a_188130_n13996.n326 a_188130_n13996.n325 0.196152
R35436 a_188130_n13996.n325 a_188130_n13996.n323 0.196152
R35437 a_188130_n13996.n315 a_188130_n13996.n314 0.196152
R35438 a_188130_n13996.n314 a_188130_n13996.n312 0.196152
R35439 a_188130_n13996.n304 a_188130_n13996.n303 0.196152
R35440 a_188130_n13996.n303 a_188130_n13996.n301 0.196152
R35441 a_188130_n13996.n294 a_188130_n13996.n279 0.196152
R35442 a_188130_n13996.n295 a_188130_n13996.n294 0.196152
R35443 a_188130_n13996.n386 a_188130_n13996.n385 0.196152
R35444 a_188130_n13996.n394 a_188130_n13996.n393 0.196152
R35445 a_188130_n13996.n402 a_188130_n13996.n401 0.196152
R35446 a_188130_n13996.n46 a_188130_n13996.n45 0.196152
R35447 a_188130_n13996.n146 a_188130_n13996.n145 0.196152
R35448 a_188130_n13996.n154 a_188130_n13996.n153 0.196152
R35449 a_188130_n13996.n54 a_188130_n13996.n52 0.196152
R35450 a_188130_n13996.n249 a_188130_n13996.n119 0.1955
R35451 a_188130_n13996.n146 a_188130_n13996.n6 0.194824
R35452 a_188130_n13996.n191 a_188130_n13996.n119 0.193
R35453 a_188130_n13996.n212 a_188130_n13996.n39 0.191241
R35454 a_188130_n13996.n235 a_188130_n13996.n228 0.190315
R35455 a_188130_n13996.n18 a_188130_n13996.n287 0.186853
R35456 a_188130_n13996.n192 a_188130_n13996.n191 0.178741
R35457 a_188130_n13996.n250 a_188130_n13996.n249 0.152583
R35458 a_188130_n13996.n381 a_188130_n13996.n23 0.1505
R35459 a_188130_n13996.n375 a_188130_n13996.n360 0.1505
R35460 a_188130_n13996.n375 a_188130_n13996.n374 0.1505
R35461 a_188130_n13996.n374 a_188130_n13996.n372 0.1505
R35462 a_188130_n13996.n372 a_188130_n13996.n370 0.1505
R35463 a_188130_n13996.n370 a_188130_n13996.n368 0.1505
R35464 a_188130_n13996.n368 a_188130_n13996.n366 0.1505
R35465 a_188130_n13996.n366 a_188130_n13996.n364 0.1505
R35466 a_188130_n13996.n364 a_188130_n13996.n362 0.1505
R35467 a_188130_n13996.n180 a_188130_n13996.n122 0.1505
R35468 a_188130_n13996.n175 a_188130_n13996.n122 0.1505
R35469 a_188130_n13996.n175 a_188130_n13996.n174 0.1505
R35470 a_188130_n13996.n174 a_188130_n13996.n172 0.1505
R35471 a_188130_n13996.n172 a_188130_n13996.n170 0.1505
R35472 a_188130_n13996.n170 a_188130_n13996.n168 0.1505
R35473 a_188130_n13996.n168 a_188130_n13996.n166 0.1505
R35474 a_188130_n13996.n166 a_188130_n13996.n164 0.1505
R35475 a_188130_n13996.n159 a_188130_n13996.n136 0.1505
R35476 a_188130_n13996.n254 a_188130_n13996.n252 0.1505
R35477 a_188130_n13996.n270 a_188130_n13996.n250 0.1505
R35478 a_188130_n13996.n270 a_188130_n13996.n269 0.1505
R35479 a_188130_n13996.n269 a_188130_n13996.n267 0.1505
R35480 a_188130_n13996.n267 a_188130_n13996.n265 0.1505
R35481 a_188130_n13996.n265 a_188130_n13996.n263 0.1505
R35482 a_188130_n13996.n263 a_188130_n13996.n261 0.1505
R35483 a_188130_n13996.n261 a_188130_n13996.n259 0.1505
R35484 a_188130_n13996.n259 a_188130_n13996.n257 0.1505
R35485 a_188130_n13996.n350 a_188130_n13996.n87 0.1505
R35486 a_188130_n13996.n345 a_188130_n13996.n87 0.1505
R35487 a_188130_n13996.n345 a_188130_n13996.n344 0.1505
R35488 a_188130_n13996.n344 a_188130_n13996.n342 0.1505
R35489 a_188130_n13996.n342 a_188130_n13996.n340 0.1505
R35490 a_188130_n13996.n340 a_188130_n13996.n338 0.1505
R35491 a_188130_n13996.n338 a_188130_n13996.n336 0.1505
R35492 a_188130_n13996.n336 a_188130_n13996.n334 0.1505
R35493 a_188130_n13996.n103 a_188130_n13996.n101 0.1505
R35494 a_188130_n13996.n362 a_188130_n13996.n0 0.149806
R35495 a_188130_n13996.n164 a_188130_n13996.n1 0.149806
R35496 a_188130_n13996.n257 a_188130_n13996.n3 0.149806
R35497 a_188130_n13996.n334 a_188130_n13996.n4 0.149806
R35498 a_188130_n13996.n24 a_188130_n13996.n23 0.145639
R35499 a_188130_n13996.n20 a_188130_n13996.n159 0.145639
R35500 a_188130_n13996.n252 a_188130_n13996.n21 0.145639
R35501 a_188130_n13996.n22 a_188130_n13996.n103 0.145639
R35502 a_188130_n13996.n181 a_188130_n13996.n120 0.1305
R35503 a_188130_n13996.n246 a_188130_n13996.n245 0.1305
R35504 a_188130_n13996.n359 a_188130_n13996.n83 0.1305
R35505 a_188130_n13996.n356 a_188130_n13996.n354 0.1305
R35506 a_188130_n13996.n247 a_188130_n13996.n106 0.1255
R35507 a_188130_n13996.n352 a_188130_n13996.n351 0.1255
R35508 a_188130_n13996.n353 a_188130_n13996.n86 0.1255
R35509 a_188130_n13996.n190 a_188130_n13996.n106 0.1205
R35510 a_188130_n13996.n210 a_188130_n13996.n86 0.1205
R35511 a_188130_n13996.n351 a_188130_n13996.n38 0.1205
R35512 a_188130_n13996.n37 a_188130_n13996.n15 0.118
R35513 a_188130_n13996.n359 a_188130_n13996.n358 0.1155
R35514 a_188130_n13996.n243 a_188130_n13996.n181 0.1155
R35515 a_188130_n13996.n245 a_188130_n13996.n244 0.1155
R35516 a_188130_n13996.n357 a_188130_n13996.n356 0.1155
R35517 a_188130_n13996.n279 a_188130_n13996.n18 0.112457
R35518 a_188130_n13996.n355 a_188130_n13996.n24 0.10675
R35519 a_188130_n13996.n22 a_188130_n13996.n105 0.10675
R35520 a_188130_n13996.n21 a_188130_n13996.n275 0.10675
R35521 a_188130_n13996.n20 a_188130_n13996.n19 0.10675
R35522 a_188130_n13996.n153 a_188130_n13996.n6 0.104486
R35523 a_188130_n13996.n4 a_188130_n13996.n101 0.102583
R35524 a_188130_n13996.n3 a_188130_n13996.n254 0.102583
R35525 a_188130_n13996.n1 a_188130_n13996.n136 0.102583
R35526 a_188130_n13996.n0 a_188130_n13996.n381 0.102583
R35527 a_188130_n13996.n276 a_188130_n13996.n2 0.0990583
R35528 a_188130_n13996.n331 a_188130_n13996.n330 0.0990583
R35529 a_188130_n13996.n326 a_188130_n13996.n319 0.0735676
R35530 a_188130_n13996.n315 a_188130_n13996.n308 0.0735676
R35531 a_188130_n13996.n304 a_188130_n13996.n297 0.0735676
R35532 a_188130_n13996.n228 a_188130_n13996.n185 0.0605
R35533 a_188130_n13996.n236 a_188130_n13996.n235 0.0605
R35534 a_188130_n13996.n63 a_188130_n13996.n59 0.0572633
R35535 a_188130_n13996.n386 a_188130_n13996.n58 0.0572633
R35536 a_188130_n13996.n394 a_188130_n13996.n57 0.0572633
R35537 a_188130_n13996.n402 a_188130_n13996.n56 0.0572633
R35538 a_188130_n13996.n46 a_188130_n13996.n42 0.0572633
R35539 a_188130_n13996.n55 a_188130_n13996.n54 0.0572633
R35540 a_188130_n13996.n235 a_188130_n13996.n184 0.0555
R35541 a_188130_n13996.n228 a_188130_n13996.n186 0.0555
R35542 a_188130_n13996.n157 a_188130_n13996.n156 0.0506333
R35543 a_188130_n13996.n161 a_188130_n13996.n50 0.0506333
R35544 a_188130_n13996.n407 a_188130_n13996.n406 0.0506333
R35545 a_188130_n13996.n406 a_188130_n13996.n398 0.0506333
R35546 a_188130_n13996.n390 a_188130_n13996.n382 0.0506333
R35547 a_188130_n13996.n68 a_188130_n13996.n67 0.0506333
R35548 a_188130_n13996.n161 a_188130_n13996.n157 0.0490667
R35549 a_188130_n13996.n407 a_188130_n13996.n50 0.0490667
R35550 a_188130_n13996.n398 a_188130_n13996.n390 0.0490667
R35551 a_188130_n13996.n382 a_188130_n13996.n68 0.0490667
R35552 CLK.n22 CLK.n21 280.079
R35553 CLK.n20 CLK.t2 231.907
R35554 CLK.n21 CLK.t14 231.361
R35555 CLK.n1 CLK.t16 212.081
R35556 CLK.n0 CLK.t9 212.081
R35557 CLK.n6 CLK.t6 212.081
R35558 CLK.n7 CLK.t1 212.081
R35559 CLK.n11 CLK.t5 212.081
R35560 CLK.n14 CLK.t18 212.081
R35561 CLK.n16 CLK.t8 212.081
R35562 CLK.n15 CLK.t3 212.081
R35563 CLK.n1 CLK 182.786
R35564 CLK.n20 CLK.t7 170.308
R35565 CLK.n18 CLK.n17 153.28
R35566 CLK.n3 CLK.n2 152
R35567 CLK.n5 CLK.n4 152
R35568 CLK.n9 CLK.n8 152
R35569 CLK.n13 CLK.n12 152
R35570 CLK.n1 CLK.t11 139.78
R35571 CLK.n0 CLK.t4 139.78
R35572 CLK.n6 CLK.t17 139.78
R35573 CLK.n7 CLK.t12 139.78
R35574 CLK.n11 CLK.t15 139.78
R35575 CLK.n14 CLK.t10 139.78
R35576 CLK.n16 CLK.t0 139.78
R35577 CLK.n15 CLK.t13 139.78
R35578 CLK.n16 CLK.n15 61.346
R35579 CLK.n21 CLK.n20 54.0627
R35580 CLK.n2 CLK.n1 30.6732
R35581 CLK.n2 CLK.n0 30.6732
R35582 CLK.n5 CLK.n0 30.6732
R35583 CLK.n6 CLK.n5 30.6732
R35584 CLK.n8 CLK.n6 30.6732
R35585 CLK.n8 CLK.n7 30.6732
R35586 CLK.n13 CLK.n11 30.6732
R35587 CLK.n14 CLK.n13 30.6732
R35588 CLK.n17 CLK.n14 30.6732
R35589 CLK.n17 CLK.n16 30.6732
R35590 CLK.n3 CLK 18.4325
R35591 CLK.n25 CLK.n24 17.2105
R35592 CLK.n4 CLK 16.3845
R35593 CLK.n19 CLK.n10 14.9687
R35594 CLK.n12 CLK 14.8485
R35595 CLK.n19 CLK.n18 14.0312
R35596 CLK CLK.n22 12.0005
R35597 CLK.n9 CLK 9.2165
R35598 CLK.n12 CLK 8.7045
R35599 CLK.n10 CLK.n9 8.4485
R35600 CLK.n4 CLK 7.1685
R35601 CLK.n22 CLK 6.13383
R35602 CLK.n24 CLK.n23 5.90819
R35603 CLK.n10 CLK 5.8885
R35604 CLK.n24 CLK 5.66204
R35605 CLK.n23 CLK 5.6005
R35606 CLK.n18 CLK 5.3765
R35607 CLK.n23 CLK 5.16973
R35608 CLK CLK.n3 5.1205
R35609 CLK.n25 CLK.n19 4.01523
R35610 CLK CLK.n25 0.2731
R35611 a_188937_n26928.n121 a_188937_n26928.n39 194.291
R35612 a_188937_n26928.n121 a_188937_n26928.n110 585
R35613 a_188937_n26928.n121 a_188937_n26928.n109 585
R35614 a_188937_n26928.n121 a_188937_n26928.n108 585
R35615 a_188937_n26928.n121 a_188937_n26928.n106 585
R35616 a_188937_n26928.n121 a_188937_n26928.n105 585
R35617 a_188937_n26928.n121 a_188937_n26928.n104 585
R35618 a_188937_n26928.n121 a_188937_n26928.n103 585
R35619 a_188937_n26928.n121 a_188937_n26928.n102 585
R35620 a_188937_n26928.n121 a_188937_n26928.n49 585
R35621 a_188937_n26928.n93 a_188937_n26928.n38 194.291
R35622 a_188937_n26928.n93 a_188937_n26928.n84 585
R35623 a_188937_n26928.n93 a_188937_n26928.n83 585
R35624 a_188937_n26928.n93 a_188937_n26928.n82 585
R35625 a_188937_n26928.n93 a_188937_n26928.n80 585
R35626 a_188937_n26928.n93 a_188937_n26928.n79 585
R35627 a_188937_n26928.n93 a_188937_n26928.n78 585
R35628 a_188937_n26928.n93 a_188937_n26928.n77 585
R35629 a_188937_n26928.n93 a_188937_n26928.n76 585
R35630 a_188937_n26928.n94 a_188937_n26928.n93 585
R35631 a_188937_n26928.n157 a_188937_n26928.n41 194.291
R35632 a_188937_n26928.n157 a_188937_n26928.n63 585
R35633 a_188937_n26928.n157 a_188937_n26928.n62 585
R35634 a_188937_n26928.n157 a_188937_n26928.n64 585
R35635 a_188937_n26928.n157 a_188937_n26928.n60 585
R35636 a_188937_n26928.n157 a_188937_n26928.n65 585
R35637 a_188937_n26928.n157 a_188937_n26928.n59 585
R35638 a_188937_n26928.n157 a_188937_n26928.n66 585
R35639 a_188937_n26928.n157 a_188937_n26928.n50 291.375
R35640 a_188937_n26928.t7 a_188937_n26928.n10 308.31
R35641 a_188937_n26928.n149 a_188937_n26928.t7 308.31
R35642 a_188937_n26928.t5 a_188937_n26928.n156 308.31
R35643 a_188937_n26928.n10 a_188937_n26928.t5 308.31
R35644 a_188937_n26928.n121 a_188937_n26928.n107 286.238
R35645 a_188937_n26928.n93 a_188937_n26928.n81 286.238
R35646 a_188937_n26928.n157 a_188937_n26928.n61 286.238
R35647 a_188937_n26928.n56 a_188937_n26928.n55 6.98494
R35648 a_188937_n26928.n58 a_188937_n26928.n57 6.98494
R35649 a_188937_n26928.t13 a_188937_n26928.n6 209.939
R35650 a_188937_n26928.n54 a_188937_n26928.t22 104.094
R35651 a_188937_n26928.n52 a_188937_n26928.t23 104.094
R35652 a_188937_n26928.n8 a_188937_n26928.t11 209.938
R35653 a_188937_n26928.t19 a_188937_n26928.n2 209.93
R35654 a_188937_n26928.n12 a_188937_n26928.t19 209.93
R35655 a_188937_n26928.t9 a_188937_n26928.n3 209.93
R35656 a_188937_n26928.n4 a_188937_n26928.t9 209.93
R35657 a_188937_n26928.n122 a_188937_n26928.t13 209.93
R35658 a_188937_n26928.t27 a_188937_n26928.n95 209.93
R35659 a_188937_n26928.n96 a_188937_n26928.t27 209.93
R35660 a_188937_n26928.n98 a_188937_n26928.t26 209.93
R35661 a_188937_n26928.t26 a_188937_n26928.n97 209.93
R35662 a_188937_n26928.t11 a_188937_n26928.n1 209.93
R35663 a_188937_n26928.n141 a_188937_n26928.t15 209.93
R35664 a_188937_n26928.t15 a_188937_n26928.n0 209.93
R35665 a_188937_n26928.t17 a_188937_n26928.n142 209.93
R35666 a_188937_n26928.n14 a_188937_n26928.t17 209.93
R35667 a_188937_n26928.n99 a_188937_n26928.t25 209.93
R35668 a_188937_n26928.t25 a_188937_n26928.n13 209.93
R35669 a_188937_n26928.t24 a_188937_n26928.n100 209.93
R35670 a_188937_n26928.n101 a_188937_n26928.t24 209.93
R35671 a_188937_n26928.n148 a_188937_n26928.n48 92.3135
R35672 a_188937_n26928.n148 a_188937_n26928.n144 185
R35673 a_188937_n26928.n148 a_188937_n26928.n20 92.3135
R35674 a_188937_n26928.n155 a_188937_n26928.n45 92.3135
R35675 a_188937_n26928.n155 a_188937_n26928.n151 185
R35676 a_188937_n26928.n155 a_188937_n26928.n17 92.3135
R35677 a_188937_n26928.n139 a_188937_n26928.n138 185
R35678 a_188937_n26928.n135 a_188937_n26928.n134 185
R35679 a_188937_n26928.n129 a_188937_n26928.n128 185
R35680 a_188937_n26928.n125 a_188937_n26928.n124 185
R35681 a_188937_n26928.n136 a_188937_n26928.t2 174.857
R35682 a_188937_n26928.n126 a_188937_n26928.t4 174.857
R35683 a_188937_n26928.n56 a_188937_n26928.n139 244.714
R35684 a_188937_n26928.n139 a_188937_n26928.n134 140.69
R35685 a_188937_n26928.n58 a_188937_n26928.n129 244.714
R35686 a_188937_n26928.n129 a_188937_n26928.n124 140.69
R35687 a_188937_n26928.n148 a_188937_n26928.n143 86.5152
R35688 a_188937_n26928.n155 a_188937_n26928.n150 86.5152
R35689 a_188937_n26928.t2 a_188937_n26928.n134 70.3453
R35690 a_188937_n26928.t4 a_188937_n26928.n124 70.3453
R35691 a_188937_n26928.n136 a_188937_n26928.n135 28.4333
R35692 a_188937_n26928.n126 a_188937_n26928.n125 28.4333
R35693 a_188937_n26928.n146 a_188937_n26928.n144 25.6005
R35694 a_188937_n26928.n153 a_188937_n26928.n151 25.6005
R35695 a_188937_n26928.n117 a_188937_n26928.n108 24.8476
R35696 a_188937_n26928.n116 a_188937_n26928.n106 24.8476
R35697 a_188937_n26928.n90 a_188937_n26928.n82 24.8476
R35698 a_188937_n26928.n89 a_188937_n26928.n80 24.8476
R35699 a_188937_n26928.n138 a_188937_n26928.n137 24.8476
R35700 a_188937_n26928.n128 a_188937_n26928.n127 24.8476
R35701 a_188937_n26928.n72 a_188937_n26928.n64 24.8476
R35702 a_188937_n26928.n71 a_188937_n26928.n60 24.8476
R35703 a_188937_n26928.n145 a_188937_n26928.n20 27.7565
R35704 a_188937_n26928.n152 a_188937_n26928.n17 27.7565
R35705 a_188937_n26928.n118 a_188937_n26928.n109 23.3417
R35706 a_188937_n26928.n115 a_188937_n26928.n105 23.3417
R35707 a_188937_n26928.n91 a_188937_n26928.n83 23.3417
R35708 a_188937_n26928.n88 a_188937_n26928.n79 23.3417
R35709 a_188937_n26928.n73 a_188937_n26928.n62 23.3417
R35710 a_188937_n26928.n70 a_188937_n26928.n65 23.3417
R35711 a_188937_n26928.n48 a_188937_n26928.n47 6.60954
R35712 a_188937_n26928.n20 a_188937_n26928.n18 6.60954
R35713 a_188937_n26928.n45 a_188937_n26928.n44 6.60954
R35714 a_188937_n26928.n17 a_188937_n26928.n15 6.60954
R35715 a_188937_n26928.n9 a_188937_n26928.n132 22.3909
R35716 a_188937_n26928.n9 a_188937_n26928.n131 22.3909
R35717 a_188937_n26928.n119 a_188937_n26928.n110 21.8358
R35718 a_188937_n26928.n114 a_188937_n26928.n104 21.8358
R35719 a_188937_n26928.n92 a_188937_n26928.n84 21.8358
R35720 a_188937_n26928.n87 a_188937_n26928.n78 21.8358
R35721 a_188937_n26928.n74 a_188937_n26928.n63 21.8358
R35722 a_188937_n26928.n69 a_188937_n26928.n59 21.8358
R35723 a_188937_n26928.n113 a_188937_n26928.n103 20.3299
R35724 a_188937_n26928.n86 a_188937_n26928.n77 20.3299
R35725 a_188937_n26928.n68 a_188937_n26928.n66 20.3299
R35726 a_188937_n26928.n3 a_188937_n26928.n49 19.0887
R35727 a_188937_n26928.n1 a_188937_n26928.n94 19.0887
R35728 a_188937_n26928.n39 a_188937_n26928.n5 6.07169
R35729 a_188937_n26928.n112 a_188937_n26928.n102 18.824
R35730 a_188937_n26928.n7 a_188937_n26928.n38 6.07169
R35731 a_188937_n26928.n85 a_188937_n26928.n76 18.824
R35732 a_188937_n26928.n11 a_188937_n26928.n41 6.07169
R35733 a_188937_n26928.n67 a_188937_n26928.n50 24.6333
R35734 a_188937_n26928.n111 a_188937_n26928.n49 17.3181
R35735 a_188937_n26928.n94 a_188937_n26928.n75 17.3181
R35736 a_188937_n26928.n50 a_188937_n26928.n2 9.76605
R35737 a_188937_n26928.n145 a_188937_n26928.n143 13.4786
R35738 a_188937_n26928.n152 a_188937_n26928.n150 13.4786
R35739 a_188937_n26928.n117 a_188937_n26928.n107 13.2799
R35740 a_188937_n26928.n116 a_188937_n26928.n107 13.2799
R35741 a_188937_n26928.n90 a_188937_n26928.n81 13.2799
R35742 a_188937_n26928.n89 a_188937_n26928.n81 13.2799
R35743 a_188937_n26928.n72 a_188937_n26928.n61 13.2799
R35744 a_188937_n26928.n71 a_188937_n26928.n61 13.2799
R35745 a_188937_n26928.n146 a_188937_n26928.n143 11.9727
R35746 a_188937_n26928.n153 a_188937_n26928.n150 11.9727
R35747 a_188937_n26928.n2 a_188937_n26928.n10 9.61161
R35748 a_188937_n26928.n8 a_188937_n26928.n51 9.47511
R35749 a_188937_n26928.n6 a_188937_n26928.n53 9.47106
R35750 a_188937_n26928.n13 a_188937_n26928.n12 9.3755
R35751 a_188937_n26928.n43 a_188937_n26928.n154 9.3005
R35752 a_188937_n26928.n16 a_188937_n26928.n153 9.3005
R35753 a_188937_n26928.n16 a_188937_n26928.n152 9.3005
R35754 a_188937_n26928.n46 a_188937_n26928.n147 9.3005
R35755 a_188937_n26928.n19 a_188937_n26928.n146 9.3005
R35756 a_188937_n26928.n19 a_188937_n26928.n145 9.3005
R35757 a_188937_n26928.n137 a_188937_n26928.n21 9.3005
R35758 a_188937_n26928.n133 a_188937_n26928.n21 9.3005
R35759 a_188937_n26928.n127 a_188937_n26928.n22 9.3005
R35760 a_188937_n26928.n123 a_188937_n26928.n22 9.3005
R35761 a_188937_n26928.n75 a_188937_n26928.n27 9.3005
R35762 a_188937_n26928.n23 a_188937_n26928.n90 9.3005
R35763 a_188937_n26928.n23 a_188937_n26928.n91 9.3005
R35764 a_188937_n26928.n24 a_188937_n26928.n92 9.3005
R35765 a_188937_n26928.n24 a_188937_n26928.n37 9.3005
R35766 a_188937_n26928.n25 a_188937_n26928.n89 9.3005
R35767 a_188937_n26928.n25 a_188937_n26928.n88 9.3005
R35768 a_188937_n26928.n26 a_188937_n26928.n87 9.3005
R35769 a_188937_n26928.n26 a_188937_n26928.n86 9.3005
R35770 a_188937_n26928.n27 a_188937_n26928.n85 9.3005
R35771 a_188937_n26928.n28 a_188937_n26928.n117 9.3005
R35772 a_188937_n26928.n28 a_188937_n26928.n118 9.3005
R35773 a_188937_n26928.n29 a_188937_n26928.n119 9.3005
R35774 a_188937_n26928.n29 a_188937_n26928.n120 9.3005
R35775 a_188937_n26928.n30 a_188937_n26928.n116 9.3005
R35776 a_188937_n26928.n30 a_188937_n26928.n115 9.3005
R35777 a_188937_n26928.n31 a_188937_n26928.n114 9.3005
R35778 a_188937_n26928.n31 a_188937_n26928.n113 9.3005
R35779 a_188937_n26928.n32 a_188937_n26928.n112 9.3005
R35780 a_188937_n26928.n32 a_188937_n26928.n111 9.3005
R35781 a_188937_n26928.n33 a_188937_n26928.n72 9.3005
R35782 a_188937_n26928.n34 a_188937_n26928.n73 9.3005
R35783 a_188937_n26928.n34 a_188937_n26928.n74 9.3005
R35784 a_188937_n26928.n42 a_188937_n26928.n40 9.3005
R35785 a_188937_n26928.n33 a_188937_n26928.n71 9.3005
R35786 a_188937_n26928.n35 a_188937_n26928.n70 9.3005
R35787 a_188937_n26928.n35 a_188937_n26928.n69 9.3005
R35788 a_188937_n26928.n36 a_188937_n26928.n68 9.3005
R35789 a_188937_n26928.n36 a_188937_n26928.n67 9.3005
R35790 a_188937_n26928.n111 a_188937_n26928.n102 8.28285
R35791 a_188937_n26928.n76 a_188937_n26928.n75 8.28285
R35792 a_188937_n26928.n1 a_188937_n26928.n140 7.04926
R35793 a_188937_n26928.n130 a_188937_n26928.n122 6.96926
R35794 a_188937_n26928.n148 a_188937_n26928.t8 6.9605
R35795 a_188937_n26928.n155 a_188937_n26928.t6 6.9605
R35796 a_188937_n26928.n39 a_188937_n26928.n120 28.1963
R35797 a_188937_n26928.n112 a_188937_n26928.n103 6.77697
R35798 a_188937_n26928.n38 a_188937_n26928.n37 28.1963
R35799 a_188937_n26928.n85 a_188937_n26928.n77 6.77697
R35800 a_188937_n26928.n41 a_188937_n26928.n40 28.1963
R35801 a_188937_n26928.n67 a_188937_n26928.n66 6.77697
R35802 a_188937_n26928.n121 a_188937_n26928.t14 5.7135
R35803 a_188937_n26928.n121 a_188937_n26928.t10 5.7135
R35804 a_188937_n26928.n93 a_188937_n26928.t16 5.7135
R35805 a_188937_n26928.n93 a_188937_n26928.t12 5.7135
R35806 a_188937_n26928.t20 a_188937_n26928.n157 5.7135
R35807 a_188937_n26928.n157 a_188937_n26928.t18 5.7135
R35808 a_188937_n26928.n21 a_188937_n26928.n136 5.33935
R35809 a_188937_n26928.n22 a_188937_n26928.n126 5.33935
R35810 a_188937_n26928.n120 a_188937_n26928.n110 5.27109
R35811 a_188937_n26928.n113 a_188937_n26928.n104 5.27109
R35812 a_188937_n26928.n37 a_188937_n26928.n84 5.27109
R35813 a_188937_n26928.n86 a_188937_n26928.n78 5.27109
R35814 a_188937_n26928.n40 a_188937_n26928.n63 5.27109
R35815 a_188937_n26928.n68 a_188937_n26928.n59 5.27109
R35816 a_188937_n26928.n130 a_188937_n26928.n57 4.5005
R35817 a_188937_n26928.n140 a_188937_n26928.n55 4.5005
R35818 a_188937_n26928.n119 a_188937_n26928.n109 3.76521
R35819 a_188937_n26928.n114 a_188937_n26928.n105 3.76521
R35820 a_188937_n26928.n92 a_188937_n26928.n83 3.76521
R35821 a_188937_n26928.n87 a_188937_n26928.n79 3.76521
R35822 a_188937_n26928.n56 a_188937_n26928.n133 27.242
R35823 a_188937_n26928.n58 a_188937_n26928.n123 27.242
R35824 a_188937_n26928.n74 a_188937_n26928.n62 3.76521
R35825 a_188937_n26928.n69 a_188937_n26928.n65 3.76521
R35826 a_188937_n26928.n9 a_188937_n26928.n130 3.716
R35827 a_188937_n26928.n52 a_188937_n26928.n51 1.75048
R35828 a_188937_n26928.n53 a_188937_n26928.n54 1.74802
R35829 a_188937_n26928.n132 a_188937_n26928.t21 3.4805
R35830 a_188937_n26928.n132 a_188937_n26928.t0 3.4805
R35831 a_188937_n26928.n131 a_188937_n26928.t1 3.4805
R35832 a_188937_n26928.n131 a_188937_n26928.t3 3.4805
R35833 a_188937_n26928.n48 a_188937_n26928.n147 27.7565
R35834 a_188937_n26928.n45 a_188937_n26928.n154 27.7565
R35835 a_188937_n26928.n140 a_188937_n26928.n9 4.01562
R35836 a_188937_n26928.n118 a_188937_n26928.n108 2.25932
R35837 a_188937_n26928.n115 a_188937_n26928.n106 2.25932
R35838 a_188937_n26928.n91 a_188937_n26928.n82 2.25932
R35839 a_188937_n26928.n88 a_188937_n26928.n80 2.25932
R35840 a_188937_n26928.n138 a_188937_n26928.n133 2.25932
R35841 a_188937_n26928.n128 a_188937_n26928.n123 2.25932
R35842 a_188937_n26928.n73 a_188937_n26928.n64 2.25932
R35843 a_188937_n26928.n70 a_188937_n26928.n60 2.25932
R35844 a_188937_n26928.n147 a_188937_n26928.n144 1.50638
R35845 a_188937_n26928.n154 a_188937_n26928.n151 1.50638
R35846 a_188937_n26928.n137 a_188937_n26928.n135 0.753441
R35847 a_188937_n26928.n127 a_188937_n26928.n125 0.753441
R35848 a_188937_n26928.n53 a_188937_n26928.n101 0.726434
R35849 a_188937_n26928.n14 a_188937_n26928.n0 0.645765
R35850 a_188937_n26928.n142 a_188937_n26928.n141 0.645765
R35851 a_188937_n26928.n101 a_188937_n26928.n13 0.645765
R35852 a_188937_n26928.n97 a_188937_n26928.n96 0.645765
R35853 a_188937_n26928.n100 a_188937_n26928.n54 2.39323
R35854 a_188937_n26928.n96 a_188937_n26928.n51 0.731421
R35855 a_188937_n26928.n100 a_188937_n26928.n99 0.645765
R35856 a_188937_n26928.n99 a_188937_n26928.n98 0.645765
R35857 a_188937_n26928.n98 a_188937_n26928.n95 0.645765
R35858 a_188937_n26928.n52 a_188937_n26928.n95 2.39569
R35859 a_188937_n26928.n47 a_188937_n26928.n10 0.658
R35860 a_188937_n26928.n36 a_188937_n26928.n2 0.649958
R35861 a_188937_n26928.n4 a_188937_n26928.n12 0.645765
R35862 a_188937_n26928.n3 a_188937_n26928.n2 0.645765
R35863 a_188937_n26928.n122 a_188937_n26928.n3 0.645765
R35864 a_188937_n26928.n1 a_188937_n26928.n0 0.645765
R35865 a_188937_n26928.n141 a_188937_n26928.n8 0.631808
R35866 a_188937_n26928.n6 a_188937_n26928.n4 0.630877
R35867 a_188937_n26928.n5 a_188937_n26928.n29 0.584196
R35868 a_188937_n26928.n7 a_188937_n26928.n24 0.584196
R35869 a_188937_n26928.n97 a_188937_n26928.n13 0.56139
R35870 a_188937_n26928.n142 a_188937_n26928.n12 0.56139
R35871 a_188937_n26928.n2 a_188937_n26928.n14 0.446618
R35872 a_188937_n26928.n57 a_188937_n26928.n22 0.411505
R35873 a_188937_n26928.n55 a_188937_n26928.n21 0.411505
R35874 a_188937_n26928.n156 a_188937_n26928.n149 0.3955
R35875 a_188937_n26928.n35 a_188937_n26928.n36 0.391804
R35876 a_188937_n26928.n33 a_188937_n26928.n35 0.391804
R35877 a_188937_n26928.n34 a_188937_n26928.n33 0.391804
R35878 a_188937_n26928.n42 a_188937_n26928.n34 0.391804
R35879 a_188937_n26928.n30 a_188937_n26928.n31 0.391804
R35880 a_188937_n26928.n28 a_188937_n26928.n30 0.391804
R35881 a_188937_n26928.n29 a_188937_n26928.n28 0.391804
R35882 a_188937_n26928.n25 a_188937_n26928.n26 0.391804
R35883 a_188937_n26928.n23 a_188937_n26928.n25 0.391804
R35884 a_188937_n26928.n24 a_188937_n26928.n23 0.391804
R35885 a_188937_n26928.n19 a_188937_n26928.n18 0.391804
R35886 a_188937_n26928.n46 a_188937_n26928.n19 0.391804
R35887 a_188937_n26928.n16 a_188937_n26928.n15 0.391804
R35888 a_188937_n26928.n43 a_188937_n26928.n16 0.391804
R35889 a_188937_n26928.n31 a_188937_n26928.n32 0.388109
R35890 a_188937_n26928.n26 a_188937_n26928.n27 0.388109
R35891 a_188937_n26928.n11 a_188937_n26928.n42 0.387101
R35892 a_188937_n26928.n156 a_188937_n26928.n15 0.368217
R35893 a_188937_n26928.n149 a_188937_n26928.n18 0.368217
R35894 a_188937_n26928.n47 a_188937_n26928.n46 0.364413
R35895 a_188937_n26928.n44 a_188937_n26928.n43 0.364413
R35896 a_188937_n26928.n10 a_188937_n26928.n44 0.363
R35897 a_188937_n26928.n6 a_188937_n26928.n5 0.363
R35898 a_188937_n26928.n8 a_188937_n26928.n7 0.363
R35899 a_188937_n26928.n32 a_188937_n26928.n3 0.358
R35900 a_188937_n26928.n1 a_188937_n26928.n27 0.358
R35901 a_188937_n26928.n12 a_188937_n26928.n11 0.353
R35902 a_157137_n26928.n152 a_157137_n26928.n43 194.291
R35903 a_157137_n26928.n152 a_157137_n26928.n93 585
R35904 a_157137_n26928.n152 a_157137_n26928.n92 585
R35905 a_157137_n26928.n152 a_157137_n26928.n91 585
R35906 a_157137_n26928.n152 a_157137_n26928.n89 585
R35907 a_157137_n26928.n152 a_157137_n26928.n88 585
R35908 a_157137_n26928.n152 a_157137_n26928.n87 585
R35909 a_157137_n26928.n152 a_157137_n26928.n86 585
R35910 a_157137_n26928.n152 a_157137_n26928.n51 291.375
R35911 a_157137_n26928.n113 a_157137_n26928.n40 194.291
R35912 a_157137_n26928.n113 a_157137_n26928.n102 585
R35913 a_157137_n26928.n113 a_157137_n26928.n101 585
R35914 a_157137_n26928.n113 a_157137_n26928.n100 585
R35915 a_157137_n26928.n113 a_157137_n26928.n98 585
R35916 a_157137_n26928.n113 a_157137_n26928.n97 585
R35917 a_157137_n26928.n113 a_157137_n26928.n96 585
R35918 a_157137_n26928.n113 a_157137_n26928.n95 585
R35919 a_157137_n26928.n113 a_157137_n26928.n94 585
R35920 a_157137_n26928.n113 a_157137_n26928.n50 585
R35921 a_157137_n26928.n157 a_157137_n26928.n39 194.291
R35922 a_157137_n26928.n157 a_157137_n26928.n65 585
R35923 a_157137_n26928.n157 a_157137_n26928.n64 585
R35924 a_157137_n26928.n157 a_157137_n26928.n66 585
R35925 a_157137_n26928.n157 a_157137_n26928.n62 585
R35926 a_157137_n26928.n157 a_157137_n26928.n67 585
R35927 a_157137_n26928.n157 a_157137_n26928.n61 585
R35928 a_157137_n26928.n157 a_157137_n26928.n68 585
R35929 a_157137_n26928.n157 a_157137_n26928.n60 585
R35930 a_157137_n26928.n157 a_157137_n26928.n156 585
R35931 a_157137_n26928.t3 a_157137_n26928.n9 308.31
R35932 a_157137_n26928.n135 a_157137_n26928.t3 308.31
R35933 a_157137_n26928.t1 a_157137_n26928.n142 308.31
R35934 a_157137_n26928.n9 a_157137_n26928.t1 308.31
R35935 a_157137_n26928.n152 a_157137_n26928.n90 286.238
R35936 a_157137_n26928.n113 a_157137_n26928.n99 286.238
R35937 a_157137_n26928.n157 a_157137_n26928.n63 286.238
R35938 a_157137_n26928.n57 a_157137_n26928.n56 6.98494
R35939 a_157137_n26928.n59 a_157137_n26928.n58 6.98494
R35940 a_157137_n26928.n55 a_157137_n26928.t23 104.094
R35941 a_157137_n26928.n4 a_157137_n26928.t13 209.939
R35942 a_157137_n26928.t15 a_157137_n26928.n6 209.938
R35943 a_157137_n26928.t22 a_157137_n26928.n53 104.094
R35944 a_157137_n26928.t11 a_157137_n26928.n14 209.93
R35945 a_157137_n26928.n10 a_157137_n26928.t11 209.93
R35946 a_157137_n26928.t7 a_157137_n26928.n128 209.93
R35947 a_157137_n26928.n2 a_157137_n26928.t7 209.93
R35948 a_157137_n26928.n1 a_157137_n26928.t15 209.93
R35949 a_157137_n26928.t5 a_157137_n26928.n0 209.93
R35950 a_157137_n26928.n85 a_157137_n26928.t5 209.93
R35951 a_157137_n26928.n15 a_157137_n26928.t9 209.93
R35952 a_157137_n26928.t9 a_157137_n26928.n12 209.93
R35953 a_157137_n26928.n155 a_157137_n26928.t27 209.93
R35954 a_157137_n26928.t27 a_157137_n26928.n154 209.93
R35955 a_157137_n26928.t25 a_157137_n26928.n84 209.93
R35956 a_157137_n26928.n153 a_157137_n26928.t25 209.93
R35957 a_157137_n26928.n114 a_157137_n26928.t24 209.93
R35958 a_157137_n26928.t24 a_157137_n26928.n11 209.93
R35959 a_157137_n26928.t26 a_157137_n26928.n115 209.93
R35960 a_157137_n26928.n116 a_157137_n26928.t26 209.93
R35961 a_157137_n26928.t13 a_157137_n26928.n127 209.93
R35962 a_157137_n26928.n134 a_157137_n26928.n49 92.3135
R35963 a_157137_n26928.n134 a_157137_n26928.n130 185
R35964 a_157137_n26928.n134 a_157137_n26928.n21 92.3135
R35965 a_157137_n26928.n141 a_157137_n26928.n46 92.3135
R35966 a_157137_n26928.n141 a_157137_n26928.n137 185
R35967 a_157137_n26928.n141 a_157137_n26928.n18 92.3135
R35968 a_157137_n26928.n125 a_157137_n26928.n124 185
R35969 a_157137_n26928.n121 a_157137_n26928.n120 185
R35970 a_157137_n26928.n75 a_157137_n26928.n74 185
R35971 a_157137_n26928.n71 a_157137_n26928.n70 185
R35972 a_157137_n26928.n122 a_157137_n26928.t18 174.857
R35973 a_157137_n26928.n72 a_157137_n26928.t20 174.857
R35974 a_157137_n26928.n57 a_157137_n26928.n125 244.714
R35975 a_157137_n26928.n125 a_157137_n26928.n120 140.69
R35976 a_157137_n26928.n59 a_157137_n26928.n75 244.714
R35977 a_157137_n26928.n75 a_157137_n26928.n70 140.69
R35978 a_157137_n26928.n134 a_157137_n26928.n129 86.5152
R35979 a_157137_n26928.n141 a_157137_n26928.n136 86.5152
R35980 a_157137_n26928.t18 a_157137_n26928.n120 70.3453
R35981 a_157137_n26928.t20 a_157137_n26928.n70 70.3453
R35982 a_157137_n26928.n122 a_157137_n26928.n121 28.4333
R35983 a_157137_n26928.n72 a_157137_n26928.n71 28.4333
R35984 a_157137_n26928.n132 a_157137_n26928.n130 25.6005
R35985 a_157137_n26928.n139 a_157137_n26928.n137 25.6005
R35986 a_157137_n26928.n148 a_157137_n26928.n91 24.8476
R35987 a_157137_n26928.n147 a_157137_n26928.n89 24.8476
R35988 a_157137_n26928.n109 a_157137_n26928.n100 24.8476
R35989 a_157137_n26928.n108 a_157137_n26928.n98 24.8476
R35990 a_157137_n26928.n124 a_157137_n26928.n123 24.8476
R35991 a_157137_n26928.n74 a_157137_n26928.n73 24.8476
R35992 a_157137_n26928.n81 a_157137_n26928.n66 24.8476
R35993 a_157137_n26928.n80 a_157137_n26928.n62 24.8476
R35994 a_157137_n26928.n131 a_157137_n26928.n21 27.7565
R35995 a_157137_n26928.n138 a_157137_n26928.n18 27.7565
R35996 a_157137_n26928.n149 a_157137_n26928.n92 23.3417
R35997 a_157137_n26928.n146 a_157137_n26928.n88 23.3417
R35998 a_157137_n26928.n110 a_157137_n26928.n101 23.3417
R35999 a_157137_n26928.n107 a_157137_n26928.n97 23.3417
R36000 a_157137_n26928.n82 a_157137_n26928.n64 23.3417
R36001 a_157137_n26928.n79 a_157137_n26928.n67 23.3417
R36002 a_157137_n26928.n49 a_157137_n26928.n48 6.60954
R36003 a_157137_n26928.n21 a_157137_n26928.n19 6.60954
R36004 a_157137_n26928.n46 a_157137_n26928.n45 6.60954
R36005 a_157137_n26928.n18 a_157137_n26928.n16 6.60954
R36006 a_157137_n26928.n8 a_157137_n26928.n117 22.3909
R36007 a_157137_n26928.n8 a_157137_n26928.n118 22.3909
R36008 a_157137_n26928.n150 a_157137_n26928.n93 21.8358
R36009 a_157137_n26928.n145 a_157137_n26928.n87 21.8358
R36010 a_157137_n26928.n111 a_157137_n26928.n102 21.8358
R36011 a_157137_n26928.n106 a_157137_n26928.n96 21.8358
R36012 a_157137_n26928.n83 a_157137_n26928.n65 21.8358
R36013 a_157137_n26928.n78 a_157137_n26928.n61 21.8358
R36014 a_157137_n26928.n144 a_157137_n26928.n86 20.3299
R36015 a_157137_n26928.n105 a_157137_n26928.n95 20.3299
R36016 a_157137_n26928.n77 a_157137_n26928.n68 20.3299
R36017 a_157137_n26928.n2 a_157137_n26928.n50 19.0887
R36018 a_157137_n26928.n156 a_157137_n26928.n1 19.0887
R36019 a_157137_n26928.n43 a_157137_n26928.n13 6.07169
R36020 a_157137_n26928.n143 a_157137_n26928.n51 24.6333
R36021 a_157137_n26928.n40 a_157137_n26928.n3 6.07169
R36022 a_157137_n26928.n104 a_157137_n26928.n94 18.824
R36023 a_157137_n26928.n5 a_157137_n26928.n39 6.07169
R36024 a_157137_n26928.n76 a_157137_n26928.n60 18.824
R36025 a_157137_n26928.n10 a_157137_n26928.n51 9.76605
R36026 a_157137_n26928.n103 a_157137_n26928.n50 17.3181
R36027 a_157137_n26928.n156 a_157137_n26928.n41 17.3181
R36028 a_157137_n26928.n131 a_157137_n26928.n129 13.4786
R36029 a_157137_n26928.n138 a_157137_n26928.n136 13.4786
R36030 a_157137_n26928.n148 a_157137_n26928.n90 13.2799
R36031 a_157137_n26928.n147 a_157137_n26928.n90 13.2799
R36032 a_157137_n26928.n109 a_157137_n26928.n99 13.2799
R36033 a_157137_n26928.n108 a_157137_n26928.n99 13.2799
R36034 a_157137_n26928.n81 a_157137_n26928.n63 13.2799
R36035 a_157137_n26928.n80 a_157137_n26928.n63 13.2799
R36036 a_157137_n26928.n132 a_157137_n26928.n129 11.9727
R36037 a_157137_n26928.n139 a_157137_n26928.n136 11.9727
R36038 a_157137_n26928.n10 a_157137_n26928.n9 9.61161
R36039 a_157137_n26928.n6 a_157137_n26928.n52 9.47511
R36040 a_157137_n26928.n4 a_157137_n26928.n54 9.47106
R36041 a_157137_n26928.n11 a_157137_n26928.n14 9.3755
R36042 a_157137_n26928.n44 a_157137_n26928.n140 9.3005
R36043 a_157137_n26928.n17 a_157137_n26928.n139 9.3005
R36044 a_157137_n26928.n17 a_157137_n26928.n138 9.3005
R36045 a_157137_n26928.n47 a_157137_n26928.n133 9.3005
R36046 a_157137_n26928.n20 a_157137_n26928.n132 9.3005
R36047 a_157137_n26928.n20 a_157137_n26928.n131 9.3005
R36048 a_157137_n26928.n123 a_157137_n26928.n22 9.3005
R36049 a_157137_n26928.n119 a_157137_n26928.n22 9.3005
R36050 a_157137_n26928.n73 a_157137_n26928.n23 9.3005
R36051 a_157137_n26928.n69 a_157137_n26928.n23 9.3005
R36052 a_157137_n26928.n28 a_157137_n26928.n103 9.3005
R36053 a_157137_n26928.n24 a_157137_n26928.n109 9.3005
R36054 a_157137_n26928.n24 a_157137_n26928.n110 9.3005
R36055 a_157137_n26928.n25 a_157137_n26928.n111 9.3005
R36056 a_157137_n26928.n25 a_157137_n26928.n112 9.3005
R36057 a_157137_n26928.n26 a_157137_n26928.n108 9.3005
R36058 a_157137_n26928.n26 a_157137_n26928.n107 9.3005
R36059 a_157137_n26928.n27 a_157137_n26928.n106 9.3005
R36060 a_157137_n26928.n27 a_157137_n26928.n105 9.3005
R36061 a_157137_n26928.n28 a_157137_n26928.n104 9.3005
R36062 a_157137_n26928.n29 a_157137_n26928.n148 9.3005
R36063 a_157137_n26928.n30 a_157137_n26928.n149 9.3005
R36064 a_157137_n26928.n30 a_157137_n26928.n150 9.3005
R36065 a_157137_n26928.n42 a_157137_n26928.n151 9.3005
R36066 a_157137_n26928.n29 a_157137_n26928.n147 9.3005
R36067 a_157137_n26928.n31 a_157137_n26928.n146 9.3005
R36068 a_157137_n26928.n31 a_157137_n26928.n145 9.3005
R36069 a_157137_n26928.n32 a_157137_n26928.n144 9.3005
R36070 a_157137_n26928.n32 a_157137_n26928.n143 9.3005
R36071 a_157137_n26928.n33 a_157137_n26928.n81 9.3005
R36072 a_157137_n26928.n33 a_157137_n26928.n82 9.3005
R36073 a_157137_n26928.n34 a_157137_n26928.n83 9.3005
R36074 a_157137_n26928.n34 a_157137_n26928.n38 9.3005
R36075 a_157137_n26928.n35 a_157137_n26928.n80 9.3005
R36076 a_157137_n26928.n35 a_157137_n26928.n79 9.3005
R36077 a_157137_n26928.n36 a_157137_n26928.n78 9.3005
R36078 a_157137_n26928.n36 a_157137_n26928.n77 9.3005
R36079 a_157137_n26928.n37 a_157137_n26928.n76 9.3005
R36080 a_157137_n26928.n37 a_157137_n26928.n41 9.3005
R36081 a_157137_n26928.n103 a_157137_n26928.n94 8.28285
R36082 a_157137_n26928.n41 a_157137_n26928.n60 8.28285
R36083 a_157137_n26928.n1 a_157137_n26928.n7 7.04926
R36084 a_157137_n26928.n127 a_157137_n26928.n126 6.96926
R36085 a_157137_n26928.n134 a_157137_n26928.t4 6.9605
R36086 a_157137_n26928.n141 a_157137_n26928.t2 6.9605
R36087 a_157137_n26928.n43 a_157137_n26928.n151 28.1963
R36088 a_157137_n26928.n143 a_157137_n26928.n86 6.77697
R36089 a_157137_n26928.n40 a_157137_n26928.n112 28.1963
R36090 a_157137_n26928.n104 a_157137_n26928.n95 6.77697
R36091 a_157137_n26928.n39 a_157137_n26928.n38 28.1963
R36092 a_157137_n26928.n76 a_157137_n26928.n68 6.77697
R36093 a_157137_n26928.n152 a_157137_n26928.t12 5.7135
R36094 a_157137_n26928.n152 a_157137_n26928.t10 5.7135
R36095 a_157137_n26928.n113 a_157137_n26928.t14 5.7135
R36096 a_157137_n26928.n113 a_157137_n26928.t8 5.7135
R36097 a_157137_n26928.n157 a_157137_n26928.t6 5.7135
R36098 a_157137_n26928.t16 a_157137_n26928.n157 5.7135
R36099 a_157137_n26928.n22 a_157137_n26928.n122 5.33935
R36100 a_157137_n26928.n23 a_157137_n26928.n72 5.33935
R36101 a_157137_n26928.n151 a_157137_n26928.n93 5.27109
R36102 a_157137_n26928.n144 a_157137_n26928.n87 5.27109
R36103 a_157137_n26928.n112 a_157137_n26928.n102 5.27109
R36104 a_157137_n26928.n105 a_157137_n26928.n96 5.27109
R36105 a_157137_n26928.n38 a_157137_n26928.n65 5.27109
R36106 a_157137_n26928.n77 a_157137_n26928.n61 5.27109
R36107 a_157137_n26928.n7 a_157137_n26928.n58 4.5005
R36108 a_157137_n26928.n126 a_157137_n26928.n56 4.5005
R36109 a_157137_n26928.n150 a_157137_n26928.n92 3.76521
R36110 a_157137_n26928.n145 a_157137_n26928.n88 3.76521
R36111 a_157137_n26928.n111 a_157137_n26928.n101 3.76521
R36112 a_157137_n26928.n106 a_157137_n26928.n97 3.76521
R36113 a_157137_n26928.n57 a_157137_n26928.n119 27.242
R36114 a_157137_n26928.n59 a_157137_n26928.n69 27.242
R36115 a_157137_n26928.n83 a_157137_n26928.n64 3.76521
R36116 a_157137_n26928.n78 a_157137_n26928.n67 3.76521
R36117 a_157137_n26928.n8 a_157137_n26928.n7 3.716
R36118 a_157137_n26928.n52 a_157137_n26928.n53 1.75048
R36119 a_157137_n26928.n54 a_157137_n26928.n55 1.74802
R36120 a_157137_n26928.n117 a_157137_n26928.t0 3.4805
R36121 a_157137_n26928.n117 a_157137_n26928.t21 3.4805
R36122 a_157137_n26928.n118 a_157137_n26928.t17 3.4805
R36123 a_157137_n26928.n118 a_157137_n26928.t19 3.4805
R36124 a_157137_n26928.n49 a_157137_n26928.n133 27.7565
R36125 a_157137_n26928.n46 a_157137_n26928.n140 27.7565
R36126 a_157137_n26928.n126 a_157137_n26928.n8 4.01562
R36127 a_157137_n26928.n149 a_157137_n26928.n91 2.25932
R36128 a_157137_n26928.n146 a_157137_n26928.n89 2.25932
R36129 a_157137_n26928.n110 a_157137_n26928.n100 2.25932
R36130 a_157137_n26928.n107 a_157137_n26928.n98 2.25932
R36131 a_157137_n26928.n124 a_157137_n26928.n119 2.25932
R36132 a_157137_n26928.n74 a_157137_n26928.n69 2.25932
R36133 a_157137_n26928.n82 a_157137_n26928.n66 2.25932
R36134 a_157137_n26928.n79 a_157137_n26928.n62 2.25932
R36135 a_157137_n26928.n133 a_157137_n26928.n130 1.50638
R36136 a_157137_n26928.n140 a_157137_n26928.n137 1.50638
R36137 a_157137_n26928.n123 a_157137_n26928.n121 0.753441
R36138 a_157137_n26928.n73 a_157137_n26928.n71 0.753441
R36139 a_157137_n26928.n54 a_157137_n26928.n116 0.726434
R36140 a_157137_n26928.n12 a_157137_n26928.n85 0.645765
R36141 a_157137_n26928.n116 a_157137_n26928.n11 0.645765
R36142 a_157137_n26928.n154 a_157137_n26928.n153 0.645765
R36143 a_157137_n26928.n115 a_157137_n26928.n55 2.39323
R36144 a_157137_n26928.n154 a_157137_n26928.n52 0.731421
R36145 a_157137_n26928.n115 a_157137_n26928.n114 0.645765
R36146 a_157137_n26928.n114 a_157137_n26928.n84 0.645765
R36147 a_157137_n26928.n155 a_157137_n26928.n84 0.645765
R36148 a_157137_n26928.n53 a_157137_n26928.n155 2.39569
R36149 a_157137_n26928.n48 a_157137_n26928.n9 0.658
R36150 a_157137_n26928.n32 a_157137_n26928.n10 0.649958
R36151 a_157137_n26928.n10 a_157137_n26928.n2 0.645765
R36152 a_157137_n26928.n128 a_157137_n26928.n14 0.645765
R36153 a_157137_n26928.n15 a_157137_n26928.n0 0.645765
R36154 a_157137_n26928.n127 a_157137_n26928.n2 0.645765
R36155 a_157137_n26928.n1 a_157137_n26928.n0 0.645765
R36156 a_157137_n26928.n85 a_157137_n26928.n6 0.631808
R36157 a_157137_n26928.n128 a_157137_n26928.n4 0.630877
R36158 a_157137_n26928.n5 a_157137_n26928.n34 0.584196
R36159 a_157137_n26928.n3 a_157137_n26928.n25 0.584196
R36160 a_157137_n26928.n14 a_157137_n26928.n12 0.56139
R36161 a_157137_n26928.n153 a_157137_n26928.n11 0.56139
R36162 a_157137_n26928.n10 a_157137_n26928.n15 0.446618
R36163 a_157137_n26928.n58 a_157137_n26928.n23 0.411505
R36164 a_157137_n26928.n56 a_157137_n26928.n22 0.411505
R36165 a_157137_n26928.n142 a_157137_n26928.n135 0.3955
R36166 a_157137_n26928.n35 a_157137_n26928.n36 0.391804
R36167 a_157137_n26928.n33 a_157137_n26928.n35 0.391804
R36168 a_157137_n26928.n34 a_157137_n26928.n33 0.391804
R36169 a_157137_n26928.n31 a_157137_n26928.n32 0.391804
R36170 a_157137_n26928.n29 a_157137_n26928.n31 0.391804
R36171 a_157137_n26928.n30 a_157137_n26928.n29 0.391804
R36172 a_157137_n26928.n42 a_157137_n26928.n30 0.391804
R36173 a_157137_n26928.n26 a_157137_n26928.n27 0.391804
R36174 a_157137_n26928.n24 a_157137_n26928.n26 0.391804
R36175 a_157137_n26928.n25 a_157137_n26928.n24 0.391804
R36176 a_157137_n26928.n20 a_157137_n26928.n19 0.391804
R36177 a_157137_n26928.n47 a_157137_n26928.n20 0.391804
R36178 a_157137_n26928.n17 a_157137_n26928.n16 0.391804
R36179 a_157137_n26928.n44 a_157137_n26928.n17 0.391804
R36180 a_157137_n26928.n36 a_157137_n26928.n37 0.388109
R36181 a_157137_n26928.n27 a_157137_n26928.n28 0.388109
R36182 a_157137_n26928.n13 a_157137_n26928.n42 0.387101
R36183 a_157137_n26928.n142 a_157137_n26928.n16 0.368217
R36184 a_157137_n26928.n135 a_157137_n26928.n19 0.368217
R36185 a_157137_n26928.n48 a_157137_n26928.n47 0.364413
R36186 a_157137_n26928.n45 a_157137_n26928.n44 0.364413
R36187 a_157137_n26928.n9 a_157137_n26928.n45 0.363
R36188 a_157137_n26928.n4 a_157137_n26928.n3 0.363
R36189 a_157137_n26928.n6 a_157137_n26928.n5 0.363
R36190 a_157137_n26928.n1 a_157137_n26928.n37 0.358
R36191 a_157137_n26928.n28 a_157137_n26928.n2 0.358
R36192 a_157137_n26928.n14 a_157137_n26928.n13 0.353
R36193 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t19 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n98 210.794
R36194 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t44 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n96 210.794
R36195 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n97 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t44 210.794
R36196 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n95 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t27 210.794
R36197 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t27 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n19 210.794
R36198 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t33 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n94 210.794
R36199 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n52 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t23 210.794
R36200 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t23 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n29 210.794
R36201 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n51 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t43 210.794
R36202 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t43 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n50 210.794
R36203 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t34 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n30 210.794
R36204 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n49 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t34 210.794
R36205 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t41 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n47 210.794
R36206 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n48 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t41 210.794
R36207 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n46 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t39 210.794
R36208 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t39 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n31 210.794
R36209 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n45 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t29 210.794
R36210 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t29 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n44 210.794
R36211 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t18 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n32 210.794
R36212 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n43 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t18 210.794
R36213 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t22 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n41 210.794
R36214 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n42 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t22 210.794
R36215 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n40 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t17 210.794
R36216 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t17 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n33 210.794
R36217 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n39 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t47 210.794
R36218 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t47 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n38 210.794
R36219 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t21 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n34 210.794
R36220 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n37 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t21 210.794
R36221 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n36 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t38 210.794
R36222 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t38 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n35 210.794
R36223 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t25 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n28 210.794
R36224 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n53 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t25 210.794
R36225 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n55 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t40 210.794
R36226 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t40 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n54 210.794
R36227 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n56 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t37 210.794
R36228 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t37 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n27 210.794
R36229 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t28 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n57 210.794
R36230 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n58 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t28 210.794
R36231 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t36 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n26 210.794
R36232 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n59 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t36 210.794
R36233 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n61 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t32 210.794
R36234 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t32 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n60 210.794
R36235 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n62 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t16 210.794
R36236 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t16 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n25 210.794
R36237 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t46 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n63 210.794
R36238 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n64 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t46 210.794
R36239 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t20 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n24 210.794
R36240 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n65 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t20 210.794
R36241 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n67 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t45 210.794
R36242 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t45 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n66 210.794
R36243 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n68 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t42 210.794
R36244 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t42 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n23 210.794
R36245 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t35 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n69 210.794
R36246 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n70 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t35 210.794
R36247 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t31 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n22 210.794
R36248 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n71 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t31 210.794
R36249 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n73 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t26 210.794
R36250 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t26 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n72 210.794
R36251 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n82 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n81 185
R36252 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n14 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n13 185
R36253 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t14 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n99 120.469
R36254 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n92 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t8 120.465
R36255 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n89 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t12 120.419
R36256 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t12 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n88 120.419
R36257 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t8 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n91 120.419
R36258 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n100 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t14 120.419
R36259 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n87 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t10 120.419
R36260 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t10 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n86 120.419
R36261 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n93 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t30 104.566
R36262 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n18 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t24 104.562
R36263 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n81 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n80 86.5152
R36264 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n15 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n14 86.5152
R36265 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n8 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n7 50.9993
R36266 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n102 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n101 47.5895
R36267 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n76 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n21 47.5893
R36268 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n85 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n84 38.0154
R36269 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n82 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n78 25.6005
R36270 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n13 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n11 25.6005
R36271 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n80 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n79 22.7786
R36272 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n16 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n15 22.7786
R36273 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n4 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n3 0.0650981
R36274 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n4 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t19 210.808
R36275 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t33 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n6 210.808
R36276 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n5 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n6 0.0650981
R36277 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n81 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t9 13.9205
R36278 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n81 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t13 13.9205
R36279 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n14 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t11 13.9205
R36280 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n14 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t15 13.9205
R36281 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n80 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n78 11.9727
R36282 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n15 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n11 11.9727
R36283 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n83 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n82 10.8064
R36284 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n13 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n12 10.8064
R36285 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n5 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n92 9.59564
R36286 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n99 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n3 9.59208
R36287 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n11 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n10 9.3005
R36288 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n78 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n77 9.3005
R36289 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n91 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n76 8.93258
R36290 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n102 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n100 8.84758
R36291 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n84 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t1 6.9605
R36292 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n84 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t0 6.9605
R36293 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n7 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t5 5.7135
R36294 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n7 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t4 5.7135
R36295 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n21 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t6 5.7135
R36296 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n21 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t3 5.7135
R36297 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n101 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t2 5.7135
R36298 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n101 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t7 5.7135
R36299 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n1 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n29 4.293
R36300 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n36 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n2 4.218
R36301 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n1 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n52 3.94612
R36302 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n35 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n2 3.87112
R36303 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n76 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n75 3.4105
R36304 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n103 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n102 3.4105
R36305 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n28 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n0 3.29712
R36306 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n53 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n1 3.29612
R36307 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n72 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n2 3.23112
R36308 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n74 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n73 3.23112
R36309 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n98 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n18 2.3168
R36310 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n103 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n0 2.31333
R36311 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n94 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n93 2.31188
R36312 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n75 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n74 2.30692
R36313 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n93 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n6 2.28563
R36314 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n94 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n19 0.645765
R36315 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n97 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n19 0.645765
R36316 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n98 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n97 0.645765
R36317 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n96 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n95 0.645765
R36318 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n88 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n87 0.645765
R36319 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n37 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n36 0.645765
R36320 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n38 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n37 0.645765
R36321 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n38 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n33 0.645765
R36322 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n42 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n33 0.645765
R36323 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n43 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n42 0.645765
R36324 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n44 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n43 0.645765
R36325 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n44 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n31 0.645765
R36326 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n48 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n31 0.645765
R36327 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n49 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n48 0.645765
R36328 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n50 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n49 0.645765
R36329 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n50 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n29 0.645765
R36330 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n35 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n34 0.645765
R36331 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n39 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n34 0.645765
R36332 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n40 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n39 0.645765
R36333 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n41 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n40 0.645765
R36334 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n41 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n32 0.645765
R36335 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n45 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n32 0.645765
R36336 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n46 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n45 0.645765
R36337 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n47 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n46 0.645765
R36338 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n47 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n30 0.645765
R36339 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n51 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n30 0.645765
R36340 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n52 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n51 0.645765
R36341 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n72 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n71 0.645765
R36342 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n71 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n70 0.645765
R36343 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n70 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n23 0.645765
R36344 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n66 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n23 0.645765
R36345 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n66 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n65 0.645765
R36346 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n65 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n64 0.645765
R36347 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n64 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n25 0.645765
R36348 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n60 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n25 0.645765
R36349 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n60 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n59 0.645765
R36350 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n59 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n58 0.645765
R36351 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n58 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n27 0.645765
R36352 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n54 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n27 0.645765
R36353 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n54 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n53 0.645765
R36354 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n73 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n22 0.645765
R36355 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n69 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n22 0.645765
R36356 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n69 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n68 0.645765
R36357 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n68 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n67 0.645765
R36358 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n67 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n24 0.645765
R36359 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n63 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n24 0.645765
R36360 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n63 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n62 0.645765
R36361 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n62 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n61 0.645765
R36362 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n61 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n26 0.645765
R36363 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n57 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n26 0.645765
R36364 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n57 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n56 0.645765
R36365 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n56 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n55 0.645765
R36366 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n55 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n28 0.645765
R36367 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n96 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n3 0.552061
R36368 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n95 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n5 0.550633
R36369 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n88 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n20 0.333133
R36370 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n90 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n89 0.333133
R36371 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n86 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n9 0.323133
R36372 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n100 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n9 0.323133
R36373 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n87 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n17 0.323133
R36374 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n91 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n90 0.313133
R36375 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n86 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n85 0.278133
R36376 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n89 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n85 0.268133
R36377 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n99 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n17 0.256274
R36378 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n92 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n20 0.252692
R36379 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n90 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n83 0.219522
R36380 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n12 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n9 0.217348
R36381 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n17 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n16 0.217348
R36382 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n79 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n20 0.216386
R36383 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n103 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n8 0.204167
R36384 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n75 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n8 0.204167
R36385 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n12 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n10 0.196152
R36386 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n16 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n10 0.196152
R36387 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n83 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n77 0.196152
R36388 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n79 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n77 0.196152
R36389 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n4 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n18 2.28913
R36390 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n74 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n2 0.4755
R36391 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n1 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n0 0.4755
R36392 a_214193_n11375.n5 a_214193_n11375.n4 7.70214
R36393 a_214193_n11375.n1 a_214193_n11375.n0 7.69294
R36394 a_214193_n11375.n5 a_214193_n11375.t2 2.81388
R36395 a_214193_n11375.t0 a_214193_n11375.n5 2.81161
R36396 a_214193_n11375.n0 a_214193_n11375.t1 2.80271
R36397 a_214193_n11375.n0 a_214193_n11375.t7 2.80044
R36398 a_214193_n11375.n2 a_214193_n11375.n1 0.522904
R36399 a_214193_n11375.n3 a_214193_n11375.n2 0.522904
R36400 a_214193_n11375.n4 a_214193_n11375.n3 0.522904
R36401 a_214193_n11375.n1 a_214193_n11375.t5 0.0535478
R36402 a_214193_n11375.n2 a_214193_n11375.t4 0.0535478
R36403 a_214193_n11375.n3 a_214193_n11375.t3 0.0535478
R36404 a_214193_n11375.n4 a_214193_n11375.t6 0.0535478
R36405 a_156122_n20028.n31 a_156122_n20028.n193 91.4185
R36406 a_156122_n20028.n56 a_156122_n20028.n193 14.3253
R36407 a_156122_n20028.n33 a_156122_n20028.n196 91.4185
R36408 a_156122_n20028.n58 a_156122_n20028.n196 14.3253
R36409 a_156122_n20028.n35 a_156122_n20028.n69 91.4185
R36410 a_156122_n20028.n60 a_156122_n20028.n69 14.3253
R36411 a_156122_n20028.n37 a_156122_n20028.n129 91.4185
R36412 a_156122_n20028.n62 a_156122_n20028.n129 14.3253
R36413 a_156122_n20028.n39 a_156122_n20028.n132 91.4185
R36414 a_156122_n20028.n64 a_156122_n20028.n132 14.3253
R36415 a_156122_n20028.n77 a_156122_n20028.n15 15.3734
R36416 a_156122_n20028.n77 a_156122_n20028.n72 185
R36417 a_156122_n20028.n77 a_156122_n20028.n23 91.4184
R36418 a_156122_n20028.n83 a_156122_n20028.n17 15.3734
R36419 a_156122_n20028.n83 a_156122_n20028.n78 185
R36420 a_156122_n20028.n83 a_156122_n20028.n25 91.4184
R36421 a_156122_n20028.n89 a_156122_n20028.n19 15.3734
R36422 a_156122_n20028.n89 a_156122_n20028.n84 185
R36423 a_156122_n20028.n89 a_156122_n20028.n27 91.4184
R36424 a_156122_n20028.n97 a_156122_n20028.n96 185
R36425 a_156122_n20028.n94 a_156122_n20028.n93 185
R36426 a_156122_n20028.n102 a_156122_n20028.n101 185
R36427 a_156122_n20028.n104 a_156122_n20028.n103 185
R36428 a_156122_n20028.n91 a_156122_n20028.n90 185
R36429 a_156122_n20028.n192 a_156122_n20028.n191 185
R36430 a_156122_n20028.n189 a_156122_n20028.n175 185
R36431 a_156122_n20028.n179 a_156122_n20028.n176 185
R36432 a_156122_n20028.n184 a_156122_n20028.n183 185
R36433 a_156122_n20028.n182 a_156122_n20028.n181 185
R36434 a_156122_n20028.n158 a_156122_n20028.n157 185
R36435 a_156122_n20028.n165 a_156122_n20028.n164 185
R36436 a_156122_n20028.n166 a_156122_n20028.n155 185
R36437 a_156122_n20028.n171 a_156122_n20028.n170 185
R36438 a_156122_n20028.n169 a_156122_n20028.n168 185
R36439 a_156122_n20028.n50 a_156122_n20028.n148 91.4187
R36440 a_156122_n20028.n149 a_156122_n20028.n148 185
R36441 a_156122_n20028.n9 a_156122_n20028.n148 15.371
R36442 a_156122_n20028.n52 a_156122_n20028.n142 91.4187
R36443 a_156122_n20028.n143 a_156122_n20028.n142 185
R36444 a_156122_n20028.n11 a_156122_n20028.n142 15.371
R36445 a_156122_n20028.n54 a_156122_n20028.n136 91.4187
R36446 a_156122_n20028.n137 a_156122_n20028.n136 185
R36447 a_156122_n20028.n13 a_156122_n20028.n136 15.371
R36448 a_156122_n20028.n116 a_156122_n20028.n115 185
R36449 a_156122_n20028.n117 a_156122_n20028.n110 185
R36450 a_156122_n20028.n126 a_156122_n20028.n125 185
R36451 a_156122_n20028.n124 a_156122_n20028.n123 185
R36452 a_156122_n20028.n119 a_156122_n20028.n118 185
R36453 a_156122_n20028.n200 a_156122_n20028.n45 91.4185
R36454 a_156122_n20028.n200 a_156122_n20028.n68 14.3253
R36455 a_156122_n20028.t27 a_156122_n20028.n95 174.857
R36456 a_156122_n20028.n180 a_156122_n20028.t21 174.857
R36457 a_156122_n20028.n167 a_156122_n20028.t0 174.857
R36458 a_156122_n20028.n120 a_156122_n20028.t20 174.857
R36459 a_156122_n20028.n96 a_156122_n20028.n93 140.69
R36460 a_156122_n20028.n102 a_156122_n20028.n93 140.69
R36461 a_156122_n20028.n103 a_156122_n20028.n102 140.69
R36462 a_156122_n20028.n103 a_156122_n20028.n90 140.69
R36463 a_156122_n20028.n29 a_156122_n20028.n90 256.962
R36464 a_156122_n20028.n40 a_156122_n20028.n192 256.962
R36465 a_156122_n20028.n192 a_156122_n20028.n175 140.69
R36466 a_156122_n20028.n179 a_156122_n20028.n175 140.69
R36467 a_156122_n20028.n183 a_156122_n20028.n179 140.69
R36468 a_156122_n20028.n183 a_156122_n20028.n182 140.69
R36469 a_156122_n20028.n48 a_156122_n20028.n157 256.962
R36470 a_156122_n20028.n165 a_156122_n20028.n157 140.69
R36471 a_156122_n20028.n166 a_156122_n20028.n165 140.69
R36472 a_156122_n20028.n170 a_156122_n20028.n166 140.69
R36473 a_156122_n20028.n170 a_156122_n20028.n169 140.69
R36474 a_156122_n20028.n116 a_156122_n20028.n43 256.962
R36475 a_156122_n20028.n117 a_156122_n20028.n116 140.69
R36476 a_156122_n20028.n125 a_156122_n20028.n117 140.69
R36477 a_156122_n20028.n125 a_156122_n20028.n124 140.69
R36478 a_156122_n20028.n124 a_156122_n20028.n118 140.69
R36479 a_156122_n20028.n96 a_156122_n20028.t27 70.3453
R36480 a_156122_n20028.n182 a_156122_n20028.t21 70.3453
R36481 a_156122_n20028.n169 a_156122_n20028.t0 70.3453
R36482 a_156122_n20028.t20 a_156122_n20028.n118 70.3453
R36483 a_156122_n20028.n97 a_156122_n20028.n95 28.4333
R36484 a_156122_n20028.n181 a_156122_n20028.n180 28.4333
R36485 a_156122_n20028.n168 a_156122_n20028.n167 28.4333
R36486 a_156122_n20028.n120 a_156122_n20028.n119 28.4333
R36487 a_156122_n20028.n15 a_156122_n20028.n14 3.21237
R36488 a_156122_n20028.n98 a_156122_n20028.n94 24.8476
R36489 a_156122_n20028.n184 a_156122_n20028.n178 24.8476
R36490 a_156122_n20028.n171 a_156122_n20028.n156 24.8476
R36491 a_156122_n20028.n123 a_156122_n20028.n122 24.8476
R36492 a_156122_n20028.n101 a_156122_n20028.n100 23.3417
R36493 a_156122_n20028.n185 a_156122_n20028.n176 23.3417
R36494 a_156122_n20028.n172 a_156122_n20028.n155 23.3417
R36495 a_156122_n20028.n126 a_156122_n20028.n111 23.3417
R36496 a_156122_n20028.n15 a_156122_n20028.n75 27.6334
R36497 a_156122_n20028.n17 a_156122_n20028.n81 27.6334
R36498 a_156122_n20028.n19 a_156122_n20028.n87 27.6334
R36499 a_156122_n20028.n104 a_156122_n20028.n92 21.8358
R36500 a_156122_n20028.n189 a_156122_n20028.n188 21.8358
R36501 a_156122_n20028.n164 a_156122_n20028.n163 21.8358
R36502 a_156122_n20028.n127 a_156122_n20028.n110 21.8358
R36503 a_156122_n20028.n75 a_156122_n20028.n72 20.3299
R36504 a_156122_n20028.n81 a_156122_n20028.n78 20.3299
R36505 a_156122_n20028.n87 a_156122_n20028.n84 20.3299
R36506 a_156122_n20028.n105 a_156122_n20028.n91 20.3299
R36507 a_156122_n20028.n191 a_156122_n20028.n190 20.3299
R36508 a_156122_n20028.n162 a_156122_n20028.n158 20.3299
R36509 a_156122_n20028.n153 a_156122_n20028.n149 20.3299
R36510 a_156122_n20028.n147 a_156122_n20028.n143 20.3299
R36511 a_156122_n20028.n141 a_156122_n20028.n137 20.3299
R36512 a_156122_n20028.n115 a_156122_n20028.n114 20.3299
R36513 a_156122_n20028.n73 a_156122_n20028.n23 24.4363
R36514 a_156122_n20028.n79 a_156122_n20028.n25 24.4363
R36515 a_156122_n20028.n85 a_156122_n20028.n27 24.4363
R36516 a_156122_n20028.n29 a_156122_n20028.n108 22.9459
R36517 a_156122_n20028.n30 a_156122_n20028.n31 9.72532
R36518 a_156122_n20028.n32 a_156122_n20028.n33 9.72532
R36519 a_156122_n20028.n34 a_156122_n20028.n35 9.72532
R36520 a_156122_n20028.n36 a_156122_n20028.n37 9.72532
R36521 a_156122_n20028.n38 a_156122_n20028.n39 9.72532
R36522 a_156122_n20028.n23 a_156122_n20028.n22 9.72509
R36523 a_156122_n20028.n25 a_156122_n20028.n24 9.72509
R36524 a_156122_n20028.n27 a_156122_n20028.n26 9.72509
R36525 a_156122_n20028.n29 a_156122_n20028.n28 11.3106
R36526 a_156122_n20028.n41 a_156122_n20028.n40 11.3108
R36527 a_156122_n20028.n48 a_156122_n20028.n47 11.3109
R36528 a_156122_n20028.n49 a_156122_n20028.n50 9.72555
R36529 a_156122_n20028.n51 a_156122_n20028.n52 9.72555
R36530 a_156122_n20028.n53 a_156122_n20028.n54 9.72555
R36531 a_156122_n20028.n42 a_156122_n20028.n43 11.3108
R36532 a_156122_n20028.n46 a_156122_n20028.n45 9.72532
R36533 a_156122_n20028.n17 a_156122_n20028.n16 3.21237
R36534 a_156122_n20028.n19 a_156122_n20028.n18 3.21237
R36535 a_156122_n20028.n8 a_156122_n20028.n9 3.21131
R36536 a_156122_n20028.n10 a_156122_n20028.n11 3.21131
R36537 a_156122_n20028.n12 a_156122_n20028.n13 3.21131
R36538 a_156122_n20028.n55 a_156122_n20028.n56 2.85029
R36539 a_156122_n20028.n57 a_156122_n20028.n58 2.85029
R36540 a_156122_n20028.n59 a_156122_n20028.n60 2.85029
R36541 a_156122_n20028.n61 a_156122_n20028.n62 2.85029
R36542 a_156122_n20028.n63 a_156122_n20028.n64 2.85029
R36543 a_156122_n20028.n68 a_156122_n20028.n7 2.85029
R36544 a_156122_n20028.n195 a_156122_n20028.n194 9.3005
R36545 a_156122_n20028.n198 a_156122_n20028.n197 9.3005
R36546 a_156122_n20028.n71 a_156122_n20028.n70 9.3005
R36547 a_156122_n20028.n131 a_156122_n20028.n130 9.3005
R36548 a_156122_n20028.n134 a_156122_n20028.n133 9.3005
R36549 a_156122_n20028.n76 a_156122_n20028.n75 9.3005
R36550 a_156122_n20028.n74 a_156122_n20028.n73 9.3005
R36551 a_156122_n20028.n82 a_156122_n20028.n81 9.3005
R36552 a_156122_n20028.n80 a_156122_n20028.n79 9.3005
R36553 a_156122_n20028.n88 a_156122_n20028.n87 9.3005
R36554 a_156122_n20028.n86 a_156122_n20028.n85 9.3005
R36555 a_156122_n20028.n99 a_156122_n20028.n98 9.3005
R36556 a_156122_n20028.n92 a_156122_n20028.n3 9.3005
R36557 a_156122_n20028.n106 a_156122_n20028.n105 9.3005
R36558 a_156122_n20028.n108 a_156122_n20028.n107 9.3005
R36559 a_156122_n20028.n100 a_156122_n20028.n3 9.3005
R36560 a_156122_n20028.n178 a_156122_n20028.n177 9.3005
R36561 a_156122_n20028.n186 a_156122_n20028.n185 9.3005
R36562 a_156122_n20028.n188 a_156122_n20028.n187 9.3005
R36563 a_156122_n20028.n190 a_156122_n20028.n66 9.3005
R36564 a_156122_n20028.n174 a_156122_n20028.n65 9.3005
R36565 a_156122_n20028.n156 a_156122_n20028.n154 9.3005
R36566 a_156122_n20028.n2 a_156122_n20028.n172 9.3005
R36567 a_156122_n20028.n163 a_156122_n20028.n2 9.3005
R36568 a_156122_n20028.n162 a_156122_n20028.n161 9.3005
R36569 a_156122_n20028.n160 a_156122_n20028.n159 9.3005
R36570 a_156122_n20028.n153 a_156122_n20028.n152 9.3005
R36571 a_156122_n20028.n151 a_156122_n20028.n150 9.3005
R36572 a_156122_n20028.n147 a_156122_n20028.n146 9.3005
R36573 a_156122_n20028.n145 a_156122_n20028.n144 9.3005
R36574 a_156122_n20028.n141 a_156122_n20028.n140 9.3005
R36575 a_156122_n20028.n139 a_156122_n20028.n138 9.3005
R36576 a_156122_n20028.n122 a_156122_n20028.n121 9.3005
R36577 a_156122_n20028.n111 a_156122_n20028.n109 9.3005
R36578 a_156122_n20028.n128 a_156122_n20028.n127 9.3005
R36579 a_156122_n20028.n114 a_156122_n20028.n67 9.3005
R36580 a_156122_n20028.n113 a_156122_n20028.n112 9.3005
R36581 a_156122_n20028.n199 a_156122_n20028.n44 9.3005
R36582 a_156122_n20028.n31 a_156122_n20028.n195 24.4362
R36583 a_156122_n20028.n33 a_156122_n20028.n198 24.4362
R36584 a_156122_n20028.n35 a_156122_n20028.n71 24.4362
R36585 a_156122_n20028.n37 a_156122_n20028.n131 24.4362
R36586 a_156122_n20028.n39 a_156122_n20028.n134 24.4362
R36587 a_156122_n20028.n40 a_156122_n20028.n174 22.9458
R36588 a_156122_n20028.n159 a_156122_n20028.n48 22.9457
R36589 a_156122_n20028.n150 a_156122_n20028.n50 24.4361
R36590 a_156122_n20028.n144 a_156122_n20028.n52 24.4361
R36591 a_156122_n20028.n138 a_156122_n20028.n54 24.4361
R36592 a_156122_n20028.n43 a_156122_n20028.n113 22.9458
R36593 a_156122_n20028.n45 a_156122_n20028.n44 24.4362
R36594 a_156122_n20028.n6 a_156122_n20028.n30 7.9105
R36595 a_156122_n20028.n6 a_156122_n20028.n32 7.9105
R36596 a_156122_n20028.n4 a_156122_n20028.n34 7.9105
R36597 a_156122_n20028.n5 a_156122_n20028.n36 7.9105
R36598 a_156122_n20028.n5 a_156122_n20028.n38 7.9105
R36599 a_156122_n20028.n1 a_156122_n20028.n14 7.9105
R36600 a_156122_n20028.n1 a_156122_n20028.n16 7.9105
R36601 a_156122_n20028.n1 a_156122_n20028.n18 7.9105
R36602 a_156122_n20028.n1 a_156122_n20028.n3 7.9105
R36603 a_156122_n20028.n1 a_156122_n20028.n28 7.9105
R36604 a_156122_n20028.n1 a_156122_n20028.n26 7.9105
R36605 a_156122_n20028.n1 a_156122_n20028.n24 7.9105
R36606 a_156122_n20028.n1 a_156122_n20028.n22 7.9105
R36607 a_156122_n20028.n0 a_156122_n20028.n47 7.9105
R36608 a_156122_n20028.n0 a_156122_n20028.n49 7.9105
R36609 a_156122_n20028.n0 a_156122_n20028.n51 7.9105
R36610 a_156122_n20028.n0 a_156122_n20028.n53 7.9105
R36611 a_156122_n20028.n0 a_156122_n20028.n12 7.9105
R36612 a_156122_n20028.n0 a_156122_n20028.n10 7.9105
R36613 a_156122_n20028.n0 a_156122_n20028.n8 7.9105
R36614 a_156122_n20028.n0 a_156122_n20028.n2 7.9105
R36615 a_156122_n20028.n5 a_156122_n20028.n63 7.9105
R36616 a_156122_n20028.n5 a_156122_n20028.n61 7.9105
R36617 a_156122_n20028.n4 a_156122_n20028.n59 7.9105
R36618 a_156122_n20028.n6 a_156122_n20028.n57 7.9105
R36619 a_156122_n20028.n6 a_156122_n20028.n55 7.9105
R36620 a_156122_n20028.n46 a_156122_n20028.n4 7.9105
R36621 a_156122_n20028.n4 a_156122_n20028.n7 7.9105
R36622 a_156122_n20028.n56 a_156122_n20028.n195 28.3048
R36623 a_156122_n20028.n58 a_156122_n20028.n198 28.3048
R36624 a_156122_n20028.n60 a_156122_n20028.n71 28.3048
R36625 a_156122_n20028.n62 a_156122_n20028.n131 28.3048
R36626 a_156122_n20028.n64 a_156122_n20028.n134 28.3048
R36627 a_156122_n20028.n73 a_156122_n20028.n72 6.77697
R36628 a_156122_n20028.n79 a_156122_n20028.n78 6.77697
R36629 a_156122_n20028.n85 a_156122_n20028.n84 6.77697
R36630 a_156122_n20028.n108 a_156122_n20028.n91 6.77697
R36631 a_156122_n20028.n191 a_156122_n20028.n174 6.77697
R36632 a_156122_n20028.n159 a_156122_n20028.n158 6.77697
R36633 a_156122_n20028.n150 a_156122_n20028.n149 6.77697
R36634 a_156122_n20028.n144 a_156122_n20028.n143 6.77697
R36635 a_156122_n20028.n138 a_156122_n20028.n137 6.77697
R36636 a_156122_n20028.n115 a_156122_n20028.n113 6.77697
R36637 a_156122_n20028.n44 a_156122_n20028.n68 28.3048
R36638 a_156122_n20028.n99 a_156122_n20028.n95 5.33935
R36639 a_156122_n20028.n180 a_156122_n20028.n177 5.33935
R36640 a_156122_n20028.n167 a_156122_n20028.n154 5.33935
R36641 a_156122_n20028.n121 a_156122_n20028.n120 5.33935
R36642 a_156122_n20028.n105 a_156122_n20028.n104 5.27109
R36643 a_156122_n20028.n190 a_156122_n20028.n189 5.27109
R36644 a_156122_n20028.n164 a_156122_n20028.n162 5.27109
R36645 a_156122_n20028.n9 a_156122_n20028.n153 27.6341
R36646 a_156122_n20028.n11 a_156122_n20028.n147 27.6341
R36647 a_156122_n20028.n13 a_156122_n20028.n141 27.6341
R36648 a_156122_n20028.n114 a_156122_n20028.n110 5.27109
R36649 a_156122_n20028.n20 a_156122_n20028.n66 4.56989
R36650 a_156122_n20028.n21 a_156122_n20028.n67 4.56989
R36651 a_156122_n20028.n20 a_156122_n20028.n41 4.5005
R36652 a_156122_n20028.n21 a_156122_n20028.n42 4.5005
R36653 a_156122_n20028.n101 a_156122_n20028.n92 3.76521
R36654 a_156122_n20028.n188 a_156122_n20028.n176 3.76521
R36655 a_156122_n20028.n163 a_156122_n20028.n155 3.76521
R36656 a_156122_n20028.n127 a_156122_n20028.n126 3.76521
R36657 a_156122_n20028.n193 a_156122_n20028.t14 3.4805
R36658 a_156122_n20028.n193 a_156122_n20028.t13 3.4805
R36659 a_156122_n20028.n196 a_156122_n20028.t15 3.4805
R36660 a_156122_n20028.n196 a_156122_n20028.t19 3.4805
R36661 a_156122_n20028.n69 a_156122_n20028.t22 3.4805
R36662 a_156122_n20028.n69 a_156122_n20028.t10 3.4805
R36663 a_156122_n20028.n129 a_156122_n20028.t12 3.4805
R36664 a_156122_n20028.n129 a_156122_n20028.t11 3.4805
R36665 a_156122_n20028.n132 a_156122_n20028.t18 3.4805
R36666 a_156122_n20028.n132 a_156122_n20028.t16 3.4805
R36667 a_156122_n20028.n77 a_156122_n20028.t1 3.4805
R36668 a_156122_n20028.n77 a_156122_n20028.t7 3.4805
R36669 a_156122_n20028.n83 a_156122_n20028.t9 3.4805
R36670 a_156122_n20028.n83 a_156122_n20028.t2 3.4805
R36671 a_156122_n20028.n89 a_156122_n20028.t24 3.4805
R36672 a_156122_n20028.n89 a_156122_n20028.t4 3.4805
R36673 a_156122_n20028.n148 a_156122_n20028.t5 3.4805
R36674 a_156122_n20028.n148 a_156122_n20028.t25 3.4805
R36675 a_156122_n20028.n142 a_156122_n20028.t26 3.4805
R36676 a_156122_n20028.n142 a_156122_n20028.t3 3.4805
R36677 a_156122_n20028.n136 a_156122_n20028.t6 3.4805
R36678 a_156122_n20028.n136 a_156122_n20028.t8 3.4805
R36679 a_156122_n20028.t23 a_156122_n20028.n200 3.4805
R36680 a_156122_n20028.n200 a_156122_n20028.t17 3.4805
R36681 a_156122_n20028.n135 a_156122_n20028.n1 2.68111
R36682 a_156122_n20028.n173 a_156122_n20028.n1 2.5834
R36683 a_156122_n20028.n20 a_156122_n20028.n173 2.26061
R36684 a_156122_n20028.n135 a_156122_n20028.n21 2.26061
R36685 a_156122_n20028.n100 a_156122_n20028.n94 2.25932
R36686 a_156122_n20028.n185 a_156122_n20028.n184 2.25932
R36687 a_156122_n20028.n172 a_156122_n20028.n171 2.25932
R36688 a_156122_n20028.n123 a_156122_n20028.n111 2.25932
R36689 a_156122_n20028.n173 a_156122_n20028.n0 1.93434
R36690 a_156122_n20028.n0 a_156122_n20028.n135 1.83663
R36691 a_156122_n20028.n6 a_156122_n20028.n20 1.83146
R36692 a_156122_n20028.n21 a_156122_n20028.n5 1.82972
R36693 a_156122_n20028.n98 a_156122_n20028.n97 0.753441
R36694 a_156122_n20028.n181 a_156122_n20028.n178 0.753441
R36695 a_156122_n20028.n168 a_156122_n20028.n156 0.753441
R36696 a_156122_n20028.n122 a_156122_n20028.n119 0.753441
R36697 a_156122_n20028.n3 a_156122_n20028.n99 0.298809
R36698 a_156122_n20028.n2 a_156122_n20028.n154 0.298809
R36699 a_156122_n20028.n140 a_156122_n20028.n12 0.274655
R36700 a_156122_n20028.n146 a_156122_n20028.n10 0.274655
R36701 a_156122_n20028.n152 a_156122_n20028.n8 0.274655
R36702 a_156122_n20028.n5 a_156122_n20028.n4 0.270315
R36703 a_156122_n20028.n18 a_156122_n20028.n88 0.26922
R36704 a_156122_n20028.n16 a_156122_n20028.n82 0.26922
R36705 a_156122_n20028.n14 a_156122_n20028.n76 0.26922
R36706 a_156122_n20028.n107 a_156122_n20028.n28 0.231176
R36707 a_156122_n20028.n86 a_156122_n20028.n26 0.231176
R36708 a_156122_n20028.n80 a_156122_n20028.n24 0.231176
R36709 a_156122_n20028.n74 a_156122_n20028.n22 0.231176
R36710 a_156122_n20028.n199 a_156122_n20028.n46 0.228459
R36711 a_156122_n20028.n112 a_156122_n20028.n42 0.228459
R36712 a_156122_n20028.n41 a_156122_n20028.n65 0.228459
R36713 a_156122_n20028.n133 a_156122_n20028.n38 0.228459
R36714 a_156122_n20028.n130 a_156122_n20028.n36 0.228459
R36715 a_156122_n20028.n70 a_156122_n20028.n34 0.228459
R36716 a_156122_n20028.n197 a_156122_n20028.n32 0.228459
R36717 a_156122_n20028.n194 a_156122_n20028.n30 0.228459
R36718 a_156122_n20028.n139 a_156122_n20028.n53 0.225742
R36719 a_156122_n20028.n145 a_156122_n20028.n51 0.225742
R36720 a_156122_n20028.n151 a_156122_n20028.n49 0.225742
R36721 a_156122_n20028.n160 a_156122_n20028.n47 0.225742
R36722 a_156122_n20028.n76 a_156122_n20028.n74 0.196152
R36723 a_156122_n20028.n82 a_156122_n20028.n80 0.196152
R36724 a_156122_n20028.n88 a_156122_n20028.n86 0.196152
R36725 a_156122_n20028.n106 a_156122_n20028.n3 0.196152
R36726 a_156122_n20028.n107 a_156122_n20028.n106 0.196152
R36727 a_156122_n20028.n187 a_156122_n20028.n186 0.196152
R36728 a_156122_n20028.n186 a_156122_n20028.n177 0.196152
R36729 a_156122_n20028.n161 a_156122_n20028.n160 0.196152
R36730 a_156122_n20028.n161 a_156122_n20028.n2 0.196152
R36731 a_156122_n20028.n152 a_156122_n20028.n151 0.196152
R36732 a_156122_n20028.n146 a_156122_n20028.n145 0.196152
R36733 a_156122_n20028.n140 a_156122_n20028.n139 0.196152
R36734 a_156122_n20028.n128 a_156122_n20028.n109 0.196152
R36735 a_156122_n20028.n121 a_156122_n20028.n109 0.196152
R36736 a_156122_n20028.n4 a_156122_n20028.n6 0.179796
R36737 a_156122_n20028.n7 a_156122_n20028.n199 0.168676
R36738 a_156122_n20028.n133 a_156122_n20028.n63 0.168676
R36739 a_156122_n20028.n130 a_156122_n20028.n61 0.168676
R36740 a_156122_n20028.n70 a_156122_n20028.n59 0.168676
R36741 a_156122_n20028.n197 a_156122_n20028.n57 0.168676
R36742 a_156122_n20028.n194 a_156122_n20028.n55 0.168676
R36743 a_156122_n20028.n66 a_156122_n20028.n65 0.158954
R36744 a_156122_n20028.n112 a_156122_n20028.n67 0.158954
R36745 a_156122_n20028.n67 a_156122_n20028.n128 0.140355
R36746 a_156122_n20028.n187 a_156122_n20028.n66 0.140355
R36747 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t35 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n95 210.794
R36748 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t32 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n99 210.794
R36749 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n98 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t23 210.794
R36750 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t23 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n97 210.794
R36751 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t39 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n20 210.794
R36752 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n96 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t39 210.794
R36753 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n53 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t36 210.794
R36754 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t36 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n30 210.794
R36755 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n52 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t22 210.794
R36756 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t22 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n51 210.794
R36757 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t46 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n31 210.794
R36758 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n50 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t46 210.794
R36759 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t21 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n48 210.794
R36760 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n49 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t21 210.794
R36761 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n47 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t18 210.794
R36762 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t18 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n32 210.794
R36763 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n46 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t42 210.794
R36764 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t42 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n45 210.794
R36765 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t31 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n33 210.794
R36766 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n44 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t31 210.794
R36767 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t25 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n42 210.794
R36768 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n43 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t25 210.794
R36769 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n41 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t47 210.794
R36770 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t47 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n34 210.794
R36771 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n40 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t44 210.794
R36772 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t44 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n39 210.794
R36773 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t38 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n35 210.794
R36774 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n38 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t38 210.794
R36775 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n37 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t37 210.794
R36776 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t37 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n36 210.794
R36777 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t28 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n29 210.794
R36778 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n54 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t28 210.794
R36779 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n56 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t20 210.794
R36780 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t20 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n55 210.794
R36781 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n57 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t17 210.794
R36782 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t17 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n28 210.794
R36783 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t41 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n58 210.794
R36784 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n59 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t41 210.794
R36785 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t16 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n27 210.794
R36786 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n60 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t16 210.794
R36787 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n62 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t45 210.794
R36788 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t45 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n61 210.794
R36789 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n63 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t30 210.794
R36790 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t30 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n26 210.794
R36791 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t27 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n64 210.794
R36792 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n65 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t27 210.794
R36793 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t19 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n25 210.794
R36794 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n66 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t19 210.794
R36795 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n68 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t43 210.794
R36796 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t43 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n67 210.794
R36797 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n69 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t40 210.794
R36798 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t40 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n24 210.794
R36799 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t26 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n70 210.794
R36800 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n71 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t26 210.794
R36801 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t34 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n23 210.794
R36802 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n72 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t34 210.794
R36803 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n74 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t29 210.794
R36804 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t29 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n73 210.794
R36805 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n15 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n14 185
R36806 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n84 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n83 185
R36807 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t2 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n100 120.469
R36808 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n93 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t0 120.465
R36809 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n87 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t4 120.419
R36810 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t4 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n22 120.419
R36811 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n91 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t6 120.419
R36812 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t6 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n90 120.419
R36813 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n101 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t2 120.419
R36814 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n79 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t0 120.419
R36815 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n94 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t33 104.566
R36816 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n19 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t24 104.562
R36817 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n16 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n15 86.5152
R36818 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n83 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n82 86.5152
R36819 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n8 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n7 50.9993
R36820 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n78 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n77 47.5895
R36821 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n102 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n9 47.5893
R36822 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n89 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n88 38.0154
R36823 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n14 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n12 25.6005
R36824 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n84 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n81 25.6005
R36825 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n17 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n16 22.7786
R36826 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n82 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n21 22.7786
R36827 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t35 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n6 210.808
R36828 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n5 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n6 0.0650981
R36829 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n4 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n3 0.0650981
R36830 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n4 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t32 210.808
R36831 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n15 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t5 13.9205
R36832 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n15 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t3 13.9205
R36833 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n83 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t1 13.9205
R36834 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n83 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t7 13.9205
R36835 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n16 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n12 11.9727
R36836 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n82 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n81 11.9727
R36837 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n14 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n13 10.8064
R36838 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n85 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n84 10.8064
R36839 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n5 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n93 9.59564
R36840 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n100 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n3 9.59208
R36841 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n81 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n80 9.3005
R36842 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n12 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n11 9.3005
R36843 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n79 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n78 8.93258
R36844 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n102 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n101 8.84758
R36845 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n88 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t9 6.9605
R36846 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n88 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t8 6.9605
R36847 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n9 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t10 5.7135
R36848 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n9 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t14 5.7135
R36849 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n7 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t12 5.7135
R36850 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n7 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t11 5.7135
R36851 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n77 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t15 5.7135
R36852 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n77 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t13 5.7135
R36853 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n1 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n30 4.293
R36854 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n37 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n2 4.218
R36855 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n1 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n53 3.94612
R36856 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n36 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n2 3.87112
R36857 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n103 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n102 3.4105
R36858 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n78 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n76 3.4105
R36859 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n29 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n0 3.29712
R36860 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n54 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n1 3.29612
R36861 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n73 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n2 3.23112
R36862 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n75 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n74 3.23112
R36863 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n99 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n19 2.3168
R36864 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n103 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n0 2.31333
R36865 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n95 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n94 2.31188
R36866 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n76 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n75 2.30692
R36867 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n94 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n6 2.28563
R36868 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n97 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n96 0.645765
R36869 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n95 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n20 0.645765
R36870 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n98 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n20 0.645765
R36871 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n99 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n98 0.645765
R36872 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n91 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n22 0.645765
R36873 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n38 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n37 0.645765
R36874 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n39 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n38 0.645765
R36875 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n39 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n34 0.645765
R36876 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n43 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n34 0.645765
R36877 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n44 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n43 0.645765
R36878 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n45 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n44 0.645765
R36879 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n45 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n32 0.645765
R36880 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n49 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n32 0.645765
R36881 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n50 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n49 0.645765
R36882 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n51 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n50 0.645765
R36883 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n51 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n30 0.645765
R36884 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n36 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n35 0.645765
R36885 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n40 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n35 0.645765
R36886 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n41 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n40 0.645765
R36887 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n42 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n41 0.645765
R36888 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n42 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n33 0.645765
R36889 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n46 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n33 0.645765
R36890 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n47 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n46 0.645765
R36891 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n48 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n47 0.645765
R36892 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n48 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n31 0.645765
R36893 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n52 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n31 0.645765
R36894 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n53 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n52 0.645765
R36895 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n73 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n72 0.645765
R36896 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n72 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n71 0.645765
R36897 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n71 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n24 0.645765
R36898 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n67 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n24 0.645765
R36899 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n67 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n66 0.645765
R36900 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n66 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n65 0.645765
R36901 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n65 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n26 0.645765
R36902 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n61 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n26 0.645765
R36903 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n61 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n60 0.645765
R36904 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n60 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n59 0.645765
R36905 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n59 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n28 0.645765
R36906 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n55 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n28 0.645765
R36907 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n55 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n54 0.645765
R36908 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n74 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n23 0.645765
R36909 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n70 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n23 0.645765
R36910 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n70 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n69 0.645765
R36911 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n69 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n68 0.645765
R36912 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n68 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n25 0.645765
R36913 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n64 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n25 0.645765
R36914 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n64 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n63 0.645765
R36915 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n63 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n62 0.645765
R36916 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n62 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n27 0.645765
R36917 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n58 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n27 0.645765
R36918 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n58 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n57 0.645765
R36919 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n57 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n56 0.645765
R36920 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n56 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n29 0.645765
R36921 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n97 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n3 0.552061
R36922 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n96 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n5 0.550633
R36923 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n90 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n86 0.333133
R36924 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n92 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n91 0.333133
R36925 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n22 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n18 0.323133
R36926 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n87 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n10 0.323133
R36927 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n101 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n10 0.323133
R36928 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n86 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n79 0.313133
R36929 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n89 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n87 0.278133
R36930 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n90 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n89 0.268133
R36931 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n100 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n18 0.256274
R36932 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n93 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n92 0.252692
R36933 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n86 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n85 0.219522
R36934 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n18 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n17 0.217348
R36935 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n13 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n10 0.217348
R36936 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n92 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n21 0.216386
R36937 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n103 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n8 0.204167
R36938 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n76 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n8 0.204167
R36939 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n85 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n80 0.196152
R36940 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n80 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n21 0.196152
R36941 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n13 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n11 0.196152
R36942 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n17 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n11 0.196152
R36943 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n4 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n19 2.28913
R36944 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n75 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n2 0.4755
R36945 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n1 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n0 0.4755
R36946 a_187922_n20028.n31 a_187922_n20028.n196 91.4185
R36947 a_187922_n20028.n56 a_187922_n20028.n196 14.3253
R36948 a_187922_n20028.n33 a_187922_n20028.n69 91.4185
R36949 a_187922_n20028.n58 a_187922_n20028.n69 14.3253
R36950 a_187922_n20028.n35 a_187922_n20028.n129 91.4185
R36951 a_187922_n20028.n60 a_187922_n20028.n129 14.3253
R36952 a_187922_n20028.n37 a_187922_n20028.n132 91.4185
R36953 a_187922_n20028.n62 a_187922_n20028.n132 14.3253
R36954 a_187922_n20028.n39 a_187922_n20028.n135 91.4185
R36955 a_187922_n20028.n64 a_187922_n20028.n135 14.3253
R36956 a_187922_n20028.n77 a_187922_n20028.n15 15.3734
R36957 a_187922_n20028.n77 a_187922_n20028.n72 185
R36958 a_187922_n20028.n77 a_187922_n20028.n23 91.4184
R36959 a_187922_n20028.n83 a_187922_n20028.n17 15.3734
R36960 a_187922_n20028.n83 a_187922_n20028.n78 185
R36961 a_187922_n20028.n83 a_187922_n20028.n25 91.4184
R36962 a_187922_n20028.n89 a_187922_n20028.n19 15.3734
R36963 a_187922_n20028.n89 a_187922_n20028.n84 185
R36964 a_187922_n20028.n89 a_187922_n20028.n27 91.4184
R36965 a_187922_n20028.n97 a_187922_n20028.n96 185
R36966 a_187922_n20028.n94 a_187922_n20028.n93 185
R36967 a_187922_n20028.n102 a_187922_n20028.n101 185
R36968 a_187922_n20028.n104 a_187922_n20028.n103 185
R36969 a_187922_n20028.n91 a_187922_n20028.n90 185
R36970 a_187922_n20028.n195 a_187922_n20028.n194 185
R36971 a_187922_n20028.n192 a_187922_n20028.n178 185
R36972 a_187922_n20028.n182 a_187922_n20028.n179 185
R36973 a_187922_n20028.n187 a_187922_n20028.n186 185
R36974 a_187922_n20028.n185 a_187922_n20028.n184 185
R36975 a_187922_n20028.n161 a_187922_n20028.n160 185
R36976 a_187922_n20028.n168 a_187922_n20028.n167 185
R36977 a_187922_n20028.n169 a_187922_n20028.n158 185
R36978 a_187922_n20028.n174 a_187922_n20028.n173 185
R36979 a_187922_n20028.n172 a_187922_n20028.n171 185
R36980 a_187922_n20028.n50 a_187922_n20028.n151 91.4187
R36981 a_187922_n20028.n152 a_187922_n20028.n151 185
R36982 a_187922_n20028.n9 a_187922_n20028.n151 15.371
R36983 a_187922_n20028.n52 a_187922_n20028.n145 91.4187
R36984 a_187922_n20028.n146 a_187922_n20028.n145 185
R36985 a_187922_n20028.n11 a_187922_n20028.n145 15.371
R36986 a_187922_n20028.n54 a_187922_n20028.n139 91.4187
R36987 a_187922_n20028.n140 a_187922_n20028.n139 185
R36988 a_187922_n20028.n13 a_187922_n20028.n139 15.371
R36989 a_187922_n20028.n116 a_187922_n20028.n115 185
R36990 a_187922_n20028.n117 a_187922_n20028.n110 185
R36991 a_187922_n20028.n126 a_187922_n20028.n125 185
R36992 a_187922_n20028.n124 a_187922_n20028.n123 185
R36993 a_187922_n20028.n119 a_187922_n20028.n118 185
R36994 a_187922_n20028.n200 a_187922_n20028.n45 91.4185
R36995 a_187922_n20028.n200 a_187922_n20028.n68 14.3253
R36996 a_187922_n20028.t24 a_187922_n20028.n95 174.857
R36997 a_187922_n20028.n183 a_187922_n20028.t15 174.857
R36998 a_187922_n20028.n170 a_187922_n20028.t4 174.857
R36999 a_187922_n20028.n120 a_187922_n20028.t14 174.857
R37000 a_187922_n20028.n96 a_187922_n20028.n93 140.69
R37001 a_187922_n20028.n102 a_187922_n20028.n93 140.69
R37002 a_187922_n20028.n103 a_187922_n20028.n102 140.69
R37003 a_187922_n20028.n103 a_187922_n20028.n90 140.69
R37004 a_187922_n20028.n29 a_187922_n20028.n90 256.962
R37005 a_187922_n20028.n40 a_187922_n20028.n195 256.962
R37006 a_187922_n20028.n195 a_187922_n20028.n178 140.69
R37007 a_187922_n20028.n182 a_187922_n20028.n178 140.69
R37008 a_187922_n20028.n186 a_187922_n20028.n182 140.69
R37009 a_187922_n20028.n186 a_187922_n20028.n185 140.69
R37010 a_187922_n20028.n48 a_187922_n20028.n160 256.962
R37011 a_187922_n20028.n168 a_187922_n20028.n160 140.69
R37012 a_187922_n20028.n169 a_187922_n20028.n168 140.69
R37013 a_187922_n20028.n173 a_187922_n20028.n169 140.69
R37014 a_187922_n20028.n173 a_187922_n20028.n172 140.69
R37015 a_187922_n20028.n116 a_187922_n20028.n43 256.962
R37016 a_187922_n20028.n117 a_187922_n20028.n116 140.69
R37017 a_187922_n20028.n125 a_187922_n20028.n117 140.69
R37018 a_187922_n20028.n125 a_187922_n20028.n124 140.69
R37019 a_187922_n20028.n124 a_187922_n20028.n118 140.69
R37020 a_187922_n20028.n96 a_187922_n20028.t24 70.3453
R37021 a_187922_n20028.n185 a_187922_n20028.t15 70.3453
R37022 a_187922_n20028.n172 a_187922_n20028.t4 70.3453
R37023 a_187922_n20028.t14 a_187922_n20028.n118 70.3453
R37024 a_187922_n20028.n97 a_187922_n20028.n95 28.4333
R37025 a_187922_n20028.n184 a_187922_n20028.n183 28.4333
R37026 a_187922_n20028.n171 a_187922_n20028.n170 28.4333
R37027 a_187922_n20028.n120 a_187922_n20028.n119 28.4333
R37028 a_187922_n20028.n15 a_187922_n20028.n14 3.21237
R37029 a_187922_n20028.n98 a_187922_n20028.n94 24.8476
R37030 a_187922_n20028.n187 a_187922_n20028.n181 24.8476
R37031 a_187922_n20028.n174 a_187922_n20028.n159 24.8476
R37032 a_187922_n20028.n123 a_187922_n20028.n122 24.8476
R37033 a_187922_n20028.n101 a_187922_n20028.n100 23.3417
R37034 a_187922_n20028.n188 a_187922_n20028.n179 23.3417
R37035 a_187922_n20028.n175 a_187922_n20028.n158 23.3417
R37036 a_187922_n20028.n126 a_187922_n20028.n111 23.3417
R37037 a_187922_n20028.n15 a_187922_n20028.n75 27.6334
R37038 a_187922_n20028.n17 a_187922_n20028.n81 27.6334
R37039 a_187922_n20028.n19 a_187922_n20028.n87 27.6334
R37040 a_187922_n20028.n104 a_187922_n20028.n92 21.8358
R37041 a_187922_n20028.n192 a_187922_n20028.n191 21.8358
R37042 a_187922_n20028.n167 a_187922_n20028.n166 21.8358
R37043 a_187922_n20028.n127 a_187922_n20028.n110 21.8358
R37044 a_187922_n20028.n75 a_187922_n20028.n72 20.3299
R37045 a_187922_n20028.n81 a_187922_n20028.n78 20.3299
R37046 a_187922_n20028.n87 a_187922_n20028.n84 20.3299
R37047 a_187922_n20028.n105 a_187922_n20028.n91 20.3299
R37048 a_187922_n20028.n194 a_187922_n20028.n193 20.3299
R37049 a_187922_n20028.n165 a_187922_n20028.n161 20.3299
R37050 a_187922_n20028.n156 a_187922_n20028.n152 20.3299
R37051 a_187922_n20028.n150 a_187922_n20028.n146 20.3299
R37052 a_187922_n20028.n144 a_187922_n20028.n140 20.3299
R37053 a_187922_n20028.n115 a_187922_n20028.n114 20.3299
R37054 a_187922_n20028.n73 a_187922_n20028.n23 24.4363
R37055 a_187922_n20028.n79 a_187922_n20028.n25 24.4363
R37056 a_187922_n20028.n85 a_187922_n20028.n27 24.4363
R37057 a_187922_n20028.n29 a_187922_n20028.n108 22.9459
R37058 a_187922_n20028.n30 a_187922_n20028.n31 9.72532
R37059 a_187922_n20028.n32 a_187922_n20028.n33 9.72532
R37060 a_187922_n20028.n34 a_187922_n20028.n35 9.72532
R37061 a_187922_n20028.n36 a_187922_n20028.n37 9.72532
R37062 a_187922_n20028.n38 a_187922_n20028.n39 9.72532
R37063 a_187922_n20028.n23 a_187922_n20028.n22 9.72509
R37064 a_187922_n20028.n25 a_187922_n20028.n24 9.72509
R37065 a_187922_n20028.n27 a_187922_n20028.n26 9.72509
R37066 a_187922_n20028.n29 a_187922_n20028.n28 11.3106
R37067 a_187922_n20028.n41 a_187922_n20028.n40 11.3108
R37068 a_187922_n20028.n48 a_187922_n20028.n47 11.3109
R37069 a_187922_n20028.n49 a_187922_n20028.n50 9.72555
R37070 a_187922_n20028.n51 a_187922_n20028.n52 9.72555
R37071 a_187922_n20028.n53 a_187922_n20028.n54 9.72555
R37072 a_187922_n20028.n42 a_187922_n20028.n43 11.3108
R37073 a_187922_n20028.n46 a_187922_n20028.n45 9.72532
R37074 a_187922_n20028.n17 a_187922_n20028.n16 3.21237
R37075 a_187922_n20028.n19 a_187922_n20028.n18 3.21237
R37076 a_187922_n20028.n8 a_187922_n20028.n9 3.21131
R37077 a_187922_n20028.n10 a_187922_n20028.n11 3.21131
R37078 a_187922_n20028.n12 a_187922_n20028.n13 3.21131
R37079 a_187922_n20028.n55 a_187922_n20028.n56 2.85029
R37080 a_187922_n20028.n57 a_187922_n20028.n58 2.85029
R37081 a_187922_n20028.n59 a_187922_n20028.n60 2.85029
R37082 a_187922_n20028.n61 a_187922_n20028.n62 2.85029
R37083 a_187922_n20028.n63 a_187922_n20028.n64 2.85029
R37084 a_187922_n20028.n68 a_187922_n20028.n6 2.85029
R37085 a_187922_n20028.n198 a_187922_n20028.n197 9.3005
R37086 a_187922_n20028.n71 a_187922_n20028.n70 9.3005
R37087 a_187922_n20028.n131 a_187922_n20028.n130 9.3005
R37088 a_187922_n20028.n134 a_187922_n20028.n133 9.3005
R37089 a_187922_n20028.n137 a_187922_n20028.n136 9.3005
R37090 a_187922_n20028.n76 a_187922_n20028.n75 9.3005
R37091 a_187922_n20028.n74 a_187922_n20028.n73 9.3005
R37092 a_187922_n20028.n82 a_187922_n20028.n81 9.3005
R37093 a_187922_n20028.n80 a_187922_n20028.n79 9.3005
R37094 a_187922_n20028.n88 a_187922_n20028.n87 9.3005
R37095 a_187922_n20028.n86 a_187922_n20028.n85 9.3005
R37096 a_187922_n20028.n99 a_187922_n20028.n98 9.3005
R37097 a_187922_n20028.n92 a_187922_n20028.n3 9.3005
R37098 a_187922_n20028.n106 a_187922_n20028.n105 9.3005
R37099 a_187922_n20028.n108 a_187922_n20028.n107 9.3005
R37100 a_187922_n20028.n100 a_187922_n20028.n3 9.3005
R37101 a_187922_n20028.n181 a_187922_n20028.n180 9.3005
R37102 a_187922_n20028.n189 a_187922_n20028.n188 9.3005
R37103 a_187922_n20028.n191 a_187922_n20028.n190 9.3005
R37104 a_187922_n20028.n193 a_187922_n20028.n66 9.3005
R37105 a_187922_n20028.n177 a_187922_n20028.n65 9.3005
R37106 a_187922_n20028.n159 a_187922_n20028.n157 9.3005
R37107 a_187922_n20028.n2 a_187922_n20028.n175 9.3005
R37108 a_187922_n20028.n166 a_187922_n20028.n2 9.3005
R37109 a_187922_n20028.n165 a_187922_n20028.n164 9.3005
R37110 a_187922_n20028.n163 a_187922_n20028.n162 9.3005
R37111 a_187922_n20028.n156 a_187922_n20028.n155 9.3005
R37112 a_187922_n20028.n154 a_187922_n20028.n153 9.3005
R37113 a_187922_n20028.n150 a_187922_n20028.n149 9.3005
R37114 a_187922_n20028.n148 a_187922_n20028.n147 9.3005
R37115 a_187922_n20028.n144 a_187922_n20028.n143 9.3005
R37116 a_187922_n20028.n142 a_187922_n20028.n141 9.3005
R37117 a_187922_n20028.n122 a_187922_n20028.n121 9.3005
R37118 a_187922_n20028.n111 a_187922_n20028.n109 9.3005
R37119 a_187922_n20028.n128 a_187922_n20028.n127 9.3005
R37120 a_187922_n20028.n114 a_187922_n20028.n67 9.3005
R37121 a_187922_n20028.n113 a_187922_n20028.n112 9.3005
R37122 a_187922_n20028.n199 a_187922_n20028.n44 9.3005
R37123 a_187922_n20028.n31 a_187922_n20028.n198 24.4362
R37124 a_187922_n20028.n33 a_187922_n20028.n71 24.4362
R37125 a_187922_n20028.n35 a_187922_n20028.n131 24.4362
R37126 a_187922_n20028.n37 a_187922_n20028.n134 24.4362
R37127 a_187922_n20028.n39 a_187922_n20028.n137 24.4362
R37128 a_187922_n20028.n40 a_187922_n20028.n177 22.9458
R37129 a_187922_n20028.n162 a_187922_n20028.n48 22.9457
R37130 a_187922_n20028.n153 a_187922_n20028.n50 24.4361
R37131 a_187922_n20028.n147 a_187922_n20028.n52 24.4361
R37132 a_187922_n20028.n141 a_187922_n20028.n54 24.4361
R37133 a_187922_n20028.n43 a_187922_n20028.n113 22.9458
R37134 a_187922_n20028.n45 a_187922_n20028.n44 24.4362
R37135 a_187922_n20028.n7 a_187922_n20028.n30 7.9105
R37136 a_187922_n20028.n4 a_187922_n20028.n32 7.9105
R37137 a_187922_n20028.n4 a_187922_n20028.n34 7.9105
R37138 a_187922_n20028.n5 a_187922_n20028.n36 7.9105
R37139 a_187922_n20028.n5 a_187922_n20028.n38 7.9105
R37140 a_187922_n20028.n1 a_187922_n20028.n14 7.9105
R37141 a_187922_n20028.n1 a_187922_n20028.n16 7.9105
R37142 a_187922_n20028.n1 a_187922_n20028.n18 7.9105
R37143 a_187922_n20028.n1 a_187922_n20028.n3 7.9105
R37144 a_187922_n20028.n1 a_187922_n20028.n28 7.9105
R37145 a_187922_n20028.n1 a_187922_n20028.n26 7.9105
R37146 a_187922_n20028.n1 a_187922_n20028.n24 7.9105
R37147 a_187922_n20028.n1 a_187922_n20028.n22 7.9105
R37148 a_187922_n20028.n0 a_187922_n20028.n47 7.9105
R37149 a_187922_n20028.n0 a_187922_n20028.n49 7.9105
R37150 a_187922_n20028.n0 a_187922_n20028.n51 7.9105
R37151 a_187922_n20028.n0 a_187922_n20028.n53 7.9105
R37152 a_187922_n20028.n0 a_187922_n20028.n12 7.9105
R37153 a_187922_n20028.n0 a_187922_n20028.n10 7.9105
R37154 a_187922_n20028.n0 a_187922_n20028.n8 7.9105
R37155 a_187922_n20028.n0 a_187922_n20028.n2 7.9105
R37156 a_187922_n20028.n5 a_187922_n20028.n63 7.9105
R37157 a_187922_n20028.n5 a_187922_n20028.n61 7.9105
R37158 a_187922_n20028.n4 a_187922_n20028.n59 7.9105
R37159 a_187922_n20028.n4 a_187922_n20028.n57 7.9105
R37160 a_187922_n20028.n7 a_187922_n20028.n55 7.9105
R37161 a_187922_n20028.n46 a_187922_n20028.n7 7.9105
R37162 a_187922_n20028.n7 a_187922_n20028.n6 7.9105
R37163 a_187922_n20028.n56 a_187922_n20028.n198 28.3048
R37164 a_187922_n20028.n58 a_187922_n20028.n71 28.3048
R37165 a_187922_n20028.n60 a_187922_n20028.n131 28.3048
R37166 a_187922_n20028.n62 a_187922_n20028.n134 28.3048
R37167 a_187922_n20028.n64 a_187922_n20028.n137 28.3048
R37168 a_187922_n20028.n73 a_187922_n20028.n72 6.77697
R37169 a_187922_n20028.n79 a_187922_n20028.n78 6.77697
R37170 a_187922_n20028.n85 a_187922_n20028.n84 6.77697
R37171 a_187922_n20028.n108 a_187922_n20028.n91 6.77697
R37172 a_187922_n20028.n194 a_187922_n20028.n177 6.77697
R37173 a_187922_n20028.n162 a_187922_n20028.n161 6.77697
R37174 a_187922_n20028.n153 a_187922_n20028.n152 6.77697
R37175 a_187922_n20028.n147 a_187922_n20028.n146 6.77697
R37176 a_187922_n20028.n141 a_187922_n20028.n140 6.77697
R37177 a_187922_n20028.n115 a_187922_n20028.n113 6.77697
R37178 a_187922_n20028.n44 a_187922_n20028.n68 28.3048
R37179 a_187922_n20028.n99 a_187922_n20028.n95 5.33935
R37180 a_187922_n20028.n183 a_187922_n20028.n180 5.33935
R37181 a_187922_n20028.n170 a_187922_n20028.n157 5.33935
R37182 a_187922_n20028.n121 a_187922_n20028.n120 5.33935
R37183 a_187922_n20028.n105 a_187922_n20028.n104 5.27109
R37184 a_187922_n20028.n193 a_187922_n20028.n192 5.27109
R37185 a_187922_n20028.n167 a_187922_n20028.n165 5.27109
R37186 a_187922_n20028.n9 a_187922_n20028.n156 27.6341
R37187 a_187922_n20028.n11 a_187922_n20028.n150 27.6341
R37188 a_187922_n20028.n13 a_187922_n20028.n144 27.6341
R37189 a_187922_n20028.n114 a_187922_n20028.n110 5.27109
R37190 a_187922_n20028.n20 a_187922_n20028.n66 4.56989
R37191 a_187922_n20028.n21 a_187922_n20028.n67 4.56989
R37192 a_187922_n20028.n20 a_187922_n20028.n41 4.5005
R37193 a_187922_n20028.n21 a_187922_n20028.n42 4.5005
R37194 a_187922_n20028.n101 a_187922_n20028.n92 3.76521
R37195 a_187922_n20028.n191 a_187922_n20028.n179 3.76521
R37196 a_187922_n20028.n166 a_187922_n20028.n158 3.76521
R37197 a_187922_n20028.n127 a_187922_n20028.n126 3.76521
R37198 a_187922_n20028.n196 a_187922_n20028.t20 3.4805
R37199 a_187922_n20028.n196 a_187922_n20028.t18 3.4805
R37200 a_187922_n20028.n69 a_187922_n20028.t13 3.4805
R37201 a_187922_n20028.n69 a_187922_n20028.t8 3.4805
R37202 a_187922_n20028.n129 a_187922_n20028.t19 3.4805
R37203 a_187922_n20028.n129 a_187922_n20028.t16 3.4805
R37204 a_187922_n20028.n132 a_187922_n20028.t11 3.4805
R37205 a_187922_n20028.n132 a_187922_n20028.t9 3.4805
R37206 a_187922_n20028.n135 a_187922_n20028.t12 3.4805
R37207 a_187922_n20028.n135 a_187922_n20028.t17 3.4805
R37208 a_187922_n20028.n77 a_187922_n20028.t26 3.4805
R37209 a_187922_n20028.n77 a_187922_n20028.t5 3.4805
R37210 a_187922_n20028.n83 a_187922_n20028.t3 3.4805
R37211 a_187922_n20028.n83 a_187922_n20028.t6 3.4805
R37212 a_187922_n20028.n89 a_187922_n20028.t25 3.4805
R37213 a_187922_n20028.n89 a_187922_n20028.t23 3.4805
R37214 a_187922_n20028.n151 a_187922_n20028.t0 3.4805
R37215 a_187922_n20028.n151 a_187922_n20028.t27 3.4805
R37216 a_187922_n20028.n145 a_187922_n20028.t22 3.4805
R37217 a_187922_n20028.n145 a_187922_n20028.t7 3.4805
R37218 a_187922_n20028.n139 a_187922_n20028.t2 3.4805
R37219 a_187922_n20028.n139 a_187922_n20028.t1 3.4805
R37220 a_187922_n20028.t21 a_187922_n20028.n200 3.4805
R37221 a_187922_n20028.n200 a_187922_n20028.t10 3.4805
R37222 a_187922_n20028.n138 a_187922_n20028.n1 2.68111
R37223 a_187922_n20028.n176 a_187922_n20028.n1 2.5834
R37224 a_187922_n20028.n20 a_187922_n20028.n176 2.26061
R37225 a_187922_n20028.n138 a_187922_n20028.n21 2.26061
R37226 a_187922_n20028.n100 a_187922_n20028.n94 2.25932
R37227 a_187922_n20028.n188 a_187922_n20028.n187 2.25932
R37228 a_187922_n20028.n175 a_187922_n20028.n174 2.25932
R37229 a_187922_n20028.n123 a_187922_n20028.n111 2.25932
R37230 a_187922_n20028.n176 a_187922_n20028.n0 1.93434
R37231 a_187922_n20028.n0 a_187922_n20028.n138 1.83663
R37232 a_187922_n20028.n7 a_187922_n20028.n20 1.83146
R37233 a_187922_n20028.n21 a_187922_n20028.n5 1.82972
R37234 a_187922_n20028.n98 a_187922_n20028.n97 0.753441
R37235 a_187922_n20028.n184 a_187922_n20028.n181 0.753441
R37236 a_187922_n20028.n171 a_187922_n20028.n159 0.753441
R37237 a_187922_n20028.n122 a_187922_n20028.n119 0.753441
R37238 a_187922_n20028.n3 a_187922_n20028.n99 0.298809
R37239 a_187922_n20028.n2 a_187922_n20028.n157 0.298809
R37240 a_187922_n20028.n143 a_187922_n20028.n12 0.274655
R37241 a_187922_n20028.n149 a_187922_n20028.n10 0.274655
R37242 a_187922_n20028.n155 a_187922_n20028.n8 0.274655
R37243 a_187922_n20028.n5 a_187922_n20028.n4 0.270315
R37244 a_187922_n20028.n18 a_187922_n20028.n88 0.26922
R37245 a_187922_n20028.n16 a_187922_n20028.n82 0.26922
R37246 a_187922_n20028.n14 a_187922_n20028.n76 0.26922
R37247 a_187922_n20028.n107 a_187922_n20028.n28 0.231176
R37248 a_187922_n20028.n86 a_187922_n20028.n26 0.231176
R37249 a_187922_n20028.n80 a_187922_n20028.n24 0.231176
R37250 a_187922_n20028.n74 a_187922_n20028.n22 0.231176
R37251 a_187922_n20028.n199 a_187922_n20028.n46 0.228459
R37252 a_187922_n20028.n112 a_187922_n20028.n42 0.228459
R37253 a_187922_n20028.n41 a_187922_n20028.n65 0.228459
R37254 a_187922_n20028.n136 a_187922_n20028.n38 0.228459
R37255 a_187922_n20028.n133 a_187922_n20028.n36 0.228459
R37256 a_187922_n20028.n130 a_187922_n20028.n34 0.228459
R37257 a_187922_n20028.n70 a_187922_n20028.n32 0.228459
R37258 a_187922_n20028.n197 a_187922_n20028.n30 0.228459
R37259 a_187922_n20028.n142 a_187922_n20028.n53 0.225742
R37260 a_187922_n20028.n148 a_187922_n20028.n51 0.225742
R37261 a_187922_n20028.n154 a_187922_n20028.n49 0.225742
R37262 a_187922_n20028.n163 a_187922_n20028.n47 0.225742
R37263 a_187922_n20028.n76 a_187922_n20028.n74 0.196152
R37264 a_187922_n20028.n82 a_187922_n20028.n80 0.196152
R37265 a_187922_n20028.n88 a_187922_n20028.n86 0.196152
R37266 a_187922_n20028.n106 a_187922_n20028.n3 0.196152
R37267 a_187922_n20028.n107 a_187922_n20028.n106 0.196152
R37268 a_187922_n20028.n190 a_187922_n20028.n189 0.196152
R37269 a_187922_n20028.n189 a_187922_n20028.n180 0.196152
R37270 a_187922_n20028.n164 a_187922_n20028.n163 0.196152
R37271 a_187922_n20028.n164 a_187922_n20028.n2 0.196152
R37272 a_187922_n20028.n155 a_187922_n20028.n154 0.196152
R37273 a_187922_n20028.n149 a_187922_n20028.n148 0.196152
R37274 a_187922_n20028.n143 a_187922_n20028.n142 0.196152
R37275 a_187922_n20028.n128 a_187922_n20028.n109 0.196152
R37276 a_187922_n20028.n121 a_187922_n20028.n109 0.196152
R37277 a_187922_n20028.n7 a_187922_n20028.n4 0.179796
R37278 a_187922_n20028.n6 a_187922_n20028.n199 0.168676
R37279 a_187922_n20028.n136 a_187922_n20028.n63 0.168676
R37280 a_187922_n20028.n133 a_187922_n20028.n61 0.168676
R37281 a_187922_n20028.n130 a_187922_n20028.n59 0.168676
R37282 a_187922_n20028.n70 a_187922_n20028.n57 0.168676
R37283 a_187922_n20028.n197 a_187922_n20028.n55 0.168676
R37284 a_187922_n20028.n66 a_187922_n20028.n65 0.158954
R37285 a_187922_n20028.n112 a_187922_n20028.n67 0.158954
R37286 a_187922_n20028.n67 a_187922_n20028.n128 0.140355
R37287 a_187922_n20028.n190 a_187922_n20028.n66 0.140355
R37288 C2S2_Amp_F_I_1.OUT.n72 C2S2_Amp_F_I_1.OUT.n66 585
R37289 C2S2_Amp_F_I_1.OUT.n72 C2S2_Amp_F_I_1.OUT.n65 585
R37290 C2S2_Amp_F_I_1.OUT.n73 C2S2_Amp_F_I_1.OUT.n72 585
R37291 C2S2_Amp_F_I_1.OUT.n85 C2S2_Amp_F_I_1.OUT.n79 585
R37292 C2S2_Amp_F_I_1.OUT.n85 C2S2_Amp_F_I_1.OUT.n78 585
R37293 C2S2_Amp_F_I_1.OUT.n86 C2S2_Amp_F_I_1.OUT.n85 585
R37294 C2S2_Amp_F_I_1.OUT.n98 C2S2_Amp_F_I_1.OUT.n92 585
R37295 C2S2_Amp_F_I_1.OUT.n98 C2S2_Amp_F_I_1.OUT.n91 585
R37296 C2S2_Amp_F_I_1.OUT.n99 C2S2_Amp_F_I_1.OUT.n98 585
R37297 C2S2_Amp_F_I_1.OUT.n111 C2S2_Amp_F_I_1.OUT.n105 585
R37298 C2S2_Amp_F_I_1.OUT.n111 C2S2_Amp_F_I_1.OUT.n104 585
R37299 C2S2_Amp_F_I_1.OUT.n112 C2S2_Amp_F_I_1.OUT.n111 585
R37300 C2S2_Amp_F_I_1.OUT.n124 C2S2_Amp_F_I_1.OUT.n118 585
R37301 C2S2_Amp_F_I_1.OUT.n124 C2S2_Amp_F_I_1.OUT.n117 585
R37302 C2S2_Amp_F_I_1.OUT.n125 C2S2_Amp_F_I_1.OUT.n124 585
R37303 C2S2_Amp_F_I_1.OUT.n137 C2S2_Amp_F_I_1.OUT.n131 585
R37304 C2S2_Amp_F_I_1.OUT.n137 C2S2_Amp_F_I_1.OUT.n130 585
R37305 C2S2_Amp_F_I_1.OUT.n138 C2S2_Amp_F_I_1.OUT.n137 585
R37306 C2S2_Amp_F_I_1.OUT.n150 C2S2_Amp_F_I_1.OUT.n144 585
R37307 C2S2_Amp_F_I_1.OUT.n150 C2S2_Amp_F_I_1.OUT.n143 585
R37308 C2S2_Amp_F_I_1.OUT.n151 C2S2_Amp_F_I_1.OUT.n150 585
R37309 C2S2_Amp_F_I_1.OUT.n163 C2S2_Amp_F_I_1.OUT.n157 585
R37310 C2S2_Amp_F_I_1.OUT.n163 C2S2_Amp_F_I_1.OUT.n156 585
R37311 C2S2_Amp_F_I_1.OUT.n164 C2S2_Amp_F_I_1.OUT.n163 585
R37312 C2S2_Amp_F_I_1.OUT.n176 C2S2_Amp_F_I_1.OUT.n170 585
R37313 C2S2_Amp_F_I_1.OUT.n176 C2S2_Amp_F_I_1.OUT.n169 585
R37314 C2S2_Amp_F_I_1.OUT.n177 C2S2_Amp_F_I_1.OUT.n176 585
R37315 C2S2_Amp_F_I_1.OUT.n189 C2S2_Amp_F_I_1.OUT.n183 585
R37316 C2S2_Amp_F_I_1.OUT.n189 C2S2_Amp_F_I_1.OUT.n182 585
R37317 C2S2_Amp_F_I_1.OUT.n190 C2S2_Amp_F_I_1.OUT.n189 585
R37318 C2S2_Amp_F_I_1.OUT.n202 C2S2_Amp_F_I_1.OUT.n196 585
R37319 C2S2_Amp_F_I_1.OUT.n202 C2S2_Amp_F_I_1.OUT.n195 585
R37320 C2S2_Amp_F_I_1.OUT.n203 C2S2_Amp_F_I_1.OUT.n202 585
R37321 C2S2_Amp_F_I_1.OUT.n215 C2S2_Amp_F_I_1.OUT.n209 585
R37322 C2S2_Amp_F_I_1.OUT.n215 C2S2_Amp_F_I_1.OUT.n208 585
R37323 C2S2_Amp_F_I_1.OUT.n216 C2S2_Amp_F_I_1.OUT.n215 585
R37324 C2S2_Amp_F_I_1.OUT.n228 C2S2_Amp_F_I_1.OUT.n222 585
R37325 C2S2_Amp_F_I_1.OUT.n228 C2S2_Amp_F_I_1.OUT.n221 585
R37326 C2S2_Amp_F_I_1.OUT.n229 C2S2_Amp_F_I_1.OUT.n228 585
R37327 C2S2_Amp_F_I_1.OUT.n241 C2S2_Amp_F_I_1.OUT.n235 585
R37328 C2S2_Amp_F_I_1.OUT.n241 C2S2_Amp_F_I_1.OUT.n234 585
R37329 C2S2_Amp_F_I_1.OUT.n242 C2S2_Amp_F_I_1.OUT.n241 585
R37330 C2S2_Amp_F_I_1.OUT.n254 C2S2_Amp_F_I_1.OUT.n248 585
R37331 C2S2_Amp_F_I_1.OUT.n254 C2S2_Amp_F_I_1.OUT.n247 585
R37332 C2S2_Amp_F_I_1.OUT.n255 C2S2_Amp_F_I_1.OUT.n254 585
R37333 C2S2_Amp_F_I_1.OUT.n267 C2S2_Amp_F_I_1.OUT.n261 585
R37334 C2S2_Amp_F_I_1.OUT.n267 C2S2_Amp_F_I_1.OUT.n260 585
R37335 C2S2_Amp_F_I_1.OUT.n268 C2S2_Amp_F_I_1.OUT.n267 585
R37336 C2S2_Amp_F_I_1.OUT.n280 C2S2_Amp_F_I_1.OUT.n274 585
R37337 C2S2_Amp_F_I_1.OUT.n280 C2S2_Amp_F_I_1.OUT.n273 585
R37338 C2S2_Amp_F_I_1.OUT.n281 C2S2_Amp_F_I_1.OUT.n280 585
R37339 C2S2_Amp_F_I_1.OUT.n293 C2S2_Amp_F_I_1.OUT.n287 585
R37340 C2S2_Amp_F_I_1.OUT.n293 C2S2_Amp_F_I_1.OUT.n286 585
R37341 C2S2_Amp_F_I_1.OUT.n294 C2S2_Amp_F_I_1.OUT.n293 585
R37342 C2S2_Amp_F_I_1.OUT.n305 C2S2_Amp_F_I_1.OUT.n304 585
R37343 C2S2_Amp_F_I_1.OUT.n304 C2S2_Amp_F_I_1.OUT.n303 585
R37344 C2S2_Amp_F_I_1.OUT.n304 C2S2_Amp_F_I_1.OUT.n300 585
R37345 C2S2_Amp_F_I_1.OUT.n58 C2S2_Amp_F_I_1.OUT.n57 585
R37346 C2S2_Amp_F_I_1.OUT.n57 C2S2_Amp_F_I_1.OUT.n56 585
R37347 C2S2_Amp_F_I_1.OUT.n57 C2S2_Amp_F_I_1.OUT.n52 585
R37348 C2S2_Amp_F_I_1.OUT.n7 C2S2_Amp_F_I_1.OUT.n5 325.69
R37349 C2S2_Amp_F_I_1.OUT.n404 C2S2_Amp_F_I_1.OUT.n402 325.69
R37350 C2S2_Amp_F_I_1.OUT.n6 C2S2_Amp_F_I_1.OUT.n5 185
R37351 C2S2_Amp_F_I_1.OUT.n14 C2S2_Amp_F_I_1.OUT.n13 185
R37352 C2S2_Amp_F_I_1.OUT.n15 C2S2_Amp_F_I_1.OUT.n3 185
R37353 C2S2_Amp_F_I_1.OUT.n24 C2S2_Amp_F_I_1.OUT.n23 185
R37354 C2S2_Amp_F_I_1.OUT.n22 C2S2_Amp_F_I_1.OUT.n21 185
R37355 C2S2_Amp_F_I_1.OUT.n17 C2S2_Amp_F_I_1.OUT.n16 185
R37356 C2S2_Amp_F_I_1.OUT.n336 C2S2_Amp_F_I_1.OUT.n334 185
R37357 C2S2_Amp_F_I_1.OUT.n335 C2S2_Amp_F_I_1.OUT.n334 185
R37358 C2S2_Amp_F_I_1.OUT.n341 C2S2_Amp_F_I_1.OUT.n334 185
R37359 C2S2_Amp_F_I_1.OUT.n349 C2S2_Amp_F_I_1.OUT.n347 185
R37360 C2S2_Amp_F_I_1.OUT.n348 C2S2_Amp_F_I_1.OUT.n347 185
R37361 C2S2_Amp_F_I_1.OUT.n354 C2S2_Amp_F_I_1.OUT.n347 185
R37362 C2S2_Amp_F_I_1.OUT.n362 C2S2_Amp_F_I_1.OUT.n360 185
R37363 C2S2_Amp_F_I_1.OUT.n361 C2S2_Amp_F_I_1.OUT.n360 185
R37364 C2S2_Amp_F_I_1.OUT.n367 C2S2_Amp_F_I_1.OUT.n360 185
R37365 C2S2_Amp_F_I_1.OUT.n375 C2S2_Amp_F_I_1.OUT.n373 185
R37366 C2S2_Amp_F_I_1.OUT.n374 C2S2_Amp_F_I_1.OUT.n373 185
R37367 C2S2_Amp_F_I_1.OUT.n380 C2S2_Amp_F_I_1.OUT.n373 185
R37368 C2S2_Amp_F_I_1.OUT.n388 C2S2_Amp_F_I_1.OUT.n386 185
R37369 C2S2_Amp_F_I_1.OUT.n387 C2S2_Amp_F_I_1.OUT.n386 185
R37370 C2S2_Amp_F_I_1.OUT.n393 C2S2_Amp_F_I_1.OUT.n386 185
R37371 C2S2_Amp_F_I_1.OUT.n403 C2S2_Amp_F_I_1.OUT.n402 185
R37372 C2S2_Amp_F_I_1.OUT.n411 C2S2_Amp_F_I_1.OUT.n410 185
R37373 C2S2_Amp_F_I_1.OUT.n412 C2S2_Amp_F_I_1.OUT.n400 185
R37374 C2S2_Amp_F_I_1.OUT.n421 C2S2_Amp_F_I_1.OUT.n420 185
R37375 C2S2_Amp_F_I_1.OUT.n419 C2S2_Amp_F_I_1.OUT.n418 185
R37376 C2S2_Amp_F_I_1.OUT.n414 C2S2_Amp_F_I_1.OUT.n413 185
R37377 C2S2_Amp_F_I_1.OUT.n18 C2S2_Amp_F_I_1.OUT.t20 174.857
R37378 C2S2_Amp_F_I_1.OUT.n415 C2S2_Amp_F_I_1.OUT.t17 174.857
R37379 C2S2_Amp_F_I_1.OUT.n14 C2S2_Amp_F_I_1.OUT.n5 140.69
R37380 C2S2_Amp_F_I_1.OUT.n15 C2S2_Amp_F_I_1.OUT.n14 140.69
R37381 C2S2_Amp_F_I_1.OUT.n23 C2S2_Amp_F_I_1.OUT.n15 140.69
R37382 C2S2_Amp_F_I_1.OUT.n23 C2S2_Amp_F_I_1.OUT.n22 140.69
R37383 C2S2_Amp_F_I_1.OUT.n22 C2S2_Amp_F_I_1.OUT.n16 140.69
R37384 C2S2_Amp_F_I_1.OUT.n411 C2S2_Amp_F_I_1.OUT.n402 140.69
R37385 C2S2_Amp_F_I_1.OUT.n412 C2S2_Amp_F_I_1.OUT.n411 140.69
R37386 C2S2_Amp_F_I_1.OUT.n420 C2S2_Amp_F_I_1.OUT.n412 140.69
R37387 C2S2_Amp_F_I_1.OUT.n420 C2S2_Amp_F_I_1.OUT.n419 140.69
R37388 C2S2_Amp_F_I_1.OUT.n419 C2S2_Amp_F_I_1.OUT.n413 140.69
R37389 C2S2_Amp_F_I_1.OUT.t20 C2S2_Amp_F_I_1.OUT.n16 70.3453
R37390 C2S2_Amp_F_I_1.OUT.t17 C2S2_Amp_F_I_1.OUT.n413 70.3453
R37391 C2S2_Amp_F_I_1.OUT.n72 C2S2_Amp_F_I_1.OUT.n71 51.669
R37392 C2S2_Amp_F_I_1.OUT.n85 C2S2_Amp_F_I_1.OUT.n84 51.669
R37393 C2S2_Amp_F_I_1.OUT.n98 C2S2_Amp_F_I_1.OUT.n97 51.669
R37394 C2S2_Amp_F_I_1.OUT.n111 C2S2_Amp_F_I_1.OUT.n110 51.669
R37395 C2S2_Amp_F_I_1.OUT.n124 C2S2_Amp_F_I_1.OUT.n123 51.669
R37396 C2S2_Amp_F_I_1.OUT.n137 C2S2_Amp_F_I_1.OUT.n136 51.669
R37397 C2S2_Amp_F_I_1.OUT.n150 C2S2_Amp_F_I_1.OUT.n149 51.669
R37398 C2S2_Amp_F_I_1.OUT.n163 C2S2_Amp_F_I_1.OUT.n162 51.669
R37399 C2S2_Amp_F_I_1.OUT.n176 C2S2_Amp_F_I_1.OUT.n175 51.669
R37400 C2S2_Amp_F_I_1.OUT.n189 C2S2_Amp_F_I_1.OUT.n188 51.669
R37401 C2S2_Amp_F_I_1.OUT.n202 C2S2_Amp_F_I_1.OUT.n201 51.669
R37402 C2S2_Amp_F_I_1.OUT.n215 C2S2_Amp_F_I_1.OUT.n214 51.669
R37403 C2S2_Amp_F_I_1.OUT.n228 C2S2_Amp_F_I_1.OUT.n227 51.669
R37404 C2S2_Amp_F_I_1.OUT.n241 C2S2_Amp_F_I_1.OUT.n240 51.669
R37405 C2S2_Amp_F_I_1.OUT.n254 C2S2_Amp_F_I_1.OUT.n253 51.669
R37406 C2S2_Amp_F_I_1.OUT.n267 C2S2_Amp_F_I_1.OUT.n266 51.669
R37407 C2S2_Amp_F_I_1.OUT.n280 C2S2_Amp_F_I_1.OUT.n279 51.669
R37408 C2S2_Amp_F_I_1.OUT.n293 C2S2_Amp_F_I_1.OUT.n292 51.669
R37409 C2S2_Amp_F_I_1.OUT.n304 C2S2_Amp_F_I_1.OUT.n297 51.669
R37410 C2S2_Amp_F_I_1.OUT.n57 C2S2_Amp_F_I_1.OUT.n49 51.669
R37411 C2S2_Amp_F_I_1.OUT.n71 C2S2_Amp_F_I_1.OUT.n70 29.812
R37412 C2S2_Amp_F_I_1.OUT.n84 C2S2_Amp_F_I_1.OUT.n83 29.812
R37413 C2S2_Amp_F_I_1.OUT.n97 C2S2_Amp_F_I_1.OUT.n96 29.812
R37414 C2S2_Amp_F_I_1.OUT.n110 C2S2_Amp_F_I_1.OUT.n109 29.812
R37415 C2S2_Amp_F_I_1.OUT.n123 C2S2_Amp_F_I_1.OUT.n122 29.812
R37416 C2S2_Amp_F_I_1.OUT.n136 C2S2_Amp_F_I_1.OUT.n135 29.812
R37417 C2S2_Amp_F_I_1.OUT.n149 C2S2_Amp_F_I_1.OUT.n148 29.812
R37418 C2S2_Amp_F_I_1.OUT.n162 C2S2_Amp_F_I_1.OUT.n161 29.812
R37419 C2S2_Amp_F_I_1.OUT.n175 C2S2_Amp_F_I_1.OUT.n174 29.812
R37420 C2S2_Amp_F_I_1.OUT.n188 C2S2_Amp_F_I_1.OUT.n187 29.812
R37421 C2S2_Amp_F_I_1.OUT.n201 C2S2_Amp_F_I_1.OUT.n200 29.812
R37422 C2S2_Amp_F_I_1.OUT.n214 C2S2_Amp_F_I_1.OUT.n213 29.812
R37423 C2S2_Amp_F_I_1.OUT.n227 C2S2_Amp_F_I_1.OUT.n226 29.812
R37424 C2S2_Amp_F_I_1.OUT.n240 C2S2_Amp_F_I_1.OUT.n239 29.812
R37425 C2S2_Amp_F_I_1.OUT.n253 C2S2_Amp_F_I_1.OUT.n252 29.812
R37426 C2S2_Amp_F_I_1.OUT.n266 C2S2_Amp_F_I_1.OUT.n265 29.812
R37427 C2S2_Amp_F_I_1.OUT.n279 C2S2_Amp_F_I_1.OUT.n278 29.812
R37428 C2S2_Amp_F_I_1.OUT.n292 C2S2_Amp_F_I_1.OUT.n291 29.812
R37429 C2S2_Amp_F_I_1.OUT.n306 C2S2_Amp_F_I_1.OUT.n297 29.812
R37430 C2S2_Amp_F_I_1.OUT.n59 C2S2_Amp_F_I_1.OUT.n49 29.812
R37431 C2S2_Amp_F_I_1.OUT.n18 C2S2_Amp_F_I_1.OUT.n17 28.4333
R37432 C2S2_Amp_F_I_1.OUT.n415 C2S2_Amp_F_I_1.OUT.n414 28.4333
R37433 C2S2_Amp_F_I_1.OUT.n343 C2S2_Amp_F_I_1.OUT.n342 27.6063
R37434 C2S2_Amp_F_I_1.OUT.n356 C2S2_Amp_F_I_1.OUT.n355 27.6063
R37435 C2S2_Amp_F_I_1.OUT.n369 C2S2_Amp_F_I_1.OUT.n368 27.6063
R37436 C2S2_Amp_F_I_1.OUT.n382 C2S2_Amp_F_I_1.OUT.n381 27.6063
R37437 C2S2_Amp_F_I_1.OUT.n395 C2S2_Amp_F_I_1.OUT.n394 27.6063
R37438 C2S2_Amp_F_I_1.OUT.n21 C2S2_Amp_F_I_1.OUT.n20 24.8476
R37439 C2S2_Amp_F_I_1.OUT.n418 C2S2_Amp_F_I_1.OUT.n417 24.8476
R37440 C2S2_Amp_F_I_1.OUT.n24 C2S2_Amp_F_I_1.OUT.n4 23.3417
R37441 C2S2_Amp_F_I_1.OUT.n421 C2S2_Amp_F_I_1.OUT.n401 23.3417
R37442 C2S2_Amp_F_I_1.OUT.n25 C2S2_Amp_F_I_1.OUT.n3 21.8358
R37443 C2S2_Amp_F_I_1.OUT.n422 C2S2_Amp_F_I_1.OUT.n400 21.8358
R37444 C2S2_Amp_F_I_1.OUT.n13 C2S2_Amp_F_I_1.OUT.n12 20.3299
R37445 C2S2_Amp_F_I_1.OUT.n342 C2S2_Amp_F_I_1.OUT.n341 20.3299
R37446 C2S2_Amp_F_I_1.OUT.n355 C2S2_Amp_F_I_1.OUT.n354 20.3299
R37447 C2S2_Amp_F_I_1.OUT.n368 C2S2_Amp_F_I_1.OUT.n367 20.3299
R37448 C2S2_Amp_F_I_1.OUT.n381 C2S2_Amp_F_I_1.OUT.n380 20.3299
R37449 C2S2_Amp_F_I_1.OUT.n394 C2S2_Amp_F_I_1.OUT.n393 20.3299
R37450 C2S2_Amp_F_I_1.OUT.n410 C2S2_Amp_F_I_1.OUT.n409 20.3299
R37451 C2S2_Amp_F_I_1.OUT.n70 C2S2_Amp_F_I_1.OUT.n66 20.3299
R37452 C2S2_Amp_F_I_1.OUT.n83 C2S2_Amp_F_I_1.OUT.n79 20.3299
R37453 C2S2_Amp_F_I_1.OUT.n96 C2S2_Amp_F_I_1.OUT.n92 20.3299
R37454 C2S2_Amp_F_I_1.OUT.n109 C2S2_Amp_F_I_1.OUT.n105 20.3299
R37455 C2S2_Amp_F_I_1.OUT.n122 C2S2_Amp_F_I_1.OUT.n118 20.3299
R37456 C2S2_Amp_F_I_1.OUT.n135 C2S2_Amp_F_I_1.OUT.n131 20.3299
R37457 C2S2_Amp_F_I_1.OUT.n148 C2S2_Amp_F_I_1.OUT.n144 20.3299
R37458 C2S2_Amp_F_I_1.OUT.n161 C2S2_Amp_F_I_1.OUT.n157 20.3299
R37459 C2S2_Amp_F_I_1.OUT.n174 C2S2_Amp_F_I_1.OUT.n170 20.3299
R37460 C2S2_Amp_F_I_1.OUT.n187 C2S2_Amp_F_I_1.OUT.n183 20.3299
R37461 C2S2_Amp_F_I_1.OUT.n200 C2S2_Amp_F_I_1.OUT.n196 20.3299
R37462 C2S2_Amp_F_I_1.OUT.n213 C2S2_Amp_F_I_1.OUT.n209 20.3299
R37463 C2S2_Amp_F_I_1.OUT.n226 C2S2_Amp_F_I_1.OUT.n222 20.3299
R37464 C2S2_Amp_F_I_1.OUT.n239 C2S2_Amp_F_I_1.OUT.n235 20.3299
R37465 C2S2_Amp_F_I_1.OUT.n252 C2S2_Amp_F_I_1.OUT.n248 20.3299
R37466 C2S2_Amp_F_I_1.OUT.n265 C2S2_Amp_F_I_1.OUT.n261 20.3299
R37467 C2S2_Amp_F_I_1.OUT.n278 C2S2_Amp_F_I_1.OUT.n274 20.3299
R37468 C2S2_Amp_F_I_1.OUT.n291 C2S2_Amp_F_I_1.OUT.n287 20.3299
R37469 C2S2_Amp_F_I_1.OUT.n306 C2S2_Amp_F_I_1.OUT.n305 20.3299
R37470 C2S2_Amp_F_I_1.OUT.n59 C2S2_Amp_F_I_1.OUT.n58 20.3299
R37471 C2S2_Amp_F_I_1.OUT.n74 C2S2_Amp_F_I_1.OUT.n73 19.1618
R37472 C2S2_Amp_F_I_1.OUT.n87 C2S2_Amp_F_I_1.OUT.n86 19.1618
R37473 C2S2_Amp_F_I_1.OUT.n100 C2S2_Amp_F_I_1.OUT.n99 19.1618
R37474 C2S2_Amp_F_I_1.OUT.n113 C2S2_Amp_F_I_1.OUT.n112 19.1618
R37475 C2S2_Amp_F_I_1.OUT.n126 C2S2_Amp_F_I_1.OUT.n125 19.1618
R37476 C2S2_Amp_F_I_1.OUT.n139 C2S2_Amp_F_I_1.OUT.n138 19.1618
R37477 C2S2_Amp_F_I_1.OUT.n152 C2S2_Amp_F_I_1.OUT.n151 19.1618
R37478 C2S2_Amp_F_I_1.OUT.n165 C2S2_Amp_F_I_1.OUT.n164 19.1618
R37479 C2S2_Amp_F_I_1.OUT.n178 C2S2_Amp_F_I_1.OUT.n177 19.1618
R37480 C2S2_Amp_F_I_1.OUT.n191 C2S2_Amp_F_I_1.OUT.n190 19.1618
R37481 C2S2_Amp_F_I_1.OUT.n204 C2S2_Amp_F_I_1.OUT.n203 19.1618
R37482 C2S2_Amp_F_I_1.OUT.n217 C2S2_Amp_F_I_1.OUT.n216 19.1618
R37483 C2S2_Amp_F_I_1.OUT.n230 C2S2_Amp_F_I_1.OUT.n229 19.1618
R37484 C2S2_Amp_F_I_1.OUT.n243 C2S2_Amp_F_I_1.OUT.n242 19.1618
R37485 C2S2_Amp_F_I_1.OUT.n256 C2S2_Amp_F_I_1.OUT.n255 19.1618
R37486 C2S2_Amp_F_I_1.OUT.n269 C2S2_Amp_F_I_1.OUT.n268 19.1618
R37487 C2S2_Amp_F_I_1.OUT.n282 C2S2_Amp_F_I_1.OUT.n281 19.1618
R37488 C2S2_Amp_F_I_1.OUT.n295 C2S2_Amp_F_I_1.OUT.n294 19.1618
R37489 C2S2_Amp_F_I_1.OUT.n300 C2S2_Amp_F_I_1.OUT.n30 19.1618
R37490 C2S2_Amp_F_I_1.OUT.n53 C2S2_Amp_F_I_1.OUT.n52 19.1618
R37491 C2S2_Amp_F_I_1.OUT.n7 C2S2_Amp_F_I_1.OUT.n0 19.1591
R37492 C2S2_Amp_F_I_1.OUT.n336 C2S2_Amp_F_I_1.OUT.n332 19.1591
R37493 C2S2_Amp_F_I_1.OUT.n349 C2S2_Amp_F_I_1.OUT.n331 19.1591
R37494 C2S2_Amp_F_I_1.OUT.n362 C2S2_Amp_F_I_1.OUT.n330 19.1591
R37495 C2S2_Amp_F_I_1.OUT.n375 C2S2_Amp_F_I_1.OUT.n329 19.1591
R37496 C2S2_Amp_F_I_1.OUT.n388 C2S2_Amp_F_I_1.OUT.n328 19.1591
R37497 C2S2_Amp_F_I_1.OUT.n404 C2S2_Amp_F_I_1.OUT.n327 19.1591
R37498 C2S2_Amp_F_I_1.OUT.n11 C2S2_Amp_F_I_1.OUT.n6 18.824
R37499 C2S2_Amp_F_I_1.OUT.n340 C2S2_Amp_F_I_1.OUT.n335 18.824
R37500 C2S2_Amp_F_I_1.OUT.n353 C2S2_Amp_F_I_1.OUT.n348 18.824
R37501 C2S2_Amp_F_I_1.OUT.n366 C2S2_Amp_F_I_1.OUT.n361 18.824
R37502 C2S2_Amp_F_I_1.OUT.n379 C2S2_Amp_F_I_1.OUT.n374 18.824
R37503 C2S2_Amp_F_I_1.OUT.n392 C2S2_Amp_F_I_1.OUT.n387 18.824
R37504 C2S2_Amp_F_I_1.OUT.n408 C2S2_Amp_F_I_1.OUT.n403 18.824
R37505 C2S2_Amp_F_I_1.OUT.n67 C2S2_Amp_F_I_1.OUT.n65 18.824
R37506 C2S2_Amp_F_I_1.OUT.n80 C2S2_Amp_F_I_1.OUT.n78 18.824
R37507 C2S2_Amp_F_I_1.OUT.n93 C2S2_Amp_F_I_1.OUT.n91 18.824
R37508 C2S2_Amp_F_I_1.OUT.n106 C2S2_Amp_F_I_1.OUT.n104 18.824
R37509 C2S2_Amp_F_I_1.OUT.n119 C2S2_Amp_F_I_1.OUT.n117 18.824
R37510 C2S2_Amp_F_I_1.OUT.n132 C2S2_Amp_F_I_1.OUT.n130 18.824
R37511 C2S2_Amp_F_I_1.OUT.n145 C2S2_Amp_F_I_1.OUT.n143 18.824
R37512 C2S2_Amp_F_I_1.OUT.n158 C2S2_Amp_F_I_1.OUT.n156 18.824
R37513 C2S2_Amp_F_I_1.OUT.n171 C2S2_Amp_F_I_1.OUT.n169 18.824
R37514 C2S2_Amp_F_I_1.OUT.n184 C2S2_Amp_F_I_1.OUT.n182 18.824
R37515 C2S2_Amp_F_I_1.OUT.n197 C2S2_Amp_F_I_1.OUT.n195 18.824
R37516 C2S2_Amp_F_I_1.OUT.n210 C2S2_Amp_F_I_1.OUT.n208 18.824
R37517 C2S2_Amp_F_I_1.OUT.n223 C2S2_Amp_F_I_1.OUT.n221 18.824
R37518 C2S2_Amp_F_I_1.OUT.n236 C2S2_Amp_F_I_1.OUT.n234 18.824
R37519 C2S2_Amp_F_I_1.OUT.n249 C2S2_Amp_F_I_1.OUT.n247 18.824
R37520 C2S2_Amp_F_I_1.OUT.n262 C2S2_Amp_F_I_1.OUT.n260 18.824
R37521 C2S2_Amp_F_I_1.OUT.n275 C2S2_Amp_F_I_1.OUT.n273 18.824
R37522 C2S2_Amp_F_I_1.OUT.n288 C2S2_Amp_F_I_1.OUT.n286 18.824
R37523 C2S2_Amp_F_I_1.OUT.n303 C2S2_Amp_F_I_1.OUT.n299 18.824
R37524 C2S2_Amp_F_I_1.OUT.n56 C2S2_Amp_F_I_1.OUT.n51 18.824
R37525 C2S2_Amp_F_I_1.OUT.n8 C2S2_Amp_F_I_1.OUT.n7 17.3181
R37526 C2S2_Amp_F_I_1.OUT.n337 C2S2_Amp_F_I_1.OUT.n336 17.3181
R37527 C2S2_Amp_F_I_1.OUT.n350 C2S2_Amp_F_I_1.OUT.n349 17.3181
R37528 C2S2_Amp_F_I_1.OUT.n363 C2S2_Amp_F_I_1.OUT.n362 17.3181
R37529 C2S2_Amp_F_I_1.OUT.n376 C2S2_Amp_F_I_1.OUT.n375 17.3181
R37530 C2S2_Amp_F_I_1.OUT.n389 C2S2_Amp_F_I_1.OUT.n388 17.3181
R37531 C2S2_Amp_F_I_1.OUT.n405 C2S2_Amp_F_I_1.OUT.n404 17.3181
R37532 C2S2_Amp_F_I_1.OUT.n73 C2S2_Amp_F_I_1.OUT.n64 17.3181
R37533 C2S2_Amp_F_I_1.OUT.n86 C2S2_Amp_F_I_1.OUT.n77 17.3181
R37534 C2S2_Amp_F_I_1.OUT.n99 C2S2_Amp_F_I_1.OUT.n90 17.3181
R37535 C2S2_Amp_F_I_1.OUT.n112 C2S2_Amp_F_I_1.OUT.n103 17.3181
R37536 C2S2_Amp_F_I_1.OUT.n125 C2S2_Amp_F_I_1.OUT.n116 17.3181
R37537 C2S2_Amp_F_I_1.OUT.n138 C2S2_Amp_F_I_1.OUT.n129 17.3181
R37538 C2S2_Amp_F_I_1.OUT.n151 C2S2_Amp_F_I_1.OUT.n142 17.3181
R37539 C2S2_Amp_F_I_1.OUT.n164 C2S2_Amp_F_I_1.OUT.n155 17.3181
R37540 C2S2_Amp_F_I_1.OUT.n177 C2S2_Amp_F_I_1.OUT.n168 17.3181
R37541 C2S2_Amp_F_I_1.OUT.n190 C2S2_Amp_F_I_1.OUT.n181 17.3181
R37542 C2S2_Amp_F_I_1.OUT.n203 C2S2_Amp_F_I_1.OUT.n194 17.3181
R37543 C2S2_Amp_F_I_1.OUT.n216 C2S2_Amp_F_I_1.OUT.n207 17.3181
R37544 C2S2_Amp_F_I_1.OUT.n229 C2S2_Amp_F_I_1.OUT.n220 17.3181
R37545 C2S2_Amp_F_I_1.OUT.n242 C2S2_Amp_F_I_1.OUT.n233 17.3181
R37546 C2S2_Amp_F_I_1.OUT.n255 C2S2_Amp_F_I_1.OUT.n246 17.3181
R37547 C2S2_Amp_F_I_1.OUT.n268 C2S2_Amp_F_I_1.OUT.n259 17.3181
R37548 C2S2_Amp_F_I_1.OUT.n281 C2S2_Amp_F_I_1.OUT.n272 17.3181
R37549 C2S2_Amp_F_I_1.OUT.n294 C2S2_Amp_F_I_1.OUT.n285 17.3181
R37550 C2S2_Amp_F_I_1.OUT.n302 C2S2_Amp_F_I_1.OUT.n300 17.3181
R37551 C2S2_Amp_F_I_1.OUT.n55 C2S2_Amp_F_I_1.OUT.n52 17.3181
R37552 C2S2_Amp_F_I_1.OUT.n343 C2S2_Amp_F_I_1.OUT.n334 15.4484
R37553 C2S2_Amp_F_I_1.OUT.n356 C2S2_Amp_F_I_1.OUT.n347 15.4484
R37554 C2S2_Amp_F_I_1.OUT.n369 C2S2_Amp_F_I_1.OUT.n360 15.4484
R37555 C2S2_Amp_F_I_1.OUT.n382 C2S2_Amp_F_I_1.OUT.n373 15.4484
R37556 C2S2_Amp_F_I_1.OUT.n395 C2S2_Amp_F_I_1.OUT.n386 15.4484
R37557 C2S2_Amp_F_I_1.OUT.n20 C2S2_Amp_F_I_1.OUT.n19 9.3005
R37558 C2S2_Amp_F_I_1.OUT.n4 C2S2_Amp_F_I_1.OUT.n2 9.3005
R37559 C2S2_Amp_F_I_1.OUT.n26 C2S2_Amp_F_I_1.OUT.n25 9.3005
R37560 C2S2_Amp_F_I_1.OUT.n12 C2S2_Amp_F_I_1.OUT.n1 9.3005
R37561 C2S2_Amp_F_I_1.OUT.n11 C2S2_Amp_F_I_1.OUT.n10 9.3005
R37562 C2S2_Amp_F_I_1.OUT.n9 C2S2_Amp_F_I_1.OUT.n8 9.3005
R37563 C2S2_Amp_F_I_1.OUT.n342 C2S2_Amp_F_I_1.OUT.n333 9.3005
R37564 C2S2_Amp_F_I_1.OUT.n340 C2S2_Amp_F_I_1.OUT.n339 9.3005
R37565 C2S2_Amp_F_I_1.OUT.n338 C2S2_Amp_F_I_1.OUT.n337 9.3005
R37566 C2S2_Amp_F_I_1.OUT.n355 C2S2_Amp_F_I_1.OUT.n346 9.3005
R37567 C2S2_Amp_F_I_1.OUT.n353 C2S2_Amp_F_I_1.OUT.n352 9.3005
R37568 C2S2_Amp_F_I_1.OUT.n351 C2S2_Amp_F_I_1.OUT.n350 9.3005
R37569 C2S2_Amp_F_I_1.OUT.n368 C2S2_Amp_F_I_1.OUT.n359 9.3005
R37570 C2S2_Amp_F_I_1.OUT.n366 C2S2_Amp_F_I_1.OUT.n365 9.3005
R37571 C2S2_Amp_F_I_1.OUT.n364 C2S2_Amp_F_I_1.OUT.n363 9.3005
R37572 C2S2_Amp_F_I_1.OUT.n381 C2S2_Amp_F_I_1.OUT.n372 9.3005
R37573 C2S2_Amp_F_I_1.OUT.n379 C2S2_Amp_F_I_1.OUT.n378 9.3005
R37574 C2S2_Amp_F_I_1.OUT.n377 C2S2_Amp_F_I_1.OUT.n376 9.3005
R37575 C2S2_Amp_F_I_1.OUT.n394 C2S2_Amp_F_I_1.OUT.n385 9.3005
R37576 C2S2_Amp_F_I_1.OUT.n392 C2S2_Amp_F_I_1.OUT.n391 9.3005
R37577 C2S2_Amp_F_I_1.OUT.n390 C2S2_Amp_F_I_1.OUT.n389 9.3005
R37578 C2S2_Amp_F_I_1.OUT.n417 C2S2_Amp_F_I_1.OUT.n416 9.3005
R37579 C2S2_Amp_F_I_1.OUT.n401 C2S2_Amp_F_I_1.OUT.n399 9.3005
R37580 C2S2_Amp_F_I_1.OUT.n423 C2S2_Amp_F_I_1.OUT.n422 9.3005
R37581 C2S2_Amp_F_I_1.OUT.n409 C2S2_Amp_F_I_1.OUT.n398 9.3005
R37582 C2S2_Amp_F_I_1.OUT.n408 C2S2_Amp_F_I_1.OUT.n407 9.3005
R37583 C2S2_Amp_F_I_1.OUT.n406 C2S2_Amp_F_I_1.OUT.n405 9.3005
R37584 C2S2_Amp_F_I_1.OUT.n64 C2S2_Amp_F_I_1.OUT.n63 9.3005
R37585 C2S2_Amp_F_I_1.OUT.n70 C2S2_Amp_F_I_1.OUT.n69 9.3005
R37586 C2S2_Amp_F_I_1.OUT.n68 C2S2_Amp_F_I_1.OUT.n67 9.3005
R37587 C2S2_Amp_F_I_1.OUT.n77 C2S2_Amp_F_I_1.OUT.n76 9.3005
R37588 C2S2_Amp_F_I_1.OUT.n83 C2S2_Amp_F_I_1.OUT.n82 9.3005
R37589 C2S2_Amp_F_I_1.OUT.n81 C2S2_Amp_F_I_1.OUT.n80 9.3005
R37590 C2S2_Amp_F_I_1.OUT.n90 C2S2_Amp_F_I_1.OUT.n89 9.3005
R37591 C2S2_Amp_F_I_1.OUT.n96 C2S2_Amp_F_I_1.OUT.n95 9.3005
R37592 C2S2_Amp_F_I_1.OUT.n94 C2S2_Amp_F_I_1.OUT.n93 9.3005
R37593 C2S2_Amp_F_I_1.OUT.n103 C2S2_Amp_F_I_1.OUT.n102 9.3005
R37594 C2S2_Amp_F_I_1.OUT.n109 C2S2_Amp_F_I_1.OUT.n108 9.3005
R37595 C2S2_Amp_F_I_1.OUT.n107 C2S2_Amp_F_I_1.OUT.n106 9.3005
R37596 C2S2_Amp_F_I_1.OUT.n116 C2S2_Amp_F_I_1.OUT.n115 9.3005
R37597 C2S2_Amp_F_I_1.OUT.n122 C2S2_Amp_F_I_1.OUT.n121 9.3005
R37598 C2S2_Amp_F_I_1.OUT.n120 C2S2_Amp_F_I_1.OUT.n119 9.3005
R37599 C2S2_Amp_F_I_1.OUT.n129 C2S2_Amp_F_I_1.OUT.n128 9.3005
R37600 C2S2_Amp_F_I_1.OUT.n135 C2S2_Amp_F_I_1.OUT.n134 9.3005
R37601 C2S2_Amp_F_I_1.OUT.n133 C2S2_Amp_F_I_1.OUT.n132 9.3005
R37602 C2S2_Amp_F_I_1.OUT.n142 C2S2_Amp_F_I_1.OUT.n141 9.3005
R37603 C2S2_Amp_F_I_1.OUT.n148 C2S2_Amp_F_I_1.OUT.n147 9.3005
R37604 C2S2_Amp_F_I_1.OUT.n146 C2S2_Amp_F_I_1.OUT.n145 9.3005
R37605 C2S2_Amp_F_I_1.OUT.n155 C2S2_Amp_F_I_1.OUT.n154 9.3005
R37606 C2S2_Amp_F_I_1.OUT.n161 C2S2_Amp_F_I_1.OUT.n160 9.3005
R37607 C2S2_Amp_F_I_1.OUT.n159 C2S2_Amp_F_I_1.OUT.n158 9.3005
R37608 C2S2_Amp_F_I_1.OUT.n168 C2S2_Amp_F_I_1.OUT.n167 9.3005
R37609 C2S2_Amp_F_I_1.OUT.n174 C2S2_Amp_F_I_1.OUT.n173 9.3005
R37610 C2S2_Amp_F_I_1.OUT.n172 C2S2_Amp_F_I_1.OUT.n171 9.3005
R37611 C2S2_Amp_F_I_1.OUT.n181 C2S2_Amp_F_I_1.OUT.n180 9.3005
R37612 C2S2_Amp_F_I_1.OUT.n187 C2S2_Amp_F_I_1.OUT.n186 9.3005
R37613 C2S2_Amp_F_I_1.OUT.n185 C2S2_Amp_F_I_1.OUT.n184 9.3005
R37614 C2S2_Amp_F_I_1.OUT.n194 C2S2_Amp_F_I_1.OUT.n193 9.3005
R37615 C2S2_Amp_F_I_1.OUT.n200 C2S2_Amp_F_I_1.OUT.n199 9.3005
R37616 C2S2_Amp_F_I_1.OUT.n198 C2S2_Amp_F_I_1.OUT.n197 9.3005
R37617 C2S2_Amp_F_I_1.OUT.n207 C2S2_Amp_F_I_1.OUT.n206 9.3005
R37618 C2S2_Amp_F_I_1.OUT.n213 C2S2_Amp_F_I_1.OUT.n212 9.3005
R37619 C2S2_Amp_F_I_1.OUT.n211 C2S2_Amp_F_I_1.OUT.n210 9.3005
R37620 C2S2_Amp_F_I_1.OUT.n220 C2S2_Amp_F_I_1.OUT.n219 9.3005
R37621 C2S2_Amp_F_I_1.OUT.n226 C2S2_Amp_F_I_1.OUT.n225 9.3005
R37622 C2S2_Amp_F_I_1.OUT.n224 C2S2_Amp_F_I_1.OUT.n223 9.3005
R37623 C2S2_Amp_F_I_1.OUT.n233 C2S2_Amp_F_I_1.OUT.n232 9.3005
R37624 C2S2_Amp_F_I_1.OUT.n239 C2S2_Amp_F_I_1.OUT.n238 9.3005
R37625 C2S2_Amp_F_I_1.OUT.n237 C2S2_Amp_F_I_1.OUT.n236 9.3005
R37626 C2S2_Amp_F_I_1.OUT.n246 C2S2_Amp_F_I_1.OUT.n245 9.3005
R37627 C2S2_Amp_F_I_1.OUT.n252 C2S2_Amp_F_I_1.OUT.n251 9.3005
R37628 C2S2_Amp_F_I_1.OUT.n250 C2S2_Amp_F_I_1.OUT.n249 9.3005
R37629 C2S2_Amp_F_I_1.OUT.n259 C2S2_Amp_F_I_1.OUT.n258 9.3005
R37630 C2S2_Amp_F_I_1.OUT.n265 C2S2_Amp_F_I_1.OUT.n264 9.3005
R37631 C2S2_Amp_F_I_1.OUT.n263 C2S2_Amp_F_I_1.OUT.n262 9.3005
R37632 C2S2_Amp_F_I_1.OUT.n272 C2S2_Amp_F_I_1.OUT.n271 9.3005
R37633 C2S2_Amp_F_I_1.OUT.n278 C2S2_Amp_F_I_1.OUT.n277 9.3005
R37634 C2S2_Amp_F_I_1.OUT.n276 C2S2_Amp_F_I_1.OUT.n275 9.3005
R37635 C2S2_Amp_F_I_1.OUT.n285 C2S2_Amp_F_I_1.OUT.n284 9.3005
R37636 C2S2_Amp_F_I_1.OUT.n291 C2S2_Amp_F_I_1.OUT.n290 9.3005
R37637 C2S2_Amp_F_I_1.OUT.n289 C2S2_Amp_F_I_1.OUT.n288 9.3005
R37638 C2S2_Amp_F_I_1.OUT.n302 C2S2_Amp_F_I_1.OUT.n301 9.3005
R37639 C2S2_Amp_F_I_1.OUT.n307 C2S2_Amp_F_I_1.OUT.n306 9.3005
R37640 C2S2_Amp_F_I_1.OUT.n299 C2S2_Amp_F_I_1.OUT.n298 9.3005
R37641 C2S2_Amp_F_I_1.OUT.n55 C2S2_Amp_F_I_1.OUT.n54 9.3005
R37642 C2S2_Amp_F_I_1.OUT.n60 C2S2_Amp_F_I_1.OUT.n59 9.3005
R37643 C2S2_Amp_F_I_1.OUT.n51 C2S2_Amp_F_I_1.OUT.n50 9.3005
R37644 C2S2_Amp_F_I_1.OUT.n8 C2S2_Amp_F_I_1.OUT.n6 8.28285
R37645 C2S2_Amp_F_I_1.OUT.n337 C2S2_Amp_F_I_1.OUT.n335 8.28285
R37646 C2S2_Amp_F_I_1.OUT.n350 C2S2_Amp_F_I_1.OUT.n348 8.28285
R37647 C2S2_Amp_F_I_1.OUT.n363 C2S2_Amp_F_I_1.OUT.n361 8.28285
R37648 C2S2_Amp_F_I_1.OUT.n376 C2S2_Amp_F_I_1.OUT.n374 8.28285
R37649 C2S2_Amp_F_I_1.OUT.n389 C2S2_Amp_F_I_1.OUT.n387 8.28285
R37650 C2S2_Amp_F_I_1.OUT.n405 C2S2_Amp_F_I_1.OUT.n403 8.28285
R37651 C2S2_Amp_F_I_1.OUT.n65 C2S2_Amp_F_I_1.OUT.n64 8.28285
R37652 C2S2_Amp_F_I_1.OUT.n78 C2S2_Amp_F_I_1.OUT.n77 8.28285
R37653 C2S2_Amp_F_I_1.OUT.n91 C2S2_Amp_F_I_1.OUT.n90 8.28285
R37654 C2S2_Amp_F_I_1.OUT.n104 C2S2_Amp_F_I_1.OUT.n103 8.28285
R37655 C2S2_Amp_F_I_1.OUT.n117 C2S2_Amp_F_I_1.OUT.n116 8.28285
R37656 C2S2_Amp_F_I_1.OUT.n130 C2S2_Amp_F_I_1.OUT.n129 8.28285
R37657 C2S2_Amp_F_I_1.OUT.n143 C2S2_Amp_F_I_1.OUT.n142 8.28285
R37658 C2S2_Amp_F_I_1.OUT.n156 C2S2_Amp_F_I_1.OUT.n155 8.28285
R37659 C2S2_Amp_F_I_1.OUT.n169 C2S2_Amp_F_I_1.OUT.n168 8.28285
R37660 C2S2_Amp_F_I_1.OUT.n182 C2S2_Amp_F_I_1.OUT.n181 8.28285
R37661 C2S2_Amp_F_I_1.OUT.n195 C2S2_Amp_F_I_1.OUT.n194 8.28285
R37662 C2S2_Amp_F_I_1.OUT.n208 C2S2_Amp_F_I_1.OUT.n207 8.28285
R37663 C2S2_Amp_F_I_1.OUT.n221 C2S2_Amp_F_I_1.OUT.n220 8.28285
R37664 C2S2_Amp_F_I_1.OUT.n234 C2S2_Amp_F_I_1.OUT.n233 8.28285
R37665 C2S2_Amp_F_I_1.OUT.n247 C2S2_Amp_F_I_1.OUT.n246 8.28285
R37666 C2S2_Amp_F_I_1.OUT.n260 C2S2_Amp_F_I_1.OUT.n259 8.28285
R37667 C2S2_Amp_F_I_1.OUT.n273 C2S2_Amp_F_I_1.OUT.n272 8.28285
R37668 C2S2_Amp_F_I_1.OUT.n286 C2S2_Amp_F_I_1.OUT.n285 8.28285
R37669 C2S2_Amp_F_I_1.OUT.n303 C2S2_Amp_F_I_1.OUT.n302 8.28285
R37670 C2S2_Amp_F_I_1.OUT.n56 C2S2_Amp_F_I_1.OUT.n55 8.28285
R37671 C2S2_Amp_F_I_1.OUT.n433 C2S2_Amp_F_I_1.OUT.n432 8.09988
R37672 C2S2_Amp_F_I_1.OUT.n427 C2S2_Amp_F_I_1.OUT.n426 8.09988
R37673 C2S2_Amp_F_I_1.OUT.n28 C2S2_Amp_F_I_1.OUT.n0 7.9105
R37674 C2S2_Amp_F_I_1.OUT.n345 C2S2_Amp_F_I_1.OUT.n332 7.9105
R37675 C2S2_Amp_F_I_1.OUT.n358 C2S2_Amp_F_I_1.OUT.n331 7.9105
R37676 C2S2_Amp_F_I_1.OUT.n371 C2S2_Amp_F_I_1.OUT.n330 7.9105
R37677 C2S2_Amp_F_I_1.OUT.n384 C2S2_Amp_F_I_1.OUT.n329 7.9105
R37678 C2S2_Amp_F_I_1.OUT.n397 C2S2_Amp_F_I_1.OUT.n328 7.9105
R37679 C2S2_Amp_F_I_1.OUT.n425 C2S2_Amp_F_I_1.OUT.n327 7.9105
R37680 C2S2_Amp_F_I_1.OUT.n75 C2S2_Amp_F_I_1.OUT.n48 7.9105
R37681 C2S2_Amp_F_I_1.OUT.n88 C2S2_Amp_F_I_1.OUT.n47 7.9105
R37682 C2S2_Amp_F_I_1.OUT.n101 C2S2_Amp_F_I_1.OUT.n46 7.9105
R37683 C2S2_Amp_F_I_1.OUT.n114 C2S2_Amp_F_I_1.OUT.n45 7.9105
R37684 C2S2_Amp_F_I_1.OUT.n127 C2S2_Amp_F_I_1.OUT.n44 7.9105
R37685 C2S2_Amp_F_I_1.OUT.n140 C2S2_Amp_F_I_1.OUT.n43 7.9105
R37686 C2S2_Amp_F_I_1.OUT.n153 C2S2_Amp_F_I_1.OUT.n42 7.9105
R37687 C2S2_Amp_F_I_1.OUT.n166 C2S2_Amp_F_I_1.OUT.n41 7.9105
R37688 C2S2_Amp_F_I_1.OUT.n179 C2S2_Amp_F_I_1.OUT.n40 7.9105
R37689 C2S2_Amp_F_I_1.OUT.n192 C2S2_Amp_F_I_1.OUT.n39 7.9105
R37690 C2S2_Amp_F_I_1.OUT.n205 C2S2_Amp_F_I_1.OUT.n38 7.9105
R37691 C2S2_Amp_F_I_1.OUT.n218 C2S2_Amp_F_I_1.OUT.n37 7.9105
R37692 C2S2_Amp_F_I_1.OUT.n231 C2S2_Amp_F_I_1.OUT.n36 7.9105
R37693 C2S2_Amp_F_I_1.OUT.n244 C2S2_Amp_F_I_1.OUT.n35 7.9105
R37694 C2S2_Amp_F_I_1.OUT.n257 C2S2_Amp_F_I_1.OUT.n34 7.9105
R37695 C2S2_Amp_F_I_1.OUT.n270 C2S2_Amp_F_I_1.OUT.n33 7.9105
R37696 C2S2_Amp_F_I_1.OUT.n283 C2S2_Amp_F_I_1.OUT.n32 7.9105
R37697 C2S2_Amp_F_I_1.OUT.n296 C2S2_Amp_F_I_1.OUT.n31 7.9105
R37698 C2S2_Amp_F_I_1.OUT.n296 C2S2_Amp_F_I_1.OUT.n295 7.9105
R37699 C2S2_Amp_F_I_1.OUT.n283 C2S2_Amp_F_I_1.OUT.n282 7.9105
R37700 C2S2_Amp_F_I_1.OUT.n270 C2S2_Amp_F_I_1.OUT.n269 7.9105
R37701 C2S2_Amp_F_I_1.OUT.n257 C2S2_Amp_F_I_1.OUT.n256 7.9105
R37702 C2S2_Amp_F_I_1.OUT.n244 C2S2_Amp_F_I_1.OUT.n243 7.9105
R37703 C2S2_Amp_F_I_1.OUT.n231 C2S2_Amp_F_I_1.OUT.n230 7.9105
R37704 C2S2_Amp_F_I_1.OUT.n218 C2S2_Amp_F_I_1.OUT.n217 7.9105
R37705 C2S2_Amp_F_I_1.OUT.n205 C2S2_Amp_F_I_1.OUT.n204 7.9105
R37706 C2S2_Amp_F_I_1.OUT.n192 C2S2_Amp_F_I_1.OUT.n191 7.9105
R37707 C2S2_Amp_F_I_1.OUT.n179 C2S2_Amp_F_I_1.OUT.n178 7.9105
R37708 C2S2_Amp_F_I_1.OUT.n166 C2S2_Amp_F_I_1.OUT.n165 7.9105
R37709 C2S2_Amp_F_I_1.OUT.n153 C2S2_Amp_F_I_1.OUT.n152 7.9105
R37710 C2S2_Amp_F_I_1.OUT.n140 C2S2_Amp_F_I_1.OUT.n139 7.9105
R37711 C2S2_Amp_F_I_1.OUT.n127 C2S2_Amp_F_I_1.OUT.n126 7.9105
R37712 C2S2_Amp_F_I_1.OUT.n114 C2S2_Amp_F_I_1.OUT.n113 7.9105
R37713 C2S2_Amp_F_I_1.OUT.n101 C2S2_Amp_F_I_1.OUT.n100 7.9105
R37714 C2S2_Amp_F_I_1.OUT.n88 C2S2_Amp_F_I_1.OUT.n87 7.9105
R37715 C2S2_Amp_F_I_1.OUT.n75 C2S2_Amp_F_I_1.OUT.n74 7.9105
R37716 C2S2_Amp_F_I_1.OUT.n425 C2S2_Amp_F_I_1.OUT.n424 7.9105
R37717 C2S2_Amp_F_I_1.OUT.n397 C2S2_Amp_F_I_1.OUT.n396 7.9105
R37718 C2S2_Amp_F_I_1.OUT.n384 C2S2_Amp_F_I_1.OUT.n383 7.9105
R37719 C2S2_Amp_F_I_1.OUT.n371 C2S2_Amp_F_I_1.OUT.n370 7.9105
R37720 C2S2_Amp_F_I_1.OUT.n358 C2S2_Amp_F_I_1.OUT.n357 7.9105
R37721 C2S2_Amp_F_I_1.OUT.n345 C2S2_Amp_F_I_1.OUT.n344 7.9105
R37722 C2S2_Amp_F_I_1.OUT.n28 C2S2_Amp_F_I_1.OUT.n27 7.9105
R37723 C2S2_Amp_F_I_1.OUT.n13 C2S2_Amp_F_I_1.OUT.n11 6.77697
R37724 C2S2_Amp_F_I_1.OUT.n341 C2S2_Amp_F_I_1.OUT.n340 6.77697
R37725 C2S2_Amp_F_I_1.OUT.n354 C2S2_Amp_F_I_1.OUT.n353 6.77697
R37726 C2S2_Amp_F_I_1.OUT.n367 C2S2_Amp_F_I_1.OUT.n366 6.77697
R37727 C2S2_Amp_F_I_1.OUT.n380 C2S2_Amp_F_I_1.OUT.n379 6.77697
R37728 C2S2_Amp_F_I_1.OUT.n393 C2S2_Amp_F_I_1.OUT.n392 6.77697
R37729 C2S2_Amp_F_I_1.OUT.n410 C2S2_Amp_F_I_1.OUT.n408 6.77697
R37730 C2S2_Amp_F_I_1.OUT.n67 C2S2_Amp_F_I_1.OUT.n66 6.77697
R37731 C2S2_Amp_F_I_1.OUT.n80 C2S2_Amp_F_I_1.OUT.n79 6.77697
R37732 C2S2_Amp_F_I_1.OUT.n93 C2S2_Amp_F_I_1.OUT.n92 6.77697
R37733 C2S2_Amp_F_I_1.OUT.n106 C2S2_Amp_F_I_1.OUT.n105 6.77697
R37734 C2S2_Amp_F_I_1.OUT.n119 C2S2_Amp_F_I_1.OUT.n118 6.77697
R37735 C2S2_Amp_F_I_1.OUT.n132 C2S2_Amp_F_I_1.OUT.n131 6.77697
R37736 C2S2_Amp_F_I_1.OUT.n145 C2S2_Amp_F_I_1.OUT.n144 6.77697
R37737 C2S2_Amp_F_I_1.OUT.n158 C2S2_Amp_F_I_1.OUT.n157 6.77697
R37738 C2S2_Amp_F_I_1.OUT.n171 C2S2_Amp_F_I_1.OUT.n170 6.77697
R37739 C2S2_Amp_F_I_1.OUT.n184 C2S2_Amp_F_I_1.OUT.n183 6.77697
R37740 C2S2_Amp_F_I_1.OUT.n197 C2S2_Amp_F_I_1.OUT.n196 6.77697
R37741 C2S2_Amp_F_I_1.OUT.n210 C2S2_Amp_F_I_1.OUT.n209 6.77697
R37742 C2S2_Amp_F_I_1.OUT.n223 C2S2_Amp_F_I_1.OUT.n222 6.77697
R37743 C2S2_Amp_F_I_1.OUT.n236 C2S2_Amp_F_I_1.OUT.n235 6.77697
R37744 C2S2_Amp_F_I_1.OUT.n249 C2S2_Amp_F_I_1.OUT.n248 6.77697
R37745 C2S2_Amp_F_I_1.OUT.n262 C2S2_Amp_F_I_1.OUT.n261 6.77697
R37746 C2S2_Amp_F_I_1.OUT.n275 C2S2_Amp_F_I_1.OUT.n274 6.77697
R37747 C2S2_Amp_F_I_1.OUT.n288 C2S2_Amp_F_I_1.OUT.n287 6.77697
R37748 C2S2_Amp_F_I_1.OUT.n305 C2S2_Amp_F_I_1.OUT.n299 6.77697
R37749 C2S2_Amp_F_I_1.OUT.n58 C2S2_Amp_F_I_1.OUT.n51 6.77697
R37750 C2S2_Amp_F_I_1.OUT.n432 C2S2_Amp_F_I_1.OUT.n431 6.14516
R37751 C2S2_Amp_F_I_1.OUT.n428 C2S2_Amp_F_I_1.OUT.n427 6.1428
R37752 C2S2_Amp_F_I_1.OUT.n72 C2S2_Amp_F_I_1.OUT.t61 5.7135
R37753 C2S2_Amp_F_I_1.OUT.n72 C2S2_Amp_F_I_1.OUT.t51 5.7135
R37754 C2S2_Amp_F_I_1.OUT.n85 C2S2_Amp_F_I_1.OUT.t28 5.7135
R37755 C2S2_Amp_F_I_1.OUT.n85 C2S2_Amp_F_I_1.OUT.t64 5.7135
R37756 C2S2_Amp_F_I_1.OUT.n98 C2S2_Amp_F_I_1.OUT.t56 5.7135
R37757 C2S2_Amp_F_I_1.OUT.n98 C2S2_Amp_F_I_1.OUT.t47 5.7135
R37758 C2S2_Amp_F_I_1.OUT.n111 C2S2_Amp_F_I_1.OUT.t48 5.7135
R37759 C2S2_Amp_F_I_1.OUT.n111 C2S2_Amp_F_I_1.OUT.t37 5.7135
R37760 C2S2_Amp_F_I_1.OUT.n124 C2S2_Amp_F_I_1.OUT.t30 5.7135
R37761 C2S2_Amp_F_I_1.OUT.n124 C2S2_Amp_F_I_1.OUT.t58 5.7135
R37762 C2S2_Amp_F_I_1.OUT.n137 C2S2_Amp_F_I_1.OUT.t44 5.7135
R37763 C2S2_Amp_F_I_1.OUT.n137 C2S2_Amp_F_I_1.OUT.t38 5.7135
R37764 C2S2_Amp_F_I_1.OUT.n150 C2S2_Amp_F_I_1.OUT.t41 5.7135
R37765 C2S2_Amp_F_I_1.OUT.n150 C2S2_Amp_F_I_1.OUT.t31 5.7135
R37766 C2S2_Amp_F_I_1.OUT.n163 C2S2_Amp_F_I_1.OUT.t26 5.7135
R37767 C2S2_Amp_F_I_1.OUT.n163 C2S2_Amp_F_I_1.OUT.t62 5.7135
R37768 C2S2_Amp_F_I_1.OUT.n176 C2S2_Amp_F_I_1.OUT.t34 5.7135
R37769 C2S2_Amp_F_I_1.OUT.n176 C2S2_Amp_F_I_1.OUT.t29 5.7135
R37770 C2S2_Amp_F_I_1.OUT.n189 C2S2_Amp_F_I_1.OUT.t45 5.7135
R37771 C2S2_Amp_F_I_1.OUT.n189 C2S2_Amp_F_I_1.OUT.t39 5.7135
R37772 C2S2_Amp_F_I_1.OUT.n202 C2S2_Amp_F_I_1.OUT.t59 5.7135
R37773 C2S2_Amp_F_I_1.OUT.n202 C2S2_Amp_F_I_1.OUT.t54 5.7135
R37774 C2S2_Amp_F_I_1.OUT.n215 C2S2_Amp_F_I_1.OUT.t27 5.7135
R37775 C2S2_Amp_F_I_1.OUT.n215 C2S2_Amp_F_I_1.OUT.t25 5.7135
R37776 C2S2_Amp_F_I_1.OUT.n228 C2S2_Amp_F_I_1.OUT.t32 5.7135
R37777 C2S2_Amp_F_I_1.OUT.n228 C2S2_Amp_F_I_1.OUT.t49 5.7135
R37778 C2S2_Amp_F_I_1.OUT.n241 C2S2_Amp_F_I_1.OUT.t52 5.7135
R37779 C2S2_Amp_F_I_1.OUT.n241 C2S2_Amp_F_I_1.OUT.t43 5.7135
R37780 C2S2_Amp_F_I_1.OUT.n254 C2S2_Amp_F_I_1.OUT.t33 5.7135
R37781 C2S2_Amp_F_I_1.OUT.n254 C2S2_Amp_F_I_1.OUT.t57 5.7135
R37782 C2S2_Amp_F_I_1.OUT.n267 C2S2_Amp_F_I_1.OUT.t46 5.7135
R37783 C2S2_Amp_F_I_1.OUT.n267 C2S2_Amp_F_I_1.OUT.t36 5.7135
R37784 C2S2_Amp_F_I_1.OUT.n280 C2S2_Amp_F_I_1.OUT.t60 5.7135
R37785 C2S2_Amp_F_I_1.OUT.n280 C2S2_Amp_F_I_1.OUT.t55 5.7135
R37786 C2S2_Amp_F_I_1.OUT.n293 C2S2_Amp_F_I_1.OUT.t40 5.7135
R37787 C2S2_Amp_F_I_1.OUT.n293 C2S2_Amp_F_I_1.OUT.t35 5.7135
R37788 C2S2_Amp_F_I_1.OUT.n304 C2S2_Amp_F_I_1.OUT.t53 5.7135
R37789 C2S2_Amp_F_I_1.OUT.n304 C2S2_Amp_F_I_1.OUT.t50 5.7135
R37790 C2S2_Amp_F_I_1.OUT.n57 C2S2_Amp_F_I_1.OUT.t63 5.7135
R37791 C2S2_Amp_F_I_1.OUT.n57 C2S2_Amp_F_I_1.OUT.t42 5.7135
R37792 C2S2_Amp_F_I_1.OUT.n19 C2S2_Amp_F_I_1.OUT.n18 5.33935
R37793 C2S2_Amp_F_I_1.OUT.n416 C2S2_Amp_F_I_1.OUT.n415 5.33935
R37794 C2S2_Amp_F_I_1.OUT.n12 C2S2_Amp_F_I_1.OUT.n3 5.27109
R37795 C2S2_Amp_F_I_1.OUT.n409 C2S2_Amp_F_I_1.OUT.n400 5.27109
R37796 C2S2_Amp_F_I_1.OUT.n309 C2S2_Amp_F_I_1.OUT.n308 4.61261
R37797 C2S2_Amp_F_I_1.OUT.n62 C2S2_Amp_F_I_1.OUT.n61 4.61261
R37798 C2S2_Amp_F_I_1.OUT.n310 C2S2_Amp_F_I_1.OUT.n30 4.5005
R37799 C2S2_Amp_F_I_1.OUT.n53 C2S2_Amp_F_I_1.OUT.n29 4.5005
R37800 C2S2_Amp_F_I_1.OUT.n25 C2S2_Amp_F_I_1.OUT.n24 3.76521
R37801 C2S2_Amp_F_I_1.OUT.n422 C2S2_Amp_F_I_1.OUT.n421 3.76521
R37802 C2S2_Amp_F_I_1.OUT.n334 C2S2_Amp_F_I_1.OUT.t18 3.4805
R37803 C2S2_Amp_F_I_1.OUT.n334 C2S2_Amp_F_I_1.OUT.t14 3.4805
R37804 C2S2_Amp_F_I_1.OUT.n347 C2S2_Amp_F_I_1.OUT.t16 3.4805
R37805 C2S2_Amp_F_I_1.OUT.n347 C2S2_Amp_F_I_1.OUT.t15 3.4805
R37806 C2S2_Amp_F_I_1.OUT.n360 C2S2_Amp_F_I_1.OUT.t23 3.4805
R37807 C2S2_Amp_F_I_1.OUT.n360 C2S2_Amp_F_I_1.OUT.t19 3.4805
R37808 C2S2_Amp_F_I_1.OUT.n373 C2S2_Amp_F_I_1.OUT.t24 3.4805
R37809 C2S2_Amp_F_I_1.OUT.n373 C2S2_Amp_F_I_1.OUT.t21 3.4805
R37810 C2S2_Amp_F_I_1.OUT.n386 C2S2_Amp_F_I_1.OUT.t22 3.4805
R37811 C2S2_Amp_F_I_1.OUT.n386 C2S2_Amp_F_I_1.OUT.t13 3.4805
R37812 C2S2_Amp_F_I_1.OUT.n71 C2S2_Amp_F_I_1.OUT.n48 3.38566
R37813 C2S2_Amp_F_I_1.OUT.n84 C2S2_Amp_F_I_1.OUT.n47 3.38566
R37814 C2S2_Amp_F_I_1.OUT.n97 C2S2_Amp_F_I_1.OUT.n46 3.38566
R37815 C2S2_Amp_F_I_1.OUT.n110 C2S2_Amp_F_I_1.OUT.n45 3.38566
R37816 C2S2_Amp_F_I_1.OUT.n123 C2S2_Amp_F_I_1.OUT.n44 3.38566
R37817 C2S2_Amp_F_I_1.OUT.n136 C2S2_Amp_F_I_1.OUT.n43 3.38566
R37818 C2S2_Amp_F_I_1.OUT.n149 C2S2_Amp_F_I_1.OUT.n42 3.38566
R37819 C2S2_Amp_F_I_1.OUT.n162 C2S2_Amp_F_I_1.OUT.n41 3.38566
R37820 C2S2_Amp_F_I_1.OUT.n175 C2S2_Amp_F_I_1.OUT.n40 3.38566
R37821 C2S2_Amp_F_I_1.OUT.n188 C2S2_Amp_F_I_1.OUT.n39 3.38566
R37822 C2S2_Amp_F_I_1.OUT.n201 C2S2_Amp_F_I_1.OUT.n38 3.38566
R37823 C2S2_Amp_F_I_1.OUT.n214 C2S2_Amp_F_I_1.OUT.n37 3.38566
R37824 C2S2_Amp_F_I_1.OUT.n227 C2S2_Amp_F_I_1.OUT.n36 3.38566
R37825 C2S2_Amp_F_I_1.OUT.n240 C2S2_Amp_F_I_1.OUT.n35 3.38566
R37826 C2S2_Amp_F_I_1.OUT.n253 C2S2_Amp_F_I_1.OUT.n34 3.38566
R37827 C2S2_Amp_F_I_1.OUT.n266 C2S2_Amp_F_I_1.OUT.n33 3.38566
R37828 C2S2_Amp_F_I_1.OUT.n279 C2S2_Amp_F_I_1.OUT.n32 3.38566
R37829 C2S2_Amp_F_I_1.OUT.n292 C2S2_Amp_F_I_1.OUT.n31 3.38566
R37830 C2S2_Amp_F_I_1.OUT.n308 C2S2_Amp_F_I_1.OUT.n297 3.38566
R37831 C2S2_Amp_F_I_1.OUT.n61 C2S2_Amp_F_I_1.OUT.n49 3.38566
R37832 C2S2_Amp_F_I_1.OUT.n344 C2S2_Amp_F_I_1.OUT.n343 3.38531
R37833 C2S2_Amp_F_I_1.OUT.n357 C2S2_Amp_F_I_1.OUT.n356 3.38531
R37834 C2S2_Amp_F_I_1.OUT.n370 C2S2_Amp_F_I_1.OUT.n369 3.38531
R37835 C2S2_Amp_F_I_1.OUT.n383 C2S2_Amp_F_I_1.OUT.n382 3.38531
R37836 C2S2_Amp_F_I_1.OUT.n396 C2S2_Amp_F_I_1.OUT.n395 3.38531
R37837 C2S2_Amp_F_I_1.OUT.n21 C2S2_Amp_F_I_1.OUT.n4 2.25932
R37838 C2S2_Amp_F_I_1.OUT.n418 C2S2_Amp_F_I_1.OUT.n401 2.25932
R37839 C2S2_Amp_F_I_1.OUT.n325 C2S2_Amp_F_I_1.OUT.n324 2.25175
R37840 C2S2_Amp_F_I_1.OUT.n326 C2S2_Amp_F_I_1.OUT.n325 2.251
R37841 C2S2_Amp_F_I_1.OUT.n309 C2S2_Amp_F_I_1.OUT.n296 1.69577
R37842 C2S2_Amp_F_I_1.OUT.n75 C2S2_Amp_F_I_1.OUT.n62 1.69435
R37843 C2S2_Amp_F_I_1.OUT.n320 C2S2_Amp_F_I_1.OUT.t7 1.67859
R37844 C2S2_Amp_F_I_1.OUT.n316 C2S2_Amp_F_I_1.OUT.t11 1.67859
R37845 C2S2_Amp_F_I_1.OUT.n313 C2S2_Amp_F_I_1.OUT.t4 1.67859
R37846 C2S2_Amp_F_I_1.OUT.n322 C2S2_Amp_F_I_1.OUT.n321 1.56415
R37847 C2S2_Amp_F_I_1.OUT.n321 C2S2_Amp_F_I_1.OUT.n320 1.56415
R37848 C2S2_Amp_F_I_1.OUT.n318 C2S2_Amp_F_I_1.OUT.n317 1.56415
R37849 C2S2_Amp_F_I_1.OUT.n317 C2S2_Amp_F_I_1.OUT.n316 1.56415
R37850 C2S2_Amp_F_I_1.OUT.n315 C2S2_Amp_F_I_1.OUT.n314 1.56415
R37851 C2S2_Amp_F_I_1.OUT.n314 C2S2_Amp_F_I_1.OUT.n313 1.56415
R37852 C2S2_Amp_F_I_1.OUT.n319 C2S2_Amp_F_I_1.OUT.n315 1.55853
R37853 C2S2_Amp_F_I_1.OUT.n426 C2S2_Amp_F_I_1.OUT.n326 1.50074
R37854 C2S2_Amp_F_I_1.OUT.n323 C2S2_Amp_F_I_1.OUT.n322 1.17065
R37855 C2S2_Amp_F_I_1.OUT.n319 C2S2_Amp_F_I_1.OUT.n318 0.947532
R37856 C2S2_Amp_F_I_1.OUT.n312 C2S2_Amp_F_I_1.OUT.n311 0.805675
R37857 C2S2_Amp_F_I_1.OUT.n20 C2S2_Amp_F_I_1.OUT.n17 0.753441
R37858 C2S2_Amp_F_I_1.OUT.n417 C2S2_Amp_F_I_1.OUT.n414 0.753441
R37859 C2S2_Amp_F_I_1.OUT.n324 C2S2_Amp_F_I_1.OUT.n323 0.634315
R37860 C2S2_Amp_F_I_1.OUT C2S2_Amp_F_I_1.OUT.n433 0.557685
R37861 C2S2_Amp_F_I_1.OUT.n427 C2S2_Amp_F_I_1.OUT.n310 0.356269
R37862 C2S2_Amp_F_I_1.OUT.n432 C2S2_Amp_F_I_1.OUT.n29 0.356269
R37863 C2S2_Amp_F_I_1.OUT.n323 C2S2_Amp_F_I_1.OUT.n319 0.22362
R37864 C2S2_Amp_F_I_1.OUT.n26 C2S2_Amp_F_I_1.OUT.n2 0.196152
R37865 C2S2_Amp_F_I_1.OUT.n19 C2S2_Amp_F_I_1.OUT.n2 0.196152
R37866 C2S2_Amp_F_I_1.OUT.n423 C2S2_Amp_F_I_1.OUT.n399 0.196152
R37867 C2S2_Amp_F_I_1.OUT.n416 C2S2_Amp_F_I_1.OUT.n399 0.196152
R37868 C2S2_Amp_F_I_1.OUT.n69 C2S2_Amp_F_I_1.OUT.n68 0.196152
R37869 C2S2_Amp_F_I_1.OUT.n82 C2S2_Amp_F_I_1.OUT.n81 0.196152
R37870 C2S2_Amp_F_I_1.OUT.n95 C2S2_Amp_F_I_1.OUT.n94 0.196152
R37871 C2S2_Amp_F_I_1.OUT.n108 C2S2_Amp_F_I_1.OUT.n107 0.196152
R37872 C2S2_Amp_F_I_1.OUT.n121 C2S2_Amp_F_I_1.OUT.n120 0.196152
R37873 C2S2_Amp_F_I_1.OUT.n134 C2S2_Amp_F_I_1.OUT.n133 0.196152
R37874 C2S2_Amp_F_I_1.OUT.n147 C2S2_Amp_F_I_1.OUT.n146 0.196152
R37875 C2S2_Amp_F_I_1.OUT.n160 C2S2_Amp_F_I_1.OUT.n159 0.196152
R37876 C2S2_Amp_F_I_1.OUT.n173 C2S2_Amp_F_I_1.OUT.n172 0.196152
R37877 C2S2_Amp_F_I_1.OUT.n186 C2S2_Amp_F_I_1.OUT.n185 0.196152
R37878 C2S2_Amp_F_I_1.OUT.n199 C2S2_Amp_F_I_1.OUT.n198 0.196152
R37879 C2S2_Amp_F_I_1.OUT.n212 C2S2_Amp_F_I_1.OUT.n211 0.196152
R37880 C2S2_Amp_F_I_1.OUT.n225 C2S2_Amp_F_I_1.OUT.n224 0.196152
R37881 C2S2_Amp_F_I_1.OUT.n238 C2S2_Amp_F_I_1.OUT.n237 0.196152
R37882 C2S2_Amp_F_I_1.OUT.n251 C2S2_Amp_F_I_1.OUT.n250 0.196152
R37883 C2S2_Amp_F_I_1.OUT.n264 C2S2_Amp_F_I_1.OUT.n263 0.196152
R37884 C2S2_Amp_F_I_1.OUT.n277 C2S2_Amp_F_I_1.OUT.n276 0.196152
R37885 C2S2_Amp_F_I_1.OUT.n290 C2S2_Amp_F_I_1.OUT.n289 0.196152
R37886 C2S2_Amp_F_I_1.OUT.n307 C2S2_Amp_F_I_1.OUT.n298 0.196152
R37887 C2S2_Amp_F_I_1.OUT.n60 C2S2_Amp_F_I_1.OUT.n50 0.196152
R37888 C2S2_Amp_F_I_1.OUT.n312 C2S2_Amp_F_I_1.OUT.t0 0.192791
R37889 C2S2_Amp_F_I_1.OUT.n10 C2S2_Amp_F_I_1.OUT.n9 0.188181
R37890 C2S2_Amp_F_I_1.OUT.n339 C2S2_Amp_F_I_1.OUT.n338 0.188181
R37891 C2S2_Amp_F_I_1.OUT.n352 C2S2_Amp_F_I_1.OUT.n351 0.188181
R37892 C2S2_Amp_F_I_1.OUT.n365 C2S2_Amp_F_I_1.OUT.n364 0.188181
R37893 C2S2_Amp_F_I_1.OUT.n378 C2S2_Amp_F_I_1.OUT.n377 0.188181
R37894 C2S2_Amp_F_I_1.OUT.n391 C2S2_Amp_F_I_1.OUT.n390 0.188181
R37895 C2S2_Amp_F_I_1.OUT.n407 C2S2_Amp_F_I_1.OUT.n406 0.188181
R37896 C2S2_Amp_F_I_1.OUT.n68 C2S2_Amp_F_I_1.OUT.n63 0.186853
R37897 C2S2_Amp_F_I_1.OUT.n81 C2S2_Amp_F_I_1.OUT.n76 0.186853
R37898 C2S2_Amp_F_I_1.OUT.n94 C2S2_Amp_F_I_1.OUT.n89 0.186853
R37899 C2S2_Amp_F_I_1.OUT.n107 C2S2_Amp_F_I_1.OUT.n102 0.186853
R37900 C2S2_Amp_F_I_1.OUT.n120 C2S2_Amp_F_I_1.OUT.n115 0.186853
R37901 C2S2_Amp_F_I_1.OUT.n133 C2S2_Amp_F_I_1.OUT.n128 0.186853
R37902 C2S2_Amp_F_I_1.OUT.n146 C2S2_Amp_F_I_1.OUT.n141 0.186853
R37903 C2S2_Amp_F_I_1.OUT.n159 C2S2_Amp_F_I_1.OUT.n154 0.186853
R37904 C2S2_Amp_F_I_1.OUT.n172 C2S2_Amp_F_I_1.OUT.n167 0.186853
R37905 C2S2_Amp_F_I_1.OUT.n185 C2S2_Amp_F_I_1.OUT.n180 0.186853
R37906 C2S2_Amp_F_I_1.OUT.n198 C2S2_Amp_F_I_1.OUT.n193 0.186853
R37907 C2S2_Amp_F_I_1.OUT.n211 C2S2_Amp_F_I_1.OUT.n206 0.186853
R37908 C2S2_Amp_F_I_1.OUT.n224 C2S2_Amp_F_I_1.OUT.n219 0.186853
R37909 C2S2_Amp_F_I_1.OUT.n237 C2S2_Amp_F_I_1.OUT.n232 0.186853
R37910 C2S2_Amp_F_I_1.OUT.n250 C2S2_Amp_F_I_1.OUT.n245 0.186853
R37911 C2S2_Amp_F_I_1.OUT.n263 C2S2_Amp_F_I_1.OUT.n258 0.186853
R37912 C2S2_Amp_F_I_1.OUT.n276 C2S2_Amp_F_I_1.OUT.n271 0.186853
R37913 C2S2_Amp_F_I_1.OUT.n289 C2S2_Amp_F_I_1.OUT.n284 0.186853
R37914 C2S2_Amp_F_I_1.OUT.n301 C2S2_Amp_F_I_1.OUT.n298 0.186853
R37915 C2S2_Amp_F_I_1.OUT.n54 C2S2_Amp_F_I_1.OUT.n50 0.186853
R37916 C2S2_Amp_F_I_1.OUT.n10 C2S2_Amp_F_I_1.OUT.n1 0.158954
R37917 C2S2_Amp_F_I_1.OUT.n339 C2S2_Amp_F_I_1.OUT.n333 0.158954
R37918 C2S2_Amp_F_I_1.OUT.n352 C2S2_Amp_F_I_1.OUT.n346 0.158954
R37919 C2S2_Amp_F_I_1.OUT.n365 C2S2_Amp_F_I_1.OUT.n359 0.158954
R37920 C2S2_Amp_F_I_1.OUT.n378 C2S2_Amp_F_I_1.OUT.n372 0.158954
R37921 C2S2_Amp_F_I_1.OUT.n391 C2S2_Amp_F_I_1.OUT.n385 0.158954
R37922 C2S2_Amp_F_I_1.OUT.n407 C2S2_Amp_F_I_1.OUT.n398 0.158954
R37923 C2S2_Amp_F_I_1.OUT.n69 C2S2_Amp_F_I_1.OUT.n48 0.138785
R37924 C2S2_Amp_F_I_1.OUT.n82 C2S2_Amp_F_I_1.OUT.n47 0.138785
R37925 C2S2_Amp_F_I_1.OUT.n95 C2S2_Amp_F_I_1.OUT.n46 0.138785
R37926 C2S2_Amp_F_I_1.OUT.n108 C2S2_Amp_F_I_1.OUT.n45 0.138785
R37927 C2S2_Amp_F_I_1.OUT.n121 C2S2_Amp_F_I_1.OUT.n44 0.138785
R37928 C2S2_Amp_F_I_1.OUT.n134 C2S2_Amp_F_I_1.OUT.n43 0.138785
R37929 C2S2_Amp_F_I_1.OUT.n147 C2S2_Amp_F_I_1.OUT.n42 0.138785
R37930 C2S2_Amp_F_I_1.OUT.n160 C2S2_Amp_F_I_1.OUT.n41 0.138785
R37931 C2S2_Amp_F_I_1.OUT.n173 C2S2_Amp_F_I_1.OUT.n40 0.138785
R37932 C2S2_Amp_F_I_1.OUT.n186 C2S2_Amp_F_I_1.OUT.n39 0.138785
R37933 C2S2_Amp_F_I_1.OUT.n199 C2S2_Amp_F_I_1.OUT.n38 0.138785
R37934 C2S2_Amp_F_I_1.OUT.n212 C2S2_Amp_F_I_1.OUT.n37 0.138785
R37935 C2S2_Amp_F_I_1.OUT.n225 C2S2_Amp_F_I_1.OUT.n36 0.138785
R37936 C2S2_Amp_F_I_1.OUT.n238 C2S2_Amp_F_I_1.OUT.n35 0.138785
R37937 C2S2_Amp_F_I_1.OUT.n251 C2S2_Amp_F_I_1.OUT.n34 0.138785
R37938 C2S2_Amp_F_I_1.OUT.n264 C2S2_Amp_F_I_1.OUT.n33 0.138785
R37939 C2S2_Amp_F_I_1.OUT.n277 C2S2_Amp_F_I_1.OUT.n32 0.138785
R37940 C2S2_Amp_F_I_1.OUT.n290 C2S2_Amp_F_I_1.OUT.n31 0.138785
R37941 C2S2_Amp_F_I_1.OUT.n308 C2S2_Amp_F_I_1.OUT.n307 0.138785
R37942 C2S2_Amp_F_I_1.OUT.n61 C2S2_Amp_F_I_1.OUT.n60 0.138785
R37943 C2S2_Amp_F_I_1.OUT.n430 C2S2_Amp_F_I_1.OUT.n429 0.136017
R37944 C2S2_Amp_F_I_1.OUT.n27 C2S2_Amp_F_I_1.OUT.n26 0.130633
R37945 C2S2_Amp_F_I_1.OUT.n424 C2S2_Amp_F_I_1.OUT.n423 0.130633
R37946 C2S2_Amp_F_I_1.OUT.n322 C2S2_Amp_F_I_1.OUT.t10 0.114939
R37947 C2S2_Amp_F_I_1.OUT.n321 C2S2_Amp_F_I_1.OUT.t12 0.114939
R37948 C2S2_Amp_F_I_1.OUT.n320 C2S2_Amp_F_I_1.OUT.t5 0.114939
R37949 C2S2_Amp_F_I_1.OUT.n318 C2S2_Amp_F_I_1.OUT.t3 0.114939
R37950 C2S2_Amp_F_I_1.OUT.n317 C2S2_Amp_F_I_1.OUT.t9 0.114939
R37951 C2S2_Amp_F_I_1.OUT.n316 C2S2_Amp_F_I_1.OUT.t1 0.114939
R37952 C2S2_Amp_F_I_1.OUT.n315 C2S2_Amp_F_I_1.OUT.t2 0.114939
R37953 C2S2_Amp_F_I_1.OUT.n314 C2S2_Amp_F_I_1.OUT.t6 0.114939
R37954 C2S2_Amp_F_I_1.OUT.n313 C2S2_Amp_F_I_1.OUT.t8 0.114939
R37955 C2S2_Amp_F_I_1.OUT.n310 C2S2_Amp_F_I_1.OUT.n309 0.112608
R37956 C2S2_Amp_F_I_1.OUT.n62 C2S2_Amp_F_I_1.OUT.n29 0.112608
R37957 C2S2_Amp_F_I_1.OUT.n433 C2S2_Amp_F_I_1.OUT.n28 0.0831025
R37958 C2S2_Amp_F_I_1.OUT.n426 C2S2_Amp_F_I_1.OUT.n425 0.0817111
R37959 C2S2_Amp_F_I_1.OUT.n431 C2S2_Amp_F_I_1.OUT.t67 0.0712169
R37960 C2S2_Amp_F_I_1.OUT.n428 C2S2_Amp_F_I_1.OUT.t68 0.0699114
R37961 C2S2_Amp_F_I_1.OUT.n429 C2S2_Amp_F_I_1.OUT.n428 0.0695639
R37962 C2S2_Amp_F_I_1.OUT.n431 C2S2_Amp_F_I_1.OUT.n430 0.0682583
R37963 C2S2_Amp_F_I_1.OUT.n425 C2S2_Amp_F_I_1.OUT.n397 0.0616
R37964 C2S2_Amp_F_I_1.OUT.n397 C2S2_Amp_F_I_1.OUT.n384 0.0616
R37965 C2S2_Amp_F_I_1.OUT.n371 C2S2_Amp_F_I_1.OUT.n358 0.0616
R37966 C2S2_Amp_F_I_1.OUT.n345 C2S2_Amp_F_I_1.OUT.n28 0.0616
R37967 C2S2_Amp_F_I_1.OUT.n384 C2S2_Amp_F_I_1.OUT.n371 0.060425
R37968 C2S2_Amp_F_I_1.OUT.n358 C2S2_Amp_F_I_1.OUT.n345 0.060425
R37969 C2S2_Amp_F_I_1.OUT.n325 C2S2_Amp_F_I_1.OUT.n312 0.0502472
R37970 C2S2_Amp_F_I_1.OUT.n296 C2S2_Amp_F_I_1.OUT.n283 0.0460758
R37971 C2S2_Amp_F_I_1.OUT.n270 C2S2_Amp_F_I_1.OUT.n257 0.0460758
R37972 C2S2_Amp_F_I_1.OUT.n257 C2S2_Amp_F_I_1.OUT.n244 0.0460758
R37973 C2S2_Amp_F_I_1.OUT.n231 C2S2_Amp_F_I_1.OUT.n218 0.0460758
R37974 C2S2_Amp_F_I_1.OUT.n205 C2S2_Amp_F_I_1.OUT.n192 0.0460758
R37975 C2S2_Amp_F_I_1.OUT.n192 C2S2_Amp_F_I_1.OUT.n179 0.0460758
R37976 C2S2_Amp_F_I_1.OUT.n166 C2S2_Amp_F_I_1.OUT.n153 0.0460758
R37977 C2S2_Amp_F_I_1.OUT.n153 C2S2_Amp_F_I_1.OUT.n140 0.0460758
R37978 C2S2_Amp_F_I_1.OUT.n127 C2S2_Amp_F_I_1.OUT.n114 0.0460758
R37979 C2S2_Amp_F_I_1.OUT.n101 C2S2_Amp_F_I_1.OUT.n88 0.0460758
R37980 C2S2_Amp_F_I_1.OUT.n88 C2S2_Amp_F_I_1.OUT.n75 0.0460758
R37981 C2S2_Amp_F_I_1.OUT.n283 C2S2_Amp_F_I_1.OUT.n270 0.0446515
R37982 C2S2_Amp_F_I_1.OUT.n244 C2S2_Amp_F_I_1.OUT.n231 0.0446515
R37983 C2S2_Amp_F_I_1.OUT.n218 C2S2_Amp_F_I_1.OUT.n205 0.0446515
R37984 C2S2_Amp_F_I_1.OUT.n179 C2S2_Amp_F_I_1.OUT.n166 0.0446515
R37985 C2S2_Amp_F_I_1.OUT.n140 C2S2_Amp_F_I_1.OUT.n127 0.0446515
R37986 C2S2_Amp_F_I_1.OUT.n114 C2S2_Amp_F_I_1.OUT.n101 0.0446515
R37987 C2S2_Amp_F_I_1.OUT.n9 C2S2_Amp_F_I_1.OUT.n0 0.0407778
R37988 C2S2_Amp_F_I_1.OUT.n338 C2S2_Amp_F_I_1.OUT.n332 0.0407778
R37989 C2S2_Amp_F_I_1.OUT.n351 C2S2_Amp_F_I_1.OUT.n331 0.0407778
R37990 C2S2_Amp_F_I_1.OUT.n364 C2S2_Amp_F_I_1.OUT.n330 0.0407778
R37991 C2S2_Amp_F_I_1.OUT.n377 C2S2_Amp_F_I_1.OUT.n329 0.0407778
R37992 C2S2_Amp_F_I_1.OUT.n390 C2S2_Amp_F_I_1.OUT.n328 0.0407778
R37993 C2S2_Amp_F_I_1.OUT.n406 C2S2_Amp_F_I_1.OUT.n327 0.0407778
R37994 C2S2_Amp_F_I_1.OUT.n74 C2S2_Amp_F_I_1.OUT.n63 0.0393889
R37995 C2S2_Amp_F_I_1.OUT.n87 C2S2_Amp_F_I_1.OUT.n76 0.0393889
R37996 C2S2_Amp_F_I_1.OUT.n100 C2S2_Amp_F_I_1.OUT.n89 0.0393889
R37997 C2S2_Amp_F_I_1.OUT.n113 C2S2_Amp_F_I_1.OUT.n102 0.0393889
R37998 C2S2_Amp_F_I_1.OUT.n126 C2S2_Amp_F_I_1.OUT.n115 0.0393889
R37999 C2S2_Amp_F_I_1.OUT.n139 C2S2_Amp_F_I_1.OUT.n128 0.0393889
R38000 C2S2_Amp_F_I_1.OUT.n152 C2S2_Amp_F_I_1.OUT.n141 0.0393889
R38001 C2S2_Amp_F_I_1.OUT.n165 C2S2_Amp_F_I_1.OUT.n154 0.0393889
R38002 C2S2_Amp_F_I_1.OUT.n178 C2S2_Amp_F_I_1.OUT.n167 0.0393889
R38003 C2S2_Amp_F_I_1.OUT.n191 C2S2_Amp_F_I_1.OUT.n180 0.0393889
R38004 C2S2_Amp_F_I_1.OUT.n204 C2S2_Amp_F_I_1.OUT.n193 0.0393889
R38005 C2S2_Amp_F_I_1.OUT.n217 C2S2_Amp_F_I_1.OUT.n206 0.0393889
R38006 C2S2_Amp_F_I_1.OUT.n230 C2S2_Amp_F_I_1.OUT.n219 0.0393889
R38007 C2S2_Amp_F_I_1.OUT.n243 C2S2_Amp_F_I_1.OUT.n232 0.0393889
R38008 C2S2_Amp_F_I_1.OUT.n256 C2S2_Amp_F_I_1.OUT.n245 0.0393889
R38009 C2S2_Amp_F_I_1.OUT.n269 C2S2_Amp_F_I_1.OUT.n258 0.0393889
R38010 C2S2_Amp_F_I_1.OUT.n282 C2S2_Amp_F_I_1.OUT.n271 0.0393889
R38011 C2S2_Amp_F_I_1.OUT.n295 C2S2_Amp_F_I_1.OUT.n284 0.0393889
R38012 C2S2_Amp_F_I_1.OUT.n301 C2S2_Amp_F_I_1.OUT.n30 0.0393889
R38013 C2S2_Amp_F_I_1.OUT.n54 C2S2_Amp_F_I_1.OUT.n53 0.0393889
R38014 C2S2_Amp_F_I_1.OUT.n324 C2S2_Amp_F_I_1.OUT.n311 0.0148923
R38015 C2S2_Amp_F_I_1.OUT.n326 C2S2_Amp_F_I_1.OUT.n311 0.0148781
R38016 C2S2_Amp_F_I_1.OUT.n27 C2S2_Amp_F_I_1.OUT.n1 0.0102222
R38017 C2S2_Amp_F_I_1.OUT.n344 C2S2_Amp_F_I_1.OUT.n333 0.0102222
R38018 C2S2_Amp_F_I_1.OUT.n357 C2S2_Amp_F_I_1.OUT.n346 0.0102222
R38019 C2S2_Amp_F_I_1.OUT.n370 C2S2_Amp_F_I_1.OUT.n359 0.0102222
R38020 C2S2_Amp_F_I_1.OUT.n383 C2S2_Amp_F_I_1.OUT.n372 0.0102222
R38021 C2S2_Amp_F_I_1.OUT.n396 C2S2_Amp_F_I_1.OUT.n385 0.0102222
R38022 C2S2_Amp_F_I_1.OUT.n424 C2S2_Amp_F_I_1.OUT.n398 0.0102222
R38023 C2S2_Amp_F_I_1.OUT.n430 C2S2_Amp_F_I_1.OUT.t66 0.00345858
R38024 C2S2_Amp_F_I_1.OUT.n429 C2S2_Amp_F_I_1.OUT.t65 0.00345858
R38025 a_220333_n26938.n152 a_220333_n26938.n43 194.291
R38026 a_220333_n26938.n152 a_220333_n26938.n93 585
R38027 a_220333_n26938.n152 a_220333_n26938.n92 585
R38028 a_220333_n26938.n152 a_220333_n26938.n91 585
R38029 a_220333_n26938.n152 a_220333_n26938.n89 585
R38030 a_220333_n26938.n152 a_220333_n26938.n88 585
R38031 a_220333_n26938.n152 a_220333_n26938.n87 585
R38032 a_220333_n26938.n152 a_220333_n26938.n86 585
R38033 a_220333_n26938.n152 a_220333_n26938.n51 291.375
R38034 a_220333_n26938.n113 a_220333_n26938.n40 194.291
R38035 a_220333_n26938.n113 a_220333_n26938.n102 585
R38036 a_220333_n26938.n113 a_220333_n26938.n101 585
R38037 a_220333_n26938.n113 a_220333_n26938.n100 585
R38038 a_220333_n26938.n113 a_220333_n26938.n98 585
R38039 a_220333_n26938.n113 a_220333_n26938.n97 585
R38040 a_220333_n26938.n113 a_220333_n26938.n96 585
R38041 a_220333_n26938.n113 a_220333_n26938.n95 585
R38042 a_220333_n26938.n113 a_220333_n26938.n94 585
R38043 a_220333_n26938.n113 a_220333_n26938.n50 585
R38044 a_220333_n26938.n157 a_220333_n26938.n39 194.291
R38045 a_220333_n26938.n157 a_220333_n26938.n65 585
R38046 a_220333_n26938.n157 a_220333_n26938.n64 585
R38047 a_220333_n26938.n157 a_220333_n26938.n66 585
R38048 a_220333_n26938.n157 a_220333_n26938.n62 585
R38049 a_220333_n26938.n157 a_220333_n26938.n67 585
R38050 a_220333_n26938.n157 a_220333_n26938.n61 585
R38051 a_220333_n26938.n157 a_220333_n26938.n68 585
R38052 a_220333_n26938.n157 a_220333_n26938.n60 585
R38053 a_220333_n26938.n157 a_220333_n26938.n156 585
R38054 a_220333_n26938.t3 a_220333_n26938.n9 308.31
R38055 a_220333_n26938.n135 a_220333_n26938.t3 308.31
R38056 a_220333_n26938.t1 a_220333_n26938.n142 308.31
R38057 a_220333_n26938.n9 a_220333_n26938.t1 308.31
R38058 a_220333_n26938.n152 a_220333_n26938.n90 286.238
R38059 a_220333_n26938.n113 a_220333_n26938.n99 286.238
R38060 a_220333_n26938.n157 a_220333_n26938.n63 286.238
R38061 a_220333_n26938.n57 a_220333_n26938.n56 6.98494
R38062 a_220333_n26938.n59 a_220333_n26938.n58 6.98494
R38063 a_220333_n26938.n55 a_220333_n26938.t22 104.094
R38064 a_220333_n26938.n4 a_220333_n26938.t9 209.939
R38065 a_220333_n26938.t11 a_220333_n26938.n6 209.938
R38066 a_220333_n26938.t26 a_220333_n26938.n53 104.094
R38067 a_220333_n26938.t13 a_220333_n26938.n14 209.93
R38068 a_220333_n26938.n10 a_220333_n26938.t13 209.93
R38069 a_220333_n26938.t7 a_220333_n26938.n128 209.93
R38070 a_220333_n26938.n2 a_220333_n26938.t7 209.93
R38071 a_220333_n26938.n1 a_220333_n26938.t11 209.93
R38072 a_220333_n26938.t15 a_220333_n26938.n0 209.93
R38073 a_220333_n26938.n85 a_220333_n26938.t15 209.93
R38074 a_220333_n26938.n15 a_220333_n26938.t5 209.93
R38075 a_220333_n26938.t5 a_220333_n26938.n12 209.93
R38076 a_220333_n26938.n155 a_220333_n26938.t25 209.93
R38077 a_220333_n26938.t25 a_220333_n26938.n154 209.93
R38078 a_220333_n26938.t24 a_220333_n26938.n84 209.93
R38079 a_220333_n26938.n153 a_220333_n26938.t24 209.93
R38080 a_220333_n26938.n114 a_220333_n26938.t27 209.93
R38081 a_220333_n26938.t27 a_220333_n26938.n11 209.93
R38082 a_220333_n26938.t23 a_220333_n26938.n115 209.93
R38083 a_220333_n26938.n116 a_220333_n26938.t23 209.93
R38084 a_220333_n26938.t9 a_220333_n26938.n127 209.93
R38085 a_220333_n26938.n134 a_220333_n26938.n49 92.3135
R38086 a_220333_n26938.n134 a_220333_n26938.n130 185
R38087 a_220333_n26938.n134 a_220333_n26938.n21 92.3135
R38088 a_220333_n26938.n141 a_220333_n26938.n46 92.3135
R38089 a_220333_n26938.n141 a_220333_n26938.n137 185
R38090 a_220333_n26938.n141 a_220333_n26938.n18 92.3135
R38091 a_220333_n26938.n125 a_220333_n26938.n124 185
R38092 a_220333_n26938.n121 a_220333_n26938.n120 185
R38093 a_220333_n26938.n75 a_220333_n26938.n74 185
R38094 a_220333_n26938.n71 a_220333_n26938.n70 185
R38095 a_220333_n26938.n122 a_220333_n26938.t20 174.857
R38096 a_220333_n26938.n72 a_220333_n26938.t0 174.857
R38097 a_220333_n26938.n57 a_220333_n26938.n125 244.714
R38098 a_220333_n26938.n125 a_220333_n26938.n120 140.69
R38099 a_220333_n26938.n59 a_220333_n26938.n75 244.714
R38100 a_220333_n26938.n75 a_220333_n26938.n70 140.69
R38101 a_220333_n26938.n134 a_220333_n26938.n129 86.5152
R38102 a_220333_n26938.n141 a_220333_n26938.n136 86.5152
R38103 a_220333_n26938.t20 a_220333_n26938.n120 70.3453
R38104 a_220333_n26938.t0 a_220333_n26938.n70 70.3453
R38105 a_220333_n26938.n122 a_220333_n26938.n121 28.4333
R38106 a_220333_n26938.n72 a_220333_n26938.n71 28.4333
R38107 a_220333_n26938.n132 a_220333_n26938.n130 25.6005
R38108 a_220333_n26938.n139 a_220333_n26938.n137 25.6005
R38109 a_220333_n26938.n148 a_220333_n26938.n91 24.8476
R38110 a_220333_n26938.n147 a_220333_n26938.n89 24.8476
R38111 a_220333_n26938.n109 a_220333_n26938.n100 24.8476
R38112 a_220333_n26938.n108 a_220333_n26938.n98 24.8476
R38113 a_220333_n26938.n124 a_220333_n26938.n123 24.8476
R38114 a_220333_n26938.n74 a_220333_n26938.n73 24.8476
R38115 a_220333_n26938.n81 a_220333_n26938.n66 24.8476
R38116 a_220333_n26938.n80 a_220333_n26938.n62 24.8476
R38117 a_220333_n26938.n131 a_220333_n26938.n21 27.7565
R38118 a_220333_n26938.n138 a_220333_n26938.n18 27.7565
R38119 a_220333_n26938.n149 a_220333_n26938.n92 23.3417
R38120 a_220333_n26938.n146 a_220333_n26938.n88 23.3417
R38121 a_220333_n26938.n110 a_220333_n26938.n101 23.3417
R38122 a_220333_n26938.n107 a_220333_n26938.n97 23.3417
R38123 a_220333_n26938.n82 a_220333_n26938.n64 23.3417
R38124 a_220333_n26938.n79 a_220333_n26938.n67 23.3417
R38125 a_220333_n26938.n49 a_220333_n26938.n48 6.60954
R38126 a_220333_n26938.n21 a_220333_n26938.n19 6.60954
R38127 a_220333_n26938.n46 a_220333_n26938.n45 6.60954
R38128 a_220333_n26938.n18 a_220333_n26938.n16 6.60954
R38129 a_220333_n26938.n8 a_220333_n26938.n117 22.3909
R38130 a_220333_n26938.n8 a_220333_n26938.n118 22.3909
R38131 a_220333_n26938.n150 a_220333_n26938.n93 21.8358
R38132 a_220333_n26938.n145 a_220333_n26938.n87 21.8358
R38133 a_220333_n26938.n111 a_220333_n26938.n102 21.8358
R38134 a_220333_n26938.n106 a_220333_n26938.n96 21.8358
R38135 a_220333_n26938.n83 a_220333_n26938.n65 21.8358
R38136 a_220333_n26938.n78 a_220333_n26938.n61 21.8358
R38137 a_220333_n26938.n144 a_220333_n26938.n86 20.3299
R38138 a_220333_n26938.n105 a_220333_n26938.n95 20.3299
R38139 a_220333_n26938.n77 a_220333_n26938.n68 20.3299
R38140 a_220333_n26938.n2 a_220333_n26938.n50 19.0887
R38141 a_220333_n26938.n156 a_220333_n26938.n1 19.0887
R38142 a_220333_n26938.n43 a_220333_n26938.n13 6.07169
R38143 a_220333_n26938.n143 a_220333_n26938.n51 24.6333
R38144 a_220333_n26938.n40 a_220333_n26938.n3 6.07169
R38145 a_220333_n26938.n104 a_220333_n26938.n94 18.824
R38146 a_220333_n26938.n5 a_220333_n26938.n39 6.07169
R38147 a_220333_n26938.n76 a_220333_n26938.n60 18.824
R38148 a_220333_n26938.n10 a_220333_n26938.n51 9.76605
R38149 a_220333_n26938.n103 a_220333_n26938.n50 17.3181
R38150 a_220333_n26938.n156 a_220333_n26938.n41 17.3181
R38151 a_220333_n26938.n131 a_220333_n26938.n129 13.4786
R38152 a_220333_n26938.n138 a_220333_n26938.n136 13.4786
R38153 a_220333_n26938.n148 a_220333_n26938.n90 13.2799
R38154 a_220333_n26938.n147 a_220333_n26938.n90 13.2799
R38155 a_220333_n26938.n109 a_220333_n26938.n99 13.2799
R38156 a_220333_n26938.n108 a_220333_n26938.n99 13.2799
R38157 a_220333_n26938.n81 a_220333_n26938.n63 13.2799
R38158 a_220333_n26938.n80 a_220333_n26938.n63 13.2799
R38159 a_220333_n26938.n132 a_220333_n26938.n129 11.9727
R38160 a_220333_n26938.n139 a_220333_n26938.n136 11.9727
R38161 a_220333_n26938.n10 a_220333_n26938.n9 9.61161
R38162 a_220333_n26938.n6 a_220333_n26938.n52 9.47511
R38163 a_220333_n26938.n4 a_220333_n26938.n54 9.47106
R38164 a_220333_n26938.n11 a_220333_n26938.n14 9.3755
R38165 a_220333_n26938.n44 a_220333_n26938.n140 9.3005
R38166 a_220333_n26938.n17 a_220333_n26938.n139 9.3005
R38167 a_220333_n26938.n17 a_220333_n26938.n138 9.3005
R38168 a_220333_n26938.n47 a_220333_n26938.n133 9.3005
R38169 a_220333_n26938.n20 a_220333_n26938.n132 9.3005
R38170 a_220333_n26938.n20 a_220333_n26938.n131 9.3005
R38171 a_220333_n26938.n123 a_220333_n26938.n22 9.3005
R38172 a_220333_n26938.n119 a_220333_n26938.n22 9.3005
R38173 a_220333_n26938.n73 a_220333_n26938.n23 9.3005
R38174 a_220333_n26938.n69 a_220333_n26938.n23 9.3005
R38175 a_220333_n26938.n28 a_220333_n26938.n103 9.3005
R38176 a_220333_n26938.n24 a_220333_n26938.n109 9.3005
R38177 a_220333_n26938.n24 a_220333_n26938.n110 9.3005
R38178 a_220333_n26938.n25 a_220333_n26938.n111 9.3005
R38179 a_220333_n26938.n25 a_220333_n26938.n112 9.3005
R38180 a_220333_n26938.n26 a_220333_n26938.n108 9.3005
R38181 a_220333_n26938.n26 a_220333_n26938.n107 9.3005
R38182 a_220333_n26938.n27 a_220333_n26938.n106 9.3005
R38183 a_220333_n26938.n27 a_220333_n26938.n105 9.3005
R38184 a_220333_n26938.n28 a_220333_n26938.n104 9.3005
R38185 a_220333_n26938.n29 a_220333_n26938.n148 9.3005
R38186 a_220333_n26938.n30 a_220333_n26938.n149 9.3005
R38187 a_220333_n26938.n30 a_220333_n26938.n150 9.3005
R38188 a_220333_n26938.n42 a_220333_n26938.n151 9.3005
R38189 a_220333_n26938.n29 a_220333_n26938.n147 9.3005
R38190 a_220333_n26938.n31 a_220333_n26938.n146 9.3005
R38191 a_220333_n26938.n31 a_220333_n26938.n145 9.3005
R38192 a_220333_n26938.n32 a_220333_n26938.n144 9.3005
R38193 a_220333_n26938.n32 a_220333_n26938.n143 9.3005
R38194 a_220333_n26938.n33 a_220333_n26938.n81 9.3005
R38195 a_220333_n26938.n33 a_220333_n26938.n82 9.3005
R38196 a_220333_n26938.n34 a_220333_n26938.n83 9.3005
R38197 a_220333_n26938.n34 a_220333_n26938.n38 9.3005
R38198 a_220333_n26938.n35 a_220333_n26938.n80 9.3005
R38199 a_220333_n26938.n35 a_220333_n26938.n79 9.3005
R38200 a_220333_n26938.n36 a_220333_n26938.n78 9.3005
R38201 a_220333_n26938.n36 a_220333_n26938.n77 9.3005
R38202 a_220333_n26938.n37 a_220333_n26938.n76 9.3005
R38203 a_220333_n26938.n37 a_220333_n26938.n41 9.3005
R38204 a_220333_n26938.n103 a_220333_n26938.n94 8.28285
R38205 a_220333_n26938.n41 a_220333_n26938.n60 8.28285
R38206 a_220333_n26938.n1 a_220333_n26938.n7 7.04926
R38207 a_220333_n26938.n127 a_220333_n26938.n126 6.96926
R38208 a_220333_n26938.n134 a_220333_n26938.t4 6.9605
R38209 a_220333_n26938.n141 a_220333_n26938.t2 6.9605
R38210 a_220333_n26938.n43 a_220333_n26938.n151 28.1963
R38211 a_220333_n26938.n143 a_220333_n26938.n86 6.77697
R38212 a_220333_n26938.n40 a_220333_n26938.n112 28.1963
R38213 a_220333_n26938.n104 a_220333_n26938.n95 6.77697
R38214 a_220333_n26938.n39 a_220333_n26938.n38 28.1963
R38215 a_220333_n26938.n76 a_220333_n26938.n68 6.77697
R38216 a_220333_n26938.n152 a_220333_n26938.t14 5.7135
R38217 a_220333_n26938.n152 a_220333_n26938.t6 5.7135
R38218 a_220333_n26938.n113 a_220333_n26938.t10 5.7135
R38219 a_220333_n26938.n113 a_220333_n26938.t8 5.7135
R38220 a_220333_n26938.t16 a_220333_n26938.n157 5.7135
R38221 a_220333_n26938.n157 a_220333_n26938.t12 5.7135
R38222 a_220333_n26938.n22 a_220333_n26938.n122 5.33935
R38223 a_220333_n26938.n23 a_220333_n26938.n72 5.33935
R38224 a_220333_n26938.n151 a_220333_n26938.n93 5.27109
R38225 a_220333_n26938.n144 a_220333_n26938.n87 5.27109
R38226 a_220333_n26938.n112 a_220333_n26938.n102 5.27109
R38227 a_220333_n26938.n105 a_220333_n26938.n96 5.27109
R38228 a_220333_n26938.n38 a_220333_n26938.n65 5.27109
R38229 a_220333_n26938.n77 a_220333_n26938.n61 5.27109
R38230 a_220333_n26938.n7 a_220333_n26938.n58 4.5005
R38231 a_220333_n26938.n126 a_220333_n26938.n56 4.5005
R38232 a_220333_n26938.n150 a_220333_n26938.n92 3.76521
R38233 a_220333_n26938.n145 a_220333_n26938.n88 3.76521
R38234 a_220333_n26938.n111 a_220333_n26938.n101 3.76521
R38235 a_220333_n26938.n106 a_220333_n26938.n97 3.76521
R38236 a_220333_n26938.n57 a_220333_n26938.n119 27.242
R38237 a_220333_n26938.n59 a_220333_n26938.n69 27.242
R38238 a_220333_n26938.n83 a_220333_n26938.n64 3.76521
R38239 a_220333_n26938.n78 a_220333_n26938.n67 3.76521
R38240 a_220333_n26938.n8 a_220333_n26938.n7 3.716
R38241 a_220333_n26938.n52 a_220333_n26938.n53 1.75048
R38242 a_220333_n26938.n54 a_220333_n26938.n55 1.74802
R38243 a_220333_n26938.n117 a_220333_n26938.t19 3.4805
R38244 a_220333_n26938.n117 a_220333_n26938.t18 3.4805
R38245 a_220333_n26938.n118 a_220333_n26938.t21 3.4805
R38246 a_220333_n26938.n118 a_220333_n26938.t17 3.4805
R38247 a_220333_n26938.n49 a_220333_n26938.n133 27.7565
R38248 a_220333_n26938.n46 a_220333_n26938.n140 27.7565
R38249 a_220333_n26938.n126 a_220333_n26938.n8 4.01562
R38250 a_220333_n26938.n149 a_220333_n26938.n91 2.25932
R38251 a_220333_n26938.n146 a_220333_n26938.n89 2.25932
R38252 a_220333_n26938.n110 a_220333_n26938.n100 2.25932
R38253 a_220333_n26938.n107 a_220333_n26938.n98 2.25932
R38254 a_220333_n26938.n124 a_220333_n26938.n119 2.25932
R38255 a_220333_n26938.n74 a_220333_n26938.n69 2.25932
R38256 a_220333_n26938.n82 a_220333_n26938.n66 2.25932
R38257 a_220333_n26938.n79 a_220333_n26938.n62 2.25932
R38258 a_220333_n26938.n133 a_220333_n26938.n130 1.50638
R38259 a_220333_n26938.n140 a_220333_n26938.n137 1.50638
R38260 a_220333_n26938.n123 a_220333_n26938.n121 0.753441
R38261 a_220333_n26938.n73 a_220333_n26938.n71 0.753441
R38262 a_220333_n26938.n54 a_220333_n26938.n116 0.726434
R38263 a_220333_n26938.n12 a_220333_n26938.n85 0.645765
R38264 a_220333_n26938.n116 a_220333_n26938.n11 0.645765
R38265 a_220333_n26938.n154 a_220333_n26938.n153 0.645765
R38266 a_220333_n26938.n115 a_220333_n26938.n55 2.39323
R38267 a_220333_n26938.n154 a_220333_n26938.n52 0.731421
R38268 a_220333_n26938.n115 a_220333_n26938.n114 0.645765
R38269 a_220333_n26938.n114 a_220333_n26938.n84 0.645765
R38270 a_220333_n26938.n155 a_220333_n26938.n84 0.645765
R38271 a_220333_n26938.n53 a_220333_n26938.n155 2.39569
R38272 a_220333_n26938.n48 a_220333_n26938.n9 0.658
R38273 a_220333_n26938.n32 a_220333_n26938.n10 0.649958
R38274 a_220333_n26938.n10 a_220333_n26938.n2 0.645765
R38275 a_220333_n26938.n128 a_220333_n26938.n14 0.645765
R38276 a_220333_n26938.n15 a_220333_n26938.n0 0.645765
R38277 a_220333_n26938.n127 a_220333_n26938.n2 0.645765
R38278 a_220333_n26938.n1 a_220333_n26938.n0 0.645765
R38279 a_220333_n26938.n85 a_220333_n26938.n6 0.631808
R38280 a_220333_n26938.n128 a_220333_n26938.n4 0.630877
R38281 a_220333_n26938.n5 a_220333_n26938.n34 0.584196
R38282 a_220333_n26938.n3 a_220333_n26938.n25 0.584196
R38283 a_220333_n26938.n14 a_220333_n26938.n12 0.56139
R38284 a_220333_n26938.n153 a_220333_n26938.n11 0.56139
R38285 a_220333_n26938.n10 a_220333_n26938.n15 0.446618
R38286 a_220333_n26938.n58 a_220333_n26938.n23 0.411505
R38287 a_220333_n26938.n56 a_220333_n26938.n22 0.411505
R38288 a_220333_n26938.n142 a_220333_n26938.n135 0.3955
R38289 a_220333_n26938.n35 a_220333_n26938.n36 0.391804
R38290 a_220333_n26938.n33 a_220333_n26938.n35 0.391804
R38291 a_220333_n26938.n34 a_220333_n26938.n33 0.391804
R38292 a_220333_n26938.n31 a_220333_n26938.n32 0.391804
R38293 a_220333_n26938.n29 a_220333_n26938.n31 0.391804
R38294 a_220333_n26938.n30 a_220333_n26938.n29 0.391804
R38295 a_220333_n26938.n42 a_220333_n26938.n30 0.391804
R38296 a_220333_n26938.n26 a_220333_n26938.n27 0.391804
R38297 a_220333_n26938.n24 a_220333_n26938.n26 0.391804
R38298 a_220333_n26938.n25 a_220333_n26938.n24 0.391804
R38299 a_220333_n26938.n20 a_220333_n26938.n19 0.391804
R38300 a_220333_n26938.n47 a_220333_n26938.n20 0.391804
R38301 a_220333_n26938.n17 a_220333_n26938.n16 0.391804
R38302 a_220333_n26938.n44 a_220333_n26938.n17 0.391804
R38303 a_220333_n26938.n36 a_220333_n26938.n37 0.388109
R38304 a_220333_n26938.n27 a_220333_n26938.n28 0.388109
R38305 a_220333_n26938.n13 a_220333_n26938.n42 0.387101
R38306 a_220333_n26938.n142 a_220333_n26938.n16 0.368217
R38307 a_220333_n26938.n135 a_220333_n26938.n19 0.368217
R38308 a_220333_n26938.n48 a_220333_n26938.n47 0.364413
R38309 a_220333_n26938.n45 a_220333_n26938.n44 0.364413
R38310 a_220333_n26938.n9 a_220333_n26938.n45 0.363
R38311 a_220333_n26938.n4 a_220333_n26938.n3 0.363
R38312 a_220333_n26938.n6 a_220333_n26938.n5 0.363
R38313 a_220333_n26938.n1 a_220333_n26938.n37 0.358
R38314 a_220333_n26938.n28 a_220333_n26938.n2 0.358
R38315 a_220333_n26938.n14 a_220333_n26938.n13 0.353
R38316 a_218222_n27786.n5 a_218222_n27786.n4 22.4024
R38317 a_218222_n27786.n3 a_218222_n27786.n2 18.9924
R38318 a_218222_n27786.n7 a_218222_n27786.n6 18.9924
R38319 a_218222_n27786.n5 a_218222_n27786.n3 3.716
R38320 a_218222_n27786.n7 a_218222_n27786.n5 3.71013
R38321 a_218222_n27786.n6 a_218222_n27786.t7 3.4805
R38322 a_218222_n27786.n6 a_218222_n27786.t9 3.4805
R38323 a_218222_n27786.n2 a_218222_n27786.t4 3.4805
R38324 a_218222_n27786.n2 a_218222_n27786.t1 3.4805
R38325 a_218222_n27786.n4 a_218222_n27786.t3 3.4805
R38326 a_218222_n27786.n4 a_218222_n27786.t6 3.4805
R38327 a_218222_n27786.n0 a_218222_n27786.t2 3.04088
R38328 a_218222_n27786.n9 a_218222_n27786.t8 3.03453
R38329 a_218222_n27786.t0 a_218222_n27786.n9 2.59519
R38330 a_218222_n27786.n0 a_218222_n27786.t5 2.59419
R38331 a_218222_n27786.n3 a_218222_n27786.n1 2.55108
R38332 a_218222_n27786.n8 a_218222_n27786.n7 2.55108
R38333 a_218222_n27786.n8 a_218222_n27786.n1 0.293114
R38334 a_218222_n27786.n1 a_218222_n27786.n0 0.078625
R38335 a_218222_n27786.n9 a_218222_n27786.n8 0.0672614
R38336 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t39 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n95 210.794
R38337 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t43 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n99 210.794
R38338 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n98 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t35 210.794
R38339 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t35 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n97 210.794
R38340 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t46 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n20 210.794
R38341 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n96 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t46 210.794
R38342 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n53 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t27 210.794
R38343 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t27 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n30 210.794
R38344 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n52 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t23 210.794
R38345 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t23 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n51 210.794
R38346 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t16 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n31 210.794
R38347 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n50 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t16 210.794
R38348 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t45 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n48 210.794
R38349 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n49 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t45 210.794
R38350 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n47 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t31 210.794
R38351 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t31 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n32 210.794
R38352 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n46 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t21 210.794
R38353 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t21 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n45 210.794
R38354 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t33 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n33 210.794
R38355 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n44 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t33 210.794
R38356 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t25 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n42 210.794
R38357 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n43 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t25 210.794
R38358 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n41 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t18 210.794
R38359 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t18 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n34 210.794
R38360 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n40 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t38 210.794
R38361 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t38 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n39 210.794
R38362 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t44 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n35 210.794
R38363 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n38 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t44 210.794
R38364 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n37 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t42 210.794
R38365 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t42 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n36 210.794
R38366 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t32 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n29 210.794
R38367 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n54 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t32 210.794
R38368 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n56 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t22 210.794
R38369 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t22 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n55 210.794
R38370 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n57 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t19 210.794
R38371 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t19 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n28 210.794
R38372 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t47 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n58 210.794
R38373 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n59 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t47 210.794
R38374 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t28 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n27 210.794
R38375 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n60 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t28 210.794
R38376 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n62 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t24 210.794
R38377 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t24 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n61 210.794
R38378 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n63 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t17 210.794
R38379 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t17 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n26 210.794
R38380 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t29 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n64 210.794
R38381 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n65 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t29 210.794
R38382 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t20 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n25 210.794
R38383 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n66 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t20 210.794
R38384 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n68 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t41 210.794
R38385 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t41 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n67 210.794
R38386 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n69 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t34 210.794
R38387 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t34 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n24 210.794
R38388 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t40 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n70 210.794
R38389 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n71 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t40 210.794
R38390 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t37 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n23 210.794
R38391 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n72 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t37 210.794
R38392 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n74 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t30 210.794
R38393 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t30 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n73 210.794
R38394 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n15 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n14 185
R38395 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n84 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n83 185
R38396 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t6 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n100 120.469
R38397 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n93 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t0 120.465
R38398 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n87 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t2 120.419
R38399 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t2 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n22 120.419
R38400 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n91 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t4 120.419
R38401 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t4 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n90 120.419
R38402 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n101 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t6 120.419
R38403 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n79 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t0 120.419
R38404 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n94 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t36 104.566
R38405 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n19 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t26 104.562
R38406 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n16 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n15 86.5152
R38407 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n83 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n82 86.5152
R38408 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n8 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n7 50.9993
R38409 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n78 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n77 47.5895
R38410 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n102 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n9 47.5893
R38411 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n89 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n88 38.0154
R38412 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n14 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n12 25.6005
R38413 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n84 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n81 25.6005
R38414 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n17 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n16 22.7786
R38415 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n82 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n21 22.7786
R38416 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t39 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n6 210.808
R38417 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n5 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n6 0.0650981
R38418 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n4 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n3 0.0650981
R38419 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n4 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t43 210.808
R38420 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n15 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t3 13.9205
R38421 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n15 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t7 13.9205
R38422 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n83 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t1 13.9205
R38423 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n83 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t5 13.9205
R38424 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n16 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n12 11.9727
R38425 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n82 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n81 11.9727
R38426 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n14 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n13 10.8064
R38427 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n85 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n84 10.8064
R38428 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n5 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n93 9.59564
R38429 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n100 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n3 9.59208
R38430 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n81 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n80 9.3005
R38431 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n12 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n11 9.3005
R38432 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n79 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n78 8.93258
R38433 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n102 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n101 8.84758
R38434 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n88 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t9 6.9605
R38435 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n88 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t8 6.9605
R38436 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n9 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t12 5.7135
R38437 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n9 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t11 5.7135
R38438 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n7 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t10 5.7135
R38439 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n7 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t13 5.7135
R38440 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n77 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t15 5.7135
R38441 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n77 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t14 5.7135
R38442 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n1 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n30 4.293
R38443 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n37 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n2 4.218
R38444 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n1 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n53 3.94612
R38445 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n36 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n2 3.87112
R38446 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n103 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n102 3.4105
R38447 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n78 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n76 3.4105
R38448 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n29 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n0 3.29712
R38449 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n54 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n1 3.29612
R38450 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n73 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n2 3.23112
R38451 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n75 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n74 3.23112
R38452 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n99 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n19 2.3168
R38453 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n103 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n0 2.31333
R38454 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n95 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n94 2.31188
R38455 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n76 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n75 2.30692
R38456 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n94 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n6 2.28563
R38457 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n97 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n96 0.645765
R38458 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n95 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n20 0.645765
R38459 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n98 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n20 0.645765
R38460 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n99 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n98 0.645765
R38461 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n91 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n22 0.645765
R38462 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n38 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n37 0.645765
R38463 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n39 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n38 0.645765
R38464 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n39 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n34 0.645765
R38465 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n43 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n34 0.645765
R38466 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n44 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n43 0.645765
R38467 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n45 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n44 0.645765
R38468 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n45 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n32 0.645765
R38469 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n49 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n32 0.645765
R38470 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n50 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n49 0.645765
R38471 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n51 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n50 0.645765
R38472 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n51 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n30 0.645765
R38473 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n36 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n35 0.645765
R38474 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n40 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n35 0.645765
R38475 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n41 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n40 0.645765
R38476 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n42 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n41 0.645765
R38477 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n42 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n33 0.645765
R38478 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n46 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n33 0.645765
R38479 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n47 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n46 0.645765
R38480 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n48 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n47 0.645765
R38481 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n48 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n31 0.645765
R38482 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n52 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n31 0.645765
R38483 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n53 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n52 0.645765
R38484 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n73 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n72 0.645765
R38485 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n72 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n71 0.645765
R38486 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n71 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n24 0.645765
R38487 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n67 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n24 0.645765
R38488 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n67 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n66 0.645765
R38489 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n66 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n65 0.645765
R38490 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n65 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n26 0.645765
R38491 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n61 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n26 0.645765
R38492 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n61 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n60 0.645765
R38493 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n60 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n59 0.645765
R38494 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n59 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n28 0.645765
R38495 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n55 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n28 0.645765
R38496 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n55 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n54 0.645765
R38497 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n74 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n23 0.645765
R38498 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n70 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n23 0.645765
R38499 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n70 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n69 0.645765
R38500 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n69 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n68 0.645765
R38501 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n68 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n25 0.645765
R38502 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n64 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n25 0.645765
R38503 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n64 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n63 0.645765
R38504 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n63 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n62 0.645765
R38505 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n62 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n27 0.645765
R38506 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n58 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n27 0.645765
R38507 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n58 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n57 0.645765
R38508 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n57 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n56 0.645765
R38509 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n56 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n29 0.645765
R38510 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n97 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n3 0.552061
R38511 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n96 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n5 0.550633
R38512 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n90 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n86 0.333133
R38513 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n92 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n91 0.333133
R38514 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n22 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n18 0.323133
R38515 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n87 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n10 0.323133
R38516 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n101 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n10 0.323133
R38517 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n86 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n79 0.313133
R38518 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n89 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n87 0.278133
R38519 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n90 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n89 0.268133
R38520 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n100 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n18 0.256274
R38521 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n93 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n92 0.252692
R38522 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n86 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n85 0.219522
R38523 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n18 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n17 0.217348
R38524 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n13 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n10 0.217348
R38525 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n92 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n21 0.216386
R38526 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n103 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n8 0.204167
R38527 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n76 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n8 0.204167
R38528 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n85 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n80 0.196152
R38529 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n80 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n21 0.196152
R38530 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n13 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n11 0.196152
R38531 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n17 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n11 0.196152
R38532 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n4 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n19 2.28913
R38533 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n75 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n2 0.4755
R38534 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n1 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n0 0.4755
R38535 1Bit_DAC_Inv_0.OUT.n1 1Bit_DAC_Inv_0.OUT.t38 57.0195
R38536 1Bit_DAC_Inv_0.OUT.n55 1Bit_DAC_Inv_0.OUT.t50 56.9568
R38537 1Bit_DAC_Inv_0.OUT.n33 1Bit_DAC_Inv_0.OUT.n32 50.4558
R38538 1Bit_DAC_Inv_0.OUT.n35 1Bit_DAC_Inv_0.OUT.n34 50.4558
R38539 1Bit_DAC_Inv_0.OUT.n52 1Bit_DAC_Inv_0.OUT.n51 50.4558
R38540 1Bit_DAC_Inv_0.OUT.n11 1Bit_DAC_Inv_0.OUT.n10 50.4558
R38541 1Bit_DAC_Inv_0.OUT.n9 1Bit_DAC_Inv_0.OUT.n8 50.4558
R38542 1Bit_DAC_Inv_0.OUT.n31 1Bit_DAC_Inv_0.OUT.n30 50.438
R38543 1Bit_DAC_Inv_0.OUT.n37 1Bit_DAC_Inv_0.OUT.n36 50.438
R38544 1Bit_DAC_Inv_0.OUT.n48 1Bit_DAC_Inv_0.OUT.n47 50.438
R38545 1Bit_DAC_Inv_0.OUT.n17 1Bit_DAC_Inv_0.OUT.n16 50.438
R38546 1Bit_DAC_Inv_0.OUT.n13 1Bit_DAC_Inv_0.OUT.n12 50.438
R38547 1Bit_DAC_Inv_0.OUT.n7 1Bit_DAC_Inv_0.OUT.n6 50.438
R38548 1Bit_DAC_Inv_0.OUT.n5 1Bit_DAC_Inv_0.OUT.n4 50.438
R38549 1Bit_DAC_Inv_0.OUT.n1 1Bit_DAC_Inv_0.OUT.n0 50.438
R38550 1Bit_DAC_Inv_0.OUT.n29 1Bit_DAC_Inv_0.OUT.n28 50.4246
R38551 1Bit_DAC_Inv_0.OUT.n40 1Bit_DAC_Inv_0.OUT.n39 50.4246
R38552 1Bit_DAC_Inv_0.OUT.n44 1Bit_DAC_Inv_0.OUT.n43 50.4246
R38553 1Bit_DAC_Inv_0.OUT.n15 1Bit_DAC_Inv_0.OUT.n14 50.4246
R38554 1Bit_DAC_Inv_0.OUT.n3 1Bit_DAC_Inv_0.OUT.n2 50.4246
R38555 1Bit_DAC_Inv_0.OUT.n38 1Bit_DAC_Inv_0.OUT.t17 25.1211
R38556 1Bit_DAC_Inv_0.OUT.n25 1Bit_DAC_Inv_0.OUT.t0 25.1211
R38557 1Bit_DAC_Inv_0.OUT.n20 1Bit_DAC_Inv_0.OUT.n18 21.23
R38558 1Bit_DAC_Inv_0.OUT.n42 1Bit_DAC_Inv_0.OUT.n41 21.179
R38559 1Bit_DAC_Inv_0.OUT.n50 1Bit_DAC_Inv_0.OUT.n49 21.179
R38560 1Bit_DAC_Inv_0.OUT.n54 1Bit_DAC_Inv_0.OUT.n53 21.179
R38561 1Bit_DAC_Inv_0.OUT.n24 1Bit_DAC_Inv_0.OUT.n23 21.179
R38562 1Bit_DAC_Inv_0.OUT.n20 1Bit_DAC_Inv_0.OUT.n19 21.179
R38563 1Bit_DAC_Inv_0.OUT.n46 1Bit_DAC_Inv_0.OUT.n45 21.1611
R38564 1Bit_DAC_Inv_0.OUT.n22 1Bit_DAC_Inv_0.OUT.n21 21.1611
R38565 1Bit_DAC_Inv_0.OUT.n28 1Bit_DAC_Inv_0.OUT.t40 6.5015
R38566 1Bit_DAC_Inv_0.OUT.n28 1Bit_DAC_Inv_0.OUT.t46 6.5015
R38567 1Bit_DAC_Inv_0.OUT.n30 1Bit_DAC_Inv_0.OUT.t43 6.5015
R38568 1Bit_DAC_Inv_0.OUT.n30 1Bit_DAC_Inv_0.OUT.t45 6.5015
R38569 1Bit_DAC_Inv_0.OUT.n36 1Bit_DAC_Inv_0.OUT.t1 6.5015
R38570 1Bit_DAC_Inv_0.OUT.n36 1Bit_DAC_Inv_0.OUT.t7 6.5015
R38571 1Bit_DAC_Inv_0.OUT.n32 1Bit_DAC_Inv_0.OUT.t49 6.5015
R38572 1Bit_DAC_Inv_0.OUT.n32 1Bit_DAC_Inv_0.OUT.t8 6.5015
R38573 1Bit_DAC_Inv_0.OUT.n34 1Bit_DAC_Inv_0.OUT.t6 6.5015
R38574 1Bit_DAC_Inv_0.OUT.n34 1Bit_DAC_Inv_0.OUT.t56 6.5015
R38575 1Bit_DAC_Inv_0.OUT.n39 1Bit_DAC_Inv_0.OUT.t9 6.5015
R38576 1Bit_DAC_Inv_0.OUT.n39 1Bit_DAC_Inv_0.OUT.t10 6.5015
R38577 1Bit_DAC_Inv_0.OUT.n43 1Bit_DAC_Inv_0.OUT.t47 6.5015
R38578 1Bit_DAC_Inv_0.OUT.n43 1Bit_DAC_Inv_0.OUT.t39 6.5015
R38579 1Bit_DAC_Inv_0.OUT.n47 1Bit_DAC_Inv_0.OUT.t52 6.5015
R38580 1Bit_DAC_Inv_0.OUT.n47 1Bit_DAC_Inv_0.OUT.t4 6.5015
R38581 1Bit_DAC_Inv_0.OUT.n51 1Bit_DAC_Inv_0.OUT.t48 6.5015
R38582 1Bit_DAC_Inv_0.OUT.n51 1Bit_DAC_Inv_0.OUT.t44 6.5015
R38583 1Bit_DAC_Inv_0.OUT.n16 1Bit_DAC_Inv_0.OUT.t21 6.5015
R38584 1Bit_DAC_Inv_0.OUT.n16 1Bit_DAC_Inv_0.OUT.t34 6.5015
R38585 1Bit_DAC_Inv_0.OUT.n14 1Bit_DAC_Inv_0.OUT.t25 6.5015
R38586 1Bit_DAC_Inv_0.OUT.n14 1Bit_DAC_Inv_0.OUT.t23 6.5015
R38587 1Bit_DAC_Inv_0.OUT.n12 1Bit_DAC_Inv_0.OUT.t26 6.5015
R38588 1Bit_DAC_Inv_0.OUT.n12 1Bit_DAC_Inv_0.OUT.t24 6.5015
R38589 1Bit_DAC_Inv_0.OUT.n6 1Bit_DAC_Inv_0.OUT.t27 6.5015
R38590 1Bit_DAC_Inv_0.OUT.n6 1Bit_DAC_Inv_0.OUT.t22 6.5015
R38591 1Bit_DAC_Inv_0.OUT.n4 1Bit_DAC_Inv_0.OUT.t29 6.5015
R38592 1Bit_DAC_Inv_0.OUT.n4 1Bit_DAC_Inv_0.OUT.t28 6.5015
R38593 1Bit_DAC_Inv_0.OUT.n10 1Bit_DAC_Inv_0.OUT.t32 6.5015
R38594 1Bit_DAC_Inv_0.OUT.n10 1Bit_DAC_Inv_0.OUT.t31 6.5015
R38595 1Bit_DAC_Inv_0.OUT.n8 1Bit_DAC_Inv_0.OUT.t20 6.5015
R38596 1Bit_DAC_Inv_0.OUT.n8 1Bit_DAC_Inv_0.OUT.t33 6.5015
R38597 1Bit_DAC_Inv_0.OUT.n2 1Bit_DAC_Inv_0.OUT.t30 6.5015
R38598 1Bit_DAC_Inv_0.OUT.n2 1Bit_DAC_Inv_0.OUT.t35 6.5015
R38599 1Bit_DAC_Inv_0.OUT.n0 1Bit_DAC_Inv_0.OUT.t37 6.5015
R38600 1Bit_DAC_Inv_0.OUT.n0 1Bit_DAC_Inv_0.OUT.t36 6.5015
R38601 1Bit_DAC_Inv_0.OUT.n41 1Bit_DAC_Inv_0.OUT.t12 3.9605
R38602 1Bit_DAC_Inv_0.OUT.n41 1Bit_DAC_Inv_0.OUT.t11 3.9605
R38603 1Bit_DAC_Inv_0.OUT.n45 1Bit_DAC_Inv_0.OUT.t15 3.9605
R38604 1Bit_DAC_Inv_0.OUT.n45 1Bit_DAC_Inv_0.OUT.t18 3.9605
R38605 1Bit_DAC_Inv_0.OUT.n49 1Bit_DAC_Inv_0.OUT.t19 3.9605
R38606 1Bit_DAC_Inv_0.OUT.n49 1Bit_DAC_Inv_0.OUT.t13 3.9605
R38607 1Bit_DAC_Inv_0.OUT.n53 1Bit_DAC_Inv_0.OUT.t16 3.9605
R38608 1Bit_DAC_Inv_0.OUT.n53 1Bit_DAC_Inv_0.OUT.t14 3.9605
R38609 1Bit_DAC_Inv_0.OUT.n23 1Bit_DAC_Inv_0.OUT.t42 3.9605
R38610 1Bit_DAC_Inv_0.OUT.n23 1Bit_DAC_Inv_0.OUT.t5 3.9605
R38611 1Bit_DAC_Inv_0.OUT.n21 1Bit_DAC_Inv_0.OUT.t53 3.9605
R38612 1Bit_DAC_Inv_0.OUT.n21 1Bit_DAC_Inv_0.OUT.t3 3.9605
R38613 1Bit_DAC_Inv_0.OUT.n19 1Bit_DAC_Inv_0.OUT.t55 3.9605
R38614 1Bit_DAC_Inv_0.OUT.n19 1Bit_DAC_Inv_0.OUT.t2 3.9605
R38615 1Bit_DAC_Inv_0.OUT.n18 1Bit_DAC_Inv_0.OUT.t51 3.9605
R38616 1Bit_DAC_Inv_0.OUT.n18 1Bit_DAC_Inv_0.OUT.t54 3.9605
R38617 1Bit_DAC_Inv_0.OUT.n29 1Bit_DAC_Inv_0.OUT.t41 3.85167
R38618 1Bit_DAC_Inv_0.OUT.n27 1Bit_DAC_Inv_0.OUT.n17 0.3013
R38619 1Bit_DAC_Inv_0.OUT.n27 1Bit_DAC_Inv_0.OUT.n26 0.2355
R38620 1Bit_DAC_Inv_0.OUT.n26 1Bit_DAC_Inv_0.OUT 0.1415
R38621 1Bit_DAC_Inv_0.OUT.n3 1Bit_DAC_Inv_0.OUT.n1 0.0631667
R38622 1Bit_DAC_Inv_0.OUT.n7 1Bit_DAC_Inv_0.OUT.n5 0.0631667
R38623 1Bit_DAC_Inv_0.OUT.n9 1Bit_DAC_Inv_0.OUT.n7 0.0631667
R38624 1Bit_DAC_Inv_0.OUT.n11 1Bit_DAC_Inv_0.OUT.n9 0.0631667
R38625 1Bit_DAC_Inv_0.OUT.n13 1Bit_DAC_Inv_0.OUT.n11 0.0631667
R38626 1Bit_DAC_Inv_0.OUT.n15 1Bit_DAC_Inv_0.OUT.n13 0.0631667
R38627 1Bit_DAC_Inv_0.OUT.n24 1Bit_DAC_Inv_0.OUT.n22 0.0631667
R38628 1Bit_DAC_Inv_0.OUT.n22 1Bit_DAC_Inv_0.OUT.n20 0.0569
R38629 1Bit_DAC_Inv_0.OUT.n25 1Bit_DAC_Inv_0.OUT.n24 0.0569
R38630 1Bit_DAC_Inv_0.OUT.n5 1Bit_DAC_Inv_0.OUT.n3 0.0506333
R38631 1Bit_DAC_Inv_0.OUT.n17 1Bit_DAC_Inv_0.OUT.n15 0.0443667
R38632 1Bit_DAC_Inv_0.OUT.n26 1Bit_DAC_Inv_0.OUT.n25 0.0349667
R38633 1Bit_DAC_Inv_0.OUT.n37 1Bit_DAC_Inv_0.OUT.n35 0.024
R38634 1Bit_DAC_Inv_0.OUT.n35 1Bit_DAC_Inv_0.OUT.n33 0.024
R38635 1Bit_DAC_Inv_0.OUT.n33 1Bit_DAC_Inv_0.OUT.n31 0.024
R38636 1Bit_DAC_Inv_0.OUT.n31 1Bit_DAC_Inv_0.OUT.n29 0.01695
R38637 1Bit_DAC_Inv_0.OUT.n44 1Bit_DAC_Inv_0.OUT.n42 0.0125
R38638 1Bit_DAC_Inv_0.OUT.n40 1Bit_DAC_Inv_0.OUT.n38 0.0125
R38639 1Bit_DAC_Inv_0.OUT 1Bit_DAC_Inv_0.OUT.n55 0.0115
R38640 1Bit_DAC_Inv_0.OUT.n55 1Bit_DAC_Inv_0.OUT.n54 0.0105
R38641 1Bit_DAC_Inv_0.OUT.n54 1Bit_DAC_Inv_0.OUT.n52 0.0105
R38642 1Bit_DAC_Inv_0.OUT.n52 1Bit_DAC_Inv_0.OUT.n50 0.0105
R38643 1Bit_DAC_Inv_0.OUT.n50 1Bit_DAC_Inv_0.OUT.n48 0.0105
R38644 1Bit_DAC_Inv_0.OUT.n48 1Bit_DAC_Inv_0.OUT.n46 0.0105
R38645 1Bit_DAC_Inv_0.OUT 1Bit_DAC_Inv_0.OUT.n27 0.01
R38646 1Bit_DAC_Inv_0.OUT.n38 1Bit_DAC_Inv_0.OUT.n37 0.009025
R38647 1Bit_DAC_Inv_0.OUT.n42 1Bit_DAC_Inv_0.OUT.n40 0.0085
R38648 1Bit_DAC_Inv_0.OUT.n46 1Bit_DAC_Inv_0.OUT.n44 0.0065
R38649 a_181475_n46496.n9 a_181475_n46496.t9 1038.79
R38650 a_181475_n46496.n1 a_181475_n46496.t12 1038.78
R38651 a_181475_n46496.n9 a_181475_n46496.t14 1038.55
R38652 a_181475_n46496.n10 a_181475_n46496.t15 1038.55
R38653 a_181475_n46496.n11 a_181475_n46496.t28 1038.55
R38654 a_181475_n46496.n12 a_181475_n46496.t8 1038.55
R38655 a_181475_n46496.n13 a_181475_n46496.t22 1038.55
R38656 a_181475_n46496.n14 a_181475_n46496.t26 1038.55
R38657 a_181475_n46496.n15 a_181475_n46496.t27 1038.55
R38658 a_181475_n46496.n16 a_181475_n46496.t7 1038.55
R38659 a_181475_n46496.n17 a_181475_n46496.t21 1038.55
R38660 a_181475_n46496.n8 a_181475_n46496.t10 1038.54
R38661 a_181475_n46496.n7 a_181475_n46496.t6 1038.54
R38662 a_181475_n46496.n6 a_181475_n46496.t24 1038.54
R38663 a_181475_n46496.n5 a_181475_n46496.t23 1038.54
R38664 a_181475_n46496.n4 a_181475_n46496.t11 1038.54
R38665 a_181475_n46496.n3 a_181475_n46496.t29 1038.54
R38666 a_181475_n46496.n2 a_181475_n46496.t25 1038.54
R38667 a_181475_n46496.n1 a_181475_n46496.t13 1038.54
R38668 a_181475_n46496.n19 a_181475_n46496.t31 1024.08
R38669 a_181475_n46496.n20 a_181475_n46496.t33 1024.08
R38670 a_181475_n46496.n21 a_181475_n46496.t18 1024.08
R38671 a_181475_n46496.n22 a_181475_n46496.t19 1024.08
R38672 a_181475_n46496.n23 a_181475_n46496.t30 1024.08
R38673 a_181475_n46496.n24 a_181475_n46496.t20 1024.08
R38674 a_181475_n46496.n25 a_181475_n46496.t17 1024.08
R38675 a_181475_n46496.n26 a_181475_n46496.t16 1024.08
R38676 a_181475_n46496.n27 a_181475_n46496.t32 1024.08
R38677 a_181475_n46496.n31 a_181475_n46496.n30 52.1388
R38678 a_181475_n46496.n33 a_181475_n46496.n32 48.672
R38679 a_181475_n46496.n32 a_181475_n46496.n0 19.8859
R38680 a_181475_n46496.n24 a_181475_n46496.n23 11.077
R38681 a_181475_n46496.n29 a_181475_n46496.n18 9.73487
R38682 a_181475_n46496.n28 a_181475_n46496.n19 7.41906
R38683 a_181475_n46496.n30 a_181475_n46496.t3 6.5015
R38684 a_181475_n46496.n30 a_181475_n46496.t2 6.5015
R38685 a_181475_n46496.t5 a_181475_n46496.n33 6.5015
R38686 a_181475_n46496.n33 a_181475_n46496.t4 6.5015
R38687 a_181475_n46496.n28 a_181475_n46496.n27 6.17675
R38688 a_181475_n46496.n18 a_181475_n46496.n8 5.65425
R38689 a_181475_n46496.n18 a_181475_n46496.n17 5.40925
R38690 a_181475_n46496.n0 a_181475_n46496.t1 3.9605
R38691 a_181475_n46496.n0 a_181475_n46496.t0 3.9605
R38692 a_181475_n46496.n31 a_181475_n46496.n29 3.62884
R38693 a_181475_n46496.n32 a_181475_n46496.n31 3.48527
R38694 a_181475_n46496.n23 a_181475_n46496.n22 0.428449
R38695 a_181475_n46496.n22 a_181475_n46496.n21 0.428449
R38696 a_181475_n46496.n21 a_181475_n46496.n20 0.428449
R38697 a_181475_n46496.n20 a_181475_n46496.n19 0.428449
R38698 a_181475_n46496.n27 a_181475_n46496.n26 0.2405
R38699 a_181475_n46496.n26 a_181475_n46496.n25 0.2405
R38700 a_181475_n46496.n25 a_181475_n46496.n24 0.2405
R38701 a_181475_n46496.n2 a_181475_n46496.n1 0.2405
R38702 a_181475_n46496.n3 a_181475_n46496.n2 0.2405
R38703 a_181475_n46496.n4 a_181475_n46496.n3 0.2405
R38704 a_181475_n46496.n5 a_181475_n46496.n4 0.2405
R38705 a_181475_n46496.n6 a_181475_n46496.n5 0.2405
R38706 a_181475_n46496.n7 a_181475_n46496.n6 0.2405
R38707 a_181475_n46496.n8 a_181475_n46496.n7 0.2405
R38708 a_181475_n46496.n10 a_181475_n46496.n9 0.2405
R38709 a_181475_n46496.n11 a_181475_n46496.n10 0.2405
R38710 a_181475_n46496.n12 a_181475_n46496.n11 0.2405
R38711 a_181475_n46496.n13 a_181475_n46496.n12 0.2405
R38712 a_181475_n46496.n14 a_181475_n46496.n13 0.2405
R38713 a_181475_n46496.n15 a_181475_n46496.n14 0.2405
R38714 a_181475_n46496.n16 a_181475_n46496.n15 0.2405
R38715 a_181475_n46496.n17 a_181475_n46496.n16 0.2405
R38716 a_181475_n46496.n29 a_181475_n46496.n28 0.1255
R38717 VREFN.n45 VREFN.t36 57.4419
R38718 VREFN.n17 VREFN.t17 57.4419
R38719 VREFN.n30 VREFN.n28 51.0245
R38720 VREFN.n2 VREFN.n0 51.0245
R38721 VREFN.n42 VREFN.n41 50.9409
R38722 VREFN.n36 VREFN.n35 50.9409
R38723 VREFN.n32 VREFN.n31 50.9409
R38724 VREFN.n14 VREFN.n13 50.9409
R38725 VREFN.n8 VREFN.n7 50.9409
R38726 VREFN.n4 VREFN.n3 50.9409
R38727 VREFN.n44 VREFN.n43 50.9305
R38728 VREFN.n40 VREFN.n39 50.9305
R38729 VREFN.n38 VREFN.n37 50.9305
R38730 VREFN.n34 VREFN.n33 50.9305
R38731 VREFN.n30 VREFN.n29 50.9305
R38732 VREFN.n16 VREFN.n15 50.9305
R38733 VREFN.n12 VREFN.n11 50.9305
R38734 VREFN.n10 VREFN.n9 50.9305
R38735 VREFN.n6 VREFN.n5 50.9305
R38736 VREFN.n2 VREFN.n1 50.9305
R38737 VREFN.n48 VREFN.t4 26.3525
R38738 VREFN.n20 VREFN.t51 26.3525
R38739 VREFN.n54 VREFN.n53 22.3124
R38740 VREFN.n50 VREFN.n49 22.3124
R38741 VREFN.n26 VREFN.n25 22.3124
R38742 VREFN.n22 VREFN.n21 22.3124
R38743 VREFN.n52 VREFN.n51 22.302
R38744 VREFN.n48 VREFN.n47 22.302
R38745 VREFN.n24 VREFN.n23 22.302
R38746 VREFN.n20 VREFN.n19 22.302
R38747 VREFN.n43 VREFN.t45 6.5015
R38748 VREFN.n43 VREFN.t42 6.5015
R38749 VREFN.n41 VREFN.t30 6.5015
R38750 VREFN.n41 VREFN.t46 6.5015
R38751 VREFN.n39 VREFN.t31 6.5015
R38752 VREFN.n39 VREFN.t33 6.5015
R38753 VREFN.n37 VREFN.t35 6.5015
R38754 VREFN.n37 VREFN.t34 6.5015
R38755 VREFN.n35 VREFN.t44 6.5015
R38756 VREFN.n35 VREFN.t41 6.5015
R38757 VREFN.n33 VREFN.t29 6.5015
R38758 VREFN.n33 VREFN.t28 6.5015
R38759 VREFN.n31 VREFN.t37 6.5015
R38760 VREFN.n31 VREFN.t32 6.5015
R38761 VREFN.n29 VREFN.t38 6.5015
R38762 VREFN.n29 VREFN.t39 6.5015
R38763 VREFN.n28 VREFN.t43 6.5015
R38764 VREFN.n28 VREFN.t40 6.5015
R38765 VREFN.n15 VREFN.t26 6.5015
R38766 VREFN.n15 VREFN.t23 6.5015
R38767 VREFN.n13 VREFN.t11 6.5015
R38768 VREFN.n13 VREFN.t27 6.5015
R38769 VREFN.n11 VREFN.t12 6.5015
R38770 VREFN.n11 VREFN.t14 6.5015
R38771 VREFN.n9 VREFN.t16 6.5015
R38772 VREFN.n9 VREFN.t15 6.5015
R38773 VREFN.n7 VREFN.t25 6.5015
R38774 VREFN.n7 VREFN.t22 6.5015
R38775 VREFN.n5 VREFN.t10 6.5015
R38776 VREFN.n5 VREFN.t9 6.5015
R38777 VREFN.n3 VREFN.t18 6.5015
R38778 VREFN.n3 VREFN.t13 6.5015
R38779 VREFN.n1 VREFN.t19 6.5015
R38780 VREFN.n1 VREFN.t20 6.5015
R38781 VREFN.n0 VREFN.t24 6.5015
R38782 VREFN.n0 VREFN.t21 6.5015
R38783 VREFN.n46 VREFN.n45 5.839
R38784 VREFN.n18 VREFN.n17 5.839
R38785 VREFN.n55 VREFN.n54 4.04735
R38786 VREFN.n27 VREFN.n26 4.04735
R38787 VREFN.n53 VREFN.t6 3.9605
R38788 VREFN.n53 VREFN.t5 3.9605
R38789 VREFN.n51 VREFN.t8 3.9605
R38790 VREFN.n51 VREFN.t7 3.9605
R38791 VREFN.n49 VREFN.t2 3.9605
R38792 VREFN.n49 VREFN.t0 3.9605
R38793 VREFN.n47 VREFN.t3 3.9605
R38794 VREFN.n47 VREFN.t1 3.9605
R38795 VREFN.n25 VREFN.t53 3.9605
R38796 VREFN.n25 VREFN.t52 3.9605
R38797 VREFN.n23 VREFN.t55 3.9605
R38798 VREFN.n23 VREFN.t54 3.9605
R38799 VREFN.n21 VREFN.t49 3.9605
R38800 VREFN.n21 VREFN.t47 3.9605
R38801 VREFN.n19 VREFN.t50 3.9605
R38802 VREFN.n19 VREFN.t48 3.9605
R38803 VREFN VREFN.n27 2.78503
R38804 VREFN.n56 VREFN.n55 2.51497
R38805 VREFN VREFN.n56 0.346688
R38806 VREFN.n50 VREFN.n48 0.0945
R38807 VREFN.n54 VREFN.n52 0.0945
R38808 VREFN.n32 VREFN.n30 0.0945
R38809 VREFN.n36 VREFN.n34 0.0945
R38810 VREFN.n40 VREFN.n38 0.0945
R38811 VREFN.n42 VREFN.n40 0.0945
R38812 VREFN.n45 VREFN.n44 0.0945
R38813 VREFN.n22 VREFN.n20 0.0945
R38814 VREFN.n26 VREFN.n24 0.0945
R38815 VREFN.n4 VREFN.n2 0.0945
R38816 VREFN.n8 VREFN.n6 0.0945
R38817 VREFN.n12 VREFN.n10 0.0945
R38818 VREFN.n14 VREFN.n12 0.0945
R38819 VREFN.n17 VREFN.n16 0.0945
R38820 VREFN.n52 VREFN.n50 0.0851
R38821 VREFN.n34 VREFN.n32 0.0851
R38822 VREFN.n38 VREFN.n36 0.0851
R38823 VREFN.n44 VREFN.n42 0.0851
R38824 VREFN.n24 VREFN.n22 0.0851
R38825 VREFN.n6 VREFN.n4 0.0851
R38826 VREFN.n10 VREFN.n8 0.0851
R38827 VREFN.n16 VREFN.n14 0.0851
R38828 VREFN.n56 VREFN 0.0295
R38829 VREFN.n46 VREFN 0.0255
R38830 VREFN.n18 VREFN 0.0255
R38831 VREFN.n55 VREFN 0.016125
R38832 VREFN.n27 VREFN 0.016125
R38833 VREFN VREFN.n46 0.00675
R38834 VREFN VREFN.n18 0.00675
R38835 a_185229_n11365.n178 a_185229_n11365.n177 815.966
R38836 a_185229_n11365.n317 a_185229_n11365.n311 585
R38837 a_185229_n11365.n317 a_185229_n11365.n310 585
R38838 a_185229_n11365.n318 a_185229_n11365.n317 585
R38839 a_185229_n11365.n303 a_185229_n11365.n297 585
R38840 a_185229_n11365.n303 a_185229_n11365.n296 585
R38841 a_185229_n11365.n304 a_185229_n11365.n303 585
R38842 a_185229_n11365.n289 a_185229_n11365.n283 585
R38843 a_185229_n11365.n289 a_185229_n11365.n282 585
R38844 a_185229_n11365.n290 a_185229_n11365.n289 585
R38845 a_185229_n11365.n275 a_185229_n11365.n269 585
R38846 a_185229_n11365.n275 a_185229_n11365.n268 585
R38847 a_185229_n11365.n276 a_185229_n11365.n275 585
R38848 a_185229_n11365.n261 a_185229_n11365.n255 585
R38849 a_185229_n11365.n261 a_185229_n11365.n254 585
R38850 a_185229_n11365.n262 a_185229_n11365.n261 585
R38851 a_185229_n11365.n247 a_185229_n11365.n241 585
R38852 a_185229_n11365.n247 a_185229_n11365.n240 585
R38853 a_185229_n11365.n248 a_185229_n11365.n247 585
R38854 a_185229_n11365.n233 a_185229_n11365.n227 585
R38855 a_185229_n11365.n233 a_185229_n11365.n226 585
R38856 a_185229_n11365.n234 a_185229_n11365.n233 585
R38857 a_185229_n11365.n219 a_185229_n11365.n213 585
R38858 a_185229_n11365.n219 a_185229_n11365.n212 585
R38859 a_185229_n11365.n220 a_185229_n11365.n219 585
R38860 a_185229_n11365.n205 a_185229_n11365.n199 585
R38861 a_185229_n11365.n205 a_185229_n11365.n198 585
R38862 a_185229_n11365.n206 a_185229_n11365.n205 585
R38863 a_185229_n11365.n191 a_185229_n11365.n185 585
R38864 a_185229_n11365.n191 a_185229_n11365.n184 585
R38865 a_185229_n11365.n192 a_185229_n11365.n191 585
R38866 a_185229_n11365.n162 a_185229_n11365.n161 585
R38867 a_185229_n11365.n159 a_185229_n11365.n158 585
R38868 a_185229_n11365.n169 a_185229_n11365.n168 585
R38869 a_185229_n11365.n171 a_185229_n11365.n170 585
R38870 a_185229_n11365.n156 a_185229_n11365.n155 585
R38871 a_185229_n11365.n177 a_185229_n11365.n176 585
R38872 a_185229_n11365.n102 a_185229_n11365.t43 433.149
R38873 a_185229_n11365.t43 a_185229_n11365.n86 433.149
R38874 a_185229_n11365.n101 a_185229_n11365.t55 433.149
R38875 a_185229_n11365.t55 a_185229_n11365.n100 433.149
R38876 a_185229_n11365.t51 a_185229_n11365.n88 433.149
R38877 a_185229_n11365.n99 a_185229_n11365.t51 433.149
R38878 a_185229_n11365.t70 a_185229_n11365.n97 433.149
R38879 a_185229_n11365.n98 a_185229_n11365.t70 433.149
R38880 a_185229_n11365.n96 a_185229_n11365.t66 433.149
R38881 a_185229_n11365.t66 a_185229_n11365.n89 433.149
R38882 a_185229_n11365.n95 a_185229_n11365.t59 433.149
R38883 a_185229_n11365.t59 a_185229_n11365.n94 433.149
R38884 a_185229_n11365.t56 a_185229_n11365.n90 433.149
R38885 a_185229_n11365.n93 a_185229_n11365.t56 433.149
R38886 a_185229_n11365.t53 a_185229_n11365.n148 433.149
R38887 a_185229_n11365.n149 a_185229_n11365.t53 433.149
R38888 a_185229_n11365.t50 a_185229_n11365.n4 433.149
R38889 a_185229_n11365.n5 a_185229_n11365.t50 433.149
R38890 a_185229_n11365.t60 a_185229_n11365.n113 433.149
R38891 a_185229_n11365.n114 a_185229_n11365.t60 433.149
R38892 a_185229_n11365.n116 a_185229_n11365.t52 433.149
R38893 a_185229_n11365.t52 a_185229_n11365.n115 433.149
R38894 a_185229_n11365.n117 a_185229_n11365.t33 433.149
R38895 a_185229_n11365.t33 a_185229_n11365.n112 433.149
R38896 a_185229_n11365.t69 a_185229_n11365.n118 433.149
R38897 a_185229_n11365.n119 a_185229_n11365.t69 433.149
R38898 a_185229_n11365.t63 a_185229_n11365.n111 433.149
R38899 a_185229_n11365.n120 a_185229_n11365.t63 433.149
R38900 a_185229_n11365.n122 a_185229_n11365.t58 433.149
R38901 a_185229_n11365.t58 a_185229_n11365.n121 433.149
R38902 a_185229_n11365.n123 a_185229_n11365.t65 433.149
R38903 a_185229_n11365.t65 a_185229_n11365.n110 433.149
R38904 a_185229_n11365.t48 a_185229_n11365.n124 433.149
R38905 a_185229_n11365.n125 a_185229_n11365.t48 433.149
R38906 a_185229_n11365.t41 a_185229_n11365.n109 433.149
R38907 a_185229_n11365.n126 a_185229_n11365.t41 433.149
R38908 a_185229_n11365.n128 a_185229_n11365.t35 433.149
R38909 a_185229_n11365.t35 a_185229_n11365.n127 433.149
R38910 a_185229_n11365.n129 a_185229_n11365.t71 433.149
R38911 a_185229_n11365.t71 a_185229_n11365.n108 433.149
R38912 a_185229_n11365.t67 a_185229_n11365.n130 433.149
R38913 a_185229_n11365.n131 a_185229_n11365.t67 433.149
R38914 a_185229_n11365.t44 a_185229_n11365.n107 433.149
R38915 a_185229_n11365.n132 a_185229_n11365.t44 433.149
R38916 a_185229_n11365.n134 a_185229_n11365.t36 433.149
R38917 a_185229_n11365.t36 a_185229_n11365.n133 433.149
R38918 a_185229_n11365.n135 a_185229_n11365.t32 433.149
R38919 a_185229_n11365.t32 a_185229_n11365.n106 433.149
R38920 a_185229_n11365.t68 a_185229_n11365.n136 433.149
R38921 a_185229_n11365.n137 a_185229_n11365.t68 433.149
R38922 a_185229_n11365.t62 a_185229_n11365.n105 433.149
R38923 a_185229_n11365.n138 a_185229_n11365.t62 433.149
R38924 a_185229_n11365.n140 a_185229_n11365.t42 433.149
R38925 a_185229_n11365.t42 a_185229_n11365.n139 433.149
R38926 a_185229_n11365.n141 a_185229_n11365.t38 433.149
R38927 a_185229_n11365.t38 a_185229_n11365.n104 433.149
R38928 a_185229_n11365.t47 a_185229_n11365.n142 433.149
R38929 a_185229_n11365.n143 a_185229_n11365.t47 433.149
R38930 a_185229_n11365.t40 a_185229_n11365.n103 433.149
R38931 a_185229_n11365.n144 a_185229_n11365.t40 433.149
R38932 a_185229_n11365.n146 a_185229_n11365.t34 433.149
R38933 a_185229_n11365.t34 a_185229_n11365.n145 433.149
R38934 a_185229_n11365.n147 a_185229_n11365.t57 433.149
R38935 a_185229_n11365.t57 a_185229_n11365.n87 433.149
R38936 a_185229_n11365.n324 a_185229_n11365.t54 433.149
R38937 a_185229_n11365.t54 a_185229_n11365.n323 433.149
R38938 a_185229_n11365.t64 a_185229_n11365.n0 433.149
R38939 a_185229_n11365.n334 a_185229_n11365.t64 433.149
R38940 a_185229_n11365.t46 a_185229_n11365.n332 433.149
R38941 a_185229_n11365.n333 a_185229_n11365.t46 433.149
R38942 a_185229_n11365.n331 a_185229_n11365.t39 433.149
R38943 a_185229_n11365.t39 a_185229_n11365.n1 433.149
R38944 a_185229_n11365.n330 a_185229_n11365.t49 433.149
R38945 a_185229_n11365.t49 a_185229_n11365.n329 433.149
R38946 a_185229_n11365.t45 a_185229_n11365.n2 433.149
R38947 a_185229_n11365.n328 a_185229_n11365.t45 433.149
R38948 a_185229_n11365.t37 a_185229_n11365.n326 433.149
R38949 a_185229_n11365.n327 a_185229_n11365.t37 433.149
R38950 a_185229_n11365.n325 a_185229_n11365.t61 433.149
R38951 a_185229_n11365.t61 a_185229_n11365.n3 433.149
R38952 a_185229_n11365.t9 a_185229_n11365.n160 384.339
R38953 a_185229_n11365.n16 a_185229_n11365.n15 325.69
R38954 a_185229_n11365.n161 a_185229_n11365.n158 230.966
R38955 a_185229_n11365.n169 a_185229_n11365.n158 230.966
R38956 a_185229_n11365.n170 a_185229_n11365.n169 230.966
R38957 a_185229_n11365.n170 a_185229_n11365.n155 230.966
R38958 a_185229_n11365.n177 a_185229_n11365.n155 230.966
R38959 a_185229_n11365.n17 a_185229_n11365.n16 185
R38960 a_185229_n11365.n12 a_185229_n11365.n11 185
R38961 a_185229_n11365.n24 a_185229_n11365.n23 185
R38962 a_185229_n11365.n25 a_185229_n11365.n9 185
R38963 a_185229_n11365.n30 a_185229_n11365.n29 185
R38964 a_185229_n11365.n28 a_185229_n11365.n27 185
R38965 a_185229_n11365.n42 a_185229_n11365.n39 185
R38966 a_185229_n11365.n44 a_185229_n11365.n39 185
R38967 a_185229_n11365.n40 a_185229_n11365.n39 185
R38968 a_185229_n11365.n49 a_185229_n11365.n39 185
R38969 a_185229_n11365.n58 a_185229_n11365.n55 185
R38970 a_185229_n11365.n60 a_185229_n11365.n55 185
R38971 a_185229_n11365.n56 a_185229_n11365.n55 185
R38972 a_185229_n11365.n65 a_185229_n11365.n55 185
R38973 a_185229_n11365.n74 a_185229_n11365.n71 185
R38974 a_185229_n11365.n76 a_185229_n11365.n71 185
R38975 a_185229_n11365.n72 a_185229_n11365.n71 185
R38976 a_185229_n11365.n81 a_185229_n11365.n71 185
R38977 a_185229_n11365.n26 a_185229_n11365.t1 174.857
R38978 a_185229_n11365.n16 a_185229_n11365.n11 140.69
R38979 a_185229_n11365.n24 a_185229_n11365.n11 140.69
R38980 a_185229_n11365.n25 a_185229_n11365.n24 140.69
R38981 a_185229_n11365.n29 a_185229_n11365.n25 140.69
R38982 a_185229_n11365.n29 a_185229_n11365.n28 140.69
R38983 a_185229_n11365.n161 a_185229_n11365.t9 115.484
R38984 a_185229_n11365.n28 a_185229_n11365.t1 70.3453
R38985 a_185229_n11365.n317 a_185229_n11365.n316 51.6891
R38986 a_185229_n11365.n303 a_185229_n11365.n302 51.6891
R38987 a_185229_n11365.n289 a_185229_n11365.n288 51.6891
R38988 a_185229_n11365.n275 a_185229_n11365.n274 51.6891
R38989 a_185229_n11365.n261 a_185229_n11365.n260 51.6891
R38990 a_185229_n11365.n247 a_185229_n11365.n246 51.6891
R38991 a_185229_n11365.n233 a_185229_n11365.n232 51.6891
R38992 a_185229_n11365.n219 a_185229_n11365.n218 51.6891
R38993 a_185229_n11365.n205 a_185229_n11365.n204 51.6891
R38994 a_185229_n11365.n191 a_185229_n11365.n190 51.6891
R38995 a_185229_n11365.n316 a_185229_n11365.n315 29.8062
R38996 a_185229_n11365.n302 a_185229_n11365.n301 29.8062
R38997 a_185229_n11365.n288 a_185229_n11365.n287 29.8062
R38998 a_185229_n11365.n274 a_185229_n11365.n273 29.8062
R38999 a_185229_n11365.n260 a_185229_n11365.n259 29.8062
R39000 a_185229_n11365.n246 a_185229_n11365.n245 29.8062
R39001 a_185229_n11365.n232 a_185229_n11365.n231 29.8062
R39002 a_185229_n11365.n218 a_185229_n11365.n217 29.8062
R39003 a_185229_n11365.n204 a_185229_n11365.n203 29.8062
R39004 a_185229_n11365.n190 a_185229_n11365.n189 29.8062
R39005 a_185229_n11365.n162 a_185229_n11365.n160 29.3167
R39006 a_185229_n11365.n27 a_185229_n11365.n26 28.4333
R39007 a_185229_n11365.n51 a_185229_n11365.n50 26.8428
R39008 a_185229_n11365.n67 a_185229_n11365.n66 26.8428
R39009 a_185229_n11365.n83 a_185229_n11365.n82 26.8428
R39010 a_185229_n11365.n163 a_185229_n11365.n159 24.8476
R39011 a_185229_n11365.n30 a_185229_n11365.n10 24.8476
R39012 a_185229_n11365.n168 a_185229_n11365.n167 23.3417
R39013 a_185229_n11365.n31 a_185229_n11365.n9 23.3417
R39014 a_185229_n11365.n171 a_185229_n11365.n157 21.8358
R39015 a_185229_n11365.n23 a_185229_n11365.n22 21.8358
R39016 a_185229_n11365.n50 a_185229_n11365.n49 21.8358
R39017 a_185229_n11365.n66 a_185229_n11365.n65 21.8358
R39018 a_185229_n11365.n82 a_185229_n11365.n81 21.8358
R39019 a_185229_n11365.n315 a_185229_n11365.n311 20.3299
R39020 a_185229_n11365.n301 a_185229_n11365.n297 20.3299
R39021 a_185229_n11365.n287 a_185229_n11365.n283 20.3299
R39022 a_185229_n11365.n273 a_185229_n11365.n269 20.3299
R39023 a_185229_n11365.n259 a_185229_n11365.n255 20.3299
R39024 a_185229_n11365.n245 a_185229_n11365.n241 20.3299
R39025 a_185229_n11365.n231 a_185229_n11365.n227 20.3299
R39026 a_185229_n11365.n217 a_185229_n11365.n213 20.3299
R39027 a_185229_n11365.n203 a_185229_n11365.n199 20.3299
R39028 a_185229_n11365.n189 a_185229_n11365.n185 20.3299
R39029 a_185229_n11365.n172 a_185229_n11365.n156 20.3299
R39030 a_185229_n11365.n21 a_185229_n11365.n12 20.3299
R39031 a_185229_n11365.n48 a_185229_n11365.n40 20.3299
R39032 a_185229_n11365.n64 a_185229_n11365.n56 20.3299
R39033 a_185229_n11365.n80 a_185229_n11365.n72 20.3299
R39034 a_185229_n11365.n319 a_185229_n11365.n318 19.1618
R39035 a_185229_n11365.n305 a_185229_n11365.n304 19.1618
R39036 a_185229_n11365.n291 a_185229_n11365.n290 19.1618
R39037 a_185229_n11365.n277 a_185229_n11365.n276 19.1618
R39038 a_185229_n11365.n263 a_185229_n11365.n262 19.1618
R39039 a_185229_n11365.n249 a_185229_n11365.n248 19.1618
R39040 a_185229_n11365.n235 a_185229_n11365.n234 19.1618
R39041 a_185229_n11365.n221 a_185229_n11365.n220 19.1618
R39042 a_185229_n11365.n207 a_185229_n11365.n206 19.1618
R39043 a_185229_n11365.n193 a_185229_n11365.n192 19.1618
R39044 a_185229_n11365.n179 a_185229_n11365.n178 19.1618
R39045 a_185229_n11365.n15 a_185229_n11365.n6 19.1618
R39046 a_185229_n11365.n42 a_185229_n11365.n37 19.1618
R39047 a_185229_n11365.n58 a_185229_n11365.n36 19.1618
R39048 a_185229_n11365.n74 a_185229_n11365.n35 19.1618
R39049 a_185229_n11365.n312 a_185229_n11365.n310 18.824
R39050 a_185229_n11365.n298 a_185229_n11365.n296 18.824
R39051 a_185229_n11365.n284 a_185229_n11365.n282 18.824
R39052 a_185229_n11365.n270 a_185229_n11365.n268 18.824
R39053 a_185229_n11365.n256 a_185229_n11365.n254 18.824
R39054 a_185229_n11365.n242 a_185229_n11365.n240 18.824
R39055 a_185229_n11365.n228 a_185229_n11365.n226 18.824
R39056 a_185229_n11365.n214 a_185229_n11365.n212 18.824
R39057 a_185229_n11365.n200 a_185229_n11365.n198 18.824
R39058 a_185229_n11365.n186 a_185229_n11365.n184 18.824
R39059 a_185229_n11365.n176 a_185229_n11365.n175 18.824
R39060 a_185229_n11365.n18 a_185229_n11365.n17 18.824
R39061 a_185229_n11365.n45 a_185229_n11365.n44 18.824
R39062 a_185229_n11365.n61 a_185229_n11365.n60 18.824
R39063 a_185229_n11365.n77 a_185229_n11365.n76 18.824
R39064 a_185229_n11365.n318 a_185229_n11365.n309 17.3181
R39065 a_185229_n11365.n304 a_185229_n11365.n295 17.3181
R39066 a_185229_n11365.n290 a_185229_n11365.n281 17.3181
R39067 a_185229_n11365.n276 a_185229_n11365.n267 17.3181
R39068 a_185229_n11365.n262 a_185229_n11365.n253 17.3181
R39069 a_185229_n11365.n248 a_185229_n11365.n239 17.3181
R39070 a_185229_n11365.n234 a_185229_n11365.n225 17.3181
R39071 a_185229_n11365.n220 a_185229_n11365.n211 17.3181
R39072 a_185229_n11365.n206 a_185229_n11365.n197 17.3181
R39073 a_185229_n11365.n192 a_185229_n11365.n183 17.3181
R39074 a_185229_n11365.n178 a_185229_n11365.n154 17.3181
R39075 a_185229_n11365.n15 a_185229_n11365.n14 17.3181
R39076 a_185229_n11365.n43 a_185229_n11365.n42 17.3181
R39077 a_185229_n11365.n59 a_185229_n11365.n58 17.3181
R39078 a_185229_n11365.n75 a_185229_n11365.n74 17.3181
R39079 a_185229_n11365.n51 a_185229_n11365.n39 16.7801
R39080 a_185229_n11365.n67 a_185229_n11365.n55 16.7801
R39081 a_185229_n11365.n83 a_185229_n11365.n71 16.7801
R39082 a_185229_n11365.n309 a_185229_n11365.n308 9.3005
R39083 a_185229_n11365.n315 a_185229_n11365.n314 9.3005
R39084 a_185229_n11365.n313 a_185229_n11365.n312 9.3005
R39085 a_185229_n11365.n295 a_185229_n11365.n294 9.3005
R39086 a_185229_n11365.n301 a_185229_n11365.n300 9.3005
R39087 a_185229_n11365.n299 a_185229_n11365.n298 9.3005
R39088 a_185229_n11365.n281 a_185229_n11365.n280 9.3005
R39089 a_185229_n11365.n287 a_185229_n11365.n286 9.3005
R39090 a_185229_n11365.n285 a_185229_n11365.n284 9.3005
R39091 a_185229_n11365.n267 a_185229_n11365.n266 9.3005
R39092 a_185229_n11365.n273 a_185229_n11365.n272 9.3005
R39093 a_185229_n11365.n271 a_185229_n11365.n270 9.3005
R39094 a_185229_n11365.n253 a_185229_n11365.n252 9.3005
R39095 a_185229_n11365.n259 a_185229_n11365.n258 9.3005
R39096 a_185229_n11365.n257 a_185229_n11365.n256 9.3005
R39097 a_185229_n11365.n239 a_185229_n11365.n238 9.3005
R39098 a_185229_n11365.n245 a_185229_n11365.n244 9.3005
R39099 a_185229_n11365.n243 a_185229_n11365.n242 9.3005
R39100 a_185229_n11365.n225 a_185229_n11365.n224 9.3005
R39101 a_185229_n11365.n231 a_185229_n11365.n230 9.3005
R39102 a_185229_n11365.n229 a_185229_n11365.n228 9.3005
R39103 a_185229_n11365.n211 a_185229_n11365.n210 9.3005
R39104 a_185229_n11365.n217 a_185229_n11365.n216 9.3005
R39105 a_185229_n11365.n215 a_185229_n11365.n214 9.3005
R39106 a_185229_n11365.n197 a_185229_n11365.n196 9.3005
R39107 a_185229_n11365.n203 a_185229_n11365.n202 9.3005
R39108 a_185229_n11365.n201 a_185229_n11365.n200 9.3005
R39109 a_185229_n11365.n183 a_185229_n11365.n182 9.3005
R39110 a_185229_n11365.n189 a_185229_n11365.n188 9.3005
R39111 a_185229_n11365.n187 a_185229_n11365.n186 9.3005
R39112 a_185229_n11365.n164 a_185229_n11365.n163 9.3005
R39113 a_185229_n11365.n167 a_185229_n11365.n166 9.3005
R39114 a_185229_n11365.n154 a_185229_n11365.n153 9.3005
R39115 a_185229_n11365.n173 a_185229_n11365.n172 9.3005
R39116 a_185229_n11365.n175 a_185229_n11365.n174 9.3005
R39117 a_185229_n11365.n165 a_185229_n11365.n157 9.3005
R39118 a_185229_n11365.n10 a_185229_n11365.n8 9.3005
R39119 a_185229_n11365.n32 a_185229_n11365.n31 9.3005
R39120 a_185229_n11365.n22 a_185229_n11365.n7 9.3005
R39121 a_185229_n11365.n21 a_185229_n11365.n20 9.3005
R39122 a_185229_n11365.n19 a_185229_n11365.n18 9.3005
R39123 a_185229_n11365.n14 a_185229_n11365.n13 9.3005
R39124 a_185229_n11365.n50 a_185229_n11365.n38 9.3005
R39125 a_185229_n11365.n48 a_185229_n11365.n47 9.3005
R39126 a_185229_n11365.n46 a_185229_n11365.n45 9.3005
R39127 a_185229_n11365.n43 a_185229_n11365.n41 9.3005
R39128 a_185229_n11365.n66 a_185229_n11365.n54 9.3005
R39129 a_185229_n11365.n64 a_185229_n11365.n63 9.3005
R39130 a_185229_n11365.n62 a_185229_n11365.n61 9.3005
R39131 a_185229_n11365.n59 a_185229_n11365.n57 9.3005
R39132 a_185229_n11365.n82 a_185229_n11365.n70 9.3005
R39133 a_185229_n11365.n80 a_185229_n11365.n79 9.3005
R39134 a_185229_n11365.n78 a_185229_n11365.n77 9.3005
R39135 a_185229_n11365.n75 a_185229_n11365.n73 9.3005
R39136 a_185229_n11365.n310 a_185229_n11365.n309 8.28285
R39137 a_185229_n11365.n296 a_185229_n11365.n295 8.28285
R39138 a_185229_n11365.n282 a_185229_n11365.n281 8.28285
R39139 a_185229_n11365.n268 a_185229_n11365.n267 8.28285
R39140 a_185229_n11365.n254 a_185229_n11365.n253 8.28285
R39141 a_185229_n11365.n240 a_185229_n11365.n239 8.28285
R39142 a_185229_n11365.n226 a_185229_n11365.n225 8.28285
R39143 a_185229_n11365.n212 a_185229_n11365.n211 8.28285
R39144 a_185229_n11365.n198 a_185229_n11365.n197 8.28285
R39145 a_185229_n11365.n184 a_185229_n11365.n183 8.28285
R39146 a_185229_n11365.n176 a_185229_n11365.n154 8.28285
R39147 a_185229_n11365.n17 a_185229_n11365.n14 8.28285
R39148 a_185229_n11365.n44 a_185229_n11365.n43 8.28285
R39149 a_185229_n11365.n60 a_185229_n11365.n59 8.28285
R39150 a_185229_n11365.n76 a_185229_n11365.n75 8.28285
R39151 a_185229_n11365.n320 a_185229_n11365.n307 7.9105
R39152 a_185229_n11365.n306 a_185229_n11365.n293 7.9105
R39153 a_185229_n11365.n292 a_185229_n11365.n279 7.9105
R39154 a_185229_n11365.n278 a_185229_n11365.n265 7.9105
R39155 a_185229_n11365.n264 a_185229_n11365.n251 7.9105
R39156 a_185229_n11365.n250 a_185229_n11365.n237 7.9105
R39157 a_185229_n11365.n236 a_185229_n11365.n223 7.9105
R39158 a_185229_n11365.n222 a_185229_n11365.n209 7.9105
R39159 a_185229_n11365.n208 a_185229_n11365.n195 7.9105
R39160 a_185229_n11365.n194 a_185229_n11365.n181 7.9105
R39161 a_185229_n11365.n180 a_185229_n11365.n152 7.9105
R39162 a_185229_n11365.n34 a_185229_n11365.n6 7.9105
R39163 a_185229_n11365.n53 a_185229_n11365.n37 7.9105
R39164 a_185229_n11365.n69 a_185229_n11365.n36 7.9105
R39165 a_185229_n11365.n85 a_185229_n11365.n35 7.9105
R39166 a_185229_n11365.n85 a_185229_n11365.n84 7.9105
R39167 a_185229_n11365.n69 a_185229_n11365.n68 7.9105
R39168 a_185229_n11365.n53 a_185229_n11365.n52 7.9105
R39169 a_185229_n11365.n34 a_185229_n11365.n33 7.9105
R39170 a_185229_n11365.n180 a_185229_n11365.n179 7.9105
R39171 a_185229_n11365.n194 a_185229_n11365.n193 7.9105
R39172 a_185229_n11365.n208 a_185229_n11365.n207 7.9105
R39173 a_185229_n11365.n222 a_185229_n11365.n221 7.9105
R39174 a_185229_n11365.n236 a_185229_n11365.n235 7.9105
R39175 a_185229_n11365.n250 a_185229_n11365.n249 7.9105
R39176 a_185229_n11365.n264 a_185229_n11365.n263 7.9105
R39177 a_185229_n11365.n278 a_185229_n11365.n277 7.9105
R39178 a_185229_n11365.n292 a_185229_n11365.n291 7.9105
R39179 a_185229_n11365.n306 a_185229_n11365.n305 7.9105
R39180 a_185229_n11365.n320 a_185229_n11365.n319 7.9105
R39181 a_185229_n11365.n312 a_185229_n11365.n311 6.77697
R39182 a_185229_n11365.n298 a_185229_n11365.n297 6.77697
R39183 a_185229_n11365.n284 a_185229_n11365.n283 6.77697
R39184 a_185229_n11365.n270 a_185229_n11365.n269 6.77697
R39185 a_185229_n11365.n256 a_185229_n11365.n255 6.77697
R39186 a_185229_n11365.n242 a_185229_n11365.n241 6.77697
R39187 a_185229_n11365.n228 a_185229_n11365.n227 6.77697
R39188 a_185229_n11365.n214 a_185229_n11365.n213 6.77697
R39189 a_185229_n11365.n200 a_185229_n11365.n199 6.77697
R39190 a_185229_n11365.n186 a_185229_n11365.n185 6.77697
R39191 a_185229_n11365.n175 a_185229_n11365.n156 6.77697
R39192 a_185229_n11365.n18 a_185229_n11365.n12 6.77697
R39193 a_185229_n11365.n45 a_185229_n11365.n40 6.77697
R39194 a_185229_n11365.n61 a_185229_n11365.n56 6.77697
R39195 a_185229_n11365.n77 a_185229_n11365.n72 6.77697
R39196 a_185229_n11365.n317 a_185229_n11365.t10 5.7135
R39197 a_185229_n11365.n317 a_185229_n11365.t21 5.7135
R39198 a_185229_n11365.n303 a_185229_n11365.t18 5.7135
R39199 a_185229_n11365.n303 a_185229_n11365.t15 5.7135
R39200 a_185229_n11365.n289 a_185229_n11365.t23 5.7135
R39201 a_185229_n11365.n289 a_185229_n11365.t20 5.7135
R39202 a_185229_n11365.n275 a_185229_n11365.t5 5.7135
R39203 a_185229_n11365.n275 a_185229_n11365.t22 5.7135
R39204 a_185229_n11365.n261 a_185229_n11365.t14 5.7135
R39205 a_185229_n11365.n261 a_185229_n11365.t8 5.7135
R39206 a_185229_n11365.n247 a_185229_n11365.t3 5.7135
R39207 a_185229_n11365.n247 a_185229_n11365.t17 5.7135
R39208 a_185229_n11365.n233 a_185229_n11365.t11 5.7135
R39209 a_185229_n11365.n233 a_185229_n11365.t7 5.7135
R39210 a_185229_n11365.n219 a_185229_n11365.t19 5.7135
R39211 a_185229_n11365.n219 a_185229_n11365.t16 5.7135
R39212 a_185229_n11365.n205 a_185229_n11365.t12 5.7135
R39213 a_185229_n11365.n205 a_185229_n11365.t4 5.7135
R39214 a_185229_n11365.n191 a_185229_n11365.t6 5.7135
R39215 a_185229_n11365.n191 a_185229_n11365.t13 5.7135
R39216 a_185229_n11365.n151 a_185229_n11365.n150 5.58552
R39217 a_185229_n11365.n322 a_185229_n11365.n321 5.58552
R39218 a_185229_n11365.n26 a_185229_n11365.n8 5.33935
R39219 a_185229_n11365.n172 a_185229_n11365.n171 5.27109
R39220 a_185229_n11365.n23 a_185229_n11365.n21 5.27109
R39221 a_185229_n11365.n49 a_185229_n11365.n48 5.27109
R39222 a_185229_n11365.n65 a_185229_n11365.n64 5.27109
R39223 a_185229_n11365.n81 a_185229_n11365.n80 5.27109
R39224 a_185229_n11365.n164 a_185229_n11365.n160 4.51911
R39225 a_185229_n11365.n151 a_185229_n11365.n85 3.82472
R39226 a_185229_n11365.n321 a_185229_n11365.n34 3.80493
R39227 a_185229_n11365.n168 a_185229_n11365.n157 3.76521
R39228 a_185229_n11365.n22 a_185229_n11365.n9 3.76521
R39229 a_185229_n11365.n52 a_185229_n11365.n51 3.75827
R39230 a_185229_n11365.n68 a_185229_n11365.n67 3.75827
R39231 a_185229_n11365.n84 a_185229_n11365.n83 3.75827
R39232 a_185229_n11365.n39 a_185229_n11365.t24 3.4805
R39233 a_185229_n11365.n39 a_185229_n11365.t31 3.4805
R39234 a_185229_n11365.n55 a_185229_n11365.t26 3.4805
R39235 a_185229_n11365.n55 a_185229_n11365.t0 3.4805
R39236 a_185229_n11365.n71 a_185229_n11365.t27 3.4805
R39237 a_185229_n11365.n71 a_185229_n11365.t28 3.4805
R39238 a_185229_n11365.n316 a_185229_n11365.n307 3.43565
R39239 a_185229_n11365.n302 a_185229_n11365.n293 3.43565
R39240 a_185229_n11365.n288 a_185229_n11365.n279 3.43565
R39241 a_185229_n11365.n274 a_185229_n11365.n265 3.43565
R39242 a_185229_n11365.n260 a_185229_n11365.n251 3.43565
R39243 a_185229_n11365.n246 a_185229_n11365.n237 3.43565
R39244 a_185229_n11365.n232 a_185229_n11365.n223 3.43565
R39245 a_185229_n11365.n218 a_185229_n11365.n209 3.43565
R39246 a_185229_n11365.n204 a_185229_n11365.n195 3.43565
R39247 a_185229_n11365.n190 a_185229_n11365.n181 3.43565
R39248 a_185229_n11365.n91 a_185229_n11365.t30 2.84983
R39249 a_185229_n11365.t2 a_185229_n11365.n336 2.83411
R39250 a_185229_n11365.n91 a_185229_n11365.t29 2.7853
R39251 a_185229_n11365.n336 a_185229_n11365.t25 2.77004
R39252 a_185229_n11365.n167 a_185229_n11365.n159 2.25932
R39253 a_185229_n11365.n31 a_185229_n11365.n30 2.25932
R39254 a_185229_n11365.n321 a_185229_n11365.n320 1.75537
R39255 a_185229_n11365.n180 a_185229_n11365.n151 1.72874
R39256 a_185229_n11365.n93 a_185229_n11365.n92 1.11019
R39257 a_185229_n11365.n335 a_185229_n11365.n334 1.09519
R39258 a_185229_n11365.n92 a_185229_n11365.n90 1.06331
R39259 a_185229_n11365.n335 a_185229_n11365.n0 1.04831
R39260 a_185229_n11365.n163 a_185229_n11365.n162 0.753441
R39261 a_185229_n11365.n27 a_185229_n11365.n10 0.753441
R39262 a_185229_n11365.n327 a_185229_n11365.n3 0.3955
R39263 a_185229_n11365.n328 a_185229_n11365.n327 0.3955
R39264 a_185229_n11365.n329 a_185229_n11365.n328 0.3955
R39265 a_185229_n11365.n329 a_185229_n11365.n1 0.3955
R39266 a_185229_n11365.n333 a_185229_n11365.n1 0.3955
R39267 a_185229_n11365.n334 a_185229_n11365.n333 0.3955
R39268 a_185229_n11365.n145 a_185229_n11365.n87 0.3955
R39269 a_185229_n11365.n145 a_185229_n11365.n144 0.3955
R39270 a_185229_n11365.n144 a_185229_n11365.n143 0.3955
R39271 a_185229_n11365.n143 a_185229_n11365.n104 0.3955
R39272 a_185229_n11365.n139 a_185229_n11365.n104 0.3955
R39273 a_185229_n11365.n139 a_185229_n11365.n138 0.3955
R39274 a_185229_n11365.n138 a_185229_n11365.n137 0.3955
R39275 a_185229_n11365.n137 a_185229_n11365.n106 0.3955
R39276 a_185229_n11365.n133 a_185229_n11365.n106 0.3955
R39277 a_185229_n11365.n133 a_185229_n11365.n132 0.3955
R39278 a_185229_n11365.n132 a_185229_n11365.n131 0.3955
R39279 a_185229_n11365.n131 a_185229_n11365.n108 0.3955
R39280 a_185229_n11365.n127 a_185229_n11365.n108 0.3955
R39281 a_185229_n11365.n127 a_185229_n11365.n126 0.3955
R39282 a_185229_n11365.n126 a_185229_n11365.n125 0.3955
R39283 a_185229_n11365.n125 a_185229_n11365.n110 0.3955
R39284 a_185229_n11365.n121 a_185229_n11365.n110 0.3955
R39285 a_185229_n11365.n121 a_185229_n11365.n120 0.3955
R39286 a_185229_n11365.n120 a_185229_n11365.n119 0.3955
R39287 a_185229_n11365.n119 a_185229_n11365.n112 0.3955
R39288 a_185229_n11365.n115 a_185229_n11365.n112 0.3955
R39289 a_185229_n11365.n115 a_185229_n11365.n114 0.3955
R39290 a_185229_n11365.n114 a_185229_n11365.n5 0.3955
R39291 a_185229_n11365.n94 a_185229_n11365.n93 0.3955
R39292 a_185229_n11365.n94 a_185229_n11365.n89 0.3955
R39293 a_185229_n11365.n98 a_185229_n11365.n89 0.3955
R39294 a_185229_n11365.n99 a_185229_n11365.n98 0.3955
R39295 a_185229_n11365.n100 a_185229_n11365.n99 0.3955
R39296 a_185229_n11365.n100 a_185229_n11365.n86 0.3955
R39297 a_185229_n11365.n95 a_185229_n11365.n90 0.3955
R39298 a_185229_n11365.n96 a_185229_n11365.n95 0.3955
R39299 a_185229_n11365.n97 a_185229_n11365.n96 0.3955
R39300 a_185229_n11365.n97 a_185229_n11365.n88 0.3955
R39301 a_185229_n11365.n101 a_185229_n11365.n88 0.3955
R39302 a_185229_n11365.n102 a_185229_n11365.n101 0.3955
R39303 a_185229_n11365.n148 a_185229_n11365.n102 0.3955
R39304 a_185229_n11365.n148 a_185229_n11365.n147 0.3955
R39305 a_185229_n11365.n147 a_185229_n11365.n146 0.3955
R39306 a_185229_n11365.n146 a_185229_n11365.n103 0.3955
R39307 a_185229_n11365.n142 a_185229_n11365.n103 0.3955
R39308 a_185229_n11365.n142 a_185229_n11365.n141 0.3955
R39309 a_185229_n11365.n141 a_185229_n11365.n140 0.3955
R39310 a_185229_n11365.n140 a_185229_n11365.n105 0.3955
R39311 a_185229_n11365.n136 a_185229_n11365.n105 0.3955
R39312 a_185229_n11365.n136 a_185229_n11365.n135 0.3955
R39313 a_185229_n11365.n135 a_185229_n11365.n134 0.3955
R39314 a_185229_n11365.n134 a_185229_n11365.n107 0.3955
R39315 a_185229_n11365.n130 a_185229_n11365.n107 0.3955
R39316 a_185229_n11365.n130 a_185229_n11365.n129 0.3955
R39317 a_185229_n11365.n129 a_185229_n11365.n128 0.3955
R39318 a_185229_n11365.n128 a_185229_n11365.n109 0.3955
R39319 a_185229_n11365.n124 a_185229_n11365.n109 0.3955
R39320 a_185229_n11365.n124 a_185229_n11365.n123 0.3955
R39321 a_185229_n11365.n123 a_185229_n11365.n122 0.3955
R39322 a_185229_n11365.n122 a_185229_n11365.n111 0.3955
R39323 a_185229_n11365.n118 a_185229_n11365.n111 0.3955
R39324 a_185229_n11365.n118 a_185229_n11365.n117 0.3955
R39325 a_185229_n11365.n117 a_185229_n11365.n116 0.3955
R39326 a_185229_n11365.n116 a_185229_n11365.n113 0.3955
R39327 a_185229_n11365.n113 a_185229_n11365.n4 0.3955
R39328 a_185229_n11365.n324 a_185229_n11365.n4 0.3955
R39329 a_185229_n11365.n325 a_185229_n11365.n324 0.3955
R39330 a_185229_n11365.n326 a_185229_n11365.n325 0.3955
R39331 a_185229_n11365.n326 a_185229_n11365.n2 0.3955
R39332 a_185229_n11365.n330 a_185229_n11365.n2 0.3955
R39333 a_185229_n11365.n331 a_185229_n11365.n330 0.3955
R39334 a_185229_n11365.n332 a_185229_n11365.n331 0.3955
R39335 a_185229_n11365.n332 a_185229_n11365.n0 0.3955
R39336 a_185229_n11365.n323 a_185229_n11365.n5 0.370955
R39337 a_185229_n11365.n149 a_185229_n11365.n87 0.351864
R39338 a_185229_n11365.n92 a_185229_n11365.n91 0.349638
R39339 a_185229_n11365.n336 a_185229_n11365.n335 0.349638
R39340 a_185229_n11365.n314 a_185229_n11365.n313 0.196152
R39341 a_185229_n11365.n300 a_185229_n11365.n299 0.196152
R39342 a_185229_n11365.n286 a_185229_n11365.n285 0.196152
R39343 a_185229_n11365.n272 a_185229_n11365.n271 0.196152
R39344 a_185229_n11365.n258 a_185229_n11365.n257 0.196152
R39345 a_185229_n11365.n244 a_185229_n11365.n243 0.196152
R39346 a_185229_n11365.n230 a_185229_n11365.n229 0.196152
R39347 a_185229_n11365.n216 a_185229_n11365.n215 0.196152
R39348 a_185229_n11365.n202 a_185229_n11365.n201 0.196152
R39349 a_185229_n11365.n188 a_185229_n11365.n187 0.196152
R39350 a_185229_n11365.n166 a_185229_n11365.n164 0.196152
R39351 a_185229_n11365.n174 a_185229_n11365.n173 0.196152
R39352 a_185229_n11365.n20 a_185229_n11365.n19 0.196152
R39353 a_185229_n11365.n20 a_185229_n11365.n7 0.196152
R39354 a_185229_n11365.n47 a_185229_n11365.n46 0.196152
R39355 a_185229_n11365.n47 a_185229_n11365.n38 0.196152
R39356 a_185229_n11365.n63 a_185229_n11365.n62 0.196152
R39357 a_185229_n11365.n63 a_185229_n11365.n54 0.196152
R39358 a_185229_n11365.n79 a_185229_n11365.n78 0.196152
R39359 a_185229_n11365.n79 a_185229_n11365.n70 0.196152
R39360 a_185229_n11365.n166 a_185229_n11365.n165 0.194824
R39361 a_185229_n11365.n313 a_185229_n11365.n308 0.186853
R39362 a_185229_n11365.n299 a_185229_n11365.n294 0.186853
R39363 a_185229_n11365.n285 a_185229_n11365.n280 0.186853
R39364 a_185229_n11365.n271 a_185229_n11365.n266 0.186853
R39365 a_185229_n11365.n257 a_185229_n11365.n252 0.186853
R39366 a_185229_n11365.n243 a_185229_n11365.n238 0.186853
R39367 a_185229_n11365.n229 a_185229_n11365.n224 0.186853
R39368 a_185229_n11365.n215 a_185229_n11365.n210 0.186853
R39369 a_185229_n11365.n201 a_185229_n11365.n196 0.186853
R39370 a_185229_n11365.n187 a_185229_n11365.n182 0.186853
R39371 a_185229_n11365.n174 a_185229_n11365.n153 0.186853
R39372 a_185229_n11365.n19 a_185229_n11365.n13 0.186853
R39373 a_185229_n11365.n46 a_185229_n11365.n41 0.186853
R39374 a_185229_n11365.n62 a_185229_n11365.n57 0.186853
R39375 a_185229_n11365.n78 a_185229_n11365.n73 0.186853
R39376 a_185229_n11365.n32 a_185229_n11365.n8 0.184196
R39377 a_185229_n11365.n150 a_185229_n11365.n86 0.166409
R39378 a_185229_n11365.n322 a_185229_n11365.n3 0.131409
R39379 a_185229_n11365.n33 a_185229_n11365.n7 0.0790024
R39380 a_185229_n11365.n52 a_185229_n11365.n38 0.0790024
R39381 a_185229_n11365.n68 a_185229_n11365.n54 0.0790024
R39382 a_185229_n11365.n84 a_185229_n11365.n70 0.0790024
R39383 a_185229_n11365.n323 a_185229_n11365.n322 0.0709545
R39384 a_185229_n11365.n314 a_185229_n11365.n307 0.0572633
R39385 a_185229_n11365.n300 a_185229_n11365.n293 0.0572633
R39386 a_185229_n11365.n286 a_185229_n11365.n279 0.0572633
R39387 a_185229_n11365.n272 a_185229_n11365.n265 0.0572633
R39388 a_185229_n11365.n258 a_185229_n11365.n251 0.0572633
R39389 a_185229_n11365.n244 a_185229_n11365.n237 0.0572633
R39390 a_185229_n11365.n230 a_185229_n11365.n223 0.0572633
R39391 a_185229_n11365.n216 a_185229_n11365.n209 0.0572633
R39392 a_185229_n11365.n202 a_185229_n11365.n195 0.0572633
R39393 a_185229_n11365.n188 a_185229_n11365.n181 0.0572633
R39394 a_185229_n11365.n173 a_185229_n11365.n152 0.0572633
R39395 a_185229_n11365.n150 a_185229_n11365.n149 0.0550455
R39396 a_185229_n11365.n208 a_185229_n11365.n194 0.0506333
R39397 a_185229_n11365.n222 a_185229_n11365.n208 0.0506333
R39398 a_185229_n11365.n250 a_185229_n11365.n236 0.0506333
R39399 a_185229_n11365.n278 a_185229_n11365.n264 0.0506333
R39400 a_185229_n11365.n292 a_185229_n11365.n278 0.0506333
R39401 a_185229_n11365.n320 a_185229_n11365.n306 0.0506333
R39402 a_185229_n11365.n194 a_185229_n11365.n180 0.0490667
R39403 a_185229_n11365.n236 a_185229_n11365.n222 0.0490667
R39404 a_185229_n11365.n264 a_185229_n11365.n250 0.0490667
R39405 a_185229_n11365.n306 a_185229_n11365.n292 0.0490667
R39406 a_185229_n11365.n165 a_185229_n11365.n152 0.0477222
R39407 a_185229_n11365.n85 a_185229_n11365.n69 0.0400789
R39408 a_185229_n11365.n53 a_185229_n11365.n34 0.0400789
R39409 a_185229_n11365.n319 a_185229_n11365.n308 0.0393889
R39410 a_185229_n11365.n305 a_185229_n11365.n294 0.0393889
R39411 a_185229_n11365.n291 a_185229_n11365.n280 0.0393889
R39412 a_185229_n11365.n277 a_185229_n11365.n266 0.0393889
R39413 a_185229_n11365.n263 a_185229_n11365.n252 0.0393889
R39414 a_185229_n11365.n249 a_185229_n11365.n238 0.0393889
R39415 a_185229_n11365.n235 a_185229_n11365.n224 0.0393889
R39416 a_185229_n11365.n221 a_185229_n11365.n210 0.0393889
R39417 a_185229_n11365.n207 a_185229_n11365.n196 0.0393889
R39418 a_185229_n11365.n193 a_185229_n11365.n182 0.0393889
R39419 a_185229_n11365.n179 a_185229_n11365.n153 0.0393889
R39420 a_185229_n11365.n13 a_185229_n11365.n6 0.0393889
R39421 a_185229_n11365.n41 a_185229_n11365.n37 0.0393889
R39422 a_185229_n11365.n57 a_185229_n11365.n36 0.0393889
R39423 a_185229_n11365.n73 a_185229_n11365.n35 0.0393889
R39424 a_185229_n11365.n69 a_185229_n11365.n53 0.0388421
R39425 a_185229_n11365.n33 a_185229_n11365.n32 0.0366111
R39426 C2S2_Amp_F_I_0.VN.t10 C2S2_Amp_F_I_0.VN.n12 428.81
R39427 C2S2_Amp_F_I_0.VN.n24 C2S2_Amp_F_I_0.VN.t10 428.81
R39428 C2S2_Amp_F_I_0.VN.t5 C2S2_Amp_F_I_0.VN.n22 428.81
R39429 C2S2_Amp_F_I_0.VN.n23 C2S2_Amp_F_I_0.VN.t5 428.81
R39430 C2S2_Amp_F_I_0.VN.n21 C2S2_Amp_F_I_0.VN.t2 428.81
R39431 C2S2_Amp_F_I_0.VN.t2 C2S2_Amp_F_I_0.VN.n13 428.81
R39432 C2S2_Amp_F_I_0.VN.n20 C2S2_Amp_F_I_0.VN.t16 428.81
R39433 C2S2_Amp_F_I_0.VN.t16 C2S2_Amp_F_I_0.VN.n19 428.81
R39434 C2S2_Amp_F_I_0.VN.t14 C2S2_Amp_F_I_0.VN.n14 428.81
R39435 C2S2_Amp_F_I_0.VN.n18 C2S2_Amp_F_I_0.VN.t14 428.81
R39436 C2S2_Amp_F_I_0.VN.t9 C2S2_Amp_F_I_0.VN.n16 428.81
R39437 C2S2_Amp_F_I_0.VN.n17 C2S2_Amp_F_I_0.VN.t9 428.81
R39438 C2S2_Amp_F_I_0.VN.n15 C2S2_Amp_F_I_0.VN.t4 213.694
R39439 C2S2_Amp_F_I_0.VN.n26 C2S2_Amp_F_I_0.VN.n11 5.65673
R39440 C2S2_Amp_F_I_0.VN.n27 C2S2_Amp_F_I_0.VN.t0 3.80966
R39441 C2S2_Amp_F_I_0.VN.n11 C2S2_Amp_F_I_0.VN.t1 3.63099
R39442 C2S2_Amp_F_I_0.VN.n26 C2S2_Amp_F_I_0.VN.n25 3.35505
R39443 C2S2_Amp_F_I_0.VN.n16 C2S2_Amp_F_I_0.VN.n15 1.82094
R39444 C2S2_Amp_F_I_0.VN.n17 C2S2_Amp_F_I_0.VN.n15 1.82094
R39445 C2S2_Amp_F_I_0.VN.n25 C2S2_Amp_F_I_0.VN.n24 1.29456
R39446 C2S2_Amp_F_I_0.VN.n25 C2S2_Amp_F_I_0.VN.n12 1.29456
R39447 C2S2_Amp_F_I_0.VN.n6 C2S2_Amp_F_I_0.VN.n2 0.653665
R39448 C2S2_Amp_F_I_0.VN.n10 C2S2_Amp_F_I_0.VN.n6 0.447
R39449 C2S2_Amp_F_I_0.VN.n18 C2S2_Amp_F_I_0.VN.n17 0.3955
R39450 C2S2_Amp_F_I_0.VN.n19 C2S2_Amp_F_I_0.VN.n18 0.3955
R39451 C2S2_Amp_F_I_0.VN.n19 C2S2_Amp_F_I_0.VN.n13 0.3955
R39452 C2S2_Amp_F_I_0.VN.n23 C2S2_Amp_F_I_0.VN.n13 0.3955
R39453 C2S2_Amp_F_I_0.VN.n24 C2S2_Amp_F_I_0.VN.n23 0.3955
R39454 C2S2_Amp_F_I_0.VN.n16 C2S2_Amp_F_I_0.VN.n14 0.3955
R39455 C2S2_Amp_F_I_0.VN.n20 C2S2_Amp_F_I_0.VN.n14 0.3955
R39456 C2S2_Amp_F_I_0.VN.n21 C2S2_Amp_F_I_0.VN.n20 0.3955
R39457 C2S2_Amp_F_I_0.VN.n22 C2S2_Amp_F_I_0.VN.n21 0.3955
R39458 C2S2_Amp_F_I_0.VN.n22 C2S2_Amp_F_I_0.VN.n12 0.3955
R39459 C2S2_Amp_F_I_0.VN.n11 C2S2_Amp_F_I_0.VN.n10 0.29378
R39460 C2S2_Amp_F_I_0.VN.n10 C2S2_Amp_F_I_0.VN.n9 0.230665
R39461 C2S2_Amp_F_I_0.VN.n6 C2S2_Amp_F_I_0.VN.n5 0.230665
R39462 C2S2_Amp_F_I_0.VN.n7 C2S2_Amp_F_I_0.VN.t17 0.230482
R39463 C2S2_Amp_F_I_0.VN.n3 C2S2_Amp_F_I_0.VN.t12 0.230482
R39464 C2S2_Amp_F_I_0.VN.n0 C2S2_Amp_F_I_0.VN.t11 0.230482
R39465 C2S2_Amp_F_I_0.VN.n8 C2S2_Amp_F_I_0.VN.n7 0.227365
R39466 C2S2_Amp_F_I_0.VN.n9 C2S2_Amp_F_I_0.VN.n8 0.227365
R39467 C2S2_Amp_F_I_0.VN.n4 C2S2_Amp_F_I_0.VN.n3 0.227365
R39468 C2S2_Amp_F_I_0.VN.n5 C2S2_Amp_F_I_0.VN.n4 0.227365
R39469 C2S2_Amp_F_I_0.VN.n1 C2S2_Amp_F_I_0.VN.n0 0.227365
R39470 C2S2_Amp_F_I_0.VN.n2 C2S2_Amp_F_I_0.VN.n1 0.227365
R39471 C2S2_Amp_F_I_0.VN C2S2_Amp_F_I_0.VN.n27 0.132871
R39472 C2S2_Amp_F_I_0.VN.n27 C2S2_Amp_F_I_0.VN.n26 0.0719985
R39473 C2S2_Amp_F_I_0.VN.n7 C2S2_Amp_F_I_0.VN.t19 0.00361634
R39474 C2S2_Amp_F_I_0.VN.n8 C2S2_Amp_F_I_0.VN.t8 0.00361634
R39475 C2S2_Amp_F_I_0.VN.n9 C2S2_Amp_F_I_0.VN.t3 0.00361634
R39476 C2S2_Amp_F_I_0.VN.n3 C2S2_Amp_F_I_0.VN.t15 0.00361634
R39477 C2S2_Amp_F_I_0.VN.n4 C2S2_Amp_F_I_0.VN.t7 0.00361634
R39478 C2S2_Amp_F_I_0.VN.n5 C2S2_Amp_F_I_0.VN.t20 0.00361634
R39479 C2S2_Amp_F_I_0.VN.n0 C2S2_Amp_F_I_0.VN.t13 0.00361634
R39480 C2S2_Amp_F_I_0.VN.n1 C2S2_Amp_F_I_0.VN.t6 0.00361634
R39481 C2S2_Amp_F_I_0.VN.n2 C2S2_Amp_F_I_0.VN.t18 0.00361634
R39482 VMID.t2 VMID.n34 428.81
R39483 VMID.n35 VMID.t2 428.81
R39484 VMID.t18 VMID.n32 428.81
R39485 VMID.n36 VMID.t18 428.81
R39486 VMID.n38 VMID.t13 428.81
R39487 VMID.t13 VMID.n37 428.81
R39488 VMID.n39 VMID.t1 428.81
R39489 VMID.t1 VMID.n31 428.81
R39490 VMID.t16 VMID.n40 428.81
R39491 VMID.n41 VMID.t16 428.81
R39492 VMID.t8 VMID.n30 428.81
R39493 VMID.n42 VMID.t8 428.81
R39494 VMID.t9 VMID.n19 428.81
R39495 VMID.n20 VMID.t9 428.81
R39496 VMID.t6 VMID.n17 428.81
R39497 VMID.n21 VMID.t6 428.81
R39498 VMID.n23 VMID.t0 428.81
R39499 VMID.t0 VMID.n22 428.81
R39500 VMID.n24 VMID.t20 428.81
R39501 VMID.t20 VMID.n16 428.81
R39502 VMID.t15 VMID.n25 428.81
R39503 VMID.n26 VMID.t15 428.81
R39504 VMID.t7 VMID.n15 428.81
R39505 VMID.n27 VMID.t7 428.81
R39506 VMID.t3 VMID.n4 428.81
R39507 VMID.n5 VMID.t3 428.81
R39508 VMID.t19 VMID.n2 428.81
R39509 VMID.n6 VMID.t19 428.81
R39510 VMID.n8 VMID.t4 428.81
R39511 VMID.t4 VMID.n7 428.81
R39512 VMID.n9 VMID.t14 428.81
R39513 VMID.t14 VMID.n1 428.81
R39514 VMID.t12 VMID.n10 428.81
R39515 VMID.n11 VMID.t12 428.81
R39516 VMID.t10 VMID.n0 428.81
R39517 VMID.n12 VMID.t10 428.81
R39518 VMID.n33 VMID.t11 213.691
R39519 VMID.n18 VMID.t17 213.691
R39520 VMID.n3 VMID.t5 213.691
R39521 VMID VMID.n43 3.42832
R39522 VMID VMID.n28 3.42832
R39523 VMID.n14 VMID.n13 3.17512
R39524 VMID.n35 VMID.n33 1.8259
R39525 VMID.n34 VMID.n33 1.8259
R39526 VMID.n20 VMID.n18 1.8259
R39527 VMID.n19 VMID.n18 1.8259
R39528 VMID.n5 VMID.n3 1.8259
R39529 VMID.n4 VMID.n3 1.8259
R39530 VMID.n43 VMID.n42 1.28956
R39531 VMID.n43 VMID.n30 1.28956
R39532 VMID.n28 VMID.n27 1.28956
R39533 VMID.n28 VMID.n15 1.28956
R39534 VMID.n13 VMID.n12 1.28956
R39535 VMID.n13 VMID.n0 1.28956
R39536 VMID.n29 VMID.n14 0.714177
R39537 VMID VMID.n44 0.519463
R39538 VMID.n42 VMID.n41 0.3955
R39539 VMID.n41 VMID.n31 0.3955
R39540 VMID.n37 VMID.n31 0.3955
R39541 VMID.n37 VMID.n36 0.3955
R39542 VMID.n36 VMID.n35 0.3955
R39543 VMID.n40 VMID.n30 0.3955
R39544 VMID.n40 VMID.n39 0.3955
R39545 VMID.n39 VMID.n38 0.3955
R39546 VMID.n38 VMID.n32 0.3955
R39547 VMID.n34 VMID.n32 0.3955
R39548 VMID.n27 VMID.n26 0.3955
R39549 VMID.n26 VMID.n16 0.3955
R39550 VMID.n22 VMID.n16 0.3955
R39551 VMID.n22 VMID.n21 0.3955
R39552 VMID.n21 VMID.n20 0.3955
R39553 VMID.n25 VMID.n15 0.3955
R39554 VMID.n25 VMID.n24 0.3955
R39555 VMID.n24 VMID.n23 0.3955
R39556 VMID.n23 VMID.n17 0.3955
R39557 VMID.n19 VMID.n17 0.3955
R39558 VMID.n12 VMID.n11 0.3955
R39559 VMID.n11 VMID.n1 0.3955
R39560 VMID.n7 VMID.n1 0.3955
R39561 VMID.n7 VMID.n6 0.3955
R39562 VMID.n6 VMID.n5 0.3955
R39563 VMID.n10 VMID.n0 0.3955
R39564 VMID.n10 VMID.n9 0.3955
R39565 VMID.n9 VMID.n8 0.3955
R39566 VMID.n8 VMID.n2 0.3955
R39567 VMID.n4 VMID.n2 0.3955
R39568 VMID.n44 VMID 0.277896
R39569 VMID.n29 VMID 0.268496
R39570 VMID.n14 VMID 0.253961
R39571 VMID VMID.n29 0.0551768
R39572 VMID.n44 VMID 0.0171143
R39573 a_150997_n11365.n1 a_150997_n11365.n0 7.70214
R39574 a_150997_n11365.n5 a_150997_n11365.n4 7.69294
R39575 a_150997_n11365.n0 a_150997_n11365.t6 2.81388
R39576 a_150997_n11365.n0 a_150997_n11365.t7 2.81161
R39577 a_150997_n11365.n5 a_150997_n11365.t1 2.80271
R39578 a_150997_n11365.t0 a_150997_n11365.n5 2.80144
R39579 a_150997_n11365.n4 a_150997_n11365.n3 0.522904
R39580 a_150997_n11365.n3 a_150997_n11365.n2 0.522904
R39581 a_150997_n11365.n2 a_150997_n11365.n1 0.522904
R39582 a_150997_n11365.n4 a_150997_n11365.t2 0.0535478
R39583 a_150997_n11365.n3 a_150997_n11365.t5 0.0535478
R39584 a_150997_n11365.n2 a_150997_n11365.t4 0.0535478
R39585 a_150997_n11365.n1 a_150997_n11365.t3 0.0535478
R39586 a_186826_n27776.n6 a_186826_n27776.n5 22.4024
R39587 a_186826_n27776.n7 a_186826_n27776.n2 18.9924
R39588 a_186826_n27776.n4 a_186826_n27776.n3 18.9924
R39589 a_186826_n27776.n7 a_186826_n27776.n6 3.716
R39590 a_186826_n27776.n6 a_186826_n27776.n4 3.71013
R39591 a_186826_n27776.n3 a_186826_n27776.t4 3.4805
R39592 a_186826_n27776.n3 a_186826_n27776.t3 3.4805
R39593 a_186826_n27776.n2 a_186826_n27776.t5 3.4805
R39594 a_186826_n27776.n2 a_186826_n27776.t6 3.4805
R39595 a_186826_n27776.n5 a_186826_n27776.t2 3.4805
R39596 a_186826_n27776.n5 a_186826_n27776.t7 3.4805
R39597 a_186826_n27776.t0 a_186826_n27776.n9 3.04188
R39598 a_186826_n27776.n0 a_186826_n27776.t8 3.03453
R39599 a_186826_n27776.n0 a_186826_n27776.t9 2.59419
R39600 a_186826_n27776.n9 a_186826_n27776.t1 2.59419
R39601 a_186826_n27776.n8 a_186826_n27776.n7 2.55108
R39602 a_186826_n27776.n4 a_186826_n27776.n1 2.55108
R39603 a_186826_n27776.n8 a_186826_n27776.n1 0.293114
R39604 a_186826_n27776.n9 a_186826_n27776.n8 0.078625
R39605 a_186826_n27776.n1 a_186826_n27776.n0 0.0672614
R39606 a_182797_n11365.n5 a_182797_n11365.n4 7.70214
R39607 a_182797_n11365.n1 a_182797_n11365.n0 7.69294
R39608 a_182797_n11365.n5 a_182797_n11365.t1 2.81388
R39609 a_182797_n11365.t0 a_182797_n11365.n5 2.81161
R39610 a_182797_n11365.n0 a_182797_n11365.t6 2.80271
R39611 a_182797_n11365.n0 a_182797_n11365.t7 2.80044
R39612 a_182797_n11365.n2 a_182797_n11365.n1 0.522904
R39613 a_182797_n11365.n3 a_182797_n11365.n2 0.522904
R39614 a_182797_n11365.n4 a_182797_n11365.n3 0.522904
R39615 a_182797_n11365.n1 a_182797_n11365.t4 0.0535478
R39616 a_182797_n11365.n2 a_182797_n11365.t5 0.0535478
R39617 a_182797_n11365.n3 a_182797_n11365.t3 0.0535478
R39618 a_182797_n11365.n4 a_182797_n11365.t2 0.0535478
R39619 C2S2_Amp_F_I_1.VN.t6 C2S2_Amp_F_I_1.VN.n14 428.81
R39620 C2S2_Amp_F_I_1.VN.n26 C2S2_Amp_F_I_1.VN.t6 428.81
R39621 C2S2_Amp_F_I_1.VN.t19 C2S2_Amp_F_I_1.VN.n24 428.81
R39622 C2S2_Amp_F_I_1.VN.n25 C2S2_Amp_F_I_1.VN.t19 428.81
R39623 C2S2_Amp_F_I_1.VN.n23 C2S2_Amp_F_I_1.VN.t14 428.81
R39624 C2S2_Amp_F_I_1.VN.t14 C2S2_Amp_F_I_1.VN.n15 428.81
R39625 C2S2_Amp_F_I_1.VN.n22 C2S2_Amp_F_I_1.VN.t10 428.81
R39626 C2S2_Amp_F_I_1.VN.t10 C2S2_Amp_F_I_1.VN.n21 428.81
R39627 C2S2_Amp_F_I_1.VN.t17 C2S2_Amp_F_I_1.VN.n16 428.81
R39628 C2S2_Amp_F_I_1.VN.n20 C2S2_Amp_F_I_1.VN.t17 428.81
R39629 C2S2_Amp_F_I_1.VN.t13 C2S2_Amp_F_I_1.VN.n18 428.81
R39630 C2S2_Amp_F_I_1.VN.n19 C2S2_Amp_F_I_1.VN.t13 428.81
R39631 C2S2_Amp_F_I_1.VN.n17 C2S2_Amp_F_I_1.VN.t2 213.694
R39632 C2S2_Amp_F_I_1.VN.n13 C2S2_Amp_F_I_1.VN.n12 5.71607
R39633 C2S2_Amp_F_I_1.VN.n12 C2S2_Amp_F_I_1.VN.t0 3.63037
R39634 C2S2_Amp_F_I_1.VN.n29 C2S2_Amp_F_I_1.VN.t1 3.58673
R39635 C2S2_Amp_F_I_1.VN.n28 C2S2_Amp_F_I_1.VN.n27 3.38152
R39636 C2S2_Amp_F_I_1.VN.n18 C2S2_Amp_F_I_1.VN.n17 1.82094
R39637 C2S2_Amp_F_I_1.VN.n19 C2S2_Amp_F_I_1.VN.n17 1.82094
R39638 C2S2_Amp_F_I_1.VN.n27 C2S2_Amp_F_I_1.VN.n26 1.29456
R39639 C2S2_Amp_F_I_1.VN.n27 C2S2_Amp_F_I_1.VN.n14 1.29456
R39640 C2S2_Amp_F_I_1.VN.n30 C2S2_Amp_F_I_1.VN.n29 0.853
R39641 C2S2_Amp_F_I_1.VN.n29 C2S2_Amp_F_I_1.VN.n28 0.853
R39642 C2S2_Amp_F_I_1.VN.n7 C2S2_Amp_F_I_1.VN.n3 0.677282
R39643 C2S2_Amp_F_I_1.VN.n11 C2S2_Amp_F_I_1.VN.n7 0.447
R39644 C2S2_Amp_F_I_1.VN.n13 C2S2_Amp_F_I_1.VN.n0 0.422647
R39645 C2S2_Amp_F_I_1.VN.n20 C2S2_Amp_F_I_1.VN.n19 0.3955
R39646 C2S2_Amp_F_I_1.VN.n21 C2S2_Amp_F_I_1.VN.n20 0.3955
R39647 C2S2_Amp_F_I_1.VN.n21 C2S2_Amp_F_I_1.VN.n15 0.3955
R39648 C2S2_Amp_F_I_1.VN.n25 C2S2_Amp_F_I_1.VN.n15 0.3955
R39649 C2S2_Amp_F_I_1.VN.n26 C2S2_Amp_F_I_1.VN.n25 0.3955
R39650 C2S2_Amp_F_I_1.VN.n18 C2S2_Amp_F_I_1.VN.n16 0.3955
R39651 C2S2_Amp_F_I_1.VN.n22 C2S2_Amp_F_I_1.VN.n16 0.3955
R39652 C2S2_Amp_F_I_1.VN.n23 C2S2_Amp_F_I_1.VN.n22 0.3955
R39653 C2S2_Amp_F_I_1.VN.n24 C2S2_Amp_F_I_1.VN.n23 0.3955
R39654 C2S2_Amp_F_I_1.VN.n24 C2S2_Amp_F_I_1.VN.n14 0.3955
R39655 C2S2_Amp_F_I_1.VN.n12 C2S2_Amp_F_I_1.VN.n11 0.315518
R39656 C2S2_Amp_F_I_1.VN.n7 C2S2_Amp_F_I_1.VN.n6 0.230783
R39657 C2S2_Amp_F_I_1.VN.n11 C2S2_Amp_F_I_1.VN.n10 0.230783
R39658 C2S2_Amp_F_I_1.VN.n1 C2S2_Amp_F_I_1.VN.t12 0.230482
R39659 C2S2_Amp_F_I_1.VN.n4 C2S2_Amp_F_I_1.VN.t5 0.230482
R39660 C2S2_Amp_F_I_1.VN.n8 C2S2_Amp_F_I_1.VN.t3 0.230482
R39661 C2S2_Amp_F_I_1.VN.n2 C2S2_Amp_F_I_1.VN.n1 0.227365
R39662 C2S2_Amp_F_I_1.VN.n3 C2S2_Amp_F_I_1.VN.n2 0.227365
R39663 C2S2_Amp_F_I_1.VN.n5 C2S2_Amp_F_I_1.VN.n4 0.227365
R39664 C2S2_Amp_F_I_1.VN.n6 C2S2_Amp_F_I_1.VN.n5 0.227365
R39665 C2S2_Amp_F_I_1.VN.n9 C2S2_Amp_F_I_1.VN.n8 0.227365
R39666 C2S2_Amp_F_I_1.VN.n10 C2S2_Amp_F_I_1.VN.n9 0.227365
R39667 C2S2_Amp_F_I_1.VN C2S2_Amp_F_I_1.VN.n30 0.155038
R39668 C2S2_Amp_F_I_1.VN.n29 C2S2_Amp_F_I_1.VN.n13 0.0505
R39669 C2S2_Amp_F_I_1.VN.n30 C2S2_Amp_F_I_1.VN.n0 0.0102064
R39670 C2S2_Amp_F_I_1.VN.n28 C2S2_Amp_F_I_1.VN.n0 0.0102064
R39671 C2S2_Amp_F_I_1.VN.n1 C2S2_Amp_F_I_1.VN.t15 0.00361634
R39672 C2S2_Amp_F_I_1.VN.n2 C2S2_Amp_F_I_1.VN.t4 0.00361634
R39673 C2S2_Amp_F_I_1.VN.n3 C2S2_Amp_F_I_1.VN.t16 0.00361634
R39674 C2S2_Amp_F_I_1.VN.n4 C2S2_Amp_F_I_1.VN.t8 0.00361634
R39675 C2S2_Amp_F_I_1.VN.n5 C2S2_Amp_F_I_1.VN.t20 0.00361634
R39676 C2S2_Amp_F_I_1.VN.n6 C2S2_Amp_F_I_1.VN.t11 0.00361634
R39677 C2S2_Amp_F_I_1.VN.n8 C2S2_Amp_F_I_1.VN.t7 0.00361634
R39678 C2S2_Amp_F_I_1.VN.n9 C2S2_Amp_F_I_1.VN.t18 0.00361634
R39679 C2S2_Amp_F_I_1.VN.n10 C2S2_Amp_F_I_1.VN.t9 0.00361634
R39680 SIG.n0 SIG.t0 2.60536
R39681 SIG SIG.n0 1.48091
R39682 SIG.n1 SIG.n0 0.714972
R39683 SIG.n1 SIG 0.0154417
R39684 SIG SIG.n1 0.00993414
C0 1Bit_Clk_ADC_0.x9.A VDD 1.4234f
C1 1Bit_Clk_ADC_0.x11.A 1Bit_Clk_ADC_0.x4.B 1.39e-21
C2 a_208326_n43908# VDD 0.287749f
C3 1Bit_Clk_ADC_0.x14.Y 1Bit_Clk_ADC_0.sky130_fd_sc_hd__nand2_4_0.Y 0.472902f
C4 C2S2_Amp_F_I_1.OUT C2S2_Amp_F_I_0.OUT 0.052781f
C5 a_232625_n27343# 1Bit_Clk_ADC_0.sky130_fd_sc_hd__nand2_4_0.Y 0.001317f
C6 1Bit_Clk_ADC_0.x3.B a_230193_n27343# 0.002101f
C7 1Bit_Clk_ADC_0.x3.A VDD 1.41412f
C8 a_230137_n27658# VDD 0.035557f
C9 a_174650_n12474# VMID 0.075988f
C10 1Bit_Clk_ADC_0.x6.B CLK 0.232183f
C11 1Bit_Clk_ADC_0.x3.Y a_231797_n27343# 0.003025f
C12 1Bit_Clk_ADC_0.x14.Y a_230965_n27658# 0.016153f
C13 a_231021_n27343# CLK 0.003368f
C14 1Bit_Clk_ADC_0.x3.Y VDD 1.14384f
C15 1Bit_Clk_ADC_0.x11.A 1Bit_Clk_ADC_0.sky130_fd_sc_hd__nand2_4_0.Y 0.007114f
C16 C2S2_Amp_F_I_0.OUT VMID 2.35681f
C17 1Bit_Clk_ADC_0.x3.B a_231797_n27343# 0.007147f
C18 a_232253_n27658# VDD 0.021076f
C19 C2S2_Amp_F_I_1.OUT C2S2_Amp_F_I_0.VN 2.28282f
C20 a_177926_n46392# VDD 0.046325f
C21 1Bit_Clk_ADC_0.x3.B VDD 2.12484f
C22 1Bit_Clk_ADC_0.x14.Y CLK 0.543823f
C23 1Bit_Clk_ADC_0.x6.B a_231021_n27343# 0.0012f
C24 a_177926_n46392# 1Bit_DAC_Inv_0.OUT 0.86117f
C25 1Bit_Clk_ADC_0.x5.A 1Bit_Clk_ADC_0.x4.B 2.64e-19
C26 1Bit_Clk_ADC_0.x14.Y a_233081_n27658# 1.5e-19
C27 1Bit_Clk_ADC_0.x11.A a_230965_n27658# 0.008179f
C28 a_230193_n27343# VDD 0.03612f
C29 a_141908_n24334# a_144392_n24334# 0.30621f
C30 1Bit_Clk_ADC_0.x9.B 1Bit_Clk_ADC_0.sky130_fd_sc_hd__nand2_4_0.Y 0.264611f
C31 1Bit_Clk_ADC_0.x6.B 1Bit_Clk_ADC_0.x14.Y 0.105891f
C32 1Bit_Clk_ADC_0.sky130_fd_sc_hd__nand2_4_0.Y OUT 0.05444f
C33 a_208326_n46392# 1Bit_DAC_0.OUT 0.441661f
C34 C2S2_Amp_F_I_0.VN VMID 1.7323f
C35 a_141908_n24334# SIG 0.36427f
C36 1Bit_Clk_ADC_0.x14.Y a_231021_n27343# 0.009615f
C37 1Bit_Clk_ADC_0.x11.A CLK 4.73e-19
C38 C2S2_Amp_F_I_0.VN OUT 0.001563f
C39 a_196466_n45150# OUT 0.799391f
C40 C2S2_Amp_F_I_0.OUT a_208326_n43908# 0.001002f
C41 1Bit_Clk_ADC_0.x3.A 1Bit_Clk_ADC_0.x4.B 0.011558f
C42 1Bit_Clk_ADC_0.x4.B a_230137_n27658# 0.184132f
C43 1Bit_Clk_ADC_0.x11.A a_233081_n27658# 7.73e-19
C44 a_231797_n27343# VDD 0.019515f
C45 a_143150_n12474# C2S2_Amp_F_I_1.VN 0.34387f
C46 1Bit_Clk_ADC_0.x9.A 1Bit_Clk_ADC_0.sky130_fd_sc_hd__nand2_4_0.Y 0.010607f
C47 1Bit_Clk_ADC_0.x3.Y 1Bit_Clk_ADC_0.x4.B 0.051718f
C48 1Bit_DAC_Inv_0.OUT VDD 1.50487f
C49 1Bit_Clk_ADC_0.x14.Y a_232625_n27343# 0.003952f
C50 1Bit_Clk_ADC_0.x11.A a_231021_n27343# 3.88e-19
C51 1Bit_DAC_0.OUT VDD 1.67622f
C52 a_175892_n24334# C2S2_Amp_F_I_0.VN 0.021836f
C53 C2S2_Amp_F_I_0.VN a_208326_n43908# 0.014343f
C54 1Bit_Clk_ADC_0.x3.B 1Bit_Clk_ADC_0.x4.B 0.291994f
C55 1Bit_Clk_ADC_0.x9.B a_233081_n27658# 0.200111f
C56 a_233081_n27658# OUT 0.080702f
C57 C2S2_Amp_F_I_1.VN VDD 0.13086f
C58 1Bit_Clk_ADC_0.x14.Y 1Bit_Clk_ADC_0.x11.A 0.261475f
C59 1Bit_Clk_ADC_0.x6.B VMID 1.22144f
C60 1Bit_Clk_ADC_0.x5.A CLK 0.067364f
C61 1Bit_Clk_ADC_0.x3.Y 1Bit_Clk_ADC_0.sky130_fd_sc_hd__nand2_4_0.Y 2.9e-19
C62 1Bit_Clk_ADC_0.x11.A a_232625_n27343# 0.003318f
C63 a_196466_n47634# OUT 0.078037f
C64 1Bit_Clk_ADC_0.x9.B a_231021_n27343# 2.87e-19
C65 1Bit_Clk_ADC_0.x3.A a_230965_n27658# 0.001508f
C66 a_230137_n27658# a_230965_n27658# 0.027461f
C67 1Bit_Clk_ADC_0.sky130_fd_sc_hd__nand2_4_0.Y a_232253_n27658# 0.239039f
C68 a_196466_n47634# VREFP 0.012483f
C69 1Bit_Clk_ADC_0.x6.B 1Bit_Clk_ADC_0.x5.A 0.623713f
C70 1Bit_Clk_ADC_0.x3.B 1Bit_Clk_ADC_0.sky130_fd_sc_hd__nand2_4_0.Y 0.266335f
C71 1Bit_Clk_ADC_0.x9.A a_233081_n27658# 0.001566f
C72 1Bit_Clk_ADC_0.x3.Y a_230965_n27658# 0.075819f
C73 a_172166_n12474# a_174650_n12474# 0.314613f
C74 1Bit_Clk_ADC_0.x14.Y 1Bit_Clk_ADC_0.x9.B 0.066398f
C75 1Bit_Clk_ADC_0.x3.A CLK 0.333547f
C76 1Bit_Clk_ADC_0.x14.Y OUT 0.002558f
C77 a_230137_n27658# CLK 0.099582f
C78 OUT VREFN 4.61068f
C79 1Bit_Clk_ADC_0.x4.B VDD 1.40209f
C80 1Bit_Clk_ADC_0.x9.B a_232625_n27343# 0.244651f
C81 a_232625_n27343# OUT 0.248997f
C82 C2S2_Amp_F_I_1.OUT a_173408_n24334# 0.350818f
C83 1Bit_Clk_ADC_0.x3.B a_230965_n27658# 0.202079f
C84 1Bit_Clk_ADC_0.x5.A 1Bit_Clk_ADC_0.x14.Y 7.77e-19
C85 VREFN VREFP 9.41687f
C86 C2S2_Amp_F_I_0.OUT VDD 0.125761p
C87 1Bit_Clk_ADC_0.x3.Y CLK 0.009765f
C88 1Bit_Clk_ADC_0.x6.B 1Bit_Clk_ADC_0.x3.A 0.014137f
C89 1Bit_Clk_ADC_0.x6.B a_230137_n27658# 0.220263f
C90 C2S2_Amp_F_I_1.OUT VMID 0.875751f
C91 1Bit_Clk_ADC_0.x11.A 1Bit_Clk_ADC_0.x9.B 0.076231f
C92 1Bit_Clk_ADC_0.x3.A a_231021_n27343# 0.067928f
C93 a_232253_n27658# CLK 1.15e-19
C94 1Bit_Clk_ADC_0.x14.Y 1Bit_Clk_ADC_0.x9.A 0.23354f
C95 1Bit_Clk_ADC_0.x11.A OUT 0.010009f
C96 1Bit_Clk_ADC_0.x3.B CLK 0.041965f
C97 a_232253_n27658# a_233081_n27658# 0.027461f
C98 1Bit_Clk_ADC_0.x6.B 1Bit_Clk_ADC_0.x3.Y 0.001169f
C99 1Bit_Clk_ADC_0.x9.A a_232625_n27343# 0.074684f
C100 1Bit_Clk_ADC_0.sky130_fd_sc_hd__nand2_4_0.Y VDD 1.13916f
C101 1Bit_Clk_ADC_0.x3.Y a_231021_n27343# 0.193553f
C102 1Bit_Clk_ADC_0.x3.A 1Bit_Clk_ADC_0.x14.Y 0.010804f
C103 1Bit_Clk_ADC_0.x14.Y a_230137_n27658# 0.021134f
C104 C2S2_Amp_F_I_0.VN VDD 5.9774f
C105 a_196466_n45150# VDD 0.067373f
C106 a_230193_n27343# CLK 0.231767f
C107 1Bit_Clk_ADC_0.x6.B 1Bit_Clk_ADC_0.x3.B 0.002721f
C108 C2S2_Amp_F_I_1.OUT a_177926_n43908# 0.001817f
C109 1Bit_Clk_ADC_0.x3.B a_231021_n27343# 0.296644f
C110 1Bit_Clk_ADC_0.x11.A 1Bit_Clk_ADC_0.x9.A 0.444517f
C111 a_230965_n27658# VDD 0.021472f
C112 1Bit_Clk_ADC_0.x14.Y 1Bit_Clk_ADC_0.x3.Y 0.11772f
C113 1Bit_Clk_ADC_0.x9.B OUT 0.737179f
C114 C2S2_Amp_F_I_1.OUT a_175892_n24334# 0.013927f
C115 C2S2_Amp_F_I_1.VN a_166066_n45150# 0.335195f
C116 1Bit_Clk_ADC_0.x6.B a_230193_n27343# 0.030731f
C117 C2S2_Amp_F_I_1.VN C2S2_Amp_F_I_0.VN 0.02f
C118 1Bit_Clk_ADC_0.x14.Y a_232253_n27658# 0.076815f
C119 a_230193_n27343# a_231021_n27343# 0.027461f
C120 1Bit_Clk_ADC_0.x3.A 1Bit_Clk_ADC_0.x11.A 5.71e-20
C121 OUT VREFP 5.91022f
C122 a_173408_n24334# a_175892_n24334# 0.30621f
C123 1Bit_Clk_ADC_0.x3.B 1Bit_Clk_ADC_0.x14.Y 0.374656f
C124 VDD CLK 1.56277f
C125 a_233081_n27658# VDD 0.009152f
C126 1Bit_Clk_ADC_0.x9.B 1Bit_Clk_ADC_0.x9.A 0.155205f
C127 1Bit_Clk_ADC_0.x11.A 1Bit_Clk_ADC_0.x3.Y 0.002138f
C128 1Bit_Clk_ADC_0.x14.Y a_230193_n27343# 0.002875f
C129 1Bit_Clk_ADC_0.x9.A OUT 0.596854f
C130 1Bit_Clk_ADC_0.x6.B a_231797_n27343# 4.38e-20
C131 a_208326_n43908# OUT 0.060961f
C132 1Bit_Clk_ADC_0.x6.B VDD 0.110476p
C133 a_231021_n27343# a_231797_n27343# 0.051797f
C134 1Bit_Clk_ADC_0.x11.A a_232253_n27658# 0.032674f
C135 a_174650_n12474# C2S2_Amp_F_I_0.VN 0.318218f
C136 1Bit_Clk_ADC_0.x4.B 1Bit_Clk_ADC_0.sky130_fd_sc_hd__nand2_4_0.Y 1.28e-19
C137 1Bit_Clk_ADC_0.x3.A 1Bit_Clk_ADC_0.x9.B 1.56e-20
C138 1Bit_Clk_ADC_0.x3.B 1Bit_Clk_ADC_0.x11.A 0.58279f
C139 a_231021_n27343# VDD 0.018306f
C140 a_141908_n24334# C2S2_Amp_F_I_1.VN 9.97e-21
C141 1Bit_Clk_ADC_0.x14.Y a_231797_n27343# 0.229759f
C142 1Bit_Clk_ADC_0.x9.B 1Bit_Clk_ADC_0.x3.Y 6.05e-20
C143 1Bit_Clk_ADC_0.x5.A 1Bit_Clk_ADC_0.x3.A 0.28721f
C144 1Bit_Clk_ADC_0.x5.A a_230137_n27658# 0.001508f
C145 C2S2_Amp_F_I_0.OUT C2S2_Amp_F_I_0.VN 0.285903p
C146 1Bit_Clk_ADC_0.x14.Y VDD 2.76658f
C147 a_231797_n27343# a_232625_n27343# 0.027461f
C148 1Bit_Clk_ADC_0.x4.B a_230965_n27658# 0.213809f
C149 VDD VREFN 1.49715f
C150 1Bit_DAC_Inv_0.OUT VREFN 22.8759f
C151 a_232625_n27343# VDD 0.010259f
C152 1Bit_Clk_ADC_0.x9.B a_232253_n27658# 0.009429f
C153 1Bit_Clk_ADC_0.x5.A 1Bit_Clk_ADC_0.x3.Y 2.39e-20
C154 1Bit_Clk_ADC_0.x3.B 1Bit_Clk_ADC_0.x9.B 0.001361f
C155 1Bit_Clk_ADC_0.x3.A 1Bit_Clk_ADC_0.x9.A 0.004063f
C156 1Bit_Clk_ADC_0.x3.B OUT 8.88e-20
C157 1Bit_DAC_0.OUT VREFN 22.9102f
C158 1Bit_Clk_ADC_0.x4.B CLK 0.419006f
C159 1Bit_Clk_ADC_0.x11.A a_231797_n27343# 0.11656f
C160 a_208326_n46392# OUT 0.731511f
C161 1Bit_Clk_ADC_0.x9.A 1Bit_Clk_ADC_0.x3.Y 0.003053f
C162 1Bit_Clk_ADC_0.x5.A 1Bit_Clk_ADC_0.x3.B 2.89e-19
C163 C2S2_Amp_F_I_1.OUT VDD 38.5169f
C164 1Bit_Clk_ADC_0.x11.A VDD 0.742348f
C165 C2S2_Amp_F_I_0.VN a_196466_n45150# 0.359531f
C166 1Bit_Clk_ADC_0.sky130_fd_sc_hd__nand2_4_0.Y a_230965_n27658# 2.43e-19
C167 a_144392_n24334# C2S2_Amp_F_I_1.VN 1.80416f
C168 a_177926_n43908# a_177926_n46392# 0.329456f
C169 1Bit_Clk_ADC_0.x6.B 1Bit_Clk_ADC_0.x4.B 0.206519f
C170 1Bit_Clk_ADC_0.x3.A 1Bit_Clk_ADC_0.x3.Y 0.300624f
C171 1Bit_Clk_ADC_0.x5.A a_230193_n27343# 0.079345f
C172 1Bit_Clk_ADC_0.x3.B 1Bit_Clk_ADC_0.x9.A 0.002027f
C173 a_231021_n27343# 1Bit_Clk_ADC_0.x4.B 0.001491f
C174 C2S2_Amp_F_I_0.OUT 1Bit_Clk_ADC_0.x6.B 2.82451f
C175 C2S2_Amp_F_I_1.OUT C2S2_Amp_F_I_1.VN 0.28569p
C176 1Bit_Clk_ADC_0.x9.B a_231797_n27343# 0.006032f
C177 VDD VMID 59.9898f
C178 a_231797_n27343# OUT 9.05e-19
C179 a_208326_n43908# a_208326_n46392# 0.30621f
C180 a_172166_n12474# VMID 0.078261f
C181 1Bit_Clk_ADC_0.sky130_fd_sc_hd__nand2_4_0.Y a_233081_n27658# 0.265834f
C182 1Bit_Clk_ADC_0.x3.A 1Bit_Clk_ADC_0.x3.B 0.058791f
C183 1Bit_Clk_ADC_0.x9.B VDD 1.24414f
C184 1Bit_Clk_ADC_0.x3.B a_230137_n27658# 0.001359f
C185 VDD OUT 17.945599f
C186 a_166066_n45150# a_166066_n47634# 0.300332f
C187 1Bit_Clk_ADC_0.x14.Y 1Bit_Clk_ADC_0.x4.B 0.094667f
C188 1Bit_DAC_Inv_0.OUT OUT 4.77363f
C189 VDD VREFP 1.87743f
C190 1Bit_Clk_ADC_0.x3.A a_230193_n27343# 0.186379f
C191 1Bit_Clk_ADC_0.x3.B 1Bit_Clk_ADC_0.x3.Y 1.03376f
C192 1Bit_Clk_ADC_0.x5.A VDD 0.73774f
C193 a_230965_n27658# CLK 0.007075f
C194 1Bit_DAC_0.OUT OUT 5.80476f
C195 1Bit_DAC_Inv_0.OUT VREFP 22.275301f
C196 a_140666_n12474# a_143150_n12474# 0.314613f
C197 C2S2_Amp_F_I_1.VN VMID 0.128417f
C198 a_196466_n45150# a_196466_n47634# 0.314613f
C199 1Bit_Clk_ADC_0.x9.A a_231797_n27343# 0.179363f
C200 a_177926_n43908# VDD 0.098147f
C201 1Bit_Clk_ADC_0.x3.B a_232253_n27658# 0.211683f
C202 1Bit_DAC_0.OUT VREFP 22.617401f
C203 1Bit_Clk_ADC_0.x3.Y a_230193_n27343# 3.83e-19
C204 VREFP GND 95.88653f
C205 VREFN GND 81.199844f
C206 OUT GND 0.103449p
C207 CLK GND 4.14803f
C208 VMID GND 0.111856p
C209 SIG GND 2.67679f
C210 VDD GND 0.707463p
C211 a_233081_n27658# GND 0.520902f
C212 a_232253_n27658# GND 0.52311f
C213 a_230965_n27658# GND 0.522503f
C214 a_230137_n27658# GND 0.533106f
C215 1Bit_Clk_ADC_0.sky130_fd_sc_hd__nand2_4_0.Y GND 0.690821f
C216 1Bit_Clk_ADC_0.x4.B GND 0.544647f
C217 1Bit_DAC_0.OUT GND 19.42917f
C218 a_196466_n47634# GND 3.749f
C219 a_208326_n46392# GND 3.11889f
C220 a_196466_n45150# GND 3.1032f
C221 a_208326_n43908# GND 3.13839f
C222 1Bit_DAC_Inv_0.OUT GND 16.557985f
C223 a_166066_n47634# GND 3.49882f
C224 a_177926_n46392# GND 3.44174f
C225 a_166066_n45150# GND 3.13081f
C226 a_177926_n43908# GND 3.29573f
C227 a_232625_n27343# GND 0.524587f
C228 a_231797_n27343# GND 0.501639f
C229 a_231021_n27343# GND 0.491501f
C230 a_230193_n27343# GND 0.52031f
C231 1Bit_Clk_ADC_0.x3.Y GND 0.615402f
C232 1Bit_Clk_ADC_0.x9.A GND 0.507131f
C233 1Bit_Clk_ADC_0.x9.B GND 1.014f
C234 1Bit_Clk_ADC_0.x11.A GND 0.961749f
C235 1Bit_Clk_ADC_0.x14.Y GND 2.370527f
C236 1Bit_Clk_ADC_0.x3.B GND 1.893877f
C237 1Bit_Clk_ADC_0.x3.A GND 0.484392f
C238 1Bit_Clk_ADC_0.x5.A GND 0.691117f
C239 1Bit_Clk_ADC_0.x6.B GND 41.9156f
C240 C2S2_Amp_F_I_0.VN GND 73.48906f
C241 a_175892_n24334# GND 3.5131f
C242 a_174650_n12474# GND 2.9871f
C243 a_173408_n24334# GND 3.29615f
C244 a_172166_n12474# GND 3.27394f
C245 C2S2_Amp_F_I_0.OUT GND 0.127025p
C246 C2S2_Amp_F_I_1.VN GND 69.36782f
C247 a_144392_n24334# GND 3.5131f
C248 a_143150_n12474# GND 2.9871f
C249 a_141908_n24334# GND 3.29148f
C250 a_140666_n12474# GND 3.27394f
C251 C2S2_Amp_F_I_1.OUT GND 0.117888p
C252 C2S2_Amp_F_I_1.VN.t1 GND 0.867778f
C253 C2S2_Amp_F_I_1.VN.t12 GND 19.0241f
C254 C2S2_Amp_F_I_1.VN.t15 GND 9.81608f
C255 C2S2_Amp_F_I_1.VN.n1 GND 9.502151f
C256 C2S2_Amp_F_I_1.VN.t4 GND 9.81608f
C257 C2S2_Amp_F_I_1.VN.n2 GND 9.375669f
C258 C2S2_Amp_F_I_1.VN.t16 GND 9.81608f
C259 C2S2_Amp_F_I_1.VN.n3 GND 10.2173f
C260 C2S2_Amp_F_I_1.VN.t5 GND 19.0241f
C261 C2S2_Amp_F_I_1.VN.t8 GND 9.81608f
C262 C2S2_Amp_F_I_1.VN.n4 GND 9.502151f
C263 C2S2_Amp_F_I_1.VN.t20 GND 9.81608f
C264 C2S2_Amp_F_I_1.VN.n5 GND 9.375669f
C265 C2S2_Amp_F_I_1.VN.t11 GND 9.81608f
C266 C2S2_Amp_F_I_1.VN.n6 GND 9.34184f
C267 C2S2_Amp_F_I_1.VN.n7 GND 2.29622f
C268 C2S2_Amp_F_I_1.VN.t3 GND 19.0241f
C269 C2S2_Amp_F_I_1.VN.t7 GND 9.81608f
C270 C2S2_Amp_F_I_1.VN.n8 GND 9.502151f
C271 C2S2_Amp_F_I_1.VN.t18 GND 9.81608f
C272 C2S2_Amp_F_I_1.VN.n9 GND 9.375669f
C273 C2S2_Amp_F_I_1.VN.t9 GND 9.81608f
C274 C2S2_Amp_F_I_1.VN.n10 GND 9.34184f
C275 C2S2_Amp_F_I_1.VN.n11 GND 1.6247f
C276 C2S2_Amp_F_I_1.VN.t0 GND 0.643635f
C277 C2S2_Amp_F_I_1.VN.n12 GND 15.079299f
C278 C2S2_Amp_F_I_1.VN.n13 GND 19.528198f
C279 C2S2_Amp_F_I_1.VN.n14 GND 0.046866f
C280 C2S2_Amp_F_I_1.VN.n15 GND 0.030462f
C281 C2S2_Amp_F_I_1.VN.n16 GND 0.030462f
C282 C2S2_Amp_F_I_1.VN.t2 GND 0.078658f
C283 C2S2_Amp_F_I_1.VN.n17 GND 0.03642f
C284 C2S2_Amp_F_I_1.VN.n18 GND 0.096176f
C285 C2S2_Amp_F_I_1.VN.t13 GND 0.078658f
C286 C2S2_Amp_F_I_1.VN.n19 GND 0.096176f
C287 C2S2_Amp_F_I_1.VN.t17 GND 0.078658f
C288 C2S2_Amp_F_I_1.VN.n20 GND 0.030462f
C289 C2S2_Amp_F_I_1.VN.n21 GND 0.030462f
C290 C2S2_Amp_F_I_1.VN.t10 GND 0.078658f
C291 C2S2_Amp_F_I_1.VN.n22 GND 0.030462f
C292 C2S2_Amp_F_I_1.VN.t14 GND 0.078658f
C293 C2S2_Amp_F_I_1.VN.n23 GND 0.030462f
C294 C2S2_Amp_F_I_1.VN.n24 GND 0.030462f
C295 C2S2_Amp_F_I_1.VN.t19 GND 0.078658f
C296 C2S2_Amp_F_I_1.VN.n25 GND 0.030462f
C297 C2S2_Amp_F_I_1.VN.t6 GND 0.078658f
C298 C2S2_Amp_F_I_1.VN.n26 GND 0.046866f
C299 C2S2_Amp_F_I_1.VN.n27 GND 1.01293f
C300 C2S2_Amp_F_I_1.VN.n28 GND 8.537971f
C301 C2S2_Amp_F_I_1.VN.n29 GND 5.25466f
C302 C2S2_Amp_F_I_1.VN.n30 GND 1.84532f
C303 a_182797_n11365.t7 GND 0.517854f
C304 a_182797_n11365.t6 GND 0.52009f
C305 a_182797_n11365.n0 GND 6.03626f
C306 a_182797_n11365.t4 GND 20.8342f
C307 a_182797_n11365.n1 GND 7.27757f
C308 a_182797_n11365.t5 GND 20.8342f
C309 a_182797_n11365.n2 GND 4.66798f
C310 a_182797_n11365.t3 GND 20.8342f
C311 a_182797_n11365.n3 GND 4.66798f
C312 a_182797_n11365.t2 GND 20.8342f
C313 a_182797_n11365.n4 GND 7.29735f
C314 a_182797_n11365.t1 GND 0.519976f
C315 a_182797_n11365.n5 GND 6.0404f
C316 a_182797_n11365.t0 GND 0.517749f
C317 a_186826_n27776.t8 GND 0.194162f
C318 a_186826_n27776.t9 GND 0.10698f
C319 a_186826_n27776.n0 GND 1.28057f
C320 a_186826_n27776.n1 GND 0.194927f
C321 a_186826_n27776.t5 GND 0.009165f
C322 a_186826_n27776.t6 GND 0.009165f
C323 a_186826_n27776.n2 GND 0.032429f
C324 a_186826_n27776.t4 GND 0.009165f
C325 a_186826_n27776.t3 GND 0.009165f
C326 a_186826_n27776.n3 GND 0.032429f
C327 a_186826_n27776.n4 GND 0.095668f
C328 a_186826_n27776.t2 GND 0.009165f
C329 a_186826_n27776.t7 GND 0.009165f
C330 a_186826_n27776.n5 GND 0.038664f
C331 a_186826_n27776.n6 GND 0.110693f
C332 a_186826_n27776.n7 GND 0.095728f
C333 a_186826_n27776.n8 GND 0.200489f
C334 a_186826_n27776.t1 GND 0.10698f
C335 a_186826_n27776.n9 GND 1.51993f
C336 a_186826_n27776.t0 GND 0.235357f
C337 a_150997_n11365.t2 GND 17.2646f
C338 a_150997_n11365.t5 GND 17.2646f
C339 a_150997_n11365.t4 GND 17.2646f
C340 a_150997_n11365.t3 GND 17.2646f
C341 a_150997_n11365.t7 GND 0.429041f
C342 a_150997_n11365.t6 GND 0.430886f
C343 a_150997_n11365.n0 GND 5.00548f
C344 a_150997_n11365.n1 GND 6.04706f
C345 a_150997_n11365.n2 GND 3.86819f
C346 a_150997_n11365.n3 GND 3.86819f
C347 a_150997_n11365.n4 GND 6.03068f
C348 a_150997_n11365.t1 GND 0.43098f
C349 a_150997_n11365.n5 GND 5.00197f
C350 a_150997_n11365.t0 GND 0.429193f
C351 VMID.n0 GND 0.028568f
C352 VMID.n1 GND 0.018576f
C353 VMID.n2 GND 0.018576f
C354 VMID.t5 GND 0.047968f
C355 VMID.n3 GND 0.022176f
C356 VMID.n4 GND 0.058729f
C357 VMID.t3 GND 0.047968f
C358 VMID.n5 GND 0.058729f
C359 VMID.t19 GND 0.047968f
C360 VMID.n6 GND 0.018576f
C361 VMID.n7 GND 0.018576f
C362 VMID.t4 GND 0.047968f
C363 VMID.n8 GND 0.018576f
C364 VMID.t14 GND 0.047968f
C365 VMID.n9 GND 0.018576f
C366 VMID.n10 GND 0.018576f
C367 VMID.t12 GND 0.047968f
C368 VMID.n11 GND 0.018576f
C369 VMID.t10 GND 0.047968f
C370 VMID.n12 GND 0.028568f
C371 VMID.n13 GND 0.394163f
C372 VMID.n14 GND 13.1926f
C373 VMID.n15 GND 0.028568f
C374 VMID.n16 GND 0.018576f
C375 VMID.n17 GND 0.018576f
C376 VMID.t17 GND 0.047968f
C377 VMID.n18 GND 0.022176f
C378 VMID.n19 GND 0.058729f
C379 VMID.t9 GND 0.047968f
C380 VMID.n20 GND 0.058729f
C381 VMID.t6 GND 0.047968f
C382 VMID.n21 GND 0.018576f
C383 VMID.n22 GND 0.018576f
C384 VMID.t0 GND 0.047968f
C385 VMID.n23 GND 0.018576f
C386 VMID.t20 GND 0.047968f
C387 VMID.n24 GND 0.018576f
C388 VMID.n25 GND 0.018576f
C389 VMID.t15 GND 0.047968f
C390 VMID.n26 GND 0.018576f
C391 VMID.t7 GND 0.047968f
C392 VMID.n27 GND 0.028568f
C393 VMID.n28 GND 0.705685f
C394 VMID.n29 GND 18.6742f
C395 VMID.n30 GND 0.028568f
C396 VMID.n31 GND 0.018576f
C397 VMID.n32 GND 0.018576f
C398 VMID.t11 GND 0.047968f
C399 VMID.n33 GND 0.022176f
C400 VMID.n34 GND 0.058729f
C401 VMID.t2 GND 0.047968f
C402 VMID.n35 GND 0.058729f
C403 VMID.t18 GND 0.047968f
C404 VMID.n36 GND 0.018576f
C405 VMID.n37 GND 0.018576f
C406 VMID.t13 GND 0.047968f
C407 VMID.n38 GND 0.018576f
C408 VMID.t1 GND 0.047968f
C409 VMID.n39 GND 0.018576f
C410 VMID.n40 GND 0.018576f
C411 VMID.t16 GND 0.047968f
C412 VMID.n41 GND 0.018576f
C413 VMID.t8 GND 0.047968f
C414 VMID.n42 GND 0.028568f
C415 VMID.n43 GND 0.705685f
C416 VMID.n44 GND 14.344799f
C417 C2S2_Amp_F_I_0.VN.t0 GND 1.19074f
C418 C2S2_Amp_F_I_0.VN.t11 GND 19.5456f
C419 C2S2_Amp_F_I_0.VN.t13 GND 10.0852f
C420 C2S2_Amp_F_I_0.VN.n0 GND 9.76265f
C421 C2S2_Amp_F_I_0.VN.t6 GND 10.0852f
C422 C2S2_Amp_F_I_0.VN.n1 GND 9.6327f
C423 C2S2_Amp_F_I_0.VN.t18 GND 10.0852f
C424 C2S2_Amp_F_I_0.VN.n2 GND 10.8794f
C425 C2S2_Amp_F_I_0.VN.t12 GND 19.5456f
C426 C2S2_Amp_F_I_0.VN.t15 GND 10.0852f
C427 C2S2_Amp_F_I_0.VN.n3 GND 9.76265f
C428 C2S2_Amp_F_I_0.VN.t7 GND 10.0852f
C429 C2S2_Amp_F_I_0.VN.n4 GND 9.6327f
C430 C2S2_Amp_F_I_0.VN.t20 GND 10.0852f
C431 C2S2_Amp_F_I_0.VN.n5 GND 9.59858f
C432 C2S2_Amp_F_I_0.VN.n6 GND 2.55186f
C433 C2S2_Amp_F_I_0.VN.t17 GND 19.5456f
C434 C2S2_Amp_F_I_0.VN.t19 GND 10.0852f
C435 C2S2_Amp_F_I_0.VN.n7 GND 9.76265f
C436 C2S2_Amp_F_I_0.VN.t8 GND 10.0852f
C437 C2S2_Amp_F_I_0.VN.n8 GND 9.6327f
C438 C2S2_Amp_F_I_0.VN.t3 GND 10.0852f
C439 C2S2_Amp_F_I_0.VN.n9 GND 9.59858f
C440 C2S2_Amp_F_I_0.VN.n10 GND 1.6291f
C441 C2S2_Amp_F_I_0.VN.t1 GND 0.661361f
C442 C2S2_Amp_F_I_0.VN.n11 GND 15.965099f
C443 C2S2_Amp_F_I_0.VN.n12 GND 0.048151f
C444 C2S2_Amp_F_I_0.VN.n13 GND 0.031297f
C445 C2S2_Amp_F_I_0.VN.n14 GND 0.031297f
C446 C2S2_Amp_F_I_0.VN.t4 GND 0.080815f
C447 C2S2_Amp_F_I_0.VN.n15 GND 0.037418f
C448 C2S2_Amp_F_I_0.VN.n16 GND 0.098813f
C449 C2S2_Amp_F_I_0.VN.t9 GND 0.080815f
C450 C2S2_Amp_F_I_0.VN.n17 GND 0.098813f
C451 C2S2_Amp_F_I_0.VN.t14 GND 0.080815f
C452 C2S2_Amp_F_I_0.VN.n18 GND 0.031297f
C453 C2S2_Amp_F_I_0.VN.n19 GND 0.031297f
C454 C2S2_Amp_F_I_0.VN.t16 GND 0.080815f
C455 C2S2_Amp_F_I_0.VN.n20 GND 0.031297f
C456 C2S2_Amp_F_I_0.VN.t2 GND 0.080815f
C457 C2S2_Amp_F_I_0.VN.n21 GND 0.031297f
C458 C2S2_Amp_F_I_0.VN.n22 GND 0.031297f
C459 C2S2_Amp_F_I_0.VN.t5 GND 0.080815f
C460 C2S2_Amp_F_I_0.VN.n23 GND 0.031297f
C461 C2S2_Amp_F_I_0.VN.t10 GND 0.080815f
C462 C2S2_Amp_F_I_0.VN.n24 GND 0.048151f
C463 C2S2_Amp_F_I_0.VN.n25 GND 0.975434f
C464 C2S2_Amp_F_I_0.VN.n26 GND 28.0714f
C465 C2S2_Amp_F_I_0.VN.n27 GND 7.58772f
C466 a_185229_n11365.n0 GND 0.150606f
C467 a_185229_n11365.n1 GND 0.104449f
C468 a_185229_n11365.n2 GND 0.104449f
C469 a_185229_n11365.n3 GND 0.103718f
C470 a_185229_n11365.n4 GND 0.104449f
C471 a_185229_n11365.t50 GND 0.269595f
C472 a_185229_n11365.n5 GND 0.103768f
C473 a_185229_n11365.n6 GND 0.033198f
C474 a_185229_n11365.n7 GND 0.010247f
C475 a_185229_n11365.n8 GND 0.195697f
C476 a_185229_n11365.n9 GND 0.004124f
C477 a_185229_n11365.n10 GND 0.003895f
C478 a_185229_n11365.n11 GND 0.01329f
C479 a_185229_n11365.n12 GND 0.004124f
C480 a_185229_n11365.n13 GND 0.011088f
C481 a_185229_n11365.n14 GND 0.003895f
C482 a_185229_n11365.n15 GND 0.014674f
C483 a_185229_n11365.n16 GND 0.023503f
C484 a_185229_n11365.n17 GND 0.004124f
C485 a_185229_n11365.n18 GND 0.003895f
C486 a_185229_n11365.n19 GND 0.010936f
C487 a_185229_n11365.n20 GND 0.01116f
C488 a_185229_n11365.n21 GND 0.003895f
C489 a_185229_n11365.n22 GND 0.003895f
C490 a_185229_n11365.n23 GND 0.004124f
C491 a_185229_n11365.n24 GND 0.01329f
C492 a_185229_n11365.n25 GND 0.01329f
C493 a_185229_n11365.t1 GND 0.019076f
C494 a_185229_n11365.n26 GND 0.031577f
C495 a_185229_n11365.n27 GND 0.004835f
C496 a_185229_n11365.n28 GND 0.009967f
C497 a_185229_n11365.n29 GND 0.01329f
C498 a_185229_n11365.n30 GND 0.004124f
C499 a_185229_n11365.n31 GND 0.003895f
C500 a_185229_n11365.n32 GND 0.01113f
C501 a_185229_n11365.n33 GND 0.020747f
C502 a_185229_n11365.n34 GND 2.57091f
C503 a_185229_n11365.n35 GND 0.033198f
C504 a_185229_n11365.n36 GND 0.033198f
C505 a_185229_n11365.n37 GND 0.033198f
C506 a_185229_n11365.n38 GND 0.010247f
C507 a_185229_n11365.t24 GND 0.04886f
C508 a_185229_n11365.t31 GND 0.04886f
C509 a_185229_n11365.n39 GND 0.104474f
C510 a_185229_n11365.n40 GND 0.004124f
C511 a_185229_n11365.n41 GND 0.011088f
C512 a_185229_n11365.n42 GND 0.006907f
C513 a_185229_n11365.n43 GND 0.003895f
C514 a_185229_n11365.n44 GND 0.004124f
C515 a_185229_n11365.n45 GND 0.003895f
C516 a_185229_n11365.n46 GND 0.010936f
C517 a_185229_n11365.n47 GND 0.01116f
C518 a_185229_n11365.n48 GND 0.003895f
C519 a_185229_n11365.n49 GND 0.004124f
C520 a_185229_n11365.n50 GND 0.009096f
C521 a_185229_n11365.n51 GND 0.007118f
C522 a_185229_n11365.n52 GND 0.178986f
C523 a_185229_n11365.n53 GND 0.427503f
C524 a_185229_n11365.n54 GND 0.010247f
C525 a_185229_n11365.t26 GND 0.04886f
C526 a_185229_n11365.t0 GND 0.04886f
C527 a_185229_n11365.n55 GND 0.104474f
C528 a_185229_n11365.n56 GND 0.004124f
C529 a_185229_n11365.n57 GND 0.011088f
C530 a_185229_n11365.n58 GND 0.006907f
C531 a_185229_n11365.n59 GND 0.003895f
C532 a_185229_n11365.n60 GND 0.004124f
C533 a_185229_n11365.n61 GND 0.003895f
C534 a_185229_n11365.n62 GND 0.010936f
C535 a_185229_n11365.n63 GND 0.01116f
C536 a_185229_n11365.n64 GND 0.003895f
C537 a_185229_n11365.n65 GND 0.004124f
C538 a_185229_n11365.n66 GND 0.009096f
C539 a_185229_n11365.n67 GND 0.007118f
C540 a_185229_n11365.n68 GND 0.178986f
C541 a_185229_n11365.n69 GND 0.427503f
C542 a_185229_n11365.n70 GND 0.010247f
C543 a_185229_n11365.t27 GND 0.04886f
C544 a_185229_n11365.t28 GND 0.04886f
C545 a_185229_n11365.n71 GND 0.104474f
C546 a_185229_n11365.n72 GND 0.004124f
C547 a_185229_n11365.n73 GND 0.011088f
C548 a_185229_n11365.n74 GND 0.006907f
C549 a_185229_n11365.n75 GND 0.003895f
C550 a_185229_n11365.n76 GND 0.004124f
C551 a_185229_n11365.n77 GND 0.003895f
C552 a_185229_n11365.n78 GND 0.010936f
C553 a_185229_n11365.n79 GND 0.01116f
C554 a_185229_n11365.n80 GND 0.003895f
C555 a_185229_n11365.n81 GND 0.004124f
C556 a_185229_n11365.n82 GND 0.009096f
C557 a_185229_n11365.n83 GND 0.007118f
C558 a_185229_n11365.n84 GND 0.178986f
C559 a_185229_n11365.n85 GND 2.76314f
C560 a_185229_n11365.n86 GND 0.103175f
C561 a_185229_n11365.n87 GND 0.103465f
C562 a_185229_n11365.n88 GND 0.104449f
C563 a_185229_n11365.n89 GND 0.104449f
C564 a_185229_n11365.n90 GND 0.150771f
C565 a_185229_n11365.t30 GND 0.932339f
C566 a_185229_n11365.t29 GND 0.833027f
C567 a_185229_n11365.n91 GND 9.08508f
C568 a_185229_n11365.n92 GND 0.609697f
C569 a_185229_n11365.t56 GND 0.269595f
C570 a_185229_n11365.n93 GND 0.154543f
C571 a_185229_n11365.n94 GND 0.104449f
C572 a_185229_n11365.t59 GND 0.269595f
C573 a_185229_n11365.n95 GND 0.104449f
C574 a_185229_n11365.t66 GND 0.269595f
C575 a_185229_n11365.n96 GND 0.104449f
C576 a_185229_n11365.n97 GND 0.104449f
C577 a_185229_n11365.t70 GND 0.269595f
C578 a_185229_n11365.n98 GND 0.104449f
C579 a_185229_n11365.t51 GND 0.269595f
C580 a_185229_n11365.n99 GND 0.104449f
C581 a_185229_n11365.n100 GND 0.104449f
C582 a_185229_n11365.t55 GND 0.269595f
C583 a_185229_n11365.n101 GND 0.104449f
C584 a_185229_n11365.t43 GND 0.269595f
C585 a_185229_n11365.n102 GND 0.104449f
C586 a_185229_n11365.n103 GND 0.104449f
C587 a_185229_n11365.n104 GND 0.104449f
C588 a_185229_n11365.n105 GND 0.104449f
C589 a_185229_n11365.n106 GND 0.104449f
C590 a_185229_n11365.n107 GND 0.104449f
C591 a_185229_n11365.n108 GND 0.104449f
C592 a_185229_n11365.n109 GND 0.104449f
C593 a_185229_n11365.n110 GND 0.104449f
C594 a_185229_n11365.n111 GND 0.104449f
C595 a_185229_n11365.n112 GND 0.104449f
C596 a_185229_n11365.n113 GND 0.104449f
C597 a_185229_n11365.t60 GND 0.269595f
C598 a_185229_n11365.n114 GND 0.104449f
C599 a_185229_n11365.n115 GND 0.104449f
C600 a_185229_n11365.t52 GND 0.269595f
C601 a_185229_n11365.n116 GND 0.104449f
C602 a_185229_n11365.t33 GND 0.269595f
C603 a_185229_n11365.n117 GND 0.104449f
C604 a_185229_n11365.n118 GND 0.104449f
C605 a_185229_n11365.t69 GND 0.269595f
C606 a_185229_n11365.n119 GND 0.104449f
C607 a_185229_n11365.t63 GND 0.269595f
C608 a_185229_n11365.n120 GND 0.104449f
C609 a_185229_n11365.n121 GND 0.104449f
C610 a_185229_n11365.t58 GND 0.269595f
C611 a_185229_n11365.n122 GND 0.104449f
C612 a_185229_n11365.t65 GND 0.269595f
C613 a_185229_n11365.n123 GND 0.104449f
C614 a_185229_n11365.n124 GND 0.104449f
C615 a_185229_n11365.t48 GND 0.269595f
C616 a_185229_n11365.n125 GND 0.104449f
C617 a_185229_n11365.t41 GND 0.269595f
C618 a_185229_n11365.n126 GND 0.104449f
C619 a_185229_n11365.n127 GND 0.104449f
C620 a_185229_n11365.t35 GND 0.269595f
C621 a_185229_n11365.n128 GND 0.104449f
C622 a_185229_n11365.t71 GND 0.269595f
C623 a_185229_n11365.n129 GND 0.104449f
C624 a_185229_n11365.n130 GND 0.104449f
C625 a_185229_n11365.t67 GND 0.269595f
C626 a_185229_n11365.n131 GND 0.104449f
C627 a_185229_n11365.t44 GND 0.269595f
C628 a_185229_n11365.n132 GND 0.104449f
C629 a_185229_n11365.n133 GND 0.104449f
C630 a_185229_n11365.t36 GND 0.269595f
C631 a_185229_n11365.n134 GND 0.104449f
C632 a_185229_n11365.t32 GND 0.269595f
C633 a_185229_n11365.n135 GND 0.104449f
C634 a_185229_n11365.n136 GND 0.104449f
C635 a_185229_n11365.t68 GND 0.269595f
C636 a_185229_n11365.n137 GND 0.104449f
C637 a_185229_n11365.t62 GND 0.269595f
C638 a_185229_n11365.n138 GND 0.104449f
C639 a_185229_n11365.n139 GND 0.104449f
C640 a_185229_n11365.t42 GND 0.269595f
C641 a_185229_n11365.n140 GND 0.104449f
C642 a_185229_n11365.t38 GND 0.269595f
C643 a_185229_n11365.n141 GND 0.104449f
C644 a_185229_n11365.n142 GND 0.104449f
C645 a_185229_n11365.t47 GND 0.269595f
C646 a_185229_n11365.n143 GND 0.104449f
C647 a_185229_n11365.t40 GND 0.269595f
C648 a_185229_n11365.n144 GND 0.104449f
C649 a_185229_n11365.n145 GND 0.104449f
C650 a_185229_n11365.t34 GND 0.269595f
C651 a_185229_n11365.n146 GND 0.104449f
C652 a_185229_n11365.t57 GND 0.269595f
C653 a_185229_n11365.n147 GND 0.104449f
C654 a_185229_n11365.n148 GND 0.104449f
C655 a_185229_n11365.t53 GND 0.269595f
C656 a_185229_n11365.n149 GND 0.107487f
C657 a_185229_n11365.n150 GND 0.110891f
C658 a_185229_n11365.n151 GND 1.82882f
C659 a_185229_n11365.n152 GND 0.02041f
C660 a_185229_n11365.n153 GND 0.011088f
C661 a_185229_n11365.n154 GND 0.003895f
C662 a_185229_n11365.n155 GND 0.01329f
C663 a_185229_n11365.n156 GND 0.004124f
C664 a_185229_n11365.n157 GND 0.003895f
C665 a_185229_n11365.n158 GND 0.01329f
C666 a_185229_n11365.n159 GND 0.004124f
C667 a_185229_n11365.n160 GND 0.032372f
C668 a_185229_n11365.t9 GND 0.024889f
C669 a_185229_n11365.n161 GND 0.009967f
C670 a_185229_n11365.n162 GND 0.005094f
C671 a_185229_n11365.n163 GND 0.003895f
C672 a_185229_n11365.n164 GND 0.189103f
C673 a_185229_n11365.n165 GND 0.010921f
C674 a_185229_n11365.n166 GND 0.011123f
C675 a_185229_n11365.n167 GND 0.003895f
C676 a_185229_n11365.n168 GND 0.004124f
C677 a_185229_n11365.n169 GND 0.01329f
C678 a_185229_n11365.n170 GND 0.01329f
C679 a_185229_n11365.n171 GND 0.004124f
C680 a_185229_n11365.n172 GND 0.003895f
C681 a_185229_n11365.n173 GND 0.010557f
C682 a_185229_n11365.n174 GND 0.010936f
C683 a_185229_n11365.n175 GND 0.003895f
C684 a_185229_n11365.n176 GND 0.004124f
C685 a_185229_n11365.n177 GND 0.026181f
C686 a_185229_n11365.n178 GND 0.011997f
C687 a_185229_n11365.n179 GND 0.033198f
C688 a_185229_n11365.n180 GND 0.621914f
C689 a_185229_n11365.n181 GND 0.200066f
C690 a_185229_n11365.n182 GND 0.011088f
C691 a_185229_n11365.n183 GND 0.003895f
C692 a_185229_n11365.t6 GND 0.04886f
C693 a_185229_n11365.n184 GND 0.004124f
C694 a_185229_n11365.n185 GND 0.004124f
C695 a_185229_n11365.n186 GND 0.003895f
C696 a_185229_n11365.n187 GND 0.010936f
C697 a_185229_n11365.n188 GND 0.010557f
C698 a_185229_n11365.n189 GND 0.009005f
C699 a_185229_n11365.n190 GND 0.008838f
C700 a_185229_n11365.t13 GND 0.04886f
C701 a_185229_n11365.n191 GND 0.100636f
C702 a_185229_n11365.n192 GND 0.006907f
C703 a_185229_n11365.n193 GND 0.033198f
C704 a_185229_n11365.n194 GND 0.342588f
C705 a_185229_n11365.n195 GND 0.200066f
C706 a_185229_n11365.n196 GND 0.011088f
C707 a_185229_n11365.n197 GND 0.003895f
C708 a_185229_n11365.t12 GND 0.04886f
C709 a_185229_n11365.n198 GND 0.004124f
C710 a_185229_n11365.n199 GND 0.004124f
C711 a_185229_n11365.n200 GND 0.003895f
C712 a_185229_n11365.n201 GND 0.010936f
C713 a_185229_n11365.n202 GND 0.010557f
C714 a_185229_n11365.n203 GND 0.009005f
C715 a_185229_n11365.n204 GND 0.008838f
C716 a_185229_n11365.t4 GND 0.04886f
C717 a_185229_n11365.n205 GND 0.100636f
C718 a_185229_n11365.n206 GND 0.006907f
C719 a_185229_n11365.n207 GND 0.033198f
C720 a_185229_n11365.n208 GND 0.347642f
C721 a_185229_n11365.n209 GND 0.200066f
C722 a_185229_n11365.n210 GND 0.011088f
C723 a_185229_n11365.n211 GND 0.003895f
C724 a_185229_n11365.t19 GND 0.04886f
C725 a_185229_n11365.n212 GND 0.004124f
C726 a_185229_n11365.n213 GND 0.004124f
C727 a_185229_n11365.n214 GND 0.003895f
C728 a_185229_n11365.n215 GND 0.010936f
C729 a_185229_n11365.n216 GND 0.010557f
C730 a_185229_n11365.n217 GND 0.009005f
C731 a_185229_n11365.n218 GND 0.008838f
C732 a_185229_n11365.t16 GND 0.04886f
C733 a_185229_n11365.n219 GND 0.100636f
C734 a_185229_n11365.n220 GND 0.006907f
C735 a_185229_n11365.n221 GND 0.033198f
C736 a_185229_n11365.n222 GND 0.342588f
C737 a_185229_n11365.n223 GND 0.200066f
C738 a_185229_n11365.n224 GND 0.011088f
C739 a_185229_n11365.n225 GND 0.003895f
C740 a_185229_n11365.t11 GND 0.04886f
C741 a_185229_n11365.n226 GND 0.004124f
C742 a_185229_n11365.n227 GND 0.004124f
C743 a_185229_n11365.n228 GND 0.003895f
C744 a_185229_n11365.n229 GND 0.010936f
C745 a_185229_n11365.n230 GND 0.010557f
C746 a_185229_n11365.n231 GND 0.009005f
C747 a_185229_n11365.n232 GND 0.008838f
C748 a_185229_n11365.t7 GND 0.04886f
C749 a_185229_n11365.n233 GND 0.100636f
C750 a_185229_n11365.n234 GND 0.006907f
C751 a_185229_n11365.n235 GND 0.033198f
C752 a_185229_n11365.n236 GND 0.342588f
C753 a_185229_n11365.n237 GND 0.200066f
C754 a_185229_n11365.n238 GND 0.011088f
C755 a_185229_n11365.n239 GND 0.003895f
C756 a_185229_n11365.t3 GND 0.04886f
C757 a_185229_n11365.n240 GND 0.004124f
C758 a_185229_n11365.n241 GND 0.004124f
C759 a_185229_n11365.n242 GND 0.003895f
C760 a_185229_n11365.n243 GND 0.010936f
C761 a_185229_n11365.n244 GND 0.010557f
C762 a_185229_n11365.n245 GND 0.009005f
C763 a_185229_n11365.n246 GND 0.008838f
C764 a_185229_n11365.t17 GND 0.04886f
C765 a_185229_n11365.n247 GND 0.100636f
C766 a_185229_n11365.n248 GND 0.006907f
C767 a_185229_n11365.n249 GND 0.033198f
C768 a_185229_n11365.n250 GND 0.342588f
C769 a_185229_n11365.n251 GND 0.200066f
C770 a_185229_n11365.n252 GND 0.011088f
C771 a_185229_n11365.n253 GND 0.003895f
C772 a_185229_n11365.t14 GND 0.04886f
C773 a_185229_n11365.n254 GND 0.004124f
C774 a_185229_n11365.n255 GND 0.004124f
C775 a_185229_n11365.n256 GND 0.003895f
C776 a_185229_n11365.n257 GND 0.010936f
C777 a_185229_n11365.n258 GND 0.010557f
C778 a_185229_n11365.n259 GND 0.009005f
C779 a_185229_n11365.n260 GND 0.008838f
C780 a_185229_n11365.t8 GND 0.04886f
C781 a_185229_n11365.n261 GND 0.100636f
C782 a_185229_n11365.n262 GND 0.006907f
C783 a_185229_n11365.n263 GND 0.033198f
C784 a_185229_n11365.n264 GND 0.342588f
C785 a_185229_n11365.n265 GND 0.200066f
C786 a_185229_n11365.n266 GND 0.011088f
C787 a_185229_n11365.n267 GND 0.003895f
C788 a_185229_n11365.t5 GND 0.04886f
C789 a_185229_n11365.n268 GND 0.004124f
C790 a_185229_n11365.n269 GND 0.004124f
C791 a_185229_n11365.n270 GND 0.003895f
C792 a_185229_n11365.n271 GND 0.010936f
C793 a_185229_n11365.n272 GND 0.010557f
C794 a_185229_n11365.n273 GND 0.009005f
C795 a_185229_n11365.n274 GND 0.008838f
C796 a_185229_n11365.t22 GND 0.04886f
C797 a_185229_n11365.n275 GND 0.100636f
C798 a_185229_n11365.n276 GND 0.006907f
C799 a_185229_n11365.n277 GND 0.033198f
C800 a_185229_n11365.n278 GND 0.347642f
C801 a_185229_n11365.n279 GND 0.200066f
C802 a_185229_n11365.n280 GND 0.011088f
C803 a_185229_n11365.n281 GND 0.003895f
C804 a_185229_n11365.t23 GND 0.04886f
C805 a_185229_n11365.n282 GND 0.004124f
C806 a_185229_n11365.n283 GND 0.004124f
C807 a_185229_n11365.n284 GND 0.003895f
C808 a_185229_n11365.n285 GND 0.010936f
C809 a_185229_n11365.n286 GND 0.010557f
C810 a_185229_n11365.n287 GND 0.009005f
C811 a_185229_n11365.n288 GND 0.008838f
C812 a_185229_n11365.t20 GND 0.04886f
C813 a_185229_n11365.n289 GND 0.100636f
C814 a_185229_n11365.n290 GND 0.006907f
C815 a_185229_n11365.n291 GND 0.033198f
C816 a_185229_n11365.n292 GND 0.342588f
C817 a_185229_n11365.n293 GND 0.200066f
C818 a_185229_n11365.n294 GND 0.011088f
C819 a_185229_n11365.n295 GND 0.003895f
C820 a_185229_n11365.t18 GND 0.04886f
C821 a_185229_n11365.n296 GND 0.004124f
C822 a_185229_n11365.n297 GND 0.004124f
C823 a_185229_n11365.n298 GND 0.003895f
C824 a_185229_n11365.n299 GND 0.010936f
C825 a_185229_n11365.n300 GND 0.010557f
C826 a_185229_n11365.n301 GND 0.009005f
C827 a_185229_n11365.n302 GND 0.008838f
C828 a_185229_n11365.t15 GND 0.04886f
C829 a_185229_n11365.n303 GND 0.100636f
C830 a_185229_n11365.n304 GND 0.006907f
C831 a_185229_n11365.n305 GND 0.033198f
C832 a_185229_n11365.n306 GND 0.342588f
C833 a_185229_n11365.n307 GND 0.200066f
C834 a_185229_n11365.n308 GND 0.011088f
C835 a_185229_n11365.n309 GND 0.003895f
C836 a_185229_n11365.t10 GND 0.04886f
C837 a_185229_n11365.n310 GND 0.004124f
C838 a_185229_n11365.n311 GND 0.004124f
C839 a_185229_n11365.n312 GND 0.003895f
C840 a_185229_n11365.n313 GND 0.010936f
C841 a_185229_n11365.n314 GND 0.010557f
C842 a_185229_n11365.n315 GND 0.009005f
C843 a_185229_n11365.n316 GND 0.008838f
C844 a_185229_n11365.t21 GND 0.04886f
C845 a_185229_n11365.n317 GND 0.100636f
C846 a_185229_n11365.n318 GND 0.006907f
C847 a_185229_n11365.n319 GND 0.033198f
C848 a_185229_n11365.n320 GND 0.790823f
C849 a_185229_n11365.n321 GND 1.82417f
C850 a_185229_n11365.n322 GND 0.110583f
C851 a_185229_n11365.n323 GND 0.106949f
C852 a_185229_n11365.t54 GND 0.269595f
C853 a_185229_n11365.n324 GND 0.104449f
C854 a_185229_n11365.t61 GND 0.269595f
C855 a_185229_n11365.n325 GND 0.104449f
C856 a_185229_n11365.n326 GND 0.104449f
C857 a_185229_n11365.t37 GND 0.269595f
C858 a_185229_n11365.n327 GND 0.104449f
C859 a_185229_n11365.t45 GND 0.269595f
C860 a_185229_n11365.n328 GND 0.104449f
C861 a_185229_n11365.n329 GND 0.104449f
C862 a_185229_n11365.t49 GND 0.269595f
C863 a_185229_n11365.n330 GND 0.104449f
C864 a_185229_n11365.t39 GND 0.269595f
C865 a_185229_n11365.n331 GND 0.104449f
C866 a_185229_n11365.n332 GND 0.104449f
C867 a_185229_n11365.t46 GND 0.269595f
C868 a_185229_n11365.n333 GND 0.104449f
C869 a_185229_n11365.t64 GND 0.269595f
C870 a_185229_n11365.n334 GND 0.154394f
C871 a_185229_n11365.n335 GND 0.607988f
C872 a_185229_n11365.t25 GND 0.829336f
C873 a_185229_n11365.n336 GND 9.19451f
C874 a_185229_n11365.t2 GND 0.929383f
C875 VREFN.t24 GND 0.013743f
C876 VREFN.t21 GND 0.013743f
C877 VREFN.n0 GND 0.037182f
C878 VREFN.t19 GND 0.013743f
C879 VREFN.t20 GND 0.013743f
C880 VREFN.n1 GND 0.037057f
C881 VREFN.n2 GND 0.133023f
C882 VREFN.t18 GND 0.013743f
C883 VREFN.t13 GND 0.013743f
C884 VREFN.n3 GND 0.037133f
C885 VREFN.n4 GND 0.065415f
C886 VREFN.t10 GND 0.013743f
C887 VREFN.t9 GND 0.013743f
C888 VREFN.n5 GND 0.037057f
C889 VREFN.n6 GND 0.064492f
C890 VREFN.t25 GND 0.013743f
C891 VREFN.t22 GND 0.013743f
C892 VREFN.n7 GND 0.037133f
C893 VREFN.n8 GND 0.065415f
C894 VREFN.t16 GND 0.013743f
C895 VREFN.t15 GND 0.013743f
C896 VREFN.n9 GND 0.037057f
C897 VREFN.n10 GND 0.064492f
C898 VREFN.t12 GND 0.013743f
C899 VREFN.t14 GND 0.013743f
C900 VREFN.n11 GND 0.037057f
C901 VREFN.n12 GND 0.065325f
C902 VREFN.t11 GND 0.013743f
C903 VREFN.t27 GND 0.013743f
C904 VREFN.n13 GND 0.037133f
C905 VREFN.n14 GND 0.065415f
C906 VREFN.t26 GND 0.013743f
C907 VREFN.t23 GND 0.013743f
C908 VREFN.n15 GND 0.037057f
C909 VREFN.n16 GND 0.064492f
C910 VREFN.t17 GND 0.055906f
C911 VREFN.n17 GND 0.123421f
C912 VREFN.n18 GND 0.129476f
C913 VREFN.t51 GND 0.064489f
C914 VREFN.t50 GND 0.013743f
C915 VREFN.t48 GND 0.013743f
C916 VREFN.n19 GND 0.048631f
C917 VREFN.n20 GND 0.116908f
C918 VREFN.t49 GND 0.013743f
C919 VREFN.t47 GND 0.013743f
C920 VREFN.n21 GND 0.0488f
C921 VREFN.n22 GND 0.052139f
C922 VREFN.t55 GND 0.013743f
C923 VREFN.t54 GND 0.013743f
C924 VREFN.n23 GND 0.048631f
C925 VREFN.n24 GND 0.051308f
C926 VREFN.t53 GND 0.013743f
C927 VREFN.t52 GND 0.013743f
C928 VREFN.n25 GND 0.0488f
C929 VREFN.n26 GND 0.153604f
C930 VREFN.n27 GND 2.7833f
C931 VREFN.t43 GND 0.013743f
C932 VREFN.t40 GND 0.013743f
C933 VREFN.n28 GND 0.037182f
C934 VREFN.t38 GND 0.013743f
C935 VREFN.t39 GND 0.013743f
C936 VREFN.n29 GND 0.037057f
C937 VREFN.n30 GND 0.133023f
C938 VREFN.t37 GND 0.013743f
C939 VREFN.t32 GND 0.013743f
C940 VREFN.n31 GND 0.037133f
C941 VREFN.n32 GND 0.065415f
C942 VREFN.t29 GND 0.013743f
C943 VREFN.t28 GND 0.013743f
C944 VREFN.n33 GND 0.037057f
C945 VREFN.n34 GND 0.064492f
C946 VREFN.t44 GND 0.013743f
C947 VREFN.t41 GND 0.013743f
C948 VREFN.n35 GND 0.037133f
C949 VREFN.n36 GND 0.065415f
C950 VREFN.t35 GND 0.013743f
C951 VREFN.t34 GND 0.013743f
C952 VREFN.n37 GND 0.037057f
C953 VREFN.n38 GND 0.064492f
C954 VREFN.t31 GND 0.013743f
C955 VREFN.t33 GND 0.013743f
C956 VREFN.n39 GND 0.037057f
C957 VREFN.n40 GND 0.065325f
C958 VREFN.t30 GND 0.013743f
C959 VREFN.t46 GND 0.013743f
C960 VREFN.n41 GND 0.037133f
C961 VREFN.n42 GND 0.065415f
C962 VREFN.t45 GND 0.013743f
C963 VREFN.t42 GND 0.013743f
C964 VREFN.n43 GND 0.037057f
C965 VREFN.n44 GND 0.064492f
C966 VREFN.t36 GND 0.055906f
C967 VREFN.n45 GND 0.123421f
C968 VREFN.n46 GND 0.129476f
C969 VREFN.t4 GND 0.064489f
C970 VREFN.t3 GND 0.013743f
C971 VREFN.t1 GND 0.013743f
C972 VREFN.n47 GND 0.048631f
C973 VREFN.n48 GND 0.116908f
C974 VREFN.t2 GND 0.013743f
C975 VREFN.t0 GND 0.013743f
C976 VREFN.n49 GND 0.0488f
C977 VREFN.n50 GND 0.052139f
C978 VREFN.t8 GND 0.013743f
C979 VREFN.t7 GND 0.013743f
C980 VREFN.n51 GND 0.048631f
C981 VREFN.n52 GND 0.051308f
C982 VREFN.t6 GND 0.013743f
C983 VREFN.t5 GND 0.013743f
C984 VREFN.n53 GND 0.0488f
C985 VREFN.n54 GND 0.153604f
C986 VREFN.n55 GND 1.02118f
C987 VREFN.n56 GND 14.304099f
C988 a_181475_n46496.t4 GND 0.105853f
C989 a_181475_n46496.t1 GND 0.105853f
C990 a_181475_n46496.t0 GND 0.105853f
C991 a_181475_n46496.n0 GND 0.355165f
C992 a_181475_n46496.t12 GND 0.156137f
C993 a_181475_n46496.t13 GND 0.156078f
C994 a_181475_n46496.n1 GND 0.460192f
C995 a_181475_n46496.t25 GND 0.156078f
C996 a_181475_n46496.n2 GND 0.202861f
C997 a_181475_n46496.t29 GND 0.156078f
C998 a_181475_n46496.n3 GND 0.202861f
C999 a_181475_n46496.t11 GND 0.156078f
C1000 a_181475_n46496.n4 GND 0.202861f
C1001 a_181475_n46496.t23 GND 0.156078f
C1002 a_181475_n46496.n5 GND 0.202861f
C1003 a_181475_n46496.t24 GND 0.156078f
C1004 a_181475_n46496.n6 GND 0.202861f
C1005 a_181475_n46496.t6 GND 0.156078f
C1006 a_181475_n46496.n7 GND 0.202861f
C1007 a_181475_n46496.t10 GND 0.156078f
C1008 a_181475_n46496.n8 GND 0.382422f
C1009 a_181475_n46496.t21 GND 0.156079f
C1010 a_181475_n46496.t7 GND 0.156079f
C1011 a_181475_n46496.t27 GND 0.156079f
C1012 a_181475_n46496.t26 GND 0.156079f
C1013 a_181475_n46496.t22 GND 0.156079f
C1014 a_181475_n46496.t8 GND 0.156079f
C1015 a_181475_n46496.t28 GND 0.156079f
C1016 a_181475_n46496.t15 GND 0.156079f
C1017 a_181475_n46496.t14 GND 0.156079f
C1018 a_181475_n46496.t9 GND 0.156122f
C1019 a_181475_n46496.n9 GND 0.400211f
C1020 a_181475_n46496.n10 GND 0.213278f
C1021 a_181475_n46496.n11 GND 0.213278f
C1022 a_181475_n46496.n12 GND 0.213278f
C1023 a_181475_n46496.n13 GND 0.213278f
C1024 a_181475_n46496.n14 GND 0.213278f
C1025 a_181475_n46496.n15 GND 0.213278f
C1026 a_181475_n46496.n16 GND 0.213278f
C1027 a_181475_n46496.n17 GND 0.324368f
C1028 a_181475_n46496.n18 GND 2.39091f
C1029 a_181475_n46496.t31 GND 0.155249f
C1030 a_181475_n46496.n19 GND 0.995725f
C1031 a_181475_n46496.t33 GND 0.155249f
C1032 a_181475_n46496.n20 GND 0.150788f
C1033 a_181475_n46496.t18 GND 0.155249f
C1034 a_181475_n46496.n21 GND 0.150788f
C1035 a_181475_n46496.t19 GND 0.155249f
C1036 a_181475_n46496.n22 GND 0.150788f
C1037 a_181475_n46496.t30 GND 0.155249f
C1038 a_181475_n46496.n23 GND 0.62113f
C1039 a_181475_n46496.t20 GND 0.155249f
C1040 a_181475_n46496.n24 GND 0.734886f
C1041 a_181475_n46496.t17 GND 0.155249f
C1042 a_181475_n46496.n25 GND 0.19898f
C1043 a_181475_n46496.t16 GND 0.155249f
C1044 a_181475_n46496.n26 GND 0.19898f
C1045 a_181475_n46496.t32 GND 0.155249f
C1046 a_181475_n46496.n27 GND 0.908992f
C1047 a_181475_n46496.n28 GND 0.928431f
C1048 a_181475_n46496.n29 GND 1.87243f
C1049 a_181475_n46496.t3 GND 0.105853f
C1050 a_181475_n46496.t2 GND 0.105853f
C1051 a_181475_n46496.n30 GND 0.318799f
C1052 a_181475_n46496.n31 GND 1.05381f
C1053 a_181475_n46496.n32 GND 1.11674f
C1054 a_181475_n46496.n33 GND 0.277395f
C1055 a_181475_n46496.t5 GND 0.105853f
C1056 1Bit_DAC_Inv_0.OUT.t38 GND 0.365303f
C1057 1Bit_DAC_Inv_0.OUT.t37 GND 0.088589f
C1058 1Bit_DAC_Inv_0.OUT.t36 GND 0.088589f
C1059 1Bit_DAC_Inv_0.OUT.n0 GND 0.24434f
C1060 1Bit_DAC_Inv_0.OUT.n1 GND 1.2488f
C1061 1Bit_DAC_Inv_0.OUT.t30 GND 0.088589f
C1062 1Bit_DAC_Inv_0.OUT.t35 GND 0.088589f
C1063 1Bit_DAC_Inv_0.OUT.n2 GND 0.24458f
C1064 1Bit_DAC_Inv_0.OUT.n3 GND 0.620479f
C1065 1Bit_DAC_Inv_0.OUT.t29 GND 0.088589f
C1066 1Bit_DAC_Inv_0.OUT.t28 GND 0.088589f
C1067 1Bit_DAC_Inv_0.OUT.n4 GND 0.24434f
C1068 1Bit_DAC_Inv_0.OUT.n5 GND 0.614814f
C1069 1Bit_DAC_Inv_0.OUT.t27 GND 0.088589f
C1070 1Bit_DAC_Inv_0.OUT.t22 GND 0.088589f
C1071 1Bit_DAC_Inv_0.OUT.n6 GND 0.24434f
C1072 1Bit_DAC_Inv_0.OUT.n7 GND 0.630921f
C1073 1Bit_DAC_Inv_0.OUT.t20 GND 0.088589f
C1074 1Bit_DAC_Inv_0.OUT.t33 GND 0.088589f
C1075 1Bit_DAC_Inv_0.OUT.n8 GND 0.244487f
C1076 1Bit_DAC_Inv_0.OUT.n9 GND 0.63131f
C1077 1Bit_DAC_Inv_0.OUT.t32 GND 0.088589f
C1078 1Bit_DAC_Inv_0.OUT.t31 GND 0.088589f
C1079 1Bit_DAC_Inv_0.OUT.n10 GND 0.244487f
C1080 1Bit_DAC_Inv_0.OUT.n11 GND 0.63131f
C1081 1Bit_DAC_Inv_0.OUT.t26 GND 0.088589f
C1082 1Bit_DAC_Inv_0.OUT.t24 GND 0.088589f
C1083 1Bit_DAC_Inv_0.OUT.n12 GND 0.24434f
C1084 1Bit_DAC_Inv_0.OUT.n13 GND 0.630921f
C1085 1Bit_DAC_Inv_0.OUT.t25 GND 0.088589f
C1086 1Bit_DAC_Inv_0.OUT.t23 GND 0.088589f
C1087 1Bit_DAC_Inv_0.OUT.n14 GND 0.24458f
C1088 1Bit_DAC_Inv_0.OUT.n15 GND 0.612426f
C1089 1Bit_DAC_Inv_0.OUT.t21 GND 0.088589f
C1090 1Bit_DAC_Inv_0.OUT.t34 GND 0.088589f
C1091 1Bit_DAC_Inv_0.OUT.n16 GND 0.24434f
C1092 1Bit_DAC_Inv_0.OUT.n17 GND 0.691268f
C1093 1Bit_DAC_Inv_0.OUT.t51 GND 0.088589f
C1094 1Bit_DAC_Inv_0.OUT.t54 GND 0.088589f
C1095 1Bit_DAC_Inv_0.OUT.n18 GND 0.31648f
C1096 1Bit_DAC_Inv_0.OUT.t55 GND 0.088589f
C1097 1Bit_DAC_Inv_0.OUT.t2 GND 0.088589f
C1098 1Bit_DAC_Inv_0.OUT.n19 GND 0.318679f
C1099 1Bit_DAC_Inv_0.OUT.n20 GND 1.02282f
C1100 1Bit_DAC_Inv_0.OUT.t53 GND 0.088589f
C1101 1Bit_DAC_Inv_0.OUT.t3 GND 0.088589f
C1102 1Bit_DAC_Inv_0.OUT.n21 GND 0.318402f
C1103 1Bit_DAC_Inv_0.OUT.n22 GND 0.480253f
C1104 1Bit_DAC_Inv_0.OUT.t42 GND 0.088589f
C1105 1Bit_DAC_Inv_0.OUT.t5 GND 0.088589f
C1106 1Bit_DAC_Inv_0.OUT.n23 GND 0.318679f
C1107 1Bit_DAC_Inv_0.OUT.n24 GND 0.480512f
C1108 1Bit_DAC_Inv_0.OUT.t0 GND 0.413331f
C1109 1Bit_DAC_Inv_0.OUT.n25 GND 0.504784f
C1110 1Bit_DAC_Inv_0.OUT.n26 GND 0.057712f
C1111 1Bit_DAC_Inv_0.OUT.n27 GND 0.159171f
C1112 1Bit_DAC_Inv_0.OUT.t41 GND 4.31233f
C1113 1Bit_DAC_Inv_0.OUT.t40 GND 0.088589f
C1114 1Bit_DAC_Inv_0.OUT.t46 GND 0.088589f
C1115 1Bit_DAC_Inv_0.OUT.n28 GND 0.244774f
C1116 1Bit_DAC_Inv_0.OUT.n29 GND 19.1831f
C1117 1Bit_DAC_Inv_0.OUT.t43 GND 0.088589f
C1118 1Bit_DAC_Inv_0.OUT.t45 GND 0.088589f
C1119 1Bit_DAC_Inv_0.OUT.n30 GND 0.244504f
C1120 1Bit_DAC_Inv_0.OUT.n31 GND 0.842028f
C1121 1Bit_DAC_Inv_0.OUT.t49 GND 0.088589f
C1122 1Bit_DAC_Inv_0.OUT.t8 GND 0.088589f
C1123 1Bit_DAC_Inv_0.OUT.n32 GND 0.244261f
C1124 1Bit_DAC_Inv_0.OUT.n33 GND 0.900257f
C1125 1Bit_DAC_Inv_0.OUT.t6 GND 0.088589f
C1126 1Bit_DAC_Inv_0.OUT.t56 GND 0.088589f
C1127 1Bit_DAC_Inv_0.OUT.n34 GND 0.244261f
C1128 1Bit_DAC_Inv_0.OUT.n35 GND 0.900257f
C1129 1Bit_DAC_Inv_0.OUT.t1 GND 0.088589f
C1130 1Bit_DAC_Inv_0.OUT.t7 GND 0.088589f
C1131 1Bit_DAC_Inv_0.OUT.n36 GND 0.244515f
C1132 1Bit_DAC_Inv_0.OUT.n37 GND 0.780115f
C1133 1Bit_DAC_Inv_0.OUT.t17 GND 0.413331f
C1134 1Bit_DAC_Inv_0.OUT.n38 GND 0.644054f
C1135 1Bit_DAC_Inv_0.OUT.t9 GND 0.088589f
C1136 1Bit_DAC_Inv_0.OUT.t10 GND 0.088589f
C1137 1Bit_DAC_Inv_0.OUT.n39 GND 0.244774f
C1138 1Bit_DAC_Inv_0.OUT.n40 GND 0.735451f
C1139 1Bit_DAC_Inv_0.OUT.t12 GND 0.088589f
C1140 1Bit_DAC_Inv_0.OUT.t11 GND 0.088589f
C1141 1Bit_DAC_Inv_0.OUT.n41 GND 0.318679f
C1142 1Bit_DAC_Inv_0.OUT.n42 GND 0.581987f
C1143 1Bit_DAC_Inv_0.OUT.t47 GND 0.088589f
C1144 1Bit_DAC_Inv_0.OUT.t39 GND 0.088589f
C1145 1Bit_DAC_Inv_0.OUT.n43 GND 0.244774f
C1146 1Bit_DAC_Inv_0.OUT.n44 GND 0.710217f
C1147 1Bit_DAC_Inv_0.OUT.t15 GND 0.088589f
C1148 1Bit_DAC_Inv_0.OUT.t18 GND 0.088589f
C1149 1Bit_DAC_Inv_0.OUT.n45 GND 0.318402f
C1150 1Bit_DAC_Inv_0.OUT.n46 GND 0.531259f
C1151 1Bit_DAC_Inv_0.OUT.t52 GND 0.088589f
C1152 1Bit_DAC_Inv_0.OUT.t4 GND 0.088589f
C1153 1Bit_DAC_Inv_0.OUT.n47 GND 0.244504f
C1154 1Bit_DAC_Inv_0.OUT.n48 GND 0.729278f
C1155 1Bit_DAC_Inv_0.OUT.t19 GND 0.088589f
C1156 1Bit_DAC_Inv_0.OUT.t13 GND 0.088589f
C1157 1Bit_DAC_Inv_0.OUT.n49 GND 0.318679f
C1158 1Bit_DAC_Inv_0.OUT.n50 GND 0.581987f
C1159 1Bit_DAC_Inv_0.OUT.t48 GND 0.088589f
C1160 1Bit_DAC_Inv_0.OUT.t44 GND 0.088589f
C1161 1Bit_DAC_Inv_0.OUT.n51 GND 0.244261f
C1162 1Bit_DAC_Inv_0.OUT.n52 GND 0.723078f
C1163 1Bit_DAC_Inv_0.OUT.t16 GND 0.088589f
C1164 1Bit_DAC_Inv_0.OUT.t14 GND 0.088589f
C1165 1Bit_DAC_Inv_0.OUT.n53 GND 0.318679f
C1166 1Bit_DAC_Inv_0.OUT.n54 GND 0.581987f
C1167 1Bit_DAC_Inv_0.OUT.t50 GND 0.364423f
C1168 1Bit_DAC_Inv_0.OUT.n55 GND 0.771236f
C1169 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n0 GND 1.66014f
C1170 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n1 GND 1.71545f
C1171 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n2 GND 1.71025f
C1172 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n3 GND 0.055365f
C1173 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n4 GND 0.223603f
C1174 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n5 GND 0.055354f
C1175 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n6 GND 0.22333f
C1176 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t10 GND 0.026782f
C1177 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t13 GND 0.026782f
C1178 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n7 GND 0.080784f
C1179 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n8 GND 0.259053f
C1180 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t12 GND 0.026782f
C1181 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t11 GND 0.026782f
C1182 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n9 GND 0.07048f
C1183 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n10 GND 0.019099f
C1184 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n11 GND 0.006117f
C1185 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n12 GND 0.00427f
C1186 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t3 GND 0.006695f
C1187 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t7 GND 0.006695f
C1188 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n13 GND 0.007096f
C1189 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n14 GND 0.00545f
C1190 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n15 GND 0.013391f
C1191 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n16 GND 0.002585f
C1192 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n17 GND 0.00996f
C1193 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n18 GND 0.016925f
C1194 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t26 GND 0.289853f
C1195 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n19 GND 0.098788f
C1196 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n20 GND 0.108669f
C1197 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t0 GND 0.126379f
C1198 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n21 GND 0.009972f
C1199 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n22 GND 0.044247f
C1200 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n23 GND 0.108669f
C1201 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n24 GND 0.108669f
C1202 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n25 GND 0.108669f
C1203 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n26 GND 0.108669f
C1204 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n27 GND 0.108669f
C1205 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n28 GND 0.108669f
C1206 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n29 GND 0.167531f
C1207 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n30 GND 0.22454f
C1208 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n31 GND 0.108669f
C1209 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n32 GND 0.108669f
C1210 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n33 GND 0.108669f
C1211 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n34 GND 0.108669f
C1212 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n35 GND 0.108669f
C1213 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n36 GND 0.176677f
C1214 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t42 GND 0.289853f
C1215 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n37 GND 0.224017f
C1216 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t44 GND 0.289853f
C1217 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n38 GND 0.108669f
C1218 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n39 GND 0.108669f
C1219 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t38 GND 0.289853f
C1220 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n40 GND 0.108669f
C1221 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t18 GND 0.289853f
C1222 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n41 GND 0.108669f
C1223 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n42 GND 0.108669f
C1224 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t25 GND 0.289853f
C1225 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n43 GND 0.108669f
C1226 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t33 GND 0.289853f
C1227 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n44 GND 0.108669f
C1228 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n45 GND 0.108669f
C1229 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t21 GND 0.289853f
C1230 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n46 GND 0.108669f
C1231 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t31 GND 0.289853f
C1232 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n47 GND 0.108669f
C1233 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n48 GND 0.108669f
C1234 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t45 GND 0.289853f
C1235 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n49 GND 0.108669f
C1236 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t16 GND 0.289853f
C1237 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n50 GND 0.108669f
C1238 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n51 GND 0.108669f
C1239 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t23 GND 0.289853f
C1240 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n52 GND 0.108669f
C1241 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t27 GND 0.289853f
C1242 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n53 GND 0.177902f
C1243 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t32 GND 0.289853f
C1244 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n54 GND 0.167528f
C1245 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n55 GND 0.108669f
C1246 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t22 GND 0.289853f
C1247 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n56 GND 0.108669f
C1248 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t19 GND 0.289853f
C1249 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n57 GND 0.108669f
C1250 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n58 GND 0.108669f
C1251 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t47 GND 0.289853f
C1252 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n59 GND 0.108669f
C1253 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t28 GND 0.289853f
C1254 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n60 GND 0.108669f
C1255 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n61 GND 0.108669f
C1256 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t24 GND 0.289853f
C1257 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n62 GND 0.108669f
C1258 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t17 GND 0.289853f
C1259 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n63 GND 0.108669f
C1260 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n64 GND 0.108669f
C1261 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t29 GND 0.289853f
C1262 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n65 GND 0.108669f
C1263 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t20 GND 0.289853f
C1264 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n66 GND 0.108669f
C1265 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n67 GND 0.108669f
C1266 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t41 GND 0.289853f
C1267 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n68 GND 0.108669f
C1268 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t34 GND 0.289853f
C1269 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n69 GND 0.108669f
C1270 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n70 GND 0.108669f
C1271 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t40 GND 0.289853f
C1272 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n71 GND 0.108669f
C1273 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t37 GND 0.289853f
C1274 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n72 GND 0.108669f
C1275 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n73 GND 0.166527f
C1276 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t30 GND 0.289853f
C1277 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n74 GND 0.166527f
C1278 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n75 GND 1.65709f
C1279 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n76 GND 0.566584f
C1280 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t15 GND 0.026782f
C1281 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t14 GND 0.026782f
C1282 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n77 GND 0.07048f
C1283 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n78 GND 0.622075f
C1284 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n79 GND 0.201345f
C1285 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n80 GND 0.006117f
C1286 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n81 GND 0.00427f
C1287 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t1 GND 0.006695f
C1288 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n82 GND 0.002585f
C1289 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t5 GND 0.006695f
C1290 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n83 GND 0.013391f
C1291 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n84 GND 0.00545f
C1292 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n85 GND 0.007072f
C1293 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n86 GND 0.019052f
C1294 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t2 GND 0.126372f
C1295 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n87 GND 0.03609f
C1296 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t9 GND 0.013391f
C1297 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t8 GND 0.013391f
C1298 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n88 GND 0.060699f
C1299 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n89 GND 0.160597f
C1300 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n90 GND 0.036089f
C1301 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t4 GND 0.126372f
C1302 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n91 GND 0.044482f
C1303 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n92 GND 0.017099f
C1304 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n93 GND 0.067599f
C1305 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t36 GND 0.289853f
C1306 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n94 GND 0.098988f
C1307 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n95 GND 0.238659f
C1308 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t39 GND 0.289858f
C1309 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t46 GND 0.289853f
C1310 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n96 GND 0.105933f
C1311 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n97 GND 0.10596f
C1312 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t35 GND 0.289853f
C1313 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n98 GND 0.108669f
C1314 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n99 GND 0.238899f
C1315 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t43 GND 0.289858f
C1316 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n100 GND 0.066709f
C1317 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.t6 GND 0.12638f
C1318 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n101 GND 0.200054f
C1319 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n102 GND 0.620464f
C1320 1Bit_Clk_ADC_0.C2S2_Fingers_Amplifier_0.constant_gm_fingers_0.Vout.n103 GND 0.569359f
C1321 a_218222_n27786.t8 GND 0.194162f
C1322 a_218222_n27786.t2 GND 0.235357f
C1323 a_218222_n27786.t5 GND 0.10698f
C1324 a_218222_n27786.n0 GND 1.51993f
C1325 a_218222_n27786.n1 GND 0.200489f
C1326 a_218222_n27786.t4 GND 0.009165f
C1327 a_218222_n27786.t1 GND 0.009165f
C1328 a_218222_n27786.n2 GND 0.032429f
C1329 a_218222_n27786.n3 GND 0.095728f
C1330 a_218222_n27786.t3 GND 0.009165f
C1331 a_218222_n27786.t6 GND 0.009165f
C1332 a_218222_n27786.n4 GND 0.038664f
C1333 a_218222_n27786.n5 GND 0.110693f
C1334 a_218222_n27786.t7 GND 0.009165f
C1335 a_218222_n27786.t9 GND 0.009165f
C1336 a_218222_n27786.n6 GND 0.032429f
C1337 a_218222_n27786.n7 GND 0.095668f
C1338 a_218222_n27786.n8 GND 0.194927f
C1339 a_218222_n27786.n9 GND 1.28053f
C1340 a_218222_n27786.t0 GND 0.107029f
C1341 a_220333_n26938.n0 GND 0.224177f
C1342 a_220333_n26938.n1 GND 0.580261f
C1343 a_220333_n26938.n2 GND 0.281977f
C1344 a_220333_n26938.n3 GND 0.060445f
C1345 a_220333_n26938.n4 GND 0.358112f
C1346 a_220333_n26938.n5 GND 0.060445f
C1347 a_220333_n26938.n6 GND 0.358203f
C1348 a_220333_n26938.n7 GND 1.26025f
C1349 a_220333_n26938.n8 GND 0.94806f
C1350 a_220333_n26938.n9 GND 0.272686f
C1351 a_220333_n26938.n10 GND 0.414211f
C1352 a_220333_n26938.n11 GND 0.361457f
C1353 a_220333_n26938.n12 GND 0.223547f
C1354 a_220333_n26938.n13 GND 0.061415f
C1355 a_220333_n26938.n14 GND 0.368761f
C1356 a_220333_n26938.n15 GND 0.220921f
C1357 a_220333_n26938.n16 GND 0.044676f
C1358 a_220333_n26938.n17 GND 0.026567f
C1359 a_220333_n26938.n18 GND 0.011146f
C1360 a_220333_n26938.n19 GND 0.044676f
C1361 a_220333_n26938.n20 GND 0.026567f
C1362 a_220333_n26938.n21 GND 0.011146f
C1363 a_220333_n26938.n22 GND 0.246237f
C1364 a_220333_n26938.n23 GND 0.246237f
C1365 a_220333_n26938.n24 GND 0.026567f
C1366 a_220333_n26938.n25 GND 0.026567f
C1367 a_220333_n26938.n26 GND 0.026567f
C1368 a_220333_n26938.n27 GND 0.026567f
C1369 a_220333_n26938.n28 GND 0.027418f
C1370 a_220333_n26938.n29 GND 0.026567f
C1371 a_220333_n26938.n30 GND 0.026567f
C1372 a_220333_n26938.n31 GND 0.026567f
C1373 a_220333_n26938.n32 GND 0.026492f
C1374 a_220333_n26938.n33 GND 0.026567f
C1375 a_220333_n26938.n34 GND 0.026567f
C1376 a_220333_n26938.n35 GND 0.026567f
C1377 a_220333_n26938.n36 GND 0.026567f
C1378 a_220333_n26938.n37 GND 0.027418f
C1379 a_220333_n26938.n38 GND 0.006751f
C1380 a_220333_n26938.n39 GND 0.009775f
C1381 a_220333_n26938.n40 GND 0.009775f
C1382 a_220333_n26938.n41 GND 0.004636f
C1383 a_220333_n26938.n42 GND 0.013284f
C1384 a_220333_n26938.n43 GND 0.009775f
C1385 a_220333_n26938.n44 GND 0.013496f
C1386 a_220333_n26938.n45 GND 0.047048f
C1387 a_220333_n26938.n46 GND 0.011146f
C1388 a_220333_n26938.n47 GND 0.013496f
C1389 a_220333_n26938.n48 GND 0.047048f
C1390 a_220333_n26938.n49 GND 0.011146f
C1391 a_220333_n26938.n50 GND 0.008165f
C1392 a_220333_n26938.n51 GND 0.009311f
C1393 a_220333_n26938.n52 GND 0.564647f
C1394 a_220333_n26938.n53 GND 0.11767f
C1395 a_220333_n26938.n54 GND 0.563925f
C1396 a_220333_n26938.n55 GND 0.117768f
C1397 a_220333_n26938.n56 GND 0.162595f
C1398 a_220333_n26938.n57 GND 0.032543f
C1399 a_220333_n26938.n58 GND 0.162595f
C1400 a_220333_n26938.n59 GND 0.032543f
C1401 a_220333_n26938.n60 GND 0.004909f
C1402 a_220333_n26938.n61 GND 0.004909f
C1403 a_220333_n26938.n62 GND 0.004909f
C1404 a_220333_n26938.n63 GND 5.41e-19
C1405 a_220333_n26938.n64 GND 0.004909f
C1406 a_220333_n26938.t12 GND 0.058156f
C1407 a_220333_n26938.n65 GND 0.004909f
C1408 a_220333_n26938.n66 GND 0.004909f
C1409 a_220333_n26938.n67 GND 0.004909f
C1410 a_220333_n26938.n68 GND 0.004909f
C1411 a_220333_n26938.n69 GND 0.00585f
C1412 a_220333_n26938.n70 GND 0.011864f
C1413 a_220333_n26938.n71 GND 0.005755f
C1414 a_220333_n26938.t0 GND 0.022705f
C1415 a_220333_n26938.n72 GND 0.037585f
C1416 a_220333_n26938.n73 GND 0.004636f
C1417 a_220333_n26938.n74 GND 0.004909f
C1418 a_220333_n26938.n75 GND 0.02808f
C1419 a_220333_n26938.n76 GND 0.004636f
C1420 a_220333_n26938.n77 GND 0.004636f
C1421 a_220333_n26938.n78 GND 0.004636f
C1422 a_220333_n26938.n79 GND 0.004636f
C1423 a_220333_n26938.n80 GND 0.009139f
C1424 a_220333_n26938.n81 GND 0.009139f
C1425 a_220333_n26938.n82 GND 0.004636f
C1426 a_220333_n26938.n83 GND 0.004636f
C1427 a_220333_n26938.n84 GND 0.240763f
C1428 a_220333_n26938.t15 GND 0.634271f
C1429 a_220333_n26938.n85 GND 0.224177f
C1430 a_220333_n26938.t14 GND 0.058156f
C1431 a_220333_n26938.n86 GND 0.004909f
C1432 a_220333_n26938.n87 GND 0.004909f
C1433 a_220333_n26938.n88 GND 0.004909f
C1434 a_220333_n26938.n89 GND 0.004909f
C1435 a_220333_n26938.n90 GND 5.41e-19
C1436 a_220333_n26938.n91 GND 0.004909f
C1437 a_220333_n26938.n92 GND 0.004909f
C1438 a_220333_n26938.n93 GND 0.004909f
C1439 a_220333_n26938.t10 GND 0.058156f
C1440 a_220333_n26938.n94 GND 0.004909f
C1441 a_220333_n26938.n95 GND 0.004909f
C1442 a_220333_n26938.n96 GND 0.004909f
C1443 a_220333_n26938.n97 GND 0.004909f
C1444 a_220333_n26938.n98 GND 0.004909f
C1445 a_220333_n26938.n99 GND 5.41e-19
C1446 a_220333_n26938.n100 GND 0.004909f
C1447 a_220333_n26938.n101 GND 0.004909f
C1448 a_220333_n26938.n102 GND 0.004909f
C1449 a_220333_n26938.n103 GND 0.004636f
C1450 a_220333_n26938.n104 GND 0.004636f
C1451 a_220333_n26938.n105 GND 0.004636f
C1452 a_220333_n26938.n106 GND 0.004636f
C1453 a_220333_n26938.n107 GND 0.004636f
C1454 a_220333_n26938.n108 GND 0.009139f
C1455 a_220333_n26938.n109 GND 0.009139f
C1456 a_220333_n26938.n110 GND 0.004636f
C1457 a_220333_n26938.n111 GND 0.004636f
C1458 a_220333_n26938.n112 GND 0.006751f
C1459 a_220333_n26938.t8 GND 0.058156f
C1460 a_220333_n26938.n113 GND 0.116585f
C1461 a_220333_n26938.t27 GND 0.634271f
C1462 a_220333_n26938.n114 GND 0.240763f
C1463 a_220333_n26938.n115 GND 0.559694f
C1464 a_220333_n26938.t23 GND 0.634271f
C1465 a_220333_n26938.n116 GND 0.23991f
C1466 a_220333_n26938.t22 GND 0.634277f
C1467 a_220333_n26938.t19 GND 0.058156f
C1468 a_220333_n26938.t18 GND 0.058156f
C1469 a_220333_n26938.n117 GND 0.245256f
C1470 a_220333_n26938.t21 GND 0.058156f
C1471 a_220333_n26938.t17 GND 0.058156f
C1472 a_220333_n26938.n118 GND 0.245256f
C1473 a_220333_n26938.n119 GND 0.00585f
C1474 a_220333_n26938.n120 GND 0.011864f
C1475 a_220333_n26938.n121 GND 0.005755f
C1476 a_220333_n26938.t20 GND 0.022705f
C1477 a_220333_n26938.n122 GND 0.037585f
C1478 a_220333_n26938.n123 GND 0.004636f
C1479 a_220333_n26938.n124 GND 0.004909f
C1480 a_220333_n26938.n125 GND 0.02808f
C1481 a_220333_n26938.n126 GND 1.25657f
C1482 a_220333_n26938.n127 GND 0.519726f
C1483 a_220333_n26938.t9 GND 0.634277f
C1484 a_220333_n26938.n128 GND 0.223919f
C1485 a_220333_n26938.t7 GND 0.634271f
C1486 a_220333_n26938.t13 GND 0.634271f
C1487 a_220333_n26938.t5 GND 0.634271f
C1488 a_220333_n26938.n129 GND 5.48e-19
C1489 a_220333_n26938.t4 GND 0.029078f
C1490 a_220333_n26938.n130 GND 0.004909f
C1491 a_220333_n26938.n131 GND 0.010014f
C1492 a_220333_n26938.n132 GND 0.009273f
C1493 a_220333_n26938.n133 GND 0.005654f
C1494 a_220333_n26938.n134 GND 0.087871f
C1495 a_220333_n26938.t3 GND 0.200999f
C1496 a_220333_n26938.n135 GND 0.081473f
C1497 a_220333_n26938.t2 GND 0.029078f
C1498 a_220333_n26938.n136 GND 5.48e-19
C1499 a_220333_n26938.n137 GND 0.004909f
C1500 a_220333_n26938.n138 GND 0.010014f
C1501 a_220333_n26938.n139 GND 0.009273f
C1502 a_220333_n26938.n140 GND 0.005654f
C1503 a_220333_n26938.n141 GND 0.087871f
C1504 a_220333_n26938.n142 GND 0.081473f
C1505 a_220333_n26938.t1 GND 0.200999f
C1506 a_220333_n26938.n143 GND 0.006121f
C1507 a_220333_n26938.n144 GND 0.004636f
C1508 a_220333_n26938.n145 GND 0.004636f
C1509 a_220333_n26938.n146 GND 0.004636f
C1510 a_220333_n26938.n147 GND 0.009139f
C1511 a_220333_n26938.n148 GND 0.009139f
C1512 a_220333_n26938.n149 GND 0.004636f
C1513 a_220333_n26938.n150 GND 0.004636f
C1514 a_220333_n26938.n151 GND 0.006751f
C1515 a_220333_n26938.t6 GND 0.058156f
C1516 a_220333_n26938.n152 GND 0.116684f
C1517 a_220333_n26938.t24 GND 0.634271f
C1518 a_220333_n26938.n153 GND 0.223547f
C1519 a_220333_n26938.n154 GND 0.239955f
C1520 a_220333_n26938.t25 GND 0.634271f
C1521 a_220333_n26938.n155 GND 0.559878f
C1522 a_220333_n26938.t26 GND 0.634276f
C1523 a_220333_n26938.t11 GND 0.634276f
C1524 a_220333_n26938.n156 GND 0.008165f
C1525 a_220333_n26938.n157 GND 0.116585f
C1526 a_220333_n26938.t16 GND 0.058156f
C1527 C2S2_Amp_F_I_1.OUT.n0 GND 0.015806f
C1528 C2S2_Amp_F_I_1.OUT.n1 GND 0.005278f
C1529 C2S2_Amp_F_I_1.OUT.n2 GND 0.005314f
C1530 C2S2_Amp_F_I_1.OUT.n3 GND 0.001964f
C1531 C2S2_Amp_F_I_1.OUT.n4 GND 0.001855f
C1532 C2S2_Amp_F_I_1.OUT.n5 GND 0.011191f
C1533 C2S2_Amp_F_I_1.OUT.n6 GND 0.001964f
C1534 C2S2_Amp_F_I_1.OUT.n7 GND 0.006986f
C1535 C2S2_Amp_F_I_1.OUT.n8 GND 0.001855f
C1536 C2S2_Amp_F_I_1.OUT.n9 GND 0.005268f
C1537 C2S2_Amp_F_I_1.OUT.n10 GND 0.005081f
C1538 C2S2_Amp_F_I_1.OUT.n11 GND 0.001855f
C1539 C2S2_Amp_F_I_1.OUT.n12 GND 0.001855f
C1540 C2S2_Amp_F_I_1.OUT.n13 GND 0.001964f
C1541 C2S2_Amp_F_I_1.OUT.n14 GND 0.006328f
C1542 C2S2_Amp_F_I_1.OUT.n15 GND 0.006328f
C1543 C2S2_Amp_F_I_1.OUT.n16 GND 0.004746f
C1544 C2S2_Amp_F_I_1.OUT.n17 GND 0.002302f
C1545 C2S2_Amp_F_I_1.OUT.t20 GND 0.009083f
C1546 C2S2_Amp_F_I_1.OUT.n18 GND 0.015035f
C1547 C2S2_Amp_F_I_1.OUT.n19 GND 0.093309f
C1548 C2S2_Amp_F_I_1.OUT.n20 GND 0.001855f
C1549 C2S2_Amp_F_I_1.OUT.n21 GND 0.001964f
C1550 C2S2_Amp_F_I_1.OUT.n22 GND 0.006328f
C1551 C2S2_Amp_F_I_1.OUT.n23 GND 0.006328f
C1552 C2S2_Amp_F_I_1.OUT.n24 GND 0.001964f
C1553 C2S2_Amp_F_I_1.OUT.n25 GND 0.001855f
C1554 C2S2_Amp_F_I_1.OUT.n26 GND 0.005122f
C1555 C2S2_Amp_F_I_1.OUT.n27 GND 0.009666f
C1556 C2S2_Amp_F_I_1.OUT.n28 GND 0.998261f
C1557 C2S2_Amp_F_I_1.OUT.n29 GND 0.063616f
C1558 C2S2_Amp_F_I_1.OUT.t68 GND 30.136301f
C1559 C2S2_Amp_F_I_1.OUT.n30 GND 0.011449f
C1560 C2S2_Amp_F_I_1.OUT.n31 GND 0.096381f
C1561 C2S2_Amp_F_I_1.OUT.n32 GND 0.096381f
C1562 C2S2_Amp_F_I_1.OUT.n33 GND 0.096381f
C1563 C2S2_Amp_F_I_1.OUT.n34 GND 0.096381f
C1564 C2S2_Amp_F_I_1.OUT.n35 GND 0.096381f
C1565 C2S2_Amp_F_I_1.OUT.n36 GND 0.096381f
C1566 C2S2_Amp_F_I_1.OUT.n37 GND 0.096381f
C1567 C2S2_Amp_F_I_1.OUT.n38 GND 0.096381f
C1568 C2S2_Amp_F_I_1.OUT.n39 GND 0.096381f
C1569 C2S2_Amp_F_I_1.OUT.n40 GND 0.096381f
C1570 C2S2_Amp_F_I_1.OUT.n41 GND 0.096381f
C1571 C2S2_Amp_F_I_1.OUT.n42 GND 0.096381f
C1572 C2S2_Amp_F_I_1.OUT.n43 GND 0.096381f
C1573 C2S2_Amp_F_I_1.OUT.n44 GND 0.096381f
C1574 C2S2_Amp_F_I_1.OUT.n45 GND 0.096381f
C1575 C2S2_Amp_F_I_1.OUT.n46 GND 0.096381f
C1576 C2S2_Amp_F_I_1.OUT.n47 GND 0.096381f
C1577 C2S2_Amp_F_I_1.OUT.n48 GND 0.096381f
C1578 C2S2_Amp_F_I_1.OUT.n49 GND 0.002959f
C1579 C2S2_Amp_F_I_1.OUT.n50 GND 0.005207f
C1580 C2S2_Amp_F_I_1.OUT.n51 GND 0.001855f
C1581 C2S2_Amp_F_I_1.OUT.t63 GND 0.023264f
C1582 C2S2_Amp_F_I_1.OUT.n52 GND 0.003289f
C1583 C2S2_Amp_F_I_1.OUT.n53 GND 0.011449f
C1584 C2S2_Amp_F_I_1.OUT.n54 GND 0.00528f
C1585 C2S2_Amp_F_I_1.OUT.n55 GND 0.001855f
C1586 C2S2_Amp_F_I_1.OUT.n56 GND 0.001964f
C1587 C2S2_Amp_F_I_1.OUT.t42 GND 0.023264f
C1588 C2S2_Amp_F_I_1.OUT.n57 GND 0.04788f
C1589 C2S2_Amp_F_I_1.OUT.n58 GND 0.001964f
C1590 C2S2_Amp_F_I_1.OUT.n59 GND 0.004288f
C1591 C2S2_Amp_F_I_1.OUT.n60 GND 0.005191f
C1592 C2S2_Amp_F_I_1.OUT.n61 GND 0.09286f
C1593 C2S2_Amp_F_I_1.OUT.n62 GND 0.038409f
C1594 C2S2_Amp_F_I_1.OUT.n63 GND 0.00528f
C1595 C2S2_Amp_F_I_1.OUT.n64 GND 0.001855f
C1596 C2S2_Amp_F_I_1.OUT.t61 GND 0.023264f
C1597 C2S2_Amp_F_I_1.OUT.n65 GND 0.001964f
C1598 C2S2_Amp_F_I_1.OUT.n66 GND 0.001964f
C1599 C2S2_Amp_F_I_1.OUT.n67 GND 0.001855f
C1600 C2S2_Amp_F_I_1.OUT.n68 GND 0.005207f
C1601 C2S2_Amp_F_I_1.OUT.n69 GND 0.005191f
C1602 C2S2_Amp_F_I_1.OUT.n70 GND 0.004288f
C1603 C2S2_Amp_F_I_1.OUT.n71 GND 0.002959f
C1604 C2S2_Amp_F_I_1.OUT.t51 GND 0.023264f
C1605 C2S2_Amp_F_I_1.OUT.n72 GND 0.04788f
C1606 C2S2_Amp_F_I_1.OUT.n73 GND 0.003289f
C1607 C2S2_Amp_F_I_1.OUT.n74 GND 0.015807f
C1608 C2S2_Amp_F_I_1.OUT.n75 GND 0.358765f
C1609 C2S2_Amp_F_I_1.OUT.n76 GND 0.00528f
C1610 C2S2_Amp_F_I_1.OUT.n77 GND 0.001855f
C1611 C2S2_Amp_F_I_1.OUT.t28 GND 0.023264f
C1612 C2S2_Amp_F_I_1.OUT.n78 GND 0.001964f
C1613 C2S2_Amp_F_I_1.OUT.n79 GND 0.001964f
C1614 C2S2_Amp_F_I_1.OUT.n80 GND 0.001855f
C1615 C2S2_Amp_F_I_1.OUT.n81 GND 0.005207f
C1616 C2S2_Amp_F_I_1.OUT.n82 GND 0.005191f
C1617 C2S2_Amp_F_I_1.OUT.n83 GND 0.004288f
C1618 C2S2_Amp_F_I_1.OUT.n84 GND 0.002959f
C1619 C2S2_Amp_F_I_1.OUT.t64 GND 0.023264f
C1620 C2S2_Amp_F_I_1.OUT.n85 GND 0.04788f
C1621 C2S2_Amp_F_I_1.OUT.n86 GND 0.003289f
C1622 C2S2_Amp_F_I_1.OUT.n87 GND 0.015807f
C1623 C2S2_Amp_F_I_1.OUT.n88 GND 0.18093f
C1624 C2S2_Amp_F_I_1.OUT.n89 GND 0.00528f
C1625 C2S2_Amp_F_I_1.OUT.n90 GND 0.001855f
C1626 C2S2_Amp_F_I_1.OUT.t56 GND 0.023264f
C1627 C2S2_Amp_F_I_1.OUT.n91 GND 0.001964f
C1628 C2S2_Amp_F_I_1.OUT.n92 GND 0.001964f
C1629 C2S2_Amp_F_I_1.OUT.n93 GND 0.001855f
C1630 C2S2_Amp_F_I_1.OUT.n94 GND 0.005207f
C1631 C2S2_Amp_F_I_1.OUT.n95 GND 0.005191f
C1632 C2S2_Amp_F_I_1.OUT.n96 GND 0.004288f
C1633 C2S2_Amp_F_I_1.OUT.n97 GND 0.002959f
C1634 C2S2_Amp_F_I_1.OUT.t47 GND 0.023264f
C1635 C2S2_Amp_F_I_1.OUT.n98 GND 0.04788f
C1636 C2S2_Amp_F_I_1.OUT.n99 GND 0.003289f
C1637 C2S2_Amp_F_I_1.OUT.n100 GND 0.015807f
C1638 C2S2_Amp_F_I_1.OUT.n101 GND 0.178282f
C1639 C2S2_Amp_F_I_1.OUT.n102 GND 0.00528f
C1640 C2S2_Amp_F_I_1.OUT.n103 GND 0.001855f
C1641 C2S2_Amp_F_I_1.OUT.t48 GND 0.023264f
C1642 C2S2_Amp_F_I_1.OUT.n104 GND 0.001964f
C1643 C2S2_Amp_F_I_1.OUT.n105 GND 0.001964f
C1644 C2S2_Amp_F_I_1.OUT.n106 GND 0.001855f
C1645 C2S2_Amp_F_I_1.OUT.n107 GND 0.005207f
C1646 C2S2_Amp_F_I_1.OUT.n108 GND 0.005191f
C1647 C2S2_Amp_F_I_1.OUT.n109 GND 0.004288f
C1648 C2S2_Amp_F_I_1.OUT.n110 GND 0.002959f
C1649 C2S2_Amp_F_I_1.OUT.t37 GND 0.023264f
C1650 C2S2_Amp_F_I_1.OUT.n111 GND 0.04788f
C1651 C2S2_Amp_F_I_1.OUT.n112 GND 0.003289f
C1652 C2S2_Amp_F_I_1.OUT.n113 GND 0.015807f
C1653 C2S2_Amp_F_I_1.OUT.n114 GND 0.178282f
C1654 C2S2_Amp_F_I_1.OUT.n115 GND 0.00528f
C1655 C2S2_Amp_F_I_1.OUT.n116 GND 0.001855f
C1656 C2S2_Amp_F_I_1.OUT.t30 GND 0.023264f
C1657 C2S2_Amp_F_I_1.OUT.n117 GND 0.001964f
C1658 C2S2_Amp_F_I_1.OUT.n118 GND 0.001964f
C1659 C2S2_Amp_F_I_1.OUT.n119 GND 0.001855f
C1660 C2S2_Amp_F_I_1.OUT.n120 GND 0.005207f
C1661 C2S2_Amp_F_I_1.OUT.n121 GND 0.005191f
C1662 C2S2_Amp_F_I_1.OUT.n122 GND 0.004288f
C1663 C2S2_Amp_F_I_1.OUT.n123 GND 0.002959f
C1664 C2S2_Amp_F_I_1.OUT.t58 GND 0.023264f
C1665 C2S2_Amp_F_I_1.OUT.n124 GND 0.04788f
C1666 C2S2_Amp_F_I_1.OUT.n125 GND 0.003289f
C1667 C2S2_Amp_F_I_1.OUT.n126 GND 0.015807f
C1668 C2S2_Amp_F_I_1.OUT.n127 GND 0.178282f
C1669 C2S2_Amp_F_I_1.OUT.n128 GND 0.00528f
C1670 C2S2_Amp_F_I_1.OUT.n129 GND 0.001855f
C1671 C2S2_Amp_F_I_1.OUT.t44 GND 0.023264f
C1672 C2S2_Amp_F_I_1.OUT.n130 GND 0.001964f
C1673 C2S2_Amp_F_I_1.OUT.n131 GND 0.001964f
C1674 C2S2_Amp_F_I_1.OUT.n132 GND 0.001855f
C1675 C2S2_Amp_F_I_1.OUT.n133 GND 0.005207f
C1676 C2S2_Amp_F_I_1.OUT.n134 GND 0.005191f
C1677 C2S2_Amp_F_I_1.OUT.n135 GND 0.004288f
C1678 C2S2_Amp_F_I_1.OUT.n136 GND 0.002959f
C1679 C2S2_Amp_F_I_1.OUT.t38 GND 0.023264f
C1680 C2S2_Amp_F_I_1.OUT.n137 GND 0.04788f
C1681 C2S2_Amp_F_I_1.OUT.n138 GND 0.003289f
C1682 C2S2_Amp_F_I_1.OUT.n139 GND 0.015807f
C1683 C2S2_Amp_F_I_1.OUT.n140 GND 0.178282f
C1684 C2S2_Amp_F_I_1.OUT.n141 GND 0.00528f
C1685 C2S2_Amp_F_I_1.OUT.n142 GND 0.001855f
C1686 C2S2_Amp_F_I_1.OUT.t41 GND 0.023264f
C1687 C2S2_Amp_F_I_1.OUT.n143 GND 0.001964f
C1688 C2S2_Amp_F_I_1.OUT.n144 GND 0.001964f
C1689 C2S2_Amp_F_I_1.OUT.n145 GND 0.001855f
C1690 C2S2_Amp_F_I_1.OUT.n146 GND 0.005207f
C1691 C2S2_Amp_F_I_1.OUT.n147 GND 0.005191f
C1692 C2S2_Amp_F_I_1.OUT.n148 GND 0.004288f
C1693 C2S2_Amp_F_I_1.OUT.n149 GND 0.002959f
C1694 C2S2_Amp_F_I_1.OUT.t31 GND 0.023264f
C1695 C2S2_Amp_F_I_1.OUT.n150 GND 0.04788f
C1696 C2S2_Amp_F_I_1.OUT.n151 GND 0.003289f
C1697 C2S2_Amp_F_I_1.OUT.n152 GND 0.015807f
C1698 C2S2_Amp_F_I_1.OUT.n153 GND 0.18093f
C1699 C2S2_Amp_F_I_1.OUT.n154 GND 0.00528f
C1700 C2S2_Amp_F_I_1.OUT.n155 GND 0.001855f
C1701 C2S2_Amp_F_I_1.OUT.t26 GND 0.023264f
C1702 C2S2_Amp_F_I_1.OUT.n156 GND 0.001964f
C1703 C2S2_Amp_F_I_1.OUT.n157 GND 0.001964f
C1704 C2S2_Amp_F_I_1.OUT.n158 GND 0.001855f
C1705 C2S2_Amp_F_I_1.OUT.n159 GND 0.005207f
C1706 C2S2_Amp_F_I_1.OUT.n160 GND 0.005191f
C1707 C2S2_Amp_F_I_1.OUT.n161 GND 0.004288f
C1708 C2S2_Amp_F_I_1.OUT.n162 GND 0.002959f
C1709 C2S2_Amp_F_I_1.OUT.t62 GND 0.023264f
C1710 C2S2_Amp_F_I_1.OUT.n163 GND 0.04788f
C1711 C2S2_Amp_F_I_1.OUT.n164 GND 0.003289f
C1712 C2S2_Amp_F_I_1.OUT.n165 GND 0.015807f
C1713 C2S2_Amp_F_I_1.OUT.n166 GND 0.178282f
C1714 C2S2_Amp_F_I_1.OUT.n167 GND 0.00528f
C1715 C2S2_Amp_F_I_1.OUT.n168 GND 0.001855f
C1716 C2S2_Amp_F_I_1.OUT.t34 GND 0.023264f
C1717 C2S2_Amp_F_I_1.OUT.n169 GND 0.001964f
C1718 C2S2_Amp_F_I_1.OUT.n170 GND 0.001964f
C1719 C2S2_Amp_F_I_1.OUT.n171 GND 0.001855f
C1720 C2S2_Amp_F_I_1.OUT.n172 GND 0.005207f
C1721 C2S2_Amp_F_I_1.OUT.n173 GND 0.005191f
C1722 C2S2_Amp_F_I_1.OUT.n174 GND 0.004288f
C1723 C2S2_Amp_F_I_1.OUT.n175 GND 0.002959f
C1724 C2S2_Amp_F_I_1.OUT.t29 GND 0.023264f
C1725 C2S2_Amp_F_I_1.OUT.n176 GND 0.04788f
C1726 C2S2_Amp_F_I_1.OUT.n177 GND 0.003289f
C1727 C2S2_Amp_F_I_1.OUT.n178 GND 0.015807f
C1728 C2S2_Amp_F_I_1.OUT.n179 GND 0.178282f
C1729 C2S2_Amp_F_I_1.OUT.n180 GND 0.00528f
C1730 C2S2_Amp_F_I_1.OUT.n181 GND 0.001855f
C1731 C2S2_Amp_F_I_1.OUT.t45 GND 0.023264f
C1732 C2S2_Amp_F_I_1.OUT.n182 GND 0.001964f
C1733 C2S2_Amp_F_I_1.OUT.n183 GND 0.001964f
C1734 C2S2_Amp_F_I_1.OUT.n184 GND 0.001855f
C1735 C2S2_Amp_F_I_1.OUT.n185 GND 0.005207f
C1736 C2S2_Amp_F_I_1.OUT.n186 GND 0.005191f
C1737 C2S2_Amp_F_I_1.OUT.n187 GND 0.004288f
C1738 C2S2_Amp_F_I_1.OUT.n188 GND 0.002959f
C1739 C2S2_Amp_F_I_1.OUT.t39 GND 0.023264f
C1740 C2S2_Amp_F_I_1.OUT.n189 GND 0.04788f
C1741 C2S2_Amp_F_I_1.OUT.n190 GND 0.003289f
C1742 C2S2_Amp_F_I_1.OUT.n191 GND 0.015807f
C1743 C2S2_Amp_F_I_1.OUT.n192 GND 0.18093f
C1744 C2S2_Amp_F_I_1.OUT.n193 GND 0.00528f
C1745 C2S2_Amp_F_I_1.OUT.n194 GND 0.001855f
C1746 C2S2_Amp_F_I_1.OUT.t59 GND 0.023264f
C1747 C2S2_Amp_F_I_1.OUT.n195 GND 0.001964f
C1748 C2S2_Amp_F_I_1.OUT.n196 GND 0.001964f
C1749 C2S2_Amp_F_I_1.OUT.n197 GND 0.001855f
C1750 C2S2_Amp_F_I_1.OUT.n198 GND 0.005207f
C1751 C2S2_Amp_F_I_1.OUT.n199 GND 0.005191f
C1752 C2S2_Amp_F_I_1.OUT.n200 GND 0.004288f
C1753 C2S2_Amp_F_I_1.OUT.n201 GND 0.002959f
C1754 C2S2_Amp_F_I_1.OUT.t54 GND 0.023264f
C1755 C2S2_Amp_F_I_1.OUT.n202 GND 0.04788f
C1756 C2S2_Amp_F_I_1.OUT.n203 GND 0.003289f
C1757 C2S2_Amp_F_I_1.OUT.n204 GND 0.015807f
C1758 C2S2_Amp_F_I_1.OUT.n205 GND 0.178282f
C1759 C2S2_Amp_F_I_1.OUT.n206 GND 0.00528f
C1760 C2S2_Amp_F_I_1.OUT.n207 GND 0.001855f
C1761 C2S2_Amp_F_I_1.OUT.t27 GND 0.023264f
C1762 C2S2_Amp_F_I_1.OUT.n208 GND 0.001964f
C1763 C2S2_Amp_F_I_1.OUT.n209 GND 0.001964f
C1764 C2S2_Amp_F_I_1.OUT.n210 GND 0.001855f
C1765 C2S2_Amp_F_I_1.OUT.n211 GND 0.005207f
C1766 C2S2_Amp_F_I_1.OUT.n212 GND 0.005191f
C1767 C2S2_Amp_F_I_1.OUT.n213 GND 0.004288f
C1768 C2S2_Amp_F_I_1.OUT.n214 GND 0.002959f
C1769 C2S2_Amp_F_I_1.OUT.t25 GND 0.023264f
C1770 C2S2_Amp_F_I_1.OUT.n215 GND 0.04788f
C1771 C2S2_Amp_F_I_1.OUT.n216 GND 0.003289f
C1772 C2S2_Amp_F_I_1.OUT.n217 GND 0.015807f
C1773 C2S2_Amp_F_I_1.OUT.n218 GND 0.178282f
C1774 C2S2_Amp_F_I_1.OUT.n219 GND 0.00528f
C1775 C2S2_Amp_F_I_1.OUT.n220 GND 0.001855f
C1776 C2S2_Amp_F_I_1.OUT.t32 GND 0.023264f
C1777 C2S2_Amp_F_I_1.OUT.n221 GND 0.001964f
C1778 C2S2_Amp_F_I_1.OUT.n222 GND 0.001964f
C1779 C2S2_Amp_F_I_1.OUT.n223 GND 0.001855f
C1780 C2S2_Amp_F_I_1.OUT.n224 GND 0.005207f
C1781 C2S2_Amp_F_I_1.OUT.n225 GND 0.005191f
C1782 C2S2_Amp_F_I_1.OUT.n226 GND 0.004288f
C1783 C2S2_Amp_F_I_1.OUT.n227 GND 0.002959f
C1784 C2S2_Amp_F_I_1.OUT.t49 GND 0.023264f
C1785 C2S2_Amp_F_I_1.OUT.n228 GND 0.04788f
C1786 C2S2_Amp_F_I_1.OUT.n229 GND 0.003289f
C1787 C2S2_Amp_F_I_1.OUT.n230 GND 0.015807f
C1788 C2S2_Amp_F_I_1.OUT.n231 GND 0.178282f
C1789 C2S2_Amp_F_I_1.OUT.n232 GND 0.00528f
C1790 C2S2_Amp_F_I_1.OUT.n233 GND 0.001855f
C1791 C2S2_Amp_F_I_1.OUT.t52 GND 0.023264f
C1792 C2S2_Amp_F_I_1.OUT.n234 GND 0.001964f
C1793 C2S2_Amp_F_I_1.OUT.n235 GND 0.001964f
C1794 C2S2_Amp_F_I_1.OUT.n236 GND 0.001855f
C1795 C2S2_Amp_F_I_1.OUT.n237 GND 0.005207f
C1796 C2S2_Amp_F_I_1.OUT.n238 GND 0.005191f
C1797 C2S2_Amp_F_I_1.OUT.n239 GND 0.004288f
C1798 C2S2_Amp_F_I_1.OUT.n240 GND 0.002959f
C1799 C2S2_Amp_F_I_1.OUT.t43 GND 0.023264f
C1800 C2S2_Amp_F_I_1.OUT.n241 GND 0.04788f
C1801 C2S2_Amp_F_I_1.OUT.n242 GND 0.003289f
C1802 C2S2_Amp_F_I_1.OUT.n243 GND 0.015807f
C1803 C2S2_Amp_F_I_1.OUT.n244 GND 0.178282f
C1804 C2S2_Amp_F_I_1.OUT.n245 GND 0.00528f
C1805 C2S2_Amp_F_I_1.OUT.n246 GND 0.001855f
C1806 C2S2_Amp_F_I_1.OUT.t33 GND 0.023264f
C1807 C2S2_Amp_F_I_1.OUT.n247 GND 0.001964f
C1808 C2S2_Amp_F_I_1.OUT.n248 GND 0.001964f
C1809 C2S2_Amp_F_I_1.OUT.n249 GND 0.001855f
C1810 C2S2_Amp_F_I_1.OUT.n250 GND 0.005207f
C1811 C2S2_Amp_F_I_1.OUT.n251 GND 0.005191f
C1812 C2S2_Amp_F_I_1.OUT.n252 GND 0.004288f
C1813 C2S2_Amp_F_I_1.OUT.n253 GND 0.002959f
C1814 C2S2_Amp_F_I_1.OUT.t57 GND 0.023264f
C1815 C2S2_Amp_F_I_1.OUT.n254 GND 0.04788f
C1816 C2S2_Amp_F_I_1.OUT.n255 GND 0.003289f
C1817 C2S2_Amp_F_I_1.OUT.n256 GND 0.015807f
C1818 C2S2_Amp_F_I_1.OUT.n257 GND 0.18093f
C1819 C2S2_Amp_F_I_1.OUT.n258 GND 0.00528f
C1820 C2S2_Amp_F_I_1.OUT.n259 GND 0.001855f
C1821 C2S2_Amp_F_I_1.OUT.t46 GND 0.023264f
C1822 C2S2_Amp_F_I_1.OUT.n260 GND 0.001964f
C1823 C2S2_Amp_F_I_1.OUT.n261 GND 0.001964f
C1824 C2S2_Amp_F_I_1.OUT.n262 GND 0.001855f
C1825 C2S2_Amp_F_I_1.OUT.n263 GND 0.005207f
C1826 C2S2_Amp_F_I_1.OUT.n264 GND 0.005191f
C1827 C2S2_Amp_F_I_1.OUT.n265 GND 0.004288f
C1828 C2S2_Amp_F_I_1.OUT.n266 GND 0.002959f
C1829 C2S2_Amp_F_I_1.OUT.t36 GND 0.023264f
C1830 C2S2_Amp_F_I_1.OUT.n267 GND 0.04788f
C1831 C2S2_Amp_F_I_1.OUT.n268 GND 0.003289f
C1832 C2S2_Amp_F_I_1.OUT.n269 GND 0.015807f
C1833 C2S2_Amp_F_I_1.OUT.n270 GND 0.178282f
C1834 C2S2_Amp_F_I_1.OUT.n271 GND 0.00528f
C1835 C2S2_Amp_F_I_1.OUT.n272 GND 0.001855f
C1836 C2S2_Amp_F_I_1.OUT.t60 GND 0.023264f
C1837 C2S2_Amp_F_I_1.OUT.n273 GND 0.001964f
C1838 C2S2_Amp_F_I_1.OUT.n274 GND 0.001964f
C1839 C2S2_Amp_F_I_1.OUT.n275 GND 0.001855f
C1840 C2S2_Amp_F_I_1.OUT.n276 GND 0.005207f
C1841 C2S2_Amp_F_I_1.OUT.n277 GND 0.005191f
C1842 C2S2_Amp_F_I_1.OUT.n278 GND 0.004288f
C1843 C2S2_Amp_F_I_1.OUT.n279 GND 0.002959f
C1844 C2S2_Amp_F_I_1.OUT.t55 GND 0.023264f
C1845 C2S2_Amp_F_I_1.OUT.n280 GND 0.04788f
C1846 C2S2_Amp_F_I_1.OUT.n281 GND 0.003289f
C1847 C2S2_Amp_F_I_1.OUT.n282 GND 0.015807f
C1848 C2S2_Amp_F_I_1.OUT.n283 GND 0.178282f
C1849 C2S2_Amp_F_I_1.OUT.n284 GND 0.00528f
C1850 C2S2_Amp_F_I_1.OUT.n285 GND 0.001855f
C1851 C2S2_Amp_F_I_1.OUT.t40 GND 0.023264f
C1852 C2S2_Amp_F_I_1.OUT.n286 GND 0.001964f
C1853 C2S2_Amp_F_I_1.OUT.n287 GND 0.001964f
C1854 C2S2_Amp_F_I_1.OUT.n288 GND 0.001855f
C1855 C2S2_Amp_F_I_1.OUT.n289 GND 0.005207f
C1856 C2S2_Amp_F_I_1.OUT.n290 GND 0.005191f
C1857 C2S2_Amp_F_I_1.OUT.n291 GND 0.004288f
C1858 C2S2_Amp_F_I_1.OUT.n292 GND 0.002959f
C1859 C2S2_Amp_F_I_1.OUT.t35 GND 0.023264f
C1860 C2S2_Amp_F_I_1.OUT.n293 GND 0.04788f
C1861 C2S2_Amp_F_I_1.OUT.n294 GND 0.003289f
C1862 C2S2_Amp_F_I_1.OUT.n295 GND 0.015807f
C1863 C2S2_Amp_F_I_1.OUT.n296 GND 0.358684f
C1864 C2S2_Amp_F_I_1.OUT.n297 GND 0.002959f
C1865 C2S2_Amp_F_I_1.OUT.n298 GND 0.005207f
C1866 C2S2_Amp_F_I_1.OUT.n299 GND 0.001855f
C1867 C2S2_Amp_F_I_1.OUT.t53 GND 0.023264f
C1868 C2S2_Amp_F_I_1.OUT.n300 GND 0.003289f
C1869 C2S2_Amp_F_I_1.OUT.n301 GND 0.00528f
C1870 C2S2_Amp_F_I_1.OUT.n302 GND 0.001855f
C1871 C2S2_Amp_F_I_1.OUT.n303 GND 0.001964f
C1872 C2S2_Amp_F_I_1.OUT.t50 GND 0.023264f
C1873 C2S2_Amp_F_I_1.OUT.n304 GND 0.04788f
C1874 C2S2_Amp_F_I_1.OUT.n305 GND 0.001964f
C1875 C2S2_Amp_F_I_1.OUT.n306 GND 0.004288f
C1876 C2S2_Amp_F_I_1.OUT.n307 GND 0.005191f
C1877 C2S2_Amp_F_I_1.OUT.n308 GND 0.09286f
C1878 C2S2_Amp_F_I_1.OUT.n309 GND 0.038489f
C1879 C2S2_Amp_F_I_1.OUT.n310 GND 0.063616f
C1880 C2S2_Amp_F_I_1.OUT.n311 GND 0.020055f
C1881 C2S2_Amp_F_I_1.OUT.t0 GND 1.19448f
C1882 C2S2_Amp_F_I_1.OUT.n312 GND 0.809395f
C1883 C2S2_Amp_F_I_1.OUT.t4 GND 18.600801f
C1884 C2S2_Amp_F_I_1.OUT.t8 GND 16.953001f
C1885 C2S2_Amp_F_I_1.OUT.n313 GND 1.88894f
C1886 C2S2_Amp_F_I_1.OUT.t6 GND 16.953001f
C1887 C2S2_Amp_F_I_1.OUT.n314 GND 1.76835f
C1888 C2S2_Amp_F_I_1.OUT.t2 GND 16.953001f
C1889 C2S2_Amp_F_I_1.OUT.n315 GND 2.22011f
C1890 C2S2_Amp_F_I_1.OUT.t11 GND 18.600801f
C1891 C2S2_Amp_F_I_1.OUT.t1 GND 16.953001f
C1892 C2S2_Amp_F_I_1.OUT.n316 GND 1.88894f
C1893 C2S2_Amp_F_I_1.OUT.t9 GND 16.953001f
C1894 C2S2_Amp_F_I_1.OUT.n317 GND 1.76835f
C1895 C2S2_Amp_F_I_1.OUT.t3 GND 16.953001f
C1896 C2S2_Amp_F_I_1.OUT.n318 GND 1.71005f
C1897 C2S2_Amp_F_I_1.OUT.n319 GND 3.55065f
C1898 C2S2_Amp_F_I_1.OUT.t7 GND 18.600801f
C1899 C2S2_Amp_F_I_1.OUT.t5 GND 16.953001f
C1900 C2S2_Amp_F_I_1.OUT.n320 GND 1.88894f
C1901 C2S2_Amp_F_I_1.OUT.t12 GND 16.953001f
C1902 C2S2_Amp_F_I_1.OUT.n321 GND 1.76835f
C1903 C2S2_Amp_F_I_1.OUT.t10 GND 16.953001f
C1904 C2S2_Amp_F_I_1.OUT.n322 GND 2.32719f
C1905 C2S2_Amp_F_I_1.OUT.n323 GND 4.41566f
C1906 C2S2_Amp_F_I_1.OUT.n324 GND 2.65543f
C1907 C2S2_Amp_F_I_1.OUT.n325 GND 0.301259f
C1908 C2S2_Amp_F_I_1.OUT.n326 GND 11.8481f
C1909 C2S2_Amp_F_I_1.OUT.n327 GND 0.015806f
C1910 C2S2_Amp_F_I_1.OUT.n328 GND 0.015806f
C1911 C2S2_Amp_F_I_1.OUT.n329 GND 0.015806f
C1912 C2S2_Amp_F_I_1.OUT.n330 GND 0.015806f
C1913 C2S2_Amp_F_I_1.OUT.n331 GND 0.015806f
C1914 C2S2_Amp_F_I_1.OUT.n332 GND 0.015806f
C1915 C2S2_Amp_F_I_1.OUT.n333 GND 0.005278f
C1916 C2S2_Amp_F_I_1.OUT.t18 GND 0.023264f
C1917 C2S2_Amp_F_I_1.OUT.t14 GND 0.023264f
C1918 C2S2_Amp_F_I_1.OUT.n334 GND 0.050651f
C1919 C2S2_Amp_F_I_1.OUT.n335 GND 0.001964f
C1920 C2S2_Amp_F_I_1.OUT.n336 GND 0.003288f
C1921 C2S2_Amp_F_I_1.OUT.n337 GND 0.001855f
C1922 C2S2_Amp_F_I_1.OUT.n338 GND 0.005268f
C1923 C2S2_Amp_F_I_1.OUT.n339 GND 0.005081f
C1924 C2S2_Amp_F_I_1.OUT.n340 GND 0.001855f
C1925 C2S2_Amp_F_I_1.OUT.n341 GND 0.001964f
C1926 C2S2_Amp_F_I_1.OUT.n342 GND 0.004222f
C1927 C2S2_Amp_F_I_1.OUT.n343 GND 0.006302f
C1928 C2S2_Amp_F_I_1.OUT.n344 GND 0.090385f
C1929 C2S2_Amp_F_I_1.OUT.n345 GND 0.342015f
C1930 C2S2_Amp_F_I_1.OUT.n346 GND 0.005278f
C1931 C2S2_Amp_F_I_1.OUT.t16 GND 0.023264f
C1932 C2S2_Amp_F_I_1.OUT.t15 GND 0.023264f
C1933 C2S2_Amp_F_I_1.OUT.n347 GND 0.050651f
C1934 C2S2_Amp_F_I_1.OUT.n348 GND 0.001964f
C1935 C2S2_Amp_F_I_1.OUT.n349 GND 0.003288f
C1936 C2S2_Amp_F_I_1.OUT.n350 GND 0.001855f
C1937 C2S2_Amp_F_I_1.OUT.n351 GND 0.005268f
C1938 C2S2_Amp_F_I_1.OUT.n352 GND 0.005081f
C1939 C2S2_Amp_F_I_1.OUT.n353 GND 0.001855f
C1940 C2S2_Amp_F_I_1.OUT.n354 GND 0.001964f
C1941 C2S2_Amp_F_I_1.OUT.n355 GND 0.004222f
C1942 C2S2_Amp_F_I_1.OUT.n356 GND 0.006302f
C1943 C2S2_Amp_F_I_1.OUT.n357 GND 0.090385f
C1944 C2S2_Amp_F_I_1.OUT.n358 GND 0.342015f
C1945 C2S2_Amp_F_I_1.OUT.n359 GND 0.005278f
C1946 C2S2_Amp_F_I_1.OUT.t23 GND 0.023264f
C1947 C2S2_Amp_F_I_1.OUT.t19 GND 0.023264f
C1948 C2S2_Amp_F_I_1.OUT.n360 GND 0.050651f
C1949 C2S2_Amp_F_I_1.OUT.n361 GND 0.001964f
C1950 C2S2_Amp_F_I_1.OUT.n362 GND 0.003288f
C1951 C2S2_Amp_F_I_1.OUT.n363 GND 0.001855f
C1952 C2S2_Amp_F_I_1.OUT.n364 GND 0.005268f
C1953 C2S2_Amp_F_I_1.OUT.n365 GND 0.005081f
C1954 C2S2_Amp_F_I_1.OUT.n366 GND 0.001855f
C1955 C2S2_Amp_F_I_1.OUT.n367 GND 0.001964f
C1956 C2S2_Amp_F_I_1.OUT.n368 GND 0.004222f
C1957 C2S2_Amp_F_I_1.OUT.n369 GND 0.006302f
C1958 C2S2_Amp_F_I_1.OUT.n370 GND 0.090385f
C1959 C2S2_Amp_F_I_1.OUT.n371 GND 0.342015f
C1960 C2S2_Amp_F_I_1.OUT.n372 GND 0.005278f
C1961 C2S2_Amp_F_I_1.OUT.t24 GND 0.023264f
C1962 C2S2_Amp_F_I_1.OUT.t21 GND 0.023264f
C1963 C2S2_Amp_F_I_1.OUT.n373 GND 0.050651f
C1964 C2S2_Amp_F_I_1.OUT.n374 GND 0.001964f
C1965 C2S2_Amp_F_I_1.OUT.n375 GND 0.003288f
C1966 C2S2_Amp_F_I_1.OUT.n376 GND 0.001855f
C1967 C2S2_Amp_F_I_1.OUT.n377 GND 0.005268f
C1968 C2S2_Amp_F_I_1.OUT.n378 GND 0.005081f
C1969 C2S2_Amp_F_I_1.OUT.n379 GND 0.001855f
C1970 C2S2_Amp_F_I_1.OUT.n380 GND 0.001964f
C1971 C2S2_Amp_F_I_1.OUT.n381 GND 0.004222f
C1972 C2S2_Amp_F_I_1.OUT.n382 GND 0.006302f
C1973 C2S2_Amp_F_I_1.OUT.n383 GND 0.090385f
C1974 C2S2_Amp_F_I_1.OUT.n384 GND 0.342015f
C1975 C2S2_Amp_F_I_1.OUT.n385 GND 0.005278f
C1976 C2S2_Amp_F_I_1.OUT.t22 GND 0.023264f
C1977 C2S2_Amp_F_I_1.OUT.t13 GND 0.023264f
C1978 C2S2_Amp_F_I_1.OUT.n386 GND 0.050651f
C1979 C2S2_Amp_F_I_1.OUT.n387 GND 0.001964f
C1980 C2S2_Amp_F_I_1.OUT.n388 GND 0.003288f
C1981 C2S2_Amp_F_I_1.OUT.n389 GND 0.001855f
C1982 C2S2_Amp_F_I_1.OUT.n390 GND 0.005268f
C1983 C2S2_Amp_F_I_1.OUT.n391 GND 0.005081f
C1984 C2S2_Amp_F_I_1.OUT.n392 GND 0.001855f
C1985 C2S2_Amp_F_I_1.OUT.n393 GND 0.001964f
C1986 C2S2_Amp_F_I_1.OUT.n394 GND 0.004222f
C1987 C2S2_Amp_F_I_1.OUT.n395 GND 0.006302f
C1988 C2S2_Amp_F_I_1.OUT.n396 GND 0.090385f
C1989 C2S2_Amp_F_I_1.OUT.n397 GND 0.345224f
C1990 C2S2_Amp_F_I_1.OUT.n398 GND 0.005278f
C1991 C2S2_Amp_F_I_1.OUT.n399 GND 0.005314f
C1992 C2S2_Amp_F_I_1.OUT.n400 GND 0.001964f
C1993 C2S2_Amp_F_I_1.OUT.n401 GND 0.001855f
C1994 C2S2_Amp_F_I_1.OUT.n402 GND 0.011191f
C1995 C2S2_Amp_F_I_1.OUT.n403 GND 0.001964f
C1996 C2S2_Amp_F_I_1.OUT.n404 GND 0.006986f
C1997 C2S2_Amp_F_I_1.OUT.n405 GND 0.001855f
C1998 C2S2_Amp_F_I_1.OUT.n406 GND 0.005268f
C1999 C2S2_Amp_F_I_1.OUT.n407 GND 0.005081f
C2000 C2S2_Amp_F_I_1.OUT.n408 GND 0.001855f
C2001 C2S2_Amp_F_I_1.OUT.n409 GND 0.001855f
C2002 C2S2_Amp_F_I_1.OUT.n410 GND 0.001964f
C2003 C2S2_Amp_F_I_1.OUT.n411 GND 0.006328f
C2004 C2S2_Amp_F_I_1.OUT.n412 GND 0.006328f
C2005 C2S2_Amp_F_I_1.OUT.n413 GND 0.004746f
C2006 C2S2_Amp_F_I_1.OUT.n414 GND 0.002302f
C2007 C2S2_Amp_F_I_1.OUT.t17 GND 0.009083f
C2008 C2S2_Amp_F_I_1.OUT.n415 GND 0.015035f
C2009 C2S2_Amp_F_I_1.OUT.n416 GND 0.093309f
C2010 C2S2_Amp_F_I_1.OUT.n417 GND 0.001855f
C2011 C2S2_Amp_F_I_1.OUT.n418 GND 0.001964f
C2012 C2S2_Amp_F_I_1.OUT.n419 GND 0.006328f
C2013 C2S2_Amp_F_I_1.OUT.n420 GND 0.006328f
C2014 C2S2_Amp_F_I_1.OUT.n421 GND 0.001964f
C2015 C2S2_Amp_F_I_1.OUT.n422 GND 0.001855f
C2016 C2S2_Amp_F_I_1.OUT.n423 GND 0.005122f
C2017 C2S2_Amp_F_I_1.OUT.n424 GND 0.009666f
C2018 C2S2_Amp_F_I_1.OUT.n425 GND 1.03451f
C2019 C2S2_Amp_F_I_1.OUT.n426 GND 21.112902f
C2020 C2S2_Amp_F_I_1.OUT.n427 GND 1.15792f
C2021 C2S2_Amp_F_I_1.OUT.n428 GND 6.29052f
C2022 C2S2_Amp_F_I_1.OUT.t65 GND 16.4295f
C2023 C2S2_Amp_F_I_1.OUT.n429 GND 14.5703f
C2024 C2S2_Amp_F_I_1.OUT.t66 GND 16.4295f
C2025 C2S2_Amp_F_I_1.OUT.n430 GND 14.542099f
C2026 C2S2_Amp_F_I_1.OUT.t67 GND 30.1756f
C2027 C2S2_Amp_F_I_1.OUT.n431 GND 6.28086f
C2028 C2S2_Amp_F_I_1.OUT.n432 GND 1.15879f
C2029 C2S2_Amp_F_I_1.OUT.n433 GND 11.395901f
C2030 a_187922_n20028.n0 GND 4.26146f
C2031 a_187922_n20028.n1 GND 4.4951f
C2032 a_187922_n20028.n2 GND 0.038056f
C2033 a_187922_n20028.n3 GND 0.038013f
C2034 a_187922_n20028.n4 GND 0.890262f
C2035 a_187922_n20028.n5 GND 1.11609f
C2036 a_187922_n20028.n6 GND 0.193483f
C2037 a_187922_n20028.n7 GND 1.11566f
C2038 a_187922_n20028.n8 GND 0.179668f
C2039 a_187922_n20028.n9 GND 0.004329f
C2040 a_187922_n20028.n10 GND 0.179668f
C2041 a_187922_n20028.n11 GND 0.004329f
C2042 a_187922_n20028.n12 GND 0.179668f
C2043 a_187922_n20028.n13 GND 0.004329f
C2044 a_187922_n20028.n14 GND 0.17961f
C2045 a_187922_n20028.n15 GND 0.00436f
C2046 a_187922_n20028.n16 GND 0.17961f
C2047 a_187922_n20028.n17 GND 0.00436f
C2048 a_187922_n20028.n18 GND 0.17961f
C2049 a_187922_n20028.n19 GND 0.00436f
C2050 a_187922_n20028.n20 GND 0.826379f
C2051 a_187922_n20028.n21 GND 0.825949f
C2052 a_187922_n20028.n22 GND 0.045044f
C2053 a_187922_n20028.n23 GND 0.00707f
C2054 a_187922_n20028.n24 GND 0.045044f
C2055 a_187922_n20028.n25 GND 0.00707f
C2056 a_187922_n20028.n26 GND 0.045044f
C2057 a_187922_n20028.n27 GND 0.00707f
C2058 a_187922_n20028.n28 GND 0.050086f
C2059 a_187922_n20028.n29 GND 0.021014f
C2060 a_187922_n20028.n30 GND 0.045069f
C2061 a_187922_n20028.n31 GND 0.007071f
C2062 a_187922_n20028.n32 GND 0.045069f
C2063 a_187922_n20028.n33 GND 0.007071f
C2064 a_187922_n20028.n34 GND 0.045069f
C2065 a_187922_n20028.n35 GND 0.007071f
C2066 a_187922_n20028.n36 GND 0.045069f
C2067 a_187922_n20028.n37 GND 0.007071f
C2068 a_187922_n20028.n38 GND 0.045069f
C2069 a_187922_n20028.n39 GND 0.007071f
C2070 a_187922_n20028.n40 GND 0.021015f
C2071 a_187922_n20028.n41 GND 0.041843f
C2072 a_187922_n20028.n42 GND 0.041843f
C2073 a_187922_n20028.n43 GND 0.021015f
C2074 a_187922_n20028.n44 GND 0.008904f
C2075 a_187922_n20028.n45 GND 0.007071f
C2076 a_187922_n20028.n46 GND 0.045069f
C2077 a_187922_n20028.n47 GND 0.050135f
C2078 a_187922_n20028.n48 GND 0.021016f
C2079 a_187922_n20028.n49 GND 0.045092f
C2080 a_187922_n20028.n50 GND 0.007071f
C2081 a_187922_n20028.n51 GND 0.045092f
C2082 a_187922_n20028.n52 GND 0.007071f
C2083 a_187922_n20028.n53 GND 0.045092f
C2084 a_187922_n20028.n54 GND 0.007071f
C2085 a_187922_n20028.n55 GND 0.193483f
C2086 a_187922_n20028.n56 GND 0.005875f
C2087 a_187922_n20028.n57 GND 0.193483f
C2088 a_187922_n20028.n58 GND 0.005875f
C2089 a_187922_n20028.n59 GND 0.193483f
C2090 a_187922_n20028.n60 GND 0.005875f
C2091 a_187922_n20028.n61 GND 0.193483f
C2092 a_187922_n20028.n62 GND 0.005875f
C2093 a_187922_n20028.n63 GND 0.193483f
C2094 a_187922_n20028.n64 GND 0.005875f
C2095 a_187922_n20028.n65 GND 0.009641f
C2096 a_187922_n20028.n66 GND 0.021086f
C2097 a_187922_n20028.n67 GND 0.021086f
C2098 a_187922_n20028.n68 GND 0.005875f
C2099 a_187922_n20028.t10 GND 0.044142f
C2100 a_187922_n20028.t13 GND 0.044142f
C2101 a_187922_n20028.t8 GND 0.044142f
C2102 a_187922_n20028.n69 GND 0.097902f
C2103 a_187922_n20028.n70 GND 0.009641f
C2104 a_187922_n20028.n71 GND 0.008904f
C2105 a_187922_n20028.t26 GND 0.044142f
C2106 a_187922_n20028.n72 GND 0.003726f
C2107 a_187922_n20028.n73 GND 0.004616f
C2108 a_187922_n20028.n74 GND 0.00993f
C2109 a_187922_n20028.n75 GND 0.008016f
C2110 a_187922_n20028.n76 GND 0.010083f
C2111 a_187922_n20028.t5 GND 0.044142f
C2112 a_187922_n20028.n77 GND 0.095491f
C2113 a_187922_n20028.t3 GND 0.044142f
C2114 a_187922_n20028.n78 GND 0.003726f
C2115 a_187922_n20028.n79 GND 0.004616f
C2116 a_187922_n20028.n80 GND 0.00993f
C2117 a_187922_n20028.n81 GND 0.008016f
C2118 a_187922_n20028.n82 GND 0.010083f
C2119 a_187922_n20028.t6 GND 0.044142f
C2120 a_187922_n20028.n83 GND 0.095491f
C2121 a_187922_n20028.t25 GND 0.044142f
C2122 a_187922_n20028.n84 GND 0.003726f
C2123 a_187922_n20028.n85 GND 0.004616f
C2124 a_187922_n20028.n86 GND 0.00993f
C2125 a_187922_n20028.n87 GND 0.008016f
C2126 a_187922_n20028.n88 GND 0.010083f
C2127 a_187922_n20028.t23 GND 0.044142f
C2128 a_187922_n20028.n89 GND 0.095491f
C2129 a_187922_n20028.n90 GND 0.021745f
C2130 a_187922_n20028.n91 GND 0.003726f
C2131 a_187922_n20028.n92 GND 0.003519f
C2132 a_187922_n20028.n93 GND 0.012007f
C2133 a_187922_n20028.n94 GND 0.003726f
C2134 a_187922_n20028.n95 GND 0.028528f
C2135 a_187922_n20028.t24 GND 0.017234f
C2136 a_187922_n20028.n96 GND 0.009005f
C2137 a_187922_n20028.n97 GND 0.004368f
C2138 a_187922_n20028.n98 GND 0.003519f
C2139 a_187922_n20028.n99 GND 0.176844f
C2140 a_187922_n20028.n100 GND 0.003519f
C2141 a_187922_n20028.n101 GND 0.003726f
C2142 a_187922_n20028.n102 GND 0.012007f
C2143 a_187922_n20028.n103 GND 0.012007f
C2144 a_187922_n20028.n104 GND 0.003726f
C2145 a_187922_n20028.n105 GND 0.003519f
C2146 a_187922_n20028.n106 GND 0.010083f
C2147 a_187922_n20028.n107 GND 0.00993f
C2148 a_187922_n20028.n108 GND 0.004377f
C2149 a_187922_n20028.n109 GND 0.010083f
C2150 a_187922_n20028.n110 GND 0.003726f
C2151 a_187922_n20028.n111 GND 0.003519f
C2152 a_187922_n20028.n112 GND 0.009641f
C2153 a_187922_n20028.n113 GND 0.004377f
C2154 a_187922_n20028.n114 GND 0.003519f
C2155 a_187922_n20028.n115 GND 0.003726f
C2156 a_187922_n20028.n116 GND 0.021745f
C2157 a_187922_n20028.n117 GND 0.012007f
C2158 a_187922_n20028.n118 GND 0.009005f
C2159 a_187922_n20028.n119 GND 0.004368f
C2160 a_187922_n20028.t14 GND 0.017234f
C2161 a_187922_n20028.n120 GND 0.028528f
C2162 a_187922_n20028.n121 GND 0.177047f
C2163 a_187922_n20028.n122 GND 0.003519f
C2164 a_187922_n20028.n123 GND 0.003726f
C2165 a_187922_n20028.n124 GND 0.012007f
C2166 a_187922_n20028.n125 GND 0.012007f
C2167 a_187922_n20028.n126 GND 0.003726f
C2168 a_187922_n20028.n127 GND 0.003519f
C2169 a_187922_n20028.n128 GND 0.009718f
C2170 a_187922_n20028.t19 GND 0.044142f
C2171 a_187922_n20028.t16 GND 0.044142f
C2172 a_187922_n20028.n129 GND 0.097902f
C2173 a_187922_n20028.n130 GND 0.009641f
C2174 a_187922_n20028.n131 GND 0.008904f
C2175 a_187922_n20028.t11 GND 0.044142f
C2176 a_187922_n20028.t9 GND 0.044142f
C2177 a_187922_n20028.n132 GND 0.097902f
C2178 a_187922_n20028.n133 GND 0.009641f
C2179 a_187922_n20028.n134 GND 0.008904f
C2180 a_187922_n20028.t12 GND 0.044142f
C2181 a_187922_n20028.t17 GND 0.044142f
C2182 a_187922_n20028.n135 GND 0.097902f
C2183 a_187922_n20028.n136 GND 0.009641f
C2184 a_187922_n20028.n137 GND 0.008904f
C2185 a_187922_n20028.n138 GND 1.30222f
C2186 a_187922_n20028.t2 GND 0.044142f
C2187 a_187922_n20028.t1 GND 0.044142f
C2188 a_187922_n20028.n139 GND 0.095463f
C2189 a_187922_n20028.n140 GND 0.003726f
C2190 a_187922_n20028.n141 GND 0.004616f
C2191 a_187922_n20028.n142 GND 0.00988f
C2192 a_187922_n20028.n143 GND 0.010083f
C2193 a_187922_n20028.n144 GND 0.008016f
C2194 a_187922_n20028.t22 GND 0.044142f
C2195 a_187922_n20028.t7 GND 0.044142f
C2196 a_187922_n20028.n145 GND 0.095463f
C2197 a_187922_n20028.n146 GND 0.003726f
C2198 a_187922_n20028.n147 GND 0.004616f
C2199 a_187922_n20028.n148 GND 0.00988f
C2200 a_187922_n20028.n149 GND 0.010083f
C2201 a_187922_n20028.n150 GND 0.008016f
C2202 a_187922_n20028.t0 GND 0.044142f
C2203 a_187922_n20028.t27 GND 0.044142f
C2204 a_187922_n20028.n151 GND 0.095463f
C2205 a_187922_n20028.n152 GND 0.003726f
C2206 a_187922_n20028.n153 GND 0.004616f
C2207 a_187922_n20028.n154 GND 0.00988f
C2208 a_187922_n20028.n155 GND 0.010083f
C2209 a_187922_n20028.n156 GND 0.008016f
C2210 a_187922_n20028.n157 GND 0.176801f
C2211 a_187922_n20028.n158 GND 0.003726f
C2212 a_187922_n20028.n159 GND 0.003519f
C2213 a_187922_n20028.n160 GND 0.021745f
C2214 a_187922_n20028.n161 GND 0.003726f
C2215 a_187922_n20028.n162 GND 0.004377f
C2216 a_187922_n20028.n163 GND 0.00988f
C2217 a_187922_n20028.n164 GND 0.010083f
C2218 a_187922_n20028.n165 GND 0.003519f
C2219 a_187922_n20028.n166 GND 0.003519f
C2220 a_187922_n20028.n167 GND 0.003726f
C2221 a_187922_n20028.n168 GND 0.012007f
C2222 a_187922_n20028.n169 GND 0.012007f
C2223 a_187922_n20028.t4 GND 0.017234f
C2224 a_187922_n20028.n170 GND 0.028528f
C2225 a_187922_n20028.n171 GND 0.004368f
C2226 a_187922_n20028.n172 GND 0.009005f
C2227 a_187922_n20028.n173 GND 0.012007f
C2228 a_187922_n20028.n174 GND 0.003726f
C2229 a_187922_n20028.n175 GND 0.003519f
C2230 a_187922_n20028.n176 GND 1.29828f
C2231 a_187922_n20028.n177 GND 0.004377f
C2232 a_187922_n20028.n178 GND 0.012007f
C2233 a_187922_n20028.n179 GND 0.003726f
C2234 a_187922_n20028.n180 GND 0.177047f
C2235 a_187922_n20028.n181 GND 0.003519f
C2236 a_187922_n20028.n182 GND 0.012007f
C2237 a_187922_n20028.t15 GND 0.017234f
C2238 a_187922_n20028.n183 GND 0.028528f
C2239 a_187922_n20028.n184 GND 0.004368f
C2240 a_187922_n20028.n185 GND 0.009005f
C2241 a_187922_n20028.n186 GND 0.012007f
C2242 a_187922_n20028.n187 GND 0.003726f
C2243 a_187922_n20028.n188 GND 0.003519f
C2244 a_187922_n20028.n189 GND 0.010083f
C2245 a_187922_n20028.n190 GND 0.009718f
C2246 a_187922_n20028.n191 GND 0.003519f
C2247 a_187922_n20028.n192 GND 0.003726f
C2248 a_187922_n20028.n193 GND 0.003519f
C2249 a_187922_n20028.n194 GND 0.003726f
C2250 a_187922_n20028.n195 GND 0.021745f
C2251 a_187922_n20028.t20 GND 0.044142f
C2252 a_187922_n20028.t18 GND 0.044142f
C2253 a_187922_n20028.n196 GND 0.097902f
C2254 a_187922_n20028.n197 GND 0.009641f
C2255 a_187922_n20028.n198 GND 0.008904f
C2256 a_187922_n20028.n199 GND 0.009641f
C2257 a_187922_n20028.n200 GND 0.097902f
C2258 a_187922_n20028.t21 GND 0.044142f
C2259 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n0 GND 1.69497f
C2260 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n1 GND 1.75144f
C2261 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n2 GND 1.74613f
C2262 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n3 GND 0.056526f
C2263 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n4 GND 0.228294f
C2264 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n5 GND 0.056515f
C2265 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n6 GND 0.228016f
C2266 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t12 GND 0.027344f
C2267 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t11 GND 0.027344f
C2268 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n7 GND 0.082479f
C2269 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n8 GND 0.264487f
C2270 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t10 GND 0.027344f
C2271 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t14 GND 0.027344f
C2272 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n9 GND 0.071959f
C2273 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n10 GND 0.0195f
C2274 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n11 GND 0.006246f
C2275 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n12 GND 0.00436f
C2276 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t5 GND 0.006836f
C2277 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t3 GND 0.006836f
C2278 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n13 GND 0.007245f
C2279 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n14 GND 0.005564f
C2280 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n15 GND 0.013672f
C2281 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n16 GND 0.002639f
C2282 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n17 GND 0.010169f
C2283 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n18 GND 0.01728f
C2284 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t24 GND 0.295934f
C2285 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n19 GND 0.100861f
C2286 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n20 GND 0.110949f
C2287 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t0 GND 0.129031f
C2288 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n21 GND 0.010182f
C2289 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n22 GND 0.045176f
C2290 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n23 GND 0.110949f
C2291 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n24 GND 0.110949f
C2292 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n25 GND 0.110949f
C2293 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n26 GND 0.110949f
C2294 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n27 GND 0.110949f
C2295 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n28 GND 0.110949f
C2296 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n29 GND 0.171046f
C2297 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n30 GND 0.22925f
C2298 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n31 GND 0.110949f
C2299 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n32 GND 0.110949f
C2300 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n33 GND 0.110949f
C2301 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n34 GND 0.110949f
C2302 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n35 GND 0.110949f
C2303 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n36 GND 0.180384f
C2304 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t37 GND 0.295934f
C2305 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n37 GND 0.228717f
C2306 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t38 GND 0.295934f
C2307 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n38 GND 0.110949f
C2308 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n39 GND 0.110949f
C2309 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t44 GND 0.295934f
C2310 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n40 GND 0.110949f
C2311 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t47 GND 0.295934f
C2312 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n41 GND 0.110949f
C2313 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n42 GND 0.110949f
C2314 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t25 GND 0.295934f
C2315 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n43 GND 0.110949f
C2316 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t31 GND 0.295934f
C2317 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n44 GND 0.110949f
C2318 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n45 GND 0.110949f
C2319 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t42 GND 0.295934f
C2320 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n46 GND 0.110949f
C2321 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t18 GND 0.295934f
C2322 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n47 GND 0.110949f
C2323 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n48 GND 0.110949f
C2324 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t21 GND 0.295934f
C2325 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n49 GND 0.110949f
C2326 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t46 GND 0.295934f
C2327 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n50 GND 0.110949f
C2328 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n51 GND 0.110949f
C2329 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t22 GND 0.295934f
C2330 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n52 GND 0.110949f
C2331 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t36 GND 0.295934f
C2332 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n53 GND 0.181634f
C2333 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t28 GND 0.295934f
C2334 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n54 GND 0.171043f
C2335 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n55 GND 0.110949f
C2336 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t20 GND 0.295934f
C2337 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n56 GND 0.110949f
C2338 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t17 GND 0.295934f
C2339 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n57 GND 0.110949f
C2340 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n58 GND 0.110949f
C2341 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t41 GND 0.295934f
C2342 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n59 GND 0.110949f
C2343 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t16 GND 0.295934f
C2344 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n60 GND 0.110949f
C2345 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n61 GND 0.110949f
C2346 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t45 GND 0.295934f
C2347 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n62 GND 0.110949f
C2348 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t30 GND 0.295934f
C2349 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n63 GND 0.110949f
C2350 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n64 GND 0.110949f
C2351 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t27 GND 0.295934f
C2352 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n65 GND 0.110949f
C2353 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t19 GND 0.295934f
C2354 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n66 GND 0.110949f
C2355 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n67 GND 0.110949f
C2356 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t43 GND 0.295934f
C2357 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n68 GND 0.110949f
C2358 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t40 GND 0.295934f
C2359 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n69 GND 0.110949f
C2360 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n70 GND 0.110949f
C2361 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t26 GND 0.295934f
C2362 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n71 GND 0.110949f
C2363 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t34 GND 0.295934f
C2364 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n72 GND 0.110949f
C2365 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n73 GND 0.170021f
C2366 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t29 GND 0.295934f
C2367 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n74 GND 0.170021f
C2368 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n75 GND 1.69185f
C2369 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n76 GND 0.57847f
C2370 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t15 GND 0.027344f
C2371 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t13 GND 0.027344f
C2372 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n77 GND 0.071959f
C2373 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n78 GND 0.635126f
C2374 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n79 GND 0.205569f
C2375 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n80 GND 0.006246f
C2376 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n81 GND 0.00436f
C2377 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t1 GND 0.006836f
C2378 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n82 GND 0.002639f
C2379 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t7 GND 0.006836f
C2380 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n83 GND 0.013672f
C2381 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n84 GND 0.005564f
C2382 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n85 GND 0.00722f
C2383 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n86 GND 0.019452f
C2384 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t4 GND 0.129023f
C2385 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n87 GND 0.036847f
C2386 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t9 GND 0.013672f
C2387 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t8 GND 0.013672f
C2388 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n88 GND 0.061972f
C2389 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n89 GND 0.163966f
C2390 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n90 GND 0.036847f
C2391 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t6 GND 0.129023f
C2392 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n91 GND 0.045416f
C2393 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n92 GND 0.017458f
C2394 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n93 GND 0.069017f
C2395 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t33 GND 0.295934f
C2396 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n94 GND 0.101064f
C2397 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n95 GND 0.243666f
C2398 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t35 GND 0.295939f
C2399 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t39 GND 0.295934f
C2400 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n96 GND 0.108156f
C2401 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n97 GND 0.108183f
C2402 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t23 GND 0.295934f
C2403 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n98 GND 0.110949f
C2404 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n99 GND 0.243911f
C2405 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t32 GND 0.295939f
C2406 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n100 GND 0.068109f
C2407 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.t2 GND 0.129031f
C2408 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n101 GND 0.204251f
C2409 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n102 GND 0.633481f
C2410 C2S2_Amp_F_I_0.constant_gm_fingers_0.Vout.n103 GND 0.581303f
C2411 a_156122_n20028.n0 GND 4.09756f
C2412 a_156122_n20028.n1 GND 4.32222f
C2413 a_156122_n20028.n2 GND 0.036592f
C2414 a_156122_n20028.n3 GND 0.03655f
C2415 a_156122_n20028.n4 GND 0.856021f
C2416 a_156122_n20028.n5 GND 1.07316f
C2417 a_156122_n20028.n6 GND 1.07275f
C2418 a_156122_n20028.n7 GND 0.186041f
C2419 a_156122_n20028.n8 GND 0.172758f
C2420 a_156122_n20028.n9 GND 0.004162f
C2421 a_156122_n20028.n10 GND 0.172758f
C2422 a_156122_n20028.n11 GND 0.004162f
C2423 a_156122_n20028.n12 GND 0.172758f
C2424 a_156122_n20028.n13 GND 0.004162f
C2425 a_156122_n20028.n14 GND 0.172702f
C2426 a_156122_n20028.n15 GND 0.004192f
C2427 a_156122_n20028.n16 GND 0.172702f
C2428 a_156122_n20028.n17 GND 0.004192f
C2429 a_156122_n20028.n18 GND 0.172702f
C2430 a_156122_n20028.n19 GND 0.004192f
C2431 a_156122_n20028.n20 GND 0.794595f
C2432 a_156122_n20028.n21 GND 0.794182f
C2433 a_156122_n20028.n22 GND 0.043311f
C2434 a_156122_n20028.n23 GND 0.006798f
C2435 a_156122_n20028.n24 GND 0.043311f
C2436 a_156122_n20028.n25 GND 0.006798f
C2437 a_156122_n20028.n26 GND 0.043311f
C2438 a_156122_n20028.n27 GND 0.006798f
C2439 a_156122_n20028.n28 GND 0.04816f
C2440 a_156122_n20028.n29 GND 0.020206f
C2441 a_156122_n20028.n30 GND 0.043336f
C2442 a_156122_n20028.n31 GND 0.006799f
C2443 a_156122_n20028.n32 GND 0.043336f
C2444 a_156122_n20028.n33 GND 0.006799f
C2445 a_156122_n20028.n34 GND 0.043336f
C2446 a_156122_n20028.n35 GND 0.006799f
C2447 a_156122_n20028.n36 GND 0.043336f
C2448 a_156122_n20028.n37 GND 0.006799f
C2449 a_156122_n20028.n38 GND 0.043336f
C2450 a_156122_n20028.n39 GND 0.006799f
C2451 a_156122_n20028.n40 GND 0.020206f
C2452 a_156122_n20028.n41 GND 0.040234f
C2453 a_156122_n20028.n42 GND 0.040234f
C2454 a_156122_n20028.n43 GND 0.020206f
C2455 a_156122_n20028.n44 GND 0.008562f
C2456 a_156122_n20028.n45 GND 0.006799f
C2457 a_156122_n20028.n46 GND 0.043336f
C2458 a_156122_n20028.n47 GND 0.048206f
C2459 a_156122_n20028.n48 GND 0.020207f
C2460 a_156122_n20028.n49 GND 0.043358f
C2461 a_156122_n20028.n50 GND 0.006799f
C2462 a_156122_n20028.n51 GND 0.043358f
C2463 a_156122_n20028.n52 GND 0.006799f
C2464 a_156122_n20028.n53 GND 0.043358f
C2465 a_156122_n20028.n54 GND 0.006799f
C2466 a_156122_n20028.n55 GND 0.186041f
C2467 a_156122_n20028.n56 GND 0.005649f
C2468 a_156122_n20028.n57 GND 0.186041f
C2469 a_156122_n20028.n58 GND 0.005649f
C2470 a_156122_n20028.n59 GND 0.186041f
C2471 a_156122_n20028.n60 GND 0.005649f
C2472 a_156122_n20028.n61 GND 0.186041f
C2473 a_156122_n20028.n62 GND 0.005649f
C2474 a_156122_n20028.n63 GND 0.186041f
C2475 a_156122_n20028.n64 GND 0.005649f
C2476 a_156122_n20028.n65 GND 0.00927f
C2477 a_156122_n20028.n66 GND 0.020275f
C2478 a_156122_n20028.n67 GND 0.020275f
C2479 a_156122_n20028.n68 GND 0.005649f
C2480 a_156122_n20028.t17 GND 0.042445f
C2481 a_156122_n20028.t22 GND 0.042445f
C2482 a_156122_n20028.t10 GND 0.042445f
C2483 a_156122_n20028.n69 GND 0.094137f
C2484 a_156122_n20028.n70 GND 0.00927f
C2485 a_156122_n20028.n71 GND 0.008562f
C2486 a_156122_n20028.t1 GND 0.042445f
C2487 a_156122_n20028.n72 GND 0.003583f
C2488 a_156122_n20028.n73 GND 0.004438f
C2489 a_156122_n20028.n74 GND 0.009548f
C2490 a_156122_n20028.n75 GND 0.007707f
C2491 a_156122_n20028.n76 GND 0.009695f
C2492 a_156122_n20028.t7 GND 0.042445f
C2493 a_156122_n20028.n77 GND 0.091818f
C2494 a_156122_n20028.t9 GND 0.042445f
C2495 a_156122_n20028.n78 GND 0.003583f
C2496 a_156122_n20028.n79 GND 0.004438f
C2497 a_156122_n20028.n80 GND 0.009548f
C2498 a_156122_n20028.n81 GND 0.007707f
C2499 a_156122_n20028.n82 GND 0.009695f
C2500 a_156122_n20028.t2 GND 0.042445f
C2501 a_156122_n20028.n83 GND 0.091818f
C2502 a_156122_n20028.t24 GND 0.042445f
C2503 a_156122_n20028.n84 GND 0.003583f
C2504 a_156122_n20028.n85 GND 0.004438f
C2505 a_156122_n20028.n86 GND 0.009548f
C2506 a_156122_n20028.n87 GND 0.007707f
C2507 a_156122_n20028.n88 GND 0.009695f
C2508 a_156122_n20028.t4 GND 0.042445f
C2509 a_156122_n20028.n89 GND 0.091818f
C2510 a_156122_n20028.n90 GND 0.020909f
C2511 a_156122_n20028.n91 GND 0.003583f
C2512 a_156122_n20028.n92 GND 0.003384f
C2513 a_156122_n20028.n93 GND 0.011545f
C2514 a_156122_n20028.n94 GND 0.003583f
C2515 a_156122_n20028.n95 GND 0.027431f
C2516 a_156122_n20028.t27 GND 0.016571f
C2517 a_156122_n20028.n96 GND 0.008659f
C2518 a_156122_n20028.n97 GND 0.0042f
C2519 a_156122_n20028.n98 GND 0.003384f
C2520 a_156122_n20028.n99 GND 0.170043f
C2521 a_156122_n20028.n100 GND 0.003384f
C2522 a_156122_n20028.n101 GND 0.003583f
C2523 a_156122_n20028.n102 GND 0.011545f
C2524 a_156122_n20028.n103 GND 0.011545f
C2525 a_156122_n20028.n104 GND 0.003583f
C2526 a_156122_n20028.n105 GND 0.003384f
C2527 a_156122_n20028.n106 GND 0.009695f
C2528 a_156122_n20028.n107 GND 0.009548f
C2529 a_156122_n20028.n108 GND 0.004209f
C2530 a_156122_n20028.n109 GND 0.009695f
C2531 a_156122_n20028.n110 GND 0.003583f
C2532 a_156122_n20028.n111 GND 0.003384f
C2533 a_156122_n20028.n112 GND 0.00927f
C2534 a_156122_n20028.n113 GND 0.004209f
C2535 a_156122_n20028.n114 GND 0.003384f
C2536 a_156122_n20028.n115 GND 0.003583f
C2537 a_156122_n20028.n116 GND 0.020909f
C2538 a_156122_n20028.n117 GND 0.011545f
C2539 a_156122_n20028.n118 GND 0.008659f
C2540 a_156122_n20028.n119 GND 0.0042f
C2541 a_156122_n20028.t20 GND 0.016571f
C2542 a_156122_n20028.n120 GND 0.027431f
C2543 a_156122_n20028.n121 GND 0.170238f
C2544 a_156122_n20028.n122 GND 0.003384f
C2545 a_156122_n20028.n123 GND 0.003583f
C2546 a_156122_n20028.n124 GND 0.011545f
C2547 a_156122_n20028.n125 GND 0.011545f
C2548 a_156122_n20028.n126 GND 0.003583f
C2549 a_156122_n20028.n127 GND 0.003384f
C2550 a_156122_n20028.n128 GND 0.009344f
C2551 a_156122_n20028.t12 GND 0.042445f
C2552 a_156122_n20028.t11 GND 0.042445f
C2553 a_156122_n20028.n129 GND 0.094137f
C2554 a_156122_n20028.n130 GND 0.00927f
C2555 a_156122_n20028.n131 GND 0.008562f
C2556 a_156122_n20028.t18 GND 0.042445f
C2557 a_156122_n20028.t16 GND 0.042445f
C2558 a_156122_n20028.n132 GND 0.094137f
C2559 a_156122_n20028.n133 GND 0.00927f
C2560 a_156122_n20028.n134 GND 0.008562f
C2561 a_156122_n20028.n135 GND 1.25213f
C2562 a_156122_n20028.t6 GND 0.042445f
C2563 a_156122_n20028.t8 GND 0.042445f
C2564 a_156122_n20028.n136 GND 0.091792f
C2565 a_156122_n20028.n137 GND 0.003583f
C2566 a_156122_n20028.n138 GND 0.004438f
C2567 a_156122_n20028.n139 GND 0.0095f
C2568 a_156122_n20028.n140 GND 0.009695f
C2569 a_156122_n20028.n141 GND 0.007708f
C2570 a_156122_n20028.t26 GND 0.042445f
C2571 a_156122_n20028.t3 GND 0.042445f
C2572 a_156122_n20028.n142 GND 0.091792f
C2573 a_156122_n20028.n143 GND 0.003583f
C2574 a_156122_n20028.n144 GND 0.004438f
C2575 a_156122_n20028.n145 GND 0.0095f
C2576 a_156122_n20028.n146 GND 0.009695f
C2577 a_156122_n20028.n147 GND 0.007708f
C2578 a_156122_n20028.t5 GND 0.042445f
C2579 a_156122_n20028.t25 GND 0.042445f
C2580 a_156122_n20028.n148 GND 0.091792f
C2581 a_156122_n20028.n149 GND 0.003583f
C2582 a_156122_n20028.n150 GND 0.004438f
C2583 a_156122_n20028.n151 GND 0.0095f
C2584 a_156122_n20028.n152 GND 0.009695f
C2585 a_156122_n20028.n153 GND 0.007708f
C2586 a_156122_n20028.n154 GND 0.170001f
C2587 a_156122_n20028.n155 GND 0.003583f
C2588 a_156122_n20028.n156 GND 0.003384f
C2589 a_156122_n20028.n157 GND 0.020909f
C2590 a_156122_n20028.n158 GND 0.003583f
C2591 a_156122_n20028.n159 GND 0.004209f
C2592 a_156122_n20028.n160 GND 0.0095f
C2593 a_156122_n20028.n161 GND 0.009695f
C2594 a_156122_n20028.n162 GND 0.003384f
C2595 a_156122_n20028.n163 GND 0.003384f
C2596 a_156122_n20028.n164 GND 0.003583f
C2597 a_156122_n20028.n165 GND 0.011545f
C2598 a_156122_n20028.n166 GND 0.011545f
C2599 a_156122_n20028.t0 GND 0.016571f
C2600 a_156122_n20028.n167 GND 0.027431f
C2601 a_156122_n20028.n168 GND 0.0042f
C2602 a_156122_n20028.n169 GND 0.008659f
C2603 a_156122_n20028.n170 GND 0.011545f
C2604 a_156122_n20028.n171 GND 0.003583f
C2605 a_156122_n20028.n172 GND 0.003384f
C2606 a_156122_n20028.n173 GND 1.24834f
C2607 a_156122_n20028.n174 GND 0.004209f
C2608 a_156122_n20028.n175 GND 0.011545f
C2609 a_156122_n20028.n176 GND 0.003583f
C2610 a_156122_n20028.n177 GND 0.170238f
C2611 a_156122_n20028.n178 GND 0.003384f
C2612 a_156122_n20028.n179 GND 0.011545f
C2613 a_156122_n20028.t21 GND 0.016571f
C2614 a_156122_n20028.n180 GND 0.027431f
C2615 a_156122_n20028.n181 GND 0.0042f
C2616 a_156122_n20028.n182 GND 0.008659f
C2617 a_156122_n20028.n183 GND 0.011545f
C2618 a_156122_n20028.n184 GND 0.003583f
C2619 a_156122_n20028.n185 GND 0.003384f
C2620 a_156122_n20028.n186 GND 0.009695f
C2621 a_156122_n20028.n187 GND 0.009344f
C2622 a_156122_n20028.n188 GND 0.003384f
C2623 a_156122_n20028.n189 GND 0.003583f
C2624 a_156122_n20028.n190 GND 0.003384f
C2625 a_156122_n20028.n191 GND 0.003583f
C2626 a_156122_n20028.n192 GND 0.020909f
C2627 a_156122_n20028.t14 GND 0.042445f
C2628 a_156122_n20028.t13 GND 0.042445f
C2629 a_156122_n20028.n193 GND 0.094137f
C2630 a_156122_n20028.n194 GND 0.00927f
C2631 a_156122_n20028.n195 GND 0.008562f
C2632 a_156122_n20028.t15 GND 0.042445f
C2633 a_156122_n20028.t19 GND 0.042445f
C2634 a_156122_n20028.n196 GND 0.094137f
C2635 a_156122_n20028.n197 GND 0.00927f
C2636 a_156122_n20028.n198 GND 0.008562f
C2637 a_156122_n20028.n199 GND 0.00927f
C2638 a_156122_n20028.n200 GND 0.094137f
C2639 a_156122_n20028.t23 GND 0.042445f
C2640 a_214193_n11375.t7 GND 0.517854f
C2641 a_214193_n11375.t1 GND 0.52009f
C2642 a_214193_n11375.n0 GND 6.03626f
C2643 a_214193_n11375.t5 GND 20.8342f
C2644 a_214193_n11375.n1 GND 7.27757f
C2645 a_214193_n11375.t4 GND 20.8342f
C2646 a_214193_n11375.n2 GND 4.66798f
C2647 a_214193_n11375.t3 GND 20.8342f
C2648 a_214193_n11375.n3 GND 4.66798f
C2649 a_214193_n11375.t6 GND 20.8342f
C2650 a_214193_n11375.n4 GND 7.29735f
C2651 a_214193_n11375.t2 GND 0.519976f
C2652 a_214193_n11375.n5 GND 6.0404f
C2653 a_214193_n11375.t0 GND 0.517749f
C2654 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n0 GND 1.69497f
C2655 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n1 GND 1.75144f
C2656 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n2 GND 1.74613f
C2657 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n3 GND 0.056526f
C2658 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n4 GND 0.228294f
C2659 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n5 GND 0.056515f
C2660 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n6 GND 0.228016f
C2661 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t5 GND 0.027344f
C2662 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t4 GND 0.027344f
C2663 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n7 GND 0.082479f
C2664 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n8 GND 0.264487f
C2665 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n9 GND 0.0195f
C2666 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n10 GND 0.006246f
C2667 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n11 GND 0.00436f
C2668 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t11 GND 0.006836f
C2669 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t15 GND 0.006836f
C2670 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n12 GND 0.007245f
C2671 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n13 GND 0.005564f
C2672 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n14 GND 0.013672f
C2673 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n15 GND 0.002639f
C2674 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n16 GND 0.010169f
C2675 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n17 GND 0.01728f
C2676 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t24 GND 0.295934f
C2677 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n18 GND 0.100861f
C2678 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n19 GND 0.110949f
C2679 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n20 GND 0.017458f
C2680 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t6 GND 0.027344f
C2681 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t3 GND 0.027344f
C2682 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n21 GND 0.071959f
C2683 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n22 GND 0.110949f
C2684 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n23 GND 0.110949f
C2685 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n24 GND 0.110949f
C2686 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n25 GND 0.110949f
C2687 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n26 GND 0.110949f
C2688 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n27 GND 0.110949f
C2689 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n28 GND 0.171046f
C2690 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n29 GND 0.22925f
C2691 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n30 GND 0.110949f
C2692 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n31 GND 0.110949f
C2693 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n32 GND 0.110949f
C2694 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n33 GND 0.110949f
C2695 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n34 GND 0.110949f
C2696 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n35 GND 0.180384f
C2697 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t38 GND 0.295934f
C2698 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n36 GND 0.228717f
C2699 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t21 GND 0.295934f
C2700 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n37 GND 0.110949f
C2701 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n38 GND 0.110949f
C2702 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t47 GND 0.295934f
C2703 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n39 GND 0.110949f
C2704 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t17 GND 0.295934f
C2705 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n40 GND 0.110949f
C2706 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n41 GND 0.110949f
C2707 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t22 GND 0.295934f
C2708 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n42 GND 0.110949f
C2709 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t18 GND 0.295934f
C2710 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n43 GND 0.110949f
C2711 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n44 GND 0.110949f
C2712 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t29 GND 0.295934f
C2713 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n45 GND 0.110949f
C2714 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t39 GND 0.295934f
C2715 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n46 GND 0.110949f
C2716 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n47 GND 0.110949f
C2717 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t41 GND 0.295934f
C2718 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n48 GND 0.110949f
C2719 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t34 GND 0.295934f
C2720 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n49 GND 0.110949f
C2721 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n50 GND 0.110949f
C2722 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t43 GND 0.295934f
C2723 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n51 GND 0.110949f
C2724 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t23 GND 0.295934f
C2725 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n52 GND 0.181634f
C2726 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t25 GND 0.295934f
C2727 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n53 GND 0.171043f
C2728 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n54 GND 0.110949f
C2729 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t40 GND 0.295934f
C2730 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n55 GND 0.110949f
C2731 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t37 GND 0.295934f
C2732 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n56 GND 0.110949f
C2733 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n57 GND 0.110949f
C2734 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t28 GND 0.295934f
C2735 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n58 GND 0.110949f
C2736 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t36 GND 0.295934f
C2737 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n59 GND 0.110949f
C2738 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n60 GND 0.110949f
C2739 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t32 GND 0.295934f
C2740 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n61 GND 0.110949f
C2741 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t16 GND 0.295934f
C2742 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n62 GND 0.110949f
C2743 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n63 GND 0.110949f
C2744 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t46 GND 0.295934f
C2745 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n64 GND 0.110949f
C2746 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t20 GND 0.295934f
C2747 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n65 GND 0.110949f
C2748 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n66 GND 0.110949f
C2749 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t45 GND 0.295934f
C2750 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n67 GND 0.110949f
C2751 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t42 GND 0.295934f
C2752 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n68 GND 0.110949f
C2753 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n69 GND 0.110949f
C2754 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t35 GND 0.295934f
C2755 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n70 GND 0.110949f
C2756 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t31 GND 0.295934f
C2757 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n71 GND 0.110949f
C2758 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n72 GND 0.170021f
C2759 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t26 GND 0.295934f
C2760 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n73 GND 0.170021f
C2761 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n74 GND 1.69185f
C2762 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n75 GND 0.57847f
C2763 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n76 GND 0.635126f
C2764 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n77 GND 0.006246f
C2765 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n78 GND 0.00436f
C2766 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t9 GND 0.006836f
C2767 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n79 GND 0.010182f
C2768 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n80 GND 0.002639f
C2769 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t13 GND 0.006836f
C2770 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n81 GND 0.013672f
C2771 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n82 GND 0.005564f
C2772 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n83 GND 0.00722f
C2773 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t1 GND 0.013672f
C2774 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t0 GND 0.013672f
C2775 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n84 GND 0.061972f
C2776 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n85 GND 0.163966f
C2777 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n86 GND 0.036847f
C2778 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t10 GND 0.129023f
C2779 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n87 GND 0.045176f
C2780 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n88 GND 0.045416f
C2781 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t12 GND 0.129023f
C2782 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n89 GND 0.036847f
C2783 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n90 GND 0.019452f
C2784 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n91 GND 0.205569f
C2785 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t8 GND 0.129031f
C2786 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n92 GND 0.069017f
C2787 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t30 GND 0.295934f
C2788 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n93 GND 0.101064f
C2789 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n94 GND 0.243666f
C2790 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t33 GND 0.295939f
C2791 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t27 GND 0.295934f
C2792 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n95 GND 0.108156f
C2793 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n96 GND 0.108183f
C2794 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t44 GND 0.295934f
C2795 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n97 GND 0.110949f
C2796 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n98 GND 0.243911f
C2797 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t19 GND 0.295939f
C2798 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n99 GND 0.068109f
C2799 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t14 GND 0.129031f
C2800 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n100 GND 0.204251f
C2801 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t2 GND 0.027344f
C2802 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.t7 GND 0.027344f
C2803 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n101 GND 0.071959f
C2804 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n102 GND 0.633481f
C2805 C2S2_Amp_F_I_1.constant_gm_fingers_0.Vout.n103 GND 0.581303f
C2806 a_157137_n26928.n0 GND 0.224177f
C2807 a_157137_n26928.n1 GND 0.580261f
C2808 a_157137_n26928.n2 GND 0.281977f
C2809 a_157137_n26928.n3 GND 0.060445f
C2810 a_157137_n26928.n4 GND 0.358112f
C2811 a_157137_n26928.n5 GND 0.060445f
C2812 a_157137_n26928.n6 GND 0.358203f
C2813 a_157137_n26928.n7 GND 1.26025f
C2814 a_157137_n26928.n8 GND 0.94806f
C2815 a_157137_n26928.n9 GND 0.272686f
C2816 a_157137_n26928.n10 GND 0.414211f
C2817 a_157137_n26928.n11 GND 0.361457f
C2818 a_157137_n26928.n12 GND 0.223547f
C2819 a_157137_n26928.n13 GND 0.061415f
C2820 a_157137_n26928.n14 GND 0.368761f
C2821 a_157137_n26928.n15 GND 0.220921f
C2822 a_157137_n26928.n16 GND 0.044676f
C2823 a_157137_n26928.n17 GND 0.026567f
C2824 a_157137_n26928.n18 GND 0.011146f
C2825 a_157137_n26928.n19 GND 0.044676f
C2826 a_157137_n26928.n20 GND 0.026567f
C2827 a_157137_n26928.n21 GND 0.011146f
C2828 a_157137_n26928.n22 GND 0.246237f
C2829 a_157137_n26928.n23 GND 0.246237f
C2830 a_157137_n26928.n24 GND 0.026567f
C2831 a_157137_n26928.n25 GND 0.026567f
C2832 a_157137_n26928.n26 GND 0.026567f
C2833 a_157137_n26928.n27 GND 0.026567f
C2834 a_157137_n26928.n28 GND 0.027418f
C2835 a_157137_n26928.n29 GND 0.026567f
C2836 a_157137_n26928.n30 GND 0.026567f
C2837 a_157137_n26928.n31 GND 0.026567f
C2838 a_157137_n26928.n32 GND 0.026492f
C2839 a_157137_n26928.n33 GND 0.026567f
C2840 a_157137_n26928.n34 GND 0.026567f
C2841 a_157137_n26928.n35 GND 0.026567f
C2842 a_157137_n26928.n36 GND 0.026567f
C2843 a_157137_n26928.n37 GND 0.027418f
C2844 a_157137_n26928.n38 GND 0.006751f
C2845 a_157137_n26928.n39 GND 0.009775f
C2846 a_157137_n26928.n40 GND 0.009775f
C2847 a_157137_n26928.n41 GND 0.004636f
C2848 a_157137_n26928.n42 GND 0.013284f
C2849 a_157137_n26928.n43 GND 0.009775f
C2850 a_157137_n26928.n44 GND 0.013496f
C2851 a_157137_n26928.n45 GND 0.047048f
C2852 a_157137_n26928.n46 GND 0.011146f
C2853 a_157137_n26928.n47 GND 0.013496f
C2854 a_157137_n26928.n48 GND 0.047048f
C2855 a_157137_n26928.n49 GND 0.011146f
C2856 a_157137_n26928.n50 GND 0.008165f
C2857 a_157137_n26928.n51 GND 0.009311f
C2858 a_157137_n26928.n52 GND 0.564647f
C2859 a_157137_n26928.n53 GND 0.11767f
C2860 a_157137_n26928.n54 GND 0.563925f
C2861 a_157137_n26928.n55 GND 0.117768f
C2862 a_157137_n26928.n56 GND 0.162595f
C2863 a_157137_n26928.n57 GND 0.032543f
C2864 a_157137_n26928.n58 GND 0.162595f
C2865 a_157137_n26928.n59 GND 0.032543f
C2866 a_157137_n26928.t6 GND 0.058156f
C2867 a_157137_n26928.n60 GND 0.004909f
C2868 a_157137_n26928.n61 GND 0.004909f
C2869 a_157137_n26928.n62 GND 0.004909f
C2870 a_157137_n26928.n63 GND 5.41e-19
C2871 a_157137_n26928.n64 GND 0.004909f
C2872 a_157137_n26928.n65 GND 0.004909f
C2873 a_157137_n26928.n66 GND 0.004909f
C2874 a_157137_n26928.n67 GND 0.004909f
C2875 a_157137_n26928.n68 GND 0.004909f
C2876 a_157137_n26928.n69 GND 0.00585f
C2877 a_157137_n26928.n70 GND 0.011864f
C2878 a_157137_n26928.n71 GND 0.005755f
C2879 a_157137_n26928.t20 GND 0.022705f
C2880 a_157137_n26928.n72 GND 0.037585f
C2881 a_157137_n26928.n73 GND 0.004636f
C2882 a_157137_n26928.n74 GND 0.004909f
C2883 a_157137_n26928.n75 GND 0.02808f
C2884 a_157137_n26928.n76 GND 0.004636f
C2885 a_157137_n26928.n77 GND 0.004636f
C2886 a_157137_n26928.n78 GND 0.004636f
C2887 a_157137_n26928.n79 GND 0.004636f
C2888 a_157137_n26928.n80 GND 0.009139f
C2889 a_157137_n26928.n81 GND 0.009139f
C2890 a_157137_n26928.n82 GND 0.004636f
C2891 a_157137_n26928.n83 GND 0.004636f
C2892 a_157137_n26928.n84 GND 0.240763f
C2893 a_157137_n26928.t5 GND 0.634271f
C2894 a_157137_n26928.n85 GND 0.224177f
C2895 a_157137_n26928.t12 GND 0.058156f
C2896 a_157137_n26928.n86 GND 0.004909f
C2897 a_157137_n26928.n87 GND 0.004909f
C2898 a_157137_n26928.n88 GND 0.004909f
C2899 a_157137_n26928.n89 GND 0.004909f
C2900 a_157137_n26928.n90 GND 5.41e-19
C2901 a_157137_n26928.n91 GND 0.004909f
C2902 a_157137_n26928.n92 GND 0.004909f
C2903 a_157137_n26928.n93 GND 0.004909f
C2904 a_157137_n26928.t14 GND 0.058156f
C2905 a_157137_n26928.n94 GND 0.004909f
C2906 a_157137_n26928.n95 GND 0.004909f
C2907 a_157137_n26928.n96 GND 0.004909f
C2908 a_157137_n26928.n97 GND 0.004909f
C2909 a_157137_n26928.n98 GND 0.004909f
C2910 a_157137_n26928.n99 GND 5.41e-19
C2911 a_157137_n26928.n100 GND 0.004909f
C2912 a_157137_n26928.n101 GND 0.004909f
C2913 a_157137_n26928.n102 GND 0.004909f
C2914 a_157137_n26928.n103 GND 0.004636f
C2915 a_157137_n26928.n104 GND 0.004636f
C2916 a_157137_n26928.n105 GND 0.004636f
C2917 a_157137_n26928.n106 GND 0.004636f
C2918 a_157137_n26928.n107 GND 0.004636f
C2919 a_157137_n26928.n108 GND 0.009139f
C2920 a_157137_n26928.n109 GND 0.009139f
C2921 a_157137_n26928.n110 GND 0.004636f
C2922 a_157137_n26928.n111 GND 0.004636f
C2923 a_157137_n26928.n112 GND 0.006751f
C2924 a_157137_n26928.t8 GND 0.058156f
C2925 a_157137_n26928.n113 GND 0.116585f
C2926 a_157137_n26928.t24 GND 0.634271f
C2927 a_157137_n26928.n114 GND 0.240763f
C2928 a_157137_n26928.n115 GND 0.559694f
C2929 a_157137_n26928.t26 GND 0.634271f
C2930 a_157137_n26928.n116 GND 0.23991f
C2931 a_157137_n26928.t23 GND 0.634277f
C2932 a_157137_n26928.t0 GND 0.058156f
C2933 a_157137_n26928.t21 GND 0.058156f
C2934 a_157137_n26928.n117 GND 0.245256f
C2935 a_157137_n26928.t17 GND 0.058156f
C2936 a_157137_n26928.t19 GND 0.058156f
C2937 a_157137_n26928.n118 GND 0.245256f
C2938 a_157137_n26928.n119 GND 0.00585f
C2939 a_157137_n26928.n120 GND 0.011864f
C2940 a_157137_n26928.n121 GND 0.005755f
C2941 a_157137_n26928.t18 GND 0.022705f
C2942 a_157137_n26928.n122 GND 0.037585f
C2943 a_157137_n26928.n123 GND 0.004636f
C2944 a_157137_n26928.n124 GND 0.004909f
C2945 a_157137_n26928.n125 GND 0.02808f
C2946 a_157137_n26928.n126 GND 1.25657f
C2947 a_157137_n26928.n127 GND 0.519726f
C2948 a_157137_n26928.t13 GND 0.634277f
C2949 a_157137_n26928.n128 GND 0.223919f
C2950 a_157137_n26928.t7 GND 0.634271f
C2951 a_157137_n26928.t11 GND 0.634271f
C2952 a_157137_n26928.t9 GND 0.634271f
C2953 a_157137_n26928.n129 GND 5.48e-19
C2954 a_157137_n26928.t4 GND 0.029078f
C2955 a_157137_n26928.n130 GND 0.004909f
C2956 a_157137_n26928.n131 GND 0.010014f
C2957 a_157137_n26928.n132 GND 0.009273f
C2958 a_157137_n26928.n133 GND 0.005654f
C2959 a_157137_n26928.n134 GND 0.087871f
C2960 a_157137_n26928.t3 GND 0.200999f
C2961 a_157137_n26928.n135 GND 0.081473f
C2962 a_157137_n26928.t2 GND 0.029078f
C2963 a_157137_n26928.n136 GND 5.48e-19
C2964 a_157137_n26928.n137 GND 0.004909f
C2965 a_157137_n26928.n138 GND 0.010014f
C2966 a_157137_n26928.n139 GND 0.009273f
C2967 a_157137_n26928.n140 GND 0.005654f
C2968 a_157137_n26928.n141 GND 0.087871f
C2969 a_157137_n26928.n142 GND 0.081473f
C2970 a_157137_n26928.t1 GND 0.200999f
C2971 a_157137_n26928.n143 GND 0.006121f
C2972 a_157137_n26928.n144 GND 0.004636f
C2973 a_157137_n26928.n145 GND 0.004636f
C2974 a_157137_n26928.n146 GND 0.004636f
C2975 a_157137_n26928.n147 GND 0.009139f
C2976 a_157137_n26928.n148 GND 0.009139f
C2977 a_157137_n26928.n149 GND 0.004636f
C2978 a_157137_n26928.n150 GND 0.004636f
C2979 a_157137_n26928.n151 GND 0.006751f
C2980 a_157137_n26928.t10 GND 0.058156f
C2981 a_157137_n26928.n152 GND 0.116684f
C2982 a_157137_n26928.t25 GND 0.634271f
C2983 a_157137_n26928.n153 GND 0.223547f
C2984 a_157137_n26928.n154 GND 0.239955f
C2985 a_157137_n26928.t27 GND 0.634271f
C2986 a_157137_n26928.n155 GND 0.559878f
C2987 a_157137_n26928.t22 GND 0.634276f
C2988 a_157137_n26928.t15 GND 0.634276f
C2989 a_157137_n26928.n156 GND 0.008165f
C2990 a_157137_n26928.n157 GND 0.116585f
C2991 a_157137_n26928.t16 GND 0.058156f
C2992 a_188937_n26928.n0 GND 0.224177f
C2993 a_188937_n26928.n1 GND 0.580261f
C2994 a_188937_n26928.n2 GND 0.414211f
C2995 a_188937_n26928.n3 GND 0.281977f
C2996 a_188937_n26928.n4 GND 0.223919f
C2997 a_188937_n26928.n5 GND 0.060445f
C2998 a_188937_n26928.n6 GND 0.358112f
C2999 a_188937_n26928.n7 GND 0.060445f
C3000 a_188937_n26928.n8 GND 0.358203f
C3001 a_188937_n26928.n9 GND 0.94806f
C3002 a_188937_n26928.n10 GND 0.272686f
C3003 a_188937_n26928.n11 GND 0.061415f
C3004 a_188937_n26928.n12 GND 0.368761f
C3005 a_188937_n26928.n13 GND 0.361457f
C3006 a_188937_n26928.n14 GND 0.220921f
C3007 a_188937_n26928.n15 GND 0.044676f
C3008 a_188937_n26928.n16 GND 0.026567f
C3009 a_188937_n26928.n17 GND 0.011146f
C3010 a_188937_n26928.n18 GND 0.044676f
C3011 a_188937_n26928.n19 GND 0.026567f
C3012 a_188937_n26928.n20 GND 0.011146f
C3013 a_188937_n26928.n21 GND 0.246237f
C3014 a_188937_n26928.n22 GND 0.246237f
C3015 a_188937_n26928.n23 GND 0.026567f
C3016 a_188937_n26928.n24 GND 0.026567f
C3017 a_188937_n26928.n25 GND 0.026567f
C3018 a_188937_n26928.n26 GND 0.026567f
C3019 a_188937_n26928.n27 GND 0.027418f
C3020 a_188937_n26928.n28 GND 0.026567f
C3021 a_188937_n26928.n29 GND 0.026567f
C3022 a_188937_n26928.n30 GND 0.026567f
C3023 a_188937_n26928.n31 GND 0.026567f
C3024 a_188937_n26928.n32 GND 0.027418f
C3025 a_188937_n26928.n33 GND 0.026567f
C3026 a_188937_n26928.n34 GND 0.026567f
C3027 a_188937_n26928.n35 GND 0.026567f
C3028 a_188937_n26928.n36 GND 0.026492f
C3029 a_188937_n26928.n37 GND 0.006751f
C3030 a_188937_n26928.n38 GND 0.009775f
C3031 a_188937_n26928.n39 GND 0.009775f
C3032 a_188937_n26928.n40 GND 0.006751f
C3033 a_188937_n26928.n41 GND 0.009775f
C3034 a_188937_n26928.n42 GND 0.013284f
C3035 a_188937_n26928.n43 GND 0.013496f
C3036 a_188937_n26928.n44 GND 0.047048f
C3037 a_188937_n26928.n45 GND 0.011146f
C3038 a_188937_n26928.n46 GND 0.013496f
C3039 a_188937_n26928.n47 GND 0.047048f
C3040 a_188937_n26928.n48 GND 0.011146f
C3041 a_188937_n26928.n49 GND 0.008165f
C3042 a_188937_n26928.n50 GND 0.009311f
C3043 a_188937_n26928.n51 GND 0.564647f
C3044 a_188937_n26928.n52 GND 0.11767f
C3045 a_188937_n26928.n53 GND 0.563925f
C3046 a_188937_n26928.n54 GND 0.117768f
C3047 a_188937_n26928.n55 GND 0.162595f
C3048 a_188937_n26928.n56 GND 0.032543f
C3049 a_188937_n26928.n57 GND 0.162595f
C3050 a_188937_n26928.n58 GND 0.032543f
C3051 a_188937_n26928.n59 GND 0.004909f
C3052 a_188937_n26928.n60 GND 0.004909f
C3053 a_188937_n26928.n61 GND 5.41e-19
C3054 a_188937_n26928.n62 GND 0.004909f
C3055 a_188937_n26928.t18 GND 0.058156f
C3056 a_188937_n26928.n63 GND 0.004909f
C3057 a_188937_n26928.n64 GND 0.004909f
C3058 a_188937_n26928.n65 GND 0.004909f
C3059 a_188937_n26928.n66 GND 0.004909f
C3060 a_188937_n26928.n67 GND 0.006121f
C3061 a_188937_n26928.n68 GND 0.004636f
C3062 a_188937_n26928.n69 GND 0.004636f
C3063 a_188937_n26928.n70 GND 0.004636f
C3064 a_188937_n26928.n71 GND 0.009139f
C3065 a_188937_n26928.n72 GND 0.009139f
C3066 a_188937_n26928.n73 GND 0.004636f
C3067 a_188937_n26928.n74 GND 0.004636f
C3068 a_188937_n26928.n75 GND 0.004636f
C3069 a_188937_n26928.t16 GND 0.058156f
C3070 a_188937_n26928.n76 GND 0.004909f
C3071 a_188937_n26928.n77 GND 0.004909f
C3072 a_188937_n26928.n78 GND 0.004909f
C3073 a_188937_n26928.n79 GND 0.004909f
C3074 a_188937_n26928.n80 GND 0.004909f
C3075 a_188937_n26928.n81 GND 5.41e-19
C3076 a_188937_n26928.n82 GND 0.004909f
C3077 a_188937_n26928.n83 GND 0.004909f
C3078 a_188937_n26928.n84 GND 0.004909f
C3079 a_188937_n26928.t12 GND 0.058156f
C3080 a_188937_n26928.n85 GND 0.004636f
C3081 a_188937_n26928.n86 GND 0.004636f
C3082 a_188937_n26928.n87 GND 0.004636f
C3083 a_188937_n26928.n88 GND 0.004636f
C3084 a_188937_n26928.n89 GND 0.009139f
C3085 a_188937_n26928.n90 GND 0.009139f
C3086 a_188937_n26928.n91 GND 0.004636f
C3087 a_188937_n26928.n92 GND 0.004636f
C3088 a_188937_n26928.n93 GND 0.116585f
C3089 a_188937_n26928.n94 GND 0.008165f
C3090 a_188937_n26928.n95 GND 0.559878f
C3091 a_188937_n26928.t23 GND 0.634276f
C3092 a_188937_n26928.t27 GND 0.63427f
C3093 a_188937_n26928.n96 GND 0.239955f
C3094 a_188937_n26928.n97 GND 0.223547f
C3095 a_188937_n26928.t26 GND 0.63427f
C3096 a_188937_n26928.n98 GND 0.240763f
C3097 a_188937_n26928.t25 GND 0.63427f
C3098 a_188937_n26928.n99 GND 0.240763f
C3099 a_188937_n26928.n100 GND 0.559693f
C3100 a_188937_n26928.t24 GND 0.63427f
C3101 a_188937_n26928.n101 GND 0.23991f
C3102 a_188937_n26928.t22 GND 0.634276f
C3103 a_188937_n26928.t19 GND 0.63427f
C3104 a_188937_n26928.t9 GND 0.63427f
C3105 a_188937_n26928.t14 GND 0.058156f
C3106 a_188937_n26928.n102 GND 0.004909f
C3107 a_188937_n26928.n103 GND 0.004909f
C3108 a_188937_n26928.n104 GND 0.004909f
C3109 a_188937_n26928.n105 GND 0.004909f
C3110 a_188937_n26928.n106 GND 0.004909f
C3111 a_188937_n26928.n107 GND 5.41e-19
C3112 a_188937_n26928.n108 GND 0.004909f
C3113 a_188937_n26928.n109 GND 0.004909f
C3114 a_188937_n26928.n110 GND 0.004909f
C3115 a_188937_n26928.n111 GND 0.004636f
C3116 a_188937_n26928.n112 GND 0.004636f
C3117 a_188937_n26928.n113 GND 0.004636f
C3118 a_188937_n26928.n114 GND 0.004636f
C3119 a_188937_n26928.n115 GND 0.004636f
C3120 a_188937_n26928.n116 GND 0.009139f
C3121 a_188937_n26928.n117 GND 0.009139f
C3122 a_188937_n26928.n118 GND 0.004636f
C3123 a_188937_n26928.n119 GND 0.004636f
C3124 a_188937_n26928.n120 GND 0.006751f
C3125 a_188937_n26928.t10 GND 0.058156f
C3126 a_188937_n26928.n121 GND 0.116585f
C3127 a_188937_n26928.t13 GND 0.634276f
C3128 a_188937_n26928.n122 GND 0.519726f
C3129 a_188937_n26928.n123 GND 0.00585f
C3130 a_188937_n26928.n124 GND 0.011864f
C3131 a_188937_n26928.n125 GND 0.005755f
C3132 a_188937_n26928.t4 GND 0.022705f
C3133 a_188937_n26928.n126 GND 0.037585f
C3134 a_188937_n26928.n127 GND 0.004636f
C3135 a_188937_n26928.n128 GND 0.004909f
C3136 a_188937_n26928.n129 GND 0.02808f
C3137 a_188937_n26928.n130 GND 1.25657f
C3138 a_188937_n26928.t1 GND 0.058156f
C3139 a_188937_n26928.t3 GND 0.058156f
C3140 a_188937_n26928.n131 GND 0.245256f
C3141 a_188937_n26928.t21 GND 0.058156f
C3142 a_188937_n26928.t0 GND 0.058156f
C3143 a_188937_n26928.n132 GND 0.245256f
C3144 a_188937_n26928.n133 GND 0.00585f
C3145 a_188937_n26928.n134 GND 0.011864f
C3146 a_188937_n26928.n135 GND 0.005755f
C3147 a_188937_n26928.t2 GND 0.022705f
C3148 a_188937_n26928.n136 GND 0.037585f
C3149 a_188937_n26928.n137 GND 0.004636f
C3150 a_188937_n26928.n138 GND 0.004909f
C3151 a_188937_n26928.n139 GND 0.02808f
C3152 a_188937_n26928.n140 GND 1.26025f
C3153 a_188937_n26928.t11 GND 0.634276f
C3154 a_188937_n26928.t15 GND 0.63427f
C3155 a_188937_n26928.n141 GND 0.224177f
C3156 a_188937_n26928.n142 GND 0.223547f
C3157 a_188937_n26928.t17 GND 0.63427f
C3158 a_188937_n26928.n143 GND 5.48e-19
C3159 a_188937_n26928.t8 GND 0.029078f
C3160 a_188937_n26928.n144 GND 0.004909f
C3161 a_188937_n26928.n145 GND 0.010014f
C3162 a_188937_n26928.n146 GND 0.009273f
C3163 a_188937_n26928.n147 GND 0.005654f
C3164 a_188937_n26928.n148 GND 0.087871f
C3165 a_188937_n26928.t7 GND 0.200999f
C3166 a_188937_n26928.n149 GND 0.081473f
C3167 a_188937_n26928.t6 GND 0.029078f
C3168 a_188937_n26928.n150 GND 5.48e-19
C3169 a_188937_n26928.n151 GND 0.004909f
C3170 a_188937_n26928.n152 GND 0.010014f
C3171 a_188937_n26928.n153 GND 0.009273f
C3172 a_188937_n26928.n154 GND 0.005654f
C3173 a_188937_n26928.n155 GND 0.087871f
C3174 a_188937_n26928.n156 GND 0.081473f
C3175 a_188937_n26928.t5 GND 0.200999f
C3176 a_188937_n26928.n157 GND 0.116684f
C3177 a_188937_n26928.t20 GND 0.058156f
C3178 a_188130_n13996.n0 GND 0.043242f
C3179 a_188130_n13996.n1 GND 0.043242f
C3180 a_188130_n13996.n2 GND 0.084714f
C3181 a_188130_n13996.n3 GND 0.03304f
C3182 a_188130_n13996.n4 GND 0.03304f
C3183 a_188130_n13996.n5 GND 0.005132f
C3184 a_188130_n13996.n6 GND 0.041278f
C3185 a_188130_n13996.n7 GND 0.065687f
C3186 a_188130_n13996.n8 GND 0.01031f
C3187 a_188130_n13996.n9 GND 0.065687f
C3188 a_188130_n13996.n10 GND 0.01031f
C3189 a_188130_n13996.n11 GND 0.065687f
C3190 a_188130_n13996.n12 GND 0.01031f
C3191 a_188130_n13996.n13 GND 0.07304f
C3192 a_188130_n13996.n14 GND 0.030644f
C3193 a_188130_n13996.n15 GND 2.89225f
C3194 a_188130_n13996.n16 GND 0.06592f
C3195 a_188130_n13996.n17 GND 0.010339f
C3196 a_188130_n13996.n18 GND 0.041899f
C3197 a_188130_n13996.n19 GND 0.023688f
C3198 a_188130_n13996.n20 GND 0.043297f
C3199 a_188130_n13996.n21 GND 0.03124f
C3200 a_188130_n13996.n22 GND 0.03124f
C3201 a_188130_n13996.n23 GND 0.01892f
C3202 a_188130_n13996.n24 GND 0.043297f
C3203 a_188130_n13996.n25 GND 0.06592f
C3204 a_188130_n13996.n26 GND 0.010339f
C3205 a_188130_n13996.n27 GND 0.06592f
C3206 a_188130_n13996.n28 GND 0.010339f
C3207 a_188130_n13996.n29 GND 0.06592f
C3208 a_188130_n13996.n30 GND 0.010339f
C3209 a_188130_n13996.n31 GND 0.06592f
C3210 a_188130_n13996.n32 GND 0.010339f
C3211 a_188130_n13996.n33 GND 0.070626f
C3212 a_188130_n13996.n34 GND 0.026553f
C3213 a_188130_n13996.n35 GND 0.06592f
C3214 a_188130_n13996.n36 GND 0.010339f
C3215 a_188130_n13996.n37 GND 2.85906f
C3216 a_188130_n13996.n38 GND 0.119184f
C3217 a_188130_n13996.n39 GND 0.492083f
C3218 a_188130_n13996.t11 GND 0.064372f
C3219 a_188130_n13996.n40 GND 0.011644f
C3220 a_188130_n13996.n41 GND 0.005434f
C3221 a_188130_n13996.n42 GND 0.263581f
C3222 a_188130_n13996.t27 GND 0.064372f
C3223 a_188130_n13996.n43 GND 0.005434f
C3224 a_188130_n13996.n44 GND 0.006774f
C3225 a_188130_n13996.n45 GND 0.014408f
C3226 a_188130_n13996.n46 GND 0.013908f
C3227 a_188130_n13996.n47 GND 0.011863f
C3228 a_188130_n13996.n48 GND 0.011644f
C3229 a_188130_n13996.t21 GND 0.064372f
C3230 a_188130_n13996.n49 GND 0.132696f
C3231 a_188130_n13996.n50 GND 0.451349f
C3232 a_188130_n13996.n51 GND 0.006774f
C3233 a_188130_n13996.n52 GND 0.014408f
C3234 a_188130_n13996.n53 GND 0.011863f
C3235 a_188130_n13996.n54 GND 0.013908f
C3236 a_188130_n13996.n55 GND 0.263581f
C3237 a_188130_n13996.n56 GND 0.263581f
C3238 a_188130_n13996.n57 GND 0.263581f
C3239 a_188130_n13996.n58 GND 0.263581f
C3240 a_188130_n13996.n59 GND 0.263581f
C3241 a_188130_n13996.t9 GND 0.064372f
C3242 a_188130_n13996.n60 GND 0.005434f
C3243 a_188130_n13996.n61 GND 0.006774f
C3244 a_188130_n13996.n62 GND 0.014408f
C3245 a_188130_n13996.n63 GND 0.013908f
C3246 a_188130_n13996.n64 GND 0.011863f
C3247 a_188130_n13996.n65 GND 0.011644f
C3248 a_188130_n13996.t31 GND 0.064372f
C3249 a_188130_n13996.n66 GND 0.132696f
C3250 a_188130_n13996.n67 GND 0.504623f
C3251 a_188130_n13996.n68 GND 0.419527f
C3252 a_188130_n13996.n69 GND 0.005434f
C3253 a_188130_n13996.n70 GND 0.005132f
C3254 a_188130_n13996.t35 GND 0.064372f
C3255 a_188130_n13996.n71 GND 0.009037f
C3256 a_188130_n13996.n72 GND 0.005132f
C3257 a_188130_n13996.n73 GND 0.005434f
C3258 a_188130_n13996.n74 GND 0.005132f
C3259 a_188130_n13996.n75 GND 0.005434f
C3260 a_188130_n13996.n76 GND 0.005434f
C3261 a_188130_n13996.n77 GND 5.99e-19
C3262 a_188130_n13996.n78 GND 0.005434f
C3263 a_188130_n13996.n79 GND 0.005434f
C3264 a_188130_n13996.n80 GND 0.005434f
C3265 a_188130_n13996.n81 GND 0.005434f
C3266 a_188130_n13996.n82 GND 0.005434f
C3267 a_188130_n13996.t29 GND 0.064372f
C3268 a_188130_n13996.n83 GND 0.125843f
C3269 a_188130_n13996.n84 GND 0.137608f
C3270 a_188130_n13996.t32 GND 0.355184f
C3271 a_188130_n13996.n85 GND 0.137608f
C3272 a_188130_n13996.n86 GND 0.030321f
C3273 a_188130_n13996.n87 GND 0.019178f
C3274 a_188130_n13996.n88 GND 0.005132f
C3275 a_188130_n13996.t25 GND 0.064372f
C3276 a_188130_n13996.n89 GND 0.009037f
C3277 a_188130_n13996.n90 GND 0.005434f
C3278 a_188130_n13996.n91 GND 0.005434f
C3279 a_188130_n13996.n92 GND 0.005434f
C3280 a_188130_n13996.n93 GND 0.005434f
C3281 a_188130_n13996.n94 GND 0.005434f
C3282 a_188130_n13996.n95 GND 5.99e-19
C3283 a_188130_n13996.n96 GND 0.005434f
C3284 a_188130_n13996.n97 GND 0.005434f
C3285 a_188130_n13996.n98 GND 0.005434f
C3286 a_188130_n13996.n99 GND 0.005434f
C3287 a_188130_n13996.n100 GND 0.005132f
C3288 a_188130_n13996.n101 GND 0.016538f
C3289 a_188130_n13996.n102 GND 0.005132f
C3290 a_188130_n13996.n103 GND 0.01892f
C3291 a_188130_n13996.n104 GND 0.005132f
C3292 a_188130_n13996.n105 GND 0.023688f
C3293 a_188130_n13996.n106 GND 0.030321f
C3294 a_188130_n13996.n107 GND 0.005132f
C3295 a_188130_n13996.t43 GND 0.064372f
C3296 a_188130_n13996.n108 GND 0.005434f
C3297 a_188130_n13996.n109 GND 0.005434f
C3298 a_188130_n13996.n110 GND 0.005434f
C3299 a_188130_n13996.n111 GND 0.005434f
C3300 a_188130_n13996.n112 GND 0.005434f
C3301 a_188130_n13996.n113 GND 5.99e-19
C3302 a_188130_n13996.n114 GND 0.005434f
C3303 a_188130_n13996.n115 GND 0.005434f
C3304 a_188130_n13996.n116 GND 0.005434f
C3305 a_188130_n13996.n117 GND 0.005434f
C3306 a_188130_n13996.n118 GND 0.005434f
C3307 a_188130_n13996.t15 GND 0.064372f
C3308 a_188130_n13996.n119 GND 0.119739f
C3309 a_188130_n13996.n120 GND 0.125843f
C3310 a_188130_n13996.n121 GND 0.137608f
C3311 a_188130_n13996.n122 GND 0.019178f
C3312 a_188130_n13996.n123 GND 0.005132f
C3313 a_188130_n13996.t13 GND 0.064372f
C3314 a_188130_n13996.n124 GND 0.009037f
C3315 a_188130_n13996.n125 GND 0.005434f
C3316 a_188130_n13996.n126 GND 0.005434f
C3317 a_188130_n13996.n127 GND 0.005434f
C3318 a_188130_n13996.n128 GND 0.005434f
C3319 a_188130_n13996.n129 GND 0.005434f
C3320 a_188130_n13996.n130 GND 5.99e-19
C3321 a_188130_n13996.n131 GND 0.005434f
C3322 a_188130_n13996.n132 GND 0.005434f
C3323 a_188130_n13996.n133 GND 0.005434f
C3324 a_188130_n13996.n134 GND 0.005434f
C3325 a_188130_n13996.n135 GND 0.005132f
C3326 a_188130_n13996.n136 GND 0.016538f
C3327 a_188130_n13996.n137 GND 0.038111f
C3328 a_188130_n13996.n138 GND 0.005434f
C3329 a_188130_n13996.n139 GND 0.017509f
C3330 a_188130_n13996.n140 GND 0.005434f
C3331 a_188130_n13996.n141 GND 0.04265f
C3332 a_188130_n13996.t7 GND 0.032791f
C3333 a_188130_n13996.n142 GND 0.013132f
C3334 a_188130_n13996.n143 GND 0.006711f
C3335 a_188130_n13996.n144 GND 0.005132f
C3336 a_188130_n13996.n145 GND 0.249138f
C3337 a_188130_n13996.n146 GND 0.014655f
C3338 a_188130_n13996.n147 GND 0.005132f
C3339 a_188130_n13996.n148 GND 0.005434f
C3340 a_188130_n13996.n149 GND 0.017509f
C3341 a_188130_n13996.n150 GND 0.017509f
C3342 a_188130_n13996.n151 GND 0.005434f
C3343 a_188130_n13996.n152 GND 0.005132f
C3344 a_188130_n13996.n153 GND 0.013908f
C3345 a_188130_n13996.n154 GND 0.014408f
C3346 a_188130_n13996.n155 GND 0.006562f
C3347 a_188130_n13996.n156 GND 0.284427f
C3348 a_188130_n13996.n157 GND 0.419527f
C3349 a_188130_n13996.n158 GND 0.005132f
C3350 a_188130_n13996.n159 GND 0.01892f
C3351 a_188130_n13996.n160 GND 0.005132f
C3352 a_188130_n13996.n161 GND 0.451349f
C3353 a_188130_n13996.n162 GND 0.005132f
C3354 a_188130_n13996.n163 GND 0.005132f
C3355 a_188130_n13996.n164 GND 0.019135f
C3356 a_188130_n13996.n165 GND 0.010115f
C3357 a_188130_n13996.n166 GND 0.019178f
C3358 a_188130_n13996.n167 GND 0.010115f
C3359 a_188130_n13996.n168 GND 0.019178f
C3360 a_188130_n13996.n169 GND 0.005132f
C3361 a_188130_n13996.n170 GND 0.019178f
C3362 a_188130_n13996.n171 GND 0.005132f
C3363 a_188130_n13996.n172 GND 0.019178f
C3364 a_188130_n13996.n173 GND 0.005132f
C3365 a_188130_n13996.n174 GND 0.019178f
C3366 a_188130_n13996.n175 GND 0.019178f
C3367 a_188130_n13996.n176 GND 0.005132f
C3368 a_188130_n13996.n177 GND 0.005434f
C3369 a_188130_n13996.t39 GND 0.064372f
C3370 a_188130_n13996.n178 GND 0.128744f
C3371 a_188130_n13996.n179 GND 0.009037f
C3372 a_188130_n13996.n180 GND 0.026434f
C3373 a_188130_n13996.n181 GND 0.030588f
C3374 a_188130_n13996.n182 GND 0.137608f
C3375 a_188130_n13996.n183 GND 0.137608f
C3376 a_188130_n13996.n184 GND 0.122514f
C3377 a_188130_n13996.n185 GND 0.122736f
C3378 a_188130_n13996.n186 GND 0.122514f
C3379 a_188130_n13996.n187 GND 0.137608f
C3380 a_188130_n13996.n188 GND 0.137608f
C3381 a_188130_n13996.n189 GND 0.137608f
C3382 a_188130_n13996.t42 GND 0.355184f
C3383 a_188130_n13996.n190 GND 0.257338f
C3384 a_188130_n13996.t6 GND 0.355362f
C3385 a_188130_n13996.n191 GND 0.371731f
C3386 a_188130_n13996.n192 GND 0.724054f
C3387 a_188130_n13996.t63 GND 0.355184f
C3388 a_188130_n13996.n193 GND 0.086163f
C3389 a_188130_n13996.t66 GND 0.355184f
C3390 a_188130_n13996.n194 GND 0.404244f
C3391 a_188130_n13996.n195 GND 0.137608f
C3392 a_188130_n13996.t59 GND 0.355184f
C3393 a_188130_n13996.n196 GND 0.131171f
C3394 a_188130_n13996.t60 GND 0.355184f
C3395 a_188130_n13996.n197 GND 0.137608f
C3396 a_188130_n13996.n198 GND 0.137608f
C3397 a_188130_n13996.t68 GND 0.355184f
C3398 a_188130_n13996.n199 GND 0.137608f
C3399 a_188130_n13996.t53 GND 0.355184f
C3400 a_188130_n13996.n200 GND 0.137608f
C3401 a_188130_n13996.n201 GND 0.137608f
C3402 a_188130_n13996.t56 GND 0.355184f
C3403 a_188130_n13996.n202 GND 0.137608f
C3404 a_188130_n13996.t61 GND 0.355184f
C3405 a_188130_n13996.n203 GND 0.137608f
C3406 a_188130_n13996.n204 GND 0.137608f
C3407 a_188130_n13996.t65 GND 0.355184f
C3408 a_188130_n13996.n205 GND 0.137608f
C3409 a_188130_n13996.t69 GND 0.355184f
C3410 a_188130_n13996.n206 GND 0.137608f
C3411 a_188130_n13996.n207 GND 0.137608f
C3412 a_188130_n13996.n208 GND 0.137608f
C3413 a_188130_n13996.n209 GND 0.137608f
C3414 a_188130_n13996.t8 GND 0.355184f
C3415 a_188130_n13996.t18 GND 0.355184f
C3416 a_188130_n13996.n210 GND 0.1254f
C3417 a_188130_n13996.n211 GND 0.26999f
C3418 a_188130_n13996.t30 GND 0.355305f
C3419 a_188130_n13996.n212 GND 0.739734f
C3420 a_188130_n13996.t51 GND 0.355184f
C3421 a_188130_n13996.n213 GND 0.086023f
C3422 a_188130_n13996.t62 GND 0.355184f
C3423 a_188130_n13996.n214 GND 0.404353f
C3424 a_188130_n13996.n215 GND 0.137608f
C3425 a_188130_n13996.t57 GND 0.355184f
C3426 a_188130_n13996.n216 GND 0.131393f
C3427 a_188130_n13996.t54 GND 0.355184f
C3428 a_188130_n13996.n217 GND 0.137608f
C3429 a_188130_n13996.n218 GND 0.137608f
C3430 a_188130_n13996.t52 GND 0.355184f
C3431 a_188130_n13996.n219 GND 0.137608f
C3432 a_188130_n13996.t49 GND 0.355184f
C3433 a_188130_n13996.n220 GND 0.137608f
C3434 a_188130_n13996.n221 GND 0.137608f
C3435 a_188130_n13996.t50 GND 0.355184f
C3436 a_188130_n13996.n222 GND 0.137608f
C3437 a_188130_n13996.t67 GND 0.355184f
C3438 a_188130_n13996.n223 GND 0.137608f
C3439 a_188130_n13996.n224 GND 0.137608f
C3440 a_188130_n13996.t64 GND 0.355184f
C3441 a_188130_n13996.n225 GND 0.137608f
C3442 a_188130_n13996.t58 GND 0.355184f
C3443 a_188130_n13996.n226 GND 0.137608f
C3444 a_188130_n13996.n227 GND 0.137608f
C3445 a_188130_n13996.t55 GND 0.355184f
C3446 a_188130_n13996.n228 GND 0.383331f
C3447 a_188130_n13996.n229 GND 0.137608f
C3448 a_188130_n13996.t40 GND 0.355184f
C3449 a_188130_n13996.n230 GND 0.137608f
C3450 a_188130_n13996.n231 GND 0.137608f
C3451 a_188130_n13996.t4 GND 0.355184f
C3452 a_188130_n13996.n232 GND 0.137608f
C3453 a_188130_n13996.t16 GND 0.355184f
C3454 a_188130_n13996.n233 GND 0.137608f
C3455 a_188130_n13996.n234 GND 0.137608f
C3456 a_188130_n13996.t22 GND 0.355185f
C3457 a_188130_n13996.n235 GND 0.383331f
C3458 a_188130_n13996.t36 GND 0.355184f
C3459 a_188130_n13996.n236 GND 0.122736f
C3460 a_188130_n13996.n237 GND 0.137608f
C3461 a_188130_n13996.t44 GND 0.355184f
C3462 a_188130_n13996.n238 GND 0.137608f
C3463 a_188130_n13996.t10 GND 0.355184f
C3464 a_188130_n13996.n239 GND 0.137608f
C3465 a_188130_n13996.n240 GND 0.137608f
C3466 a_188130_n13996.t20 GND 0.355184f
C3467 a_188130_n13996.n241 GND 0.137608f
C3468 a_188130_n13996.t26 GND 0.355184f
C3469 a_188130_n13996.n242 GND 0.137608f
C3470 a_188130_n13996.n243 GND 0.125178f
C3471 a_188130_n13996.t38 GND 0.355184f
C3472 a_188130_n13996.n244 GND 0.125178f
C3473 a_188130_n13996.n245 GND 0.030321f
C3474 a_188130_n13996.t12 GND 0.355184f
C3475 a_188130_n13996.n246 GND 0.125843f
C3476 a_188130_n13996.n247 GND 0.125622f
C3477 a_188130_n13996.t14 GND 0.355184f
C3478 a_188130_n13996.n248 GND 0.128951f
C3479 a_188130_n13996.n249 GND 0.027258f
C3480 a_188130_n13996.n250 GND 0.023104f
C3481 a_188130_n13996.n251 GND 0.005132f
C3482 a_188130_n13996.n252 GND 0.01892f
C3483 a_188130_n13996.n253 GND 0.005132f
C3484 a_188130_n13996.n254 GND 0.016538f
C3485 a_188130_n13996.n255 GND 0.005132f
C3486 a_188130_n13996.n256 GND 0.005132f
C3487 a_188130_n13996.n257 GND 0.019135f
C3488 a_188130_n13996.n258 GND 0.010115f
C3489 a_188130_n13996.n259 GND 0.019178f
C3490 a_188130_n13996.n260 GND 0.010115f
C3491 a_188130_n13996.n261 GND 0.019178f
C3492 a_188130_n13996.n262 GND 0.005132f
C3493 a_188130_n13996.n263 GND 0.019178f
C3494 a_188130_n13996.n264 GND 0.005132f
C3495 a_188130_n13996.n265 GND 0.019178f
C3496 a_188130_n13996.n266 GND 0.005132f
C3497 a_188130_n13996.n267 GND 0.019178f
C3498 a_188130_n13996.n268 GND 0.005132f
C3499 a_188130_n13996.n269 GND 0.019178f
C3500 a_188130_n13996.n270 GND 0.019178f
C3501 a_188130_n13996.n271 GND 0.005132f
C3502 a_188130_n13996.n272 GND 0.009037f
C3503 a_188130_n13996.n273 GND 0.128744f
C3504 a_188130_n13996.n274 GND 0.009037f
C3505 a_188130_n13996.n275 GND 0.023688f
C3506 a_188130_n13996.n276 GND 1.29341f
C3507 a_188130_n13996.n277 GND 0.031711f
C3508 a_188130_n13996.n278 GND 0.005434f
C3509 a_188130_n13996.n279 GND 0.013534f
C3510 a_188130_n13996.n280 GND 0.005132f
C3511 a_188130_n13996.n281 GND 0.017509f
C3512 a_188130_n13996.n282 GND 0.005434f
C3513 a_188130_n13996.n283 GND 0.041602f
C3514 a_188130_n13996.t2 GND 0.025132f
C3515 a_188130_n13996.n284 GND 0.013132f
C3516 a_188130_n13996.n285 GND 0.00637f
C3517 a_188130_n13996.n286 GND 0.005132f
C3518 a_188130_n13996.n287 GND 0.257889f
C3519 a_188130_n13996.n288 GND 0.005132f
C3520 a_188130_n13996.n289 GND 0.005434f
C3521 a_188130_n13996.n290 GND 0.017509f
C3522 a_188130_n13996.n291 GND 0.017509f
C3523 a_188130_n13996.n292 GND 0.005434f
C3524 a_188130_n13996.n293 GND 0.005132f
C3525 a_188130_n13996.n294 GND 0.014703f
C3526 a_188130_n13996.n295 GND 0.014481f
C3527 a_188130_n13996.n296 GND 0.006383f
C3528 a_188130_n13996.n297 GND 0.235578f
C3529 a_188130_n13996.t1 GND 0.064372f
C3530 a_188130_n13996.n298 GND 0.005434f
C3531 a_188130_n13996.n299 GND 0.005434f
C3532 a_188130_n13996.n300 GND 0.006731f
C3533 a_188130_n13996.n301 GND 0.014481f
C3534 a_188130_n13996.n302 GND 0.005132f
C3535 a_188130_n13996.n303 GND 0.014703f
C3536 a_188130_n13996.n304 GND 0.013534f
C3537 a_188130_n13996.n305 GND 0.011983f
C3538 a_188130_n13996.n306 GND 0.00956f
C3539 a_188130_n13996.t47 GND 0.064372f
C3540 a_188130_n13996.n307 GND 0.138f
C3541 a_188130_n13996.n308 GND 0.235578f
C3542 a_188130_n13996.t46 GND 0.064372f
C3543 a_188130_n13996.n309 GND 0.005434f
C3544 a_188130_n13996.n310 GND 0.005434f
C3545 a_188130_n13996.n311 GND 0.006731f
C3546 a_188130_n13996.n312 GND 0.014481f
C3547 a_188130_n13996.n313 GND 0.005132f
C3548 a_188130_n13996.n314 GND 0.014703f
C3549 a_188130_n13996.n315 GND 0.013534f
C3550 a_188130_n13996.n316 GND 0.011983f
C3551 a_188130_n13996.n317 GND 0.00956f
C3552 a_188130_n13996.t0 GND 0.064372f
C3553 a_188130_n13996.n318 GND 0.138f
C3554 a_188130_n13996.n319 GND 0.235578f
C3555 a_188130_n13996.t48 GND 0.064372f
C3556 a_188130_n13996.n320 GND 0.005434f
C3557 a_188130_n13996.n321 GND 0.005434f
C3558 a_188130_n13996.n322 GND 0.006731f
C3559 a_188130_n13996.n323 GND 0.014481f
C3560 a_188130_n13996.n324 GND 0.005132f
C3561 a_188130_n13996.n325 GND 0.014703f
C3562 a_188130_n13996.n326 GND 0.013534f
C3563 a_188130_n13996.n327 GND 0.011983f
C3564 a_188130_n13996.n328 GND 0.00956f
C3565 a_188130_n13996.t3 GND 0.064372f
C3566 a_188130_n13996.n329 GND 0.138f
C3567 a_188130_n13996.n330 GND 1.29287f
C3568 a_188130_n13996.n331 GND 0.084714f
C3569 a_188130_n13996.n332 GND 0.005132f
C3570 a_188130_n13996.n333 GND 0.005132f
C3571 a_188130_n13996.n334 GND 0.019135f
C3572 a_188130_n13996.n335 GND 0.010115f
C3573 a_188130_n13996.n336 GND 0.019178f
C3574 a_188130_n13996.n337 GND 0.010115f
C3575 a_188130_n13996.n338 GND 0.019178f
C3576 a_188130_n13996.n339 GND 0.005132f
C3577 a_188130_n13996.n340 GND 0.019178f
C3578 a_188130_n13996.n341 GND 0.005132f
C3579 a_188130_n13996.n342 GND 0.019178f
C3580 a_188130_n13996.n343 GND 0.005132f
C3581 a_188130_n13996.n344 GND 0.019178f
C3582 a_188130_n13996.n345 GND 0.019178f
C3583 a_188130_n13996.n346 GND 0.005132f
C3584 a_188130_n13996.n347 GND 0.005434f
C3585 a_188130_n13996.t19 GND 0.064372f
C3586 a_188130_n13996.n348 GND 0.128744f
C3587 a_188130_n13996.n349 GND 0.009037f
C3588 a_188130_n13996.n350 GND 0.026434f
C3589 a_188130_n13996.n351 GND 0.030588f
C3590 a_188130_n13996.n352 GND 0.125622f
C3591 a_188130_n13996.t24 GND 0.355184f
C3592 a_188130_n13996.n353 GND 0.125622f
C3593 a_188130_n13996.t28 GND 0.355184f
C3594 a_188130_n13996.n354 GND 0.125843f
C3595 a_188130_n13996.n355 GND 0.023688f
C3596 a_188130_n13996.n356 GND 0.030321f
C3597 a_188130_n13996.n357 GND 0.125178f
C3598 a_188130_n13996.t34 GND 0.355184f
C3599 a_188130_n13996.n358 GND 0.125178f
C3600 a_188130_n13996.n359 GND 0.030588f
C3601 a_188130_n13996.n360 GND 0.026434f
C3602 a_188130_n13996.n361 GND 0.005132f
C3603 a_188130_n13996.n362 GND 0.019135f
C3604 a_188130_n13996.n363 GND 0.010115f
C3605 a_188130_n13996.n364 GND 0.019178f
C3606 a_188130_n13996.n365 GND 0.010115f
C3607 a_188130_n13996.n366 GND 0.019178f
C3608 a_188130_n13996.n367 GND 0.005132f
C3609 a_188130_n13996.n368 GND 0.019178f
C3610 a_188130_n13996.n369 GND 0.005132f
C3611 a_188130_n13996.n370 GND 0.019178f
C3612 a_188130_n13996.n371 GND 0.005132f
C3613 a_188130_n13996.n372 GND 0.019178f
C3614 a_188130_n13996.n373 GND 0.005132f
C3615 a_188130_n13996.n374 GND 0.019178f
C3616 a_188130_n13996.n375 GND 0.019178f
C3617 a_188130_n13996.n376 GND 0.005132f
C3618 a_188130_n13996.n377 GND 0.009037f
C3619 a_188130_n13996.n378 GND 0.128744f
C3620 a_188130_n13996.n379 GND 0.005434f
C3621 a_188130_n13996.n380 GND 0.005132f
C3622 a_188130_n13996.n381 GND 0.016538f
C3623 a_188130_n13996.n382 GND 0.451349f
C3624 a_188130_n13996.t41 GND 0.064372f
C3625 a_188130_n13996.n383 GND 0.005434f
C3626 a_188130_n13996.n384 GND 0.006774f
C3627 a_188130_n13996.n385 GND 0.014408f
C3628 a_188130_n13996.n386 GND 0.013908f
C3629 a_188130_n13996.n387 GND 0.011863f
C3630 a_188130_n13996.n388 GND 0.011644f
C3631 a_188130_n13996.t33 GND 0.064372f
C3632 a_188130_n13996.n389 GND 0.132696f
C3633 a_188130_n13996.n390 GND 0.451349f
C3634 a_188130_n13996.t17 GND 0.064372f
C3635 a_188130_n13996.n391 GND 0.005434f
C3636 a_188130_n13996.n392 GND 0.006774f
C3637 a_188130_n13996.n393 GND 0.014408f
C3638 a_188130_n13996.n394 GND 0.013908f
C3639 a_188130_n13996.n395 GND 0.011863f
C3640 a_188130_n13996.n396 GND 0.011644f
C3641 a_188130_n13996.t5 GND 0.064372f
C3642 a_188130_n13996.n397 GND 0.132696f
C3643 a_188130_n13996.n398 GND 0.451349f
C3644 a_188130_n13996.t37 GND 0.064372f
C3645 a_188130_n13996.n399 GND 0.005434f
C3646 a_188130_n13996.n400 GND 0.006774f
C3647 a_188130_n13996.n401 GND 0.014408f
C3648 a_188130_n13996.n402 GND 0.013908f
C3649 a_188130_n13996.n403 GND 0.011863f
C3650 a_188130_n13996.n404 GND 0.011644f
C3651 a_188130_n13996.t23 GND 0.064372f
C3652 a_188130_n13996.n405 GND 0.132696f
C3653 a_188130_n13996.n406 GND 0.458009f
C3654 a_188130_n13996.n407 GND 0.451349f
C3655 a_188130_n13996.n408 GND 0.132696f
C3656 a_188130_n13996.t45 GND 0.064372f
C3657 a_219318_n20038.n0 GND 4.24325f
C3658 a_219318_n20038.n1 GND 4.4759f
C3659 a_219318_n20038.n2 GND 0.037893f
C3660 a_219318_n20038.n3 GND 0.03785f
C3661 a_219318_n20038.n4 GND 1.11132f
C3662 a_219318_n20038.n5 GND 0.886457f
C3663 a_219318_n20038.n6 GND 1.11089f
C3664 a_219318_n20038.n7 GND 0.178901f
C3665 a_219318_n20038.n8 GND 0.00431f
C3666 a_219318_n20038.n9 GND 0.178901f
C3667 a_219318_n20038.n10 GND 0.00431f
C3668 a_219318_n20038.n11 GND 0.178901f
C3669 a_219318_n20038.n12 GND 0.00431f
C3670 a_219318_n20038.n13 GND 0.178842f
C3671 a_219318_n20038.n14 GND 0.004341f
C3672 a_219318_n20038.n15 GND 0.178842f
C3673 a_219318_n20038.n16 GND 0.004341f
C3674 a_219318_n20038.n17 GND 0.178842f
C3675 a_219318_n20038.n18 GND 0.004341f
C3676 a_219318_n20038.n19 GND 0.822848f
C3677 a_219318_n20038.n20 GND 0.822419f
C3678 a_219318_n20038.n21 GND 0.044851f
C3679 a_219318_n20038.n22 GND 0.00704f
C3680 a_219318_n20038.n23 GND 0.044851f
C3681 a_219318_n20038.n24 GND 0.00704f
C3682 a_219318_n20038.n25 GND 0.044851f
C3683 a_219318_n20038.n26 GND 0.00704f
C3684 a_219318_n20038.n27 GND 0.049872f
C3685 a_219318_n20038.n28 GND 0.020924f
C3686 a_219318_n20038.n29 GND 0.041664f
C3687 a_219318_n20038.n30 GND 0.020925f
C3688 a_219318_n20038.n31 GND 0.044876f
C3689 a_219318_n20038.n32 GND 0.00704f
C3690 a_219318_n20038.n33 GND 0.044876f
C3691 a_219318_n20038.n34 GND 0.00704f
C3692 a_219318_n20038.n35 GND 0.044876f
C3693 a_219318_n20038.n36 GND 0.00704f
C3694 a_219318_n20038.n37 GND 0.044876f
C3695 a_219318_n20038.n38 GND 0.00704f
C3696 a_219318_n20038.n39 GND 0.044876f
C3697 a_219318_n20038.n40 GND 0.00704f
C3698 a_219318_n20038.n41 GND 0.044876f
C3699 a_219318_n20038.n42 GND 0.00704f
C3700 a_219318_n20038.n43 GND 0.020925f
C3701 a_219318_n20038.n44 GND 0.041664f
C3702 a_219318_n20038.n45 GND 0.04992f
C3703 a_219318_n20038.n46 GND 0.020926f
C3704 a_219318_n20038.n47 GND 0.0449f
C3705 a_219318_n20038.n48 GND 0.007041f
C3706 a_219318_n20038.n49 GND 0.0449f
C3707 a_219318_n20038.n50 GND 0.007041f
C3708 a_219318_n20038.n51 GND 0.004596f
C3709 a_219318_n20038.n52 GND 0.007041f
C3710 a_219318_n20038.n53 GND 0.0449f
C3711 a_219318_n20038.n54 GND 0.020996f
C3712 a_219318_n20038.n55 GND 0.192656f
C3713 a_219318_n20038.n56 GND 0.00585f
C3714 a_219318_n20038.n57 GND 0.192656f
C3715 a_219318_n20038.n58 GND 0.00585f
C3716 a_219318_n20038.n59 GND 0.192656f
C3717 a_219318_n20038.n60 GND 0.00585f
C3718 a_219318_n20038.n61 GND 0.192656f
C3719 a_219318_n20038.n62 GND 0.00585f
C3720 a_219318_n20038.n63 GND 0.192656f
C3721 a_219318_n20038.n64 GND 0.00585f
C3722 a_219318_n20038.n65 GND 0.192656f
C3723 a_219318_n20038.n66 GND 0.00585f
C3724 a_219318_n20038.n67 GND 0.0096f
C3725 a_219318_n20038.n68 GND 0.020996f
C3726 a_219318_n20038.t20 GND 0.043954f
C3727 a_219318_n20038.n69 GND 0.00371f
C3728 a_219318_n20038.n70 GND 0.007982f
C3729 a_219318_n20038.n71 GND 0.01004f
C3730 a_219318_n20038.t22 GND 0.043954f
C3731 a_219318_n20038.t21 GND 0.043954f
C3732 a_219318_n20038.n72 GND 0.095056f
C3733 a_219318_n20038.n73 GND 0.00371f
C3734 a_219318_n20038.n74 GND 0.004596f
C3735 a_219318_n20038.n75 GND 0.009838f
C3736 a_219318_n20038.n76 GND 0.01004f
C3737 a_219318_n20038.n77 GND 0.007982f
C3738 a_219318_n20038.t4 GND 0.043954f
C3739 a_219318_n20038.n78 GND 0.00371f
C3740 a_219318_n20038.n79 GND 0.004596f
C3741 a_219318_n20038.n80 GND 0.009888f
C3742 a_219318_n20038.n81 GND 0.007981f
C3743 a_219318_n20038.n82 GND 0.01004f
C3744 a_219318_n20038.t1 GND 0.043954f
C3745 a_219318_n20038.n83 GND 0.095083f
C3746 a_219318_n20038.n84 GND 0.01004f
C3747 a_219318_n20038.n85 GND 0.00371f
C3748 a_219318_n20038.n86 GND 0.003504f
C3749 a_219318_n20038.n87 GND 0.0096f
C3750 a_219318_n20038.n88 GND 0.004358f
C3751 a_219318_n20038.n89 GND 0.003504f
C3752 a_219318_n20038.n90 GND 0.00371f
C3753 a_219318_n20038.n91 GND 0.021652f
C3754 a_219318_n20038.n92 GND 0.011955f
C3755 a_219318_n20038.n93 GND 0.008967f
C3756 a_219318_n20038.n94 GND 0.00435f
C3757 a_219318_n20038.t0 GND 0.01716f
C3758 a_219318_n20038.n95 GND 0.028406f
C3759 a_219318_n20038.n96 GND 0.176291f
C3760 a_219318_n20038.n97 GND 0.003504f
C3761 a_219318_n20038.n98 GND 0.00371f
C3762 a_219318_n20038.n99 GND 0.011955f
C3763 a_219318_n20038.n100 GND 0.011955f
C3764 a_219318_n20038.n101 GND 0.00371f
C3765 a_219318_n20038.n102 GND 0.003504f
C3766 a_219318_n20038.n103 GND 0.009676f
C3767 a_219318_n20038.t14 GND 0.043954f
C3768 a_219318_n20038.n104 GND 0.00371f
C3769 a_219318_n20038.n105 GND 0.004596f
C3770 a_219318_n20038.n106 GND 0.009888f
C3771 a_219318_n20038.n107 GND 0.007981f
C3772 a_219318_n20038.n108 GND 0.01004f
C3773 a_219318_n20038.t2 GND 0.043954f
C3774 a_219318_n20038.n109 GND 0.095083f
C3775 a_219318_n20038.t11 GND 0.043954f
C3776 a_219318_n20038.n110 GND 0.00371f
C3777 a_219318_n20038.n111 GND 0.004596f
C3778 a_219318_n20038.n112 GND 0.009888f
C3779 a_219318_n20038.n113 GND 0.007981f
C3780 a_219318_n20038.n114 GND 0.01004f
C3781 a_219318_n20038.t17 GND 0.043954f
C3782 a_219318_n20038.n115 GND 0.095083f
C3783 a_219318_n20038.n116 GND 0.021652f
C3784 a_219318_n20038.n117 GND 0.00371f
C3785 a_219318_n20038.n118 GND 0.003504f
C3786 a_219318_n20038.n119 GND 0.011955f
C3787 a_219318_n20038.n120 GND 0.00371f
C3788 a_219318_n20038.n121 GND 0.028406f
C3789 a_219318_n20038.t15 GND 0.01716f
C3790 a_219318_n20038.n122 GND 0.008967f
C3791 a_219318_n20038.n123 GND 0.00435f
C3792 a_219318_n20038.n124 GND 0.003504f
C3793 a_219318_n20038.n125 GND 0.176089f
C3794 a_219318_n20038.n126 GND 0.003504f
C3795 a_219318_n20038.n127 GND 0.00371f
C3796 a_219318_n20038.n128 GND 0.011955f
C3797 a_219318_n20038.n129 GND 0.011955f
C3798 a_219318_n20038.n130 GND 0.00371f
C3799 a_219318_n20038.n131 GND 0.003504f
C3800 a_219318_n20038.n132 GND 0.01004f
C3801 a_219318_n20038.n133 GND 0.009888f
C3802 a_219318_n20038.n134 GND 0.004358f
C3803 a_219318_n20038.n135 GND 1.29665f
C3804 a_219318_n20038.n136 GND 0.004358f
C3805 a_219318_n20038.n137 GND 0.011955f
C3806 a_219318_n20038.n138 GND 0.00371f
C3807 a_219318_n20038.n139 GND 0.176291f
C3808 a_219318_n20038.n140 GND 0.003504f
C3809 a_219318_n20038.n141 GND 0.011955f
C3810 a_219318_n20038.t12 GND 0.01716f
C3811 a_219318_n20038.n142 GND 0.028406f
C3812 a_219318_n20038.n143 GND 0.00435f
C3813 a_219318_n20038.n144 GND 0.008967f
C3814 a_219318_n20038.n145 GND 0.011955f
C3815 a_219318_n20038.n146 GND 0.00371f
C3816 a_219318_n20038.n147 GND 0.003504f
C3817 a_219318_n20038.n148 GND 0.01004f
C3818 a_219318_n20038.n149 GND 0.009676f
C3819 a_219318_n20038.n150 GND 0.003504f
C3820 a_219318_n20038.n151 GND 0.00371f
C3821 a_219318_n20038.n152 GND 0.003504f
C3822 a_219318_n20038.n153 GND 0.00371f
C3823 a_219318_n20038.n154 GND 0.021652f
C3824 a_219318_n20038.t16 GND 0.043954f
C3825 a_219318_n20038.t26 GND 0.043954f
C3826 a_219318_n20038.n155 GND 0.097484f
C3827 a_219318_n20038.n156 GND 0.0096f
C3828 a_219318_n20038.n157 GND 0.008866f
C3829 a_219318_n20038.t10 GND 0.043954f
C3830 a_219318_n20038.t27 GND 0.043954f
C3831 a_219318_n20038.n158 GND 0.097484f
C3832 a_219318_n20038.n159 GND 0.0096f
C3833 a_219318_n20038.n160 GND 0.008866f
C3834 a_219318_n20038.t8 GND 0.043954f
C3835 a_219318_n20038.t7 GND 0.043954f
C3836 a_219318_n20038.n161 GND 0.097484f
C3837 a_219318_n20038.n162 GND 0.0096f
C3838 a_219318_n20038.n163 GND 0.008866f
C3839 a_219318_n20038.t13 GND 0.043954f
C3840 a_219318_n20038.t5 GND 0.043954f
C3841 a_219318_n20038.n164 GND 0.097484f
C3842 a_219318_n20038.n165 GND 0.0096f
C3843 a_219318_n20038.n166 GND 0.008866f
C3844 a_219318_n20038.t6 GND 0.043954f
C3845 a_219318_n20038.t9 GND 0.043954f
C3846 a_219318_n20038.n167 GND 0.097484f
C3847 a_219318_n20038.n168 GND 0.0096f
C3848 a_219318_n20038.n169 GND 0.008866f
C3849 a_219318_n20038.t25 GND 0.043954f
C3850 a_219318_n20038.t3 GND 0.043954f
C3851 a_219318_n20038.n170 GND 0.097484f
C3852 a_219318_n20038.n171 GND 0.0096f
C3853 a_219318_n20038.n172 GND 0.008866f
C3854 a_219318_n20038.n173 GND 1.29273f
C3855 a_219318_n20038.n174 GND 0.176046f
C3856 a_219318_n20038.n175 GND 0.00371f
C3857 a_219318_n20038.n176 GND 0.003504f
C3858 a_219318_n20038.n177 GND 0.021652f
C3859 a_219318_n20038.n178 GND 0.00371f
C3860 a_219318_n20038.n179 GND 0.004358f
C3861 a_219318_n20038.n180 GND 0.009838f
C3862 a_219318_n20038.n181 GND 0.01004f
C3863 a_219318_n20038.n182 GND 0.003504f
C3864 a_219318_n20038.n183 GND 0.003504f
C3865 a_219318_n20038.n184 GND 0.00371f
C3866 a_219318_n20038.n185 GND 0.011955f
C3867 a_219318_n20038.n186 GND 0.011955f
C3868 a_219318_n20038.t23 GND 0.01716f
C3869 a_219318_n20038.n187 GND 0.028406f
C3870 a_219318_n20038.n188 GND 0.00435f
C3871 a_219318_n20038.n189 GND 0.008967f
C3872 a_219318_n20038.n190 GND 0.011955f
C3873 a_219318_n20038.n191 GND 0.00371f
C3874 a_219318_n20038.n192 GND 0.003504f
C3875 a_219318_n20038.t19 GND 0.043954f
C3876 a_219318_n20038.t18 GND 0.043954f
C3877 a_219318_n20038.n193 GND 0.095056f
C3878 a_219318_n20038.n194 GND 0.00371f
C3879 a_219318_n20038.n195 GND 0.004596f
C3880 a_219318_n20038.n196 GND 0.009838f
C3881 a_219318_n20038.n197 GND 0.01004f
C3882 a_219318_n20038.n198 GND 0.007982f
C3883 a_219318_n20038.n199 GND 0.009838f
C3884 a_219318_n20038.n200 GND 0.095056f
C3885 a_219318_n20038.t24 GND 0.043954f
C3886 VREFP.t44 GND 0.061503f
C3887 VREFP.t52 GND 0.015089f
C3888 VREFP.t50 GND 0.015089f
C3889 VREFP.n0 GND 0.040781f
C3890 VREFP.n1 GND 0.145665f
C3891 VREFP.t53 GND 0.015089f
C3892 VREFP.t54 GND 0.015089f
C3893 VREFP.n2 GND 0.040865f
C3894 VREFP.n3 GND 0.072232f
C3895 VREFP.t41 GND 0.015089f
C3896 VREFP.t55 GND 0.015089f
C3897 VREFP.n4 GND 0.040781f
C3898 VREFP.n5 GND 0.072133f
C3899 VREFP.t43 GND 0.015089f
C3900 VREFP.t42 GND 0.015089f
C3901 VREFP.n6 GND 0.040781f
C3902 VREFP.n7 GND 0.071219f
C3903 VREFP.t51 GND 0.015089f
C3904 VREFP.t49 GND 0.015089f
C3905 VREFP.n8 GND 0.040865f
C3906 VREFP.n9 GND 0.072232f
C3907 VREFP.t38 GND 0.015089f
C3908 VREFP.t37 GND 0.015089f
C3909 VREFP.n10 GND 0.040781f
C3910 VREFP.n11 GND 0.071219f
C3911 VREFP.t45 GND 0.015089f
C3912 VREFP.t39 GND 0.015089f
C3913 VREFP.n12 GND 0.040865f
C3914 VREFP.n13 GND 0.072232f
C3915 VREFP.t46 GND 0.015089f
C3916 VREFP.t40 GND 0.015089f
C3917 VREFP.n14 GND 0.040781f
C3918 VREFP.n15 GND 0.072133f
C3919 VREFP.t48 GND 0.015089f
C3920 VREFP.t47 GND 0.015089f
C3921 VREFP.n16 GND 0.040781f
C3922 VREFP.n17 GND 0.158624f
C3923 VREFP.t23 GND 0.015089f
C3924 VREFP.t22 GND 0.015089f
C3925 VREFP.n18 GND 0.054092f
C3926 VREFP.t26 GND 0.015089f
C3927 VREFP.t24 GND 0.015089f
C3928 VREFP.n19 GND 0.053395f
C3929 VREFP.n20 GND 0.109318f
C3930 VREFP.t27 GND 0.015089f
C3931 VREFP.t25 GND 0.015089f
C3932 VREFP.n21 GND 0.05358f
C3933 VREFP.n22 GND 0.057246f
C3934 VREFP.t20 GND 0.015089f
C3935 VREFP.t28 GND 0.015089f
C3936 VREFP.n23 GND 0.053395f
C3937 VREFP.n24 GND 0.057248f
C3938 VREFP.t21 GND 0.070551f
C3939 VREFP.n25 GND 0.180661f
C3940 VREFP.n26 GND 0.174567f
C3941 VREFP.n27 GND 0.058754f
C3942 VREFP.t3 GND 0.015089f
C3943 VREFP.t0 GND 0.015089f
C3944 VREFP.n28 GND 0.054092f
C3945 VREFP.t2 GND 0.015089f
C3946 VREFP.t32 GND 0.015089f
C3947 VREFP.n29 GND 0.053395f
C3948 VREFP.n30 GND 0.109318f
C3949 VREFP.t1 GND 0.015089f
C3950 VREFP.t34 GND 0.015089f
C3951 VREFP.n31 GND 0.05358f
C3952 VREFP.n32 GND 0.057246f
C3953 VREFP.t35 GND 0.015089f
C3954 VREFP.t36 GND 0.015089f
C3955 VREFP.n33 GND 0.053395f
C3956 VREFP.n34 GND 0.057248f
C3957 VREFP.t33 GND 0.070551f
C3958 VREFP.n35 GND 0.122365f
C3959 VREFP.t10 GND 0.061438f
C3960 VREFP.n36 GND 0.078448f
C3961 VREFP.t11 GND 0.015089f
C3962 VREFP.t19 GND 0.015089f
C3963 VREFP.n37 GND 0.040781f
C3964 VREFP.n38 GND 0.066929f
C3965 VREFP.t9 GND 0.015089f
C3966 VREFP.t18 GND 0.015089f
C3967 VREFP.n39 GND 0.040865f
C3968 VREFP.n40 GND 0.072424f
C3969 VREFP.t12 GND 0.015089f
C3970 VREFP.t5 GND 0.015089f
C3971 VREFP.n41 GND 0.040781f
C3972 VREFP.n42 GND 0.072316f
C3973 VREFP.t7 GND 0.015089f
C3974 VREFP.t13 GND 0.015089f
C3975 VREFP.n43 GND 0.040781f
C3976 VREFP.n44 GND 0.071411f
C3977 VREFP.t15 GND 0.015089f
C3978 VREFP.t30 GND 0.015089f
C3979 VREFP.n45 GND 0.040865f
C3980 VREFP.n46 GND 0.072424f
C3981 VREFP.t4 GND 0.015089f
C3982 VREFP.t17 GND 0.015089f
C3983 VREFP.n47 GND 0.040781f
C3984 VREFP.n48 GND 0.065255f
C3985 VREFP.n49 GND 0.00742f
C3986 VREFP.t6 GND 0.015089f
C3987 VREFP.t16 GND 0.015089f
C3988 VREFP.n50 GND 0.040865f
C3989 VREFP.n51 GND 0.070433f
C3990 VREFP.t31 GND 0.015089f
C3991 VREFP.t8 GND 0.015089f
C3992 VREFP.n52 GND 0.040781f
C3993 VREFP.n53 GND 0.072316f
C3994 VREFP.t14 GND 0.015089f
C3995 VREFP.t29 GND 0.015089f
C3996 VREFP.n54 GND 0.040781f
C3997 VREFP.n55 GND 0.159109f
C3998 VREFP.n56 GND 0.173651f
C3999 VREFP.n57 GND 0.527876f
C4000 VREFP.n58 GND 15.450299f
C4001 1Bit_DAC_0.OUT.t36 GND 0.307164f
C4002 1Bit_DAC_0.OUT.t32 GND 0.07449f
C4003 1Bit_DAC_0.OUT.t37 GND 0.07449f
C4004 1Bit_DAC_0.OUT.n0 GND 0.205453f
C4005 1Bit_DAC_0.OUT.n1 GND 1.05005f
C4006 1Bit_DAC_0.OUT.t56 GND 0.07449f
C4007 1Bit_DAC_0.OUT.t40 GND 0.07449f
C4008 1Bit_DAC_0.OUT.n2 GND 0.205655f
C4009 1Bit_DAC_0.OUT.n3 GND 0.521729f
C4010 1Bit_DAC_0.OUT.t38 GND 0.07449f
C4011 1Bit_DAC_0.OUT.t50 GND 0.07449f
C4012 1Bit_DAC_0.OUT.n4 GND 0.205453f
C4013 1Bit_DAC_0.OUT.n5 GND 0.516965f
C4014 1Bit_DAC_0.OUT.t48 GND 0.07449f
C4015 1Bit_DAC_0.OUT.t45 GND 0.07449f
C4016 1Bit_DAC_0.OUT.n6 GND 0.205453f
C4017 1Bit_DAC_0.OUT.n7 GND 0.530509f
C4018 1Bit_DAC_0.OUT.t44 GND 0.07449f
C4019 1Bit_DAC_0.OUT.t41 GND 0.07449f
C4020 1Bit_DAC_0.OUT.n8 GND 0.205576f
C4021 1Bit_DAC_0.OUT.n9 GND 0.530836f
C4022 1Bit_DAC_0.OUT.t53 GND 0.07449f
C4023 1Bit_DAC_0.OUT.t51 GND 0.07449f
C4024 1Bit_DAC_0.OUT.n10 GND 0.205576f
C4025 1Bit_DAC_0.OUT.n11 GND 0.530836f
C4026 1Bit_DAC_0.OUT.t52 GND 0.07449f
C4027 1Bit_DAC_0.OUT.t30 GND 0.07449f
C4028 1Bit_DAC_0.OUT.n12 GND 0.205453f
C4029 1Bit_DAC_0.OUT.n13 GND 0.530509f
C4030 1Bit_DAC_0.OUT.t39 GND 0.07449f
C4031 1Bit_DAC_0.OUT.t31 GND 0.07449f
C4032 1Bit_DAC_0.OUT.n14 GND 0.205655f
C4033 1Bit_DAC_0.OUT.n15 GND 0.514957f
C4034 1Bit_DAC_0.OUT.t33 GND 0.07449f
C4035 1Bit_DAC_0.OUT.t43 GND 0.07449f
C4036 1Bit_DAC_0.OUT.n16 GND 0.205453f
C4037 1Bit_DAC_0.OUT.n17 GND 0.513579f
C4038 1Bit_DAC_0.OUT.t26 GND 0.07449f
C4039 1Bit_DAC_0.OUT.t7 GND 0.07449f
C4040 1Bit_DAC_0.OUT.n18 GND 0.266112f
C4041 1Bit_DAC_0.OUT.t5 GND 0.07449f
C4042 1Bit_DAC_0.OUT.t17 GND 0.07449f
C4043 1Bit_DAC_0.OUT.n19 GND 0.267961f
C4044 1Bit_DAC_0.OUT.n20 GND 0.860037f
C4045 1Bit_DAC_0.OUT.t23 GND 0.07449f
C4046 1Bit_DAC_0.OUT.t4 GND 0.07449f
C4047 1Bit_DAC_0.OUT.n21 GND 0.267728f
C4048 1Bit_DAC_0.OUT.n22 GND 0.40382f
C4049 1Bit_DAC_0.OUT.t3 GND 0.07449f
C4050 1Bit_DAC_0.OUT.t25 GND 0.07449f
C4051 1Bit_DAC_0.OUT.n23 GND 0.267961f
C4052 1Bit_DAC_0.OUT.n24 GND 0.404038f
C4053 1Bit_DAC_0.OUT.t6 GND 0.347549f
C4054 1Bit_DAC_0.OUT.n25 GND 0.424447f
C4055 1Bit_DAC_0.OUT.n26 GND 0.216698f
C4056 1Bit_DAC_0.OUT.t2 GND 0.07449f
C4057 1Bit_DAC_0.OUT.t0 GND 0.07449f
C4058 1Bit_DAC_0.OUT.n27 GND 0.206276f
C4059 1Bit_DAC_0.OUT.t28 GND 4.85035f
C4060 1Bit_DAC_0.OUT.t12 GND 0.07449f
C4061 1Bit_DAC_0.OUT.t8 GND 0.07449f
C4062 1Bit_DAC_0.OUT.n28 GND 0.205818f
C4063 1Bit_DAC_0.OUT.n29 GND 24.4948f
C4064 1Bit_DAC_0.OUT.n30 GND 0.810859f
C4065 1Bit_DAC_0.OUT.t13 GND 0.07449f
C4066 1Bit_DAC_0.OUT.t19 GND 0.07449f
C4067 1Bit_DAC_0.OUT.n31 GND 0.205386f
C4068 1Bit_DAC_0.OUT.n32 GND 0.73234f
C4069 1Bit_DAC_0.OUT.t20 GND 0.07449f
C4070 1Bit_DAC_0.OUT.t27 GND 0.07449f
C4071 1Bit_DAC_0.OUT.n33 GND 0.205386f
C4072 1Bit_DAC_0.OUT.n34 GND 0.755174f
C4073 1Bit_DAC_0.OUT.t22 GND 0.07449f
C4074 1Bit_DAC_0.OUT.t16 GND 0.07449f
C4075 1Bit_DAC_0.OUT.n35 GND 0.2056f
C4076 1Bit_DAC_0.OUT.n36 GND 0.652299f
C4077 1Bit_DAC_0.OUT.t42 GND 0.347549f
C4078 1Bit_DAC_0.OUT.n37 GND 0.508644f
C4079 1Bit_DAC_0.OUT.t18 GND 0.07449f
C4080 1Bit_DAC_0.OUT.t10 GND 0.07449f
C4081 1Bit_DAC_0.OUT.n38 GND 0.205818f
C4082 1Bit_DAC_0.OUT.n39 GND 0.584996f
C4083 1Bit_DAC_0.OUT.t34 GND 0.07449f
C4084 1Bit_DAC_0.OUT.t35 GND 0.07449f
C4085 1Bit_DAC_0.OUT.n40 GND 0.267961f
C4086 1Bit_DAC_0.OUT.n41 GND 0.457761f
C4087 1Bit_DAC_0.OUT.t21 GND 0.07449f
C4088 1Bit_DAC_0.OUT.t15 GND 0.07449f
C4089 1Bit_DAC_0.OUT.n42 GND 0.205818f
C4090 1Bit_DAC_0.OUT.n43 GND 0.566937f
C4091 1Bit_DAC_0.OUT.t47 GND 0.07449f
C4092 1Bit_DAC_0.OUT.t54 GND 0.07449f
C4093 1Bit_DAC_0.OUT.n44 GND 0.267728f
C4094 1Bit_DAC_0.OUT.n45 GND 0.421427f
C4095 1Bit_DAC_0.OUT.t1 GND 0.07449f
C4096 1Bit_DAC_0.OUT.t24 GND 0.07449f
C4097 1Bit_DAC_0.OUT.n46 GND 0.205591f
C4098 1Bit_DAC_0.OUT.n47 GND 0.579805f
C4099 1Bit_DAC_0.OUT.t55 GND 0.07449f
C4100 1Bit_DAC_0.OUT.t46 GND 0.07449f
C4101 1Bit_DAC_0.OUT.n48 GND 0.267961f
C4102 1Bit_DAC_0.OUT.n49 GND 0.457761f
C4103 1Bit_DAC_0.OUT.t9 GND 0.07449f
C4104 1Bit_DAC_0.OUT.t14 GND 0.07449f
C4105 1Bit_DAC_0.OUT.n50 GND 0.205386f
C4106 1Bit_DAC_0.OUT.n51 GND 0.574592f
C4107 1Bit_DAC_0.OUT.t29 GND 0.07449f
C4108 1Bit_DAC_0.OUT.t49 GND 0.07449f
C4109 1Bit_DAC_0.OUT.n52 GND 0.267961f
C4110 1Bit_DAC_0.OUT.n53 GND 0.457761f
C4111 1Bit_DAC_0.OUT.t11 GND 0.306424f
C4112 1Bit_DAC_0.OUT.n54 GND 0.613505f
C4113 a_155026_n27776.t9 GND 0.194162f
C4114 a_155026_n27776.t3 GND 0.10698f
C4115 a_155026_n27776.n0 GND 1.28057f
C4116 a_155026_n27776.n1 GND 0.194927f
C4117 a_155026_n27776.t8 GND 0.009165f
C4118 a_155026_n27776.t7 GND 0.009165f
C4119 a_155026_n27776.n2 GND 0.032429f
C4120 a_155026_n27776.t5 GND 0.009165f
C4121 a_155026_n27776.t4 GND 0.009165f
C4122 a_155026_n27776.n3 GND 0.032429f
C4123 a_155026_n27776.n4 GND 0.095668f
C4124 a_155026_n27776.t6 GND 0.009165f
C4125 a_155026_n27776.t1 GND 0.009165f
C4126 a_155026_n27776.n5 GND 0.038664f
C4127 a_155026_n27776.n6 GND 0.110693f
C4128 a_155026_n27776.n7 GND 0.095728f
C4129 a_155026_n27776.n8 GND 0.200489f
C4130 a_155026_n27776.t2 GND 0.235357f
C4131 a_155026_n27776.n9 GND 1.51988f
C4132 a_155026_n27776.t0 GND 0.107029f
C4133 a_216435_n47946.t2 GND 0.105281f
C4134 a_216435_n47946.t0 GND 0.105281f
C4135 a_216435_n47946.t1 GND 0.105281f
C4136 a_216435_n47946.n0 GND 0.353246f
C4137 a_216435_n47946.t14 GND 0.155234f
C4138 a_216435_n47946.n1 GND 0.5096f
C4139 a_216435_n47946.t13 GND 0.155235f
C4140 a_216435_n47946.t16 GND 0.155235f
C4141 a_216435_n47946.t17 GND 0.155235f
C4142 a_216435_n47946.t26 GND 0.155235f
C4143 a_216435_n47946.t10 GND 0.155235f
C4144 a_216435_n47946.t21 GND 0.155235f
C4145 a_216435_n47946.t23 GND 0.155235f
C4146 a_216435_n47946.t8 GND 0.155235f
C4147 a_216435_n47946.t9 GND 0.155235f
C4148 a_216435_n47946.t20 GND 0.155235f
C4149 a_216435_n47946.t24 GND 0.155234f
C4150 a_216435_n47946.n2 GND 0.201765f
C4151 a_216435_n47946.t25 GND 0.155234f
C4152 a_216435_n47946.n3 GND 0.201765f
C4153 a_216435_n47946.t29 GND 0.155234f
C4154 a_216435_n47946.n4 GND 0.201765f
C4155 a_216435_n47946.t12 GND 0.155234f
C4156 a_216435_n47946.n5 GND 0.201765f
C4157 a_216435_n47946.t22 GND 0.155234f
C4158 a_216435_n47946.n6 GND 0.201765f
C4159 a_216435_n47946.t6 GND 0.155234f
C4160 a_216435_n47946.n7 GND 0.201765f
C4161 a_216435_n47946.t7 GND 0.155234f
C4162 a_216435_n47946.n8 GND 0.201765f
C4163 a_216435_n47946.t11 GND 0.155234f
C4164 a_216435_n47946.n9 GND 0.758672f
C4165 a_216435_n47946.n10 GND 0.71824f
C4166 a_216435_n47946.n11 GND 0.212126f
C4167 a_216435_n47946.n12 GND 0.212126f
C4168 a_216435_n47946.n13 GND 0.212126f
C4169 a_216435_n47946.n14 GND 0.212126f
C4170 a_216435_n47946.n15 GND 0.212126f
C4171 a_216435_n47946.n16 GND 0.212126f
C4172 a_216435_n47946.n17 GND 0.212126f
C4173 a_216435_n47946.n18 GND 0.212126f
C4174 a_216435_n47946.n19 GND 0.364999f
C4175 a_216435_n47946.n20 GND 0.775383f
C4176 a_216435_n47946.t30 GND 0.154452f
C4177 a_216435_n47946.t31 GND 0.15441f
C4178 a_216435_n47946.n21 GND 0.235971f
C4179 a_216435_n47946.t15 GND 0.15441f
C4180 a_216435_n47946.n22 GND 0.142572f
C4181 a_216435_n47946.t19 GND 0.15441f
C4182 a_216435_n47946.n23 GND 0.26826f
C4183 a_216435_n47946.t28 GND 0.154456f
C4184 a_216435_n47946.t32 GND 0.15441f
C4185 a_216435_n47946.n24 GND 0.259537f
C4186 a_216435_n47946.t33 GND 0.15441f
C4187 a_216435_n47946.n25 GND 0.149974f
C4188 a_216435_n47946.t18 GND 0.15441f
C4189 a_216435_n47946.n26 GND 0.149974f
C4190 a_216435_n47946.t27 GND 0.15441f
C4191 a_216435_n47946.n27 GND 0.240839f
C4192 a_216435_n47946.n28 GND 1.99327f
C4193 a_216435_n47946.n29 GND 1.55098f
C4194 a_216435_n47946.t4 GND 0.105281f
C4195 a_216435_n47946.t3 GND 0.105281f
C4196 a_216435_n47946.n30 GND 0.317077f
C4197 a_216435_n47946.n31 GND 1.04451f
C4198 a_216435_n47946.n32 GND 1.11071f
C4199 a_216435_n47946.n33 GND 0.275896f
C4200 a_216435_n47946.t5 GND 0.105281f
C4201 OUT.t11 GND 0.001508f
C4202 OUT.t9 GND 0.001508f
C4203 OUT.n0 GND 0.003259f
C4204 OUT.t8 GND 0.001508f
C4205 OUT.t10 GND 0.001508f
C4206 OUT.n1 GND 0.00496f
C4207 OUT.n2 GND 0.013781f
C4208 OUT.t2 GND 0.001508f
C4209 OUT.t3 GND 0.001508f
C4210 OUT.n3 GND 0.00458f
C4211 OUT.t0 GND 0.001508f
C4212 OUT.t1 GND 0.001508f
C4213 OUT.n4 GND 0.003353f
C4214 OUT.n5 GND 0.014922f
C4215 OUT.n6 GND 0.001002f
C4216 OUT.t5 GND 9.8e-19
C4217 OUT.t7 GND 9.8e-19
C4218 OUT.n7 GND 0.002445f
C4219 OUT.t4 GND 9.8e-19
C4220 OUT.t6 GND 9.8e-19
C4221 OUT.n8 GND 0.001961f
C4222 OUT.n9 GND 0.004521f
C4223 OUT.n10 GND 0.009217f
C4224 OUT.t73 GND 0.001383f
C4225 OUT.t20 GND 0.002346f
C4226 OUT.t37 GND 0.001383f
C4227 OUT.t60 GND 0.002346f
C4228 OUT.n11 GND 0.003162f
C4229 OUT.n12 GND 0.001285f
C4230 OUT.n13 GND 0.001548f
C4231 OUT.n14 GND 0.003384f
C4232 OUT.t57 GND 0.001383f
C4233 OUT.t83 GND 0.002346f
C4234 OUT.t18 GND 0.001383f
C4235 OUT.t46 GND 0.002346f
C4236 OUT.n15 GND 0.003937f
C4237 OUT.n16 GND 0.004158f
C4238 OUT.n17 GND 0.001568f
C4239 OUT.n18 GND 0.00266f
C4240 OUT.n19 GND 0.033342f
C4241 OUT.n20 GND 0.002179f
C4242 OUT.n21 GND 0.024579f
C4243 OUT.n22 GND 0.234645f
C4244 OUT.n23 GND 0.307797f
C4245 OUT.t40 GND 0.01359f
C4246 OUT.t80 GND 0.01359f
C4247 OUT.t78 GND 0.01359f
C4248 OUT.t49 GND 0.01359f
C4249 OUT.t42 GND 0.01359f
C4250 OUT.t81 GND 0.01359f
C4251 OUT.t54 GND 0.01359f
C4252 OUT.t22 GND 0.01359f
C4253 OUT.t21 GND 0.01359f
C4254 OUT.t15 GND 0.01359f
C4255 OUT.t38 GND 0.01359f
C4256 OUT.t29 GND 0.01359f
C4257 OUT.t25 GND 0.01357f
C4258 OUT.t59 GND 0.013522f
C4259 OUT.t62 GND 0.013518f
C4260 OUT.n24 GND 0.020659f
C4261 OUT.t19 GND 0.013518f
C4262 OUT.n25 GND 0.012482f
C4263 OUT.t26 GND 0.013518f
C4264 OUT.n26 GND 0.023486f
C4265 OUT.t56 GND 0.013522f
C4266 OUT.t64 GND 0.013518f
C4267 OUT.n27 GND 0.022722f
C4268 OUT.t66 GND 0.013518f
C4269 OUT.n28 GND 0.01313f
C4270 OUT.t23 GND 0.013518f
C4271 OUT.n29 GND 0.01313f
C4272 OUT.t55 GND 0.013518f
C4273 OUT.n30 GND 0.021085f
C4274 OUT.n31 GND 0.187142f
C4275 OUT.n32 GND 0.15263f
C4276 OUT.t31 GND 0.013658f
C4277 OUT.n33 GND 0.053999f
C4278 OUT.n34 GND 0.030235f
C4279 OUT.n35 GND 0.025429f
C4280 OUT.n36 GND 0.035776f
C4281 OUT.n37 GND 0.035776f
C4282 OUT.n38 GND 0.018571f
C4283 OUT.n39 GND 0.018571f
C4284 OUT.n40 GND 0.018571f
C4285 OUT.n41 GND 0.018571f
C4286 OUT.n42 GND 0.018571f
C4287 OUT.n43 GND 0.018571f
C4288 OUT.n44 GND 0.018571f
C4289 OUT.n45 GND 0.018571f
C4290 OUT.n46 GND 0.06288f
C4291 OUT.t85 GND 0.01359f
C4292 OUT.n47 GND 0.06642f
C4293 OUT.t76 GND 0.01359f
C4294 OUT.n48 GND 0.017664f
C4295 OUT.t75 GND 0.01359f
C4296 OUT.n49 GND 0.017664f
C4297 OUT.t45 GND 0.01359f
C4298 OUT.n50 GND 0.017664f
C4299 OUT.t86 GND 0.01359f
C4300 OUT.n51 GND 0.017664f
C4301 OUT.t58 GND 0.01359f
C4302 OUT.n52 GND 0.017664f
C4303 OUT.t53 GND 0.01359f
C4304 OUT.n53 GND 0.017664f
C4305 OUT.t52 GND 0.01359f
C4306 OUT.n54 GND 0.017664f
C4307 OUT.t17 GND 0.01359f
C4308 OUT.n55 GND 0.034869f
C4309 OUT.t67 GND 0.01359f
C4310 OUT.n56 GND 0.034869f
C4311 OUT.t34 GND 0.01359f
C4312 OUT.n57 GND 0.029514f
C4313 OUT.n58 GND 12.909201f
C4314 OUT.t50 GND 0.013595f
C4315 OUT.t14 GND 0.01359f
C4316 OUT.n59 GND 0.051293f
C4317 OUT.t35 GND 0.013596f
C4318 OUT.t36 GND 0.01359f
C4319 OUT.n60 GND 0.040071f
C4320 OUT.t69 GND 0.01359f
C4321 OUT.n61 GND 0.017664f
C4322 OUT.t74 GND 0.01359f
C4323 OUT.n62 GND 0.017664f
C4324 OUT.t33 GND 0.01359f
C4325 OUT.n63 GND 0.017664f
C4326 OUT.t65 GND 0.01359f
C4327 OUT.n64 GND 0.017664f
C4328 OUT.t68 GND 0.01359f
C4329 OUT.n65 GND 0.017664f
C4330 OUT.t24 GND 0.01359f
C4331 OUT.n66 GND 0.017664f
C4332 OUT.t32 GND 0.01359f
C4333 OUT.n67 GND 0.033299f
C4334 OUT.t61 GND 0.01359f
C4335 OUT.t27 GND 0.01359f
C4336 OUT.t71 GND 0.01359f
C4337 OUT.t70 GND 0.01359f
C4338 OUT.t63 GND 0.01359f
C4339 OUT.t28 GND 0.01359f
C4340 OUT.t72 GND 0.01359f
C4341 OUT.t41 GND 0.01359f
C4342 OUT.t39 GND 0.01359f
C4343 OUT.t30 GND 0.013594f
C4344 OUT.n68 GND 0.034848f
C4345 OUT.n69 GND 0.018571f
C4346 OUT.n70 GND 0.018571f
C4347 OUT.n71 GND 0.018571f
C4348 OUT.n72 GND 0.018571f
C4349 OUT.n73 GND 0.018571f
C4350 OUT.n74 GND 0.018571f
C4351 OUT.n75 GND 0.018571f
C4352 OUT.n76 GND 0.028244f
C4353 OUT.n77 GND 0.218282f
C4354 OUT.n78 GND 0.194929f
C4355 OUT.n79 GND 0.059213f
C4356 OUT.n80 GND 0.012289f
C4357 OUT.n81 GND 0.082396f
C4358 OUT.t87 GND 0.01359f
C4359 OUT.t16 GND 0.013595f
C4360 OUT.n82 GND 0.045727f
C4361 OUT.n83 GND 0.005376f
C4362 OUT.n84 GND 0.042175f
C4363 OUT.t79 GND 0.013523f
C4364 OUT.t13 GND 0.013518f
C4365 OUT.n85 GND 0.023379f
C4366 OUT.t47 GND 0.013518f
C4367 OUT.n86 GND 0.01313f
C4368 OUT.t48 GND 0.013518f
C4369 OUT.n87 GND 0.01313f
C4370 OUT.t77 GND 0.013518f
C4371 OUT.n88 GND 0.054085f
C4372 OUT.t51 GND 0.013518f
C4373 OUT.n89 GND 0.06399f
C4374 OUT.t44 GND 0.013518f
C4375 OUT.n90 GND 0.017326f
C4376 OUT.t43 GND 0.013518f
C4377 OUT.n91 GND 0.017326f
C4378 OUT.t84 GND 0.013518f
C4379 OUT.n92 GND 0.065032f
C4380 OUT.t12 GND 0.013518f
C4381 OUT.n93 GND 0.079231f
C4382 OUT.n94 GND 0.007084f
C4383 OUT.t82 GND 0.013606f
C4384 OUT.n95 GND 0.086585f
C4385 OUT.n96 GND 0.007821f
C4386 OUT.n97 GND 3.77453f
C4387 OUT.n98 GND 20.748f
C4388 1Bit_Clk_ADC_0.x3.B.n0 GND 0.013359f
C4389 1Bit_Clk_ADC_0.x3.B.t6 GND 0.00748f
C4390 1Bit_Clk_ADC_0.x3.B.t7 GND 0.00748f
C4391 1Bit_Clk_ADC_0.x3.B.n1 GND 0.018657f
C4392 1Bit_Clk_ADC_0.x3.B.t4 GND 0.00748f
C4393 1Bit_Clk_ADC_0.x3.B.t5 GND 0.00748f
C4394 1Bit_Clk_ADC_0.x3.B.n2 GND 0.014961f
C4395 1Bit_Clk_ADC_0.x3.B.n3 GND 0.036229f
C4396 1Bit_Clk_ADC_0.x3.B.t21 GND 0.017902f
C4397 1Bit_Clk_ADC_0.x3.B.t16 GND 0.010549f
C4398 1Bit_Clk_ADC_0.x3.B.n4 GND 0.037964f
C4399 1Bit_Clk_ADC_0.x3.B.t35 GND 0.017902f
C4400 1Bit_Clk_ADC_0.x3.B.t26 GND 0.010549f
C4401 1Bit_Clk_ADC_0.x3.B.t28 GND 0.017902f
C4402 1Bit_Clk_ADC_0.x3.B.t22 GND 0.010549f
C4403 1Bit_Clk_ADC_0.x3.B.n5 GND 0.025817f
C4404 1Bit_Clk_ADC_0.x3.B.t14 GND 0.017902f
C4405 1Bit_Clk_ADC_0.x3.B.t32 GND 0.010549f
C4406 1Bit_Clk_ADC_0.x3.B.n6 GND 0.024129f
C4407 1Bit_Clk_ADC_0.x3.B.n7 GND 0.011815f
C4408 1Bit_Clk_ADC_0.x3.B.n8 GND 0.009803f
C4409 1Bit_Clk_ADC_0.x3.B.n9 GND 0.009803f
C4410 1Bit_Clk_ADC_0.x3.B.n10 GND 0.011815f
C4411 1Bit_Clk_ADC_0.x3.B.n11 GND 0.025817f
C4412 1Bit_Clk_ADC_0.x3.B.n12 GND 0.011815f
C4413 1Bit_Clk_ADC_0.x3.B.n13 GND 0.00341f
C4414 1Bit_Clk_ADC_0.x3.B.n14 GND 0.085699f
C4415 1Bit_Clk_ADC_0.x3.B.t27 GND 0.010549f
C4416 1Bit_Clk_ADC_0.x3.B.t12 GND 0.017902f
C4417 1Bit_Clk_ADC_0.x3.B.t34 GND 0.010549f
C4418 1Bit_Clk_ADC_0.x3.B.t18 GND 0.017902f
C4419 1Bit_Clk_ADC_0.x3.B.n15 GND 0.025817f
C4420 1Bit_Clk_ADC_0.x3.B.t33 GND 0.010549f
C4421 1Bit_Clk_ADC_0.x3.B.t17 GND 0.017902f
C4422 1Bit_Clk_ADC_0.x3.B.t13 GND 0.010549f
C4423 1Bit_Clk_ADC_0.x3.B.t20 GND 0.017902f
C4424 1Bit_Clk_ADC_0.x3.B.n16 GND 0.024129f
C4425 1Bit_Clk_ADC_0.x3.B.n17 GND 0.011935f
C4426 1Bit_Clk_ADC_0.x3.B.n18 GND 0.025817f
C4427 1Bit_Clk_ADC_0.x3.B.n19 GND 0.011815f
C4428 1Bit_Clk_ADC_0.x3.B.n20 GND 0.009803f
C4429 1Bit_Clk_ADC_0.x3.B.n21 GND 0.009803f
C4430 1Bit_Clk_ADC_0.x3.B.n22 GND 0.011815f
C4431 1Bit_Clk_ADC_0.x3.B.n23 GND 0.040098f
C4432 1Bit_Clk_ADC_0.x3.B.t29 GND 0.010549f
C4433 1Bit_Clk_ADC_0.x3.B.t15 GND 0.017902f
C4434 1Bit_Clk_ADC_0.x3.B.t19 GND 0.010549f
C4435 1Bit_Clk_ADC_0.x3.B.t25 GND 0.017902f
C4436 1Bit_Clk_ADC_0.x3.B.n24 GND 0.025817f
C4437 1Bit_Clk_ADC_0.x3.B.t24 GND 0.010549f
C4438 1Bit_Clk_ADC_0.x3.B.t31 GND 0.017902f
C4439 1Bit_Clk_ADC_0.x3.B.n25 GND 0.024129f
C4440 1Bit_Clk_ADC_0.x3.B.n26 GND 0.011815f
C4441 1Bit_Clk_ADC_0.x3.B.n27 GND 0.009164f
C4442 1Bit_Clk_ADC_0.x3.B.n28 GND 0.00959f
C4443 1Bit_Clk_ADC_0.x3.B.n29 GND 0.011815f
C4444 1Bit_Clk_ADC_0.x3.B.n30 GND 0.025817f
C4445 1Bit_Clk_ADC_0.x3.B.t23 GND 0.010549f
C4446 1Bit_Clk_ADC_0.x3.B.t30 GND 0.017902f
C4447 1Bit_Clk_ADC_0.x3.B.n31 GND 0.012134f
C4448 1Bit_Clk_ADC_0.x3.B.n32 GND 0.037834f
C4449 1Bit_Clk_ADC_0.x3.B.n33 GND 0.011815f
C4450 1Bit_Clk_ADC_0.x3.B.n34 GND 0.002451f
C4451 1Bit_Clk_ADC_0.x3.B.n35 GND 0.019516f
C4452 1Bit_Clk_ADC_0.x3.B.n36 GND 0.212334f
C4453 1Bit_Clk_ADC_0.x3.B.n37 GND 0.201584f
C4454 1Bit_Clk_ADC_0.x3.B.n38 GND 0.020768f
C4455 1Bit_Clk_ADC_0.x3.B.t8 GND 0.011508f
C4456 1Bit_Clk_ADC_0.x3.B.t9 GND 0.011508f
C4457 1Bit_Clk_ADC_0.x3.B.n39 GND 0.024865f
C4458 1Bit_Clk_ADC_0.x3.B.t10 GND 0.011508f
C4459 1Bit_Clk_ADC_0.x3.B.t11 GND 0.011508f
C4460 1Bit_Clk_ADC_0.x3.B.n40 GND 0.037845f
C4461 1Bit_Clk_ADC_0.x3.B.n41 GND 0.105155f
C4462 1Bit_Clk_ADC_0.x3.B.n42 GND 0.020869f
C4463 1Bit_Clk_ADC_0.x3.B.t2 GND 0.011508f
C4464 1Bit_Clk_ADC_0.x3.B.t0 GND 0.011508f
C4465 1Bit_Clk_ADC_0.x3.B.n43 GND 0.025583f
C4466 1Bit_Clk_ADC_0.x3.B.t1 GND 0.011508f
C4467 1Bit_Clk_ADC_0.x3.B.t3 GND 0.011508f
C4468 1Bit_Clk_ADC_0.x3.B.n44 GND 0.034943f
C4469 1Bit_Clk_ADC_0.x3.B.n45 GND 0.113861f
C4470 1Bit_Clk_ADC_0.x14.Y.t1 GND 0.02612f
C4471 1Bit_Clk_ADC_0.x14.Y.n0 GND 0.008403f
C4472 1Bit_Clk_ADC_0.x14.Y.t12 GND 0.015406f
C4473 1Bit_Clk_ADC_0.x14.Y.t16 GND 0.026143f
C4474 1Bit_Clk_ADC_0.x14.Y.t5 GND 0.015406f
C4475 1Bit_Clk_ADC_0.x14.Y.t10 GND 0.026143f
C4476 1Bit_Clk_ADC_0.x14.Y.n1 GND 0.035237f
C4477 1Bit_Clk_ADC_0.x14.Y.n2 GND 0.017254f
C4478 1Bit_Clk_ADC_0.x14.Y.n3 GND 0.037702f
C4479 1Bit_Clk_ADC_0.x14.Y.t7 GND 0.015406f
C4480 1Bit_Clk_ADC_0.x14.Y.t14 GND 0.026143f
C4481 1Bit_Clk_ADC_0.x14.Y.t3 GND 0.015406f
C4482 1Bit_Clk_ADC_0.x14.Y.t9 GND 0.026143f
C4483 1Bit_Clk_ADC_0.x14.Y.n4 GND 0.043864f
C4484 1Bit_Clk_ADC_0.x14.Y.n5 GND 0.046329f
C4485 1Bit_Clk_ADC_0.x14.Y.n6 GND 0.017855f
C4486 1Bit_Clk_ADC_0.x14.Y.n7 GND 0.039956f
C4487 1Bit_Clk_ADC_0.x14.Y.t6 GND 0.026143f
C4488 1Bit_Clk_ADC_0.x14.Y.t18 GND 0.015406f
C4489 1Bit_Clk_ADC_0.x14.Y.t17 GND 0.026143f
C4490 1Bit_Clk_ADC_0.x14.Y.t13 GND 0.015406f
C4491 1Bit_Clk_ADC_0.x14.Y.n8 GND 0.037702f
C4492 1Bit_Clk_ADC_0.x14.Y.t8 GND 0.026143f
C4493 1Bit_Clk_ADC_0.x14.Y.t4 GND 0.015406f
C4494 1Bit_Clk_ADC_0.x14.Y.n9 GND 0.035237f
C4495 1Bit_Clk_ADC_0.x14.Y.n10 GND 0.017254f
C4496 1Bit_Clk_ADC_0.x14.Y.n11 GND 0.017254f
C4497 1Bit_Clk_ADC_0.x14.Y.n12 GND 0.037702f
C4498 1Bit_Clk_ADC_0.x14.Y.t15 GND 0.026143f
C4499 1Bit_Clk_ADC_0.x14.Y.t11 GND 0.015406f
C4500 1Bit_Clk_ADC_0.x14.Y.n13 GND 0.01772f
C4501 1Bit_Clk_ADC_0.x14.Y.n14 GND 0.05525f
C4502 1Bit_Clk_ADC_0.x14.Y.n15 GND 0.017254f
C4503 1Bit_Clk_ADC_0.x14.Y.n16 GND 0.012293f
C4504 1Bit_Clk_ADC_0.x14.Y.n17 GND 0.083147f
C4505 1Bit_Clk_ADC_0.x14.Y.n18 GND 1.373f
C4506 1Bit_Clk_ADC_0.x14.Y.n19 GND 0.092533f
C4507 1Bit_Clk_ADC_0.x14.Y.t0 GND 0.014117f
C4508 1Bit_Clk_ADC_0.x14.Y.t2 GND 0.014117f
C4509 1Bit_Clk_ADC_0.x14.Y.n20 GND 0.030892f
C4510 a_219526_n14006.n0 GND 0.005132f
C4511 a_219526_n14006.n1 GND 0.041278f
C4512 a_219526_n14006.n2 GND 0.043242f
C4513 a_219526_n14006.n3 GND 0.03304f
C4514 a_219526_n14006.n4 GND 0.03304f
C4515 a_219526_n14006.n5 GND 0.043242f
C4516 a_219526_n14006.n6 GND 0.065687f
C4517 a_219526_n14006.n7 GND 0.01031f
C4518 a_219526_n14006.n8 GND 0.065687f
C4519 a_219526_n14006.n9 GND 0.01031f
C4520 a_219526_n14006.n10 GND 0.065687f
C4521 a_219526_n14006.n11 GND 0.01031f
C4522 a_219526_n14006.n12 GND 0.07304f
C4523 a_219526_n14006.n13 GND 0.030644f
C4524 a_219526_n14006.n14 GND 2.85905f
C4525 a_219526_n14006.n15 GND 2.89225f
C4526 a_219526_n14006.n16 GND 0.06592f
C4527 a_219526_n14006.n17 GND 0.010339f
C4528 a_219526_n14006.n18 GND 0.041899f
C4529 a_219526_n14006.n19 GND 0.06592f
C4530 a_219526_n14006.n20 GND 0.010339f
C4531 a_219526_n14006.n21 GND 0.06592f
C4532 a_219526_n14006.n22 GND 0.010339f
C4533 a_219526_n14006.n23 GND 0.06592f
C4534 a_219526_n14006.n24 GND 0.010339f
C4535 a_219526_n14006.n25 GND 0.06592f
C4536 a_219526_n14006.n26 GND 0.010339f
C4537 a_219526_n14006.n27 GND 0.06592f
C4538 a_219526_n14006.n28 GND 0.010339f
C4539 a_219526_n14006.n29 GND 0.070626f
C4540 a_219526_n14006.n30 GND 0.026553f
C4541 a_219526_n14006.n31 GND 0.01892f
C4542 a_219526_n14006.n32 GND 0.043297f
C4543 a_219526_n14006.n33 GND 0.005132f
C4544 a_219526_n14006.n34 GND 0.03124f
C4545 a_219526_n14006.n35 GND 0.03124f
C4546 a_219526_n14006.n36 GND 0.005132f
C4547 a_219526_n14006.n37 GND 0.043297f
C4548 a_219526_n14006.t2 GND 0.355305f
C4549 a_219526_n14006.n38 GND 0.492082f
C4550 a_219526_n14006.t7 GND 0.064372f
C4551 a_219526_n14006.n39 GND 0.005434f
C4552 a_219526_n14006.n40 GND 0.005434f
C4553 a_219526_n14006.n41 GND 0.005434f
C4554 a_219526_n14006.n42 GND 5.99e-19
C4555 a_219526_n14006.n43 GND 0.005434f
C4556 a_219526_n14006.n44 GND 0.005434f
C4557 a_219526_n14006.n45 GND 0.009037f
C4558 a_219526_n14006.n46 GND 0.005434f
C4559 a_219526_n14006.n47 GND 0.005434f
C4560 a_219526_n14006.n48 GND 0.005434f
C4561 a_219526_n14006.n49 GND 0.005434f
C4562 a_219526_n14006.n50 GND 0.005434f
C4563 a_219526_n14006.n51 GND 0.125843f
C4564 a_219526_n14006.n52 GND 0.137608f
C4565 a_219526_n14006.t12 GND 0.355184f
C4566 a_219526_n14006.n53 GND 0.137608f
C4567 a_219526_n14006.t40 GND 0.355184f
C4568 a_219526_n14006.n54 GND 0.125843f
C4569 a_219526_n14006.n55 GND 0.005132f
C4570 a_219526_n14006.n56 GND 0.01892f
C4571 a_219526_n14006.n57 GND 0.005132f
C4572 a_219526_n14006.n58 GND 0.016538f
C4573 a_219526_n14006.n59 GND 0.263581f
C4574 a_219526_n14006.t19 GND 0.064372f
C4575 a_219526_n14006.n60 GND 0.005434f
C4576 a_219526_n14006.n61 GND 0.006774f
C4577 a_219526_n14006.n62 GND 0.014408f
C4578 a_219526_n14006.n63 GND 0.013908f
C4579 a_219526_n14006.n64 GND 0.011863f
C4580 a_219526_n14006.n65 GND 0.011644f
C4581 a_219526_n14006.t13 GND 0.064372f
C4582 a_219526_n14006.n66 GND 0.132696f
C4583 a_219526_n14006.n67 GND 0.451349f
C4584 a_219526_n14006.n68 GND 0.235578f
C4585 a_219526_n14006.t43 GND 0.064372f
C4586 a_219526_n14006.n69 GND 0.005434f
C4587 a_219526_n14006.n70 GND 0.005434f
C4588 a_219526_n14006.n71 GND 0.006731f
C4589 a_219526_n14006.n72 GND 0.014481f
C4590 a_219526_n14006.n73 GND 0.005132f
C4591 a_219526_n14006.n74 GND 0.014703f
C4592 a_219526_n14006.n75 GND 0.013534f
C4593 a_219526_n14006.n76 GND 0.011983f
C4594 a_219526_n14006.n77 GND 0.00956f
C4595 a_219526_n14006.t48 GND 0.064372f
C4596 a_219526_n14006.n78 GND 0.138f
C4597 a_219526_n14006.n79 GND 0.030321f
C4598 a_219526_n14006.n80 GND 0.005132f
C4599 a_219526_n14006.t25 GND 0.064372f
C4600 a_219526_n14006.n81 GND 0.005434f
C4601 a_219526_n14006.n82 GND 0.005434f
C4602 a_219526_n14006.n83 GND 0.005132f
C4603 a_219526_n14006.n84 GND 0.01892f
C4604 a_219526_n14006.n85 GND 0.016538f
C4605 a_219526_n14006.n86 GND 0.005132f
C4606 a_219526_n14006.n87 GND 0.005434f
C4607 a_219526_n14006.n88 GND 0.005434f
C4608 a_219526_n14006.n89 GND 0.005434f
C4609 a_219526_n14006.n90 GND 5.99e-19
C4610 a_219526_n14006.n91 GND 0.005434f
C4611 a_219526_n14006.n92 GND 0.005434f
C4612 a_219526_n14006.n93 GND 0.005434f
C4613 a_219526_n14006.n94 GND 0.005434f
C4614 a_219526_n14006.n95 GND 0.005434f
C4615 a_219526_n14006.t15 GND 0.064372f
C4616 a_219526_n14006.n96 GND 0.131393f
C4617 a_219526_n14006.t65 GND 0.355184f
C4618 a_219526_n14006.n97 GND 0.137608f
C4619 a_219526_n14006.n98 GND 0.137608f
C4620 a_219526_n14006.n99 GND 0.137608f
C4621 a_219526_n14006.n100 GND 0.38333f
C4622 a_219526_n14006.n101 GND 0.137608f
C4623 a_219526_n14006.n102 GND 0.137608f
C4624 a_219526_n14006.n103 GND 0.137608f
C4625 a_219526_n14006.n104 GND 0.131171f
C4626 a_219526_n14006.t59 GND 0.355184f
C4627 a_219526_n14006.n105 GND 0.086162f
C4628 a_219526_n14006.t20 GND 0.355362f
C4629 a_219526_n14006.n106 GND 0.027258f
C4630 a_219526_n14006.n107 GND 0.125621f
C4631 a_219526_n14006.t17 GND 0.064372f
C4632 a_219526_n14006.n108 GND 0.005434f
C4633 a_219526_n14006.n109 GND 0.005434f
C4634 a_219526_n14006.n110 GND 0.005434f
C4635 a_219526_n14006.n111 GND 0.005434f
C4636 a_219526_n14006.n112 GND 0.005434f
C4637 a_219526_n14006.n113 GND 5.99e-19
C4638 a_219526_n14006.n114 GND 0.005434f
C4639 a_219526_n14006.n115 GND 0.005434f
C4640 a_219526_n14006.n116 GND 0.005434f
C4641 a_219526_n14006.n117 GND 0.005434f
C4642 a_219526_n14006.n118 GND 0.005434f
C4643 a_219526_n14006.t37 GND 0.064372f
C4644 a_219526_n14006.n119 GND 0.023104f
C4645 a_219526_n14006.n120 GND 0.005132f
C4646 a_219526_n14006.n121 GND 0.01892f
C4647 a_219526_n14006.n122 GND 0.005132f
C4648 a_219526_n14006.n123 GND 0.016538f
C4649 a_219526_n14006.n124 GND 0.235578f
C4650 a_219526_n14006.n125 GND 0.235578f
C4651 a_219526_n14006.t42 GND 0.064372f
C4652 a_219526_n14006.n126 GND 0.005434f
C4653 a_219526_n14006.n127 GND 0.005434f
C4654 a_219526_n14006.n128 GND 0.006731f
C4655 a_219526_n14006.n129 GND 0.014481f
C4656 a_219526_n14006.n130 GND 0.005132f
C4657 a_219526_n14006.n131 GND 0.014703f
C4658 a_219526_n14006.n132 GND 0.013534f
C4659 a_219526_n14006.n133 GND 0.011983f
C4660 a_219526_n14006.n134 GND 0.00956f
C4661 a_219526_n14006.t44 GND 0.064372f
C4662 a_219526_n14006.n135 GND 0.138f
C4663 a_219526_n14006.t46 GND 0.064372f
C4664 a_219526_n14006.n136 GND 0.005434f
C4665 a_219526_n14006.n137 GND 0.005434f
C4666 a_219526_n14006.n138 GND 0.006731f
C4667 a_219526_n14006.n139 GND 0.014481f
C4668 a_219526_n14006.n140 GND 0.005132f
C4669 a_219526_n14006.n141 GND 0.014703f
C4670 a_219526_n14006.n142 GND 0.013534f
C4671 a_219526_n14006.n143 GND 0.011983f
C4672 a_219526_n14006.n144 GND 0.00956f
C4673 a_219526_n14006.t45 GND 0.064372f
C4674 a_219526_n14006.n145 GND 0.138f
C4675 a_219526_n14006.n146 GND 0.031711f
C4676 a_219526_n14006.n147 GND 0.005434f
C4677 a_219526_n14006.n148 GND 0.013534f
C4678 a_219526_n14006.n149 GND 0.005132f
C4679 a_219526_n14006.n150 GND 0.017509f
C4680 a_219526_n14006.n151 GND 0.005434f
C4681 a_219526_n14006.n152 GND 0.041602f
C4682 a_219526_n14006.t47 GND 0.025132f
C4683 a_219526_n14006.n153 GND 0.013132f
C4684 a_219526_n14006.n154 GND 0.00637f
C4685 a_219526_n14006.n155 GND 0.005132f
C4686 a_219526_n14006.n156 GND 0.257889f
C4687 a_219526_n14006.n157 GND 0.005132f
C4688 a_219526_n14006.n158 GND 0.005434f
C4689 a_219526_n14006.n159 GND 0.017509f
C4690 a_219526_n14006.n160 GND 0.017509f
C4691 a_219526_n14006.n161 GND 0.005434f
C4692 a_219526_n14006.n162 GND 0.005132f
C4693 a_219526_n14006.n163 GND 0.014703f
C4694 a_219526_n14006.n164 GND 0.014481f
C4695 a_219526_n14006.n165 GND 0.006383f
C4696 a_219526_n14006.n166 GND 1.29341f
C4697 a_219526_n14006.n167 GND 0.038111f
C4698 a_219526_n14006.n168 GND 0.005434f
C4699 a_219526_n14006.n169 GND 0.017509f
C4700 a_219526_n14006.n170 GND 0.005434f
C4701 a_219526_n14006.n171 GND 0.042649f
C4702 a_219526_n14006.t21 GND 0.032791f
C4703 a_219526_n14006.n172 GND 0.013132f
C4704 a_219526_n14006.n173 GND 0.006711f
C4705 a_219526_n14006.n174 GND 0.005132f
C4706 a_219526_n14006.n175 GND 0.249137f
C4707 a_219526_n14006.n176 GND 0.014655f
C4708 a_219526_n14006.n177 GND 0.005132f
C4709 a_219526_n14006.n178 GND 0.005434f
C4710 a_219526_n14006.n179 GND 0.017509f
C4711 a_219526_n14006.n180 GND 0.017509f
C4712 a_219526_n14006.n181 GND 0.005434f
C4713 a_219526_n14006.n182 GND 0.005132f
C4714 a_219526_n14006.n183 GND 0.013908f
C4715 a_219526_n14006.n184 GND 0.014408f
C4716 a_219526_n14006.n185 GND 0.006562f
C4717 a_219526_n14006.n186 GND 0.284426f
C4718 a_219526_n14006.n187 GND 0.263581f
C4719 a_219526_n14006.n188 GND 0.263581f
C4720 a_219526_n14006.n189 GND 0.263581f
C4721 a_219526_n14006.n190 GND 0.263581f
C4722 a_219526_n14006.t1 GND 0.064372f
C4723 a_219526_n14006.n191 GND 0.005434f
C4724 a_219526_n14006.n192 GND 0.006774f
C4725 a_219526_n14006.n193 GND 0.014408f
C4726 a_219526_n14006.n194 GND 0.013908f
C4727 a_219526_n14006.n195 GND 0.011863f
C4728 a_219526_n14006.n196 GND 0.011644f
C4729 a_219526_n14006.t23 GND 0.064372f
C4730 a_219526_n14006.n197 GND 0.132696f
C4731 a_219526_n14006.n198 GND 0.451349f
C4732 a_219526_n14006.t39 GND 0.064372f
C4733 a_219526_n14006.n199 GND 0.005434f
C4734 a_219526_n14006.n200 GND 0.006774f
C4735 a_219526_n14006.n201 GND 0.014408f
C4736 a_219526_n14006.n202 GND 0.013908f
C4737 a_219526_n14006.n203 GND 0.011863f
C4738 a_219526_n14006.n204 GND 0.011644f
C4739 a_219526_n14006.t35 GND 0.064372f
C4740 a_219526_n14006.n205 GND 0.132696f
C4741 a_219526_n14006.n206 GND 0.458008f
C4742 a_219526_n14006.t11 GND 0.064372f
C4743 a_219526_n14006.n207 GND 0.005434f
C4744 a_219526_n14006.n208 GND 0.006774f
C4745 a_219526_n14006.n209 GND 0.014408f
C4746 a_219526_n14006.n210 GND 0.013908f
C4747 a_219526_n14006.n211 GND 0.011863f
C4748 a_219526_n14006.n212 GND 0.011644f
C4749 a_219526_n14006.t5 GND 0.064372f
C4750 a_219526_n14006.n213 GND 0.132696f
C4751 a_219526_n14006.n214 GND 0.451349f
C4752 a_219526_n14006.t33 GND 0.064372f
C4753 a_219526_n14006.n215 GND 0.005434f
C4754 a_219526_n14006.n216 GND 0.006774f
C4755 a_219526_n14006.n217 GND 0.014408f
C4756 a_219526_n14006.n218 GND 0.013908f
C4757 a_219526_n14006.n219 GND 0.011863f
C4758 a_219526_n14006.n220 GND 0.011644f
C4759 a_219526_n14006.t29 GND 0.064372f
C4760 a_219526_n14006.n221 GND 0.132696f
C4761 a_219526_n14006.n222 GND 0.451349f
C4762 a_219526_n14006.n223 GND 0.005434f
C4763 a_219526_n14006.n224 GND 0.005132f
C4764 a_219526_n14006.t31 GND 0.064372f
C4765 a_219526_n14006.n225 GND 0.009037f
C4766 a_219526_n14006.n226 GND 0.005132f
C4767 a_219526_n14006.n227 GND 0.005434f
C4768 a_219526_n14006.n228 GND 0.005132f
C4769 a_219526_n14006.n229 GND 0.005434f
C4770 a_219526_n14006.n230 GND 0.005434f
C4771 a_219526_n14006.n231 GND 5.99e-19
C4772 a_219526_n14006.n232 GND 0.005434f
C4773 a_219526_n14006.n233 GND 0.005434f
C4774 a_219526_n14006.n234 GND 0.005434f
C4775 a_219526_n14006.n235 GND 0.005434f
C4776 a_219526_n14006.n236 GND 0.005434f
C4777 a_219526_n14006.t27 GND 0.064372f
C4778 a_219526_n14006.n237 GND 0.125177f
C4779 a_219526_n14006.t36 GND 0.355184f
C4780 a_219526_n14006.n238 GND 0.128951f
C4781 a_219526_n14006.n239 GND 0.023688f
C4782 a_219526_n14006.n240 GND 0.137608f
C4783 a_219526_n14006.n241 GND 0.137608f
C4784 a_219526_n14006.n242 GND 0.137608f
C4785 a_219526_n14006.n243 GND 0.137608f
C4786 a_219526_n14006.n244 GND 0.137608f
C4787 a_219526_n14006.t18 GND 0.355184f
C4788 a_219526_n14006.n245 GND 0.137608f
C4789 a_219526_n14006.t22 GND 0.355184f
C4790 a_219526_n14006.n246 GND 0.137608f
C4791 a_219526_n14006.n247 GND 0.137608f
C4792 a_219526_n14006.t0 GND 0.355184f
C4793 a_219526_n14006.n248 GND 0.122514f
C4794 a_219526_n14006.t34 GND 0.355184f
C4795 a_219526_n14006.n249 GND 0.38333f
C4796 a_219526_n14006.n250 GND 0.122736f
C4797 a_219526_n14006.t38 GND 0.355184f
C4798 a_219526_n14006.n251 GND 0.137608f
C4799 a_219526_n14006.t4 GND 0.355184f
C4800 a_219526_n14006.n252 GND 0.137608f
C4801 a_219526_n14006.n253 GND 0.137608f
C4802 a_219526_n14006.t10 GND 0.355184f
C4803 a_219526_n14006.n254 GND 0.137608f
C4804 a_219526_n14006.t28 GND 0.355184f
C4805 a_219526_n14006.n255 GND 0.137608f
C4806 a_219526_n14006.n256 GND 0.137608f
C4807 a_219526_n14006.t32 GND 0.355184f
C4808 a_219526_n14006.n257 GND 0.137608f
C4809 a_219526_n14006.t26 GND 0.355184f
C4810 a_219526_n14006.n258 GND 0.125177f
C4811 a_219526_n14006.n259 GND 0.030321f
C4812 a_219526_n14006.n260 GND 0.125843f
C4813 a_219526_n14006.t30 GND 0.355184f
C4814 a_219526_n14006.n261 GND 0.125843f
C4815 a_219526_n14006.n262 GND 0.030588f
C4816 a_219526_n14006.n263 GND 0.026434f
C4817 a_219526_n14006.n264 GND 0.005132f
C4818 a_219526_n14006.n265 GND 0.019135f
C4819 a_219526_n14006.n266 GND 0.010115f
C4820 a_219526_n14006.n267 GND 0.019178f
C4821 a_219526_n14006.n268 GND 0.010115f
C4822 a_219526_n14006.n269 GND 0.019178f
C4823 a_219526_n14006.n270 GND 0.005132f
C4824 a_219526_n14006.n271 GND 0.019178f
C4825 a_219526_n14006.n272 GND 0.005132f
C4826 a_219526_n14006.n273 GND 0.019178f
C4827 a_219526_n14006.n274 GND 0.005132f
C4828 a_219526_n14006.n275 GND 0.019178f
C4829 a_219526_n14006.n276 GND 0.005132f
C4830 a_219526_n14006.n277 GND 0.019178f
C4831 a_219526_n14006.n278 GND 0.019178f
C4832 a_219526_n14006.n279 GND 0.005132f
C4833 a_219526_n14006.n280 GND 0.009037f
C4834 a_219526_n14006.n281 GND 0.128744f
C4835 a_219526_n14006.n282 GND 0.005434f
C4836 a_219526_n14006.n283 GND 0.005132f
C4837 a_219526_n14006.n284 GND 0.016538f
C4838 a_219526_n14006.n285 GND 0.451349f
C4839 a_219526_n14006.n286 GND 0.419526f
C4840 a_219526_n14006.n287 GND 0.084714f
C4841 a_219526_n14006.n288 GND 0.005132f
C4842 a_219526_n14006.n289 GND 0.005132f
C4843 a_219526_n14006.n290 GND 0.019135f
C4844 a_219526_n14006.n291 GND 0.010115f
C4845 a_219526_n14006.n292 GND 0.019178f
C4846 a_219526_n14006.n293 GND 0.010115f
C4847 a_219526_n14006.n294 GND 0.019178f
C4848 a_219526_n14006.n295 GND 0.005132f
C4849 a_219526_n14006.n296 GND 0.019178f
C4850 a_219526_n14006.n297 GND 0.005132f
C4851 a_219526_n14006.n298 GND 0.019178f
C4852 a_219526_n14006.n299 GND 0.005132f
C4853 a_219526_n14006.n300 GND 0.019178f
C4854 a_219526_n14006.n301 GND 0.005132f
C4855 a_219526_n14006.n302 GND 0.019178f
C4856 a_219526_n14006.n303 GND 0.019178f
C4857 a_219526_n14006.n304 GND 0.005132f
C4858 a_219526_n14006.n305 GND 0.009037f
C4859 a_219526_n14006.n306 GND 0.128744f
C4860 a_219526_n14006.n307 GND 0.009037f
C4861 a_219526_n14006.n308 GND 0.023688f
C4862 a_219526_n14006.n309 GND 0.030321f
C4863 a_219526_n14006.n310 GND 0.257338f
C4864 a_219526_n14006.t16 GND 0.355184f
C4865 a_219526_n14006.n311 GND 0.119739f
C4866 a_219526_n14006.n312 GND 0.37173f
C4867 a_219526_n14006.n313 GND 0.724053f
C4868 a_219526_n14006.t61 GND 0.355184f
C4869 a_219526_n14006.n314 GND 0.404244f
C4870 a_219526_n14006.t51 GND 0.355184f
C4871 a_219526_n14006.n315 GND 0.137608f
C4872 a_219526_n14006.n316 GND 0.137608f
C4873 a_219526_n14006.t54 GND 0.355184f
C4874 a_219526_n14006.n317 GND 0.137608f
C4875 a_219526_n14006.t56 GND 0.355184f
C4876 a_219526_n14006.n318 GND 0.137608f
C4877 a_219526_n14006.n319 GND 0.137608f
C4878 a_219526_n14006.t53 GND 0.355184f
C4879 a_219526_n14006.n320 GND 0.137608f
C4880 a_219526_n14006.t55 GND 0.355184f
C4881 a_219526_n14006.n321 GND 0.137608f
C4882 a_219526_n14006.n322 GND 0.137608f
C4883 a_219526_n14006.t64 GND 0.355184f
C4884 a_219526_n14006.n323 GND 0.137608f
C4885 a_219526_n14006.t67 GND 0.355184f
C4886 a_219526_n14006.n324 GND 0.137608f
C4887 a_219526_n14006.n325 GND 0.122736f
C4888 a_219526_n14006.t50 GND 0.355184f
C4889 a_219526_n14006.n326 GND 0.137608f
C4890 a_219526_n14006.t52 GND 0.355184f
C4891 a_219526_n14006.n327 GND 0.137608f
C4892 a_219526_n14006.n328 GND 0.137608f
C4893 a_219526_n14006.t69 GND 0.355184f
C4894 a_219526_n14006.n329 GND 0.122514f
C4895 a_219526_n14006.t58 GND 0.355184f
C4896 a_219526_n14006.n330 GND 0.137608f
C4897 a_219526_n14006.n331 GND 0.137608f
C4898 a_219526_n14006.t60 GND 0.355184f
C4899 a_219526_n14006.n332 GND 0.137608f
C4900 a_219526_n14006.t63 GND 0.355184f
C4901 a_219526_n14006.n333 GND 0.137608f
C4902 a_219526_n14006.n334 GND 0.137608f
C4903 a_219526_n14006.t66 GND 0.355184f
C4904 a_219526_n14006.n335 GND 0.137608f
C4905 a_219526_n14006.t49 GND 0.355184f
C4906 a_219526_n14006.n336 GND 0.137608f
C4907 a_219526_n14006.n337 GND 0.137608f
C4908 a_219526_n14006.t57 GND 0.355184f
C4909 a_219526_n14006.n338 GND 0.137608f
C4910 a_219526_n14006.t62 GND 0.355184f
C4911 a_219526_n14006.n339 GND 0.137608f
C4912 a_219526_n14006.n340 GND 0.404353f
C4913 a_219526_n14006.t68 GND 0.355184f
C4914 a_219526_n14006.n341 GND 0.086023f
C4915 a_219526_n14006.n342 GND 0.739733f
C4916 a_219526_n14006.t8 GND 0.355184f
C4917 a_219526_n14006.n343 GND 0.26999f
C4918 a_219526_n14006.n344 GND 0.125399f
C4919 a_219526_n14006.t14 GND 0.355184f
C4920 a_219526_n14006.n345 GND 0.119184f
C4921 a_219526_n14006.n346 GND 0.125621f
C4922 a_219526_n14006.t24 GND 0.355184f
C4923 a_219526_n14006.n347 GND 0.125621f
C4924 a_219526_n14006.n348 GND 0.030588f
C4925 a_219526_n14006.n349 GND 0.026434f
C4926 a_219526_n14006.n350 GND 0.005132f
C4927 a_219526_n14006.n351 GND 0.005132f
C4928 a_219526_n14006.n352 GND 0.019135f
C4929 a_219526_n14006.n353 GND 0.010115f
C4930 a_219526_n14006.n354 GND 0.019178f
C4931 a_219526_n14006.n355 GND 0.010115f
C4932 a_219526_n14006.n356 GND 0.019178f
C4933 a_219526_n14006.n357 GND 0.005132f
C4934 a_219526_n14006.n358 GND 0.019178f
C4935 a_219526_n14006.n359 GND 0.005132f
C4936 a_219526_n14006.n360 GND 0.019178f
C4937 a_219526_n14006.n361 GND 0.005132f
C4938 a_219526_n14006.n362 GND 0.019178f
C4939 a_219526_n14006.n363 GND 0.005132f
C4940 a_219526_n14006.n364 GND 0.019178f
C4941 a_219526_n14006.n365 GND 0.019178f
C4942 a_219526_n14006.n366 GND 0.005132f
C4943 a_219526_n14006.n367 GND 0.009037f
C4944 a_219526_n14006.n368 GND 0.128744f
C4945 a_219526_n14006.n369 GND 0.009037f
C4946 a_219526_n14006.n370 GND 0.023688f
C4947 a_219526_n14006.n371 GND 1.29287f
C4948 a_219526_n14006.n372 GND 0.084714f
C4949 a_219526_n14006.n373 GND 0.263581f
C4950 a_219526_n14006.t9 GND 0.064372f
C4951 a_219526_n14006.n374 GND 0.005434f
C4952 a_219526_n14006.n375 GND 0.006774f
C4953 a_219526_n14006.n376 GND 0.014408f
C4954 a_219526_n14006.n377 GND 0.013908f
C4955 a_219526_n14006.n378 GND 0.011863f
C4956 a_219526_n14006.n379 GND 0.011644f
C4957 a_219526_n14006.t3 GND 0.064372f
C4958 a_219526_n14006.n380 GND 0.132696f
C4959 a_219526_n14006.n381 GND 0.504622f
C4960 a_219526_n14006.n382 GND 0.419526f
C4961 a_219526_n14006.n383 GND 0.451349f
C4962 a_219526_n14006.n384 GND 0.005132f
C4963 a_219526_n14006.n385 GND 0.005132f
C4964 a_219526_n14006.n386 GND 0.019135f
C4965 a_219526_n14006.n387 GND 0.010115f
C4966 a_219526_n14006.n388 GND 0.019178f
C4967 a_219526_n14006.n389 GND 0.010115f
C4968 a_219526_n14006.n390 GND 0.019178f
C4969 a_219526_n14006.n391 GND 0.005132f
C4970 a_219526_n14006.n392 GND 0.019178f
C4971 a_219526_n14006.n393 GND 0.005132f
C4972 a_219526_n14006.n394 GND 0.019178f
C4973 a_219526_n14006.n395 GND 0.005132f
C4974 a_219526_n14006.n396 GND 0.019178f
C4975 a_219526_n14006.n397 GND 0.005132f
C4976 a_219526_n14006.n398 GND 0.019178f
C4977 a_219526_n14006.n399 GND 0.005132f
C4978 a_219526_n14006.n400 GND 0.019178f
C4979 a_219526_n14006.n401 GND 0.026434f
C4980 a_219526_n14006.n402 GND 0.030588f
C4981 a_219526_n14006.n403 GND 0.125177f
C4982 a_219526_n14006.t6 GND 0.355184f
C4983 a_219526_n14006.n404 GND 0.125177f
C4984 a_219526_n14006.n405 GND 0.030321f
C4985 a_219526_n14006.n406 GND 0.023688f
C4986 a_219526_n14006.n407 GND 0.009037f
C4987 a_219526_n14006.n408 GND 0.128744f
C4988 a_219526_n14006.t41 GND 0.064372f
C4989 a_216625_n11375.n0 GND 0.150606f
C4990 a_216625_n11375.n1 GND 0.104449f
C4991 a_216625_n11375.n2 GND 0.104449f
C4992 a_216625_n11375.n3 GND 0.103718f
C4993 a_216625_n11375.n4 GND 0.104449f
C4994 a_216625_n11375.t35 GND 0.269595f
C4995 a_216625_n11375.n5 GND 0.103768f
C4996 a_216625_n11375.n6 GND 0.033198f
C4997 a_216625_n11375.n7 GND 0.010247f
C4998 a_216625_n11375.n8 GND 0.195697f
C4999 a_216625_n11375.n9 GND 0.004124f
C5000 a_216625_n11375.n10 GND 0.003895f
C5001 a_216625_n11375.n11 GND 0.01329f
C5002 a_216625_n11375.n12 GND 0.004124f
C5003 a_216625_n11375.n13 GND 0.011088f
C5004 a_216625_n11375.n14 GND 0.003895f
C5005 a_216625_n11375.n15 GND 0.014674f
C5006 a_216625_n11375.n16 GND 0.023503f
C5007 a_216625_n11375.n17 GND 0.004124f
C5008 a_216625_n11375.n18 GND 0.003895f
C5009 a_216625_n11375.n19 GND 0.010936f
C5010 a_216625_n11375.n20 GND 0.01116f
C5011 a_216625_n11375.n21 GND 0.003895f
C5012 a_216625_n11375.n22 GND 0.003895f
C5013 a_216625_n11375.n23 GND 0.004124f
C5014 a_216625_n11375.n24 GND 0.01329f
C5015 a_216625_n11375.n25 GND 0.01329f
C5016 a_216625_n11375.t7 GND 0.019076f
C5017 a_216625_n11375.n26 GND 0.031577f
C5018 a_216625_n11375.n27 GND 0.004835f
C5019 a_216625_n11375.n28 GND 0.009967f
C5020 a_216625_n11375.n29 GND 0.01329f
C5021 a_216625_n11375.n30 GND 0.004124f
C5022 a_216625_n11375.n31 GND 0.003895f
C5023 a_216625_n11375.n32 GND 0.01113f
C5024 a_216625_n11375.n33 GND 0.020747f
C5025 a_216625_n11375.n34 GND 2.57091f
C5026 a_216625_n11375.n35 GND 0.033198f
C5027 a_216625_n11375.n36 GND 0.033198f
C5028 a_216625_n11375.n37 GND 0.033198f
C5029 a_216625_n11375.n38 GND 0.010247f
C5030 a_216625_n11375.t8 GND 0.04886f
C5031 a_216625_n11375.t13 GND 0.04886f
C5032 a_216625_n11375.n39 GND 0.104474f
C5033 a_216625_n11375.n40 GND 0.004124f
C5034 a_216625_n11375.n41 GND 0.011088f
C5035 a_216625_n11375.n42 GND 0.006907f
C5036 a_216625_n11375.n43 GND 0.003895f
C5037 a_216625_n11375.n44 GND 0.004124f
C5038 a_216625_n11375.n45 GND 0.003895f
C5039 a_216625_n11375.n46 GND 0.010936f
C5040 a_216625_n11375.n47 GND 0.01116f
C5041 a_216625_n11375.n48 GND 0.003895f
C5042 a_216625_n11375.n49 GND 0.004124f
C5043 a_216625_n11375.n50 GND 0.009096f
C5044 a_216625_n11375.n51 GND 0.007118f
C5045 a_216625_n11375.n52 GND 0.178986f
C5046 a_216625_n11375.n53 GND 0.427503f
C5047 a_216625_n11375.n54 GND 0.010247f
C5048 a_216625_n11375.t26 GND 0.04886f
C5049 a_216625_n11375.t23 GND 0.04886f
C5050 a_216625_n11375.n55 GND 0.104474f
C5051 a_216625_n11375.n56 GND 0.004124f
C5052 a_216625_n11375.n57 GND 0.011088f
C5053 a_216625_n11375.n58 GND 0.006907f
C5054 a_216625_n11375.n59 GND 0.003895f
C5055 a_216625_n11375.n60 GND 0.004124f
C5056 a_216625_n11375.n61 GND 0.003895f
C5057 a_216625_n11375.n62 GND 0.010936f
C5058 a_216625_n11375.n63 GND 0.01116f
C5059 a_216625_n11375.n64 GND 0.003895f
C5060 a_216625_n11375.n65 GND 0.004124f
C5061 a_216625_n11375.n66 GND 0.009096f
C5062 a_216625_n11375.n67 GND 0.007118f
C5063 a_216625_n11375.n68 GND 0.178986f
C5064 a_216625_n11375.n69 GND 0.427503f
C5065 a_216625_n11375.n70 GND 0.010247f
C5066 a_216625_n11375.t24 GND 0.04886f
C5067 a_216625_n11375.t22 GND 0.04886f
C5068 a_216625_n11375.n71 GND 0.104474f
C5069 a_216625_n11375.n72 GND 0.004124f
C5070 a_216625_n11375.n73 GND 0.011088f
C5071 a_216625_n11375.n74 GND 0.006907f
C5072 a_216625_n11375.n75 GND 0.003895f
C5073 a_216625_n11375.n76 GND 0.004124f
C5074 a_216625_n11375.n77 GND 0.003895f
C5075 a_216625_n11375.n78 GND 0.010936f
C5076 a_216625_n11375.n79 GND 0.01116f
C5077 a_216625_n11375.n80 GND 0.003895f
C5078 a_216625_n11375.n81 GND 0.004124f
C5079 a_216625_n11375.n82 GND 0.009096f
C5080 a_216625_n11375.n83 GND 0.007118f
C5081 a_216625_n11375.n84 GND 0.178986f
C5082 a_216625_n11375.n85 GND 2.76314f
C5083 a_216625_n11375.n86 GND 0.103175f
C5084 a_216625_n11375.n87 GND 0.103465f
C5085 a_216625_n11375.n88 GND 0.104449f
C5086 a_216625_n11375.n89 GND 0.104449f
C5087 a_216625_n11375.n90 GND 0.150771f
C5088 a_216625_n11375.t31 GND 0.932339f
C5089 a_216625_n11375.t10 GND 0.833027f
C5090 a_216625_n11375.n91 GND 9.08508f
C5091 a_216625_n11375.n92 GND 0.609697f
C5092 a_216625_n11375.t62 GND 0.269595f
C5093 a_216625_n11375.n93 GND 0.154543f
C5094 a_216625_n11375.n94 GND 0.104449f
C5095 a_216625_n11375.t44 GND 0.269595f
C5096 a_216625_n11375.n95 GND 0.104449f
C5097 a_216625_n11375.t32 GND 0.269595f
C5098 a_216625_n11375.n96 GND 0.104449f
C5099 a_216625_n11375.n97 GND 0.104449f
C5100 a_216625_n11375.t37 GND 0.269595f
C5101 a_216625_n11375.n98 GND 0.104449f
C5102 a_216625_n11375.t45 GND 0.269595f
C5103 a_216625_n11375.n99 GND 0.104449f
C5104 a_216625_n11375.n100 GND 0.104449f
C5105 a_216625_n11375.t50 GND 0.269595f
C5106 a_216625_n11375.n101 GND 0.104449f
C5107 a_216625_n11375.t66 GND 0.269595f
C5108 a_216625_n11375.n102 GND 0.104449f
C5109 a_216625_n11375.n103 GND 0.104449f
C5110 a_216625_n11375.n104 GND 0.104449f
C5111 a_216625_n11375.n105 GND 0.104449f
C5112 a_216625_n11375.n106 GND 0.104449f
C5113 a_216625_n11375.n107 GND 0.104449f
C5114 a_216625_n11375.n108 GND 0.104449f
C5115 a_216625_n11375.n109 GND 0.104449f
C5116 a_216625_n11375.n110 GND 0.104449f
C5117 a_216625_n11375.n111 GND 0.104449f
C5118 a_216625_n11375.n112 GND 0.104449f
C5119 a_216625_n11375.n113 GND 0.104449f
C5120 a_216625_n11375.t52 GND 0.269595f
C5121 a_216625_n11375.n114 GND 0.104449f
C5122 a_216625_n11375.n115 GND 0.104449f
C5123 a_216625_n11375.t47 GND 0.269595f
C5124 a_216625_n11375.n116 GND 0.104449f
C5125 a_216625_n11375.t43 GND 0.269595f
C5126 a_216625_n11375.n117 GND 0.104449f
C5127 a_216625_n11375.n118 GND 0.104449f
C5128 a_216625_n11375.t34 GND 0.269595f
C5129 a_216625_n11375.n119 GND 0.104449f
C5130 a_216625_n11375.t70 GND 0.269595f
C5131 a_216625_n11375.n120 GND 0.104449f
C5132 a_216625_n11375.n121 GND 0.104449f
C5133 a_216625_n11375.t49 GND 0.269595f
C5134 a_216625_n11375.n122 GND 0.104449f
C5135 a_216625_n11375.t48 GND 0.269595f
C5136 a_216625_n11375.n123 GND 0.104449f
C5137 a_216625_n11375.n124 GND 0.104449f
C5138 a_216625_n11375.t40 GND 0.269595f
C5139 a_216625_n11375.n125 GND 0.104449f
C5140 a_216625_n11375.t68 GND 0.269595f
C5141 a_216625_n11375.n126 GND 0.104449f
C5142 a_216625_n11375.n127 GND 0.104449f
C5143 a_216625_n11375.t64 GND 0.269595f
C5144 a_216625_n11375.n128 GND 0.104449f
C5145 a_216625_n11375.t60 GND 0.269595f
C5146 a_216625_n11375.n129 GND 0.104449f
C5147 a_216625_n11375.n130 GND 0.104449f
C5148 a_216625_n11375.t57 GND 0.269595f
C5149 a_216625_n11375.n131 GND 0.104449f
C5150 a_216625_n11375.t51 GND 0.269595f
C5151 a_216625_n11375.n132 GND 0.104449f
C5152 a_216625_n11375.n133 GND 0.104449f
C5153 a_216625_n11375.t46 GND 0.269595f
C5154 a_216625_n11375.n134 GND 0.104449f
C5155 a_216625_n11375.t42 GND 0.269595f
C5156 a_216625_n11375.n135 GND 0.104449f
C5157 a_216625_n11375.n136 GND 0.104449f
C5158 a_216625_n11375.t56 GND 0.269595f
C5159 a_216625_n11375.n137 GND 0.104449f
C5160 a_216625_n11375.t55 GND 0.269595f
C5161 a_216625_n11375.n138 GND 0.104449f
C5162 a_216625_n11375.n139 GND 0.104449f
C5163 a_216625_n11375.t63 GND 0.269595f
C5164 a_216625_n11375.n140 GND 0.104449f
C5165 a_216625_n11375.t59 GND 0.269595f
C5166 a_216625_n11375.n141 GND 0.104449f
C5167 a_216625_n11375.n142 GND 0.104449f
C5168 a_216625_n11375.t53 GND 0.269595f
C5169 a_216625_n11375.n143 GND 0.104449f
C5170 a_216625_n11375.t33 GND 0.269595f
C5171 a_216625_n11375.n144 GND 0.104449f
C5172 a_216625_n11375.n145 GND 0.104449f
C5173 a_216625_n11375.t67 GND 0.269595f
C5174 a_216625_n11375.n146 GND 0.104449f
C5175 a_216625_n11375.t58 GND 0.269595f
C5176 a_216625_n11375.n147 GND 0.104449f
C5177 a_216625_n11375.n148 GND 0.104449f
C5178 a_216625_n11375.t38 GND 0.269595f
C5179 a_216625_n11375.n149 GND 0.107487f
C5180 a_216625_n11375.n150 GND 0.110891f
C5181 a_216625_n11375.n151 GND 1.82882f
C5182 a_216625_n11375.n152 GND 0.02041f
C5183 a_216625_n11375.n153 GND 0.011088f
C5184 a_216625_n11375.n154 GND 0.003895f
C5185 a_216625_n11375.n155 GND 0.01329f
C5186 a_216625_n11375.n156 GND 0.004124f
C5187 a_216625_n11375.n157 GND 0.003895f
C5188 a_216625_n11375.n158 GND 0.01329f
C5189 a_216625_n11375.n159 GND 0.004124f
C5190 a_216625_n11375.n160 GND 0.032372f
C5191 a_216625_n11375.t20 GND 0.024889f
C5192 a_216625_n11375.n161 GND 0.009967f
C5193 a_216625_n11375.n162 GND 0.005094f
C5194 a_216625_n11375.n163 GND 0.003895f
C5195 a_216625_n11375.n164 GND 0.189103f
C5196 a_216625_n11375.n165 GND 0.010921f
C5197 a_216625_n11375.n166 GND 0.011123f
C5198 a_216625_n11375.n167 GND 0.003895f
C5199 a_216625_n11375.n168 GND 0.004124f
C5200 a_216625_n11375.n169 GND 0.01329f
C5201 a_216625_n11375.n170 GND 0.01329f
C5202 a_216625_n11375.n171 GND 0.004124f
C5203 a_216625_n11375.n172 GND 0.003895f
C5204 a_216625_n11375.n173 GND 0.010557f
C5205 a_216625_n11375.n174 GND 0.010936f
C5206 a_216625_n11375.n175 GND 0.003895f
C5207 a_216625_n11375.n176 GND 0.004124f
C5208 a_216625_n11375.n177 GND 0.026181f
C5209 a_216625_n11375.n178 GND 0.011997f
C5210 a_216625_n11375.n179 GND 0.033198f
C5211 a_216625_n11375.n180 GND 0.621914f
C5212 a_216625_n11375.n181 GND 0.200066f
C5213 a_216625_n11375.n182 GND 0.011088f
C5214 a_216625_n11375.n183 GND 0.003895f
C5215 a_216625_n11375.t16 GND 0.04886f
C5216 a_216625_n11375.n184 GND 0.004124f
C5217 a_216625_n11375.n185 GND 0.004124f
C5218 a_216625_n11375.n186 GND 0.003895f
C5219 a_216625_n11375.n187 GND 0.010936f
C5220 a_216625_n11375.n188 GND 0.010557f
C5221 a_216625_n11375.n189 GND 0.009005f
C5222 a_216625_n11375.n190 GND 0.008838f
C5223 a_216625_n11375.t2 GND 0.04886f
C5224 a_216625_n11375.n191 GND 0.100636f
C5225 a_216625_n11375.n192 GND 0.006907f
C5226 a_216625_n11375.n193 GND 0.033198f
C5227 a_216625_n11375.n194 GND 0.342588f
C5228 a_216625_n11375.n195 GND 0.200066f
C5229 a_216625_n11375.n196 GND 0.011088f
C5230 a_216625_n11375.n197 GND 0.003895f
C5231 a_216625_n11375.t3 GND 0.04886f
C5232 a_216625_n11375.n198 GND 0.004124f
C5233 a_216625_n11375.n199 GND 0.004124f
C5234 a_216625_n11375.n200 GND 0.003895f
C5235 a_216625_n11375.n201 GND 0.010936f
C5236 a_216625_n11375.n202 GND 0.010557f
C5237 a_216625_n11375.n203 GND 0.009005f
C5238 a_216625_n11375.n204 GND 0.008838f
C5239 a_216625_n11375.t21 GND 0.04886f
C5240 a_216625_n11375.n205 GND 0.100636f
C5241 a_216625_n11375.n206 GND 0.006907f
C5242 a_216625_n11375.n207 GND 0.033198f
C5243 a_216625_n11375.n208 GND 0.347642f
C5244 a_216625_n11375.n209 GND 0.200066f
C5245 a_216625_n11375.n210 GND 0.011088f
C5246 a_216625_n11375.n211 GND 0.003895f
C5247 a_216625_n11375.t9 GND 0.04886f
C5248 a_216625_n11375.n212 GND 0.004124f
C5249 a_216625_n11375.n213 GND 0.004124f
C5250 a_216625_n11375.n214 GND 0.003895f
C5251 a_216625_n11375.n215 GND 0.010936f
C5252 a_216625_n11375.n216 GND 0.010557f
C5253 a_216625_n11375.n217 GND 0.009005f
C5254 a_216625_n11375.n218 GND 0.008838f
C5255 a_216625_n11375.t4 GND 0.04886f
C5256 a_216625_n11375.n219 GND 0.100636f
C5257 a_216625_n11375.n220 GND 0.006907f
C5258 a_216625_n11375.n221 GND 0.033198f
C5259 a_216625_n11375.n222 GND 0.342588f
C5260 a_216625_n11375.n223 GND 0.200066f
C5261 a_216625_n11375.n224 GND 0.011088f
C5262 a_216625_n11375.n225 GND 0.003895f
C5263 a_216625_n11375.t17 GND 0.04886f
C5264 a_216625_n11375.n226 GND 0.004124f
C5265 a_216625_n11375.n227 GND 0.004124f
C5266 a_216625_n11375.n228 GND 0.003895f
C5267 a_216625_n11375.n229 GND 0.010936f
C5268 a_216625_n11375.n230 GND 0.010557f
C5269 a_216625_n11375.n231 GND 0.009005f
C5270 a_216625_n11375.n232 GND 0.008838f
C5271 a_216625_n11375.t15 GND 0.04886f
C5272 a_216625_n11375.n233 GND 0.100636f
C5273 a_216625_n11375.n234 GND 0.006907f
C5274 a_216625_n11375.n235 GND 0.033198f
C5275 a_216625_n11375.n236 GND 0.342588f
C5276 a_216625_n11375.n237 GND 0.200066f
C5277 a_216625_n11375.n238 GND 0.011088f
C5278 a_216625_n11375.n239 GND 0.003895f
C5279 a_216625_n11375.t6 GND 0.04886f
C5280 a_216625_n11375.n240 GND 0.004124f
C5281 a_216625_n11375.n241 GND 0.004124f
C5282 a_216625_n11375.n242 GND 0.003895f
C5283 a_216625_n11375.n243 GND 0.010936f
C5284 a_216625_n11375.n244 GND 0.010557f
C5285 a_216625_n11375.n245 GND 0.009005f
C5286 a_216625_n11375.n246 GND 0.008838f
C5287 a_216625_n11375.t18 GND 0.04886f
C5288 a_216625_n11375.n247 GND 0.100636f
C5289 a_216625_n11375.n248 GND 0.006907f
C5290 a_216625_n11375.n249 GND 0.033198f
C5291 a_216625_n11375.n250 GND 0.342588f
C5292 a_216625_n11375.n251 GND 0.200066f
C5293 a_216625_n11375.n252 GND 0.011088f
C5294 a_216625_n11375.n253 GND 0.003895f
C5295 a_216625_n11375.t28 GND 0.04886f
C5296 a_216625_n11375.n254 GND 0.004124f
C5297 a_216625_n11375.n255 GND 0.004124f
C5298 a_216625_n11375.n256 GND 0.003895f
C5299 a_216625_n11375.n257 GND 0.010936f
C5300 a_216625_n11375.n258 GND 0.010557f
C5301 a_216625_n11375.n259 GND 0.009005f
C5302 a_216625_n11375.n260 GND 0.008838f
C5303 a_216625_n11375.t29 GND 0.04886f
C5304 a_216625_n11375.n261 GND 0.100636f
C5305 a_216625_n11375.n262 GND 0.006907f
C5306 a_216625_n11375.n263 GND 0.033198f
C5307 a_216625_n11375.n264 GND 0.342588f
C5308 a_216625_n11375.n265 GND 0.200066f
C5309 a_216625_n11375.n266 GND 0.011088f
C5310 a_216625_n11375.n267 GND 0.003895f
C5311 a_216625_n11375.t27 GND 0.04886f
C5312 a_216625_n11375.n268 GND 0.004124f
C5313 a_216625_n11375.n269 GND 0.004124f
C5314 a_216625_n11375.n270 GND 0.003895f
C5315 a_216625_n11375.n271 GND 0.010936f
C5316 a_216625_n11375.n272 GND 0.010557f
C5317 a_216625_n11375.n273 GND 0.009005f
C5318 a_216625_n11375.n274 GND 0.008838f
C5319 a_216625_n11375.t11 GND 0.04886f
C5320 a_216625_n11375.n275 GND 0.100636f
C5321 a_216625_n11375.n276 GND 0.006907f
C5322 a_216625_n11375.n277 GND 0.033198f
C5323 a_216625_n11375.n278 GND 0.347642f
C5324 a_216625_n11375.n279 GND 0.200066f
C5325 a_216625_n11375.n280 GND 0.011088f
C5326 a_216625_n11375.n281 GND 0.003895f
C5327 a_216625_n11375.t14 GND 0.04886f
C5328 a_216625_n11375.n282 GND 0.004124f
C5329 a_216625_n11375.n283 GND 0.004124f
C5330 a_216625_n11375.n284 GND 0.003895f
C5331 a_216625_n11375.n285 GND 0.010936f
C5332 a_216625_n11375.n286 GND 0.010557f
C5333 a_216625_n11375.n287 GND 0.009005f
C5334 a_216625_n11375.n288 GND 0.008838f
C5335 a_216625_n11375.t5 GND 0.04886f
C5336 a_216625_n11375.n289 GND 0.100636f
C5337 a_216625_n11375.n290 GND 0.006907f
C5338 a_216625_n11375.n291 GND 0.033198f
C5339 a_216625_n11375.n292 GND 0.342588f
C5340 a_216625_n11375.n293 GND 0.200066f
C5341 a_216625_n11375.n294 GND 0.011088f
C5342 a_216625_n11375.n295 GND 0.003895f
C5343 a_216625_n11375.t19 GND 0.04886f
C5344 a_216625_n11375.n296 GND 0.004124f
C5345 a_216625_n11375.n297 GND 0.004124f
C5346 a_216625_n11375.n298 GND 0.003895f
C5347 a_216625_n11375.n299 GND 0.010936f
C5348 a_216625_n11375.n300 GND 0.010557f
C5349 a_216625_n11375.n301 GND 0.009005f
C5350 a_216625_n11375.n302 GND 0.008838f
C5351 a_216625_n11375.t1 GND 0.04886f
C5352 a_216625_n11375.n303 GND 0.100636f
C5353 a_216625_n11375.n304 GND 0.006907f
C5354 a_216625_n11375.n305 GND 0.033198f
C5355 a_216625_n11375.n306 GND 0.342588f
C5356 a_216625_n11375.n307 GND 0.200066f
C5357 a_216625_n11375.n308 GND 0.011088f
C5358 a_216625_n11375.n309 GND 0.003895f
C5359 a_216625_n11375.t25 GND 0.04886f
C5360 a_216625_n11375.n310 GND 0.004124f
C5361 a_216625_n11375.n311 GND 0.004124f
C5362 a_216625_n11375.n312 GND 0.003895f
C5363 a_216625_n11375.n313 GND 0.010936f
C5364 a_216625_n11375.n314 GND 0.010557f
C5365 a_216625_n11375.n315 GND 0.009005f
C5366 a_216625_n11375.n316 GND 0.008838f
C5367 a_216625_n11375.t30 GND 0.04886f
C5368 a_216625_n11375.n317 GND 0.100636f
C5369 a_216625_n11375.n318 GND 0.006907f
C5370 a_216625_n11375.n319 GND 0.033198f
C5371 a_216625_n11375.n320 GND 0.790823f
C5372 a_216625_n11375.n321 GND 1.82417f
C5373 a_216625_n11375.n322 GND 0.110583f
C5374 a_216625_n11375.n323 GND 0.106949f
C5375 a_216625_n11375.t39 GND 0.269595f
C5376 a_216625_n11375.n324 GND 0.104449f
C5377 a_216625_n11375.t65 GND 0.269595f
C5378 a_216625_n11375.n325 GND 0.104449f
C5379 a_216625_n11375.n326 GND 0.104449f
C5380 a_216625_n11375.t69 GND 0.269595f
C5381 a_216625_n11375.n327 GND 0.104449f
C5382 a_216625_n11375.t41 GND 0.269595f
C5383 a_216625_n11375.n328 GND 0.104449f
C5384 a_216625_n11375.n329 GND 0.104449f
C5385 a_216625_n11375.t54 GND 0.269595f
C5386 a_216625_n11375.n330 GND 0.104449f
C5387 a_216625_n11375.t61 GND 0.269595f
C5388 a_216625_n11375.n331 GND 0.104449f
C5389 a_216625_n11375.n332 GND 0.104449f
C5390 a_216625_n11375.t71 GND 0.269595f
C5391 a_216625_n11375.n333 GND 0.104449f
C5392 a_216625_n11375.t36 GND 0.269595f
C5393 a_216625_n11375.n334 GND 0.154394f
C5394 a_216625_n11375.n335 GND 0.607988f
C5395 a_216625_n11375.t12 GND 0.829336f
C5396 a_216625_n11375.n336 GND 9.19451f
C5397 a_216625_n11375.t0 GND 0.929383f
C5398 VDD.n0 GND 2.06594f
C5399 VDD.n1 GND 1.88886f
C5400 VDD.n3 GND 1.88886f
C5401 VDD.n5 GND 0.335437f
C5402 VDD.n6 GND 0.005467f
C5403 VDD.n7 GND 0.002367f
C5404 VDD.n8 GND 8.53e-19
C5405 VDD.n9 GND 0.00291f
C5406 VDD.n10 GND 9.03e-19
C5407 VDD.n11 GND 0.007088f
C5408 VDD.t125 GND 0.00545f
C5409 VDD.n12 GND 0.002183f
C5410 VDD.n13 GND 0.001115f
C5411 VDD.n14 GND 8.53e-19
C5412 VDD.n15 GND 0.041407f
C5413 VDD.n16 GND 0.002444f
C5414 VDD.n17 GND 8.53e-19
C5415 VDD.n18 GND 9.03e-19
C5416 VDD.n19 GND 0.00291f
C5417 VDD.n20 GND 0.006447f
C5418 VDD.n21 GND 9.03e-19
C5419 VDD.n22 GND 0.00116f
C5420 VDD.n23 GND 0.002806f
C5421 VDD.n24 GND 0.018731f
C5422 VDD.n25 GND 0.12073f
C5423 VDD.n26 GND 0.018612f
C5424 VDD.n27 GND 0.011119f
C5425 VDD.n28 GND 0.001062f
C5426 VDD.n29 GND 0.001706f
C5427 VDD.n31 GND 0.247293f
C5428 VDD.n32 GND 0.001706f
C5429 VDD.n33 GND 0.001706f
C5430 VDD.n35 GND 0.003712f
C5431 VDD.n36 GND 0.001706f
C5432 VDD.n37 GND 0.001706f
C5433 VDD.n38 GND 0.188724f
C5434 VDD.n39 GND 0.001706f
C5435 VDD.n40 GND 0.074839f
C5436 VDD.n41 GND 0.001706f
C5437 VDD.n42 GND 0.003712f
C5438 VDD.n43 GND 0.001706f
C5439 VDD.n44 GND 0.003712f
C5440 VDD.n45 GND 0.001706f
C5441 VDD.n46 GND 0.001706f
C5442 VDD.t121 GND 0.073754f
C5443 VDD.n47 GND 0.001706f
C5444 VDD.n48 GND 0.001706f
C5445 VDD.n49 GND 0.147508f
C5446 VDD.n50 GND 0.001706f
C5447 VDD.n51 GND 0.001706f
C5448 VDD.n52 GND 0.003714f
C5449 VDD.n53 GND 0.001706f
C5450 VDD.n54 GND 0.001706f
C5451 VDD.n55 GND 0.001706f
C5452 VDD.n57 GND 0.001706f
C5453 VDD.n58 GND 0.001003f
C5454 VDD.n60 GND 0.001706f
C5455 VDD.n61 GND 0.001706f
C5456 VDD.n62 GND 0.001062f
C5457 VDD.n63 GND 0.001003f
C5458 VDD.n64 GND 0.001149f
C5459 VDD.n65 GND 0.001704f
C5460 VDD.n66 GND 0.001706f
C5461 VDD.n68 GND 0.001706f
C5462 VDD.n69 GND 0.001706f
C5463 VDD.n70 GND 0.001706f
C5464 VDD.n71 GND 0.001706f
C5465 VDD.n72 GND 0.001706f
C5466 VDD.n73 GND 0.001706f
C5467 VDD.n75 GND 0.001706f
C5468 VDD.n76 GND 0.003714f
C5469 VDD.n77 GND 0.003712f
C5470 VDD.n78 GND 0.003712f
C5471 VDD.n79 GND 0.001706f
C5472 VDD.n80 GND 0.001706f
C5473 VDD.n81 GND 0.001706f
C5474 VDD.n82 GND 0.001706f
C5475 VDD.n83 GND 0.001706f
C5476 VDD.n84 GND 0.001706f
C5477 VDD.t105 GND 0.073754f
C5478 VDD.n85 GND 0.001706f
C5479 VDD.n86 GND 0.001706f
C5480 VDD.n87 GND 0.001706f
C5481 VDD.n88 GND 0.087854f
C5482 VDD.n89 GND 0.001706f
C5483 VDD.n90 GND 0.001706f
C5484 VDD.n91 GND 0.147508f
C5485 VDD.n92 GND 0.001706f
C5486 VDD.n93 GND 0.001706f
C5487 VDD.n94 GND 0.001706f
C5488 VDD.n95 GND 0.001706f
C5489 VDD.n96 GND 0.001706f
C5490 VDD.t31 GND 0.073754f
C5491 VDD.n97 GND 0.001706f
C5492 VDD.n98 GND 0.001706f
C5493 VDD.n99 GND 0.001706f
C5494 VDD.n100 GND 0.103039f
C5495 VDD.n101 GND 0.001706f
C5496 VDD.n102 GND 0.001706f
C5497 VDD.n103 GND 0.147508f
C5498 VDD.n104 GND 0.001706f
C5499 VDD.n105 GND 0.001706f
C5500 VDD.n106 GND 0.001706f
C5501 VDD.n107 GND 0.001706f
C5502 VDD.n108 GND 0.001706f
C5503 VDD.t29 GND 0.073754f
C5504 VDD.n109 GND 0.001706f
C5505 VDD.n110 GND 0.001706f
C5506 VDD.n111 GND 0.001706f
C5507 VDD.n112 GND 0.118224f
C5508 VDD.n113 GND 0.001706f
C5509 VDD.n114 GND 0.001706f
C5510 VDD.n115 GND 0.147508f
C5511 VDD.n116 GND 0.001706f
C5512 VDD.n117 GND 0.001706f
C5513 VDD.n118 GND 0.001706f
C5514 VDD.n119 GND 0.001706f
C5515 VDD.n120 GND 0.001706f
C5516 VDD.t343 GND 0.073754f
C5517 VDD.n121 GND 0.001706f
C5518 VDD.n122 GND 0.001706f
C5519 VDD.n123 GND 0.001706f
C5520 VDD.n124 GND 0.133408f
C5521 VDD.n125 GND 0.001706f
C5522 VDD.n126 GND 0.001706f
C5523 VDD.n127 GND 0.146424f
C5524 VDD.n128 GND 0.001706f
C5525 VDD.n129 GND 0.001706f
C5526 VDD.n130 GND 0.001706f
C5527 VDD.t123 GND 0.073754f
C5528 VDD.n131 GND 0.001706f
C5529 VDD.n132 GND 0.001706f
C5530 VDD.n133 GND 0.147508f
C5531 VDD.n134 GND 0.001706f
C5532 VDD.n135 GND 0.003714f
C5533 VDD.n136 GND 0.003714f
C5534 VDD.n137 GND 0.003712f
C5535 VDD.n138 GND 0.003712f
C5536 VDD.n139 GND 0.229939f
C5537 VDD.n140 GND 0.003714f
C5538 VDD.n141 GND 0.001706f
C5539 VDD.n142 GND 0.001706f
C5540 VDD.n143 GND 0.001704f
C5541 VDD.n144 GND 0.001706f
C5542 VDD.n145 GND 0.001062f
C5543 VDD.t705 GND 0.010699f
C5544 VDD.t706 GND 0.010699f
C5545 VDD.n146 GND 0.032273f
C5546 VDD.n147 GND 0.107301f
C5547 VDD.n148 GND 0.005784f
C5548 VDD.n149 GND 0.005969f
C5549 VDD.n150 GND 8.53e-19
C5550 VDD.n151 GND 0.002183f
C5551 VDD.n152 GND 8.78e-19
C5552 VDD.n153 GND 0.004516f
C5553 VDD.n154 GND 0.004516f
C5554 VDD.n155 GND 0.001062f
C5555 VDD.t252 GND 0.001455f
C5556 VDD.n156 GND 0.005656f
C5557 VDD.n157 GND 8.78e-19
C5558 VDD.n158 GND 0.001115f
C5559 VDD.n159 GND 0.00636f
C5560 VDD.n160 GND 0.041968f
C5561 VDD.n161 GND 0.001022f
C5562 VDD.n162 GND 0.001706f
C5563 VDD.n163 GND 0.001706f
C5564 VDD.n164 GND 0.001706f
C5565 VDD.n166 GND 0.001706f
C5566 VDD.n167 GND 0.001706f
C5567 VDD.n168 GND 0.001706f
C5568 VDD.n169 GND 0.001706f
C5569 VDD.n170 GND 0.001706f
C5570 VDD.n172 GND 0.001706f
C5571 VDD.n174 GND 0.001706f
C5572 VDD.n175 GND 0.001706f
C5573 VDD.n176 GND 0.00173f
C5574 VDD.n177 GND 0.002023f
C5575 VDD.n178 GND 0.001706f
C5576 VDD.n180 GND 0.001706f
C5577 VDD.n181 GND 0.001706f
C5578 VDD.n182 GND 0.001706f
C5579 VDD.n183 GND 0.001706f
C5580 VDD.n184 GND 0.003714f
C5581 VDD.n185 GND 0.001706f
C5582 VDD.n186 GND 0.001706f
C5583 VDD.n187 GND 0.001706f
C5584 VDD.n188 GND 0.001062f
C5585 VDD.n189 GND 0.004516f
C5586 VDD.n190 GND 0.005656f
C5587 VDD.n191 GND 8.53e-19
C5588 VDD.n192 GND 0.006434f
C5589 VDD.n193 GND 9.03e-19
C5590 VDD.t253 GND 0.010699f
C5591 VDD.t254 GND 0.010699f
C5592 VDD.n194 GND 0.032273f
C5593 VDD.n195 GND 0.229486f
C5594 VDD.n196 GND 0.586149f
C5595 VDD.n197 GND 0.107744f
C5596 VDD.n198 GND 0.030806f
C5597 VDD.n199 GND 0.025832f
C5598 VDD.n200 GND 0.005784f
C5599 VDD.n201 GND 0.001162f
C5600 VDD.n202 GND 0.0023f
C5601 VDD.n203 GND 0.004516f
C5602 VDD.n204 GND 0.00173f
C5603 VDD.n205 GND 0.001706f
C5604 VDD.n206 GND 0.001706f
C5605 VDD.n207 GND 0.001706f
C5606 VDD.n208 GND 0.003714f
C5607 VDD.n209 GND 0.003714f
C5608 VDD.n211 GND 0.001706f
C5609 VDD.n213 GND 0.001706f
C5610 VDD.n214 GND 0.001706f
C5611 VDD.n215 GND 0.001706f
C5612 VDD.n216 GND 0.001706f
C5613 VDD.n217 GND 0.001706f
C5614 VDD.n219 GND 0.001706f
C5615 VDD.n220 GND 0.001706f
C5616 VDD.n221 GND 0.001706f
C5617 VDD.n222 GND 0.004516f
C5618 VDD.n223 GND 0.001003f
C5619 VDD.n225 GND 0.001706f
C5620 VDD.n227 GND 0.001706f
C5621 VDD.n228 GND 0.001062f
C5622 VDD.n229 GND 0.002023f
C5623 VDD.n230 GND 0.004516f
C5624 VDD.n231 GND 0.005969f
C5625 VDD.n232 GND 8.53e-19
C5626 VDD.n233 GND 9.03e-19
C5627 VDD.n234 GND 0.00291f
C5628 VDD.t122 GND 0.001455f
C5629 VDD.n235 GND 0.002183f
C5630 VDD.n236 GND 8.78e-19
C5631 VDD.n237 GND 8.78e-19
C5632 VDD.n238 GND 0.001115f
C5633 VDD.n239 GND 0.00636f
C5634 VDD.n240 GND 0.041968f
C5635 VDD.n241 GND 0.001022f
C5636 VDD.n242 GND 0.001645f
C5637 VDD.n243 GND 0.001706f
C5638 VDD.n244 GND 0.001706f
C5639 VDD.n246 GND 0.001706f
C5640 VDD.n248 GND 0.001706f
C5641 VDD.n249 GND 0.001706f
C5642 VDD.n250 GND 0.001706f
C5643 VDD.n251 GND 0.001706f
C5644 VDD.n252 GND 0.001706f
C5645 VDD.n254 GND 0.003714f
C5646 VDD.n255 GND 0.003712f
C5647 VDD.n256 GND 0.003712f
C5648 VDD.n257 GND 0.001706f
C5649 VDD.n258 GND 0.001706f
C5650 VDD.n259 GND 0.001706f
C5651 VDD.n260 GND 0.001706f
C5652 VDD.n261 GND 0.001706f
C5653 VDD.n262 GND 0.001706f
C5654 VDD.n263 GND 0.001706f
C5655 VDD.n264 GND 0.001706f
C5656 VDD.n265 GND 0.001706f
C5657 VDD.n266 GND 0.001706f
C5658 VDD.n267 GND 0.001706f
C5659 VDD.n268 GND 0.001706f
C5660 VDD.n269 GND 0.001706f
C5661 VDD.n270 GND 0.001706f
C5662 VDD.n271 GND 0.001706f
C5663 VDD.n272 GND 0.001706f
C5664 VDD.n273 GND 0.001706f
C5665 VDD.n274 GND 0.001706f
C5666 VDD.n275 GND 0.001706f
C5667 VDD.n276 GND 0.001706f
C5668 VDD.n277 GND 0.001706f
C5669 VDD.n278 GND 0.001706f
C5670 VDD.n279 GND 0.001706f
C5671 VDD.n280 GND 0.001706f
C5672 VDD.n281 GND 0.001706f
C5673 VDD.n282 GND 0.001706f
C5674 VDD.n283 GND 0.001706f
C5675 VDD.n284 GND 0.001706f
C5676 VDD.n285 GND 0.001706f
C5677 VDD.n286 GND 0.001706f
C5678 VDD.n287 GND 0.001706f
C5679 VDD.n288 GND 0.001706f
C5680 VDD.n289 GND 0.001706f
C5681 VDD.n290 GND 0.003712f
C5682 VDD.n292 GND 0.003714f
C5683 VDD.n293 GND 0.003714f
C5684 VDD.n294 GND 0.001706f
C5685 VDD.n295 GND 0.001706f
C5686 VDD.n296 GND 0.001706f
C5687 VDD.n298 GND 0.001706f
C5688 VDD.n300 GND 0.001706f
C5689 VDD.n301 GND 0.001706f
C5690 VDD.n302 GND 0.001706f
C5691 VDD.n303 GND 0.001645f
C5692 VDD.n304 GND 0.001706f
C5693 VDD.n306 GND 0.001706f
C5694 VDD.n307 GND 0.001062f
C5695 VDD.n308 GND 0.001003f
C5696 VDD.n309 GND 0.004516f
C5697 VDD.n310 GND 0.004516f
C5698 VDD.n311 GND 8.53e-19
C5699 VDD.n312 GND 9.03e-19
C5700 VDD.n313 GND 0.00291f
C5701 VDD.n314 GND 0.006434f
C5702 VDD.n315 GND 9.03e-19
C5703 VDD.n316 GND 0.001162f
C5704 VDD.n317 GND 0.0023f
C5705 VDD.n318 GND 0.025832f
C5706 VDD.n319 GND 0.033011f
C5707 VDD.n320 GND 0.172693f
C5708 VDD.t106 GND 0.010699f
C5709 VDD.t32 GND 0.010699f
C5710 VDD.n321 GND 0.032325f
C5711 VDD.n322 GND 0.102342f
C5712 VDD.t30 GND 0.010699f
C5713 VDD.t344 GND 0.010699f
C5714 VDD.n323 GND 0.032325f
C5715 VDD.n324 GND 0.102988f
C5716 VDD.n325 GND 0.005467f
C5717 VDD.n326 GND 0.002367f
C5718 VDD.n327 GND 8.53e-19
C5719 VDD.n328 GND 0.00291f
C5720 VDD.n329 GND 9.03e-19
C5721 VDD.n330 GND 0.007088f
C5722 VDD.t124 GND 0.00545f
C5723 VDD.n331 GND 0.002183f
C5724 VDD.n332 GND 0.001115f
C5725 VDD.n333 GND 8.53e-19
C5726 VDD.n334 GND 0.041407f
C5727 VDD.n335 GND 0.002444f
C5728 VDD.n336 GND 8.53e-19
C5729 VDD.n337 GND 9.03e-19
C5730 VDD.n338 GND 0.00291f
C5731 VDD.n339 GND 0.006447f
C5732 VDD.n340 GND 9.03e-19
C5733 VDD.n341 GND 0.00116f
C5734 VDD.n342 GND 0.002806f
C5735 VDD.n343 GND 0.018731f
C5736 VDD.n344 GND 0.052956f
C5737 VDD.n345 GND 0.192513f
C5738 VDD.n346 GND 0.031168f
C5739 VDD.n347 GND 0.017532f
C5740 VDD.n348 GND 0.00102f
C5741 VDD.n350 GND 0.001706f
C5742 VDD.n351 GND 0.001706f
C5743 VDD.n352 GND 0.001706f
C5744 VDD.n353 GND 0.001706f
C5745 VDD.n354 GND 0.001706f
C5746 VDD.n355 GND 0.001706f
C5747 VDD.n356 GND 0.001706f
C5748 VDD.n357 GND 0.001706f
C5749 VDD.n358 GND 0.001706f
C5750 VDD.n359 GND 0.001706f
C5751 VDD.n360 GND 0.001706f
C5752 VDD.n361 GND 0.001706f
C5753 VDD.n362 GND 0.001706f
C5754 VDD.n363 GND 0.001706f
C5755 VDD.n364 GND 0.001706f
C5756 VDD.n365 GND 0.001706f
C5757 VDD.n366 GND 0.001706f
C5758 VDD.n367 GND 0.001706f
C5759 VDD.n368 GND 0.001706f
C5760 VDD.n369 GND 0.001706f
C5761 VDD.n370 GND 0.001706f
C5762 VDD.n371 GND 0.001706f
C5763 VDD.n372 GND 0.001706f
C5764 VDD.n373 GND 0.001706f
C5765 VDD.n374 GND 0.001706f
C5766 VDD.n375 GND 0.001706f
C5767 VDD.n376 GND 0.001706f
C5768 VDD.n377 GND 0.001706f
C5769 VDD.n378 GND 0.001706f
C5770 VDD.n379 GND 0.001706f
C5771 VDD.n380 GND 0.001706f
C5772 VDD.n381 GND 0.001706f
C5773 VDD.n382 GND 0.003712f
C5774 VDD.n383 GND 0.003714f
C5775 VDD.n384 GND 0.003714f
C5776 VDD.n386 GND 0.001706f
C5777 VDD.n387 GND 0.001706f
C5778 VDD.n388 GND 0.001706f
C5779 VDD.n389 GND 0.001706f
C5780 VDD.n390 GND 0.001706f
C5781 VDD.n392 GND 0.001706f
C5782 VDD.n393 GND 0.001706f
C5783 VDD.n394 GND 0.001706f
C5784 VDD.n395 GND 0.001547f
C5785 VDD.n396 GND 0.001706f
C5786 VDD.n398 GND 0.001706f
C5787 VDD.n399 GND 0.001062f
C5788 VDD.n400 GND 0.001003f
C5789 VDD.n401 GND 0.011119f
C5790 VDD.n402 GND 0.018664f
C5791 VDD.n403 GND 0.001003f
C5792 VDD.n404 GND 0.001149f
C5793 VDD.n405 GND 0.001706f
C5794 VDD.n407 GND 0.001706f
C5795 VDD.n409 GND 0.001706f
C5796 VDD.n410 GND 0.001706f
C5797 VDD.n411 GND 0.001706f
C5798 VDD.n412 GND 0.001706f
C5799 VDD.n413 GND 0.001706f
C5800 VDD.n415 GND 0.001706f
C5801 VDD.n417 GND 0.001706f
C5802 VDD.n418 GND 0.001706f
C5803 VDD.n419 GND 0.003714f
C5804 VDD.n420 GND 0.003712f
C5805 VDD.n421 GND 0.003712f
C5806 VDD.n422 GND 0.188724f
C5807 VDD.n423 GND 0.003712f
C5808 VDD.n424 GND 0.003712f
C5809 VDD.n425 GND 0.001706f
C5810 VDD.n426 GND 0.001706f
C5811 VDD.n427 GND 0.001706f
C5812 VDD.n428 GND 0.074839f
C5813 VDD.n429 GND 0.001706f
C5814 VDD.n430 GND 0.001706f
C5815 VDD.n431 GND 0.001706f
C5816 VDD.n432 GND 0.001706f
C5817 VDD.n433 GND 0.001706f
C5818 VDD.n434 GND 0.147508f
C5819 VDD.n435 GND 0.001706f
C5820 VDD.n436 GND 0.001706f
C5821 VDD.n437 GND 0.001706f
C5822 VDD.n438 GND 0.001706f
C5823 VDD.n439 GND 0.001706f
C5824 VDD.n440 GND 0.087854f
C5825 VDD.n441 GND 0.001706f
C5826 VDD.n442 GND 0.001706f
C5827 VDD.n443 GND 0.001706f
C5828 VDD.n444 GND 0.001706f
C5829 VDD.n445 GND 0.001706f
C5830 VDD.n446 GND 0.147508f
C5831 VDD.n447 GND 0.001706f
C5832 VDD.n448 GND 0.001706f
C5833 VDD.n449 GND 0.001706f
C5834 VDD.n450 GND 0.001706f
C5835 VDD.n451 GND 0.001706f
C5836 VDD.n452 GND 0.103039f
C5837 VDD.n453 GND 0.001706f
C5838 VDD.n454 GND 0.001706f
C5839 VDD.n455 GND 0.001706f
C5840 VDD.n456 GND 0.001706f
C5841 VDD.n457 GND 0.001706f
C5842 VDD.n458 GND 0.147508f
C5843 VDD.n459 GND 0.001706f
C5844 VDD.n460 GND 0.001706f
C5845 VDD.n461 GND 0.001706f
C5846 VDD.n462 GND 0.001706f
C5847 VDD.n463 GND 0.001706f
C5848 VDD.n464 GND 0.118224f
C5849 VDD.n465 GND 0.001706f
C5850 VDD.n466 GND 0.001706f
C5851 VDD.n467 GND 0.001706f
C5852 VDD.n468 GND 0.001706f
C5853 VDD.n469 GND 0.001706f
C5854 VDD.n470 GND 0.147508f
C5855 VDD.n471 GND 0.001706f
C5856 VDD.n472 GND 0.001706f
C5857 VDD.n473 GND 0.001706f
C5858 VDD.n474 GND 0.001706f
C5859 VDD.n475 GND 0.001706f
C5860 VDD.n476 GND 0.133408f
C5861 VDD.n477 GND 0.001706f
C5862 VDD.n478 GND 0.001706f
C5863 VDD.n479 GND 0.001706f
C5864 VDD.n480 GND 0.001706f
C5865 VDD.n481 GND 0.001706f
C5866 VDD.n482 GND 0.146424f
C5867 VDD.n483 GND 0.001706f
C5868 VDD.n484 GND 0.001706f
C5869 VDD.n485 GND 0.001706f
C5870 VDD.n486 GND 0.001706f
C5871 VDD.n487 GND 0.001706f
C5872 VDD.n488 GND 0.147508f
C5873 VDD.n489 GND 0.001706f
C5874 VDD.n490 GND 0.001706f
C5875 VDD.n491 GND 0.003712f
C5876 VDD.n492 GND 0.003714f
C5877 VDD.n493 GND 0.003714f
C5878 VDD.n495 GND 0.001706f
C5879 VDD.n496 GND 0.001706f
C5880 VDD.n497 GND 0.001706f
C5881 VDD.n498 GND 0.001706f
C5882 VDD.n499 GND 0.001706f
C5883 VDD.n500 GND 0.001706f
C5884 VDD.n502 GND 0.001706f
C5885 VDD.n503 GND 0.001706f
C5886 VDD.n504 GND 0.001547f
C5887 VDD.n505 GND 0.00102f
C5888 VDD.n506 GND 0.017479f
C5889 VDD.n507 GND 3.28559f
C5890 VDD.n508 GND 21.755f
C5891 VDD.n509 GND 0.007272f
C5892 VDD.n510 GND 0.007272f
C5893 VDD.n511 GND 0.002244f
C5894 VDD.t160 GND 0.010699f
C5895 VDD.t96 GND 0.010699f
C5896 VDD.n512 GND 0.022031f
C5897 VDD.n513 GND 9.03e-19
C5898 VDD.n514 GND 0.001516f
C5899 VDD.n515 GND 8.53e-19
C5900 VDD.n516 GND 0.002454f
C5901 VDD.n517 GND 0.002363f
C5902 VDD.n518 GND 8.53e-19
C5903 VDD.n519 GND 9.03e-19
C5904 VDD.n520 GND 0.001972f
C5905 VDD.n521 GND 0.001783f
C5906 VDD.n522 GND 0.044032f
C5907 VDD.n523 GND 0.05786f
C5908 VDD.n524 GND 0.072213f
C5909 VDD.n525 GND 0.007272f
C5910 VDD.n526 GND 0.007272f
C5911 VDD.n527 GND 0.002244f
C5912 VDD.n528 GND 0.002384f
C5913 VDD.n529 GND 9.03e-19
C5914 VDD.n530 GND 8.53e-19
C5915 VDD.n531 GND 0.005733f
C5916 VDD.n532 GND 9.03e-19
C5917 VDD.n533 GND 0.00263f
C5918 VDD.n534 GND 8.53e-19
C5919 VDD.n535 GND 0.002454f
C5920 VDD.n536 GND 0.002363f
C5921 VDD.n537 GND 8.53e-19
C5922 VDD.n538 GND 8.53e-19
C5923 VDD.n539 GND 9.03e-19
C5924 VDD.n540 GND 0.00291f
C5925 VDD.n541 GND 0.00291f
C5926 VDD.n542 GND 0.002183f
C5927 VDD.n543 GND 0.001115f
C5928 VDD.t229 GND 0.00545f
C5929 VDD.n544 GND 0.007088f
C5930 VDD.n545 GND 0.041407f
C5931 VDD.n546 GND 8.53e-19
C5932 VDD.n547 GND 9.03e-19
C5933 VDD.n548 GND 0.00291f
C5934 VDD.n549 GND 0.00291f
C5935 VDD.n550 GND 9.03e-19
C5936 VDD.n551 GND 8.53e-19
C5937 VDD.n552 GND 0.002437f
C5938 VDD.n553 GND 0.004543f
C5939 VDD.n554 GND 0.047272f
C5940 VDD.n555 GND 0.002244f
C5941 VDD.t378 GND 0.010699f
C5942 VDD.t17 GND 0.010699f
C5943 VDD.n556 GND 0.022031f
C5944 VDD.n557 GND 9.03e-19
C5945 VDD.n558 GND 0.001516f
C5946 VDD.n559 GND 8.53e-19
C5947 VDD.n560 GND 0.002454f
C5948 VDD.n561 GND 0.002363f
C5949 VDD.n562 GND 8.53e-19
C5950 VDD.n563 GND 9.03e-19
C5951 VDD.n564 GND 0.001972f
C5952 VDD.n565 GND 0.001783f
C5953 VDD.n566 GND 0.044032f
C5954 VDD.n567 GND 0.05786f
C5955 VDD.n568 GND 0.069098f
C5956 VDD.n569 GND 0.043713f
C5957 VDD.n570 GND 0.001512f
C5958 VDD.n571 GND 0.002407f
C5959 VDD.n572 GND 8.53e-19
C5960 VDD.t51 GND 0.010699f
C5961 VDD.n573 GND 0.001985f
C5962 VDD.n574 GND 0.002355f
C5963 VDD.n575 GND 0.001972f
C5964 VDD.n576 GND 9.03e-19
C5965 VDD.t84 GND 0.010699f
C5966 VDD.n577 GND 0.022036f
C5967 VDD.n578 GND 9.03e-19
C5968 VDD.n579 GND 8.53e-19
C5969 VDD.n580 GND 0.002417f
C5970 VDD.n581 GND 0.007268f
C5971 VDD.n582 GND 0.065607f
C5972 VDD.n583 GND 0.06968f
C5973 VDD.n584 GND 0.043713f
C5974 VDD.n585 GND 0.004453f
C5975 VDD.n586 GND 0.002626f
C5976 VDD.n587 GND 0.002407f
C5977 VDD.n588 GND 8.53e-19
C5978 VDD.n589 GND 0.00291f
C5979 VDD.n590 GND 9.03e-19
C5980 VDD.n591 GND 0.041407f
C5981 VDD.n592 GND 8.53e-19
C5982 VDD.n593 GND 0.00291f
C5983 VDD.t308 GND 0.00545f
C5984 VDD.n594 GND 0.007088f
C5985 VDD.n595 GND 0.001115f
C5986 VDD.n596 GND 0.002183f
C5987 VDD.n597 GND 0.00291f
C5988 VDD.n598 GND 9.03e-19
C5989 VDD.n599 GND 8.53e-19
C5990 VDD.n600 GND 0.002444f
C5991 VDD.n601 GND 0.002355f
C5992 VDD.n602 GND 8.53e-19
C5993 VDD.n603 GND 9.03e-19
C5994 VDD.n604 GND 0.002355f
C5995 VDD.n605 GND 8.53e-19
C5996 VDD.n606 GND 9.03e-19
C5997 VDD.n607 GND 0.00291f
C5998 VDD.n608 GND 0.005733f
C5999 VDD.n609 GND 9.03e-19
C6000 VDD.n610 GND 8.53e-19
C6001 VDD.n611 GND 0.002417f
C6002 VDD.n612 GND 0.007268f
C6003 VDD.n613 GND 0.047272f
C6004 VDD.n614 GND 0.001512f
C6005 VDD.n615 GND 0.002407f
C6006 VDD.n616 GND 8.53e-19
C6007 VDD.t147 GND 0.010699f
C6008 VDD.n617 GND 0.001985f
C6009 VDD.n618 GND 0.002355f
C6010 VDD.n619 GND 0.001972f
C6011 VDD.n620 GND 9.03e-19
C6012 VDD.t110 GND 0.010699f
C6013 VDD.n621 GND 0.022036f
C6014 VDD.n622 GND 9.03e-19
C6015 VDD.n623 GND 8.53e-19
C6016 VDD.n624 GND 0.002417f
C6017 VDD.n625 GND 0.007268f
C6018 VDD.n626 GND 0.05786f
C6019 VDD.n627 GND 0.068374f
C6020 VDD.n628 GND 0.043713f
C6021 VDD.n629 GND 0.001512f
C6022 VDD.n630 GND 0.002407f
C6023 VDD.n631 GND 8.53e-19
C6024 VDD.t100 GND 0.010699f
C6025 VDD.n632 GND 0.001985f
C6026 VDD.n633 GND 0.002355f
C6027 VDD.n634 GND 0.001972f
C6028 VDD.n635 GND 9.03e-19
C6029 VDD.t101 GND 0.010699f
C6030 VDD.n636 GND 0.022036f
C6031 VDD.n637 GND 9.03e-19
C6032 VDD.n638 GND 8.53e-19
C6033 VDD.n639 GND 0.002417f
C6034 VDD.n640 GND 0.007268f
C6035 VDD.n641 GND 0.05786f
C6036 VDD.n642 GND 0.043713f
C6037 VDD.n643 GND 0.001512f
C6038 VDD.n644 GND 0.002407f
C6039 VDD.n645 GND 8.53e-19
C6040 VDD.t513 GND 0.010699f
C6041 VDD.n646 GND 0.001985f
C6042 VDD.n647 GND 0.002355f
C6043 VDD.n648 GND 0.001972f
C6044 VDD.n649 GND 9.03e-19
C6045 VDD.t359 GND 0.010699f
C6046 VDD.n650 GND 0.022036f
C6047 VDD.n651 GND 9.03e-19
C6048 VDD.n652 GND 8.53e-19
C6049 VDD.n653 GND 0.002417f
C6050 VDD.n654 GND 0.007268f
C6051 VDD.n655 GND 0.075015f
C6052 VDD.n656 GND 0.043713f
C6053 VDD.n657 GND 0.001512f
C6054 VDD.n658 GND 0.002407f
C6055 VDD.n659 GND 8.53e-19
C6056 VDD.t286 GND 0.010699f
C6057 VDD.n660 GND 0.001985f
C6058 VDD.n661 GND 0.002355f
C6059 VDD.n662 GND 0.001972f
C6060 VDD.n663 GND 9.03e-19
C6061 VDD.t109 GND 0.010699f
C6062 VDD.n664 GND 0.022036f
C6063 VDD.n665 GND 9.03e-19
C6064 VDD.n666 GND 8.53e-19
C6065 VDD.n667 GND 0.002417f
C6066 VDD.n668 GND 0.007268f
C6067 VDD.n669 GND 0.075015f
C6068 VDD.n670 GND 0.043713f
C6069 VDD.n671 GND 0.001512f
C6070 VDD.n672 GND 0.002407f
C6071 VDD.n673 GND 8.53e-19
C6072 VDD.t82 GND 0.010699f
C6073 VDD.n674 GND 0.001985f
C6074 VDD.n675 GND 0.002355f
C6075 VDD.n676 GND 0.001972f
C6076 VDD.n677 GND 9.03e-19
C6077 VDD.t194 GND 0.010699f
C6078 VDD.n678 GND 0.022036f
C6079 VDD.n679 GND 9.03e-19
C6080 VDD.n680 GND 8.53e-19
C6081 VDD.n681 GND 0.002417f
C6082 VDD.n682 GND 0.007268f
C6083 VDD.n683 GND 0.05786f
C6084 VDD.n684 GND 0.043713f
C6085 VDD.n685 GND 0.043713f
C6086 VDD.n686 GND 0.043713f
C6087 VDD.n687 GND 0.043713f
C6088 VDD.n688 GND 0.001512f
C6089 VDD.n689 GND 0.002407f
C6090 VDD.n690 GND 8.53e-19
C6091 VDD.t309 GND 0.010699f
C6092 VDD.n691 GND 0.001985f
C6093 VDD.n692 GND 0.002355f
C6094 VDD.n693 GND 0.001972f
C6095 VDD.n694 GND 9.03e-19
C6096 VDD.t361 GND 0.010699f
C6097 VDD.n695 GND 0.022036f
C6098 VDD.n696 GND 9.03e-19
C6099 VDD.n697 GND 8.53e-19
C6100 VDD.n698 GND 0.002417f
C6101 VDD.n699 GND 0.007268f
C6102 VDD.n700 GND 0.05786f
C6103 VDD.n701 GND 0.001512f
C6104 VDD.n702 GND 0.002407f
C6105 VDD.n703 GND 8.53e-19
C6106 VDD.t197 GND 0.010699f
C6107 VDD.n704 GND 0.001985f
C6108 VDD.n705 GND 0.002355f
C6109 VDD.n706 GND 0.001972f
C6110 VDD.n707 GND 9.03e-19
C6111 VDD.t196 GND 0.010699f
C6112 VDD.n708 GND 0.022036f
C6113 VDD.n709 GND 9.03e-19
C6114 VDD.n710 GND 8.53e-19
C6115 VDD.n711 GND 0.002417f
C6116 VDD.n712 GND 0.007268f
C6117 VDD.n713 GND 0.076121f
C6118 VDD.n714 GND 0.001512f
C6119 VDD.n715 GND 0.002407f
C6120 VDD.n716 GND 8.53e-19
C6121 VDD.t53 GND 0.010699f
C6122 VDD.n717 GND 0.001985f
C6123 VDD.n718 GND 0.002355f
C6124 VDD.n719 GND 0.001972f
C6125 VDD.n720 GND 9.03e-19
C6126 VDD.t512 GND 0.010699f
C6127 VDD.n721 GND 0.022036f
C6128 VDD.n722 GND 9.03e-19
C6129 VDD.n723 GND 8.53e-19
C6130 VDD.n724 GND 0.002417f
C6131 VDD.n725 GND 0.007268f
C6132 VDD.n726 GND 0.075015f
C6133 VDD.n727 GND 0.001512f
C6134 VDD.n728 GND 0.002407f
C6135 VDD.n729 GND 8.53e-19
C6136 VDD.t285 GND 0.010699f
C6137 VDD.n730 GND 0.001985f
C6138 VDD.n731 GND 0.002355f
C6139 VDD.n732 GND 0.001972f
C6140 VDD.n733 GND 9.03e-19
C6141 VDD.t149 GND 0.010699f
C6142 VDD.n734 GND 0.022036f
C6143 VDD.n735 GND 9.03e-19
C6144 VDD.n736 GND 8.53e-19
C6145 VDD.n737 GND 0.002417f
C6146 VDD.n738 GND 0.007268f
C6147 VDD.n739 GND 0.05786f
C6148 VDD.n740 GND 0.060777f
C6149 VDD.n741 GND 1.36913f
C6150 VDD.n742 GND 0.007272f
C6151 VDD.n743 GND 0.002244f
C6152 VDD.t88 GND 0.010699f
C6153 VDD.t335 GND 0.010699f
C6154 VDD.n744 GND 0.022031f
C6155 VDD.n745 GND 9.03e-19
C6156 VDD.n746 GND 0.001516f
C6157 VDD.n747 GND 8.53e-19
C6158 VDD.n748 GND 0.002454f
C6159 VDD.n749 GND 0.002363f
C6160 VDD.n750 GND 8.53e-19
C6161 VDD.n751 GND 9.03e-19
C6162 VDD.n752 GND 0.001972f
C6163 VDD.n753 GND 0.001783f
C6164 VDD.n754 GND 0.044032f
C6165 VDD.n755 GND 0.076121f
C6166 VDD.n756 GND 0.007272f
C6167 VDD.n757 GND 0.002244f
C6168 VDD.t92 GND 0.010699f
C6169 VDD.t94 GND 0.010699f
C6170 VDD.n758 GND 0.022031f
C6171 VDD.n759 GND 9.03e-19
C6172 VDD.n760 GND 0.001516f
C6173 VDD.n761 GND 8.53e-19
C6174 VDD.n762 GND 0.002454f
C6175 VDD.n763 GND 0.002363f
C6176 VDD.n764 GND 8.53e-19
C6177 VDD.n765 GND 9.03e-19
C6178 VDD.n766 GND 0.001972f
C6179 VDD.n767 GND 0.001783f
C6180 VDD.n768 GND 0.044032f
C6181 VDD.n769 GND 0.075015f
C6182 VDD.n770 GND 0.007272f
C6183 VDD.n771 GND 0.002244f
C6184 VDD.t178 GND 0.010699f
C6185 VDD.t227 GND 0.010699f
C6186 VDD.n772 GND 0.022031f
C6187 VDD.n773 GND 9.03e-19
C6188 VDD.n774 GND 0.001516f
C6189 VDD.n775 GND 8.53e-19
C6190 VDD.n776 GND 0.002454f
C6191 VDD.n777 GND 0.002363f
C6192 VDD.n778 GND 8.53e-19
C6193 VDD.n779 GND 9.03e-19
C6194 VDD.n780 GND 0.001972f
C6195 VDD.n781 GND 0.001783f
C6196 VDD.n782 GND 0.044032f
C6197 VDD.n783 GND 0.056753f
C6198 VDD.n784 GND 0.007272f
C6199 VDD.n785 GND 0.007272f
C6200 VDD.n786 GND 0.007272f
C6201 VDD.n787 GND 0.007272f
C6202 VDD.n788 GND 0.002244f
C6203 VDD.t112 GND 0.010699f
C6204 VDD.t519 GND 0.010699f
C6205 VDD.n789 GND 0.022031f
C6206 VDD.n790 GND 9.03e-19
C6207 VDD.n791 GND 0.001516f
C6208 VDD.n792 GND 8.53e-19
C6209 VDD.n793 GND 0.002454f
C6210 VDD.n794 GND 0.002363f
C6211 VDD.n795 GND 8.53e-19
C6212 VDD.n796 GND 9.03e-19
C6213 VDD.n797 GND 0.001972f
C6214 VDD.n798 GND 0.001783f
C6215 VDD.n799 GND 0.044032f
C6216 VDD.n800 GND 0.05786f
C6217 VDD.n801 GND 0.002244f
C6218 VDD.t90 GND 0.010699f
C6219 VDD.t466 GND 0.010699f
C6220 VDD.n802 GND 0.022031f
C6221 VDD.n803 GND 9.03e-19
C6222 VDD.n804 GND 0.001516f
C6223 VDD.n805 GND 8.53e-19
C6224 VDD.n806 GND 0.002454f
C6225 VDD.n807 GND 0.002363f
C6226 VDD.n808 GND 8.53e-19
C6227 VDD.n809 GND 9.03e-19
C6228 VDD.n810 GND 0.001972f
C6229 VDD.n811 GND 0.001783f
C6230 VDD.n812 GND 0.044032f
C6231 VDD.n813 GND 0.076121f
C6232 VDD.n814 GND 0.002244f
C6233 VDD.t332 GND 0.010699f
C6234 VDD.t465 GND 0.010699f
C6235 VDD.n815 GND 0.022031f
C6236 VDD.n816 GND 9.03e-19
C6237 VDD.n817 GND 0.001516f
C6238 VDD.n818 GND 8.53e-19
C6239 VDD.n819 GND 0.002454f
C6240 VDD.n820 GND 0.002363f
C6241 VDD.n821 GND 8.53e-19
C6242 VDD.n822 GND 9.03e-19
C6243 VDD.n823 GND 0.001972f
C6244 VDD.n824 GND 0.001783f
C6245 VDD.n825 GND 0.044032f
C6246 VDD.n826 GND 0.075015f
C6247 VDD.n827 GND 0.002244f
C6248 VDD.t267 GND 0.010699f
C6249 VDD.t259 GND 0.010699f
C6250 VDD.n828 GND 0.022031f
C6251 VDD.n829 GND 9.03e-19
C6252 VDD.n830 GND 0.001516f
C6253 VDD.n831 GND 8.53e-19
C6254 VDD.n832 GND 0.002454f
C6255 VDD.n833 GND 0.002363f
C6256 VDD.n834 GND 8.53e-19
C6257 VDD.n835 GND 9.03e-19
C6258 VDD.n836 GND 0.001972f
C6259 VDD.n837 GND 0.001783f
C6260 VDD.n838 GND 0.044032f
C6261 VDD.n839 GND 0.05786f
C6262 VDD.n840 GND 0.062709f
C6263 VDD.n841 GND 0.00991f
C6264 VDD.n842 GND 0.001706f
C6265 VDD.n843 GND 0.012142f
C6266 VDD.n844 GND 0.001706f
C6267 VDD.n845 GND 0.001706f
C6268 VDD.n846 GND 0.119161f
C6269 VDD.n847 GND 0.001706f
C6270 VDD.t701 GND 0.117408f
C6271 VDD.n848 GND 0.001706f
C6272 VDD.n849 GND 0.001706f
C6273 VDD.n850 GND 8.53e-19
C6274 VDD.n851 GND 9.03e-19
C6275 VDD.n852 GND 0.010359f
C6276 VDD.n853 GND 0.010359f
C6277 VDD.n854 GND 9.03e-19
C6278 VDD.n855 GND 8.78e-19
C6279 VDD.n856 GND 0.001706f
C6280 VDD.n857 GND 0.001706f
C6281 VDD.n858 GND 0.026285f
C6282 VDD.n859 GND 0.001706f
C6283 VDD.n860 GND 0.001706f
C6284 VDD.n861 GND 8.53e-19
C6285 VDD.n862 GND 9.03e-19
C6286 VDD.n863 GND 0.021453f
C6287 VDD.n864 GND 0.013609f
C6288 VDD.n865 GND 0.508412f
C6289 VDD.n866 GND 0.004436f
C6290 VDD.n867 GND 0.002626f
C6291 VDD.n868 GND 0.002407f
C6292 VDD.n869 GND 8.53e-19
C6293 VDD.n870 GND 0.00291f
C6294 VDD.n871 GND 9.03e-19
C6295 VDD.n872 GND 0.041407f
C6296 VDD.n873 GND 8.53e-19
C6297 VDD.n874 GND 0.00291f
C6298 VDD.t80 GND 0.00545f
C6299 VDD.n875 GND 0.007088f
C6300 VDD.n876 GND 0.001115f
C6301 VDD.n877 GND 0.002183f
C6302 VDD.n878 GND 0.00291f
C6303 VDD.n879 GND 9.03e-19
C6304 VDD.n880 GND 8.53e-19
C6305 VDD.n881 GND 0.002385f
C6306 VDD.n882 GND 0.002421f
C6307 VDD.n883 GND 8.53e-19
C6308 VDD.n884 GND 9.03e-19
C6309 VDD.n885 GND 0.002366f
C6310 VDD.n886 GND 8.53e-19
C6311 VDD.n887 GND 9.03e-19
C6312 VDD.n888 GND 0.00291f
C6313 VDD.n889 GND 0.005733f
C6314 VDD.n890 GND 9.03e-19
C6315 VDD.n891 GND 8.53e-19
C6316 VDD.n892 GND 0.002417f
C6317 VDD.n893 GND 0.007268f
C6318 VDD.n894 GND 0.050371f
C6319 VDD.n895 GND 0.044305f
C6320 VDD.n896 GND 0.001512f
C6321 VDD.n897 GND 0.002407f
C6322 VDD.n898 GND 8.53e-19
C6323 VDD.t296 GND 0.010699f
C6324 VDD.n899 GND 0.001399f
C6325 VDD.n900 GND 0.002366f
C6326 VDD.n901 GND 0.001972f
C6327 VDD.n902 GND 9.03e-19
C6328 VDD.t7 GND 0.010699f
C6329 VDD.n903 GND 0.02202f
C6330 VDD.n904 GND 9.03e-19
C6331 VDD.n905 GND 8.53e-19
C6332 VDD.n906 GND 0.002417f
C6333 VDD.n907 GND 0.007268f
C6334 VDD.n908 GND 0.062508f
C6335 VDD.n909 GND 0.115599f
C6336 VDD.n910 GND 0.044305f
C6337 VDD.n911 GND 0.001512f
C6338 VDD.n912 GND 0.002407f
C6339 VDD.n913 GND 8.53e-19
C6340 VDD.t175 GND 0.010699f
C6341 VDD.n914 GND 0.001399f
C6342 VDD.n915 GND 0.002366f
C6343 VDD.n916 GND 0.001972f
C6344 VDD.n917 GND 9.03e-19
C6345 VDD.t78 GND 0.010699f
C6346 VDD.n918 GND 0.02202f
C6347 VDD.n919 GND 9.03e-19
C6348 VDD.n920 GND 8.53e-19
C6349 VDD.n921 GND 0.002417f
C6350 VDD.n922 GND 0.007268f
C6351 VDD.n923 GND 0.063726f
C6352 VDD.n924 GND 0.044305f
C6353 VDD.n925 GND 0.001512f
C6354 VDD.n926 GND 0.002407f
C6355 VDD.n927 GND 8.53e-19
C6356 VDD.t5 GND 0.010699f
C6357 VDD.n928 GND 0.001399f
C6358 VDD.n929 GND 0.002366f
C6359 VDD.n930 GND 0.001972f
C6360 VDD.n931 GND 9.03e-19
C6361 VDD.t98 GND 0.010699f
C6362 VDD.n932 GND 0.02202f
C6363 VDD.n933 GND 9.03e-19
C6364 VDD.n934 GND 8.53e-19
C6365 VDD.n935 GND 0.002417f
C6366 VDD.n936 GND 0.007268f
C6367 VDD.n937 GND 0.081987f
C6368 VDD.n938 GND 0.044305f
C6369 VDD.n939 GND 0.001512f
C6370 VDD.n940 GND 0.002407f
C6371 VDD.n941 GND 8.53e-19
C6372 VDD.t543 GND 0.010699f
C6373 VDD.n942 GND 0.001399f
C6374 VDD.n943 GND 0.002366f
C6375 VDD.n944 GND 0.001972f
C6376 VDD.n945 GND 9.03e-19
C6377 VDD.t349 GND 0.010699f
C6378 VDD.n946 GND 0.02202f
C6379 VDD.n947 GND 9.03e-19
C6380 VDD.n948 GND 8.53e-19
C6381 VDD.n949 GND 0.002417f
C6382 VDD.n950 GND 0.007268f
C6383 VDD.n951 GND 0.081987f
C6384 VDD.n952 GND 0.044305f
C6385 VDD.n953 GND 0.001512f
C6386 VDD.n954 GND 0.002407f
C6387 VDD.n955 GND 8.53e-19
C6388 VDD.t453 GND 0.010699f
C6389 VDD.n956 GND 0.001399f
C6390 VDD.n957 GND 0.002366f
C6391 VDD.n958 GND 0.001972f
C6392 VDD.n959 GND 9.03e-19
C6393 VDD.t471 GND 0.010699f
C6394 VDD.n960 GND 0.02202f
C6395 VDD.n961 GND 9.03e-19
C6396 VDD.n962 GND 8.53e-19
C6397 VDD.n963 GND 0.002417f
C6398 VDD.n964 GND 0.007268f
C6399 VDD.n965 GND 0.081987f
C6400 VDD.n966 GND 0.044305f
C6401 VDD.n967 GND 0.001512f
C6402 VDD.n968 GND 0.002407f
C6403 VDD.n969 GND 8.53e-19
C6404 VDD.t469 GND 0.010699f
C6405 VDD.n970 GND 0.001399f
C6406 VDD.n971 GND 0.002366f
C6407 VDD.n972 GND 0.001972f
C6408 VDD.n973 GND 9.03e-19
C6409 VDD.t499 GND 0.010699f
C6410 VDD.n974 GND 0.02202f
C6411 VDD.n975 GND 9.03e-19
C6412 VDD.n976 GND 8.53e-19
C6413 VDD.n977 GND 0.002417f
C6414 VDD.n978 GND 0.007268f
C6415 VDD.n979 GND 0.081987f
C6416 VDD.n980 GND 0.044305f
C6417 VDD.n981 GND 0.001512f
C6418 VDD.n982 GND 0.002407f
C6419 VDD.n983 GND 8.53e-19
C6420 VDD.t243 GND 0.010699f
C6421 VDD.n984 GND 0.001399f
C6422 VDD.n985 GND 0.002366f
C6423 VDD.n986 GND 0.001972f
C6424 VDD.n987 GND 9.03e-19
C6425 VDD.t535 GND 0.010699f
C6426 VDD.n988 GND 0.02202f
C6427 VDD.n989 GND 9.03e-19
C6428 VDD.n990 GND 8.53e-19
C6429 VDD.n991 GND 0.002417f
C6430 VDD.n992 GND 0.007268f
C6431 VDD.n993 GND 0.063726f
C6432 VDD.n994 GND 0.044305f
C6433 VDD.n995 GND 0.044305f
C6434 VDD.n996 GND 0.044305f
C6435 VDD.n997 GND 0.044305f
C6436 VDD.n998 GND 0.044305f
C6437 VDD.n999 GND 0.044305f
C6438 VDD.n1000 GND 0.044305f
C6439 VDD.n1001 GND 0.044305f
C6440 VDD.n1002 GND 0.044305f
C6441 VDD.n1003 GND 0.044305f
C6442 VDD.n1004 GND 0.044305f
C6443 VDD.n1005 GND 0.044305f
C6444 VDD.n1006 GND 0.004436f
C6445 VDD.n1007 GND 0.002626f
C6446 VDD.n1008 GND 0.002407f
C6447 VDD.n1009 GND 8.53e-19
C6448 VDD.n1010 GND 0.00291f
C6449 VDD.n1011 GND 9.03e-19
C6450 VDD.n1012 GND 0.041407f
C6451 VDD.n1013 GND 8.53e-19
C6452 VDD.n1014 GND 0.00291f
C6453 VDD.t517 GND 0.00545f
C6454 VDD.n1015 GND 0.007088f
C6455 VDD.n1016 GND 0.001115f
C6456 VDD.n1017 GND 0.002183f
C6457 VDD.n1018 GND 0.00291f
C6458 VDD.n1019 GND 9.03e-19
C6459 VDD.n1020 GND 8.53e-19
C6460 VDD.n1021 GND 0.002385f
C6461 VDD.n1022 GND 0.002421f
C6462 VDD.n1023 GND 8.53e-19
C6463 VDD.n1024 GND 9.03e-19
C6464 VDD.n1025 GND 0.002366f
C6465 VDD.n1026 GND 8.53e-19
C6466 VDD.n1027 GND 9.03e-19
C6467 VDD.n1028 GND 0.00291f
C6468 VDD.n1029 GND 0.005733f
C6469 VDD.n1030 GND 9.03e-19
C6470 VDD.n1031 GND 8.53e-19
C6471 VDD.n1032 GND 0.002417f
C6472 VDD.n1033 GND 0.007268f
C6473 VDD.n1034 GND 0.051588f
C6474 VDD.n1035 GND 0.001512f
C6475 VDD.n1036 GND 0.002407f
C6476 VDD.n1037 GND 8.53e-19
C6477 VDD.t37 GND 0.010699f
C6478 VDD.n1038 GND 0.001399f
C6479 VDD.n1039 GND 0.002366f
C6480 VDD.n1040 GND 0.001972f
C6481 VDD.n1041 GND 9.03e-19
C6482 VDD.t127 GND 0.010699f
C6483 VDD.n1042 GND 0.02202f
C6484 VDD.n1043 GND 9.03e-19
C6485 VDD.n1044 GND 8.53e-19
C6486 VDD.n1045 GND 0.002417f
C6487 VDD.n1046 GND 0.007268f
C6488 VDD.n1047 GND 0.062508f
C6489 VDD.n1048 GND 0.113942f
C6490 VDD.n1049 GND 0.001512f
C6491 VDD.n1050 GND 0.002407f
C6492 VDD.n1051 GND 8.53e-19
C6493 VDD.t539 GND 0.010699f
C6494 VDD.n1052 GND 0.001399f
C6495 VDD.n1053 GND 0.002366f
C6496 VDD.n1054 GND 0.001972f
C6497 VDD.n1055 GND 9.03e-19
C6498 VDD.t222 GND 0.010699f
C6499 VDD.n1056 GND 0.02202f
C6500 VDD.n1057 GND 9.03e-19
C6501 VDD.n1058 GND 8.53e-19
C6502 VDD.n1059 GND 0.002417f
C6503 VDD.n1060 GND 0.007268f
C6504 VDD.n1061 GND 0.063726f
C6505 VDD.n1062 GND 0.001512f
C6506 VDD.n1063 GND 0.002407f
C6507 VDD.n1064 GND 8.53e-19
C6508 VDD.t502 GND 0.010699f
C6509 VDD.n1065 GND 0.001399f
C6510 VDD.n1066 GND 0.002366f
C6511 VDD.n1067 GND 0.001972f
C6512 VDD.n1068 GND 9.03e-19
C6513 VDD.t358 GND 0.010699f
C6514 VDD.n1069 GND 0.02202f
C6515 VDD.n1070 GND 9.03e-19
C6516 VDD.n1071 GND 8.53e-19
C6517 VDD.n1072 GND 0.002417f
C6518 VDD.n1073 GND 0.007268f
C6519 VDD.n1074 GND 0.081987f
C6520 VDD.n1075 GND 0.001512f
C6521 VDD.n1076 GND 0.002407f
C6522 VDD.n1077 GND 8.53e-19
C6523 VDD.t337 GND 0.010699f
C6524 VDD.n1078 GND 0.001399f
C6525 VDD.n1079 GND 0.002366f
C6526 VDD.n1080 GND 0.001972f
C6527 VDD.n1081 GND 9.03e-19
C6528 VDD.t249 GND 0.010699f
C6529 VDD.n1082 GND 0.02202f
C6530 VDD.n1083 GND 9.03e-19
C6531 VDD.n1084 GND 8.53e-19
C6532 VDD.n1085 GND 0.002417f
C6533 VDD.n1086 GND 0.007268f
C6534 VDD.n1087 GND 0.081987f
C6535 VDD.n1088 GND 0.001512f
C6536 VDD.n1089 GND 0.002407f
C6537 VDD.n1090 GND 8.53e-19
C6538 VDD.t272 GND 0.010699f
C6539 VDD.n1091 GND 0.001399f
C6540 VDD.n1092 GND 0.002366f
C6541 VDD.n1093 GND 0.001972f
C6542 VDD.n1094 GND 9.03e-19
C6543 VDD.t190 GND 0.010699f
C6544 VDD.n1095 GND 0.02202f
C6545 VDD.n1096 GND 9.03e-19
C6546 VDD.n1097 GND 8.53e-19
C6547 VDD.n1098 GND 0.002417f
C6548 VDD.n1099 GND 0.007268f
C6549 VDD.n1100 GND 0.083204f
C6550 VDD.n1101 GND 0.001512f
C6551 VDD.n1102 GND 0.002407f
C6552 VDD.n1103 GND 8.53e-19
C6553 VDD.t455 GND 0.010699f
C6554 VDD.n1104 GND 0.001399f
C6555 VDD.n1105 GND 0.002366f
C6556 VDD.n1106 GND 0.001972f
C6557 VDD.n1107 GND 9.03e-19
C6558 VDD.t347 GND 0.010699f
C6559 VDD.n1108 GND 0.02202f
C6560 VDD.n1109 GND 9.03e-19
C6561 VDD.n1110 GND 8.53e-19
C6562 VDD.n1111 GND 0.002417f
C6563 VDD.n1112 GND 0.007268f
C6564 VDD.n1113 GND 0.081987f
C6565 VDD.n1114 GND 0.001512f
C6566 VDD.n1115 GND 0.002407f
C6567 VDD.n1116 GND 8.53e-19
C6568 VDD.t247 GND 0.010699f
C6569 VDD.n1117 GND 0.001399f
C6570 VDD.n1118 GND 0.002366f
C6571 VDD.n1119 GND 0.001972f
C6572 VDD.n1120 GND 9.03e-19
C6573 VDD.t251 GND 0.010699f
C6574 VDD.n1121 GND 0.02202f
C6575 VDD.n1122 GND 9.03e-19
C6576 VDD.n1123 GND 8.53e-19
C6577 VDD.n1124 GND 0.002417f
C6578 VDD.n1125 GND 0.007268f
C6579 VDD.n1126 GND 0.062508f
C6580 VDD.n1127 GND 0.06242f
C6581 VDD.n1128 GND 0.001512f
C6582 VDD.n1129 GND 0.002407f
C6583 VDD.n1130 GND 8.53e-19
C6584 VDD.t35 GND 0.010699f
C6585 VDD.n1131 GND 0.001399f
C6586 VDD.n1132 GND 0.002366f
C6587 VDD.n1133 GND 0.001972f
C6588 VDD.n1134 GND 9.03e-19
C6589 VDD.t325 GND 0.010699f
C6590 VDD.n1135 GND 0.02202f
C6591 VDD.n1136 GND 9.03e-19
C6592 VDD.n1137 GND 8.53e-19
C6593 VDD.n1138 GND 0.002417f
C6594 VDD.n1139 GND 0.007268f
C6595 VDD.n1140 GND 0.063726f
C6596 VDD.n1141 GND 0.001512f
C6597 VDD.n1142 GND 0.002407f
C6598 VDD.n1143 GND 8.53e-19
C6599 VDD.t13 GND 0.010699f
C6600 VDD.n1144 GND 0.001399f
C6601 VDD.n1145 GND 0.002366f
C6602 VDD.n1146 GND 0.001972f
C6603 VDD.n1147 GND 9.03e-19
C6604 VDD.t241 GND 0.010699f
C6605 VDD.n1148 GND 0.02202f
C6606 VDD.n1149 GND 9.03e-19
C6607 VDD.n1150 GND 8.53e-19
C6608 VDD.n1151 GND 0.002417f
C6609 VDD.n1152 GND 0.007268f
C6610 VDD.n1153 GND 0.081987f
C6611 VDD.n1154 GND 0.001512f
C6612 VDD.n1155 GND 0.002407f
C6613 VDD.n1156 GND 8.53e-19
C6614 VDD.t385 GND 0.010699f
C6615 VDD.n1157 GND 0.001399f
C6616 VDD.n1158 GND 0.002366f
C6617 VDD.n1159 GND 0.001972f
C6618 VDD.n1160 GND 9.03e-19
C6619 VDD.t293 GND 0.010699f
C6620 VDD.n1161 GND 0.02202f
C6621 VDD.n1162 GND 9.03e-19
C6622 VDD.n1163 GND 8.53e-19
C6623 VDD.n1164 GND 0.002417f
C6624 VDD.n1165 GND 0.007268f
C6625 VDD.n1166 GND 0.081987f
C6626 VDD.n1167 GND 0.001512f
C6627 VDD.n1168 GND 0.002407f
C6628 VDD.n1169 GND 8.53e-19
C6629 VDD.t351 GND 0.010699f
C6630 VDD.n1170 GND 0.001399f
C6631 VDD.n1171 GND 0.002366f
C6632 VDD.n1172 GND 0.001972f
C6633 VDD.n1173 GND 9.03e-19
C6634 VDD.t11 GND 0.010699f
C6635 VDD.n1174 GND 0.02202f
C6636 VDD.n1175 GND 9.03e-19
C6637 VDD.n1176 GND 8.53e-19
C6638 VDD.n1177 GND 0.002417f
C6639 VDD.n1178 GND 0.007268f
C6640 VDD.n1179 GND 0.081987f
C6641 VDD.n1180 GND 0.001512f
C6642 VDD.n1181 GND 0.002407f
C6643 VDD.n1182 GND 8.53e-19
C6644 VDD.t702 GND 0.010699f
C6645 VDD.n1183 GND 0.001399f
C6646 VDD.n1184 GND 0.002366f
C6647 VDD.n1185 GND 0.001972f
C6648 VDD.n1186 GND 9.03e-19
C6649 VDD.t274 GND 0.010699f
C6650 VDD.n1187 GND 0.02202f
C6651 VDD.n1188 GND 9.03e-19
C6652 VDD.n1189 GND 8.53e-19
C6653 VDD.n1190 GND 0.002417f
C6654 VDD.n1191 GND 0.007268f
C6655 VDD.n1192 GND 0.062508f
C6656 VDD.n1193 GND 0.06242f
C6657 VDD.n1194 GND 0.506755f
C6658 VDD.n1195 GND 0.859285f
C6659 VDD.n1196 GND 0.010271f
C6660 VDD.n1197 GND 0.017055f
C6661 VDD.n1198 GND 9.03e-19
C6662 VDD.n1199 GND 8.78e-19
C6663 VDD.n1200 GND 0.001706f
C6664 VDD.n1201 GND 0.001706f
C6665 VDD.t34 GND 0.117408f
C6666 VDD.n1202 GND 0.001706f
C6667 VDD.n1203 GND 0.001706f
C6668 VDD.n1204 GND 0.001706f
C6669 VDD.t89 GND 0.117408f
C6670 VDD.n1205 GND 0.001706f
C6671 VDD.n1206 GND 0.001706f
C6672 VDD.n1207 GND 0.001706f
C6673 VDD.n1208 GND 8.53e-19
C6674 VDD.n1209 GND 9.03e-19
C6675 VDD.n1210 GND 0.010359f
C6676 VDD.n1211 GND 0.010359f
C6677 VDD.n1212 GND 8.78e-19
C6678 VDD.n1213 GND 8.53e-19
C6679 VDD.n1214 GND 0.001706f
C6680 VDD.n1215 GND 0.001706f
C6681 VDD.t324 GND 0.117408f
C6682 VDD.n1216 GND 0.119161f
C6683 VDD.n1217 GND 0.001706f
C6684 VDD.n1218 GND 8.53e-19
C6685 VDD.n1219 GND 9.03e-19
C6686 VDD.n1220 GND 0.002444f
C6687 VDD.n1221 GND 8.53e-19
C6688 VDD.n1222 GND 0.001706f
C6689 VDD.t195 GND 0.117408f
C6690 VDD.n1223 GND 0.001706f
C6691 VDD.n1224 GND 0.001706f
C6692 VDD.n1225 GND 0.001706f
C6693 VDD.t246 GND 0.117408f
C6694 VDD.n1226 GND 0.001706f
C6695 VDD.n1227 GND 0.001706f
C6696 VDD.n1228 GND 0.001706f
C6697 VDD.n1229 GND 8.53e-19
C6698 VDD.n1230 GND 0.001706f
C6699 VDD.n1231 GND 0.001706f
C6700 VDD.n1232 GND 0.06659f
C6701 VDD.n1233 GND 0.001706f
C6702 VDD.n1234 GND 0.001706f
C6703 VDD.t250 GND 0.117408f
C6704 VDD.n1235 GND 0.001706f
C6705 VDD.n1236 GND 0.001706f
C6706 VDD.n1237 GND 0.012142f
C6707 VDD.n1238 GND 0.00133f
C6708 VDD.n1239 GND 0.001706f
C6709 VDD.n1240 GND 0.001706f
C6710 VDD.n1241 GND 0.049066f
C6711 VDD.n1242 GND 0.001706f
C6712 VDD.n1243 GND 0.001706f
C6713 VDD.n1244 GND 0.110399f
C6714 VDD.n1245 GND 0.001706f
C6715 VDD.n1246 GND 0.001706f
C6716 VDD.n1247 GND 8.53e-19
C6717 VDD.n1248 GND 9.03e-19
C6718 VDD.n1249 GND 0.002444f
C6719 VDD.n1250 GND 9.03e-19
C6720 VDD.n1251 GND 8.53e-19
C6721 VDD.n1252 GND 0.001706f
C6722 VDD.n1253 GND 9.03e-19
C6723 VDD.n1254 GND 9.03e-19
C6724 VDD.n1255 GND 8.53e-19
C6725 VDD.n1256 GND 0.002444f
C6726 VDD.n1257 GND 0.002444f
C6727 VDD.n1258 GND 0.002444f
C6728 VDD.n1259 GND 8.53e-19
C6729 VDD.n1260 GND 0.001706f
C6730 VDD.n1261 GND 0.119161f
C6731 VDD.n1262 GND 0.001706f
C6732 VDD.n1263 GND 0.001706f
C6733 VDD.n1264 GND 0.001706f
C6734 VDD.t146 GND 0.117408f
C6735 VDD.n1265 GND 0.001706f
C6736 VDD.n1266 GND 0.001706f
C6737 VDD.n1267 GND 0.001706f
C6738 VDD.n1268 GND 0.001706f
C6739 VDD.n1269 GND 0.001706f
C6740 VDD.n1270 GND 0.001706f
C6741 VDD.n1271 GND 0.001706f
C6742 VDD.n1272 GND 0.001706f
C6743 VDD.n1273 GND 0.091123f
C6744 VDD.n1274 GND 0.001706f
C6745 VDD.n1275 GND 0.001706f
C6746 VDD.t16 GND 0.117408f
C6747 VDD.n1276 GND 0.001706f
C6748 VDD.n1277 GND 0.001706f
C6749 VDD.n1278 GND 0.001706f
C6750 VDD.n1279 GND 0.001706f
C6751 VDD.n1280 GND 0.001706f
C6752 VDD.n1281 GND 0.001706f
C6753 VDD.n1282 GND 0.001706f
C6754 VDD.n1283 GND 0.001706f
C6755 VDD.n1284 GND 0.001706f
C6756 VDD.n1285 GND 0.001706f
C6757 VDD.n1286 GND 0.052571f
C6758 VDD.n1287 GND 0.001706f
C6759 VDD.n1288 GND 0.001706f
C6760 VDD.t228 GND 0.117408f
C6761 VDD.n1289 GND 0.001706f
C6762 VDD.n1290 GND 0.003727f
C6763 VDD.n1291 GND 0.003727f
C6764 VDD.n1292 GND 0.014019f
C6765 VDD.n1293 GND 0.003723f
C6766 VDD.n1294 GND 0.003723f
C6767 VDD.n1295 GND 0.187503f
C6768 VDD.n1296 GND 0.003727f
C6769 VDD.n1297 GND 0.001706f
C6770 VDD.n1298 GND 0.001706f
C6771 VDD.n1313 GND 0.003727f
C6772 VDD.n1314 GND 0.075352f
C6773 VDD.n1315 GND 0.001706f
C6774 VDD.n1316 GND 0.001706f
C6775 VDD.n1317 GND 0.031543f
C6776 VDD.n1318 GND 0.001706f
C6777 VDD.n1319 GND 0.070094f
C6778 VDD.n1320 GND 0.001706f
C6779 VDD.n1321 GND 0.001706f
C6780 VDD.n1322 GND 0.001706f
C6781 VDD.n1323 GND 0.108646f
C6782 VDD.n1324 GND 0.001706f
C6783 VDD.n1325 GND 0.001706f
C6784 VDD.n1326 GND 0.119161f
C6785 VDD.n1327 GND 0.001706f
C6786 VDD.n1328 GND 0.001706f
C6787 VDD.n1329 GND 0.012142f
C6788 VDD.n1330 GND 0.024533f
C6789 VDD.n1331 GND 0.001706f
C6790 VDD.n1332 GND 0.001706f
C6791 VDD.n1333 GND 0.063085f
C6792 VDD.n1334 GND 0.001706f
C6793 VDD.n1335 GND 0.001706f
C6794 VDD.n1336 GND 9.03e-19
C6795 VDD.n1337 GND 0.001706f
C6796 VDD.n1338 GND 0.001706f
C6797 VDD.n1339 GND 0.101637f
C6798 VDD.n1340 GND 0.001706f
C6799 VDD.n1341 GND 0.001706f
C6800 VDD.t240 GND 0.117408f
C6801 VDD.n1342 GND 0.001706f
C6802 VDD.n1343 GND 0.001706f
C6803 VDD.n1344 GND 8.53e-19
C6804 VDD.n1345 GND 9.03e-19
C6805 VDD.n1346 GND 0.010359f
C6806 VDD.n1347 GND 9.03e-19
C6807 VDD.n1348 GND 8.53e-19
C6808 VDD.n1349 GND 0.010359f
C6809 VDD.n1350 GND 9.03e-19
C6810 VDD.n1351 GND 8.53e-19
C6811 VDD.n1352 GND 0.001706f
C6812 VDD.n1353 GND 8.78e-19
C6813 VDD.n1354 GND 8.53e-19
C6814 VDD.n1355 GND 9.03e-19
C6815 VDD.n1356 GND 0.001706f
C6816 VDD.n1357 GND 0.001706f
C6817 VDD.t464 GND 0.117408f
C6818 VDD.n1358 GND 0.057828f
C6819 VDD.n1359 GND 0.001706f
C6820 VDD.n1360 GND 9.03e-19
C6821 VDD.n1361 GND 0.018487f
C6822 VDD.n1362 GND 8.53e-19
C6823 VDD.n1363 GND 0.001706f
C6824 VDD.n1364 GND 0.119161f
C6825 VDD.n1365 GND 0.001706f
C6826 VDD.n1366 GND 0.001706f
C6827 VDD.n1367 GND 0.001706f
C6828 VDD.n1368 GND 0.001706f
C6829 VDD.n1369 GND 0.001706f
C6830 VDD.n1370 GND 0.021028f
C6831 VDD.n1371 GND 0.001706f
C6832 VDD.t12 GND 0.117408f
C6833 VDD.n1372 GND 0.001706f
C6834 VDD.n1373 GND 0.001706f
C6835 VDD.n1374 GND 0.001706f
C6836 VDD.n1375 GND 8.53e-19
C6837 VDD.n1376 GND 9.03e-19
C6838 VDD.n1377 GND 0.010359f
C6839 VDD.n1378 GND 9.03e-19
C6840 VDD.n1379 GND 8.53e-19
C6841 VDD.n1380 GND 0.010359f
C6842 VDD.n1381 GND 9.03e-19
C6843 VDD.n1382 GND 8.53e-19
C6844 VDD.n1383 GND 9.03e-19
C6845 VDD.n1384 GND 0.010359f
C6846 VDD.n1385 GND 0.010359f
C6847 VDD.n1386 GND 8.53e-19
C6848 VDD.n1387 GND 0.001706f
C6849 VDD.n1388 GND 8.53e-19
C6850 VDD.n1389 GND 9.03e-19
C6851 VDD.t292 GND 0.117408f
C6852 VDD.t148 GND 0.117408f
C6853 VDD.n1390 GND 0.099885f
C6854 VDD.n1391 GND 0.001706f
C6855 VDD.n1392 GND 0.001706f
C6856 VDD.n1393 GND 8.53e-19
C6857 VDD.n1394 GND 9.03e-19
C6858 VDD.n1395 GND 0.018487f
C6859 VDD.n1396 GND 8.53e-19
C6860 VDD.n1397 GND 0.001706f
C6861 VDD.t384 GND 0.117408f
C6862 VDD.n1398 GND 0.001706f
C6863 VDD.n1399 GND 0.001706f
C6864 VDD.n1400 GND 0.001706f
C6865 VDD.t266 GND 0.117408f
C6866 VDD.n1401 GND 0.001706f
C6867 VDD.n1402 GND 0.001706f
C6868 VDD.n1403 GND 0.001706f
C6869 VDD.n1404 GND 8.53e-19
C6870 VDD.n1405 GND 9.03e-19
C6871 VDD.n1406 GND 0.010359f
C6872 VDD.n1407 GND 0.010359f
C6873 VDD.n1408 GND 9.03e-19
C6874 VDD.n1409 GND 0.010359f
C6875 VDD.n1410 GND 8.53e-19
C6876 VDD.n1411 GND 0.001706f
C6877 VDD.n1412 GND 0.119161f
C6878 VDD.n1413 GND 0.001706f
C6879 VDD.n1414 GND 0.001706f
C6880 VDD.t193 GND 0.117408f
C6881 VDD.n1415 GND 0.001706f
C6882 VDD.n1416 GND 0.001706f
C6883 VDD.n1417 GND 0.001706f
C6884 VDD.n1418 GND 0.001706f
C6885 VDD.n1419 GND 0.001706f
C6886 VDD.n1420 GND 0.001706f
C6887 VDD.n1421 GND 0.001706f
C6888 VDD.n1422 GND 0.001706f
C6889 VDD.n1423 GND 0.05958f
C6890 VDD.n1424 GND 0.001706f
C6891 VDD.n1425 GND 0.001706f
C6892 VDD.n1426 GND 0.098132f
C6893 VDD.n1427 GND 0.001706f
C6894 VDD.n1428 GND 0.001706f
C6895 VDD.n1429 GND 0.119161f
C6896 VDD.n1430 GND 0.001706f
C6897 VDD.n1431 GND 0.001706f
C6898 VDD.n1432 GND 0.001706f
C6899 VDD.n1433 GND 0.038552f
C6900 VDD.n1434 GND 0.001706f
C6901 VDD.t81 GND 0.117408f
C6902 VDD.n1435 GND 0.001706f
C6903 VDD.n1436 GND 0.001706f
C6904 VDD.n1437 GND 0.001706f
C6905 VDD.n1438 GND 8.53e-19
C6906 VDD.n1439 GND 9.03e-19
C6907 VDD.n1440 GND 0.010359f
C6908 VDD.n1441 GND 9.03e-19
C6909 VDD.n1442 GND 8.53e-19
C6910 VDD.n1443 GND 0.010359f
C6911 VDD.n1444 GND 9.03e-19
C6912 VDD.n1445 GND 0.010359f
C6913 VDD.n1446 GND 0.010359f
C6914 VDD.n1447 GND 8.53e-19
C6915 VDD.n1448 GND 0.001706f
C6916 VDD.n1449 GND 0.119161f
C6917 VDD.n1450 GND 0.001706f
C6918 VDD.n1451 GND 0.001706f
C6919 VDD.n1452 GND 8.53e-19
C6920 VDD.n1453 GND 9.03e-19
C6921 VDD.n1454 GND 8.53e-19
C6922 VDD.n1455 GND 0.001706f
C6923 VDD.t93 GND 0.117408f
C6924 VDD.n1456 GND 0.001706f
C6925 VDD.n1457 GND 0.001706f
C6926 VDD.t350 GND 0.117408f
C6927 VDD.n1458 GND 0.001706f
C6928 VDD.n1459 GND 0.001706f
C6929 VDD.n1460 GND 0.001003f
C6930 VDD.n1461 GND 0.012142f
C6931 VDD.n1462 GND 0.001706f
C6932 VDD.n1463 GND 0.077104f
C6933 VDD.n1464 GND 0.001706f
C6934 VDD.t91 GND 0.117408f
C6935 VDD.n1465 GND 0.094628f
C6936 VDD.n1466 GND 0.001706f
C6937 VDD.n1467 GND 0.001706f
C6938 VDD.n1468 GND 0.001706f
C6939 VDD.n1469 GND 0.014019f
C6940 VDD.n1470 GND 0.001706f
C6941 VDD.n1471 GND 0.012142f
C6942 VDD.n1472 GND 0.035047f
C6943 VDD.n1473 GND 0.001706f
C6944 VDD.t334 GND 0.117408f
C6945 VDD.n1474 GND 0.001706f
C6946 VDD.n1475 GND 0.001706f
C6947 VDD.n1476 GND 9.03e-19
C6948 VDD.n1477 GND 0.014037f
C6949 VDD.n1478 GND 0.010359f
C6950 VDD.n1479 GND 9.03e-19
C6951 VDD.n1480 GND 8.53e-19
C6952 VDD.n1481 GND 0.001706f
C6953 VDD.n1482 GND 8.53e-19
C6954 VDD.n1483 GND 9.03e-19
C6955 VDD.t87 GND 0.117408f
C6956 VDD.t534 GND 0.117408f
C6957 VDD.n1484 GND 0.085866f
C6958 VDD.n1485 GND 0.001706f
C6959 VDD.n1486 GND 0.001706f
C6960 VDD.n1487 GND 8.53e-19
C6961 VDD.n1488 GND 9.03e-19
C6962 VDD.n1489 GND 0.002444f
C6963 VDD.n1490 GND 8.53e-19
C6964 VDD.n1491 GND 0.001706f
C6965 VDD.t95 GND 0.117408f
C6966 VDD.n1492 GND 0.001706f
C6967 VDD.n1493 GND 0.001706f
C6968 VDD.n1494 GND 0.001706f
C6969 VDD.t242 GND 0.117408f
C6970 VDD.n1495 GND 0.001706f
C6971 VDD.n1496 GND 0.001706f
C6972 VDD.n1497 GND 0.001706f
C6973 VDD.n1498 GND 0.001706f
C6974 VDD.n1499 GND 0.001706f
C6975 VDD.n1500 GND 0.119161f
C6976 VDD.n1501 GND 0.001706f
C6977 VDD.n1502 GND 0.001706f
C6978 VDD.t498 GND 0.117408f
C6979 VDD.n1503 GND 0.001706f
C6980 VDD.n1504 GND 0.001706f
C6981 VDD.n1505 GND 0.001706f
C6982 VDD.n1506 GND 0.001229f
C6983 VDD.n1507 GND 0.001706f
C6984 VDD.n1508 GND 0.012142f
C6985 VDD.n1509 GND 0.001706f
C6986 VDD.n1510 GND 0.073599f
C6987 VDD.n1511 GND 0.001706f
C6988 VDD.n1512 GND 0.001706f
C6989 VDD.n1513 GND 0.112151f
C6990 VDD.n1514 GND 0.001706f
C6991 VDD.n1515 GND 0.001706f
C6992 VDD.n1516 GND 0.010514f
C6993 VDD.n1517 GND 0.001706f
C6994 VDD.n1518 GND 0.001706f
C6995 VDD.n1519 GND 0.001706f
C6996 VDD.n1520 GND 0.049066f
C6997 VDD.n1521 GND 0.001706f
C6998 VDD.t468 GND 0.117408f
C6999 VDD.n1522 GND 0.001706f
C7000 VDD.n1523 GND 0.001706f
C7001 VDD.n1524 GND 0.001706f
C7002 VDD.n1525 GND 0.001706f
C7003 VDD.n1526 GND 0.001706f
C7004 VDD.n1527 GND 0.087618f
C7005 VDD.n1528 GND 0.001706f
C7006 VDD.n1529 GND 0.001706f
C7007 VDD.t470 GND 0.117408f
C7008 VDD.n1530 GND 0.001706f
C7009 VDD.n1531 GND 0.001706f
C7010 VDD.n1532 GND 0.001706f
C7011 VDD.n1533 GND 0.001706f
C7012 VDD.n1534 GND 0.001706f
C7013 VDD.n1535 GND 0.001706f
C7014 VDD.n1536 GND 8.53e-19
C7015 VDD.n1537 GND 9.03e-19
C7016 VDD.n1538 GND 0.005502f
C7017 VDD.n1539 GND 8.53e-19
C7018 VDD.n1540 GND 0.001706f
C7019 VDD.n1541 GND 0.001706f
C7020 VDD.n1542 GND 0.003723f
C7021 VDD.n1543 GND 0.003723f
C7022 VDD.n1544 GND 0.108646f
C7023 VDD.n1545 GND 0.003723f
C7024 VDD.n1546 GND 0.001706f
C7025 VDD.n1547 GND 0.001706f
C7026 VDD.n1548 GND 0.078856f
C7027 VDD.n1549 GND 0.003727f
C7028 VDD.n1557 GND 0.18575f
C7029 VDD.n1566 GND 0.001706f
C7030 VDD.n1567 GND 0.001706f
C7031 VDD.n1568 GND 0.001706f
C7032 VDD.n1569 GND 0.001706f
C7033 VDD.n1570 GND 0.001706f
C7034 VDD.n1571 GND 0.183998f
C7035 VDD.n1572 GND 0.001706f
C7036 VDD.n1573 GND 0.001706f
C7037 VDD.n1574 GND 0.001706f
C7038 VDD.n1575 GND 0.001706f
C7039 VDD.n1576 GND 0.22255f
C7040 VDD.t542 GND 0.119161f
C7041 VDD.n1577 GND 0.001706f
C7042 VDD.n1578 GND 0.001706f
C7043 VDD.n1579 GND 0.001706f
C7044 VDD.n1580 GND 0.238321f
C7045 VDD.n1581 GND 0.001706f
C7046 VDD.n1582 GND 0.001706f
C7047 VDD.n1583 GND 0.001706f
C7048 VDD.t4 GND 0.119161f
C7049 VDD.n1584 GND 0.001706f
C7050 VDD.n1585 GND 0.001706f
C7051 VDD.n1586 GND 0.001706f
C7052 VDD.t77 GND 0.119161f
C7053 VDD.n1587 GND 0.001706f
C7054 VDD.n1588 GND 0.001706f
C7055 VDD.n1589 GND 0.001706f
C7056 VDD.t174 GND 0.119161f
C7057 VDD.n1590 GND 0.176989f
C7058 VDD.n1591 GND 0.001706f
C7059 VDD.n1592 GND 0.001706f
C7060 VDD.n1593 GND 0.001706f
C7061 VDD.n1594 GND 0.138437f
C7062 VDD.n1595 GND 0.001706f
C7063 VDD.n1596 GND 0.001706f
C7064 VDD.n1597 GND 0.001706f
C7065 VDD.n1598 GND 0.176989f
C7066 VDD.t6 GND 0.119161f
C7067 VDD.n1599 GND 0.001706f
C7068 VDD.n1600 GND 0.001706f
C7069 VDD.n1601 GND 0.001706f
C7070 VDD.n1602 GND 0.215541f
C7071 VDD.n1603 GND 0.001706f
C7072 VDD.n1604 GND 0.003781f
C7073 VDD.n1605 GND 0.003781f
C7074 VDD.n1606 GND 0.315425f
C7075 VDD.t79 GND 0.119161f
C7076 VDD.n1607 GND 0.003781f
C7077 VDD.n1608 GND 0.001706f
C7078 VDD.n1609 GND 0.001706f
C7079 VDD.n1617 GND 0.001706f
C7080 VDD.n1618 GND 0.001706f
C7081 VDD.n1619 GND 0.001706f
C7082 VDD.n1620 GND 0.001706f
C7083 VDD.n1621 GND 0.001706f
C7084 VDD.n1622 GND 0.001706f
C7085 VDD.n1623 GND 0.001706f
C7086 VDD.n1624 GND 0.001706f
C7087 VDD.n1625 GND 0.001706f
C7088 VDD.n1626 GND 0.001706f
C7089 VDD.n1627 GND 0.001706f
C7090 VDD.n1628 GND 0.001706f
C7091 VDD.n1629 GND 0.001706f
C7092 VDD.n1630 GND 0.001706f
C7093 VDD.n1631 GND 0.001706f
C7094 VDD.n1632 GND 0.001706f
C7095 VDD.n1633 GND 0.001706f
C7096 VDD.n1634 GND 0.001706f
C7097 VDD.n1635 GND 0.001706f
C7098 VDD.n1636 GND 0.001706f
C7099 VDD.n1637 GND 0.001706f
C7100 VDD.n1638 GND 0.001706f
C7101 VDD.n1639 GND 0.001706f
C7102 VDD.n1640 GND 0.001706f
C7103 VDD.n1641 GND 0.001706f
C7104 VDD.n1642 GND 0.001706f
C7105 VDD.n1643 GND 0.001706f
C7106 VDD.n1644 GND 0.001706f
C7107 VDD.n1645 GND 0.003795f
C7108 VDD.n1646 GND 0.003795f
C7109 VDD.n1647 GND 0.403043f
C7110 VDD.n1649 GND 0.003795f
C7111 VDD.n1650 GND 0.003795f
C7112 VDD.n1651 GND 0.003781f
C7113 VDD.n1652 GND 0.001706f
C7114 VDD.n1653 GND 0.001706f
C7115 VDD.n1654 GND 0.141941f
C7116 VDD.n1655 GND 0.001706f
C7117 VDD.n1656 GND 0.001706f
C7118 VDD.n1657 GND 0.001706f
C7119 VDD.n1658 GND 0.001706f
C7120 VDD.n1659 GND 0.001706f
C7121 VDD.t295 GND 0.119161f
C7122 VDD.n1660 GND 0.180493f
C7123 VDD.n1661 GND 0.001706f
C7124 VDD.n1662 GND 0.001706f
C7125 VDD.n1663 GND 0.001706f
C7126 VDD.n1664 GND 0.001706f
C7127 VDD.n1665 GND 0.001706f
C7128 VDD.n1666 GND 0.219045f
C7129 VDD.n1667 GND 0.001706f
C7130 VDD.n1668 GND 0.001706f
C7131 VDD.n1669 GND 0.001706f
C7132 VDD.n1670 GND 0.001706f
C7133 VDD.n1671 GND 0.001706f
C7134 VDD.n1672 GND 0.138437f
C7135 VDD.n1673 GND 0.238321f
C7136 VDD.n1674 GND 0.001706f
C7137 VDD.n1675 GND 0.001706f
C7138 VDD.n1676 GND 0.001706f
C7139 VDD.n1677 GND 0.001706f
C7140 VDD.n1678 GND 0.001706f
C7141 VDD.n1679 GND 0.219045f
C7142 VDD.n1680 GND 0.001706f
C7143 VDD.n1681 GND 0.001706f
C7144 VDD.n1682 GND 0.001706f
C7145 VDD.n1683 GND 0.001706f
C7146 VDD.n1684 GND 0.001706f
C7147 VDD.n1685 GND 0.215541f
C7148 VDD.n1686 GND 0.180493f
C7149 VDD.n1687 GND 0.001706f
C7150 VDD.n1688 GND 0.001706f
C7151 VDD.n1689 GND 0.001706f
C7152 VDD.n1690 GND 0.001706f
C7153 VDD.n1691 GND 0.001706f
C7154 VDD.n1692 GND 0.141941f
C7155 VDD.n1693 GND 0.001706f
C7156 VDD.n1694 GND 0.001706f
C7157 VDD.n1695 GND 0.001706f
C7158 VDD.n1696 GND 0.001706f
C7159 VDD.n1697 GND 0.001706f
C7160 VDD.t97 GND 0.119161f
C7161 VDD.n1698 GND 0.134932f
C7162 VDD.n1699 GND 0.001706f
C7163 VDD.n1700 GND 0.001706f
C7164 VDD.n1701 GND 0.001706f
C7165 VDD.n1702 GND 0.001706f
C7166 VDD.n1703 GND 0.001706f
C7167 VDD.n1704 GND 0.001706f
C7168 VDD.n1705 GND 0.173484f
C7169 VDD.n1706 GND 0.001706f
C7170 VDD.n1707 GND 0.001706f
C7171 VDD.n1708 GND 0.001706f
C7172 VDD.n1709 GND 9.17e-19
C7173 VDD.n1710 GND 9.03e-19
C7174 VDD.n1711 GND 0.002444f
C7175 VDD.n1712 GND 9.03e-19
C7176 VDD.n1713 GND 0.002444f
C7177 VDD.n1714 GND 8.53e-19
C7178 VDD.n1715 GND 0.001706f
C7179 VDD.n1716 GND 9.03e-19
C7180 VDD.n1717 GND 0.002313f
C7181 VDD.n1718 GND 8.53e-19
C7182 VDD.n1719 GND 9.03e-19
C7183 VDD.n1720 GND 8.53e-19
C7184 VDD.n1721 GND 0.002444f
C7185 VDD.n1722 GND 0.002444f
C7186 VDD.n1723 GND 8.53e-19
C7187 VDD.n1724 GND 9.03e-19
C7188 VDD.n1725 GND 0.001706f
C7189 VDD.n1726 GND 0.001706f
C7190 VDD.n1727 GND 9.03e-19
C7191 VDD.n1728 GND 8.53e-19
C7192 VDD.n1729 GND 0.002444f
C7193 VDD.n1730 GND 0.002444f
C7194 VDD.n1731 GND 8.53e-19
C7195 VDD.n1732 GND 9.03e-19
C7196 VDD.n1733 GND 8.53e-19
C7197 VDD.n1734 GND 0.001706f
C7198 VDD.n1735 GND 9.03e-19
C7199 VDD.n1736 GND 8.53e-19
C7200 VDD.n1737 GND 0.002444f
C7201 VDD.n1738 GND 0.005502f
C7202 VDD.n1739 GND 8.53e-19
C7203 VDD.n1740 GND 9.03e-19
C7204 VDD.n1741 GND 0.001706f
C7205 VDD.n1742 GND 0.001706f
C7206 VDD.n1743 GND 0.001029f
C7207 VDD.n1744 GND 0.001706f
C7208 VDD.n1745 GND 0.001706f
C7209 VDD.n1746 GND 0.001706f
C7210 VDD.n1747 GND 0.001706f
C7211 VDD.n1748 GND 0.001706f
C7212 VDD.n1749 GND 0.001706f
C7213 VDD.t348 GND 0.119161f
C7214 VDD.n1750 GND 0.212036f
C7215 VDD.n1751 GND 0.001706f
C7216 VDD.n1752 GND 0.001706f
C7217 VDD.n1753 GND 0.001706f
C7218 VDD.n1754 GND 0.001706f
C7219 VDD.n1755 GND 9.03e-19
C7220 VDD.n1756 GND 9.17e-19
C7221 VDD.n1757 GND 0.001029f
C7222 VDD.n1758 GND 0.001706f
C7223 VDD.n1759 GND 0.001706f
C7224 VDD.n1760 GND 0.120913f
C7225 VDD.t452 GND 0.117408f
C7226 VDD.n1761 GND 0.001706f
C7227 VDD.n1762 GND 0.001706f
C7228 VDD.n1763 GND 0.001706f
C7229 VDD.n1764 GND 0.001706f
C7230 VDD.n1765 GND 0.001706f
C7231 VDD.n1766 GND 0.001706f
C7232 VDD.n1767 GND 0.001706f
C7233 VDD.n1768 GND 0.001706f
C7234 VDD.n1769 GND 0.001706f
C7235 VDD.n1770 GND 0.001706f
C7236 VDD.n1771 GND 0.001706f
C7237 VDD.n1772 GND 0.001706f
C7238 VDD.n1773 GND 0.001706f
C7239 VDD.n1774 GND 0.001706f
C7240 VDD.n1775 GND 0.001706f
C7241 VDD.n1776 GND 0.001706f
C7242 VDD.n1777 GND 0.001706f
C7243 VDD.n1778 GND 0.001706f
C7244 VDD.n1779 GND 0.001706f
C7245 VDD.n1780 GND 0.001706f
C7246 VDD.n1781 GND 0.001706f
C7247 VDD.n1782 GND 0.001706f
C7248 VDD.n1783 GND 0.001706f
C7249 VDD.n1784 GND 0.001706f
C7250 VDD.n1785 GND 0.001706f
C7251 VDD.n1786 GND 0.001706f
C7252 VDD.n1787 GND 0.001706f
C7253 VDD.n1788 GND 0.001706f
C7254 VDD.n1789 GND 0.003727f
C7255 VDD.n1790 GND 0.003723f
C7256 VDD.n1791 GND 0.003723f
C7257 VDD.n1792 GND 0.012266f
C7258 VDD.n1793 GND 0.003723f
C7259 VDD.n1794 GND 0.001706f
C7260 VDD.n1795 GND 0.003723f
C7261 VDD.n1796 GND 0.003727f
C7262 VDD.n1797 GND 0.003727f
C7263 VDD.n1798 GND 0.001706f
C7264 VDD.n1799 GND 0.001706f
C7265 VDD.n1800 GND 0.001706f
C7266 VDD.n1801 GND 0.001706f
C7267 VDD.n1802 GND 0.001706f
C7268 VDD.n1803 GND 0.001706f
C7269 VDD.n1804 GND 0.001706f
C7270 VDD.n1805 GND 0.001706f
C7271 VDD.n1806 GND 0.001706f
C7272 VDD.n1807 GND 0.001706f
C7273 VDD.n1808 GND 0.001706f
C7274 VDD.n1809 GND 0.001706f
C7275 VDD.n1810 GND 0.001706f
C7276 VDD.n1811 GND 0.001706f
C7277 VDD.n1812 GND 0.001706f
C7278 VDD.n1813 GND 0.001706f
C7279 VDD.n1814 GND 0.001706f
C7280 VDD.n1815 GND 0.001706f
C7281 VDD.n1816 GND 0.001706f
C7282 VDD.n1817 GND 0.001706f
C7283 VDD.n1818 GND 0.001706f
C7284 VDD.n1819 GND 0.001706f
C7285 VDD.n1820 GND 0.001706f
C7286 VDD.n1821 GND 0.001706f
C7287 VDD.n1822 GND 0.001706f
C7288 VDD.n1823 GND 0.001706f
C7289 VDD.n1824 GND 0.001706f
C7290 VDD.n1825 GND 0.001706f
C7291 VDD.n1826 GND 0.001706f
C7292 VDD.n1827 GND 0.003727f
C7293 VDD.n1828 GND 0.003727f
C7294 VDD.n1829 GND 0.119161f
C7295 VDD.n1831 GND 0.003727f
C7296 VDD.n1832 GND 0.003727f
C7297 VDD.n1833 GND 0.003723f
C7298 VDD.n1834 GND 0.001706f
C7299 VDD.n1835 GND 0.001706f
C7300 VDD.n1836 GND 0.001706f
C7301 VDD.t50 GND 0.117408f
C7302 VDD.n1837 GND 0.033295f
C7303 VDD.n1838 GND 0.001706f
C7304 VDD.n1839 GND 0.001706f
C7305 VDD.n1840 GND 0.001706f
C7306 VDD.n1841 GND 0.001706f
C7307 VDD.n1842 GND 0.001706f
C7308 VDD.n1843 GND 0.001706f
C7309 VDD.t83 GND 0.117408f
C7310 VDD.n1844 GND 0.071847f
C7311 VDD.n1845 GND 0.070094f
C7312 VDD.n1846 GND 0.001706f
C7313 VDD.n1847 GND 9.03e-19
C7314 VDD.n1848 GND 9.03e-19
C7315 VDD.n1849 GND 8.53e-19
C7316 VDD.n1850 GND 0.002444f
C7317 VDD.n1851 GND 0.002444f
C7318 VDD.n1852 GND 0.002444f
C7319 VDD.n1853 GND 9.03e-19
C7320 VDD.n1854 GND 8.53e-19
C7321 VDD.n1855 GND 0.001706f
C7322 VDD.n1856 GND 9.03e-19
C7323 VDD.n1857 GND 8.53e-19
C7324 VDD.n1858 GND 0.002444f
C7325 VDD.n1859 GND 0.002444f
C7326 VDD.n1860 GND 8.53e-19
C7327 VDD.n1861 GND 9.03e-19
C7328 VDD.n1862 GND 0.001706f
C7329 VDD.n1863 GND 0.031543f
C7330 VDD.t99 GND 0.117408f
C7331 VDD.n1864 GND 0.110399f
C7332 VDD.n1865 GND 0.001706f
C7333 VDD.n1866 GND 0.001706f
C7334 VDD.n1867 GND 0.001706f
C7335 VDD.n1868 GND 0.001706f
C7336 VDD.n1869 GND 0.001706f
C7337 VDD.n1870 GND 0.001706f
C7338 VDD.n1871 GND 0.050818f
C7339 VDD.n1872 GND 0.001706f
C7340 VDD.n1873 GND 0.001706f
C7341 VDD.n1874 GND 0.001706f
C7342 VDD.n1875 GND 0.001706f
C7343 VDD.n1876 GND 0.001706f
C7344 VDD.n1877 GND 0.001706f
C7345 VDD.n1878 GND 0.08937f
C7346 VDD.n1879 GND 0.001706f
C7347 VDD.n1880 GND 0.001706f
C7348 VDD.n1881 GND 0.001706f
C7349 VDD.n1882 GND 0.001706f
C7350 VDD.n1883 GND 0.001706f
C7351 VDD.n1884 GND 0.119161f
C7352 VDD.n1885 GND 0.001706f
C7353 VDD.n1886 GND 0.001706f
C7354 VDD.n1887 GND 0.001706f
C7355 VDD.n1888 GND 0.001706f
C7356 VDD.n1889 GND 0.001706f
C7357 VDD.n1890 GND 0.02979f
C7358 VDD.n1891 GND 0.001706f
C7359 VDD.n1892 GND 0.001706f
C7360 VDD.n1893 GND 0.001706f
C7361 VDD.n1894 GND 0.001706f
C7362 VDD.n1895 GND 0.001706f
C7363 VDD.n1896 GND 0.001706f
C7364 VDD.n1897 GND 0.068342f
C7365 VDD.n1898 GND 0.001706f
C7366 VDD.n1899 GND 0.009463f
C7367 VDD.n1900 GND 0.004145f
C7368 VDD.n1901 GND 0.001229f
C7369 VDD.n1902 GND 0.001706f
C7370 VDD.n1903 GND 0.001706f
C7371 VDD.n1904 GND 0.001706f
C7372 VDD.n1905 GND 0.008762f
C7373 VDD.n1906 GND 0.001706f
C7374 VDD.n1907 GND 0.001706f
C7375 VDD.n1908 GND 0.001706f
C7376 VDD.n1909 GND 0.001706f
C7377 VDD.n1910 GND 0.001706f
C7378 VDD.n1911 GND 0.001706f
C7379 VDD.n1912 GND 0.047314f
C7380 VDD.n1913 GND 0.091123f
C7381 VDD.n1914 GND 0.001706f
C7382 VDD.n1915 GND 9.03e-19
C7383 VDD.n1916 GND 9.03e-19
C7384 VDD.n1917 GND 8.53e-19
C7385 VDD.n1918 GND 0.002444f
C7386 VDD.n1919 GND 0.002444f
C7387 VDD.n1920 GND 0.003712f
C7388 VDD.n1921 GND 9.03e-19
C7389 VDD.n1922 GND 8.53e-19
C7390 VDD.n1923 GND 0.001706f
C7391 VDD.n1924 GND 9.03e-19
C7392 VDD.n1925 GND 8.53e-19
C7393 VDD.n1926 GND 0.002444f
C7394 VDD.n1927 GND 0.002444f
C7395 VDD.n1928 GND 8.53e-19
C7396 VDD.n1929 GND 9.03e-19
C7397 VDD.n1930 GND 0.001706f
C7398 VDD.n1931 GND 0.052571f
C7399 VDD.n1932 GND 0.001706f
C7400 VDD.n1933 GND 0.001706f
C7401 VDD.n1934 GND 0.001706f
C7402 VDD.n1935 GND 9.03e-19
C7403 VDD.n1936 GND 8.53e-19
C7404 VDD.n1937 GND 0.010359f
C7405 VDD.n1938 GND 0.010359f
C7406 VDD.n1939 GND 8.53e-19
C7407 VDD.n1940 GND 0.001129f
C7408 VDD.n1941 GND 0.001706f
C7409 VDD.n1942 GND 0.106894f
C7410 VDD.n1943 GND 0.001706f
C7411 VDD.n1944 GND 0.001706f
C7412 VDD.n1945 GND 0.119161f
C7413 VDD.n1946 GND 0.001706f
C7414 VDD.n1947 GND 0.001706f
C7415 VDD.n1948 GND 0.001706f
C7416 VDD.n1949 GND 0.001706f
C7417 VDD.n1950 GND 0.001706f
C7418 VDD.n1951 GND 0.001706f
C7419 VDD.n1952 GND 0.001706f
C7420 VDD.t273 GND 0.117408f
C7421 VDD.n1953 GND 0.001706f
C7422 VDD.n1954 GND 0.001706f
C7423 VDD.n1955 GND 0.043809f
C7424 VDD.n1956 GND 0.001706f
C7425 VDD.n1957 GND 8.53e-19
C7426 VDD.n1958 GND 9.03e-19
C7427 VDD.n1959 GND 8.53e-19
C7428 VDD.n1960 GND 9.03e-19
C7429 VDD.n1961 GND 0.010215f
C7430 VDD.n1962 GND 0.010359f
C7431 VDD.n1963 GND 0.006187f
C7432 VDD.n1964 GND 0.009208f
C7433 VDD.n1965 GND 0.098305f
C7434 VDD.n1966 GND 1.00116f
C7435 VDD.n1967 GND 0.098017f
C7436 VDD.n1968 GND 0.005467f
C7437 VDD.n1969 GND 0.010359f
C7438 VDD.n1970 GND 8.53e-19
C7439 VDD.n1971 GND 0.001706f
C7440 VDD.n1972 GND 9.03e-19
C7441 VDD.n1973 GND 8.53e-19
C7442 VDD.n1974 GND 9.03e-19
C7443 VDD.n1975 GND 8.53e-19
C7444 VDD.n1976 GND 9.03e-19
C7445 VDD.n1977 GND 8.53e-19
C7446 VDD.n1978 GND 0.010359f
C7447 VDD.n1979 GND 0.010359f
C7448 VDD.n1980 GND 8.53e-19
C7449 VDD.n1981 GND 9.03e-19
C7450 VDD.n1982 GND 0.001706f
C7451 VDD.n1983 GND 0.064837f
C7452 VDD.n1984 GND 0.001706f
C7453 VDD.n1985 GND 0.011071f
C7454 VDD.n1986 GND 0.005301f
C7455 VDD.n1987 GND 0.001706f
C7456 VDD.n1988 GND 0.001706f
C7457 VDD.n1989 GND 0.001706f
C7458 VDD.n1990 GND 0.001003f
C7459 VDD.n1991 GND 0.001706f
C7460 VDD.n1992 GND 0.082361f
C7461 VDD.n1993 GND 0.056076f
C7462 VDD.n1994 GND 0.001706f
C7463 VDD.n1995 GND 9.03e-19
C7464 VDD.n1996 GND 9.03e-19
C7465 VDD.n1997 GND 8.53e-19
C7466 VDD.n1998 GND 0.018487f
C7467 VDD.n1999 GND 0.018487f
C7468 VDD.n2000 GND 0.018487f
C7469 VDD.n2001 GND 9.03e-19
C7470 VDD.n2002 GND 8.53e-19
C7471 VDD.n2003 GND 0.001706f
C7472 VDD.n2004 GND 9.03e-19
C7473 VDD.n2005 GND 8.53e-19
C7474 VDD.n2006 GND 0.018487f
C7475 VDD.n2007 GND 0.018487f
C7476 VDD.n2008 GND 8.53e-19
C7477 VDD.n2009 GND 9.03e-19
C7478 VDD.n2010 GND 0.001706f
C7479 VDD.n2011 GND 0.017524f
C7480 VDD.n2012 GND 0.001706f
C7481 VDD.n2013 GND 0.001706f
C7482 VDD.n2014 GND 8.53e-19
C7483 VDD.n2015 GND 9.03e-19
C7484 VDD.n2016 GND 0.001706f
C7485 VDD.n2017 GND 0.001706f
C7486 VDD.n2018 GND 9.03e-19
C7487 VDD.n2019 GND 8.53e-19
C7488 VDD.n2020 GND 0.010359f
C7489 VDD.n2021 GND 0.010359f
C7490 VDD.n2022 GND 8.53e-19
C7491 VDD.n2023 GND 9.03e-19
C7492 VDD.n2024 GND 0.001706f
C7493 VDD.n2025 GND 0.103389f
C7494 VDD.n2026 GND 0.001706f
C7495 VDD.n2027 GND 0.001706f
C7496 VDD.n2028 GND 0.001706f
C7497 VDD.n2029 GND 0.001706f
C7498 VDD.n2030 GND 0.001706f
C7499 VDD.t10 GND 0.119161f
C7500 VDD.n2031 GND 0.001706f
C7501 VDD.n2032 GND 0.001706f
C7502 VDD.n2033 GND 0.001706f
C7503 VDD.n2034 GND 0.001706f
C7504 VDD.n2035 GND 0.001706f
C7505 VDD.n2036 GND 0.001706f
C7506 VDD.n2037 GND 0.001706f
C7507 VDD.n2038 GND 0.001706f
C7508 VDD.n2039 GND 0.001706f
C7509 VDD.n2040 GND 0.001706f
C7510 VDD.n2041 GND 0.001706f
C7511 VDD.n2042 GND 0.001706f
C7512 VDD.n2043 GND 0.001706f
C7513 VDD.n2044 GND 0.001706f
C7514 VDD.n2045 GND 0.040304f
C7515 VDD.n2046 GND 0.001706f
C7516 VDD.n2047 GND 0.001706f
C7517 VDD.n2048 GND 0.001706f
C7518 VDD.n2049 GND 0.001706f
C7519 VDD.n2050 GND 0.001706f
C7520 VDD.n2051 GND 0.078856f
C7521 VDD.n2052 GND 0.001706f
C7522 VDD.n2053 GND 0.001706f
C7523 VDD.n2054 GND 0.001706f
C7524 VDD.n2055 GND 0.001706f
C7525 VDD.n2056 GND 0.001706f
C7526 VDD.n2057 GND 0.001706f
C7527 VDD.n2058 GND 0.022781f
C7528 VDD.n2059 GND 0.001706f
C7529 VDD.n2060 GND 9.03e-19
C7530 VDD.n2061 GND 9.03e-19
C7531 VDD.n2062 GND 8.53e-19
C7532 VDD.n2063 GND 0.010359f
C7533 VDD.n2064 GND 0.010359f
C7534 VDD.n2065 GND 0.010359f
C7535 VDD.n2066 GND 8.53e-19
C7536 VDD.n2067 GND 9.03e-19
C7537 VDD.n2068 GND 8.53e-19
C7538 VDD.n2069 GND 9.03e-19
C7539 VDD.n2070 GND 8.53e-19
C7540 VDD.n2071 GND 0.010359f
C7541 VDD.n2072 GND 0.010359f
C7542 VDD.n2073 GND 8.53e-19
C7543 VDD.n2074 GND 8.78e-19
C7544 VDD.n2075 GND 8.78e-19
C7545 VDD.n2076 GND 0.001706f
C7546 VDD.n2077 GND 0.061333f
C7547 VDD.n2078 GND 0.080609f
C7548 VDD.n2079 GND 0.001706f
C7549 VDD.n2080 GND 9.03e-19
C7550 VDD.n2081 GND 9.03e-19
C7551 VDD.n2082 GND 8.53e-19
C7552 VDD.n2083 GND 0.018487f
C7553 VDD.n2084 GND 0.018487f
C7554 VDD.n2085 GND 9.03e-19
C7555 VDD.n2086 GND 8.53e-19
C7556 VDD.n2087 GND 0.018487f
C7557 VDD.n2088 GND 0.018487f
C7558 VDD.n2089 GND 8.53e-19
C7559 VDD.n2090 GND 9.03e-19
C7560 VDD.n2091 GND 0.001706f
C7561 VDD.n2092 GND 0.042057f
C7562 VDD.n2093 GND 0.001706f
C7563 VDD.n2094 GND 0.001706f
C7564 VDD.n2095 GND 0.003505f
C7565 VDD.n2096 GND 0.001706f
C7566 VDD.n2097 GND 9.03e-19
C7567 VDD.n2098 GND 8.53e-19
C7568 VDD.n2099 GND 0.010359f
C7569 VDD.n2100 GND 0.010359f
C7570 VDD.n2101 GND 8.53e-19
C7571 VDD.n2102 GND 9.03e-19
C7572 VDD.n2103 GND 0.001706f
C7573 VDD.n2104 GND 0.117408f
C7574 VDD.n2105 GND 0.001706f
C7575 VDD.n2106 GND 0.001706f
C7576 VDD.n2107 GND 0.001706f
C7577 VDD.n2108 GND 0.001706f
C7578 VDD.n2109 GND 0.001706f
C7579 VDD.n2110 GND 0.001706f
C7580 VDD.t52 GND 0.117408f
C7581 VDD.n2111 GND 0.019276f
C7582 VDD.n2112 GND 0.119161f
C7583 VDD.n2113 GND 0.001706f
C7584 VDD.n2114 GND 9.03e-19
C7585 VDD.n2115 GND 8.53e-19
C7586 VDD.n2116 GND 0.018487f
C7587 VDD.n2117 GND 0.018487f
C7588 VDD.n2118 GND 8.53e-19
C7589 VDD.n2119 GND 8.53e-19
C7590 VDD.n2120 GND 9.03e-19
C7591 VDD.n2121 GND 0.001706f
C7592 VDD.n2122 GND 0.084113f
C7593 VDD.n2123 GND 0.001706f
C7594 VDD.n2124 GND 9.03e-19
C7595 VDD.n2125 GND 8.53e-19
C7596 VDD.n2126 GND 0.010359f
C7597 VDD.n2127 GND 0.010359f
C7598 VDD.n2128 GND 8.53e-19
C7599 VDD.n2129 GND 9.03e-19
C7600 VDD.n2130 GND 0.001706f
C7601 VDD.n2131 GND 0.0368f
C7602 VDD.n2132 GND 0.001706f
C7603 VDD.n2133 GND 0.001706f
C7604 VDD.n2134 GND 9.03e-19
C7605 VDD.n2135 GND 0.005814f
C7606 VDD.n2136 GND 0.012142f
C7607 VDD.n2137 GND 0.011785f
C7608 VDD.n2138 GND 0.001706f
C7609 VDD.n2139 GND 0.075352f
C7610 VDD.n2140 GND 0.001706f
C7611 VDD.n2141 GND 0.001706f
C7612 VDD.n2142 GND 0.001706f
C7613 VDD.n2143 GND 0.001706f
C7614 VDD.n2144 GND 0.001706f
C7615 VDD.n2145 GND 0.113904f
C7616 VDD.n2146 GND 0.001706f
C7617 VDD.n2147 GND 0.001706f
C7618 VDD.n2148 GND 0.007589f
C7619 VDD.n2149 GND 0.001706f
C7620 VDD.n2150 GND 0.012142f
C7621 VDD.n2151 GND 0.010624f
C7622 VDD.n2152 GND 0.001706f
C7623 VDD.n2153 GND 0.015771f
C7624 VDD.n2154 GND 0.001706f
C7625 VDD.n2155 GND 0.001706f
C7626 VDD.n2156 GND 0.001706f
C7627 VDD.n2157 GND 0.001706f
C7628 VDD.n2158 GND 8.53e-19
C7629 VDD.n2159 GND 9.03e-19
C7630 VDD.n2160 GND 0.010359f
C7631 VDD.n2161 GND 8.53e-19
C7632 VDD.n2162 GND 0.001706f
C7633 VDD.n2163 GND 9.03e-19
C7634 VDD.n2164 GND 9.03e-19
C7635 VDD.n2165 GND 8.53e-19
C7636 VDD.n2166 GND 0.010359f
C7637 VDD.n2167 GND 9.03e-19
C7638 VDD.n2168 GND 9.03e-19
C7639 VDD.n2169 GND 8.53e-19
C7640 VDD.n2170 GND 0.010359f
C7641 VDD.n2171 GND 0.010359f
C7642 VDD.n2172 GND 0.014703f
C7643 VDD.n2173 GND 0.002444f
C7644 VDD.t454 GND 0.117408f
C7645 VDD.n2174 GND 0.010514f
C7646 VDD.n2175 GND 0.001706f
C7647 VDD.n2176 GND 9.03e-19
C7648 VDD.n2177 GND 0.002444f
C7649 VDD.n2178 GND 8.53e-19
C7650 VDD.n2179 GND 0.001706f
C7651 VDD.n2180 GND 9.03e-19
C7652 VDD.n2181 GND 0.002444f
C7653 VDD.n2182 GND 9.17e-19
C7654 VDD.n2183 GND 0.001706f
C7655 VDD.n2184 GND 0.001706f
C7656 VDD.n2185 GND 0.001706f
C7657 VDD.n2186 GND 0.001706f
C7658 VDD.t336 GND 0.119161f
C7659 VDD.n2187 GND 0.183998f
C7660 VDD.n2188 GND 0.001706f
C7661 VDD.n2189 GND 0.001706f
C7662 VDD.n2190 GND 0.001706f
C7663 VDD.n2191 GND 0.001706f
C7664 VDD.n2192 GND 9.03e-19
C7665 VDD.n2193 GND 0.002444f
C7666 VDD.n2194 GND 8.53e-19
C7667 VDD.n2195 GND 9.03e-19
C7668 VDD.n2196 GND 0.002444f
C7669 VDD.n2197 GND 8.53e-19
C7670 VDD.n2198 GND 9.03e-19
C7671 VDD.n2199 GND 0.001706f
C7672 VDD.n2200 GND 0.001706f
C7673 VDD.n2201 GND 9.03e-19
C7674 VDD.n2202 GND 8.53e-19
C7675 VDD.n2203 GND 0.005502f
C7676 VDD.n2204 GND 9.17e-19
C7677 VDD.n2205 GND 0.001029f
C7678 VDD.n2206 GND 0.001706f
C7679 VDD.n2207 GND 0.001706f
C7680 VDD.n2208 GND 0.001706f
C7681 VDD.n2209 GND 0.001706f
C7682 VDD.n2210 GND 0.001706f
C7683 VDD.n2211 GND 0.001706f
C7684 VDD.n2212 GND 0.001706f
C7685 VDD.t248 GND 0.119161f
C7686 VDD.n2213 GND 0.001706f
C7687 VDD.n2214 GND 0.001706f
C7688 VDD.n2215 GND 0.001706f
C7689 VDD.n2216 GND 0.238321f
C7690 VDD.n2217 GND 0.001706f
C7691 VDD.n2218 GND 0.001706f
C7692 VDD.n2219 GND 0.001706f
C7693 VDD.n2220 GND 0.001706f
C7694 VDD.n2221 GND 0.001706f
C7695 VDD.n2222 GND 0.001706f
C7696 VDD.t538 GND 0.119161f
C7697 VDD.n2223 GND 0.001706f
C7698 VDD.n2224 GND 0.001706f
C7699 VDD.n2225 GND 0.001706f
C7700 VDD.n2226 GND 0.176989f
C7701 VDD.n2227 GND 0.001706f
C7702 VDD.n2228 GND 0.001706f
C7703 VDD.n2229 GND 0.001706f
C7704 VDD.n2230 GND 0.138437f
C7705 VDD.n2231 GND 0.001706f
C7706 VDD.n2232 GND 0.001706f
C7707 VDD.n2233 GND 0.001706f
C7708 VDD.t36 GND 0.119161f
C7709 VDD.n2234 GND 0.001706f
C7710 VDD.n2235 GND 0.001706f
C7711 VDD.n2236 GND 0.001706f
C7712 VDD.n2237 GND 0.215541f
C7713 VDD.n2238 GND 0.001706f
C7714 VDD.n2239 GND 0.003781f
C7715 VDD.n2240 GND 0.003781f
C7716 VDD.t516 GND 0.119161f
C7717 VDD.n2241 GND 0.001706f
C7718 VDD.n2242 GND 0.003781f
C7719 VDD.n2250 GND 0.001706f
C7720 VDD.n2251 GND 0.001706f
C7721 VDD.n2252 GND 0.001706f
C7722 VDD.n2253 GND 0.001706f
C7723 VDD.n2254 GND 0.001706f
C7724 VDD.n2255 GND 0.001706f
C7725 VDD.n2256 GND 0.001706f
C7726 VDD.n2257 GND 0.001706f
C7727 VDD.n2258 GND 0.001706f
C7728 VDD.n2259 GND 0.001706f
C7729 VDD.n2260 GND 0.001706f
C7730 VDD.n2261 GND 0.001706f
C7731 VDD.n2262 GND 0.001706f
C7732 VDD.n2263 GND 0.001706f
C7733 VDD.n2264 GND 0.001706f
C7734 VDD.n2265 GND 0.001706f
C7735 VDD.n2266 GND 0.001706f
C7736 VDD.n2267 GND 0.001706f
C7737 VDD.n2268 GND 0.001706f
C7738 VDD.n2269 GND 0.001706f
C7739 VDD.n2270 GND 0.001706f
C7740 VDD.n2271 GND 0.001706f
C7741 VDD.n2272 GND 0.001706f
C7742 VDD.n2273 GND 0.001706f
C7743 VDD.n2274 GND 0.003781f
C7744 VDD.n2275 GND 0.003795f
C7745 VDD.n2276 GND 0.003795f
C7746 VDD.n2277 GND 0.001706f
C7747 VDD.n2278 GND 0.001706f
C7748 VDD.n2279 GND 0.001706f
C7749 VDD.n2280 GND 0.001706f
C7750 VDD.n2281 GND 0.001706f
C7751 VDD.n2282 GND 0.001706f
C7752 VDD.n2283 GND 0.001706f
C7753 VDD.n2284 GND 0.001706f
C7754 VDD.n2285 GND 0.001706f
C7755 VDD.n2286 GND 0.001706f
C7756 VDD.n2287 GND 0.001706f
C7757 VDD.n2288 GND 0.001706f
C7758 VDD.n2289 GND 0.001706f
C7759 VDD.n2290 GND 0.001706f
C7760 VDD.n2291 GND 0.001706f
C7761 VDD.n2292 GND 0.001706f
C7762 VDD.n2293 GND 0.001706f
C7763 VDD.n2294 GND 0.001706f
C7764 VDD.n2295 GND 0.001706f
C7765 VDD.n2296 GND 0.001706f
C7766 VDD.n2297 GND 0.001706f
C7767 VDD.n2298 GND 0.001706f
C7768 VDD.n2299 GND 0.001706f
C7769 VDD.n2300 GND 0.001706f
C7770 VDD.n2301 GND 0.001706f
C7771 VDD.n2302 GND 0.001706f
C7772 VDD.n2303 GND 0.001706f
C7773 VDD.n2304 GND 0.001706f
C7774 VDD.n2305 GND 0.003795f
C7775 VDD.n2306 GND 0.003795f
C7776 VDD.n2308 GND 0.382015f
C7777 VDD.n2309 GND 0.315425f
C7778 VDD.n2310 GND 0.141941f
C7779 VDD.n2311 GND 0.001706f
C7780 VDD.n2312 GND 0.001706f
C7781 VDD.n2313 GND 0.001706f
C7782 VDD.n2314 GND 0.001706f
C7783 VDD.n2315 GND 0.001706f
C7784 VDD.n2316 GND 0.180493f
C7785 VDD.t126 GND 0.119161f
C7786 VDD.n2317 GND 0.176989f
C7787 VDD.n2318 GND 0.219045f
C7788 VDD.n2319 GND 0.001706f
C7789 VDD.n2320 GND 0.001706f
C7790 VDD.n2321 GND 0.001706f
C7791 VDD.n2322 GND 0.001706f
C7792 VDD.n2323 GND 0.001706f
C7793 VDD.n2324 GND 0.238321f
C7794 VDD.n2325 GND 0.138437f
C7795 VDD.t221 GND 0.119161f
C7796 VDD.n2326 GND 0.219045f
C7797 VDD.n2327 GND 0.001706f
C7798 VDD.n2328 GND 0.001706f
C7799 VDD.n2329 GND 0.001706f
C7800 VDD.n2330 GND 0.001706f
C7801 VDD.n2331 GND 0.001706f
C7802 VDD.n2332 GND 0.180493f
C7803 VDD.n2333 GND 0.215541f
C7804 VDD.t357 GND 0.119161f
C7805 VDD.n2334 GND 0.141941f
C7806 VDD.n2335 GND 0.001706f
C7807 VDD.n2336 GND 0.001706f
C7808 VDD.n2337 GND 0.001706f
C7809 VDD.n2338 GND 0.001706f
C7810 VDD.n2339 GND 0.001706f
C7811 VDD.n2340 GND 0.134932f
C7812 VDD.t501 GND 0.119161f
C7813 VDD.n2341 GND 0.22255f
C7814 VDD.n2342 GND 0.173484f
C7815 VDD.n2343 GND 0.001706f
C7816 VDD.n2344 GND 0.001706f
C7817 VDD.n2345 GND 0.001706f
C7818 VDD.n2346 GND 0.001706f
C7819 VDD.n2347 GND 0.001706f
C7820 VDD.n2348 GND 0.212036f
C7821 VDD.n2349 GND 0.001706f
C7822 VDD.n2350 GND 0.001706f
C7823 VDD.n2351 GND 0.001706f
C7824 VDD.n2352 GND 0.001706f
C7825 VDD.n2353 GND 0.001706f
C7826 VDD.n2354 GND 0.001029f
C7827 VDD.n2355 GND 0.001706f
C7828 VDD.n2356 GND 0.001706f
C7829 VDD.n2357 GND 9.03e-19
C7830 VDD.n2358 GND 8.53e-19
C7831 VDD.n2359 GND 0.005502f
C7832 VDD.n2360 GND 0.002444f
C7833 VDD.n2361 GND 8.53e-19
C7834 VDD.n2362 GND 9.03e-19
C7835 VDD.n2363 GND 0.001706f
C7836 VDD.n2364 GND 0.001706f
C7837 VDD.n2365 GND 9.03e-19
C7838 VDD.n2366 GND 8.53e-19
C7839 VDD.n2367 GND 9.03e-19
C7840 VDD.n2368 GND 8.53e-19
C7841 VDD.n2369 GND 0.002444f
C7842 VDD.n2370 GND 0.002444f
C7843 VDD.n2371 GND 8.53e-19
C7844 VDD.n2372 GND 9.03e-19
C7845 VDD.n2373 GND 8.53e-19
C7846 VDD.n2374 GND 0.001706f
C7847 VDD.n2375 GND 9.03e-19
C7848 VDD.n2376 GND 8.53e-19
C7849 VDD.n2377 GND 0.002444f
C7850 VDD.n2378 GND 0.002375f
C7851 VDD.n2379 GND 8.53e-19
C7852 VDD.n2380 GND 9.03e-19
C7853 VDD.n2381 GND 0.001706f
C7854 VDD.n2382 GND 0.087618f
C7855 VDD.n2383 GND 0.001706f
C7856 VDD.t111 GND 0.117408f
C7857 VDD.n2384 GND 0.054323f
C7858 VDD.n2385 GND 0.001706f
C7859 VDD.n2386 GND 0.001706f
C7860 VDD.n2387 GND 0.001706f
C7861 VDD.n2388 GND 0.001706f
C7862 VDD.n2389 GND 0.001706f
C7863 VDD.n2390 GND 0.001706f
C7864 VDD.n2391 GND 0.001706f
C7865 VDD.n2392 GND 0.001706f
C7866 VDD.n2393 GND 0.001706f
C7867 VDD.n2394 GND 0.001706f
C7868 VDD.n2395 GND 0.001706f
C7869 VDD.t346 GND 0.117408f
C7870 VDD.n2396 GND 0.02979f
C7871 VDD.n2397 GND 0.001706f
C7872 VDD.n2398 GND 0.001706f
C7873 VDD.n2399 GND 0.001706f
C7874 VDD.n2400 GND 0.001706f
C7875 VDD.n2401 GND 0.001706f
C7876 VDD.t271 GND 0.117408f
C7877 VDD.n2402 GND 0.068342f
C7878 VDD.n2403 GND 0.001706f
C7879 VDD.n2404 GND 0.001706f
C7880 VDD.n2405 GND 0.001706f
C7881 VDD.n2406 GND 0.001706f
C7882 VDD.n2407 GND 0.001706f
C7883 VDD.n2408 GND 0.001706f
C7884 VDD.n2409 GND 0.001706f
C7885 VDD.n2410 GND 0.001706f
C7886 VDD.n2411 GND 0.001706f
C7887 VDD.n2412 GND 0.001706f
C7888 VDD.n2413 GND 0.001706f
C7889 VDD.n2414 GND 0.001706f
C7890 VDD.n2415 GND 0.001706f
C7891 VDD.n2416 GND 0.001706f
C7892 VDD.n2417 GND 0.001706f
C7893 VDD.n2418 GND 0.001706f
C7894 VDD.n2419 GND 0.001706f
C7895 VDD.n2420 GND 0.001706f
C7896 VDD.n2421 GND 0.001706f
C7897 VDD.n2422 GND 0.001706f
C7898 VDD.n2423 GND 0.001706f
C7899 VDD.n2424 GND 0.001706f
C7900 VDD.n2425 GND 0.001706f
C7901 VDD.n2426 GND 0.001706f
C7902 VDD.n2427 GND 0.001706f
C7903 VDD.n2428 GND 0.001706f
C7904 VDD.n2429 GND 0.001706f
C7905 VDD.n2430 GND 0.001706f
C7906 VDD.n2431 GND 0.001706f
C7907 VDD.n2432 GND 0.003727f
C7908 VDD.n2433 GND 0.003723f
C7909 VDD.n2434 GND 0.001706f
C7910 VDD.n2435 GND 0.001706f
C7911 VDD.t189 GND 0.117408f
C7912 VDD.n2436 GND 0.106894f
C7913 VDD.n2437 GND 0.001706f
C7914 VDD.n2438 GND 0.001706f
C7915 VDD.n2439 GND 0.003723f
C7916 VDD.n2440 GND 0.003727f
C7917 VDD.n2441 GND 0.003727f
C7918 VDD.n2442 GND 0.001706f
C7919 VDD.n2443 GND 0.001706f
C7920 VDD.n2444 GND 0.001706f
C7921 VDD.n2445 GND 0.001706f
C7922 VDD.n2446 GND 0.001706f
C7923 VDD.n2447 GND 0.001706f
C7924 VDD.n2448 GND 0.001706f
C7925 VDD.n2449 GND 0.001706f
C7926 VDD.n2450 GND 0.001706f
C7927 VDD.n2451 GND 0.001706f
C7928 VDD.n2452 GND 0.001706f
C7929 VDD.n2453 GND 0.001706f
C7930 VDD.n2454 GND 0.001706f
C7931 VDD.n2455 GND 0.001706f
C7932 VDD.n2456 GND 0.001706f
C7933 VDD.n2457 GND 0.001706f
C7934 VDD.n2458 GND 0.001706f
C7935 VDD.n2459 GND 0.001706f
C7936 VDD.n2460 GND 0.001706f
C7937 VDD.n2461 GND 0.001706f
C7938 VDD.n2462 GND 0.001706f
C7939 VDD.n2463 GND 0.001706f
C7940 VDD.n2464 GND 0.001706f
C7941 VDD.n2465 GND 0.001706f
C7942 VDD.n2466 GND 0.001706f
C7943 VDD.n2467 GND 0.001706f
C7944 VDD.n2468 GND 0.001706f
C7945 VDD.n2469 GND 0.001706f
C7946 VDD.n2470 GND 0.001706f
C7947 VDD.n2472 GND 0.119161f
C7948 VDD.n2474 GND 0.001706f
C7949 VDD.n2475 GND 0.001706f
C7950 VDD.n2476 GND 0.003727f
C7951 VDD.n2477 GND 0.003723f
C7952 VDD.n2478 GND 0.003723f
C7953 VDD.n2479 GND 0.119161f
C7954 VDD.n2480 GND 0.003723f
C7955 VDD.n2481 GND 0.003723f
C7956 VDD.n2482 GND 0.001706f
C7957 VDD.n2483 GND 0.001706f
C7958 VDD.n2484 GND 0.001706f
C7959 VDD.n2485 GND 0.08937f
C7960 VDD.n2486 GND 0.001706f
C7961 VDD.n2487 GND 0.001706f
C7962 VDD.n2488 GND 0.001706f
C7963 VDD.n2489 GND 0.001706f
C7964 VDD.n2490 GND 0.001706f
C7965 VDD.n2491 GND 0.050818f
C7966 VDD.n2492 GND 0.001706f
C7967 VDD.n2493 GND 0.001706f
C7968 VDD.n2494 GND 0.001706f
C7969 VDD.n2495 GND 0.001706f
C7970 VDD.n2496 GND 0.001706f
C7971 VDD.n2497 GND 0.012266f
C7972 VDD.n2498 GND 0.119161f
C7973 VDD.n2499 GND 0.001706f
C7974 VDD.n2500 GND 9.03e-19
C7975 VDD.n2501 GND 8.53e-19
C7976 VDD.n2502 GND 0.002444f
C7977 VDD.n2503 GND 0.002444f
C7978 VDD.n2504 GND 8.53e-19
C7979 VDD.n2505 GND 9.03e-19
C7980 VDD.n2506 GND 0.001706f
C7981 VDD.n2507 GND 0.028038f
C7982 VDD.t360 GND 0.117408f
C7983 VDD.n2508 GND 0.092875f
C7984 VDD.n2509 GND 0.001706f
C7985 VDD.n2510 GND 0.00133f
C7986 VDD.n2511 GND 0.003632f
C7987 VDD.n2512 GND 0.008749f
C7988 VDD.n2513 GND 0.001706f
C7989 VDD.n2514 GND 0.071847f
C7990 VDD.n2515 GND 0.001706f
C7991 VDD.n2516 GND 0.001706f
C7992 VDD.n2517 GND 0.001706f
C7993 VDD.n2518 GND 0.001129f
C7994 VDD.n2519 GND 0.001706f
C7995 VDD.n2520 GND 0.033295f
C7996 VDD.n2521 GND 0.105142f
C7997 VDD.n2522 GND 0.001706f
C7998 VDD.n2523 GND 9.03e-19
C7999 VDD.n2524 GND 8.53e-19
C8000 VDD.n2525 GND 0.002444f
C8001 VDD.n2526 GND 0.002316f
C8002 VDD.n2527 GND 8.53e-19
C8003 VDD.n2528 GND 9.03e-19
C8004 VDD.n2529 GND 0.001706f
C8005 VDD.n2530 GND 0.007009f
C8006 VDD.n2531 GND 0.001706f
C8007 VDD.n2532 GND 9.03e-19
C8008 VDD.n2533 GND 8.53e-19
C8009 VDD.n2534 GND 0.010359f
C8010 VDD.n2535 GND 0.010359f
C8011 VDD.n2536 GND 8.53e-19
C8012 VDD.n2537 GND 9.03e-19
C8013 VDD.n2538 GND 0.001706f
C8014 VDD.n2539 GND 0.09638f
C8015 VDD.n2540 GND 0.045561f
C8016 VDD.n2541 GND 0.001706f
C8017 VDD.n2542 GND 8.78e-19
C8018 VDD.n2543 GND 8.53e-19
C8019 VDD.n2544 GND 0.01746f
C8020 VDD.n2545 GND 0.102225f
C8021 VDD.n2546 GND 0.601507f
C8022 VDD.n2547 GND 0.102225f
C8023 VDD.n2548 GND 0.014122f
C8024 VDD.n2549 GND 8.53e-19
C8025 VDD.n2550 GND 8.78e-19
C8026 VDD.n2551 GND 8.78e-19
C8027 VDD.n2552 GND 0.001706f
C8028 VDD.n2553 GND 0.115656f
C8029 VDD.n2554 GND 0.001706f
C8030 VDD.n2555 GND 8.78e-19
C8031 VDD.n2556 GND 8.53e-19
C8032 VDD.n2557 GND 0.010359f
C8033 VDD.n2558 GND 0.010359f
C8034 VDD.n2559 GND 8.53e-19
C8035 VDD.n2560 GND 9.03e-19
C8036 VDD.n2561 GND 0.001706f
C8037 VDD.n2562 GND 0.005257f
C8038 VDD.n2563 GND 0.001706f
C8039 VDD.n2564 GND 0.008303f
C8040 VDD.n2565 GND 0.072346f
C8041 VDD.n2566 GND 1.79982f
C8042 VDD.n2567 GND 0.073151f
C8043 VDD.n2568 GND 0.002244f
C8044 VDD.t333 GND 0.010699f
C8045 VDD.t377 GND 0.010699f
C8046 VDD.n2569 GND 0.022031f
C8047 VDD.n2570 GND 9.03e-19
C8048 VDD.n2571 GND 0.001516f
C8049 VDD.n2572 GND 8.53e-19
C8050 VDD.n2573 GND 0.002454f
C8051 VDD.n2574 GND 0.002363f
C8052 VDD.n2575 GND 8.53e-19
C8053 VDD.n2576 GND 9.03e-19
C8054 VDD.n2577 GND 0.001972f
C8055 VDD.n2578 GND 0.001783f
C8056 VDD.n2579 GND 0.044032f
C8057 VDD.n2580 GND 2.75612f
C8058 VDD.n2581 GND 26.0199f
C8059 VDD.n2582 GND 7.64969f
C8060 VDD.n2585 GND 1.88886f
C8061 VDD.n2586 GND 1.88886f
C8062 VDD.n2587 GND 1.88886f
C8063 VDD.n2589 GND 1.88886f
C8064 VDD.n2592 GND 2.36108f
C8065 VDD.n2593 GND 2.36108f
C8066 VDD.n2596 GND 1.88886f
C8067 VDD.n2597 GND 1.77081f
C8068 VDD.n2599 GND 0.335437f
C8069 VDD.n2600 GND 0.005467f
C8070 VDD.n2601 GND 0.002367f
C8071 VDD.n2602 GND 8.53e-19
C8072 VDD.n2603 GND 0.00291f
C8073 VDD.n2604 GND 9.03e-19
C8074 VDD.n2605 GND 0.007088f
C8075 VDD.t345 GND 0.00545f
C8076 VDD.n2606 GND 0.002183f
C8077 VDD.n2607 GND 0.001115f
C8078 VDD.n2608 GND 8.53e-19
C8079 VDD.n2609 GND 0.041407f
C8080 VDD.n2610 GND 0.002444f
C8081 VDD.n2611 GND 8.53e-19
C8082 VDD.n2612 GND 9.03e-19
C8083 VDD.n2613 GND 0.00291f
C8084 VDD.n2614 GND 0.006447f
C8085 VDD.n2615 GND 9.03e-19
C8086 VDD.n2616 GND 0.00116f
C8087 VDD.n2617 GND 0.002806f
C8088 VDD.n2618 GND 0.018731f
C8089 VDD.n2619 GND 0.12073f
C8090 VDD.n2620 GND 0.018612f
C8091 VDD.n2621 GND 0.011119f
C8092 VDD.n2622 GND 0.001062f
C8093 VDD.n2623 GND 0.001706f
C8094 VDD.n2625 GND 0.247293f
C8095 VDD.n2626 GND 0.001706f
C8096 VDD.n2627 GND 0.001706f
C8097 VDD.n2629 GND 0.003712f
C8098 VDD.n2630 GND 0.001706f
C8099 VDD.n2631 GND 0.001706f
C8100 VDD.n2632 GND 0.188724f
C8101 VDD.n2633 GND 0.001706f
C8102 VDD.n2634 GND 0.074839f
C8103 VDD.n2635 GND 0.001706f
C8104 VDD.n2636 GND 0.003712f
C8105 VDD.n2637 GND 0.001706f
C8106 VDD.n2638 GND 0.003712f
C8107 VDD.n2639 GND 0.001706f
C8108 VDD.n2640 GND 0.001706f
C8109 VDD.t75 GND 0.073754f
C8110 VDD.n2641 GND 0.001706f
C8111 VDD.n2642 GND 0.001706f
C8112 VDD.n2643 GND 0.147508f
C8113 VDD.n2644 GND 0.001706f
C8114 VDD.n2645 GND 0.001706f
C8115 VDD.n2646 GND 0.003714f
C8116 VDD.n2647 GND 0.001706f
C8117 VDD.n2648 GND 0.001706f
C8118 VDD.n2649 GND 0.001706f
C8119 VDD.n2651 GND 0.001706f
C8120 VDD.n2652 GND 0.001003f
C8121 VDD.n2654 GND 0.001706f
C8122 VDD.n2655 GND 0.001706f
C8123 VDD.n2656 GND 0.001062f
C8124 VDD.n2657 GND 0.001003f
C8125 VDD.n2658 GND 0.001149f
C8126 VDD.n2659 GND 0.001704f
C8127 VDD.n2660 GND 0.001706f
C8128 VDD.n2662 GND 0.001706f
C8129 VDD.n2663 GND 0.001706f
C8130 VDD.n2664 GND 0.001706f
C8131 VDD.n2665 GND 0.001706f
C8132 VDD.n2666 GND 0.001706f
C8133 VDD.n2667 GND 0.001706f
C8134 VDD.n2669 GND 0.001706f
C8135 VDD.n2670 GND 0.003714f
C8136 VDD.n2671 GND 0.003712f
C8137 VDD.n2672 GND 0.003712f
C8138 VDD.n2673 GND 0.001706f
C8139 VDD.n2674 GND 0.001706f
C8140 VDD.n2675 GND 0.001706f
C8141 VDD.n2676 GND 0.001706f
C8142 VDD.n2677 GND 0.001706f
C8143 VDD.n2678 GND 0.001706f
C8144 VDD.t67 GND 0.073754f
C8145 VDD.n2679 GND 0.001706f
C8146 VDD.n2680 GND 0.001706f
C8147 VDD.n2681 GND 0.001706f
C8148 VDD.n2682 GND 0.087854f
C8149 VDD.n2683 GND 0.001706f
C8150 VDD.n2684 GND 0.001706f
C8151 VDD.n2685 GND 0.147508f
C8152 VDD.n2686 GND 0.001706f
C8153 VDD.n2687 GND 0.001706f
C8154 VDD.n2688 GND 0.001706f
C8155 VDD.n2689 GND 0.001706f
C8156 VDD.n2690 GND 0.001706f
C8157 VDD.t503 GND 0.073754f
C8158 VDD.n2691 GND 0.001706f
C8159 VDD.n2692 GND 0.001706f
C8160 VDD.n2693 GND 0.001706f
C8161 VDD.n2694 GND 0.103039f
C8162 VDD.n2695 GND 0.001706f
C8163 VDD.n2696 GND 0.001706f
C8164 VDD.n2697 GND 0.147508f
C8165 VDD.n2698 GND 0.001706f
C8166 VDD.n2699 GND 0.001706f
C8167 VDD.n2700 GND 0.001706f
C8168 VDD.n2701 GND 0.001706f
C8169 VDD.n2702 GND 0.001706f
C8170 VDD.t505 GND 0.073754f
C8171 VDD.n2703 GND 0.001706f
C8172 VDD.n2704 GND 0.001706f
C8173 VDD.n2705 GND 0.001706f
C8174 VDD.n2706 GND 0.118224f
C8175 VDD.n2707 GND 0.001706f
C8176 VDD.n2708 GND 0.001706f
C8177 VDD.n2709 GND 0.147508f
C8178 VDD.n2710 GND 0.001706f
C8179 VDD.n2711 GND 0.001706f
C8180 VDD.n2712 GND 0.001706f
C8181 VDD.n2713 GND 0.001706f
C8182 VDD.n2714 GND 0.001706f
C8183 VDD.t63 GND 0.073754f
C8184 VDD.n2715 GND 0.001706f
C8185 VDD.n2716 GND 0.001706f
C8186 VDD.n2717 GND 0.001706f
C8187 VDD.n2718 GND 0.133408f
C8188 VDD.n2719 GND 0.001706f
C8189 VDD.n2720 GND 0.001706f
C8190 VDD.n2721 GND 0.146424f
C8191 VDD.n2722 GND 0.001706f
C8192 VDD.n2723 GND 0.001706f
C8193 VDD.n2724 GND 0.001706f
C8194 VDD.t73 GND 0.073754f
C8195 VDD.n2725 GND 0.001706f
C8196 VDD.n2726 GND 0.001706f
C8197 VDD.n2727 GND 0.147508f
C8198 VDD.n2728 GND 0.001706f
C8199 VDD.n2729 GND 0.003714f
C8200 VDD.n2730 GND 0.003714f
C8201 VDD.n2731 GND 0.003712f
C8202 VDD.n2732 GND 0.003712f
C8203 VDD.n2733 GND 0.229939f
C8204 VDD.n2734 GND 0.003714f
C8205 VDD.n2735 GND 0.001706f
C8206 VDD.n2736 GND 0.001706f
C8207 VDD.n2737 GND 0.001704f
C8208 VDD.n2738 GND 0.001706f
C8209 VDD.n2739 GND 0.001062f
C8210 VDD.t506 GND 0.010699f
C8211 VDD.t69 GND 0.010699f
C8212 VDD.n2740 GND 0.032273f
C8213 VDD.n2741 GND 0.107301f
C8214 VDD.n2742 GND 0.005784f
C8215 VDD.n2743 GND 0.005969f
C8216 VDD.n2744 GND 8.53e-19
C8217 VDD.n2745 GND 0.002183f
C8218 VDD.n2746 GND 8.78e-19
C8219 VDD.n2747 GND 0.004516f
C8220 VDD.n2748 GND 0.004516f
C8221 VDD.n2749 GND 0.001062f
C8222 VDD.t74 GND 0.001455f
C8223 VDD.n2750 GND 0.005656f
C8224 VDD.n2751 GND 8.78e-19
C8225 VDD.n2752 GND 0.001115f
C8226 VDD.n2753 GND 0.00636f
C8227 VDD.n2754 GND 0.041968f
C8228 VDD.n2755 GND 0.001022f
C8229 VDD.n2756 GND 0.001706f
C8230 VDD.n2757 GND 0.001706f
C8231 VDD.n2758 GND 0.001706f
C8232 VDD.n2760 GND 0.001706f
C8233 VDD.n2761 GND 0.001706f
C8234 VDD.n2762 GND 0.001706f
C8235 VDD.n2763 GND 0.001706f
C8236 VDD.n2764 GND 0.001706f
C8237 VDD.n2766 GND 0.001706f
C8238 VDD.n2768 GND 0.001706f
C8239 VDD.n2769 GND 0.001706f
C8240 VDD.n2770 GND 0.00173f
C8241 VDD.n2771 GND 0.002023f
C8242 VDD.n2772 GND 0.001706f
C8243 VDD.n2774 GND 0.001706f
C8244 VDD.n2775 GND 0.001706f
C8245 VDD.n2776 GND 0.001706f
C8246 VDD.n2777 GND 0.001706f
C8247 VDD.n2778 GND 0.003714f
C8248 VDD.n2779 GND 0.001706f
C8249 VDD.n2780 GND 0.001706f
C8250 VDD.n2781 GND 0.001706f
C8251 VDD.n2782 GND 0.001062f
C8252 VDD.n2783 GND 0.004516f
C8253 VDD.n2784 GND 0.005656f
C8254 VDD.n2785 GND 8.53e-19
C8255 VDD.n2786 GND 0.006434f
C8256 VDD.n2787 GND 9.03e-19
C8257 VDD.t68 GND 0.010699f
C8258 VDD.t504 GND 0.010699f
C8259 VDD.n2788 GND 0.032273f
C8260 VDD.n2789 GND 0.229486f
C8261 VDD.n2790 GND 0.586149f
C8262 VDD.n2791 GND 0.107744f
C8263 VDD.n2792 GND 0.030806f
C8264 VDD.n2793 GND 0.025832f
C8265 VDD.n2794 GND 0.005784f
C8266 VDD.n2795 GND 0.001162f
C8267 VDD.n2796 GND 0.0023f
C8268 VDD.n2797 GND 0.004516f
C8269 VDD.n2798 GND 0.00173f
C8270 VDD.n2799 GND 0.001706f
C8271 VDD.n2800 GND 0.001706f
C8272 VDD.n2801 GND 0.001706f
C8273 VDD.n2802 GND 0.003714f
C8274 VDD.n2803 GND 0.003714f
C8275 VDD.n2805 GND 0.001706f
C8276 VDD.n2807 GND 0.001706f
C8277 VDD.n2808 GND 0.001706f
C8278 VDD.n2809 GND 0.001706f
C8279 VDD.n2810 GND 0.001706f
C8280 VDD.n2811 GND 0.001706f
C8281 VDD.n2813 GND 0.001706f
C8282 VDD.n2814 GND 0.001706f
C8283 VDD.n2815 GND 0.001706f
C8284 VDD.n2816 GND 0.004516f
C8285 VDD.n2817 GND 0.001003f
C8286 VDD.n2819 GND 0.001706f
C8287 VDD.n2821 GND 0.001706f
C8288 VDD.n2822 GND 0.001062f
C8289 VDD.n2823 GND 0.002023f
C8290 VDD.n2824 GND 0.004516f
C8291 VDD.n2825 GND 0.005969f
C8292 VDD.n2826 GND 8.53e-19
C8293 VDD.n2827 GND 9.03e-19
C8294 VDD.n2828 GND 0.00291f
C8295 VDD.t76 GND 0.001455f
C8296 VDD.n2829 GND 0.002183f
C8297 VDD.n2830 GND 8.78e-19
C8298 VDD.n2831 GND 8.78e-19
C8299 VDD.n2832 GND 0.001115f
C8300 VDD.n2833 GND 0.00636f
C8301 VDD.n2834 GND 0.041968f
C8302 VDD.n2835 GND 0.001022f
C8303 VDD.n2836 GND 0.001645f
C8304 VDD.n2837 GND 0.001706f
C8305 VDD.n2838 GND 0.001706f
C8306 VDD.n2840 GND 0.001706f
C8307 VDD.n2842 GND 0.001706f
C8308 VDD.n2843 GND 0.001706f
C8309 VDD.n2844 GND 0.001706f
C8310 VDD.n2845 GND 0.001706f
C8311 VDD.n2846 GND 0.001706f
C8312 VDD.n2848 GND 0.003714f
C8313 VDD.n2849 GND 0.003712f
C8314 VDD.n2850 GND 0.003712f
C8315 VDD.n2851 GND 0.001706f
C8316 VDD.n2852 GND 0.001706f
C8317 VDD.n2853 GND 0.001706f
C8318 VDD.n2854 GND 0.001706f
C8319 VDD.n2855 GND 0.001706f
C8320 VDD.n2856 GND 0.001706f
C8321 VDD.n2857 GND 0.001706f
C8322 VDD.n2858 GND 0.001706f
C8323 VDD.n2859 GND 0.001706f
C8324 VDD.n2860 GND 0.001706f
C8325 VDD.n2861 GND 0.001706f
C8326 VDD.n2862 GND 0.001706f
C8327 VDD.n2863 GND 0.001706f
C8328 VDD.n2864 GND 0.001706f
C8329 VDD.n2865 GND 0.001706f
C8330 VDD.n2866 GND 0.001706f
C8331 VDD.n2867 GND 0.001706f
C8332 VDD.n2868 GND 0.001706f
C8333 VDD.n2869 GND 0.001706f
C8334 VDD.n2870 GND 0.001706f
C8335 VDD.n2871 GND 0.001706f
C8336 VDD.n2872 GND 0.001706f
C8337 VDD.n2873 GND 0.001706f
C8338 VDD.n2874 GND 0.001706f
C8339 VDD.n2875 GND 0.001706f
C8340 VDD.n2876 GND 0.001706f
C8341 VDD.n2877 GND 0.001706f
C8342 VDD.n2878 GND 0.001706f
C8343 VDD.n2879 GND 0.001706f
C8344 VDD.n2880 GND 0.001706f
C8345 VDD.n2881 GND 0.001706f
C8346 VDD.n2882 GND 0.001706f
C8347 VDD.n2883 GND 0.001706f
C8348 VDD.n2884 GND 0.003712f
C8349 VDD.n2886 GND 0.003714f
C8350 VDD.n2887 GND 0.003714f
C8351 VDD.n2888 GND 0.001706f
C8352 VDD.n2889 GND 0.001706f
C8353 VDD.n2890 GND 0.001706f
C8354 VDD.n2892 GND 0.001706f
C8355 VDD.n2894 GND 0.001706f
C8356 VDD.n2895 GND 0.001706f
C8357 VDD.n2896 GND 0.001706f
C8358 VDD.n2897 GND 0.001645f
C8359 VDD.n2898 GND 0.001706f
C8360 VDD.n2900 GND 0.001706f
C8361 VDD.n2901 GND 0.001062f
C8362 VDD.n2902 GND 0.001003f
C8363 VDD.n2903 GND 0.004516f
C8364 VDD.n2904 GND 0.004516f
C8365 VDD.n2905 GND 8.53e-19
C8366 VDD.n2906 GND 9.03e-19
C8367 VDD.n2907 GND 0.00291f
C8368 VDD.n2908 GND 0.006434f
C8369 VDD.n2909 GND 9.03e-19
C8370 VDD.n2910 GND 0.001162f
C8371 VDD.n2911 GND 0.0023f
C8372 VDD.n2912 GND 0.025832f
C8373 VDD.n2913 GND 0.033011f
C8374 VDD.n2914 GND 0.172693f
C8375 VDD.t549 GND 0.010699f
C8376 VDD.t715 GND 0.010699f
C8377 VDD.n2915 GND 0.032325f
C8378 VDD.n2916 GND 0.102342f
C8379 VDD.t544 GND 0.010699f
C8380 VDD.t64 GND 0.010699f
C8381 VDD.n2917 GND 0.032325f
C8382 VDD.n2918 GND 0.102988f
C8383 VDD.n2919 GND 0.005467f
C8384 VDD.n2920 GND 0.002367f
C8385 VDD.n2921 GND 8.53e-19
C8386 VDD.n2922 GND 0.00291f
C8387 VDD.n2923 GND 9.03e-19
C8388 VDD.n2924 GND 0.007088f
C8389 VDD.t533 GND 0.00545f
C8390 VDD.n2925 GND 0.002183f
C8391 VDD.n2926 GND 0.001115f
C8392 VDD.n2927 GND 8.53e-19
C8393 VDD.n2928 GND 0.041407f
C8394 VDD.n2929 GND 0.002444f
C8395 VDD.n2930 GND 8.53e-19
C8396 VDD.n2931 GND 9.03e-19
C8397 VDD.n2932 GND 0.00291f
C8398 VDD.n2933 GND 0.006447f
C8399 VDD.n2934 GND 9.03e-19
C8400 VDD.n2935 GND 0.00116f
C8401 VDD.n2936 GND 0.002806f
C8402 VDD.n2937 GND 0.018731f
C8403 VDD.n2938 GND 0.052956f
C8404 VDD.n2939 GND 0.192513f
C8405 VDD.n2940 GND 0.031168f
C8406 VDD.n2941 GND 0.017532f
C8407 VDD.n2942 GND 0.00102f
C8408 VDD.n2944 GND 0.001706f
C8409 VDD.n2945 GND 0.001706f
C8410 VDD.n2946 GND 0.001706f
C8411 VDD.n2947 GND 0.001706f
C8412 VDD.n2948 GND 0.001706f
C8413 VDD.n2949 GND 0.001706f
C8414 VDD.n2950 GND 0.001706f
C8415 VDD.n2951 GND 0.001706f
C8416 VDD.n2952 GND 0.001706f
C8417 VDD.n2953 GND 0.001706f
C8418 VDD.n2954 GND 0.001706f
C8419 VDD.n2955 GND 0.001706f
C8420 VDD.n2956 GND 0.001706f
C8421 VDD.n2957 GND 0.001706f
C8422 VDD.n2958 GND 0.001706f
C8423 VDD.n2959 GND 0.001706f
C8424 VDD.n2960 GND 0.001706f
C8425 VDD.n2961 GND 0.001706f
C8426 VDD.n2962 GND 0.001706f
C8427 VDD.n2963 GND 0.001706f
C8428 VDD.n2964 GND 0.001706f
C8429 VDD.n2965 GND 0.001706f
C8430 VDD.n2966 GND 0.001706f
C8431 VDD.n2967 GND 0.001706f
C8432 VDD.n2968 GND 0.001706f
C8433 VDD.n2969 GND 0.001706f
C8434 VDD.n2970 GND 0.001706f
C8435 VDD.n2971 GND 0.001706f
C8436 VDD.n2972 GND 0.001706f
C8437 VDD.n2973 GND 0.001706f
C8438 VDD.n2974 GND 0.001706f
C8439 VDD.n2975 GND 0.001706f
C8440 VDD.n2976 GND 0.003712f
C8441 VDD.n2977 GND 0.003714f
C8442 VDD.n2978 GND 0.003714f
C8443 VDD.n2980 GND 0.001706f
C8444 VDD.n2981 GND 0.001706f
C8445 VDD.n2982 GND 0.001706f
C8446 VDD.n2983 GND 0.001706f
C8447 VDD.n2984 GND 0.001706f
C8448 VDD.n2986 GND 0.001706f
C8449 VDD.n2987 GND 0.001706f
C8450 VDD.n2988 GND 0.001706f
C8451 VDD.n2989 GND 0.001547f
C8452 VDD.n2990 GND 0.001706f
C8453 VDD.n2992 GND 0.001706f
C8454 VDD.n2993 GND 0.001062f
C8455 VDD.n2994 GND 0.001003f
C8456 VDD.n2995 GND 0.011119f
C8457 VDD.n2996 GND 0.018664f
C8458 VDD.n2997 GND 0.001003f
C8459 VDD.n2998 GND 0.001149f
C8460 VDD.n2999 GND 0.001706f
C8461 VDD.n3001 GND 0.001706f
C8462 VDD.n3003 GND 0.001706f
C8463 VDD.n3004 GND 0.001706f
C8464 VDD.n3005 GND 0.001706f
C8465 VDD.n3006 GND 0.001706f
C8466 VDD.n3007 GND 0.001706f
C8467 VDD.n3009 GND 0.001706f
C8468 VDD.n3011 GND 0.001706f
C8469 VDD.n3012 GND 0.001706f
C8470 VDD.n3013 GND 0.003714f
C8471 VDD.n3014 GND 0.003712f
C8472 VDD.n3015 GND 0.003712f
C8473 VDD.n3016 GND 0.188724f
C8474 VDD.n3017 GND 0.003712f
C8475 VDD.n3018 GND 0.003712f
C8476 VDD.n3019 GND 0.001706f
C8477 VDD.n3020 GND 0.001706f
C8478 VDD.n3021 GND 0.001706f
C8479 VDD.n3022 GND 0.074839f
C8480 VDD.n3023 GND 0.001706f
C8481 VDD.n3024 GND 0.001706f
C8482 VDD.n3025 GND 0.001706f
C8483 VDD.n3026 GND 0.001706f
C8484 VDD.n3027 GND 0.001706f
C8485 VDD.n3028 GND 0.147508f
C8486 VDD.n3029 GND 0.001706f
C8487 VDD.n3030 GND 0.001706f
C8488 VDD.n3031 GND 0.001706f
C8489 VDD.n3032 GND 0.001706f
C8490 VDD.n3033 GND 0.001706f
C8491 VDD.n3034 GND 0.087854f
C8492 VDD.n3035 GND 0.001706f
C8493 VDD.n3036 GND 0.001706f
C8494 VDD.n3037 GND 0.001706f
C8495 VDD.n3038 GND 0.001706f
C8496 VDD.n3039 GND 0.001706f
C8497 VDD.n3040 GND 0.147508f
C8498 VDD.n3041 GND 0.001706f
C8499 VDD.n3042 GND 0.001706f
C8500 VDD.n3043 GND 0.001706f
C8501 VDD.n3044 GND 0.001706f
C8502 VDD.n3045 GND 0.001706f
C8503 VDD.n3046 GND 0.103039f
C8504 VDD.n3047 GND 0.001706f
C8505 VDD.n3048 GND 0.001706f
C8506 VDD.n3049 GND 0.001706f
C8507 VDD.n3050 GND 0.001706f
C8508 VDD.n3051 GND 0.001706f
C8509 VDD.n3052 GND 0.147508f
C8510 VDD.n3053 GND 0.001706f
C8511 VDD.n3054 GND 0.001706f
C8512 VDD.n3055 GND 0.001706f
C8513 VDD.n3056 GND 0.001706f
C8514 VDD.n3057 GND 0.001706f
C8515 VDD.n3058 GND 0.118224f
C8516 VDD.n3059 GND 0.001706f
C8517 VDD.n3060 GND 0.001706f
C8518 VDD.n3061 GND 0.001706f
C8519 VDD.n3062 GND 0.001706f
C8520 VDD.n3063 GND 0.001706f
C8521 VDD.n3064 GND 0.147508f
C8522 VDD.n3065 GND 0.001706f
C8523 VDD.n3066 GND 0.001706f
C8524 VDD.n3067 GND 0.001706f
C8525 VDD.n3068 GND 0.001706f
C8526 VDD.n3069 GND 0.001706f
C8527 VDD.n3070 GND 0.133408f
C8528 VDD.n3071 GND 0.001706f
C8529 VDD.n3072 GND 0.001706f
C8530 VDD.n3073 GND 0.001706f
C8531 VDD.n3074 GND 0.001706f
C8532 VDD.n3075 GND 0.001706f
C8533 VDD.n3076 GND 0.146424f
C8534 VDD.n3077 GND 0.001706f
C8535 VDD.n3078 GND 0.001706f
C8536 VDD.n3079 GND 0.001706f
C8537 VDD.n3080 GND 0.001706f
C8538 VDD.n3081 GND 0.001706f
C8539 VDD.n3082 GND 0.147508f
C8540 VDD.n3083 GND 0.001706f
C8541 VDD.n3084 GND 0.001706f
C8542 VDD.n3085 GND 0.003712f
C8543 VDD.n3086 GND 0.003714f
C8544 VDD.n3087 GND 0.003714f
C8545 VDD.n3089 GND 0.001706f
C8546 VDD.n3090 GND 0.001706f
C8547 VDD.n3091 GND 0.001706f
C8548 VDD.n3092 GND 0.001706f
C8549 VDD.n3093 GND 0.001706f
C8550 VDD.n3094 GND 0.001706f
C8551 VDD.n3096 GND 0.001706f
C8552 VDD.n3097 GND 0.001706f
C8553 VDD.n3098 GND 0.001547f
C8554 VDD.n3099 GND 0.00102f
C8555 VDD.n3100 GND 0.017479f
C8556 VDD.n3101 GND 3.28559f
C8557 VDD.n3102 GND 21.755f
C8558 VDD.n3103 GND 0.007272f
C8559 VDD.n3104 GND 0.007272f
C8560 VDD.n3105 GND 0.002244f
C8561 VDD.t430 GND 0.010699f
C8562 VDD.t422 GND 0.010699f
C8563 VDD.n3106 GND 0.022031f
C8564 VDD.n3107 GND 9.03e-19
C8565 VDD.n3108 GND 0.001516f
C8566 VDD.n3109 GND 8.53e-19
C8567 VDD.n3110 GND 0.002454f
C8568 VDD.n3111 GND 0.002363f
C8569 VDD.n3112 GND 8.53e-19
C8570 VDD.n3113 GND 9.03e-19
C8571 VDD.n3114 GND 0.001972f
C8572 VDD.n3115 GND 0.001783f
C8573 VDD.n3116 GND 0.044032f
C8574 VDD.n3117 GND 0.05786f
C8575 VDD.n3118 GND 0.072213f
C8576 VDD.n3119 GND 0.007272f
C8577 VDD.n3120 GND 0.007272f
C8578 VDD.n3121 GND 0.002244f
C8579 VDD.n3122 GND 0.002384f
C8580 VDD.n3123 GND 9.03e-19
C8581 VDD.n3124 GND 8.53e-19
C8582 VDD.n3125 GND 0.005733f
C8583 VDD.n3126 GND 9.03e-19
C8584 VDD.n3127 GND 0.00263f
C8585 VDD.n3128 GND 8.53e-19
C8586 VDD.n3129 GND 0.002454f
C8587 VDD.n3130 GND 0.002363f
C8588 VDD.n3131 GND 8.53e-19
C8589 VDD.n3132 GND 8.53e-19
C8590 VDD.n3133 GND 9.03e-19
C8591 VDD.n3134 GND 0.00291f
C8592 VDD.n3135 GND 0.00291f
C8593 VDD.n3136 GND 0.002183f
C8594 VDD.n3137 GND 0.001115f
C8595 VDD.t449 GND 0.00545f
C8596 VDD.n3138 GND 0.007088f
C8597 VDD.n3139 GND 0.041407f
C8598 VDD.n3140 GND 8.53e-19
C8599 VDD.n3141 GND 9.03e-19
C8600 VDD.n3142 GND 0.00291f
C8601 VDD.n3143 GND 0.00291f
C8602 VDD.n3144 GND 9.03e-19
C8603 VDD.n3145 GND 8.53e-19
C8604 VDD.n3146 GND 0.002437f
C8605 VDD.n3147 GND 0.004543f
C8606 VDD.n3148 GND 0.047272f
C8607 VDD.n3149 GND 0.002244f
C8608 VDD.t425 GND 0.010699f
C8609 VDD.t416 GND 0.010699f
C8610 VDD.n3150 GND 0.022031f
C8611 VDD.n3151 GND 9.03e-19
C8612 VDD.n3152 GND 0.001516f
C8613 VDD.n3153 GND 8.53e-19
C8614 VDD.n3154 GND 0.002454f
C8615 VDD.n3155 GND 0.002363f
C8616 VDD.n3156 GND 8.53e-19
C8617 VDD.n3157 GND 9.03e-19
C8618 VDD.n3158 GND 0.001972f
C8619 VDD.n3159 GND 0.001783f
C8620 VDD.n3160 GND 0.044032f
C8621 VDD.n3161 GND 0.05786f
C8622 VDD.n3162 GND 0.069098f
C8623 VDD.n3163 GND 0.043713f
C8624 VDD.n3164 GND 0.001512f
C8625 VDD.n3165 GND 0.002407f
C8626 VDD.n3166 GND 8.53e-19
C8627 VDD.t401 GND 0.010699f
C8628 VDD.n3167 GND 0.001985f
C8629 VDD.n3168 GND 0.002355f
C8630 VDD.n3169 GND 0.001972f
C8631 VDD.n3170 GND 9.03e-19
C8632 VDD.t393 GND 0.010699f
C8633 VDD.n3171 GND 0.022036f
C8634 VDD.n3172 GND 9.03e-19
C8635 VDD.n3173 GND 8.53e-19
C8636 VDD.n3174 GND 0.002417f
C8637 VDD.n3175 GND 0.007268f
C8638 VDD.n3176 GND 0.065607f
C8639 VDD.n3177 GND 0.06968f
C8640 VDD.n3178 GND 0.043713f
C8641 VDD.n3179 GND 0.004453f
C8642 VDD.n3180 GND 0.002626f
C8643 VDD.n3181 GND 0.002407f
C8644 VDD.n3182 GND 8.53e-19
C8645 VDD.n3183 GND 0.00291f
C8646 VDD.n3184 GND 9.03e-19
C8647 VDD.n3185 GND 0.041407f
C8648 VDD.n3186 GND 8.53e-19
C8649 VDD.n3187 GND 0.00291f
C8650 VDD.t403 GND 0.00545f
C8651 VDD.n3188 GND 0.007088f
C8652 VDD.n3189 GND 0.001115f
C8653 VDD.n3190 GND 0.002183f
C8654 VDD.n3191 GND 0.00291f
C8655 VDD.n3192 GND 9.03e-19
C8656 VDD.n3193 GND 8.53e-19
C8657 VDD.n3194 GND 0.002444f
C8658 VDD.n3195 GND 0.002355f
C8659 VDD.n3196 GND 8.53e-19
C8660 VDD.n3197 GND 9.03e-19
C8661 VDD.n3198 GND 0.002355f
C8662 VDD.n3199 GND 8.53e-19
C8663 VDD.n3200 GND 9.03e-19
C8664 VDD.n3201 GND 0.00291f
C8665 VDD.n3202 GND 0.005733f
C8666 VDD.n3203 GND 9.03e-19
C8667 VDD.n3204 GND 8.53e-19
C8668 VDD.n3205 GND 0.002417f
C8669 VDD.n3206 GND 0.007268f
C8670 VDD.n3207 GND 0.047272f
C8671 VDD.n3208 GND 0.001512f
C8672 VDD.n3209 GND 0.002407f
C8673 VDD.n3210 GND 8.53e-19
C8674 VDD.t439 GND 0.010699f
C8675 VDD.n3211 GND 0.001985f
C8676 VDD.n3212 GND 0.002355f
C8677 VDD.n3213 GND 0.001972f
C8678 VDD.n3214 GND 9.03e-19
C8679 VDD.t426 GND 0.010699f
C8680 VDD.n3215 GND 0.022036f
C8681 VDD.n3216 GND 9.03e-19
C8682 VDD.n3217 GND 8.53e-19
C8683 VDD.n3218 GND 0.002417f
C8684 VDD.n3219 GND 0.007268f
C8685 VDD.n3220 GND 0.05786f
C8686 VDD.n3221 GND 0.068374f
C8687 VDD.n3222 GND 0.043713f
C8688 VDD.n3223 GND 0.001512f
C8689 VDD.n3224 GND 0.002407f
C8690 VDD.n3225 GND 8.53e-19
C8691 VDD.t443 GND 0.010699f
C8692 VDD.n3226 GND 0.001985f
C8693 VDD.n3227 GND 0.002355f
C8694 VDD.n3228 GND 0.001972f
C8695 VDD.n3229 GND 9.03e-19
C8696 VDD.t436 GND 0.010699f
C8697 VDD.n3230 GND 0.022036f
C8698 VDD.n3231 GND 9.03e-19
C8699 VDD.n3232 GND 8.53e-19
C8700 VDD.n3233 GND 0.002417f
C8701 VDD.n3234 GND 0.007268f
C8702 VDD.n3235 GND 0.05786f
C8703 VDD.n3236 GND 0.043713f
C8704 VDD.n3237 GND 0.001512f
C8705 VDD.n3238 GND 0.002407f
C8706 VDD.n3239 GND 8.53e-19
C8707 VDD.t391 GND 0.010699f
C8708 VDD.n3240 GND 0.001985f
C8709 VDD.n3241 GND 0.002355f
C8710 VDD.n3242 GND 0.001972f
C8711 VDD.n3243 GND 9.03e-19
C8712 VDD.t423 GND 0.010699f
C8713 VDD.n3244 GND 0.022036f
C8714 VDD.n3245 GND 9.03e-19
C8715 VDD.n3246 GND 8.53e-19
C8716 VDD.n3247 GND 0.002417f
C8717 VDD.n3248 GND 0.007268f
C8718 VDD.n3249 GND 0.075015f
C8719 VDD.n3250 GND 0.043713f
C8720 VDD.n3251 GND 0.001512f
C8721 VDD.n3252 GND 0.002407f
C8722 VDD.n3253 GND 8.53e-19
C8723 VDD.t412 GND 0.010699f
C8724 VDD.n3254 GND 0.001985f
C8725 VDD.n3255 GND 0.002355f
C8726 VDD.n3256 GND 0.001972f
C8727 VDD.n3257 GND 9.03e-19
C8728 VDD.t404 GND 0.010699f
C8729 VDD.n3258 GND 0.022036f
C8730 VDD.n3259 GND 9.03e-19
C8731 VDD.n3260 GND 8.53e-19
C8732 VDD.n3261 GND 0.002417f
C8733 VDD.n3262 GND 0.007268f
C8734 VDD.n3263 GND 0.075015f
C8735 VDD.n3264 GND 0.043713f
C8736 VDD.n3265 GND 0.001512f
C8737 VDD.n3266 GND 0.002407f
C8738 VDD.n3267 GND 8.53e-19
C8739 VDD.t399 GND 0.010699f
C8740 VDD.n3268 GND 0.001985f
C8741 VDD.n3269 GND 0.002355f
C8742 VDD.n3270 GND 0.001972f
C8743 VDD.n3271 GND 9.03e-19
C8744 VDD.t446 GND 0.010699f
C8745 VDD.n3272 GND 0.022036f
C8746 VDD.n3273 GND 9.03e-19
C8747 VDD.n3274 GND 8.53e-19
C8748 VDD.n3275 GND 0.002417f
C8749 VDD.n3276 GND 0.007268f
C8750 VDD.n3277 GND 0.05786f
C8751 VDD.n3278 GND 0.043713f
C8752 VDD.n3279 GND 0.043713f
C8753 VDD.n3280 GND 0.043713f
C8754 VDD.n3281 GND 0.043713f
C8755 VDD.n3282 GND 0.001512f
C8756 VDD.n3283 GND 0.002407f
C8757 VDD.n3284 GND 8.53e-19
C8758 VDD.t397 GND 0.010699f
C8759 VDD.n3285 GND 0.001985f
C8760 VDD.n3286 GND 0.002355f
C8761 VDD.n3287 GND 0.001972f
C8762 VDD.n3288 GND 9.03e-19
C8763 VDD.t450 GND 0.010699f
C8764 VDD.n3289 GND 0.022036f
C8765 VDD.n3290 GND 9.03e-19
C8766 VDD.n3291 GND 8.53e-19
C8767 VDD.n3292 GND 0.002417f
C8768 VDD.n3293 GND 0.007268f
C8769 VDD.n3294 GND 0.05786f
C8770 VDD.n3295 GND 0.001512f
C8771 VDD.n3296 GND 0.002407f
C8772 VDD.n3297 GND 8.53e-19
C8773 VDD.t407 GND 0.010699f
C8774 VDD.n3298 GND 0.001985f
C8775 VDD.n3299 GND 0.002355f
C8776 VDD.n3300 GND 0.001972f
C8777 VDD.n3301 GND 9.03e-19
C8778 VDD.t441 GND 0.010699f
C8779 VDD.n3302 GND 0.022036f
C8780 VDD.n3303 GND 9.03e-19
C8781 VDD.n3304 GND 8.53e-19
C8782 VDD.n3305 GND 0.002417f
C8783 VDD.n3306 GND 0.007268f
C8784 VDD.n3307 GND 0.076121f
C8785 VDD.n3308 GND 0.001512f
C8786 VDD.n3309 GND 0.002407f
C8787 VDD.n3310 GND 8.53e-19
C8788 VDD.t418 GND 0.010699f
C8789 VDD.n3311 GND 0.001985f
C8790 VDD.n3312 GND 0.002355f
C8791 VDD.n3313 GND 0.001972f
C8792 VDD.n3314 GND 9.03e-19
C8793 VDD.t417 GND 0.010699f
C8794 VDD.n3315 GND 0.022036f
C8795 VDD.n3316 GND 9.03e-19
C8796 VDD.n3317 GND 8.53e-19
C8797 VDD.n3318 GND 0.002417f
C8798 VDD.n3319 GND 0.007268f
C8799 VDD.n3320 GND 0.075015f
C8800 VDD.n3321 GND 0.001512f
C8801 VDD.n3322 GND 0.002407f
C8802 VDD.n3323 GND 8.53e-19
C8803 VDD.t447 GND 0.010699f
C8804 VDD.n3324 GND 0.001985f
C8805 VDD.n3325 GND 0.002355f
C8806 VDD.n3326 GND 0.001972f
C8807 VDD.n3327 GND 9.03e-19
C8808 VDD.t435 GND 0.010699f
C8809 VDD.n3328 GND 0.022036f
C8810 VDD.n3329 GND 9.03e-19
C8811 VDD.n3330 GND 8.53e-19
C8812 VDD.n3331 GND 0.002417f
C8813 VDD.n3332 GND 0.007268f
C8814 VDD.n3333 GND 0.05786f
C8815 VDD.n3334 GND 0.060777f
C8816 VDD.n3335 GND 1.36913f
C8817 VDD.n3336 GND 0.007272f
C8818 VDD.n3337 GND 0.002244f
C8819 VDD.t440 GND 0.010699f
C8820 VDD.t414 GND 0.010699f
C8821 VDD.n3338 GND 0.022031f
C8822 VDD.n3339 GND 9.03e-19
C8823 VDD.n3340 GND 0.001516f
C8824 VDD.n3341 GND 8.53e-19
C8825 VDD.n3342 GND 0.002454f
C8826 VDD.n3343 GND 0.002363f
C8827 VDD.n3344 GND 8.53e-19
C8828 VDD.n3345 GND 9.03e-19
C8829 VDD.n3346 GND 0.001972f
C8830 VDD.n3347 GND 0.001783f
C8831 VDD.n3348 GND 0.044032f
C8832 VDD.n3349 GND 0.076121f
C8833 VDD.n3350 GND 0.007272f
C8834 VDD.n3351 GND 0.002244f
C8835 VDD.t406 GND 0.010699f
C8836 VDD.t389 GND 0.010699f
C8837 VDD.n3352 GND 0.022031f
C8838 VDD.n3353 GND 9.03e-19
C8839 VDD.n3354 GND 0.001516f
C8840 VDD.n3355 GND 8.53e-19
C8841 VDD.n3356 GND 0.002454f
C8842 VDD.n3357 GND 0.002363f
C8843 VDD.n3358 GND 8.53e-19
C8844 VDD.n3359 GND 9.03e-19
C8845 VDD.n3360 GND 0.001972f
C8846 VDD.n3361 GND 0.001783f
C8847 VDD.n3362 GND 0.044032f
C8848 VDD.n3363 GND 0.075015f
C8849 VDD.n3364 GND 0.007272f
C8850 VDD.n3365 GND 0.002244f
C8851 VDD.t445 GND 0.010699f
C8852 VDD.t432 GND 0.010699f
C8853 VDD.n3366 GND 0.022031f
C8854 VDD.n3367 GND 9.03e-19
C8855 VDD.n3368 GND 0.001516f
C8856 VDD.n3369 GND 8.53e-19
C8857 VDD.n3370 GND 0.002454f
C8858 VDD.n3371 GND 0.002363f
C8859 VDD.n3372 GND 8.53e-19
C8860 VDD.n3373 GND 9.03e-19
C8861 VDD.n3374 GND 0.001972f
C8862 VDD.n3375 GND 0.001783f
C8863 VDD.n3376 GND 0.044032f
C8864 VDD.n3377 GND 0.056753f
C8865 VDD.n3378 GND 0.007272f
C8866 VDD.n3379 GND 0.007272f
C8867 VDD.n3380 GND 0.007272f
C8868 VDD.n3381 GND 0.007272f
C8869 VDD.n3382 GND 0.002244f
C8870 VDD.t444 GND 0.010699f
C8871 VDD.t438 GND 0.010699f
C8872 VDD.n3383 GND 0.022031f
C8873 VDD.n3384 GND 9.03e-19
C8874 VDD.n3385 GND 0.001516f
C8875 VDD.n3386 GND 8.53e-19
C8876 VDD.n3387 GND 0.002454f
C8877 VDD.n3388 GND 0.002363f
C8878 VDD.n3389 GND 8.53e-19
C8879 VDD.n3390 GND 9.03e-19
C8880 VDD.n3391 GND 0.001972f
C8881 VDD.n3392 GND 0.001783f
C8882 VDD.n3393 GND 0.044032f
C8883 VDD.n3394 GND 0.05786f
C8884 VDD.n3395 GND 0.002244f
C8885 VDD.t395 GND 0.010699f
C8886 VDD.t428 GND 0.010699f
C8887 VDD.n3396 GND 0.022031f
C8888 VDD.n3397 GND 9.03e-19
C8889 VDD.n3398 GND 0.001516f
C8890 VDD.n3399 GND 8.53e-19
C8891 VDD.n3400 GND 0.002454f
C8892 VDD.n3401 GND 0.002363f
C8893 VDD.n3402 GND 8.53e-19
C8894 VDD.n3403 GND 9.03e-19
C8895 VDD.n3404 GND 0.001972f
C8896 VDD.n3405 GND 0.001783f
C8897 VDD.n3406 GND 0.044032f
C8898 VDD.n3407 GND 0.076121f
C8899 VDD.n3408 GND 0.002244f
C8900 VDD.t411 GND 0.010699f
C8901 VDD.t409 GND 0.010699f
C8902 VDD.n3409 GND 0.022031f
C8903 VDD.n3410 GND 9.03e-19
C8904 VDD.n3411 GND 0.001516f
C8905 VDD.n3412 GND 8.53e-19
C8906 VDD.n3413 GND 0.002454f
C8907 VDD.n3414 GND 0.002363f
C8908 VDD.n3415 GND 8.53e-19
C8909 VDD.n3416 GND 9.03e-19
C8910 VDD.n3417 GND 0.001972f
C8911 VDD.n3418 GND 0.001783f
C8912 VDD.n3419 GND 0.044032f
C8913 VDD.n3420 GND 0.075015f
C8914 VDD.n3421 GND 0.002244f
C8915 VDD.t434 GND 0.010699f
C8916 VDD.t420 GND 0.010699f
C8917 VDD.n3422 GND 0.022031f
C8918 VDD.n3423 GND 9.03e-19
C8919 VDD.n3424 GND 0.001516f
C8920 VDD.n3425 GND 8.53e-19
C8921 VDD.n3426 GND 0.002454f
C8922 VDD.n3427 GND 0.002363f
C8923 VDD.n3428 GND 8.53e-19
C8924 VDD.n3429 GND 9.03e-19
C8925 VDD.n3430 GND 0.001972f
C8926 VDD.n3431 GND 0.001783f
C8927 VDD.n3432 GND 0.044032f
C8928 VDD.n3433 GND 0.05786f
C8929 VDD.n3434 GND 0.062709f
C8930 VDD.n3435 GND 0.00991f
C8931 VDD.n3436 GND 0.001706f
C8932 VDD.n3437 GND 0.012142f
C8933 VDD.n3438 GND 0.001706f
C8934 VDD.n3439 GND 0.001706f
C8935 VDD.n3440 GND 0.119161f
C8936 VDD.n3441 GND 0.001706f
C8937 VDD.t589 GND 0.117408f
C8938 VDD.n3442 GND 0.001706f
C8939 VDD.n3443 GND 0.001706f
C8940 VDD.n3444 GND 8.53e-19
C8941 VDD.n3445 GND 9.03e-19
C8942 VDD.n3446 GND 0.010359f
C8943 VDD.n3447 GND 0.010359f
C8944 VDD.n3448 GND 9.03e-19
C8945 VDD.n3449 GND 8.78e-19
C8946 VDD.n3450 GND 0.001706f
C8947 VDD.n3451 GND 0.001706f
C8948 VDD.n3452 GND 0.026285f
C8949 VDD.n3453 GND 0.001706f
C8950 VDD.n3454 GND 0.001706f
C8951 VDD.n3455 GND 8.53e-19
C8952 VDD.n3456 GND 9.03e-19
C8953 VDD.n3457 GND 0.021453f
C8954 VDD.n3458 GND 0.013609f
C8955 VDD.n3459 GND 0.508412f
C8956 VDD.n3460 GND 0.004436f
C8957 VDD.n3461 GND 0.002626f
C8958 VDD.n3462 GND 0.002407f
C8959 VDD.n3463 GND 8.53e-19
C8960 VDD.n3464 GND 0.00291f
C8961 VDD.n3465 GND 9.03e-19
C8962 VDD.n3466 GND 0.041407f
C8963 VDD.n3467 GND 8.53e-19
C8964 VDD.n3468 GND 0.00291f
C8965 VDD.t646 GND 0.00545f
C8966 VDD.n3469 GND 0.007088f
C8967 VDD.n3470 GND 0.001115f
C8968 VDD.n3471 GND 0.002183f
C8969 VDD.n3472 GND 0.00291f
C8970 VDD.n3473 GND 9.03e-19
C8971 VDD.n3474 GND 8.53e-19
C8972 VDD.n3475 GND 0.002385f
C8973 VDD.n3476 GND 0.002421f
C8974 VDD.n3477 GND 8.53e-19
C8975 VDD.n3478 GND 9.03e-19
C8976 VDD.n3479 GND 0.002366f
C8977 VDD.n3480 GND 8.53e-19
C8978 VDD.n3481 GND 9.03e-19
C8979 VDD.n3482 GND 0.00291f
C8980 VDD.n3483 GND 0.005733f
C8981 VDD.n3484 GND 9.03e-19
C8982 VDD.n3485 GND 8.53e-19
C8983 VDD.n3486 GND 0.002417f
C8984 VDD.n3487 GND 0.007268f
C8985 VDD.n3488 GND 0.050371f
C8986 VDD.n3489 GND 0.044305f
C8987 VDD.n3490 GND 0.001512f
C8988 VDD.n3491 GND 0.002407f
C8989 VDD.n3492 GND 8.53e-19
C8990 VDD.t640 GND 0.010699f
C8991 VDD.n3493 GND 0.001399f
C8992 VDD.n3494 GND 0.002366f
C8993 VDD.n3495 GND 0.001972f
C8994 VDD.n3496 GND 9.03e-19
C8995 VDD.t622 GND 0.010699f
C8996 VDD.n3497 GND 0.02202f
C8997 VDD.n3498 GND 9.03e-19
C8998 VDD.n3499 GND 8.53e-19
C8999 VDD.n3500 GND 0.002417f
C9000 VDD.n3501 GND 0.007268f
C9001 VDD.n3502 GND 0.062508f
C9002 VDD.n3503 GND 0.115599f
C9003 VDD.n3504 GND 0.044305f
C9004 VDD.n3505 GND 0.001512f
C9005 VDD.n3506 GND 0.002407f
C9006 VDD.n3507 GND 8.53e-19
C9007 VDD.t610 GND 0.010699f
C9008 VDD.n3508 GND 0.001399f
C9009 VDD.n3509 GND 0.002366f
C9010 VDD.n3510 GND 0.001972f
C9011 VDD.n3511 GND 9.03e-19
C9012 VDD.t660 GND 0.010699f
C9013 VDD.n3512 GND 0.02202f
C9014 VDD.n3513 GND 9.03e-19
C9015 VDD.n3514 GND 8.53e-19
C9016 VDD.n3515 GND 0.002417f
C9017 VDD.n3516 GND 0.007268f
C9018 VDD.n3517 GND 0.063726f
C9019 VDD.n3518 GND 0.044305f
C9020 VDD.n3519 GND 0.001512f
C9021 VDD.n3520 GND 0.002407f
C9022 VDD.n3521 GND 8.53e-19
C9023 VDD.t650 GND 0.010699f
C9024 VDD.n3522 GND 0.001399f
C9025 VDD.n3523 GND 0.002366f
C9026 VDD.n3524 GND 0.001972f
C9027 VDD.n3525 GND 9.03e-19
C9028 VDD.t632 GND 0.010699f
C9029 VDD.n3526 GND 0.02202f
C9030 VDD.n3527 GND 9.03e-19
C9031 VDD.n3528 GND 8.53e-19
C9032 VDD.n3529 GND 0.002417f
C9033 VDD.n3530 GND 0.007268f
C9034 VDD.n3531 GND 0.081987f
C9035 VDD.n3532 GND 0.044305f
C9036 VDD.n3533 GND 0.001512f
C9037 VDD.n3534 GND 0.002407f
C9038 VDD.n3535 GND 8.53e-19
C9039 VDD.t612 GND 0.010699f
C9040 VDD.n3536 GND 0.001399f
C9041 VDD.n3537 GND 0.002366f
C9042 VDD.n3538 GND 0.001972f
C9043 VDD.n3539 GND 9.03e-19
C9044 VDD.t606 GND 0.010699f
C9045 VDD.n3540 GND 0.02202f
C9046 VDD.n3541 GND 9.03e-19
C9047 VDD.n3542 GND 8.53e-19
C9048 VDD.n3543 GND 0.002417f
C9049 VDD.n3544 GND 0.007268f
C9050 VDD.n3545 GND 0.081987f
C9051 VDD.n3546 GND 0.044305f
C9052 VDD.n3547 GND 0.001512f
C9053 VDD.n3548 GND 0.002407f
C9054 VDD.n3549 GND 8.53e-19
C9055 VDD.t654 GND 0.010699f
C9056 VDD.n3550 GND 0.001399f
C9057 VDD.n3551 GND 0.002366f
C9058 VDD.n3552 GND 0.001972f
C9059 VDD.n3553 GND 9.03e-19
C9060 VDD.t644 GND 0.010699f
C9061 VDD.n3554 GND 0.02202f
C9062 VDD.n3555 GND 9.03e-19
C9063 VDD.n3556 GND 8.53e-19
C9064 VDD.n3557 GND 0.002417f
C9065 VDD.n3558 GND 0.007268f
C9066 VDD.n3559 GND 0.081987f
C9067 VDD.n3560 GND 0.044305f
C9068 VDD.n3561 GND 0.001512f
C9069 VDD.n3562 GND 0.002407f
C9070 VDD.n3563 GND 8.53e-19
C9071 VDD.t626 GND 0.010699f
C9072 VDD.n3564 GND 0.001399f
C9073 VDD.n3565 GND 0.002366f
C9074 VDD.n3566 GND 0.001972f
C9075 VDD.n3567 GND 9.03e-19
C9076 VDD.t604 GND 0.010699f
C9077 VDD.n3568 GND 0.02202f
C9078 VDD.n3569 GND 9.03e-19
C9079 VDD.n3570 GND 8.53e-19
C9080 VDD.n3571 GND 0.002417f
C9081 VDD.n3572 GND 0.007268f
C9082 VDD.n3573 GND 0.081987f
C9083 VDD.n3574 GND 0.044305f
C9084 VDD.n3575 GND 0.001512f
C9085 VDD.n3576 GND 0.002407f
C9086 VDD.n3577 GND 8.53e-19
C9087 VDD.t638 GND 0.010699f
C9088 VDD.n3578 GND 0.001399f
C9089 VDD.n3579 GND 0.002366f
C9090 VDD.n3580 GND 0.001972f
C9091 VDD.n3581 GND 9.03e-19
C9092 VDD.t594 GND 0.010699f
C9093 VDD.n3582 GND 0.02202f
C9094 VDD.n3583 GND 9.03e-19
C9095 VDD.n3584 GND 8.53e-19
C9096 VDD.n3585 GND 0.002417f
C9097 VDD.n3586 GND 0.007268f
C9098 VDD.n3587 GND 0.063726f
C9099 VDD.n3588 GND 0.044305f
C9100 VDD.n3589 GND 0.044305f
C9101 VDD.n3590 GND 0.044305f
C9102 VDD.n3591 GND 0.044305f
C9103 VDD.n3592 GND 0.044305f
C9104 VDD.n3593 GND 0.044305f
C9105 VDD.n3594 GND 0.044305f
C9106 VDD.n3595 GND 0.044305f
C9107 VDD.n3596 GND 0.044305f
C9108 VDD.n3597 GND 0.044305f
C9109 VDD.n3598 GND 0.044305f
C9110 VDD.n3599 GND 0.044305f
C9111 VDD.n3600 GND 0.004436f
C9112 VDD.n3601 GND 0.002626f
C9113 VDD.n3602 GND 0.002407f
C9114 VDD.n3603 GND 8.53e-19
C9115 VDD.n3604 GND 0.00291f
C9116 VDD.n3605 GND 9.03e-19
C9117 VDD.n3606 GND 0.041407f
C9118 VDD.n3607 GND 8.53e-19
C9119 VDD.n3608 GND 0.00291f
C9120 VDD.t624 GND 0.00545f
C9121 VDD.n3609 GND 0.007088f
C9122 VDD.n3610 GND 0.001115f
C9123 VDD.n3611 GND 0.002183f
C9124 VDD.n3612 GND 0.00291f
C9125 VDD.n3613 GND 9.03e-19
C9126 VDD.n3614 GND 8.53e-19
C9127 VDD.n3615 GND 0.002385f
C9128 VDD.n3616 GND 0.002421f
C9129 VDD.n3617 GND 8.53e-19
C9130 VDD.n3618 GND 9.03e-19
C9131 VDD.n3619 GND 0.002366f
C9132 VDD.n3620 GND 8.53e-19
C9133 VDD.n3621 GND 9.03e-19
C9134 VDD.n3622 GND 0.00291f
C9135 VDD.n3623 GND 0.005733f
C9136 VDD.n3624 GND 9.03e-19
C9137 VDD.n3625 GND 8.53e-19
C9138 VDD.n3626 GND 0.002417f
C9139 VDD.n3627 GND 0.007268f
C9140 VDD.n3628 GND 0.051588f
C9141 VDD.n3629 GND 0.001512f
C9142 VDD.n3630 GND 0.002407f
C9143 VDD.n3631 GND 8.53e-19
C9144 VDD.t642 GND 0.010699f
C9145 VDD.n3632 GND 0.001399f
C9146 VDD.n3633 GND 0.002366f
C9147 VDD.n3634 GND 0.001972f
C9148 VDD.n3635 GND 9.03e-19
C9149 VDD.t666 GND 0.010699f
C9150 VDD.n3636 GND 0.02202f
C9151 VDD.n3637 GND 9.03e-19
C9152 VDD.n3638 GND 8.53e-19
C9153 VDD.n3639 GND 0.002417f
C9154 VDD.n3640 GND 0.007268f
C9155 VDD.n3641 GND 0.062508f
C9156 VDD.n3642 GND 0.113942f
C9157 VDD.n3643 GND 0.001512f
C9158 VDD.n3644 GND 0.002407f
C9159 VDD.n3645 GND 8.53e-19
C9160 VDD.t668 GND 0.010699f
C9161 VDD.n3646 GND 0.001399f
C9162 VDD.n3647 GND 0.002366f
C9163 VDD.n3648 GND 0.001972f
C9164 VDD.n3649 GND 9.03e-19
C9165 VDD.t662 GND 0.010699f
C9166 VDD.n3650 GND 0.02202f
C9167 VDD.n3651 GND 9.03e-19
C9168 VDD.n3652 GND 8.53e-19
C9169 VDD.n3653 GND 0.002417f
C9170 VDD.n3654 GND 0.007268f
C9171 VDD.n3655 GND 0.063726f
C9172 VDD.n3656 GND 0.001512f
C9173 VDD.n3657 GND 0.002407f
C9174 VDD.n3658 GND 8.53e-19
C9175 VDD.t634 GND 0.010699f
C9176 VDD.n3659 GND 0.001399f
C9177 VDD.n3660 GND 0.002366f
C9178 VDD.n3661 GND 0.001972f
C9179 VDD.n3662 GND 9.03e-19
C9180 VDD.t596 GND 0.010699f
C9181 VDD.n3663 GND 0.02202f
C9182 VDD.n3664 GND 9.03e-19
C9183 VDD.n3665 GND 8.53e-19
C9184 VDD.n3666 GND 0.002417f
C9185 VDD.n3667 GND 0.007268f
C9186 VDD.n3668 GND 0.081987f
C9187 VDD.n3669 GND 0.001512f
C9188 VDD.n3670 GND 0.002407f
C9189 VDD.n3671 GND 8.53e-19
C9190 VDD.t614 GND 0.010699f
C9191 VDD.n3672 GND 0.001399f
C9192 VDD.n3673 GND 0.002366f
C9193 VDD.n3674 GND 0.001972f
C9194 VDD.n3675 GND 9.03e-19
C9195 VDD.t652 GND 0.010699f
C9196 VDD.n3676 GND 0.02202f
C9197 VDD.n3677 GND 9.03e-19
C9198 VDD.n3678 GND 8.53e-19
C9199 VDD.n3679 GND 0.002417f
C9200 VDD.n3680 GND 0.007268f
C9201 VDD.n3681 GND 0.081987f
C9202 VDD.n3682 GND 0.001512f
C9203 VDD.n3683 GND 0.002407f
C9204 VDD.n3684 GND 8.53e-19
C9205 VDD.t656 GND 0.010699f
C9206 VDD.n3685 GND 0.001399f
C9207 VDD.n3686 GND 0.002366f
C9208 VDD.n3687 GND 0.001972f
C9209 VDD.n3688 GND 9.03e-19
C9210 VDD.t636 GND 0.010699f
C9211 VDD.n3689 GND 0.02202f
C9212 VDD.n3690 GND 9.03e-19
C9213 VDD.n3691 GND 8.53e-19
C9214 VDD.n3692 GND 0.002417f
C9215 VDD.n3693 GND 0.007268f
C9216 VDD.n3694 GND 0.083204f
C9217 VDD.n3695 GND 0.001512f
C9218 VDD.n3696 GND 0.002407f
C9219 VDD.n3697 GND 8.53e-19
C9220 VDD.t616 GND 0.010699f
C9221 VDD.n3698 GND 0.001399f
C9222 VDD.n3699 GND 0.002366f
C9223 VDD.n3700 GND 0.001972f
C9224 VDD.n3701 GND 9.03e-19
C9225 VDD.t600 GND 0.010699f
C9226 VDD.n3702 GND 0.02202f
C9227 VDD.n3703 GND 9.03e-19
C9228 VDD.n3704 GND 8.53e-19
C9229 VDD.n3705 GND 0.002417f
C9230 VDD.n3706 GND 0.007268f
C9231 VDD.n3707 GND 0.081987f
C9232 VDD.n3708 GND 0.001512f
C9233 VDD.n3709 GND 0.002407f
C9234 VDD.n3710 GND 8.53e-19
C9235 VDD.t602 GND 0.010699f
C9236 VDD.n3711 GND 0.001399f
C9237 VDD.n3712 GND 0.002366f
C9238 VDD.n3713 GND 0.001972f
C9239 VDD.n3714 GND 9.03e-19
C9240 VDD.t628 GND 0.010699f
C9241 VDD.n3715 GND 0.02202f
C9242 VDD.n3716 GND 9.03e-19
C9243 VDD.n3717 GND 8.53e-19
C9244 VDD.n3718 GND 0.002417f
C9245 VDD.n3719 GND 0.007268f
C9246 VDD.n3720 GND 0.062508f
C9247 VDD.n3721 GND 0.06242f
C9248 VDD.n3722 GND 0.001512f
C9249 VDD.n3723 GND 0.002407f
C9250 VDD.n3724 GND 8.53e-19
C9251 VDD.t664 GND 0.010699f
C9252 VDD.n3725 GND 0.001399f
C9253 VDD.n3726 GND 0.002366f
C9254 VDD.n3727 GND 0.001972f
C9255 VDD.n3728 GND 9.03e-19
C9256 VDD.t620 GND 0.010699f
C9257 VDD.n3729 GND 0.02202f
C9258 VDD.n3730 GND 9.03e-19
C9259 VDD.n3731 GND 8.53e-19
C9260 VDD.n3732 GND 0.002417f
C9261 VDD.n3733 GND 0.007268f
C9262 VDD.n3734 GND 0.063726f
C9263 VDD.n3735 GND 0.001512f
C9264 VDD.n3736 GND 0.002407f
C9265 VDD.n3737 GND 8.53e-19
C9266 VDD.t598 GND 0.010699f
C9267 VDD.n3738 GND 0.001399f
C9268 VDD.n3739 GND 0.002366f
C9269 VDD.n3740 GND 0.001972f
C9270 VDD.n3741 GND 9.03e-19
C9271 VDD.t592 GND 0.010699f
C9272 VDD.n3742 GND 0.02202f
C9273 VDD.n3743 GND 9.03e-19
C9274 VDD.n3744 GND 8.53e-19
C9275 VDD.n3745 GND 0.002417f
C9276 VDD.n3746 GND 0.007268f
C9277 VDD.n3747 GND 0.081987f
C9278 VDD.n3748 GND 0.001512f
C9279 VDD.n3749 GND 0.002407f
C9280 VDD.n3750 GND 8.53e-19
C9281 VDD.t618 GND 0.010699f
C9282 VDD.n3751 GND 0.001399f
C9283 VDD.n3752 GND 0.002366f
C9284 VDD.n3753 GND 0.001972f
C9285 VDD.n3754 GND 9.03e-19
C9286 VDD.t608 GND 0.010699f
C9287 VDD.n3755 GND 0.02202f
C9288 VDD.n3756 GND 9.03e-19
C9289 VDD.n3757 GND 8.53e-19
C9290 VDD.n3758 GND 0.002417f
C9291 VDD.n3759 GND 0.007268f
C9292 VDD.n3760 GND 0.081987f
C9293 VDD.n3761 GND 0.001512f
C9294 VDD.n3762 GND 0.002407f
C9295 VDD.n3763 GND 8.53e-19
C9296 VDD.t648 GND 0.010699f
C9297 VDD.n3764 GND 0.001399f
C9298 VDD.n3765 GND 0.002366f
C9299 VDD.n3766 GND 0.001972f
C9300 VDD.n3767 GND 9.03e-19
C9301 VDD.t630 GND 0.010699f
C9302 VDD.n3768 GND 0.02202f
C9303 VDD.n3769 GND 9.03e-19
C9304 VDD.n3770 GND 8.53e-19
C9305 VDD.n3771 GND 0.002417f
C9306 VDD.n3772 GND 0.007268f
C9307 VDD.n3773 GND 0.081987f
C9308 VDD.n3774 GND 0.001512f
C9309 VDD.n3775 GND 0.002407f
C9310 VDD.n3776 GND 8.53e-19
C9311 VDD.t590 GND 0.010699f
C9312 VDD.n3777 GND 0.001399f
C9313 VDD.n3778 GND 0.002366f
C9314 VDD.n3779 GND 0.001972f
C9315 VDD.n3780 GND 9.03e-19
C9316 VDD.t658 GND 0.010699f
C9317 VDD.n3781 GND 0.02202f
C9318 VDD.n3782 GND 9.03e-19
C9319 VDD.n3783 GND 8.53e-19
C9320 VDD.n3784 GND 0.002417f
C9321 VDD.n3785 GND 0.007268f
C9322 VDD.n3786 GND 0.062508f
C9323 VDD.n3787 GND 0.06242f
C9324 VDD.n3788 GND 0.506755f
C9325 VDD.n3789 GND 0.859285f
C9326 VDD.n3790 GND 0.010271f
C9327 VDD.n3791 GND 0.017055f
C9328 VDD.n3792 GND 9.03e-19
C9329 VDD.n3793 GND 8.78e-19
C9330 VDD.n3794 GND 0.001706f
C9331 VDD.n3795 GND 0.001706f
C9332 VDD.t663 GND 0.117408f
C9333 VDD.n3796 GND 0.001706f
C9334 VDD.n3797 GND 0.001706f
C9335 VDD.n3798 GND 0.001706f
C9336 VDD.t394 GND 0.117408f
C9337 VDD.n3799 GND 0.001706f
C9338 VDD.n3800 GND 0.001706f
C9339 VDD.n3801 GND 0.001706f
C9340 VDD.n3802 GND 8.53e-19
C9341 VDD.n3803 GND 9.03e-19
C9342 VDD.n3804 GND 0.010359f
C9343 VDD.n3805 GND 0.010359f
C9344 VDD.n3806 GND 8.78e-19
C9345 VDD.n3807 GND 8.53e-19
C9346 VDD.n3808 GND 0.001706f
C9347 VDD.n3809 GND 0.001706f
C9348 VDD.t619 GND 0.117408f
C9349 VDD.n3810 GND 0.119161f
C9350 VDD.n3811 GND 0.001706f
C9351 VDD.n3812 GND 8.53e-19
C9352 VDD.n3813 GND 9.03e-19
C9353 VDD.n3814 GND 0.002444f
C9354 VDD.n3815 GND 8.53e-19
C9355 VDD.n3816 GND 0.001706f
C9356 VDD.t427 GND 0.117408f
C9357 VDD.n3817 GND 0.001706f
C9358 VDD.n3818 GND 0.001706f
C9359 VDD.n3819 GND 0.001706f
C9360 VDD.t601 GND 0.117408f
C9361 VDD.n3820 GND 0.001706f
C9362 VDD.n3821 GND 0.001706f
C9363 VDD.n3822 GND 0.001706f
C9364 VDD.n3823 GND 8.53e-19
C9365 VDD.n3824 GND 0.001706f
C9366 VDD.n3825 GND 0.001706f
C9367 VDD.n3826 GND 0.06659f
C9368 VDD.n3827 GND 0.001706f
C9369 VDD.n3828 GND 0.001706f
C9370 VDD.t627 GND 0.117408f
C9371 VDD.n3829 GND 0.001706f
C9372 VDD.n3830 GND 0.001706f
C9373 VDD.n3831 GND 0.012142f
C9374 VDD.n3832 GND 0.00133f
C9375 VDD.n3833 GND 0.001706f
C9376 VDD.n3834 GND 0.001706f
C9377 VDD.n3835 GND 0.049066f
C9378 VDD.n3836 GND 0.001706f
C9379 VDD.n3837 GND 0.001706f
C9380 VDD.n3838 GND 0.110399f
C9381 VDD.n3839 GND 0.001706f
C9382 VDD.n3840 GND 0.001706f
C9383 VDD.n3841 GND 8.53e-19
C9384 VDD.n3842 GND 9.03e-19
C9385 VDD.n3843 GND 0.002444f
C9386 VDD.n3844 GND 9.03e-19
C9387 VDD.n3845 GND 8.53e-19
C9388 VDD.n3846 GND 0.001706f
C9389 VDD.n3847 GND 9.03e-19
C9390 VDD.n3848 GND 9.03e-19
C9391 VDD.n3849 GND 8.53e-19
C9392 VDD.n3850 GND 0.002444f
C9393 VDD.n3851 GND 0.002444f
C9394 VDD.n3852 GND 0.002444f
C9395 VDD.n3853 GND 8.53e-19
C9396 VDD.n3854 GND 0.001706f
C9397 VDD.n3855 GND 0.119161f
C9398 VDD.n3856 GND 0.001706f
C9399 VDD.n3857 GND 0.001706f
C9400 VDD.n3858 GND 0.001706f
C9401 VDD.t424 GND 0.117408f
C9402 VDD.n3859 GND 0.001706f
C9403 VDD.n3860 GND 0.001706f
C9404 VDD.n3861 GND 0.001706f
C9405 VDD.n3862 GND 0.001706f
C9406 VDD.n3863 GND 0.001706f
C9407 VDD.n3864 GND 0.001706f
C9408 VDD.n3865 GND 0.001706f
C9409 VDD.n3866 GND 0.001706f
C9410 VDD.n3867 GND 0.091123f
C9411 VDD.n3868 GND 0.001706f
C9412 VDD.n3869 GND 0.001706f
C9413 VDD.t415 GND 0.117408f
C9414 VDD.n3870 GND 0.001706f
C9415 VDD.n3871 GND 0.001706f
C9416 VDD.n3872 GND 0.001706f
C9417 VDD.n3873 GND 0.001706f
C9418 VDD.n3874 GND 0.001706f
C9419 VDD.n3875 GND 0.001706f
C9420 VDD.n3876 GND 0.001706f
C9421 VDD.n3877 GND 0.001706f
C9422 VDD.n3878 GND 0.001706f
C9423 VDD.n3879 GND 0.001706f
C9424 VDD.n3880 GND 0.052571f
C9425 VDD.n3881 GND 0.001706f
C9426 VDD.n3882 GND 0.001706f
C9427 VDD.t402 GND 0.117408f
C9428 VDD.n3883 GND 0.001706f
C9429 VDD.n3884 GND 0.003727f
C9430 VDD.n3885 GND 0.003727f
C9431 VDD.n3886 GND 0.014019f
C9432 VDD.n3887 GND 0.003723f
C9433 VDD.n3888 GND 0.003723f
C9434 VDD.n3889 GND 0.187503f
C9435 VDD.n3890 GND 0.003727f
C9436 VDD.n3891 GND 0.001706f
C9437 VDD.n3892 GND 0.001706f
C9438 VDD.n3907 GND 0.003727f
C9439 VDD.n3908 GND 0.075352f
C9440 VDD.n3909 GND 0.001706f
C9441 VDD.n3910 GND 0.001706f
C9442 VDD.n3911 GND 0.031543f
C9443 VDD.n3912 GND 0.001706f
C9444 VDD.n3913 GND 0.070094f
C9445 VDD.n3914 GND 0.001706f
C9446 VDD.n3915 GND 0.001706f
C9447 VDD.n3916 GND 0.001706f
C9448 VDD.n3917 GND 0.108646f
C9449 VDD.n3918 GND 0.001706f
C9450 VDD.n3919 GND 0.001706f
C9451 VDD.n3920 GND 0.119161f
C9452 VDD.n3921 GND 0.001706f
C9453 VDD.n3922 GND 0.001706f
C9454 VDD.n3923 GND 0.012142f
C9455 VDD.n3924 GND 0.024533f
C9456 VDD.n3925 GND 0.001706f
C9457 VDD.n3926 GND 0.001706f
C9458 VDD.n3927 GND 0.063085f
C9459 VDD.n3928 GND 0.001706f
C9460 VDD.n3929 GND 0.001706f
C9461 VDD.n3930 GND 9.03e-19
C9462 VDD.n3931 GND 0.001706f
C9463 VDD.n3932 GND 0.001706f
C9464 VDD.n3933 GND 0.101637f
C9465 VDD.n3934 GND 0.001706f
C9466 VDD.n3935 GND 0.001706f
C9467 VDD.t591 GND 0.117408f
C9468 VDD.n3936 GND 0.001706f
C9469 VDD.n3937 GND 0.001706f
C9470 VDD.n3938 GND 8.53e-19
C9471 VDD.n3939 GND 9.03e-19
C9472 VDD.n3940 GND 0.010359f
C9473 VDD.n3941 GND 9.03e-19
C9474 VDD.n3942 GND 8.53e-19
C9475 VDD.n3943 GND 0.010359f
C9476 VDD.n3944 GND 9.03e-19
C9477 VDD.n3945 GND 8.53e-19
C9478 VDD.n3946 GND 0.001706f
C9479 VDD.n3947 GND 8.78e-19
C9480 VDD.n3948 GND 8.53e-19
C9481 VDD.n3949 GND 9.03e-19
C9482 VDD.n3950 GND 0.001706f
C9483 VDD.n3951 GND 0.001706f
C9484 VDD.t408 GND 0.117408f
C9485 VDD.n3952 GND 0.057828f
C9486 VDD.n3953 GND 0.001706f
C9487 VDD.n3954 GND 9.03e-19
C9488 VDD.n3955 GND 0.018487f
C9489 VDD.n3956 GND 8.53e-19
C9490 VDD.n3957 GND 0.001706f
C9491 VDD.n3958 GND 0.119161f
C9492 VDD.n3959 GND 0.001706f
C9493 VDD.n3960 GND 0.001706f
C9494 VDD.n3961 GND 0.001706f
C9495 VDD.n3962 GND 0.001706f
C9496 VDD.n3963 GND 0.001706f
C9497 VDD.n3964 GND 0.021028f
C9498 VDD.n3965 GND 0.001706f
C9499 VDD.t597 GND 0.117408f
C9500 VDD.n3966 GND 0.001706f
C9501 VDD.n3967 GND 0.001706f
C9502 VDD.n3968 GND 0.001706f
C9503 VDD.n3969 GND 8.53e-19
C9504 VDD.n3970 GND 9.03e-19
C9505 VDD.n3971 GND 0.010359f
C9506 VDD.n3972 GND 9.03e-19
C9507 VDD.n3973 GND 8.53e-19
C9508 VDD.n3974 GND 0.010359f
C9509 VDD.n3975 GND 9.03e-19
C9510 VDD.n3976 GND 8.53e-19
C9511 VDD.n3977 GND 9.03e-19
C9512 VDD.n3978 GND 0.010359f
C9513 VDD.n3979 GND 0.010359f
C9514 VDD.n3980 GND 8.53e-19
C9515 VDD.n3981 GND 0.001706f
C9516 VDD.n3982 GND 8.53e-19
C9517 VDD.n3983 GND 9.03e-19
C9518 VDD.t607 GND 0.117408f
C9519 VDD.t419 GND 0.117408f
C9520 VDD.n3984 GND 0.099885f
C9521 VDD.n3985 GND 0.001706f
C9522 VDD.n3986 GND 0.001706f
C9523 VDD.n3987 GND 8.53e-19
C9524 VDD.n3988 GND 9.03e-19
C9525 VDD.n3989 GND 0.018487f
C9526 VDD.n3990 GND 8.53e-19
C9527 VDD.n3991 GND 0.001706f
C9528 VDD.t617 GND 0.117408f
C9529 VDD.n3992 GND 0.001706f
C9530 VDD.n3993 GND 0.001706f
C9531 VDD.n3994 GND 0.001706f
C9532 VDD.t433 GND 0.117408f
C9533 VDD.n3995 GND 0.001706f
C9534 VDD.n3996 GND 0.001706f
C9535 VDD.n3997 GND 0.001706f
C9536 VDD.n3998 GND 8.53e-19
C9537 VDD.n3999 GND 9.03e-19
C9538 VDD.n4000 GND 0.010359f
C9539 VDD.n4001 GND 0.010359f
C9540 VDD.n4002 GND 9.03e-19
C9541 VDD.n4003 GND 0.010359f
C9542 VDD.n4004 GND 8.53e-19
C9543 VDD.n4005 GND 0.001706f
C9544 VDD.n4006 GND 0.119161f
C9545 VDD.n4007 GND 0.001706f
C9546 VDD.n4008 GND 0.001706f
C9547 VDD.t431 GND 0.117408f
C9548 VDD.n4009 GND 0.001706f
C9549 VDD.n4010 GND 0.001706f
C9550 VDD.n4011 GND 0.001706f
C9551 VDD.n4012 GND 0.001706f
C9552 VDD.n4013 GND 0.001706f
C9553 VDD.n4014 GND 0.001706f
C9554 VDD.n4015 GND 0.001706f
C9555 VDD.n4016 GND 0.001706f
C9556 VDD.n4017 GND 0.05958f
C9557 VDD.n4018 GND 0.001706f
C9558 VDD.n4019 GND 0.001706f
C9559 VDD.n4020 GND 0.098132f
C9560 VDD.n4021 GND 0.001706f
C9561 VDD.n4022 GND 0.001706f
C9562 VDD.n4023 GND 0.119161f
C9563 VDD.n4024 GND 0.001706f
C9564 VDD.n4025 GND 0.001706f
C9565 VDD.n4026 GND 0.001706f
C9566 VDD.n4027 GND 0.038552f
C9567 VDD.n4028 GND 0.001706f
C9568 VDD.t398 GND 0.117408f
C9569 VDD.n4029 GND 0.001706f
C9570 VDD.n4030 GND 0.001706f
C9571 VDD.n4031 GND 0.001706f
C9572 VDD.n4032 GND 8.53e-19
C9573 VDD.n4033 GND 9.03e-19
C9574 VDD.n4034 GND 0.010359f
C9575 VDD.n4035 GND 9.03e-19
C9576 VDD.n4036 GND 8.53e-19
C9577 VDD.n4037 GND 0.010359f
C9578 VDD.n4038 GND 9.03e-19
C9579 VDD.n4039 GND 0.010359f
C9580 VDD.n4040 GND 0.010359f
C9581 VDD.n4041 GND 8.53e-19
C9582 VDD.n4042 GND 0.001706f
C9583 VDD.n4043 GND 0.119161f
C9584 VDD.n4044 GND 0.001706f
C9585 VDD.n4045 GND 0.001706f
C9586 VDD.n4046 GND 8.53e-19
C9587 VDD.n4047 GND 9.03e-19
C9588 VDD.n4048 GND 8.53e-19
C9589 VDD.n4049 GND 0.001706f
C9590 VDD.t388 GND 0.117408f
C9591 VDD.n4050 GND 0.001706f
C9592 VDD.n4051 GND 0.001706f
C9593 VDD.t647 GND 0.117408f
C9594 VDD.n4052 GND 0.001706f
C9595 VDD.n4053 GND 0.001706f
C9596 VDD.n4054 GND 0.001003f
C9597 VDD.n4055 GND 0.012142f
C9598 VDD.n4056 GND 0.001706f
C9599 VDD.n4057 GND 0.077104f
C9600 VDD.n4058 GND 0.001706f
C9601 VDD.t405 GND 0.117408f
C9602 VDD.n4059 GND 0.094628f
C9603 VDD.n4060 GND 0.001706f
C9604 VDD.n4061 GND 0.001706f
C9605 VDD.n4062 GND 0.001706f
C9606 VDD.n4063 GND 0.014019f
C9607 VDD.n4064 GND 0.001706f
C9608 VDD.n4065 GND 0.012142f
C9609 VDD.n4066 GND 0.035047f
C9610 VDD.n4067 GND 0.001706f
C9611 VDD.t413 GND 0.117408f
C9612 VDD.n4068 GND 0.001706f
C9613 VDD.n4069 GND 0.001706f
C9614 VDD.n4070 GND 9.03e-19
C9615 VDD.n4071 GND 0.014037f
C9616 VDD.n4072 GND 0.010359f
C9617 VDD.n4073 GND 9.03e-19
C9618 VDD.n4074 GND 8.53e-19
C9619 VDD.n4075 GND 0.001706f
C9620 VDD.n4076 GND 8.53e-19
C9621 VDD.n4077 GND 9.03e-19
C9622 VDD.t390 GND 0.117408f
C9623 VDD.t593 GND 0.117408f
C9624 VDD.n4078 GND 0.085866f
C9625 VDD.n4079 GND 0.001706f
C9626 VDD.n4080 GND 0.001706f
C9627 VDD.n4081 GND 8.53e-19
C9628 VDD.n4082 GND 9.03e-19
C9629 VDD.n4083 GND 0.002444f
C9630 VDD.n4084 GND 8.53e-19
C9631 VDD.n4085 GND 0.001706f
C9632 VDD.t421 GND 0.117408f
C9633 VDD.n4086 GND 0.001706f
C9634 VDD.n4087 GND 0.001706f
C9635 VDD.n4088 GND 0.001706f
C9636 VDD.t637 GND 0.117408f
C9637 VDD.n4089 GND 0.001706f
C9638 VDD.n4090 GND 0.001706f
C9639 VDD.n4091 GND 0.001706f
C9640 VDD.n4092 GND 0.001706f
C9641 VDD.n4093 GND 0.001706f
C9642 VDD.n4094 GND 0.119161f
C9643 VDD.n4095 GND 0.001706f
C9644 VDD.n4096 GND 0.001706f
C9645 VDD.t603 GND 0.117408f
C9646 VDD.n4097 GND 0.001706f
C9647 VDD.n4098 GND 0.001706f
C9648 VDD.n4099 GND 0.001706f
C9649 VDD.n4100 GND 0.001229f
C9650 VDD.n4101 GND 0.001706f
C9651 VDD.n4102 GND 0.012142f
C9652 VDD.n4103 GND 0.001706f
C9653 VDD.n4104 GND 0.073599f
C9654 VDD.n4105 GND 0.001706f
C9655 VDD.n4106 GND 0.001706f
C9656 VDD.n4107 GND 0.112151f
C9657 VDD.n4108 GND 0.001706f
C9658 VDD.n4109 GND 0.001706f
C9659 VDD.n4110 GND 0.010514f
C9660 VDD.n4111 GND 0.001706f
C9661 VDD.n4112 GND 0.001706f
C9662 VDD.n4113 GND 0.001706f
C9663 VDD.n4114 GND 0.049066f
C9664 VDD.n4115 GND 0.001706f
C9665 VDD.t625 GND 0.117408f
C9666 VDD.n4116 GND 0.001706f
C9667 VDD.n4117 GND 0.001706f
C9668 VDD.n4118 GND 0.001706f
C9669 VDD.n4119 GND 0.001706f
C9670 VDD.n4120 GND 0.001706f
C9671 VDD.n4121 GND 0.087618f
C9672 VDD.n4122 GND 0.001706f
C9673 VDD.n4123 GND 0.001706f
C9674 VDD.t643 GND 0.117408f
C9675 VDD.n4124 GND 0.001706f
C9676 VDD.n4125 GND 0.001706f
C9677 VDD.n4126 GND 0.001706f
C9678 VDD.n4127 GND 0.001706f
C9679 VDD.n4128 GND 0.001706f
C9680 VDD.n4129 GND 0.001706f
C9681 VDD.n4130 GND 8.53e-19
C9682 VDD.n4131 GND 9.03e-19
C9683 VDD.n4132 GND 0.005502f
C9684 VDD.n4133 GND 8.53e-19
C9685 VDD.n4134 GND 0.001706f
C9686 VDD.n4135 GND 0.001706f
C9687 VDD.n4136 GND 0.003723f
C9688 VDD.n4137 GND 0.003723f
C9689 VDD.n4138 GND 0.108646f
C9690 VDD.n4139 GND 0.003723f
C9691 VDD.n4140 GND 0.001706f
C9692 VDD.n4141 GND 0.001706f
C9693 VDD.n4142 GND 0.078856f
C9694 VDD.n4143 GND 0.003727f
C9695 VDD.n4151 GND 0.18575f
C9696 VDD.n4160 GND 0.001706f
C9697 VDD.n4161 GND 0.001706f
C9698 VDD.n4162 GND 0.001706f
C9699 VDD.n4163 GND 0.001706f
C9700 VDD.n4164 GND 0.001706f
C9701 VDD.n4165 GND 0.183998f
C9702 VDD.n4166 GND 0.001706f
C9703 VDD.n4167 GND 0.001706f
C9704 VDD.n4168 GND 0.001706f
C9705 VDD.n4169 GND 0.001706f
C9706 VDD.n4170 GND 0.22255f
C9707 VDD.t611 GND 0.119161f
C9708 VDD.n4171 GND 0.001706f
C9709 VDD.n4172 GND 0.001706f
C9710 VDD.n4173 GND 0.001706f
C9711 VDD.n4174 GND 0.238321f
C9712 VDD.n4175 GND 0.001706f
C9713 VDD.n4176 GND 0.001706f
C9714 VDD.n4177 GND 0.001706f
C9715 VDD.t649 GND 0.119161f
C9716 VDD.n4178 GND 0.001706f
C9717 VDD.n4179 GND 0.001706f
C9718 VDD.n4180 GND 0.001706f
C9719 VDD.t659 GND 0.119161f
C9720 VDD.n4181 GND 0.001706f
C9721 VDD.n4182 GND 0.001706f
C9722 VDD.n4183 GND 0.001706f
C9723 VDD.t609 GND 0.119161f
C9724 VDD.n4184 GND 0.176989f
C9725 VDD.n4185 GND 0.001706f
C9726 VDD.n4186 GND 0.001706f
C9727 VDD.n4187 GND 0.001706f
C9728 VDD.n4188 GND 0.138437f
C9729 VDD.n4189 GND 0.001706f
C9730 VDD.n4190 GND 0.001706f
C9731 VDD.n4191 GND 0.001706f
C9732 VDD.n4192 GND 0.176989f
C9733 VDD.t621 GND 0.119161f
C9734 VDD.n4193 GND 0.001706f
C9735 VDD.n4194 GND 0.001706f
C9736 VDD.n4195 GND 0.001706f
C9737 VDD.n4196 GND 0.215541f
C9738 VDD.n4197 GND 0.001706f
C9739 VDD.n4198 GND 0.003781f
C9740 VDD.n4199 GND 0.003781f
C9741 VDD.n4200 GND 0.315425f
C9742 VDD.t645 GND 0.119161f
C9743 VDD.n4201 GND 0.003781f
C9744 VDD.n4202 GND 0.001706f
C9745 VDD.n4203 GND 0.001706f
C9746 VDD.n4211 GND 0.001706f
C9747 VDD.n4212 GND 0.001706f
C9748 VDD.n4213 GND 0.001706f
C9749 VDD.n4214 GND 0.001706f
C9750 VDD.n4215 GND 0.001706f
C9751 VDD.n4216 GND 0.001706f
C9752 VDD.n4217 GND 0.001706f
C9753 VDD.n4218 GND 0.001706f
C9754 VDD.n4219 GND 0.001706f
C9755 VDD.n4220 GND 0.001706f
C9756 VDD.n4221 GND 0.001706f
C9757 VDD.n4222 GND 0.001706f
C9758 VDD.n4223 GND 0.001706f
C9759 VDD.n4224 GND 0.001706f
C9760 VDD.n4225 GND 0.001706f
C9761 VDD.n4226 GND 0.001706f
C9762 VDD.n4227 GND 0.001706f
C9763 VDD.n4228 GND 0.001706f
C9764 VDD.n4229 GND 0.001706f
C9765 VDD.n4230 GND 0.001706f
C9766 VDD.n4231 GND 0.001706f
C9767 VDD.n4232 GND 0.001706f
C9768 VDD.n4233 GND 0.001706f
C9769 VDD.n4234 GND 0.001706f
C9770 VDD.n4235 GND 0.001706f
C9771 VDD.n4236 GND 0.001706f
C9772 VDD.n4237 GND 0.001706f
C9773 VDD.n4238 GND 0.001706f
C9774 VDD.n4239 GND 0.003795f
C9775 VDD.n4240 GND 0.003795f
C9776 VDD.n4241 GND 0.403043f
C9777 VDD.n4243 GND 0.003795f
C9778 VDD.n4244 GND 0.003795f
C9779 VDD.n4245 GND 0.003781f
C9780 VDD.n4246 GND 0.001706f
C9781 VDD.n4247 GND 0.001706f
C9782 VDD.n4248 GND 0.141941f
C9783 VDD.n4249 GND 0.001706f
C9784 VDD.n4250 GND 0.001706f
C9785 VDD.n4251 GND 0.001706f
C9786 VDD.n4252 GND 0.001706f
C9787 VDD.n4253 GND 0.001706f
C9788 VDD.t639 GND 0.119161f
C9789 VDD.n4254 GND 0.180493f
C9790 VDD.n4255 GND 0.001706f
C9791 VDD.n4256 GND 0.001706f
C9792 VDD.n4257 GND 0.001706f
C9793 VDD.n4258 GND 0.001706f
C9794 VDD.n4259 GND 0.001706f
C9795 VDD.n4260 GND 0.219045f
C9796 VDD.n4261 GND 0.001706f
C9797 VDD.n4262 GND 0.001706f
C9798 VDD.n4263 GND 0.001706f
C9799 VDD.n4264 GND 0.001706f
C9800 VDD.n4265 GND 0.001706f
C9801 VDD.n4266 GND 0.138437f
C9802 VDD.n4267 GND 0.238321f
C9803 VDD.n4268 GND 0.001706f
C9804 VDD.n4269 GND 0.001706f
C9805 VDD.n4270 GND 0.001706f
C9806 VDD.n4271 GND 0.001706f
C9807 VDD.n4272 GND 0.001706f
C9808 VDD.n4273 GND 0.219045f
C9809 VDD.n4274 GND 0.001706f
C9810 VDD.n4275 GND 0.001706f
C9811 VDD.n4276 GND 0.001706f
C9812 VDD.n4277 GND 0.001706f
C9813 VDD.n4278 GND 0.001706f
C9814 VDD.n4279 GND 0.215541f
C9815 VDD.n4280 GND 0.180493f
C9816 VDD.n4281 GND 0.001706f
C9817 VDD.n4282 GND 0.001706f
C9818 VDD.n4283 GND 0.001706f
C9819 VDD.n4284 GND 0.001706f
C9820 VDD.n4285 GND 0.001706f
C9821 VDD.n4286 GND 0.141941f
C9822 VDD.n4287 GND 0.001706f
C9823 VDD.n4288 GND 0.001706f
C9824 VDD.n4289 GND 0.001706f
C9825 VDD.n4290 GND 0.001706f
C9826 VDD.n4291 GND 0.001706f
C9827 VDD.t631 GND 0.119161f
C9828 VDD.n4292 GND 0.134932f
C9829 VDD.n4293 GND 0.001706f
C9830 VDD.n4294 GND 0.001706f
C9831 VDD.n4295 GND 0.001706f
C9832 VDD.n4296 GND 0.001706f
C9833 VDD.n4297 GND 0.001706f
C9834 VDD.n4298 GND 0.001706f
C9835 VDD.n4299 GND 0.173484f
C9836 VDD.n4300 GND 0.001706f
C9837 VDD.n4301 GND 0.001706f
C9838 VDD.n4302 GND 0.001706f
C9839 VDD.n4303 GND 9.17e-19
C9840 VDD.n4304 GND 9.03e-19
C9841 VDD.n4305 GND 0.002444f
C9842 VDD.n4306 GND 9.03e-19
C9843 VDD.n4307 GND 0.002444f
C9844 VDD.n4308 GND 8.53e-19
C9845 VDD.n4309 GND 0.001706f
C9846 VDD.n4310 GND 9.03e-19
C9847 VDD.n4311 GND 0.002313f
C9848 VDD.n4312 GND 8.53e-19
C9849 VDD.n4313 GND 9.03e-19
C9850 VDD.n4314 GND 8.53e-19
C9851 VDD.n4315 GND 0.002444f
C9852 VDD.n4316 GND 0.002444f
C9853 VDD.n4317 GND 8.53e-19
C9854 VDD.n4318 GND 9.03e-19
C9855 VDD.n4319 GND 0.001706f
C9856 VDD.n4320 GND 0.001706f
C9857 VDD.n4321 GND 9.03e-19
C9858 VDD.n4322 GND 8.53e-19
C9859 VDD.n4323 GND 0.002444f
C9860 VDD.n4324 GND 0.002444f
C9861 VDD.n4325 GND 8.53e-19
C9862 VDD.n4326 GND 9.03e-19
C9863 VDD.n4327 GND 8.53e-19
C9864 VDD.n4328 GND 0.001706f
C9865 VDD.n4329 GND 9.03e-19
C9866 VDD.n4330 GND 8.53e-19
C9867 VDD.n4331 GND 0.002444f
C9868 VDD.n4332 GND 0.005502f
C9869 VDD.n4333 GND 8.53e-19
C9870 VDD.n4334 GND 9.03e-19
C9871 VDD.n4335 GND 0.001706f
C9872 VDD.n4336 GND 0.001706f
C9873 VDD.n4337 GND 0.001029f
C9874 VDD.n4338 GND 0.001706f
C9875 VDD.n4339 GND 0.001706f
C9876 VDD.n4340 GND 0.001706f
C9877 VDD.n4341 GND 0.001706f
C9878 VDD.n4342 GND 0.001706f
C9879 VDD.n4343 GND 0.001706f
C9880 VDD.t605 GND 0.119161f
C9881 VDD.n4344 GND 0.212036f
C9882 VDD.n4345 GND 0.001706f
C9883 VDD.n4346 GND 0.001706f
C9884 VDD.n4347 GND 0.001706f
C9885 VDD.n4348 GND 0.001706f
C9886 VDD.n4349 GND 9.03e-19
C9887 VDD.n4350 GND 9.17e-19
C9888 VDD.n4351 GND 0.001029f
C9889 VDD.n4352 GND 0.001706f
C9890 VDD.n4353 GND 0.001706f
C9891 VDD.n4354 GND 0.120913f
C9892 VDD.t653 GND 0.117408f
C9893 VDD.n4355 GND 0.001706f
C9894 VDD.n4356 GND 0.001706f
C9895 VDD.n4357 GND 0.001706f
C9896 VDD.n4358 GND 0.001706f
C9897 VDD.n4359 GND 0.001706f
C9898 VDD.n4360 GND 0.001706f
C9899 VDD.n4361 GND 0.001706f
C9900 VDD.n4362 GND 0.001706f
C9901 VDD.n4363 GND 0.001706f
C9902 VDD.n4364 GND 0.001706f
C9903 VDD.n4365 GND 0.001706f
C9904 VDD.n4366 GND 0.001706f
C9905 VDD.n4367 GND 0.001706f
C9906 VDD.n4368 GND 0.001706f
C9907 VDD.n4369 GND 0.001706f
C9908 VDD.n4370 GND 0.001706f
C9909 VDD.n4371 GND 0.001706f
C9910 VDD.n4372 GND 0.001706f
C9911 VDD.n4373 GND 0.001706f
C9912 VDD.n4374 GND 0.001706f
C9913 VDD.n4375 GND 0.001706f
C9914 VDD.n4376 GND 0.001706f
C9915 VDD.n4377 GND 0.001706f
C9916 VDD.n4378 GND 0.001706f
C9917 VDD.n4379 GND 0.001706f
C9918 VDD.n4380 GND 0.001706f
C9919 VDD.n4381 GND 0.001706f
C9920 VDD.n4382 GND 0.001706f
C9921 VDD.n4383 GND 0.003727f
C9922 VDD.n4384 GND 0.003723f
C9923 VDD.n4385 GND 0.003723f
C9924 VDD.n4386 GND 0.012266f
C9925 VDD.n4387 GND 0.003723f
C9926 VDD.n4388 GND 0.001706f
C9927 VDD.n4389 GND 0.003723f
C9928 VDD.n4390 GND 0.003727f
C9929 VDD.n4391 GND 0.003727f
C9930 VDD.n4392 GND 0.001706f
C9931 VDD.n4393 GND 0.001706f
C9932 VDD.n4394 GND 0.001706f
C9933 VDD.n4395 GND 0.001706f
C9934 VDD.n4396 GND 0.001706f
C9935 VDD.n4397 GND 0.001706f
C9936 VDD.n4398 GND 0.001706f
C9937 VDD.n4399 GND 0.001706f
C9938 VDD.n4400 GND 0.001706f
C9939 VDD.n4401 GND 0.001706f
C9940 VDD.n4402 GND 0.001706f
C9941 VDD.n4403 GND 0.001706f
C9942 VDD.n4404 GND 0.001706f
C9943 VDD.n4405 GND 0.001706f
C9944 VDD.n4406 GND 0.001706f
C9945 VDD.n4407 GND 0.001706f
C9946 VDD.n4408 GND 0.001706f
C9947 VDD.n4409 GND 0.001706f
C9948 VDD.n4410 GND 0.001706f
C9949 VDD.n4411 GND 0.001706f
C9950 VDD.n4412 GND 0.001706f
C9951 VDD.n4413 GND 0.001706f
C9952 VDD.n4414 GND 0.001706f
C9953 VDD.n4415 GND 0.001706f
C9954 VDD.n4416 GND 0.001706f
C9955 VDD.n4417 GND 0.001706f
C9956 VDD.n4418 GND 0.001706f
C9957 VDD.n4419 GND 0.001706f
C9958 VDD.n4420 GND 0.001706f
C9959 VDD.n4421 GND 0.003727f
C9960 VDD.n4422 GND 0.003727f
C9961 VDD.n4423 GND 0.119161f
C9962 VDD.n4425 GND 0.003727f
C9963 VDD.n4426 GND 0.003727f
C9964 VDD.n4427 GND 0.003723f
C9965 VDD.n4428 GND 0.001706f
C9966 VDD.n4429 GND 0.001706f
C9967 VDD.n4430 GND 0.001706f
C9968 VDD.t400 GND 0.117408f
C9969 VDD.n4431 GND 0.033295f
C9970 VDD.n4432 GND 0.001706f
C9971 VDD.n4433 GND 0.001706f
C9972 VDD.n4434 GND 0.001706f
C9973 VDD.n4435 GND 0.001706f
C9974 VDD.n4436 GND 0.001706f
C9975 VDD.n4437 GND 0.001706f
C9976 VDD.t392 GND 0.117408f
C9977 VDD.n4438 GND 0.071847f
C9978 VDD.n4439 GND 0.070094f
C9979 VDD.n4440 GND 0.001706f
C9980 VDD.n4441 GND 9.03e-19
C9981 VDD.n4442 GND 9.03e-19
C9982 VDD.n4443 GND 8.53e-19
C9983 VDD.n4444 GND 0.002444f
C9984 VDD.n4445 GND 0.002444f
C9985 VDD.n4446 GND 0.002444f
C9986 VDD.n4447 GND 9.03e-19
C9987 VDD.n4448 GND 8.53e-19
C9988 VDD.n4449 GND 0.001706f
C9989 VDD.n4450 GND 9.03e-19
C9990 VDD.n4451 GND 8.53e-19
C9991 VDD.n4452 GND 0.002444f
C9992 VDD.n4453 GND 0.002444f
C9993 VDD.n4454 GND 8.53e-19
C9994 VDD.n4455 GND 9.03e-19
C9995 VDD.n4456 GND 0.001706f
C9996 VDD.n4457 GND 0.031543f
C9997 VDD.t429 GND 0.117408f
C9998 VDD.n4458 GND 0.110399f
C9999 VDD.n4459 GND 0.001706f
C10000 VDD.n4460 GND 0.001706f
C10001 VDD.n4461 GND 0.001706f
C10002 VDD.n4462 GND 0.001706f
C10003 VDD.n4463 GND 0.001706f
C10004 VDD.n4464 GND 0.001706f
C10005 VDD.n4465 GND 0.050818f
C10006 VDD.n4466 GND 0.001706f
C10007 VDD.n4467 GND 0.001706f
C10008 VDD.n4468 GND 0.001706f
C10009 VDD.n4469 GND 0.001706f
C10010 VDD.n4470 GND 0.001706f
C10011 VDD.n4471 GND 0.001706f
C10012 VDD.n4472 GND 0.08937f
C10013 VDD.n4473 GND 0.001706f
C10014 VDD.n4474 GND 0.001706f
C10015 VDD.n4475 GND 0.001706f
C10016 VDD.n4476 GND 0.001706f
C10017 VDD.n4477 GND 0.001706f
C10018 VDD.n4478 GND 0.119161f
C10019 VDD.n4479 GND 0.001706f
C10020 VDD.n4480 GND 0.001706f
C10021 VDD.n4481 GND 0.001706f
C10022 VDD.n4482 GND 0.001706f
C10023 VDD.n4483 GND 0.001706f
C10024 VDD.n4484 GND 0.02979f
C10025 VDD.n4485 GND 0.001706f
C10026 VDD.n4486 GND 0.001706f
C10027 VDD.n4487 GND 0.001706f
C10028 VDD.n4488 GND 0.001706f
C10029 VDD.n4489 GND 0.001706f
C10030 VDD.n4490 GND 0.001706f
C10031 VDD.n4491 GND 0.068342f
C10032 VDD.n4492 GND 0.001706f
C10033 VDD.n4493 GND 0.009463f
C10034 VDD.n4494 GND 0.004145f
C10035 VDD.n4495 GND 0.001229f
C10036 VDD.n4496 GND 0.001706f
C10037 VDD.n4497 GND 0.001706f
C10038 VDD.n4498 GND 0.001706f
C10039 VDD.n4499 GND 0.008762f
C10040 VDD.n4500 GND 0.001706f
C10041 VDD.n4501 GND 0.001706f
C10042 VDD.n4502 GND 0.001706f
C10043 VDD.n4503 GND 0.001706f
C10044 VDD.n4504 GND 0.001706f
C10045 VDD.n4505 GND 0.001706f
C10046 VDD.n4506 GND 0.047314f
C10047 VDD.n4507 GND 0.091123f
C10048 VDD.n4508 GND 0.001706f
C10049 VDD.n4509 GND 9.03e-19
C10050 VDD.n4510 GND 9.03e-19
C10051 VDD.n4511 GND 8.53e-19
C10052 VDD.n4512 GND 0.002444f
C10053 VDD.n4513 GND 0.002444f
C10054 VDD.n4514 GND 0.003712f
C10055 VDD.n4515 GND 9.03e-19
C10056 VDD.n4516 GND 8.53e-19
C10057 VDD.n4517 GND 0.001706f
C10058 VDD.n4518 GND 9.03e-19
C10059 VDD.n4519 GND 8.53e-19
C10060 VDD.n4520 GND 0.002444f
C10061 VDD.n4521 GND 0.002444f
C10062 VDD.n4522 GND 8.53e-19
C10063 VDD.n4523 GND 9.03e-19
C10064 VDD.n4524 GND 0.001706f
C10065 VDD.n4525 GND 0.052571f
C10066 VDD.n4526 GND 0.001706f
C10067 VDD.n4527 GND 0.001706f
C10068 VDD.n4528 GND 0.001706f
C10069 VDD.n4529 GND 9.03e-19
C10070 VDD.n4530 GND 8.53e-19
C10071 VDD.n4531 GND 0.010359f
C10072 VDD.n4532 GND 0.010359f
C10073 VDD.n4533 GND 8.53e-19
C10074 VDD.n4534 GND 0.001129f
C10075 VDD.n4535 GND 0.001706f
C10076 VDD.n4536 GND 0.106894f
C10077 VDD.n4537 GND 0.001706f
C10078 VDD.n4538 GND 0.001706f
C10079 VDD.n4539 GND 0.119161f
C10080 VDD.n4540 GND 0.001706f
C10081 VDD.n4541 GND 0.001706f
C10082 VDD.n4542 GND 0.001706f
C10083 VDD.n4543 GND 0.001706f
C10084 VDD.n4544 GND 0.001706f
C10085 VDD.n4545 GND 0.001706f
C10086 VDD.n4546 GND 0.001706f
C10087 VDD.t657 GND 0.117408f
C10088 VDD.n4547 GND 0.001706f
C10089 VDD.n4548 GND 0.001706f
C10090 VDD.n4549 GND 0.043809f
C10091 VDD.n4550 GND 0.001706f
C10092 VDD.n4551 GND 8.53e-19
C10093 VDD.n4552 GND 9.03e-19
C10094 VDD.n4553 GND 8.53e-19
C10095 VDD.n4554 GND 9.03e-19
C10096 VDD.n4555 GND 0.010215f
C10097 VDD.n4556 GND 0.010359f
C10098 VDD.n4557 GND 0.006187f
C10099 VDD.n4558 GND 0.009208f
C10100 VDD.n4559 GND 0.098305f
C10101 VDD.n4560 GND 1.00116f
C10102 VDD.n4561 GND 0.098017f
C10103 VDD.n4562 GND 0.005467f
C10104 VDD.n4563 GND 0.010359f
C10105 VDD.n4564 GND 8.53e-19
C10106 VDD.n4565 GND 0.001706f
C10107 VDD.n4566 GND 9.03e-19
C10108 VDD.n4567 GND 8.53e-19
C10109 VDD.n4568 GND 9.03e-19
C10110 VDD.n4569 GND 8.53e-19
C10111 VDD.n4570 GND 9.03e-19
C10112 VDD.n4571 GND 8.53e-19
C10113 VDD.n4572 GND 0.010359f
C10114 VDD.n4573 GND 0.010359f
C10115 VDD.n4574 GND 8.53e-19
C10116 VDD.n4575 GND 9.03e-19
C10117 VDD.n4576 GND 0.001706f
C10118 VDD.n4577 GND 0.064837f
C10119 VDD.n4578 GND 0.001706f
C10120 VDD.n4579 GND 0.011071f
C10121 VDD.n4580 GND 0.005301f
C10122 VDD.n4581 GND 0.001706f
C10123 VDD.n4582 GND 0.001706f
C10124 VDD.n4583 GND 0.001706f
C10125 VDD.n4584 GND 0.001003f
C10126 VDD.n4585 GND 0.001706f
C10127 VDD.n4586 GND 0.082361f
C10128 VDD.n4587 GND 0.056076f
C10129 VDD.n4588 GND 0.001706f
C10130 VDD.n4589 GND 9.03e-19
C10131 VDD.n4590 GND 9.03e-19
C10132 VDD.n4591 GND 8.53e-19
C10133 VDD.n4592 GND 0.018487f
C10134 VDD.n4593 GND 0.018487f
C10135 VDD.n4594 GND 0.018487f
C10136 VDD.n4595 GND 9.03e-19
C10137 VDD.n4596 GND 8.53e-19
C10138 VDD.n4597 GND 0.001706f
C10139 VDD.n4598 GND 9.03e-19
C10140 VDD.n4599 GND 8.53e-19
C10141 VDD.n4600 GND 0.018487f
C10142 VDD.n4601 GND 0.018487f
C10143 VDD.n4602 GND 8.53e-19
C10144 VDD.n4603 GND 9.03e-19
C10145 VDD.n4604 GND 0.001706f
C10146 VDD.n4605 GND 0.017524f
C10147 VDD.n4606 GND 0.001706f
C10148 VDD.n4607 GND 0.001706f
C10149 VDD.n4608 GND 8.53e-19
C10150 VDD.n4609 GND 9.03e-19
C10151 VDD.n4610 GND 0.001706f
C10152 VDD.n4611 GND 0.001706f
C10153 VDD.n4612 GND 9.03e-19
C10154 VDD.n4613 GND 8.53e-19
C10155 VDD.n4614 GND 0.010359f
C10156 VDD.n4615 GND 0.010359f
C10157 VDD.n4616 GND 8.53e-19
C10158 VDD.n4617 GND 9.03e-19
C10159 VDD.n4618 GND 0.001706f
C10160 VDD.n4619 GND 0.103389f
C10161 VDD.n4620 GND 0.001706f
C10162 VDD.n4621 GND 0.001706f
C10163 VDD.n4622 GND 0.001706f
C10164 VDD.n4623 GND 0.001706f
C10165 VDD.n4624 GND 0.001706f
C10166 VDD.t629 GND 0.119161f
C10167 VDD.n4625 GND 0.001706f
C10168 VDD.n4626 GND 0.001706f
C10169 VDD.n4627 GND 0.001706f
C10170 VDD.n4628 GND 0.001706f
C10171 VDD.n4629 GND 0.001706f
C10172 VDD.n4630 GND 0.001706f
C10173 VDD.n4631 GND 0.001706f
C10174 VDD.n4632 GND 0.001706f
C10175 VDD.n4633 GND 0.001706f
C10176 VDD.n4634 GND 0.001706f
C10177 VDD.n4635 GND 0.001706f
C10178 VDD.n4636 GND 0.001706f
C10179 VDD.n4637 GND 0.001706f
C10180 VDD.n4638 GND 0.001706f
C10181 VDD.n4639 GND 0.040304f
C10182 VDD.n4640 GND 0.001706f
C10183 VDD.n4641 GND 0.001706f
C10184 VDD.n4642 GND 0.001706f
C10185 VDD.n4643 GND 0.001706f
C10186 VDD.n4644 GND 0.001706f
C10187 VDD.n4645 GND 0.078856f
C10188 VDD.n4646 GND 0.001706f
C10189 VDD.n4647 GND 0.001706f
C10190 VDD.n4648 GND 0.001706f
C10191 VDD.n4649 GND 0.001706f
C10192 VDD.n4650 GND 0.001706f
C10193 VDD.n4651 GND 0.001706f
C10194 VDD.n4652 GND 0.022781f
C10195 VDD.n4653 GND 0.001706f
C10196 VDD.n4654 GND 9.03e-19
C10197 VDD.n4655 GND 9.03e-19
C10198 VDD.n4656 GND 8.53e-19
C10199 VDD.n4657 GND 0.010359f
C10200 VDD.n4658 GND 0.010359f
C10201 VDD.n4659 GND 0.010359f
C10202 VDD.n4660 GND 8.53e-19
C10203 VDD.n4661 GND 9.03e-19
C10204 VDD.n4662 GND 8.53e-19
C10205 VDD.n4663 GND 9.03e-19
C10206 VDD.n4664 GND 8.53e-19
C10207 VDD.n4665 GND 0.010359f
C10208 VDD.n4666 GND 0.010359f
C10209 VDD.n4667 GND 8.53e-19
C10210 VDD.n4668 GND 8.78e-19
C10211 VDD.n4669 GND 8.78e-19
C10212 VDD.n4670 GND 0.001706f
C10213 VDD.n4671 GND 0.061333f
C10214 VDD.n4672 GND 0.080609f
C10215 VDD.n4673 GND 0.001706f
C10216 VDD.n4674 GND 9.03e-19
C10217 VDD.n4675 GND 9.03e-19
C10218 VDD.n4676 GND 8.53e-19
C10219 VDD.n4677 GND 0.018487f
C10220 VDD.n4678 GND 0.018487f
C10221 VDD.n4679 GND 9.03e-19
C10222 VDD.n4680 GND 8.53e-19
C10223 VDD.n4681 GND 0.018487f
C10224 VDD.n4682 GND 0.018487f
C10225 VDD.n4683 GND 8.53e-19
C10226 VDD.n4684 GND 9.03e-19
C10227 VDD.n4685 GND 0.001706f
C10228 VDD.n4686 GND 0.042057f
C10229 VDD.n4687 GND 0.001706f
C10230 VDD.n4688 GND 0.001706f
C10231 VDD.n4689 GND 0.003505f
C10232 VDD.n4690 GND 0.001706f
C10233 VDD.n4691 GND 9.03e-19
C10234 VDD.n4692 GND 8.53e-19
C10235 VDD.n4693 GND 0.010359f
C10236 VDD.n4694 GND 0.010359f
C10237 VDD.n4695 GND 8.53e-19
C10238 VDD.n4696 GND 9.03e-19
C10239 VDD.n4697 GND 0.001706f
C10240 VDD.n4698 GND 0.117408f
C10241 VDD.n4699 GND 0.001706f
C10242 VDD.n4700 GND 0.001706f
C10243 VDD.n4701 GND 0.001706f
C10244 VDD.n4702 GND 0.001706f
C10245 VDD.n4703 GND 0.001706f
C10246 VDD.n4704 GND 0.001706f
C10247 VDD.t410 GND 0.117408f
C10248 VDD.n4705 GND 0.019276f
C10249 VDD.n4706 GND 0.119161f
C10250 VDD.n4707 GND 0.001706f
C10251 VDD.n4708 GND 9.03e-19
C10252 VDD.n4709 GND 8.53e-19
C10253 VDD.n4710 GND 0.018487f
C10254 VDD.n4711 GND 0.018487f
C10255 VDD.n4712 GND 8.53e-19
C10256 VDD.n4713 GND 8.53e-19
C10257 VDD.n4714 GND 9.03e-19
C10258 VDD.n4715 GND 0.001706f
C10259 VDD.n4716 GND 0.084113f
C10260 VDD.n4717 GND 0.001706f
C10261 VDD.n4718 GND 9.03e-19
C10262 VDD.n4719 GND 8.53e-19
C10263 VDD.n4720 GND 0.010359f
C10264 VDD.n4721 GND 0.010359f
C10265 VDD.n4722 GND 8.53e-19
C10266 VDD.n4723 GND 9.03e-19
C10267 VDD.n4724 GND 0.001706f
C10268 VDD.n4725 GND 0.0368f
C10269 VDD.n4726 GND 0.001706f
C10270 VDD.n4727 GND 0.001706f
C10271 VDD.n4728 GND 9.03e-19
C10272 VDD.n4729 GND 0.005814f
C10273 VDD.n4730 GND 0.012142f
C10274 VDD.n4731 GND 0.011785f
C10275 VDD.n4732 GND 0.001706f
C10276 VDD.n4733 GND 0.075352f
C10277 VDD.n4734 GND 0.001706f
C10278 VDD.n4735 GND 0.001706f
C10279 VDD.n4736 GND 0.001706f
C10280 VDD.n4737 GND 0.001706f
C10281 VDD.n4738 GND 0.001706f
C10282 VDD.n4739 GND 0.113904f
C10283 VDD.n4740 GND 0.001706f
C10284 VDD.n4741 GND 0.001706f
C10285 VDD.n4742 GND 0.007589f
C10286 VDD.n4743 GND 0.001706f
C10287 VDD.n4744 GND 0.012142f
C10288 VDD.n4745 GND 0.010624f
C10289 VDD.n4746 GND 0.001706f
C10290 VDD.n4747 GND 0.015771f
C10291 VDD.n4748 GND 0.001706f
C10292 VDD.n4749 GND 0.001706f
C10293 VDD.n4750 GND 0.001706f
C10294 VDD.n4751 GND 0.001706f
C10295 VDD.n4752 GND 8.53e-19
C10296 VDD.n4753 GND 9.03e-19
C10297 VDD.n4754 GND 0.010359f
C10298 VDD.n4755 GND 8.53e-19
C10299 VDD.n4756 GND 0.001706f
C10300 VDD.n4757 GND 9.03e-19
C10301 VDD.n4758 GND 9.03e-19
C10302 VDD.n4759 GND 8.53e-19
C10303 VDD.n4760 GND 0.010359f
C10304 VDD.n4761 GND 9.03e-19
C10305 VDD.n4762 GND 9.03e-19
C10306 VDD.n4763 GND 8.53e-19
C10307 VDD.n4764 GND 0.010359f
C10308 VDD.n4765 GND 0.010359f
C10309 VDD.n4766 GND 0.014703f
C10310 VDD.n4767 GND 0.002444f
C10311 VDD.t615 GND 0.117408f
C10312 VDD.n4768 GND 0.010514f
C10313 VDD.n4769 GND 0.001706f
C10314 VDD.n4770 GND 9.03e-19
C10315 VDD.n4771 GND 0.002444f
C10316 VDD.n4772 GND 8.53e-19
C10317 VDD.n4773 GND 0.001706f
C10318 VDD.n4774 GND 9.03e-19
C10319 VDD.n4775 GND 0.002444f
C10320 VDD.n4776 GND 9.17e-19
C10321 VDD.n4777 GND 0.001706f
C10322 VDD.n4778 GND 0.001706f
C10323 VDD.n4779 GND 0.001706f
C10324 VDD.n4780 GND 0.001706f
C10325 VDD.t613 GND 0.119161f
C10326 VDD.n4781 GND 0.183998f
C10327 VDD.n4782 GND 0.001706f
C10328 VDD.n4783 GND 0.001706f
C10329 VDD.n4784 GND 0.001706f
C10330 VDD.n4785 GND 0.001706f
C10331 VDD.n4786 GND 9.03e-19
C10332 VDD.n4787 GND 0.002444f
C10333 VDD.n4788 GND 8.53e-19
C10334 VDD.n4789 GND 9.03e-19
C10335 VDD.n4790 GND 0.002444f
C10336 VDD.n4791 GND 8.53e-19
C10337 VDD.n4792 GND 9.03e-19
C10338 VDD.n4793 GND 0.001706f
C10339 VDD.n4794 GND 0.001706f
C10340 VDD.n4795 GND 9.03e-19
C10341 VDD.n4796 GND 8.53e-19
C10342 VDD.n4797 GND 0.005502f
C10343 VDD.n4798 GND 9.17e-19
C10344 VDD.n4799 GND 0.001029f
C10345 VDD.n4800 GND 0.001706f
C10346 VDD.n4801 GND 0.001706f
C10347 VDD.n4802 GND 0.001706f
C10348 VDD.n4803 GND 0.001706f
C10349 VDD.n4804 GND 0.001706f
C10350 VDD.n4805 GND 0.001706f
C10351 VDD.n4806 GND 0.001706f
C10352 VDD.t651 GND 0.119161f
C10353 VDD.n4807 GND 0.001706f
C10354 VDD.n4808 GND 0.001706f
C10355 VDD.n4809 GND 0.001706f
C10356 VDD.n4810 GND 0.238321f
C10357 VDD.n4811 GND 0.001706f
C10358 VDD.n4812 GND 0.001706f
C10359 VDD.n4813 GND 0.001706f
C10360 VDD.n4814 GND 0.001706f
C10361 VDD.n4815 GND 0.001706f
C10362 VDD.n4816 GND 0.001706f
C10363 VDD.t667 GND 0.119161f
C10364 VDD.n4817 GND 0.001706f
C10365 VDD.n4818 GND 0.001706f
C10366 VDD.n4819 GND 0.001706f
C10367 VDD.n4820 GND 0.176989f
C10368 VDD.n4821 GND 0.001706f
C10369 VDD.n4822 GND 0.001706f
C10370 VDD.n4823 GND 0.001706f
C10371 VDD.n4824 GND 0.138437f
C10372 VDD.n4825 GND 0.001706f
C10373 VDD.n4826 GND 0.001706f
C10374 VDD.n4827 GND 0.001706f
C10375 VDD.t641 GND 0.119161f
C10376 VDD.n4828 GND 0.001706f
C10377 VDD.n4829 GND 0.001706f
C10378 VDD.n4830 GND 0.001706f
C10379 VDD.n4831 GND 0.215541f
C10380 VDD.n4832 GND 0.001706f
C10381 VDD.n4833 GND 0.003781f
C10382 VDD.n4834 GND 0.003781f
C10383 VDD.t623 GND 0.119161f
C10384 VDD.n4835 GND 0.001706f
C10385 VDD.n4836 GND 0.003781f
C10386 VDD.n4844 GND 0.001706f
C10387 VDD.n4845 GND 0.001706f
C10388 VDD.n4846 GND 0.001706f
C10389 VDD.n4847 GND 0.001706f
C10390 VDD.n4848 GND 0.001706f
C10391 VDD.n4849 GND 0.001706f
C10392 VDD.n4850 GND 0.001706f
C10393 VDD.n4851 GND 0.001706f
C10394 VDD.n4852 GND 0.001706f
C10395 VDD.n4853 GND 0.001706f
C10396 VDD.n4854 GND 0.001706f
C10397 VDD.n4855 GND 0.001706f
C10398 VDD.n4856 GND 0.001706f
C10399 VDD.n4857 GND 0.001706f
C10400 VDD.n4858 GND 0.001706f
C10401 VDD.n4859 GND 0.001706f
C10402 VDD.n4860 GND 0.001706f
C10403 VDD.n4861 GND 0.001706f
C10404 VDD.n4862 GND 0.001706f
C10405 VDD.n4863 GND 0.001706f
C10406 VDD.n4864 GND 0.001706f
C10407 VDD.n4865 GND 0.001706f
C10408 VDD.n4866 GND 0.001706f
C10409 VDD.n4867 GND 0.001706f
C10410 VDD.n4868 GND 0.003781f
C10411 VDD.n4869 GND 0.003795f
C10412 VDD.n4870 GND 0.003795f
C10413 VDD.n4871 GND 0.001706f
C10414 VDD.n4872 GND 0.001706f
C10415 VDD.n4873 GND 0.001706f
C10416 VDD.n4874 GND 0.001706f
C10417 VDD.n4875 GND 0.001706f
C10418 VDD.n4876 GND 0.001706f
C10419 VDD.n4877 GND 0.001706f
C10420 VDD.n4878 GND 0.001706f
C10421 VDD.n4879 GND 0.001706f
C10422 VDD.n4880 GND 0.001706f
C10423 VDD.n4881 GND 0.001706f
C10424 VDD.n4882 GND 0.001706f
C10425 VDD.n4883 GND 0.001706f
C10426 VDD.n4884 GND 0.001706f
C10427 VDD.n4885 GND 0.001706f
C10428 VDD.n4886 GND 0.001706f
C10429 VDD.n4887 GND 0.001706f
C10430 VDD.n4888 GND 0.001706f
C10431 VDD.n4889 GND 0.001706f
C10432 VDD.n4890 GND 0.001706f
C10433 VDD.n4891 GND 0.001706f
C10434 VDD.n4892 GND 0.001706f
C10435 VDD.n4893 GND 0.001706f
C10436 VDD.n4894 GND 0.001706f
C10437 VDD.n4895 GND 0.001706f
C10438 VDD.n4896 GND 0.001706f
C10439 VDD.n4897 GND 0.001706f
C10440 VDD.n4898 GND 0.001706f
C10441 VDD.n4899 GND 0.003795f
C10442 VDD.n4900 GND 0.003795f
C10443 VDD.n4902 GND 0.382015f
C10444 VDD.n4903 GND 0.315425f
C10445 VDD.n4904 GND 0.141941f
C10446 VDD.n4905 GND 0.001706f
C10447 VDD.n4906 GND 0.001706f
C10448 VDD.n4907 GND 0.001706f
C10449 VDD.n4908 GND 0.001706f
C10450 VDD.n4909 GND 0.001706f
C10451 VDD.n4910 GND 0.180493f
C10452 VDD.t665 GND 0.119161f
C10453 VDD.n4911 GND 0.176989f
C10454 VDD.n4912 GND 0.219045f
C10455 VDD.n4913 GND 0.001706f
C10456 VDD.n4914 GND 0.001706f
C10457 VDD.n4915 GND 0.001706f
C10458 VDD.n4916 GND 0.001706f
C10459 VDD.n4917 GND 0.001706f
C10460 VDD.n4918 GND 0.238321f
C10461 VDD.n4919 GND 0.138437f
C10462 VDD.t661 GND 0.119161f
C10463 VDD.n4920 GND 0.219045f
C10464 VDD.n4921 GND 0.001706f
C10465 VDD.n4922 GND 0.001706f
C10466 VDD.n4923 GND 0.001706f
C10467 VDD.n4924 GND 0.001706f
C10468 VDD.n4925 GND 0.001706f
C10469 VDD.n4926 GND 0.180493f
C10470 VDD.n4927 GND 0.215541f
C10471 VDD.t595 GND 0.119161f
C10472 VDD.n4928 GND 0.141941f
C10473 VDD.n4929 GND 0.001706f
C10474 VDD.n4930 GND 0.001706f
C10475 VDD.n4931 GND 0.001706f
C10476 VDD.n4932 GND 0.001706f
C10477 VDD.n4933 GND 0.001706f
C10478 VDD.n4934 GND 0.134932f
C10479 VDD.t633 GND 0.119161f
C10480 VDD.n4935 GND 0.22255f
C10481 VDD.n4936 GND 0.173484f
C10482 VDD.n4937 GND 0.001706f
C10483 VDD.n4938 GND 0.001706f
C10484 VDD.n4939 GND 0.001706f
C10485 VDD.n4940 GND 0.001706f
C10486 VDD.n4941 GND 0.001706f
C10487 VDD.n4942 GND 0.212036f
C10488 VDD.n4943 GND 0.001706f
C10489 VDD.n4944 GND 0.001706f
C10490 VDD.n4945 GND 0.001706f
C10491 VDD.n4946 GND 0.001706f
C10492 VDD.n4947 GND 0.001706f
C10493 VDD.n4948 GND 0.001029f
C10494 VDD.n4949 GND 0.001706f
C10495 VDD.n4950 GND 0.001706f
C10496 VDD.n4951 GND 9.03e-19
C10497 VDD.n4952 GND 8.53e-19
C10498 VDD.n4953 GND 0.005502f
C10499 VDD.n4954 GND 0.002444f
C10500 VDD.n4955 GND 8.53e-19
C10501 VDD.n4956 GND 9.03e-19
C10502 VDD.n4957 GND 0.001706f
C10503 VDD.n4958 GND 0.001706f
C10504 VDD.n4959 GND 9.03e-19
C10505 VDD.n4960 GND 8.53e-19
C10506 VDD.n4961 GND 9.03e-19
C10507 VDD.n4962 GND 8.53e-19
C10508 VDD.n4963 GND 0.002444f
C10509 VDD.n4964 GND 0.002444f
C10510 VDD.n4965 GND 8.53e-19
C10511 VDD.n4966 GND 9.03e-19
C10512 VDD.n4967 GND 8.53e-19
C10513 VDD.n4968 GND 0.001706f
C10514 VDD.n4969 GND 9.03e-19
C10515 VDD.n4970 GND 8.53e-19
C10516 VDD.n4971 GND 0.002444f
C10517 VDD.n4972 GND 0.002375f
C10518 VDD.n4973 GND 8.53e-19
C10519 VDD.n4974 GND 9.03e-19
C10520 VDD.n4975 GND 0.001706f
C10521 VDD.n4976 GND 0.087618f
C10522 VDD.n4977 GND 0.001706f
C10523 VDD.t396 GND 0.117408f
C10524 VDD.n4978 GND 0.054323f
C10525 VDD.n4979 GND 0.001706f
C10526 VDD.n4980 GND 0.001706f
C10527 VDD.n4981 GND 0.001706f
C10528 VDD.n4982 GND 0.001706f
C10529 VDD.n4983 GND 0.001706f
C10530 VDD.n4984 GND 0.001706f
C10531 VDD.n4985 GND 0.001706f
C10532 VDD.n4986 GND 0.001706f
C10533 VDD.n4987 GND 0.001706f
C10534 VDD.n4988 GND 0.001706f
C10535 VDD.n4989 GND 0.001706f
C10536 VDD.t599 GND 0.117408f
C10537 VDD.n4990 GND 0.02979f
C10538 VDD.n4991 GND 0.001706f
C10539 VDD.n4992 GND 0.001706f
C10540 VDD.n4993 GND 0.001706f
C10541 VDD.n4994 GND 0.001706f
C10542 VDD.n4995 GND 0.001706f
C10543 VDD.t655 GND 0.117408f
C10544 VDD.n4996 GND 0.068342f
C10545 VDD.n4997 GND 0.001706f
C10546 VDD.n4998 GND 0.001706f
C10547 VDD.n4999 GND 0.001706f
C10548 VDD.n5000 GND 0.001706f
C10549 VDD.n5001 GND 0.001706f
C10550 VDD.n5002 GND 0.001706f
C10551 VDD.n5003 GND 0.001706f
C10552 VDD.n5004 GND 0.001706f
C10553 VDD.n5005 GND 0.001706f
C10554 VDD.n5006 GND 0.001706f
C10555 VDD.n5007 GND 0.001706f
C10556 VDD.n5008 GND 0.001706f
C10557 VDD.n5009 GND 0.001706f
C10558 VDD.n5010 GND 0.001706f
C10559 VDD.n5011 GND 0.001706f
C10560 VDD.n5012 GND 0.001706f
C10561 VDD.n5013 GND 0.001706f
C10562 VDD.n5014 GND 0.001706f
C10563 VDD.n5015 GND 0.001706f
C10564 VDD.n5016 GND 0.001706f
C10565 VDD.n5017 GND 0.001706f
C10566 VDD.n5018 GND 0.001706f
C10567 VDD.n5019 GND 0.001706f
C10568 VDD.n5020 GND 0.001706f
C10569 VDD.n5021 GND 0.001706f
C10570 VDD.n5022 GND 0.001706f
C10571 VDD.n5023 GND 0.001706f
C10572 VDD.n5024 GND 0.001706f
C10573 VDD.n5025 GND 0.001706f
C10574 VDD.n5026 GND 0.003727f
C10575 VDD.n5027 GND 0.003723f
C10576 VDD.n5028 GND 0.001706f
C10577 VDD.n5029 GND 0.001706f
C10578 VDD.t635 GND 0.117408f
C10579 VDD.n5030 GND 0.106894f
C10580 VDD.n5031 GND 0.001706f
C10581 VDD.n5032 GND 0.001706f
C10582 VDD.n5033 GND 0.003723f
C10583 VDD.n5034 GND 0.003727f
C10584 VDD.n5035 GND 0.003727f
C10585 VDD.n5036 GND 0.001706f
C10586 VDD.n5037 GND 0.001706f
C10587 VDD.n5038 GND 0.001706f
C10588 VDD.n5039 GND 0.001706f
C10589 VDD.n5040 GND 0.001706f
C10590 VDD.n5041 GND 0.001706f
C10591 VDD.n5042 GND 0.001706f
C10592 VDD.n5043 GND 0.001706f
C10593 VDD.n5044 GND 0.001706f
C10594 VDD.n5045 GND 0.001706f
C10595 VDD.n5046 GND 0.001706f
C10596 VDD.n5047 GND 0.001706f
C10597 VDD.n5048 GND 0.001706f
C10598 VDD.n5049 GND 0.001706f
C10599 VDD.n5050 GND 0.001706f
C10600 VDD.n5051 GND 0.001706f
C10601 VDD.n5052 GND 0.001706f
C10602 VDD.n5053 GND 0.001706f
C10603 VDD.n5054 GND 0.001706f
C10604 VDD.n5055 GND 0.001706f
C10605 VDD.n5056 GND 0.001706f
C10606 VDD.n5057 GND 0.001706f
C10607 VDD.n5058 GND 0.001706f
C10608 VDD.n5059 GND 0.001706f
C10609 VDD.n5060 GND 0.001706f
C10610 VDD.n5061 GND 0.001706f
C10611 VDD.n5062 GND 0.001706f
C10612 VDD.n5063 GND 0.001706f
C10613 VDD.n5064 GND 0.001706f
C10614 VDD.n5066 GND 0.119161f
C10615 VDD.n5068 GND 0.001706f
C10616 VDD.n5069 GND 0.001706f
C10617 VDD.n5070 GND 0.003727f
C10618 VDD.n5071 GND 0.003723f
C10619 VDD.n5072 GND 0.003723f
C10620 VDD.n5073 GND 0.119161f
C10621 VDD.n5074 GND 0.003723f
C10622 VDD.n5075 GND 0.003723f
C10623 VDD.n5076 GND 0.001706f
C10624 VDD.n5077 GND 0.001706f
C10625 VDD.n5078 GND 0.001706f
C10626 VDD.n5079 GND 0.08937f
C10627 VDD.n5080 GND 0.001706f
C10628 VDD.n5081 GND 0.001706f
C10629 VDD.n5082 GND 0.001706f
C10630 VDD.n5083 GND 0.001706f
C10631 VDD.n5084 GND 0.001706f
C10632 VDD.n5085 GND 0.050818f
C10633 VDD.n5086 GND 0.001706f
C10634 VDD.n5087 GND 0.001706f
C10635 VDD.n5088 GND 0.001706f
C10636 VDD.n5089 GND 0.001706f
C10637 VDD.n5090 GND 0.001706f
C10638 VDD.n5091 GND 0.012266f
C10639 VDD.n5092 GND 0.119161f
C10640 VDD.n5093 GND 0.001706f
C10641 VDD.n5094 GND 9.03e-19
C10642 VDD.n5095 GND 8.53e-19
C10643 VDD.n5096 GND 0.002444f
C10644 VDD.n5097 GND 0.002444f
C10645 VDD.n5098 GND 8.53e-19
C10646 VDD.n5099 GND 9.03e-19
C10647 VDD.n5100 GND 0.001706f
C10648 VDD.n5101 GND 0.028038f
C10649 VDD.t437 GND 0.117408f
C10650 VDD.n5102 GND 0.092875f
C10651 VDD.n5103 GND 0.001706f
C10652 VDD.n5104 GND 0.00133f
C10653 VDD.n5105 GND 0.003632f
C10654 VDD.n5106 GND 0.008749f
C10655 VDD.n5107 GND 0.001706f
C10656 VDD.n5108 GND 0.071847f
C10657 VDD.n5109 GND 0.001706f
C10658 VDD.n5110 GND 0.001706f
C10659 VDD.n5111 GND 0.001706f
C10660 VDD.n5112 GND 0.001129f
C10661 VDD.n5113 GND 0.001706f
C10662 VDD.n5114 GND 0.033295f
C10663 VDD.n5115 GND 0.105142f
C10664 VDD.n5116 GND 0.001706f
C10665 VDD.n5117 GND 9.03e-19
C10666 VDD.n5118 GND 8.53e-19
C10667 VDD.n5119 GND 0.002444f
C10668 VDD.n5120 GND 0.002316f
C10669 VDD.n5121 GND 8.53e-19
C10670 VDD.n5122 GND 9.03e-19
C10671 VDD.n5123 GND 0.001706f
C10672 VDD.n5124 GND 0.007009f
C10673 VDD.n5125 GND 0.001706f
C10674 VDD.n5126 GND 9.03e-19
C10675 VDD.n5127 GND 8.53e-19
C10676 VDD.n5128 GND 0.010359f
C10677 VDD.n5129 GND 0.010359f
C10678 VDD.n5130 GND 8.53e-19
C10679 VDD.n5131 GND 9.03e-19
C10680 VDD.n5132 GND 0.001706f
C10681 VDD.n5133 GND 0.09638f
C10682 VDD.n5134 GND 0.045561f
C10683 VDD.n5135 GND 0.001706f
C10684 VDD.n5136 GND 8.78e-19
C10685 VDD.n5137 GND 8.53e-19
C10686 VDD.n5138 GND 0.01746f
C10687 VDD.n5139 GND 0.102225f
C10688 VDD.n5140 GND 0.601507f
C10689 VDD.n5141 GND 0.102225f
C10690 VDD.n5142 GND 0.014122f
C10691 VDD.n5143 GND 8.53e-19
C10692 VDD.n5144 GND 8.78e-19
C10693 VDD.n5145 GND 8.78e-19
C10694 VDD.n5146 GND 0.001706f
C10695 VDD.n5147 GND 0.115656f
C10696 VDD.n5148 GND 0.001706f
C10697 VDD.n5149 GND 8.78e-19
C10698 VDD.n5150 GND 8.53e-19
C10699 VDD.n5151 GND 0.010359f
C10700 VDD.n5152 GND 0.010359f
C10701 VDD.n5153 GND 8.53e-19
C10702 VDD.n5154 GND 9.03e-19
C10703 VDD.n5155 GND 0.001706f
C10704 VDD.n5156 GND 0.005257f
C10705 VDD.n5157 GND 0.001706f
C10706 VDD.n5158 GND 0.008303f
C10707 VDD.n5159 GND 0.072346f
C10708 VDD.n5160 GND 1.79982f
C10709 VDD.n5161 GND 0.073151f
C10710 VDD.n5162 GND 0.002244f
C10711 VDD.t448 GND 0.010699f
C10712 VDD.t442 GND 0.010699f
C10713 VDD.n5163 GND 0.022031f
C10714 VDD.n5164 GND 9.03e-19
C10715 VDD.n5165 GND 0.001516f
C10716 VDD.n5166 GND 8.53e-19
C10717 VDD.n5167 GND 0.002454f
C10718 VDD.n5168 GND 0.002363f
C10719 VDD.n5169 GND 8.53e-19
C10720 VDD.n5170 GND 9.03e-19
C10721 VDD.n5171 GND 0.001972f
C10722 VDD.n5172 GND 0.001783f
C10723 VDD.n5173 GND 0.044032f
C10724 VDD.n5174 GND 2.75612f
C10725 VDD.n5175 GND 26.0199f
C10726 VDD.n5176 GND 7.64969f
C10727 VDD.n5177 GND 44.5653f
C10728 VDD.n5180 GND 1.88886f
C10729 VDD.n5182 GND 2.36108f
C10730 VDD.n5183 GND 1.88886f
C10731 VDD.n5187 GND 0.009297f
C10732 VDD.n5188 GND 0.096908f
C10733 VDD.n5189 GND 0.028852f
C10734 VDD.n5190 GND 0.033745f
C10735 VDD.n5191 GND 0.007454f
C10736 VDD.n5192 GND 0.042542f
C10737 VDD.n5193 GND 0.171595f
C10738 VDD.t205 GND 0.13687f
C10739 VDD.n5194 GND 0.04235f
C10740 VDD.n5195 GND 0.04235f
C10741 VDD.n5196 GND 0.118283f
C10742 VDD.n5197 GND 0.003537f
C10743 VDD.n5198 GND 0.018938f
C10744 VDD.n5199 GND 0.010918f
C10745 VDD.t116 GND 0.053019f
C10746 VDD.n5200 GND 0.075161f
C10747 VDD.n5201 GND 0.005291f
C10748 VDD.n5202 GND 0.024537f
C10749 VDD.n5203 GND 0.024537f
C10750 VDD.n5204 GND 0.024537f
C10751 VDD.t485 GND 0.012174f
C10752 VDD.t714 GND 0.012174f
C10753 VDD.n5205 GND 0.036626f
C10754 VDD.n5206 GND 0.076059f
C10755 VDD.t60 GND 0.053019f
C10756 VDD.n5207 GND 0.078027f
C10757 VDD.n5208 GND 0.013734f
C10758 VDD.n5209 GND 0.021265f
C10759 VDD.n5210 GND 0.153284f
C10760 VDD.t59 GND 0.149993f
C10761 VDD.t484 GND 0.076393f
C10762 VDD.n5211 GND 0.050928f
C10763 VDD.t713 GND 0.076393f
C10764 VDD.t115 GND 0.149993f
C10765 VDD.n5212 GND 0.153284f
C10766 VDD.n5213 GND 0.021239f
C10767 VDD.n5214 GND 0.013724f
C10768 VDD.n5215 GND 0.020807f
C10769 VDD.n5216 GND 0.111635f
C10770 VDD.n5217 GND 0.023282f
C10771 VDD.n5218 GND 0.009355f
C10772 VDD.n5219 GND 0.004824f
C10773 VDD.n5220 GND 0.007693f
C10774 VDD.n5221 GND 0.02997f
C10775 VDD.n5222 GND 0.028855f
C10776 VDD.n5223 GND 0.034976f
C10777 VDD.n5224 GND 0.0157f
C10778 VDD.t379 GND 0.101857f
C10779 VDD.t478 GND 0.101857f
C10780 VDD.t55 GND 0.101857f
C10781 VDD.t477 GND 0.101857f
C10782 VDD.t54 GND 0.101857f
C10783 VDD.t480 GND 0.101857f
C10784 VDD.t367 GND 0.101857f
C10785 VDD.t56 GND 0.101857f
C10786 VDD.t380 GND 0.101857f
C10787 VDD.t474 GND 0.101857f
C10788 VDD.t307 GND 0.101857f
C10789 VDD.t42 GND 0.101857f
C10790 VDD.t366 GND 0.101857f
C10791 VDD.t721 GND 0.101857f
C10792 VDD.t365 GND 0.101857f
C10793 VDD.t720 GND 0.101857f
C10794 VDD.t719 GND 0.101857f
C10795 VDD.t716 GND 0.149993f
C10796 VDD.n5225 GND 0.171595f
C10797 VDD.n5226 GND 0.030514f
C10798 VDD.n5227 GND 0.04235f
C10799 VDD.n5228 GND 0.03395f
C10800 VDD.n5229 GND 0.042542f
C10801 VDD.n5230 GND 0.137931f
C10802 VDD.n5231 GND 0.137931f
C10803 VDD.t518 GND 0.13687f
C10804 VDD.t514 GND 0.101857f
C10805 VDD.t451 GND 0.101857f
C10806 VDD.t522 GND 0.101857f
C10807 VDD.t72 GND 0.101857f
C10808 VDD.t472 GND 0.101857f
C10809 VDD.t289 GND 0.101857f
C10810 VDD.t171 GND 0.101857f
C10811 VDD.t192 GND 0.101857f
C10812 VDD.t457 GND 0.149993f
C10813 VDD.t294 GND 0.101857f
C10814 VDD.t456 GND 0.101857f
C10815 VDD.t386 GND 0.101857f
C10816 VDD.t140 GND 0.101857f
C10817 VDD.t515 GND 0.101857f
C10818 VDD.t707 GND 0.101857f
C10819 VDD.t136 GND 0.101857f
C10820 VDD.t137 GND 0.101857f
C10821 VDD.n5232 GND 0.010398f
C10822 VDD.n5233 GND 0.028852f
C10823 VDD.n5234 GND 0.02734f
C10824 VDD.n5235 GND 0.019507f
C10825 VDD.n5236 GND 0.016007f
C10826 VDD.n5237 GND 0.031248f
C10827 VDD.n5238 GND 0.04235f
C10828 VDD.n5239 GND 0.04235f
C10829 VDD.t26 GND 0.101857f
C10830 VDD.n5240 GND 0.04235f
C10831 VDD.n5241 GND 0.004829f
C10832 VDD.n5242 GND 0.009557f
C10833 VDD.n5243 GND 0.018741f
C10834 VDD.n5244 GND 0.037374f
C10835 VDD.n5245 GND 0.131519f
C10836 VDD.n5246 GND 0.009129f
C10837 VDD.n5247 GND 3.57288f
C10838 VDD.n5248 GND 0.02734f
C10839 VDD.n5249 GND 0.010398f
C10840 VDD.n5250 GND 0.04235f
C10841 VDD.n5251 GND 0.04235f
C10842 VDD.n5252 GND 0.04235f
C10843 VDD.n5253 GND 0.137931f
C10844 VDD.n5254 GND 0.009557f
C10845 VDD.n5255 GND 0.028852f
C10846 VDD.n5256 GND 0.009355f
C10847 VDD.n5257 GND 0.04235f
C10848 VDD.n5258 GND 0.04235f
C10849 VDD.n5259 GND 0.010918f
C10850 VDD.t482 GND 0.053019f
C10851 VDD.n5260 GND 0.075161f
C10852 VDD.n5261 GND 0.005291f
C10853 VDD.n5262 GND 0.024537f
C10854 VDD.n5263 GND 0.024537f
C10855 VDD.n5264 GND 0.024537f
C10856 VDD.t554 GND 0.012174f
C10857 VDD.t718 GND 0.012174f
C10858 VDD.n5265 GND 0.036626f
C10859 VDD.n5266 GND 0.076059f
C10860 VDD.t700 GND 0.053019f
C10861 VDD.n5267 GND 0.078027f
C10862 VDD.n5268 GND 0.013734f
C10863 VDD.n5269 GND 0.021265f
C10864 VDD.n5270 GND 0.153284f
C10865 VDD.t699 GND 0.149993f
C10866 VDD.t553 GND 0.076393f
C10867 VDD.n5271 GND 0.050928f
C10868 VDD.t717 GND 0.076393f
C10869 VDD.t481 GND 0.149993f
C10870 VDD.n5272 GND 0.153284f
C10871 VDD.n5273 GND 0.021239f
C10872 VDD.n5274 GND 0.013724f
C10873 VDD.n5275 GND 0.020807f
C10874 VDD.n5276 GND 0.004824f
C10875 VDD.n5277 GND 0.007693f
C10876 VDD.n5278 GND 0.02997f
C10877 VDD.n5279 GND 0.028855f
C10878 VDD.n5280 GND 0.034976f
C10879 VDD.n5281 GND 0.0157f
C10880 VDD.n5282 GND 0.030514f
C10881 VDD.n5283 GND 0.171595f
C10882 VDD.t387 GND 0.149993f
C10883 VDD.t383 GND 0.101857f
C10884 VDD.t328 GND 0.101857f
C10885 VDD.t722 GND 0.101857f
C10886 VDD.t711 GND 0.101857f
C10887 VDD.t697 GND 0.101857f
C10888 VDD.t270 GND 0.101857f
C10889 VDD.t545 GND 0.101857f
C10890 VDD.t209 GND 0.101857f
C10891 VDD.t548 GND 0.13687f
C10892 VDD.t500 GND 0.101857f
C10893 VDD.t372 GND 0.101857f
C10894 VDD.t33 GND 0.101857f
C10895 VDD.t354 GND 0.101857f
C10896 VDD.t467 GND 0.101857f
C10897 VDD.t532 GND 0.101857f
C10898 VDD.t312 GND 0.101857f
C10899 VDD.t191 GND 0.101857f
C10900 VDD.t355 GND 0.101857f
C10901 VDD.n5284 GND 0.04235f
C10902 VDD.n5285 GND 0.042542f
C10903 VDD.n5286 GND 0.03395f
C10904 VDD.n5287 GND 0.018937f
C10905 VDD.n5288 GND 0.043609f
C10906 VDD.n5289 GND 0.004829f
C10907 VDD.n5290 GND 0.007454f
C10908 VDD.n5291 GND 0.028852f
C10909 VDD.n5292 GND 0.028852f
C10910 VDD.n5293 GND 0.043609f
C10911 VDD.n5294 GND 0.018741f
C10912 VDD.n5295 GND 0.033745f
C10913 VDD.n5296 GND 0.042542f
C10914 VDD.n5297 GND 0.137931f
C10915 VDD.t487 GND 0.13687f
C10916 VDD.t486 GND 0.101857f
C10917 VDD.t204 GND 0.101857f
C10918 VDD.t712 GND 0.101857f
C10919 VDD.t206 GND 0.101857f
C10920 VDD.t102 GND 0.101857f
C10921 VDD.t113 GND 0.101857f
C10922 VDD.t114 GND 0.101857f
C10923 VDD.t58 GND 0.101857f
C10924 VDD.t483 GND 0.101857f
C10925 VDD.t460 GND 0.101857f
C10926 VDD.t461 GND 0.101857f
C10927 VDD.t103 GND 0.101857f
C10928 VDD.t117 GND 0.101857f
C10929 VDD.t104 GND 0.101857f
C10930 VDD.t552 GND 0.101857f
C10931 VDD.t57 GND 0.101857f
C10932 VDD.t488 GND 0.101857f
C10933 VDD.t120 GND 0.149993f
C10934 VDD.n5298 GND 0.171595f
C10935 VDD.n5299 GND 0.031248f
C10936 VDD.n5300 GND 0.016007f
C10937 VDD.n5301 GND 0.019507f
C10938 VDD.n5302 GND 59.7783f
C10939 VDD.n5303 GND 14.829801f
C10940 VDD.n5304 GND 1.18054f
C10941 VDD.n5305 GND 1.18054f
C10942 VDD.n5307 GND 1.84102f
C10943 VDD.n5308 GND 1.18201f
C10944 VDD.n5309 GND 19.153f
C10945 VDD.n5310 GND 0.017341f
C10946 VDD.n5311 GND 0.016003f
C10947 VDD.t521 GND 0.001992f
C10948 VDD.t682 GND 0.001992f
C10949 VDD.n5312 GND 0.004276f
C10950 VDD.n5313 GND 0.004876f
C10951 VDD.t688 GND 0.001992f
C10952 VDD.t692 GND 0.001992f
C10953 VDD.n5314 GND 0.004276f
C10954 VDD.n5315 GND 0.004587f
C10955 VDD.n5316 GND 0.003825f
C10956 VDD.t70 GND 0.041005f
C10957 VDD.n5317 GND 0.002318f
C10958 VDD.t463 GND 0.001992f
C10959 VDD.t258 GND 0.001992f
C10960 VDD.n5318 GND 0.004276f
C10961 VDD.n5319 GND 0.006366f
C10962 VDD.t497 GND 0.007944f
C10963 VDD.n5320 GND 0.003825f
C10964 VDD.t491 GND 0.001992f
C10965 VDD.t493 GND 0.001992f
C10966 VDD.n5321 GND 0.004276f
C10967 VDD.n5322 GND 0.00683f
C10968 VDD.n5323 GND 0.006517f
C10969 VDD.n5324 GND 0.002689f
C10970 VDD.n5325 GND 0.001482f
C10971 VDD.t531 GND 0.001992f
C10972 VDD.t525 GND 0.001992f
C10973 VDD.n5326 GND 0.004276f
C10974 VDD.n5327 GND 0.004876f
C10975 VDD.t133 GND 0.007946f
C10976 VDD.n5328 GND 0.00386f
C10977 VDD.t224 GND 0.001992f
C10978 VDD.t291 GND 0.001992f
C10979 VDD.n5329 GND 0.004276f
C10980 VDD.n5330 GND 0.005816f
C10981 VDD.n5331 GND 0.004887f
C10982 VDD.t709 GND 0.006973f
C10983 VDD.n5332 GND 0.006035f
C10984 VDD.t244 GND 0.022412f
C10985 VDD.n5333 GND 0.001167f
C10986 VDD.t281 GND 0.001992f
C10987 VDD.t321 GND 0.001992f
C10988 VDD.n5334 GND 0.004276f
C10989 VDD.n5335 GND 0.004876f
C10990 VDD.n5336 GND 0.006517f
C10991 VDD.t288 GND 0.001992f
C10992 VDD.t186 GND 0.001992f
C10993 VDD.n5337 GND 0.004276f
C10994 VDD.n5338 GND 0.003228f
C10995 VDD.t306 GND 0.007944f
C10996 VDD.n5339 GND 0.011336f
C10997 VDD.t556 GND 0.007505f
C10998 VDD.n5340 GND 0.007735f
C10999 VDD.t118 GND 0.050253f
C11000 VDD.t550 GND 0.02789f
C11001 VDD.t475 GND 0.017099f
C11002 VDD.n5341 GND 7.65e-19
C11003 VDD.t369 GND 0.001992f
C11004 VDD.t304 GND 0.001992f
C11005 VDD.n5342 GND 0.004276f
C11006 VDD.n5343 GND 0.004876f
C11007 VDD.t119 GND 0.007779f
C11008 VDD.t551 GND 0.001992f
C11009 VDD.t476 GND 0.001992f
C11010 VDD.n5344 GND 0.004276f
C11011 VDD.n5345 GND 0.005392f
C11012 VDD.n5346 GND 0.013433f
C11013 VDD.n5347 GND 0.024211f
C11014 VDD.n5348 GND 0.006517f
C11015 VDD.t300 GND 0.001992f
C11016 VDD.t302 GND 0.001992f
C11017 VDD.n5349 GND 0.004276f
C11018 VDD.n5350 GND 0.003825f
C11019 VDD.n5351 GND 0.006517f
C11020 VDD.n5352 GND 0.001894f
C11021 VDD.n5353 GND 0.004876f
C11022 VDD.n5354 GND 0.001279f
C11023 VDD.n5355 GND 0.001982f
C11024 VDD.n5356 GND 0.006517f
C11025 VDD.n5357 GND 0.006517f
C11026 VDD.n5358 GND 0.001342f
C11027 VDD.n5359 GND 0.003693f
C11028 VDD.n5360 GND 0.01207f
C11029 VDD.t368 GND 0.024736f
C11030 VDD.t303 GND 0.02789f
C11031 VDD.t299 GND 0.02789f
C11032 VDD.t301 GND 0.02789f
C11033 VDD.t305 GND 0.02457f
C11034 VDD.t338 GND 0.02789f
C11035 VDD.t185 GND 0.02789f
C11036 VDD.t287 GND 0.02789f
C11037 VDD.t555 GND 0.024404f
C11038 VDD.n5361 GND 0.027337f
C11039 VDD.n5362 GND -3.69e-19
C11040 VDD.n5363 GND 0.003188f
C11041 VDD.n5364 GND 0.004887f
C11042 VDD.n5365 GND 0.006517f
C11043 VDD.n5366 GND 0.006517f
C11044 VDD.n5367 GND 0.001586f
C11045 VDD.n5368 GND 0.004876f
C11046 VDD.n5369 GND 0.001781f
C11047 VDD.t339 GND 0.001992f
C11048 VDD.t245 GND 0.001992f
C11049 VDD.n5370 GND 0.004276f
C11050 VDD.n5371 GND 0.004876f
C11051 VDD.n5372 GND 0.00148f
C11052 VDD.n5373 GND 0.006517f
C11053 VDD.n5374 GND 0.006517f
C11054 VDD.n5375 GND 0.003825f
C11055 VDD.t459 GND 0.007944f
C11056 VDD.n5376 GND 0.011143f
C11057 VDD.n5377 GND 0.001894f
C11058 VDD.n5378 GND 0.006517f
C11059 VDD.n5379 GND 0.006517f
C11060 VDD.n5380 GND 9.41e-19
C11061 VDD.n5381 GND 0.004573f
C11062 VDD.n5382 GND 0.012076f
C11063 VDD.t280 GND 0.019424f
C11064 VDD.t320 GND 0.02789f
C11065 VDD.t458 GND 0.02457f
C11066 VDD.t708 GND 0.030712f
C11067 VDD.t132 GND 0.026396f
C11068 VDD.t290 GND 0.02789f
C11069 VDD.t223 GND 0.019424f
C11070 VDD.n5383 GND 0.012076f
C11071 VDD.n5384 GND 0.004573f
C11072 VDD.n5385 GND 9.53e-19
C11073 VDD.n5386 GND 0.006517f
C11074 VDD.n5387 GND 0.006517f
C11075 VDD.n5388 GND 0.006517f
C11076 VDD.n5389 GND 0.001894f
C11077 VDD.n5390 GND 0.011616f
C11078 VDD.t529 GND 0.007505f
C11079 VDD.n5391 GND 0.008879f
C11080 VDD.n5392 GND 0.001541f
C11081 VDD.n5393 GND 0.004887f
C11082 VDD.n5394 GND 0.006517f
C11083 VDD.n5395 GND 0.006517f
C11084 VDD.t527 GND 0.001992f
C11085 VDD.t495 GND 0.001992f
C11086 VDD.n5396 GND 0.004276f
C11087 VDD.n5397 GND 0.004876f
C11088 VDD.n5398 GND 0.00148f
C11089 VDD.n5399 GND 0.001781f
C11090 VDD.n5400 GND 0.006517f
C11091 VDD.n5401 GND 0.006517f
C11092 VDD.n5402 GND 0.002464f
C11093 VDD.n5403 GND 0.001182f
C11094 VDD.n5404 GND 0.027171f
C11095 VDD.t528 GND 0.014111f
C11096 VDD.t530 GND 0.02789f
C11097 VDD.t524 GND 0.02789f
C11098 VDD.t526 GND 0.02789f
C11099 VDD.t494 GND 0.02789f
C11100 VDD.t490 GND 0.01876f
C11101 VDD.t496 GND 0.02457f
C11102 VDD.t492 GND 0.023076f
C11103 VDD.n5405 GND 0.012064f
C11104 VDD.n5406 GND 0.001237f
C11105 VDD.n5407 GND 3.93e-19
C11106 VDD.n5408 GND 0.006517f
C11107 VDD.n5409 GND 0.006517f
C11108 VDD.n5410 GND 0.002312f
C11109 VDD.n5411 GND 0.011256f
C11110 VDD.t71 GND 0.007586f
C11111 VDD.n5412 GND 0.007772f
C11112 VDD.n5413 GND 0.001116f
C11113 VDD.n5414 GND 0.004887f
C11114 VDD.n5415 GND 0.006517f
C11115 VDD.n5416 GND 0.003896f
C11116 VDD.n5417 GND 0.00148f
C11117 VDD.n5418 GND 0.001743f
C11118 VDD.n5419 GND 0.006517f
C11119 VDD.n5420 GND 0.006517f
C11120 VDD.n5421 GND 0.001664f
C11121 VDD.n5422 GND 0.001045f
C11122 VDD.n5423 GND 0.012064f
C11123 VDD.t462 GND 0.016103f
C11124 VDD.t257 GND 0.02789f
C11125 VDD.t520 GND 0.02789f
C11126 VDD.t681 GND 0.02789f
C11127 VDD.t687 GND 0.02789f
C11128 VDD.t691 GND 0.016767f
C11129 VDD.t546 GND 0.017645f
C11130 VDD.t150 GND 0.027f
C11131 VDD.t685 GND 0.021748f
C11132 VDD.n5424 GND 0.012076f
C11133 VDD.n5425 GND 0.004447f
C11134 VDD.t151 GND 0.006281f
C11135 VDD.n5426 GND 0.004887f
C11136 VDD.t547 GND 0.005799f
C11137 VDD.n5427 GND 0.009833f
C11138 VDD.n5428 GND 0.00386f
C11139 VDD.n5429 GND 0.006517f
C11140 VDD.n5430 GND 0.001681f
C11141 VDD.n5431 GND 0.011335f
C11142 VDD.t686 GND 0.007944f
C11143 VDD.n5432 GND 0.010892f
C11144 VDD.n5433 GND 0.001154f
C11145 VDD.n5434 GND 0.006517f
C11146 VDD.n5435 GND 0.004887f
C11147 VDD.n5436 GND 0.001279f
C11148 VDD.n5437 GND 0.001982f
C11149 VDD.n5438 GND 0.002678f
C11150 VDD.n5439 GND 0.014647f
C11151 VDD.n5440 GND 0.017761f
C11152 VDD.n5441 GND 0.019448f
C11153 VDD.n5442 GND 0.001411f
C11154 VDD.t578 GND 0.001992f
C11155 VDD.t572 GND 0.001992f
C11156 VDD.n5443 GND 0.004276f
C11157 VDD.n5444 GND 0.001393f
C11158 VDD.t576 GND 0.007586f
C11159 VDD.n5445 GND 0.007772f
C11160 VDD.n5446 GND 0.001894f
C11161 VDD.n5447 GND 0.006517f
C11162 VDD.t684 GND 0.001992f
C11163 VDD.t690 GND 0.001992f
C11164 VDD.n5448 GND 0.004276f
C11165 VDD.t696 GND 0.007946f
C11166 VDD.n5449 GND 0.00386f
C11167 VDD.n5450 GND 0.010061f
C11168 VDD.n5451 GND 0.001894f
C11169 VDD.n5452 GND 0.00603f
C11170 VDD.n5453 GND 0.006517f
C11171 VDD.n5454 GND 0.006517f
C11172 VDD.n5455 GND 0.004887f
C11173 VDD.t694 GND 0.006973f
C11174 VDD.n5456 GND 0.006387f
C11175 VDD.n5457 GND 0.001355f
C11176 VDD.n5458 GND 0.004887f
C11177 VDD.n5459 GND 0.006517f
C11178 VDD.n5460 GND 0.004887f
C11179 VDD.n5461 GND 0.004416f
C11180 VDD.t310 GND 0.00858f
C11181 VDD.n5462 GND 9.66e-19
C11182 VDD.t15 GND 0.001992f
C11183 VDD.t382 GND 0.001992f
C11184 VDD.n5463 GND 0.004276f
C11185 VDD.n5464 GND 0.004876f
C11186 VDD.n5465 GND 0.006517f
C11187 VDD.t582 GND 0.007586f
C11188 VDD.t586 GND 0.001992f
C11189 VDD.t588 GND 0.001992f
C11190 VDD.n5466 GND 0.004276f
C11191 VDD.n5467 GND 0.006967f
C11192 VDD.n5468 GND 0.006517f
C11193 VDD.n5469 GND 0.002515f
C11194 VDD.n5470 GND 6.27e-20
C11195 VDD.t277 GND 0.001992f
C11196 VDD.t541 GND 0.001992f
C11197 VDD.n5471 GND 0.004276f
C11198 VDD.n5472 GND 0.004876f
C11199 VDD.n5473 GND 0.006517f
C11200 VDD.t220 GND 0.001992f
C11201 VDD.t135 GND 0.001992f
C11202 VDD.n5474 GND 0.004276f
C11203 VDD.n5475 GND 0.003153f
C11204 VDD.n5476 GND 0.006517f
C11205 VDD.n5477 GND 0.0021f
C11206 VDD.t672 GND 0.001992f
C11207 VDD.t108 GND 0.001992f
C11208 VDD.n5478 GND 0.004276f
C11209 VDD.n5479 GND 0.006827f
C11210 VDD.t239 GND 0.007795f
C11211 VDD.n5480 GND 0.009297f
C11212 VDD.t674 GND 0.007586f
C11213 VDD.n5481 GND 0.007741f
C11214 VDD.n5482 GND 0.006517f
C11215 VDD.t235 GND 0.001992f
C11216 VDD.t237 GND 0.001992f
C11217 VDD.n5483 GND 0.004276f
C11218 VDD.n5484 GND 0.001982f
C11219 VDD.n5485 GND 0.024211f
C11220 VDD.t563 GND 0.077668f
C11221 VDD.t567 GND 0.025287f
C11222 VDD.t569 GND 0.018815f
C11223 VDD.t238 GND 0.022277f
C11224 VDD.t236 GND 0.025287f
C11225 VDD.t234 GND 0.025287f
C11226 VDD.t232 GND 0.025287f
C11227 VDD.t565 GND 0.019116f
C11228 VDD.n5486 GND 0.010777f
C11229 VDD.t568 GND 0.001992f
C11230 VDD.t570 GND 0.001992f
C11231 VDD.n5487 GND 0.004276f
C11232 VDD.t564 GND 0.007779f
C11233 VDD.n5488 GND 0.013433f
C11234 VDD.n5489 GND 0.005392f
C11235 VDD.n5490 GND 0.001041f
C11236 VDD.n5491 GND 0.006452f
C11237 VDD.t566 GND 0.001992f
C11238 VDD.t233 GND 0.001992f
C11239 VDD.n5492 GND 0.004276f
C11240 VDD.n5493 GND 0.004876f
C11241 VDD.n5494 GND 0.001066f
C11242 VDD.n5495 GND 0.006517f
C11243 VDD.n5496 GND 0.006517f
C11244 VDD.n5497 GND 0.006517f
C11245 VDD.n5498 GND 0.001279f
C11246 VDD.n5499 GND 0.004876f
C11247 VDD.n5500 GND 0.002271f
C11248 VDD.n5501 GND 0.003668f
C11249 VDD.n5502 GND 0.003825f
C11250 VDD.n5503 GND 0.006517f
C11251 VDD.t676 GND 0.001992f
C11252 VDD.t670 GND 0.001992f
C11253 VDD.n5504 GND 0.004276f
C11254 VDD.n5505 GND 0.004876f
C11255 VDD.n5506 GND 0.001681f
C11256 VDD.n5507 GND 0.001367f
C11257 VDD.n5508 GND 0.006517f
C11258 VDD.n5509 GND 0.004887f
C11259 VDD.n5510 GND 0.003152f
C11260 VDD.n5511 GND 0.001369f
C11261 VDD.n5512 GND 0.02461f
C11262 VDD.t673 GND 0.038081f
C11263 VDD.t675 GND 0.025287f
C11264 VDD.t669 GND 0.025287f
C11265 VDD.t671 GND 0.017009f
C11266 VDD.t187 GND 0.022277f
C11267 VDD.t134 GND 0.025287f
C11268 VDD.t219 GND 0.025287f
C11269 VDD.t107 GND 0.020922f
C11270 VDD.n5513 GND 0.010762f
C11271 VDD.n5514 GND -9.33e-19
C11272 VDD.n5515 GND 0.004283f
C11273 VDD.n5516 GND 0.006517f
C11274 VDD.n5517 GND 0.006517f
C11275 VDD.n5518 GND 0.006517f
C11276 VDD.n5519 GND 0.001279f
C11277 VDD.n5520 GND 0.004876f
C11278 VDD.n5521 GND 0.002183f
C11279 VDD.t188 GND 0.007795f
C11280 VDD.t353 GND 0.007795f
C11281 VDD.n5522 GND 0.009574f
C11282 VDD.n5523 GND 0.009587f
C11283 VDD.n5524 GND 0.001192f
C11284 VDD.n5525 GND 0.003825f
C11285 VDD.n5526 GND 0.002267f
C11286 VDD.n5527 GND 0.006517f
C11287 VDD.t66 GND 0.001992f
C11288 VDD.t584 GND 0.001992f
C11289 VDD.n5528 GND 0.004276f
C11290 VDD.n5529 GND 0.004876f
C11291 VDD.n5530 GND 0.001982f
C11292 VDD.n5531 GND 0.001279f
C11293 VDD.n5532 GND 0.006517f
C11294 VDD.n5533 GND 0.005879f
C11295 VDD.n5534 GND 0.002145f
C11296 VDD.n5535 GND 0.006452f
C11297 VDD.n5536 GND 0.012282f
C11298 VDD.t352 GND 0.017159f
C11299 VDD.t276 GND 0.025287f
C11300 VDD.t540 GND 0.025287f
C11301 VDD.t65 GND 0.025287f
C11302 VDD.t583 GND 0.023029f
C11303 VDD.t581 GND 0.044252f
C11304 VDD.t587 GND 0.025287f
C11305 VDD.t585 GND 0.014901f
C11306 VDD.n5537 GND 0.010762f
C11307 VDD.n5538 GND 0.001914f
C11308 VDD.n5539 GND 0.002081f
C11309 VDD.n5540 GND 0.006517f
C11310 VDD.n5541 GND 0.006517f
C11311 VDD.n5542 GND 0.001651f
C11312 VDD.n5543 GND 0.001367f
C11313 VDD.n5544 GND 0.007772f
C11314 VDD.t311 GND 0.007795f
C11315 VDD.n5545 GND 0.009612f
C11316 VDD.n5546 GND 0.001442f
C11317 VDD.n5547 GND 0.004887f
C11318 VDD.n5548 GND 0.002267f
C11319 VDD.n5549 GND 0.004179f
C11320 VDD.n5550 GND 0.006517f
C11321 VDD.t173 GND 0.001992f
C11322 VDD.t574 GND 0.001992f
C11323 VDD.n5551 GND 0.004276f
C11324 VDD.n5552 GND 0.004876f
C11325 VDD.n5553 GND 0.001982f
C11326 VDD.n5554 GND 0.001279f
C11327 VDD.n5555 GND 0.006517f
C11328 VDD.n5556 GND 0.005879f
C11329 VDD.n5557 GND 0.001242f
C11330 VDD.n5558 GND 0.006452f
C11331 VDD.n5559 GND 0.010777f
C11332 VDD.t14 GND 0.021223f
C11333 VDD.t381 GND 0.025287f
C11334 VDD.t172 GND 0.025287f
C11335 VDD.t573 GND 0.025287f
C11336 VDD.t577 GND 0.021223f
C11337 VDD.t695 GND 0.023932f
C11338 VDD.t689 GND 0.025287f
C11339 VDD.t683 GND 0.025287f
C11340 VDD.t693 GND 0.050273f
C11341 VDD.t575 GND 0.050273f
C11342 VDD.t571 GND 0.016708f
C11343 VDD.n5560 GND 0.010762f
C11344 VDD.n5561 GND -3.48e-19
C11345 VDD.n5562 GND 0.006095f
C11346 VDD.n5563 GND 0.003529f
C11347 VDD.n5564 GND 0.003099f
C11348 VDD.n5565 GND 0.003652f
C11349 VDD.n5566 GND 0.229687f
C11350 VDD.n5567 GND 2.98545f
C11351 VDD.n5568 GND 0.335437f
C11352 VDD.n5569 GND 0.005467f
C11353 VDD.n5570 GND 0.002367f
C11354 VDD.n5571 GND 8.53e-19
C11355 VDD.n5572 GND 0.00291f
C11356 VDD.n5573 GND 9.03e-19
C11357 VDD.n5574 GND 0.007088f
C11358 VDD.t710 GND 0.00545f
C11359 VDD.n5575 GND 0.002183f
C11360 VDD.n5576 GND 0.001115f
C11361 VDD.n5577 GND 8.53e-19
C11362 VDD.n5578 GND 0.041407f
C11363 VDD.n5579 GND 0.002444f
C11364 VDD.n5580 GND 8.53e-19
C11365 VDD.n5581 GND 9.03e-19
C11366 VDD.n5582 GND 0.00291f
C11367 VDD.n5583 GND 0.006447f
C11368 VDD.n5584 GND 9.03e-19
C11369 VDD.n5585 GND 0.00116f
C11370 VDD.n5586 GND 0.002806f
C11371 VDD.n5587 GND 0.018731f
C11372 VDD.n5588 GND 0.12073f
C11373 VDD.n5589 GND 0.018612f
C11374 VDD.n5590 GND 0.011119f
C11375 VDD.n5591 GND 0.001062f
C11376 VDD.n5592 GND 0.001706f
C11377 VDD.n5594 GND 0.247293f
C11378 VDD.n5595 GND 0.001706f
C11379 VDD.n5596 GND 0.001706f
C11380 VDD.n5598 GND 0.003712f
C11381 VDD.n5599 GND 0.001706f
C11382 VDD.n5600 GND 0.001706f
C11383 VDD.n5601 GND 0.188724f
C11384 VDD.n5602 GND 0.001706f
C11385 VDD.n5603 GND 0.074839f
C11386 VDD.n5604 GND 0.001706f
C11387 VDD.n5605 GND 0.003712f
C11388 VDD.n5606 GND 0.001706f
C11389 VDD.n5607 GND 0.003712f
C11390 VDD.n5608 GND 0.001706f
C11391 VDD.n5609 GND 0.001706f
C11392 VDD.t161 GND 0.073754f
C11393 VDD.n5610 GND 0.001706f
C11394 VDD.n5611 GND 0.001706f
C11395 VDD.n5612 GND 0.147508f
C11396 VDD.n5613 GND 0.001706f
C11397 VDD.n5614 GND 0.001706f
C11398 VDD.n5615 GND 0.003714f
C11399 VDD.n5616 GND 0.001706f
C11400 VDD.n5617 GND 0.001706f
C11401 VDD.n5618 GND 0.001706f
C11402 VDD.n5620 GND 0.001706f
C11403 VDD.n5621 GND 0.001003f
C11404 VDD.n5623 GND 0.001706f
C11405 VDD.n5624 GND 0.001706f
C11406 VDD.n5625 GND 0.001062f
C11407 VDD.n5626 GND 0.001003f
C11408 VDD.n5627 GND 0.001149f
C11409 VDD.n5628 GND 0.001704f
C11410 VDD.n5629 GND 0.001706f
C11411 VDD.n5631 GND 0.001706f
C11412 VDD.n5632 GND 0.001706f
C11413 VDD.n5633 GND 0.001706f
C11414 VDD.n5634 GND 0.001706f
C11415 VDD.n5635 GND 0.001706f
C11416 VDD.n5636 GND 0.001706f
C11417 VDD.n5638 GND 0.001706f
C11418 VDD.n5639 GND 0.003714f
C11419 VDD.n5640 GND 0.003712f
C11420 VDD.n5641 GND 0.003712f
C11421 VDD.n5642 GND 0.001706f
C11422 VDD.n5643 GND 0.001706f
C11423 VDD.n5644 GND 0.001706f
C11424 VDD.n5645 GND 0.001706f
C11425 VDD.n5646 GND 0.001706f
C11426 VDD.n5647 GND 0.001706f
C11427 VDD.t163 GND 0.073754f
C11428 VDD.n5648 GND 0.001706f
C11429 VDD.n5649 GND 0.001706f
C11430 VDD.n5650 GND 0.001706f
C11431 VDD.n5651 GND 0.087854f
C11432 VDD.n5652 GND 0.001706f
C11433 VDD.n5653 GND 0.001706f
C11434 VDD.n5654 GND 0.147508f
C11435 VDD.n5655 GND 0.001706f
C11436 VDD.n5656 GND 0.001706f
C11437 VDD.n5657 GND 0.001706f
C11438 VDD.n5658 GND 0.001706f
C11439 VDD.n5659 GND 0.001706f
C11440 VDD.t200 GND 0.073754f
C11441 VDD.n5660 GND 0.001706f
C11442 VDD.n5661 GND 0.001706f
C11443 VDD.n5662 GND 0.001706f
C11444 VDD.n5663 GND 0.103039f
C11445 VDD.n5664 GND 0.001706f
C11446 VDD.n5665 GND 0.001706f
C11447 VDD.n5666 GND 0.147508f
C11448 VDD.n5667 GND 0.001706f
C11449 VDD.n5668 GND 0.001706f
C11450 VDD.n5669 GND 0.001706f
C11451 VDD.n5670 GND 0.001706f
C11452 VDD.n5671 GND 0.001706f
C11453 VDD.t210 GND 0.073754f
C11454 VDD.n5672 GND 0.001706f
C11455 VDD.n5673 GND 0.001706f
C11456 VDD.n5674 GND 0.001706f
C11457 VDD.n5675 GND 0.118224f
C11458 VDD.n5676 GND 0.001706f
C11459 VDD.n5677 GND 0.001706f
C11460 VDD.n5678 GND 0.147508f
C11461 VDD.n5679 GND 0.001706f
C11462 VDD.n5680 GND 0.001706f
C11463 VDD.n5681 GND 0.001706f
C11464 VDD.n5682 GND 0.001706f
C11465 VDD.n5683 GND 0.001706f
C11466 VDD.t212 GND 0.073754f
C11467 VDD.n5684 GND 0.001706f
C11468 VDD.n5685 GND 0.001706f
C11469 VDD.n5686 GND 0.001706f
C11470 VDD.n5687 GND 0.133408f
C11471 VDD.n5688 GND 0.001706f
C11472 VDD.n5689 GND 0.001706f
C11473 VDD.n5690 GND 0.146424f
C11474 VDD.n5691 GND 0.001706f
C11475 VDD.n5692 GND 0.001706f
C11476 VDD.n5693 GND 0.001706f
C11477 VDD.t198 GND 0.073754f
C11478 VDD.n5694 GND 0.001706f
C11479 VDD.n5695 GND 0.001706f
C11480 VDD.n5696 GND 0.147508f
C11481 VDD.n5697 GND 0.001706f
C11482 VDD.n5698 GND 0.003714f
C11483 VDD.n5699 GND 0.003714f
C11484 VDD.n5700 GND 0.003712f
C11485 VDD.n5701 GND 0.003712f
C11486 VDD.n5702 GND 0.229939f
C11487 VDD.n5703 GND 0.003714f
C11488 VDD.n5704 GND 0.001706f
C11489 VDD.n5705 GND 0.001706f
C11490 VDD.n5706 GND 0.001704f
C11491 VDD.n5707 GND 0.001706f
C11492 VDD.n5708 GND 0.001062f
C11493 VDD.t211 GND 0.010699f
C11494 VDD.t213 GND 0.010699f
C11495 VDD.n5709 GND 0.032273f
C11496 VDD.n5710 GND 0.107301f
C11497 VDD.n5711 GND 0.005784f
C11498 VDD.n5712 GND 0.005969f
C11499 VDD.n5713 GND 8.53e-19
C11500 VDD.n5714 GND 0.002183f
C11501 VDD.n5715 GND 8.78e-19
C11502 VDD.n5716 GND 0.004516f
C11503 VDD.n5717 GND 0.004516f
C11504 VDD.n5718 GND 0.001062f
C11505 VDD.t199 GND 0.001455f
C11506 VDD.n5719 GND 0.005656f
C11507 VDD.n5720 GND 8.78e-19
C11508 VDD.n5721 GND 0.001115f
C11509 VDD.n5722 GND 0.00636f
C11510 VDD.n5723 GND 0.041968f
C11511 VDD.n5724 GND 0.001022f
C11512 VDD.n5725 GND 0.001706f
C11513 VDD.n5726 GND 0.001706f
C11514 VDD.n5727 GND 0.001706f
C11515 VDD.n5729 GND 0.001706f
C11516 VDD.n5730 GND 0.001706f
C11517 VDD.n5731 GND 0.001706f
C11518 VDD.n5732 GND 0.001706f
C11519 VDD.n5733 GND 0.001706f
C11520 VDD.n5735 GND 0.001706f
C11521 VDD.n5737 GND 0.001706f
C11522 VDD.n5738 GND 0.001706f
C11523 VDD.n5739 GND 0.00173f
C11524 VDD.n5740 GND 0.002023f
C11525 VDD.n5741 GND 0.001706f
C11526 VDD.n5743 GND 0.001706f
C11527 VDD.n5744 GND 0.001706f
C11528 VDD.n5745 GND 0.001706f
C11529 VDD.n5746 GND 0.001706f
C11530 VDD.n5747 GND 0.003714f
C11531 VDD.n5748 GND 0.001706f
C11532 VDD.n5749 GND 0.001706f
C11533 VDD.n5750 GND 0.001706f
C11534 VDD.n5751 GND 0.001062f
C11535 VDD.n5752 GND 0.004516f
C11536 VDD.n5753 GND 0.005656f
C11537 VDD.n5754 GND 8.53e-19
C11538 VDD.n5755 GND 0.006434f
C11539 VDD.n5756 GND 9.03e-19
C11540 VDD.t164 GND 0.010699f
C11541 VDD.t201 GND 0.010699f
C11542 VDD.n5757 GND 0.032273f
C11543 VDD.n5758 GND 0.229486f
C11544 VDD.n5759 GND 0.586149f
C11545 VDD.n5760 GND 0.107744f
C11546 VDD.n5761 GND 0.030806f
C11547 VDD.n5762 GND 0.025832f
C11548 VDD.n5763 GND 0.005784f
C11549 VDD.n5764 GND 0.001162f
C11550 VDD.n5765 GND 0.0023f
C11551 VDD.n5766 GND 0.004516f
C11552 VDD.n5767 GND 0.00173f
C11553 VDD.n5768 GND 0.001706f
C11554 VDD.n5769 GND 0.001706f
C11555 VDD.n5770 GND 0.001706f
C11556 VDD.n5771 GND 0.003714f
C11557 VDD.n5772 GND 0.003714f
C11558 VDD.n5774 GND 0.001706f
C11559 VDD.n5776 GND 0.001706f
C11560 VDD.n5777 GND 0.001706f
C11561 VDD.n5778 GND 0.001706f
C11562 VDD.n5779 GND 0.001706f
C11563 VDD.n5780 GND 0.001706f
C11564 VDD.n5782 GND 0.001706f
C11565 VDD.n5783 GND 0.001706f
C11566 VDD.n5784 GND 0.001706f
C11567 VDD.n5785 GND 0.004516f
C11568 VDD.n5786 GND 0.001003f
C11569 VDD.n5788 GND 0.001706f
C11570 VDD.n5790 GND 0.001706f
C11571 VDD.n5791 GND 0.001062f
C11572 VDD.n5792 GND 0.002023f
C11573 VDD.n5793 GND 0.004516f
C11574 VDD.n5794 GND 0.005969f
C11575 VDD.n5795 GND 8.53e-19
C11576 VDD.n5796 GND 9.03e-19
C11577 VDD.n5797 GND 0.00291f
C11578 VDD.t162 GND 0.001455f
C11579 VDD.n5798 GND 0.002183f
C11580 VDD.n5799 GND 8.78e-19
C11581 VDD.n5800 GND 8.78e-19
C11582 VDD.n5801 GND 0.001115f
C11583 VDD.n5802 GND 0.00636f
C11584 VDD.n5803 GND 0.041968f
C11585 VDD.n5804 GND 0.001022f
C11586 VDD.n5805 GND 0.001645f
C11587 VDD.n5806 GND 0.001706f
C11588 VDD.n5807 GND 0.001706f
C11589 VDD.n5809 GND 0.001706f
C11590 VDD.n5811 GND 0.001706f
C11591 VDD.n5812 GND 0.001706f
C11592 VDD.n5813 GND 0.001706f
C11593 VDD.n5814 GND 0.001706f
C11594 VDD.n5815 GND 0.001706f
C11595 VDD.n5817 GND 0.003714f
C11596 VDD.n5818 GND 0.003712f
C11597 VDD.n5819 GND 0.003712f
C11598 VDD.n5820 GND 0.001706f
C11599 VDD.n5821 GND 0.001706f
C11600 VDD.n5822 GND 0.001706f
C11601 VDD.n5823 GND 0.001706f
C11602 VDD.n5824 GND 0.001706f
C11603 VDD.n5825 GND 0.001706f
C11604 VDD.n5826 GND 0.001706f
C11605 VDD.n5827 GND 0.001706f
C11606 VDD.n5828 GND 0.001706f
C11607 VDD.n5829 GND 0.001706f
C11608 VDD.n5830 GND 0.001706f
C11609 VDD.n5831 GND 0.001706f
C11610 VDD.n5832 GND 0.001706f
C11611 VDD.n5833 GND 0.001706f
C11612 VDD.n5834 GND 0.001706f
C11613 VDD.n5835 GND 0.001706f
C11614 VDD.n5836 GND 0.001706f
C11615 VDD.n5837 GND 0.001706f
C11616 VDD.n5838 GND 0.001706f
C11617 VDD.n5839 GND 0.001706f
C11618 VDD.n5840 GND 0.001706f
C11619 VDD.n5841 GND 0.001706f
C11620 VDD.n5842 GND 0.001706f
C11621 VDD.n5843 GND 0.001706f
C11622 VDD.n5844 GND 0.001706f
C11623 VDD.n5845 GND 0.001706f
C11624 VDD.n5846 GND 0.001706f
C11625 VDD.n5847 GND 0.001706f
C11626 VDD.n5848 GND 0.001706f
C11627 VDD.n5849 GND 0.001706f
C11628 VDD.n5850 GND 0.001706f
C11629 VDD.n5851 GND 0.001706f
C11630 VDD.n5852 GND 0.001706f
C11631 VDD.n5853 GND 0.003712f
C11632 VDD.n5855 GND 0.003714f
C11633 VDD.n5856 GND 0.003714f
C11634 VDD.n5857 GND 0.001706f
C11635 VDD.n5858 GND 0.001706f
C11636 VDD.n5859 GND 0.001706f
C11637 VDD.n5861 GND 0.001706f
C11638 VDD.n5863 GND 0.001706f
C11639 VDD.n5864 GND 0.001706f
C11640 VDD.n5865 GND 0.001706f
C11641 VDD.n5866 GND 0.001645f
C11642 VDD.n5867 GND 0.001706f
C11643 VDD.n5869 GND 0.001706f
C11644 VDD.n5870 GND 0.001062f
C11645 VDD.n5871 GND 0.001003f
C11646 VDD.n5872 GND 0.004516f
C11647 VDD.n5873 GND 0.004516f
C11648 VDD.n5874 GND 8.53e-19
C11649 VDD.n5875 GND 9.03e-19
C11650 VDD.n5876 GND 0.00291f
C11651 VDD.n5877 GND 0.006434f
C11652 VDD.n5878 GND 9.03e-19
C11653 VDD.n5879 GND 0.001162f
C11654 VDD.n5880 GND 0.0023f
C11655 VDD.n5881 GND 0.025832f
C11656 VDD.n5882 GND 0.033011f
C11657 VDD.n5883 GND 0.172693f
C11658 VDD.t356 GND 0.010699f
C11659 VDD.t473 GND 0.010699f
C11660 VDD.n5884 GND 0.032325f
C11661 VDD.n5885 GND 0.102342f
C11662 VDD.t278 GND 0.010699f
C11663 VDD.t362 GND 0.010699f
C11664 VDD.n5886 GND 0.032325f
C11665 VDD.n5887 GND 0.102988f
C11666 VDD.n5888 GND 0.005467f
C11667 VDD.n5889 GND 0.002367f
C11668 VDD.n5890 GND 8.53e-19
C11669 VDD.n5891 GND 0.00291f
C11670 VDD.n5892 GND 9.03e-19
C11671 VDD.n5893 GND 0.007088f
C11672 VDD.t698 GND 0.00545f
C11673 VDD.n5894 GND 0.002183f
C11674 VDD.n5895 GND 0.001115f
C11675 VDD.n5896 GND 8.53e-19
C11676 VDD.n5897 GND 0.041407f
C11677 VDD.n5898 GND 0.002444f
C11678 VDD.n5899 GND 8.53e-19
C11679 VDD.n5900 GND 9.03e-19
C11680 VDD.n5901 GND 0.00291f
C11681 VDD.n5902 GND 0.006447f
C11682 VDD.n5903 GND 9.03e-19
C11683 VDD.n5904 GND 0.00116f
C11684 VDD.n5905 GND 0.002806f
C11685 VDD.n5906 GND 0.018731f
C11686 VDD.n5907 GND 0.052956f
C11687 VDD.n5908 GND 0.192513f
C11688 VDD.n5909 GND 0.031168f
C11689 VDD.n5910 GND 0.017532f
C11690 VDD.n5911 GND 0.00102f
C11691 VDD.n5913 GND 0.001706f
C11692 VDD.n5914 GND 0.001706f
C11693 VDD.n5915 GND 0.001706f
C11694 VDD.n5916 GND 0.001706f
C11695 VDD.n5917 GND 0.001706f
C11696 VDD.n5918 GND 0.001706f
C11697 VDD.n5919 GND 0.001706f
C11698 VDD.n5920 GND 0.001706f
C11699 VDD.n5921 GND 0.001706f
C11700 VDD.n5922 GND 0.001706f
C11701 VDD.n5923 GND 0.001706f
C11702 VDD.n5924 GND 0.001706f
C11703 VDD.n5925 GND 0.001706f
C11704 VDD.n5926 GND 0.001706f
C11705 VDD.n5927 GND 0.001706f
C11706 VDD.n5928 GND 0.001706f
C11707 VDD.n5929 GND 0.001706f
C11708 VDD.n5930 GND 0.001706f
C11709 VDD.n5931 GND 0.001706f
C11710 VDD.n5932 GND 0.001706f
C11711 VDD.n5933 GND 0.001706f
C11712 VDD.n5934 GND 0.001706f
C11713 VDD.n5935 GND 0.001706f
C11714 VDD.n5936 GND 0.001706f
C11715 VDD.n5937 GND 0.001706f
C11716 VDD.n5938 GND 0.001706f
C11717 VDD.n5939 GND 0.001706f
C11718 VDD.n5940 GND 0.001706f
C11719 VDD.n5941 GND 0.001706f
C11720 VDD.n5942 GND 0.001706f
C11721 VDD.n5943 GND 0.001706f
C11722 VDD.n5944 GND 0.001706f
C11723 VDD.n5945 GND 0.003712f
C11724 VDD.n5946 GND 0.003714f
C11725 VDD.n5947 GND 0.003714f
C11726 VDD.n5949 GND 0.001706f
C11727 VDD.n5950 GND 0.001706f
C11728 VDD.n5951 GND 0.001706f
C11729 VDD.n5952 GND 0.001706f
C11730 VDD.n5953 GND 0.001706f
C11731 VDD.n5955 GND 0.001706f
C11732 VDD.n5956 GND 0.001706f
C11733 VDD.n5957 GND 0.001706f
C11734 VDD.n5958 GND 0.001547f
C11735 VDD.n5959 GND 0.001706f
C11736 VDD.n5961 GND 0.001706f
C11737 VDD.n5962 GND 0.001062f
C11738 VDD.n5963 GND 0.001003f
C11739 VDD.n5964 GND 0.011119f
C11740 VDD.n5965 GND 0.018664f
C11741 VDD.n5966 GND 0.001003f
C11742 VDD.n5967 GND 0.001149f
C11743 VDD.n5968 GND 0.001706f
C11744 VDD.n5970 GND 0.001706f
C11745 VDD.n5972 GND 0.001706f
C11746 VDD.n5973 GND 0.001706f
C11747 VDD.n5974 GND 0.001706f
C11748 VDD.n5975 GND 0.001706f
C11749 VDD.n5976 GND 0.001706f
C11750 VDD.n5978 GND 0.001706f
C11751 VDD.n5980 GND 0.001706f
C11752 VDD.n5981 GND 0.001706f
C11753 VDD.n5982 GND 0.003714f
C11754 VDD.n5983 GND 0.003712f
C11755 VDD.n5984 GND 0.003712f
C11756 VDD.n5985 GND 0.188724f
C11757 VDD.n5986 GND 0.003712f
C11758 VDD.n5987 GND 0.003712f
C11759 VDD.n5988 GND 0.001706f
C11760 VDD.n5989 GND 0.001706f
C11761 VDD.n5990 GND 0.001706f
C11762 VDD.n5991 GND 0.074839f
C11763 VDD.n5992 GND 0.001706f
C11764 VDD.n5993 GND 0.001706f
C11765 VDD.n5994 GND 0.001706f
C11766 VDD.n5995 GND 0.001706f
C11767 VDD.n5996 GND 0.001706f
C11768 VDD.n5997 GND 0.147508f
C11769 VDD.n5998 GND 0.001706f
C11770 VDD.n5999 GND 0.001706f
C11771 VDD.n6000 GND 0.001706f
C11772 VDD.n6001 GND 0.001706f
C11773 VDD.n6002 GND 0.001706f
C11774 VDD.n6003 GND 0.087854f
C11775 VDD.n6004 GND 0.001706f
C11776 VDD.n6005 GND 0.001706f
C11777 VDD.n6006 GND 0.001706f
C11778 VDD.n6007 GND 0.001706f
C11779 VDD.n6008 GND 0.001706f
C11780 VDD.n6009 GND 0.147508f
C11781 VDD.n6010 GND 0.001706f
C11782 VDD.n6011 GND 0.001706f
C11783 VDD.n6012 GND 0.001706f
C11784 VDD.n6013 GND 0.001706f
C11785 VDD.n6014 GND 0.001706f
C11786 VDD.n6015 GND 0.103039f
C11787 VDD.n6016 GND 0.001706f
C11788 VDD.n6017 GND 0.001706f
C11789 VDD.n6018 GND 0.001706f
C11790 VDD.n6019 GND 0.001706f
C11791 VDD.n6020 GND 0.001706f
C11792 VDD.n6021 GND 0.147508f
C11793 VDD.n6022 GND 0.001706f
C11794 VDD.n6023 GND 0.001706f
C11795 VDD.n6024 GND 0.001706f
C11796 VDD.n6025 GND 0.001706f
C11797 VDD.n6026 GND 0.001706f
C11798 VDD.n6027 GND 0.118224f
C11799 VDD.n6028 GND 0.001706f
C11800 VDD.n6029 GND 0.001706f
C11801 VDD.n6030 GND 0.001706f
C11802 VDD.n6031 GND 0.001706f
C11803 VDD.n6032 GND 0.001706f
C11804 VDD.n6033 GND 0.147508f
C11805 VDD.n6034 GND 0.001706f
C11806 VDD.n6035 GND 0.001706f
C11807 VDD.n6036 GND 0.001706f
C11808 VDD.n6037 GND 0.001706f
C11809 VDD.n6038 GND 0.001706f
C11810 VDD.n6039 GND 0.133408f
C11811 VDD.n6040 GND 0.001706f
C11812 VDD.n6041 GND 0.001706f
C11813 VDD.n6042 GND 0.001706f
C11814 VDD.n6043 GND 0.001706f
C11815 VDD.n6044 GND 0.001706f
C11816 VDD.n6045 GND 0.146424f
C11817 VDD.n6046 GND 0.001706f
C11818 VDD.n6047 GND 0.001706f
C11819 VDD.n6048 GND 0.001706f
C11820 VDD.n6049 GND 0.001706f
C11821 VDD.n6050 GND 0.001706f
C11822 VDD.n6051 GND 0.147508f
C11823 VDD.n6052 GND 0.001706f
C11824 VDD.n6053 GND 0.001706f
C11825 VDD.n6054 GND 0.003712f
C11826 VDD.n6055 GND 0.003714f
C11827 VDD.n6056 GND 0.003714f
C11828 VDD.n6058 GND 0.001706f
C11829 VDD.n6059 GND 0.001706f
C11830 VDD.n6060 GND 0.001706f
C11831 VDD.n6061 GND 0.001706f
C11832 VDD.n6062 GND 0.001706f
C11833 VDD.n6063 GND 0.001706f
C11834 VDD.n6065 GND 0.001706f
C11835 VDD.n6066 GND 0.001706f
C11836 VDD.n6067 GND 0.001547f
C11837 VDD.n6068 GND 0.00102f
C11838 VDD.n6069 GND 0.017479f
C11839 VDD.n6070 GND 3.28559f
C11840 VDD.n6071 GND 21.312302f
C11841 VDD.n6072 GND 0.007272f
C11842 VDD.n6073 GND 0.007272f
C11843 VDD.n6074 GND 0.002244f
C11844 VDD.t279 GND 0.010699f
C11845 VDD.t489 GND 0.010699f
C11846 VDD.n6075 GND 0.022031f
C11847 VDD.n6076 GND 9.03e-19
C11848 VDD.n6077 GND 0.001516f
C11849 VDD.n6078 GND 8.53e-19
C11850 VDD.n6079 GND 0.002454f
C11851 VDD.n6080 GND 0.002363f
C11852 VDD.n6081 GND 8.53e-19
C11853 VDD.n6082 GND 9.03e-19
C11854 VDD.n6083 GND 0.001972f
C11855 VDD.n6084 GND 0.001783f
C11856 VDD.n6085 GND 0.044032f
C11857 VDD.n6086 GND 0.05786f
C11858 VDD.n6087 GND 0.072213f
C11859 VDD.n6088 GND 0.007272f
C11860 VDD.n6089 GND 0.007272f
C11861 VDD.n6090 GND 0.002244f
C11862 VDD.n6091 GND 0.002384f
C11863 VDD.n6092 GND 9.03e-19
C11864 VDD.n6093 GND 8.53e-19
C11865 VDD.n6094 GND 0.005733f
C11866 VDD.n6095 GND 9.03e-19
C11867 VDD.n6096 GND 0.00263f
C11868 VDD.n6097 GND 8.53e-19
C11869 VDD.n6098 GND 0.002454f
C11870 VDD.n6099 GND 0.002363f
C11871 VDD.n6100 GND 8.53e-19
C11872 VDD.n6101 GND 8.53e-19
C11873 VDD.n6102 GND 9.03e-19
C11874 VDD.n6103 GND 0.00291f
C11875 VDD.n6104 GND 0.00291f
C11876 VDD.n6105 GND 0.002183f
C11877 VDD.n6106 GND 0.001115f
C11878 VDD.t153 GND 0.00545f
C11879 VDD.n6107 GND 0.007088f
C11880 VDD.n6108 GND 0.041407f
C11881 VDD.n6109 GND 8.53e-19
C11882 VDD.n6110 GND 9.03e-19
C11883 VDD.n6111 GND 0.00291f
C11884 VDD.n6112 GND 0.00291f
C11885 VDD.n6113 GND 9.03e-19
C11886 VDD.n6114 GND 8.53e-19
C11887 VDD.n6115 GND 0.002437f
C11888 VDD.n6116 GND 0.004543f
C11889 VDD.n6117 GND 0.047272f
C11890 VDD.n6118 GND 0.002244f
C11891 VDD.t260 GND 0.010699f
C11892 VDD.t315 GND 0.010699f
C11893 VDD.n6119 GND 0.022031f
C11894 VDD.n6120 GND 9.03e-19
C11895 VDD.n6121 GND 0.001516f
C11896 VDD.n6122 GND 8.53e-19
C11897 VDD.n6123 GND 0.002454f
C11898 VDD.n6124 GND 0.002363f
C11899 VDD.n6125 GND 8.53e-19
C11900 VDD.n6126 GND 9.03e-19
C11901 VDD.n6127 GND 0.001972f
C11902 VDD.n6128 GND 0.001783f
C11903 VDD.n6129 GND 0.044032f
C11904 VDD.n6130 GND 0.05786f
C11905 VDD.n6131 GND 0.069098f
C11906 VDD.n6132 GND 0.043713f
C11907 VDD.n6133 GND 0.001512f
C11908 VDD.n6134 GND 0.002407f
C11909 VDD.n6135 GND 8.53e-19
C11910 VDD.t331 GND 0.010699f
C11911 VDD.n6136 GND 0.001985f
C11912 VDD.n6137 GND 0.002355f
C11913 VDD.n6138 GND 0.001972f
C11914 VDD.n6139 GND 9.03e-19
C11915 VDD.t261 GND 0.010699f
C11916 VDD.n6140 GND 0.022036f
C11917 VDD.n6141 GND 9.03e-19
C11918 VDD.n6142 GND 8.53e-19
C11919 VDD.n6143 GND 0.002417f
C11920 VDD.n6144 GND 0.007268f
C11921 VDD.n6145 GND 0.065607f
C11922 VDD.n6146 GND 0.06968f
C11923 VDD.n6147 GND 0.043713f
C11924 VDD.n6148 GND 0.004453f
C11925 VDD.n6149 GND 0.002626f
C11926 VDD.n6150 GND 0.002407f
C11927 VDD.n6151 GND 8.53e-19
C11928 VDD.n6152 GND 0.00291f
C11929 VDD.n6153 GND 9.03e-19
C11930 VDD.n6154 GND 0.041407f
C11931 VDD.n6155 GND 8.53e-19
C11932 VDD.n6156 GND 0.00291f
C11933 VDD.t680 GND 0.00545f
C11934 VDD.n6157 GND 0.007088f
C11935 VDD.n6158 GND 0.001115f
C11936 VDD.n6159 GND 0.002183f
C11937 VDD.n6160 GND 0.00291f
C11938 VDD.n6161 GND 9.03e-19
C11939 VDD.n6162 GND 8.53e-19
C11940 VDD.n6163 GND 0.002444f
C11941 VDD.n6164 GND 0.002355f
C11942 VDD.n6165 GND 8.53e-19
C11943 VDD.n6166 GND 9.03e-19
C11944 VDD.n6167 GND 0.002355f
C11945 VDD.n6168 GND 8.53e-19
C11946 VDD.n6169 GND 9.03e-19
C11947 VDD.n6170 GND 0.00291f
C11948 VDD.n6171 GND 0.005733f
C11949 VDD.n6172 GND 9.03e-19
C11950 VDD.n6173 GND 8.53e-19
C11951 VDD.n6174 GND 0.002417f
C11952 VDD.n6175 GND 0.007268f
C11953 VDD.n6176 GND 0.047272f
C11954 VDD.n6177 GND 0.001512f
C11955 VDD.n6178 GND 0.002407f
C11956 VDD.n6179 GND 8.53e-19
C11957 VDD.t23 GND 0.010699f
C11958 VDD.n6180 GND 0.001985f
C11959 VDD.n6181 GND 0.002355f
C11960 VDD.n6182 GND 0.001972f
C11961 VDD.n6183 GND 9.03e-19
C11962 VDD.t479 GND 0.010699f
C11963 VDD.n6184 GND 0.022036f
C11964 VDD.n6185 GND 9.03e-19
C11965 VDD.n6186 GND 8.53e-19
C11966 VDD.n6187 GND 0.002417f
C11967 VDD.n6188 GND 0.007268f
C11968 VDD.n6189 GND 0.05786f
C11969 VDD.n6190 GND 0.068374f
C11970 VDD.n6191 GND 0.043713f
C11971 VDD.n6192 GND 0.001512f
C11972 VDD.n6193 GND 0.002407f
C11973 VDD.n6194 GND 8.53e-19
C11974 VDD.t39 GND 0.010699f
C11975 VDD.n6195 GND 0.001985f
C11976 VDD.n6196 GND 0.002355f
C11977 VDD.n6197 GND 0.001972f
C11978 VDD.n6198 GND 9.03e-19
C11979 VDD.t44 GND 0.010699f
C11980 VDD.n6199 GND 0.022036f
C11981 VDD.n6200 GND 9.03e-19
C11982 VDD.n6201 GND 8.53e-19
C11983 VDD.n6202 GND 0.002417f
C11984 VDD.n6203 GND 0.007268f
C11985 VDD.n6204 GND 0.05786f
C11986 VDD.n6205 GND 0.043713f
C11987 VDD.n6206 GND 0.001512f
C11988 VDD.n6207 GND 0.002407f
C11989 VDD.n6208 GND 8.53e-19
C11990 VDD.t340 GND 0.010699f
C11991 VDD.n6209 GND 0.001985f
C11992 VDD.n6210 GND 0.002355f
C11993 VDD.n6211 GND 0.001972f
C11994 VDD.n6212 GND 9.03e-19
C11995 VDD.t143 GND 0.010699f
C11996 VDD.n6213 GND 0.022036f
C11997 VDD.n6214 GND 9.03e-19
C11998 VDD.n6215 GND 8.53e-19
C11999 VDD.n6216 GND 0.002417f
C12000 VDD.n6217 GND 0.007268f
C12001 VDD.n6218 GND 0.075015f
C12002 VDD.n6219 GND 0.043713f
C12003 VDD.n6220 GND 0.001512f
C12004 VDD.n6221 GND 0.002407f
C12005 VDD.n6222 GND 8.53e-19
C12006 VDD.t45 GND 0.010699f
C12007 VDD.n6223 GND 0.001985f
C12008 VDD.n6224 GND 0.002355f
C12009 VDD.n6225 GND 0.001972f
C12010 VDD.n6226 GND 9.03e-19
C12011 VDD.t263 GND 0.010699f
C12012 VDD.n6227 GND 0.022036f
C12013 VDD.n6228 GND 9.03e-19
C12014 VDD.n6229 GND 8.53e-19
C12015 VDD.n6230 GND 0.002417f
C12016 VDD.n6231 GND 0.007268f
C12017 VDD.n6232 GND 0.075015f
C12018 VDD.n6233 GND 0.043713f
C12019 VDD.n6234 GND 0.001512f
C12020 VDD.n6235 GND 0.002407f
C12021 VDD.n6236 GND 8.53e-19
C12022 VDD.t231 GND 0.010699f
C12023 VDD.n6237 GND 0.001985f
C12024 VDD.n6238 GND 0.002355f
C12025 VDD.n6239 GND 0.001972f
C12026 VDD.n6240 GND 9.03e-19
C12027 VDD.t49 GND 0.010699f
C12028 VDD.n6241 GND 0.022036f
C12029 VDD.n6242 GND 9.03e-19
C12030 VDD.n6243 GND 8.53e-19
C12031 VDD.n6244 GND 0.002417f
C12032 VDD.n6245 GND 0.007268f
C12033 VDD.n6246 GND 0.05786f
C12034 VDD.n6247 GND 0.043713f
C12035 VDD.n6248 GND 0.043713f
C12036 VDD.n6249 GND 0.043713f
C12037 VDD.n6250 GND 0.043713f
C12038 VDD.n6251 GND 0.001512f
C12039 VDD.n6252 GND 0.002407f
C12040 VDD.n6253 GND 8.53e-19
C12041 VDD.t47 GND 0.010699f
C12042 VDD.n6254 GND 0.001985f
C12043 VDD.n6255 GND 0.002355f
C12044 VDD.n6256 GND 0.001972f
C12045 VDD.n6257 GND 9.03e-19
C12046 VDD.t313 GND 0.010699f
C12047 VDD.n6258 GND 0.022036f
C12048 VDD.n6259 GND 9.03e-19
C12049 VDD.n6260 GND 8.53e-19
C12050 VDD.n6261 GND 0.002417f
C12051 VDD.n6262 GND 0.007268f
C12052 VDD.n6263 GND 0.05786f
C12053 VDD.n6264 GND 0.001512f
C12054 VDD.n6265 GND 0.002407f
C12055 VDD.n6266 GND 8.53e-19
C12056 VDD.t166 GND 0.010699f
C12057 VDD.n6267 GND 0.001985f
C12058 VDD.n6268 GND 0.002355f
C12059 VDD.n6269 GND 0.001972f
C12060 VDD.n6270 GND 9.03e-19
C12061 VDD.t217 GND 0.010699f
C12062 VDD.n6271 GND 0.022036f
C12063 VDD.n6272 GND 9.03e-19
C12064 VDD.n6273 GND 8.53e-19
C12065 VDD.n6274 GND 0.002417f
C12066 VDD.n6275 GND 0.007268f
C12067 VDD.n6276 GND 0.076121f
C12068 VDD.n6277 GND 0.001512f
C12069 VDD.n6278 GND 0.002407f
C12070 VDD.n6279 GND 8.53e-19
C12071 VDD.t679 GND 0.010699f
C12072 VDD.n6280 GND 0.001985f
C12073 VDD.n6281 GND 0.002355f
C12074 VDD.n6282 GND 0.001972f
C12075 VDD.n6283 GND 9.03e-19
C12076 VDD.t511 GND 0.010699f
C12077 VDD.n6284 GND 0.022036f
C12078 VDD.n6285 GND 9.03e-19
C12079 VDD.n6286 GND 8.53e-19
C12080 VDD.n6287 GND 0.002417f
C12081 VDD.n6288 GND 0.007268f
C12082 VDD.n6289 GND 0.075015f
C12083 VDD.n6290 GND 0.001512f
C12084 VDD.n6291 GND 0.002407f
C12085 VDD.n6292 GND 8.53e-19
C12086 VDD.t275 GND 0.010699f
C12087 VDD.n6293 GND 0.001985f
C12088 VDD.n6294 GND 0.002355f
C12089 VDD.n6295 GND 0.001972f
C12090 VDD.n6296 GND 9.03e-19
C12091 VDD.t677 GND 0.010699f
C12092 VDD.n6297 GND 0.022036f
C12093 VDD.n6298 GND 9.03e-19
C12094 VDD.n6299 GND 8.53e-19
C12095 VDD.n6300 GND 0.002417f
C12096 VDD.n6301 GND 0.007268f
C12097 VDD.n6302 GND 0.05786f
C12098 VDD.n6303 GND 0.060777f
C12099 VDD.n6304 GND 1.36913f
C12100 VDD.n6305 GND 0.007272f
C12101 VDD.n6306 GND 0.002244f
C12102 VDD.t145 GND 0.010699f
C12103 VDD.t3 GND 0.010699f
C12104 VDD.n6307 GND 0.022031f
C12105 VDD.n6308 GND 9.03e-19
C12106 VDD.n6309 GND 0.001516f
C12107 VDD.n6310 GND 8.53e-19
C12108 VDD.n6311 GND 0.002454f
C12109 VDD.n6312 GND 0.002363f
C12110 VDD.n6313 GND 8.53e-19
C12111 VDD.n6314 GND 9.03e-19
C12112 VDD.n6315 GND 0.001972f
C12113 VDD.n6316 GND 0.001783f
C12114 VDD.n6317 GND 0.044032f
C12115 VDD.n6318 GND 0.076121f
C12116 VDD.n6319 GND 0.007272f
C12117 VDD.n6320 GND 0.002244f
C12118 VDD.t1 GND 0.010699f
C12119 VDD.t678 GND 0.010699f
C12120 VDD.n6321 GND 0.022031f
C12121 VDD.n6322 GND 9.03e-19
C12122 VDD.n6323 GND 0.001516f
C12123 VDD.n6324 GND 8.53e-19
C12124 VDD.n6325 GND 0.002454f
C12125 VDD.n6326 GND 0.002363f
C12126 VDD.n6327 GND 8.53e-19
C12127 VDD.n6328 GND 9.03e-19
C12128 VDD.n6329 GND 0.001972f
C12129 VDD.n6330 GND 0.001783f
C12130 VDD.n6331 GND 0.044032f
C12131 VDD.n6332 GND 0.075015f
C12132 VDD.n6333 GND 0.007272f
C12133 VDD.n6334 GND 0.002244f
C12134 VDD.t537 GND 0.010699f
C12135 VDD.t282 GND 0.010699f
C12136 VDD.n6335 GND 0.022031f
C12137 VDD.n6336 GND 9.03e-19
C12138 VDD.n6337 GND 0.001516f
C12139 VDD.n6338 GND 8.53e-19
C12140 VDD.n6339 GND 0.002454f
C12141 VDD.n6340 GND 0.002363f
C12142 VDD.n6341 GND 8.53e-19
C12143 VDD.n6342 GND 9.03e-19
C12144 VDD.n6343 GND 0.001972f
C12145 VDD.n6344 GND 0.001783f
C12146 VDD.n6345 GND 0.044032f
C12147 VDD.n6346 GND 0.056753f
C12148 VDD.n6347 GND 0.007272f
C12149 VDD.n6348 GND 0.007272f
C12150 VDD.n6349 GND 0.007272f
C12151 VDD.n6350 GND 0.007272f
C12152 VDD.n6351 GND 0.002244f
C12153 VDD.t523 GND 0.010699f
C12154 VDD.t62 GND 0.010699f
C12155 VDD.n6352 GND 0.022031f
C12156 VDD.n6353 GND 9.03e-19
C12157 VDD.n6354 GND 0.001516f
C12158 VDD.n6355 GND 8.53e-19
C12159 VDD.n6356 GND 0.002454f
C12160 VDD.n6357 GND 0.002363f
C12161 VDD.n6358 GND 8.53e-19
C12162 VDD.n6359 GND 9.03e-19
C12163 VDD.n6360 GND 0.001972f
C12164 VDD.n6361 GND 0.001783f
C12165 VDD.n6362 GND 0.044032f
C12166 VDD.n6363 GND 0.05786f
C12167 VDD.n6364 GND 0.002244f
C12168 VDD.t536 GND 0.010699f
C12169 VDD.t218 GND 0.010699f
C12170 VDD.n6365 GND 0.022031f
C12171 VDD.n6366 GND 9.03e-19
C12172 VDD.n6367 GND 0.001516f
C12173 VDD.n6368 GND 8.53e-19
C12174 VDD.n6369 GND 0.002454f
C12175 VDD.n6370 GND 0.002363f
C12176 VDD.n6371 GND 8.53e-19
C12177 VDD.n6372 GND 9.03e-19
C12178 VDD.n6373 GND 0.001972f
C12179 VDD.n6374 GND 0.001783f
C12180 VDD.n6375 GND 0.044032f
C12181 VDD.n6376 GND 0.076121f
C12182 VDD.n6377 GND 0.002244f
C12183 VDD.t580 GND 0.010699f
C12184 VDD.t25 GND 0.010699f
C12185 VDD.n6378 GND 0.022031f
C12186 VDD.n6379 GND 9.03e-19
C12187 VDD.n6380 GND 0.001516f
C12188 VDD.n6381 GND 8.53e-19
C12189 VDD.n6382 GND 0.002454f
C12190 VDD.n6383 GND 0.002363f
C12191 VDD.n6384 GND 8.53e-19
C12192 VDD.n6385 GND 9.03e-19
C12193 VDD.n6386 GND 0.001972f
C12194 VDD.n6387 GND 0.001783f
C12195 VDD.n6388 GND 0.044032f
C12196 VDD.n6389 GND 0.075015f
C12197 VDD.n6390 GND 0.002244f
C12198 VDD.t19 GND 0.010699f
C12199 VDD.t142 GND 0.010699f
C12200 VDD.n6391 GND 0.022031f
C12201 VDD.n6392 GND 9.03e-19
C12202 VDD.n6393 GND 0.001516f
C12203 VDD.n6394 GND 8.53e-19
C12204 VDD.n6395 GND 0.002454f
C12205 VDD.n6396 GND 0.002363f
C12206 VDD.n6397 GND 8.53e-19
C12207 VDD.n6398 GND 9.03e-19
C12208 VDD.n6399 GND 0.001972f
C12209 VDD.n6400 GND 0.001783f
C12210 VDD.n6401 GND 0.044032f
C12211 VDD.n6402 GND 0.05786f
C12212 VDD.n6403 GND 0.062709f
C12213 VDD.n6404 GND 0.00991f
C12214 VDD.n6405 GND 0.001706f
C12215 VDD.n6406 GND 0.012142f
C12216 VDD.n6407 GND 0.001706f
C12217 VDD.n6408 GND 0.001706f
C12218 VDD.n6409 GND 0.119161f
C12219 VDD.n6410 GND 0.001706f
C12220 VDD.t176 GND 0.117408f
C12221 VDD.n6411 GND 0.001706f
C12222 VDD.n6412 GND 0.001706f
C12223 VDD.n6413 GND 8.53e-19
C12224 VDD.n6414 GND 9.03e-19
C12225 VDD.n6415 GND 0.010359f
C12226 VDD.n6416 GND 0.010359f
C12227 VDD.n6417 GND 9.03e-19
C12228 VDD.n6418 GND 8.78e-19
C12229 VDD.n6419 GND 0.001706f
C12230 VDD.n6420 GND 0.001706f
C12231 VDD.n6421 GND 0.026285f
C12232 VDD.n6422 GND 0.001706f
C12233 VDD.n6423 GND 0.001706f
C12234 VDD.n6424 GND 8.53e-19
C12235 VDD.n6425 GND 9.03e-19
C12236 VDD.n6426 GND 0.021453f
C12237 VDD.n6427 GND 0.013609f
C12238 VDD.n6428 GND 0.508412f
C12239 VDD.n6429 GND 0.004436f
C12240 VDD.n6430 GND 0.002626f
C12241 VDD.n6431 GND 0.002407f
C12242 VDD.n6432 GND 8.53e-19
C12243 VDD.n6433 GND 0.00291f
C12244 VDD.n6434 GND 9.03e-19
C12245 VDD.n6435 GND 0.041407f
C12246 VDD.n6436 GND 8.53e-19
C12247 VDD.n6437 GND 0.00291f
C12248 VDD.t256 GND 0.00545f
C12249 VDD.n6438 GND 0.007088f
C12250 VDD.n6439 GND 0.001115f
C12251 VDD.n6440 GND 0.002183f
C12252 VDD.n6441 GND 0.00291f
C12253 VDD.n6442 GND 9.03e-19
C12254 VDD.n6443 GND 8.53e-19
C12255 VDD.n6444 GND 0.002385f
C12256 VDD.n6445 GND 0.002421f
C12257 VDD.n6446 GND 8.53e-19
C12258 VDD.n6447 GND 9.03e-19
C12259 VDD.n6448 GND 0.002366f
C12260 VDD.n6449 GND 8.53e-19
C12261 VDD.n6450 GND 9.03e-19
C12262 VDD.n6451 GND 0.00291f
C12263 VDD.n6452 GND 0.005733f
C12264 VDD.n6453 GND 9.03e-19
C12265 VDD.n6454 GND 8.53e-19
C12266 VDD.n6455 GND 0.002417f
C12267 VDD.n6456 GND 0.007268f
C12268 VDD.n6457 GND 0.050371f
C12269 VDD.n6458 GND 0.044305f
C12270 VDD.n6459 GND 0.001512f
C12271 VDD.n6460 GND 0.002407f
C12272 VDD.n6461 GND 8.53e-19
C12273 VDD.t203 GND 0.010699f
C12274 VDD.n6462 GND 0.001399f
C12275 VDD.n6463 GND 0.002366f
C12276 VDD.n6464 GND 0.001972f
C12277 VDD.n6465 GND 9.03e-19
C12278 VDD.t159 GND 0.010699f
C12279 VDD.n6466 GND 0.02202f
C12280 VDD.n6467 GND 9.03e-19
C12281 VDD.n6468 GND 8.53e-19
C12282 VDD.n6469 GND 0.002417f
C12283 VDD.n6470 GND 0.007268f
C12284 VDD.n6471 GND 0.062508f
C12285 VDD.n6472 GND 0.115599f
C12286 VDD.n6473 GND 0.044305f
C12287 VDD.n6474 GND 0.001512f
C12288 VDD.n6475 GND 0.002407f
C12289 VDD.n6476 GND 8.53e-19
C12290 VDD.t9 GND 0.010699f
C12291 VDD.n6477 GND 0.001399f
C12292 VDD.n6478 GND 0.002366f
C12293 VDD.n6479 GND 0.001972f
C12294 VDD.n6480 GND 9.03e-19
C12295 VDD.t558 GND 0.010699f
C12296 VDD.n6481 GND 0.02202f
C12297 VDD.n6482 GND 9.03e-19
C12298 VDD.n6483 GND 8.53e-19
C12299 VDD.n6484 GND 0.002417f
C12300 VDD.n6485 GND 0.007268f
C12301 VDD.n6486 GND 0.063726f
C12302 VDD.n6487 GND 0.044305f
C12303 VDD.n6488 GND 0.001512f
C12304 VDD.n6489 GND 0.002407f
C12305 VDD.n6490 GND 8.53e-19
C12306 VDD.t265 GND 0.010699f
C12307 VDD.n6491 GND 0.001399f
C12308 VDD.n6492 GND 0.002366f
C12309 VDD.n6493 GND 0.001972f
C12310 VDD.n6494 GND 9.03e-19
C12311 VDD.t157 GND 0.010699f
C12312 VDD.n6495 GND 0.02202f
C12313 VDD.n6496 GND 9.03e-19
C12314 VDD.n6497 GND 8.53e-19
C12315 VDD.n6498 GND 0.002417f
C12316 VDD.n6499 GND 0.007268f
C12317 VDD.n6500 GND 0.081987f
C12318 VDD.n6501 GND 0.044305f
C12319 VDD.n6502 GND 0.001512f
C12320 VDD.n6503 GND 0.002407f
C12321 VDD.n6504 GND 8.53e-19
C12322 VDD.t139 GND 0.010699f
C12323 VDD.n6505 GND 0.001399f
C12324 VDD.n6506 GND 0.002366f
C12325 VDD.n6507 GND 0.001972f
C12326 VDD.n6508 GND 9.03e-19
C12327 VDD.t208 GND 0.010699f
C12328 VDD.n6509 GND 0.02202f
C12329 VDD.n6510 GND 9.03e-19
C12330 VDD.n6511 GND 8.53e-19
C12331 VDD.n6512 GND 0.002417f
C12332 VDD.n6513 GND 0.007268f
C12333 VDD.n6514 GND 0.081987f
C12334 VDD.n6515 GND 0.044305f
C12335 VDD.n6516 GND 0.001512f
C12336 VDD.n6517 GND 0.002407f
C12337 VDD.n6518 GND 8.53e-19
C12338 VDD.t374 GND 0.010699f
C12339 VDD.n6519 GND 0.001399f
C12340 VDD.n6520 GND 0.002366f
C12341 VDD.n6521 GND 0.001972f
C12342 VDD.n6522 GND 9.03e-19
C12343 VDD.t376 GND 0.010699f
C12344 VDD.n6523 GND 0.02202f
C12345 VDD.n6524 GND 9.03e-19
C12346 VDD.n6525 GND 8.53e-19
C12347 VDD.n6526 GND 0.002417f
C12348 VDD.n6527 GND 0.007268f
C12349 VDD.n6528 GND 0.081987f
C12350 VDD.n6529 GND 0.044305f
C12351 VDD.n6530 GND 0.001512f
C12352 VDD.n6531 GND 0.002407f
C12353 VDD.n6532 GND 8.53e-19
C12354 VDD.t168 GND 0.010699f
C12355 VDD.n6533 GND 0.001399f
C12356 VDD.n6534 GND 0.002366f
C12357 VDD.n6535 GND 0.001972f
C12358 VDD.n6536 GND 9.03e-19
C12359 VDD.t562 GND 0.010699f
C12360 VDD.n6537 GND 0.02202f
C12361 VDD.n6538 GND 9.03e-19
C12362 VDD.n6539 GND 8.53e-19
C12363 VDD.n6540 GND 0.002417f
C12364 VDD.n6541 GND 0.007268f
C12365 VDD.n6542 GND 0.081987f
C12366 VDD.n6543 GND 0.044305f
C12367 VDD.n6544 GND 0.001512f
C12368 VDD.n6545 GND 0.002407f
C12369 VDD.n6546 GND 8.53e-19
C12370 VDD.t86 GND 0.010699f
C12371 VDD.n6547 GND 0.001399f
C12372 VDD.n6548 GND 0.002366f
C12373 VDD.n6549 GND 0.001972f
C12374 VDD.n6550 GND 9.03e-19
C12375 VDD.t28 GND 0.010699f
C12376 VDD.n6551 GND 0.02202f
C12377 VDD.n6552 GND 9.03e-19
C12378 VDD.n6553 GND 8.53e-19
C12379 VDD.n6554 GND 0.002417f
C12380 VDD.n6555 GND 0.007268f
C12381 VDD.n6556 GND 0.063726f
C12382 VDD.n6557 GND 0.044305f
C12383 VDD.n6558 GND 0.044305f
C12384 VDD.n6559 GND 0.044305f
C12385 VDD.n6560 GND 0.044305f
C12386 VDD.n6561 GND 0.044305f
C12387 VDD.n6562 GND 0.044305f
C12388 VDD.n6563 GND 0.044305f
C12389 VDD.n6564 GND 0.044305f
C12390 VDD.n6565 GND 0.044305f
C12391 VDD.n6566 GND 0.044305f
C12392 VDD.n6567 GND 0.044305f
C12393 VDD.n6568 GND 0.044305f
C12394 VDD.n6569 GND 0.004436f
C12395 VDD.n6570 GND 0.002626f
C12396 VDD.n6571 GND 0.002407f
C12397 VDD.n6572 GND 8.53e-19
C12398 VDD.n6573 GND 0.00291f
C12399 VDD.n6574 GND 9.03e-19
C12400 VDD.n6575 GND 0.041407f
C12401 VDD.n6576 GND 8.53e-19
C12402 VDD.n6577 GND 0.00291f
C12403 VDD.t180 GND 0.00545f
C12404 VDD.n6578 GND 0.007088f
C12405 VDD.n6579 GND 0.001115f
C12406 VDD.n6580 GND 0.002183f
C12407 VDD.n6581 GND 0.00291f
C12408 VDD.n6582 GND 9.03e-19
C12409 VDD.n6583 GND 8.53e-19
C12410 VDD.n6584 GND 0.002385f
C12411 VDD.n6585 GND 0.002421f
C12412 VDD.n6586 GND 8.53e-19
C12413 VDD.n6587 GND 9.03e-19
C12414 VDD.n6588 GND 0.002366f
C12415 VDD.n6589 GND 8.53e-19
C12416 VDD.n6590 GND 9.03e-19
C12417 VDD.n6591 GND 0.00291f
C12418 VDD.n6592 GND 0.005733f
C12419 VDD.n6593 GND 9.03e-19
C12420 VDD.n6594 GND 8.53e-19
C12421 VDD.n6595 GND 0.002417f
C12422 VDD.n6596 GND 0.007268f
C12423 VDD.n6597 GND 0.051588f
C12424 VDD.n6598 GND 0.001512f
C12425 VDD.n6599 GND 0.002407f
C12426 VDD.n6600 GND 8.53e-19
C12427 VDD.t284 GND 0.010699f
C12428 VDD.n6601 GND 0.001399f
C12429 VDD.n6602 GND 0.002366f
C12430 VDD.n6603 GND 0.001972f
C12431 VDD.n6604 GND 9.03e-19
C12432 VDD.t170 GND 0.010699f
C12433 VDD.n6605 GND 0.02202f
C12434 VDD.n6606 GND 9.03e-19
C12435 VDD.n6607 GND 8.53e-19
C12436 VDD.n6608 GND 0.002417f
C12437 VDD.n6609 GND 0.007268f
C12438 VDD.n6610 GND 0.062508f
C12439 VDD.n6611 GND 0.113942f
C12440 VDD.n6612 GND 0.001512f
C12441 VDD.n6613 GND 0.002407f
C12442 VDD.n6614 GND 8.53e-19
C12443 VDD.t131 GND 0.010699f
C12444 VDD.n6615 GND 0.001399f
C12445 VDD.n6616 GND 0.002366f
C12446 VDD.n6617 GND 0.001972f
C12447 VDD.n6618 GND 9.03e-19
C12448 VDD.t510 GND 0.010699f
C12449 VDD.n6619 GND 0.02202f
C12450 VDD.n6620 GND 9.03e-19
C12451 VDD.n6621 GND 8.53e-19
C12452 VDD.n6622 GND 0.002417f
C12453 VDD.n6623 GND 0.007268f
C12454 VDD.n6624 GND 0.063726f
C12455 VDD.n6625 GND 0.001512f
C12456 VDD.n6626 GND 0.002407f
C12457 VDD.n6627 GND 8.53e-19
C12458 VDD.t269 GND 0.010699f
C12459 VDD.n6628 GND 0.001399f
C12460 VDD.n6629 GND 0.002366f
C12461 VDD.n6630 GND 0.001972f
C12462 VDD.n6631 GND 9.03e-19
C12463 VDD.t323 GND 0.010699f
C12464 VDD.n6632 GND 0.02202f
C12465 VDD.n6633 GND 9.03e-19
C12466 VDD.n6634 GND 8.53e-19
C12467 VDD.n6635 GND 0.002417f
C12468 VDD.n6636 GND 0.007268f
C12469 VDD.n6637 GND 0.081987f
C12470 VDD.n6638 GND 0.001512f
C12471 VDD.n6639 GND 0.002407f
C12472 VDD.n6640 GND 8.53e-19
C12473 VDD.t319 GND 0.010699f
C12474 VDD.n6641 GND 0.001399f
C12475 VDD.n6642 GND 0.002366f
C12476 VDD.n6643 GND 0.001972f
C12477 VDD.n6644 GND 9.03e-19
C12478 VDD.t508 GND 0.010699f
C12479 VDD.n6645 GND 0.02202f
C12480 VDD.n6646 GND 9.03e-19
C12481 VDD.n6647 GND 8.53e-19
C12482 VDD.n6648 GND 0.002417f
C12483 VDD.n6649 GND 0.007268f
C12484 VDD.n6650 GND 0.081987f
C12485 VDD.n6651 GND 0.001512f
C12486 VDD.n6652 GND 0.002407f
C12487 VDD.n6653 GND 8.53e-19
C12488 VDD.t215 GND 0.010699f
C12489 VDD.n6654 GND 0.001399f
C12490 VDD.n6655 GND 0.002366f
C12491 VDD.n6656 GND 0.001972f
C12492 VDD.n6657 GND 9.03e-19
C12493 VDD.t342 GND 0.010699f
C12494 VDD.n6658 GND 0.02202f
C12495 VDD.n6659 GND 9.03e-19
C12496 VDD.n6660 GND 8.53e-19
C12497 VDD.n6661 GND 0.002417f
C12498 VDD.n6662 GND 0.007268f
C12499 VDD.n6663 GND 0.083204f
C12500 VDD.n6664 GND 0.001512f
C12501 VDD.n6665 GND 0.002407f
C12502 VDD.n6666 GND 8.53e-19
C12503 VDD.t182 GND 0.010699f
C12504 VDD.n6667 GND 0.001399f
C12505 VDD.n6668 GND 0.002366f
C12506 VDD.n6669 GND 0.001972f
C12507 VDD.n6670 GND 9.03e-19
C12508 VDD.t41 GND 0.010699f
C12509 VDD.n6671 GND 0.02202f
C12510 VDD.n6672 GND 9.03e-19
C12511 VDD.n6673 GND 8.53e-19
C12512 VDD.n6674 GND 0.002417f
C12513 VDD.n6675 GND 0.007268f
C12514 VDD.n6676 GND 0.081987f
C12515 VDD.n6677 GND 0.001512f
C12516 VDD.n6678 GND 0.002407f
C12517 VDD.n6679 GND 8.53e-19
C12518 VDD.t560 GND 0.010699f
C12519 VDD.n6680 GND 0.001399f
C12520 VDD.n6681 GND 0.002366f
C12521 VDD.n6682 GND 0.001972f
C12522 VDD.n6683 GND 9.03e-19
C12523 VDD.t330 GND 0.010699f
C12524 VDD.n6684 GND 0.02202f
C12525 VDD.n6685 GND 9.03e-19
C12526 VDD.n6686 GND 8.53e-19
C12527 VDD.n6687 GND 0.002417f
C12528 VDD.n6688 GND 0.007268f
C12529 VDD.n6689 GND 0.062508f
C12530 VDD.n6690 GND 0.06242f
C12531 VDD.n6691 GND 0.001512f
C12532 VDD.n6692 GND 0.002407f
C12533 VDD.n6693 GND 8.53e-19
C12534 VDD.t129 GND 0.010699f
C12535 VDD.n6694 GND 0.001399f
C12536 VDD.n6695 GND 0.002366f
C12537 VDD.n6696 GND 0.001972f
C12538 VDD.n6697 GND 9.03e-19
C12539 VDD.t371 GND 0.010699f
C12540 VDD.n6698 GND 0.02202f
C12541 VDD.n6699 GND 9.03e-19
C12542 VDD.n6700 GND 8.53e-19
C12543 VDD.n6701 GND 0.002417f
C12544 VDD.n6702 GND 0.007268f
C12545 VDD.n6703 GND 0.063726f
C12546 VDD.n6704 GND 0.001512f
C12547 VDD.n6705 GND 0.002407f
C12548 VDD.n6706 GND 8.53e-19
C12549 VDD.t184 GND 0.010699f
C12550 VDD.n6707 GND 0.001399f
C12551 VDD.n6708 GND 0.002366f
C12552 VDD.n6709 GND 0.001972f
C12553 VDD.n6710 GND 9.03e-19
C12554 VDD.t226 GND 0.010699f
C12555 VDD.n6711 GND 0.02202f
C12556 VDD.n6712 GND 9.03e-19
C12557 VDD.n6713 GND 8.53e-19
C12558 VDD.n6714 GND 0.002417f
C12559 VDD.n6715 GND 0.007268f
C12560 VDD.n6716 GND 0.081987f
C12561 VDD.n6717 GND 0.001512f
C12562 VDD.n6718 GND 0.002407f
C12563 VDD.n6719 GND 8.53e-19
C12564 VDD.t364 GND 0.010699f
C12565 VDD.n6720 GND 0.001399f
C12566 VDD.n6721 GND 0.002366f
C12567 VDD.n6722 GND 0.001972f
C12568 VDD.n6723 GND 9.03e-19
C12569 VDD.t327 GND 0.010699f
C12570 VDD.n6724 GND 0.02202f
C12571 VDD.n6725 GND 9.03e-19
C12572 VDD.n6726 GND 8.53e-19
C12573 VDD.n6727 GND 0.002417f
C12574 VDD.n6728 GND 0.007268f
C12575 VDD.n6729 GND 0.081987f
C12576 VDD.n6730 GND 0.001512f
C12577 VDD.n6731 GND 0.002407f
C12578 VDD.n6732 GND 8.53e-19
C12579 VDD.t704 GND 0.010699f
C12580 VDD.n6733 GND 0.001399f
C12581 VDD.n6734 GND 0.002366f
C12582 VDD.n6735 GND 0.001972f
C12583 VDD.n6736 GND 9.03e-19
C12584 VDD.t317 GND 0.010699f
C12585 VDD.n6737 GND 0.02202f
C12586 VDD.n6738 GND 9.03e-19
C12587 VDD.n6739 GND 8.53e-19
C12588 VDD.n6740 GND 0.002417f
C12589 VDD.n6741 GND 0.007268f
C12590 VDD.n6742 GND 0.081987f
C12591 VDD.n6743 GND 0.001512f
C12592 VDD.n6744 GND 0.002407f
C12593 VDD.n6745 GND 8.53e-19
C12594 VDD.t177 GND 0.010699f
C12595 VDD.n6746 GND 0.001399f
C12596 VDD.n6747 GND 0.002366f
C12597 VDD.n6748 GND 0.001972f
C12598 VDD.n6749 GND 9.03e-19
C12599 VDD.t155 GND 0.010699f
C12600 VDD.n6750 GND 0.02202f
C12601 VDD.n6751 GND 9.03e-19
C12602 VDD.n6752 GND 8.53e-19
C12603 VDD.n6753 GND 0.002417f
C12604 VDD.n6754 GND 0.007268f
C12605 VDD.n6755 GND 0.062508f
C12606 VDD.n6756 GND 0.06242f
C12607 VDD.n6757 GND 0.506755f
C12608 VDD.n6758 GND 0.859285f
C12609 VDD.n6759 GND 0.010271f
C12610 VDD.n6760 GND 0.017055f
C12611 VDD.n6761 GND 9.03e-19
C12612 VDD.n6762 GND 8.78e-19
C12613 VDD.n6763 GND 0.001706f
C12614 VDD.n6764 GND 0.001706f
C12615 VDD.t128 GND 0.117408f
C12616 VDD.n6765 GND 0.001706f
C12617 VDD.n6766 GND 0.001706f
C12618 VDD.n6767 GND 0.001706f
C12619 VDD.t165 GND 0.117408f
C12620 VDD.n6768 GND 0.001706f
C12621 VDD.n6769 GND 0.001706f
C12622 VDD.n6770 GND 0.001706f
C12623 VDD.n6771 GND 8.53e-19
C12624 VDD.n6772 GND 9.03e-19
C12625 VDD.n6773 GND 0.010359f
C12626 VDD.n6774 GND 0.010359f
C12627 VDD.n6775 GND 8.78e-19
C12628 VDD.n6776 GND 8.53e-19
C12629 VDD.n6777 GND 0.001706f
C12630 VDD.n6778 GND 0.001706f
C12631 VDD.t370 GND 0.117408f
C12632 VDD.n6779 GND 0.119161f
C12633 VDD.n6780 GND 0.001706f
C12634 VDD.n6781 GND 8.53e-19
C12635 VDD.n6782 GND 9.03e-19
C12636 VDD.n6783 GND 0.002444f
C12637 VDD.n6784 GND 8.53e-19
C12638 VDD.n6785 GND 0.001706f
C12639 VDD.t216 GND 0.117408f
C12640 VDD.n6786 GND 0.001706f
C12641 VDD.n6787 GND 0.001706f
C12642 VDD.n6788 GND 0.001706f
C12643 VDD.t559 GND 0.117408f
C12644 VDD.n6789 GND 0.001706f
C12645 VDD.n6790 GND 0.001706f
C12646 VDD.n6791 GND 0.001706f
C12647 VDD.n6792 GND 8.53e-19
C12648 VDD.n6793 GND 0.001706f
C12649 VDD.n6794 GND 0.001706f
C12650 VDD.n6795 GND 0.06659f
C12651 VDD.n6796 GND 0.001706f
C12652 VDD.n6797 GND 0.001706f
C12653 VDD.t329 GND 0.117408f
C12654 VDD.n6798 GND 0.001706f
C12655 VDD.n6799 GND 0.001706f
C12656 VDD.n6800 GND 0.012142f
C12657 VDD.n6801 GND 0.00133f
C12658 VDD.n6802 GND 0.001706f
C12659 VDD.n6803 GND 0.001706f
C12660 VDD.n6804 GND 0.049066f
C12661 VDD.n6805 GND 0.001706f
C12662 VDD.n6806 GND 0.001706f
C12663 VDD.n6807 GND 0.110399f
C12664 VDD.n6808 GND 0.001706f
C12665 VDD.n6809 GND 0.001706f
C12666 VDD.n6810 GND 8.53e-19
C12667 VDD.n6811 GND 9.03e-19
C12668 VDD.n6812 GND 0.002444f
C12669 VDD.n6813 GND 9.03e-19
C12670 VDD.n6814 GND 8.53e-19
C12671 VDD.n6815 GND 0.001706f
C12672 VDD.n6816 GND 9.03e-19
C12673 VDD.n6817 GND 9.03e-19
C12674 VDD.n6818 GND 8.53e-19
C12675 VDD.n6819 GND 0.002444f
C12676 VDD.n6820 GND 0.002444f
C12677 VDD.n6821 GND 0.002444f
C12678 VDD.n6822 GND 8.53e-19
C12679 VDD.n6823 GND 0.001706f
C12680 VDD.n6824 GND 0.119161f
C12681 VDD.n6825 GND 0.001706f
C12682 VDD.n6826 GND 0.001706f
C12683 VDD.n6827 GND 0.001706f
C12684 VDD.t22 GND 0.117408f
C12685 VDD.n6828 GND 0.001706f
C12686 VDD.n6829 GND 0.001706f
C12687 VDD.n6830 GND 0.001706f
C12688 VDD.n6831 GND 0.001706f
C12689 VDD.n6832 GND 0.001706f
C12690 VDD.n6833 GND 0.001706f
C12691 VDD.n6834 GND 0.001706f
C12692 VDD.n6835 GND 0.001706f
C12693 VDD.n6836 GND 0.091123f
C12694 VDD.n6837 GND 0.001706f
C12695 VDD.n6838 GND 0.001706f
C12696 VDD.t314 GND 0.117408f
C12697 VDD.n6839 GND 0.001706f
C12698 VDD.n6840 GND 0.001706f
C12699 VDD.n6841 GND 0.001706f
C12700 VDD.n6842 GND 0.001706f
C12701 VDD.n6843 GND 0.001706f
C12702 VDD.n6844 GND 0.001706f
C12703 VDD.n6845 GND 0.001706f
C12704 VDD.n6846 GND 0.001706f
C12705 VDD.n6847 GND 0.001706f
C12706 VDD.n6848 GND 0.001706f
C12707 VDD.n6849 GND 0.052571f
C12708 VDD.n6850 GND 0.001706f
C12709 VDD.n6851 GND 0.001706f
C12710 VDD.t152 GND 0.117408f
C12711 VDD.n6852 GND 0.001706f
C12712 VDD.n6853 GND 0.003727f
C12713 VDD.n6854 GND 0.003727f
C12714 VDD.n6855 GND 0.014019f
C12715 VDD.n6856 GND 0.003723f
C12716 VDD.n6857 GND 0.003723f
C12717 VDD.n6858 GND 0.187503f
C12718 VDD.n6859 GND 0.003727f
C12719 VDD.n6860 GND 0.001706f
C12720 VDD.n6861 GND 0.001706f
C12721 VDD.n6876 GND 0.003727f
C12722 VDD.n6877 GND 0.075352f
C12723 VDD.n6878 GND 0.001706f
C12724 VDD.n6879 GND 0.001706f
C12725 VDD.n6880 GND 0.031543f
C12726 VDD.n6881 GND 0.001706f
C12727 VDD.n6882 GND 0.070094f
C12728 VDD.n6883 GND 0.001706f
C12729 VDD.n6884 GND 0.001706f
C12730 VDD.n6885 GND 0.001706f
C12731 VDD.n6886 GND 0.108646f
C12732 VDD.n6887 GND 0.001706f
C12733 VDD.n6888 GND 0.001706f
C12734 VDD.n6889 GND 0.119161f
C12735 VDD.n6890 GND 0.001706f
C12736 VDD.n6891 GND 0.001706f
C12737 VDD.n6892 GND 0.012142f
C12738 VDD.n6893 GND 0.024533f
C12739 VDD.n6894 GND 0.001706f
C12740 VDD.n6895 GND 0.001706f
C12741 VDD.n6896 GND 0.063085f
C12742 VDD.n6897 GND 0.001706f
C12743 VDD.n6898 GND 0.001706f
C12744 VDD.n6899 GND 9.03e-19
C12745 VDD.n6900 GND 0.001706f
C12746 VDD.n6901 GND 0.001706f
C12747 VDD.n6902 GND 0.101637f
C12748 VDD.n6903 GND 0.001706f
C12749 VDD.n6904 GND 0.001706f
C12750 VDD.t225 GND 0.117408f
C12751 VDD.n6905 GND 0.001706f
C12752 VDD.n6906 GND 0.001706f
C12753 VDD.n6907 GND 8.53e-19
C12754 VDD.n6908 GND 9.03e-19
C12755 VDD.n6909 GND 0.010359f
C12756 VDD.n6910 GND 9.03e-19
C12757 VDD.n6911 GND 8.53e-19
C12758 VDD.n6912 GND 0.010359f
C12759 VDD.n6913 GND 9.03e-19
C12760 VDD.n6914 GND 8.53e-19
C12761 VDD.n6915 GND 0.001706f
C12762 VDD.n6916 GND 8.78e-19
C12763 VDD.n6917 GND 8.53e-19
C12764 VDD.n6918 GND 9.03e-19
C12765 VDD.n6919 GND 0.001706f
C12766 VDD.n6920 GND 0.001706f
C12767 VDD.t24 GND 0.117408f
C12768 VDD.n6921 GND 0.057828f
C12769 VDD.n6922 GND 0.001706f
C12770 VDD.n6923 GND 9.03e-19
C12771 VDD.n6924 GND 0.018487f
C12772 VDD.n6925 GND 8.53e-19
C12773 VDD.n6926 GND 0.001706f
C12774 VDD.n6927 GND 0.119161f
C12775 VDD.n6928 GND 0.001706f
C12776 VDD.n6929 GND 0.001706f
C12777 VDD.n6930 GND 0.001706f
C12778 VDD.n6931 GND 0.001706f
C12779 VDD.n6932 GND 0.001706f
C12780 VDD.n6933 GND 0.021028f
C12781 VDD.n6934 GND 0.001706f
C12782 VDD.t183 GND 0.117408f
C12783 VDD.n6935 GND 0.001706f
C12784 VDD.n6936 GND 0.001706f
C12785 VDD.n6937 GND 0.001706f
C12786 VDD.n6938 GND 8.53e-19
C12787 VDD.n6939 GND 9.03e-19
C12788 VDD.n6940 GND 0.010359f
C12789 VDD.n6941 GND 9.03e-19
C12790 VDD.n6942 GND 8.53e-19
C12791 VDD.n6943 GND 0.010359f
C12792 VDD.n6944 GND 9.03e-19
C12793 VDD.n6945 GND 8.53e-19
C12794 VDD.n6946 GND 9.03e-19
C12795 VDD.n6947 GND 0.010359f
C12796 VDD.n6948 GND 0.010359f
C12797 VDD.n6949 GND 8.53e-19
C12798 VDD.n6950 GND 0.001706f
C12799 VDD.n6951 GND 8.53e-19
C12800 VDD.n6952 GND 9.03e-19
C12801 VDD.t326 GND 0.117408f
C12802 VDD.t141 GND 0.117408f
C12803 VDD.n6953 GND 0.099885f
C12804 VDD.n6954 GND 0.001706f
C12805 VDD.n6955 GND 0.001706f
C12806 VDD.n6956 GND 8.53e-19
C12807 VDD.n6957 GND 9.03e-19
C12808 VDD.n6958 GND 0.018487f
C12809 VDD.n6959 GND 8.53e-19
C12810 VDD.n6960 GND 0.001706f
C12811 VDD.t363 GND 0.117408f
C12812 VDD.n6961 GND 0.001706f
C12813 VDD.n6962 GND 0.001706f
C12814 VDD.n6963 GND 0.001706f
C12815 VDD.t18 GND 0.117408f
C12816 VDD.n6964 GND 0.001706f
C12817 VDD.n6965 GND 0.001706f
C12818 VDD.n6966 GND 0.001706f
C12819 VDD.n6967 GND 8.53e-19
C12820 VDD.n6968 GND 9.03e-19
C12821 VDD.n6969 GND 0.010359f
C12822 VDD.n6970 GND 0.010359f
C12823 VDD.n6971 GND 9.03e-19
C12824 VDD.n6972 GND 0.010359f
C12825 VDD.n6973 GND 8.53e-19
C12826 VDD.n6974 GND 0.001706f
C12827 VDD.n6975 GND 0.119161f
C12828 VDD.n6976 GND 0.001706f
C12829 VDD.n6977 GND 0.001706f
C12830 VDD.t48 GND 0.117408f
C12831 VDD.n6978 GND 0.001706f
C12832 VDD.n6979 GND 0.001706f
C12833 VDD.n6980 GND 0.001706f
C12834 VDD.n6981 GND 0.001706f
C12835 VDD.n6982 GND 0.001706f
C12836 VDD.n6983 GND 0.001706f
C12837 VDD.n6984 GND 0.001706f
C12838 VDD.n6985 GND 0.001706f
C12839 VDD.n6986 GND 0.05958f
C12840 VDD.n6987 GND 0.001706f
C12841 VDD.n6988 GND 0.001706f
C12842 VDD.n6989 GND 0.098132f
C12843 VDD.n6990 GND 0.001706f
C12844 VDD.n6991 GND 0.001706f
C12845 VDD.n6992 GND 0.119161f
C12846 VDD.n6993 GND 0.001706f
C12847 VDD.n6994 GND 0.001706f
C12848 VDD.n6995 GND 0.001706f
C12849 VDD.n6996 GND 0.038552f
C12850 VDD.n6997 GND 0.001706f
C12851 VDD.t230 GND 0.117408f
C12852 VDD.n6998 GND 0.001706f
C12853 VDD.n6999 GND 0.001706f
C12854 VDD.n7000 GND 0.001706f
C12855 VDD.n7001 GND 8.53e-19
C12856 VDD.n7002 GND 9.03e-19
C12857 VDD.n7003 GND 0.010359f
C12858 VDD.n7004 GND 9.03e-19
C12859 VDD.n7005 GND 8.53e-19
C12860 VDD.n7006 GND 0.010359f
C12861 VDD.n7007 GND 9.03e-19
C12862 VDD.n7008 GND 0.010359f
C12863 VDD.n7009 GND 0.010359f
C12864 VDD.n7010 GND 8.53e-19
C12865 VDD.n7011 GND 0.001706f
C12866 VDD.n7012 GND 0.119161f
C12867 VDD.n7013 GND 0.001706f
C12868 VDD.n7014 GND 0.001706f
C12869 VDD.n7015 GND 8.53e-19
C12870 VDD.n7016 GND 9.03e-19
C12871 VDD.n7017 GND 8.53e-19
C12872 VDD.n7018 GND 0.001706f
C12873 VDD.t262 GND 0.117408f
C12874 VDD.n7019 GND 0.001706f
C12875 VDD.n7020 GND 0.001706f
C12876 VDD.t703 GND 0.117408f
C12877 VDD.n7021 GND 0.001706f
C12878 VDD.n7022 GND 0.001706f
C12879 VDD.n7023 GND 0.001003f
C12880 VDD.n7024 GND 0.012142f
C12881 VDD.n7025 GND 0.001706f
C12882 VDD.n7026 GND 0.077104f
C12883 VDD.n7027 GND 0.001706f
C12884 VDD.t0 GND 0.117408f
C12885 VDD.n7028 GND 0.094628f
C12886 VDD.n7029 GND 0.001706f
C12887 VDD.n7030 GND 0.001706f
C12888 VDD.n7031 GND 0.001706f
C12889 VDD.n7032 GND 0.014019f
C12890 VDD.n7033 GND 0.001706f
C12891 VDD.n7034 GND 0.012142f
C12892 VDD.n7035 GND 0.035047f
C12893 VDD.n7036 GND 0.001706f
C12894 VDD.t2 GND 0.117408f
C12895 VDD.n7037 GND 0.001706f
C12896 VDD.n7038 GND 0.001706f
C12897 VDD.n7039 GND 9.03e-19
C12898 VDD.n7040 GND 0.014037f
C12899 VDD.n7041 GND 0.010359f
C12900 VDD.n7042 GND 9.03e-19
C12901 VDD.n7043 GND 8.53e-19
C12902 VDD.n7044 GND 0.001706f
C12903 VDD.n7045 GND 8.53e-19
C12904 VDD.n7046 GND 9.03e-19
C12905 VDD.t144 GND 0.117408f
C12906 VDD.t27 GND 0.117408f
C12907 VDD.n7047 GND 0.085866f
C12908 VDD.n7048 GND 0.001706f
C12909 VDD.n7049 GND 0.001706f
C12910 VDD.n7050 GND 8.53e-19
C12911 VDD.n7051 GND 9.03e-19
C12912 VDD.n7052 GND 0.002444f
C12913 VDD.n7053 GND 8.53e-19
C12914 VDD.n7054 GND 0.001706f
C12915 VDD.t43 GND 0.117408f
C12916 VDD.n7055 GND 0.001706f
C12917 VDD.n7056 GND 0.001706f
C12918 VDD.n7057 GND 0.001706f
C12919 VDD.t85 GND 0.117408f
C12920 VDD.n7058 GND 0.001706f
C12921 VDD.n7059 GND 0.001706f
C12922 VDD.n7060 GND 0.001706f
C12923 VDD.n7061 GND 0.001706f
C12924 VDD.n7062 GND 0.001706f
C12925 VDD.n7063 GND 0.119161f
C12926 VDD.n7064 GND 0.001706f
C12927 VDD.n7065 GND 0.001706f
C12928 VDD.t561 GND 0.117408f
C12929 VDD.n7066 GND 0.001706f
C12930 VDD.n7067 GND 0.001706f
C12931 VDD.n7068 GND 0.001706f
C12932 VDD.n7069 GND 0.001229f
C12933 VDD.n7070 GND 0.001706f
C12934 VDD.n7071 GND 0.012142f
C12935 VDD.n7072 GND 0.001706f
C12936 VDD.n7073 GND 0.073599f
C12937 VDD.n7074 GND 0.001706f
C12938 VDD.n7075 GND 0.001706f
C12939 VDD.n7076 GND 0.112151f
C12940 VDD.n7077 GND 0.001706f
C12941 VDD.n7078 GND 0.001706f
C12942 VDD.n7079 GND 0.010514f
C12943 VDD.n7080 GND 0.001706f
C12944 VDD.n7081 GND 0.001706f
C12945 VDD.n7082 GND 0.001706f
C12946 VDD.n7083 GND 0.049066f
C12947 VDD.n7084 GND 0.001706f
C12948 VDD.t167 GND 0.117408f
C12949 VDD.n7085 GND 0.001706f
C12950 VDD.n7086 GND 0.001706f
C12951 VDD.n7087 GND 0.001706f
C12952 VDD.n7088 GND 0.001706f
C12953 VDD.n7089 GND 0.001706f
C12954 VDD.n7090 GND 0.087618f
C12955 VDD.n7091 GND 0.001706f
C12956 VDD.n7092 GND 0.001706f
C12957 VDD.t375 GND 0.117408f
C12958 VDD.n7093 GND 0.001706f
C12959 VDD.n7094 GND 0.001706f
C12960 VDD.n7095 GND 0.001706f
C12961 VDD.n7096 GND 0.001706f
C12962 VDD.n7097 GND 0.001706f
C12963 VDD.n7098 GND 0.001706f
C12964 VDD.n7099 GND 8.53e-19
C12965 VDD.n7100 GND 9.03e-19
C12966 VDD.n7101 GND 0.005502f
C12967 VDD.n7102 GND 8.53e-19
C12968 VDD.n7103 GND 0.001706f
C12969 VDD.n7104 GND 0.001706f
C12970 VDD.n7105 GND 0.003723f
C12971 VDD.n7106 GND 0.003723f
C12972 VDD.n7107 GND 0.108646f
C12973 VDD.n7108 GND 0.003723f
C12974 VDD.n7109 GND 0.001706f
C12975 VDD.n7110 GND 0.001706f
C12976 VDD.n7111 GND 0.078856f
C12977 VDD.n7112 GND 0.003727f
C12978 VDD.n7120 GND 0.18575f
C12979 VDD.n7129 GND 0.001706f
C12980 VDD.n7130 GND 0.001706f
C12981 VDD.n7131 GND 0.001706f
C12982 VDD.n7132 GND 0.001706f
C12983 VDD.n7133 GND 0.001706f
C12984 VDD.n7134 GND 0.183998f
C12985 VDD.n7135 GND 0.001706f
C12986 VDD.n7136 GND 0.001706f
C12987 VDD.n7137 GND 0.001706f
C12988 VDD.n7138 GND 0.001706f
C12989 VDD.n7139 GND 0.22255f
C12990 VDD.t138 GND 0.119161f
C12991 VDD.n7140 GND 0.001706f
C12992 VDD.n7141 GND 0.001706f
C12993 VDD.n7142 GND 0.001706f
C12994 VDD.n7143 GND 0.238321f
C12995 VDD.n7144 GND 0.001706f
C12996 VDD.n7145 GND 0.001706f
C12997 VDD.n7146 GND 0.001706f
C12998 VDD.t264 GND 0.119161f
C12999 VDD.n7147 GND 0.001706f
C13000 VDD.n7148 GND 0.001706f
C13001 VDD.n7149 GND 0.001706f
C13002 VDD.t557 GND 0.119161f
C13003 VDD.n7150 GND 0.001706f
C13004 VDD.n7151 GND 0.001706f
C13005 VDD.n7152 GND 0.001706f
C13006 VDD.t8 GND 0.119161f
C13007 VDD.n7153 GND 0.176989f
C13008 VDD.n7154 GND 0.001706f
C13009 VDD.n7155 GND 0.001706f
C13010 VDD.n7156 GND 0.001706f
C13011 VDD.n7157 GND 0.138437f
C13012 VDD.n7158 GND 0.001706f
C13013 VDD.n7159 GND 0.001706f
C13014 VDD.n7160 GND 0.001706f
C13015 VDD.n7161 GND 0.176989f
C13016 VDD.t158 GND 0.119161f
C13017 VDD.n7162 GND 0.001706f
C13018 VDD.n7163 GND 0.001706f
C13019 VDD.n7164 GND 0.001706f
C13020 VDD.n7165 GND 0.215541f
C13021 VDD.n7166 GND 0.001706f
C13022 VDD.n7167 GND 0.003781f
C13023 VDD.n7168 GND 0.003781f
C13024 VDD.n7169 GND 0.315425f
C13025 VDD.t255 GND 0.119161f
C13026 VDD.n7170 GND 0.003781f
C13027 VDD.n7171 GND 0.001706f
C13028 VDD.n7172 GND 0.001706f
C13029 VDD.n7180 GND 0.001706f
C13030 VDD.n7181 GND 0.001706f
C13031 VDD.n7182 GND 0.001706f
C13032 VDD.n7183 GND 0.001706f
C13033 VDD.n7184 GND 0.001706f
C13034 VDD.n7185 GND 0.001706f
C13035 VDD.n7186 GND 0.001706f
C13036 VDD.n7187 GND 0.001706f
C13037 VDD.n7188 GND 0.001706f
C13038 VDD.n7189 GND 0.001706f
C13039 VDD.n7190 GND 0.001706f
C13040 VDD.n7191 GND 0.001706f
C13041 VDD.n7192 GND 0.001706f
C13042 VDD.n7193 GND 0.001706f
C13043 VDD.n7194 GND 0.001706f
C13044 VDD.n7195 GND 0.001706f
C13045 VDD.n7196 GND 0.001706f
C13046 VDD.n7197 GND 0.001706f
C13047 VDD.n7198 GND 0.001706f
C13048 VDD.n7199 GND 0.001706f
C13049 VDD.n7200 GND 0.001706f
C13050 VDD.n7201 GND 0.001706f
C13051 VDD.n7202 GND 0.001706f
C13052 VDD.n7203 GND 0.001706f
C13053 VDD.n7204 GND 0.001706f
C13054 VDD.n7205 GND 0.001706f
C13055 VDD.n7206 GND 0.001706f
C13056 VDD.n7207 GND 0.001706f
C13057 VDD.n7208 GND 0.003795f
C13058 VDD.n7209 GND 0.003795f
C13059 VDD.n7210 GND 0.403043f
C13060 VDD.n7212 GND 0.003795f
C13061 VDD.n7213 GND 0.003795f
C13062 VDD.n7214 GND 0.003781f
C13063 VDD.n7215 GND 0.001706f
C13064 VDD.n7216 GND 0.001706f
C13065 VDD.n7217 GND 0.141941f
C13066 VDD.n7218 GND 0.001706f
C13067 VDD.n7219 GND 0.001706f
C13068 VDD.n7220 GND 0.001706f
C13069 VDD.n7221 GND 0.001706f
C13070 VDD.n7222 GND 0.001706f
C13071 VDD.t202 GND 0.119161f
C13072 VDD.n7223 GND 0.180493f
C13073 VDD.n7224 GND 0.001706f
C13074 VDD.n7225 GND 0.001706f
C13075 VDD.n7226 GND 0.001706f
C13076 VDD.n7227 GND 0.001706f
C13077 VDD.n7228 GND 0.001706f
C13078 VDD.n7229 GND 0.219045f
C13079 VDD.n7230 GND 0.001706f
C13080 VDD.n7231 GND 0.001706f
C13081 VDD.n7232 GND 0.001706f
C13082 VDD.n7233 GND 0.001706f
C13083 VDD.n7234 GND 0.001706f
C13084 VDD.n7235 GND 0.138437f
C13085 VDD.n7236 GND 0.238321f
C13086 VDD.n7237 GND 0.001706f
C13087 VDD.n7238 GND 0.001706f
C13088 VDD.n7239 GND 0.001706f
C13089 VDD.n7240 GND 0.001706f
C13090 VDD.n7241 GND 0.001706f
C13091 VDD.n7242 GND 0.219045f
C13092 VDD.n7243 GND 0.001706f
C13093 VDD.n7244 GND 0.001706f
C13094 VDD.n7245 GND 0.001706f
C13095 VDD.n7246 GND 0.001706f
C13096 VDD.n7247 GND 0.001706f
C13097 VDD.n7248 GND 0.215541f
C13098 VDD.n7249 GND 0.180493f
C13099 VDD.n7250 GND 0.001706f
C13100 VDD.n7251 GND 0.001706f
C13101 VDD.n7252 GND 0.001706f
C13102 VDD.n7253 GND 0.001706f
C13103 VDD.n7254 GND 0.001706f
C13104 VDD.n7255 GND 0.141941f
C13105 VDD.n7256 GND 0.001706f
C13106 VDD.n7257 GND 0.001706f
C13107 VDD.n7258 GND 0.001706f
C13108 VDD.n7259 GND 0.001706f
C13109 VDD.n7260 GND 0.001706f
C13110 VDD.t156 GND 0.119161f
C13111 VDD.n7261 GND 0.134932f
C13112 VDD.n7262 GND 0.001706f
C13113 VDD.n7263 GND 0.001706f
C13114 VDD.n7264 GND 0.001706f
C13115 VDD.n7265 GND 0.001706f
C13116 VDD.n7266 GND 0.001706f
C13117 VDD.n7267 GND 0.001706f
C13118 VDD.n7268 GND 0.173484f
C13119 VDD.n7269 GND 0.001706f
C13120 VDD.n7270 GND 0.001706f
C13121 VDD.n7271 GND 0.001706f
C13122 VDD.n7272 GND 9.17e-19
C13123 VDD.n7273 GND 9.03e-19
C13124 VDD.n7274 GND 0.002444f
C13125 VDD.n7275 GND 9.03e-19
C13126 VDD.n7276 GND 0.002444f
C13127 VDD.n7277 GND 8.53e-19
C13128 VDD.n7278 GND 0.001706f
C13129 VDD.n7279 GND 9.03e-19
C13130 VDD.n7280 GND 0.002313f
C13131 VDD.n7281 GND 8.53e-19
C13132 VDD.n7282 GND 9.03e-19
C13133 VDD.n7283 GND 8.53e-19
C13134 VDD.n7284 GND 0.002444f
C13135 VDD.n7285 GND 0.002444f
C13136 VDD.n7286 GND 8.53e-19
C13137 VDD.n7287 GND 9.03e-19
C13138 VDD.n7288 GND 0.001706f
C13139 VDD.n7289 GND 0.001706f
C13140 VDD.n7290 GND 9.03e-19
C13141 VDD.n7291 GND 8.53e-19
C13142 VDD.n7292 GND 0.002444f
C13143 VDD.n7293 GND 0.002444f
C13144 VDD.n7294 GND 8.53e-19
C13145 VDD.n7295 GND 9.03e-19
C13146 VDD.n7296 GND 8.53e-19
C13147 VDD.n7297 GND 0.001706f
C13148 VDD.n7298 GND 9.03e-19
C13149 VDD.n7299 GND 8.53e-19
C13150 VDD.n7300 GND 0.002444f
C13151 VDD.n7301 GND 0.005502f
C13152 VDD.n7302 GND 8.53e-19
C13153 VDD.n7303 GND 9.03e-19
C13154 VDD.n7304 GND 0.001706f
C13155 VDD.n7305 GND 0.001706f
C13156 VDD.n7306 GND 0.001029f
C13157 VDD.n7307 GND 0.001706f
C13158 VDD.n7308 GND 0.001706f
C13159 VDD.n7309 GND 0.001706f
C13160 VDD.n7310 GND 0.001706f
C13161 VDD.n7311 GND 0.001706f
C13162 VDD.n7312 GND 0.001706f
C13163 VDD.t207 GND 0.119161f
C13164 VDD.n7313 GND 0.212036f
C13165 VDD.n7314 GND 0.001706f
C13166 VDD.n7315 GND 0.001706f
C13167 VDD.n7316 GND 0.001706f
C13168 VDD.n7317 GND 0.001706f
C13169 VDD.n7318 GND 9.03e-19
C13170 VDD.n7319 GND 9.17e-19
C13171 VDD.n7320 GND 0.001029f
C13172 VDD.n7321 GND 0.001706f
C13173 VDD.n7322 GND 0.001706f
C13174 VDD.n7323 GND 0.120913f
C13175 VDD.t373 GND 0.117408f
C13176 VDD.n7324 GND 0.001706f
C13177 VDD.n7325 GND 0.001706f
C13178 VDD.n7326 GND 0.001706f
C13179 VDD.n7327 GND 0.001706f
C13180 VDD.n7328 GND 0.001706f
C13181 VDD.n7329 GND 0.001706f
C13182 VDD.n7330 GND 0.001706f
C13183 VDD.n7331 GND 0.001706f
C13184 VDD.n7332 GND 0.001706f
C13185 VDD.n7333 GND 0.001706f
C13186 VDD.n7334 GND 0.001706f
C13187 VDD.n7335 GND 0.001706f
C13188 VDD.n7336 GND 0.001706f
C13189 VDD.n7337 GND 0.001706f
C13190 VDD.n7338 GND 0.001706f
C13191 VDD.n7339 GND 0.001706f
C13192 VDD.n7340 GND 0.001706f
C13193 VDD.n7341 GND 0.001706f
C13194 VDD.n7342 GND 0.001706f
C13195 VDD.n7343 GND 0.001706f
C13196 VDD.n7344 GND 0.001706f
C13197 VDD.n7345 GND 0.001706f
C13198 VDD.n7346 GND 0.001706f
C13199 VDD.n7347 GND 0.001706f
C13200 VDD.n7348 GND 0.001706f
C13201 VDD.n7349 GND 0.001706f
C13202 VDD.n7350 GND 0.001706f
C13203 VDD.n7351 GND 0.001706f
C13204 VDD.n7352 GND 0.003727f
C13205 VDD.n7353 GND 0.003723f
C13206 VDD.n7354 GND 0.003723f
C13207 VDD.n7355 GND 0.012266f
C13208 VDD.n7356 GND 0.003723f
C13209 VDD.n7357 GND 0.001706f
C13210 VDD.n7358 GND 0.003723f
C13211 VDD.n7359 GND 0.003727f
C13212 VDD.n7360 GND 0.003727f
C13213 VDD.n7361 GND 0.001706f
C13214 VDD.n7362 GND 0.001706f
C13215 VDD.n7363 GND 0.001706f
C13216 VDD.n7364 GND 0.001706f
C13217 VDD.n7365 GND 0.001706f
C13218 VDD.n7366 GND 0.001706f
C13219 VDD.n7367 GND 0.001706f
C13220 VDD.n7368 GND 0.001706f
C13221 VDD.n7369 GND 0.001706f
C13222 VDD.n7370 GND 0.001706f
C13223 VDD.n7371 GND 0.001706f
C13224 VDD.n7372 GND 0.001706f
C13225 VDD.n7373 GND 0.001706f
C13226 VDD.n7374 GND 0.001706f
C13227 VDD.n7375 GND 0.001706f
C13228 VDD.n7376 GND 0.001706f
C13229 VDD.n7377 GND 0.001706f
C13230 VDD.n7378 GND 0.001706f
C13231 VDD.n7379 GND 0.001706f
C13232 VDD.n7380 GND 0.001706f
C13233 VDD.n7381 GND 0.001706f
C13234 VDD.n7382 GND 0.001706f
C13235 VDD.n7383 GND 0.001706f
C13236 VDD.n7384 GND 0.001706f
C13237 VDD.n7385 GND 0.001706f
C13238 VDD.n7386 GND 0.001706f
C13239 VDD.n7387 GND 0.001706f
C13240 VDD.n7388 GND 0.001706f
C13241 VDD.n7389 GND 0.001706f
C13242 VDD.n7390 GND 0.003727f
C13243 VDD.n7391 GND 0.003727f
C13244 VDD.n7392 GND 0.119161f
C13245 VDD.n7394 GND 0.003727f
C13246 VDD.n7395 GND 0.003727f
C13247 VDD.n7396 GND 0.003723f
C13248 VDD.n7397 GND 0.001706f
C13249 VDD.n7398 GND 0.001706f
C13250 VDD.n7399 GND 0.001706f
C13251 VDD.t297 GND 0.117408f
C13252 VDD.n7400 GND 0.033295f
C13253 VDD.n7401 GND 0.001706f
C13254 VDD.n7402 GND 0.001706f
C13255 VDD.n7403 GND 0.001706f
C13256 VDD.n7404 GND 0.001706f
C13257 VDD.n7405 GND 0.001706f
C13258 VDD.n7406 GND 0.001706f
C13259 VDD.t20 GND 0.117408f
C13260 VDD.n7407 GND 0.071847f
C13261 VDD.n7408 GND 0.070094f
C13262 VDD.n7409 GND 0.001706f
C13263 VDD.n7410 GND 9.03e-19
C13264 VDD.n7411 GND 9.03e-19
C13265 VDD.n7412 GND 8.53e-19
C13266 VDD.n7413 GND 0.002444f
C13267 VDD.n7414 GND 0.002444f
C13268 VDD.n7415 GND 0.002444f
C13269 VDD.n7416 GND 9.03e-19
C13270 VDD.n7417 GND 8.53e-19
C13271 VDD.n7418 GND 0.001706f
C13272 VDD.n7419 GND 9.03e-19
C13273 VDD.n7420 GND 8.53e-19
C13274 VDD.n7421 GND 0.002444f
C13275 VDD.n7422 GND 0.002444f
C13276 VDD.n7423 GND 8.53e-19
C13277 VDD.n7424 GND 9.03e-19
C13278 VDD.n7425 GND 0.001706f
C13279 VDD.n7426 GND 0.031543f
C13280 VDD.t38 GND 0.117408f
C13281 VDD.n7427 GND 0.110399f
C13282 VDD.n7428 GND 0.001706f
C13283 VDD.n7429 GND 0.001706f
C13284 VDD.n7430 GND 0.001706f
C13285 VDD.n7431 GND 0.001706f
C13286 VDD.n7432 GND 0.001706f
C13287 VDD.n7433 GND 0.001706f
C13288 VDD.n7434 GND 0.050818f
C13289 VDD.n7435 GND 0.001706f
C13290 VDD.n7436 GND 0.001706f
C13291 VDD.n7437 GND 0.001706f
C13292 VDD.n7438 GND 0.001706f
C13293 VDD.n7439 GND 0.001706f
C13294 VDD.n7440 GND 0.001706f
C13295 VDD.n7441 GND 0.08937f
C13296 VDD.n7442 GND 0.001706f
C13297 VDD.n7443 GND 0.001706f
C13298 VDD.n7444 GND 0.001706f
C13299 VDD.n7445 GND 0.001706f
C13300 VDD.n7446 GND 0.001706f
C13301 VDD.n7447 GND 0.119161f
C13302 VDD.n7448 GND 0.001706f
C13303 VDD.n7449 GND 0.001706f
C13304 VDD.n7450 GND 0.001706f
C13305 VDD.n7451 GND 0.001706f
C13306 VDD.n7452 GND 0.001706f
C13307 VDD.n7453 GND 0.02979f
C13308 VDD.n7454 GND 0.001706f
C13309 VDD.n7455 GND 0.001706f
C13310 VDD.n7456 GND 0.001706f
C13311 VDD.n7457 GND 0.001706f
C13312 VDD.n7458 GND 0.001706f
C13313 VDD.n7459 GND 0.001706f
C13314 VDD.n7460 GND 0.068342f
C13315 VDD.n7461 GND 0.001706f
C13316 VDD.n7462 GND 0.009463f
C13317 VDD.n7463 GND 0.004145f
C13318 VDD.n7464 GND 0.001229f
C13319 VDD.n7465 GND 0.001706f
C13320 VDD.n7466 GND 0.001706f
C13321 VDD.n7467 GND 0.001706f
C13322 VDD.n7468 GND 0.008762f
C13323 VDD.n7469 GND 0.001706f
C13324 VDD.n7470 GND 0.001706f
C13325 VDD.n7471 GND 0.001706f
C13326 VDD.n7472 GND 0.001706f
C13327 VDD.n7473 GND 0.001706f
C13328 VDD.n7474 GND 0.001706f
C13329 VDD.n7475 GND 0.047314f
C13330 VDD.n7476 GND 0.091123f
C13331 VDD.n7477 GND 0.001706f
C13332 VDD.n7478 GND 9.03e-19
C13333 VDD.n7479 GND 9.03e-19
C13334 VDD.n7480 GND 8.53e-19
C13335 VDD.n7481 GND 0.002444f
C13336 VDD.n7482 GND 0.002444f
C13337 VDD.n7483 GND 0.003712f
C13338 VDD.n7484 GND 9.03e-19
C13339 VDD.n7485 GND 8.53e-19
C13340 VDD.n7486 GND 0.001706f
C13341 VDD.n7487 GND 9.03e-19
C13342 VDD.n7488 GND 8.53e-19
C13343 VDD.n7489 GND 0.002444f
C13344 VDD.n7490 GND 0.002444f
C13345 VDD.n7491 GND 8.53e-19
C13346 VDD.n7492 GND 9.03e-19
C13347 VDD.n7493 GND 0.001706f
C13348 VDD.n7494 GND 0.052571f
C13349 VDD.n7495 GND 0.001706f
C13350 VDD.n7496 GND 0.001706f
C13351 VDD.n7497 GND 0.001706f
C13352 VDD.n7498 GND 9.03e-19
C13353 VDD.n7499 GND 8.53e-19
C13354 VDD.n7500 GND 0.010359f
C13355 VDD.n7501 GND 0.010359f
C13356 VDD.n7502 GND 8.53e-19
C13357 VDD.n7503 GND 0.001129f
C13358 VDD.n7504 GND 0.001706f
C13359 VDD.n7505 GND 0.106894f
C13360 VDD.n7506 GND 0.001706f
C13361 VDD.n7507 GND 0.001706f
C13362 VDD.n7508 GND 0.119161f
C13363 VDD.n7509 GND 0.001706f
C13364 VDD.n7510 GND 0.001706f
C13365 VDD.n7511 GND 0.001706f
C13366 VDD.n7512 GND 0.001706f
C13367 VDD.n7513 GND 0.001706f
C13368 VDD.n7514 GND 0.001706f
C13369 VDD.n7515 GND 0.001706f
C13370 VDD.t154 GND 0.117408f
C13371 VDD.n7516 GND 0.001706f
C13372 VDD.n7517 GND 0.001706f
C13373 VDD.n7518 GND 0.043809f
C13374 VDD.n7519 GND 0.001706f
C13375 VDD.n7520 GND 8.53e-19
C13376 VDD.n7521 GND 9.03e-19
C13377 VDD.n7522 GND 8.53e-19
C13378 VDD.n7523 GND 9.03e-19
C13379 VDD.n7524 GND 0.010215f
C13380 VDD.n7525 GND 0.010359f
C13381 VDD.n7526 GND 0.006187f
C13382 VDD.n7527 GND 0.009208f
C13383 VDD.n7528 GND 0.098305f
C13384 VDD.n7529 GND 1.00116f
C13385 VDD.n7530 GND 0.098017f
C13386 VDD.n7531 GND 0.005467f
C13387 VDD.n7532 GND 0.010359f
C13388 VDD.n7533 GND 8.53e-19
C13389 VDD.n7534 GND 0.001706f
C13390 VDD.n7535 GND 9.03e-19
C13391 VDD.n7536 GND 8.53e-19
C13392 VDD.n7537 GND 9.03e-19
C13393 VDD.n7538 GND 8.53e-19
C13394 VDD.n7539 GND 9.03e-19
C13395 VDD.n7540 GND 8.53e-19
C13396 VDD.n7541 GND 0.010359f
C13397 VDD.n7542 GND 0.010359f
C13398 VDD.n7543 GND 8.53e-19
C13399 VDD.n7544 GND 9.03e-19
C13400 VDD.n7545 GND 0.001706f
C13401 VDD.n7546 GND 0.064837f
C13402 VDD.n7547 GND 0.001706f
C13403 VDD.n7548 GND 0.011071f
C13404 VDD.n7549 GND 0.005301f
C13405 VDD.n7550 GND 0.001706f
C13406 VDD.n7551 GND 0.001706f
C13407 VDD.n7552 GND 0.001706f
C13408 VDD.n7553 GND 0.001003f
C13409 VDD.n7554 GND 0.001706f
C13410 VDD.n7555 GND 0.082361f
C13411 VDD.n7556 GND 0.056076f
C13412 VDD.n7557 GND 0.001706f
C13413 VDD.n7558 GND 9.03e-19
C13414 VDD.n7559 GND 9.03e-19
C13415 VDD.n7560 GND 8.53e-19
C13416 VDD.n7561 GND 0.018487f
C13417 VDD.n7562 GND 0.018487f
C13418 VDD.n7563 GND 0.018487f
C13419 VDD.n7564 GND 9.03e-19
C13420 VDD.n7565 GND 8.53e-19
C13421 VDD.n7566 GND 0.001706f
C13422 VDD.n7567 GND 9.03e-19
C13423 VDD.n7568 GND 8.53e-19
C13424 VDD.n7569 GND 0.018487f
C13425 VDD.n7570 GND 0.018487f
C13426 VDD.n7571 GND 8.53e-19
C13427 VDD.n7572 GND 9.03e-19
C13428 VDD.n7573 GND 0.001706f
C13429 VDD.n7574 GND 0.017524f
C13430 VDD.n7575 GND 0.001706f
C13431 VDD.n7576 GND 0.001706f
C13432 VDD.n7577 GND 8.53e-19
C13433 VDD.n7578 GND 9.03e-19
C13434 VDD.n7579 GND 0.001706f
C13435 VDD.n7580 GND 0.001706f
C13436 VDD.n7581 GND 9.03e-19
C13437 VDD.n7582 GND 8.53e-19
C13438 VDD.n7583 GND 0.010359f
C13439 VDD.n7584 GND 0.010359f
C13440 VDD.n7585 GND 8.53e-19
C13441 VDD.n7586 GND 9.03e-19
C13442 VDD.n7587 GND 0.001706f
C13443 VDD.n7588 GND 0.103389f
C13444 VDD.n7589 GND 0.001706f
C13445 VDD.n7590 GND 0.001706f
C13446 VDD.n7591 GND 0.001706f
C13447 VDD.n7592 GND 0.001706f
C13448 VDD.n7593 GND 0.001706f
C13449 VDD.t316 GND 0.119161f
C13450 VDD.n7594 GND 0.001706f
C13451 VDD.n7595 GND 0.001706f
C13452 VDD.n7596 GND 0.001706f
C13453 VDD.n7597 GND 0.001706f
C13454 VDD.n7598 GND 0.001706f
C13455 VDD.n7599 GND 0.001706f
C13456 VDD.n7600 GND 0.001706f
C13457 VDD.n7601 GND 0.001706f
C13458 VDD.n7602 GND 0.001706f
C13459 VDD.n7603 GND 0.001706f
C13460 VDD.n7604 GND 0.001706f
C13461 VDD.n7605 GND 0.001706f
C13462 VDD.n7606 GND 0.001706f
C13463 VDD.n7607 GND 0.001706f
C13464 VDD.n7608 GND 0.040304f
C13465 VDD.n7609 GND 0.001706f
C13466 VDD.n7610 GND 0.001706f
C13467 VDD.n7611 GND 0.001706f
C13468 VDD.n7612 GND 0.001706f
C13469 VDD.n7613 GND 0.001706f
C13470 VDD.n7614 GND 0.078856f
C13471 VDD.n7615 GND 0.001706f
C13472 VDD.n7616 GND 0.001706f
C13473 VDD.n7617 GND 0.001706f
C13474 VDD.n7618 GND 0.001706f
C13475 VDD.n7619 GND 0.001706f
C13476 VDD.n7620 GND 0.001706f
C13477 VDD.n7621 GND 0.022781f
C13478 VDD.n7622 GND 0.001706f
C13479 VDD.n7623 GND 9.03e-19
C13480 VDD.n7624 GND 9.03e-19
C13481 VDD.n7625 GND 8.53e-19
C13482 VDD.n7626 GND 0.010359f
C13483 VDD.n7627 GND 0.010359f
C13484 VDD.n7628 GND 0.010359f
C13485 VDD.n7629 GND 8.53e-19
C13486 VDD.n7630 GND 9.03e-19
C13487 VDD.n7631 GND 8.53e-19
C13488 VDD.n7632 GND 9.03e-19
C13489 VDD.n7633 GND 8.53e-19
C13490 VDD.n7634 GND 0.010359f
C13491 VDD.n7635 GND 0.010359f
C13492 VDD.n7636 GND 8.53e-19
C13493 VDD.n7637 GND 8.78e-19
C13494 VDD.n7638 GND 8.78e-19
C13495 VDD.n7639 GND 0.001706f
C13496 VDD.n7640 GND 0.061333f
C13497 VDD.n7641 GND 0.080609f
C13498 VDD.n7642 GND 0.001706f
C13499 VDD.n7643 GND 9.03e-19
C13500 VDD.n7644 GND 9.03e-19
C13501 VDD.n7645 GND 8.53e-19
C13502 VDD.n7646 GND 0.018487f
C13503 VDD.n7647 GND 0.018487f
C13504 VDD.n7648 GND 9.03e-19
C13505 VDD.n7649 GND 8.53e-19
C13506 VDD.n7650 GND 0.018487f
C13507 VDD.n7651 GND 0.018487f
C13508 VDD.n7652 GND 8.53e-19
C13509 VDD.n7653 GND 9.03e-19
C13510 VDD.n7654 GND 0.001706f
C13511 VDD.n7655 GND 0.042057f
C13512 VDD.n7656 GND 0.001706f
C13513 VDD.n7657 GND 0.001706f
C13514 VDD.n7658 GND 0.003505f
C13515 VDD.n7659 GND 0.001706f
C13516 VDD.n7660 GND 9.03e-19
C13517 VDD.n7661 GND 8.53e-19
C13518 VDD.n7662 GND 0.010359f
C13519 VDD.n7663 GND 0.010359f
C13520 VDD.n7664 GND 8.53e-19
C13521 VDD.n7665 GND 9.03e-19
C13522 VDD.n7666 GND 0.001706f
C13523 VDD.n7667 GND 0.117408f
C13524 VDD.n7668 GND 0.001706f
C13525 VDD.n7669 GND 0.001706f
C13526 VDD.n7670 GND 0.001706f
C13527 VDD.n7671 GND 0.001706f
C13528 VDD.n7672 GND 0.001706f
C13529 VDD.n7673 GND 0.001706f
C13530 VDD.t579 GND 0.117408f
C13531 VDD.n7674 GND 0.019276f
C13532 VDD.n7675 GND 0.119161f
C13533 VDD.n7676 GND 0.001706f
C13534 VDD.n7677 GND 9.03e-19
C13535 VDD.n7678 GND 8.53e-19
C13536 VDD.n7679 GND 0.018487f
C13537 VDD.n7680 GND 0.018487f
C13538 VDD.n7681 GND 8.53e-19
C13539 VDD.n7682 GND 8.53e-19
C13540 VDD.n7683 GND 9.03e-19
C13541 VDD.n7684 GND 0.001706f
C13542 VDD.n7685 GND 0.084113f
C13543 VDD.n7686 GND 0.001706f
C13544 VDD.n7687 GND 9.03e-19
C13545 VDD.n7688 GND 8.53e-19
C13546 VDD.n7689 GND 0.010359f
C13547 VDD.n7690 GND 0.010359f
C13548 VDD.n7691 GND 8.53e-19
C13549 VDD.n7692 GND 9.03e-19
C13550 VDD.n7693 GND 0.001706f
C13551 VDD.n7694 GND 0.0368f
C13552 VDD.n7695 GND 0.001706f
C13553 VDD.n7696 GND 0.001706f
C13554 VDD.n7697 GND 9.03e-19
C13555 VDD.n7698 GND 0.005814f
C13556 VDD.n7699 GND 0.012142f
C13557 VDD.n7700 GND 0.011785f
C13558 VDD.n7701 GND 0.001706f
C13559 VDD.n7702 GND 0.075352f
C13560 VDD.n7703 GND 0.001706f
C13561 VDD.n7704 GND 0.001706f
C13562 VDD.n7705 GND 0.001706f
C13563 VDD.n7706 GND 0.001706f
C13564 VDD.n7707 GND 0.001706f
C13565 VDD.n7708 GND 0.113904f
C13566 VDD.n7709 GND 0.001706f
C13567 VDD.n7710 GND 0.001706f
C13568 VDD.n7711 GND 0.007589f
C13569 VDD.n7712 GND 0.001706f
C13570 VDD.n7713 GND 0.012142f
C13571 VDD.n7714 GND 0.010624f
C13572 VDD.n7715 GND 0.001706f
C13573 VDD.n7716 GND 0.015771f
C13574 VDD.n7717 GND 0.001706f
C13575 VDD.n7718 GND 0.001706f
C13576 VDD.n7719 GND 0.001706f
C13577 VDD.n7720 GND 0.001706f
C13578 VDD.n7721 GND 8.53e-19
C13579 VDD.n7722 GND 9.03e-19
C13580 VDD.n7723 GND 0.010359f
C13581 VDD.n7724 GND 8.53e-19
C13582 VDD.n7725 GND 0.001706f
C13583 VDD.n7726 GND 9.03e-19
C13584 VDD.n7727 GND 9.03e-19
C13585 VDD.n7728 GND 8.53e-19
C13586 VDD.n7729 GND 0.010359f
C13587 VDD.n7730 GND 9.03e-19
C13588 VDD.n7731 GND 9.03e-19
C13589 VDD.n7732 GND 8.53e-19
C13590 VDD.n7733 GND 0.010359f
C13591 VDD.n7734 GND 0.010359f
C13592 VDD.n7735 GND 0.014703f
C13593 VDD.n7736 GND 0.002444f
C13594 VDD.t181 GND 0.117408f
C13595 VDD.n7737 GND 0.010514f
C13596 VDD.n7738 GND 0.001706f
C13597 VDD.n7739 GND 9.03e-19
C13598 VDD.n7740 GND 0.002444f
C13599 VDD.n7741 GND 8.53e-19
C13600 VDD.n7742 GND 0.001706f
C13601 VDD.n7743 GND 9.03e-19
C13602 VDD.n7744 GND 0.002444f
C13603 VDD.n7745 GND 9.17e-19
C13604 VDD.n7746 GND 0.001706f
C13605 VDD.n7747 GND 0.001706f
C13606 VDD.n7748 GND 0.001706f
C13607 VDD.n7749 GND 0.001706f
C13608 VDD.t318 GND 0.119161f
C13609 VDD.n7750 GND 0.183998f
C13610 VDD.n7751 GND 0.001706f
C13611 VDD.n7752 GND 0.001706f
C13612 VDD.n7753 GND 0.001706f
C13613 VDD.n7754 GND 0.001706f
C13614 VDD.n7755 GND 9.03e-19
C13615 VDD.n7756 GND 0.002444f
C13616 VDD.n7757 GND 8.53e-19
C13617 VDD.n7758 GND 9.03e-19
C13618 VDD.n7759 GND 0.002444f
C13619 VDD.n7760 GND 8.53e-19
C13620 VDD.n7761 GND 9.03e-19
C13621 VDD.n7762 GND 0.001706f
C13622 VDD.n7763 GND 0.001706f
C13623 VDD.n7764 GND 9.03e-19
C13624 VDD.n7765 GND 8.53e-19
C13625 VDD.n7766 GND 0.005502f
C13626 VDD.n7767 GND 9.17e-19
C13627 VDD.n7768 GND 0.001029f
C13628 VDD.n7769 GND 0.001706f
C13629 VDD.n7770 GND 0.001706f
C13630 VDD.n7771 GND 0.001706f
C13631 VDD.n7772 GND 0.001706f
C13632 VDD.n7773 GND 0.001706f
C13633 VDD.n7774 GND 0.001706f
C13634 VDD.n7775 GND 0.001706f
C13635 VDD.t507 GND 0.119161f
C13636 VDD.n7776 GND 0.001706f
C13637 VDD.n7777 GND 0.001706f
C13638 VDD.n7778 GND 0.001706f
C13639 VDD.n7779 GND 0.238321f
C13640 VDD.n7780 GND 0.001706f
C13641 VDD.n7781 GND 0.001706f
C13642 VDD.n7782 GND 0.001706f
C13643 VDD.n7783 GND 0.001706f
C13644 VDD.n7784 GND 0.001706f
C13645 VDD.n7785 GND 0.001706f
C13646 VDD.t130 GND 0.119161f
C13647 VDD.n7786 GND 0.001706f
C13648 VDD.n7787 GND 0.001706f
C13649 VDD.n7788 GND 0.001706f
C13650 VDD.n7789 GND 0.176989f
C13651 VDD.n7790 GND 0.001706f
C13652 VDD.n7791 GND 0.001706f
C13653 VDD.n7792 GND 0.001706f
C13654 VDD.n7793 GND 0.138437f
C13655 VDD.n7794 GND 0.001706f
C13656 VDD.n7795 GND 0.001706f
C13657 VDD.n7796 GND 0.001706f
C13658 VDD.t283 GND 0.119161f
C13659 VDD.n7797 GND 0.001706f
C13660 VDD.n7798 GND 0.001706f
C13661 VDD.n7799 GND 0.001706f
C13662 VDD.n7800 GND 0.215541f
C13663 VDD.n7801 GND 0.001706f
C13664 VDD.n7802 GND 0.003781f
C13665 VDD.n7803 GND 0.003781f
C13666 VDD.t179 GND 0.119161f
C13667 VDD.n7804 GND 0.001706f
C13668 VDD.n7805 GND 0.003781f
C13669 VDD.n7813 GND 0.001706f
C13670 VDD.n7814 GND 0.001706f
C13671 VDD.n7815 GND 0.001706f
C13672 VDD.n7816 GND 0.001706f
C13673 VDD.n7817 GND 0.001706f
C13674 VDD.n7818 GND 0.001706f
C13675 VDD.n7819 GND 0.001706f
C13676 VDD.n7820 GND 0.001706f
C13677 VDD.n7821 GND 0.001706f
C13678 VDD.n7822 GND 0.001706f
C13679 VDD.n7823 GND 0.001706f
C13680 VDD.n7824 GND 0.001706f
C13681 VDD.n7825 GND 0.001706f
C13682 VDD.n7826 GND 0.001706f
C13683 VDD.n7827 GND 0.001706f
C13684 VDD.n7828 GND 0.001706f
C13685 VDD.n7829 GND 0.001706f
C13686 VDD.n7830 GND 0.001706f
C13687 VDD.n7831 GND 0.001706f
C13688 VDD.n7832 GND 0.001706f
C13689 VDD.n7833 GND 0.001706f
C13690 VDD.n7834 GND 0.001706f
C13691 VDD.n7835 GND 0.001706f
C13692 VDD.n7836 GND 0.001706f
C13693 VDD.n7837 GND 0.003781f
C13694 VDD.n7838 GND 0.003795f
C13695 VDD.n7839 GND 0.003795f
C13696 VDD.n7840 GND 0.001706f
C13697 VDD.n7841 GND 0.001706f
C13698 VDD.n7842 GND 0.001706f
C13699 VDD.n7843 GND 0.001706f
C13700 VDD.n7844 GND 0.001706f
C13701 VDD.n7845 GND 0.001706f
C13702 VDD.n7846 GND 0.001706f
C13703 VDD.n7847 GND 0.001706f
C13704 VDD.n7848 GND 0.001706f
C13705 VDD.n7849 GND 0.001706f
C13706 VDD.n7850 GND 0.001706f
C13707 VDD.n7851 GND 0.001706f
C13708 VDD.n7852 GND 0.001706f
C13709 VDD.n7853 GND 0.001706f
C13710 VDD.n7854 GND 0.001706f
C13711 VDD.n7855 GND 0.001706f
C13712 VDD.n7856 GND 0.001706f
C13713 VDD.n7857 GND 0.001706f
C13714 VDD.n7858 GND 0.001706f
C13715 VDD.n7859 GND 0.001706f
C13716 VDD.n7860 GND 0.001706f
C13717 VDD.n7861 GND 0.001706f
C13718 VDD.n7862 GND 0.001706f
C13719 VDD.n7863 GND 0.001706f
C13720 VDD.n7864 GND 0.001706f
C13721 VDD.n7865 GND 0.001706f
C13722 VDD.n7866 GND 0.001706f
C13723 VDD.n7867 GND 0.001706f
C13724 VDD.n7868 GND 0.003795f
C13725 VDD.n7869 GND 0.003795f
C13726 VDD.n7871 GND 0.382015f
C13727 VDD.n7872 GND 0.315425f
C13728 VDD.n7873 GND 0.141941f
C13729 VDD.n7874 GND 0.001706f
C13730 VDD.n7875 GND 0.001706f
C13731 VDD.n7876 GND 0.001706f
C13732 VDD.n7877 GND 0.001706f
C13733 VDD.n7878 GND 0.001706f
C13734 VDD.n7879 GND 0.180493f
C13735 VDD.t169 GND 0.119161f
C13736 VDD.n7880 GND 0.176989f
C13737 VDD.n7881 GND 0.219045f
C13738 VDD.n7882 GND 0.001706f
C13739 VDD.n7883 GND 0.001706f
C13740 VDD.n7884 GND 0.001706f
C13741 VDD.n7885 GND 0.001706f
C13742 VDD.n7886 GND 0.001706f
C13743 VDD.n7887 GND 0.238321f
C13744 VDD.n7888 GND 0.138437f
C13745 VDD.t509 GND 0.119161f
C13746 VDD.n7889 GND 0.219045f
C13747 VDD.n7890 GND 0.001706f
C13748 VDD.n7891 GND 0.001706f
C13749 VDD.n7892 GND 0.001706f
C13750 VDD.n7893 GND 0.001706f
C13751 VDD.n7894 GND 0.001706f
C13752 VDD.n7895 GND 0.180493f
C13753 VDD.n7896 GND 0.215541f
C13754 VDD.t322 GND 0.119161f
C13755 VDD.n7897 GND 0.141941f
C13756 VDD.n7898 GND 0.001706f
C13757 VDD.n7899 GND 0.001706f
C13758 VDD.n7900 GND 0.001706f
C13759 VDD.n7901 GND 0.001706f
C13760 VDD.n7902 GND 0.001706f
C13761 VDD.n7903 GND 0.134932f
C13762 VDD.t268 GND 0.119161f
C13763 VDD.n7904 GND 0.22255f
C13764 VDD.n7905 GND 0.173484f
C13765 VDD.n7906 GND 0.001706f
C13766 VDD.n7907 GND 0.001706f
C13767 VDD.n7908 GND 0.001706f
C13768 VDD.n7909 GND 0.001706f
C13769 VDD.n7910 GND 0.001706f
C13770 VDD.n7911 GND 0.212036f
C13771 VDD.n7912 GND 0.001706f
C13772 VDD.n7913 GND 0.001706f
C13773 VDD.n7914 GND 0.001706f
C13774 VDD.n7915 GND 0.001706f
C13775 VDD.n7916 GND 0.001706f
C13776 VDD.n7917 GND 0.001029f
C13777 VDD.n7918 GND 0.001706f
C13778 VDD.n7919 GND 0.001706f
C13779 VDD.n7920 GND 9.03e-19
C13780 VDD.n7921 GND 8.53e-19
C13781 VDD.n7922 GND 0.005502f
C13782 VDD.n7923 GND 0.002444f
C13783 VDD.n7924 GND 8.53e-19
C13784 VDD.n7925 GND 9.03e-19
C13785 VDD.n7926 GND 0.001706f
C13786 VDD.n7927 GND 0.001706f
C13787 VDD.n7928 GND 9.03e-19
C13788 VDD.n7929 GND 8.53e-19
C13789 VDD.n7930 GND 9.03e-19
C13790 VDD.n7931 GND 8.53e-19
C13791 VDD.n7932 GND 0.002444f
C13792 VDD.n7933 GND 0.002444f
C13793 VDD.n7934 GND 8.53e-19
C13794 VDD.n7935 GND 9.03e-19
C13795 VDD.n7936 GND 8.53e-19
C13796 VDD.n7937 GND 0.001706f
C13797 VDD.n7938 GND 9.03e-19
C13798 VDD.n7939 GND 8.53e-19
C13799 VDD.n7940 GND 0.002444f
C13800 VDD.n7941 GND 0.002375f
C13801 VDD.n7942 GND 8.53e-19
C13802 VDD.n7943 GND 9.03e-19
C13803 VDD.n7944 GND 0.001706f
C13804 VDD.n7945 GND 0.087618f
C13805 VDD.n7946 GND 0.001706f
C13806 VDD.t46 GND 0.117408f
C13807 VDD.n7947 GND 0.054323f
C13808 VDD.n7948 GND 0.001706f
C13809 VDD.n7949 GND 0.001706f
C13810 VDD.n7950 GND 0.001706f
C13811 VDD.n7951 GND 0.001706f
C13812 VDD.n7952 GND 0.001706f
C13813 VDD.n7953 GND 0.001706f
C13814 VDD.n7954 GND 0.001706f
C13815 VDD.n7955 GND 0.001706f
C13816 VDD.n7956 GND 0.001706f
C13817 VDD.n7957 GND 0.001706f
C13818 VDD.n7958 GND 0.001706f
C13819 VDD.t40 GND 0.117408f
C13820 VDD.n7959 GND 0.02979f
C13821 VDD.n7960 GND 0.001706f
C13822 VDD.n7961 GND 0.001706f
C13823 VDD.n7962 GND 0.001706f
C13824 VDD.n7963 GND 0.001706f
C13825 VDD.n7964 GND 0.001706f
C13826 VDD.t214 GND 0.117408f
C13827 VDD.n7965 GND 0.068342f
C13828 VDD.n7966 GND 0.001706f
C13829 VDD.n7967 GND 0.001706f
C13830 VDD.n7968 GND 0.001706f
C13831 VDD.n7969 GND 0.001706f
C13832 VDD.n7970 GND 0.001706f
C13833 VDD.n7971 GND 0.001706f
C13834 VDD.n7972 GND 0.001706f
C13835 VDD.n7973 GND 0.001706f
C13836 VDD.n7974 GND 0.001706f
C13837 VDD.n7975 GND 0.001706f
C13838 VDD.n7976 GND 0.001706f
C13839 VDD.n7977 GND 0.001706f
C13840 VDD.n7978 GND 0.001706f
C13841 VDD.n7979 GND 0.001706f
C13842 VDD.n7980 GND 0.001706f
C13843 VDD.n7981 GND 0.001706f
C13844 VDD.n7982 GND 0.001706f
C13845 VDD.n7983 GND 0.001706f
C13846 VDD.n7984 GND 0.001706f
C13847 VDD.n7985 GND 0.001706f
C13848 VDD.n7986 GND 0.001706f
C13849 VDD.n7987 GND 0.001706f
C13850 VDD.n7988 GND 0.001706f
C13851 VDD.n7989 GND 0.001706f
C13852 VDD.n7990 GND 0.001706f
C13853 VDD.n7991 GND 0.001706f
C13854 VDD.n7992 GND 0.001706f
C13855 VDD.n7993 GND 0.001706f
C13856 VDD.n7994 GND 0.001706f
C13857 VDD.n7995 GND 0.003727f
C13858 VDD.n7996 GND 0.003723f
C13859 VDD.n7997 GND 0.001706f
C13860 VDD.n7998 GND 0.001706f
C13861 VDD.t341 GND 0.117408f
C13862 VDD.n7999 GND 0.106894f
C13863 VDD.n8000 GND 0.001706f
C13864 VDD.n8001 GND 0.001706f
C13865 VDD.n8002 GND 0.003723f
C13866 VDD.n8003 GND 0.003727f
C13867 VDD.n8004 GND 0.003727f
C13868 VDD.n8005 GND 0.001706f
C13869 VDD.n8006 GND 0.001706f
C13870 VDD.n8007 GND 0.001706f
C13871 VDD.n8008 GND 0.001706f
C13872 VDD.n8009 GND 0.001706f
C13873 VDD.n8010 GND 0.001706f
C13874 VDD.n8011 GND 0.001706f
C13875 VDD.n8012 GND 0.001706f
C13876 VDD.n8013 GND 0.001706f
C13877 VDD.n8014 GND 0.001706f
C13878 VDD.n8015 GND 0.001706f
C13879 VDD.n8016 GND 0.001706f
C13880 VDD.n8017 GND 0.001706f
C13881 VDD.n8018 GND 0.001706f
C13882 VDD.n8019 GND 0.001706f
C13883 VDD.n8020 GND 0.001706f
C13884 VDD.n8021 GND 0.001706f
C13885 VDD.n8022 GND 0.001706f
C13886 VDD.n8023 GND 0.001706f
C13887 VDD.n8024 GND 0.001706f
C13888 VDD.n8025 GND 0.001706f
C13889 VDD.n8026 GND 0.001706f
C13890 VDD.n8027 GND 0.001706f
C13891 VDD.n8028 GND 0.001706f
C13892 VDD.n8029 GND 0.001706f
C13893 VDD.n8030 GND 0.001706f
C13894 VDD.n8031 GND 0.001706f
C13895 VDD.n8032 GND 0.001706f
C13896 VDD.n8033 GND 0.001706f
C13897 VDD.n8035 GND 0.119161f
C13898 VDD.n8037 GND 0.001706f
C13899 VDD.n8038 GND 0.001706f
C13900 VDD.n8039 GND 0.003727f
C13901 VDD.n8040 GND 0.003723f
C13902 VDD.n8041 GND 0.003723f
C13903 VDD.n8042 GND 0.119161f
C13904 VDD.n8043 GND 0.003723f
C13905 VDD.n8044 GND 0.003723f
C13906 VDD.n8045 GND 0.001706f
C13907 VDD.n8046 GND 0.001706f
C13908 VDD.n8047 GND 0.001706f
C13909 VDD.n8048 GND 0.08937f
C13910 VDD.n8049 GND 0.001706f
C13911 VDD.n8050 GND 0.001706f
C13912 VDD.n8051 GND 0.001706f
C13913 VDD.n8052 GND 0.001706f
C13914 VDD.n8053 GND 0.001706f
C13915 VDD.n8054 GND 0.050818f
C13916 VDD.n8055 GND 0.001706f
C13917 VDD.n8056 GND 0.001706f
C13918 VDD.n8057 GND 0.001706f
C13919 VDD.n8058 GND 0.001706f
C13920 VDD.n8059 GND 0.001706f
C13921 VDD.n8060 GND 0.012266f
C13922 VDD.n8061 GND 0.119161f
C13923 VDD.n8062 GND 0.001706f
C13924 VDD.n8063 GND 9.03e-19
C13925 VDD.n8064 GND 8.53e-19
C13926 VDD.n8065 GND 0.002444f
C13927 VDD.n8066 GND 0.002444f
C13928 VDD.n8067 GND 8.53e-19
C13929 VDD.n8068 GND 9.03e-19
C13930 VDD.n8069 GND 0.001706f
C13931 VDD.n8070 GND 0.028038f
C13932 VDD.t61 GND 0.117408f
C13933 VDD.n8071 GND 0.092875f
C13934 VDD.n8072 GND 0.001706f
C13935 VDD.n8073 GND 0.00133f
C13936 VDD.n8074 GND 0.003632f
C13937 VDD.n8075 GND 0.008749f
C13938 VDD.n8076 GND 0.001706f
C13939 VDD.n8077 GND 0.071847f
C13940 VDD.n8078 GND 0.001706f
C13941 VDD.n8079 GND 0.001706f
C13942 VDD.n8080 GND 0.001706f
C13943 VDD.n8081 GND 0.001129f
C13944 VDD.n8082 GND 0.001706f
C13945 VDD.n8083 GND 0.033295f
C13946 VDD.n8084 GND 0.105142f
C13947 VDD.n8085 GND 0.001706f
C13948 VDD.n8086 GND 9.03e-19
C13949 VDD.n8087 GND 8.53e-19
C13950 VDD.n8088 GND 0.002444f
C13951 VDD.n8089 GND 0.002316f
C13952 VDD.n8090 GND 8.53e-19
C13953 VDD.n8091 GND 9.03e-19
C13954 VDD.n8092 GND 0.001706f
C13955 VDD.n8093 GND 0.007009f
C13956 VDD.n8094 GND 0.001706f
C13957 VDD.n8095 GND 9.03e-19
C13958 VDD.n8096 GND 8.53e-19
C13959 VDD.n8097 GND 0.010359f
C13960 VDD.n8098 GND 0.010359f
C13961 VDD.n8099 GND 8.53e-19
C13962 VDD.n8100 GND 9.03e-19
C13963 VDD.n8101 GND 0.001706f
C13964 VDD.n8102 GND 0.09638f
C13965 VDD.n8103 GND 0.045561f
C13966 VDD.n8104 GND 0.001706f
C13967 VDD.n8105 GND 8.78e-19
C13968 VDD.n8106 GND 8.53e-19
C13969 VDD.n8107 GND 0.01746f
C13970 VDD.n8108 GND 0.102225f
C13971 VDD.n8109 GND 0.601507f
C13972 VDD.n8110 GND 0.102225f
C13973 VDD.n8111 GND 0.014122f
C13974 VDD.n8112 GND 8.53e-19
C13975 VDD.n8113 GND 8.78e-19
C13976 VDD.n8114 GND 8.78e-19
C13977 VDD.n8115 GND 0.001706f
C13978 VDD.n8116 GND 0.115656f
C13979 VDD.n8117 GND 0.001706f
C13980 VDD.n8118 GND 8.78e-19
C13981 VDD.n8119 GND 8.53e-19
C13982 VDD.n8120 GND 0.010359f
C13983 VDD.n8121 GND 0.010359f
C13984 VDD.n8122 GND 8.53e-19
C13985 VDD.n8123 GND 9.03e-19
C13986 VDD.n8124 GND 0.001706f
C13987 VDD.n8125 GND 0.005257f
C13988 VDD.n8126 GND 0.001706f
C13989 VDD.n8127 GND 0.008303f
C13990 VDD.n8128 GND 0.072346f
C13991 VDD.n8129 GND 1.79982f
C13992 VDD.n8130 GND 0.073151f
C13993 VDD.n8131 GND 0.002244f
C13994 VDD.t298 GND 0.010699f
C13995 VDD.t21 GND 0.010699f
C13996 VDD.n8132 GND 0.022031f
C13997 VDD.n8133 GND 9.03e-19
C13998 VDD.n8134 GND 0.001516f
C13999 VDD.n8135 GND 8.53e-19
C14000 VDD.n8136 GND 0.002454f
C14001 VDD.n8137 GND 0.002363f
C14002 VDD.n8138 GND 8.53e-19
C14003 VDD.n8139 GND 9.03e-19
C14004 VDD.n8140 GND 0.001972f
C14005 VDD.n8141 GND 0.001783f
C14006 VDD.n8142 GND 0.044032f
C14007 VDD.n8143 GND 2.75612f
C14008 VDD.n8144 GND 26.031f
C14009 VDD.n8145 GND 7.66073f
C14010 VDD.n8146 GND 2.36108f
C14011 VDD.n8147 GND 1.88886f
C14012 VDD.n8148 GND 2.36108f
C14013 VDD.n8150 GND 1.88886f
C14014 VDD.n8151 GND 43.9751f
C14015 VDD.n8152 GND 43.9751f
C14016 VDD.n8154 GND 1.88886f
C14017 VDD.n8155 GND 44.5653f
C14018 VDD.n8157 GND 1.47567f
C14019 a_153429_n11365.n0 GND 0.147031f
C14020 a_153429_n11365.n1 GND 0.101858f
C14021 a_153429_n11365.n2 GND 0.101858f
C14022 a_153429_n11365.n3 GND 0.100615f
C14023 a_153429_n11365.n4 GND 0.101858f
C14024 a_153429_n11365.n5 GND 0.10814f
C14025 a_153429_n11365.n6 GND 0.101858f
C14026 a_153429_n11365.n7 GND 0.101858f
C14027 a_153429_n11365.n8 GND 0.101858f
C14028 a_153429_n11365.n9 GND 0.101858f
C14029 a_153429_n11365.n10 GND 0.101858f
C14030 a_153429_n11365.n11 GND 0.101858f
C14031 a_153429_n11365.n12 GND 0.101858f
C14032 a_153429_n11365.n13 GND 0.101858f
C14033 a_153429_n11365.n14 GND 0.101858f
C14034 a_153429_n11365.n15 GND 0.101858f
C14035 a_153429_n11365.n16 GND 0.101858f
C14036 a_153429_n11365.n17 GND 0.101858f
C14037 a_153429_n11365.n18 GND 0.101858f
C14038 a_153429_n11365.n19 GND 0.101858f
C14039 a_153429_n11365.n20 GND 0.101858f
C14040 a_153429_n11365.t31 GND 0.906218f
C14041 a_153429_n11365.t29 GND 0.808763f
C14042 a_153429_n11365.n21 GND 8.96654f
C14043 a_153429_n11365.n22 GND 0.592907f
C14044 a_153429_n11365.n23 GND 0.150564f
C14045 a_153429_n11365.t54 GND 0.262908f
C14046 a_153429_n11365.n24 GND 0.14687f
C14047 a_153429_n11365.t33 GND 0.262908f
C14048 a_153429_n11365.n25 GND 0.101858f
C14049 a_153429_n11365.n26 GND 0.101858f
C14050 a_153429_n11365.t45 GND 0.262908f
C14051 a_153429_n11365.n27 GND 0.101858f
C14052 a_153429_n11365.t35 GND 0.262908f
C14053 a_153429_n11365.n28 GND 0.101858f
C14054 a_153429_n11365.n29 GND 0.101858f
C14055 a_153429_n11365.t32 GND 0.262908f
C14056 a_153429_n11365.n30 GND 0.101858f
C14057 a_153429_n11365.t68 GND 0.262908f
C14058 a_153429_n11365.n31 GND 0.101858f
C14059 a_153429_n11365.n32 GND 0.101858f
C14060 a_153429_n11365.t49 GND 0.262908f
C14061 a_153429_n11365.n33 GND 0.101146f
C14062 a_153429_n11365.n34 GND 0.032375f
C14063 a_153429_n11365.n35 GND 0.009993f
C14064 a_153429_n11365.n36 GND 0.190843f
C14065 a_153429_n11365.n37 GND 0.004022f
C14066 a_153429_n11365.n38 GND 0.003799f
C14067 a_153429_n11365.n39 GND 0.01296f
C14068 a_153429_n11365.n40 GND 0.004022f
C14069 a_153429_n11365.n41 GND 0.010813f
C14070 a_153429_n11365.n42 GND 0.003799f
C14071 a_153429_n11365.n43 GND 0.014311f
C14072 a_153429_n11365.n44 GND 0.02292f
C14073 a_153429_n11365.n45 GND 0.004022f
C14074 a_153429_n11365.n46 GND 0.003799f
C14075 a_153429_n11365.n47 GND 0.010665f
C14076 a_153429_n11365.n48 GND 0.010883f
C14077 a_153429_n11365.n49 GND 0.003799f
C14078 a_153429_n11365.n50 GND 0.003799f
C14079 a_153429_n11365.n51 GND 0.004022f
C14080 a_153429_n11365.n52 GND 0.01296f
C14081 a_153429_n11365.n53 GND 0.01296f
C14082 a_153429_n11365.t4 GND 0.018603f
C14083 a_153429_n11365.n54 GND 0.030794f
C14084 a_153429_n11365.n55 GND 0.004715f
C14085 a_153429_n11365.n56 GND 0.00972f
C14086 a_153429_n11365.n57 GND 0.01296f
C14087 a_153429_n11365.n58 GND 0.004022f
C14088 a_153429_n11365.n59 GND 0.003799f
C14089 a_153429_n11365.n60 GND 0.010853f
C14090 a_153429_n11365.n61 GND 0.020232f
C14091 a_153429_n11365.n62 GND 2.50714f
C14092 a_153429_n11365.n63 GND 0.032375f
C14093 a_153429_n11365.n64 GND 0.032375f
C14094 a_153429_n11365.n65 GND 0.032375f
C14095 a_153429_n11365.n66 GND 0.009993f
C14096 a_153429_n11365.t2 GND 0.047648f
C14097 a_153429_n11365.t0 GND 0.047648f
C14098 a_153429_n11365.n67 GND 0.101882f
C14099 a_153429_n11365.n68 GND 0.004022f
C14100 a_153429_n11365.n69 GND 0.010813f
C14101 a_153429_n11365.n70 GND 0.006736f
C14102 a_153429_n11365.n71 GND 0.003799f
C14103 a_153429_n11365.n72 GND 0.004022f
C14104 a_153429_n11365.n73 GND 0.003799f
C14105 a_153429_n11365.n74 GND 0.010665f
C14106 a_153429_n11365.n75 GND 0.010883f
C14107 a_153429_n11365.n76 GND 0.003799f
C14108 a_153429_n11365.n77 GND 0.004022f
C14109 a_153429_n11365.n78 GND 0.00887f
C14110 a_153429_n11365.n79 GND 0.006942f
C14111 a_153429_n11365.n80 GND 0.174546f
C14112 a_153429_n11365.n81 GND 0.416899f
C14113 a_153429_n11365.n82 GND 0.009993f
C14114 a_153429_n11365.t3 GND 0.047648f
C14115 a_153429_n11365.t27 GND 0.047648f
C14116 a_153429_n11365.n83 GND 0.101882f
C14117 a_153429_n11365.n84 GND 0.004022f
C14118 a_153429_n11365.n85 GND 0.010813f
C14119 a_153429_n11365.n86 GND 0.006736f
C14120 a_153429_n11365.n87 GND 0.003799f
C14121 a_153429_n11365.n88 GND 0.004022f
C14122 a_153429_n11365.n89 GND 0.003799f
C14123 a_153429_n11365.n90 GND 0.010665f
C14124 a_153429_n11365.n91 GND 0.010883f
C14125 a_153429_n11365.n92 GND 0.003799f
C14126 a_153429_n11365.n93 GND 0.004022f
C14127 a_153429_n11365.n94 GND 0.00887f
C14128 a_153429_n11365.n95 GND 0.006942f
C14129 a_153429_n11365.n96 GND 0.174546f
C14130 a_153429_n11365.n97 GND 0.416899f
C14131 a_153429_n11365.n98 GND 0.009993f
C14132 a_153429_n11365.t30 GND 0.047648f
C14133 a_153429_n11365.t28 GND 0.047648f
C14134 a_153429_n11365.n99 GND 0.101882f
C14135 a_153429_n11365.n100 GND 0.004022f
C14136 a_153429_n11365.n101 GND 0.010813f
C14137 a_153429_n11365.n102 GND 0.006736f
C14138 a_153429_n11365.n103 GND 0.003799f
C14139 a_153429_n11365.n104 GND 0.004022f
C14140 a_153429_n11365.n105 GND 0.003799f
C14141 a_153429_n11365.n106 GND 0.010665f
C14142 a_153429_n11365.n107 GND 0.010883f
C14143 a_153429_n11365.n108 GND 0.003799f
C14144 a_153429_n11365.n109 GND 0.004022f
C14145 a_153429_n11365.n110 GND 0.00887f
C14146 a_153429_n11365.n111 GND 0.006942f
C14147 a_153429_n11365.n112 GND 0.174546f
C14148 a_153429_n11365.n113 GND 2.69459f
C14149 a_153429_n11365.n114 GND 1.78345f
C14150 a_153429_n11365.n115 GND 0.019904f
C14151 a_153429_n11365.n116 GND 0.010813f
C14152 a_153429_n11365.n117 GND 0.003799f
C14153 a_153429_n11365.n118 GND 0.01296f
C14154 a_153429_n11365.n119 GND 0.004022f
C14155 a_153429_n11365.n120 GND 0.003799f
C14156 a_153429_n11365.n121 GND 0.01296f
C14157 a_153429_n11365.n122 GND 0.004022f
C14158 a_153429_n11365.n123 GND 0.031569f
C14159 a_153429_n11365.t10 GND 0.024272f
C14160 a_153429_n11365.n124 GND 0.00972f
C14161 a_153429_n11365.n125 GND 0.004967f
C14162 a_153429_n11365.n126 GND 0.003799f
C14163 a_153429_n11365.n127 GND 0.184412f
C14164 a_153429_n11365.n128 GND 0.01065f
C14165 a_153429_n11365.n129 GND 0.010847f
C14166 a_153429_n11365.n130 GND 0.003799f
C14167 a_153429_n11365.n131 GND 0.004022f
C14168 a_153429_n11365.n132 GND 0.01296f
C14169 a_153429_n11365.n133 GND 0.01296f
C14170 a_153429_n11365.n134 GND 0.004022f
C14171 a_153429_n11365.n135 GND 0.003799f
C14172 a_153429_n11365.n136 GND 0.010295f
C14173 a_153429_n11365.n137 GND 0.010665f
C14174 a_153429_n11365.n138 GND 0.003799f
C14175 a_153429_n11365.n139 GND 0.004022f
C14176 a_153429_n11365.n140 GND 0.025532f
C14177 a_153429_n11365.n141 GND 0.011699f
C14178 a_153429_n11365.n142 GND 0.032375f
C14179 a_153429_n11365.n143 GND 0.606487f
C14180 a_153429_n11365.n144 GND 0.195103f
C14181 a_153429_n11365.n145 GND 0.010813f
C14182 a_153429_n11365.n146 GND 0.003799f
C14183 a_153429_n11365.t7 GND 0.047648f
C14184 a_153429_n11365.n147 GND 0.004022f
C14185 a_153429_n11365.n148 GND 0.004022f
C14186 a_153429_n11365.n149 GND 0.003799f
C14187 a_153429_n11365.n150 GND 0.010665f
C14188 a_153429_n11365.n151 GND 0.010295f
C14189 a_153429_n11365.n152 GND 0.008781f
C14190 a_153429_n11365.n153 GND 0.008619f
C14191 a_153429_n11365.t23 GND 0.047648f
C14192 a_153429_n11365.n154 GND 0.09814f
C14193 a_153429_n11365.n155 GND 0.006736f
C14194 a_153429_n11365.n156 GND 0.032375f
C14195 a_153429_n11365.n157 GND 0.334089f
C14196 a_153429_n11365.n158 GND 0.195103f
C14197 a_153429_n11365.n159 GND 0.010813f
C14198 a_153429_n11365.n160 GND 0.003799f
C14199 a_153429_n11365.t20 GND 0.047648f
C14200 a_153429_n11365.n161 GND 0.004022f
C14201 a_153429_n11365.n162 GND 0.004022f
C14202 a_153429_n11365.n163 GND 0.003799f
C14203 a_153429_n11365.n164 GND 0.010665f
C14204 a_153429_n11365.n165 GND 0.010295f
C14205 a_153429_n11365.n166 GND 0.008781f
C14206 a_153429_n11365.n167 GND 0.008619f
C14207 a_153429_n11365.t6 GND 0.047648f
C14208 a_153429_n11365.n168 GND 0.09814f
C14209 a_153429_n11365.n169 GND 0.006736f
C14210 a_153429_n11365.n170 GND 0.032375f
C14211 a_153429_n11365.n171 GND 0.339019f
C14212 a_153429_n11365.n172 GND 0.195103f
C14213 a_153429_n11365.n173 GND 0.010813f
C14214 a_153429_n11365.n174 GND 0.003799f
C14215 a_153429_n11365.t17 GND 0.047648f
C14216 a_153429_n11365.n175 GND 0.004022f
C14217 a_153429_n11365.n176 GND 0.004022f
C14218 a_153429_n11365.n177 GND 0.003799f
C14219 a_153429_n11365.n178 GND 0.010665f
C14220 a_153429_n11365.n179 GND 0.010295f
C14221 a_153429_n11365.n180 GND 0.008781f
C14222 a_153429_n11365.n181 GND 0.008619f
C14223 a_153429_n11365.t14 GND 0.047648f
C14224 a_153429_n11365.n182 GND 0.09814f
C14225 a_153429_n11365.n183 GND 0.006736f
C14226 a_153429_n11365.n184 GND 0.032375f
C14227 a_153429_n11365.n185 GND 0.334089f
C14228 a_153429_n11365.n186 GND 0.195103f
C14229 a_153429_n11365.n187 GND 0.010813f
C14230 a_153429_n11365.n188 GND 0.003799f
C14231 a_153429_n11365.t12 GND 0.047648f
C14232 a_153429_n11365.n189 GND 0.004022f
C14233 a_153429_n11365.n190 GND 0.004022f
C14234 a_153429_n11365.n191 GND 0.003799f
C14235 a_153429_n11365.n192 GND 0.010665f
C14236 a_153429_n11365.n193 GND 0.010295f
C14237 a_153429_n11365.n194 GND 0.008781f
C14238 a_153429_n11365.n195 GND 0.008619f
C14239 a_153429_n11365.t9 GND 0.047648f
C14240 a_153429_n11365.n196 GND 0.09814f
C14241 a_153429_n11365.n197 GND 0.006736f
C14242 a_153429_n11365.n198 GND 0.032375f
C14243 a_153429_n11365.n199 GND 0.334089f
C14244 a_153429_n11365.n200 GND 0.195103f
C14245 a_153429_n11365.n201 GND 0.010813f
C14246 a_153429_n11365.n202 GND 0.003799f
C14247 a_153429_n11365.t24 GND 0.047648f
C14248 a_153429_n11365.n203 GND 0.004022f
C14249 a_153429_n11365.n204 GND 0.004022f
C14250 a_153429_n11365.n205 GND 0.003799f
C14251 a_153429_n11365.n206 GND 0.010665f
C14252 a_153429_n11365.n207 GND 0.010295f
C14253 a_153429_n11365.n208 GND 0.008781f
C14254 a_153429_n11365.n209 GND 0.008619f
C14255 a_153429_n11365.t25 GND 0.047648f
C14256 a_153429_n11365.n210 GND 0.09814f
C14257 a_153429_n11365.n211 GND 0.006736f
C14258 a_153429_n11365.n212 GND 0.032375f
C14259 a_153429_n11365.n213 GND 0.334089f
C14260 a_153429_n11365.n214 GND 0.195103f
C14261 a_153429_n11365.n215 GND 0.010813f
C14262 a_153429_n11365.n216 GND 0.003799f
C14263 a_153429_n11365.t19 GND 0.047648f
C14264 a_153429_n11365.n217 GND 0.004022f
C14265 a_153429_n11365.n218 GND 0.004022f
C14266 a_153429_n11365.n219 GND 0.003799f
C14267 a_153429_n11365.n220 GND 0.010665f
C14268 a_153429_n11365.n221 GND 0.010295f
C14269 a_153429_n11365.n222 GND 0.008781f
C14270 a_153429_n11365.n223 GND 0.008619f
C14271 a_153429_n11365.t16 GND 0.047648f
C14272 a_153429_n11365.n224 GND 0.09814f
C14273 a_153429_n11365.n225 GND 0.006736f
C14274 a_153429_n11365.n226 GND 0.032375f
C14275 a_153429_n11365.n227 GND 0.334089f
C14276 a_153429_n11365.n228 GND 0.195103f
C14277 a_153429_n11365.n229 GND 0.010813f
C14278 a_153429_n11365.n230 GND 0.003799f
C14279 a_153429_n11365.t15 GND 0.047648f
C14280 a_153429_n11365.n231 GND 0.004022f
C14281 a_153429_n11365.n232 GND 0.004022f
C14282 a_153429_n11365.n233 GND 0.003799f
C14283 a_153429_n11365.n234 GND 0.010665f
C14284 a_153429_n11365.n235 GND 0.010295f
C14285 a_153429_n11365.n236 GND 0.008781f
C14286 a_153429_n11365.n237 GND 0.008619f
C14287 a_153429_n11365.t13 GND 0.047648f
C14288 a_153429_n11365.n238 GND 0.09814f
C14289 a_153429_n11365.n239 GND 0.006736f
C14290 a_153429_n11365.n240 GND 0.032375f
C14291 a_153429_n11365.n241 GND 0.339019f
C14292 a_153429_n11365.n242 GND 0.195103f
C14293 a_153429_n11365.n243 GND 0.010813f
C14294 a_153429_n11365.n244 GND 0.003799f
C14295 a_153429_n11365.t22 GND 0.047648f
C14296 a_153429_n11365.n245 GND 0.004022f
C14297 a_153429_n11365.n246 GND 0.004022f
C14298 a_153429_n11365.n247 GND 0.003799f
C14299 a_153429_n11365.n248 GND 0.010665f
C14300 a_153429_n11365.n249 GND 0.010295f
C14301 a_153429_n11365.n250 GND 0.008781f
C14302 a_153429_n11365.n251 GND 0.008619f
C14303 a_153429_n11365.t8 GND 0.047648f
C14304 a_153429_n11365.n252 GND 0.09814f
C14305 a_153429_n11365.n253 GND 0.006736f
C14306 a_153429_n11365.n254 GND 0.032375f
C14307 a_153429_n11365.n255 GND 0.334089f
C14308 a_153429_n11365.n256 GND 0.195103f
C14309 a_153429_n11365.n257 GND 0.010813f
C14310 a_153429_n11365.n258 GND 0.003799f
C14311 a_153429_n11365.t26 GND 0.047648f
C14312 a_153429_n11365.n259 GND 0.004022f
C14313 a_153429_n11365.n260 GND 0.004022f
C14314 a_153429_n11365.n261 GND 0.003799f
C14315 a_153429_n11365.n262 GND 0.010665f
C14316 a_153429_n11365.n263 GND 0.010295f
C14317 a_153429_n11365.n264 GND 0.008781f
C14318 a_153429_n11365.n265 GND 0.008619f
C14319 a_153429_n11365.t21 GND 0.047648f
C14320 a_153429_n11365.n266 GND 0.09814f
C14321 a_153429_n11365.n267 GND 0.006736f
C14322 a_153429_n11365.n268 GND 0.032375f
C14323 a_153429_n11365.n269 GND 0.334089f
C14324 a_153429_n11365.n270 GND 0.195103f
C14325 a_153429_n11365.n271 GND 0.010813f
C14326 a_153429_n11365.n272 GND 0.003799f
C14327 a_153429_n11365.t18 GND 0.047648f
C14328 a_153429_n11365.n273 GND 0.004022f
C14329 a_153429_n11365.n274 GND 0.004022f
C14330 a_153429_n11365.n275 GND 0.003799f
C14331 a_153429_n11365.n276 GND 0.010665f
C14332 a_153429_n11365.n277 GND 0.010295f
C14333 a_153429_n11365.n278 GND 0.008781f
C14334 a_153429_n11365.n279 GND 0.008619f
C14335 a_153429_n11365.t11 GND 0.047648f
C14336 a_153429_n11365.n280 GND 0.09814f
C14337 a_153429_n11365.n281 GND 0.006736f
C14338 a_153429_n11365.n282 GND 0.032375f
C14339 a_153429_n11365.n283 GND 0.771206f
C14340 a_153429_n11365.n284 GND 1.77892f
C14341 a_153429_n11365.n285 GND 0.10784f
C14342 a_153429_n11365.t40 GND 0.262908f
C14343 a_153429_n11365.n286 GND 0.104296f
C14344 a_153429_n11365.n287 GND 0.101194f
C14345 a_153429_n11365.t59 GND 0.262908f
C14346 a_153429_n11365.n288 GND 0.101858f
C14347 a_153429_n11365.t48 GND 0.262908f
C14348 a_153429_n11365.n289 GND 0.101858f
C14349 a_153429_n11365.n290 GND 0.101858f
C14350 a_153429_n11365.t38 GND 0.262908f
C14351 a_153429_n11365.n291 GND 0.101858f
C14352 a_153429_n11365.t66 GND 0.262908f
C14353 a_153429_n11365.n292 GND 0.101858f
C14354 a_153429_n11365.n293 GND 0.101858f
C14355 a_153429_n11365.t58 GND 0.262908f
C14356 a_153429_n11365.n294 GND 0.101858f
C14357 a_153429_n11365.t52 GND 0.262908f
C14358 a_153429_n11365.n295 GND 0.101858f
C14359 a_153429_n11365.n296 GND 0.101858f
C14360 a_153429_n11365.t65 GND 0.262908f
C14361 a_153429_n11365.n297 GND 0.101858f
C14362 a_153429_n11365.t55 GND 0.262908f
C14363 a_153429_n11365.n298 GND 0.101858f
C14364 a_153429_n11365.n299 GND 0.101858f
C14365 a_153429_n11365.t34 GND 0.262908f
C14366 a_153429_n11365.n300 GND 0.101858f
C14367 a_153429_n11365.t70 GND 0.262908f
C14368 a_153429_n11365.n301 GND 0.101858f
C14369 a_153429_n11365.n302 GND 0.101858f
C14370 a_153429_n11365.t67 GND 0.262908f
C14371 a_153429_n11365.n303 GND 0.101858f
C14372 a_153429_n11365.t62 GND 0.262908f
C14373 a_153429_n11365.n304 GND 0.101858f
C14374 a_153429_n11365.n305 GND 0.101858f
C14375 a_153429_n11365.t57 GND 0.262908f
C14376 a_153429_n11365.n306 GND 0.101858f
C14377 a_153429_n11365.t51 GND 0.262908f
C14378 a_153429_n11365.n307 GND 0.101858f
C14379 a_153429_n11365.n308 GND 0.101858f
C14380 a_153429_n11365.t42 GND 0.262908f
C14381 a_153429_n11365.n309 GND 0.101858f
C14382 a_153429_n11365.t37 GND 0.262908f
C14383 a_153429_n11365.n310 GND 0.101858f
C14384 a_153429_n11365.n311 GND 0.101858f
C14385 a_153429_n11365.t71 GND 0.262908f
C14386 a_153429_n11365.n312 GND 0.101858f
C14387 a_153429_n11365.t69 GND 0.262908f
C14388 a_153429_n11365.n313 GND 0.101858f
C14389 a_153429_n11365.n314 GND 0.101858f
C14390 a_153429_n11365.t47 GND 0.262908f
C14391 a_153429_n11365.n315 GND 0.101858f
C14392 a_153429_n11365.t64 GND 0.262908f
C14393 a_153429_n11365.n316 GND 0.101858f
C14394 a_153429_n11365.n317 GND 0.101858f
C14395 a_153429_n11365.t53 GND 0.262908f
C14396 a_153429_n11365.n318 GND 0.101858f
C14397 a_153429_n11365.t44 GND 0.262908f
C14398 a_153429_n11365.n319 GND 0.101858f
C14399 a_153429_n11365.n320 GND 0.101858f
C14400 a_153429_n11365.t39 GND 0.262908f
C14401 a_153429_n11365.n321 GND 0.101858f
C14402 a_153429_n11365.t63 GND 0.262908f
C14403 a_153429_n11365.n322 GND 0.100899f
C14404 a_153429_n11365.n323 GND 0.104821f
C14405 a_153429_n11365.t60 GND 0.262908f
C14406 a_153429_n11365.n324 GND 0.101858f
C14407 a_153429_n11365.t50 GND 0.262908f
C14408 a_153429_n11365.n325 GND 0.101858f
C14409 a_153429_n11365.n326 GND 0.101858f
C14410 a_153429_n11365.t41 GND 0.262908f
C14411 a_153429_n11365.n327 GND 0.101858f
C14412 a_153429_n11365.t36 GND 0.262908f
C14413 a_153429_n11365.n328 GND 0.101858f
C14414 a_153429_n11365.n329 GND 0.101858f
C14415 a_153429_n11365.t61 GND 0.262908f
C14416 a_153429_n11365.n330 GND 0.101858f
C14417 a_153429_n11365.t56 GND 0.262908f
C14418 a_153429_n11365.n331 GND 0.101858f
C14419 a_153429_n11365.n332 GND 0.101858f
C14420 a_153429_n11365.t46 GND 0.262908f
C14421 a_153429_n11365.n333 GND 0.101858f
C14422 a_153429_n11365.t43 GND 0.262908f
C14423 a_153429_n11365.n334 GND 0.15071f
C14424 a_153429_n11365.n335 GND 0.594573f
C14425 a_153429_n11365.t5 GND 0.812363f
C14426 a_153429_n11365.n336 GND 8.85972f
C14427 a_153429_n11365.t1 GND 0.909211f
C14428 a_156330_n13996.n0 GND 0.777917f
C14429 a_156330_n13996.n1 GND 1.18353f
C14430 a_156330_n13996.n2 GND 1.24966f
C14431 a_156330_n13996.n3 GND 0.552541f
C14432 a_156330_n13996.n4 GND 0.552541f
C14433 a_156330_n13996.n5 GND 0.905006f
C14434 a_156330_n13996.n6 GND 0.820308f
C14435 a_156330_n13996.n7 GND 0.552541f
C14436 a_156330_n13996.n8 GND 0.552541f
C14437 a_156330_n13996.n9 GND 0.552541f
C14438 a_156330_n13996.t68 GND 0.356545f
C14439 a_156330_n13996.n10 GND 0.682063f
C14440 a_156330_n13996.n11 GND 0.27627f
C14441 a_156330_n13996.n12 GND 1.64606f
C14442 a_156330_n13996.n13 GND 1.68345f
C14443 a_156330_n13996.n14 GND 1.4598f
C14444 a_156330_n13996.n15 GND 0.06876f
C14445 a_156330_n13996.n16 GND 0.153971f
C14446 a_156330_n13996.n17 GND 0.194469f
C14447 a_156330_n13996.n18 GND 0.194469f
C14448 a_156330_n13996.n19 GND 0.93221f
C14449 a_156330_n13996.n20 GND 0.011902f
C14450 a_156330_n13996.n21 GND 0.076964f
C14451 a_156330_n13996.n22 GND 0.011902f
C14452 a_156330_n13996.n23 GND 7.62712f
C14453 a_156330_n13996.t16 GND 0.356545f
C14454 a_156330_n13996.t30 GND 0.356545f
C14455 a_156330_n13996.n24 GND 0.010861f
C14456 a_156330_n13996.n25 GND 0.010861f
C14457 a_156330_n13996.n26 GND 0.086352f
C14458 a_156330_n13996.n27 GND 7.29562f
C14459 a_156330_n13996.n28 GND 0.010345f
C14460 a_156330_n13996.n29 GND 0.010345f
C14461 a_156330_n13996.n30 GND 0.010345f
C14462 a_156330_n13996.n31 GND 1.38286f
C14463 a_156330_n13996.n32 GND 1.3834f
C14464 a_156330_n13996.t47 GND 0.064619f
C14465 a_156330_n13996.t1 GND 0.064619f
C14466 a_156330_n13996.t2 GND 0.064619f
C14467 a_156330_n13996.n33 GND 0.229545f
C14468 a_156330_n13996.t33 GND 0.064619f
C14469 a_156330_n13996.n34 GND 0.005455f
C14470 a_156330_n13996.n35 GND 0.005455f
C14471 a_156330_n13996.n36 GND 0.005455f
C14472 a_156330_n13996.n37 GND 0.005455f
C14473 a_156330_n13996.n38 GND 6.01e-19
C14474 a_156330_n13996.n39 GND 0.005455f
C14475 a_156330_n13996.n40 GND 0.005455f
C14476 a_156330_n13996.n41 GND 0.005455f
C14477 a_156330_n13996.n42 GND 0.005455f
C14478 a_156330_n13996.n43 GND 0.005455f
C14479 a_156330_n13996.t23 GND 0.064619f
C14480 a_156330_n13996.t6 GND 0.356545f
C14481 a_156330_n13996.t25 GND 0.064619f
C14482 a_156330_n13996.n44 GND 0.005455f
C14483 a_156330_n13996.n45 GND 0.005455f
C14484 a_156330_n13996.n46 GND 0.005455f
C14485 a_156330_n13996.n47 GND 0.005455f
C14486 a_156330_n13996.n48 GND 6.01e-19
C14487 a_156330_n13996.n49 GND 0.005455f
C14488 a_156330_n13996.n50 GND 0.005455f
C14489 a_156330_n13996.n51 GND 0.005455f
C14490 a_156330_n13996.n52 GND 0.005152f
C14491 a_156330_n13996.t43 GND 0.071771f
C14492 a_156330_n13996.t21 GND 0.064619f
C14493 a_156330_n13996.n53 GND 0.005455f
C14494 a_156330_n13996.n54 GND 0.006801f
C14495 a_156330_n13996.n55 GND 0.005152f
C14496 a_156330_n13996.n56 GND 0.005455f
C14497 a_156330_n13996.n57 GND 0.005455f
C14498 a_156330_n13996.n58 GND 0.005455f
C14499 a_156330_n13996.n59 GND 6.01e-19
C14500 a_156330_n13996.n60 GND 0.005455f
C14501 a_156330_n13996.n61 GND 0.005455f
C14502 a_156330_n13996.n62 GND 0.005455f
C14503 a_156330_n13996.t35 GND 0.064619f
C14504 a_156330_n13996.t37 GND 0.064619f
C14505 a_156330_n13996.n63 GND 0.005455f
C14506 a_156330_n13996.n64 GND 6.01e-19
C14507 a_156330_n13996.n65 GND 0.005455f
C14508 a_156330_n13996.t27 GND 0.064619f
C14509 a_156330_n13996.t42 GND 0.356724f
C14510 a_156330_n13996.t34 GND 0.356545f
C14511 a_156330_n13996.t14 GND 0.356545f
C14512 a_156330_n13996.t8 GND 0.356545f
C14513 a_156330_n13996.t4 GND 0.356545f
C14514 a_156330_n13996.t40 GND 0.356545f
C14515 a_156330_n13996.t10 GND 0.356545f
C14516 a_156330_n13996.t12 GND 0.356545f
C14517 a_156330_n13996.t18 GND 0.356545f
C14518 a_156330_n13996.t28 GND 0.356545f
C14519 a_156330_n13996.t64 GND 0.356545f
C14520 a_156330_n13996.t22 GND 0.356545f
C14521 a_156330_n13996.t44 GND 0.356666f
C14522 a_156330_n13996.t57 GND 0.356545f
C14523 a_156330_n13996.t54 GND 0.356545f
C14524 a_156330_n13996.t49 GND 0.356545f
C14525 a_156330_n13996.t67 GND 0.356545f
C14526 a_156330_n13996.t53 GND 0.356545f
C14527 a_156330_n13996.t62 GND 0.356545f
C14528 a_156330_n13996.t60 GND 0.356545f
C14529 a_156330_n13996.t59 GND 0.356545f
C14530 a_156330_n13996.t56 GND 0.356545f
C14531 a_156330_n13996.t50 GND 0.356545f
C14532 a_156330_n13996.t51 GND 0.356545f
C14533 a_156330_n13996.t66 GND 0.356545f
C14534 a_156330_n13996.t63 GND 0.356545f
C14535 a_156330_n13996.t61 GND 0.356545f
C14536 a_156330_n13996.t58 GND 0.356545f
C14537 a_156330_n13996.t69 GND 0.356545f
C14538 a_156330_n13996.t55 GND 0.356545f
C14539 a_156330_n13996.t52 GND 0.356545f
C14540 a_156330_n13996.t65 GND 0.356545f
C14541 a_156330_n13996.n66 GND 0.086493f
C14542 a_156330_n13996.t36 GND 0.356545f
C14543 a_156330_n13996.t46 GND 0.064619f
C14544 a_156330_n13996.t48 GND 0.064619f
C14545 a_156330_n13996.n67 GND 0.229545f
C14546 a_156330_n13996.t3 GND 0.07282f
C14547 a_156330_n13996.n68 GND 0.007799f
C14548 a_156330_n13996.n69 GND 0.010154f
C14549 a_156330_n13996.n70 GND 0.010154f
C14550 a_156330_n13996.n71 GND 0.007799f
C14551 a_156330_n13996.n72 GND 0.130706f
C14552 a_156330_n13996.t26 GND 0.356545f
C14553 a_156330_n13996.t20 GND 0.356545f
C14554 a_156330_n13996.n73 GND 0.005152f
C14555 a_156330_n13996.n74 GND 0.005152f
C14556 a_156330_n13996.n75 GND 0.010154f
C14557 a_156330_n13996.n76 GND 0.010154f
C14558 a_156330_n13996.n77 GND 0.005152f
C14559 a_156330_n13996.n78 GND 0.005152f
C14560 a_156330_n13996.n79 GND 0.007501f
C14561 a_156330_n13996.n80 GND 0.12965f
C14562 a_156330_n13996.t15 GND 0.064619f
C14563 a_156330_n13996.t9 GND 0.064619f
C14564 a_156330_n13996.n81 GND 0.16888f
C14565 a_156330_n13996.t5 GND 0.064619f
C14566 a_156330_n13996.t41 GND 0.064619f
C14567 a_156330_n13996.n82 GND 0.16888f
C14568 a_156330_n13996.t29 GND 0.064619f
C14569 a_156330_n13996.t31 GND 0.064619f
C14570 a_156330_n13996.n83 GND 0.16888f
C14571 a_156330_n13996.t19 GND 0.064619f
C14572 a_156330_n13996.t13 GND 0.064619f
C14573 a_156330_n13996.n84 GND 0.16888f
C14574 a_156330_n13996.t11 GND 0.064619f
C14575 a_156330_n13996.t7 GND 0.064619f
C14576 a_156330_n13996.n85 GND 0.16888f
C14577 a_156330_n13996.n86 GND 0.006801f
C14578 a_156330_n13996.t17 GND 0.064619f
C14579 a_156330_n13996.t45 GND 0.064619f
C14580 a_156330_n13996.n87 GND 0.16888f
C14581 a_156330_n13996.n88 GND 0.005152f
C14582 a_156330_n13996.n89 GND 0.005152f
C14583 a_156330_n13996.n90 GND 0.010154f
C14584 a_156330_n13996.n91 GND 0.010154f
C14585 a_156330_n13996.n92 GND 0.005152f
C14586 a_156330_n13996.n93 GND 0.005152f
C14587 a_156330_n13996.n94 GND 0.007501f
C14588 a_156330_n13996.t39 GND 0.064619f
C14589 a_156330_n13996.n95 GND 0.12965f
C14590 a_156330_n13996.t24 GND 0.356545f
C14591 a_156330_n13996.t38 GND 0.356545f
C14592 a_156330_n13996.t32 GND 0.356545f
C14593 a_156330_n13996.n96 GND 0.006801f
C14594 a_156330_n13996.n97 GND 0.005152f
C14595 a_156330_n13996.n98 GND 0.005152f
C14596 a_156330_n13996.n99 GND 0.005152f
C14597 a_156330_n13996.n100 GND 0.010154f
C14598 a_156330_n13996.n101 GND 0.010154f
C14599 a_156330_n13996.n102 GND 0.005152f
C14600 a_156330_n13996.n103 GND 0.005152f
C14601 a_156330_n13996.n104 GND 0.005152f
C14602 a_156330_n13996.n105 GND 0.005152f
C14603 a_156330_n13996.n106 GND 0.005152f
C14604 a_156330_n13996.n107 GND 0.009072f
C14605 a_156330_n13996.n108 GND 0.129348f
C14606 a_156330_n13996.n109 GND 0.229544f
C14607 a_156330_n13996.t0 GND 0.064619f
.ends

