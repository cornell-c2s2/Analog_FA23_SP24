magic
tech sky130A
magscale 1 2
timestamp 1711205355
<< checkpaint >>
rect 8842 209802 11784 209908
rect 8842 209696 12522 209802
rect 8842 209590 13260 209696
rect 8842 1404 13998 209590
rect 8842 1356 14312 1404
rect 8842 1308 14810 1356
rect 8842 -1390 15308 1308
rect 9580 -1496 15308 -1390
rect 10318 -1602 15308 -1496
rect 11056 -1708 15308 -1602
rect 11440 -1756 15308 -1708
rect 11754 -1804 15308 -1756
rect 12252 -1852 15308 -1804
<< error_s >>
rect 10284 208510 10342 208516
rect 10284 208476 10296 208510
rect 10284 208470 10342 208476
rect 11022 208404 11080 208410
rect 11022 208370 11034 208404
rect 11022 208364 11080 208370
rect 11760 208298 11818 208304
rect 11760 208264 11772 208298
rect 11760 208258 11818 208264
rect 10284 195582 10342 195588
rect 10284 195548 10296 195582
rect 10284 195542 10342 195548
rect 10284 195474 10342 195480
rect 11022 195476 11080 195482
rect 10284 195440 10296 195474
rect 11022 195442 11034 195476
rect 10284 195434 10342 195440
rect 11022 195436 11080 195442
rect 11022 195368 11080 195374
rect 11760 195370 11818 195376
rect 11022 195334 11034 195368
rect 11760 195336 11772 195370
rect 11022 195328 11080 195334
rect 11760 195330 11818 195336
rect 11760 195262 11818 195268
rect 11760 195228 11772 195262
rect 11760 195222 11818 195228
rect 10284 182546 10342 182552
rect 10284 182512 10296 182546
rect 10284 182506 10342 182512
rect 10284 182438 10342 182444
rect 11022 182440 11080 182446
rect 10284 182404 10296 182438
rect 11022 182406 11034 182440
rect 10284 182398 10342 182404
rect 11022 182400 11080 182406
rect 11022 182332 11080 182338
rect 11760 182334 11818 182340
rect 11022 182298 11034 182332
rect 11760 182300 11772 182334
rect 11022 182292 11080 182298
rect 11760 182294 11818 182300
rect 11760 182226 11818 182232
rect 11760 182192 11772 182226
rect 11760 182186 11818 182192
rect 10284 169510 10342 169516
rect 10284 169476 10296 169510
rect 10284 169470 10342 169476
rect 10284 169402 10342 169408
rect 11022 169404 11080 169410
rect 10284 169368 10296 169402
rect 11022 169370 11034 169404
rect 10284 169362 10342 169368
rect 11022 169364 11080 169370
rect 11022 169296 11080 169302
rect 11760 169298 11818 169304
rect 11022 169262 11034 169296
rect 11760 169264 11772 169298
rect 11022 169256 11080 169262
rect 11760 169258 11818 169264
rect 11760 169190 11818 169196
rect 11760 169156 11772 169190
rect 11760 169150 11818 169156
rect 10284 156474 10342 156480
rect 10284 156440 10296 156474
rect 10284 156434 10342 156440
rect 10284 156366 10342 156372
rect 11022 156368 11080 156374
rect 10284 156332 10296 156366
rect 11022 156334 11034 156368
rect 10284 156326 10342 156332
rect 11022 156328 11080 156334
rect 11022 156260 11080 156266
rect 11760 156262 11818 156268
rect 11022 156226 11034 156260
rect 11760 156228 11772 156262
rect 11022 156220 11080 156226
rect 11760 156222 11818 156228
rect 11760 156154 11818 156160
rect 11760 156120 11772 156154
rect 11760 156114 11818 156120
rect 10284 143438 10342 143444
rect 10284 143404 10296 143438
rect 10284 143398 10342 143404
rect 10284 143330 10342 143336
rect 11022 143332 11080 143338
rect 10284 143296 10296 143330
rect 11022 143298 11034 143332
rect 10284 143290 10342 143296
rect 11022 143292 11080 143298
rect 11022 143224 11080 143230
rect 11760 143226 11818 143232
rect 11022 143190 11034 143224
rect 11760 143192 11772 143226
rect 11022 143184 11080 143190
rect 11760 143186 11818 143192
rect 11760 143118 11818 143124
rect 11760 143084 11772 143118
rect 11760 143078 11818 143084
rect 10284 130402 10342 130408
rect 10284 130368 10296 130402
rect 10284 130362 10342 130368
rect 10284 130294 10342 130300
rect 11022 130296 11080 130302
rect 10284 130260 10296 130294
rect 11022 130262 11034 130296
rect 10284 130254 10342 130260
rect 11022 130256 11080 130262
rect 11022 130188 11080 130194
rect 11760 130190 11818 130196
rect 11022 130154 11034 130188
rect 11760 130156 11772 130190
rect 11022 130148 11080 130154
rect 11760 130150 11818 130156
rect 11760 130082 11818 130088
rect 11760 130048 11772 130082
rect 11760 130042 11818 130048
rect 10284 117366 10342 117372
rect 10284 117332 10296 117366
rect 10284 117326 10342 117332
rect 10284 117258 10342 117264
rect 11022 117260 11080 117266
rect 10284 117224 10296 117258
rect 11022 117226 11034 117260
rect 10284 117218 10342 117224
rect 11022 117220 11080 117226
rect 11022 117152 11080 117158
rect 11760 117154 11818 117160
rect 11022 117118 11034 117152
rect 11760 117120 11772 117154
rect 11022 117112 11080 117118
rect 11760 117114 11818 117120
rect 11760 117046 11818 117052
rect 11760 117012 11772 117046
rect 11760 117006 11818 117012
rect 10284 104330 10342 104336
rect 10284 104296 10296 104330
rect 10284 104290 10342 104296
rect 10284 104222 10342 104228
rect 11022 104224 11080 104230
rect 10284 104188 10296 104222
rect 11022 104190 11034 104224
rect 10284 104182 10342 104188
rect 11022 104184 11080 104190
rect 11022 104116 11080 104122
rect 11760 104118 11818 104124
rect 11022 104082 11034 104116
rect 11760 104084 11772 104118
rect 11022 104076 11080 104082
rect 11760 104078 11818 104084
rect 11760 104010 11818 104016
rect 11760 103976 11772 104010
rect 11760 103970 11818 103976
rect 10284 91294 10342 91300
rect 10284 91260 10296 91294
rect 10284 91254 10342 91260
rect 10284 91186 10342 91192
rect 11022 91188 11080 91194
rect 10284 91152 10296 91186
rect 11022 91154 11034 91188
rect 10284 91146 10342 91152
rect 11022 91148 11080 91154
rect 11022 91080 11080 91086
rect 11760 91082 11818 91088
rect 11022 91046 11034 91080
rect 11760 91048 11772 91082
rect 11022 91040 11080 91046
rect 11760 91042 11818 91048
rect 11760 90974 11818 90980
rect 11760 90940 11772 90974
rect 11760 90934 11818 90940
rect 10284 78258 10342 78264
rect 10284 78224 10296 78258
rect 10284 78218 10342 78224
rect 10284 78150 10342 78156
rect 11022 78152 11080 78158
rect 10284 78116 10296 78150
rect 11022 78118 11034 78152
rect 10284 78110 10342 78116
rect 11022 78112 11080 78118
rect 11022 78044 11080 78050
rect 11760 78046 11818 78052
rect 11022 78010 11034 78044
rect 11760 78012 11772 78046
rect 11022 78004 11080 78010
rect 11760 78006 11818 78012
rect 11760 77938 11818 77944
rect 11760 77904 11772 77938
rect 11760 77898 11818 77904
rect 10284 65222 10342 65228
rect 10284 65188 10296 65222
rect 10284 65182 10342 65188
rect 10284 65114 10342 65120
rect 11022 65116 11080 65122
rect 10284 65080 10296 65114
rect 11022 65082 11034 65116
rect 10284 65074 10342 65080
rect 11022 65076 11080 65082
rect 11022 65008 11080 65014
rect 11760 65010 11818 65016
rect 11022 64974 11034 65008
rect 11760 64976 11772 65010
rect 11022 64968 11080 64974
rect 11760 64970 11818 64976
rect 11760 64902 11818 64908
rect 11760 64868 11772 64902
rect 11760 64862 11818 64868
rect 10138 53069 10172 53087
rect 9915 52931 9973 52937
rect 9915 52897 9927 52931
rect 9915 52891 9973 52897
rect 9915 46421 9973 46427
rect 9915 46387 9927 46421
rect 9915 46381 9973 46387
rect 9915 46313 9973 46319
rect 9915 46279 9927 46313
rect 9915 46273 9973 46279
rect 9915 39803 9973 39809
rect 9915 39769 9927 39803
rect 9915 39763 9973 39769
rect 9915 39695 9973 39701
rect 9915 39661 9927 39695
rect 9915 39655 9973 39661
rect 9915 33185 9973 33191
rect 9915 33151 9927 33185
rect 9915 33145 9973 33151
rect 9915 33077 9973 33083
rect 9915 33043 9927 33077
rect 9915 33037 9973 33043
rect 9915 26567 9973 26573
rect 9915 26533 9927 26567
rect 9915 26527 9973 26533
rect 9915 26459 9973 26465
rect 9915 26425 9927 26459
rect 9915 26419 9973 26425
rect 9915 19949 9973 19955
rect 9915 19915 9927 19949
rect 9915 19909 9973 19915
rect 9915 19841 9973 19847
rect 9915 19807 9927 19841
rect 9915 19801 9973 19807
rect 9915 13331 9973 13337
rect 9915 13297 9927 13331
rect 9915 13291 9973 13297
rect 9915 13223 9973 13229
rect 9915 13189 9927 13223
rect 9915 13183 9973 13189
rect 9915 6713 9973 6719
rect 9915 6679 9927 6713
rect 9915 6673 9973 6679
rect 9915 6605 9973 6611
rect 9915 6571 9927 6605
rect 9915 6565 9973 6571
rect 1272 717 1303 749
rect 2782 669 2812 701
rect 9769 606 9782 619
rect 3594 573 3625 605
rect 5104 525 5134 557
rect 5916 429 5947 461
rect 7426 381 7456 413
rect 8238 285 8269 317
rect 9733 285 9786 606
rect 9915 95 9973 101
rect 9735 7 9748 41
rect 9769 -27 9782 75
rect 9915 61 9927 95
rect 9915 55 9973 61
rect 10102 -41 10172 53069
rect 10454 52963 10488 52981
rect 10876 52963 10910 52981
rect 10454 52927 10524 52963
rect 10471 52893 10542 52927
rect 10284 52186 10342 52192
rect 10284 52152 10296 52186
rect 10284 52146 10342 52152
rect 10284 52078 10342 52084
rect 10284 52044 10296 52078
rect 10284 52038 10342 52044
rect 10284 39150 10342 39156
rect 10284 39116 10296 39150
rect 10284 39110 10342 39116
rect 10284 39042 10342 39048
rect 10284 39008 10296 39042
rect 10284 39002 10342 39008
rect 10284 26114 10342 26120
rect 10284 26080 10296 26114
rect 10284 26074 10342 26080
rect 10284 26006 10342 26012
rect 10284 25972 10296 26006
rect 10284 25966 10342 25972
rect 10284 13078 10342 13084
rect 10284 13044 10296 13078
rect 10284 13038 10342 13044
rect 10284 12970 10342 12976
rect 10284 12936 10296 12970
rect 10284 12930 10342 12936
rect 10284 42 10342 48
rect 10284 8 10296 42
rect 10284 2 10342 8
rect 10102 -77 10155 -41
rect 10471 -94 10541 52893
rect 10653 52825 10711 52831
rect 10653 52791 10665 52825
rect 10653 52785 10711 52791
rect 10653 46315 10711 46321
rect 10653 46281 10665 46315
rect 10653 46275 10711 46281
rect 10653 46207 10711 46213
rect 10653 46173 10665 46207
rect 10653 46167 10711 46173
rect 10653 39697 10711 39703
rect 10653 39663 10665 39697
rect 10653 39657 10711 39663
rect 10653 39589 10711 39595
rect 10653 39555 10665 39589
rect 10653 39549 10711 39555
rect 10653 33079 10711 33085
rect 10653 33045 10665 33079
rect 10653 33039 10711 33045
rect 10653 32971 10711 32977
rect 10653 32937 10665 32971
rect 10653 32931 10711 32937
rect 10653 26461 10711 26467
rect 10653 26427 10665 26461
rect 10653 26421 10711 26427
rect 10653 26353 10711 26359
rect 10653 26319 10665 26353
rect 10653 26313 10711 26319
rect 10653 19843 10711 19849
rect 10653 19809 10665 19843
rect 10653 19803 10711 19809
rect 10653 19735 10711 19741
rect 10653 19701 10665 19735
rect 10653 19695 10711 19701
rect 10653 13225 10711 13231
rect 10653 13191 10665 13225
rect 10653 13185 10711 13191
rect 10653 13117 10711 13123
rect 10653 13083 10665 13117
rect 10653 13077 10711 13083
rect 10653 6607 10711 6613
rect 10653 6573 10665 6607
rect 10653 6567 10711 6573
rect 10653 6499 10711 6505
rect 10653 6465 10665 6499
rect 10653 6459 10711 6465
rect 10653 -11 10711 -5
rect 10653 -45 10665 -11
rect 10653 -51 10711 -45
rect 10471 -130 10524 -94
rect 10840 -147 10910 52963
rect 11192 52857 11226 52875
rect 11614 52857 11648 52875
rect 11192 52821 11262 52857
rect 11209 52787 11280 52821
rect 11022 52080 11080 52086
rect 11022 52046 11034 52080
rect 11022 52040 11080 52046
rect 11022 51972 11080 51978
rect 11022 51938 11034 51972
rect 11022 51932 11080 51938
rect 11022 39044 11080 39050
rect 11022 39010 11034 39044
rect 11022 39004 11080 39010
rect 11022 38936 11080 38942
rect 11022 38902 11034 38936
rect 11022 38896 11080 38902
rect 11022 26008 11080 26014
rect 11022 25974 11034 26008
rect 11022 25968 11080 25974
rect 11022 25900 11080 25906
rect 11022 25866 11034 25900
rect 11022 25860 11080 25866
rect 11022 12972 11080 12978
rect 11022 12938 11034 12972
rect 11022 12932 11080 12938
rect 11022 12864 11080 12870
rect 11022 12830 11034 12864
rect 11022 12824 11080 12830
rect 11022 -64 11080 -58
rect 11022 -98 11034 -64
rect 11022 -104 11080 -98
rect 10840 -183 10893 -147
rect 11209 -200 11279 52787
rect 11391 52719 11449 52725
rect 11391 52685 11403 52719
rect 11391 52679 11449 52685
rect 11391 46209 11449 46215
rect 11391 46175 11403 46209
rect 11391 46169 11449 46175
rect 11391 46101 11449 46107
rect 11391 46067 11403 46101
rect 11391 46061 11449 46067
rect 11391 39591 11449 39597
rect 11391 39557 11403 39591
rect 11391 39551 11449 39557
rect 11391 39483 11449 39489
rect 11391 39449 11403 39483
rect 11391 39443 11449 39449
rect 11391 32973 11449 32979
rect 11391 32939 11403 32973
rect 11391 32933 11449 32939
rect 11391 32865 11449 32871
rect 11391 32831 11403 32865
rect 11391 32825 11449 32831
rect 11391 26355 11449 26361
rect 11391 26321 11403 26355
rect 11391 26315 11449 26321
rect 11391 26247 11449 26253
rect 11391 26213 11403 26247
rect 11391 26207 11449 26213
rect 11391 19737 11449 19743
rect 11391 19703 11403 19737
rect 11391 19697 11449 19703
rect 11391 19629 11449 19635
rect 11391 19595 11403 19629
rect 11391 19589 11449 19595
rect 11391 13119 11449 13125
rect 11391 13085 11403 13119
rect 11391 13079 11449 13085
rect 11391 13011 11449 13017
rect 11391 12977 11403 13011
rect 11391 12971 11449 12977
rect 11391 6501 11449 6507
rect 11391 6467 11403 6501
rect 11391 6461 11449 6467
rect 11391 6393 11449 6399
rect 11391 6359 11403 6393
rect 11391 6353 11449 6359
rect 11391 -117 11449 -111
rect 11391 -151 11403 -117
rect 11391 -157 11449 -151
rect 11209 -236 11262 -200
rect 11578 -253 11648 52857
rect 11930 52751 11964 52769
rect 11930 52715 12000 52751
rect 11947 52681 12018 52715
rect 11760 51974 11818 51980
rect 11760 51940 11772 51974
rect 11760 51934 11818 51940
rect 11760 51866 11818 51872
rect 11760 51832 11772 51866
rect 11760 51826 11818 51832
rect 11760 38938 11818 38944
rect 11760 38904 11772 38938
rect 11760 38898 11818 38904
rect 11760 38830 11818 38836
rect 11760 38796 11772 38830
rect 11760 38790 11818 38796
rect 11760 25902 11818 25908
rect 11760 25868 11772 25902
rect 11760 25862 11818 25868
rect 11760 25794 11818 25800
rect 11760 25760 11772 25794
rect 11760 25754 11818 25760
rect 11760 12866 11818 12872
rect 11760 12832 11772 12866
rect 11760 12826 11818 12832
rect 11760 12758 11818 12764
rect 11760 12724 11772 12758
rect 11760 12718 11818 12724
rect 11760 -170 11818 -164
rect 11760 -204 11772 -170
rect 11760 -210 11818 -204
rect 11578 -289 11631 -253
rect 11947 -306 12017 52681
rect 12129 52613 12187 52619
rect 12129 52579 12141 52613
rect 12129 52573 12187 52579
rect 12129 46103 12187 46109
rect 12129 46069 12141 46103
rect 12129 46063 12187 46069
rect 12129 45995 12187 46001
rect 12129 45961 12141 45995
rect 12129 45955 12187 45961
rect 12129 39485 12187 39491
rect 12129 39451 12141 39485
rect 12129 39445 12187 39451
rect 12129 39377 12187 39383
rect 12129 39343 12141 39377
rect 12129 39337 12187 39343
rect 12129 32867 12187 32873
rect 12129 32833 12141 32867
rect 12129 32827 12187 32833
rect 12129 32759 12187 32765
rect 12129 32725 12141 32759
rect 12129 32719 12187 32725
rect 12129 26249 12187 26255
rect 12129 26215 12141 26249
rect 12129 26209 12187 26215
rect 12129 26141 12187 26147
rect 12129 26107 12141 26141
rect 12129 26101 12187 26107
rect 12129 19631 12187 19637
rect 12129 19597 12141 19631
rect 12129 19591 12187 19597
rect 12129 19523 12187 19529
rect 12129 19489 12141 19523
rect 12129 19483 12187 19489
rect 12129 13013 12187 13019
rect 12129 12979 12141 13013
rect 12129 12973 12187 12979
rect 12129 12905 12187 12911
rect 12129 12871 12141 12905
rect 12129 12865 12187 12871
rect 12129 6395 12187 6401
rect 12129 6361 12141 6395
rect 12129 6355 12187 6361
rect 12129 6287 12187 6293
rect 12129 6253 12141 6287
rect 12129 6247 12187 6253
rect 12129 -223 12187 -217
rect 12129 -257 12141 -223
rect 12129 -263 12187 -257
rect 11947 -342 12000 -306
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
rect 0 -1600 200 -1400
rect 0 -2000 200 -1800
rect 0 -2400 200 -2200
rect 0 -2800 200 -2600
rect 0 -3200 200 -3000
rect 0 -3600 200 -3400
rect 0 -4000 200 -3800
rect 0 -4400 200 -4200
rect 0 -4800 200 -4600
rect 0 -5200 200 -5000
rect 0 -5600 200 -5400
rect 0 -6000 200 -5800
rect 0 -6400 200 -6200
rect 0 -6800 200 -6600
rect 0 -7200 200 -7000
rect 0 -7600 200 -7400
rect 0 -8000 200 -7800
rect 0 -8400 200 -8200
rect 0 -8800 200 -8600
use sky130_fd_sc_hd__or2_1  x1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 13052 0 1 -496
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  x2
timestamp 1701704242
transform 1 0 13550 0 1 -544
box -38 -48 498 592
use sky130_fd_sc_hd__inv_1  x7 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 12738 0 1 -448
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  x11
timestamp 1701704242
transform 1 0 0 0 1 600
box -38 -48 498 592
use sky130_fd_sc_hd__inv_1  x20
timestamp 1701704242
transform 1 0 498 0 1 552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_4  x21 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 812 0 1 504
box -38 -48 498 592
use sky130_fd_sc_hd__inv_16  x22 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 1310 0 1 456
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_1  x27
timestamp 1701704242
transform 1 0 2820 0 1 408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_4  x28
timestamp 1701704242
transform 1 0 3134 0 1 360
box -38 -48 498 592
use sky130_fd_sc_hd__inv_16  x29
timestamp 1701704242
transform 1 0 3632 0 1 312
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_1  x34
timestamp 1701704242
transform 1 0 5142 0 1 264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_4  x35
timestamp 1701704242
transform 1 0 5456 0 1 216
box -38 -48 498 592
use sky130_fd_sc_hd__inv_16  x36
timestamp 1701704242
transform 1 0 5954 0 1 168
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_1  x41
timestamp 1701704242
transform 1 0 7464 0 1 120
box -38 -48 314 592
use sky130_fd_sc_hd__inv_4  x42
timestamp 1701704242
transform 1 0 7778 0 1 72
box -38 -48 498 592
use sky130_fd_sc_hd__inv_16  x43
timestamp 1701704242
transform 1 0 8276 0 1 24
box -38 -48 1510 592
use sky130_fd_pr__nfet_01v8_HZDS57  XM3
timestamp 0
transform 1 0 9944 0 1 26496
box -211 -26573 211 26573
use sky130_fd_pr__pfet_01v8_VCZ8PW  XM4
timestamp 0
transform 1 0 10313 0 1 104259
box -211 -104389 211 104389
use sky130_fd_pr__nfet_01v8_HZDS57  XM5
timestamp 0
transform 1 0 10682 0 1 26390
box -211 -26573 211 26573
use sky130_fd_pr__pfet_01v8_VCZ8PW  XM6
timestamp 0
transform 1 0 11051 0 1 104153
box -211 -104389 211 104389
use sky130_fd_pr__nfet_01v8_HZDS57  XM7
timestamp 0
transform 1 0 11420 0 1 26284
box -211 -26573 211 26573
use sky130_fd_pr__pfet_01v8_VCZ8PW  XM8
timestamp 0
transform 1 0 11789 0 1 104047
box -211 -104389 211 104389
use sky130_fd_pr__nfet_01v8_HZDS57  XM9
timestamp 0
transform 1 0 12158 0 1 26178
box -211 -26573 211 26573
use sky130_fd_pr__pfet_01v8_VCZ8PW  XM10
timestamp 0
transform 1 0 12527 0 1 103941
box -211 -104389 211 104389
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 I14
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 I13
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 I12
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 I11
port 3 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 256 0 0 0 I10
port 4 nsew
flabel metal1 0 -2000 200 -1800 0 FreeSans 256 0 0 0 I9
port 5 nsew
flabel metal1 0 -2400 200 -2200 0 FreeSans 256 0 0 0 I8
port 6 nsew
flabel metal1 0 -2800 200 -2600 0 FreeSans 256 0 0 0 I7
port 7 nsew
flabel metal1 0 -3200 200 -3000 0 FreeSans 256 0 0 0 I6
port 8 nsew
flabel metal1 0 -3600 200 -3400 0 FreeSans 256 0 0 0 I5
port 9 nsew
flabel metal1 0 -4000 200 -3800 0 FreeSans 256 0 0 0 I4
port 10 nsew
flabel metal1 0 -4400 200 -4200 0 FreeSans 256 0 0 0 I3
port 11 nsew
flabel metal1 0 -4800 200 -4600 0 FreeSans 256 0 0 0 I2
port 12 nsew
flabel metal1 0 -5200 200 -5000 0 FreeSans 256 0 0 0 I1
port 13 nsew
flabel metal1 0 -5600 200 -5400 0 FreeSans 256 0 0 0 I0
port 14 nsew
flabel metal1 0 -6000 200 -5800 0 FreeSans 256 0 0 0 A4
port 15 nsew
flabel metal1 0 -6400 200 -6200 0 FreeSans 256 0 0 0 A3
port 16 nsew
flabel metal1 0 -6800 200 -6600 0 FreeSans 256 0 0 0 A2
port 17 nsew
flabel metal1 0 -7200 200 -7000 0 FreeSans 256 0 0 0 A1
port 18 nsew
flabel metal1 0 -7600 200 -7400 0 FreeSans 256 0 0 0 VDD
port 19 nsew
flabel metal1 0 -8000 200 -7800 0 FreeSans 256 0 0 0 GND
port 20 nsew
flabel metal1 0 -8400 200 -8200 0 FreeSans 256 0 0 0 I15
port 21 nsew
flabel metal1 0 -8800 200 -8600 0 FreeSans 256 0 0 0 EI
port 22 nsew
<< end >>
