magic
tech sky130A
magscale 1 2
timestamp 1714790421
<< pwell >>
rect -739 -6154 739 6154
<< psubdiff >>
rect -703 6084 -607 6118
rect 607 6084 703 6118
rect -703 6022 -669 6084
rect 669 6022 703 6084
rect -703 -6084 -669 -6022
rect 669 -6084 703 -6022
rect -703 -6118 -607 -6084
rect 607 -6118 703 -6084
<< psubdiffcont >>
rect -607 6084 607 6118
rect -703 -6022 -669 6022
rect 669 -6022 703 6022
rect -607 -6118 607 -6084
<< xpolycontact >>
rect -573 5556 573 5988
rect -573 4582 573 5014
rect -573 4046 573 4478
rect -573 3072 573 3504
rect -573 2536 573 2968
rect -573 1562 573 1994
rect -573 1026 573 1458
rect -573 52 573 484
rect -573 -484 573 -52
rect -573 -1458 573 -1026
rect -573 -1994 573 -1562
rect -573 -2968 573 -2536
rect -573 -3504 573 -3072
rect -573 -4478 573 -4046
rect -573 -5014 573 -4582
rect -573 -5988 573 -5556
<< xpolyres >>
rect -573 5014 573 5556
rect -573 3504 573 4046
rect -573 1994 573 2536
rect -573 484 573 1026
rect -573 -1026 573 -484
rect -573 -2536 573 -1994
rect -573 -4046 573 -3504
rect -573 -5556 573 -5014
<< locali >>
rect -703 6084 -607 6118
rect 607 6084 703 6118
rect -703 6022 -669 6084
rect 669 6022 703 6084
rect -703 -6084 -669 -6022
rect 669 -6084 703 -6022
rect -703 -6118 -607 -6084
rect 607 -6118 703 -6084
<< viali >>
rect -557 5573 557 5970
rect -557 4600 557 4997
rect -557 4063 557 4460
rect -557 3090 557 3487
rect -557 2553 557 2950
rect -557 1580 557 1977
rect -557 1043 557 1440
rect -557 70 557 467
rect -557 -467 557 -70
rect -557 -1440 557 -1043
rect -557 -1977 557 -1580
rect -557 -2950 557 -2553
rect -557 -3487 557 -3090
rect -557 -4460 557 -4063
rect -557 -4997 557 -4600
rect -557 -5970 557 -5573
<< metal1 >>
rect -569 5970 569 5976
rect -569 5573 -557 5970
rect 557 5573 569 5970
rect -569 5567 569 5573
rect -569 4997 569 5003
rect -569 4600 -557 4997
rect 557 4600 569 4997
rect -569 4594 569 4600
rect -569 4460 569 4466
rect -569 4063 -557 4460
rect 557 4063 569 4460
rect -569 4057 569 4063
rect -569 3487 569 3493
rect -569 3090 -557 3487
rect 557 3090 569 3487
rect -569 3084 569 3090
rect -569 2950 569 2956
rect -569 2553 -557 2950
rect 557 2553 569 2950
rect -569 2547 569 2553
rect -569 1977 569 1983
rect -569 1580 -557 1977
rect 557 1580 569 1977
rect -569 1574 569 1580
rect -569 1440 569 1446
rect -569 1043 -557 1440
rect 557 1043 569 1440
rect -569 1037 569 1043
rect -569 467 569 473
rect -569 70 -557 467
rect 557 70 569 467
rect -569 64 569 70
rect -569 -70 569 -64
rect -569 -467 -557 -70
rect 557 -467 569 -70
rect -569 -473 569 -467
rect -569 -1043 569 -1037
rect -569 -1440 -557 -1043
rect 557 -1440 569 -1043
rect -569 -1446 569 -1440
rect -569 -1580 569 -1574
rect -569 -1977 -557 -1580
rect 557 -1977 569 -1580
rect -569 -1983 569 -1977
rect -569 -2553 569 -2547
rect -569 -2950 -557 -2553
rect 557 -2950 569 -2553
rect -569 -2956 569 -2950
rect -569 -3090 569 -3084
rect -569 -3487 -557 -3090
rect 557 -3487 569 -3090
rect -569 -3493 569 -3487
rect -569 -4063 569 -4057
rect -569 -4460 -557 -4063
rect 557 -4460 569 -4063
rect -569 -4466 569 -4460
rect -569 -4600 569 -4594
rect -569 -4997 -557 -4600
rect 557 -4997 569 -4600
rect -569 -5003 569 -4997
rect -569 -5573 569 -5567
rect -569 -5970 -557 -5573
rect 557 -5970 569 -5573
rect -569 -5976 569 -5970
<< properties >>
string FIXED_BBOX -686 -6101 686 6101
string gencell sky130_fd_pr__res_xhigh_po_5p73
string library sky130
string parameters w 5.730 l 2.865 m 8 nx 1 wmin 5.730 lmin 0.50 rho 2000 val 1.065k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 5.730 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
