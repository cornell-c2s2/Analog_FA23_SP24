magic
tech sky130A
magscale 1 2
timestamp 1717026683
<< pwell >>
rect 165900 -47800 178524 -41354
rect 196300 -42700 196900 -41400
rect 197496 -47798 208300 -47600
rect 197496 -48100 208300 -48098
<< viali >>
rect 140696 -24498 140796 -24398
rect 141796 -24498 141896 -24398
rect 142896 -24498 142996 -24398
rect 143996 -24498 144096 -24398
rect 145096 -24498 145196 -24398
rect 146196 -24498 146296 -24398
rect 172296 -24498 172396 -24398
rect 173396 -24498 173496 -24398
rect 174496 -24498 174596 -24398
rect 175596 -24498 175696 -24398
rect 176696 -24498 176796 -24398
rect 177796 -24498 177896 -24398
rect 167196 -47798 167296 -47698
rect 168196 -47798 168296 -47698
rect 169296 -47798 169396 -47698
rect 170396 -47798 170496 -47698
rect 171496 -47798 171596 -47698
rect 172596 -47798 172696 -47698
rect 173696 -47798 173796 -47698
rect 174796 -47798 174896 -47698
rect 175896 -47798 175996 -47698
rect 176996 -47798 177096 -47698
rect 197596 -47798 197696 -47698
rect 198596 -47798 198696 -47698
rect 199696 -47798 199796 -47698
rect 200796 -47798 200896 -47698
rect 201896 -47798 201996 -47698
rect 202996 -47798 203096 -47698
rect 204096 -47798 204196 -47698
rect 205196 -47798 205296 -47698
rect 206296 -47798 206396 -47698
rect 207396 -47798 207496 -47698
<< metal1 >>
rect 140600 -12500 143000 -12000
rect 143200 -12500 145500 -12000
rect 145790 -12200 145800 -12100
rect 145900 -12200 145910 -12100
rect 145990 -12200 146000 -12100
rect 146100 -12200 146110 -12100
rect 146190 -12200 146200 -12100
rect 146300 -12200 146310 -12100
rect 146390 -12200 146400 -12100
rect 146500 -12200 146510 -12100
rect 146590 -12200 146600 -12100
rect 146700 -12200 146710 -12100
rect 145790 -12400 145800 -12300
rect 145900 -12400 145910 -12300
rect 145990 -12400 146000 -12300
rect 146100 -12400 146110 -12300
rect 146190 -12400 146200 -12300
rect 146300 -12400 146310 -12300
rect 146390 -12400 146400 -12300
rect 146500 -12400 146510 -12300
rect 146590 -12400 146600 -12300
rect 146700 -12400 146710 -12300
rect 172100 -12500 174500 -12000
rect 174700 -12500 177000 -12000
rect 177190 -12200 177200 -12100
rect 177300 -12200 177310 -12100
rect 177390 -12200 177400 -12100
rect 177500 -12200 177510 -12100
rect 177590 -12200 177600 -12100
rect 177700 -12200 177710 -12100
rect 177790 -12200 177800 -12100
rect 177900 -12200 177910 -12100
rect 177990 -12200 178000 -12100
rect 178100 -12200 178110 -12100
rect 177390 -12400 177400 -12300
rect 177500 -12400 177510 -12300
rect 177590 -12400 177600 -12300
rect 177700 -12400 177710 -12300
rect 177790 -12400 177800 -12300
rect 177900 -12400 177910 -12300
rect 177990 -12400 178000 -12300
rect 178100 -12400 178110 -12300
rect 140684 -23898 140908 -23892
rect 140684 -24098 140696 -23898
rect 140896 -24098 140908 -23898
rect 140684 -24104 140908 -24098
rect 141084 -23898 141308 -23892
rect 141084 -24098 141096 -23898
rect 141296 -24098 141308 -23898
rect 141084 -24104 141308 -24098
rect 141484 -23898 141708 -23892
rect 141484 -24098 141496 -23898
rect 141696 -24098 141708 -23898
rect 141484 -24104 141708 -24098
rect 141900 -24300 144300 -23900
rect 144400 -24300 146800 -23900
rect 172190 -24100 172200 -24000
rect 172300 -24100 172310 -24000
rect 172390 -24100 172400 -24000
rect 172500 -24100 172510 -24000
rect 172590 -24100 172600 -24000
rect 172700 -24100 172710 -24000
rect 172790 -24100 172800 -24000
rect 172900 -24100 172910 -24000
rect 172990 -24100 173000 -24000
rect 173100 -24200 173110 -24100
rect 172190 -24300 172200 -24200
rect 172300 -24300 172310 -24200
rect 172390 -24300 172400 -24200
rect 172500 -24300 172510 -24200
rect 172590 -24300 172600 -24200
rect 172700 -24300 172710 -24200
rect 172790 -24300 172800 -24200
rect 172900 -24300 172910 -24200
rect 172990 -24300 173000 -24200
rect 173400 -24300 175800 -23900
rect 175900 -24300 178300 -23900
rect 140684 -24398 140808 -24392
rect 141784 -24398 141908 -24392
rect 142884 -24398 143008 -24392
rect 143984 -24398 144108 -24392
rect 145084 -24398 145208 -24392
rect 146184 -24398 146308 -24392
rect 172284 -24398 172408 -24392
rect 173384 -24398 173508 -24392
rect 174484 -24398 174608 -24392
rect 175584 -24398 175708 -24392
rect 176684 -24398 176808 -24392
rect 177784 -24398 177908 -24392
rect 140496 -24498 140696 -24398
rect 140796 -24498 141796 -24398
rect 141896 -24498 142896 -24398
rect 142996 -24498 143996 -24398
rect 144096 -24498 145096 -24398
rect 145196 -24498 146196 -24398
rect 146296 -24498 148796 -24398
rect 172096 -24498 172296 -24398
rect 172396 -24498 173396 -24398
rect 173496 -24498 174496 -24398
rect 174596 -24498 175596 -24398
rect 175696 -24498 176696 -24398
rect 176796 -24498 177796 -24398
rect 177896 -24498 180496 -24398
rect 140496 -24598 148496 -24498
rect 148596 -24598 148696 -24498
rect 148796 -24598 148806 -24498
rect 172096 -24598 180496 -24498
rect 180696 -24598 180706 -24398
rect 166090 -41700 166100 -41600
rect 166200 -41700 166210 -41600
rect 166290 -41700 166300 -41600
rect 166400 -41700 166410 -41600
rect 166090 -41900 166100 -41800
rect 166200 -41900 166210 -41800
rect 166290 -41900 166300 -41800
rect 166400 -41900 166410 -41800
rect 166090 -42100 166100 -42000
rect 166200 -42100 166210 -42000
rect 166290 -42100 166300 -42000
rect 166400 -42100 166410 -42000
rect 166090 -42300 166100 -42200
rect 166200 -42300 166210 -42200
rect 166290 -42300 166300 -42200
rect 166400 -42300 166410 -42200
rect 166090 -42500 166100 -42400
rect 166200 -42500 166210 -42400
rect 166290 -42500 166300 -42400
rect 166400 -42500 166410 -42400
rect 166100 -45100 166500 -42800
rect 177900 -43900 178400 -41500
rect 166100 -47600 166500 -45300
rect 177900 -46400 178400 -44000
rect 183686 -45198 183696 -45098
rect 183796 -45198 183806 -45098
rect 183886 -45198 183896 -45098
rect 183996 -45198 184006 -45098
rect 196424 -45100 196924 -42750
rect 208324 -43900 208724 -41500
rect 177990 -46700 178000 -46600
rect 178100 -46700 178110 -46600
rect 178190 -46700 178200 -46600
rect 178300 -46700 178310 -46600
rect 177990 -46900 178000 -46800
rect 178100 -46900 178110 -46800
rect 178190 -46900 178200 -46800
rect 178300 -46900 178310 -46800
rect 171990 -47300 172000 -47000
rect 172300 -47300 172310 -47000
rect 177990 -47100 178000 -47000
rect 178100 -47100 178110 -47000
rect 178190 -47100 178200 -47000
rect 178300 -47100 178310 -47000
rect 177990 -47300 178000 -47200
rect 178100 -47300 178110 -47200
rect 178190 -47300 178200 -47200
rect 178300 -47300 178310 -47200
rect 167184 -47698 167308 -47692
rect 168184 -47698 168308 -47692
rect 169284 -47698 169408 -47692
rect 170384 -47698 170508 -47692
rect 171484 -47698 171608 -47692
rect 172000 -47698 172300 -47300
rect 177990 -47500 178000 -47400
rect 178100 -47500 178110 -47400
rect 178190 -47500 178200 -47400
rect 178300 -47500 178310 -47400
rect 196424 -47600 196924 -45300
rect 208324 -46400 208724 -44000
rect 214770 -45198 214796 -45098
rect 214896 -45198 214996 -45098
rect 215096 -45118 215196 -45098
rect 215096 -45198 215646 -45118
rect 214770 -45218 215646 -45198
rect 208390 -46700 208400 -46600
rect 208500 -46700 208510 -46600
rect 208590 -46700 208600 -46600
rect 208700 -46700 208710 -46600
rect 208390 -46900 208400 -46800
rect 208500 -46900 208510 -46800
rect 208590 -46900 208600 -46800
rect 208700 -46900 208710 -46800
rect 202390 -47300 202400 -47000
rect 202700 -47300 202710 -47000
rect 208390 -47100 208400 -47000
rect 208500 -47100 208510 -47000
rect 208590 -47100 208600 -47000
rect 208700 -47100 208710 -47000
rect 208390 -47300 208400 -47200
rect 208500 -47300 208510 -47200
rect 208590 -47300 208600 -47200
rect 208700 -47300 208710 -47200
rect 172584 -47698 172708 -47692
rect 173684 -47698 173808 -47692
rect 174784 -47698 174908 -47692
rect 175884 -47698 176008 -47692
rect 176984 -47698 177108 -47692
rect 197584 -47698 197708 -47692
rect 198584 -47698 198708 -47692
rect 199684 -47698 199808 -47692
rect 200784 -47698 200908 -47692
rect 201884 -47698 202008 -47692
rect 202400 -47698 202700 -47300
rect 208390 -47500 208400 -47400
rect 208500 -47500 208510 -47400
rect 208590 -47500 208600 -47400
rect 208700 -47500 208710 -47400
rect 202984 -47698 203108 -47692
rect 204084 -47698 204208 -47692
rect 205184 -47698 205308 -47692
rect 206284 -47698 206408 -47692
rect 207384 -47698 207508 -47692
rect 166500 -47798 167196 -47698
rect 167296 -47798 168196 -47698
rect 168296 -47798 169296 -47698
rect 169396 -47798 170396 -47698
rect 170496 -47798 171496 -47698
rect 171596 -47798 172596 -47698
rect 172696 -47798 173696 -47698
rect 173796 -47798 174796 -47698
rect 174896 -47798 175896 -47698
rect 175996 -47798 176996 -47698
rect 177096 -47798 178300 -47698
rect 196900 -47700 197596 -47698
rect 166500 -47898 178300 -47798
rect 196400 -47798 197596 -47700
rect 197696 -47798 198596 -47698
rect 198696 -47798 199696 -47698
rect 199796 -47798 200796 -47698
rect 200896 -47798 201896 -47698
rect 201996 -47798 202996 -47698
rect 203096 -47798 204096 -47698
rect 204196 -47798 205196 -47698
rect 205296 -47798 206296 -47698
rect 206396 -47798 207396 -47698
rect 207496 -47798 208700 -47698
rect 196400 -47898 208700 -47798
rect 172000 -47900 172300 -47898
rect 202400 -47900 202700 -47898
rect 185486 -48098 185496 -47998
rect 185596 -48098 185606 -47998
rect 185786 -48098 185796 -47998
rect 185896 -48098 185906 -47998
rect 217086 -48098 217096 -47998
rect 217196 -48098 217206 -47998
rect 217286 -48098 217296 -47998
rect 217396 -48098 217406 -47998
<< via1 >>
rect 145800 -12200 145900 -12100
rect 146000 -12200 146100 -12100
rect 146200 -12200 146300 -12100
rect 146400 -12200 146500 -12100
rect 146600 -12200 146700 -12100
rect 145800 -12400 145900 -12300
rect 146000 -12400 146100 -12300
rect 146200 -12400 146300 -12300
rect 146400 -12400 146500 -12300
rect 146600 -12400 146700 -12300
rect 177200 -12200 177300 -12100
rect 177400 -12200 177500 -12100
rect 177600 -12200 177700 -12100
rect 177800 -12200 177900 -12100
rect 178000 -12200 178100 -12100
rect 177200 -12400 177300 -12300
rect 177400 -12400 177500 -12300
rect 177600 -12400 177700 -12300
rect 177800 -12400 177900 -12300
rect 178000 -12400 178100 -12300
rect 140696 -24098 140896 -23898
rect 141096 -24098 141296 -23898
rect 141496 -24098 141696 -23898
rect 172200 -24100 172300 -24000
rect 172400 -24100 172500 -24000
rect 172600 -24100 172700 -24000
rect 172800 -24100 172900 -24000
rect 173000 -24100 173100 -24000
rect 172200 -24300 172300 -24200
rect 172400 -24300 172500 -24200
rect 172600 -24300 172700 -24200
rect 172800 -24300 172900 -24200
rect 173000 -24300 173100 -24200
rect 148496 -24598 148596 -24498
rect 148696 -24598 148796 -24498
rect 180496 -24598 180696 -24398
rect 166100 -41700 166200 -41600
rect 166300 -41700 166400 -41600
rect 166100 -41900 166200 -41800
rect 166300 -41900 166400 -41800
rect 166100 -42100 166200 -42000
rect 166300 -42100 166400 -42000
rect 166100 -42300 166200 -42200
rect 166300 -42300 166400 -42200
rect 166100 -42500 166200 -42400
rect 166300 -42500 166400 -42400
rect 196500 -41700 196600 -41600
rect 196700 -41700 196800 -41600
rect 196500 -41900 196600 -41800
rect 196700 -41900 196800 -41800
rect 196500 -42100 196600 -42000
rect 196700 -42100 196800 -42000
rect 196500 -42300 196600 -42200
rect 196700 -42300 196800 -42200
rect 196500 -42500 196600 -42400
rect 196700 -42500 196800 -42400
rect 183696 -45198 183796 -45098
rect 183896 -45198 183996 -45098
rect 178000 -46700 178100 -46600
rect 178200 -46700 178300 -46600
rect 178000 -46900 178100 -46800
rect 178200 -46900 178300 -46800
rect 172000 -47300 172300 -47000
rect 178000 -47100 178100 -47000
rect 178200 -47100 178300 -47000
rect 178000 -47300 178100 -47200
rect 178200 -47300 178300 -47200
rect 178000 -47500 178100 -47400
rect 178200 -47500 178300 -47400
rect 214796 -45198 214896 -45098
rect 214996 -45198 215096 -45098
rect 208400 -46700 208500 -46600
rect 208600 -46700 208700 -46600
rect 208400 -46900 208500 -46800
rect 208600 -46900 208700 -46800
rect 202400 -47300 202700 -47000
rect 208400 -47100 208500 -47000
rect 208600 -47100 208700 -47000
rect 208400 -47300 208500 -47200
rect 208600 -47300 208700 -47200
rect 208400 -47500 208500 -47400
rect 208600 -47500 208700 -47400
rect 185496 -48098 185596 -47998
rect 185796 -48098 185896 -47998
rect 217096 -48098 217196 -47998
rect 217296 -48098 217396 -47998
<< metal2 >>
rect 145700 -12100 146900 -12000
rect 145700 -12200 145800 -12100
rect 145900 -12200 146000 -12100
rect 146100 -12200 146200 -12100
rect 146300 -12200 146400 -12100
rect 146500 -12200 146600 -12100
rect 146700 -12200 146900 -12100
rect 145700 -12300 146900 -12200
rect 145700 -12400 145800 -12300
rect 145900 -12400 146000 -12300
rect 146100 -12400 146200 -12300
rect 146300 -12400 146400 -12300
rect 146500 -12400 146600 -12300
rect 146700 -12400 146900 -12300
rect 145700 -12500 146900 -12400
rect 177200 -12100 177300 -12090
rect 177400 -12100 177500 -12090
rect 177300 -12200 177400 -12102
rect 177600 -12100 177700 -12090
rect 177500 -12200 177600 -12102
rect 177800 -12100 177900 -12090
rect 177700 -12200 177800 -12102
rect 178000 -12100 178100 -12090
rect 177900 -12200 178000 -12102
rect 178100 -12200 178200 -12102
rect 177200 -12300 178200 -12200
rect 177300 -12400 177400 -12300
rect 177500 -12400 177600 -12300
rect 177700 -12400 177800 -12300
rect 177900 -12400 178000 -12300
rect 178100 -12400 178200 -12300
rect 145896 -16298 146896 -12500
rect 145896 -16498 146296 -16298
rect 146496 -16498 146696 -16298
rect 145896 -16698 146896 -16498
rect 145896 -16898 146296 -16698
rect 146496 -16898 146696 -16698
rect 140696 -23898 140896 -23888
rect 140696 -24108 140896 -24098
rect 141096 -23898 141296 -23888
rect 141096 -24108 141296 -24098
rect 141496 -23898 141696 -23888
rect 141496 -24108 141696 -24098
rect 145896 -40498 146896 -16898
rect 177200 -16298 178200 -12400
rect 177200 -16498 177396 -16298
rect 177596 -16498 177796 -16298
rect 177996 -16498 178200 -16298
rect 177200 -16698 178200 -16498
rect 177200 -16898 177396 -16698
rect 177596 -16898 177796 -16698
rect 177996 -16898 178200 -16698
rect 177200 -17100 178200 -16898
rect 178700 -16298 179696 -15998
rect 178700 -16498 178896 -16298
rect 179096 -16498 179296 -16298
rect 179496 -16498 179696 -16298
rect 178700 -16698 179696 -16498
rect 178700 -16898 178896 -16698
rect 179096 -16898 179296 -16698
rect 179496 -16898 179696 -16698
rect 172096 -17698 173096 -17398
rect 172096 -17898 172296 -17698
rect 172496 -17898 172696 -17698
rect 172896 -17898 173096 -17698
rect 172096 -18098 173096 -17898
rect 178700 -17900 179696 -16898
rect 172096 -18298 172296 -18098
rect 172496 -18298 172696 -18098
rect 172896 -18298 173096 -18098
rect 172096 -23900 173096 -18298
rect 172096 -24000 173200 -23900
rect 172096 -24100 172200 -24000
rect 172300 -24100 172400 -24000
rect 172500 -24100 172600 -24000
rect 172700 -24100 172800 -24000
rect 172900 -24100 173000 -24000
rect 173100 -24100 173200 -24000
rect 172096 -24200 173200 -24100
rect 172096 -24300 172200 -24200
rect 172300 -24300 172400 -24200
rect 172500 -24300 172600 -24200
rect 172700 -24300 172800 -24200
rect 172900 -24300 173000 -24200
rect 173100 -24300 173200 -24200
rect 172096 -24400 173200 -24300
rect 148496 -24498 148596 -24488
rect 148496 -24608 148596 -24598
rect 148696 -24498 148796 -24488
rect 148696 -24608 148796 -24598
rect 172096 -25898 173096 -24400
rect 172096 -26098 172296 -25898
rect 172496 -26098 172696 -25898
rect 172896 -26098 173096 -25898
rect 172096 -26198 173096 -26098
rect 145896 -40698 146096 -40498
rect 146296 -40698 146496 -40498
rect 146696 -40698 146896 -40498
rect 145896 -40798 146896 -40698
rect 166000 -40300 166400 -40291
rect 166000 -41500 166400 -40700
rect 178696 -40498 179696 -17900
rect 197496 -17698 198496 -17498
rect 197496 -17898 197696 -17698
rect 197896 -17898 198096 -17698
rect 198296 -17898 198496 -17698
rect 197496 -18098 198496 -17898
rect 197496 -18298 197696 -18098
rect 197896 -18298 198096 -18098
rect 198296 -18298 198496 -18098
rect 180496 -24398 180696 -24388
rect 180496 -24608 180696 -24598
rect 197496 -25898 198496 -18298
rect 197496 -26098 197696 -25898
rect 197896 -26098 198096 -25898
rect 198296 -26098 198496 -25898
rect 197696 -26108 197896 -26098
rect 198096 -26108 198296 -26098
rect 235496 -26898 236096 -26698
rect 235696 -27098 235896 -26898
rect 196405 -40300 196795 -40294
rect 178696 -40698 178896 -40498
rect 179096 -40698 179296 -40498
rect 179496 -40698 179696 -40498
rect 178696 -40898 179696 -40698
rect 196400 -40303 196800 -40300
rect 196400 -40693 196405 -40303
rect 196795 -40693 196800 -40303
rect 196400 -41500 196800 -40693
rect 166000 -41600 166500 -41500
rect 166000 -41700 166100 -41600
rect 166200 -41700 166300 -41600
rect 166400 -41700 166500 -41600
rect 166000 -41800 166500 -41700
rect 166000 -41900 166100 -41800
rect 166200 -41900 166300 -41800
rect 166400 -41900 166500 -41800
rect 166000 -42000 166500 -41900
rect 166000 -42100 166100 -42000
rect 166200 -42100 166300 -42000
rect 166400 -42100 166500 -42000
rect 166000 -42200 166500 -42100
rect 166000 -42300 166100 -42200
rect 166200 -42300 166300 -42200
rect 166400 -42300 166500 -42200
rect 166000 -42400 166500 -42300
rect 166000 -42500 166100 -42400
rect 166200 -42500 166300 -42400
rect 166400 -42500 166500 -42400
rect 166000 -42600 166500 -42500
rect 196400 -41600 196900 -41500
rect 196400 -41700 196500 -41600
rect 196600 -41700 196700 -41600
rect 196800 -41700 196900 -41600
rect 196400 -41800 196900 -41700
rect 196400 -41900 196500 -41800
rect 196600 -41900 196700 -41800
rect 196800 -41900 196900 -41800
rect 196400 -42000 196900 -41900
rect 196400 -42100 196500 -42000
rect 196600 -42100 196700 -42000
rect 196800 -42100 196900 -42000
rect 196400 -42200 196900 -42100
rect 196400 -42300 196500 -42200
rect 196600 -42300 196700 -42200
rect 196800 -42300 196900 -42200
rect 196400 -42400 196900 -42300
rect 196400 -42500 196500 -42400
rect 196600 -42500 196700 -42400
rect 196800 -42500 196900 -42400
rect 196400 -42600 196900 -42500
rect 186696 -44098 186896 -44088
rect 186496 -44298 186696 -44098
rect 186496 -44498 186896 -44298
rect 186496 -44698 186696 -44498
rect 186496 -44898 186896 -44698
rect 183696 -45098 183796 -45088
rect 183696 -45208 183796 -45198
rect 183896 -45098 183996 -45088
rect 183896 -45208 183996 -45198
rect 186496 -45098 186696 -44898
rect 235496 -44298 236096 -27098
rect 235696 -44498 235896 -44298
rect 235496 -44698 236096 -44498
rect 235696 -44898 235896 -44698
rect 186496 -45698 186896 -45098
rect 214796 -45098 215196 -44998
rect 214896 -45198 214996 -45098
rect 215096 -45198 215196 -45098
rect 214796 -45208 215096 -45198
rect 214796 -45398 214996 -45208
rect 214796 -45608 214996 -45598
rect 178000 -46300 178200 -46290
rect 220496 -46298 220696 -46288
rect 177900 -46500 178000 -46300
rect 178200 -46500 178400 -46300
rect 177900 -46600 178400 -46500
rect 177900 -46900 178000 -46600
rect 178300 -46700 178400 -46600
rect 178200 -46800 178400 -46700
rect 178100 -46900 178200 -46800
rect 178300 -46900 178400 -46800
rect 172000 -47000 172300 -46990
rect 172000 -47310 172300 -47300
rect 177900 -47000 178400 -46900
rect 208300 -46600 208800 -46500
rect 220496 -46508 220696 -46498
rect 235496 -46498 236096 -44898
rect 177900 -47100 178000 -47000
rect 178100 -47100 178200 -47000
rect 178300 -47100 178400 -47000
rect 177900 -47200 178400 -47100
rect 177900 -47300 178000 -47200
rect 178100 -47300 178200 -47200
rect 178300 -47300 178400 -47200
rect 177900 -47400 178400 -47300
rect 202400 -47000 202700 -46990
rect 202400 -47310 202700 -47300
rect 208300 -47100 208400 -46600
rect 208700 -46700 208800 -46600
rect 208600 -46800 208800 -46700
rect 208500 -46900 208600 -46800
rect 208700 -46900 208800 -46800
rect 208600 -47000 208800 -46900
rect 220496 -46698 220696 -46688
rect 235696 -46698 235896 -46498
rect 235496 -46798 236096 -46698
rect 220496 -46908 220696 -46898
rect 208700 -47100 208800 -47000
rect 208300 -47200 208800 -47100
rect 208300 -47300 208400 -47200
rect 208500 -47300 208600 -47200
rect 208700 -47300 208800 -47200
rect 177900 -47500 178000 -47400
rect 178100 -47500 178200 -47400
rect 178300 -47500 178400 -47400
rect 208300 -47400 208800 -47300
rect 187096 -47498 187296 -47488
rect 177900 -47600 178400 -47500
rect 180896 -51098 181296 -47498
rect 186896 -47698 187096 -47498
rect 208300 -47500 208400 -47400
rect 208500 -47500 208600 -47400
rect 208700 -47500 208800 -47400
rect 208300 -47600 208800 -47500
rect 185496 -47998 185596 -47988
rect 185496 -48108 185596 -48098
rect 185796 -47998 185896 -47988
rect 185796 -48108 185896 -48098
rect 186896 -48698 187296 -47698
rect 186896 -48898 187096 -48698
rect 187096 -48908 187296 -48898
rect 180896 -51298 181096 -51098
rect 214896 -51098 215296 -47498
rect 217096 -47998 217196 -47988
rect 217096 -48108 217196 -48098
rect 217296 -47998 217396 -47988
rect 217296 -48108 217396 -48098
rect 219496 -48698 219896 -47698
rect 219496 -48898 219696 -48698
rect 219696 -48908 219896 -48898
rect 214896 -51298 215096 -51098
rect 181096 -51308 181296 -51298
rect 215096 -51308 215296 -51298
<< via2 >>
rect 146296 -16498 146496 -16298
rect 146696 -16498 146896 -16298
rect 146296 -16898 146496 -16698
rect 146696 -16898 146896 -16698
rect 140696 -24098 140896 -23898
rect 141096 -24098 141296 -23898
rect 141496 -24098 141696 -23898
rect 177396 -16498 177596 -16298
rect 177796 -16498 177996 -16298
rect 177396 -16898 177596 -16698
rect 177796 -16898 177996 -16698
rect 178896 -16498 179096 -16298
rect 179296 -16498 179496 -16298
rect 178896 -16898 179096 -16698
rect 179296 -16898 179496 -16698
rect 172296 -17898 172496 -17698
rect 172696 -17898 172896 -17698
rect 172296 -18298 172496 -18098
rect 172696 -18298 172896 -18098
rect 148496 -24598 148596 -24498
rect 148696 -24598 148796 -24498
rect 172296 -26098 172496 -25898
rect 172696 -26098 172896 -25898
rect 146096 -40698 146296 -40498
rect 146496 -40698 146696 -40498
rect 166000 -40700 166400 -40300
rect 197696 -17898 197896 -17698
rect 198096 -17898 198296 -17698
rect 197696 -18298 197896 -18098
rect 198096 -18298 198296 -18098
rect 180496 -24598 180696 -24398
rect 197696 -26098 197896 -25898
rect 198096 -26098 198296 -25898
rect 235496 -27098 235696 -26898
rect 235896 -27098 236096 -26898
rect 178896 -40698 179096 -40498
rect 179296 -40698 179496 -40498
rect 196405 -40693 196795 -40303
rect 186696 -44298 186896 -44098
rect 186696 -44698 186896 -44498
rect 183696 -45198 183796 -45098
rect 183896 -45198 183996 -45098
rect 186696 -45098 186896 -44898
rect 235496 -44498 235696 -44298
rect 235896 -44498 236096 -44298
rect 235496 -44898 235696 -44698
rect 235896 -44898 236096 -44698
rect 214796 -45598 214996 -45398
rect 178000 -46500 178200 -46300
rect 220496 -46498 220696 -46298
rect 178000 -46700 178100 -46600
rect 178100 -46700 178200 -46600
rect 178000 -46800 178200 -46700
rect 172000 -47300 172300 -47000
rect 202400 -47300 202700 -47000
rect 208400 -46700 208500 -46600
rect 208500 -46700 208600 -46600
rect 208400 -46800 208600 -46700
rect 208400 -47000 208600 -46900
rect 220496 -46898 220696 -46698
rect 235496 -46698 235696 -46498
rect 235896 -46698 236096 -46498
rect 208400 -47100 208500 -47000
rect 208500 -47100 208600 -47000
rect 187096 -47698 187296 -47498
rect 185496 -48098 185596 -47998
rect 185796 -48098 185896 -47998
rect 187096 -48898 187296 -48698
rect 181096 -51298 181296 -51098
rect 217096 -48098 217196 -47998
rect 217296 -48098 217396 -47998
rect 219696 -48898 219896 -48698
rect 215096 -51298 215296 -51098
<< metal3 >>
rect 170086 -15098 170096 -14698
rect 170496 -15098 170506 -14698
rect 170686 -15098 170696 -14698
rect 171096 -15098 171106 -14698
rect 201686 -15098 201696 -14698
rect 202096 -15098 202106 -14698
rect 202286 -15098 202296 -14698
rect 202696 -15098 202706 -14698
rect 227286 -15098 227296 -14698
rect 227696 -15098 227706 -14698
rect 227886 -15098 227896 -14698
rect 228296 -15098 228306 -14698
rect 145686 -16503 145906 -16293
rect 145996 -16298 146096 -16098
rect 146196 -16298 148996 -16098
rect 178700 -16100 179696 -16098
rect 145996 -16498 146296 -16298
rect 146496 -16498 146696 -16298
rect 146896 -16498 148996 -16298
rect 145686 -16903 145906 -16693
rect 145996 -16698 148996 -16498
rect 145996 -16898 146296 -16698
rect 146496 -16898 146696 -16698
rect 146896 -16898 148996 -16698
rect 145996 -17098 148996 -16898
rect 177200 -16298 179696 -16100
rect 177200 -16498 177396 -16298
rect 177596 -16498 177796 -16298
rect 177996 -16498 178896 -16298
rect 179096 -16498 179296 -16298
rect 179496 -16498 179696 -16298
rect 177200 -16698 179696 -16498
rect 177200 -16898 177396 -16698
rect 177596 -16898 177796 -16698
rect 177996 -16898 178896 -16698
rect 179096 -16898 179296 -16698
rect 179496 -16898 179696 -16698
rect 177200 -17098 179696 -16898
rect 201796 -17098 207596 -16098
rect 177200 -17100 178800 -17098
rect 201796 -17498 202796 -17098
rect 159696 -17698 173596 -17498
rect 159696 -17898 172296 -17698
rect 172496 -17898 172696 -17698
rect 172896 -17898 173596 -17698
rect 159696 -18098 173596 -17898
rect 159696 -18298 172296 -18098
rect 172496 -18298 172696 -18098
rect 172896 -18298 173596 -18098
rect 159696 -18498 173596 -18298
rect 191496 -17698 202796 -17498
rect 191496 -17898 197696 -17698
rect 197896 -17898 198096 -17698
rect 198296 -17898 202796 -17698
rect 191496 -18098 202796 -17898
rect 191496 -18298 197696 -18098
rect 197896 -18298 198096 -18098
rect 198296 -18298 202796 -18098
rect 191496 -18498 202796 -18298
rect 140696 -23893 141696 -23298
rect 140686 -23898 141706 -23893
rect 140686 -24098 140696 -23898
rect 140896 -24098 141096 -23898
rect 141296 -24098 141496 -23898
rect 141696 -24098 141706 -23898
rect 140686 -24103 141706 -24098
rect 140696 -24298 141696 -24103
rect 148486 -24598 148496 -24298
rect 148796 -24598 148806 -24298
rect 148486 -24603 148606 -24598
rect 148686 -24603 148806 -24598
rect 180386 -24698 180396 -24298
rect 180796 -24698 180806 -24298
rect 167296 -26098 170496 -25698
rect 170896 -25898 174296 -25698
rect 170896 -26098 172296 -25898
rect 172496 -26098 172696 -25898
rect 172896 -26098 174296 -25898
rect 174696 -26098 177896 -25698
rect 178296 -26098 178496 -25698
rect 197496 -25898 200896 -25698
rect 197496 -26098 197696 -25898
rect 197896 -26098 198096 -25898
rect 198296 -26098 200896 -25898
rect 201296 -26098 204496 -25698
rect 204896 -26098 208296 -25698
rect 208696 -26098 208702 -25698
rect 172286 -26103 172506 -26098
rect 172686 -26103 172906 -26098
rect 173086 -26103 173306 -26098
rect 197686 -26103 197906 -26098
rect 198086 -26103 198306 -26098
rect 233696 -26893 236096 -26698
rect 233696 -26898 236106 -26893
rect 233696 -27098 235496 -26898
rect 235696 -27098 235896 -26898
rect 236096 -27098 236106 -26898
rect 233696 -27103 236106 -27098
rect 233696 -27298 236096 -27103
rect 228296 -29698 229296 -27598
rect 235096 -27698 236096 -27298
rect 165995 -40298 166405 -40295
rect 166891 -40298 167301 -40293
rect 145768 -40299 177096 -40298
rect 145768 -40300 168697 -40299
rect 145768 -40498 166000 -40300
rect 145768 -40698 146096 -40498
rect 146296 -40698 146496 -40498
rect 146696 -40698 166000 -40498
rect 146086 -40703 146306 -40698
rect 146486 -40703 146706 -40698
rect 165995 -40700 166000 -40698
rect 166400 -40697 168697 -40300
rect 169095 -40697 172497 -40299
rect 172895 -40697 176297 -40299
rect 176695 -40697 177096 -40299
rect 166400 -40698 177096 -40697
rect 178496 -40303 198896 -40298
rect 178496 -40498 196405 -40303
rect 178496 -40698 178896 -40498
rect 179096 -40698 179296 -40498
rect 179496 -40693 196405 -40498
rect 196795 -40693 198896 -40303
rect 179496 -40698 198896 -40693
rect 199296 -40698 202696 -40298
rect 203096 -40698 206296 -40298
rect 206696 -40698 208696 -40298
rect 166400 -40700 166405 -40698
rect 165995 -40705 166405 -40700
rect 166891 -40703 167301 -40698
rect 178886 -40703 179106 -40698
rect 179286 -40703 179506 -40698
rect 179386 -42798 179396 -42398
rect 179796 -42798 179806 -42398
rect 184086 -43498 184096 -43098
rect 184496 -43498 185496 -43098
rect 185896 -43498 185902 -43098
rect 215686 -43298 215696 -42898
rect 216096 -43298 217096 -42898
rect 217496 -43298 217502 -42898
rect 185486 -43503 185606 -43498
rect 185686 -43503 185815 -43498
rect 186686 -44098 186906 -44093
rect 186596 -44298 186696 -44098
rect 186896 -44298 236396 -44098
rect 186596 -44498 235496 -44298
rect 235696 -44498 235896 -44298
rect 236096 -44498 236396 -44298
rect 186596 -44698 186696 -44498
rect 186896 -44698 236396 -44498
rect 186596 -44898 235496 -44698
rect 235696 -44898 235896 -44698
rect 236096 -44898 236396 -44698
rect 179396 -45093 183996 -44998
rect 179396 -45098 184006 -45093
rect 186596 -45098 186696 -44898
rect 186896 -45098 236396 -44898
rect 179386 -45198 179396 -45098
rect 179496 -45198 179596 -45098
rect 179696 -45198 183696 -45098
rect 183796 -45198 183896 -45098
rect 183996 -45198 184006 -45098
rect 186686 -45103 186906 -45098
rect 183686 -45203 183806 -45198
rect 183886 -45203 184006 -45198
rect 214786 -45398 215006 -45393
rect 210596 -45498 214796 -45398
rect 210586 -45598 210596 -45498
rect 210696 -45598 210796 -45498
rect 210896 -45598 214796 -45498
rect 214996 -45598 215006 -45398
rect 214786 -45603 215006 -45598
rect 177990 -46298 178210 -46295
rect 220486 -46298 220706 -46293
rect 177900 -46300 181296 -46298
rect 177900 -46500 178000 -46300
rect 178200 -46498 181296 -46300
rect 220486 -46498 220496 -46298
rect 220696 -46498 236296 -46298
rect 178200 -46500 183496 -46498
rect 177900 -46600 183496 -46500
rect 177900 -46800 178000 -46600
rect 178200 -46800 183496 -46600
rect 177900 -46898 183496 -46800
rect 208300 -46600 215696 -46498
rect 220486 -46503 235496 -46498
rect 208300 -46800 208400 -46600
rect 208600 -46698 215696 -46600
rect 220596 -46693 235496 -46503
rect 220486 -46698 235496 -46693
rect 235696 -46698 235896 -46498
rect 236096 -46698 236296 -46498
rect 208600 -46800 217496 -46698
rect 208300 -46898 217496 -46800
rect 220486 -46898 220496 -46698
rect 220696 -46898 236296 -46698
rect 178600 -46900 178800 -46898
rect 208300 -46900 217491 -46898
rect 171990 -47000 172310 -46995
rect 171990 -47300 172000 -47000
rect 172300 -47300 172310 -47000
rect 171990 -47305 172310 -47300
rect 202390 -47000 202710 -46995
rect 202390 -47300 202400 -47000
rect 202700 -47300 202710 -47000
rect 208300 -47098 208400 -46900
rect 208390 -47100 208400 -47098
rect 208600 -46968 217491 -46900
rect 220486 -46903 220706 -46898
rect 208600 -47098 215696 -46968
rect 208600 -47100 208610 -47098
rect 208390 -47105 208610 -47100
rect 202390 -47305 202710 -47300
rect 187086 -47498 187306 -47493
rect 185896 -47698 187096 -47498
rect 187296 -47698 187306 -47498
rect 187086 -47703 187306 -47698
rect 185486 -47998 185606 -47993
rect 185486 -48098 185496 -47998
rect 185596 -48098 185606 -47998
rect 185486 -48103 185606 -48098
rect 185786 -47998 185906 -47993
rect 185786 -48098 185796 -47998
rect 185896 -48098 185906 -47998
rect 185786 -48103 185906 -48098
rect 217086 -47998 217206 -47993
rect 217086 -48098 217096 -47998
rect 217196 -48098 217206 -47998
rect 217086 -48103 217206 -48098
rect 217286 -47998 217406 -47993
rect 217286 -48098 217296 -47998
rect 217396 -48098 217406 -47998
rect 217286 -48103 217406 -48098
rect 179496 -48698 220896 -48498
rect 179496 -48898 187096 -48698
rect 187296 -48898 219696 -48698
rect 219896 -48898 220896 -48698
rect 179496 -50098 220896 -48898
rect 180886 -51298 180896 -50898
rect 181296 -51298 181306 -50898
rect 214886 -51298 214896 -50898
rect 215296 -51298 215306 -50898
rect 181086 -51303 181306 -51298
rect 215086 -51303 215306 -51298
<< via3 >>
rect 170096 -15098 170496 -14698
rect 170696 -15098 171096 -14698
rect 201696 -15098 202096 -14698
rect 202296 -15098 202696 -14698
rect 227296 -15098 227696 -14698
rect 227896 -15098 228296 -14698
rect 148496 -24498 148796 -24298
rect 148496 -24598 148596 -24498
rect 148596 -24598 148696 -24498
rect 148696 -24598 148796 -24498
rect 180396 -24398 180796 -24298
rect 180396 -24598 180496 -24398
rect 180496 -24598 180696 -24398
rect 180696 -24598 180796 -24398
rect 180396 -24698 180796 -24598
rect 170496 -26098 170896 -25698
rect 174296 -26098 174696 -25698
rect 177896 -26098 178296 -25698
rect 200896 -26098 201296 -25698
rect 204496 -26098 204896 -25698
rect 208296 -26098 208696 -25698
rect 168697 -40697 169095 -40299
rect 172497 -40697 172895 -40299
rect 176297 -40697 176695 -40299
rect 198896 -40698 199296 -40298
rect 202696 -40698 203096 -40298
rect 206296 -40698 206696 -40298
rect 179396 -42798 179796 -42398
rect 184096 -43498 184496 -43098
rect 185496 -43498 185896 -43098
rect 215696 -43298 216096 -42898
rect 217096 -43298 217496 -42898
rect 179396 -45198 179496 -45098
rect 179596 -45198 179696 -45098
rect 210596 -45598 210696 -45498
rect 210796 -45598 210896 -45498
rect 172000 -47300 172300 -47000
rect 202400 -47300 202700 -47000
rect 185496 -48098 185596 -47998
rect 185796 -48098 185896 -47998
rect 217096 -48098 217196 -47998
rect 217296 -48098 217396 -47998
rect 180896 -51098 181296 -50898
rect 180896 -51298 181096 -51098
rect 181096 -51298 181296 -51098
rect 214896 -51098 215296 -50898
rect 214896 -51298 215096 -51098
rect 215096 -51298 215296 -51098
<< metal4 >>
rect 166696 -3898 169896 -3698
rect 166696 -4298 166896 -3898
rect 167296 -4298 167696 -3898
rect 168096 -4298 168496 -3898
rect 168896 -4298 169296 -3898
rect 169696 -4298 169896 -3898
rect 166696 -4698 169896 -4298
rect 166696 -5098 166896 -4698
rect 167296 -5098 167696 -4698
rect 168096 -5098 168496 -4698
rect 168896 -5098 169296 -4698
rect 169696 -5098 169896 -4698
rect 166696 -5498 169896 -5098
rect 166696 -5898 166896 -5498
rect 167296 -5898 167696 -5498
rect 168096 -5898 168496 -5498
rect 168896 -5898 169296 -5498
rect 169696 -5898 169896 -5498
rect 166696 -6298 169896 -5898
rect 166696 -6698 166896 -6298
rect 167296 -6698 167696 -6298
rect 168096 -6698 168496 -6298
rect 168896 -6698 169296 -6298
rect 169696 -6698 169896 -6298
rect 166696 -7098 169896 -6698
rect 166696 -7498 166896 -7098
rect 167296 -7498 167696 -7098
rect 168096 -7498 168496 -7098
rect 168896 -7498 169296 -7098
rect 169696 -7498 169896 -7098
rect 166696 -7698 169896 -7498
rect 198496 -3898 201696 -3698
rect 198496 -4298 198696 -3898
rect 199096 -4298 199496 -3898
rect 199896 -4298 200296 -3898
rect 200696 -4298 201096 -3898
rect 201496 -4298 201696 -3898
rect 198496 -4698 201696 -4298
rect 198496 -5098 198696 -4698
rect 199096 -5098 199496 -4698
rect 199896 -5098 200296 -4698
rect 200696 -5098 201096 -4698
rect 201496 -5098 201696 -4698
rect 198496 -5498 201696 -5098
rect 198496 -5898 198696 -5498
rect 199096 -5898 199496 -5498
rect 199896 -5898 200296 -5498
rect 200696 -5898 201096 -5498
rect 201496 -5898 201696 -5498
rect 198496 -6298 201696 -5898
rect 198496 -6698 198696 -6298
rect 199096 -6698 199496 -6298
rect 199896 -6698 200296 -6298
rect 200696 -6698 201096 -6298
rect 201496 -6698 201696 -6298
rect 198496 -7098 201696 -6698
rect 198496 -7498 198696 -7098
rect 199096 -7498 199496 -7098
rect 199896 -7498 200296 -7098
rect 200696 -7498 201096 -7098
rect 201496 -7498 201696 -7098
rect 198496 -7698 201696 -7498
rect 229896 -3898 233096 -3698
rect 229896 -4298 230096 -3898
rect 230496 -4298 230896 -3898
rect 231296 -4298 231696 -3898
rect 232096 -4298 232496 -3898
rect 232896 -4298 233096 -3898
rect 229896 -4698 233096 -4298
rect 229896 -5098 230096 -4698
rect 230496 -5098 230896 -4698
rect 231296 -5098 231696 -4698
rect 232096 -5098 232496 -4698
rect 232896 -5098 233096 -4698
rect 229896 -5498 233096 -5098
rect 229896 -5898 230096 -5498
rect 230496 -5898 230896 -5498
rect 231296 -5898 231696 -5498
rect 232096 -5898 232496 -5498
rect 232896 -5898 233096 -5498
rect 229896 -6298 233096 -5898
rect 229896 -6698 230096 -6298
rect 230496 -6698 230896 -6298
rect 231296 -6698 231696 -6298
rect 232096 -6698 232496 -6298
rect 232896 -6698 233096 -6298
rect 229896 -7098 233096 -6698
rect 229896 -7498 230096 -7098
rect 230496 -7498 230896 -7098
rect 231296 -7498 231696 -7098
rect 232096 -7498 232496 -7098
rect 232896 -7498 233096 -7098
rect 229896 -7698 233096 -7498
rect 166696 -15298 169696 -7698
rect 170095 -14698 170497 -14697
rect 170095 -15098 170096 -14698
rect 170496 -15098 170497 -14698
rect 170095 -15099 170497 -15098
rect 170695 -14698 171097 -14697
rect 170695 -15098 170696 -14698
rect 171096 -15098 171097 -14698
rect 170695 -15099 171097 -15098
rect 198496 -15298 201496 -7698
rect 201695 -14698 202097 -14697
rect 201695 -15098 201696 -14698
rect 202096 -15098 202097 -14698
rect 201695 -15099 202097 -15098
rect 202295 -14698 202697 -14697
rect 202295 -15098 202296 -14698
rect 202696 -15098 202697 -14698
rect 202295 -15099 202697 -15098
rect 227295 -14698 227697 -14697
rect 227295 -15098 227296 -14698
rect 227696 -15098 227697 -14698
rect 227295 -15099 227697 -15098
rect 227895 -14698 228297 -14697
rect 227895 -15098 227896 -14698
rect 228296 -15098 228297 -14698
rect 227895 -15099 228297 -15098
rect 148495 -24298 148797 -24297
rect 148495 -24598 148496 -24298
rect 148796 -24598 148797 -24298
rect 148495 -24599 148797 -24598
rect 180395 -24298 180797 -24297
rect 180395 -24698 180396 -24298
rect 180796 -24698 180797 -24298
rect 180395 -24699 180797 -24698
rect 170495 -25698 170897 -25697
rect 170495 -26098 170496 -25698
rect 170896 -26098 170897 -25698
rect 170495 -26099 170897 -26098
rect 174295 -25698 174697 -25697
rect 174295 -26098 174296 -25698
rect 174696 -26098 174697 -25698
rect 174295 -26099 174697 -26098
rect 177895 -25698 178297 -25697
rect 177895 -26098 177896 -25698
rect 178296 -26098 178297 -25698
rect 177895 -26099 178297 -26098
rect 200895 -25698 201297 -25697
rect 200895 -26098 200896 -25698
rect 201296 -26098 201297 -25698
rect 200895 -26099 201297 -26098
rect 204495 -25698 204897 -25697
rect 204495 -26098 204496 -25698
rect 204896 -26098 204897 -25698
rect 204495 -26099 204897 -26098
rect 208295 -25698 208697 -25697
rect 208295 -26098 208296 -25698
rect 208696 -26098 208697 -25698
rect 208295 -26099 208697 -26098
rect 170496 -26298 170896 -26099
rect 174296 -26298 174696 -26099
rect 177896 -26298 178296 -26099
rect 200896 -26298 201296 -26099
rect 204496 -26298 204896 -26099
rect 208296 -26298 208696 -26099
rect 168696 -40299 169096 -39898
rect 168696 -40697 168697 -40299
rect 169095 -40697 169096 -40299
rect 168696 -40698 169096 -40697
rect 172496 -40299 172896 -39898
rect 172496 -40697 172497 -40299
rect 172895 -40697 172896 -40299
rect 172496 -40698 172896 -40697
rect 176296 -40299 176696 -39898
rect 198896 -40297 199296 -39898
rect 202696 -40297 203096 -39898
rect 206296 -40297 206696 -39898
rect 176296 -40697 176297 -40299
rect 176695 -40697 176696 -40299
rect 176296 -40698 176696 -40697
rect 198895 -40298 199297 -40297
rect 198895 -40698 198896 -40298
rect 199296 -40698 199297 -40298
rect 198895 -40699 199297 -40698
rect 202695 -40298 203097 -40297
rect 202695 -40698 202696 -40298
rect 203096 -40698 203097 -40298
rect 202695 -40699 203097 -40698
rect 206295 -40298 206697 -40297
rect 206295 -40698 206296 -40298
rect 206696 -40698 206697 -40298
rect 206295 -40699 206697 -40698
rect 229896 -41103 232896 -7698
rect 229696 -41303 232896 -41103
rect 148496 -44098 153296 -41498
rect 179395 -42398 179797 -42397
rect 179395 -42798 179396 -42398
rect 179796 -42798 179797 -42398
rect 179395 -42799 179797 -42798
rect 148496 -44498 149496 -44098
rect 149896 -44498 150296 -44098
rect 150696 -44498 151096 -44098
rect 151496 -44498 151896 -44098
rect 152296 -44498 153296 -44098
rect 148496 -44898 153296 -44498
rect 148496 -45298 149496 -44898
rect 149896 -45298 150296 -44898
rect 150696 -45298 151096 -44898
rect 151496 -45298 151896 -44898
rect 152296 -45298 153296 -44898
rect 179396 -45097 179796 -42799
rect 179395 -45098 179796 -45097
rect 179395 -45198 179396 -45098
rect 179496 -45198 179596 -45098
rect 179696 -45198 179796 -45098
rect 179395 -45199 179796 -45198
rect 148496 -45698 153296 -45298
rect 179396 -45398 179796 -45199
rect 180296 -43098 185096 -41698
rect 229696 -41703 229895 -41303
rect 230295 -41703 230695 -41303
rect 231095 -41703 231495 -41303
rect 231895 -41703 232295 -41303
rect 232695 -41703 232896 -41303
rect 180296 -43498 184096 -43098
rect 184496 -43498 185096 -43098
rect 180296 -44098 185096 -43498
rect 185495 -43098 185897 -43097
rect 185495 -43498 185496 -43098
rect 185896 -43498 185897 -43098
rect 185495 -43499 185897 -43498
rect 180296 -44498 181296 -44098
rect 181696 -44498 182096 -44098
rect 182496 -44498 182896 -44098
rect 183296 -44498 183696 -44098
rect 184096 -44498 185096 -44098
rect 180296 -44898 185096 -44498
rect 180296 -45298 181296 -44898
rect 181696 -45298 182096 -44898
rect 182496 -45298 182896 -44898
rect 183296 -45298 183696 -44898
rect 184096 -45298 185096 -44898
rect 148496 -46098 149496 -45698
rect 149896 -46098 150296 -45698
rect 150696 -46098 151096 -45698
rect 151496 -46098 151896 -45698
rect 152296 -46098 153296 -45698
rect 148496 -46498 153296 -46098
rect 148496 -46898 149496 -46498
rect 149896 -46898 150296 -46498
rect 150696 -46898 151096 -46498
rect 151496 -46898 151896 -46498
rect 152296 -46898 153296 -46498
rect 148496 -47298 153296 -46898
rect 180296 -45698 185096 -45298
rect 180296 -46098 181296 -45698
rect 181696 -46098 182096 -45698
rect 182496 -46098 182896 -45698
rect 183296 -46098 183696 -45698
rect 184096 -46098 185096 -45698
rect 180296 -46498 185096 -46098
rect 180296 -46898 181296 -46498
rect 181696 -46898 182096 -46498
rect 182496 -46898 182896 -46498
rect 183296 -46898 183696 -46498
rect 184096 -46898 185096 -46498
rect 148496 -47698 149496 -47298
rect 149896 -47698 150296 -47298
rect 150696 -47698 151096 -47298
rect 151496 -47698 151896 -47298
rect 152296 -47698 153296 -47298
rect 171999 -47000 172301 -46999
rect 171999 -47300 172000 -47000
rect 172300 -47300 172301 -47000
rect 171999 -47301 172301 -47300
rect 180296 -47298 185096 -46898
rect 148496 -47898 153296 -47698
rect 180296 -47698 181296 -47298
rect 181696 -47698 182096 -47298
rect 182496 -47698 182896 -47298
rect 183296 -47698 183696 -47298
rect 184096 -47698 185096 -47298
rect 180296 -47898 185096 -47698
rect 185496 -47997 185896 -43499
rect 210596 -45197 210996 -42798
rect 210595 -45299 210996 -45197
rect 210596 -45497 210996 -45299
rect 210595 -45498 210996 -45497
rect 210595 -45598 210596 -45498
rect 210696 -45598 210796 -45498
rect 210896 -45598 210996 -45498
rect 210595 -45599 210996 -45598
rect 210596 -45698 210996 -45599
rect 211696 -42898 216496 -41898
rect 229696 -42103 232896 -41703
rect 229696 -42503 229895 -42103
rect 230295 -42503 230695 -42103
rect 231095 -42503 231495 -42103
rect 231895 -42503 232295 -42103
rect 232695 -42503 232896 -42103
rect 229696 -42798 232896 -42503
rect 211696 -43298 215696 -42898
rect 216096 -43298 216496 -42898
rect 211696 -44098 216496 -43298
rect 217095 -42898 217497 -42897
rect 217095 -43298 217096 -42898
rect 217496 -43298 217497 -42898
rect 217095 -43299 217497 -43298
rect 211696 -44498 212696 -44098
rect 213096 -44498 213496 -44098
rect 213896 -44498 214296 -44098
rect 214696 -44498 215096 -44098
rect 215496 -44498 216496 -44098
rect 211696 -44898 216496 -44498
rect 211696 -45298 212696 -44898
rect 213096 -45298 213496 -44898
rect 213896 -45298 214296 -44898
rect 214696 -45298 215096 -44898
rect 215496 -45298 216496 -44898
rect 211696 -45698 216496 -45298
rect 211696 -46098 212696 -45698
rect 213096 -46098 213496 -45698
rect 213896 -46098 214296 -45698
rect 214696 -46098 215096 -45698
rect 215496 -46098 216496 -45698
rect 211696 -46498 216496 -46098
rect 211696 -46898 212696 -46498
rect 213096 -46898 213496 -46498
rect 213896 -46898 214296 -46498
rect 214696 -46898 215096 -46498
rect 215496 -46898 216496 -46498
rect 202399 -47000 202701 -46999
rect 202399 -47300 202400 -47000
rect 202700 -47300 202701 -47000
rect 202399 -47301 202701 -47300
rect 211696 -47298 216496 -46898
rect 211696 -47698 212696 -47298
rect 213096 -47698 213496 -47298
rect 213896 -47698 214296 -47298
rect 214696 -47698 215096 -47298
rect 215496 -47698 216496 -47298
rect 211696 -47898 216496 -47698
rect 217096 -47997 217496 -43299
rect 185495 -47998 185897 -47997
rect 185495 -48098 185496 -47998
rect 185596 -48098 185796 -47998
rect 185896 -48098 185897 -47998
rect 185495 -48099 185597 -48098
rect 185795 -48099 185897 -48098
rect 217095 -47998 217496 -47997
rect 217095 -48098 217096 -47998
rect 217196 -48098 217296 -47998
rect 217396 -48098 217496 -47998
rect 217095 -48099 217197 -48098
rect 217295 -48099 217397 -48098
rect 180895 -50898 181297 -50897
rect 180895 -51298 180896 -50898
rect 181296 -51298 181297 -50898
rect 180895 -51299 181297 -51298
rect 214895 -50898 215297 -50897
rect 214895 -51298 214896 -50898
rect 215296 -51298 215297 -50898
rect 214895 -51299 215297 -51298
<< via4 >>
rect 166896 -4298 167296 -3898
rect 167696 -4298 168096 -3898
rect 168496 -4298 168896 -3898
rect 169296 -4298 169696 -3898
rect 166896 -5098 167296 -4698
rect 167696 -5098 168096 -4698
rect 168496 -5098 168896 -4698
rect 169296 -5098 169696 -4698
rect 166896 -5898 167296 -5498
rect 167696 -5898 168096 -5498
rect 168496 -5898 168896 -5498
rect 169296 -5898 169696 -5498
rect 166896 -6698 167296 -6298
rect 167696 -6698 168096 -6298
rect 168496 -6698 168896 -6298
rect 169296 -6698 169696 -6298
rect 166896 -7498 167296 -7098
rect 167696 -7498 168096 -7098
rect 168496 -7498 168896 -7098
rect 169296 -7498 169696 -7098
rect 198696 -4298 199096 -3898
rect 199496 -4298 199896 -3898
rect 200296 -4298 200696 -3898
rect 201096 -4298 201496 -3898
rect 198696 -5098 199096 -4698
rect 199496 -5098 199896 -4698
rect 200296 -5098 200696 -4698
rect 201096 -5098 201496 -4698
rect 198696 -5898 199096 -5498
rect 199496 -5898 199896 -5498
rect 200296 -5898 200696 -5498
rect 201096 -5898 201496 -5498
rect 198696 -6698 199096 -6298
rect 199496 -6698 199896 -6298
rect 200296 -6698 200696 -6298
rect 201096 -6698 201496 -6298
rect 198696 -7498 199096 -7098
rect 199496 -7498 199896 -7098
rect 200296 -7498 200696 -7098
rect 201096 -7498 201496 -7098
rect 230096 -4298 230496 -3898
rect 230896 -4298 231296 -3898
rect 231696 -4298 232096 -3898
rect 232496 -4298 232896 -3898
rect 230096 -5098 230496 -4698
rect 230896 -5098 231296 -4698
rect 231696 -5098 232096 -4698
rect 232496 -5098 232896 -4698
rect 230096 -5898 230496 -5498
rect 230896 -5898 231296 -5498
rect 231696 -5898 232096 -5498
rect 232496 -5898 232896 -5498
rect 230096 -6698 230496 -6298
rect 230896 -6698 231296 -6298
rect 231696 -6698 232096 -6298
rect 232496 -6698 232896 -6298
rect 230096 -7498 230496 -7098
rect 230896 -7498 231296 -7098
rect 231696 -7498 232096 -7098
rect 232496 -7498 232896 -7098
rect 170096 -15098 170496 -14698
rect 170696 -15098 171096 -14698
rect 201696 -15098 202096 -14698
rect 202296 -15098 202696 -14698
rect 227296 -15098 227696 -14698
rect 227896 -15098 228296 -14698
rect 179396 -42798 179796 -42398
rect 149496 -44498 149896 -44098
rect 150296 -44498 150696 -44098
rect 151096 -44498 151496 -44098
rect 151896 -44498 152296 -44098
rect 149496 -45298 149896 -44898
rect 150296 -45298 150696 -44898
rect 151096 -45298 151496 -44898
rect 151896 -45298 152296 -44898
rect 229895 -41703 230295 -41303
rect 230695 -41703 231095 -41303
rect 231495 -41703 231895 -41303
rect 232295 -41703 232695 -41303
rect 210596 -42798 210996 -42398
rect 181296 -44498 181696 -44098
rect 182096 -44498 182496 -44098
rect 182896 -44498 183296 -44098
rect 183696 -44498 184096 -44098
rect 181296 -45298 181696 -44898
rect 182096 -45298 182496 -44898
rect 182896 -45298 183296 -44898
rect 183696 -45298 184096 -44898
rect 149496 -46098 149896 -45698
rect 150296 -46098 150696 -45698
rect 151096 -46098 151496 -45698
rect 151896 -46098 152296 -45698
rect 149496 -46898 149896 -46498
rect 150296 -46898 150696 -46498
rect 151096 -46898 151496 -46498
rect 151896 -46898 152296 -46498
rect 181296 -46098 181696 -45698
rect 182096 -46098 182496 -45698
rect 182896 -46098 183296 -45698
rect 183696 -46098 184096 -45698
rect 181296 -46898 181696 -46498
rect 182096 -46898 182496 -46498
rect 182896 -46898 183296 -46498
rect 183696 -46898 184096 -46498
rect 149496 -47698 149896 -47298
rect 150296 -47698 150696 -47298
rect 151096 -47698 151496 -47298
rect 151896 -47698 152296 -47298
rect 172000 -47300 172300 -47000
rect 181296 -47698 181696 -47298
rect 182096 -47698 182496 -47298
rect 182896 -47698 183296 -47298
rect 183696 -47698 184096 -47298
rect 229895 -42503 230295 -42103
rect 230695 -42503 231095 -42103
rect 231495 -42503 231895 -42103
rect 232295 -42503 232695 -42103
rect 212696 -44498 213096 -44098
rect 213496 -44498 213896 -44098
rect 214296 -44498 214696 -44098
rect 215096 -44498 215496 -44098
rect 212696 -45298 213096 -44898
rect 213496 -45298 213896 -44898
rect 214296 -45298 214696 -44898
rect 215096 -45298 215496 -44898
rect 212696 -46098 213096 -45698
rect 213496 -46098 213896 -45698
rect 214296 -46098 214696 -45698
rect 215096 -46098 215496 -45698
rect 212696 -46898 213096 -46498
rect 213496 -46898 213896 -46498
rect 214296 -46898 214696 -46498
rect 215096 -46898 215496 -46498
rect 202400 -47300 202700 -47000
rect 212696 -47698 213096 -47298
rect 213496 -47698 213896 -47298
rect 214296 -47698 214696 -47298
rect 215096 -47698 215496 -47298
rect 180896 -51298 181296 -50898
rect 214896 -51298 215296 -50898
<< metal5 >>
rect 166696 -3898 233096 -3698
rect 166696 -4298 166896 -3898
rect 167296 -4298 167696 -3898
rect 168096 -4298 168496 -3898
rect 168896 -4298 169296 -3898
rect 169696 -4298 198696 -3898
rect 199096 -4298 199496 -3898
rect 199896 -4298 200296 -3898
rect 200696 -4298 201096 -3898
rect 201496 -4298 230096 -3898
rect 230496 -4298 230896 -3898
rect 231296 -4298 231696 -3898
rect 232096 -4298 232496 -3898
rect 232896 -4298 233096 -3898
rect 166696 -4698 233096 -4298
rect 166696 -5098 166896 -4698
rect 167296 -5098 167696 -4698
rect 168096 -5098 168496 -4698
rect 168896 -5098 169296 -4698
rect 169696 -5098 198696 -4698
rect 199096 -5098 199496 -4698
rect 199896 -5098 200296 -4698
rect 200696 -5098 201096 -4698
rect 201496 -5098 230096 -4698
rect 230496 -5098 230896 -4698
rect 231296 -5098 231696 -4698
rect 232096 -5098 232496 -4698
rect 232896 -5098 233096 -4698
rect 166696 -5498 233096 -5098
rect 166696 -5898 166896 -5498
rect 167296 -5898 167696 -5498
rect 168096 -5898 168496 -5498
rect 168896 -5898 169296 -5498
rect 169696 -5898 198696 -5498
rect 199096 -5898 199496 -5498
rect 199896 -5898 200296 -5498
rect 200696 -5898 201096 -5498
rect 201496 -5898 230096 -5498
rect 230496 -5898 230896 -5498
rect 231296 -5898 231696 -5498
rect 232096 -5898 232496 -5498
rect 232896 -5898 233096 -5498
rect 166696 -6298 233096 -5898
rect 166696 -6698 166896 -6298
rect 167296 -6698 167696 -6298
rect 168096 -6698 168496 -6298
rect 168896 -6698 169296 -6298
rect 169696 -6698 198696 -6298
rect 199096 -6698 199496 -6298
rect 199896 -6698 200296 -6298
rect 200696 -6698 201096 -6298
rect 201496 -6698 230096 -6298
rect 230496 -6698 230896 -6298
rect 231296 -6698 231696 -6298
rect 232096 -6698 232496 -6298
rect 232896 -6698 233096 -6298
rect 166696 -7098 233096 -6698
rect 166696 -7498 166896 -7098
rect 167296 -7498 167696 -7098
rect 168096 -7498 168496 -7098
rect 168896 -7498 169296 -7098
rect 169696 -7498 198696 -7098
rect 199096 -7498 199496 -7098
rect 199896 -7498 200296 -7098
rect 200696 -7498 201096 -7098
rect 201496 -7498 230096 -7098
rect 230496 -7498 230896 -7098
rect 231296 -7498 231696 -7098
rect 232096 -7498 232496 -7098
rect 232896 -7498 233096 -7098
rect 166696 -7698 233096 -7498
rect 169596 -14698 228896 -13598
rect 169596 -15098 170096 -14698
rect 170496 -15098 170696 -14698
rect 171096 -15098 201696 -14698
rect 202096 -15098 202296 -14698
rect 202696 -15098 227296 -14698
rect 227696 -15098 227896 -14698
rect 228296 -15098 228896 -14698
rect 169596 -15198 228896 -15098
rect 179396 -41303 232896 -40798
rect 179396 -41703 229895 -41303
rect 230295 -41703 230695 -41303
rect 231095 -41703 231495 -41303
rect 231895 -41703 232295 -41303
rect 232695 -41703 232896 -41303
rect 179396 -42103 232896 -41703
rect 179396 -42374 229895 -42103
rect 179372 -42398 229895 -42374
rect 179372 -42798 179396 -42398
rect 179796 -42798 210596 -42398
rect 210996 -42503 229895 -42398
rect 230295 -42503 230695 -42103
rect 231095 -42503 231495 -42103
rect 231895 -42503 232295 -42103
rect 232695 -42503 232896 -42103
rect 210996 -42798 232896 -42503
rect 179372 -42822 179820 -42798
rect 210572 -42822 211020 -42798
rect 148496 -44098 216496 -43898
rect 148496 -44498 149496 -44098
rect 149896 -44498 150296 -44098
rect 150696 -44498 151096 -44098
rect 151496 -44498 151896 -44098
rect 152296 -44498 181296 -44098
rect 181696 -44498 182096 -44098
rect 182496 -44498 182896 -44098
rect 183296 -44498 183696 -44098
rect 184096 -44498 212696 -44098
rect 213096 -44498 213496 -44098
rect 213896 -44498 214296 -44098
rect 214696 -44498 215096 -44098
rect 215496 -44498 216496 -44098
rect 148496 -44898 216496 -44498
rect 148496 -45298 149496 -44898
rect 149896 -45298 150296 -44898
rect 150696 -45298 151096 -44898
rect 151496 -45298 151896 -44898
rect 152296 -45298 181296 -44898
rect 181696 -45298 182096 -44898
rect 182496 -45298 182896 -44898
rect 183296 -45298 183696 -44898
rect 184096 -45298 212696 -44898
rect 213096 -45298 213496 -44898
rect 213896 -45298 214296 -44898
rect 214696 -45298 215096 -44898
rect 215496 -45298 216496 -44898
rect 148496 -45698 216496 -45298
rect 148496 -46098 149496 -45698
rect 149896 -46098 150296 -45698
rect 150696 -46098 151096 -45698
rect 151496 -46098 151896 -45698
rect 152296 -46098 181296 -45698
rect 181696 -46098 182096 -45698
rect 182496 -46098 182896 -45698
rect 183296 -46098 183696 -45698
rect 184096 -46098 212696 -45698
rect 213096 -46098 213496 -45698
rect 213896 -46098 214296 -45698
rect 214696 -46098 215096 -45698
rect 215496 -46098 216496 -45698
rect 148496 -46498 216496 -46098
rect 148496 -46898 149496 -46498
rect 149896 -46898 150296 -46498
rect 150696 -46898 151096 -46498
rect 151496 -46898 151896 -46498
rect 152296 -46898 181296 -46498
rect 181696 -46898 182096 -46498
rect 182496 -46898 182896 -46498
rect 183296 -46898 183696 -46498
rect 184096 -46898 212696 -46498
rect 213096 -46898 213496 -46498
rect 213896 -46898 214296 -46498
rect 214696 -46898 215096 -46498
rect 215496 -46898 216496 -46498
rect 148496 -47000 216496 -46898
rect 148496 -47298 172000 -47000
rect 148496 -47698 149496 -47298
rect 149896 -47698 150296 -47298
rect 150696 -47698 151096 -47298
rect 151496 -47698 151896 -47298
rect 152296 -47300 172000 -47298
rect 172300 -47298 202400 -47000
rect 172300 -47300 181296 -47298
rect 152296 -47698 181296 -47300
rect 181696 -47698 182096 -47298
rect 182496 -47698 182896 -47298
rect 183296 -47698 183696 -47298
rect 184096 -47300 202400 -47298
rect 202700 -47298 216496 -47000
rect 202700 -47300 212696 -47298
rect 184096 -47698 212696 -47300
rect 213096 -47698 213496 -47298
rect 213896 -47698 214296 -47298
rect 214696 -47698 215096 -47298
rect 215496 -47698 216496 -47298
rect 148496 -47898 216496 -47698
rect 179496 -50898 220896 -50698
rect 179496 -51298 180896 -50898
rect 181296 -51298 214896 -50898
rect 215296 -51298 220896 -50898
rect 179496 -52298 220896 -51298
use 1Bit_Clk_ADC  1Bit_Clk_ADC_0
timestamp 1717026683
transform 1 0 228796 0 1 -26798
box -22500 -15300 5388 23160
use 1Bit_DAC  1Bit_DAC_0
timestamp 1716868724
transform -1 0 222101 0 1 -45318
box 1490 -2780 7005 210
use 1Bit_DAC_Inv  1Bit_DAC_Inv_0
timestamp 1716868724
transform -1 0 188101 0 1 -45318
box 1490 -2780 7005 210
use C2S2_Amp_F_I  C2S2_Amp_F_I_0
timestamp 1716868724
transform 1 0 145104 0 1 -704888
box 29796 662788 57684 701260
use C2S2_Amp_F_I  C2S2_Amp_F_I_1
timestamp 1716868724
transform 1 0 113304 0 1 -704888
box 29796 662788 57684 701260
use sky130_fd_pr__cap_mim_m3_1_Z67P85  sky130_fd_pr__cap_mim_m3_1_Z67P85_0
timestamp 1716868724
transform 1 0 172804 0 1 -33178
box -5508 -6920 5508 6920
use sky130_fd_pr__cap_mim_m3_1_Z67P85  sky130_fd_pr__cap_mim_m3_1_Z67P85_1
timestamp 1716868724
transform 1 0 203004 0 1 -33178
box -5508 -6920 5508 6920
use sky130_fd_pr__res_xhigh_po_5p73_UF8E3R  sky130_fd_pr__res_xhigh_po_5p73_UF8E3R_0
timestamp 1716868724
transform 1 0 175223 0 1 -18188
box -3223 -6312 3223 6312
use sky130_fd_pr__res_xhigh_po_5p73_UF8E3R  sky130_fd_pr__res_xhigh_po_5p73_UF8E3R_1
timestamp 1716868724
transform 1 0 143723 0 1 -18188
box -3223 -6312 3223 6312
use sky130_fd_pr__res_xhigh_po_5p73_UF8E3R  sky130_fd_pr__res_xhigh_po_5p73_UF8E3R_2
timestamp 1716868724
transform 0 -1 172212 1 0 -44577
box -3223 -6312 3223 6312
use sky130_fd_pr__res_xhigh_po_5p73_UF8E3R  sky130_fd_pr__res_xhigh_po_5p73_UF8E3R_3
timestamp 1716868724
transform 0 -1 202612 1 0 -44577
box -3223 -6312 3223 6312
use sky130_fd_pr__cap_mim_m3_1_QPPWMY  XC1
timestamp 1716868724
transform 1 0 139404 0 1 -55212
box 0 0 1 1
use sky130_fd_pr__cap_mim_m3_1_QPPWMY  XC3
timestamp 1716868724
transform 1 0 135892 0 1 -17032
box 0 0 1 1
<< labels >>
rlabel metal5 166696 -7698 233096 -3698 1 VDD
port 2 n
rlabel metal5 179496 -52298 220896 -50698 1 VREFN
port 4 n
rlabel metal3 179496 -50098 220896 -48498 1 VREFP
port 3 n
rlabel metal3 140696 -24298 141696 -23298 1 SIG
port 5 n
rlabel metal3 235096 -27698 236096 -26698 1 OUT
port 6 n
rlabel metal5 169696 -15098 228696 -13698 1 VMID
port 7 n
rlabel metal3 228296 -29698 229296 -28698 1 CLK
port 8 n
rlabel metal5 148496 -47898 216496 -43898 1 GND
port 1 n
<< end >>
