magic
tech sky130A
magscale 1 2
timestamp 1717119771
<< metal1 >>
rect -30 20 20 10240
rect 180 10190 1070 10230
rect 180 10140 230 10190
rect 380 10140 430 10190
rect 570 10140 620 10190
rect 770 10140 820 10190
rect 960 10140 1010 10190
rect 70 6400 80 6460
rect 140 6400 150 6460
rect 260 6400 270 6460
rect 330 6400 340 6460
rect 460 6400 470 6460
rect 530 6400 540 6460
rect 650 6400 660 6460
rect 720 6400 730 6460
rect 850 6400 860 6460
rect 920 6400 930 6460
rect 1050 6400 1060 6460
rect 1120 6400 1130 6460
rect 60 6235 70 6295
rect 130 6235 140 6295
rect 260 6235 270 6295
rect 330 6235 340 6295
rect 460 6235 470 6295
rect 530 6235 540 6295
rect 650 6235 660 6295
rect 720 6235 730 6295
rect 850 6235 860 6295
rect 920 6235 930 6295
rect 1050 6235 1060 6295
rect 1120 6235 1130 6295
rect 60 6035 70 6095
rect 130 6035 140 6095
rect 260 6035 270 6095
rect 330 6035 340 6095
rect 460 6035 470 6095
rect 530 6035 540 6095
rect 650 6035 660 6095
rect 720 6035 730 6095
rect 850 6035 860 6095
rect 920 6035 930 6095
rect 1050 6035 1060 6095
rect 1120 6035 1130 6095
rect 60 5845 70 5905
rect 130 5845 140 5905
rect 260 5845 270 5905
rect 330 5845 340 5905
rect 460 5845 470 5905
rect 530 5845 540 5905
rect 650 5845 660 5905
rect 720 5845 730 5905
rect 850 5845 860 5905
rect 920 5845 930 5905
rect 1050 5845 1060 5905
rect 1120 5845 1130 5905
rect 60 5665 70 5725
rect 130 5665 140 5725
rect 260 5665 270 5725
rect 330 5665 340 5725
rect 460 5665 470 5725
rect 530 5665 540 5725
rect 650 5665 660 5725
rect 720 5665 730 5725
rect 850 5665 860 5725
rect 920 5665 930 5725
rect 1050 5665 1060 5725
rect 1120 5665 1130 5725
rect 60 5465 70 5525
rect 130 5465 140 5525
rect 260 5465 270 5525
rect 330 5465 340 5525
rect 460 5465 470 5525
rect 530 5465 540 5525
rect 650 5465 660 5525
rect 720 5465 730 5525
rect 850 5465 860 5525
rect 920 5465 930 5525
rect 1050 5465 1060 5525
rect 1120 5465 1130 5525
rect 60 5275 70 5335
rect 130 5275 140 5335
rect 260 5275 270 5335
rect 330 5275 340 5335
rect 460 5275 470 5335
rect 530 5275 540 5335
rect 650 5275 660 5335
rect 720 5275 730 5335
rect 850 5275 860 5335
rect 920 5275 930 5335
rect 1050 5275 1060 5335
rect 1120 5275 1130 5335
rect 60 5115 70 5175
rect 130 5115 140 5175
rect 260 5115 270 5175
rect 330 5115 340 5175
rect 460 5115 470 5175
rect 530 5115 540 5175
rect 650 5115 660 5175
rect 720 5115 730 5175
rect 850 5115 860 5175
rect 920 5115 930 5175
rect 1050 5115 1060 5175
rect 1120 5115 1130 5175
rect 60 4925 70 4985
rect 130 4925 140 4985
rect 260 4925 270 4985
rect 330 4925 340 4985
rect 460 4925 470 4985
rect 530 4925 540 4985
rect 650 4925 660 4985
rect 720 4925 730 4985
rect 850 4925 860 4985
rect 920 4925 930 4985
rect 1050 4925 1060 4985
rect 1120 4925 1130 4985
rect 60 4750 70 4810
rect 130 4750 140 4810
rect 260 4750 270 4810
rect 330 4750 340 4810
rect 460 4750 470 4810
rect 530 4750 540 4810
rect 650 4750 660 4810
rect 720 4750 730 4810
rect 850 4750 860 4810
rect 920 4750 930 4810
rect 1050 4750 1060 4810
rect 1120 4750 1130 4810
rect 60 4610 70 4670
rect 130 4610 140 4670
rect 260 4610 270 4670
rect 330 4610 340 4670
rect 460 4610 470 4670
rect 530 4610 540 4670
rect 650 4610 660 4670
rect 720 4610 730 4670
rect 850 4610 860 4670
rect 920 4610 930 4670
rect 1050 4610 1060 4670
rect 1120 4610 1130 4670
rect 180 120 230 170
rect 370 120 430 170
rect 570 120 630 170
rect 760 120 820 170
rect 960 120 1020 170
rect 120 80 1020 120
rect 1180 20 1230 10240
rect -30 -30 1230 20
<< via1 >>
rect 80 6400 140 6460
rect 270 6400 330 6460
rect 470 6400 530 6460
rect 660 6400 720 6460
rect 860 6400 920 6460
rect 1060 6400 1120 6460
rect 70 6235 130 6295
rect 270 6235 330 6295
rect 470 6235 530 6295
rect 660 6235 720 6295
rect 860 6235 920 6295
rect 1060 6235 1120 6295
rect 70 6035 130 6095
rect 270 6035 330 6095
rect 470 6035 530 6095
rect 660 6035 720 6095
rect 860 6035 920 6095
rect 1060 6035 1120 6095
rect 70 5845 130 5905
rect 270 5845 330 5905
rect 470 5845 530 5905
rect 660 5845 720 5905
rect 860 5845 920 5905
rect 1060 5845 1120 5905
rect 70 5665 130 5725
rect 270 5665 330 5725
rect 470 5665 530 5725
rect 660 5665 720 5725
rect 860 5665 920 5725
rect 1060 5665 1120 5725
rect 70 5465 130 5525
rect 270 5465 330 5525
rect 470 5465 530 5525
rect 660 5465 720 5525
rect 860 5465 920 5525
rect 1060 5465 1120 5525
rect 70 5275 130 5335
rect 270 5275 330 5335
rect 470 5275 530 5335
rect 660 5275 720 5335
rect 860 5275 920 5335
rect 1060 5275 1120 5335
rect 70 5115 130 5175
rect 270 5115 330 5175
rect 470 5115 530 5175
rect 660 5115 720 5175
rect 860 5115 920 5175
rect 1060 5115 1120 5175
rect 70 4925 130 4985
rect 270 4925 330 4985
rect 470 4925 530 4985
rect 660 4925 720 4985
rect 860 4925 920 4985
rect 1060 4925 1120 4985
rect 70 4750 130 4810
rect 270 4750 330 4810
rect 470 4750 530 4810
rect 660 4750 720 4810
rect 860 4750 920 4810
rect 1060 4750 1120 4810
rect 70 4610 130 4670
rect 270 4610 330 4670
rect 470 4610 530 4670
rect 660 4610 720 4670
rect 860 4610 920 4670
rect 1060 4610 1120 4670
<< metal2 >>
rect 80 6460 140 6470
rect 80 6390 140 6400
rect 270 6460 330 6470
rect 270 6390 330 6400
rect 470 6460 530 6470
rect 470 6390 530 6400
rect 660 6460 720 6470
rect 660 6390 720 6400
rect 860 6460 920 6470
rect 860 6390 920 6400
rect 1060 6460 1120 6470
rect 1060 6390 1120 6400
rect 70 6295 130 6305
rect 70 6225 130 6235
rect 270 6295 330 6305
rect 270 6225 330 6235
rect 470 6295 530 6305
rect 470 6225 530 6235
rect 660 6295 720 6305
rect 660 6225 720 6235
rect 860 6295 920 6305
rect 860 6225 920 6235
rect 1060 6295 1120 6305
rect 1060 6225 1120 6235
rect 70 6095 130 6105
rect 70 6025 130 6035
rect 270 6095 330 6105
rect 270 6025 330 6035
rect 470 6095 530 6105
rect 470 6025 530 6035
rect 660 6095 720 6105
rect 660 6025 720 6035
rect 860 6095 920 6105
rect 860 6025 920 6035
rect 1060 6095 1120 6105
rect 1060 6025 1120 6035
rect 70 5905 130 5915
rect 70 5835 130 5845
rect 270 5905 330 5915
rect 270 5835 330 5845
rect 470 5905 530 5915
rect 470 5835 530 5845
rect 660 5905 720 5915
rect 660 5835 720 5845
rect 860 5905 920 5915
rect 860 5835 920 5845
rect 1060 5905 1120 5915
rect 1060 5835 1120 5845
rect 70 5725 130 5735
rect 70 5655 130 5665
rect 270 5725 330 5735
rect 270 5655 330 5665
rect 470 5725 530 5735
rect 470 5655 530 5665
rect 660 5725 720 5735
rect 660 5655 720 5665
rect 860 5725 920 5735
rect 860 5655 920 5665
rect 1060 5725 1120 5735
rect 1060 5655 1120 5665
rect 70 5525 130 5535
rect 70 5455 130 5465
rect 270 5525 330 5535
rect 270 5455 330 5465
rect 470 5525 530 5535
rect 470 5455 530 5465
rect 660 5525 720 5535
rect 660 5455 720 5465
rect 860 5525 920 5535
rect 860 5455 920 5465
rect 1060 5525 1120 5535
rect 1060 5455 1120 5465
rect 70 5335 130 5345
rect 70 5265 130 5275
rect 270 5335 330 5345
rect 270 5265 330 5275
rect 470 5335 530 5345
rect 470 5265 530 5275
rect 660 5335 720 5345
rect 660 5265 720 5275
rect 860 5335 920 5345
rect 860 5265 920 5275
rect 1060 5335 1120 5345
rect 1060 5265 1120 5275
rect 70 5175 130 5185
rect 70 5105 130 5115
rect 270 5175 330 5185
rect 270 5105 330 5115
rect 470 5175 530 5185
rect 470 5105 530 5115
rect 660 5175 720 5185
rect 660 5105 720 5115
rect 860 5175 920 5185
rect 860 5105 920 5115
rect 1060 5175 1120 5185
rect 1060 5105 1120 5115
rect 70 4985 130 4995
rect 70 4915 130 4925
rect 270 4985 330 4995
rect 270 4915 330 4925
rect 470 4985 530 4995
rect 470 4915 530 4925
rect 660 4985 720 4995
rect 660 4915 720 4925
rect 860 4985 920 4995
rect 860 4915 920 4925
rect 1060 4985 1120 4995
rect 1060 4915 1120 4925
rect 70 4810 130 4820
rect 70 4740 130 4750
rect 270 4810 330 4820
rect 270 4740 330 4750
rect 470 4810 530 4820
rect 470 4740 530 4750
rect 660 4810 720 4820
rect 660 4740 720 4750
rect 860 4810 920 4820
rect 860 4740 920 4750
rect 1060 4810 1120 4820
rect 1060 4740 1120 4750
rect 70 4670 130 4680
rect 70 4600 130 4610
rect 270 4670 330 4680
rect 270 4600 330 4610
rect 470 4670 530 4680
rect 470 4600 530 4610
rect 660 4670 720 4680
rect 660 4600 720 4610
rect 860 4670 920 4680
rect 860 4600 920 4610
rect 1060 4670 1120 4680
rect 1060 4600 1120 4610
<< via2 >>
rect 80 6400 140 6460
rect 270 6400 330 6460
rect 470 6400 530 6460
rect 660 6400 720 6460
rect 860 6400 920 6460
rect 1060 6400 1120 6460
rect 70 6235 130 6295
rect 270 6235 330 6295
rect 470 6235 530 6295
rect 660 6235 720 6295
rect 860 6235 920 6295
rect 1060 6235 1120 6295
rect 70 6035 130 6095
rect 270 6035 330 6095
rect 470 6035 530 6095
rect 660 6035 720 6095
rect 860 6035 920 6095
rect 1060 6035 1120 6095
rect 70 5845 130 5905
rect 270 5845 330 5905
rect 470 5845 530 5905
rect 660 5845 720 5905
rect 860 5845 920 5905
rect 1060 5845 1120 5905
rect 70 5665 130 5725
rect 270 5665 330 5725
rect 470 5665 530 5725
rect 660 5665 720 5725
rect 860 5665 920 5725
rect 1060 5665 1120 5725
rect 70 5465 130 5525
rect 270 5465 330 5525
rect 470 5465 530 5525
rect 660 5465 720 5525
rect 860 5465 920 5525
rect 1060 5465 1120 5525
rect 70 5275 130 5335
rect 270 5275 330 5335
rect 470 5275 530 5335
rect 660 5275 720 5335
rect 860 5275 920 5335
rect 1060 5275 1120 5335
rect 70 5115 130 5175
rect 270 5115 330 5175
rect 470 5115 530 5175
rect 660 5115 720 5175
rect 860 5115 920 5175
rect 1060 5115 1120 5175
rect 70 4925 130 4985
rect 270 4925 330 4985
rect 470 4925 530 4985
rect 660 4925 720 4985
rect 860 4925 920 4985
rect 1060 4925 1120 4985
rect 70 4750 130 4810
rect 270 4750 330 4810
rect 470 4750 530 4810
rect 660 4750 720 4810
rect 860 4750 920 4810
rect 1060 4750 1120 4810
rect 70 4610 130 4670
rect 270 4610 330 4670
rect 470 4610 530 4670
rect 660 4610 720 4670
rect 860 4610 920 4670
rect 1060 4610 1120 4670
<< metal3 >>
rect 40 6460 1150 6490
rect 40 6400 80 6460
rect 140 6400 270 6460
rect 330 6400 470 6460
rect 530 6400 660 6460
rect 720 6400 860 6460
rect 920 6400 1060 6460
rect 1120 6400 1150 6460
rect 40 6295 1150 6400
rect 40 6235 70 6295
rect 130 6235 270 6295
rect 330 6235 470 6295
rect 530 6235 660 6295
rect 720 6235 860 6295
rect 920 6235 1060 6295
rect 1120 6235 1150 6295
rect 40 6095 1150 6235
rect 40 6035 70 6095
rect 130 6035 270 6095
rect 330 6035 470 6095
rect 530 6035 660 6095
rect 720 6035 860 6095
rect 920 6035 1060 6095
rect 1120 6035 1150 6095
rect 40 5905 1150 6035
rect 40 5845 70 5905
rect 130 5845 270 5905
rect 330 5845 470 5905
rect 530 5845 660 5905
rect 720 5845 860 5905
rect 920 5845 1060 5905
rect 1120 5845 1150 5905
rect 40 5725 1150 5845
rect 40 5665 70 5725
rect 130 5665 270 5725
rect 330 5665 470 5725
rect 530 5665 660 5725
rect 720 5665 860 5725
rect 920 5665 1060 5725
rect 1120 5665 1150 5725
rect 40 5525 1150 5665
rect 40 5465 70 5525
rect 130 5465 270 5525
rect 330 5465 470 5525
rect 530 5465 660 5525
rect 720 5465 860 5525
rect 920 5465 1060 5525
rect 1120 5465 1150 5525
rect 40 5335 1150 5465
rect 40 5275 70 5335
rect 130 5275 270 5335
rect 330 5275 470 5335
rect 530 5275 660 5335
rect 720 5275 860 5335
rect 920 5275 1060 5335
rect 1120 5275 1150 5335
rect 40 5175 1150 5275
rect 40 5115 70 5175
rect 130 5115 270 5175
rect 330 5115 470 5175
rect 530 5115 660 5175
rect 720 5115 860 5175
rect 920 5115 1060 5175
rect 1120 5115 1150 5175
rect 40 4985 1150 5115
rect 40 4925 70 4985
rect 130 4925 270 4985
rect 330 4925 470 4985
rect 530 4925 660 4985
rect 720 4925 860 4985
rect 920 4925 1060 4985
rect 1120 4925 1150 4985
rect 40 4810 1150 4925
rect 40 4750 70 4810
rect 130 4750 270 4810
rect 330 4750 470 4810
rect 530 4750 660 4810
rect 720 4750 860 4810
rect 920 4750 1060 4810
rect 1120 4750 1150 4810
rect 40 4670 1150 4750
rect 40 4610 70 4670
rect 130 4610 270 4670
rect 330 4610 470 4670
rect 530 4610 660 4670
rect 720 4610 860 4670
rect 920 4610 1060 4670
rect 1120 4610 1150 4670
rect 40 4560 1150 4610
use sky130_fd_pr__nfet_01v8_UXPKRJ  sky130_fd_pr__nfet_01v8_UXPKRJ_0
timestamp 1717119771
transform 1 0 597 0 1 5150
box -657 -5210 657 5210
<< end >>
