magic
tech sky130A
magscale 1 2
timestamp 1716868724
<< metal3 >>
rect -1750 1672 1749 1700
rect -1750 1608 1665 1672
rect 1729 1608 1749 1672
rect -1750 1592 1749 1608
rect -1750 1528 1665 1592
rect 1729 1528 1749 1592
rect -1750 1512 1749 1528
rect -1750 1448 1665 1512
rect 1729 1448 1749 1512
rect -1750 1432 1749 1448
rect -1750 1368 1665 1432
rect 1729 1368 1749 1432
rect -1750 1352 1749 1368
rect -1750 1288 1665 1352
rect 1729 1288 1749 1352
rect -1750 1272 1749 1288
rect -1750 1208 1665 1272
rect 1729 1208 1749 1272
rect -1750 1192 1749 1208
rect -1750 1128 1665 1192
rect 1729 1128 1749 1192
rect -1750 1112 1749 1128
rect -1750 1048 1665 1112
rect 1729 1048 1749 1112
rect -1750 1032 1749 1048
rect -1750 968 1665 1032
rect 1729 968 1749 1032
rect -1750 952 1749 968
rect -1750 888 1665 952
rect 1729 888 1749 952
rect -1750 872 1749 888
rect -1750 808 1665 872
rect 1729 808 1749 872
rect -1750 792 1749 808
rect -1750 728 1665 792
rect 1729 728 1749 792
rect -1750 712 1749 728
rect -1750 648 1665 712
rect 1729 648 1749 712
rect -1750 632 1749 648
rect -1750 568 1665 632
rect 1729 568 1749 632
rect -1750 552 1749 568
rect -1750 488 1665 552
rect 1729 488 1749 552
rect -1750 472 1749 488
rect -1750 408 1665 472
rect 1729 408 1749 472
rect -1750 392 1749 408
rect -1750 328 1665 392
rect 1729 328 1749 392
rect -1750 312 1749 328
rect -1750 248 1665 312
rect 1729 248 1749 312
rect -1750 232 1749 248
rect -1750 168 1665 232
rect 1729 168 1749 232
rect -1750 152 1749 168
rect -1750 88 1665 152
rect 1729 88 1749 152
rect -1750 72 1749 88
rect -1750 8 1665 72
rect 1729 8 1749 72
rect -1750 -8 1749 8
rect -1750 -72 1665 -8
rect 1729 -72 1749 -8
rect -1750 -88 1749 -72
rect -1750 -152 1665 -88
rect 1729 -152 1749 -88
rect -1750 -168 1749 -152
rect -1750 -232 1665 -168
rect 1729 -232 1749 -168
rect -1750 -248 1749 -232
rect -1750 -312 1665 -248
rect 1729 -312 1749 -248
rect -1750 -328 1749 -312
rect -1750 -392 1665 -328
rect 1729 -392 1749 -328
rect -1750 -408 1749 -392
rect -1750 -472 1665 -408
rect 1729 -472 1749 -408
rect -1750 -488 1749 -472
rect -1750 -552 1665 -488
rect 1729 -552 1749 -488
rect -1750 -568 1749 -552
rect -1750 -632 1665 -568
rect 1729 -632 1749 -568
rect -1750 -648 1749 -632
rect -1750 -712 1665 -648
rect 1729 -712 1749 -648
rect -1750 -728 1749 -712
rect -1750 -792 1665 -728
rect 1729 -792 1749 -728
rect -1750 -808 1749 -792
rect -1750 -872 1665 -808
rect 1729 -872 1749 -808
rect -1750 -888 1749 -872
rect -1750 -952 1665 -888
rect 1729 -952 1749 -888
rect -1750 -968 1749 -952
rect -1750 -1032 1665 -968
rect 1729 -1032 1749 -968
rect -1750 -1048 1749 -1032
rect -1750 -1112 1665 -1048
rect 1729 -1112 1749 -1048
rect -1750 -1128 1749 -1112
rect -1750 -1192 1665 -1128
rect 1729 -1192 1749 -1128
rect -1750 -1208 1749 -1192
rect -1750 -1272 1665 -1208
rect 1729 -1272 1749 -1208
rect -1750 -1288 1749 -1272
rect -1750 -1352 1665 -1288
rect 1729 -1352 1749 -1288
rect -1750 -1368 1749 -1352
rect -1750 -1432 1665 -1368
rect 1729 -1432 1749 -1368
rect -1750 -1448 1749 -1432
rect -1750 -1512 1665 -1448
rect 1729 -1512 1749 -1448
rect -1750 -1528 1749 -1512
rect -1750 -1592 1665 -1528
rect 1729 -1592 1749 -1528
rect -1750 -1608 1749 -1592
rect -1750 -1672 1665 -1608
rect 1729 -1672 1749 -1608
rect -1750 -1700 1749 -1672
<< via3 >>
rect 1665 1608 1729 1672
rect 1665 1528 1729 1592
rect 1665 1448 1729 1512
rect 1665 1368 1729 1432
rect 1665 1288 1729 1352
rect 1665 1208 1729 1272
rect 1665 1128 1729 1192
rect 1665 1048 1729 1112
rect 1665 968 1729 1032
rect 1665 888 1729 952
rect 1665 808 1729 872
rect 1665 728 1729 792
rect 1665 648 1729 712
rect 1665 568 1729 632
rect 1665 488 1729 552
rect 1665 408 1729 472
rect 1665 328 1729 392
rect 1665 248 1729 312
rect 1665 168 1729 232
rect 1665 88 1729 152
rect 1665 8 1729 72
rect 1665 -72 1729 -8
rect 1665 -152 1729 -88
rect 1665 -232 1729 -168
rect 1665 -312 1729 -248
rect 1665 -392 1729 -328
rect 1665 -472 1729 -408
rect 1665 -552 1729 -488
rect 1665 -632 1729 -568
rect 1665 -712 1729 -648
rect 1665 -792 1729 -728
rect 1665 -872 1729 -808
rect 1665 -952 1729 -888
rect 1665 -1032 1729 -968
rect 1665 -1112 1729 -1048
rect 1665 -1192 1729 -1128
rect 1665 -1272 1729 -1208
rect 1665 -1352 1729 -1288
rect 1665 -1432 1729 -1368
rect 1665 -1512 1729 -1448
rect 1665 -1592 1729 -1528
rect 1665 -1672 1729 -1608
<< mimcap >>
rect -1650 1552 1550 1600
rect -1650 -1552 -1602 1552
rect 1502 -1552 1550 1552
rect -1650 -1600 1550 -1552
<< mimcapcontact >>
rect -1602 -1552 1502 1552
<< metal4 >>
rect 1649 1672 1745 1688
rect 1649 1608 1665 1672
rect 1729 1608 1745 1672
rect 1649 1592 1745 1608
rect -1611 1552 1511 1561
rect -1611 -1552 -1602 1552
rect 1502 -1552 1511 1552
rect -1611 -1561 1511 -1552
rect 1649 1528 1665 1592
rect 1729 1528 1745 1592
rect 1649 1512 1745 1528
rect 1649 1448 1665 1512
rect 1729 1448 1745 1512
rect 1649 1432 1745 1448
rect 1649 1368 1665 1432
rect 1729 1368 1745 1432
rect 1649 1352 1745 1368
rect 1649 1288 1665 1352
rect 1729 1288 1745 1352
rect 1649 1272 1745 1288
rect 1649 1208 1665 1272
rect 1729 1208 1745 1272
rect 1649 1192 1745 1208
rect 1649 1128 1665 1192
rect 1729 1128 1745 1192
rect 1649 1112 1745 1128
rect 1649 1048 1665 1112
rect 1729 1048 1745 1112
rect 1649 1032 1745 1048
rect 1649 968 1665 1032
rect 1729 968 1745 1032
rect 1649 952 1745 968
rect 1649 888 1665 952
rect 1729 888 1745 952
rect 1649 872 1745 888
rect 1649 808 1665 872
rect 1729 808 1745 872
rect 1649 792 1745 808
rect 1649 728 1665 792
rect 1729 728 1745 792
rect 1649 712 1745 728
rect 1649 648 1665 712
rect 1729 648 1745 712
rect 1649 632 1745 648
rect 1649 568 1665 632
rect 1729 568 1745 632
rect 1649 552 1745 568
rect 1649 488 1665 552
rect 1729 488 1745 552
rect 1649 472 1745 488
rect 1649 408 1665 472
rect 1729 408 1745 472
rect 1649 392 1745 408
rect 1649 328 1665 392
rect 1729 328 1745 392
rect 1649 312 1745 328
rect 1649 248 1665 312
rect 1729 248 1745 312
rect 1649 232 1745 248
rect 1649 168 1665 232
rect 1729 168 1745 232
rect 1649 152 1745 168
rect 1649 88 1665 152
rect 1729 88 1745 152
rect 1649 72 1745 88
rect 1649 8 1665 72
rect 1729 8 1745 72
rect 1649 -8 1745 8
rect 1649 -72 1665 -8
rect 1729 -72 1745 -8
rect 1649 -88 1745 -72
rect 1649 -152 1665 -88
rect 1729 -152 1745 -88
rect 1649 -168 1745 -152
rect 1649 -232 1665 -168
rect 1729 -232 1745 -168
rect 1649 -248 1745 -232
rect 1649 -312 1665 -248
rect 1729 -312 1745 -248
rect 1649 -328 1745 -312
rect 1649 -392 1665 -328
rect 1729 -392 1745 -328
rect 1649 -408 1745 -392
rect 1649 -472 1665 -408
rect 1729 -472 1745 -408
rect 1649 -488 1745 -472
rect 1649 -552 1665 -488
rect 1729 -552 1745 -488
rect 1649 -568 1745 -552
rect 1649 -632 1665 -568
rect 1729 -632 1745 -568
rect 1649 -648 1745 -632
rect 1649 -712 1665 -648
rect 1729 -712 1745 -648
rect 1649 -728 1745 -712
rect 1649 -792 1665 -728
rect 1729 -792 1745 -728
rect 1649 -808 1745 -792
rect 1649 -872 1665 -808
rect 1729 -872 1745 -808
rect 1649 -888 1745 -872
rect 1649 -952 1665 -888
rect 1729 -952 1745 -888
rect 1649 -968 1745 -952
rect 1649 -1032 1665 -968
rect 1729 -1032 1745 -968
rect 1649 -1048 1745 -1032
rect 1649 -1112 1665 -1048
rect 1729 -1112 1745 -1048
rect 1649 -1128 1745 -1112
rect 1649 -1192 1665 -1128
rect 1729 -1192 1745 -1128
rect 1649 -1208 1745 -1192
rect 1649 -1272 1665 -1208
rect 1729 -1272 1745 -1208
rect 1649 -1288 1745 -1272
rect 1649 -1352 1665 -1288
rect 1729 -1352 1745 -1288
rect 1649 -1368 1745 -1352
rect 1649 -1432 1665 -1368
rect 1729 -1432 1745 -1368
rect 1649 -1448 1745 -1432
rect 1649 -1512 1665 -1448
rect 1729 -1512 1745 -1448
rect 1649 -1528 1745 -1512
rect 1649 -1592 1665 -1528
rect 1729 -1592 1745 -1528
rect 1649 -1608 1745 -1592
rect 1649 -1672 1665 -1608
rect 1729 -1672 1745 -1608
rect 1649 -1688 1745 -1672
<< properties >>
string FIXED_BBOX -1750 -1700 1650 1700
<< end >>
