** sch_path: /foss/designs/Analog_FA23_SP24/PTAT/xschem/PTAT_v0p0p0.sch
.subckt PTAT_v0p0p0 VDD VOUT VSS
*.PININFO VSS:I VDD:I VOUT:O
XM1 net1 net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt L=1 W=19 nf=1 m=1
XM2 net2 net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt L=1 W=19 nf=1 m=1
XM3 VOUT net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt L=1 W=19 nf=1 m=1
XM4 net1 net1 VSS VSS sky130_fd_pr__nfet_01v8_lvt L=0.6 W=4 nf=1 m=1
XM5 net2 net1 net3 VSS sky130_fd_pr__nfet_01v8_lvt L=0.6 W=4 nf=1 m=20
XM6 net2 net2 net1 VSS sky130_fd_pr__nfet_01v8_lvt L=0.15 W=0.42 nf=1 m=1
XM7 VOUT VOUT VSS VSS sky130_fd_pr__nfet_01v8_lvt L=0.6 W=4 nf=1 m=1
XR1 VSS net3 VSS sky130_fd_pr__res_xhigh_po_5p73 L=85.94 mult=1 m=1
XR2 VSS net3 VSS sky130_fd_pr__res_xhigh_po_5p73 L=85.94 mult=1 m=1
.ends
.end
