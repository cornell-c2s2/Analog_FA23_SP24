magic
tech sky130A
magscale 1 2
timestamp 1709395973
<< pwell >>
rect 3450 -2700 4650 -2600
<< metal1 >>
rect 0 0 200 200
rect 2500 -50 3450 50
rect 3550 -50 4500 50
rect 4800 -50 6800 50
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
rect 2650 -1250 6700 -1150
rect 0 -1600 200 -1400
rect 3450 -1500 5850 -1400
rect 0 -2000 200 -1800
rect 3440 -2700 3450 -2600
rect 3550 -2700 4600 -2600
rect 4700 -2700 5850 -2600
<< via1 >>
rect 3450 -50 3550 50
rect 3450 -2700 3550 -2600
<< metal2 >>
rect 3450 50 3550 60
rect 3450 -2600 3550 -50
rect 3450 -2710 3550 -2700
use sky130_fd_pr__pfet_01v8_BDZ9JN  XM1
timestamp 1709390584
transform 1 0 3579 0 1 -581
box -1079 -719 1079 719
use sky130_fd_pr__nfet_01v8_KBNS5F  XM2
timestamp 1709392794
transform 1 0 4049 0 1 -2040
box -599 -710 599 710
use sky130_fd_pr__pfet_01v8_BDZ9JN  XM3
timestamp 1709390584
transform 1 0 5729 0 1 -581
box -1079 -719 1079 719
use sky130_fd_pr__nfet_01v8_KBNS5F  XM4
timestamp 1709392794
transform 1 0 5249 0 1 -2040
box -599 -710 599 710
use sky130_fd_pr__nfet_01v8_MMMA4V  XM5
timestamp 1709390584
transform 1 0 1896 0 1 -2040
box -296 -710 296 710
use sky130_fd_pr__pfet_01v8_3HZ9VM  XM8
timestamp 1709390584
transform 1 0 1921 0 1 -581
box -296 -719 296 719
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 VREF_P
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 VDD
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 OUT
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 VIN
port 3 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 256 0 0 0 VSS
port 4 nsew
flabel metal1 0 -2000 200 -1800 0 FreeSans 256 0 0 0 VREF_N
port 5 nsew
<< end >>
