magic
tech sky130A
timestamp 1714085375
<< pwell >>
rect -128 -126 128 126
<< nmos >>
rect -30 -21 30 21
<< ndiff >>
rect -59 15 -30 21
rect -59 -15 -53 15
rect -36 -15 -30 15
rect -59 -21 -30 -15
rect 30 15 59 21
rect 30 -15 36 15
rect 53 -15 59 15
rect 30 -21 59 -15
<< ndiffc >>
rect -53 -15 -36 15
rect 36 -15 53 15
<< psubdiff >>
rect -110 91 -62 108
rect 62 91 110 108
rect -110 60 -93 91
rect 93 60 110 91
rect -110 -91 -93 -60
rect 93 -91 110 -60
rect -110 -108 -62 -91
rect 62 -108 110 -91
<< psubdiffcont >>
rect -62 91 62 108
rect -110 -60 -93 60
rect 93 -60 110 60
rect -62 -108 62 -91
<< poly >>
rect -30 57 30 65
rect -30 40 -22 57
rect 22 40 30 57
rect -30 21 30 40
rect -30 -40 30 -21
rect -30 -57 -22 -40
rect 22 -57 30 -40
rect -30 -65 30 -57
<< polycont >>
rect -22 40 22 57
rect -22 -57 22 -40
<< locali >>
rect -110 91 -62 108
rect 62 91 110 108
rect -110 60 -93 91
rect 93 60 110 91
rect -30 40 -22 57
rect 22 40 30 57
rect -53 15 -36 23
rect -53 -23 -36 -15
rect 36 15 53 23
rect 36 -23 53 -15
rect -30 -57 -22 -40
rect 22 -57 30 -40
rect -110 -91 -93 -60
rect 93 -91 110 -60
rect -110 -108 -62 -91
rect 62 -108 110 -91
<< viali >>
rect -22 40 22 57
rect -53 -15 -36 15
rect 36 -15 53 15
rect -22 -57 22 -40
<< metal1 >>
rect -28 57 28 60
rect -28 40 -22 57
rect 22 40 28 57
rect -28 37 28 40
rect -56 15 -33 21
rect -56 -15 -53 15
rect -36 -15 -33 15
rect -56 -21 -33 -15
rect 33 15 56 21
rect 33 -15 36 15
rect 53 -15 56 15
rect 33 -21 56 -15
rect -28 -40 28 -37
rect -28 -57 -22 -40
rect 22 -57 28 -40
rect -28 -60 28 -57
<< properties >>
string FIXED_BBOX -101 -99 101 99
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.42 l 0.6 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
