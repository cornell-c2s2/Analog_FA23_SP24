** sch_path: /foss/designs/Analog_FA23_SP24/ComparatorLayout/class_AB_v2_sym.sch
.subckt class_AB_v2_sym VDD IB VSS VIP VIN VON VOP CLK
*.PININFO VDD:B IB:I VSS:B VIP:I VIN:I VON:O VOP:O CLK:I
XM17 net3 VIP VIR VSS sky130_fd_pr__nfet_01v8_lvt L=0.6 W=4 nf=1 m=1
XM12 IB IB VSS VSS sky130_fd_pr__nfet_01v8_lvt L=0.6 W=4 nf=1 m=1
XM15 net2 VIN VIR VSS sky130_fd_pr__nfet_01v8_lvt L=0.6 W=4 nf=1 m=1
XM13 VIR IB VSS VSS sky130_fd_pr__nfet_01v8_lvt L=0.6 W=4 nf=1 m=2
XM6 VON VOP VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4 nf=1 m=1
XM7 VOP VON VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4 nf=1 m=1
XM10 VOP VON net1 VSS sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 nf=1 m=1
XM11 VON VOP net1 VSS sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 nf=1 m=1
XM1 net1 CLK VSS VSS sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 nf=1 m=1
XM2 VOP CLK VON VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4 nf=1 m=1
XM5 net2 VIP net2 net2 sky130_fd_pr__nfet_01v8_lvt L=0.15 W=2 nf=1 m=1
XM8 net3 VIN net3 net3 sky130_fd_pr__nfet_01v8_lvt L=0.15 W=2 nf=1 m=1
XM9 net2 CLK VOP VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4 nf=1 m=1
XM14 net3 CLK VON VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=4 nf=1 m=1
XM3 VDD CLK net3 VSS sky130_fd_pr__nfet_01v8_lvt L=0.6 W=4 nf=1 m=1
XM4 VDD CLK net2 VSS sky130_fd_pr__nfet_01v8_lvt L=0.6 W=4 nf=1 m=1
.ends
.end
