magic
tech sky130A
magscale 1 2
timestamp 1716868724
<< pwell >>
rect -3223 -6312 3223 6312
<< psubdiff >>
rect -3187 6242 -3091 6276
rect 3091 6242 3187 6276
rect -3187 6180 -3153 6242
rect 3153 6180 3187 6242
rect -3187 -6242 -3153 -6180
rect 3153 -6242 3187 -6180
rect -3187 -6276 -3091 -6242
rect 3091 -6276 3187 -6242
<< psubdiffcont >>
rect -3091 6242 3091 6276
rect -3187 -6180 -3153 6180
rect 3153 -6180 3187 6180
rect -3091 -6276 3091 -6242
<< xpolycontact >>
rect -3057 5714 -1911 6146
rect -3057 -6146 -1911 -5714
rect -1815 5714 -669 6146
rect -1815 -6146 -669 -5714
rect -573 5714 573 6146
rect -573 -6146 573 -5714
rect 669 5714 1815 6146
rect 669 -6146 1815 -5714
rect 1911 5714 3057 6146
rect 1911 -6146 3057 -5714
<< xpolyres >>
rect -3057 -5714 -1911 5714
rect -1815 -5714 -669 5714
rect -573 -5714 573 5714
rect 669 -5714 1815 5714
rect 1911 -5714 3057 5714
<< locali >>
rect -3187 6242 -3091 6276
rect 3091 6242 3187 6276
rect -3187 6180 -3153 6242
rect 3153 6180 3187 6242
rect -3187 -6242 -3153 -6180
rect 3153 -6242 3187 -6180
rect -3187 -6276 -3091 -6242
rect 3091 -6276 3187 -6242
<< viali >>
rect -3041 5731 -1927 6128
rect -1799 5731 -685 6128
rect -557 5731 557 6128
rect 685 5731 1799 6128
rect 1927 5731 3041 6128
rect -3041 -6128 -1927 -5731
rect -1799 -6128 -685 -5731
rect -557 -6128 557 -5731
rect 685 -6128 1799 -5731
rect 1927 -6128 3041 -5731
<< metal1 >>
rect -3053 6128 -1915 6134
rect -3053 5731 -3041 6128
rect -1927 5731 -1915 6128
rect -3053 5725 -1915 5731
rect -1811 6128 -673 6134
rect -1811 5731 -1799 6128
rect -685 5731 -673 6128
rect -1811 5725 -673 5731
rect -569 6128 569 6134
rect -569 5731 -557 6128
rect 557 5731 569 6128
rect -569 5725 569 5731
rect 673 6128 1811 6134
rect 673 5731 685 6128
rect 1799 5731 1811 6128
rect 673 5725 1811 5731
rect 1915 6128 3053 6134
rect 1915 5731 1927 6128
rect 3041 5731 3053 6128
rect 1915 5725 3053 5731
rect -3053 -5731 -1915 -5725
rect -3053 -6128 -3041 -5731
rect -1927 -6128 -1915 -5731
rect -3053 -6134 -1915 -6128
rect -1811 -5731 -673 -5725
rect -1811 -6128 -1799 -5731
rect -685 -6128 -673 -5731
rect -1811 -6134 -673 -6128
rect -569 -5731 569 -5725
rect -569 -6128 -557 -5731
rect 557 -6128 569 -5731
rect -569 -6134 569 -6128
rect 673 -5731 1811 -5725
rect 673 -6128 685 -5731
rect 1799 -6128 1811 -5731
rect 673 -6134 1811 -6128
rect 1915 -5731 3053 -5725
rect 1915 -6128 1927 -5731
rect 3041 -6128 3053 -5731
rect 1915 -6134 3053 -6128
<< properties >>
string FIXED_BBOX -3170 -6259 3170 6259
string gencell sky130_fd_pr__res_xhigh_po_5p73
string library sky130
string parameters w 5.73 l 57.3 m 1 nx 5 wmin 5.730 lmin 0.50 rho 2000 val 20.065k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 5.730 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
