magic
tech sky130A
magscale 1 2
timestamp 1712038425
<< error_s >>
rect 2404 -346 2462 -340
rect 2404 -380 2416 -346
rect 2404 -386 2462 -380
rect 772 -417 818 -405
rect 1300 -417 1346 -405
rect 1504 -417 1550 -405
rect 2032 -417 2078 -405
rect 772 -451 778 -417
rect 1300 -451 1306 -417
rect 1504 -451 1510 -417
rect 2032 -451 2038 -417
rect 772 -463 818 -451
rect 1300 -463 1346 -451
rect 1504 -463 1550 -451
rect 2032 -463 2078 -451
rect 992 -862 1038 -850
rect 1302 -862 1348 -850
rect 1506 -862 1552 -850
rect 1816 -862 1862 -850
rect 992 -896 998 -862
rect 1302 -896 1308 -862
rect 1506 -896 1512 -862
rect 1816 -896 1822 -862
rect 2296 -874 2354 -868
rect 992 -908 1038 -896
rect 1302 -908 1348 -896
rect 1506 -908 1552 -896
rect 1816 -908 1862 -896
rect 2296 -908 2308 -874
rect 2296 -914 2354 -908
rect 992 -1178 1038 -1166
rect 1302 -1178 1348 -1166
rect 1506 -1178 1552 -1166
rect 1816 -1178 1862 -1166
rect 716 -1188 774 -1182
rect 716 -1222 728 -1188
rect 992 -1212 998 -1178
rect 1302 -1212 1308 -1178
rect 1506 -1212 1512 -1178
rect 1816 -1212 1822 -1178
rect 2082 -1188 2140 -1182
rect 716 -1228 774 -1222
rect 992 -1224 1038 -1212
rect 1302 -1224 1348 -1212
rect 1506 -1224 1552 -1212
rect 1816 -1224 1862 -1212
rect 2082 -1222 2094 -1188
rect 2082 -1228 2140 -1222
rect 716 -1698 774 -1692
rect 2082 -1698 2140 -1692
rect 716 -1732 728 -1698
rect 2082 -1732 2094 -1698
rect 716 -1738 774 -1732
rect 2082 -1738 2140 -1732
<< nwell >>
rect 350 -300 600 -210
rect 380 -410 390 -330
rect 370 -420 390 -410
rect 380 -870 390 -420
rect 450 -870 470 -850
rect 490 -870 560 -330
rect 380 -920 560 -870
rect 380 -930 390 -920
rect 450 -930 470 -920
<< locali >>
rect 310 -280 640 -240
<< viali >>
rect 860 -280 1990 -240
rect 2210 -280 2600 -240
rect 330 -1010 620 -970
rect 2230 -1020 2530 -970
<< metal1 >>
rect -1000 0 -800 200
rect -1000 -400 -800 -200
rect 770 -220 2620 -210
rect 770 -240 2530 -220
rect 770 -280 860 -240
rect 1990 -280 2160 -240
rect 770 -300 2160 -280
rect 2230 -300 2530 -280
rect 2600 -300 2620 -220
rect 380 -320 460 -310
rect 380 -380 390 -320
rect 450 -380 460 -320
rect 380 -390 460 -380
rect 490 -390 500 -330
rect 560 -390 570 -330
rect 850 -350 2000 -300
rect 850 -390 1270 -350
rect 860 -400 1270 -390
rect 1580 -400 2000 -350
rect 260 -530 380 -420
rect 260 -590 270 -530
rect 330 -590 380 -530
rect 570 -530 700 -430
rect 570 -590 620 -530
rect 680 -590 700 -530
rect -1000 -800 -800 -600
rect 260 -640 380 -590
rect 260 -700 270 -640
rect 330 -700 380 -640
rect 420 -600 500 -590
rect 420 -660 430 -600
rect 490 -660 500 -600
rect 420 -670 500 -660
rect 570 -650 700 -590
rect 260 -750 380 -700
rect 260 -810 270 -750
rect 330 -810 380 -750
rect 260 -830 380 -810
rect 570 -710 620 -650
rect 680 -710 700 -650
rect 570 -750 700 -710
rect 570 -810 620 -750
rect 680 -810 700 -750
rect 570 -820 700 -810
rect 2140 -460 2280 -430
rect 2140 -540 2160 -460
rect 2230 -540 2280 -460
rect 2140 -590 2280 -540
rect 2140 -670 2160 -590
rect 2230 -670 2280 -590
rect 2140 -710 2280 -670
rect 2140 -790 2160 -710
rect 2230 -790 2280 -710
rect 2140 -820 2280 -790
rect 2480 -460 2620 -430
rect 2480 -540 2530 -460
rect 2600 -540 2620 -460
rect 2480 -590 2620 -540
rect 2480 -670 2530 -590
rect 2600 -670 2620 -590
rect 2480 -710 2620 -670
rect 2480 -790 2530 -710
rect 2600 -790 2620 -710
rect 2480 -820 2620 -790
rect 600 -830 700 -820
rect 2510 -830 2620 -820
rect 380 -920 390 -860
rect 450 -920 460 -860
rect 380 -930 460 -920
rect 500 -920 510 -860
rect 570 -920 580 -860
rect 500 -930 580 -920
rect 230 -950 340 -940
rect -1000 -1200 -800 -1000
rect 230 -1010 270 -950
rect 330 -960 340 -950
rect 610 -960 630 -950
rect 330 -970 630 -960
rect 620 -1010 630 -970
rect 690 -1010 710 -950
rect 230 -1020 710 -1010
rect 2140 -1020 2160 -960
rect 2220 -970 2540 -960
rect 2220 -1020 2230 -970
rect 2530 -1020 2540 -970
rect 2600 -1020 2620 -960
rect 2140 -1030 2620 -1020
rect -1000 -1600 -800 -1400
rect -1000 -2000 -800 -1800
rect 1220 -2130 1700 -1950
<< via1 >>
rect 2530 -240 2600 -220
rect 2160 -280 2210 -240
rect 2210 -280 2230 -240
rect 2530 -280 2600 -240
rect 2160 -300 2230 -280
rect 2530 -300 2600 -280
rect 390 -380 450 -320
rect 500 -390 560 -330
rect 270 -590 330 -530
rect 620 -590 680 -530
rect 270 -700 330 -640
rect 430 -660 490 -600
rect 270 -810 330 -750
rect 620 -710 680 -650
rect 620 -810 680 -750
rect 2160 -540 2230 -460
rect 2160 -670 2230 -590
rect 2160 -790 2230 -710
rect 2530 -540 2600 -460
rect 2530 -670 2600 -590
rect 2530 -790 2600 -710
rect 390 -920 450 -860
rect 510 -920 570 -860
rect 270 -1010 330 -950
rect 630 -1010 690 -950
rect 2160 -1020 2220 -960
rect 2540 -1020 2600 -960
<< metal2 >>
rect 250 -530 340 -140
rect 370 -320 460 -310
rect 370 -380 390 -320
rect 450 -380 460 -320
rect 370 -390 460 -380
rect 490 -320 570 -310
rect 490 -390 500 -320
rect 560 -390 570 -320
rect 500 -400 560 -390
rect 250 -590 270 -530
rect 330 -590 340 -530
rect 250 -640 340 -590
rect 250 -700 270 -640
rect 330 -700 340 -640
rect 420 -600 490 -590
rect 420 -660 430 -600
rect 420 -670 490 -660
rect 250 -750 340 -700
rect 250 -810 270 -750
rect 330 -810 340 -750
rect 250 -950 340 -810
rect 520 -850 560 -400
rect 610 -530 700 -140
rect 610 -590 620 -530
rect 680 -590 700 -530
rect 610 -650 700 -590
rect 610 -710 620 -650
rect 680 -710 700 -650
rect 610 -750 700 -710
rect 610 -810 620 -750
rect 680 -810 700 -750
rect 380 -860 470 -850
rect 380 -920 390 -860
rect 450 -920 470 -860
rect 380 -930 470 -920
rect 500 -860 580 -850
rect 500 -920 510 -860
rect 570 -920 580 -860
rect 500 -930 580 -920
rect 250 -960 270 -950
rect 230 -1010 270 -960
rect 330 -960 340 -950
rect 610 -950 700 -810
rect 610 -960 630 -950
rect 330 -1010 630 -960
rect 690 -960 700 -950
rect 2150 -240 2240 -140
rect 2150 -300 2160 -240
rect 2230 -300 2240 -240
rect 2150 -460 2240 -300
rect 2150 -540 2160 -460
rect 2230 -540 2240 -460
rect 2150 -590 2240 -540
rect 2150 -670 2160 -590
rect 2230 -670 2240 -590
rect 2150 -710 2240 -670
rect 2150 -790 2160 -710
rect 2230 -790 2240 -710
rect 2150 -960 2240 -790
rect 2520 -220 2610 -140
rect 2520 -300 2530 -220
rect 2600 -300 2610 -220
rect 2520 -460 2610 -300
rect 2520 -540 2530 -460
rect 2600 -540 2610 -460
rect 2520 -590 2610 -540
rect 2520 -670 2530 -590
rect 2600 -670 2610 -590
rect 2520 -710 2610 -670
rect 2520 -790 2530 -710
rect 2600 -790 2610 -710
rect 2520 -960 2610 -790
rect 690 -1010 710 -960
rect 230 -1020 710 -1010
rect 2140 -1020 2160 -960
rect 2220 -1020 2540 -960
rect 2600 -1020 2620 -960
rect 2140 -1030 2620 -1020
<< via2 >>
rect 390 -380 450 -320
rect 500 -330 560 -320
rect 500 -380 560 -330
rect 430 -660 490 -600
rect 390 -920 450 -860
rect 510 -920 570 -860
<< metal3 >>
rect -50 -320 570 -310
rect -50 -380 390 -320
rect 450 -380 500 -320
rect 560 -380 570 -320
rect -50 -400 570 -380
rect -60 -600 510 -580
rect -60 -660 430 -600
rect 490 -660 510 -600
rect -60 -680 510 -660
rect -60 -860 580 -850
rect -60 -920 390 -860
rect 450 -920 510 -860
rect 570 -920 580 -860
rect -60 -930 580 -920
use sky130_fd_sc_hd__inv_4  x1 pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 1228 0 -1 -1458
box -38 -48 498 592
use sky130_fd_sc_hd__inv_4  x2
timestamp 1701704242
transform 1 0 1228 0 1 -2622
box -38 -48 498 592
use sky130_fd_pr__nfet_01v8_648S5X  XM1
timestamp 1712020331
transform 0 1 1170 -1 0 -879
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_648S5X  XM2
timestamp 1712020331
transform 0 1 1170 -1 0 -1195
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_648S5X  XM3
timestamp 1712020331
transform 0 1 1684 -1 0 -879
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_648S5X  XM4
timestamp 1712020331
transform 0 1 1684 -1 0 -1195
box -211 -310 211 310
use sky130_fd_pr__pfet_01v8_6QB8WZ  XM5
timestamp 1712020331
transform 0 1 1059 -1 0 -434
box -226 -419 226 419
use sky130_fd_pr__pfet_01v8_6QB8WZ  XM6
timestamp 1712020331
transform 0 1 1791 -1 0 -434
box -226 -419 226 419
use sky130_fd_pr__pfet_01v8_E3L9V7  XM7
timestamp 1712036258
transform 1 0 472 0 1 -627
box -275 -419 275 419
use sky130_fd_pr__pfet_01v8_EDASV7  XM8
timestamp 1712022236
transform 1 0 2379 0 1 -627
box -275 -419 275 419
use sky130_fd_pr__nfet_01v8_4WSMTB  XM9
timestamp 1712022658
transform 1 0 745 0 1 -1460
box -221 -410 221 410
use sky130_fd_pr__nfet_01v8_XJSMYS  XM10
timestamp 1712022658
transform 1 0 2111 0 1 -1460
box -221 -410 221 410
<< labels >>
flabel metal1 -1000 0 -800 200 0 FreeSans 256 0 0 0 VDD
port 0 nsew
flabel metal1 -1000 -400 -800 -200 0 FreeSans 256 0 0 0 !S
port 1 nsew
flabel metal1 -1000 -800 -800 -600 0 FreeSans 256 0 0 0 !R
port 2 nsew
flabel metal1 -1000 -1600 -800 -1400 0 FreeSans 256 0 0 0 Q
port 4 nsew
flabel metal1 -1000 -2000 -800 -1800 0 FreeSans 256 0 0 0 GND
port 5 nsew
flabel metal1 -1000 -1200 -800 -1000 0 FreeSans 256 0 0 0 !Q
port 3 nsew
<< end >>
