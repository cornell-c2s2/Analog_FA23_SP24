magic
tech sky130A
magscale 1 2
timestamp 1713142632
<< pwell >>
rect -3223 -5970 3223 5970
<< psubdiff >>
rect -3187 5900 -3091 5934
rect 3091 5900 3187 5934
rect -3187 5838 -3153 5900
rect 3153 5838 3187 5900
rect -3187 -5900 -3153 -5838
rect 3153 -5900 3187 -5838
rect -3187 -5934 -3091 -5900
rect 3091 -5934 3187 -5900
<< psubdiffcont >>
rect -3091 5900 3091 5934
rect -3187 -5838 -3153 5838
rect 3153 -5838 3187 5838
rect -3091 -5934 3091 -5900
<< xpolycontact >>
rect 1911 5372 3057 5804
rect -3057 -5804 -1911 -5372
<< xpolyres >>
rect -3057 4122 -669 5268
rect -3057 -5372 -1911 4122
rect -1815 -4122 -669 4122
rect -573 4122 1815 5268
rect -573 -4122 573 4122
rect -1815 -5268 573 -4122
rect 669 -4122 1815 4122
rect 1911 -4122 3057 5372
rect 669 -5268 3057 -4122
<< locali >>
rect -3187 5900 -3091 5934
rect 3091 5900 3187 5934
rect -3187 5838 -3153 5900
rect 3153 5838 3187 5900
rect -3187 -5900 -3153 -5838
rect 3153 -5900 3187 -5838
rect -3187 -5934 -3091 -5900
rect 3091 -5934 3187 -5900
<< properties >>
string FIXED_BBOX -3170 -5917 3170 5917
string gencell sky130_fd_pr__res_xhigh_po_5p73
string library sky130
string parameters w 5.73 l 52.68 m 1 nx 5 wmin 5.730 lmin 0.50 rho 2000 val 100.002k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 5.730 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 1 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
