magic
tech sky130A
magscale 1 2
timestamp 1715803913
<< pwell >>
rect -5086 -862 5086 862
<< psubdiff >>
rect -5050 792 5050 826
rect -5050 730 -5016 792
rect 5016 730 5050 792
rect -5050 -792 -5016 -730
rect 5016 -792 5050 -730
rect -5050 -826 5050 -792
<< psubdiffcont >>
rect -5050 -730 -5016 730
rect 5016 -730 5050 730
<< xpolycontact >>
rect -4920 264 -3774 696
rect -4920 -696 -3774 -264
rect -3678 264 -2532 696
rect -3678 -696 -2532 -264
rect -2436 264 -1290 696
rect -2436 -696 -1290 -264
rect -1194 264 -48 696
rect -1194 -696 -48 -264
rect 48 264 1194 696
rect 48 -696 1194 -264
rect 1290 264 2436 696
rect 1290 -696 2436 -264
rect 2532 264 3678 696
rect 2532 -696 3678 -264
rect 3774 264 4920 696
rect 3774 -696 4920 -264
<< xpolyres >>
rect -4920 -264 -3774 264
rect -3678 -264 -2532 264
rect -2436 -264 -1290 264
rect -1194 -264 -48 264
rect 48 -264 1194 264
rect 1290 -264 2436 264
rect 2532 -264 3678 264
rect 3774 -264 4920 264
<< locali >>
rect -5050 792 5050 826
rect -5050 730 -5016 792
rect 5016 730 5050 792
rect -5050 -792 -5016 -730
rect 5016 -792 5050 -730
rect -5050 -826 5050 -792
<< viali >>
rect -4904 281 -3790 678
rect -3662 281 -2548 678
rect -2420 281 -1306 678
rect -1178 281 -64 678
rect 64 281 1178 678
rect 1306 281 2420 678
rect 2548 281 3662 678
rect 3790 281 4904 678
rect -4904 -678 -3790 -281
rect -3662 -678 -2548 -281
rect -2420 -678 -1306 -281
rect -1178 -678 -64 -281
rect 64 -678 1178 -281
rect 1306 -678 2420 -281
rect 2548 -678 3662 -281
rect 3790 -678 4904 -281
<< metal1 >>
rect -4916 678 -3778 684
rect -4916 281 -4904 678
rect -3790 281 -3778 678
rect -4916 275 -3778 281
rect -3674 678 -2536 684
rect -3674 281 -3662 678
rect -2548 281 -2536 678
rect -3674 275 -2536 281
rect -2432 678 -1294 684
rect -2432 281 -2420 678
rect -1306 281 -1294 678
rect -2432 275 -1294 281
rect -1190 678 -52 684
rect -1190 281 -1178 678
rect -64 281 -52 678
rect -1190 275 -52 281
rect 52 678 1190 684
rect 52 281 64 678
rect 1178 281 1190 678
rect 52 275 1190 281
rect 1294 678 2432 684
rect 1294 281 1306 678
rect 2420 281 2432 678
rect 1294 275 2432 281
rect 2536 678 3674 684
rect 2536 281 2548 678
rect 3662 281 3674 678
rect 2536 275 3674 281
rect 3778 678 4916 684
rect 3778 281 3790 678
rect 4904 281 4916 678
rect 3778 275 4916 281
rect -4916 -281 -3778 -275
rect -4916 -678 -4904 -281
rect -3790 -678 -3778 -281
rect -4916 -684 -3778 -678
rect -3674 -281 -2536 -275
rect -3674 -678 -3662 -281
rect -2548 -678 -2536 -281
rect -3674 -684 -2536 -678
rect -2432 -281 -1294 -275
rect -2432 -678 -2420 -281
rect -1306 -678 -1294 -281
rect -2432 -684 -1294 -678
rect -1190 -281 -52 -275
rect -1190 -678 -1178 -281
rect -64 -678 -52 -281
rect -1190 -684 -52 -678
rect 52 -281 1190 -275
rect 52 -678 64 -281
rect 1178 -678 1190 -281
rect 52 -684 1190 -678
rect 1294 -281 2432 -275
rect 1294 -678 1306 -281
rect 2420 -678 2432 -281
rect 1294 -684 2432 -678
rect 2536 -281 3674 -275
rect 2536 -678 2548 -281
rect 3662 -678 3674 -281
rect 2536 -684 3674 -678
rect 3778 -281 4916 -275
rect 3778 -678 3790 -281
rect 4904 -678 4916 -281
rect 3778 -684 4916 -678
<< properties >>
string FIXED_BBOX -5033 -809 5033 809
string gencell sky130_fd_pr__res_xhigh_po_5p73
string library sky130
string parameters w 5.73 l 2.8 m 1 nx 8 wmin 5.730 lmin 0.50 rho 2000 val 1.043k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 5.730 guard 1 glc 1 grc 1 gtc 0 gbc 0 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>
